magic
tech scmos
timestamp 1555071769 
<< pdiffusion >>
rect 1 -10 7 -4
rect 8 -10 14 -4
rect 15 -10 21 -4
rect 71 -10 77 -4
rect 92 -10 95 -4
rect 99 -10 105 -4
rect 106 -10 112 -4
rect 113 -10 116 -4
rect 176 -10 182 -4
rect 183 -10 186 -4
rect 190 -10 196 -4
rect 197 -10 200 -4
rect 1 -23 7 -17
rect 8 -23 14 -17
rect 15 -23 21 -17
rect 57 -23 60 -17
rect 64 -23 70 -17
rect 71 -23 77 -17
rect 78 -23 81 -17
rect 85 -23 91 -17
rect 92 -23 95 -17
rect 99 -23 105 -17
rect 106 -23 112 -17
rect 113 -23 119 -17
rect 127 -23 130 -17
rect 176 -23 179 -17
rect 183 -23 189 -17
rect 197 -23 203 -17
rect 204 -23 207 -17
rect 1 -42 7 -36
rect 8 -42 14 -36
rect 43 -42 49 -36
rect 50 -42 53 -36
rect 57 -42 60 -36
rect 64 -42 70 -36
rect 71 -42 77 -36
rect 78 -42 84 -36
rect 85 -42 91 -36
rect 92 -42 98 -36
rect 99 -42 105 -36
rect 106 -42 112 -36
rect 113 -42 119 -36
rect 120 -42 123 -36
rect 127 -42 130 -36
rect 134 -42 140 -36
rect 141 -42 144 -36
rect 148 -42 154 -36
rect 155 -42 158 -36
rect 169 -42 172 -36
rect 176 -42 182 -36
rect 183 -42 186 -36
rect 1 -63 7 -57
rect 29 -63 32 -57
rect 36 -63 39 -57
rect 43 -63 49 -57
rect 50 -63 53 -57
rect 57 -63 60 -57
rect 64 -63 70 -57
rect 71 -63 77 -57
rect 78 -63 84 -57
rect 85 -63 88 -57
rect 92 -63 95 -57
rect 99 -63 105 -57
rect 106 -63 112 -57
rect 113 -63 116 -57
rect 120 -63 123 -57
rect 127 -63 133 -57
rect 134 -63 140 -57
rect 141 -63 144 -57
rect 148 -63 151 -57
rect 155 -63 161 -57
rect 162 -63 165 -57
rect 169 -63 172 -57
rect 176 -63 179 -57
rect 183 -63 189 -57
rect 190 -63 193 -57
rect 50 -92 56 -86
rect 64 -92 70 -86
rect 71 -92 74 -86
rect 78 -92 81 -86
rect 85 -92 91 -86
rect 92 -92 95 -86
rect 99 -92 105 -86
rect 106 -92 112 -86
rect 113 -92 116 -86
rect 120 -92 123 -86
rect 127 -92 133 -86
rect 134 -92 137 -86
rect 141 -92 147 -86
rect 148 -92 154 -86
rect 155 -92 158 -86
rect 162 -92 165 -86
rect 169 -92 172 -86
rect 176 -92 179 -86
rect 183 -92 186 -86
rect 190 -92 196 -86
rect 197 -92 200 -86
rect 204 -92 207 -86
rect 211 -92 214 -86
rect 218 -92 221 -86
rect 225 -92 228 -86
rect 232 -92 235 -86
rect 239 -92 245 -86
rect 246 -92 252 -86
rect 1 -121 4 -115
rect 8 -121 11 -115
rect 15 -121 21 -115
rect 22 -121 25 -115
rect 29 -121 32 -115
rect 36 -121 42 -115
rect 43 -121 49 -115
rect 50 -121 53 -115
rect 57 -121 60 -115
rect 64 -121 70 -115
rect 71 -121 77 -115
rect 78 -121 84 -115
rect 85 -121 91 -115
rect 92 -121 95 -115
rect 99 -121 105 -115
rect 106 -121 109 -115
rect 113 -121 119 -115
rect 120 -121 126 -115
rect 127 -121 130 -115
rect 134 -121 137 -115
rect 141 -121 147 -115
rect 148 -121 154 -115
rect 155 -121 161 -115
rect 162 -121 165 -115
rect 169 -121 172 -115
rect 176 -121 179 -115
rect 183 -121 186 -115
rect 190 -121 193 -115
rect 197 -121 200 -115
rect 204 -121 207 -115
rect 211 -121 214 -115
rect 218 -121 221 -115
rect 225 -121 228 -115
rect 232 -121 235 -115
rect 239 -121 242 -115
rect 246 -121 249 -115
rect 253 -121 259 -115
rect 1 -166 4 -160
rect 8 -166 11 -160
rect 15 -166 21 -160
rect 22 -166 28 -160
rect 29 -166 35 -160
rect 36 -166 42 -160
rect 43 -166 49 -160
rect 50 -166 53 -160
rect 57 -166 63 -160
rect 64 -166 67 -160
rect 71 -166 74 -160
rect 78 -166 84 -160
rect 85 -166 91 -160
rect 92 -166 98 -160
rect 99 -166 102 -160
rect 106 -166 112 -160
rect 113 -166 119 -160
rect 120 -166 123 -160
rect 127 -166 130 -160
rect 134 -166 140 -160
rect 141 -166 144 -160
rect 148 -166 151 -160
rect 155 -166 161 -160
rect 162 -166 165 -160
rect 169 -166 172 -160
rect 176 -166 179 -160
rect 183 -166 189 -160
rect 190 -166 193 -160
rect 197 -166 200 -160
rect 204 -166 207 -160
rect 211 -166 214 -160
rect 218 -166 221 -160
rect 225 -166 228 -160
rect 232 -166 235 -160
rect 239 -166 242 -160
rect 246 -166 249 -160
rect 253 -166 256 -160
rect 260 -166 263 -160
rect 267 -166 270 -160
rect 274 -166 280 -160
rect 22 -197 25 -191
rect 29 -197 32 -191
rect 36 -197 42 -191
rect 43 -197 49 -191
rect 50 -197 53 -191
rect 57 -197 60 -191
rect 64 -197 70 -191
rect 71 -197 74 -191
rect 78 -197 84 -191
rect 85 -197 88 -191
rect 92 -197 98 -191
rect 99 -197 105 -191
rect 106 -197 112 -191
rect 113 -197 119 -191
rect 120 -197 123 -191
rect 127 -197 133 -191
rect 134 -197 140 -191
rect 141 -197 147 -191
rect 148 -197 154 -191
rect 155 -197 158 -191
rect 162 -197 165 -191
rect 169 -197 172 -191
rect 176 -197 179 -191
rect 183 -197 189 -191
rect 190 -197 196 -191
rect 197 -197 200 -191
rect 204 -197 207 -191
rect 211 -197 214 -191
rect 218 -197 221 -191
rect 225 -197 228 -191
rect 232 -197 235 -191
rect 239 -197 242 -191
rect 246 -197 249 -191
rect 253 -197 256 -191
rect 260 -197 263 -191
rect 281 -197 287 -191
rect 29 -232 35 -226
rect 36 -232 39 -226
rect 43 -232 49 -226
rect 50 -232 53 -226
rect 57 -232 60 -226
rect 64 -232 67 -226
rect 71 -232 77 -226
rect 78 -232 84 -226
rect 85 -232 88 -226
rect 92 -232 98 -226
rect 99 -232 102 -226
rect 106 -232 109 -226
rect 113 -232 119 -226
rect 120 -232 123 -226
rect 127 -232 130 -226
rect 134 -232 140 -226
rect 141 -232 144 -226
rect 148 -232 154 -226
rect 155 -232 161 -226
rect 162 -232 165 -226
rect 169 -232 172 -226
rect 176 -232 182 -226
rect 183 -232 186 -226
rect 190 -232 196 -226
rect 197 -232 200 -226
rect 204 -232 207 -226
rect 211 -232 214 -226
rect 218 -232 221 -226
rect 225 -232 228 -226
rect 232 -232 235 -226
rect 239 -232 242 -226
rect 246 -232 249 -226
rect 253 -232 256 -226
rect 260 -232 266 -226
rect 267 -232 273 -226
rect 274 -232 280 -226
rect 281 -232 284 -226
rect 288 -232 291 -226
rect 15 -263 18 -257
rect 22 -263 28 -257
rect 29 -263 32 -257
rect 36 -263 39 -257
rect 43 -263 49 -257
rect 50 -263 56 -257
rect 57 -263 60 -257
rect 64 -263 67 -257
rect 71 -263 74 -257
rect 78 -263 81 -257
rect 85 -263 88 -257
rect 92 -263 95 -257
rect 99 -263 105 -257
rect 106 -263 112 -257
rect 113 -263 119 -257
rect 120 -263 123 -257
rect 127 -263 130 -257
rect 134 -263 140 -257
rect 141 -263 144 -257
rect 148 -263 151 -257
rect 155 -263 158 -257
rect 162 -263 165 -257
rect 169 -263 175 -257
rect 176 -263 182 -257
rect 183 -263 186 -257
rect 190 -263 196 -257
rect 197 -263 200 -257
rect 204 -263 207 -257
rect 211 -263 214 -257
rect 218 -263 221 -257
rect 225 -263 228 -257
rect 232 -263 235 -257
rect 239 -263 242 -257
rect 246 -263 249 -257
rect 253 -263 256 -257
rect 281 -263 284 -257
rect 288 -263 294 -257
rect 64 -290 67 -284
rect 71 -290 74 -284
rect 78 -290 84 -284
rect 85 -290 91 -284
rect 92 -290 98 -284
rect 99 -290 105 -284
rect 106 -290 109 -284
rect 113 -290 119 -284
rect 120 -290 123 -284
rect 127 -290 130 -284
rect 134 -290 137 -284
rect 141 -290 144 -284
rect 148 -290 151 -284
rect 155 -290 158 -284
rect 162 -290 168 -284
rect 169 -290 172 -284
rect 183 -290 189 -284
rect 190 -290 196 -284
rect 197 -290 200 -284
rect 204 -290 210 -284
rect 239 -290 242 -284
rect 246 -290 252 -284
rect 253 -290 256 -284
rect 50 -313 53 -307
rect 57 -313 63 -307
rect 64 -313 67 -307
rect 71 -313 77 -307
rect 78 -313 84 -307
rect 85 -313 91 -307
rect 92 -313 98 -307
rect 99 -313 105 -307
rect 106 -313 112 -307
rect 113 -313 119 -307
rect 120 -313 123 -307
rect 127 -313 130 -307
rect 134 -313 140 -307
rect 141 -313 144 -307
rect 148 -313 151 -307
rect 155 -313 158 -307
rect 162 -313 165 -307
rect 169 -313 172 -307
rect 176 -313 179 -307
rect 218 -313 221 -307
rect 225 -313 231 -307
rect 232 -313 238 -307
rect 239 -313 242 -307
rect 36 -342 39 -336
rect 43 -342 46 -336
rect 50 -342 53 -336
rect 57 -342 63 -336
rect 64 -342 67 -336
rect 71 -342 74 -336
rect 78 -342 84 -336
rect 85 -342 91 -336
rect 92 -342 98 -336
rect 99 -342 105 -336
rect 106 -342 109 -336
rect 113 -342 119 -336
rect 120 -342 123 -336
rect 127 -342 133 -336
rect 134 -342 140 -336
rect 141 -342 147 -336
rect 148 -342 151 -336
rect 155 -342 161 -336
rect 162 -342 165 -336
rect 169 -342 172 -336
rect 176 -342 179 -336
rect 183 -342 186 -336
rect 190 -342 193 -336
rect 197 -342 200 -336
rect 204 -342 207 -336
rect 211 -342 217 -336
rect 218 -342 221 -336
rect 57 -369 60 -363
rect 64 -369 67 -363
rect 71 -369 74 -363
rect 78 -369 81 -363
rect 85 -369 88 -363
rect 92 -369 98 -363
rect 99 -369 105 -363
rect 106 -369 112 -363
rect 113 -369 119 -363
rect 120 -369 123 -363
rect 127 -369 130 -363
rect 134 -369 137 -363
rect 141 -369 147 -363
rect 148 -369 151 -363
rect 155 -369 161 -363
rect 162 -369 165 -363
rect 169 -369 175 -363
rect 176 -369 179 -363
rect 183 -369 186 -363
rect 190 -369 196 -363
rect 197 -369 200 -363
rect 71 -392 74 -386
rect 78 -392 81 -386
rect 85 -392 88 -386
rect 92 -392 98 -386
rect 99 -392 105 -386
rect 106 -392 109 -386
rect 113 -392 119 -386
rect 120 -392 126 -386
rect 127 -392 130 -386
rect 134 -392 140 -386
rect 141 -392 144 -386
rect 148 -392 151 -386
rect 155 -392 158 -386
rect 162 -392 165 -386
rect 169 -392 175 -386
rect 78 -413 84 -407
rect 85 -413 88 -407
rect 92 -413 95 -407
rect 99 -413 105 -407
rect 106 -413 109 -407
rect 113 -413 119 -407
rect 120 -413 123 -407
rect 127 -413 133 -407
rect 141 -413 147 -407
rect 155 -413 158 -407
rect 162 -413 168 -407
rect 169 -413 175 -407
rect 85 -426 91 -420
rect 92 -426 95 -420
rect 113 -426 119 -420
rect 120 -426 123 -420
rect 162 -426 165 -420
rect 169 -426 175 -420
<< polysilicon >>
rect 75 -11 76 -9
rect 93 -5 94 -3
rect 93 -11 94 -9
rect 100 -5 101 -3
rect 103 -5 104 -3
rect 107 -11 108 -9
rect 114 -5 115 -3
rect 114 -11 115 -9
rect 177 -5 178 -3
rect 184 -5 185 -3
rect 184 -11 185 -9
rect 191 -5 192 -3
rect 191 -11 192 -9
rect 198 -5 199 -3
rect 198 -11 199 -9
rect 58 -18 59 -16
rect 58 -24 59 -22
rect 68 -18 69 -16
rect 65 -24 66 -22
rect 75 -18 76 -16
rect 79 -18 80 -16
rect 79 -24 80 -22
rect 89 -18 90 -16
rect 93 -18 94 -16
rect 93 -24 94 -22
rect 100 -18 101 -16
rect 107 -18 108 -16
rect 117 -18 118 -16
rect 128 -18 129 -16
rect 128 -24 129 -22
rect 177 -18 178 -16
rect 177 -24 178 -22
rect 184 -18 185 -16
rect 198 -24 199 -22
rect 205 -18 206 -16
rect 205 -24 206 -22
rect 44 -43 45 -41
rect 51 -37 52 -35
rect 51 -43 52 -41
rect 58 -37 59 -35
rect 58 -43 59 -41
rect 65 -37 66 -35
rect 65 -43 66 -41
rect 72 -43 73 -41
rect 79 -37 80 -35
rect 79 -43 80 -41
rect 86 -37 87 -35
rect 86 -43 87 -41
rect 93 -37 94 -35
rect 96 -37 97 -35
rect 100 -37 101 -35
rect 103 -43 104 -41
rect 107 -37 108 -35
rect 107 -43 108 -41
rect 110 -43 111 -41
rect 117 -37 118 -35
rect 114 -43 115 -41
rect 117 -43 118 -41
rect 121 -37 122 -35
rect 121 -43 122 -41
rect 128 -37 129 -35
rect 128 -43 129 -41
rect 138 -43 139 -41
rect 142 -37 143 -35
rect 142 -43 143 -41
rect 149 -37 150 -35
rect 152 -43 153 -41
rect 156 -37 157 -35
rect 156 -43 157 -41
rect 170 -37 171 -35
rect 170 -43 171 -41
rect 180 -37 181 -35
rect 177 -43 178 -41
rect 184 -37 185 -35
rect 184 -43 185 -41
rect 30 -58 31 -56
rect 30 -64 31 -62
rect 37 -58 38 -56
rect 37 -64 38 -62
rect 47 -64 48 -62
rect 51 -58 52 -56
rect 51 -64 52 -62
rect 58 -58 59 -56
rect 58 -64 59 -62
rect 68 -58 69 -56
rect 75 -58 76 -56
rect 72 -64 73 -62
rect 75 -64 76 -62
rect 79 -58 80 -56
rect 79 -64 80 -62
rect 82 -64 83 -62
rect 86 -58 87 -56
rect 86 -64 87 -62
rect 93 -58 94 -56
rect 93 -64 94 -62
rect 103 -58 104 -56
rect 100 -64 101 -62
rect 107 -58 108 -56
rect 114 -58 115 -56
rect 114 -64 115 -62
rect 121 -58 122 -56
rect 121 -64 122 -62
rect 131 -58 132 -56
rect 128 -64 129 -62
rect 131 -64 132 -62
rect 135 -64 136 -62
rect 138 -64 139 -62
rect 142 -58 143 -56
rect 142 -64 143 -62
rect 149 -58 150 -56
rect 149 -64 150 -62
rect 156 -58 157 -56
rect 159 -58 160 -56
rect 163 -58 164 -56
rect 163 -64 164 -62
rect 170 -58 171 -56
rect 170 -64 171 -62
rect 177 -58 178 -56
rect 177 -64 178 -62
rect 184 -58 185 -56
rect 187 -64 188 -62
rect 191 -58 192 -56
rect 191 -64 192 -62
rect 54 -87 55 -85
rect 51 -93 52 -91
rect 65 -87 66 -85
rect 68 -87 69 -85
rect 72 -87 73 -85
rect 72 -93 73 -91
rect 79 -87 80 -85
rect 79 -93 80 -91
rect 86 -87 87 -85
rect 89 -87 90 -85
rect 86 -93 87 -91
rect 89 -93 90 -91
rect 93 -87 94 -85
rect 93 -93 94 -91
rect 100 -87 101 -85
rect 103 -93 104 -91
rect 107 -87 108 -85
rect 110 -87 111 -85
rect 114 -87 115 -85
rect 114 -93 115 -91
rect 121 -87 122 -85
rect 121 -93 122 -91
rect 128 -87 129 -85
rect 131 -87 132 -85
rect 131 -93 132 -91
rect 135 -87 136 -85
rect 135 -93 136 -91
rect 142 -87 143 -85
rect 142 -93 143 -91
rect 145 -93 146 -91
rect 152 -87 153 -85
rect 152 -93 153 -91
rect 156 -87 157 -85
rect 156 -93 157 -91
rect 163 -87 164 -85
rect 163 -93 164 -91
rect 170 -87 171 -85
rect 170 -93 171 -91
rect 177 -87 178 -85
rect 177 -93 178 -91
rect 184 -87 185 -85
rect 184 -93 185 -91
rect 191 -93 192 -91
rect 194 -93 195 -91
rect 198 -87 199 -85
rect 198 -93 199 -91
rect 205 -87 206 -85
rect 205 -93 206 -91
rect 212 -87 213 -85
rect 212 -93 213 -91
rect 219 -87 220 -85
rect 219 -93 220 -91
rect 226 -87 227 -85
rect 226 -93 227 -91
rect 233 -87 234 -85
rect 233 -93 234 -91
rect 243 -87 244 -85
rect 247 -87 248 -85
rect 247 -93 248 -91
rect 250 -93 251 -91
rect 2 -116 3 -114
rect 2 -122 3 -120
rect 9 -116 10 -114
rect 9 -122 10 -120
rect 19 -122 20 -120
rect 23 -116 24 -114
rect 23 -122 24 -120
rect 30 -116 31 -114
rect 30 -122 31 -120
rect 37 -122 38 -120
rect 40 -122 41 -120
rect 44 -116 45 -114
rect 47 -116 48 -114
rect 51 -116 52 -114
rect 51 -122 52 -120
rect 58 -116 59 -114
rect 58 -122 59 -120
rect 68 -116 69 -114
rect 68 -122 69 -120
rect 75 -116 76 -114
rect 82 -116 83 -114
rect 79 -122 80 -120
rect 82 -122 83 -120
rect 86 -116 87 -114
rect 89 -122 90 -120
rect 93 -116 94 -114
rect 93 -122 94 -120
rect 100 -116 101 -114
rect 100 -122 101 -120
rect 107 -116 108 -114
rect 107 -122 108 -120
rect 114 -116 115 -114
rect 117 -116 118 -114
rect 114 -122 115 -120
rect 121 -116 122 -114
rect 124 -116 125 -114
rect 121 -122 122 -120
rect 128 -116 129 -114
rect 128 -122 129 -120
rect 135 -116 136 -114
rect 135 -122 136 -120
rect 145 -116 146 -114
rect 145 -122 146 -120
rect 149 -116 150 -114
rect 149 -122 150 -120
rect 152 -122 153 -120
rect 156 -116 157 -114
rect 159 -116 160 -114
rect 159 -122 160 -120
rect 163 -116 164 -114
rect 163 -122 164 -120
rect 170 -116 171 -114
rect 170 -122 171 -120
rect 177 -116 178 -114
rect 177 -122 178 -120
rect 184 -116 185 -114
rect 184 -122 185 -120
rect 191 -116 192 -114
rect 191 -122 192 -120
rect 198 -116 199 -114
rect 198 -122 199 -120
rect 205 -116 206 -114
rect 205 -122 206 -120
rect 212 -116 213 -114
rect 212 -122 213 -120
rect 219 -116 220 -114
rect 219 -122 220 -120
rect 226 -116 227 -114
rect 226 -122 227 -120
rect 233 -116 234 -114
rect 233 -122 234 -120
rect 240 -116 241 -114
rect 240 -122 241 -120
rect 247 -116 248 -114
rect 247 -122 248 -120
rect 254 -116 255 -114
rect 2 -161 3 -159
rect 2 -167 3 -165
rect 9 -161 10 -159
rect 9 -167 10 -165
rect 19 -161 20 -159
rect 26 -167 27 -165
rect 30 -161 31 -159
rect 33 -161 34 -159
rect 40 -161 41 -159
rect 40 -167 41 -165
rect 47 -161 48 -159
rect 47 -167 48 -165
rect 51 -161 52 -159
rect 51 -167 52 -165
rect 58 -161 59 -159
rect 58 -167 59 -165
rect 65 -161 66 -159
rect 65 -167 66 -165
rect 72 -161 73 -159
rect 72 -167 73 -165
rect 79 -167 80 -165
rect 82 -167 83 -165
rect 86 -161 87 -159
rect 89 -161 90 -159
rect 86 -167 87 -165
rect 89 -167 90 -165
rect 96 -167 97 -165
rect 100 -161 101 -159
rect 100 -167 101 -165
rect 107 -161 108 -159
rect 107 -167 108 -165
rect 110 -167 111 -165
rect 114 -161 115 -159
rect 117 -161 118 -159
rect 114 -167 115 -165
rect 117 -167 118 -165
rect 121 -161 122 -159
rect 121 -167 122 -165
rect 128 -161 129 -159
rect 128 -167 129 -165
rect 135 -161 136 -159
rect 138 -161 139 -159
rect 135 -167 136 -165
rect 138 -167 139 -165
rect 142 -161 143 -159
rect 142 -167 143 -165
rect 149 -161 150 -159
rect 149 -167 150 -165
rect 156 -161 157 -159
rect 159 -167 160 -165
rect 163 -161 164 -159
rect 163 -167 164 -165
rect 170 -161 171 -159
rect 170 -167 171 -165
rect 177 -161 178 -159
rect 177 -167 178 -165
rect 187 -161 188 -159
rect 184 -167 185 -165
rect 191 -161 192 -159
rect 191 -167 192 -165
rect 198 -161 199 -159
rect 198 -167 199 -165
rect 205 -161 206 -159
rect 205 -167 206 -165
rect 212 -161 213 -159
rect 212 -167 213 -165
rect 219 -161 220 -159
rect 219 -167 220 -165
rect 226 -161 227 -159
rect 226 -167 227 -165
rect 233 -161 234 -159
rect 233 -167 234 -165
rect 240 -161 241 -159
rect 240 -167 241 -165
rect 247 -161 248 -159
rect 247 -167 248 -165
rect 254 -161 255 -159
rect 254 -167 255 -165
rect 261 -161 262 -159
rect 261 -167 262 -165
rect 268 -161 269 -159
rect 268 -167 269 -165
rect 275 -161 276 -159
rect 275 -167 276 -165
rect 23 -192 24 -190
rect 23 -198 24 -196
rect 30 -192 31 -190
rect 30 -198 31 -196
rect 40 -192 41 -190
rect 37 -198 38 -196
rect 44 -192 45 -190
rect 44 -198 45 -196
rect 47 -198 48 -196
rect 51 -192 52 -190
rect 51 -198 52 -196
rect 58 -192 59 -190
rect 58 -198 59 -196
rect 65 -192 66 -190
rect 68 -198 69 -196
rect 72 -192 73 -190
rect 72 -198 73 -196
rect 82 -192 83 -190
rect 86 -192 87 -190
rect 86 -198 87 -196
rect 93 -198 94 -196
rect 96 -198 97 -196
rect 103 -192 104 -190
rect 103 -198 104 -196
rect 107 -192 108 -190
rect 107 -198 108 -196
rect 110 -198 111 -196
rect 114 -192 115 -190
rect 117 -198 118 -196
rect 121 -192 122 -190
rect 121 -198 122 -196
rect 128 -192 129 -190
rect 128 -198 129 -196
rect 135 -192 136 -190
rect 138 -192 139 -190
rect 135 -198 136 -196
rect 142 -198 143 -196
rect 145 -198 146 -196
rect 149 -192 150 -190
rect 152 -192 153 -190
rect 149 -198 150 -196
rect 152 -198 153 -196
rect 156 -192 157 -190
rect 156 -198 157 -196
rect 163 -192 164 -190
rect 163 -198 164 -196
rect 170 -192 171 -190
rect 170 -198 171 -196
rect 177 -192 178 -190
rect 177 -198 178 -196
rect 187 -192 188 -190
rect 187 -198 188 -196
rect 194 -192 195 -190
rect 194 -198 195 -196
rect 198 -192 199 -190
rect 198 -198 199 -196
rect 205 -192 206 -190
rect 205 -198 206 -196
rect 212 -192 213 -190
rect 212 -198 213 -196
rect 219 -192 220 -190
rect 219 -198 220 -196
rect 226 -192 227 -190
rect 226 -198 227 -196
rect 233 -192 234 -190
rect 233 -198 234 -196
rect 240 -192 241 -190
rect 240 -198 241 -196
rect 247 -192 248 -190
rect 247 -198 248 -196
rect 254 -192 255 -190
rect 254 -198 255 -196
rect 261 -192 262 -190
rect 261 -198 262 -196
rect 282 -198 283 -196
rect 30 -227 31 -225
rect 37 -227 38 -225
rect 37 -233 38 -231
rect 44 -227 45 -225
rect 51 -227 52 -225
rect 51 -233 52 -231
rect 58 -227 59 -225
rect 58 -233 59 -231
rect 65 -227 66 -225
rect 65 -233 66 -231
rect 75 -233 76 -231
rect 82 -227 83 -225
rect 79 -233 80 -231
rect 86 -227 87 -225
rect 86 -233 87 -231
rect 93 -227 94 -225
rect 96 -227 97 -225
rect 93 -233 94 -231
rect 100 -227 101 -225
rect 100 -233 101 -231
rect 107 -227 108 -225
rect 107 -233 108 -231
rect 114 -227 115 -225
rect 117 -227 118 -225
rect 114 -233 115 -231
rect 117 -233 118 -231
rect 121 -227 122 -225
rect 121 -233 122 -231
rect 128 -227 129 -225
rect 128 -233 129 -231
rect 135 -227 136 -225
rect 138 -227 139 -225
rect 142 -227 143 -225
rect 142 -233 143 -231
rect 149 -227 150 -225
rect 152 -227 153 -225
rect 159 -227 160 -225
rect 156 -233 157 -231
rect 159 -233 160 -231
rect 163 -227 164 -225
rect 163 -233 164 -231
rect 170 -227 171 -225
rect 170 -233 171 -231
rect 177 -227 178 -225
rect 180 -227 181 -225
rect 184 -227 185 -225
rect 184 -233 185 -231
rect 191 -227 192 -225
rect 194 -227 195 -225
rect 191 -233 192 -231
rect 198 -227 199 -225
rect 198 -233 199 -231
rect 205 -227 206 -225
rect 205 -233 206 -231
rect 212 -227 213 -225
rect 212 -233 213 -231
rect 219 -227 220 -225
rect 219 -233 220 -231
rect 226 -227 227 -225
rect 226 -233 227 -231
rect 233 -227 234 -225
rect 233 -233 234 -231
rect 240 -227 241 -225
rect 240 -233 241 -231
rect 247 -227 248 -225
rect 247 -233 248 -231
rect 254 -227 255 -225
rect 254 -233 255 -231
rect 261 -227 262 -225
rect 264 -227 265 -225
rect 261 -233 262 -231
rect 264 -233 265 -231
rect 271 -227 272 -225
rect 278 -227 279 -225
rect 275 -233 276 -231
rect 282 -227 283 -225
rect 282 -233 283 -231
rect 289 -227 290 -225
rect 289 -233 290 -231
rect 16 -258 17 -256
rect 16 -264 17 -262
rect 26 -264 27 -262
rect 30 -258 31 -256
rect 30 -264 31 -262
rect 37 -258 38 -256
rect 37 -264 38 -262
rect 44 -258 45 -256
rect 44 -264 45 -262
rect 47 -264 48 -262
rect 51 -264 52 -262
rect 54 -264 55 -262
rect 58 -258 59 -256
rect 58 -264 59 -262
rect 65 -258 66 -256
rect 65 -264 66 -262
rect 72 -258 73 -256
rect 72 -264 73 -262
rect 79 -258 80 -256
rect 79 -264 80 -262
rect 86 -258 87 -256
rect 86 -264 87 -262
rect 93 -258 94 -256
rect 93 -264 94 -262
rect 103 -258 104 -256
rect 100 -264 101 -262
rect 103 -264 104 -262
rect 107 -258 108 -256
rect 107 -264 108 -262
rect 114 -258 115 -256
rect 117 -258 118 -256
rect 114 -264 115 -262
rect 117 -264 118 -262
rect 121 -258 122 -256
rect 121 -264 122 -262
rect 128 -258 129 -256
rect 128 -264 129 -262
rect 135 -258 136 -256
rect 135 -264 136 -262
rect 142 -258 143 -256
rect 142 -264 143 -262
rect 149 -258 150 -256
rect 149 -264 150 -262
rect 156 -258 157 -256
rect 156 -264 157 -262
rect 163 -258 164 -256
rect 163 -264 164 -262
rect 170 -258 171 -256
rect 173 -258 174 -256
rect 173 -264 174 -262
rect 177 -258 178 -256
rect 180 -258 181 -256
rect 177 -264 178 -262
rect 180 -264 181 -262
rect 184 -258 185 -256
rect 184 -264 185 -262
rect 191 -258 192 -256
rect 191 -264 192 -262
rect 198 -258 199 -256
rect 198 -264 199 -262
rect 205 -258 206 -256
rect 205 -264 206 -262
rect 212 -258 213 -256
rect 212 -264 213 -262
rect 219 -258 220 -256
rect 219 -264 220 -262
rect 226 -258 227 -256
rect 226 -264 227 -262
rect 233 -258 234 -256
rect 233 -264 234 -262
rect 240 -258 241 -256
rect 240 -264 241 -262
rect 247 -258 248 -256
rect 247 -264 248 -262
rect 254 -258 255 -256
rect 254 -264 255 -262
rect 282 -258 283 -256
rect 282 -264 283 -262
rect 289 -264 290 -262
rect 65 -285 66 -283
rect 65 -291 66 -289
rect 72 -285 73 -283
rect 72 -291 73 -289
rect 82 -291 83 -289
rect 86 -285 87 -283
rect 89 -285 90 -283
rect 86 -291 87 -289
rect 89 -291 90 -289
rect 93 -285 94 -283
rect 96 -285 97 -283
rect 96 -291 97 -289
rect 103 -285 104 -283
rect 103 -291 104 -289
rect 107 -285 108 -283
rect 107 -291 108 -289
rect 114 -291 115 -289
rect 117 -291 118 -289
rect 121 -285 122 -283
rect 121 -291 122 -289
rect 128 -285 129 -283
rect 128 -291 129 -289
rect 135 -285 136 -283
rect 135 -291 136 -289
rect 142 -285 143 -283
rect 142 -291 143 -289
rect 149 -285 150 -283
rect 149 -291 150 -289
rect 156 -285 157 -283
rect 156 -291 157 -289
rect 166 -285 167 -283
rect 163 -291 164 -289
rect 170 -285 171 -283
rect 170 -291 171 -289
rect 184 -291 185 -289
rect 191 -285 192 -283
rect 194 -285 195 -283
rect 191 -291 192 -289
rect 194 -291 195 -289
rect 198 -285 199 -283
rect 198 -291 199 -289
rect 205 -285 206 -283
rect 208 -285 209 -283
rect 205 -291 206 -289
rect 240 -285 241 -283
rect 240 -291 241 -289
rect 247 -285 248 -283
rect 250 -291 251 -289
rect 254 -285 255 -283
rect 254 -291 255 -289
rect 51 -308 52 -306
rect 51 -314 52 -312
rect 61 -314 62 -312
rect 65 -308 66 -306
rect 65 -314 66 -312
rect 75 -308 76 -306
rect 72 -314 73 -312
rect 75 -314 76 -312
rect 82 -308 83 -306
rect 86 -308 87 -306
rect 89 -308 90 -306
rect 89 -314 90 -312
rect 96 -308 97 -306
rect 93 -314 94 -312
rect 103 -308 104 -306
rect 100 -314 101 -312
rect 107 -308 108 -306
rect 110 -308 111 -306
rect 107 -314 108 -312
rect 114 -308 115 -306
rect 117 -308 118 -306
rect 114 -314 115 -312
rect 117 -314 118 -312
rect 121 -308 122 -306
rect 121 -314 122 -312
rect 128 -308 129 -306
rect 128 -314 129 -312
rect 138 -308 139 -306
rect 135 -314 136 -312
rect 138 -314 139 -312
rect 142 -308 143 -306
rect 142 -314 143 -312
rect 149 -308 150 -306
rect 149 -314 150 -312
rect 156 -308 157 -306
rect 156 -314 157 -312
rect 163 -308 164 -306
rect 163 -314 164 -312
rect 170 -308 171 -306
rect 170 -314 171 -312
rect 177 -308 178 -306
rect 177 -314 178 -312
rect 219 -308 220 -306
rect 219 -314 220 -312
rect 226 -314 227 -312
rect 233 -308 234 -306
rect 233 -314 234 -312
rect 236 -314 237 -312
rect 240 -308 241 -306
rect 240 -314 241 -312
rect 37 -337 38 -335
rect 37 -343 38 -341
rect 44 -337 45 -335
rect 44 -343 45 -341
rect 51 -337 52 -335
rect 51 -343 52 -341
rect 61 -337 62 -335
rect 58 -343 59 -341
rect 65 -337 66 -335
rect 65 -343 66 -341
rect 72 -337 73 -335
rect 72 -343 73 -341
rect 79 -337 80 -335
rect 79 -343 80 -341
rect 86 -337 87 -335
rect 89 -337 90 -335
rect 93 -337 94 -335
rect 96 -337 97 -335
rect 93 -343 94 -341
rect 96 -343 97 -341
rect 100 -337 101 -335
rect 100 -343 101 -341
rect 103 -343 104 -341
rect 107 -337 108 -335
rect 107 -343 108 -341
rect 117 -337 118 -335
rect 114 -343 115 -341
rect 117 -343 118 -341
rect 121 -337 122 -335
rect 121 -343 122 -341
rect 128 -337 129 -335
rect 131 -337 132 -335
rect 131 -343 132 -341
rect 135 -337 136 -335
rect 138 -337 139 -335
rect 138 -343 139 -341
rect 142 -337 143 -335
rect 142 -343 143 -341
rect 145 -343 146 -341
rect 149 -337 150 -335
rect 149 -343 150 -341
rect 159 -337 160 -335
rect 156 -343 157 -341
rect 163 -337 164 -335
rect 163 -343 164 -341
rect 170 -337 171 -335
rect 170 -343 171 -341
rect 177 -337 178 -335
rect 177 -343 178 -341
rect 184 -337 185 -335
rect 184 -343 185 -341
rect 191 -337 192 -335
rect 191 -343 192 -341
rect 198 -337 199 -335
rect 198 -343 199 -341
rect 205 -337 206 -335
rect 205 -343 206 -341
rect 212 -343 213 -341
rect 215 -343 216 -341
rect 219 -337 220 -335
rect 219 -343 220 -341
rect 58 -364 59 -362
rect 58 -370 59 -368
rect 65 -364 66 -362
rect 65 -370 66 -368
rect 72 -364 73 -362
rect 72 -370 73 -368
rect 79 -364 80 -362
rect 79 -370 80 -368
rect 86 -364 87 -362
rect 86 -370 87 -368
rect 96 -364 97 -362
rect 103 -364 104 -362
rect 100 -370 101 -368
rect 110 -364 111 -362
rect 107 -370 108 -368
rect 114 -370 115 -368
rect 117 -370 118 -368
rect 121 -364 122 -362
rect 121 -370 122 -368
rect 128 -364 129 -362
rect 128 -370 129 -368
rect 135 -364 136 -362
rect 135 -370 136 -368
rect 142 -364 143 -362
rect 142 -370 143 -368
rect 145 -370 146 -368
rect 149 -364 150 -362
rect 149 -370 150 -368
rect 156 -370 157 -368
rect 163 -364 164 -362
rect 163 -370 164 -368
rect 170 -364 171 -362
rect 177 -364 178 -362
rect 177 -370 178 -368
rect 184 -364 185 -362
rect 184 -370 185 -368
rect 194 -364 195 -362
rect 198 -364 199 -362
rect 198 -370 199 -368
rect 72 -387 73 -385
rect 72 -393 73 -391
rect 79 -387 80 -385
rect 79 -393 80 -391
rect 86 -387 87 -385
rect 86 -393 87 -391
rect 93 -387 94 -385
rect 96 -387 97 -385
rect 100 -387 101 -385
rect 103 -387 104 -385
rect 100 -393 101 -391
rect 107 -387 108 -385
rect 107 -393 108 -391
rect 114 -393 115 -391
rect 117 -393 118 -391
rect 121 -387 122 -385
rect 124 -387 125 -385
rect 121 -393 122 -391
rect 128 -387 129 -385
rect 128 -393 129 -391
rect 138 -387 139 -385
rect 138 -393 139 -391
rect 142 -387 143 -385
rect 142 -393 143 -391
rect 149 -387 150 -385
rect 149 -393 150 -391
rect 156 -387 157 -385
rect 156 -393 157 -391
rect 163 -387 164 -385
rect 163 -393 164 -391
rect 170 -387 171 -385
rect 173 -387 174 -385
rect 170 -393 171 -391
rect 79 -408 80 -406
rect 86 -408 87 -406
rect 86 -414 87 -412
rect 93 -408 94 -406
rect 93 -414 94 -412
rect 100 -414 101 -412
rect 107 -408 108 -406
rect 107 -414 108 -412
rect 117 -408 118 -406
rect 117 -414 118 -412
rect 121 -408 122 -406
rect 121 -414 122 -412
rect 128 -408 129 -406
rect 131 -408 132 -406
rect 142 -408 143 -406
rect 145 -408 146 -406
rect 156 -408 157 -406
rect 156 -414 157 -412
rect 163 -408 164 -406
rect 173 -408 174 -406
rect 89 -427 90 -425
rect 93 -421 94 -419
rect 93 -427 94 -425
rect 117 -427 118 -425
rect 121 -421 122 -419
rect 121 -427 122 -425
rect 163 -421 164 -419
rect 163 -427 164 -425
rect 170 -427 171 -425
<< metal1 >>
rect 93 0 104 1
rect 177 0 185 1
rect 191 0 199 1
rect 100 -2 115 -1
rect 58 -13 69 -12
rect 79 -13 90 -12
rect 93 -13 108 -12
rect 117 -13 129 -12
rect 184 -13 192 -12
rect 198 -13 206 -12
rect 93 -15 101 -14
rect 107 -15 115 -14
rect 177 -15 185 -14
rect 79 -26 87 -25
rect 93 -26 108 -25
rect 142 -26 150 -25
rect 170 -26 178 -25
rect 180 -26 185 -25
rect 198 -26 206 -25
rect 51 -28 94 -27
rect 96 -28 157 -27
rect 65 -30 80 -29
rect 100 -30 122 -29
rect 58 -32 66 -31
rect 58 -34 118 -33
rect 44 -45 52 -44
rect 58 -45 80 -44
rect 86 -45 115 -44
rect 138 -45 150 -44
rect 159 -45 192 -44
rect 30 -47 80 -46
rect 103 -47 122 -46
rect 142 -47 164 -46
rect 170 -47 178 -46
rect 37 -49 104 -48
rect 107 -49 129 -48
rect 152 -49 171 -48
rect 51 -51 66 -50
rect 68 -51 87 -50
rect 107 -51 115 -50
rect 117 -51 178 -50
rect 58 -53 73 -52
rect 75 -53 94 -52
rect 110 -53 143 -52
rect 121 -55 132 -54
rect 30 -66 73 -65
rect 82 -66 185 -65
rect 187 -66 220 -65
rect 233 -66 244 -65
rect 37 -68 66 -67
rect 72 -68 139 -67
rect 152 -68 157 -67
rect 163 -68 206 -67
rect 47 -70 76 -69
rect 93 -70 111 -69
rect 131 -70 171 -69
rect 177 -70 248 -69
rect 51 -72 80 -71
rect 93 -72 122 -71
rect 128 -72 171 -71
rect 191 -72 227 -71
rect 54 -74 69 -73
rect 79 -74 87 -73
rect 100 -74 150 -73
rect 58 -76 90 -75
rect 114 -76 132 -75
rect 135 -76 213 -75
rect 86 -78 164 -77
rect 100 -80 115 -79
rect 128 -80 199 -79
rect 107 -82 136 -81
rect 142 -82 178 -81
rect 121 -84 143 -83
rect 2 -95 101 -94
rect 114 -95 132 -94
rect 142 -95 220 -94
rect 233 -95 251 -94
rect 9 -97 52 -96
rect 58 -97 76 -96
rect 79 -97 87 -96
rect 107 -97 115 -96
rect 124 -97 129 -96
rect 145 -97 206 -96
rect 212 -97 234 -96
rect 240 -97 255 -96
rect 23 -99 45 -98
rect 47 -99 90 -98
rect 145 -99 220 -98
rect 30 -101 104 -100
rect 152 -101 178 -100
rect 184 -101 206 -100
rect 51 -103 69 -102
rect 72 -103 150 -102
rect 184 -103 248 -102
rect 86 -105 94 -104
rect 135 -105 178 -104
rect 191 -105 227 -104
rect 82 -107 192 -106
rect 194 -107 213 -106
rect 93 -109 118 -108
rect 121 -109 136 -108
rect 198 -109 227 -108
rect 121 -111 248 -110
rect 159 -113 199 -112
rect 2 -124 41 -123
rect 58 -124 66 -123
rect 79 -124 206 -123
rect 212 -124 269 -123
rect 2 -126 52 -125
rect 86 -126 220 -125
rect 9 -128 83 -127
rect 89 -128 255 -127
rect 19 -130 38 -129
rect 47 -130 90 -129
rect 93 -130 143 -129
rect 149 -130 227 -129
rect 19 -132 41 -131
rect 51 -132 59 -131
rect 100 -132 213 -131
rect 219 -132 241 -131
rect 23 -134 34 -133
rect 100 -134 108 -133
rect 114 -134 234 -133
rect 30 -136 69 -135
rect 72 -136 115 -135
rect 117 -136 234 -135
rect 9 -138 31 -137
rect 107 -138 129 -137
rect 135 -138 206 -137
rect 226 -138 276 -137
rect 121 -140 171 -139
rect 187 -140 248 -139
rect 121 -142 146 -141
rect 149 -142 164 -141
rect 128 -144 178 -143
rect 135 -146 171 -145
rect 177 -146 192 -145
rect 138 -148 248 -147
rect 152 -150 241 -149
rect 156 -152 192 -151
rect 159 -154 262 -153
rect 163 -156 199 -155
rect 184 -158 199 -157
rect 2 -169 87 -168
rect 96 -169 143 -168
rect 149 -169 157 -168
rect 159 -169 199 -168
rect 9 -171 48 -170
rect 58 -171 66 -170
rect 82 -171 90 -170
rect 100 -171 104 -170
rect 107 -171 115 -170
rect 117 -171 234 -170
rect 23 -173 153 -172
rect 170 -173 199 -172
rect 212 -173 234 -172
rect 26 -175 73 -174
rect 79 -175 83 -174
rect 128 -175 139 -174
rect 149 -175 269 -174
rect 40 -177 45 -176
rect 51 -177 59 -176
rect 65 -177 115 -176
rect 128 -177 255 -176
rect 30 -179 41 -178
rect 51 -179 108 -178
rect 135 -179 206 -178
rect 212 -179 227 -178
rect 254 -179 276 -178
rect 72 -181 111 -180
rect 135 -181 262 -180
rect 86 -183 139 -182
rect 163 -183 171 -182
rect 184 -183 227 -182
rect 163 -185 178 -184
rect 187 -185 262 -184
rect 177 -187 195 -186
rect 191 -189 206 -188
rect 23 -200 83 -199
rect 93 -200 153 -199
rect 184 -200 195 -199
rect 282 -200 290 -199
rect 37 -202 59 -201
rect 68 -202 104 -201
rect 110 -202 164 -201
rect 187 -202 206 -201
rect 278 -202 283 -201
rect 37 -204 73 -203
rect 100 -204 129 -203
rect 135 -204 157 -203
rect 191 -204 234 -203
rect 44 -206 241 -205
rect 51 -208 97 -207
rect 117 -208 122 -207
rect 135 -208 146 -207
rect 152 -208 255 -207
rect 44 -210 52 -209
rect 58 -210 94 -209
rect 114 -210 122 -209
rect 138 -210 234 -209
rect 254 -210 272 -209
rect 65 -212 97 -211
rect 117 -212 171 -211
rect 198 -212 206 -211
rect 219 -212 241 -211
rect 86 -214 129 -213
rect 142 -214 227 -213
rect 86 -216 160 -215
rect 180 -216 227 -215
rect 107 -218 143 -217
rect 149 -218 171 -217
rect 194 -218 220 -217
rect 47 -220 108 -219
rect 149 -220 164 -219
rect 198 -220 262 -219
rect 247 -222 262 -221
rect 247 -224 265 -223
rect 16 -235 45 -234
rect 58 -235 76 -234
rect 93 -235 129 -234
rect 156 -235 255 -234
rect 275 -235 290 -234
rect 30 -237 118 -236
rect 128 -237 136 -236
rect 159 -237 234 -236
rect 240 -237 265 -236
rect 37 -239 115 -238
rect 173 -239 185 -238
rect 219 -239 234 -238
rect 240 -239 262 -238
rect 37 -241 80 -240
rect 93 -241 118 -240
rect 184 -241 199 -240
rect 205 -241 220 -240
rect 247 -241 255 -240
rect 58 -243 101 -242
rect 103 -243 143 -242
rect 163 -243 206 -242
rect 65 -245 80 -244
rect 107 -245 164 -244
rect 177 -245 199 -244
rect 51 -247 66 -246
rect 72 -247 87 -246
rect 107 -247 150 -246
rect 180 -247 248 -246
rect 86 -249 115 -248
rect 121 -249 143 -248
rect 121 -251 192 -250
rect 170 -253 192 -252
rect 156 -255 171 -254
rect 26 -266 45 -265
rect 47 -266 66 -265
rect 86 -266 104 -265
rect 114 -266 206 -265
rect 208 -266 227 -265
rect 282 -266 290 -265
rect 16 -268 87 -267
rect 89 -268 129 -267
rect 135 -268 185 -267
rect 191 -268 213 -267
rect 30 -270 97 -269
rect 103 -270 143 -269
rect 170 -270 178 -269
rect 180 -270 220 -269
rect 37 -272 108 -271
rect 128 -272 157 -271
rect 173 -272 248 -271
rect 51 -274 192 -273
rect 194 -274 241 -273
rect 54 -276 73 -275
rect 93 -276 108 -275
rect 135 -276 164 -275
rect 205 -276 234 -275
rect 240 -276 248 -275
rect 58 -278 118 -277
rect 149 -278 157 -277
rect 65 -280 94 -279
rect 100 -280 143 -279
rect 149 -280 167 -279
rect 72 -282 80 -281
rect 51 -293 115 -292
rect 117 -293 122 -292
rect 138 -293 206 -292
rect 219 -293 234 -292
rect 250 -293 255 -292
rect 65 -295 83 -294
rect 107 -295 122 -294
rect 142 -295 178 -294
rect 184 -295 195 -294
rect 65 -297 115 -296
rect 117 -297 143 -296
rect 156 -297 164 -296
rect 191 -297 199 -296
rect 72 -299 104 -298
rect 149 -299 164 -298
rect 75 -301 87 -300
rect 89 -301 108 -300
rect 110 -301 150 -300
rect 82 -303 87 -302
rect 96 -303 157 -302
rect 89 -305 97 -304
rect 103 -305 136 -304
rect 44 -316 90 -315
rect 96 -316 136 -315
rect 159 -316 171 -315
rect 177 -316 206 -315
rect 226 -316 234 -315
rect 236 -316 241 -315
rect 51 -318 90 -317
rect 107 -318 129 -317
rect 138 -318 171 -317
rect 51 -320 94 -319
rect 107 -320 122 -319
rect 128 -320 157 -319
rect 61 -322 66 -321
rect 72 -322 118 -321
rect 138 -322 192 -321
rect 61 -324 76 -323
rect 79 -324 199 -323
rect 65 -326 87 -325
rect 93 -326 101 -325
rect 114 -326 164 -325
rect 37 -328 101 -327
rect 117 -328 122 -327
rect 135 -328 164 -327
rect 72 -330 143 -329
rect 149 -330 178 -329
rect 131 -332 150 -331
rect 142 -334 185 -333
rect 37 -345 80 -344
rect 100 -345 164 -344
rect 194 -345 199 -344
rect 215 -345 220 -344
rect 44 -347 118 -346
rect 135 -347 143 -346
rect 145 -347 206 -346
rect 58 -349 94 -348
rect 110 -349 213 -348
rect 51 -351 59 -350
rect 72 -351 139 -350
rect 149 -351 164 -350
rect 177 -351 199 -350
rect 72 -353 97 -352
rect 114 -353 171 -352
rect 177 -353 192 -352
rect 79 -355 108 -354
rect 149 -355 157 -354
rect 170 -355 185 -354
rect 86 -357 143 -356
rect 96 -359 104 -358
rect 131 -359 185 -358
rect 103 -361 129 -360
rect 58 -372 125 -371
rect 135 -372 143 -371
rect 145 -372 185 -371
rect 65 -374 108 -373
rect 138 -374 150 -373
rect 156 -374 199 -373
rect 72 -376 101 -375
rect 103 -376 129 -375
rect 142 -376 164 -375
rect 170 -376 178 -375
rect 72 -378 97 -377
rect 100 -378 108 -377
rect 114 -378 157 -377
rect 79 -380 118 -379
rect 121 -380 129 -379
rect 149 -380 174 -379
rect 79 -382 94 -381
rect 121 -382 164 -381
rect 79 -395 101 -394
rect 114 -395 129 -394
rect 131 -395 150 -394
rect 170 -395 174 -394
rect 72 -397 129 -396
rect 145 -397 157 -396
rect 86 -399 139 -398
rect 79 -401 87 -400
rect 93 -401 108 -400
rect 121 -401 143 -400
rect 117 -403 122 -402
rect 142 -403 164 -402
rect 107 -405 118 -404
rect 156 -405 164 -404
rect 93 -416 101 -415
rect 117 -416 122 -415
rect 156 -416 164 -415
rect 86 -418 94 -417
rect 107 -418 122 -417
rect 89 -429 94 -428
rect 117 -429 122 -428
rect 163 -429 171 -428
<< m2contact >>
rect 93 0 94 1
rect 103 0 104 1
rect 177 0 178 1
rect 184 0 185 1
rect 191 0 192 1
rect 198 0 199 1
rect 100 -2 101 -1
rect 114 -2 115 -1
rect 58 -13 59 -12
rect 68 -13 69 -12
rect 79 -13 80 -12
rect 89 -13 90 -12
rect 93 -13 94 -12
rect 107 -13 108 -12
rect 117 -13 118 -12
rect 128 -13 129 -12
rect 184 -13 185 -12
rect 191 -13 192 -12
rect 198 -13 199 -12
rect 205 -13 206 -12
rect 93 -15 94 -14
rect 100 -15 101 -14
rect 107 -15 108 -14
rect 114 -15 115 -14
rect 177 -15 178 -14
rect 184 -15 185 -14
rect 79 -26 80 -25
rect 86 -26 87 -25
rect 93 -26 94 -25
rect 107 -26 108 -25
rect 142 -26 143 -25
rect 149 -26 150 -25
rect 170 -26 171 -25
rect 177 -26 178 -25
rect 180 -26 181 -25
rect 184 -26 185 -25
rect 198 -26 199 -25
rect 205 -26 206 -25
rect 51 -28 52 -27
rect 93 -28 94 -27
rect 96 -28 97 -27
rect 156 -28 157 -27
rect 65 -30 66 -29
rect 79 -30 80 -29
rect 100 -30 101 -29
rect 121 -30 122 -29
rect 58 -32 59 -31
rect 65 -32 66 -31
rect 58 -34 59 -33
rect 117 -34 118 -33
rect 44 -45 45 -44
rect 51 -45 52 -44
rect 58 -45 59 -44
rect 79 -45 80 -44
rect 86 -45 87 -44
rect 114 -45 115 -44
rect 138 -45 139 -44
rect 149 -45 150 -44
rect 159 -45 160 -44
rect 191 -45 192 -44
rect 30 -47 31 -46
rect 79 -47 80 -46
rect 103 -47 104 -46
rect 121 -47 122 -46
rect 142 -47 143 -46
rect 163 -47 164 -46
rect 170 -47 171 -46
rect 177 -47 178 -46
rect 37 -49 38 -48
rect 103 -49 104 -48
rect 107 -49 108 -48
rect 128 -49 129 -48
rect 152 -49 153 -48
rect 170 -49 171 -48
rect 51 -51 52 -50
rect 65 -51 66 -50
rect 68 -51 69 -50
rect 86 -51 87 -50
rect 107 -51 108 -50
rect 114 -51 115 -50
rect 117 -51 118 -50
rect 177 -51 178 -50
rect 58 -53 59 -52
rect 72 -53 73 -52
rect 75 -53 76 -52
rect 93 -53 94 -52
rect 110 -53 111 -52
rect 142 -53 143 -52
rect 121 -55 122 -54
rect 131 -55 132 -54
rect 30 -66 31 -65
rect 72 -66 73 -65
rect 82 -66 83 -65
rect 184 -66 185 -65
rect 187 -66 188 -65
rect 219 -66 220 -65
rect 233 -66 234 -65
rect 243 -66 244 -65
rect 37 -68 38 -67
rect 65 -68 66 -67
rect 72 -68 73 -67
rect 138 -68 139 -67
rect 152 -68 153 -67
rect 156 -68 157 -67
rect 163 -68 164 -67
rect 205 -68 206 -67
rect 47 -70 48 -69
rect 75 -70 76 -69
rect 93 -70 94 -69
rect 110 -70 111 -69
rect 131 -70 132 -69
rect 170 -70 171 -69
rect 177 -70 178 -69
rect 247 -70 248 -69
rect 51 -72 52 -71
rect 79 -72 80 -71
rect 93 -72 94 -71
rect 121 -72 122 -71
rect 128 -72 129 -71
rect 170 -72 171 -71
rect 191 -72 192 -71
rect 226 -72 227 -71
rect 54 -74 55 -73
rect 68 -74 69 -73
rect 79 -74 80 -73
rect 86 -74 87 -73
rect 100 -74 101 -73
rect 149 -74 150 -73
rect 58 -76 59 -75
rect 89 -76 90 -75
rect 114 -76 115 -75
rect 131 -76 132 -75
rect 135 -76 136 -75
rect 212 -76 213 -75
rect 86 -78 87 -77
rect 163 -78 164 -77
rect 100 -80 101 -79
rect 114 -80 115 -79
rect 128 -80 129 -79
rect 198 -80 199 -79
rect 107 -82 108 -81
rect 135 -82 136 -81
rect 142 -82 143 -81
rect 177 -82 178 -81
rect 121 -84 122 -83
rect 142 -84 143 -83
rect 2 -95 3 -94
rect 100 -95 101 -94
rect 114 -95 115 -94
rect 131 -95 132 -94
rect 142 -95 143 -94
rect 219 -95 220 -94
rect 233 -95 234 -94
rect 250 -95 251 -94
rect 9 -97 10 -96
rect 51 -97 52 -96
rect 58 -97 59 -96
rect 75 -97 76 -96
rect 79 -97 80 -96
rect 86 -97 87 -96
rect 107 -97 108 -96
rect 114 -97 115 -96
rect 124 -97 125 -96
rect 128 -97 129 -96
rect 145 -97 146 -96
rect 205 -97 206 -96
rect 212 -97 213 -96
rect 233 -97 234 -96
rect 240 -97 241 -96
rect 254 -97 255 -96
rect 23 -99 24 -98
rect 44 -99 45 -98
rect 47 -99 48 -98
rect 89 -99 90 -98
rect 145 -99 146 -98
rect 219 -99 220 -98
rect 30 -101 31 -100
rect 103 -101 104 -100
rect 152 -101 153 -100
rect 177 -101 178 -100
rect 184 -101 185 -100
rect 205 -101 206 -100
rect 51 -103 52 -102
rect 68 -103 69 -102
rect 72 -103 73 -102
rect 149 -103 150 -102
rect 184 -103 185 -102
rect 247 -103 248 -102
rect 86 -105 87 -104
rect 93 -105 94 -104
rect 135 -105 136 -104
rect 177 -105 178 -104
rect 191 -105 192 -104
rect 226 -105 227 -104
rect 82 -107 83 -106
rect 191 -107 192 -106
rect 194 -107 195 -106
rect 212 -107 213 -106
rect 93 -109 94 -108
rect 117 -109 118 -108
rect 121 -109 122 -108
rect 135 -109 136 -108
rect 198 -109 199 -108
rect 226 -109 227 -108
rect 121 -111 122 -110
rect 247 -111 248 -110
rect 159 -113 160 -112
rect 198 -113 199 -112
rect 2 -124 3 -123
rect 40 -124 41 -123
rect 58 -124 59 -123
rect 65 -124 66 -123
rect 79 -124 80 -123
rect 205 -124 206 -123
rect 212 -124 213 -123
rect 268 -124 269 -123
rect 2 -126 3 -125
rect 51 -126 52 -125
rect 86 -126 87 -125
rect 219 -126 220 -125
rect 9 -128 10 -127
rect 82 -128 83 -127
rect 89 -128 90 -127
rect 254 -128 255 -127
rect 19 -130 20 -129
rect 37 -130 38 -129
rect 47 -130 48 -129
rect 89 -130 90 -129
rect 93 -130 94 -129
rect 142 -130 143 -129
rect 149 -130 150 -129
rect 226 -130 227 -129
rect 19 -132 20 -131
rect 40 -132 41 -131
rect 51 -132 52 -131
rect 58 -132 59 -131
rect 100 -132 101 -131
rect 212 -132 213 -131
rect 219 -132 220 -131
rect 240 -132 241 -131
rect 23 -134 24 -133
rect 33 -134 34 -133
rect 100 -134 101 -133
rect 107 -134 108 -133
rect 114 -134 115 -133
rect 233 -134 234 -133
rect 30 -136 31 -135
rect 68 -136 69 -135
rect 72 -136 73 -135
rect 114 -136 115 -135
rect 117 -136 118 -135
rect 233 -136 234 -135
rect 9 -138 10 -137
rect 30 -138 31 -137
rect 107 -138 108 -137
rect 128 -138 129 -137
rect 135 -138 136 -137
rect 205 -138 206 -137
rect 226 -138 227 -137
rect 275 -138 276 -137
rect 121 -140 122 -139
rect 170 -140 171 -139
rect 187 -140 188 -139
rect 247 -140 248 -139
rect 121 -142 122 -141
rect 145 -142 146 -141
rect 149 -142 150 -141
rect 163 -142 164 -141
rect 128 -144 129 -143
rect 177 -144 178 -143
rect 135 -146 136 -145
rect 170 -146 171 -145
rect 177 -146 178 -145
rect 191 -146 192 -145
rect 138 -148 139 -147
rect 247 -148 248 -147
rect 152 -150 153 -149
rect 240 -150 241 -149
rect 156 -152 157 -151
rect 191 -152 192 -151
rect 159 -154 160 -153
rect 261 -154 262 -153
rect 163 -156 164 -155
rect 198 -156 199 -155
rect 184 -158 185 -157
rect 198 -158 199 -157
rect 2 -169 3 -168
rect 86 -169 87 -168
rect 96 -169 97 -168
rect 142 -169 143 -168
rect 149 -169 150 -168
rect 156 -169 157 -168
rect 159 -169 160 -168
rect 198 -169 199 -168
rect 9 -171 10 -170
rect 47 -171 48 -170
rect 58 -171 59 -170
rect 65 -171 66 -170
rect 82 -171 83 -170
rect 89 -171 90 -170
rect 100 -171 101 -170
rect 103 -171 104 -170
rect 107 -171 108 -170
rect 114 -171 115 -170
rect 117 -171 118 -170
rect 233 -171 234 -170
rect 23 -173 24 -172
rect 152 -173 153 -172
rect 170 -173 171 -172
rect 198 -173 199 -172
rect 212 -173 213 -172
rect 233 -173 234 -172
rect 26 -175 27 -174
rect 72 -175 73 -174
rect 79 -175 80 -174
rect 82 -175 83 -174
rect 128 -175 129 -174
rect 138 -175 139 -174
rect 149 -175 150 -174
rect 268 -175 269 -174
rect 40 -177 41 -176
rect 44 -177 45 -176
rect 51 -177 52 -176
rect 58 -177 59 -176
rect 65 -177 66 -176
rect 114 -177 115 -176
rect 128 -177 129 -176
rect 254 -177 255 -176
rect 30 -179 31 -178
rect 40 -179 41 -178
rect 51 -179 52 -178
rect 107 -179 108 -178
rect 135 -179 136 -178
rect 205 -179 206 -178
rect 212 -179 213 -178
rect 226 -179 227 -178
rect 254 -179 255 -178
rect 275 -179 276 -178
rect 72 -181 73 -180
rect 110 -181 111 -180
rect 135 -181 136 -180
rect 261 -181 262 -180
rect 86 -183 87 -182
rect 138 -183 139 -182
rect 163 -183 164 -182
rect 170 -183 171 -182
rect 184 -183 185 -182
rect 226 -183 227 -182
rect 163 -185 164 -184
rect 177 -185 178 -184
rect 187 -185 188 -184
rect 261 -185 262 -184
rect 177 -187 178 -186
rect 194 -187 195 -186
rect 191 -189 192 -188
rect 205 -189 206 -188
rect 23 -200 24 -199
rect 82 -200 83 -199
rect 93 -200 94 -199
rect 152 -200 153 -199
rect 184 -200 185 -199
rect 194 -200 195 -199
rect 282 -200 283 -199
rect 289 -200 290 -199
rect 37 -202 38 -201
rect 58 -202 59 -201
rect 68 -202 69 -201
rect 103 -202 104 -201
rect 110 -202 111 -201
rect 163 -202 164 -201
rect 187 -202 188 -201
rect 205 -202 206 -201
rect 278 -202 279 -201
rect 282 -202 283 -201
rect 37 -204 38 -203
rect 72 -204 73 -203
rect 100 -204 101 -203
rect 128 -204 129 -203
rect 135 -204 136 -203
rect 156 -204 157 -203
rect 191 -204 192 -203
rect 233 -204 234 -203
rect 44 -206 45 -205
rect 240 -206 241 -205
rect 51 -208 52 -207
rect 96 -208 97 -207
rect 117 -208 118 -207
rect 121 -208 122 -207
rect 135 -208 136 -207
rect 145 -208 146 -207
rect 152 -208 153 -207
rect 254 -208 255 -207
rect 44 -210 45 -209
rect 51 -210 52 -209
rect 58 -210 59 -209
rect 93 -210 94 -209
rect 114 -210 115 -209
rect 121 -210 122 -209
rect 138 -210 139 -209
rect 233 -210 234 -209
rect 254 -210 255 -209
rect 271 -210 272 -209
rect 65 -212 66 -211
rect 96 -212 97 -211
rect 117 -212 118 -211
rect 170 -212 171 -211
rect 198 -212 199 -211
rect 205 -212 206 -211
rect 219 -212 220 -211
rect 240 -212 241 -211
rect 86 -214 87 -213
rect 128 -214 129 -213
rect 142 -214 143 -213
rect 226 -214 227 -213
rect 86 -216 87 -215
rect 159 -216 160 -215
rect 180 -216 181 -215
rect 226 -216 227 -215
rect 107 -218 108 -217
rect 142 -218 143 -217
rect 149 -218 150 -217
rect 170 -218 171 -217
rect 194 -218 195 -217
rect 219 -218 220 -217
rect 47 -220 48 -219
rect 107 -220 108 -219
rect 149 -220 150 -219
rect 163 -220 164 -219
rect 198 -220 199 -219
rect 261 -220 262 -219
rect 247 -222 248 -221
rect 261 -222 262 -221
rect 247 -224 248 -223
rect 264 -224 265 -223
rect 16 -235 17 -234
rect 44 -235 45 -234
rect 58 -235 59 -234
rect 75 -235 76 -234
rect 93 -235 94 -234
rect 128 -235 129 -234
rect 156 -235 157 -234
rect 254 -235 255 -234
rect 275 -235 276 -234
rect 289 -235 290 -234
rect 30 -237 31 -236
rect 117 -237 118 -236
rect 128 -237 129 -236
rect 135 -237 136 -236
rect 159 -237 160 -236
rect 233 -237 234 -236
rect 240 -237 241 -236
rect 264 -237 265 -236
rect 37 -239 38 -238
rect 114 -239 115 -238
rect 173 -239 174 -238
rect 184 -239 185 -238
rect 219 -239 220 -238
rect 233 -239 234 -238
rect 240 -239 241 -238
rect 261 -239 262 -238
rect 37 -241 38 -240
rect 79 -241 80 -240
rect 93 -241 94 -240
rect 117 -241 118 -240
rect 184 -241 185 -240
rect 198 -241 199 -240
rect 205 -241 206 -240
rect 219 -241 220 -240
rect 247 -241 248 -240
rect 254 -241 255 -240
rect 58 -243 59 -242
rect 100 -243 101 -242
rect 103 -243 104 -242
rect 142 -243 143 -242
rect 163 -243 164 -242
rect 205 -243 206 -242
rect 65 -245 66 -244
rect 79 -245 80 -244
rect 107 -245 108 -244
rect 163 -245 164 -244
rect 177 -245 178 -244
rect 198 -245 199 -244
rect 51 -247 52 -246
rect 65 -247 66 -246
rect 72 -247 73 -246
rect 86 -247 87 -246
rect 107 -247 108 -246
rect 149 -247 150 -246
rect 180 -247 181 -246
rect 247 -247 248 -246
rect 86 -249 87 -248
rect 114 -249 115 -248
rect 121 -249 122 -248
rect 142 -249 143 -248
rect 121 -251 122 -250
rect 191 -251 192 -250
rect 170 -253 171 -252
rect 191 -253 192 -252
rect 156 -255 157 -254
rect 170 -255 171 -254
rect 26 -266 27 -265
rect 44 -266 45 -265
rect 47 -266 48 -265
rect 65 -266 66 -265
rect 86 -266 87 -265
rect 103 -266 104 -265
rect 114 -266 115 -265
rect 205 -266 206 -265
rect 208 -266 209 -265
rect 226 -266 227 -265
rect 282 -266 283 -265
rect 289 -266 290 -265
rect 16 -268 17 -267
rect 86 -268 87 -267
rect 89 -268 90 -267
rect 128 -268 129 -267
rect 135 -268 136 -267
rect 184 -268 185 -267
rect 191 -268 192 -267
rect 212 -268 213 -267
rect 30 -270 31 -269
rect 96 -270 97 -269
rect 103 -270 104 -269
rect 142 -270 143 -269
rect 170 -270 171 -269
rect 177 -270 178 -269
rect 180 -270 181 -269
rect 219 -270 220 -269
rect 37 -272 38 -271
rect 107 -272 108 -271
rect 128 -272 129 -271
rect 156 -272 157 -271
rect 173 -272 174 -271
rect 247 -272 248 -271
rect 51 -274 52 -273
rect 191 -274 192 -273
rect 194 -274 195 -273
rect 240 -274 241 -273
rect 54 -276 55 -275
rect 72 -276 73 -275
rect 93 -276 94 -275
rect 107 -276 108 -275
rect 135 -276 136 -275
rect 163 -276 164 -275
rect 205 -276 206 -275
rect 233 -276 234 -275
rect 240 -276 241 -275
rect 247 -276 248 -275
rect 58 -278 59 -277
rect 117 -278 118 -277
rect 149 -278 150 -277
rect 156 -278 157 -277
rect 65 -280 66 -279
rect 93 -280 94 -279
rect 100 -280 101 -279
rect 142 -280 143 -279
rect 149 -280 150 -279
rect 166 -280 167 -279
rect 72 -282 73 -281
rect 79 -282 80 -281
rect 51 -293 52 -292
rect 114 -293 115 -292
rect 117 -293 118 -292
rect 121 -293 122 -292
rect 138 -293 139 -292
rect 205 -293 206 -292
rect 219 -293 220 -292
rect 233 -293 234 -292
rect 250 -293 251 -292
rect 254 -293 255 -292
rect 65 -295 66 -294
rect 82 -295 83 -294
rect 107 -295 108 -294
rect 121 -295 122 -294
rect 142 -295 143 -294
rect 177 -295 178 -294
rect 184 -295 185 -294
rect 194 -295 195 -294
rect 65 -297 66 -296
rect 114 -297 115 -296
rect 117 -297 118 -296
rect 142 -297 143 -296
rect 156 -297 157 -296
rect 163 -297 164 -296
rect 191 -297 192 -296
rect 198 -297 199 -296
rect 72 -299 73 -298
rect 103 -299 104 -298
rect 149 -299 150 -298
rect 163 -299 164 -298
rect 75 -301 76 -300
rect 86 -301 87 -300
rect 89 -301 90 -300
rect 107 -301 108 -300
rect 110 -301 111 -300
rect 149 -301 150 -300
rect 82 -303 83 -302
rect 86 -303 87 -302
rect 96 -303 97 -302
rect 156 -303 157 -302
rect 89 -305 90 -304
rect 96 -305 97 -304
rect 103 -305 104 -304
rect 135 -305 136 -304
rect 44 -316 45 -315
rect 89 -316 90 -315
rect 96 -316 97 -315
rect 135 -316 136 -315
rect 159 -316 160 -315
rect 170 -316 171 -315
rect 177 -316 178 -315
rect 205 -316 206 -315
rect 226 -316 227 -315
rect 233 -316 234 -315
rect 236 -316 237 -315
rect 240 -316 241 -315
rect 51 -318 52 -317
rect 89 -318 90 -317
rect 107 -318 108 -317
rect 128 -318 129 -317
rect 138 -318 139 -317
rect 170 -318 171 -317
rect 51 -320 52 -319
rect 93 -320 94 -319
rect 107 -320 108 -319
rect 121 -320 122 -319
rect 128 -320 129 -319
rect 156 -320 157 -319
rect 61 -322 62 -321
rect 65 -322 66 -321
rect 72 -322 73 -321
rect 117 -322 118 -321
rect 138 -322 139 -321
rect 191 -322 192 -321
rect 61 -324 62 -323
rect 75 -324 76 -323
rect 79 -324 80 -323
rect 198 -324 199 -323
rect 65 -326 66 -325
rect 86 -326 87 -325
rect 93 -326 94 -325
rect 100 -326 101 -325
rect 114 -326 115 -325
rect 163 -326 164 -325
rect 37 -328 38 -327
rect 100 -328 101 -327
rect 117 -328 118 -327
rect 121 -328 122 -327
rect 135 -328 136 -327
rect 163 -328 164 -327
rect 72 -330 73 -329
rect 142 -330 143 -329
rect 149 -330 150 -329
rect 177 -330 178 -329
rect 131 -332 132 -331
rect 149 -332 150 -331
rect 142 -334 143 -333
rect 184 -334 185 -333
rect 37 -345 38 -344
rect 79 -345 80 -344
rect 100 -345 101 -344
rect 163 -345 164 -344
rect 194 -345 195 -344
rect 198 -345 199 -344
rect 215 -345 216 -344
rect 219 -345 220 -344
rect 44 -347 45 -346
rect 117 -347 118 -346
rect 135 -347 136 -346
rect 142 -347 143 -346
rect 145 -347 146 -346
rect 205 -347 206 -346
rect 58 -349 59 -348
rect 93 -349 94 -348
rect 110 -349 111 -348
rect 212 -349 213 -348
rect 51 -351 52 -350
rect 58 -351 59 -350
rect 72 -351 73 -350
rect 138 -351 139 -350
rect 149 -351 150 -350
rect 163 -351 164 -350
rect 177 -351 178 -350
rect 198 -351 199 -350
rect 72 -353 73 -352
rect 96 -353 97 -352
rect 114 -353 115 -352
rect 170 -353 171 -352
rect 177 -353 178 -352
rect 191 -353 192 -352
rect 79 -355 80 -354
rect 107 -355 108 -354
rect 149 -355 150 -354
rect 156 -355 157 -354
rect 170 -355 171 -354
rect 184 -355 185 -354
rect 86 -357 87 -356
rect 142 -357 143 -356
rect 96 -359 97 -358
rect 103 -359 104 -358
rect 131 -359 132 -358
rect 184 -359 185 -358
rect 103 -361 104 -360
rect 128 -361 129 -360
rect 58 -372 59 -371
rect 124 -372 125 -371
rect 135 -372 136 -371
rect 142 -372 143 -371
rect 145 -372 146 -371
rect 184 -372 185 -371
rect 65 -374 66 -373
rect 107 -374 108 -373
rect 138 -374 139 -373
rect 149 -374 150 -373
rect 156 -374 157 -373
rect 198 -374 199 -373
rect 72 -376 73 -375
rect 100 -376 101 -375
rect 103 -376 104 -375
rect 128 -376 129 -375
rect 142 -376 143 -375
rect 163 -376 164 -375
rect 170 -376 171 -375
rect 177 -376 178 -375
rect 72 -378 73 -377
rect 96 -378 97 -377
rect 100 -378 101 -377
rect 107 -378 108 -377
rect 114 -378 115 -377
rect 156 -378 157 -377
rect 79 -380 80 -379
rect 117 -380 118 -379
rect 121 -380 122 -379
rect 128 -380 129 -379
rect 149 -380 150 -379
rect 173 -380 174 -379
rect 79 -382 80 -381
rect 93 -382 94 -381
rect 121 -382 122 -381
rect 163 -382 164 -381
rect 79 -395 80 -394
rect 100 -395 101 -394
rect 114 -395 115 -394
rect 128 -395 129 -394
rect 131 -395 132 -394
rect 149 -395 150 -394
rect 170 -395 171 -394
rect 173 -395 174 -394
rect 72 -397 73 -396
rect 128 -397 129 -396
rect 145 -397 146 -396
rect 156 -397 157 -396
rect 86 -399 87 -398
rect 138 -399 139 -398
rect 79 -401 80 -400
rect 86 -401 87 -400
rect 93 -401 94 -400
rect 107 -401 108 -400
rect 121 -401 122 -400
rect 142 -401 143 -400
rect 117 -403 118 -402
rect 121 -403 122 -402
rect 142 -403 143 -402
rect 163 -403 164 -402
rect 107 -405 108 -404
rect 117 -405 118 -404
rect 156 -405 157 -404
rect 163 -405 164 -404
rect 93 -416 94 -415
rect 100 -416 101 -415
rect 117 -416 118 -415
rect 121 -416 122 -415
rect 156 -416 157 -415
rect 163 -416 164 -415
rect 86 -418 87 -417
rect 93 -418 94 -417
rect 107 -418 108 -417
rect 121 -418 122 -417
rect 89 -429 90 -428
rect 93 -429 94 -428
rect 117 -429 118 -428
rect 121 -429 122 -428
rect 163 -429 164 -428
rect 170 -429 171 -428
<< metal2 >>
rect 93 -3 94 1
rect 103 -3 104 1
rect 177 -3 178 1
rect 184 -3 185 1
rect 191 -3 192 1
rect 198 -3 199 1
rect 100 -3 101 -1
rect 114 -3 115 -1
rect 58 -16 59 -12
rect 68 -16 69 -12
rect 75 -13 76 -11
rect 75 -16 76 -12
rect 75 -13 76 -11
rect 75 -16 76 -12
rect 79 -16 80 -12
rect 89 -16 90 -12
rect 93 -13 94 -11
rect 107 -13 108 -11
rect 117 -16 118 -12
rect 128 -16 129 -12
rect 184 -13 185 -11
rect 191 -13 192 -11
rect 198 -13 199 -11
rect 205 -16 206 -12
rect 93 -16 94 -14
rect 100 -16 101 -14
rect 107 -16 108 -14
rect 114 -15 115 -11
rect 177 -16 178 -14
rect 184 -16 185 -14
rect 79 -26 80 -24
rect 86 -35 87 -25
rect 93 -26 94 -24
rect 107 -35 108 -25
rect 128 -26 129 -24
rect 128 -35 129 -25
rect 128 -26 129 -24
rect 128 -35 129 -25
rect 142 -35 143 -25
rect 149 -35 150 -25
rect 170 -35 171 -25
rect 177 -26 178 -24
rect 180 -35 181 -25
rect 184 -35 185 -25
rect 198 -26 199 -24
rect 205 -26 206 -24
rect 51 -35 52 -27
rect 93 -35 94 -27
rect 96 -35 97 -27
rect 156 -35 157 -27
rect 65 -30 66 -24
rect 79 -35 80 -29
rect 100 -35 101 -29
rect 121 -35 122 -29
rect 58 -32 59 -24
rect 65 -35 66 -31
rect 58 -35 59 -33
rect 117 -35 118 -33
rect 44 -45 45 -43
rect 51 -45 52 -43
rect 58 -45 59 -43
rect 79 -45 80 -43
rect 86 -45 87 -43
rect 114 -45 115 -43
rect 138 -45 139 -43
rect 149 -56 150 -44
rect 156 -45 157 -43
rect 156 -56 157 -44
rect 156 -45 157 -43
rect 156 -56 157 -44
rect 159 -56 160 -44
rect 191 -56 192 -44
rect 30 -56 31 -46
rect 79 -56 80 -46
rect 103 -47 104 -43
rect 121 -47 122 -43
rect 142 -47 143 -43
rect 163 -56 164 -46
rect 170 -47 171 -43
rect 177 -47 178 -43
rect 184 -47 185 -43
rect 184 -56 185 -46
rect 184 -47 185 -43
rect 184 -56 185 -46
rect 37 -56 38 -48
rect 103 -56 104 -48
rect 107 -49 108 -43
rect 128 -49 129 -43
rect 152 -49 153 -43
rect 170 -56 171 -48
rect 51 -56 52 -50
rect 65 -51 66 -43
rect 68 -56 69 -50
rect 86 -56 87 -50
rect 107 -56 108 -50
rect 114 -56 115 -50
rect 117 -51 118 -43
rect 177 -56 178 -50
rect 58 -56 59 -52
rect 72 -53 73 -43
rect 75 -56 76 -52
rect 93 -56 94 -52
rect 110 -53 111 -43
rect 142 -56 143 -52
rect 121 -56 122 -54
rect 131 -56 132 -54
rect 30 -66 31 -64
rect 72 -66 73 -64
rect 82 -66 83 -64
rect 184 -85 185 -65
rect 187 -66 188 -64
rect 219 -85 220 -65
rect 233 -85 234 -65
rect 243 -85 244 -65
rect 37 -68 38 -64
rect 65 -85 66 -67
rect 72 -85 73 -67
rect 138 -68 139 -64
rect 152 -85 153 -67
rect 156 -85 157 -67
rect 163 -68 164 -64
rect 205 -85 206 -67
rect 47 -70 48 -64
rect 75 -70 76 -64
rect 93 -70 94 -64
rect 110 -85 111 -69
rect 131 -70 132 -64
rect 170 -70 171 -64
rect 177 -70 178 -64
rect 247 -85 248 -69
rect 51 -72 52 -64
rect 79 -72 80 -64
rect 93 -85 94 -71
rect 121 -72 122 -64
rect 128 -72 129 -64
rect 170 -85 171 -71
rect 191 -72 192 -64
rect 226 -85 227 -71
rect 54 -85 55 -73
rect 68 -85 69 -73
rect 79 -85 80 -73
rect 86 -74 87 -64
rect 100 -74 101 -64
rect 149 -74 150 -64
rect 58 -76 59 -64
rect 89 -85 90 -75
rect 114 -76 115 -64
rect 131 -85 132 -75
rect 135 -76 136 -64
rect 212 -85 213 -75
rect 86 -85 87 -77
rect 163 -85 164 -77
rect 100 -85 101 -79
rect 114 -85 115 -79
rect 128 -85 129 -79
rect 198 -85 199 -79
rect 107 -85 108 -81
rect 135 -85 136 -81
rect 142 -82 143 -64
rect 177 -85 178 -81
rect 121 -85 122 -83
rect 142 -85 143 -83
rect 2 -114 3 -94
rect 100 -114 101 -94
rect 114 -95 115 -93
rect 131 -95 132 -93
rect 142 -95 143 -93
rect 219 -95 220 -93
rect 233 -95 234 -93
rect 250 -95 251 -93
rect 9 -114 10 -96
rect 51 -97 52 -93
rect 58 -114 59 -96
rect 75 -114 76 -96
rect 79 -97 80 -93
rect 86 -97 87 -93
rect 107 -114 108 -96
rect 114 -114 115 -96
rect 124 -114 125 -96
rect 128 -114 129 -96
rect 145 -97 146 -93
rect 205 -97 206 -93
rect 212 -97 213 -93
rect 233 -114 234 -96
rect 240 -114 241 -96
rect 254 -114 255 -96
rect 23 -114 24 -98
rect 44 -114 45 -98
rect 47 -114 48 -98
rect 89 -99 90 -93
rect 145 -114 146 -98
rect 219 -114 220 -98
rect 30 -114 31 -100
rect 103 -101 104 -93
rect 152 -101 153 -93
rect 177 -101 178 -93
rect 184 -101 185 -93
rect 205 -114 206 -100
rect 51 -114 52 -102
rect 68 -114 69 -102
rect 72 -103 73 -93
rect 149 -114 150 -102
rect 156 -103 157 -93
rect 156 -114 157 -102
rect 156 -103 157 -93
rect 156 -114 157 -102
rect 163 -103 164 -93
rect 163 -114 164 -102
rect 163 -103 164 -93
rect 163 -114 164 -102
rect 170 -103 171 -93
rect 170 -114 171 -102
rect 170 -103 171 -93
rect 170 -114 171 -102
rect 184 -114 185 -102
rect 247 -103 248 -93
rect 86 -114 87 -104
rect 93 -105 94 -93
rect 135 -105 136 -93
rect 177 -114 178 -104
rect 191 -105 192 -93
rect 226 -105 227 -93
rect 82 -114 83 -106
rect 191 -114 192 -106
rect 194 -107 195 -93
rect 212 -114 213 -106
rect 93 -114 94 -108
rect 117 -114 118 -108
rect 121 -109 122 -93
rect 135 -114 136 -108
rect 198 -109 199 -93
rect 226 -114 227 -108
rect 121 -114 122 -110
rect 247 -114 248 -110
rect 159 -114 160 -112
rect 198 -114 199 -112
rect 2 -124 3 -122
rect 40 -124 41 -122
rect 58 -124 59 -122
rect 65 -159 66 -123
rect 79 -124 80 -122
rect 205 -124 206 -122
rect 212 -124 213 -122
rect 268 -159 269 -123
rect 2 -159 3 -125
rect 51 -126 52 -122
rect 86 -159 87 -125
rect 219 -126 220 -122
rect 9 -128 10 -122
rect 82 -128 83 -122
rect 89 -128 90 -122
rect 254 -159 255 -127
rect 19 -130 20 -122
rect 37 -130 38 -122
rect 47 -159 48 -129
rect 89 -159 90 -129
rect 93 -130 94 -122
rect 142 -159 143 -129
rect 149 -130 150 -122
rect 226 -130 227 -122
rect 19 -159 20 -131
rect 40 -159 41 -131
rect 51 -159 52 -131
rect 58 -159 59 -131
rect 100 -132 101 -122
rect 212 -159 213 -131
rect 219 -159 220 -131
rect 240 -132 241 -122
rect 23 -134 24 -122
rect 33 -159 34 -133
rect 100 -159 101 -133
rect 107 -134 108 -122
rect 114 -134 115 -122
rect 233 -134 234 -122
rect 30 -136 31 -122
rect 68 -136 69 -122
rect 72 -159 73 -135
rect 114 -159 115 -135
rect 117 -159 118 -135
rect 233 -159 234 -135
rect 9 -159 10 -137
rect 30 -159 31 -137
rect 107 -159 108 -137
rect 128 -138 129 -122
rect 135 -138 136 -122
rect 205 -159 206 -137
rect 226 -159 227 -137
rect 275 -159 276 -137
rect 121 -140 122 -122
rect 170 -140 171 -122
rect 187 -159 188 -139
rect 247 -140 248 -122
rect 121 -159 122 -141
rect 145 -142 146 -122
rect 149 -159 150 -141
rect 163 -142 164 -122
rect 128 -159 129 -143
rect 177 -144 178 -122
rect 135 -159 136 -145
rect 170 -159 171 -145
rect 177 -159 178 -145
rect 191 -146 192 -122
rect 138 -159 139 -147
rect 247 -159 248 -147
rect 152 -150 153 -122
rect 240 -159 241 -149
rect 156 -159 157 -151
rect 191 -159 192 -151
rect 159 -154 160 -122
rect 261 -159 262 -153
rect 163 -159 164 -155
rect 198 -156 199 -122
rect 184 -158 185 -122
rect 198 -159 199 -157
rect 2 -169 3 -167
rect 86 -169 87 -167
rect 96 -169 97 -167
rect 142 -169 143 -167
rect 149 -169 150 -167
rect 156 -190 157 -168
rect 159 -169 160 -167
rect 198 -169 199 -167
rect 219 -169 220 -167
rect 219 -190 220 -168
rect 219 -169 220 -167
rect 219 -190 220 -168
rect 240 -169 241 -167
rect 240 -190 241 -168
rect 240 -169 241 -167
rect 240 -190 241 -168
rect 247 -169 248 -167
rect 247 -190 248 -168
rect 247 -169 248 -167
rect 247 -190 248 -168
rect 9 -171 10 -167
rect 47 -171 48 -167
rect 58 -171 59 -167
rect 65 -171 66 -167
rect 82 -171 83 -167
rect 89 -171 90 -167
rect 100 -171 101 -167
rect 103 -190 104 -170
rect 107 -171 108 -167
rect 114 -171 115 -167
rect 117 -171 118 -167
rect 233 -171 234 -167
rect 23 -190 24 -172
rect 152 -190 153 -172
rect 170 -173 171 -167
rect 198 -190 199 -172
rect 212 -173 213 -167
rect 233 -190 234 -172
rect 26 -175 27 -167
rect 72 -175 73 -167
rect 79 -175 80 -167
rect 82 -190 83 -174
rect 121 -175 122 -167
rect 121 -190 122 -174
rect 121 -175 122 -167
rect 121 -190 122 -174
rect 128 -175 129 -167
rect 138 -175 139 -167
rect 149 -190 150 -174
rect 268 -175 269 -167
rect 40 -177 41 -167
rect 44 -190 45 -176
rect 51 -177 52 -167
rect 58 -190 59 -176
rect 65 -190 66 -176
rect 114 -190 115 -176
rect 128 -190 129 -176
rect 254 -177 255 -167
rect 30 -190 31 -178
rect 40 -190 41 -178
rect 51 -190 52 -178
rect 107 -190 108 -178
rect 135 -179 136 -167
rect 205 -179 206 -167
rect 212 -190 213 -178
rect 226 -179 227 -167
rect 254 -190 255 -178
rect 275 -179 276 -167
rect 72 -190 73 -180
rect 110 -181 111 -167
rect 135 -190 136 -180
rect 261 -181 262 -167
rect 86 -190 87 -182
rect 138 -190 139 -182
rect 163 -183 164 -167
rect 170 -190 171 -182
rect 184 -183 185 -167
rect 226 -190 227 -182
rect 163 -190 164 -184
rect 177 -185 178 -167
rect 187 -190 188 -184
rect 261 -190 262 -184
rect 177 -190 178 -186
rect 194 -190 195 -186
rect 191 -189 192 -167
rect 205 -190 206 -188
rect 23 -200 24 -198
rect 82 -225 83 -199
rect 93 -200 94 -198
rect 152 -200 153 -198
rect 177 -200 178 -198
rect 177 -225 178 -199
rect 177 -200 178 -198
rect 177 -225 178 -199
rect 184 -225 185 -199
rect 194 -200 195 -198
rect 212 -200 213 -198
rect 212 -225 213 -199
rect 212 -200 213 -198
rect 212 -225 213 -199
rect 282 -200 283 -198
rect 289 -225 290 -199
rect 30 -202 31 -198
rect 30 -225 31 -201
rect 30 -202 31 -198
rect 30 -225 31 -201
rect 37 -202 38 -198
rect 58 -202 59 -198
rect 68 -202 69 -198
rect 103 -202 104 -198
rect 110 -202 111 -198
rect 163 -202 164 -198
rect 187 -202 188 -198
rect 205 -202 206 -198
rect 278 -225 279 -201
rect 282 -225 283 -201
rect 37 -225 38 -203
rect 72 -204 73 -198
rect 100 -225 101 -203
rect 128 -204 129 -198
rect 135 -204 136 -198
rect 156 -204 157 -198
rect 191 -225 192 -203
rect 233 -204 234 -198
rect 44 -206 45 -198
rect 240 -206 241 -198
rect 51 -208 52 -198
rect 96 -208 97 -198
rect 117 -208 118 -198
rect 121 -208 122 -198
rect 135 -225 136 -207
rect 145 -208 146 -198
rect 152 -225 153 -207
rect 254 -208 255 -198
rect 44 -225 45 -209
rect 51 -225 52 -209
rect 58 -225 59 -209
rect 93 -225 94 -209
rect 114 -225 115 -209
rect 121 -225 122 -209
rect 138 -225 139 -209
rect 233 -225 234 -209
rect 254 -225 255 -209
rect 271 -225 272 -209
rect 65 -225 66 -211
rect 96 -225 97 -211
rect 117 -225 118 -211
rect 170 -212 171 -198
rect 198 -212 199 -198
rect 205 -225 206 -211
rect 219 -212 220 -198
rect 240 -225 241 -211
rect 86 -214 87 -198
rect 128 -225 129 -213
rect 142 -214 143 -198
rect 226 -214 227 -198
rect 86 -225 87 -215
rect 159 -225 160 -215
rect 180 -225 181 -215
rect 226 -225 227 -215
rect 107 -218 108 -198
rect 142 -225 143 -217
rect 149 -218 150 -198
rect 170 -225 171 -217
rect 194 -225 195 -217
rect 219 -225 220 -217
rect 47 -220 48 -198
rect 107 -225 108 -219
rect 149 -225 150 -219
rect 163 -225 164 -219
rect 198 -225 199 -219
rect 261 -220 262 -198
rect 247 -222 248 -198
rect 261 -225 262 -221
rect 247 -225 248 -223
rect 264 -225 265 -223
rect 16 -256 17 -234
rect 44 -256 45 -234
rect 58 -235 59 -233
rect 75 -235 76 -233
rect 93 -235 94 -233
rect 128 -235 129 -233
rect 156 -235 157 -233
rect 254 -235 255 -233
rect 275 -235 276 -233
rect 289 -235 290 -233
rect 30 -256 31 -236
rect 117 -237 118 -233
rect 128 -256 129 -236
rect 135 -256 136 -236
rect 159 -237 160 -233
rect 233 -237 234 -233
rect 240 -237 241 -233
rect 264 -237 265 -233
rect 282 -237 283 -233
rect 282 -256 283 -236
rect 282 -237 283 -233
rect 282 -256 283 -236
rect 37 -239 38 -233
rect 114 -239 115 -233
rect 173 -256 174 -238
rect 184 -239 185 -233
rect 212 -239 213 -233
rect 212 -256 213 -238
rect 212 -239 213 -233
rect 212 -256 213 -238
rect 219 -239 220 -233
rect 233 -256 234 -238
rect 240 -256 241 -238
rect 261 -239 262 -233
rect 37 -256 38 -240
rect 79 -241 80 -233
rect 93 -256 94 -240
rect 117 -256 118 -240
rect 184 -256 185 -240
rect 198 -241 199 -233
rect 205 -241 206 -233
rect 219 -256 220 -240
rect 226 -241 227 -233
rect 226 -256 227 -240
rect 226 -241 227 -233
rect 226 -256 227 -240
rect 247 -241 248 -233
rect 254 -256 255 -240
rect 58 -256 59 -242
rect 100 -243 101 -233
rect 103 -256 104 -242
rect 142 -243 143 -233
rect 163 -243 164 -233
rect 205 -256 206 -242
rect 65 -245 66 -233
rect 79 -256 80 -244
rect 107 -245 108 -233
rect 163 -256 164 -244
rect 177 -256 178 -244
rect 198 -256 199 -244
rect 51 -247 52 -233
rect 65 -256 66 -246
rect 72 -256 73 -246
rect 86 -247 87 -233
rect 107 -256 108 -246
rect 149 -256 150 -246
rect 180 -256 181 -246
rect 247 -256 248 -246
rect 86 -256 87 -248
rect 114 -256 115 -248
rect 121 -249 122 -233
rect 142 -256 143 -248
rect 121 -256 122 -250
rect 191 -251 192 -233
rect 170 -253 171 -233
rect 191 -256 192 -252
rect 156 -256 157 -254
rect 170 -256 171 -254
rect 26 -266 27 -264
rect 44 -266 45 -264
rect 47 -266 48 -264
rect 65 -266 66 -264
rect 86 -266 87 -264
rect 103 -266 104 -264
rect 114 -266 115 -264
rect 205 -266 206 -264
rect 208 -283 209 -265
rect 226 -266 227 -264
rect 254 -266 255 -264
rect 254 -283 255 -265
rect 254 -266 255 -264
rect 254 -283 255 -265
rect 282 -266 283 -264
rect 289 -266 290 -264
rect 16 -268 17 -264
rect 86 -283 87 -267
rect 89 -283 90 -267
rect 128 -268 129 -264
rect 135 -268 136 -264
rect 184 -268 185 -264
rect 191 -268 192 -264
rect 212 -268 213 -264
rect 30 -270 31 -264
rect 96 -283 97 -269
rect 103 -283 104 -269
rect 142 -270 143 -264
rect 170 -283 171 -269
rect 177 -270 178 -264
rect 180 -270 181 -264
rect 219 -270 220 -264
rect 37 -272 38 -264
rect 107 -272 108 -264
rect 121 -272 122 -264
rect 121 -283 122 -271
rect 121 -272 122 -264
rect 121 -283 122 -271
rect 128 -283 129 -271
rect 156 -272 157 -264
rect 173 -272 174 -264
rect 247 -272 248 -264
rect 51 -274 52 -264
rect 191 -283 192 -273
rect 194 -283 195 -273
rect 240 -274 241 -264
rect 54 -276 55 -264
rect 72 -276 73 -264
rect 93 -276 94 -264
rect 107 -283 108 -275
rect 135 -283 136 -275
rect 163 -276 164 -264
rect 198 -276 199 -264
rect 198 -283 199 -275
rect 198 -276 199 -264
rect 198 -283 199 -275
rect 205 -283 206 -275
rect 233 -276 234 -264
rect 240 -283 241 -275
rect 247 -283 248 -275
rect 58 -278 59 -264
rect 117 -278 118 -264
rect 149 -278 150 -264
rect 156 -283 157 -277
rect 65 -283 66 -279
rect 93 -283 94 -279
rect 100 -280 101 -264
rect 142 -283 143 -279
rect 149 -283 150 -279
rect 166 -283 167 -279
rect 72 -283 73 -281
rect 79 -282 80 -264
rect 51 -306 52 -292
rect 114 -293 115 -291
rect 117 -293 118 -291
rect 121 -293 122 -291
rect 128 -293 129 -291
rect 128 -306 129 -292
rect 128 -293 129 -291
rect 128 -306 129 -292
rect 138 -306 139 -292
rect 205 -293 206 -291
rect 219 -306 220 -292
rect 233 -306 234 -292
rect 240 -293 241 -291
rect 240 -306 241 -292
rect 240 -293 241 -291
rect 240 -306 241 -292
rect 250 -293 251 -291
rect 254 -293 255 -291
rect 65 -295 66 -291
rect 82 -295 83 -291
rect 107 -295 108 -291
rect 121 -306 122 -294
rect 142 -295 143 -291
rect 177 -306 178 -294
rect 184 -295 185 -291
rect 194 -295 195 -291
rect 65 -306 66 -296
rect 114 -306 115 -296
rect 117 -306 118 -296
rect 142 -306 143 -296
rect 156 -297 157 -291
rect 163 -297 164 -291
rect 170 -297 171 -291
rect 170 -306 171 -296
rect 170 -297 171 -291
rect 170 -306 171 -296
rect 191 -297 192 -291
rect 198 -297 199 -291
rect 72 -299 73 -291
rect 103 -299 104 -291
rect 149 -299 150 -291
rect 163 -306 164 -298
rect 75 -306 76 -300
rect 86 -301 87 -291
rect 89 -301 90 -291
rect 107 -306 108 -300
rect 110 -306 111 -300
rect 149 -306 150 -300
rect 82 -306 83 -302
rect 86 -306 87 -302
rect 96 -303 97 -291
rect 156 -306 157 -302
rect 89 -306 90 -304
rect 96 -306 97 -304
rect 103 -306 104 -304
rect 135 -305 136 -291
rect 44 -335 45 -315
rect 89 -316 90 -314
rect 96 -335 97 -315
rect 135 -316 136 -314
rect 159 -335 160 -315
rect 170 -316 171 -314
rect 177 -316 178 -314
rect 205 -335 206 -315
rect 219 -316 220 -314
rect 219 -335 220 -315
rect 219 -316 220 -314
rect 219 -335 220 -315
rect 226 -316 227 -314
rect 233 -316 234 -314
rect 236 -316 237 -314
rect 240 -316 241 -314
rect 51 -318 52 -314
rect 89 -335 90 -317
rect 107 -318 108 -314
rect 128 -318 129 -314
rect 138 -318 139 -314
rect 170 -335 171 -317
rect 51 -335 52 -319
rect 93 -320 94 -314
rect 107 -335 108 -319
rect 121 -320 122 -314
rect 128 -335 129 -319
rect 156 -320 157 -314
rect 61 -322 62 -314
rect 65 -322 66 -314
rect 72 -322 73 -314
rect 117 -322 118 -314
rect 138 -335 139 -321
rect 191 -335 192 -321
rect 61 -335 62 -323
rect 75 -324 76 -314
rect 79 -335 80 -323
rect 198 -335 199 -323
rect 65 -335 66 -325
rect 86 -335 87 -325
rect 93 -335 94 -325
rect 100 -326 101 -314
rect 114 -326 115 -314
rect 163 -326 164 -314
rect 37 -335 38 -327
rect 100 -335 101 -327
rect 117 -335 118 -327
rect 121 -335 122 -327
rect 135 -335 136 -327
rect 163 -335 164 -327
rect 72 -335 73 -329
rect 142 -330 143 -314
rect 149 -330 150 -314
rect 177 -335 178 -329
rect 131 -335 132 -331
rect 149 -335 150 -331
rect 142 -335 143 -333
rect 184 -335 185 -333
rect 37 -345 38 -343
rect 79 -345 80 -343
rect 100 -345 101 -343
rect 163 -345 164 -343
rect 194 -362 195 -344
rect 198 -345 199 -343
rect 215 -345 216 -343
rect 219 -345 220 -343
rect 44 -347 45 -343
rect 117 -347 118 -343
rect 121 -347 122 -343
rect 121 -362 122 -346
rect 121 -347 122 -343
rect 121 -362 122 -346
rect 135 -362 136 -346
rect 142 -347 143 -343
rect 145 -347 146 -343
rect 205 -347 206 -343
rect 58 -349 59 -343
rect 93 -349 94 -343
rect 110 -362 111 -348
rect 212 -349 213 -343
rect 51 -351 52 -343
rect 58 -362 59 -350
rect 65 -351 66 -343
rect 65 -362 66 -350
rect 65 -351 66 -343
rect 65 -362 66 -350
rect 72 -351 73 -343
rect 138 -351 139 -343
rect 149 -351 150 -343
rect 163 -362 164 -350
rect 177 -351 178 -343
rect 198 -362 199 -350
rect 72 -362 73 -352
rect 96 -353 97 -343
rect 114 -353 115 -343
rect 170 -353 171 -343
rect 177 -362 178 -352
rect 191 -353 192 -343
rect 79 -362 80 -354
rect 107 -355 108 -343
rect 149 -362 150 -354
rect 156 -355 157 -343
rect 170 -362 171 -354
rect 184 -355 185 -343
rect 86 -362 87 -356
rect 142 -362 143 -356
rect 96 -362 97 -358
rect 103 -359 104 -343
rect 131 -359 132 -343
rect 184 -362 185 -358
rect 103 -362 104 -360
rect 128 -362 129 -360
rect 58 -372 59 -370
rect 124 -385 125 -371
rect 135 -372 136 -370
rect 142 -372 143 -370
rect 145 -372 146 -370
rect 184 -372 185 -370
rect 65 -374 66 -370
rect 107 -374 108 -370
rect 138 -385 139 -373
rect 149 -374 150 -370
rect 156 -374 157 -370
rect 198 -374 199 -370
rect 72 -376 73 -370
rect 100 -376 101 -370
rect 103 -385 104 -375
rect 128 -376 129 -370
rect 142 -385 143 -375
rect 163 -376 164 -370
rect 170 -385 171 -375
rect 177 -376 178 -370
rect 72 -385 73 -377
rect 96 -385 97 -377
rect 100 -385 101 -377
rect 107 -385 108 -377
rect 114 -378 115 -370
rect 156 -385 157 -377
rect 79 -380 80 -370
rect 117 -380 118 -370
rect 121 -380 122 -370
rect 128 -385 129 -379
rect 149 -385 150 -379
rect 173 -385 174 -379
rect 79 -385 80 -381
rect 93 -385 94 -381
rect 121 -385 122 -381
rect 163 -385 164 -381
rect 86 -384 87 -370
rect 86 -385 87 -383
rect 86 -384 87 -370
rect 86 -385 87 -383
rect 79 -395 80 -393
rect 100 -395 101 -393
rect 114 -395 115 -393
rect 128 -395 129 -393
rect 131 -406 132 -394
rect 149 -395 150 -393
rect 170 -395 171 -393
rect 173 -406 174 -394
rect 72 -397 73 -393
rect 128 -406 129 -396
rect 145 -406 146 -396
rect 156 -397 157 -393
rect 86 -399 87 -393
rect 138 -399 139 -393
rect 79 -406 80 -400
rect 86 -406 87 -400
rect 93 -406 94 -400
rect 107 -401 108 -393
rect 121 -401 122 -393
rect 142 -401 143 -393
rect 117 -403 118 -393
rect 121 -406 122 -402
rect 142 -406 143 -402
rect 163 -403 164 -393
rect 107 -406 108 -404
rect 117 -406 118 -404
rect 156 -406 157 -404
rect 163 -406 164 -404
rect 93 -416 94 -414
rect 100 -416 101 -414
rect 117 -416 118 -414
rect 121 -416 122 -414
rect 156 -416 157 -414
rect 163 -419 164 -415
rect 86 -418 87 -414
rect 93 -419 94 -417
rect 107 -418 108 -414
rect 121 -419 122 -417
rect 89 -429 90 -427
rect 93 -429 94 -427
rect 117 -429 118 -427
rect 121 -429 122 -427
rect 163 -429 164 -427
rect 170 -429 171 -427
<< labels >>
rlabel pdiffusion 3 -8 3 -8 0 cellNo=35
rlabel pdiffusion 10 -8 10 -8 0 cellNo=64
rlabel pdiffusion 17 -8 17 -8 0 cellNo=147
rlabel pdiffusion 73 -8 73 -8 0 cellNo=61
rlabel pdiffusion 94 -8 94 -8 0 feedthrough
rlabel pdiffusion 101 -8 101 -8 0 cellNo=105
rlabel pdiffusion 108 -8 108 -8 0 cellNo=155
rlabel pdiffusion 115 -8 115 -8 0 feedthrough
rlabel pdiffusion 178 -8 178 -8 0 cellNo=59
rlabel pdiffusion 185 -8 185 -8 0 feedthrough
rlabel pdiffusion 192 -8 192 -8 0 cellNo=177
rlabel pdiffusion 199 -8 199 -8 0 feedthrough
rlabel pdiffusion 3 -21 3 -21 0 cellNo=62
rlabel pdiffusion 10 -21 10 -21 0 cellNo=106
rlabel pdiffusion 17 -21 17 -21 0 cellNo=109
rlabel pdiffusion 59 -21 59 -21 0 feedthrough
rlabel pdiffusion 66 -21 66 -21 0 cellNo=88
rlabel pdiffusion 73 -21 73 -21 0 cellNo=128
rlabel pdiffusion 80 -21 80 -21 0 feedthrough
rlabel pdiffusion 87 -21 87 -21 0 cellNo=63
rlabel pdiffusion 94 -21 94 -21 0 feedthrough
rlabel pdiffusion 101 -21 101 -21 0 cellNo=46
rlabel pdiffusion 108 -21 108 -21 0 cellNo=10
rlabel pdiffusion 115 -21 115 -21 0 cellNo=164
rlabel pdiffusion 129 -21 129 -21 0 feedthrough
rlabel pdiffusion 178 -21 178 -21 0 feedthrough
rlabel pdiffusion 185 -21 185 -21 0 cellNo=110
rlabel pdiffusion 199 -21 199 -21 0 cellNo=29
rlabel pdiffusion 206 -21 206 -21 0 feedthrough
rlabel pdiffusion 3 -40 3 -40 0 cellNo=67
rlabel pdiffusion 10 -40 10 -40 0 cellNo=157
rlabel pdiffusion 45 -40 45 -40 0 cellNo=32
rlabel pdiffusion 52 -40 52 -40 0 feedthrough
rlabel pdiffusion 59 -40 59 -40 0 feedthrough
rlabel pdiffusion 66 -40 66 -40 0 cellNo=122
rlabel pdiffusion 73 -40 73 -40 0 cellNo=24
rlabel pdiffusion 80 -40 80 -40 0 cellNo=85
rlabel pdiffusion 87 -40 87 -40 0 cellNo=4
rlabel pdiffusion 94 -40 94 -40 0 cellNo=76
rlabel pdiffusion 101 -40 101 -40 0 cellNo=48
rlabel pdiffusion 108 -40 108 -40 0 cellNo=38
rlabel pdiffusion 115 -40 115 -40 0 cellNo=143
rlabel pdiffusion 122 -40 122 -40 0 feedthrough
rlabel pdiffusion 129 -40 129 -40 0 feedthrough
rlabel pdiffusion 136 -40 136 -40 0 cellNo=99
rlabel pdiffusion 143 -40 143 -40 0 feedthrough
rlabel pdiffusion 150 -40 150 -40 0 cellNo=170
rlabel pdiffusion 157 -40 157 -40 0 feedthrough
rlabel pdiffusion 171 -40 171 -40 0 feedthrough
rlabel pdiffusion 178 -40 178 -40 0 cellNo=131
rlabel pdiffusion 185 -40 185 -40 0 feedthrough
rlabel pdiffusion 3 -61 3 -61 0 cellNo=108
rlabel pdiffusion 31 -61 31 -61 0 feedthrough
rlabel pdiffusion 38 -61 38 -61 0 feedthrough
rlabel pdiffusion 45 -61 45 -61 0 cellNo=28
rlabel pdiffusion 52 -61 52 -61 0 feedthrough
rlabel pdiffusion 59 -61 59 -61 0 feedthrough
rlabel pdiffusion 66 -61 66 -61 0 cellNo=23
rlabel pdiffusion 73 -61 73 -61 0 cellNo=93
rlabel pdiffusion 80 -61 80 -61 0 cellNo=44
rlabel pdiffusion 87 -61 87 -61 0 feedthrough
rlabel pdiffusion 94 -61 94 -61 0 feedthrough
rlabel pdiffusion 101 -61 101 -61 0 cellNo=19
rlabel pdiffusion 108 -61 108 -61 0 cellNo=94
rlabel pdiffusion 115 -61 115 -61 0 feedthrough
rlabel pdiffusion 122 -61 122 -61 0 feedthrough
rlabel pdiffusion 129 -61 129 -61 0 cellNo=104
rlabel pdiffusion 136 -61 136 -61 0 cellNo=34
rlabel pdiffusion 143 -61 143 -61 0 feedthrough
rlabel pdiffusion 150 -61 150 -61 0 feedthrough
rlabel pdiffusion 157 -61 157 -61 0 cellNo=15
rlabel pdiffusion 164 -61 164 -61 0 feedthrough
rlabel pdiffusion 171 -61 171 -61 0 feedthrough
rlabel pdiffusion 178 -61 178 -61 0 feedthrough
rlabel pdiffusion 185 -61 185 -61 0 cellNo=45
rlabel pdiffusion 192 -61 192 -61 0 feedthrough
rlabel pdiffusion 52 -90 52 -90 0 cellNo=102
rlabel pdiffusion 66 -90 66 -90 0 cellNo=141
rlabel pdiffusion 73 -90 73 -90 0 feedthrough
rlabel pdiffusion 80 -90 80 -90 0 feedthrough
rlabel pdiffusion 87 -90 87 -90 0 cellNo=101
rlabel pdiffusion 94 -90 94 -90 0 feedthrough
rlabel pdiffusion 101 -90 101 -90 0 cellNo=148
rlabel pdiffusion 108 -90 108 -90 0 cellNo=43
rlabel pdiffusion 115 -90 115 -90 0 feedthrough
rlabel pdiffusion 122 -90 122 -90 0 feedthrough
rlabel pdiffusion 129 -90 129 -90 0 cellNo=97
rlabel pdiffusion 136 -90 136 -90 0 feedthrough
rlabel pdiffusion 143 -90 143 -90 0 cellNo=60
rlabel pdiffusion 150 -90 150 -90 0 cellNo=144
rlabel pdiffusion 157 -90 157 -90 0 feedthrough
rlabel pdiffusion 164 -90 164 -90 0 feedthrough
rlabel pdiffusion 171 -90 171 -90 0 feedthrough
rlabel pdiffusion 178 -90 178 -90 0 feedthrough
rlabel pdiffusion 185 -90 185 -90 0 feedthrough
rlabel pdiffusion 192 -90 192 -90 0 cellNo=50
rlabel pdiffusion 199 -90 199 -90 0 feedthrough
rlabel pdiffusion 206 -90 206 -90 0 feedthrough
rlabel pdiffusion 213 -90 213 -90 0 feedthrough
rlabel pdiffusion 220 -90 220 -90 0 feedthrough
rlabel pdiffusion 227 -90 227 -90 0 feedthrough
rlabel pdiffusion 234 -90 234 -90 0 feedthrough
rlabel pdiffusion 241 -90 241 -90 0 cellNo=2
rlabel pdiffusion 248 -90 248 -90 0 cellNo=54
rlabel pdiffusion 3 -119 3 -119 0 feedthrough
rlabel pdiffusion 10 -119 10 -119 0 feedthrough
rlabel pdiffusion 17 -119 17 -119 0 cellNo=21
rlabel pdiffusion 24 -119 24 -119 0 feedthrough
rlabel pdiffusion 31 -119 31 -119 0 feedthrough
rlabel pdiffusion 38 -119 38 -119 0 cellNo=71
rlabel pdiffusion 45 -119 45 -119 0 cellNo=1
rlabel pdiffusion 52 -119 52 -119 0 feedthrough
rlabel pdiffusion 59 -119 59 -119 0 feedthrough
rlabel pdiffusion 66 -119 66 -119 0 cellNo=75
rlabel pdiffusion 73 -119 73 -119 0 cellNo=22
rlabel pdiffusion 80 -119 80 -119 0 cellNo=162
rlabel pdiffusion 87 -119 87 -119 0 cellNo=47
rlabel pdiffusion 94 -119 94 -119 0 feedthrough
rlabel pdiffusion 101 -119 101 -119 0 cellNo=57
rlabel pdiffusion 108 -119 108 -119 0 feedthrough
rlabel pdiffusion 115 -119 115 -119 0 cellNo=118
rlabel pdiffusion 122 -119 122 -119 0 cellNo=136
rlabel pdiffusion 129 -119 129 -119 0 feedthrough
rlabel pdiffusion 136 -119 136 -119 0 feedthrough
rlabel pdiffusion 143 -119 143 -119 0 cellNo=56
rlabel pdiffusion 150 -119 150 -119 0 cellNo=53
rlabel pdiffusion 157 -119 157 -119 0 cellNo=42
rlabel pdiffusion 164 -119 164 -119 0 feedthrough
rlabel pdiffusion 171 -119 171 -119 0 feedthrough
rlabel pdiffusion 178 -119 178 -119 0 feedthrough
rlabel pdiffusion 185 -119 185 -119 0 feedthrough
rlabel pdiffusion 192 -119 192 -119 0 feedthrough
rlabel pdiffusion 199 -119 199 -119 0 feedthrough
rlabel pdiffusion 206 -119 206 -119 0 feedthrough
rlabel pdiffusion 213 -119 213 -119 0 feedthrough
rlabel pdiffusion 220 -119 220 -119 0 feedthrough
rlabel pdiffusion 227 -119 227 -119 0 feedthrough
rlabel pdiffusion 234 -119 234 -119 0 feedthrough
rlabel pdiffusion 241 -119 241 -119 0 feedthrough
rlabel pdiffusion 248 -119 248 -119 0 feedthrough
rlabel pdiffusion 255 -119 255 -119 0 cellNo=74
rlabel pdiffusion 3 -164 3 -164 0 feedthrough
rlabel pdiffusion 10 -164 10 -164 0 feedthrough
rlabel pdiffusion 17 -164 17 -164 0 cellNo=156
rlabel pdiffusion 24 -164 24 -164 0 cellNo=127
rlabel pdiffusion 31 -164 31 -164 0 cellNo=89
rlabel pdiffusion 38 -164 38 -164 0 cellNo=8
rlabel pdiffusion 45 -164 45 -164 0 cellNo=95
rlabel pdiffusion 52 -164 52 -164 0 feedthrough
rlabel pdiffusion 59 -164 59 -164 0 cellNo=112
rlabel pdiffusion 66 -164 66 -164 0 feedthrough
rlabel pdiffusion 73 -164 73 -164 0 feedthrough
rlabel pdiffusion 80 -164 80 -164 0 cellNo=163
rlabel pdiffusion 87 -164 87 -164 0 cellNo=152
rlabel pdiffusion 94 -164 94 -164 0 cellNo=31
rlabel pdiffusion 101 -164 101 -164 0 feedthrough
rlabel pdiffusion 108 -164 108 -164 0 cellNo=33
rlabel pdiffusion 115 -164 115 -164 0 cellNo=70
rlabel pdiffusion 122 -164 122 -164 0 feedthrough
rlabel pdiffusion 129 -164 129 -164 0 feedthrough
rlabel pdiffusion 136 -164 136 -164 0 cellNo=9
rlabel pdiffusion 143 -164 143 -164 0 feedthrough
rlabel pdiffusion 150 -164 150 -164 0 feedthrough
rlabel pdiffusion 157 -164 157 -164 0 cellNo=39
rlabel pdiffusion 164 -164 164 -164 0 feedthrough
rlabel pdiffusion 171 -164 171 -164 0 feedthrough
rlabel pdiffusion 178 -164 178 -164 0 feedthrough
rlabel pdiffusion 185 -164 185 -164 0 cellNo=3
rlabel pdiffusion 192 -164 192 -164 0 feedthrough
rlabel pdiffusion 199 -164 199 -164 0 feedthrough
rlabel pdiffusion 206 -164 206 -164 0 feedthrough
rlabel pdiffusion 213 -164 213 -164 0 feedthrough
rlabel pdiffusion 220 -164 220 -164 0 feedthrough
rlabel pdiffusion 227 -164 227 -164 0 feedthrough
rlabel pdiffusion 234 -164 234 -164 0 feedthrough
rlabel pdiffusion 241 -164 241 -164 0 feedthrough
rlabel pdiffusion 248 -164 248 -164 0 feedthrough
rlabel pdiffusion 255 -164 255 -164 0 feedthrough
rlabel pdiffusion 262 -164 262 -164 0 feedthrough
rlabel pdiffusion 269 -164 269 -164 0 feedthrough
rlabel pdiffusion 276 -164 276 -164 0 cellNo=180
rlabel pdiffusion 24 -195 24 -195 0 feedthrough
rlabel pdiffusion 31 -195 31 -195 0 feedthrough
rlabel pdiffusion 38 -195 38 -195 0 cellNo=121
rlabel pdiffusion 45 -195 45 -195 0 cellNo=30
rlabel pdiffusion 52 -195 52 -195 0 feedthrough
rlabel pdiffusion 59 -195 59 -195 0 feedthrough
rlabel pdiffusion 66 -195 66 -195 0 cellNo=150
rlabel pdiffusion 73 -195 73 -195 0 feedthrough
rlabel pdiffusion 80 -195 80 -195 0 cellNo=72
rlabel pdiffusion 87 -195 87 -195 0 feedthrough
rlabel pdiffusion 94 -195 94 -195 0 cellNo=86
rlabel pdiffusion 101 -195 101 -195 0 cellNo=149
rlabel pdiffusion 108 -195 108 -195 0 cellNo=5
rlabel pdiffusion 115 -195 115 -195 0 cellNo=27
rlabel pdiffusion 122 -195 122 -195 0 feedthrough
rlabel pdiffusion 129 -195 129 -195 0 cellNo=98
rlabel pdiffusion 136 -195 136 -195 0 cellNo=37
rlabel pdiffusion 143 -195 143 -195 0 cellNo=81
rlabel pdiffusion 150 -195 150 -195 0 cellNo=153
rlabel pdiffusion 157 -195 157 -195 0 feedthrough
rlabel pdiffusion 164 -195 164 -195 0 feedthrough
rlabel pdiffusion 171 -195 171 -195 0 feedthrough
rlabel pdiffusion 178 -195 178 -195 0 feedthrough
rlabel pdiffusion 185 -195 185 -195 0 cellNo=176
rlabel pdiffusion 192 -195 192 -195 0 cellNo=160
rlabel pdiffusion 199 -195 199 -195 0 feedthrough
rlabel pdiffusion 206 -195 206 -195 0 feedthrough
rlabel pdiffusion 213 -195 213 -195 0 feedthrough
rlabel pdiffusion 220 -195 220 -195 0 feedthrough
rlabel pdiffusion 227 -195 227 -195 0 feedthrough
rlabel pdiffusion 234 -195 234 -195 0 feedthrough
rlabel pdiffusion 241 -195 241 -195 0 feedthrough
rlabel pdiffusion 248 -195 248 -195 0 feedthrough
rlabel pdiffusion 255 -195 255 -195 0 feedthrough
rlabel pdiffusion 262 -195 262 -195 0 feedthrough
rlabel pdiffusion 283 -195 283 -195 0 cellNo=91
rlabel pdiffusion 31 -230 31 -230 0 cellNo=175
rlabel pdiffusion 38 -230 38 -230 0 feedthrough
rlabel pdiffusion 45 -230 45 -230 0 cellNo=167
rlabel pdiffusion 52 -230 52 -230 0 feedthrough
rlabel pdiffusion 59 -230 59 -230 0 feedthrough
rlabel pdiffusion 66 -230 66 -230 0 feedthrough
rlabel pdiffusion 73 -230 73 -230 0 cellNo=79
rlabel pdiffusion 80 -230 80 -230 0 cellNo=139
rlabel pdiffusion 87 -230 87 -230 0 feedthrough
rlabel pdiffusion 94 -230 94 -230 0 cellNo=138
rlabel pdiffusion 101 -230 101 -230 0 feedthrough
rlabel pdiffusion 108 -230 108 -230 0 feedthrough
rlabel pdiffusion 115 -230 115 -230 0 cellNo=87
rlabel pdiffusion 122 -230 122 -230 0 feedthrough
rlabel pdiffusion 129 -230 129 -230 0 feedthrough
rlabel pdiffusion 136 -230 136 -230 0 cellNo=14
rlabel pdiffusion 143 -230 143 -230 0 feedthrough
rlabel pdiffusion 150 -230 150 -230 0 cellNo=142
rlabel pdiffusion 157 -230 157 -230 0 cellNo=165
rlabel pdiffusion 164 -230 164 -230 0 feedthrough
rlabel pdiffusion 171 -230 171 -230 0 feedthrough
rlabel pdiffusion 178 -230 178 -230 0 cellNo=55
rlabel pdiffusion 185 -230 185 -230 0 feedthrough
rlabel pdiffusion 192 -230 192 -230 0 cellNo=17
rlabel pdiffusion 199 -230 199 -230 0 feedthrough
rlabel pdiffusion 206 -230 206 -230 0 feedthrough
rlabel pdiffusion 213 -230 213 -230 0 feedthrough
rlabel pdiffusion 220 -230 220 -230 0 feedthrough
rlabel pdiffusion 227 -230 227 -230 0 feedthrough
rlabel pdiffusion 234 -230 234 -230 0 feedthrough
rlabel pdiffusion 241 -230 241 -230 0 feedthrough
rlabel pdiffusion 248 -230 248 -230 0 feedthrough
rlabel pdiffusion 255 -230 255 -230 0 feedthrough
rlabel pdiffusion 262 -230 262 -230 0 cellNo=146
rlabel pdiffusion 269 -230 269 -230 0 cellNo=100
rlabel pdiffusion 276 -230 276 -230 0 cellNo=12
rlabel pdiffusion 283 -230 283 -230 0 feedthrough
rlabel pdiffusion 290 -230 290 -230 0 feedthrough
rlabel pdiffusion 17 -261 17 -261 0 feedthrough
rlabel pdiffusion 24 -261 24 -261 0 cellNo=18
rlabel pdiffusion 31 -261 31 -261 0 feedthrough
rlabel pdiffusion 38 -261 38 -261 0 feedthrough
rlabel pdiffusion 45 -261 45 -261 0 cellNo=171
rlabel pdiffusion 52 -261 52 -261 0 cellNo=83
rlabel pdiffusion 59 -261 59 -261 0 feedthrough
rlabel pdiffusion 66 -261 66 -261 0 feedthrough
rlabel pdiffusion 73 -261 73 -261 0 feedthrough
rlabel pdiffusion 80 -261 80 -261 0 feedthrough
rlabel pdiffusion 87 -261 87 -261 0 feedthrough
rlabel pdiffusion 94 -261 94 -261 0 feedthrough
rlabel pdiffusion 101 -261 101 -261 0 cellNo=179
rlabel pdiffusion 108 -261 108 -261 0 cellNo=130
rlabel pdiffusion 115 -261 115 -261 0 cellNo=166
rlabel pdiffusion 122 -261 122 -261 0 feedthrough
rlabel pdiffusion 129 -261 129 -261 0 feedthrough
rlabel pdiffusion 136 -261 136 -261 0 cellNo=40
rlabel pdiffusion 143 -261 143 -261 0 feedthrough
rlabel pdiffusion 150 -261 150 -261 0 feedthrough
rlabel pdiffusion 157 -261 157 -261 0 feedthrough
rlabel pdiffusion 164 -261 164 -261 0 feedthrough
rlabel pdiffusion 171 -261 171 -261 0 cellNo=36
rlabel pdiffusion 178 -261 178 -261 0 cellNo=137
rlabel pdiffusion 185 -261 185 -261 0 feedthrough
rlabel pdiffusion 192 -261 192 -261 0 cellNo=78
rlabel pdiffusion 199 -261 199 -261 0 feedthrough
rlabel pdiffusion 206 -261 206 -261 0 feedthrough
rlabel pdiffusion 213 -261 213 -261 0 feedthrough
rlabel pdiffusion 220 -261 220 -261 0 feedthrough
rlabel pdiffusion 227 -261 227 -261 0 feedthrough
rlabel pdiffusion 234 -261 234 -261 0 feedthrough
rlabel pdiffusion 241 -261 241 -261 0 feedthrough
rlabel pdiffusion 248 -261 248 -261 0 feedthrough
rlabel pdiffusion 255 -261 255 -261 0 feedthrough
rlabel pdiffusion 283 -261 283 -261 0 feedthrough
rlabel pdiffusion 290 -261 290 -261 0 cellNo=120
rlabel pdiffusion 66 -288 66 -288 0 feedthrough
rlabel pdiffusion 73 -288 73 -288 0 feedthrough
rlabel pdiffusion 80 -288 80 -288 0 cellNo=25
rlabel pdiffusion 87 -288 87 -288 0 cellNo=84
rlabel pdiffusion 94 -288 94 -288 0 cellNo=119
rlabel pdiffusion 101 -288 101 -288 0 cellNo=69
rlabel pdiffusion 108 -288 108 -288 0 feedthrough
rlabel pdiffusion 115 -288 115 -288 0 cellNo=151
rlabel pdiffusion 122 -288 122 -288 0 feedthrough
rlabel pdiffusion 129 -288 129 -288 0 feedthrough
rlabel pdiffusion 136 -288 136 -288 0 feedthrough
rlabel pdiffusion 143 -288 143 -288 0 feedthrough
rlabel pdiffusion 150 -288 150 -288 0 feedthrough
rlabel pdiffusion 157 -288 157 -288 0 feedthrough
rlabel pdiffusion 164 -288 164 -288 0 cellNo=111
rlabel pdiffusion 171 -288 171 -288 0 feedthrough
rlabel pdiffusion 185 -288 185 -288 0 cellNo=161
rlabel pdiffusion 192 -288 192 -288 0 cellNo=159
rlabel pdiffusion 199 -288 199 -288 0 feedthrough
rlabel pdiffusion 206 -288 206 -288 0 cellNo=20
rlabel pdiffusion 241 -288 241 -288 0 feedthrough
rlabel pdiffusion 248 -288 248 -288 0 cellNo=107
rlabel pdiffusion 255 -288 255 -288 0 feedthrough
rlabel pdiffusion 52 -311 52 -311 0 feedthrough
rlabel pdiffusion 59 -311 59 -311 0 cellNo=41
rlabel pdiffusion 66 -311 66 -311 0 feedthrough
rlabel pdiffusion 73 -311 73 -311 0 cellNo=116
rlabel pdiffusion 80 -311 80 -311 0 cellNo=115
rlabel pdiffusion 87 -311 87 -311 0 cellNo=169
rlabel pdiffusion 94 -311 94 -311 0 cellNo=11
rlabel pdiffusion 101 -311 101 -311 0 cellNo=80
rlabel pdiffusion 108 -311 108 -311 0 cellNo=134
rlabel pdiffusion 115 -311 115 -311 0 cellNo=133
rlabel pdiffusion 122 -311 122 -311 0 feedthrough
rlabel pdiffusion 129 -311 129 -311 0 feedthrough
rlabel pdiffusion 136 -311 136 -311 0 cellNo=77
rlabel pdiffusion 143 -311 143 -311 0 feedthrough
rlabel pdiffusion 150 -311 150 -311 0 feedthrough
rlabel pdiffusion 157 -311 157 -311 0 feedthrough
rlabel pdiffusion 164 -311 164 -311 0 feedthrough
rlabel pdiffusion 171 -311 171 -311 0 feedthrough
rlabel pdiffusion 178 -311 178 -311 0 feedthrough
rlabel pdiffusion 220 -311 220 -311 0 feedthrough
rlabel pdiffusion 227 -311 227 -311 0 cellNo=6
rlabel pdiffusion 234 -311 234 -311 0 cellNo=51
rlabel pdiffusion 241 -311 241 -311 0 feedthrough
rlabel pdiffusion 38 -340 38 -340 0 feedthrough
rlabel pdiffusion 45 -340 45 -340 0 feedthrough
rlabel pdiffusion 52 -340 52 -340 0 feedthrough
rlabel pdiffusion 59 -340 59 -340 0 cellNo=123
rlabel pdiffusion 66 -340 66 -340 0 feedthrough
rlabel pdiffusion 73 -340 73 -340 0 feedthrough
rlabel pdiffusion 80 -340 80 -340 0 cellNo=49
rlabel pdiffusion 87 -340 87 -340 0 cellNo=168
rlabel pdiffusion 94 -340 94 -340 0 cellNo=124
rlabel pdiffusion 101 -340 101 -340 0 cellNo=92
rlabel pdiffusion 108 -340 108 -340 0 feedthrough
rlabel pdiffusion 115 -340 115 -340 0 cellNo=16
rlabel pdiffusion 122 -340 122 -340 0 feedthrough
rlabel pdiffusion 129 -340 129 -340 0 cellNo=126
rlabel pdiffusion 136 -340 136 -340 0 cellNo=68
rlabel pdiffusion 143 -340 143 -340 0 cellNo=7
rlabel pdiffusion 150 -340 150 -340 0 feedthrough
rlabel pdiffusion 157 -340 157 -340 0 cellNo=129
rlabel pdiffusion 164 -340 164 -340 0 feedthrough
rlabel pdiffusion 171 -340 171 -340 0 feedthrough
rlabel pdiffusion 178 -340 178 -340 0 feedthrough
rlabel pdiffusion 185 -340 185 -340 0 feedthrough
rlabel pdiffusion 192 -340 192 -340 0 feedthrough
rlabel pdiffusion 199 -340 199 -340 0 feedthrough
rlabel pdiffusion 206 -340 206 -340 0 feedthrough
rlabel pdiffusion 213 -340 213 -340 0 cellNo=145
rlabel pdiffusion 220 -340 220 -340 0 feedthrough
rlabel pdiffusion 59 -367 59 -367 0 feedthrough
rlabel pdiffusion 66 -367 66 -367 0 feedthrough
rlabel pdiffusion 73 -367 73 -367 0 feedthrough
rlabel pdiffusion 80 -367 80 -367 0 feedthrough
rlabel pdiffusion 87 -367 87 -367 0 feedthrough
rlabel pdiffusion 94 -367 94 -367 0 cellNo=52
rlabel pdiffusion 101 -367 101 -367 0 cellNo=82
rlabel pdiffusion 108 -367 108 -367 0 cellNo=172
rlabel pdiffusion 115 -367 115 -367 0 cellNo=173
rlabel pdiffusion 122 -367 122 -367 0 feedthrough
rlabel pdiffusion 129 -367 129 -367 0 feedthrough
rlabel pdiffusion 136 -367 136 -367 0 feedthrough
rlabel pdiffusion 143 -367 143 -367 0 cellNo=132
rlabel pdiffusion 150 -367 150 -367 0 feedthrough
rlabel pdiffusion 157 -367 157 -367 0 cellNo=13
rlabel pdiffusion 164 -367 164 -367 0 feedthrough
rlabel pdiffusion 171 -367 171 -367 0 cellNo=174
rlabel pdiffusion 178 -367 178 -367 0 feedthrough
rlabel pdiffusion 185 -367 185 -367 0 feedthrough
rlabel pdiffusion 192 -367 192 -367 0 cellNo=66
rlabel pdiffusion 199 -367 199 -367 0 feedthrough
rlabel pdiffusion 73 -390 73 -390 0 feedthrough
rlabel pdiffusion 80 -390 80 -390 0 feedthrough
rlabel pdiffusion 87 -390 87 -390 0 feedthrough
rlabel pdiffusion 94 -390 94 -390 0 cellNo=26
rlabel pdiffusion 101 -390 101 -390 0 cellNo=65
rlabel pdiffusion 108 -390 108 -390 0 feedthrough
rlabel pdiffusion 115 -390 115 -390 0 cellNo=113
rlabel pdiffusion 122 -390 122 -390 0 cellNo=158
rlabel pdiffusion 129 -390 129 -390 0 feedthrough
rlabel pdiffusion 136 -390 136 -390 0 cellNo=90
rlabel pdiffusion 143 -390 143 -390 0 feedthrough
rlabel pdiffusion 150 -390 150 -390 0 feedthrough
rlabel pdiffusion 157 -390 157 -390 0 feedthrough
rlabel pdiffusion 164 -390 164 -390 0 feedthrough
rlabel pdiffusion 171 -390 171 -390 0 cellNo=135
rlabel pdiffusion 80 -411 80 -411 0 cellNo=125
rlabel pdiffusion 87 -411 87 -411 0 feedthrough
rlabel pdiffusion 94 -411 94 -411 0 feedthrough
rlabel pdiffusion 101 -411 101 -411 0 cellNo=154
rlabel pdiffusion 108 -411 108 -411 0 feedthrough
rlabel pdiffusion 115 -411 115 -411 0 cellNo=140
rlabel pdiffusion 122 -411 122 -411 0 feedthrough
rlabel pdiffusion 129 -411 129 -411 0 cellNo=73
rlabel pdiffusion 143 -411 143 -411 0 cellNo=103
rlabel pdiffusion 157 -411 157 -411 0 feedthrough
rlabel pdiffusion 164 -411 164 -411 0 cellNo=114
rlabel pdiffusion 171 -411 171 -411 0 cellNo=178
rlabel pdiffusion 87 -424 87 -424 0 cellNo=58
rlabel pdiffusion 94 -424 94 -424 0 feedthrough
rlabel pdiffusion 115 -424 115 -424 0 cellNo=117
rlabel pdiffusion 122 -424 122 -424 0 feedthrough
rlabel pdiffusion 164 -424 164 -424 0 feedthrough
rlabel pdiffusion 171 -424 171 -424 0 cellNo=96
rlabel polysilicon 75 -10 75 -10 0 4
rlabel polysilicon 93 -4 93 -4 0 1
rlabel polysilicon 93 -10 93 -10 0 3
rlabel polysilicon 100 -4 100 -4 0 1
rlabel polysilicon 103 -4 103 -4 0 2
rlabel polysilicon 107 -10 107 -10 0 3
rlabel polysilicon 114 -4 114 -4 0 1
rlabel polysilicon 114 -10 114 -10 0 3
rlabel polysilicon 177 -4 177 -4 0 1
rlabel polysilicon 184 -4 184 -4 0 1
rlabel polysilicon 184 -10 184 -10 0 3
rlabel polysilicon 191 -4 191 -4 0 1
rlabel polysilicon 191 -10 191 -10 0 3
rlabel polysilicon 198 -4 198 -4 0 1
rlabel polysilicon 198 -10 198 -10 0 3
rlabel polysilicon 58 -17 58 -17 0 1
rlabel polysilicon 58 -23 58 -23 0 3
rlabel polysilicon 68 -17 68 -17 0 2
rlabel polysilicon 65 -23 65 -23 0 3
rlabel polysilicon 75 -17 75 -17 0 2
rlabel polysilicon 79 -17 79 -17 0 1
rlabel polysilicon 79 -23 79 -23 0 3
rlabel polysilicon 89 -17 89 -17 0 2
rlabel polysilicon 93 -17 93 -17 0 1
rlabel polysilicon 93 -23 93 -23 0 3
rlabel polysilicon 100 -17 100 -17 0 1
rlabel polysilicon 107 -17 107 -17 0 1
rlabel polysilicon 117 -17 117 -17 0 2
rlabel polysilicon 128 -17 128 -17 0 1
rlabel polysilicon 128 -23 128 -23 0 3
rlabel polysilicon 177 -17 177 -17 0 1
rlabel polysilicon 177 -23 177 -23 0 3
rlabel polysilicon 184 -17 184 -17 0 1
rlabel polysilicon 198 -23 198 -23 0 3
rlabel polysilicon 205 -17 205 -17 0 1
rlabel polysilicon 205 -23 205 -23 0 3
rlabel polysilicon 44 -42 44 -42 0 3
rlabel polysilicon 51 -36 51 -36 0 1
rlabel polysilicon 51 -42 51 -42 0 3
rlabel polysilicon 58 -36 58 -36 0 1
rlabel polysilicon 58 -42 58 -42 0 3
rlabel polysilicon 65 -36 65 -36 0 1
rlabel polysilicon 65 -42 65 -42 0 3
rlabel polysilicon 72 -42 72 -42 0 3
rlabel polysilicon 79 -36 79 -36 0 1
rlabel polysilicon 79 -42 79 -42 0 3
rlabel polysilicon 86 -36 86 -36 0 1
rlabel polysilicon 86 -42 86 -42 0 3
rlabel polysilicon 93 -36 93 -36 0 1
rlabel polysilicon 96 -36 96 -36 0 2
rlabel polysilicon 100 -36 100 -36 0 1
rlabel polysilicon 103 -42 103 -42 0 4
rlabel polysilicon 107 -36 107 -36 0 1
rlabel polysilicon 107 -42 107 -42 0 3
rlabel polysilicon 110 -42 110 -42 0 4
rlabel polysilicon 117 -36 117 -36 0 2
rlabel polysilicon 114 -42 114 -42 0 3
rlabel polysilicon 117 -42 117 -42 0 4
rlabel polysilicon 121 -36 121 -36 0 1
rlabel polysilicon 121 -42 121 -42 0 3
rlabel polysilicon 128 -36 128 -36 0 1
rlabel polysilicon 128 -42 128 -42 0 3
rlabel polysilicon 138 -42 138 -42 0 4
rlabel polysilicon 142 -36 142 -36 0 1
rlabel polysilicon 142 -42 142 -42 0 3
rlabel polysilicon 149 -36 149 -36 0 1
rlabel polysilicon 152 -42 152 -42 0 4
rlabel polysilicon 156 -36 156 -36 0 1
rlabel polysilicon 156 -42 156 -42 0 3
rlabel polysilicon 170 -36 170 -36 0 1
rlabel polysilicon 170 -42 170 -42 0 3
rlabel polysilicon 180 -36 180 -36 0 2
rlabel polysilicon 177 -42 177 -42 0 3
rlabel polysilicon 184 -36 184 -36 0 1
rlabel polysilicon 184 -42 184 -42 0 3
rlabel polysilicon 30 -57 30 -57 0 1
rlabel polysilicon 30 -63 30 -63 0 3
rlabel polysilicon 37 -57 37 -57 0 1
rlabel polysilicon 37 -63 37 -63 0 3
rlabel polysilicon 47 -63 47 -63 0 4
rlabel polysilicon 51 -57 51 -57 0 1
rlabel polysilicon 51 -63 51 -63 0 3
rlabel polysilicon 58 -57 58 -57 0 1
rlabel polysilicon 58 -63 58 -63 0 3
rlabel polysilicon 68 -57 68 -57 0 2
rlabel polysilicon 75 -57 75 -57 0 2
rlabel polysilicon 72 -63 72 -63 0 3
rlabel polysilicon 75 -63 75 -63 0 4
rlabel polysilicon 79 -57 79 -57 0 1
rlabel polysilicon 79 -63 79 -63 0 3
rlabel polysilicon 82 -63 82 -63 0 4
rlabel polysilicon 86 -57 86 -57 0 1
rlabel polysilicon 86 -63 86 -63 0 3
rlabel polysilicon 93 -57 93 -57 0 1
rlabel polysilicon 93 -63 93 -63 0 3
rlabel polysilicon 103 -57 103 -57 0 2
rlabel polysilicon 100 -63 100 -63 0 3
rlabel polysilicon 107 -57 107 -57 0 1
rlabel polysilicon 114 -57 114 -57 0 1
rlabel polysilicon 114 -63 114 -63 0 3
rlabel polysilicon 121 -57 121 -57 0 1
rlabel polysilicon 121 -63 121 -63 0 3
rlabel polysilicon 131 -57 131 -57 0 2
rlabel polysilicon 128 -63 128 -63 0 3
rlabel polysilicon 131 -63 131 -63 0 4
rlabel polysilicon 135 -63 135 -63 0 3
rlabel polysilicon 138 -63 138 -63 0 4
rlabel polysilicon 142 -57 142 -57 0 1
rlabel polysilicon 142 -63 142 -63 0 3
rlabel polysilicon 149 -57 149 -57 0 1
rlabel polysilicon 149 -63 149 -63 0 3
rlabel polysilicon 156 -57 156 -57 0 1
rlabel polysilicon 159 -57 159 -57 0 2
rlabel polysilicon 163 -57 163 -57 0 1
rlabel polysilicon 163 -63 163 -63 0 3
rlabel polysilicon 170 -57 170 -57 0 1
rlabel polysilicon 170 -63 170 -63 0 3
rlabel polysilicon 177 -57 177 -57 0 1
rlabel polysilicon 177 -63 177 -63 0 3
rlabel polysilicon 184 -57 184 -57 0 1
rlabel polysilicon 187 -63 187 -63 0 4
rlabel polysilicon 191 -57 191 -57 0 1
rlabel polysilicon 191 -63 191 -63 0 3
rlabel polysilicon 54 -86 54 -86 0 2
rlabel polysilicon 51 -92 51 -92 0 3
rlabel polysilicon 65 -86 65 -86 0 1
rlabel polysilicon 68 -86 68 -86 0 2
rlabel polysilicon 72 -86 72 -86 0 1
rlabel polysilicon 72 -92 72 -92 0 3
rlabel polysilicon 79 -86 79 -86 0 1
rlabel polysilicon 79 -92 79 -92 0 3
rlabel polysilicon 86 -86 86 -86 0 1
rlabel polysilicon 89 -86 89 -86 0 2
rlabel polysilicon 86 -92 86 -92 0 3
rlabel polysilicon 89 -92 89 -92 0 4
rlabel polysilicon 93 -86 93 -86 0 1
rlabel polysilicon 93 -92 93 -92 0 3
rlabel polysilicon 100 -86 100 -86 0 1
rlabel polysilicon 103 -92 103 -92 0 4
rlabel polysilicon 107 -86 107 -86 0 1
rlabel polysilicon 110 -86 110 -86 0 2
rlabel polysilicon 114 -86 114 -86 0 1
rlabel polysilicon 114 -92 114 -92 0 3
rlabel polysilicon 121 -86 121 -86 0 1
rlabel polysilicon 121 -92 121 -92 0 3
rlabel polysilicon 128 -86 128 -86 0 1
rlabel polysilicon 131 -86 131 -86 0 2
rlabel polysilicon 131 -92 131 -92 0 4
rlabel polysilicon 135 -86 135 -86 0 1
rlabel polysilicon 135 -92 135 -92 0 3
rlabel polysilicon 142 -86 142 -86 0 1
rlabel polysilicon 142 -92 142 -92 0 3
rlabel polysilicon 145 -92 145 -92 0 4
rlabel polysilicon 152 -86 152 -86 0 2
rlabel polysilicon 152 -92 152 -92 0 4
rlabel polysilicon 156 -86 156 -86 0 1
rlabel polysilicon 156 -92 156 -92 0 3
rlabel polysilicon 163 -86 163 -86 0 1
rlabel polysilicon 163 -92 163 -92 0 3
rlabel polysilicon 170 -86 170 -86 0 1
rlabel polysilicon 170 -92 170 -92 0 3
rlabel polysilicon 177 -86 177 -86 0 1
rlabel polysilicon 177 -92 177 -92 0 3
rlabel polysilicon 184 -86 184 -86 0 1
rlabel polysilicon 184 -92 184 -92 0 3
rlabel polysilicon 191 -92 191 -92 0 3
rlabel polysilicon 194 -92 194 -92 0 4
rlabel polysilicon 198 -86 198 -86 0 1
rlabel polysilicon 198 -92 198 -92 0 3
rlabel polysilicon 205 -86 205 -86 0 1
rlabel polysilicon 205 -92 205 -92 0 3
rlabel polysilicon 212 -86 212 -86 0 1
rlabel polysilicon 212 -92 212 -92 0 3
rlabel polysilicon 219 -86 219 -86 0 1
rlabel polysilicon 219 -92 219 -92 0 3
rlabel polysilicon 226 -86 226 -86 0 1
rlabel polysilicon 226 -92 226 -92 0 3
rlabel polysilicon 233 -86 233 -86 0 1
rlabel polysilicon 233 -92 233 -92 0 3
rlabel polysilicon 243 -86 243 -86 0 2
rlabel polysilicon 247 -86 247 -86 0 1
rlabel polysilicon 247 -92 247 -92 0 3
rlabel polysilicon 250 -92 250 -92 0 4
rlabel polysilicon 2 -115 2 -115 0 1
rlabel polysilicon 2 -121 2 -121 0 3
rlabel polysilicon 9 -115 9 -115 0 1
rlabel polysilicon 9 -121 9 -121 0 3
rlabel polysilicon 19 -121 19 -121 0 4
rlabel polysilicon 23 -115 23 -115 0 1
rlabel polysilicon 23 -121 23 -121 0 3
rlabel polysilicon 30 -115 30 -115 0 1
rlabel polysilicon 30 -121 30 -121 0 3
rlabel polysilicon 37 -121 37 -121 0 3
rlabel polysilicon 40 -121 40 -121 0 4
rlabel polysilicon 44 -115 44 -115 0 1
rlabel polysilicon 47 -115 47 -115 0 2
rlabel polysilicon 51 -115 51 -115 0 1
rlabel polysilicon 51 -121 51 -121 0 3
rlabel polysilicon 58 -115 58 -115 0 1
rlabel polysilicon 58 -121 58 -121 0 3
rlabel polysilicon 68 -115 68 -115 0 2
rlabel polysilicon 68 -121 68 -121 0 4
rlabel polysilicon 75 -115 75 -115 0 2
rlabel polysilicon 82 -115 82 -115 0 2
rlabel polysilicon 79 -121 79 -121 0 3
rlabel polysilicon 82 -121 82 -121 0 4
rlabel polysilicon 86 -115 86 -115 0 1
rlabel polysilicon 89 -121 89 -121 0 4
rlabel polysilicon 93 -115 93 -115 0 1
rlabel polysilicon 93 -121 93 -121 0 3
rlabel polysilicon 100 -115 100 -115 0 1
rlabel polysilicon 100 -121 100 -121 0 3
rlabel polysilicon 107 -115 107 -115 0 1
rlabel polysilicon 107 -121 107 -121 0 3
rlabel polysilicon 114 -115 114 -115 0 1
rlabel polysilicon 117 -115 117 -115 0 2
rlabel polysilicon 114 -121 114 -121 0 3
rlabel polysilicon 121 -115 121 -115 0 1
rlabel polysilicon 124 -115 124 -115 0 2
rlabel polysilicon 121 -121 121 -121 0 3
rlabel polysilicon 128 -115 128 -115 0 1
rlabel polysilicon 128 -121 128 -121 0 3
rlabel polysilicon 135 -115 135 -115 0 1
rlabel polysilicon 135 -121 135 -121 0 3
rlabel polysilicon 145 -115 145 -115 0 2
rlabel polysilicon 145 -121 145 -121 0 4
rlabel polysilicon 149 -115 149 -115 0 1
rlabel polysilicon 149 -121 149 -121 0 3
rlabel polysilicon 152 -121 152 -121 0 4
rlabel polysilicon 156 -115 156 -115 0 1
rlabel polysilicon 159 -115 159 -115 0 2
rlabel polysilicon 159 -121 159 -121 0 4
rlabel polysilicon 163 -115 163 -115 0 1
rlabel polysilicon 163 -121 163 -121 0 3
rlabel polysilicon 170 -115 170 -115 0 1
rlabel polysilicon 170 -121 170 -121 0 3
rlabel polysilicon 177 -115 177 -115 0 1
rlabel polysilicon 177 -121 177 -121 0 3
rlabel polysilicon 184 -115 184 -115 0 1
rlabel polysilicon 184 -121 184 -121 0 3
rlabel polysilicon 191 -115 191 -115 0 1
rlabel polysilicon 191 -121 191 -121 0 3
rlabel polysilicon 198 -115 198 -115 0 1
rlabel polysilicon 198 -121 198 -121 0 3
rlabel polysilicon 205 -115 205 -115 0 1
rlabel polysilicon 205 -121 205 -121 0 3
rlabel polysilicon 212 -115 212 -115 0 1
rlabel polysilicon 212 -121 212 -121 0 3
rlabel polysilicon 219 -115 219 -115 0 1
rlabel polysilicon 219 -121 219 -121 0 3
rlabel polysilicon 226 -115 226 -115 0 1
rlabel polysilicon 226 -121 226 -121 0 3
rlabel polysilicon 233 -115 233 -115 0 1
rlabel polysilicon 233 -121 233 -121 0 3
rlabel polysilicon 240 -115 240 -115 0 1
rlabel polysilicon 240 -121 240 -121 0 3
rlabel polysilicon 247 -115 247 -115 0 1
rlabel polysilicon 247 -121 247 -121 0 3
rlabel polysilicon 254 -115 254 -115 0 1
rlabel polysilicon 2 -160 2 -160 0 1
rlabel polysilicon 2 -166 2 -166 0 3
rlabel polysilicon 9 -160 9 -160 0 1
rlabel polysilicon 9 -166 9 -166 0 3
rlabel polysilicon 19 -160 19 -160 0 2
rlabel polysilicon 26 -166 26 -166 0 4
rlabel polysilicon 30 -160 30 -160 0 1
rlabel polysilicon 33 -160 33 -160 0 2
rlabel polysilicon 40 -160 40 -160 0 2
rlabel polysilicon 40 -166 40 -166 0 4
rlabel polysilicon 47 -160 47 -160 0 2
rlabel polysilicon 47 -166 47 -166 0 4
rlabel polysilicon 51 -160 51 -160 0 1
rlabel polysilicon 51 -166 51 -166 0 3
rlabel polysilicon 58 -160 58 -160 0 1
rlabel polysilicon 58 -166 58 -166 0 3
rlabel polysilicon 65 -160 65 -160 0 1
rlabel polysilicon 65 -166 65 -166 0 3
rlabel polysilicon 72 -160 72 -160 0 1
rlabel polysilicon 72 -166 72 -166 0 3
rlabel polysilicon 79 -166 79 -166 0 3
rlabel polysilicon 82 -166 82 -166 0 4
rlabel polysilicon 86 -160 86 -160 0 1
rlabel polysilicon 89 -160 89 -160 0 2
rlabel polysilicon 86 -166 86 -166 0 3
rlabel polysilicon 89 -166 89 -166 0 4
rlabel polysilicon 96 -166 96 -166 0 4
rlabel polysilicon 100 -160 100 -160 0 1
rlabel polysilicon 100 -166 100 -166 0 3
rlabel polysilicon 107 -160 107 -160 0 1
rlabel polysilicon 107 -166 107 -166 0 3
rlabel polysilicon 110 -166 110 -166 0 4
rlabel polysilicon 114 -160 114 -160 0 1
rlabel polysilicon 117 -160 117 -160 0 2
rlabel polysilicon 114 -166 114 -166 0 3
rlabel polysilicon 117 -166 117 -166 0 4
rlabel polysilicon 121 -160 121 -160 0 1
rlabel polysilicon 121 -166 121 -166 0 3
rlabel polysilicon 128 -160 128 -160 0 1
rlabel polysilicon 128 -166 128 -166 0 3
rlabel polysilicon 135 -160 135 -160 0 1
rlabel polysilicon 138 -160 138 -160 0 2
rlabel polysilicon 135 -166 135 -166 0 3
rlabel polysilicon 138 -166 138 -166 0 4
rlabel polysilicon 142 -160 142 -160 0 1
rlabel polysilicon 142 -166 142 -166 0 3
rlabel polysilicon 149 -160 149 -160 0 1
rlabel polysilicon 149 -166 149 -166 0 3
rlabel polysilicon 156 -160 156 -160 0 1
rlabel polysilicon 159 -166 159 -166 0 4
rlabel polysilicon 163 -160 163 -160 0 1
rlabel polysilicon 163 -166 163 -166 0 3
rlabel polysilicon 170 -160 170 -160 0 1
rlabel polysilicon 170 -166 170 -166 0 3
rlabel polysilicon 177 -160 177 -160 0 1
rlabel polysilicon 177 -166 177 -166 0 3
rlabel polysilicon 187 -160 187 -160 0 2
rlabel polysilicon 184 -166 184 -166 0 3
rlabel polysilicon 191 -160 191 -160 0 1
rlabel polysilicon 191 -166 191 -166 0 3
rlabel polysilicon 198 -160 198 -160 0 1
rlabel polysilicon 198 -166 198 -166 0 3
rlabel polysilicon 205 -160 205 -160 0 1
rlabel polysilicon 205 -166 205 -166 0 3
rlabel polysilicon 212 -160 212 -160 0 1
rlabel polysilicon 212 -166 212 -166 0 3
rlabel polysilicon 219 -160 219 -160 0 1
rlabel polysilicon 219 -166 219 -166 0 3
rlabel polysilicon 226 -160 226 -160 0 1
rlabel polysilicon 226 -166 226 -166 0 3
rlabel polysilicon 233 -160 233 -160 0 1
rlabel polysilicon 233 -166 233 -166 0 3
rlabel polysilicon 240 -160 240 -160 0 1
rlabel polysilicon 240 -166 240 -166 0 3
rlabel polysilicon 247 -160 247 -160 0 1
rlabel polysilicon 247 -166 247 -166 0 3
rlabel polysilicon 254 -160 254 -160 0 1
rlabel polysilicon 254 -166 254 -166 0 3
rlabel polysilicon 261 -160 261 -160 0 1
rlabel polysilicon 261 -166 261 -166 0 3
rlabel polysilicon 268 -160 268 -160 0 1
rlabel polysilicon 268 -166 268 -166 0 3
rlabel polysilicon 275 -160 275 -160 0 1
rlabel polysilicon 275 -166 275 -166 0 3
rlabel polysilicon 23 -191 23 -191 0 1
rlabel polysilicon 23 -197 23 -197 0 3
rlabel polysilicon 30 -191 30 -191 0 1
rlabel polysilicon 30 -197 30 -197 0 3
rlabel polysilicon 40 -191 40 -191 0 2
rlabel polysilicon 37 -197 37 -197 0 3
rlabel polysilicon 44 -191 44 -191 0 1
rlabel polysilicon 44 -197 44 -197 0 3
rlabel polysilicon 47 -197 47 -197 0 4
rlabel polysilicon 51 -191 51 -191 0 1
rlabel polysilicon 51 -197 51 -197 0 3
rlabel polysilicon 58 -191 58 -191 0 1
rlabel polysilicon 58 -197 58 -197 0 3
rlabel polysilicon 65 -191 65 -191 0 1
rlabel polysilicon 68 -197 68 -197 0 4
rlabel polysilicon 72 -191 72 -191 0 1
rlabel polysilicon 72 -197 72 -197 0 3
rlabel polysilicon 82 -191 82 -191 0 2
rlabel polysilicon 86 -191 86 -191 0 1
rlabel polysilicon 86 -197 86 -197 0 3
rlabel polysilicon 93 -197 93 -197 0 3
rlabel polysilicon 96 -197 96 -197 0 4
rlabel polysilicon 103 -191 103 -191 0 2
rlabel polysilicon 103 -197 103 -197 0 4
rlabel polysilicon 107 -191 107 -191 0 1
rlabel polysilicon 107 -197 107 -197 0 3
rlabel polysilicon 110 -197 110 -197 0 4
rlabel polysilicon 114 -191 114 -191 0 1
rlabel polysilicon 117 -197 117 -197 0 4
rlabel polysilicon 121 -191 121 -191 0 1
rlabel polysilicon 121 -197 121 -197 0 3
rlabel polysilicon 128 -191 128 -191 0 1
rlabel polysilicon 128 -197 128 -197 0 3
rlabel polysilicon 135 -191 135 -191 0 1
rlabel polysilicon 138 -191 138 -191 0 2
rlabel polysilicon 135 -197 135 -197 0 3
rlabel polysilicon 142 -197 142 -197 0 3
rlabel polysilicon 145 -197 145 -197 0 4
rlabel polysilicon 149 -191 149 -191 0 1
rlabel polysilicon 152 -191 152 -191 0 2
rlabel polysilicon 149 -197 149 -197 0 3
rlabel polysilicon 152 -197 152 -197 0 4
rlabel polysilicon 156 -191 156 -191 0 1
rlabel polysilicon 156 -197 156 -197 0 3
rlabel polysilicon 163 -191 163 -191 0 1
rlabel polysilicon 163 -197 163 -197 0 3
rlabel polysilicon 170 -191 170 -191 0 1
rlabel polysilicon 170 -197 170 -197 0 3
rlabel polysilicon 177 -191 177 -191 0 1
rlabel polysilicon 177 -197 177 -197 0 3
rlabel polysilicon 187 -191 187 -191 0 2
rlabel polysilicon 187 -197 187 -197 0 4
rlabel polysilicon 194 -191 194 -191 0 2
rlabel polysilicon 194 -197 194 -197 0 4
rlabel polysilicon 198 -191 198 -191 0 1
rlabel polysilicon 198 -197 198 -197 0 3
rlabel polysilicon 205 -191 205 -191 0 1
rlabel polysilicon 205 -197 205 -197 0 3
rlabel polysilicon 212 -191 212 -191 0 1
rlabel polysilicon 212 -197 212 -197 0 3
rlabel polysilicon 219 -191 219 -191 0 1
rlabel polysilicon 219 -197 219 -197 0 3
rlabel polysilicon 226 -191 226 -191 0 1
rlabel polysilicon 226 -197 226 -197 0 3
rlabel polysilicon 233 -191 233 -191 0 1
rlabel polysilicon 233 -197 233 -197 0 3
rlabel polysilicon 240 -191 240 -191 0 1
rlabel polysilicon 240 -197 240 -197 0 3
rlabel polysilicon 247 -191 247 -191 0 1
rlabel polysilicon 247 -197 247 -197 0 3
rlabel polysilicon 254 -191 254 -191 0 1
rlabel polysilicon 254 -197 254 -197 0 3
rlabel polysilicon 261 -191 261 -191 0 1
rlabel polysilicon 261 -197 261 -197 0 3
rlabel polysilicon 282 -197 282 -197 0 3
rlabel polysilicon 30 -226 30 -226 0 1
rlabel polysilicon 37 -226 37 -226 0 1
rlabel polysilicon 37 -232 37 -232 0 3
rlabel polysilicon 44 -226 44 -226 0 1
rlabel polysilicon 51 -226 51 -226 0 1
rlabel polysilicon 51 -232 51 -232 0 3
rlabel polysilicon 58 -226 58 -226 0 1
rlabel polysilicon 58 -232 58 -232 0 3
rlabel polysilicon 65 -226 65 -226 0 1
rlabel polysilicon 65 -232 65 -232 0 3
rlabel polysilicon 75 -232 75 -232 0 4
rlabel polysilicon 82 -226 82 -226 0 2
rlabel polysilicon 79 -232 79 -232 0 3
rlabel polysilicon 86 -226 86 -226 0 1
rlabel polysilicon 86 -232 86 -232 0 3
rlabel polysilicon 93 -226 93 -226 0 1
rlabel polysilicon 96 -226 96 -226 0 2
rlabel polysilicon 93 -232 93 -232 0 3
rlabel polysilicon 100 -226 100 -226 0 1
rlabel polysilicon 100 -232 100 -232 0 3
rlabel polysilicon 107 -226 107 -226 0 1
rlabel polysilicon 107 -232 107 -232 0 3
rlabel polysilicon 114 -226 114 -226 0 1
rlabel polysilicon 117 -226 117 -226 0 2
rlabel polysilicon 114 -232 114 -232 0 3
rlabel polysilicon 117 -232 117 -232 0 4
rlabel polysilicon 121 -226 121 -226 0 1
rlabel polysilicon 121 -232 121 -232 0 3
rlabel polysilicon 128 -226 128 -226 0 1
rlabel polysilicon 128 -232 128 -232 0 3
rlabel polysilicon 135 -226 135 -226 0 1
rlabel polysilicon 138 -226 138 -226 0 2
rlabel polysilicon 142 -226 142 -226 0 1
rlabel polysilicon 142 -232 142 -232 0 3
rlabel polysilicon 149 -226 149 -226 0 1
rlabel polysilicon 152 -226 152 -226 0 2
rlabel polysilicon 159 -226 159 -226 0 2
rlabel polysilicon 156 -232 156 -232 0 3
rlabel polysilicon 159 -232 159 -232 0 4
rlabel polysilicon 163 -226 163 -226 0 1
rlabel polysilicon 163 -232 163 -232 0 3
rlabel polysilicon 170 -226 170 -226 0 1
rlabel polysilicon 170 -232 170 -232 0 3
rlabel polysilicon 177 -226 177 -226 0 1
rlabel polysilicon 180 -226 180 -226 0 2
rlabel polysilicon 184 -226 184 -226 0 1
rlabel polysilicon 184 -232 184 -232 0 3
rlabel polysilicon 191 -226 191 -226 0 1
rlabel polysilicon 194 -226 194 -226 0 2
rlabel polysilicon 191 -232 191 -232 0 3
rlabel polysilicon 198 -226 198 -226 0 1
rlabel polysilicon 198 -232 198 -232 0 3
rlabel polysilicon 205 -226 205 -226 0 1
rlabel polysilicon 205 -232 205 -232 0 3
rlabel polysilicon 212 -226 212 -226 0 1
rlabel polysilicon 212 -232 212 -232 0 3
rlabel polysilicon 219 -226 219 -226 0 1
rlabel polysilicon 219 -232 219 -232 0 3
rlabel polysilicon 226 -226 226 -226 0 1
rlabel polysilicon 226 -232 226 -232 0 3
rlabel polysilicon 233 -226 233 -226 0 1
rlabel polysilicon 233 -232 233 -232 0 3
rlabel polysilicon 240 -226 240 -226 0 1
rlabel polysilicon 240 -232 240 -232 0 3
rlabel polysilicon 247 -226 247 -226 0 1
rlabel polysilicon 247 -232 247 -232 0 3
rlabel polysilicon 254 -226 254 -226 0 1
rlabel polysilicon 254 -232 254 -232 0 3
rlabel polysilicon 261 -226 261 -226 0 1
rlabel polysilicon 264 -226 264 -226 0 2
rlabel polysilicon 261 -232 261 -232 0 3
rlabel polysilicon 264 -232 264 -232 0 4
rlabel polysilicon 271 -226 271 -226 0 2
rlabel polysilicon 278 -226 278 -226 0 2
rlabel polysilicon 275 -232 275 -232 0 3
rlabel polysilicon 282 -226 282 -226 0 1
rlabel polysilicon 282 -232 282 -232 0 3
rlabel polysilicon 289 -226 289 -226 0 1
rlabel polysilicon 289 -232 289 -232 0 3
rlabel polysilicon 16 -257 16 -257 0 1
rlabel polysilicon 16 -263 16 -263 0 3
rlabel polysilicon 26 -263 26 -263 0 4
rlabel polysilicon 30 -257 30 -257 0 1
rlabel polysilicon 30 -263 30 -263 0 3
rlabel polysilicon 37 -257 37 -257 0 1
rlabel polysilicon 37 -263 37 -263 0 3
rlabel polysilicon 44 -257 44 -257 0 1
rlabel polysilicon 44 -263 44 -263 0 3
rlabel polysilicon 47 -263 47 -263 0 4
rlabel polysilicon 51 -263 51 -263 0 3
rlabel polysilicon 54 -263 54 -263 0 4
rlabel polysilicon 58 -257 58 -257 0 1
rlabel polysilicon 58 -263 58 -263 0 3
rlabel polysilicon 65 -257 65 -257 0 1
rlabel polysilicon 65 -263 65 -263 0 3
rlabel polysilicon 72 -257 72 -257 0 1
rlabel polysilicon 72 -263 72 -263 0 3
rlabel polysilicon 79 -257 79 -257 0 1
rlabel polysilicon 79 -263 79 -263 0 3
rlabel polysilicon 86 -257 86 -257 0 1
rlabel polysilicon 86 -263 86 -263 0 3
rlabel polysilicon 93 -257 93 -257 0 1
rlabel polysilicon 93 -263 93 -263 0 3
rlabel polysilicon 103 -257 103 -257 0 2
rlabel polysilicon 100 -263 100 -263 0 3
rlabel polysilicon 103 -263 103 -263 0 4
rlabel polysilicon 107 -257 107 -257 0 1
rlabel polysilicon 107 -263 107 -263 0 3
rlabel polysilicon 114 -257 114 -257 0 1
rlabel polysilicon 117 -257 117 -257 0 2
rlabel polysilicon 114 -263 114 -263 0 3
rlabel polysilicon 117 -263 117 -263 0 4
rlabel polysilicon 121 -257 121 -257 0 1
rlabel polysilicon 121 -263 121 -263 0 3
rlabel polysilicon 128 -257 128 -257 0 1
rlabel polysilicon 128 -263 128 -263 0 3
rlabel polysilicon 135 -257 135 -257 0 1
rlabel polysilicon 135 -263 135 -263 0 3
rlabel polysilicon 142 -257 142 -257 0 1
rlabel polysilicon 142 -263 142 -263 0 3
rlabel polysilicon 149 -257 149 -257 0 1
rlabel polysilicon 149 -263 149 -263 0 3
rlabel polysilicon 156 -257 156 -257 0 1
rlabel polysilicon 156 -263 156 -263 0 3
rlabel polysilicon 163 -257 163 -257 0 1
rlabel polysilicon 163 -263 163 -263 0 3
rlabel polysilicon 170 -257 170 -257 0 1
rlabel polysilicon 173 -257 173 -257 0 2
rlabel polysilicon 173 -263 173 -263 0 4
rlabel polysilicon 177 -257 177 -257 0 1
rlabel polysilicon 180 -257 180 -257 0 2
rlabel polysilicon 177 -263 177 -263 0 3
rlabel polysilicon 180 -263 180 -263 0 4
rlabel polysilicon 184 -257 184 -257 0 1
rlabel polysilicon 184 -263 184 -263 0 3
rlabel polysilicon 191 -257 191 -257 0 1
rlabel polysilicon 191 -263 191 -263 0 3
rlabel polysilicon 198 -257 198 -257 0 1
rlabel polysilicon 198 -263 198 -263 0 3
rlabel polysilicon 205 -257 205 -257 0 1
rlabel polysilicon 205 -263 205 -263 0 3
rlabel polysilicon 212 -257 212 -257 0 1
rlabel polysilicon 212 -263 212 -263 0 3
rlabel polysilicon 219 -257 219 -257 0 1
rlabel polysilicon 219 -263 219 -263 0 3
rlabel polysilicon 226 -257 226 -257 0 1
rlabel polysilicon 226 -263 226 -263 0 3
rlabel polysilicon 233 -257 233 -257 0 1
rlabel polysilicon 233 -263 233 -263 0 3
rlabel polysilicon 240 -257 240 -257 0 1
rlabel polysilicon 240 -263 240 -263 0 3
rlabel polysilicon 247 -257 247 -257 0 1
rlabel polysilicon 247 -263 247 -263 0 3
rlabel polysilicon 254 -257 254 -257 0 1
rlabel polysilicon 254 -263 254 -263 0 3
rlabel polysilicon 282 -257 282 -257 0 1
rlabel polysilicon 282 -263 282 -263 0 3
rlabel polysilicon 289 -263 289 -263 0 3
rlabel polysilicon 65 -284 65 -284 0 1
rlabel polysilicon 65 -290 65 -290 0 3
rlabel polysilicon 72 -284 72 -284 0 1
rlabel polysilicon 72 -290 72 -290 0 3
rlabel polysilicon 82 -290 82 -290 0 4
rlabel polysilicon 86 -284 86 -284 0 1
rlabel polysilicon 89 -284 89 -284 0 2
rlabel polysilicon 86 -290 86 -290 0 3
rlabel polysilicon 89 -290 89 -290 0 4
rlabel polysilicon 93 -284 93 -284 0 1
rlabel polysilicon 96 -284 96 -284 0 2
rlabel polysilicon 96 -290 96 -290 0 4
rlabel polysilicon 103 -284 103 -284 0 2
rlabel polysilicon 103 -290 103 -290 0 4
rlabel polysilicon 107 -284 107 -284 0 1
rlabel polysilicon 107 -290 107 -290 0 3
rlabel polysilicon 114 -290 114 -290 0 3
rlabel polysilicon 117 -290 117 -290 0 4
rlabel polysilicon 121 -284 121 -284 0 1
rlabel polysilicon 121 -290 121 -290 0 3
rlabel polysilicon 128 -284 128 -284 0 1
rlabel polysilicon 128 -290 128 -290 0 3
rlabel polysilicon 135 -284 135 -284 0 1
rlabel polysilicon 135 -290 135 -290 0 3
rlabel polysilicon 142 -284 142 -284 0 1
rlabel polysilicon 142 -290 142 -290 0 3
rlabel polysilicon 149 -284 149 -284 0 1
rlabel polysilicon 149 -290 149 -290 0 3
rlabel polysilicon 156 -284 156 -284 0 1
rlabel polysilicon 156 -290 156 -290 0 3
rlabel polysilicon 166 -284 166 -284 0 2
rlabel polysilicon 163 -290 163 -290 0 3
rlabel polysilicon 170 -284 170 -284 0 1
rlabel polysilicon 170 -290 170 -290 0 3
rlabel polysilicon 184 -290 184 -290 0 3
rlabel polysilicon 191 -284 191 -284 0 1
rlabel polysilicon 194 -284 194 -284 0 2
rlabel polysilicon 191 -290 191 -290 0 3
rlabel polysilicon 194 -290 194 -290 0 4
rlabel polysilicon 198 -284 198 -284 0 1
rlabel polysilicon 198 -290 198 -290 0 3
rlabel polysilicon 205 -284 205 -284 0 1
rlabel polysilicon 208 -284 208 -284 0 2
rlabel polysilicon 205 -290 205 -290 0 3
rlabel polysilicon 240 -284 240 -284 0 1
rlabel polysilicon 240 -290 240 -290 0 3
rlabel polysilicon 247 -284 247 -284 0 1
rlabel polysilicon 250 -290 250 -290 0 4
rlabel polysilicon 254 -284 254 -284 0 1
rlabel polysilicon 254 -290 254 -290 0 3
rlabel polysilicon 51 -307 51 -307 0 1
rlabel polysilicon 51 -313 51 -313 0 3
rlabel polysilicon 61 -313 61 -313 0 4
rlabel polysilicon 65 -307 65 -307 0 1
rlabel polysilicon 65 -313 65 -313 0 3
rlabel polysilicon 75 -307 75 -307 0 2
rlabel polysilicon 72 -313 72 -313 0 3
rlabel polysilicon 75 -313 75 -313 0 4
rlabel polysilicon 82 -307 82 -307 0 2
rlabel polysilicon 86 -307 86 -307 0 1
rlabel polysilicon 89 -307 89 -307 0 2
rlabel polysilicon 89 -313 89 -313 0 4
rlabel polysilicon 96 -307 96 -307 0 2
rlabel polysilicon 93 -313 93 -313 0 3
rlabel polysilicon 103 -307 103 -307 0 2
rlabel polysilicon 100 -313 100 -313 0 3
rlabel polysilicon 107 -307 107 -307 0 1
rlabel polysilicon 110 -307 110 -307 0 2
rlabel polysilicon 107 -313 107 -313 0 3
rlabel polysilicon 114 -307 114 -307 0 1
rlabel polysilicon 117 -307 117 -307 0 2
rlabel polysilicon 114 -313 114 -313 0 3
rlabel polysilicon 117 -313 117 -313 0 4
rlabel polysilicon 121 -307 121 -307 0 1
rlabel polysilicon 121 -313 121 -313 0 3
rlabel polysilicon 128 -307 128 -307 0 1
rlabel polysilicon 128 -313 128 -313 0 3
rlabel polysilicon 138 -307 138 -307 0 2
rlabel polysilicon 135 -313 135 -313 0 3
rlabel polysilicon 138 -313 138 -313 0 4
rlabel polysilicon 142 -307 142 -307 0 1
rlabel polysilicon 142 -313 142 -313 0 3
rlabel polysilicon 149 -307 149 -307 0 1
rlabel polysilicon 149 -313 149 -313 0 3
rlabel polysilicon 156 -307 156 -307 0 1
rlabel polysilicon 156 -313 156 -313 0 3
rlabel polysilicon 163 -307 163 -307 0 1
rlabel polysilicon 163 -313 163 -313 0 3
rlabel polysilicon 170 -307 170 -307 0 1
rlabel polysilicon 170 -313 170 -313 0 3
rlabel polysilicon 177 -307 177 -307 0 1
rlabel polysilicon 177 -313 177 -313 0 3
rlabel polysilicon 219 -307 219 -307 0 1
rlabel polysilicon 219 -313 219 -313 0 3
rlabel polysilicon 226 -313 226 -313 0 3
rlabel polysilicon 233 -307 233 -307 0 1
rlabel polysilicon 233 -313 233 -313 0 3
rlabel polysilicon 236 -313 236 -313 0 4
rlabel polysilicon 240 -307 240 -307 0 1
rlabel polysilicon 240 -313 240 -313 0 3
rlabel polysilicon 37 -336 37 -336 0 1
rlabel polysilicon 37 -342 37 -342 0 3
rlabel polysilicon 44 -336 44 -336 0 1
rlabel polysilicon 44 -342 44 -342 0 3
rlabel polysilicon 51 -336 51 -336 0 1
rlabel polysilicon 51 -342 51 -342 0 3
rlabel polysilicon 61 -336 61 -336 0 2
rlabel polysilicon 58 -342 58 -342 0 3
rlabel polysilicon 65 -336 65 -336 0 1
rlabel polysilicon 65 -342 65 -342 0 3
rlabel polysilicon 72 -336 72 -336 0 1
rlabel polysilicon 72 -342 72 -342 0 3
rlabel polysilicon 79 -336 79 -336 0 1
rlabel polysilicon 79 -342 79 -342 0 3
rlabel polysilicon 86 -336 86 -336 0 1
rlabel polysilicon 89 -336 89 -336 0 2
rlabel polysilicon 93 -336 93 -336 0 1
rlabel polysilicon 96 -336 96 -336 0 2
rlabel polysilicon 93 -342 93 -342 0 3
rlabel polysilicon 96 -342 96 -342 0 4
rlabel polysilicon 100 -336 100 -336 0 1
rlabel polysilicon 100 -342 100 -342 0 3
rlabel polysilicon 103 -342 103 -342 0 4
rlabel polysilicon 107 -336 107 -336 0 1
rlabel polysilicon 107 -342 107 -342 0 3
rlabel polysilicon 117 -336 117 -336 0 2
rlabel polysilicon 114 -342 114 -342 0 3
rlabel polysilicon 117 -342 117 -342 0 4
rlabel polysilicon 121 -336 121 -336 0 1
rlabel polysilicon 121 -342 121 -342 0 3
rlabel polysilicon 128 -336 128 -336 0 1
rlabel polysilicon 131 -336 131 -336 0 2
rlabel polysilicon 131 -342 131 -342 0 4
rlabel polysilicon 135 -336 135 -336 0 1
rlabel polysilicon 138 -336 138 -336 0 2
rlabel polysilicon 138 -342 138 -342 0 4
rlabel polysilicon 142 -336 142 -336 0 1
rlabel polysilicon 142 -342 142 -342 0 3
rlabel polysilicon 145 -342 145 -342 0 4
rlabel polysilicon 149 -336 149 -336 0 1
rlabel polysilicon 149 -342 149 -342 0 3
rlabel polysilicon 159 -336 159 -336 0 2
rlabel polysilicon 156 -342 156 -342 0 3
rlabel polysilicon 163 -336 163 -336 0 1
rlabel polysilicon 163 -342 163 -342 0 3
rlabel polysilicon 170 -336 170 -336 0 1
rlabel polysilicon 170 -342 170 -342 0 3
rlabel polysilicon 177 -336 177 -336 0 1
rlabel polysilicon 177 -342 177 -342 0 3
rlabel polysilicon 184 -336 184 -336 0 1
rlabel polysilicon 184 -342 184 -342 0 3
rlabel polysilicon 191 -336 191 -336 0 1
rlabel polysilicon 191 -342 191 -342 0 3
rlabel polysilicon 198 -336 198 -336 0 1
rlabel polysilicon 198 -342 198 -342 0 3
rlabel polysilicon 205 -336 205 -336 0 1
rlabel polysilicon 205 -342 205 -342 0 3
rlabel polysilicon 212 -342 212 -342 0 3
rlabel polysilicon 215 -342 215 -342 0 4
rlabel polysilicon 219 -336 219 -336 0 1
rlabel polysilicon 219 -342 219 -342 0 3
rlabel polysilicon 58 -363 58 -363 0 1
rlabel polysilicon 58 -369 58 -369 0 3
rlabel polysilicon 65 -363 65 -363 0 1
rlabel polysilicon 65 -369 65 -369 0 3
rlabel polysilicon 72 -363 72 -363 0 1
rlabel polysilicon 72 -369 72 -369 0 3
rlabel polysilicon 79 -363 79 -363 0 1
rlabel polysilicon 79 -369 79 -369 0 3
rlabel polysilicon 86 -363 86 -363 0 1
rlabel polysilicon 86 -369 86 -369 0 3
rlabel polysilicon 96 -363 96 -363 0 2
rlabel polysilicon 103 -363 103 -363 0 2
rlabel polysilicon 100 -369 100 -369 0 3
rlabel polysilicon 110 -363 110 -363 0 2
rlabel polysilicon 107 -369 107 -369 0 3
rlabel polysilicon 114 -369 114 -369 0 3
rlabel polysilicon 117 -369 117 -369 0 4
rlabel polysilicon 121 -363 121 -363 0 1
rlabel polysilicon 121 -369 121 -369 0 3
rlabel polysilicon 128 -363 128 -363 0 1
rlabel polysilicon 128 -369 128 -369 0 3
rlabel polysilicon 135 -363 135 -363 0 1
rlabel polysilicon 135 -369 135 -369 0 3
rlabel polysilicon 142 -363 142 -363 0 1
rlabel polysilicon 142 -369 142 -369 0 3
rlabel polysilicon 145 -369 145 -369 0 4
rlabel polysilicon 149 -363 149 -363 0 1
rlabel polysilicon 149 -369 149 -369 0 3
rlabel polysilicon 156 -369 156 -369 0 3
rlabel polysilicon 163 -363 163 -363 0 1
rlabel polysilicon 163 -369 163 -369 0 3
rlabel polysilicon 170 -363 170 -363 0 1
rlabel polysilicon 177 -363 177 -363 0 1
rlabel polysilicon 177 -369 177 -369 0 3
rlabel polysilicon 184 -363 184 -363 0 1
rlabel polysilicon 184 -369 184 -369 0 3
rlabel polysilicon 194 -363 194 -363 0 2
rlabel polysilicon 198 -363 198 -363 0 1
rlabel polysilicon 198 -369 198 -369 0 3
rlabel polysilicon 72 -386 72 -386 0 1
rlabel polysilicon 72 -392 72 -392 0 3
rlabel polysilicon 79 -386 79 -386 0 1
rlabel polysilicon 79 -392 79 -392 0 3
rlabel polysilicon 86 -386 86 -386 0 1
rlabel polysilicon 86 -392 86 -392 0 3
rlabel polysilicon 93 -386 93 -386 0 1
rlabel polysilicon 96 -386 96 -386 0 2
rlabel polysilicon 100 -386 100 -386 0 1
rlabel polysilicon 103 -386 103 -386 0 2
rlabel polysilicon 100 -392 100 -392 0 3
rlabel polysilicon 107 -386 107 -386 0 1
rlabel polysilicon 107 -392 107 -392 0 3
rlabel polysilicon 114 -392 114 -392 0 3
rlabel polysilicon 117 -392 117 -392 0 4
rlabel polysilicon 121 -386 121 -386 0 1
rlabel polysilicon 124 -386 124 -386 0 2
rlabel polysilicon 121 -392 121 -392 0 3
rlabel polysilicon 128 -386 128 -386 0 1
rlabel polysilicon 128 -392 128 -392 0 3
rlabel polysilicon 138 -386 138 -386 0 2
rlabel polysilicon 138 -392 138 -392 0 4
rlabel polysilicon 142 -386 142 -386 0 1
rlabel polysilicon 142 -392 142 -392 0 3
rlabel polysilicon 149 -386 149 -386 0 1
rlabel polysilicon 149 -392 149 -392 0 3
rlabel polysilicon 156 -386 156 -386 0 1
rlabel polysilicon 156 -392 156 -392 0 3
rlabel polysilicon 163 -386 163 -386 0 1
rlabel polysilicon 163 -392 163 -392 0 3
rlabel polysilicon 170 -386 170 -386 0 1
rlabel polysilicon 173 -386 173 -386 0 2
rlabel polysilicon 170 -392 170 -392 0 3
rlabel polysilicon 79 -407 79 -407 0 1
rlabel polysilicon 86 -407 86 -407 0 1
rlabel polysilicon 86 -413 86 -413 0 3
rlabel polysilicon 93 -407 93 -407 0 1
rlabel polysilicon 93 -413 93 -413 0 3
rlabel polysilicon 100 -413 100 -413 0 3
rlabel polysilicon 107 -407 107 -407 0 1
rlabel polysilicon 107 -413 107 -413 0 3
rlabel polysilicon 117 -407 117 -407 0 2
rlabel polysilicon 117 -413 117 -413 0 4
rlabel polysilicon 121 -407 121 -407 0 1
rlabel polysilicon 121 -413 121 -413 0 3
rlabel polysilicon 128 -407 128 -407 0 1
rlabel polysilicon 131 -407 131 -407 0 2
rlabel polysilicon 142 -407 142 -407 0 1
rlabel polysilicon 145 -407 145 -407 0 2
rlabel polysilicon 156 -407 156 -407 0 1
rlabel polysilicon 156 -413 156 -413 0 3
rlabel polysilicon 163 -407 163 -407 0 1
rlabel polysilicon 173 -407 173 -407 0 2
rlabel polysilicon 89 -426 89 -426 0 4
rlabel polysilicon 93 -420 93 -420 0 1
rlabel polysilicon 93 -426 93 -426 0 3
rlabel polysilicon 117 -426 117 -426 0 4
rlabel polysilicon 121 -420 121 -420 0 1
rlabel polysilicon 121 -426 121 -426 0 3
rlabel polysilicon 163 -420 163 -420 0 1
rlabel polysilicon 163 -426 163 -426 0 3
rlabel polysilicon 170 -426 170 -426 0 3
rlabel metal2 93 1 93 1 0 net=531
rlabel metal2 177 1 177 1 0 net=287
rlabel metal2 191 1 191 1 0 net=515
rlabel metal2 100 -1 100 -1 0 net=419
rlabel metal2 58 -12 58 -12 0 net=491
rlabel metal2 75 -12 75 -12 0 net=88
rlabel metal2 75 -12 75 -12 0 net=88
rlabel metal2 79 -12 79 -12 0 net=571
rlabel metal2 93 -12 93 -12 0 net=532
rlabel metal2 117 -12 117 -12 0 net=293
rlabel metal2 184 -12 184 -12 0 net=288
rlabel metal2 198 -12 198 -12 0 net=517
rlabel metal2 93 -14 93 -14 0 net=201
rlabel metal2 107 -14 107 -14 0 net=420
rlabel metal2 177 -14 177 -14 0 net=597
rlabel metal2 79 -25 79 -25 0 net=572
rlabel metal2 93 -25 93 -25 0 net=202
rlabel metal2 128 -25 128 -25 0 net=295
rlabel metal2 128 -25 128 -25 0 net=295
rlabel metal2 142 -25 142 -25 0 net=533
rlabel metal2 170 -25 170 -25 0 net=599
rlabel metal2 180 -25 180 -25 0 net=543
rlabel metal2 198 -25 198 -25 0 net=518
rlabel metal2 51 -27 51 -27 0 net=639
rlabel metal2 96 -27 96 -27 0 net=595
rlabel metal2 65 -29 65 -29 0 net=26
rlabel metal2 100 -29 100 -29 0 net=255
rlabel metal2 58 -31 58 -31 0 net=492
rlabel metal2 58 -33 58 -33 0 net=385
rlabel metal2 44 -44 44 -44 0 net=640
rlabel metal2 58 -44 58 -44 0 net=386
rlabel metal2 86 -44 86 -44 0 net=29
rlabel metal2 138 -44 138 -44 0 net=495
rlabel metal2 156 -44 156 -44 0 net=596
rlabel metal2 156 -44 156 -44 0 net=596
rlabel metal2 159 -44 159 -44 0 net=629
rlabel metal2 30 -46 30 -46 0 net=635
rlabel metal2 103 -46 103 -46 0 net=256
rlabel metal2 142 -46 142 -46 0 net=535
rlabel metal2 170 -46 170 -46 0 net=600
rlabel metal2 184 -46 184 -46 0 net=544
rlabel metal2 184 -46 184 -46 0 net=544
rlabel metal2 37 -48 37 -48 0 net=583
rlabel metal2 107 -48 107 -48 0 net=296
rlabel metal2 152 -48 152 -48 0 net=567
rlabel metal2 51 -50 51 -50 0 net=477
rlabel metal2 68 -50 68 -50 0 net=455
rlabel metal2 107 -50 107 -50 0 net=257
rlabel metal2 117 -50 117 -50 0 net=429
rlabel metal2 58 -52 58 -52 0 net=291
rlabel metal2 75 -52 75 -52 0 net=445
rlabel metal2 110 -52 110 -52 0 net=407
rlabel metal2 121 -54 121 -54 0 net=249
rlabel metal2 30 -65 30 -65 0 net=636
rlabel metal2 82 -65 82 -65 0 net=447
rlabel metal2 187 -65 187 -65 0 net=627
rlabel metal2 233 -65 233 -65 0 net=655
rlabel metal2 37 -67 37 -67 0 net=584
rlabel metal2 72 -67 72 -67 0 net=329
rlabel metal2 152 -67 152 -67 0 net=357
rlabel metal2 163 -67 163 -67 0 net=537
rlabel metal2 47 -69 47 -69 0 net=57
rlabel metal2 93 -69 93 -69 0 net=446
rlabel metal2 131 -69 131 -69 0 net=568
rlabel metal2 177 -69 177 -69 0 net=430
rlabel metal2 51 -71 51 -71 0 net=478
rlabel metal2 93 -71 93 -71 0 net=251
rlabel metal2 128 -71 128 -71 0 net=389
rlabel metal2 191 -71 191 -71 0 net=631
rlabel metal2 54 -73 54 -73 0 net=123
rlabel metal2 79 -73 79 -73 0 net=457
rlabel metal2 100 -73 100 -73 0 net=496
rlabel metal2 58 -75 58 -75 0 net=292
rlabel metal2 114 -75 114 -75 0 net=258
rlabel metal2 135 -75 135 -75 0 net=559
rlabel metal2 86 -77 86 -77 0 net=359
rlabel metal2 100 -79 100 -79 0 net=253
rlabel metal2 128 -79 128 -79 0 net=521
rlabel metal2 107 -81 107 -81 0 net=281
rlabel metal2 142 -81 142 -81 0 net=409
rlabel metal2 121 -83 121 -83 0 net=321
rlabel metal2 2 -94 2 -94 0 net=633
rlabel metal2 114 -94 114 -94 0 net=254
rlabel metal2 142 -94 142 -94 0 net=628
rlabel metal2 233 -94 233 -94 0 net=656
rlabel metal2 9 -96 9 -96 0 net=603
rlabel metal2 58 -96 58 -96 0 net=307
rlabel metal2 79 -96 79 -96 0 net=458
rlabel metal2 107 -96 107 -96 0 net=339
rlabel metal2 124 -96 124 -96 0 net=305
rlabel metal2 145 -96 145 -96 0 net=538
rlabel metal2 212 -96 212 -96 0 net=561
rlabel metal2 240 -96 240 -96 0 net=549
rlabel metal2 23 -98 23 -98 0 net=511
rlabel metal2 47 -98 47 -98 0 net=165
rlabel metal2 145 -98 145 -98 0 net=489
rlabel metal2 30 -100 30 -100 0 net=453
rlabel metal2 152 -100 152 -100 0 net=410
rlabel metal2 184 -100 184 -100 0 net=449
rlabel metal2 51 -102 51 -102 0 net=393
rlabel metal2 72 -102 72 -102 0 net=330
rlabel metal2 156 -102 156 -102 0 net=358
rlabel metal2 156 -102 156 -102 0 net=358
rlabel metal2 163 -102 163 -102 0 net=361
rlabel metal2 163 -102 163 -102 0 net=361
rlabel metal2 170 -102 170 -102 0 net=391
rlabel metal2 170 -102 170 -102 0 net=391
rlabel metal2 184 -102 184 -102 0 net=411
rlabel metal2 86 -104 86 -104 0 net=252
rlabel metal2 135 -104 135 -104 0 net=283
rlabel metal2 191 -104 191 -104 0 net=632
rlabel metal2 82 -106 82 -106 0 net=421
rlabel metal2 194 -106 194 -106 0 net=643
rlabel metal2 93 -108 93 -108 0 net=259
rlabel metal2 121 -108 121 -108 0 net=323
rlabel metal2 198 -108 198 -108 0 net=523
rlabel metal2 121 -110 121 -110 0 net=591
rlabel metal2 159 -112 159 -112 0 net=439
rlabel metal2 2 -123 2 -123 0 net=634
rlabel metal2 58 -123 58 -123 0 net=309
rlabel metal2 79 -123 79 -123 0 net=450
rlabel metal2 212 -123 212 -123 0 net=645
rlabel metal2 2 -125 2 -125 0 net=395
rlabel metal2 86 -125 86 -125 0 net=490
rlabel metal2 9 -127 9 -127 0 net=604
rlabel metal2 89 -127 89 -127 0 net=575
rlabel metal2 19 -129 19 -129 0 net=177
rlabel metal2 47 -129 47 -129 0 net=99
rlabel metal2 93 -129 93 -129 0 net=261
rlabel metal2 149 -129 149 -129 0 net=524
rlabel metal2 19 -131 19 -131 0 net=40
rlabel metal2 51 -131 51 -131 0 net=381
rlabel metal2 100 -131 100 -131 0 net=585
rlabel metal2 219 -131 219 -131 0 net=551
rlabel metal2 23 -133 23 -133 0 net=512
rlabel metal2 100 -133 100 -133 0 net=341
rlabel metal2 114 -133 114 -133 0 net=562
rlabel metal2 30 -135 30 -135 0 net=454
rlabel metal2 72 -135 72 -135 0 net=299
rlabel metal2 117 -135 117 -135 0 net=509
rlabel metal2 9 -137 9 -137 0 net=317
rlabel metal2 107 -137 107 -137 0 net=306
rlabel metal2 135 -137 135 -137 0 net=325
rlabel metal2 226 -137 226 -137 0 net=469
rlabel metal2 121 -139 121 -139 0 net=392
rlabel metal2 187 -139 187 -139 0 net=592
rlabel metal2 121 -141 121 -141 0 net=245
rlabel metal2 149 -141 149 -141 0 net=363
rlabel metal2 128 -143 128 -143 0 net=285
rlabel metal2 135 -145 135 -145 0 net=497
rlabel metal2 177 -145 177 -145 0 net=423
rlabel metal2 138 -147 138 -147 0 net=613
rlabel metal2 152 -149 152 -149 0 net=607
rlabel metal2 156 -151 156 -151 0 net=563
rlabel metal2 159 -153 159 -153 0 net=625
rlabel metal2 163 -155 163 -155 0 net=441
rlabel metal2 184 -157 184 -157 0 net=413
rlabel metal2 2 -168 2 -168 0 net=396
rlabel metal2 96 -168 96 -168 0 net=262
rlabel metal2 149 -168 149 -168 0 net=365
rlabel metal2 159 -168 159 -168 0 net=414
rlabel metal2 219 -168 219 -168 0 net=553
rlabel metal2 219 -168 219 -168 0 net=553
rlabel metal2 240 -168 240 -168 0 net=609
rlabel metal2 240 -168 240 -168 0 net=609
rlabel metal2 247 -168 247 -168 0 net=615
rlabel metal2 247 -168 247 -168 0 net=615
rlabel metal2 9 -170 9 -170 0 net=318
rlabel metal2 58 -170 58 -170 0 net=310
rlabel metal2 82 -170 82 -170 0 net=66
rlabel metal2 100 -170 100 -170 0 net=342
rlabel metal2 107 -170 107 -170 0 net=72
rlabel metal2 117 -170 117 -170 0 net=510
rlabel metal2 23 -172 23 -172 0 net=289
rlabel metal2 170 -172 170 -172 0 net=499
rlabel metal2 212 -172 212 -172 0 net=587
rlabel metal2 26 -174 26 -174 0 net=300
rlabel metal2 79 -174 79 -174 0 net=169
rlabel metal2 121 -174 121 -174 0 net=247
rlabel metal2 121 -174 121 -174 0 net=247
rlabel metal2 128 -174 128 -174 0 net=286
rlabel metal2 149 -174 149 -174 0 net=646
rlabel metal2 40 -176 40 -176 0 net=142
rlabel metal2 51 -176 51 -176 0 net=383
rlabel metal2 65 -176 65 -176 0 net=21
rlabel metal2 128 -176 128 -176 0 net=576
rlabel metal2 30 -178 30 -178 0 net=233
rlabel metal2 51 -178 51 -178 0 net=185
rlabel metal2 135 -178 135 -178 0 net=326
rlabel metal2 212 -178 212 -178 0 net=471
rlabel metal2 254 -178 254 -178 0 net=651
rlabel metal2 72 -180 72 -180 0 net=401
rlabel metal2 135 -180 135 -180 0 net=626
rlabel metal2 86 -182 86 -182 0 net=187
rlabel metal2 163 -182 163 -182 0 net=443
rlabel metal2 184 -182 184 -182 0 net=573
rlabel metal2 163 -184 163 -184 0 net=425
rlabel metal2 187 -184 187 -184 0 net=349
rlabel metal2 177 -186 177 -186 0 net=513
rlabel metal2 191 -188 191 -188 0 net=565
rlabel metal2 23 -199 23 -199 0 net=290
rlabel metal2 93 -199 93 -199 0 net=115
rlabel metal2 177 -199 177 -199 0 net=514
rlabel metal2 177 -199 177 -199 0 net=514
rlabel metal2 184 -199 184 -199 0 net=405
rlabel metal2 212 -199 212 -199 0 net=473
rlabel metal2 212 -199 212 -199 0 net=473
rlabel metal2 282 -199 282 -199 0 net=611
rlabel metal2 30 -201 30 -201 0 net=234
rlabel metal2 30 -201 30 -201 0 net=234
rlabel metal2 37 -201 37 -201 0 net=384
rlabel metal2 68 -201 68 -201 0 net=30
rlabel metal2 110 -201 110 -201 0 net=426
rlabel metal2 187 -201 187 -201 0 net=566
rlabel metal2 278 -201 278 -201 0 net=483
rlabel metal2 37 -203 37 -203 0 net=403
rlabel metal2 100 -203 100 -203 0 net=215
rlabel metal2 135 -203 135 -203 0 net=366
rlabel metal2 191 -203 191 -203 0 net=588
rlabel metal2 44 -205 44 -205 0 net=610
rlabel metal2 51 -207 51 -207 0 net=186
rlabel metal2 117 -207 117 -207 0 net=248
rlabel metal2 135 -207 135 -207 0 net=58
rlabel metal2 152 -207 152 -207 0 net=652
rlabel metal2 44 -209 44 -209 0 net=331
rlabel metal2 58 -209 58 -209 0 net=519
rlabel metal2 114 -209 114 -209 0 net=229
rlabel metal2 138 -209 138 -209 0 net=461
rlabel metal2 254 -209 254 -209 0 net=657
rlabel metal2 65 -211 65 -211 0 net=373
rlabel metal2 117 -211 117 -211 0 net=444
rlabel metal2 198 -211 198 -211 0 net=501
rlabel metal2 219 -211 219 -211 0 net=555
rlabel metal2 86 -213 86 -213 0 net=189
rlabel metal2 142 -213 142 -213 0 net=574
rlabel metal2 86 -215 86 -215 0 net=219
rlabel metal2 180 -215 180 -215 0 net=545
rlabel metal2 107 -217 107 -217 0 net=371
rlabel metal2 149 -217 149 -217 0 net=569
rlabel metal2 194 -217 194 -217 0 net=479
rlabel metal2 47 -219 47 -219 0 net=269
rlabel metal2 149 -219 149 -219 0 net=397
rlabel metal2 198 -219 198 -219 0 net=351
rlabel metal2 247 -221 247 -221 0 net=616
rlabel metal2 247 -223 247 -223 0 net=577
rlabel metal2 16 -234 16 -234 0 net=601
rlabel metal2 58 -234 58 -234 0 net=520
rlabel metal2 93 -234 93 -234 0 net=190
rlabel metal2 156 -234 156 -234 0 net=658
rlabel metal2 275 -234 275 -234 0 net=612
rlabel metal2 30 -236 30 -236 0 net=467
rlabel metal2 128 -236 128 -236 0 net=235
rlabel metal2 159 -236 159 -236 0 net=462
rlabel metal2 240 -236 240 -236 0 net=556
rlabel metal2 282 -236 282 -236 0 net=485
rlabel metal2 282 -236 282 -236 0 net=485
rlabel metal2 37 -238 37 -238 0 net=404
rlabel metal2 173 -238 173 -238 0 net=406
rlabel metal2 212 -238 212 -238 0 net=475
rlabel metal2 212 -238 212 -238 0 net=475
rlabel metal2 219 -238 219 -238 0 net=481
rlabel metal2 240 -238 240 -238 0 net=557
rlabel metal2 37 -240 37 -240 0 net=379
rlabel metal2 93 -240 93 -240 0 net=191
rlabel metal2 184 -240 184 -240 0 net=353
rlabel metal2 205 -240 205 -240 0 net=503
rlabel metal2 226 -240 226 -240 0 net=547
rlabel metal2 226 -240 226 -240 0 net=547
rlabel metal2 247 -240 247 -240 0 net=579
rlabel metal2 58 -242 58 -242 0 net=217
rlabel metal2 103 -242 103 -242 0 net=372
rlabel metal2 163 -242 163 -242 0 net=399
rlabel metal2 65 -244 65 -244 0 net=375
rlabel metal2 107 -244 107 -244 0 net=271
rlabel metal2 177 -244 177 -244 0 net=527
rlabel metal2 51 -246 51 -246 0 net=333
rlabel metal2 72 -246 72 -246 0 net=221
rlabel metal2 107 -246 107 -246 0 net=539
rlabel metal2 180 -246 180 -246 0 net=589
rlabel metal2 86 -248 86 -248 0 net=311
rlabel metal2 121 -248 121 -248 0 net=231
rlabel metal2 121 -250 121 -250 0 net=367
rlabel metal2 170 -252 170 -252 0 net=570
rlabel metal2 156 -254 156 -254 0 net=263
rlabel metal2 26 -265 26 -265 0 net=122
rlabel metal2 47 -265 47 -265 0 net=334
rlabel metal2 86 -265 86 -265 0 net=312
rlabel metal2 114 -265 114 -265 0 net=400
rlabel metal2 208 -265 208 -265 0 net=548
rlabel metal2 254 -265 254 -265 0 net=581
rlabel metal2 254 -265 254 -265 0 net=581
rlabel metal2 282 -265 282 -265 0 net=486
rlabel metal2 16 -267 16 -267 0 net=602
rlabel metal2 89 -267 89 -267 0 net=236
rlabel metal2 135 -267 135 -267 0 net=354
rlabel metal2 191 -267 191 -267 0 net=476
rlabel metal2 30 -269 30 -269 0 net=468
rlabel metal2 103 -269 103 -269 0 net=232
rlabel metal2 170 -269 170 -269 0 net=505
rlabel metal2 180 -269 180 -269 0 net=504
rlabel metal2 37 -271 37 -271 0 net=380
rlabel metal2 121 -271 121 -271 0 net=369
rlabel metal2 121 -271 121 -271 0 net=369
rlabel metal2 128 -271 128 -271 0 net=265
rlabel metal2 173 -271 173 -271 0 net=590
rlabel metal2 51 -273 51 -273 0 net=53
rlabel metal2 194 -273 194 -273 0 net=558
rlabel metal2 54 -275 54 -275 0 net=222
rlabel metal2 93 -275 93 -275 0 net=193
rlabel metal2 135 -275 135 -275 0 net=273
rlabel metal2 198 -275 198 -275 0 net=529
rlabel metal2 198 -275 198 -275 0 net=529
rlabel metal2 205 -275 205 -275 0 net=482
rlabel metal2 240 -275 240 -275 0 net=435
rlabel metal2 58 -277 58 -277 0 net=218
rlabel metal2 149 -277 149 -277 0 net=541
rlabel metal2 65 -279 65 -279 0 net=313
rlabel metal2 100 -279 100 -279 0 net=619
rlabel metal2 149 -279 149 -279 0 net=415
rlabel metal2 72 -281 72 -281 0 net=377
rlabel metal2 51 -292 51 -292 0 net=593
rlabel metal2 117 -292 117 -292 0 net=370
rlabel metal2 128 -292 128 -292 0 net=267
rlabel metal2 128 -292 128 -292 0 net=267
rlabel metal2 138 -292 138 -292 0 net=140
rlabel metal2 219 -292 219 -292 0 net=647
rlabel metal2 240 -292 240 -292 0 net=437
rlabel metal2 240 -292 240 -292 0 net=437
rlabel metal2 250 -292 250 -292 0 net=582
rlabel metal2 65 -294 65 -294 0 net=314
rlabel metal2 107 -294 107 -294 0 net=195
rlabel metal2 142 -294 142 -294 0 net=621
rlabel metal2 184 -294 184 -294 0 net=91
rlabel metal2 65 -296 65 -296 0 net=297
rlabel metal2 117 -296 117 -296 0 net=301
rlabel metal2 156 -296 156 -296 0 net=542
rlabel metal2 170 -296 170 -296 0 net=507
rlabel metal2 170 -296 170 -296 0 net=507
rlabel metal2 191 -296 191 -296 0 net=530
rlabel metal2 72 -298 72 -298 0 net=378
rlabel metal2 149 -298 149 -298 0 net=417
rlabel metal2 75 -300 75 -300 0 net=10
rlabel metal2 89 -300 89 -300 0 net=11
rlabel metal2 110 -300 110 -300 0 net=343
rlabel metal2 82 -302 82 -302 0 net=90
rlabel metal2 96 -302 96 -302 0 net=319
rlabel metal2 89 -304 89 -304 0 net=147
rlabel metal2 103 -304 103 -304 0 net=274
rlabel metal2 44 -315 44 -315 0 net=387
rlabel metal2 96 -315 96 -315 0 net=12
rlabel metal2 159 -315 159 -315 0 net=508
rlabel metal2 177 -315 177 -315 0 net=623
rlabel metal2 219 -315 219 -315 0 net=649
rlabel metal2 219 -315 219 -315 0 net=649
rlabel metal2 226 -315 226 -315 0 net=114
rlabel metal2 236 -315 236 -315 0 net=438
rlabel metal2 51 -317 51 -317 0 net=594
rlabel metal2 107 -317 107 -317 0 net=268
rlabel metal2 138 -317 138 -317 0 net=327
rlabel metal2 51 -319 51 -319 0 net=237
rlabel metal2 107 -319 107 -319 0 net=197
rlabel metal2 128 -319 128 -319 0 net=320
rlabel metal2 61 -321 61 -321 0 net=298
rlabel metal2 72 -321 72 -321 0 net=136
rlabel metal2 138 -321 138 -321 0 net=431
rlabel metal2 61 -323 61 -323 0 net=156
rlabel metal2 79 -323 79 -323 0 net=617
rlabel metal2 65 -325 65 -325 0 net=223
rlabel metal2 93 -325 93 -325 0 net=128
rlabel metal2 114 -325 114 -325 0 net=418
rlabel metal2 37 -327 37 -327 0 net=605
rlabel metal2 117 -327 117 -327 0 net=207
rlabel metal2 135 -327 135 -327 0 net=315
rlabel metal2 72 -329 72 -329 0 net=303
rlabel metal2 149 -329 149 -329 0 net=345
rlabel metal2 131 -331 131 -331 0 net=275
rlabel metal2 142 -333 142 -333 0 net=459
rlabel metal2 37 -344 37 -344 0 net=606
rlabel metal2 100 -344 100 -344 0 net=316
rlabel metal2 194 -344 194 -344 0 net=618
rlabel metal2 215 -344 215 -344 0 net=650
rlabel metal2 44 -346 44 -346 0 net=388
rlabel metal2 121 -346 121 -346 0 net=209
rlabel metal2 121 -346 121 -346 0 net=209
rlabel metal2 135 -346 135 -346 0 net=487
rlabel metal2 145 -346 145 -346 0 net=624
rlabel metal2 58 -348 58 -348 0 net=22
rlabel metal2 110 -348 110 -348 0 net=135
rlabel metal2 51 -350 51 -350 0 net=239
rlabel metal2 65 -350 65 -350 0 net=225
rlabel metal2 65 -350 65 -350 0 net=225
rlabel metal2 72 -350 72 -350 0 net=304
rlabel metal2 149 -350 149 -350 0 net=277
rlabel metal2 177 -350 177 -350 0 net=347
rlabel metal2 72 -352 72 -352 0 net=637
rlabel metal2 114 -352 114 -352 0 net=328
rlabel metal2 177 -352 177 -352 0 net=433
rlabel metal2 79 -354 79 -354 0 net=199
rlabel metal2 149 -354 149 -354 0 net=427
rlabel metal2 170 -354 170 -354 0 net=460
rlabel metal2 86 -356 86 -356 0 net=181
rlabel metal2 96 -358 96 -358 0 net=51
rlabel metal2 131 -358 131 -358 0 net=653
rlabel metal2 103 -360 103 -360 0 net=227
rlabel metal2 58 -371 58 -371 0 net=240
rlabel metal2 135 -371 135 -371 0 net=488
rlabel metal2 145 -371 145 -371 0 net=654
rlabel metal2 65 -373 65 -373 0 net=226
rlabel metal2 138 -373 138 -373 0 net=428
rlabel metal2 156 -373 156 -373 0 net=348
rlabel metal2 72 -375 72 -375 0 net=638
rlabel metal2 103 -375 103 -375 0 net=228
rlabel metal2 142 -375 142 -375 0 net=279
rlabel metal2 170 -375 170 -375 0 net=434
rlabel metal2 72 -377 72 -377 0 net=493
rlabel metal2 100 -377 100 -377 0 net=463
rlabel metal2 114 -377 114 -377 0 net=451
rlabel metal2 79 -379 79 -379 0 net=200
rlabel metal2 121 -379 121 -379 0 net=211
rlabel metal2 149 -379 149 -379 0 net=355
rlabel metal2 79 -381 79 -381 0 net=213
rlabel metal2 121 -381 121 -381 0 net=525
rlabel metal2 86 -383 86 -383 0 net=183
rlabel metal2 86 -383 86 -383 0 net=183
rlabel metal2 79 -394 79 -394 0 net=214
rlabel metal2 114 -394 114 -394 0 net=212
rlabel metal2 131 -394 131 -394 0 net=356
rlabel metal2 170 -394 170 -394 0 net=86
rlabel metal2 72 -396 72 -396 0 net=494
rlabel metal2 145 -396 145 -396 0 net=452
rlabel metal2 86 -398 86 -398 0 net=184
rlabel metal2 79 -400 79 -400 0 net=241
rlabel metal2 93 -400 93 -400 0 net=465
rlabel metal2 121 -400 121 -400 0 net=280
rlabel metal2 117 -402 117 -402 0 net=641
rlabel metal2 142 -402 142 -402 0 net=526
rlabel metal2 107 -404 107 -404 0 net=203
rlabel metal2 156 -404 156 -404 0 net=335
rlabel metal2 93 -415 93 -415 0 net=466
rlabel metal2 117 -415 117 -415 0 net=642
rlabel metal2 156 -415 156 -415 0 net=337
rlabel metal2 86 -417 86 -417 0 net=243
rlabel metal2 107 -417 107 -417 0 net=205
rlabel metal2 89 -428 89 -428 0 net=244
rlabel metal2 117 -428 117 -428 0 net=206
rlabel metal2 163 -428 163 -428 0 net=338
<< end >>
