magic
tech scmos
timestamp 1555071775 
<< pdiffusion >>
rect 1 -10 7 -4
rect 8 -10 14 -4
rect 15 -10 21 -4
rect 22 -10 28 -4
rect 29 -10 35 -4
rect 36 -10 42 -4
rect 43 -10 49 -4
rect 50 -10 56 -4
rect 57 -10 63 -4
rect 64 -10 70 -4
rect 106 -10 112 -4
rect 176 -10 179 -4
rect 183 -10 189 -4
rect 190 -10 196 -4
rect 197 -10 200 -4
rect 204 -10 210 -4
rect 211 -10 217 -4
rect 218 -10 224 -4
rect 225 -10 231 -4
rect 232 -10 235 -4
rect 239 -10 245 -4
rect 246 -10 249 -4
rect 253 -10 256 -4
rect 274 -10 280 -4
rect 281 -10 284 -4
rect 288 -10 291 -4
rect 295 -10 301 -4
rect 302 -10 308 -4
rect 1 -29 7 -23
rect 8 -29 14 -23
rect 15 -29 21 -23
rect 22 -29 28 -23
rect 29 -29 35 -23
rect 36 -29 42 -23
rect 43 -29 49 -23
rect 50 -29 56 -23
rect 141 -29 144 -23
rect 148 -29 151 -23
rect 155 -29 161 -23
rect 162 -29 168 -23
rect 169 -29 175 -23
rect 176 -29 182 -23
rect 183 -29 186 -23
rect 190 -29 196 -23
rect 197 -29 200 -23
rect 204 -29 210 -23
rect 211 -29 217 -23
rect 218 -29 221 -23
rect 239 -29 242 -23
rect 246 -29 252 -23
rect 253 -29 259 -23
rect 260 -29 266 -23
rect 267 -29 270 -23
rect 274 -29 277 -23
rect 281 -29 287 -23
rect 288 -29 294 -23
rect 295 -29 298 -23
rect 302 -29 308 -23
rect 309 -29 312 -23
rect 316 -29 322 -23
rect 1 -42 7 -36
rect 8 -42 14 -36
rect 15 -42 21 -36
rect 22 -42 28 -36
rect 29 -42 35 -36
rect 36 -42 42 -36
rect 43 -42 49 -36
rect 50 -42 56 -36
rect 78 -42 84 -36
rect 134 -42 137 -36
rect 141 -42 147 -36
rect 148 -42 154 -36
rect 155 -42 158 -36
rect 169 -42 175 -36
rect 183 -42 186 -36
rect 190 -42 196 -36
rect 211 -42 217 -36
rect 218 -42 224 -36
rect 225 -42 231 -36
rect 232 -42 235 -36
rect 239 -42 245 -36
rect 246 -42 252 -36
rect 253 -42 256 -36
rect 260 -42 263 -36
rect 267 -42 273 -36
rect 274 -42 277 -36
rect 281 -42 284 -36
rect 288 -42 294 -36
rect 295 -42 298 -36
rect 302 -42 308 -36
rect 309 -42 315 -36
rect 316 -42 319 -36
rect 323 -42 326 -36
rect 330 -42 336 -36
rect 477 -42 483 -36
rect 484 -42 487 -36
rect 575 -42 581 -36
rect 582 -42 585 -36
rect 1 -65 7 -59
rect 8 -65 14 -59
rect 15 -65 21 -59
rect 22 -65 28 -59
rect 29 -65 35 -59
rect 36 -65 42 -59
rect 43 -65 49 -59
rect 50 -65 56 -59
rect 78 -65 84 -59
rect 141 -65 147 -59
rect 148 -65 151 -59
rect 155 -65 158 -59
rect 169 -65 172 -59
rect 176 -65 182 -59
rect 183 -65 189 -59
rect 190 -65 196 -59
rect 197 -65 203 -59
rect 204 -65 207 -59
rect 211 -65 217 -59
rect 218 -65 221 -59
rect 225 -65 228 -59
rect 232 -65 238 -59
rect 239 -65 245 -59
rect 246 -65 252 -59
rect 253 -65 256 -59
rect 260 -65 263 -59
rect 267 -65 270 -59
rect 274 -65 277 -59
rect 281 -65 287 -59
rect 288 -65 291 -59
rect 295 -65 298 -59
rect 302 -65 308 -59
rect 309 -65 315 -59
rect 316 -65 322 -59
rect 323 -65 326 -59
rect 337 -65 343 -59
rect 344 -65 347 -59
rect 351 -65 354 -59
rect 358 -65 364 -59
rect 463 -65 469 -59
rect 470 -65 473 -59
rect 477 -65 480 -59
rect 575 -65 578 -59
rect 1 -88 7 -82
rect 8 -88 14 -82
rect 15 -88 21 -82
rect 22 -88 28 -82
rect 29 -88 35 -82
rect 36 -88 42 -82
rect 43 -88 49 -82
rect 120 -88 126 -82
rect 134 -88 140 -82
rect 141 -88 144 -82
rect 148 -88 151 -82
rect 155 -88 161 -82
rect 162 -88 168 -82
rect 169 -88 172 -82
rect 176 -88 179 -82
rect 183 -88 189 -82
rect 190 -88 196 -82
rect 197 -88 203 -82
rect 204 -88 210 -82
rect 211 -88 214 -82
rect 218 -88 221 -82
rect 225 -88 228 -82
rect 232 -88 235 -82
rect 239 -88 245 -82
rect 246 -88 249 -82
rect 253 -88 256 -82
rect 260 -88 263 -82
rect 267 -88 273 -82
rect 274 -88 280 -82
rect 281 -88 284 -82
rect 288 -88 294 -82
rect 295 -88 298 -82
rect 302 -88 308 -82
rect 309 -88 315 -82
rect 316 -88 319 -82
rect 323 -88 329 -82
rect 337 -88 340 -82
rect 344 -88 350 -82
rect 351 -88 354 -82
rect 470 -88 476 -82
rect 477 -88 480 -82
rect 484 -88 487 -82
rect 575 -88 578 -82
rect 1 -119 7 -113
rect 8 -119 14 -113
rect 15 -119 21 -113
rect 22 -119 28 -113
rect 29 -119 35 -113
rect 36 -119 42 -113
rect 106 -119 109 -113
rect 120 -119 126 -113
rect 127 -119 133 -113
rect 134 -119 137 -113
rect 141 -119 147 -113
rect 148 -119 154 -113
rect 155 -119 158 -113
rect 162 -119 165 -113
rect 169 -119 175 -113
rect 176 -119 182 -113
rect 183 -119 186 -113
rect 190 -119 193 -113
rect 197 -119 200 -113
rect 204 -119 210 -113
rect 211 -119 217 -113
rect 218 -119 224 -113
rect 225 -119 228 -113
rect 232 -119 235 -113
rect 239 -119 245 -113
rect 246 -119 252 -113
rect 253 -119 259 -113
rect 260 -119 263 -113
rect 267 -119 270 -113
rect 274 -119 280 -113
rect 281 -119 284 -113
rect 288 -119 291 -113
rect 295 -119 298 -113
rect 302 -119 305 -113
rect 309 -119 312 -113
rect 316 -119 322 -113
rect 323 -119 326 -113
rect 330 -119 333 -113
rect 337 -119 343 -113
rect 344 -119 347 -113
rect 351 -119 354 -113
rect 358 -119 361 -113
rect 365 -119 368 -113
rect 372 -119 375 -113
rect 379 -119 382 -113
rect 393 -119 399 -113
rect 421 -119 424 -113
rect 477 -119 483 -113
rect 484 -119 487 -113
rect 491 -119 494 -113
rect 575 -119 581 -113
rect 582 -119 585 -113
rect 589 -119 592 -113
rect 1 -158 7 -152
rect 8 -158 14 -152
rect 15 -158 21 -152
rect 22 -158 28 -152
rect 29 -158 35 -152
rect 64 -158 67 -152
rect 71 -158 74 -152
rect 78 -158 84 -152
rect 85 -158 88 -152
rect 92 -158 95 -152
rect 99 -158 105 -152
rect 106 -158 109 -152
rect 113 -158 119 -152
rect 120 -158 126 -152
rect 127 -158 133 -152
rect 134 -158 137 -152
rect 141 -158 147 -152
rect 148 -158 151 -152
rect 155 -158 158 -152
rect 162 -158 168 -152
rect 169 -158 172 -152
rect 176 -158 179 -152
rect 183 -158 186 -152
rect 190 -158 193 -152
rect 197 -158 200 -152
rect 204 -158 210 -152
rect 211 -158 217 -152
rect 218 -158 224 -152
rect 225 -158 231 -152
rect 232 -158 238 -152
rect 239 -158 245 -152
rect 246 -158 249 -152
rect 253 -158 256 -152
rect 260 -158 266 -152
rect 267 -158 270 -152
rect 274 -158 277 -152
rect 281 -158 287 -152
rect 288 -158 291 -152
rect 295 -158 301 -152
rect 302 -158 305 -152
rect 309 -158 312 -152
rect 316 -158 319 -152
rect 323 -158 326 -152
rect 330 -158 336 -152
rect 337 -158 340 -152
rect 344 -158 347 -152
rect 351 -158 357 -152
rect 358 -158 361 -152
rect 365 -158 368 -152
rect 372 -158 375 -152
rect 379 -158 382 -152
rect 386 -158 392 -152
rect 393 -158 396 -152
rect 400 -158 403 -152
rect 407 -158 413 -152
rect 414 -158 417 -152
rect 421 -158 424 -152
rect 428 -158 431 -152
rect 435 -158 438 -152
rect 442 -158 445 -152
rect 498 -158 501 -152
rect 589 -158 592 -152
rect 1 -207 7 -201
rect 8 -207 14 -201
rect 15 -207 21 -201
rect 22 -207 28 -201
rect 29 -207 35 -201
rect 78 -207 81 -201
rect 85 -207 88 -201
rect 92 -207 98 -201
rect 99 -207 102 -201
rect 106 -207 109 -201
rect 113 -207 116 -201
rect 120 -207 126 -201
rect 127 -207 130 -201
rect 134 -207 137 -201
rect 141 -207 147 -201
rect 148 -207 151 -201
rect 155 -207 161 -201
rect 162 -207 168 -201
rect 169 -207 175 -201
rect 176 -207 182 -201
rect 183 -207 189 -201
rect 190 -207 196 -201
rect 197 -207 203 -201
rect 204 -207 207 -201
rect 211 -207 217 -201
rect 218 -207 224 -201
rect 225 -207 231 -201
rect 232 -207 238 -201
rect 239 -207 245 -201
rect 246 -207 249 -201
rect 253 -207 256 -201
rect 260 -207 263 -201
rect 267 -207 270 -201
rect 274 -207 280 -201
rect 281 -207 284 -201
rect 288 -207 294 -201
rect 295 -207 301 -201
rect 302 -207 305 -201
rect 309 -207 312 -201
rect 316 -207 322 -201
rect 323 -207 326 -201
rect 330 -207 333 -201
rect 337 -207 340 -201
rect 344 -207 347 -201
rect 351 -207 354 -201
rect 358 -207 361 -201
rect 365 -207 368 -201
rect 372 -207 375 -201
rect 379 -207 382 -201
rect 386 -207 389 -201
rect 393 -207 396 -201
rect 400 -207 403 -201
rect 407 -207 410 -201
rect 414 -207 417 -201
rect 421 -207 427 -201
rect 428 -207 431 -201
rect 435 -207 438 -201
rect 442 -207 445 -201
rect 449 -207 455 -201
rect 456 -207 462 -201
rect 463 -207 466 -201
rect 505 -207 508 -201
rect 589 -207 592 -201
rect 1 -248 7 -242
rect 8 -248 14 -242
rect 15 -248 21 -242
rect 22 -248 28 -242
rect 113 -248 116 -242
rect 120 -248 126 -242
rect 127 -248 130 -242
rect 134 -248 137 -242
rect 141 -248 144 -242
rect 148 -248 151 -242
rect 155 -248 161 -242
rect 162 -248 165 -242
rect 169 -248 175 -242
rect 176 -248 179 -242
rect 183 -248 186 -242
rect 190 -248 193 -242
rect 197 -248 200 -242
rect 204 -248 210 -242
rect 211 -248 217 -242
rect 218 -248 224 -242
rect 225 -248 231 -242
rect 232 -248 238 -242
rect 239 -248 245 -242
rect 246 -248 249 -242
rect 253 -248 256 -242
rect 260 -248 266 -242
rect 267 -248 270 -242
rect 274 -248 280 -242
rect 281 -248 284 -242
rect 288 -248 294 -242
rect 295 -248 301 -242
rect 302 -248 305 -242
rect 309 -248 312 -242
rect 316 -248 322 -242
rect 323 -248 326 -242
rect 330 -248 333 -242
rect 337 -248 340 -242
rect 344 -248 350 -242
rect 351 -248 354 -242
rect 358 -248 361 -242
rect 365 -248 371 -242
rect 372 -248 375 -242
rect 379 -248 385 -242
rect 386 -248 389 -242
rect 393 -248 396 -242
rect 400 -248 403 -242
rect 407 -248 410 -242
rect 414 -248 417 -242
rect 421 -248 424 -242
rect 428 -248 431 -242
rect 435 -248 438 -242
rect 442 -248 445 -242
rect 449 -248 452 -242
rect 456 -248 462 -242
rect 463 -248 469 -242
rect 505 -248 511 -242
rect 561 -248 567 -242
rect 568 -248 574 -242
rect 589 -248 592 -242
rect 596 -248 602 -242
rect 645 -248 651 -242
rect 1 -289 7 -283
rect 8 -289 14 -283
rect 15 -289 21 -283
rect 64 -289 70 -283
rect 71 -289 77 -283
rect 78 -289 81 -283
rect 85 -289 88 -283
rect 92 -289 95 -283
rect 99 -289 105 -283
rect 106 -289 109 -283
rect 113 -289 119 -283
rect 120 -289 126 -283
rect 127 -289 130 -283
rect 134 -289 137 -283
rect 141 -289 144 -283
rect 148 -289 151 -283
rect 155 -289 158 -283
rect 162 -289 165 -283
rect 169 -289 175 -283
rect 176 -289 179 -283
rect 183 -289 189 -283
rect 190 -289 196 -283
rect 197 -289 203 -283
rect 204 -289 210 -283
rect 211 -289 217 -283
rect 218 -289 221 -283
rect 225 -289 228 -283
rect 232 -289 238 -283
rect 239 -289 245 -283
rect 246 -289 249 -283
rect 253 -289 259 -283
rect 260 -289 263 -283
rect 267 -289 270 -283
rect 274 -289 277 -283
rect 281 -289 287 -283
rect 288 -289 294 -283
rect 295 -289 301 -283
rect 302 -289 308 -283
rect 309 -289 315 -283
rect 316 -289 322 -283
rect 323 -289 329 -283
rect 330 -289 333 -283
rect 337 -289 343 -283
rect 344 -289 347 -283
rect 351 -289 354 -283
rect 358 -289 361 -283
rect 365 -289 368 -283
rect 372 -289 375 -283
rect 379 -289 385 -283
rect 386 -289 389 -283
rect 393 -289 399 -283
rect 400 -289 403 -283
rect 407 -289 410 -283
rect 414 -289 417 -283
rect 421 -289 424 -283
rect 428 -289 431 -283
rect 435 -289 438 -283
rect 442 -289 445 -283
rect 449 -289 452 -283
rect 456 -289 459 -283
rect 463 -289 466 -283
rect 470 -289 473 -283
rect 477 -289 480 -283
rect 484 -289 487 -283
rect 491 -289 494 -283
rect 498 -289 504 -283
rect 505 -289 508 -283
rect 519 -289 522 -283
rect 526 -289 529 -283
rect 561 -289 564 -283
rect 610 -289 613 -283
rect 645 -289 648 -283
rect 1 -338 7 -332
rect 8 -338 14 -332
rect 71 -338 77 -332
rect 78 -338 81 -332
rect 85 -338 88 -332
rect 92 -338 95 -332
rect 99 -338 102 -332
rect 106 -338 109 -332
rect 113 -338 116 -332
rect 120 -338 123 -332
rect 127 -338 133 -332
rect 134 -338 137 -332
rect 141 -338 144 -332
rect 148 -338 154 -332
rect 155 -338 161 -332
rect 162 -338 168 -332
rect 169 -338 172 -332
rect 176 -338 179 -332
rect 183 -338 189 -332
rect 190 -338 193 -332
rect 197 -338 200 -332
rect 204 -338 207 -332
rect 211 -338 214 -332
rect 218 -338 224 -332
rect 225 -338 231 -332
rect 232 -338 238 -332
rect 239 -338 242 -332
rect 246 -338 249 -332
rect 253 -338 256 -332
rect 260 -338 266 -332
rect 267 -338 273 -332
rect 274 -338 277 -332
rect 281 -338 287 -332
rect 288 -338 291 -332
rect 295 -338 298 -332
rect 302 -338 305 -332
rect 309 -338 315 -332
rect 316 -338 319 -332
rect 323 -338 329 -332
rect 330 -338 333 -332
rect 337 -338 343 -332
rect 344 -338 350 -332
rect 351 -338 354 -332
rect 358 -338 364 -332
rect 365 -338 371 -332
rect 372 -338 375 -332
rect 379 -338 382 -332
rect 386 -338 392 -332
rect 393 -338 396 -332
rect 400 -338 403 -332
rect 407 -338 413 -332
rect 414 -338 417 -332
rect 421 -338 427 -332
rect 428 -338 431 -332
rect 435 -338 438 -332
rect 442 -338 445 -332
rect 449 -338 452 -332
rect 456 -338 459 -332
rect 463 -338 466 -332
rect 470 -338 473 -332
rect 477 -338 480 -332
rect 484 -338 487 -332
rect 491 -338 494 -332
rect 498 -338 501 -332
rect 505 -338 508 -332
rect 512 -338 518 -332
rect 519 -338 522 -332
rect 526 -338 529 -332
rect 533 -338 536 -332
rect 540 -338 546 -332
rect 547 -338 550 -332
rect 554 -338 560 -332
rect 561 -338 564 -332
rect 603 -338 606 -332
rect 645 -338 651 -332
rect 652 -338 655 -332
rect 659 -338 662 -332
rect 673 -338 676 -332
rect 680 -338 686 -332
rect 1 -389 7 -383
rect 29 -389 35 -383
rect 43 -389 46 -383
rect 50 -389 53 -383
rect 57 -389 60 -383
rect 64 -389 70 -383
rect 71 -389 74 -383
rect 78 -389 81 -383
rect 85 -389 88 -383
rect 92 -389 95 -383
rect 99 -389 102 -383
rect 106 -389 112 -383
rect 113 -389 116 -383
rect 120 -389 123 -383
rect 127 -389 130 -383
rect 134 -389 140 -383
rect 141 -389 144 -383
rect 148 -389 154 -383
rect 155 -389 161 -383
rect 162 -389 168 -383
rect 169 -389 172 -383
rect 176 -389 179 -383
rect 183 -389 186 -383
rect 190 -389 193 -383
rect 197 -389 200 -383
rect 204 -389 207 -383
rect 211 -389 217 -383
rect 218 -389 224 -383
rect 225 -389 231 -383
rect 232 -389 238 -383
rect 239 -389 245 -383
rect 246 -389 249 -383
rect 253 -389 256 -383
rect 260 -389 263 -383
rect 267 -389 270 -383
rect 274 -389 280 -383
rect 281 -389 284 -383
rect 288 -389 294 -383
rect 295 -389 298 -383
rect 302 -389 305 -383
rect 309 -389 312 -383
rect 316 -389 319 -383
rect 323 -389 329 -383
rect 330 -389 336 -383
rect 337 -389 343 -383
rect 344 -389 347 -383
rect 351 -389 357 -383
rect 358 -389 364 -383
rect 365 -389 368 -383
rect 372 -389 375 -383
rect 379 -389 382 -383
rect 386 -389 392 -383
rect 393 -389 396 -383
rect 400 -389 403 -383
rect 407 -389 410 -383
rect 414 -389 417 -383
rect 421 -389 427 -383
rect 428 -389 431 -383
rect 435 -389 438 -383
rect 442 -389 445 -383
rect 449 -389 455 -383
rect 456 -389 462 -383
rect 463 -389 466 -383
rect 470 -389 473 -383
rect 477 -389 480 -383
rect 484 -389 487 -383
rect 491 -389 494 -383
rect 498 -389 501 -383
rect 505 -389 508 -383
rect 512 -389 515 -383
rect 519 -389 525 -383
rect 526 -389 529 -383
rect 533 -389 536 -383
rect 540 -389 543 -383
rect 547 -389 550 -383
rect 554 -389 557 -383
rect 561 -389 567 -383
rect 568 -389 571 -383
rect 575 -389 578 -383
rect 582 -389 585 -383
rect 589 -389 592 -383
rect 596 -389 599 -383
rect 603 -389 606 -383
rect 610 -389 613 -383
rect 617 -389 620 -383
rect 624 -389 627 -383
rect 631 -389 634 -383
rect 638 -389 644 -383
rect 645 -389 648 -383
rect 652 -389 655 -383
rect 659 -389 665 -383
rect 666 -389 669 -383
rect 673 -389 679 -383
rect 680 -389 683 -383
rect 687 -389 690 -383
rect 1 -446 4 -440
rect 8 -446 14 -440
rect 15 -446 18 -440
rect 22 -446 25 -440
rect 29 -446 35 -440
rect 36 -446 39 -440
rect 43 -446 46 -440
rect 50 -446 53 -440
rect 57 -446 60 -440
rect 64 -446 67 -440
rect 71 -446 74 -440
rect 78 -446 81 -440
rect 85 -446 91 -440
rect 92 -446 95 -440
rect 99 -446 102 -440
rect 106 -446 109 -440
rect 113 -446 119 -440
rect 120 -446 123 -440
rect 127 -446 130 -440
rect 134 -446 140 -440
rect 141 -446 147 -440
rect 148 -446 151 -440
rect 155 -446 161 -440
rect 162 -446 165 -440
rect 169 -446 172 -440
rect 176 -446 182 -440
rect 183 -446 189 -440
rect 190 -446 193 -440
rect 197 -446 203 -440
rect 204 -446 207 -440
rect 211 -446 217 -440
rect 218 -446 221 -440
rect 225 -446 228 -440
rect 232 -446 238 -440
rect 239 -446 245 -440
rect 246 -446 249 -440
rect 253 -446 256 -440
rect 260 -446 263 -440
rect 267 -446 270 -440
rect 274 -446 277 -440
rect 281 -446 287 -440
rect 288 -446 294 -440
rect 295 -446 298 -440
rect 302 -446 308 -440
rect 309 -446 312 -440
rect 316 -446 319 -440
rect 323 -446 329 -440
rect 330 -446 333 -440
rect 337 -446 343 -440
rect 344 -446 347 -440
rect 351 -446 354 -440
rect 358 -446 361 -440
rect 365 -446 371 -440
rect 372 -446 378 -440
rect 379 -446 382 -440
rect 386 -446 389 -440
rect 393 -446 399 -440
rect 400 -446 406 -440
rect 407 -446 413 -440
rect 414 -446 417 -440
rect 421 -446 424 -440
rect 428 -446 431 -440
rect 435 -446 441 -440
rect 442 -446 445 -440
rect 449 -446 452 -440
rect 456 -446 459 -440
rect 463 -446 469 -440
rect 470 -446 473 -440
rect 477 -446 480 -440
rect 484 -446 487 -440
rect 491 -446 494 -440
rect 498 -446 501 -440
rect 505 -446 511 -440
rect 512 -446 515 -440
rect 519 -446 522 -440
rect 526 -446 529 -440
rect 533 -446 536 -440
rect 540 -446 543 -440
rect 547 -446 550 -440
rect 554 -446 560 -440
rect 561 -446 564 -440
rect 568 -446 571 -440
rect 575 -446 578 -440
rect 582 -446 585 -440
rect 589 -446 592 -440
rect 596 -446 599 -440
rect 603 -446 606 -440
rect 610 -446 613 -440
rect 617 -446 620 -440
rect 624 -446 630 -440
rect 631 -446 637 -440
rect 638 -446 641 -440
rect 645 -446 651 -440
rect 652 -446 655 -440
rect 659 -446 665 -440
rect 666 -446 669 -440
rect 8 -503 11 -497
rect 15 -503 18 -497
rect 22 -503 25 -497
rect 29 -503 32 -497
rect 36 -503 39 -497
rect 43 -503 46 -497
rect 50 -503 53 -497
rect 57 -503 63 -497
rect 64 -503 70 -497
rect 71 -503 74 -497
rect 78 -503 81 -497
rect 85 -503 88 -497
rect 92 -503 98 -497
rect 99 -503 102 -497
rect 106 -503 112 -497
rect 113 -503 119 -497
rect 120 -503 123 -497
rect 127 -503 133 -497
rect 134 -503 140 -497
rect 141 -503 144 -497
rect 148 -503 154 -497
rect 155 -503 161 -497
rect 162 -503 168 -497
rect 169 -503 172 -497
rect 176 -503 179 -497
rect 183 -503 186 -497
rect 190 -503 193 -497
rect 197 -503 203 -497
rect 204 -503 210 -497
rect 211 -503 217 -497
rect 218 -503 221 -497
rect 225 -503 228 -497
rect 232 -503 235 -497
rect 239 -503 245 -497
rect 246 -503 249 -497
rect 253 -503 256 -497
rect 260 -503 266 -497
rect 267 -503 273 -497
rect 274 -503 277 -497
rect 281 -503 284 -497
rect 288 -503 291 -497
rect 295 -503 298 -497
rect 302 -503 305 -497
rect 309 -503 312 -497
rect 316 -503 319 -497
rect 323 -503 326 -497
rect 330 -503 336 -497
rect 337 -503 340 -497
rect 344 -503 347 -497
rect 351 -503 357 -497
rect 358 -503 361 -497
rect 365 -503 371 -497
rect 372 -503 375 -497
rect 379 -503 385 -497
rect 386 -503 392 -497
rect 393 -503 399 -497
rect 400 -503 403 -497
rect 407 -503 410 -497
rect 414 -503 420 -497
rect 421 -503 424 -497
rect 428 -503 431 -497
rect 435 -503 441 -497
rect 442 -503 445 -497
rect 449 -503 452 -497
rect 456 -503 459 -497
rect 463 -503 466 -497
rect 470 -503 473 -497
rect 477 -503 483 -497
rect 484 -503 487 -497
rect 491 -503 494 -497
rect 498 -503 501 -497
rect 505 -503 511 -497
rect 512 -503 515 -497
rect 519 -503 522 -497
rect 526 -503 529 -497
rect 533 -503 536 -497
rect 540 -503 543 -497
rect 547 -503 550 -497
rect 554 -503 557 -497
rect 561 -503 564 -497
rect 568 -503 571 -497
rect 575 -503 578 -497
rect 582 -503 585 -497
rect 589 -503 595 -497
rect 596 -503 599 -497
rect 603 -503 609 -497
rect 610 -503 616 -497
rect 617 -503 620 -497
rect 624 -503 630 -497
rect 631 -503 634 -497
rect 638 -503 641 -497
rect 645 -503 648 -497
rect 652 -503 655 -497
rect 659 -503 662 -497
rect 666 -503 672 -497
rect 1 -560 7 -554
rect 8 -560 11 -554
rect 15 -560 18 -554
rect 22 -560 25 -554
rect 29 -560 32 -554
rect 36 -560 39 -554
rect 43 -560 46 -554
rect 50 -560 53 -554
rect 57 -560 63 -554
rect 64 -560 67 -554
rect 71 -560 77 -554
rect 78 -560 84 -554
rect 85 -560 88 -554
rect 92 -560 95 -554
rect 99 -560 105 -554
rect 106 -560 109 -554
rect 113 -560 119 -554
rect 120 -560 123 -554
rect 127 -560 133 -554
rect 134 -560 137 -554
rect 141 -560 147 -554
rect 148 -560 154 -554
rect 155 -560 158 -554
rect 162 -560 165 -554
rect 169 -560 172 -554
rect 176 -560 182 -554
rect 183 -560 186 -554
rect 190 -560 196 -554
rect 197 -560 200 -554
rect 204 -560 210 -554
rect 211 -560 214 -554
rect 218 -560 221 -554
rect 225 -560 228 -554
rect 232 -560 235 -554
rect 239 -560 245 -554
rect 246 -560 249 -554
rect 253 -560 256 -554
rect 260 -560 263 -554
rect 267 -560 270 -554
rect 274 -560 280 -554
rect 281 -560 287 -554
rect 288 -560 294 -554
rect 295 -560 298 -554
rect 302 -560 305 -554
rect 309 -560 315 -554
rect 316 -560 322 -554
rect 323 -560 326 -554
rect 330 -560 333 -554
rect 337 -560 343 -554
rect 344 -560 350 -554
rect 351 -560 357 -554
rect 358 -560 364 -554
rect 365 -560 368 -554
rect 372 -560 378 -554
rect 379 -560 382 -554
rect 386 -560 389 -554
rect 393 -560 396 -554
rect 400 -560 406 -554
rect 407 -560 410 -554
rect 414 -560 417 -554
rect 421 -560 427 -554
rect 428 -560 431 -554
rect 435 -560 438 -554
rect 442 -560 445 -554
rect 449 -560 452 -554
rect 456 -560 462 -554
rect 463 -560 466 -554
rect 470 -560 473 -554
rect 477 -560 483 -554
rect 484 -560 487 -554
rect 491 -560 494 -554
rect 498 -560 504 -554
rect 505 -560 508 -554
rect 512 -560 515 -554
rect 519 -560 522 -554
rect 526 -560 529 -554
rect 533 -560 536 -554
rect 540 -560 543 -554
rect 547 -560 550 -554
rect 554 -560 557 -554
rect 561 -560 564 -554
rect 568 -560 571 -554
rect 575 -560 578 -554
rect 582 -560 585 -554
rect 589 -560 592 -554
rect 596 -560 599 -554
rect 603 -560 606 -554
rect 610 -560 613 -554
rect 617 -560 623 -554
rect 624 -560 630 -554
rect 631 -560 634 -554
rect 638 -560 641 -554
rect 645 -560 648 -554
rect 652 -560 655 -554
rect 659 -560 662 -554
rect 666 -560 672 -554
rect 673 -560 676 -554
rect 680 -560 686 -554
rect 687 -560 690 -554
rect 1 -617 4 -611
rect 8 -617 11 -611
rect 15 -617 21 -611
rect 22 -617 25 -611
rect 29 -617 32 -611
rect 36 -617 42 -611
rect 43 -617 49 -611
rect 50 -617 53 -611
rect 57 -617 60 -611
rect 64 -617 67 -611
rect 71 -617 77 -611
rect 78 -617 81 -611
rect 85 -617 91 -611
rect 92 -617 98 -611
rect 99 -617 105 -611
rect 106 -617 109 -611
rect 113 -617 119 -611
rect 120 -617 123 -611
rect 127 -617 133 -611
rect 134 -617 137 -611
rect 141 -617 144 -611
rect 148 -617 151 -611
rect 155 -617 161 -611
rect 162 -617 168 -611
rect 169 -617 175 -611
rect 176 -617 182 -611
rect 183 -617 189 -611
rect 190 -617 193 -611
rect 197 -617 200 -611
rect 204 -617 207 -611
rect 211 -617 214 -611
rect 218 -617 221 -611
rect 225 -617 228 -611
rect 232 -617 238 -611
rect 239 -617 245 -611
rect 246 -617 249 -611
rect 253 -617 256 -611
rect 260 -617 266 -611
rect 267 -617 270 -611
rect 274 -617 280 -611
rect 281 -617 284 -611
rect 288 -617 291 -611
rect 295 -617 298 -611
rect 302 -617 308 -611
rect 309 -617 312 -611
rect 316 -617 319 -611
rect 323 -617 326 -611
rect 330 -617 333 -611
rect 337 -617 340 -611
rect 344 -617 347 -611
rect 351 -617 357 -611
rect 358 -617 361 -611
rect 365 -617 371 -611
rect 372 -617 375 -611
rect 379 -617 385 -611
rect 386 -617 392 -611
rect 393 -617 399 -611
rect 400 -617 403 -611
rect 407 -617 410 -611
rect 414 -617 417 -611
rect 421 -617 424 -611
rect 428 -617 431 -611
rect 435 -617 438 -611
rect 442 -617 445 -611
rect 449 -617 455 -611
rect 456 -617 459 -611
rect 463 -617 469 -611
rect 470 -617 476 -611
rect 477 -617 480 -611
rect 484 -617 487 -611
rect 491 -617 497 -611
rect 498 -617 501 -611
rect 505 -617 508 -611
rect 512 -617 515 -611
rect 519 -617 522 -611
rect 526 -617 529 -611
rect 533 -617 536 -611
rect 540 -617 543 -611
rect 547 -617 550 -611
rect 554 -617 557 -611
rect 561 -617 564 -611
rect 568 -617 571 -611
rect 575 -617 578 -611
rect 582 -617 585 -611
rect 589 -617 592 -611
rect 596 -617 599 -611
rect 603 -617 609 -611
rect 610 -617 613 -611
rect 617 -617 620 -611
rect 624 -617 627 -611
rect 631 -617 634 -611
rect 638 -617 641 -611
rect 645 -617 648 -611
rect 652 -617 658 -611
rect 659 -617 662 -611
rect 673 -617 679 -611
rect 687 -617 693 -611
rect 1 -690 4 -684
rect 8 -690 11 -684
rect 15 -690 21 -684
rect 22 -690 25 -684
rect 29 -690 32 -684
rect 36 -690 39 -684
rect 43 -690 46 -684
rect 50 -690 56 -684
rect 57 -690 63 -684
rect 64 -690 67 -684
rect 71 -690 74 -684
rect 78 -690 84 -684
rect 85 -690 91 -684
rect 92 -690 98 -684
rect 99 -690 105 -684
rect 106 -690 109 -684
rect 113 -690 116 -684
rect 120 -690 123 -684
rect 127 -690 130 -684
rect 134 -690 140 -684
rect 141 -690 147 -684
rect 148 -690 151 -684
rect 155 -690 158 -684
rect 162 -690 168 -684
rect 169 -690 172 -684
rect 176 -690 179 -684
rect 183 -690 189 -684
rect 190 -690 196 -684
rect 197 -690 200 -684
rect 204 -690 207 -684
rect 211 -690 217 -684
rect 218 -690 221 -684
rect 225 -690 231 -684
rect 232 -690 238 -684
rect 239 -690 245 -684
rect 246 -690 249 -684
rect 253 -690 256 -684
rect 260 -690 263 -684
rect 267 -690 270 -684
rect 274 -690 280 -684
rect 281 -690 287 -684
rect 288 -690 291 -684
rect 295 -690 301 -684
rect 302 -690 305 -684
rect 309 -690 312 -684
rect 316 -690 319 -684
rect 323 -690 326 -684
rect 330 -690 333 -684
rect 337 -690 340 -684
rect 344 -690 350 -684
rect 351 -690 354 -684
rect 358 -690 364 -684
rect 365 -690 371 -684
rect 372 -690 378 -684
rect 379 -690 382 -684
rect 386 -690 389 -684
rect 393 -690 396 -684
rect 400 -690 403 -684
rect 407 -690 413 -684
rect 414 -690 417 -684
rect 421 -690 427 -684
rect 428 -690 431 -684
rect 435 -690 438 -684
rect 442 -690 445 -684
rect 449 -690 455 -684
rect 456 -690 462 -684
rect 463 -690 469 -684
rect 470 -690 473 -684
rect 477 -690 480 -684
rect 484 -690 487 -684
rect 491 -690 494 -684
rect 498 -690 501 -684
rect 505 -690 508 -684
rect 512 -690 515 -684
rect 519 -690 522 -684
rect 526 -690 529 -684
rect 533 -690 536 -684
rect 540 -690 543 -684
rect 547 -690 550 -684
rect 554 -690 557 -684
rect 561 -690 564 -684
rect 568 -690 571 -684
rect 575 -690 578 -684
rect 582 -690 585 -684
rect 589 -690 592 -684
rect 596 -690 599 -684
rect 603 -690 606 -684
rect 610 -690 613 -684
rect 617 -690 620 -684
rect 624 -690 627 -684
rect 631 -690 634 -684
rect 638 -690 641 -684
rect 645 -690 648 -684
rect 652 -690 655 -684
rect 659 -690 662 -684
rect 666 -690 669 -684
rect 673 -690 679 -684
rect 680 -690 686 -684
rect 687 -690 690 -684
rect 694 -690 697 -684
rect 701 -690 704 -684
rect 715 -690 721 -684
rect 729 -690 732 -684
rect 1 -757 4 -751
rect 8 -757 11 -751
rect 15 -757 18 -751
rect 22 -757 25 -751
rect 29 -757 32 -751
rect 36 -757 42 -751
rect 43 -757 46 -751
rect 50 -757 53 -751
rect 57 -757 60 -751
rect 64 -757 67 -751
rect 71 -757 74 -751
rect 78 -757 84 -751
rect 85 -757 91 -751
rect 92 -757 95 -751
rect 99 -757 105 -751
rect 106 -757 109 -751
rect 113 -757 116 -751
rect 120 -757 126 -751
rect 127 -757 130 -751
rect 134 -757 137 -751
rect 141 -757 144 -751
rect 148 -757 151 -751
rect 155 -757 158 -751
rect 162 -757 165 -751
rect 169 -757 172 -751
rect 176 -757 179 -751
rect 183 -757 186 -751
rect 190 -757 193 -751
rect 197 -757 203 -751
rect 204 -757 207 -751
rect 211 -757 214 -751
rect 218 -757 221 -751
rect 225 -757 231 -751
rect 232 -757 238 -751
rect 239 -757 242 -751
rect 246 -757 252 -751
rect 253 -757 256 -751
rect 260 -757 263 -751
rect 267 -757 270 -751
rect 274 -757 280 -751
rect 281 -757 287 -751
rect 288 -757 294 -751
rect 295 -757 298 -751
rect 302 -757 305 -751
rect 309 -757 312 -751
rect 316 -757 319 -751
rect 323 -757 329 -751
rect 330 -757 333 -751
rect 337 -757 343 -751
rect 344 -757 347 -751
rect 351 -757 354 -751
rect 358 -757 364 -751
rect 365 -757 368 -751
rect 372 -757 375 -751
rect 379 -757 385 -751
rect 386 -757 392 -751
rect 393 -757 399 -751
rect 400 -757 403 -751
rect 407 -757 413 -751
rect 414 -757 417 -751
rect 421 -757 424 -751
rect 428 -757 434 -751
rect 435 -757 438 -751
rect 442 -757 445 -751
rect 449 -757 455 -751
rect 456 -757 459 -751
rect 463 -757 466 -751
rect 470 -757 473 -751
rect 477 -757 480 -751
rect 484 -757 490 -751
rect 491 -757 497 -751
rect 498 -757 501 -751
rect 505 -757 508 -751
rect 512 -757 515 -751
rect 519 -757 522 -751
rect 526 -757 532 -751
rect 533 -757 536 -751
rect 540 -757 546 -751
rect 547 -757 550 -751
rect 554 -757 557 -751
rect 561 -757 567 -751
rect 568 -757 571 -751
rect 575 -757 578 -751
rect 582 -757 588 -751
rect 589 -757 592 -751
rect 596 -757 599 -751
rect 603 -757 606 -751
rect 610 -757 613 -751
rect 617 -757 620 -751
rect 624 -757 627 -751
rect 631 -757 634 -751
rect 638 -757 641 -751
rect 645 -757 648 -751
rect 652 -757 655 -751
rect 659 -757 662 -751
rect 666 -757 669 -751
rect 673 -757 676 -751
rect 680 -757 683 -751
rect 687 -757 690 -751
rect 694 -757 697 -751
rect 701 -757 704 -751
rect 708 -757 714 -751
rect 715 -757 718 -751
rect 722 -757 725 -751
rect 729 -757 735 -751
rect 736 -757 742 -751
rect 743 -757 746 -751
rect 750 -757 756 -751
rect 799 -757 805 -751
rect 806 -757 809 -751
rect 1 -834 4 -828
rect 8 -834 11 -828
rect 15 -834 18 -828
rect 22 -834 28 -828
rect 29 -834 35 -828
rect 36 -834 39 -828
rect 43 -834 46 -828
rect 50 -834 56 -828
rect 57 -834 60 -828
rect 64 -834 67 -828
rect 71 -834 74 -828
rect 78 -834 84 -828
rect 85 -834 91 -828
rect 92 -834 95 -828
rect 99 -834 102 -828
rect 106 -834 112 -828
rect 113 -834 116 -828
rect 120 -834 126 -828
rect 127 -834 130 -828
rect 134 -834 140 -828
rect 141 -834 147 -828
rect 148 -834 151 -828
rect 155 -834 158 -828
rect 162 -834 168 -828
rect 169 -834 172 -828
rect 176 -834 179 -828
rect 183 -834 186 -828
rect 190 -834 196 -828
rect 197 -834 203 -828
rect 204 -834 207 -828
rect 211 -834 217 -828
rect 218 -834 224 -828
rect 225 -834 228 -828
rect 232 -834 235 -828
rect 239 -834 245 -828
rect 246 -834 249 -828
rect 253 -834 256 -828
rect 260 -834 266 -828
rect 267 -834 270 -828
rect 274 -834 277 -828
rect 281 -834 287 -828
rect 288 -834 294 -828
rect 295 -834 301 -828
rect 302 -834 305 -828
rect 309 -834 312 -828
rect 316 -834 319 -828
rect 323 -834 326 -828
rect 330 -834 336 -828
rect 337 -834 340 -828
rect 344 -834 347 -828
rect 351 -834 354 -828
rect 358 -834 361 -828
rect 365 -834 368 -828
rect 372 -834 375 -828
rect 379 -834 385 -828
rect 386 -834 392 -828
rect 393 -834 396 -828
rect 400 -834 406 -828
rect 407 -834 410 -828
rect 414 -834 420 -828
rect 421 -834 424 -828
rect 428 -834 434 -828
rect 435 -834 441 -828
rect 442 -834 445 -828
rect 449 -834 452 -828
rect 456 -834 462 -828
rect 463 -834 466 -828
rect 470 -834 473 -828
rect 477 -834 480 -828
rect 484 -834 490 -828
rect 491 -834 497 -828
rect 498 -834 501 -828
rect 505 -834 508 -828
rect 512 -834 515 -828
rect 519 -834 525 -828
rect 526 -834 532 -828
rect 533 -834 536 -828
rect 540 -834 543 -828
rect 547 -834 550 -828
rect 554 -834 557 -828
rect 561 -834 564 -828
rect 568 -834 571 -828
rect 575 -834 578 -828
rect 582 -834 585 -828
rect 589 -834 592 -828
rect 596 -834 599 -828
rect 603 -834 606 -828
rect 610 -834 613 -828
rect 617 -834 620 -828
rect 624 -834 627 -828
rect 631 -834 634 -828
rect 638 -834 641 -828
rect 645 -834 648 -828
rect 652 -834 655 -828
rect 659 -834 662 -828
rect 666 -834 669 -828
rect 673 -834 676 -828
rect 680 -834 683 -828
rect 687 -834 690 -828
rect 694 -834 697 -828
rect 701 -834 704 -828
rect 708 -834 711 -828
rect 715 -834 718 -828
rect 722 -834 725 -828
rect 729 -834 732 -828
rect 736 -834 739 -828
rect 743 -834 746 -828
rect 750 -834 753 -828
rect 757 -834 760 -828
rect 764 -834 767 -828
rect 771 -834 774 -828
rect 778 -834 781 -828
rect 785 -834 788 -828
rect 792 -834 795 -828
rect 799 -834 805 -828
rect 806 -834 809 -828
rect 8 -921 11 -915
rect 15 -921 18 -915
rect 22 -921 25 -915
rect 29 -921 32 -915
rect 36 -921 39 -915
rect 43 -921 46 -915
rect 50 -921 53 -915
rect 57 -921 60 -915
rect 64 -921 70 -915
rect 71 -921 77 -915
rect 78 -921 81 -915
rect 85 -921 91 -915
rect 92 -921 95 -915
rect 99 -921 102 -915
rect 106 -921 109 -915
rect 113 -921 116 -915
rect 120 -921 123 -915
rect 127 -921 133 -915
rect 134 -921 137 -915
rect 141 -921 144 -915
rect 148 -921 154 -915
rect 155 -921 161 -915
rect 162 -921 165 -915
rect 169 -921 175 -915
rect 176 -921 182 -915
rect 183 -921 186 -915
rect 190 -921 196 -915
rect 197 -921 203 -915
rect 204 -921 207 -915
rect 211 -921 214 -915
rect 218 -921 224 -915
rect 225 -921 231 -915
rect 232 -921 238 -915
rect 239 -921 245 -915
rect 246 -921 249 -915
rect 253 -921 256 -915
rect 260 -921 263 -915
rect 267 -921 270 -915
rect 274 -921 280 -915
rect 281 -921 287 -915
rect 288 -921 291 -915
rect 295 -921 298 -915
rect 302 -921 305 -915
rect 309 -921 312 -915
rect 316 -921 319 -915
rect 323 -921 326 -915
rect 330 -921 333 -915
rect 337 -921 340 -915
rect 344 -921 350 -915
rect 351 -921 354 -915
rect 358 -921 361 -915
rect 365 -921 371 -915
rect 372 -921 375 -915
rect 379 -921 385 -915
rect 386 -921 389 -915
rect 393 -921 399 -915
rect 400 -921 403 -915
rect 407 -921 413 -915
rect 414 -921 420 -915
rect 421 -921 424 -915
rect 428 -921 431 -915
rect 435 -921 438 -915
rect 442 -921 445 -915
rect 449 -921 455 -915
rect 456 -921 462 -915
rect 463 -921 469 -915
rect 470 -921 473 -915
rect 477 -921 480 -915
rect 484 -921 490 -915
rect 491 -921 494 -915
rect 498 -921 504 -915
rect 505 -921 508 -915
rect 512 -921 515 -915
rect 519 -921 522 -915
rect 526 -921 529 -915
rect 533 -921 536 -915
rect 540 -921 543 -915
rect 547 -921 550 -915
rect 554 -921 557 -915
rect 561 -921 564 -915
rect 568 -921 571 -915
rect 575 -921 581 -915
rect 582 -921 585 -915
rect 589 -921 592 -915
rect 596 -921 599 -915
rect 603 -921 606 -915
rect 610 -921 613 -915
rect 617 -921 620 -915
rect 624 -921 627 -915
rect 631 -921 634 -915
rect 638 -921 641 -915
rect 645 -921 648 -915
rect 652 -921 655 -915
rect 659 -921 662 -915
rect 666 -921 669 -915
rect 673 -921 676 -915
rect 680 -921 683 -915
rect 687 -921 690 -915
rect 694 -921 697 -915
rect 701 -921 704 -915
rect 708 -921 711 -915
rect 715 -921 718 -915
rect 722 -921 725 -915
rect 729 -921 732 -915
rect 736 -921 739 -915
rect 743 -921 746 -915
rect 750 -921 753 -915
rect 757 -921 760 -915
rect 764 -921 767 -915
rect 771 -921 777 -915
rect 778 -921 784 -915
rect 785 -921 788 -915
rect 792 -921 798 -915
rect 8 -998 11 -992
rect 15 -998 18 -992
rect 22 -998 25 -992
rect 29 -998 32 -992
rect 36 -998 39 -992
rect 43 -998 46 -992
rect 50 -998 53 -992
rect 57 -998 60 -992
rect 64 -998 67 -992
rect 71 -998 77 -992
rect 78 -998 84 -992
rect 85 -998 88 -992
rect 92 -998 98 -992
rect 99 -998 105 -992
rect 106 -998 109 -992
rect 113 -998 119 -992
rect 120 -998 123 -992
rect 127 -998 130 -992
rect 134 -998 137 -992
rect 141 -998 144 -992
rect 148 -998 151 -992
rect 155 -998 161 -992
rect 162 -998 165 -992
rect 169 -998 172 -992
rect 176 -998 179 -992
rect 183 -998 186 -992
rect 190 -998 193 -992
rect 197 -998 203 -992
rect 204 -998 207 -992
rect 211 -998 214 -992
rect 218 -998 224 -992
rect 225 -998 228 -992
rect 232 -998 238 -992
rect 239 -998 245 -992
rect 246 -998 249 -992
rect 253 -998 259 -992
rect 260 -998 263 -992
rect 267 -998 270 -992
rect 274 -998 277 -992
rect 281 -998 287 -992
rect 288 -998 291 -992
rect 295 -998 298 -992
rect 302 -998 305 -992
rect 309 -998 315 -992
rect 316 -998 322 -992
rect 323 -998 326 -992
rect 330 -998 333 -992
rect 337 -998 340 -992
rect 344 -998 350 -992
rect 351 -998 357 -992
rect 358 -998 364 -992
rect 365 -998 371 -992
rect 372 -998 378 -992
rect 379 -998 382 -992
rect 386 -998 392 -992
rect 393 -998 399 -992
rect 400 -998 403 -992
rect 407 -998 410 -992
rect 414 -998 420 -992
rect 421 -998 427 -992
rect 428 -998 434 -992
rect 435 -998 438 -992
rect 442 -998 448 -992
rect 449 -998 455 -992
rect 456 -998 459 -992
rect 463 -998 469 -992
rect 470 -998 476 -992
rect 477 -998 480 -992
rect 484 -998 487 -992
rect 491 -998 494 -992
rect 498 -998 501 -992
rect 505 -998 508 -992
rect 512 -998 515 -992
rect 519 -998 522 -992
rect 526 -998 529 -992
rect 533 -998 539 -992
rect 540 -998 543 -992
rect 547 -998 550 -992
rect 554 -998 557 -992
rect 561 -998 564 -992
rect 568 -998 571 -992
rect 575 -998 578 -992
rect 582 -998 585 -992
rect 589 -998 592 -992
rect 596 -998 599 -992
rect 603 -998 606 -992
rect 610 -998 613 -992
rect 617 -998 620 -992
rect 624 -998 627 -992
rect 631 -998 634 -992
rect 638 -998 641 -992
rect 645 -998 648 -992
rect 652 -998 655 -992
rect 659 -998 662 -992
rect 666 -998 669 -992
rect 673 -998 676 -992
rect 680 -998 683 -992
rect 687 -998 690 -992
rect 694 -998 697 -992
rect 701 -998 704 -992
rect 708 -998 711 -992
rect 715 -998 718 -992
rect 722 -998 725 -992
rect 729 -998 732 -992
rect 736 -998 742 -992
rect 743 -998 749 -992
rect 750 -998 756 -992
rect 757 -998 760 -992
rect 22 -1073 25 -1067
rect 29 -1073 35 -1067
rect 36 -1073 39 -1067
rect 43 -1073 46 -1067
rect 50 -1073 53 -1067
rect 57 -1073 63 -1067
rect 64 -1073 67 -1067
rect 71 -1073 77 -1067
rect 78 -1073 81 -1067
rect 85 -1073 91 -1067
rect 92 -1073 95 -1067
rect 99 -1073 105 -1067
rect 106 -1073 112 -1067
rect 113 -1073 116 -1067
rect 120 -1073 123 -1067
rect 127 -1073 130 -1067
rect 134 -1073 137 -1067
rect 141 -1073 144 -1067
rect 148 -1073 154 -1067
rect 155 -1073 158 -1067
rect 162 -1073 168 -1067
rect 169 -1073 172 -1067
rect 176 -1073 182 -1067
rect 183 -1073 186 -1067
rect 190 -1073 196 -1067
rect 197 -1073 203 -1067
rect 204 -1073 207 -1067
rect 211 -1073 214 -1067
rect 218 -1073 221 -1067
rect 225 -1073 228 -1067
rect 232 -1073 235 -1067
rect 239 -1073 245 -1067
rect 246 -1073 252 -1067
rect 253 -1073 256 -1067
rect 260 -1073 263 -1067
rect 267 -1073 270 -1067
rect 274 -1073 280 -1067
rect 281 -1073 284 -1067
rect 288 -1073 291 -1067
rect 295 -1073 298 -1067
rect 302 -1073 305 -1067
rect 309 -1073 315 -1067
rect 316 -1073 319 -1067
rect 323 -1073 326 -1067
rect 330 -1073 336 -1067
rect 337 -1073 340 -1067
rect 344 -1073 347 -1067
rect 351 -1073 354 -1067
rect 358 -1073 361 -1067
rect 365 -1073 368 -1067
rect 372 -1073 375 -1067
rect 379 -1073 382 -1067
rect 386 -1073 389 -1067
rect 393 -1073 396 -1067
rect 400 -1073 406 -1067
rect 407 -1073 413 -1067
rect 414 -1073 420 -1067
rect 421 -1073 427 -1067
rect 428 -1073 431 -1067
rect 435 -1073 441 -1067
rect 442 -1073 445 -1067
rect 449 -1073 455 -1067
rect 456 -1073 459 -1067
rect 463 -1073 466 -1067
rect 470 -1073 476 -1067
rect 477 -1073 483 -1067
rect 484 -1073 487 -1067
rect 491 -1073 497 -1067
rect 498 -1073 501 -1067
rect 505 -1073 511 -1067
rect 512 -1073 515 -1067
rect 519 -1073 525 -1067
rect 526 -1073 529 -1067
rect 533 -1073 539 -1067
rect 540 -1073 546 -1067
rect 547 -1073 550 -1067
rect 554 -1073 557 -1067
rect 561 -1073 567 -1067
rect 568 -1073 571 -1067
rect 575 -1073 578 -1067
rect 582 -1073 585 -1067
rect 589 -1073 592 -1067
rect 596 -1073 599 -1067
rect 603 -1073 606 -1067
rect 610 -1073 613 -1067
rect 617 -1073 620 -1067
rect 624 -1073 627 -1067
rect 631 -1073 634 -1067
rect 638 -1073 641 -1067
rect 645 -1073 648 -1067
rect 652 -1073 655 -1067
rect 659 -1073 662 -1067
rect 666 -1073 669 -1067
rect 673 -1073 676 -1067
rect 680 -1073 683 -1067
rect 687 -1073 693 -1067
rect 694 -1073 697 -1067
rect 701 -1073 704 -1067
rect 708 -1073 711 -1067
rect 715 -1073 721 -1067
rect 722 -1073 725 -1067
rect 729 -1073 732 -1067
rect 736 -1073 739 -1067
rect 8 -1134 11 -1128
rect 15 -1134 18 -1128
rect 22 -1134 25 -1128
rect 29 -1134 35 -1128
rect 36 -1134 39 -1128
rect 43 -1134 49 -1128
rect 50 -1134 53 -1128
rect 57 -1134 60 -1128
rect 64 -1134 70 -1128
rect 71 -1134 74 -1128
rect 78 -1134 84 -1128
rect 85 -1134 88 -1128
rect 92 -1134 98 -1128
rect 99 -1134 102 -1128
rect 106 -1134 109 -1128
rect 113 -1134 116 -1128
rect 120 -1134 126 -1128
rect 127 -1134 130 -1128
rect 134 -1134 137 -1128
rect 141 -1134 147 -1128
rect 148 -1134 151 -1128
rect 155 -1134 161 -1128
rect 162 -1134 168 -1128
rect 169 -1134 175 -1128
rect 176 -1134 182 -1128
rect 183 -1134 189 -1128
rect 190 -1134 196 -1128
rect 197 -1134 203 -1128
rect 204 -1134 207 -1128
rect 211 -1134 217 -1128
rect 218 -1134 221 -1128
rect 225 -1134 228 -1128
rect 232 -1134 235 -1128
rect 239 -1134 245 -1128
rect 246 -1134 252 -1128
rect 253 -1134 256 -1128
rect 260 -1134 263 -1128
rect 267 -1134 270 -1128
rect 274 -1134 280 -1128
rect 281 -1134 284 -1128
rect 288 -1134 291 -1128
rect 295 -1134 298 -1128
rect 302 -1134 305 -1128
rect 309 -1134 315 -1128
rect 316 -1134 319 -1128
rect 323 -1134 326 -1128
rect 330 -1134 336 -1128
rect 337 -1134 340 -1128
rect 344 -1134 350 -1128
rect 351 -1134 354 -1128
rect 358 -1134 364 -1128
rect 365 -1134 371 -1128
rect 372 -1134 378 -1128
rect 379 -1134 385 -1128
rect 386 -1134 392 -1128
rect 393 -1134 399 -1128
rect 400 -1134 403 -1128
rect 407 -1134 410 -1128
rect 414 -1134 417 -1128
rect 421 -1134 427 -1128
rect 428 -1134 434 -1128
rect 435 -1134 438 -1128
rect 442 -1134 445 -1128
rect 449 -1134 452 -1128
rect 456 -1134 459 -1128
rect 463 -1134 466 -1128
rect 470 -1134 473 -1128
rect 477 -1134 480 -1128
rect 484 -1134 487 -1128
rect 491 -1134 494 -1128
rect 498 -1134 501 -1128
rect 505 -1134 511 -1128
rect 512 -1134 515 -1128
rect 519 -1134 525 -1128
rect 526 -1134 529 -1128
rect 533 -1134 536 -1128
rect 540 -1134 543 -1128
rect 547 -1134 550 -1128
rect 554 -1134 557 -1128
rect 561 -1134 564 -1128
rect 568 -1134 571 -1128
rect 575 -1134 578 -1128
rect 582 -1134 585 -1128
rect 589 -1134 592 -1128
rect 596 -1134 599 -1128
rect 603 -1134 606 -1128
rect 610 -1134 613 -1128
rect 617 -1134 620 -1128
rect 624 -1134 627 -1128
rect 631 -1134 634 -1128
rect 638 -1134 641 -1128
rect 645 -1134 648 -1128
rect 652 -1134 655 -1128
rect 659 -1134 662 -1128
rect 666 -1134 669 -1128
rect 673 -1134 679 -1128
rect 680 -1134 686 -1128
rect 687 -1134 690 -1128
rect 694 -1134 697 -1128
rect 701 -1134 704 -1128
rect 708 -1134 711 -1128
rect 1 -1191 4 -1185
rect 8 -1191 11 -1185
rect 15 -1191 21 -1185
rect 22 -1191 28 -1185
rect 29 -1191 32 -1185
rect 36 -1191 39 -1185
rect 43 -1191 46 -1185
rect 50 -1191 53 -1185
rect 57 -1191 60 -1185
rect 64 -1191 70 -1185
rect 71 -1191 77 -1185
rect 78 -1191 81 -1185
rect 85 -1191 91 -1185
rect 92 -1191 95 -1185
rect 99 -1191 105 -1185
rect 106 -1191 112 -1185
rect 113 -1191 119 -1185
rect 120 -1191 123 -1185
rect 127 -1191 130 -1185
rect 134 -1191 137 -1185
rect 141 -1191 147 -1185
rect 148 -1191 154 -1185
rect 155 -1191 161 -1185
rect 162 -1191 165 -1185
rect 169 -1191 175 -1185
rect 176 -1191 179 -1185
rect 183 -1191 186 -1185
rect 190 -1191 196 -1185
rect 197 -1191 200 -1185
rect 204 -1191 210 -1185
rect 211 -1191 217 -1185
rect 218 -1191 221 -1185
rect 225 -1191 228 -1185
rect 232 -1191 238 -1185
rect 239 -1191 242 -1185
rect 246 -1191 249 -1185
rect 253 -1191 256 -1185
rect 260 -1191 263 -1185
rect 267 -1191 270 -1185
rect 274 -1191 280 -1185
rect 281 -1191 284 -1185
rect 288 -1191 291 -1185
rect 295 -1191 298 -1185
rect 302 -1191 308 -1185
rect 309 -1191 312 -1185
rect 316 -1191 322 -1185
rect 323 -1191 329 -1185
rect 330 -1191 336 -1185
rect 337 -1191 343 -1185
rect 344 -1191 350 -1185
rect 351 -1191 354 -1185
rect 358 -1191 361 -1185
rect 365 -1191 368 -1185
rect 372 -1191 375 -1185
rect 379 -1191 382 -1185
rect 386 -1191 392 -1185
rect 393 -1191 396 -1185
rect 400 -1191 403 -1185
rect 407 -1191 410 -1185
rect 414 -1191 417 -1185
rect 421 -1191 424 -1185
rect 428 -1191 431 -1185
rect 435 -1191 441 -1185
rect 442 -1191 448 -1185
rect 449 -1191 455 -1185
rect 456 -1191 459 -1185
rect 463 -1191 469 -1185
rect 470 -1191 473 -1185
rect 477 -1191 480 -1185
rect 484 -1191 487 -1185
rect 491 -1191 494 -1185
rect 498 -1191 501 -1185
rect 505 -1191 508 -1185
rect 512 -1191 515 -1185
rect 519 -1191 522 -1185
rect 526 -1191 532 -1185
rect 533 -1191 536 -1185
rect 540 -1191 546 -1185
rect 547 -1191 550 -1185
rect 554 -1191 557 -1185
rect 561 -1191 564 -1185
rect 568 -1191 571 -1185
rect 575 -1191 578 -1185
rect 582 -1191 585 -1185
rect 589 -1191 592 -1185
rect 596 -1191 599 -1185
rect 603 -1191 606 -1185
rect 610 -1191 613 -1185
rect 617 -1191 620 -1185
rect 624 -1191 627 -1185
rect 631 -1191 634 -1185
rect 638 -1191 641 -1185
rect 645 -1191 648 -1185
rect 652 -1191 658 -1185
rect 659 -1191 662 -1185
rect 666 -1191 672 -1185
rect 673 -1191 679 -1185
rect 680 -1191 683 -1185
rect 687 -1191 690 -1185
rect 701 -1191 704 -1185
rect 708 -1191 711 -1185
rect 1 -1262 4 -1256
rect 8 -1262 11 -1256
rect 15 -1262 18 -1256
rect 22 -1262 25 -1256
rect 29 -1262 32 -1256
rect 36 -1262 39 -1256
rect 43 -1262 49 -1256
rect 50 -1262 56 -1256
rect 57 -1262 63 -1256
rect 64 -1262 67 -1256
rect 71 -1262 77 -1256
rect 78 -1262 81 -1256
rect 85 -1262 88 -1256
rect 92 -1262 95 -1256
rect 99 -1262 105 -1256
rect 106 -1262 112 -1256
rect 113 -1262 116 -1256
rect 120 -1262 126 -1256
rect 127 -1262 130 -1256
rect 134 -1262 137 -1256
rect 141 -1262 147 -1256
rect 148 -1262 151 -1256
rect 155 -1262 158 -1256
rect 162 -1262 168 -1256
rect 169 -1262 172 -1256
rect 176 -1262 182 -1256
rect 183 -1262 189 -1256
rect 190 -1262 196 -1256
rect 197 -1262 203 -1256
rect 204 -1262 207 -1256
rect 211 -1262 217 -1256
rect 218 -1262 224 -1256
rect 225 -1262 231 -1256
rect 232 -1262 238 -1256
rect 239 -1262 242 -1256
rect 246 -1262 252 -1256
rect 253 -1262 259 -1256
rect 260 -1262 263 -1256
rect 267 -1262 273 -1256
rect 274 -1262 277 -1256
rect 281 -1262 284 -1256
rect 288 -1262 291 -1256
rect 295 -1262 298 -1256
rect 302 -1262 308 -1256
rect 309 -1262 315 -1256
rect 316 -1262 319 -1256
rect 323 -1262 329 -1256
rect 330 -1262 336 -1256
rect 337 -1262 340 -1256
rect 344 -1262 347 -1256
rect 351 -1262 357 -1256
rect 358 -1262 361 -1256
rect 365 -1262 368 -1256
rect 372 -1262 375 -1256
rect 379 -1262 385 -1256
rect 386 -1262 389 -1256
rect 393 -1262 399 -1256
rect 400 -1262 403 -1256
rect 407 -1262 410 -1256
rect 414 -1262 417 -1256
rect 421 -1262 424 -1256
rect 428 -1262 434 -1256
rect 435 -1262 438 -1256
rect 442 -1262 445 -1256
rect 449 -1262 455 -1256
rect 456 -1262 462 -1256
rect 463 -1262 466 -1256
rect 470 -1262 473 -1256
rect 477 -1262 480 -1256
rect 484 -1262 487 -1256
rect 491 -1262 497 -1256
rect 498 -1262 501 -1256
rect 505 -1262 508 -1256
rect 512 -1262 518 -1256
rect 519 -1262 522 -1256
rect 526 -1262 529 -1256
rect 533 -1262 536 -1256
rect 540 -1262 543 -1256
rect 547 -1262 550 -1256
rect 554 -1262 557 -1256
rect 561 -1262 564 -1256
rect 568 -1262 571 -1256
rect 575 -1262 578 -1256
rect 582 -1262 585 -1256
rect 589 -1262 592 -1256
rect 596 -1262 599 -1256
rect 603 -1262 606 -1256
rect 610 -1262 613 -1256
rect 617 -1262 620 -1256
rect 624 -1262 627 -1256
rect 631 -1262 634 -1256
rect 638 -1262 641 -1256
rect 645 -1262 648 -1256
rect 652 -1262 655 -1256
rect 659 -1262 662 -1256
rect 666 -1262 669 -1256
rect 673 -1262 676 -1256
rect 680 -1262 683 -1256
rect 687 -1262 690 -1256
rect 694 -1262 697 -1256
rect 701 -1262 707 -1256
rect 708 -1262 714 -1256
rect 715 -1262 718 -1256
rect 1 -1333 4 -1327
rect 8 -1333 11 -1327
rect 15 -1333 21 -1327
rect 22 -1333 25 -1327
rect 29 -1333 35 -1327
rect 36 -1333 42 -1327
rect 43 -1333 46 -1327
rect 50 -1333 53 -1327
rect 57 -1333 60 -1327
rect 64 -1333 67 -1327
rect 71 -1333 77 -1327
rect 78 -1333 84 -1327
rect 85 -1333 88 -1327
rect 92 -1333 95 -1327
rect 99 -1333 102 -1327
rect 106 -1333 109 -1327
rect 113 -1333 116 -1327
rect 120 -1333 123 -1327
rect 127 -1333 133 -1327
rect 134 -1333 140 -1327
rect 141 -1333 144 -1327
rect 148 -1333 154 -1327
rect 155 -1333 158 -1327
rect 162 -1333 165 -1327
rect 169 -1333 175 -1327
rect 176 -1333 182 -1327
rect 183 -1333 186 -1327
rect 190 -1333 193 -1327
rect 197 -1333 200 -1327
rect 204 -1333 210 -1327
rect 211 -1333 214 -1327
rect 218 -1333 221 -1327
rect 225 -1333 228 -1327
rect 232 -1333 238 -1327
rect 239 -1333 242 -1327
rect 246 -1333 249 -1327
rect 253 -1333 256 -1327
rect 260 -1333 263 -1327
rect 267 -1333 270 -1327
rect 274 -1333 277 -1327
rect 281 -1333 287 -1327
rect 288 -1333 291 -1327
rect 295 -1333 301 -1327
rect 302 -1333 308 -1327
rect 309 -1333 312 -1327
rect 316 -1333 319 -1327
rect 323 -1333 329 -1327
rect 330 -1333 333 -1327
rect 337 -1333 343 -1327
rect 344 -1333 347 -1327
rect 351 -1333 357 -1327
rect 358 -1333 364 -1327
rect 365 -1333 371 -1327
rect 372 -1333 378 -1327
rect 379 -1333 385 -1327
rect 386 -1333 392 -1327
rect 393 -1333 399 -1327
rect 400 -1333 403 -1327
rect 407 -1333 413 -1327
rect 414 -1333 417 -1327
rect 421 -1333 427 -1327
rect 428 -1333 431 -1327
rect 435 -1333 438 -1327
rect 442 -1333 445 -1327
rect 449 -1333 455 -1327
rect 456 -1333 459 -1327
rect 463 -1333 469 -1327
rect 470 -1333 476 -1327
rect 477 -1333 483 -1327
rect 484 -1333 487 -1327
rect 491 -1333 494 -1327
rect 498 -1333 504 -1327
rect 505 -1333 508 -1327
rect 512 -1333 515 -1327
rect 519 -1333 522 -1327
rect 526 -1333 529 -1327
rect 533 -1333 536 -1327
rect 540 -1333 543 -1327
rect 547 -1333 550 -1327
rect 554 -1333 557 -1327
rect 561 -1333 564 -1327
rect 568 -1333 571 -1327
rect 575 -1333 578 -1327
rect 582 -1333 585 -1327
rect 589 -1333 592 -1327
rect 596 -1333 599 -1327
rect 603 -1333 606 -1327
rect 610 -1333 613 -1327
rect 617 -1333 620 -1327
rect 624 -1333 627 -1327
rect 631 -1333 634 -1327
rect 638 -1333 641 -1327
rect 645 -1333 651 -1327
rect 652 -1333 655 -1327
rect 659 -1333 665 -1327
rect 666 -1333 672 -1327
rect 673 -1333 676 -1327
rect 680 -1333 683 -1327
rect 701 -1333 704 -1327
rect 29 -1392 35 -1386
rect 36 -1392 39 -1386
rect 43 -1392 46 -1386
rect 50 -1392 53 -1386
rect 57 -1392 60 -1386
rect 64 -1392 67 -1386
rect 71 -1392 74 -1386
rect 78 -1392 81 -1386
rect 85 -1392 88 -1386
rect 92 -1392 95 -1386
rect 99 -1392 105 -1386
rect 106 -1392 109 -1386
rect 113 -1392 116 -1386
rect 120 -1392 126 -1386
rect 127 -1392 130 -1386
rect 134 -1392 140 -1386
rect 141 -1392 147 -1386
rect 148 -1392 151 -1386
rect 155 -1392 161 -1386
rect 162 -1392 165 -1386
rect 169 -1392 172 -1386
rect 176 -1392 179 -1386
rect 183 -1392 189 -1386
rect 190 -1392 196 -1386
rect 197 -1392 203 -1386
rect 204 -1392 210 -1386
rect 211 -1392 214 -1386
rect 218 -1392 224 -1386
rect 225 -1392 228 -1386
rect 232 -1392 238 -1386
rect 239 -1392 245 -1386
rect 246 -1392 252 -1386
rect 253 -1392 256 -1386
rect 260 -1392 263 -1386
rect 267 -1392 270 -1386
rect 274 -1392 277 -1386
rect 281 -1392 287 -1386
rect 288 -1392 291 -1386
rect 295 -1392 298 -1386
rect 302 -1392 305 -1386
rect 309 -1392 312 -1386
rect 316 -1392 319 -1386
rect 323 -1392 326 -1386
rect 330 -1392 333 -1386
rect 337 -1392 340 -1386
rect 344 -1392 350 -1386
rect 351 -1392 354 -1386
rect 358 -1392 364 -1386
rect 365 -1392 371 -1386
rect 372 -1392 375 -1386
rect 379 -1392 385 -1386
rect 386 -1392 392 -1386
rect 393 -1392 396 -1386
rect 400 -1392 406 -1386
rect 407 -1392 410 -1386
rect 414 -1392 420 -1386
rect 421 -1392 427 -1386
rect 428 -1392 434 -1386
rect 435 -1392 438 -1386
rect 442 -1392 445 -1386
rect 449 -1392 452 -1386
rect 456 -1392 462 -1386
rect 463 -1392 469 -1386
rect 470 -1392 473 -1386
rect 477 -1392 483 -1386
rect 484 -1392 487 -1386
rect 491 -1392 494 -1386
rect 498 -1392 501 -1386
rect 505 -1392 508 -1386
rect 512 -1392 515 -1386
rect 519 -1392 522 -1386
rect 526 -1392 529 -1386
rect 533 -1392 536 -1386
rect 540 -1392 543 -1386
rect 547 -1392 550 -1386
rect 554 -1392 557 -1386
rect 561 -1392 564 -1386
rect 568 -1392 571 -1386
rect 575 -1392 578 -1386
rect 582 -1392 585 -1386
rect 589 -1392 592 -1386
rect 596 -1392 602 -1386
rect 603 -1392 606 -1386
rect 610 -1392 613 -1386
rect 617 -1392 623 -1386
rect 624 -1392 627 -1386
rect 631 -1392 637 -1386
rect 638 -1392 641 -1386
rect 645 -1392 648 -1386
rect 652 -1392 658 -1386
rect 659 -1392 662 -1386
rect 666 -1392 669 -1386
rect 701 -1392 707 -1386
rect 36 -1451 39 -1445
rect 43 -1451 46 -1445
rect 50 -1451 53 -1445
rect 57 -1451 60 -1445
rect 64 -1451 67 -1445
rect 71 -1451 74 -1445
rect 78 -1451 81 -1445
rect 85 -1451 88 -1445
rect 92 -1451 95 -1445
rect 99 -1451 105 -1445
rect 106 -1451 109 -1445
rect 113 -1451 119 -1445
rect 120 -1451 126 -1445
rect 127 -1451 130 -1445
rect 134 -1451 140 -1445
rect 141 -1451 147 -1445
rect 148 -1451 151 -1445
rect 155 -1451 161 -1445
rect 162 -1451 165 -1445
rect 169 -1451 172 -1445
rect 176 -1451 179 -1445
rect 183 -1451 189 -1445
rect 190 -1451 193 -1445
rect 197 -1451 203 -1445
rect 204 -1451 207 -1445
rect 211 -1451 217 -1445
rect 218 -1451 221 -1445
rect 225 -1451 231 -1445
rect 232 -1451 238 -1445
rect 239 -1451 245 -1445
rect 246 -1451 249 -1445
rect 253 -1451 256 -1445
rect 260 -1451 263 -1445
rect 267 -1451 273 -1445
rect 274 -1451 277 -1445
rect 281 -1451 284 -1445
rect 288 -1451 291 -1445
rect 295 -1451 298 -1445
rect 302 -1451 305 -1445
rect 309 -1451 312 -1445
rect 316 -1451 319 -1445
rect 323 -1451 329 -1445
rect 330 -1451 333 -1445
rect 337 -1451 340 -1445
rect 344 -1451 347 -1445
rect 351 -1451 357 -1445
rect 358 -1451 364 -1445
rect 365 -1451 371 -1445
rect 372 -1451 378 -1445
rect 379 -1451 382 -1445
rect 386 -1451 392 -1445
rect 393 -1451 399 -1445
rect 400 -1451 403 -1445
rect 407 -1451 410 -1445
rect 414 -1451 417 -1445
rect 421 -1451 424 -1445
rect 428 -1451 431 -1445
rect 435 -1451 441 -1445
rect 442 -1451 448 -1445
rect 449 -1451 455 -1445
rect 456 -1451 459 -1445
rect 463 -1451 469 -1445
rect 470 -1451 473 -1445
rect 477 -1451 483 -1445
rect 484 -1451 487 -1445
rect 491 -1451 494 -1445
rect 498 -1451 501 -1445
rect 505 -1451 508 -1445
rect 512 -1451 515 -1445
rect 519 -1451 522 -1445
rect 526 -1451 529 -1445
rect 533 -1451 536 -1445
rect 540 -1451 543 -1445
rect 547 -1451 553 -1445
rect 554 -1451 557 -1445
rect 561 -1451 567 -1445
rect 568 -1451 574 -1445
rect 575 -1451 578 -1445
rect 582 -1451 585 -1445
rect 589 -1451 592 -1445
rect 596 -1451 599 -1445
rect 603 -1451 606 -1445
rect 645 -1451 651 -1445
rect 701 -1451 707 -1445
rect 708 -1451 714 -1445
rect 15 -1504 18 -1498
rect 22 -1504 28 -1498
rect 29 -1504 32 -1498
rect 36 -1504 39 -1498
rect 43 -1504 49 -1498
rect 50 -1504 56 -1498
rect 57 -1504 60 -1498
rect 64 -1504 67 -1498
rect 71 -1504 74 -1498
rect 78 -1504 81 -1498
rect 85 -1504 91 -1498
rect 92 -1504 95 -1498
rect 99 -1504 102 -1498
rect 106 -1504 112 -1498
rect 113 -1504 116 -1498
rect 120 -1504 126 -1498
rect 127 -1504 130 -1498
rect 134 -1504 137 -1498
rect 141 -1504 144 -1498
rect 148 -1504 154 -1498
rect 155 -1504 161 -1498
rect 162 -1504 168 -1498
rect 169 -1504 175 -1498
rect 176 -1504 182 -1498
rect 183 -1504 189 -1498
rect 190 -1504 193 -1498
rect 197 -1504 200 -1498
rect 204 -1504 210 -1498
rect 211 -1504 214 -1498
rect 218 -1504 221 -1498
rect 225 -1504 231 -1498
rect 232 -1504 238 -1498
rect 239 -1504 245 -1498
rect 246 -1504 252 -1498
rect 253 -1504 256 -1498
rect 260 -1504 263 -1498
rect 267 -1504 273 -1498
rect 274 -1504 277 -1498
rect 281 -1504 284 -1498
rect 288 -1504 294 -1498
rect 295 -1504 298 -1498
rect 302 -1504 308 -1498
rect 309 -1504 315 -1498
rect 316 -1504 322 -1498
rect 323 -1504 329 -1498
rect 330 -1504 333 -1498
rect 337 -1504 340 -1498
rect 344 -1504 347 -1498
rect 351 -1504 354 -1498
rect 358 -1504 361 -1498
rect 365 -1504 371 -1498
rect 372 -1504 375 -1498
rect 379 -1504 382 -1498
rect 386 -1504 389 -1498
rect 393 -1504 396 -1498
rect 400 -1504 403 -1498
rect 407 -1504 410 -1498
rect 414 -1504 417 -1498
rect 421 -1504 427 -1498
rect 428 -1504 434 -1498
rect 435 -1504 438 -1498
rect 442 -1504 445 -1498
rect 449 -1504 452 -1498
rect 456 -1504 459 -1498
rect 463 -1504 466 -1498
rect 470 -1504 473 -1498
rect 477 -1504 483 -1498
rect 484 -1504 487 -1498
rect 491 -1504 494 -1498
rect 498 -1504 501 -1498
rect 505 -1504 508 -1498
rect 512 -1504 515 -1498
rect 519 -1504 522 -1498
rect 526 -1504 529 -1498
rect 533 -1504 536 -1498
rect 540 -1504 543 -1498
rect 547 -1504 550 -1498
rect 554 -1504 557 -1498
rect 561 -1504 567 -1498
rect 568 -1504 571 -1498
rect 575 -1504 581 -1498
rect 582 -1504 585 -1498
rect 589 -1504 592 -1498
rect 50 -1553 53 -1547
rect 57 -1553 63 -1547
rect 64 -1553 67 -1547
rect 71 -1553 77 -1547
rect 78 -1553 81 -1547
rect 85 -1553 88 -1547
rect 92 -1553 98 -1547
rect 99 -1553 105 -1547
rect 106 -1553 112 -1547
rect 113 -1553 116 -1547
rect 120 -1553 123 -1547
rect 127 -1553 130 -1547
rect 134 -1553 137 -1547
rect 141 -1553 144 -1547
rect 148 -1553 154 -1547
rect 155 -1553 161 -1547
rect 162 -1553 165 -1547
rect 169 -1553 175 -1547
rect 176 -1553 179 -1547
rect 183 -1553 186 -1547
rect 190 -1553 196 -1547
rect 197 -1553 203 -1547
rect 204 -1553 207 -1547
rect 211 -1553 214 -1547
rect 218 -1553 224 -1547
rect 225 -1553 231 -1547
rect 232 -1553 238 -1547
rect 239 -1553 245 -1547
rect 246 -1553 249 -1547
rect 253 -1553 256 -1547
rect 260 -1553 263 -1547
rect 267 -1553 270 -1547
rect 274 -1553 277 -1547
rect 281 -1553 287 -1547
rect 288 -1553 294 -1547
rect 295 -1553 298 -1547
rect 302 -1553 305 -1547
rect 309 -1553 312 -1547
rect 316 -1553 319 -1547
rect 323 -1553 329 -1547
rect 330 -1553 333 -1547
rect 337 -1553 340 -1547
rect 344 -1553 347 -1547
rect 351 -1553 354 -1547
rect 358 -1553 361 -1547
rect 365 -1553 371 -1547
rect 372 -1553 375 -1547
rect 379 -1553 385 -1547
rect 386 -1553 392 -1547
rect 393 -1553 396 -1547
rect 400 -1553 403 -1547
rect 407 -1553 410 -1547
rect 414 -1553 420 -1547
rect 421 -1553 427 -1547
rect 428 -1553 431 -1547
rect 435 -1553 438 -1547
rect 442 -1553 445 -1547
rect 449 -1553 452 -1547
rect 456 -1553 459 -1547
rect 463 -1553 466 -1547
rect 470 -1553 476 -1547
rect 477 -1553 480 -1547
rect 484 -1553 490 -1547
rect 491 -1553 494 -1547
rect 498 -1553 504 -1547
rect 505 -1553 508 -1547
rect 512 -1553 515 -1547
rect 519 -1553 522 -1547
rect 526 -1553 529 -1547
rect 582 -1553 588 -1547
rect 589 -1553 592 -1547
rect 71 -1590 77 -1584
rect 78 -1590 81 -1584
rect 127 -1590 130 -1584
rect 134 -1590 137 -1584
rect 141 -1590 147 -1584
rect 148 -1590 154 -1584
rect 155 -1590 161 -1584
rect 162 -1590 165 -1584
rect 169 -1590 172 -1584
rect 176 -1590 182 -1584
rect 183 -1590 189 -1584
rect 190 -1590 196 -1584
rect 197 -1590 203 -1584
rect 204 -1590 210 -1584
rect 211 -1590 214 -1584
rect 218 -1590 224 -1584
rect 225 -1590 231 -1584
rect 232 -1590 235 -1584
rect 239 -1590 245 -1584
rect 246 -1590 249 -1584
rect 253 -1590 256 -1584
rect 260 -1590 263 -1584
rect 267 -1590 273 -1584
rect 274 -1590 277 -1584
rect 281 -1590 287 -1584
rect 288 -1590 291 -1584
rect 295 -1590 298 -1584
rect 302 -1590 305 -1584
rect 309 -1590 315 -1584
rect 316 -1590 322 -1584
rect 323 -1590 326 -1584
rect 330 -1590 333 -1584
rect 337 -1590 343 -1584
rect 344 -1590 350 -1584
rect 351 -1590 354 -1584
rect 358 -1590 361 -1584
rect 365 -1590 371 -1584
rect 372 -1590 375 -1584
rect 379 -1590 385 -1584
rect 386 -1590 392 -1584
rect 393 -1590 396 -1584
rect 400 -1590 403 -1584
rect 421 -1590 427 -1584
rect 428 -1590 431 -1584
rect 435 -1590 438 -1584
rect 463 -1590 466 -1584
rect 470 -1590 473 -1584
rect 484 -1590 490 -1584
rect 491 -1590 494 -1584
rect 505 -1590 511 -1584
rect 512 -1590 515 -1584
rect 29 -1623 35 -1617
rect 71 -1623 74 -1617
rect 78 -1623 84 -1617
rect 85 -1623 91 -1617
rect 92 -1623 95 -1617
rect 99 -1623 105 -1617
rect 113 -1623 116 -1617
rect 120 -1623 126 -1617
rect 127 -1623 133 -1617
rect 134 -1623 137 -1617
rect 141 -1623 144 -1617
rect 148 -1623 154 -1617
rect 155 -1623 158 -1617
rect 162 -1623 165 -1617
rect 169 -1623 175 -1617
rect 176 -1623 182 -1617
rect 190 -1623 196 -1617
rect 197 -1623 203 -1617
rect 204 -1623 207 -1617
rect 211 -1623 217 -1617
rect 218 -1623 221 -1617
rect 225 -1623 228 -1617
rect 232 -1623 238 -1617
rect 239 -1623 245 -1617
rect 246 -1623 252 -1617
rect 253 -1623 256 -1617
rect 260 -1623 266 -1617
rect 267 -1623 273 -1617
rect 274 -1623 280 -1617
rect 281 -1623 287 -1617
rect 288 -1623 291 -1617
rect 295 -1623 301 -1617
rect 302 -1623 305 -1617
rect 309 -1623 312 -1617
rect 316 -1623 319 -1617
rect 323 -1623 326 -1617
rect 330 -1623 336 -1617
rect 337 -1623 343 -1617
rect 344 -1623 347 -1617
rect 351 -1623 354 -1617
rect 358 -1623 361 -1617
rect 365 -1623 368 -1617
rect 379 -1623 385 -1617
rect 386 -1623 389 -1617
rect 393 -1623 396 -1617
rect 442 -1623 445 -1617
rect 463 -1623 469 -1617
rect 470 -1623 473 -1617
rect 484 -1623 490 -1617
rect 491 -1623 494 -1617
rect 29 -1652 35 -1646
rect 36 -1652 39 -1646
rect 43 -1652 46 -1646
rect 50 -1652 53 -1646
rect 57 -1652 63 -1646
rect 64 -1652 67 -1646
rect 71 -1652 74 -1646
rect 78 -1652 81 -1646
rect 85 -1652 88 -1646
rect 92 -1652 98 -1646
rect 99 -1652 102 -1646
rect 106 -1652 112 -1646
rect 113 -1652 119 -1646
rect 120 -1652 126 -1646
rect 127 -1652 133 -1646
rect 134 -1652 140 -1646
rect 141 -1652 147 -1646
rect 148 -1652 151 -1646
rect 155 -1652 158 -1646
rect 162 -1652 165 -1646
rect 169 -1652 172 -1646
rect 176 -1652 179 -1646
rect 183 -1652 189 -1646
rect 190 -1652 193 -1646
rect 197 -1652 203 -1646
rect 204 -1652 210 -1646
rect 211 -1652 217 -1646
rect 218 -1652 224 -1646
rect 225 -1652 231 -1646
rect 232 -1652 238 -1646
rect 239 -1652 245 -1646
rect 246 -1652 249 -1646
rect 253 -1652 256 -1646
rect 260 -1652 263 -1646
rect 267 -1652 273 -1646
rect 274 -1652 280 -1646
rect 281 -1652 287 -1646
rect 288 -1652 291 -1646
rect 295 -1652 298 -1646
rect 302 -1652 308 -1646
rect 309 -1652 312 -1646
rect 316 -1652 319 -1646
rect 323 -1652 329 -1646
rect 330 -1652 333 -1646
rect 337 -1652 340 -1646
rect 344 -1652 347 -1646
rect 351 -1652 354 -1646
rect 358 -1652 361 -1646
rect 365 -1652 368 -1646
rect 372 -1652 375 -1646
rect 379 -1652 382 -1646
rect 386 -1652 389 -1646
rect 393 -1652 399 -1646
rect 400 -1652 406 -1646
rect 1 -1687 7 -1681
rect 15 -1687 21 -1681
rect 22 -1687 25 -1681
rect 29 -1687 35 -1681
rect 78 -1687 84 -1681
rect 99 -1687 105 -1681
rect 106 -1687 109 -1681
rect 113 -1687 119 -1681
rect 120 -1687 123 -1681
rect 127 -1687 133 -1681
rect 134 -1687 137 -1681
rect 141 -1687 147 -1681
rect 148 -1687 151 -1681
rect 155 -1687 158 -1681
rect 162 -1687 165 -1681
rect 169 -1687 175 -1681
rect 176 -1687 182 -1681
rect 183 -1687 189 -1681
rect 190 -1687 196 -1681
rect 197 -1687 200 -1681
rect 204 -1687 210 -1681
rect 211 -1687 217 -1681
rect 218 -1687 224 -1681
rect 225 -1687 231 -1681
rect 232 -1687 235 -1681
rect 239 -1687 245 -1681
rect 246 -1687 249 -1681
rect 253 -1687 259 -1681
rect 260 -1687 266 -1681
rect 267 -1687 270 -1681
rect 274 -1687 280 -1681
rect 281 -1687 287 -1681
rect 288 -1687 294 -1681
rect 295 -1687 298 -1681
rect 302 -1687 305 -1681
rect 309 -1687 312 -1681
rect 316 -1687 322 -1681
rect 323 -1687 326 -1681
rect 330 -1687 333 -1681
rect 337 -1687 340 -1681
rect 344 -1687 350 -1681
rect 351 -1687 354 -1681
rect 358 -1687 364 -1681
rect 365 -1687 371 -1681
rect 372 -1687 375 -1681
rect 379 -1687 382 -1681
rect 386 -1687 392 -1681
rect 393 -1687 396 -1681
rect 400 -1687 403 -1681
rect 1 -1710 7 -1704
rect 8 -1710 11 -1704
rect 15 -1710 21 -1704
rect 29 -1710 35 -1704
rect 78 -1710 84 -1704
rect 85 -1710 91 -1704
rect 92 -1710 98 -1704
rect 99 -1710 105 -1704
rect 113 -1710 119 -1704
rect 120 -1710 126 -1704
rect 127 -1710 133 -1704
rect 134 -1710 137 -1704
rect 141 -1710 147 -1704
rect 148 -1710 154 -1704
rect 155 -1710 158 -1704
rect 162 -1710 165 -1704
rect 169 -1710 172 -1704
rect 176 -1710 179 -1704
rect 183 -1710 189 -1704
rect 190 -1710 196 -1704
rect 197 -1710 203 -1704
rect 204 -1710 207 -1704
rect 211 -1710 214 -1704
rect 218 -1710 224 -1704
rect 225 -1710 231 -1704
rect 232 -1710 235 -1704
rect 239 -1710 245 -1704
rect 253 -1710 259 -1704
rect 274 -1710 280 -1704
rect 281 -1710 287 -1704
rect 288 -1710 294 -1704
rect 295 -1710 301 -1704
rect 302 -1710 308 -1704
rect 309 -1710 312 -1704
rect 316 -1710 322 -1704
rect 323 -1710 326 -1704
rect 351 -1710 357 -1704
<< polysilicon >>
rect 107 -11 108 -9
rect 110 -11 111 -9
rect 177 -5 178 -3
rect 177 -11 178 -9
rect 187 -5 188 -3
rect 191 -11 192 -9
rect 194 -11 195 -9
rect 198 -5 199 -3
rect 198 -11 199 -9
rect 205 -5 206 -3
rect 208 -5 209 -3
rect 208 -11 209 -9
rect 215 -5 216 -3
rect 215 -11 216 -9
rect 222 -5 223 -3
rect 219 -11 220 -9
rect 226 -11 227 -9
rect 233 -5 234 -3
rect 233 -11 234 -9
rect 240 -5 241 -3
rect 243 -5 244 -3
rect 247 -5 248 -3
rect 247 -11 248 -9
rect 254 -5 255 -3
rect 254 -11 255 -9
rect 275 -5 276 -3
rect 282 -5 283 -3
rect 282 -11 283 -9
rect 289 -5 290 -3
rect 289 -11 290 -9
rect 299 -5 300 -3
rect 299 -11 300 -9
rect 303 -11 304 -9
rect 142 -24 143 -22
rect 142 -30 143 -28
rect 149 -24 150 -22
rect 149 -30 150 -28
rect 159 -24 160 -22
rect 163 -24 164 -22
rect 170 -24 171 -22
rect 177 -30 178 -28
rect 180 -30 181 -28
rect 184 -24 185 -22
rect 184 -30 185 -28
rect 194 -24 195 -22
rect 191 -30 192 -28
rect 198 -24 199 -22
rect 198 -30 199 -28
rect 208 -24 209 -22
rect 212 -30 213 -28
rect 219 -24 220 -22
rect 219 -30 220 -28
rect 240 -24 241 -22
rect 240 -30 241 -28
rect 247 -24 248 -22
rect 257 -30 258 -28
rect 264 -24 265 -22
rect 268 -24 269 -22
rect 268 -30 269 -28
rect 275 -24 276 -22
rect 275 -30 276 -28
rect 285 -30 286 -28
rect 289 -24 290 -22
rect 292 -24 293 -22
rect 289 -30 290 -28
rect 296 -24 297 -22
rect 296 -30 297 -28
rect 303 -30 304 -28
rect 310 -24 311 -22
rect 310 -30 311 -28
rect 320 -30 321 -28
rect 82 -43 83 -41
rect 135 -37 136 -35
rect 135 -43 136 -41
rect 145 -37 146 -35
rect 149 -37 150 -35
rect 152 -37 153 -35
rect 149 -43 150 -41
rect 152 -43 153 -41
rect 156 -37 157 -35
rect 156 -43 157 -41
rect 173 -43 174 -41
rect 184 -37 185 -35
rect 184 -43 185 -41
rect 194 -43 195 -41
rect 212 -43 213 -41
rect 222 -43 223 -41
rect 226 -37 227 -35
rect 229 -43 230 -41
rect 233 -37 234 -35
rect 233 -43 234 -41
rect 243 -37 244 -35
rect 247 -37 248 -35
rect 247 -43 248 -41
rect 250 -43 251 -41
rect 254 -37 255 -35
rect 254 -43 255 -41
rect 261 -37 262 -35
rect 261 -43 262 -41
rect 268 -43 269 -41
rect 275 -37 276 -35
rect 275 -43 276 -41
rect 282 -37 283 -35
rect 282 -43 283 -41
rect 292 -37 293 -35
rect 292 -43 293 -41
rect 296 -37 297 -35
rect 296 -43 297 -41
rect 303 -37 304 -35
rect 310 -43 311 -41
rect 317 -37 318 -35
rect 317 -43 318 -41
rect 324 -37 325 -35
rect 324 -43 325 -41
rect 334 -43 335 -41
rect 478 -37 479 -35
rect 485 -37 486 -35
rect 485 -43 486 -41
rect 579 -37 580 -35
rect 583 -37 584 -35
rect 583 -43 584 -41
rect 79 -60 80 -58
rect 142 -66 143 -64
rect 149 -60 150 -58
rect 149 -66 150 -64
rect 156 -60 157 -58
rect 156 -66 157 -64
rect 170 -60 171 -58
rect 170 -66 171 -64
rect 177 -60 178 -58
rect 177 -66 178 -64
rect 184 -60 185 -58
rect 194 -60 195 -58
rect 198 -66 199 -64
rect 205 -60 206 -58
rect 205 -66 206 -64
rect 212 -60 213 -58
rect 215 -60 216 -58
rect 219 -60 220 -58
rect 219 -66 220 -64
rect 226 -60 227 -58
rect 226 -66 227 -64
rect 233 -60 234 -58
rect 236 -66 237 -64
rect 240 -60 241 -58
rect 243 -60 244 -58
rect 240 -66 241 -64
rect 247 -60 248 -58
rect 247 -66 248 -64
rect 254 -60 255 -58
rect 254 -66 255 -64
rect 261 -60 262 -58
rect 261 -66 262 -64
rect 268 -60 269 -58
rect 268 -66 269 -64
rect 275 -60 276 -58
rect 275 -66 276 -64
rect 282 -60 283 -58
rect 289 -60 290 -58
rect 289 -66 290 -64
rect 296 -60 297 -58
rect 296 -66 297 -64
rect 306 -66 307 -64
rect 310 -66 311 -64
rect 317 -60 318 -58
rect 320 -60 321 -58
rect 320 -66 321 -64
rect 324 -60 325 -58
rect 324 -66 325 -64
rect 338 -60 339 -58
rect 341 -60 342 -58
rect 345 -60 346 -58
rect 345 -66 346 -64
rect 352 -60 353 -58
rect 352 -66 353 -64
rect 362 -60 363 -58
rect 467 -60 468 -58
rect 471 -60 472 -58
rect 471 -66 472 -64
rect 478 -60 479 -58
rect 478 -66 479 -64
rect 576 -60 577 -58
rect 576 -66 577 -64
rect 121 -89 122 -87
rect 138 -83 139 -81
rect 142 -83 143 -81
rect 142 -89 143 -87
rect 149 -83 150 -81
rect 149 -89 150 -87
rect 159 -89 160 -87
rect 163 -83 164 -81
rect 166 -83 167 -81
rect 166 -89 167 -87
rect 170 -83 171 -81
rect 170 -89 171 -87
rect 177 -83 178 -81
rect 177 -89 178 -87
rect 187 -89 188 -87
rect 194 -89 195 -87
rect 198 -83 199 -81
rect 201 -89 202 -87
rect 205 -83 206 -81
rect 205 -89 206 -87
rect 212 -83 213 -81
rect 212 -89 213 -87
rect 219 -83 220 -81
rect 219 -89 220 -87
rect 226 -83 227 -81
rect 226 -89 227 -87
rect 233 -83 234 -81
rect 233 -89 234 -87
rect 240 -83 241 -81
rect 243 -83 244 -81
rect 240 -89 241 -87
rect 243 -89 244 -87
rect 247 -83 248 -81
rect 247 -89 248 -87
rect 254 -83 255 -81
rect 254 -89 255 -87
rect 261 -83 262 -81
rect 261 -89 262 -87
rect 268 -83 269 -81
rect 271 -89 272 -87
rect 275 -83 276 -81
rect 278 -83 279 -81
rect 282 -83 283 -81
rect 282 -89 283 -87
rect 289 -83 290 -81
rect 296 -83 297 -81
rect 296 -89 297 -87
rect 303 -83 304 -81
rect 310 -89 311 -87
rect 317 -83 318 -81
rect 317 -89 318 -87
rect 324 -83 325 -81
rect 324 -89 325 -87
rect 338 -83 339 -81
rect 338 -89 339 -87
rect 345 -83 346 -81
rect 345 -89 346 -87
rect 348 -89 349 -87
rect 352 -83 353 -81
rect 352 -89 353 -87
rect 471 -83 472 -81
rect 474 -83 475 -81
rect 478 -83 479 -81
rect 478 -89 479 -87
rect 485 -83 486 -81
rect 485 -89 486 -87
rect 576 -83 577 -81
rect 576 -89 577 -87
rect 107 -114 108 -112
rect 107 -120 108 -118
rect 121 -114 122 -112
rect 124 -120 125 -118
rect 128 -114 129 -112
rect 135 -114 136 -112
rect 135 -120 136 -118
rect 142 -114 143 -112
rect 145 -114 146 -112
rect 145 -120 146 -118
rect 152 -114 153 -112
rect 156 -114 157 -112
rect 156 -120 157 -118
rect 163 -114 164 -112
rect 163 -120 164 -118
rect 170 -120 171 -118
rect 173 -120 174 -118
rect 180 -114 181 -112
rect 184 -114 185 -112
rect 184 -120 185 -118
rect 191 -114 192 -112
rect 191 -120 192 -118
rect 198 -114 199 -112
rect 198 -120 199 -118
rect 205 -120 206 -118
rect 208 -120 209 -118
rect 212 -114 213 -112
rect 219 -114 220 -112
rect 222 -114 223 -112
rect 219 -120 220 -118
rect 222 -120 223 -118
rect 226 -114 227 -112
rect 226 -120 227 -118
rect 233 -114 234 -112
rect 233 -120 234 -118
rect 243 -114 244 -112
rect 240 -120 241 -118
rect 243 -120 244 -118
rect 250 -114 251 -112
rect 254 -114 255 -112
rect 257 -114 258 -112
rect 257 -120 258 -118
rect 261 -114 262 -112
rect 261 -120 262 -118
rect 268 -114 269 -112
rect 268 -120 269 -118
rect 275 -114 276 -112
rect 275 -120 276 -118
rect 278 -120 279 -118
rect 282 -114 283 -112
rect 282 -120 283 -118
rect 289 -114 290 -112
rect 289 -120 290 -118
rect 296 -114 297 -112
rect 296 -120 297 -118
rect 303 -114 304 -112
rect 303 -120 304 -118
rect 310 -114 311 -112
rect 310 -120 311 -118
rect 317 -114 318 -112
rect 320 -114 321 -112
rect 324 -114 325 -112
rect 324 -120 325 -118
rect 331 -114 332 -112
rect 331 -120 332 -118
rect 338 -114 339 -112
rect 341 -114 342 -112
rect 345 -114 346 -112
rect 345 -120 346 -118
rect 352 -114 353 -112
rect 352 -120 353 -118
rect 359 -114 360 -112
rect 359 -120 360 -118
rect 366 -114 367 -112
rect 366 -120 367 -118
rect 373 -114 374 -112
rect 373 -120 374 -118
rect 380 -114 381 -112
rect 380 -120 381 -118
rect 397 -114 398 -112
rect 394 -120 395 -118
rect 422 -114 423 -112
rect 422 -120 423 -118
rect 478 -114 479 -112
rect 481 -114 482 -112
rect 478 -120 479 -118
rect 485 -114 486 -112
rect 485 -120 486 -118
rect 492 -114 493 -112
rect 492 -120 493 -118
rect 576 -114 577 -112
rect 576 -120 577 -118
rect 583 -114 584 -112
rect 583 -120 584 -118
rect 590 -114 591 -112
rect 590 -120 591 -118
rect 65 -153 66 -151
rect 65 -159 66 -157
rect 72 -153 73 -151
rect 72 -159 73 -157
rect 79 -159 80 -157
rect 86 -153 87 -151
rect 86 -159 87 -157
rect 93 -153 94 -151
rect 93 -159 94 -157
rect 100 -153 101 -151
rect 103 -159 104 -157
rect 107 -153 108 -151
rect 107 -159 108 -157
rect 114 -153 115 -151
rect 114 -159 115 -157
rect 121 -159 122 -157
rect 124 -159 125 -157
rect 128 -153 129 -151
rect 131 -153 132 -151
rect 128 -159 129 -157
rect 131 -159 132 -157
rect 135 -153 136 -151
rect 135 -159 136 -157
rect 142 -159 143 -157
rect 145 -159 146 -157
rect 149 -153 150 -151
rect 149 -159 150 -157
rect 156 -153 157 -151
rect 156 -159 157 -157
rect 163 -159 164 -157
rect 166 -159 167 -157
rect 170 -153 171 -151
rect 170 -159 171 -157
rect 177 -153 178 -151
rect 177 -159 178 -157
rect 184 -153 185 -151
rect 184 -159 185 -157
rect 191 -153 192 -151
rect 191 -159 192 -157
rect 198 -153 199 -151
rect 198 -159 199 -157
rect 205 -153 206 -151
rect 208 -153 209 -151
rect 208 -159 209 -157
rect 212 -153 213 -151
rect 212 -159 213 -157
rect 219 -153 220 -151
rect 222 -153 223 -151
rect 226 -153 227 -151
rect 229 -153 230 -151
rect 226 -159 227 -157
rect 233 -153 234 -151
rect 236 -153 237 -151
rect 233 -159 234 -157
rect 240 -153 241 -151
rect 243 -153 244 -151
rect 240 -159 241 -157
rect 243 -159 244 -157
rect 247 -153 248 -151
rect 247 -159 248 -157
rect 254 -153 255 -151
rect 254 -159 255 -157
rect 261 -153 262 -151
rect 264 -153 265 -151
rect 261 -159 262 -157
rect 264 -159 265 -157
rect 268 -153 269 -151
rect 268 -159 269 -157
rect 275 -153 276 -151
rect 275 -159 276 -157
rect 285 -153 286 -151
rect 289 -153 290 -151
rect 289 -159 290 -157
rect 299 -153 300 -151
rect 299 -159 300 -157
rect 303 -153 304 -151
rect 303 -159 304 -157
rect 310 -153 311 -151
rect 310 -159 311 -157
rect 317 -153 318 -151
rect 317 -159 318 -157
rect 324 -153 325 -151
rect 324 -159 325 -157
rect 334 -153 335 -151
rect 331 -159 332 -157
rect 338 -153 339 -151
rect 338 -159 339 -157
rect 345 -153 346 -151
rect 345 -159 346 -157
rect 352 -153 353 -151
rect 352 -159 353 -157
rect 359 -153 360 -151
rect 359 -159 360 -157
rect 366 -153 367 -151
rect 366 -159 367 -157
rect 373 -153 374 -151
rect 373 -159 374 -157
rect 380 -153 381 -151
rect 380 -159 381 -157
rect 387 -153 388 -151
rect 387 -159 388 -157
rect 394 -153 395 -151
rect 394 -159 395 -157
rect 401 -153 402 -151
rect 401 -159 402 -157
rect 408 -159 409 -157
rect 415 -153 416 -151
rect 415 -159 416 -157
rect 422 -153 423 -151
rect 422 -159 423 -157
rect 429 -153 430 -151
rect 429 -159 430 -157
rect 436 -153 437 -151
rect 436 -159 437 -157
rect 443 -153 444 -151
rect 443 -159 444 -157
rect 499 -153 500 -151
rect 499 -159 500 -157
rect 590 -153 591 -151
rect 590 -159 591 -157
rect 12 -208 13 -206
rect 19 -202 20 -200
rect 26 -202 27 -200
rect 79 -202 80 -200
rect 79 -208 80 -206
rect 86 -202 87 -200
rect 86 -208 87 -206
rect 93 -202 94 -200
rect 100 -202 101 -200
rect 100 -208 101 -206
rect 107 -202 108 -200
rect 107 -208 108 -206
rect 114 -202 115 -200
rect 114 -208 115 -206
rect 121 -202 122 -200
rect 128 -202 129 -200
rect 128 -208 129 -206
rect 135 -202 136 -200
rect 135 -208 136 -206
rect 142 -202 143 -200
rect 145 -208 146 -206
rect 149 -202 150 -200
rect 149 -208 150 -206
rect 156 -202 157 -200
rect 159 -202 160 -200
rect 156 -208 157 -206
rect 163 -202 164 -200
rect 166 -208 167 -206
rect 170 -202 171 -200
rect 173 -208 174 -206
rect 177 -202 178 -200
rect 180 -202 181 -200
rect 184 -208 185 -206
rect 191 -202 192 -200
rect 191 -208 192 -206
rect 198 -208 199 -206
rect 201 -208 202 -206
rect 205 -202 206 -200
rect 205 -208 206 -206
rect 212 -202 213 -200
rect 212 -208 213 -206
rect 215 -208 216 -206
rect 219 -202 220 -200
rect 219 -208 220 -206
rect 222 -208 223 -206
rect 226 -202 227 -200
rect 226 -208 227 -206
rect 236 -202 237 -200
rect 236 -208 237 -206
rect 240 -202 241 -200
rect 243 -202 244 -200
rect 240 -208 241 -206
rect 243 -208 244 -206
rect 247 -202 248 -200
rect 247 -208 248 -206
rect 254 -202 255 -200
rect 254 -208 255 -206
rect 261 -202 262 -200
rect 261 -208 262 -206
rect 268 -202 269 -200
rect 268 -208 269 -206
rect 275 -202 276 -200
rect 278 -202 279 -200
rect 275 -208 276 -206
rect 278 -208 279 -206
rect 282 -202 283 -200
rect 282 -208 283 -206
rect 289 -202 290 -200
rect 292 -208 293 -206
rect 296 -202 297 -200
rect 299 -202 300 -200
rect 296 -208 297 -206
rect 303 -202 304 -200
rect 303 -208 304 -206
rect 310 -202 311 -200
rect 310 -208 311 -206
rect 317 -202 318 -200
rect 320 -202 321 -200
rect 317 -208 318 -206
rect 324 -202 325 -200
rect 324 -208 325 -206
rect 331 -202 332 -200
rect 331 -208 332 -206
rect 338 -202 339 -200
rect 338 -208 339 -206
rect 345 -202 346 -200
rect 345 -208 346 -206
rect 352 -202 353 -200
rect 352 -208 353 -206
rect 359 -202 360 -200
rect 359 -208 360 -206
rect 366 -202 367 -200
rect 366 -208 367 -206
rect 373 -202 374 -200
rect 373 -208 374 -206
rect 380 -202 381 -200
rect 380 -208 381 -206
rect 387 -202 388 -200
rect 387 -208 388 -206
rect 394 -202 395 -200
rect 394 -208 395 -206
rect 401 -202 402 -200
rect 401 -208 402 -206
rect 408 -202 409 -200
rect 408 -208 409 -206
rect 415 -202 416 -200
rect 415 -208 416 -206
rect 422 -202 423 -200
rect 429 -202 430 -200
rect 429 -208 430 -206
rect 436 -202 437 -200
rect 436 -208 437 -206
rect 443 -202 444 -200
rect 443 -208 444 -206
rect 453 -208 454 -206
rect 460 -202 461 -200
rect 464 -202 465 -200
rect 464 -208 465 -206
rect 506 -202 507 -200
rect 506 -208 507 -206
rect 590 -202 591 -200
rect 590 -208 591 -206
rect 12 -243 13 -241
rect 114 -243 115 -241
rect 114 -249 115 -247
rect 124 -249 125 -247
rect 128 -243 129 -241
rect 128 -249 129 -247
rect 135 -243 136 -241
rect 135 -249 136 -247
rect 142 -243 143 -241
rect 142 -249 143 -247
rect 149 -243 150 -241
rect 149 -249 150 -247
rect 156 -243 157 -241
rect 156 -249 157 -247
rect 159 -249 160 -247
rect 163 -243 164 -241
rect 163 -249 164 -247
rect 170 -249 171 -247
rect 177 -243 178 -241
rect 177 -249 178 -247
rect 184 -243 185 -241
rect 184 -249 185 -247
rect 191 -243 192 -241
rect 191 -249 192 -247
rect 198 -243 199 -241
rect 198 -249 199 -247
rect 208 -249 209 -247
rect 212 -243 213 -241
rect 215 -243 216 -241
rect 222 -243 223 -241
rect 219 -249 220 -247
rect 222 -249 223 -247
rect 226 -243 227 -241
rect 229 -249 230 -247
rect 236 -243 237 -241
rect 236 -249 237 -247
rect 240 -243 241 -241
rect 243 -243 244 -241
rect 240 -249 241 -247
rect 243 -249 244 -247
rect 247 -243 248 -241
rect 247 -249 248 -247
rect 254 -243 255 -241
rect 254 -249 255 -247
rect 261 -243 262 -241
rect 264 -243 265 -241
rect 268 -243 269 -241
rect 268 -249 269 -247
rect 275 -243 276 -241
rect 278 -243 279 -241
rect 275 -249 276 -247
rect 278 -249 279 -247
rect 282 -243 283 -241
rect 282 -249 283 -247
rect 289 -243 290 -241
rect 292 -243 293 -241
rect 296 -243 297 -241
rect 303 -243 304 -241
rect 303 -249 304 -247
rect 310 -243 311 -241
rect 310 -249 311 -247
rect 317 -243 318 -241
rect 320 -243 321 -241
rect 317 -249 318 -247
rect 320 -249 321 -247
rect 324 -243 325 -241
rect 324 -249 325 -247
rect 331 -243 332 -241
rect 331 -249 332 -247
rect 338 -243 339 -241
rect 338 -249 339 -247
rect 345 -243 346 -241
rect 348 -243 349 -241
rect 348 -249 349 -247
rect 352 -243 353 -241
rect 352 -249 353 -247
rect 359 -243 360 -241
rect 359 -249 360 -247
rect 366 -243 367 -241
rect 366 -249 367 -247
rect 373 -243 374 -241
rect 373 -249 374 -247
rect 383 -243 384 -241
rect 380 -249 381 -247
rect 387 -243 388 -241
rect 387 -249 388 -247
rect 394 -243 395 -241
rect 394 -249 395 -247
rect 401 -243 402 -241
rect 401 -249 402 -247
rect 408 -243 409 -241
rect 408 -249 409 -247
rect 415 -243 416 -241
rect 415 -249 416 -247
rect 422 -243 423 -241
rect 422 -249 423 -247
rect 429 -243 430 -241
rect 429 -249 430 -247
rect 436 -243 437 -241
rect 436 -249 437 -247
rect 443 -243 444 -241
rect 443 -249 444 -247
rect 450 -243 451 -241
rect 450 -249 451 -247
rect 460 -243 461 -241
rect 464 -249 465 -247
rect 509 -243 510 -241
rect 506 -249 507 -247
rect 562 -243 563 -241
rect 562 -249 563 -247
rect 572 -243 573 -241
rect 590 -243 591 -241
rect 590 -249 591 -247
rect 597 -249 598 -247
rect 600 -249 601 -247
rect 646 -249 647 -247
rect 65 -284 66 -282
rect 75 -290 76 -288
rect 79 -284 80 -282
rect 79 -290 80 -288
rect 86 -284 87 -282
rect 86 -290 87 -288
rect 93 -284 94 -282
rect 93 -290 94 -288
rect 103 -290 104 -288
rect 107 -284 108 -282
rect 107 -290 108 -288
rect 114 -284 115 -282
rect 117 -290 118 -288
rect 121 -284 122 -282
rect 128 -284 129 -282
rect 128 -290 129 -288
rect 135 -284 136 -282
rect 135 -290 136 -288
rect 142 -284 143 -282
rect 142 -290 143 -288
rect 149 -284 150 -282
rect 149 -290 150 -288
rect 156 -284 157 -282
rect 156 -290 157 -288
rect 163 -284 164 -282
rect 163 -290 164 -288
rect 170 -284 171 -282
rect 173 -284 174 -282
rect 173 -290 174 -288
rect 177 -284 178 -282
rect 177 -290 178 -288
rect 184 -284 185 -282
rect 187 -284 188 -282
rect 187 -290 188 -288
rect 194 -284 195 -282
rect 194 -290 195 -288
rect 201 -284 202 -282
rect 198 -290 199 -288
rect 205 -284 206 -282
rect 208 -284 209 -282
rect 212 -290 213 -288
rect 219 -284 220 -282
rect 219 -290 220 -288
rect 226 -284 227 -282
rect 226 -290 227 -288
rect 233 -284 234 -282
rect 236 -284 237 -282
rect 236 -290 237 -288
rect 243 -284 244 -282
rect 240 -290 241 -288
rect 247 -284 248 -282
rect 247 -290 248 -288
rect 257 -284 258 -282
rect 254 -290 255 -288
rect 257 -290 258 -288
rect 261 -284 262 -282
rect 261 -290 262 -288
rect 268 -284 269 -282
rect 268 -290 269 -288
rect 275 -284 276 -282
rect 275 -290 276 -288
rect 282 -290 283 -288
rect 289 -284 290 -282
rect 292 -284 293 -282
rect 289 -290 290 -288
rect 296 -284 297 -282
rect 299 -284 300 -282
rect 303 -284 304 -282
rect 303 -290 304 -288
rect 313 -284 314 -282
rect 317 -284 318 -282
rect 320 -284 321 -282
rect 320 -290 321 -288
rect 324 -284 325 -282
rect 327 -284 328 -282
rect 324 -290 325 -288
rect 331 -284 332 -282
rect 331 -290 332 -288
rect 338 -284 339 -282
rect 341 -290 342 -288
rect 345 -284 346 -282
rect 345 -290 346 -288
rect 352 -284 353 -282
rect 352 -290 353 -288
rect 359 -284 360 -282
rect 359 -290 360 -288
rect 366 -284 367 -282
rect 366 -290 367 -288
rect 373 -284 374 -282
rect 373 -290 374 -288
rect 383 -284 384 -282
rect 387 -284 388 -282
rect 387 -290 388 -288
rect 394 -290 395 -288
rect 401 -284 402 -282
rect 401 -290 402 -288
rect 408 -284 409 -282
rect 408 -290 409 -288
rect 415 -284 416 -282
rect 415 -290 416 -288
rect 422 -284 423 -282
rect 422 -290 423 -288
rect 429 -284 430 -282
rect 429 -290 430 -288
rect 436 -284 437 -282
rect 436 -290 437 -288
rect 443 -284 444 -282
rect 443 -290 444 -288
rect 450 -284 451 -282
rect 450 -290 451 -288
rect 457 -284 458 -282
rect 457 -290 458 -288
rect 464 -284 465 -282
rect 464 -290 465 -288
rect 471 -284 472 -282
rect 471 -290 472 -288
rect 478 -284 479 -282
rect 478 -290 479 -288
rect 485 -284 486 -282
rect 485 -290 486 -288
rect 492 -284 493 -282
rect 492 -290 493 -288
rect 499 -284 500 -282
rect 502 -284 503 -282
rect 506 -284 507 -282
rect 506 -290 507 -288
rect 520 -284 521 -282
rect 520 -290 521 -288
rect 527 -284 528 -282
rect 527 -290 528 -288
rect 562 -284 563 -282
rect 562 -290 563 -288
rect 611 -284 612 -282
rect 611 -290 612 -288
rect 646 -284 647 -282
rect 646 -290 647 -288
rect 72 -339 73 -337
rect 79 -333 80 -331
rect 79 -339 80 -337
rect 86 -333 87 -331
rect 86 -339 87 -337
rect 93 -333 94 -331
rect 93 -339 94 -337
rect 100 -333 101 -331
rect 100 -339 101 -337
rect 107 -333 108 -331
rect 107 -339 108 -337
rect 114 -333 115 -331
rect 114 -339 115 -337
rect 121 -333 122 -331
rect 121 -339 122 -337
rect 128 -333 129 -331
rect 128 -339 129 -337
rect 135 -333 136 -331
rect 135 -339 136 -337
rect 142 -333 143 -331
rect 142 -339 143 -337
rect 152 -333 153 -331
rect 152 -339 153 -337
rect 156 -339 157 -337
rect 163 -333 164 -331
rect 163 -339 164 -337
rect 170 -333 171 -331
rect 170 -339 171 -337
rect 177 -333 178 -331
rect 177 -339 178 -337
rect 184 -339 185 -337
rect 191 -333 192 -331
rect 191 -339 192 -337
rect 198 -333 199 -331
rect 198 -339 199 -337
rect 205 -333 206 -331
rect 205 -339 206 -337
rect 212 -333 213 -331
rect 212 -339 213 -337
rect 219 -333 220 -331
rect 219 -339 220 -337
rect 226 -333 227 -331
rect 229 -333 230 -331
rect 226 -339 227 -337
rect 233 -333 234 -331
rect 233 -339 234 -337
rect 236 -339 237 -337
rect 240 -333 241 -331
rect 240 -339 241 -337
rect 247 -333 248 -331
rect 247 -339 248 -337
rect 254 -333 255 -331
rect 254 -339 255 -337
rect 264 -333 265 -331
rect 264 -339 265 -337
rect 271 -339 272 -337
rect 275 -333 276 -331
rect 275 -339 276 -337
rect 282 -333 283 -331
rect 285 -339 286 -337
rect 289 -333 290 -331
rect 289 -339 290 -337
rect 296 -333 297 -331
rect 296 -339 297 -337
rect 303 -333 304 -331
rect 303 -339 304 -337
rect 313 -333 314 -331
rect 313 -339 314 -337
rect 317 -333 318 -331
rect 317 -339 318 -337
rect 324 -333 325 -331
rect 324 -339 325 -337
rect 327 -339 328 -337
rect 331 -333 332 -331
rect 331 -339 332 -337
rect 338 -333 339 -331
rect 341 -339 342 -337
rect 345 -333 346 -331
rect 348 -333 349 -331
rect 348 -339 349 -337
rect 352 -333 353 -331
rect 352 -339 353 -337
rect 359 -333 360 -331
rect 359 -339 360 -337
rect 362 -339 363 -337
rect 366 -333 367 -331
rect 369 -333 370 -331
rect 366 -339 367 -337
rect 373 -333 374 -331
rect 373 -339 374 -337
rect 380 -333 381 -331
rect 380 -339 381 -337
rect 387 -333 388 -331
rect 390 -333 391 -331
rect 394 -333 395 -331
rect 394 -339 395 -337
rect 401 -333 402 -331
rect 401 -339 402 -337
rect 408 -333 409 -331
rect 411 -339 412 -337
rect 415 -333 416 -331
rect 415 -339 416 -337
rect 422 -333 423 -331
rect 425 -333 426 -331
rect 422 -339 423 -337
rect 429 -333 430 -331
rect 429 -339 430 -337
rect 436 -333 437 -331
rect 436 -339 437 -337
rect 443 -333 444 -331
rect 443 -339 444 -337
rect 450 -333 451 -331
rect 450 -339 451 -337
rect 457 -333 458 -331
rect 457 -339 458 -337
rect 464 -333 465 -331
rect 464 -339 465 -337
rect 471 -333 472 -331
rect 471 -339 472 -337
rect 478 -333 479 -331
rect 478 -339 479 -337
rect 485 -333 486 -331
rect 485 -339 486 -337
rect 492 -333 493 -331
rect 492 -339 493 -337
rect 499 -333 500 -331
rect 499 -339 500 -337
rect 506 -333 507 -331
rect 506 -339 507 -337
rect 516 -333 517 -331
rect 520 -333 521 -331
rect 520 -339 521 -337
rect 527 -333 528 -331
rect 527 -339 528 -337
rect 534 -333 535 -331
rect 534 -339 535 -337
rect 541 -333 542 -331
rect 544 -333 545 -331
rect 541 -339 542 -337
rect 544 -339 545 -337
rect 548 -333 549 -331
rect 548 -339 549 -337
rect 555 -333 556 -331
rect 558 -339 559 -337
rect 562 -333 563 -331
rect 562 -339 563 -337
rect 604 -333 605 -331
rect 604 -339 605 -337
rect 649 -333 650 -331
rect 649 -339 650 -337
rect 653 -333 654 -331
rect 653 -339 654 -337
rect 660 -333 661 -331
rect 660 -339 661 -337
rect 674 -333 675 -331
rect 674 -339 675 -337
rect 681 -333 682 -331
rect 30 -390 31 -388
rect 44 -384 45 -382
rect 44 -390 45 -388
rect 51 -384 52 -382
rect 51 -390 52 -388
rect 58 -384 59 -382
rect 58 -390 59 -388
rect 68 -384 69 -382
rect 72 -384 73 -382
rect 72 -390 73 -388
rect 79 -384 80 -382
rect 79 -390 80 -388
rect 86 -384 87 -382
rect 86 -390 87 -388
rect 93 -384 94 -382
rect 93 -390 94 -388
rect 100 -384 101 -382
rect 100 -390 101 -388
rect 107 -384 108 -382
rect 110 -384 111 -382
rect 114 -384 115 -382
rect 114 -390 115 -388
rect 121 -384 122 -382
rect 121 -390 122 -388
rect 128 -384 129 -382
rect 128 -390 129 -388
rect 135 -384 136 -382
rect 138 -384 139 -382
rect 138 -390 139 -388
rect 142 -384 143 -382
rect 142 -390 143 -388
rect 152 -384 153 -382
rect 152 -390 153 -388
rect 156 -384 157 -382
rect 159 -384 160 -382
rect 159 -390 160 -388
rect 166 -384 167 -382
rect 166 -390 167 -388
rect 170 -384 171 -382
rect 170 -390 171 -388
rect 177 -384 178 -382
rect 177 -390 178 -388
rect 184 -384 185 -382
rect 184 -390 185 -388
rect 191 -384 192 -382
rect 191 -390 192 -388
rect 198 -384 199 -382
rect 198 -390 199 -388
rect 205 -384 206 -382
rect 205 -390 206 -388
rect 215 -384 216 -382
rect 212 -390 213 -388
rect 215 -390 216 -388
rect 219 -384 220 -382
rect 222 -384 223 -382
rect 222 -390 223 -388
rect 229 -384 230 -382
rect 233 -384 234 -382
rect 236 -384 237 -382
rect 236 -390 237 -388
rect 240 -384 241 -382
rect 243 -384 244 -382
rect 240 -390 241 -388
rect 247 -384 248 -382
rect 247 -390 248 -388
rect 254 -384 255 -382
rect 254 -390 255 -388
rect 261 -384 262 -382
rect 261 -390 262 -388
rect 268 -384 269 -382
rect 268 -390 269 -388
rect 278 -390 279 -388
rect 282 -384 283 -382
rect 282 -390 283 -388
rect 292 -384 293 -382
rect 289 -390 290 -388
rect 292 -390 293 -388
rect 296 -384 297 -382
rect 296 -390 297 -388
rect 303 -384 304 -382
rect 303 -390 304 -388
rect 310 -384 311 -382
rect 310 -390 311 -388
rect 317 -384 318 -382
rect 317 -390 318 -388
rect 324 -384 325 -382
rect 327 -384 328 -382
rect 324 -390 325 -388
rect 331 -384 332 -382
rect 334 -384 335 -382
rect 334 -390 335 -388
rect 338 -384 339 -382
rect 341 -384 342 -382
rect 341 -390 342 -388
rect 345 -384 346 -382
rect 345 -390 346 -388
rect 352 -390 353 -388
rect 355 -390 356 -388
rect 362 -384 363 -382
rect 359 -390 360 -388
rect 366 -384 367 -382
rect 366 -390 367 -388
rect 373 -384 374 -382
rect 373 -390 374 -388
rect 380 -384 381 -382
rect 380 -390 381 -388
rect 387 -384 388 -382
rect 390 -384 391 -382
rect 387 -390 388 -388
rect 394 -384 395 -382
rect 394 -390 395 -388
rect 401 -384 402 -382
rect 401 -390 402 -388
rect 408 -384 409 -382
rect 408 -390 409 -388
rect 415 -384 416 -382
rect 415 -390 416 -388
rect 422 -384 423 -382
rect 425 -384 426 -382
rect 429 -384 430 -382
rect 429 -390 430 -388
rect 436 -384 437 -382
rect 436 -390 437 -388
rect 443 -384 444 -382
rect 443 -390 444 -388
rect 450 -384 451 -382
rect 450 -390 451 -388
rect 460 -384 461 -382
rect 460 -390 461 -388
rect 464 -384 465 -382
rect 464 -390 465 -388
rect 471 -384 472 -382
rect 471 -390 472 -388
rect 478 -384 479 -382
rect 478 -390 479 -388
rect 485 -384 486 -382
rect 485 -390 486 -388
rect 492 -384 493 -382
rect 492 -390 493 -388
rect 499 -384 500 -382
rect 499 -390 500 -388
rect 506 -384 507 -382
rect 506 -390 507 -388
rect 513 -384 514 -382
rect 513 -390 514 -388
rect 523 -384 524 -382
rect 527 -384 528 -382
rect 527 -390 528 -388
rect 534 -384 535 -382
rect 534 -390 535 -388
rect 541 -384 542 -382
rect 541 -390 542 -388
rect 548 -384 549 -382
rect 548 -390 549 -388
rect 555 -384 556 -382
rect 555 -390 556 -388
rect 562 -384 563 -382
rect 569 -384 570 -382
rect 569 -390 570 -388
rect 576 -384 577 -382
rect 576 -390 577 -388
rect 583 -384 584 -382
rect 583 -390 584 -388
rect 590 -384 591 -382
rect 590 -390 591 -388
rect 597 -384 598 -382
rect 597 -390 598 -388
rect 604 -384 605 -382
rect 604 -390 605 -388
rect 611 -384 612 -382
rect 611 -390 612 -388
rect 618 -384 619 -382
rect 618 -390 619 -388
rect 625 -384 626 -382
rect 625 -390 626 -388
rect 632 -384 633 -382
rect 632 -390 633 -388
rect 639 -384 640 -382
rect 642 -384 643 -382
rect 646 -384 647 -382
rect 646 -390 647 -388
rect 653 -384 654 -382
rect 653 -390 654 -388
rect 660 -384 661 -382
rect 667 -384 668 -382
rect 667 -390 668 -388
rect 674 -390 675 -388
rect 681 -384 682 -382
rect 681 -390 682 -388
rect 688 -384 689 -382
rect 688 -390 689 -388
rect 2 -441 3 -439
rect 2 -447 3 -445
rect 9 -447 10 -445
rect 16 -441 17 -439
rect 16 -447 17 -445
rect 23 -441 24 -439
rect 23 -447 24 -445
rect 33 -447 34 -445
rect 37 -441 38 -439
rect 37 -447 38 -445
rect 44 -441 45 -439
rect 44 -447 45 -445
rect 51 -441 52 -439
rect 51 -447 52 -445
rect 58 -441 59 -439
rect 58 -447 59 -445
rect 65 -441 66 -439
rect 65 -447 66 -445
rect 72 -441 73 -439
rect 72 -447 73 -445
rect 79 -441 80 -439
rect 79 -447 80 -445
rect 86 -441 87 -439
rect 86 -447 87 -445
rect 93 -441 94 -439
rect 93 -447 94 -445
rect 100 -441 101 -439
rect 100 -447 101 -445
rect 107 -441 108 -439
rect 107 -447 108 -445
rect 114 -441 115 -439
rect 114 -447 115 -445
rect 121 -441 122 -439
rect 121 -447 122 -445
rect 128 -441 129 -439
rect 128 -447 129 -445
rect 135 -441 136 -439
rect 138 -447 139 -445
rect 145 -441 146 -439
rect 142 -447 143 -445
rect 145 -447 146 -445
rect 149 -441 150 -439
rect 149 -447 150 -445
rect 159 -441 160 -439
rect 159 -447 160 -445
rect 163 -441 164 -439
rect 163 -447 164 -445
rect 170 -441 171 -439
rect 170 -447 171 -445
rect 177 -441 178 -439
rect 180 -441 181 -439
rect 177 -447 178 -445
rect 180 -447 181 -445
rect 184 -441 185 -439
rect 187 -441 188 -439
rect 184 -447 185 -445
rect 187 -447 188 -445
rect 191 -441 192 -439
rect 191 -447 192 -445
rect 198 -441 199 -439
rect 198 -447 199 -445
rect 205 -441 206 -439
rect 205 -447 206 -445
rect 215 -441 216 -439
rect 215 -447 216 -445
rect 219 -441 220 -439
rect 219 -447 220 -445
rect 226 -441 227 -439
rect 226 -447 227 -445
rect 233 -441 234 -439
rect 236 -441 237 -439
rect 233 -447 234 -445
rect 236 -447 237 -445
rect 240 -441 241 -439
rect 243 -447 244 -445
rect 247 -441 248 -439
rect 247 -447 248 -445
rect 254 -441 255 -439
rect 254 -447 255 -445
rect 261 -441 262 -439
rect 261 -447 262 -445
rect 268 -441 269 -439
rect 268 -447 269 -445
rect 275 -441 276 -439
rect 275 -447 276 -445
rect 282 -441 283 -439
rect 285 -441 286 -439
rect 282 -447 283 -445
rect 285 -447 286 -445
rect 289 -441 290 -439
rect 289 -447 290 -445
rect 292 -447 293 -445
rect 296 -441 297 -439
rect 296 -447 297 -445
rect 303 -441 304 -439
rect 310 -441 311 -439
rect 310 -447 311 -445
rect 317 -441 318 -439
rect 317 -447 318 -445
rect 324 -441 325 -439
rect 327 -441 328 -439
rect 331 -441 332 -439
rect 331 -447 332 -445
rect 338 -441 339 -439
rect 341 -441 342 -439
rect 345 -441 346 -439
rect 345 -447 346 -445
rect 352 -441 353 -439
rect 352 -447 353 -445
rect 359 -441 360 -439
rect 359 -447 360 -445
rect 369 -441 370 -439
rect 366 -447 367 -445
rect 369 -447 370 -445
rect 373 -441 374 -439
rect 376 -441 377 -439
rect 373 -447 374 -445
rect 376 -447 377 -445
rect 380 -441 381 -439
rect 380 -447 381 -445
rect 387 -441 388 -439
rect 387 -447 388 -445
rect 397 -441 398 -439
rect 397 -447 398 -445
rect 401 -441 402 -439
rect 404 -441 405 -439
rect 404 -447 405 -445
rect 408 -441 409 -439
rect 415 -441 416 -439
rect 415 -447 416 -445
rect 422 -441 423 -439
rect 422 -447 423 -445
rect 429 -441 430 -439
rect 429 -447 430 -445
rect 436 -441 437 -439
rect 439 -441 440 -439
rect 436 -447 437 -445
rect 443 -441 444 -439
rect 443 -447 444 -445
rect 450 -441 451 -439
rect 450 -447 451 -445
rect 457 -441 458 -439
rect 457 -447 458 -445
rect 467 -441 468 -439
rect 464 -447 465 -445
rect 471 -441 472 -439
rect 471 -447 472 -445
rect 478 -441 479 -439
rect 478 -447 479 -445
rect 485 -441 486 -439
rect 485 -447 486 -445
rect 492 -441 493 -439
rect 492 -447 493 -445
rect 499 -441 500 -439
rect 499 -447 500 -445
rect 509 -447 510 -445
rect 513 -441 514 -439
rect 513 -447 514 -445
rect 520 -441 521 -439
rect 520 -447 521 -445
rect 527 -441 528 -439
rect 527 -447 528 -445
rect 534 -441 535 -439
rect 534 -447 535 -445
rect 541 -441 542 -439
rect 541 -447 542 -445
rect 548 -441 549 -439
rect 548 -447 549 -445
rect 558 -441 559 -439
rect 558 -447 559 -445
rect 562 -441 563 -439
rect 562 -447 563 -445
rect 569 -441 570 -439
rect 569 -447 570 -445
rect 576 -441 577 -439
rect 576 -447 577 -445
rect 583 -441 584 -439
rect 583 -447 584 -445
rect 590 -441 591 -439
rect 590 -447 591 -445
rect 597 -441 598 -439
rect 597 -447 598 -445
rect 604 -441 605 -439
rect 604 -447 605 -445
rect 611 -441 612 -439
rect 611 -447 612 -445
rect 618 -441 619 -439
rect 618 -447 619 -445
rect 625 -441 626 -439
rect 628 -441 629 -439
rect 625 -447 626 -445
rect 632 -441 633 -439
rect 632 -447 633 -445
rect 635 -447 636 -445
rect 639 -441 640 -439
rect 639 -447 640 -445
rect 649 -441 650 -439
rect 646 -447 647 -445
rect 653 -441 654 -439
rect 653 -447 654 -445
rect 663 -441 664 -439
rect 663 -447 664 -445
rect 667 -441 668 -439
rect 667 -447 668 -445
rect 9 -498 10 -496
rect 9 -504 10 -502
rect 16 -498 17 -496
rect 16 -504 17 -502
rect 23 -498 24 -496
rect 23 -504 24 -502
rect 30 -498 31 -496
rect 30 -504 31 -502
rect 37 -498 38 -496
rect 37 -504 38 -502
rect 44 -498 45 -496
rect 44 -504 45 -502
rect 51 -498 52 -496
rect 51 -504 52 -502
rect 58 -498 59 -496
rect 65 -498 66 -496
rect 68 -504 69 -502
rect 72 -498 73 -496
rect 72 -504 73 -502
rect 79 -498 80 -496
rect 79 -504 80 -502
rect 86 -498 87 -496
rect 86 -504 87 -502
rect 93 -504 94 -502
rect 100 -498 101 -496
rect 100 -504 101 -502
rect 107 -498 108 -496
rect 110 -498 111 -496
rect 107 -504 108 -502
rect 114 -498 115 -496
rect 121 -498 122 -496
rect 121 -504 122 -502
rect 128 -498 129 -496
rect 131 -498 132 -496
rect 138 -498 139 -496
rect 135 -504 136 -502
rect 142 -498 143 -496
rect 142 -504 143 -502
rect 149 -504 150 -502
rect 152 -504 153 -502
rect 156 -498 157 -496
rect 156 -504 157 -502
rect 159 -504 160 -502
rect 163 -498 164 -496
rect 166 -498 167 -496
rect 163 -504 164 -502
rect 170 -498 171 -496
rect 170 -504 171 -502
rect 177 -498 178 -496
rect 177 -504 178 -502
rect 184 -498 185 -496
rect 184 -504 185 -502
rect 191 -498 192 -496
rect 191 -504 192 -502
rect 201 -498 202 -496
rect 198 -504 199 -502
rect 208 -498 209 -496
rect 205 -504 206 -502
rect 208 -504 209 -502
rect 212 -498 213 -496
rect 215 -498 216 -496
rect 212 -504 213 -502
rect 215 -504 216 -502
rect 219 -498 220 -496
rect 219 -504 220 -502
rect 226 -498 227 -496
rect 226 -504 227 -502
rect 233 -498 234 -496
rect 233 -504 234 -502
rect 243 -498 244 -496
rect 240 -504 241 -502
rect 243 -504 244 -502
rect 247 -498 248 -496
rect 247 -504 248 -502
rect 254 -498 255 -496
rect 254 -504 255 -502
rect 264 -498 265 -496
rect 271 -504 272 -502
rect 275 -498 276 -496
rect 275 -504 276 -502
rect 282 -498 283 -496
rect 282 -504 283 -502
rect 289 -498 290 -496
rect 289 -504 290 -502
rect 296 -498 297 -496
rect 296 -504 297 -502
rect 303 -498 304 -496
rect 303 -504 304 -502
rect 310 -498 311 -496
rect 310 -504 311 -502
rect 317 -498 318 -496
rect 317 -504 318 -502
rect 324 -498 325 -496
rect 324 -504 325 -502
rect 331 -504 332 -502
rect 338 -498 339 -496
rect 338 -504 339 -502
rect 345 -498 346 -496
rect 345 -504 346 -502
rect 352 -498 353 -496
rect 355 -498 356 -496
rect 355 -504 356 -502
rect 359 -498 360 -496
rect 359 -504 360 -502
rect 366 -498 367 -496
rect 369 -504 370 -502
rect 373 -498 374 -496
rect 373 -504 374 -502
rect 380 -498 381 -496
rect 383 -504 384 -502
rect 387 -498 388 -496
rect 390 -498 391 -496
rect 390 -504 391 -502
rect 397 -498 398 -496
rect 394 -504 395 -502
rect 397 -504 398 -502
rect 401 -498 402 -496
rect 401 -504 402 -502
rect 408 -498 409 -496
rect 408 -504 409 -502
rect 415 -498 416 -496
rect 418 -498 419 -496
rect 415 -504 416 -502
rect 422 -498 423 -496
rect 422 -504 423 -502
rect 429 -498 430 -496
rect 429 -504 430 -502
rect 436 -498 437 -496
rect 436 -504 437 -502
rect 443 -498 444 -496
rect 443 -504 444 -502
rect 450 -498 451 -496
rect 450 -504 451 -502
rect 457 -498 458 -496
rect 457 -504 458 -502
rect 464 -498 465 -496
rect 464 -504 465 -502
rect 471 -498 472 -496
rect 471 -504 472 -502
rect 478 -504 479 -502
rect 485 -498 486 -496
rect 485 -504 486 -502
rect 492 -498 493 -496
rect 492 -504 493 -502
rect 499 -498 500 -496
rect 499 -504 500 -502
rect 509 -498 510 -496
rect 513 -498 514 -496
rect 513 -504 514 -502
rect 520 -498 521 -496
rect 520 -504 521 -502
rect 527 -498 528 -496
rect 527 -504 528 -502
rect 534 -498 535 -496
rect 534 -504 535 -502
rect 541 -498 542 -496
rect 541 -504 542 -502
rect 548 -498 549 -496
rect 548 -504 549 -502
rect 555 -498 556 -496
rect 555 -504 556 -502
rect 562 -498 563 -496
rect 562 -504 563 -502
rect 569 -498 570 -496
rect 569 -504 570 -502
rect 576 -498 577 -496
rect 576 -504 577 -502
rect 583 -498 584 -496
rect 583 -504 584 -502
rect 590 -504 591 -502
rect 597 -498 598 -496
rect 597 -504 598 -502
rect 604 -504 605 -502
rect 614 -498 615 -496
rect 611 -504 612 -502
rect 614 -504 615 -502
rect 618 -498 619 -496
rect 618 -504 619 -502
rect 625 -504 626 -502
rect 628 -504 629 -502
rect 632 -498 633 -496
rect 632 -504 633 -502
rect 639 -498 640 -496
rect 639 -504 640 -502
rect 646 -498 647 -496
rect 646 -504 647 -502
rect 653 -498 654 -496
rect 653 -504 654 -502
rect 660 -498 661 -496
rect 660 -504 661 -502
rect 670 -504 671 -502
rect 5 -555 6 -553
rect 9 -555 10 -553
rect 9 -561 10 -559
rect 16 -555 17 -553
rect 16 -561 17 -559
rect 23 -555 24 -553
rect 23 -561 24 -559
rect 30 -555 31 -553
rect 30 -561 31 -559
rect 37 -555 38 -553
rect 37 -561 38 -559
rect 44 -555 45 -553
rect 44 -561 45 -559
rect 51 -555 52 -553
rect 51 -561 52 -559
rect 58 -555 59 -553
rect 61 -555 62 -553
rect 65 -555 66 -553
rect 65 -561 66 -559
rect 72 -555 73 -553
rect 72 -561 73 -559
rect 75 -561 76 -559
rect 82 -555 83 -553
rect 82 -561 83 -559
rect 86 -555 87 -553
rect 93 -555 94 -553
rect 93 -561 94 -559
rect 100 -555 101 -553
rect 100 -561 101 -559
rect 107 -555 108 -553
rect 107 -561 108 -559
rect 114 -555 115 -553
rect 117 -555 118 -553
rect 114 -561 115 -559
rect 117 -561 118 -559
rect 121 -555 122 -553
rect 121 -561 122 -559
rect 128 -555 129 -553
rect 131 -555 132 -553
rect 128 -561 129 -559
rect 131 -561 132 -559
rect 135 -555 136 -553
rect 135 -561 136 -559
rect 142 -561 143 -559
rect 149 -555 150 -553
rect 149 -561 150 -559
rect 156 -555 157 -553
rect 156 -561 157 -559
rect 163 -555 164 -553
rect 163 -561 164 -559
rect 170 -555 171 -553
rect 170 -561 171 -559
rect 180 -555 181 -553
rect 177 -561 178 -559
rect 180 -561 181 -559
rect 184 -555 185 -553
rect 184 -561 185 -559
rect 194 -561 195 -559
rect 198 -555 199 -553
rect 198 -561 199 -559
rect 205 -555 206 -553
rect 208 -555 209 -553
rect 205 -561 206 -559
rect 212 -555 213 -553
rect 212 -561 213 -559
rect 219 -555 220 -553
rect 219 -561 220 -559
rect 226 -555 227 -553
rect 226 -561 227 -559
rect 233 -555 234 -553
rect 233 -561 234 -559
rect 240 -555 241 -553
rect 243 -555 244 -553
rect 243 -561 244 -559
rect 247 -555 248 -553
rect 247 -561 248 -559
rect 254 -555 255 -553
rect 254 -561 255 -559
rect 261 -555 262 -553
rect 261 -561 262 -559
rect 268 -555 269 -553
rect 268 -561 269 -559
rect 275 -555 276 -553
rect 278 -555 279 -553
rect 278 -561 279 -559
rect 285 -555 286 -553
rect 282 -561 283 -559
rect 285 -561 286 -559
rect 292 -555 293 -553
rect 289 -561 290 -559
rect 292 -561 293 -559
rect 296 -555 297 -553
rect 296 -561 297 -559
rect 303 -555 304 -553
rect 303 -561 304 -559
rect 310 -555 311 -553
rect 313 -555 314 -553
rect 310 -561 311 -559
rect 313 -561 314 -559
rect 317 -555 318 -553
rect 317 -561 318 -559
rect 320 -561 321 -559
rect 324 -555 325 -553
rect 324 -561 325 -559
rect 331 -555 332 -553
rect 331 -561 332 -559
rect 341 -555 342 -553
rect 341 -561 342 -559
rect 345 -555 346 -553
rect 348 -555 349 -553
rect 345 -561 346 -559
rect 355 -555 356 -553
rect 352 -561 353 -559
rect 355 -561 356 -559
rect 362 -555 363 -553
rect 359 -561 360 -559
rect 366 -555 367 -553
rect 366 -561 367 -559
rect 376 -555 377 -553
rect 373 -561 374 -559
rect 376 -561 377 -559
rect 380 -555 381 -553
rect 380 -561 381 -559
rect 387 -555 388 -553
rect 387 -561 388 -559
rect 394 -555 395 -553
rect 394 -561 395 -559
rect 401 -555 402 -553
rect 401 -561 402 -559
rect 404 -561 405 -559
rect 408 -555 409 -553
rect 408 -561 409 -559
rect 415 -555 416 -553
rect 415 -561 416 -559
rect 425 -561 426 -559
rect 429 -555 430 -553
rect 429 -561 430 -559
rect 436 -555 437 -553
rect 436 -561 437 -559
rect 443 -555 444 -553
rect 443 -561 444 -559
rect 450 -555 451 -553
rect 450 -561 451 -559
rect 457 -561 458 -559
rect 460 -561 461 -559
rect 464 -555 465 -553
rect 464 -561 465 -559
rect 471 -555 472 -553
rect 471 -561 472 -559
rect 478 -555 479 -553
rect 478 -561 479 -559
rect 485 -555 486 -553
rect 485 -561 486 -559
rect 492 -555 493 -553
rect 492 -561 493 -559
rect 499 -555 500 -553
rect 502 -555 503 -553
rect 506 -555 507 -553
rect 506 -561 507 -559
rect 513 -555 514 -553
rect 513 -561 514 -559
rect 520 -555 521 -553
rect 520 -561 521 -559
rect 527 -555 528 -553
rect 527 -561 528 -559
rect 534 -555 535 -553
rect 534 -561 535 -559
rect 541 -555 542 -553
rect 541 -561 542 -559
rect 548 -555 549 -553
rect 548 -561 549 -559
rect 555 -555 556 -553
rect 555 -561 556 -559
rect 562 -555 563 -553
rect 562 -561 563 -559
rect 569 -555 570 -553
rect 569 -561 570 -559
rect 576 -555 577 -553
rect 576 -561 577 -559
rect 583 -555 584 -553
rect 583 -561 584 -559
rect 590 -555 591 -553
rect 590 -561 591 -559
rect 597 -555 598 -553
rect 597 -561 598 -559
rect 604 -555 605 -553
rect 604 -561 605 -559
rect 611 -555 612 -553
rect 611 -561 612 -559
rect 618 -555 619 -553
rect 618 -561 619 -559
rect 628 -555 629 -553
rect 625 -561 626 -559
rect 632 -555 633 -553
rect 632 -561 633 -559
rect 639 -555 640 -553
rect 639 -561 640 -559
rect 646 -555 647 -553
rect 646 -561 647 -559
rect 653 -555 654 -553
rect 653 -561 654 -559
rect 656 -561 657 -559
rect 660 -555 661 -553
rect 660 -561 661 -559
rect 667 -555 668 -553
rect 667 -561 668 -559
rect 670 -561 671 -559
rect 674 -555 675 -553
rect 674 -561 675 -559
rect 681 -555 682 -553
rect 684 -561 685 -559
rect 688 -555 689 -553
rect 688 -561 689 -559
rect 2 -612 3 -610
rect 2 -618 3 -616
rect 9 -612 10 -610
rect 9 -618 10 -616
rect 19 -612 20 -610
rect 23 -612 24 -610
rect 23 -618 24 -616
rect 30 -612 31 -610
rect 30 -618 31 -616
rect 40 -612 41 -610
rect 44 -618 45 -616
rect 51 -612 52 -610
rect 51 -618 52 -616
rect 58 -612 59 -610
rect 58 -618 59 -616
rect 65 -612 66 -610
rect 65 -618 66 -616
rect 75 -618 76 -616
rect 79 -612 80 -610
rect 79 -618 80 -616
rect 86 -618 87 -616
rect 93 -612 94 -610
rect 96 -612 97 -610
rect 93 -618 94 -616
rect 100 -612 101 -610
rect 103 -612 104 -610
rect 100 -618 101 -616
rect 107 -612 108 -610
rect 107 -618 108 -616
rect 114 -612 115 -610
rect 114 -618 115 -616
rect 117 -618 118 -616
rect 121 -612 122 -610
rect 121 -618 122 -616
rect 128 -612 129 -610
rect 131 -612 132 -610
rect 128 -618 129 -616
rect 135 -612 136 -610
rect 135 -618 136 -616
rect 142 -612 143 -610
rect 142 -618 143 -616
rect 149 -612 150 -610
rect 149 -618 150 -616
rect 156 -618 157 -616
rect 159 -618 160 -616
rect 163 -612 164 -610
rect 163 -618 164 -616
rect 166 -618 167 -616
rect 170 -612 171 -610
rect 173 -618 174 -616
rect 177 -612 178 -610
rect 180 -612 181 -610
rect 177 -618 178 -616
rect 184 -612 185 -610
rect 187 -612 188 -610
rect 187 -618 188 -616
rect 191 -612 192 -610
rect 191 -618 192 -616
rect 198 -612 199 -610
rect 198 -618 199 -616
rect 205 -612 206 -610
rect 205 -618 206 -616
rect 212 -612 213 -610
rect 212 -618 213 -616
rect 219 -612 220 -610
rect 219 -618 220 -616
rect 226 -612 227 -610
rect 226 -618 227 -616
rect 233 -612 234 -610
rect 236 -612 237 -610
rect 243 -612 244 -610
rect 240 -618 241 -616
rect 243 -618 244 -616
rect 247 -612 248 -610
rect 247 -618 248 -616
rect 254 -612 255 -610
rect 254 -618 255 -616
rect 264 -612 265 -610
rect 268 -612 269 -610
rect 268 -618 269 -616
rect 275 -612 276 -610
rect 278 -618 279 -616
rect 282 -612 283 -610
rect 282 -618 283 -616
rect 289 -612 290 -610
rect 289 -618 290 -616
rect 296 -612 297 -610
rect 296 -618 297 -616
rect 303 -612 304 -610
rect 306 -612 307 -610
rect 310 -612 311 -610
rect 310 -618 311 -616
rect 317 -612 318 -610
rect 317 -618 318 -616
rect 324 -612 325 -610
rect 324 -618 325 -616
rect 331 -612 332 -610
rect 331 -618 332 -616
rect 338 -612 339 -610
rect 338 -618 339 -616
rect 345 -612 346 -610
rect 345 -618 346 -616
rect 355 -618 356 -616
rect 359 -612 360 -610
rect 359 -618 360 -616
rect 366 -612 367 -610
rect 369 -612 370 -610
rect 366 -618 367 -616
rect 369 -618 370 -616
rect 373 -612 374 -610
rect 373 -618 374 -616
rect 380 -612 381 -610
rect 383 -612 384 -610
rect 380 -618 381 -616
rect 383 -618 384 -616
rect 387 -612 388 -610
rect 387 -618 388 -616
rect 390 -618 391 -616
rect 397 -612 398 -610
rect 394 -618 395 -616
rect 401 -612 402 -610
rect 401 -618 402 -616
rect 408 -612 409 -610
rect 408 -618 409 -616
rect 415 -612 416 -610
rect 415 -618 416 -616
rect 422 -612 423 -610
rect 422 -618 423 -616
rect 429 -612 430 -610
rect 429 -618 430 -616
rect 436 -612 437 -610
rect 436 -618 437 -616
rect 443 -612 444 -610
rect 443 -618 444 -616
rect 450 -612 451 -610
rect 453 -618 454 -616
rect 457 -612 458 -610
rect 457 -618 458 -616
rect 464 -612 465 -610
rect 467 -612 468 -610
rect 464 -618 465 -616
rect 471 -612 472 -610
rect 474 -612 475 -610
rect 474 -618 475 -616
rect 478 -612 479 -610
rect 478 -618 479 -616
rect 485 -612 486 -610
rect 485 -618 486 -616
rect 492 -618 493 -616
rect 495 -618 496 -616
rect 499 -612 500 -610
rect 499 -618 500 -616
rect 506 -612 507 -610
rect 506 -618 507 -616
rect 513 -612 514 -610
rect 513 -618 514 -616
rect 520 -612 521 -610
rect 520 -618 521 -616
rect 527 -612 528 -610
rect 527 -618 528 -616
rect 534 -612 535 -610
rect 534 -618 535 -616
rect 541 -612 542 -610
rect 541 -618 542 -616
rect 548 -612 549 -610
rect 548 -618 549 -616
rect 555 -612 556 -610
rect 555 -618 556 -616
rect 562 -612 563 -610
rect 562 -618 563 -616
rect 569 -612 570 -610
rect 569 -618 570 -616
rect 576 -612 577 -610
rect 576 -618 577 -616
rect 583 -612 584 -610
rect 583 -618 584 -616
rect 590 -612 591 -610
rect 590 -618 591 -616
rect 597 -612 598 -610
rect 597 -618 598 -616
rect 604 -612 605 -610
rect 611 -612 612 -610
rect 611 -618 612 -616
rect 618 -612 619 -610
rect 618 -618 619 -616
rect 625 -612 626 -610
rect 625 -618 626 -616
rect 632 -612 633 -610
rect 632 -618 633 -616
rect 639 -612 640 -610
rect 639 -618 640 -616
rect 646 -612 647 -610
rect 646 -618 647 -616
rect 653 -612 654 -610
rect 656 -612 657 -610
rect 653 -618 654 -616
rect 660 -612 661 -610
rect 660 -618 661 -616
rect 677 -612 678 -610
rect 688 -612 689 -610
rect 2 -685 3 -683
rect 2 -691 3 -689
rect 9 -685 10 -683
rect 9 -691 10 -689
rect 16 -685 17 -683
rect 19 -691 20 -689
rect 23 -685 24 -683
rect 23 -691 24 -689
rect 30 -685 31 -683
rect 30 -691 31 -689
rect 37 -685 38 -683
rect 37 -691 38 -689
rect 44 -685 45 -683
rect 44 -691 45 -689
rect 54 -685 55 -683
rect 61 -685 62 -683
rect 65 -685 66 -683
rect 65 -691 66 -689
rect 72 -685 73 -683
rect 72 -691 73 -689
rect 79 -685 80 -683
rect 82 -691 83 -689
rect 89 -685 90 -683
rect 89 -691 90 -689
rect 93 -685 94 -683
rect 96 -685 97 -683
rect 93 -691 94 -689
rect 100 -691 101 -689
rect 103 -691 104 -689
rect 107 -685 108 -683
rect 107 -691 108 -689
rect 114 -685 115 -683
rect 114 -691 115 -689
rect 121 -685 122 -683
rect 121 -691 122 -689
rect 128 -685 129 -683
rect 128 -691 129 -689
rect 135 -685 136 -683
rect 138 -691 139 -689
rect 142 -685 143 -683
rect 145 -685 146 -683
rect 142 -691 143 -689
rect 149 -685 150 -683
rect 149 -691 150 -689
rect 156 -685 157 -683
rect 156 -691 157 -689
rect 163 -685 164 -683
rect 166 -685 167 -683
rect 166 -691 167 -689
rect 170 -685 171 -683
rect 170 -691 171 -689
rect 177 -685 178 -683
rect 177 -691 178 -689
rect 184 -685 185 -683
rect 184 -691 185 -689
rect 187 -691 188 -689
rect 191 -685 192 -683
rect 194 -685 195 -683
rect 191 -691 192 -689
rect 198 -685 199 -683
rect 198 -691 199 -689
rect 205 -685 206 -683
rect 205 -691 206 -689
rect 212 -685 213 -683
rect 212 -691 213 -689
rect 215 -691 216 -689
rect 219 -685 220 -683
rect 219 -691 220 -689
rect 229 -685 230 -683
rect 226 -691 227 -689
rect 233 -685 234 -683
rect 233 -691 234 -689
rect 236 -691 237 -689
rect 240 -685 241 -683
rect 243 -685 244 -683
rect 240 -691 241 -689
rect 243 -691 244 -689
rect 247 -685 248 -683
rect 247 -691 248 -689
rect 254 -685 255 -683
rect 254 -691 255 -689
rect 261 -685 262 -683
rect 261 -691 262 -689
rect 268 -685 269 -683
rect 268 -691 269 -689
rect 278 -685 279 -683
rect 278 -691 279 -689
rect 282 -685 283 -683
rect 285 -685 286 -683
rect 289 -685 290 -683
rect 289 -691 290 -689
rect 299 -685 300 -683
rect 296 -691 297 -689
rect 299 -691 300 -689
rect 303 -685 304 -683
rect 303 -691 304 -689
rect 310 -685 311 -683
rect 310 -691 311 -689
rect 317 -685 318 -683
rect 317 -691 318 -689
rect 324 -685 325 -683
rect 324 -691 325 -689
rect 331 -685 332 -683
rect 331 -691 332 -689
rect 338 -685 339 -683
rect 338 -691 339 -689
rect 345 -685 346 -683
rect 348 -685 349 -683
rect 345 -691 346 -689
rect 348 -691 349 -689
rect 352 -685 353 -683
rect 352 -691 353 -689
rect 359 -691 360 -689
rect 362 -691 363 -689
rect 366 -685 367 -683
rect 369 -685 370 -683
rect 366 -691 367 -689
rect 369 -691 370 -689
rect 376 -685 377 -683
rect 373 -691 374 -689
rect 376 -691 377 -689
rect 380 -685 381 -683
rect 380 -691 381 -689
rect 387 -685 388 -683
rect 387 -691 388 -689
rect 394 -685 395 -683
rect 394 -691 395 -689
rect 401 -685 402 -683
rect 401 -691 402 -689
rect 411 -685 412 -683
rect 408 -691 409 -689
rect 411 -691 412 -689
rect 415 -685 416 -683
rect 415 -691 416 -689
rect 422 -685 423 -683
rect 425 -685 426 -683
rect 422 -691 423 -689
rect 429 -685 430 -683
rect 429 -691 430 -689
rect 436 -685 437 -683
rect 436 -691 437 -689
rect 443 -685 444 -683
rect 443 -691 444 -689
rect 453 -685 454 -683
rect 450 -691 451 -689
rect 453 -691 454 -689
rect 457 -685 458 -683
rect 457 -691 458 -689
rect 460 -691 461 -689
rect 464 -685 465 -683
rect 464 -691 465 -689
rect 467 -691 468 -689
rect 471 -685 472 -683
rect 471 -691 472 -689
rect 478 -685 479 -683
rect 478 -691 479 -689
rect 485 -685 486 -683
rect 485 -691 486 -689
rect 492 -685 493 -683
rect 492 -691 493 -689
rect 499 -685 500 -683
rect 499 -691 500 -689
rect 506 -685 507 -683
rect 506 -691 507 -689
rect 513 -685 514 -683
rect 513 -691 514 -689
rect 520 -685 521 -683
rect 520 -691 521 -689
rect 527 -685 528 -683
rect 527 -691 528 -689
rect 534 -685 535 -683
rect 534 -691 535 -689
rect 541 -685 542 -683
rect 541 -691 542 -689
rect 548 -685 549 -683
rect 548 -691 549 -689
rect 555 -685 556 -683
rect 555 -691 556 -689
rect 562 -685 563 -683
rect 562 -691 563 -689
rect 569 -685 570 -683
rect 569 -691 570 -689
rect 576 -685 577 -683
rect 576 -691 577 -689
rect 583 -685 584 -683
rect 583 -691 584 -689
rect 590 -685 591 -683
rect 590 -691 591 -689
rect 597 -685 598 -683
rect 597 -691 598 -689
rect 604 -685 605 -683
rect 604 -691 605 -689
rect 611 -685 612 -683
rect 611 -691 612 -689
rect 618 -685 619 -683
rect 618 -691 619 -689
rect 625 -685 626 -683
rect 625 -691 626 -689
rect 632 -685 633 -683
rect 632 -691 633 -689
rect 639 -685 640 -683
rect 639 -691 640 -689
rect 646 -685 647 -683
rect 646 -691 647 -689
rect 653 -685 654 -683
rect 653 -691 654 -689
rect 660 -685 661 -683
rect 660 -691 661 -689
rect 667 -685 668 -683
rect 667 -691 668 -689
rect 677 -685 678 -683
rect 674 -691 675 -689
rect 681 -685 682 -683
rect 688 -685 689 -683
rect 688 -691 689 -689
rect 695 -685 696 -683
rect 695 -691 696 -689
rect 702 -685 703 -683
rect 702 -691 703 -689
rect 716 -685 717 -683
rect 719 -685 720 -683
rect 730 -685 731 -683
rect 730 -691 731 -689
rect 2 -752 3 -750
rect 2 -758 3 -756
rect 9 -752 10 -750
rect 9 -758 10 -756
rect 16 -752 17 -750
rect 16 -758 17 -756
rect 23 -752 24 -750
rect 23 -758 24 -756
rect 30 -752 31 -750
rect 30 -758 31 -756
rect 40 -752 41 -750
rect 44 -752 45 -750
rect 44 -758 45 -756
rect 51 -752 52 -750
rect 51 -758 52 -756
rect 58 -752 59 -750
rect 58 -758 59 -756
rect 65 -752 66 -750
rect 65 -758 66 -756
rect 72 -752 73 -750
rect 72 -758 73 -756
rect 79 -752 80 -750
rect 79 -758 80 -756
rect 89 -752 90 -750
rect 86 -758 87 -756
rect 89 -758 90 -756
rect 93 -752 94 -750
rect 93 -758 94 -756
rect 100 -752 101 -750
rect 100 -758 101 -756
rect 103 -758 104 -756
rect 107 -752 108 -750
rect 107 -758 108 -756
rect 114 -752 115 -750
rect 114 -758 115 -756
rect 124 -752 125 -750
rect 121 -758 122 -756
rect 124 -758 125 -756
rect 128 -752 129 -750
rect 128 -758 129 -756
rect 135 -752 136 -750
rect 135 -758 136 -756
rect 142 -752 143 -750
rect 142 -758 143 -756
rect 149 -752 150 -750
rect 149 -758 150 -756
rect 156 -752 157 -750
rect 156 -758 157 -756
rect 163 -752 164 -750
rect 163 -758 164 -756
rect 170 -752 171 -750
rect 170 -758 171 -756
rect 177 -752 178 -750
rect 177 -758 178 -756
rect 184 -752 185 -750
rect 184 -758 185 -756
rect 191 -752 192 -750
rect 191 -758 192 -756
rect 198 -752 199 -750
rect 201 -752 202 -750
rect 198 -758 199 -756
rect 205 -752 206 -750
rect 205 -758 206 -756
rect 212 -752 213 -750
rect 212 -758 213 -756
rect 219 -752 220 -750
rect 219 -758 220 -756
rect 226 -752 227 -750
rect 226 -758 227 -756
rect 229 -758 230 -756
rect 233 -758 234 -756
rect 236 -758 237 -756
rect 240 -752 241 -750
rect 240 -758 241 -756
rect 247 -752 248 -750
rect 247 -758 248 -756
rect 250 -758 251 -756
rect 254 -752 255 -750
rect 254 -758 255 -756
rect 261 -752 262 -750
rect 261 -758 262 -756
rect 268 -752 269 -750
rect 268 -758 269 -756
rect 278 -752 279 -750
rect 282 -752 283 -750
rect 292 -752 293 -750
rect 296 -752 297 -750
rect 296 -758 297 -756
rect 303 -752 304 -750
rect 303 -758 304 -756
rect 310 -752 311 -750
rect 310 -758 311 -756
rect 317 -752 318 -750
rect 317 -758 318 -756
rect 324 -752 325 -750
rect 327 -752 328 -750
rect 327 -758 328 -756
rect 331 -752 332 -750
rect 331 -758 332 -756
rect 341 -752 342 -750
rect 338 -758 339 -756
rect 341 -758 342 -756
rect 345 -752 346 -750
rect 345 -758 346 -756
rect 352 -752 353 -750
rect 352 -758 353 -756
rect 362 -752 363 -750
rect 359 -758 360 -756
rect 362 -758 363 -756
rect 366 -752 367 -750
rect 366 -758 367 -756
rect 373 -752 374 -750
rect 373 -758 374 -756
rect 380 -752 381 -750
rect 380 -758 381 -756
rect 383 -758 384 -756
rect 387 -752 388 -750
rect 387 -758 388 -756
rect 390 -758 391 -756
rect 397 -758 398 -756
rect 401 -752 402 -750
rect 401 -758 402 -756
rect 408 -752 409 -750
rect 408 -758 409 -756
rect 411 -758 412 -756
rect 415 -752 416 -750
rect 415 -758 416 -756
rect 422 -752 423 -750
rect 422 -758 423 -756
rect 429 -752 430 -750
rect 432 -752 433 -750
rect 436 -752 437 -750
rect 436 -758 437 -756
rect 443 -752 444 -750
rect 443 -758 444 -756
rect 450 -752 451 -750
rect 453 -752 454 -750
rect 450 -758 451 -756
rect 453 -758 454 -756
rect 457 -752 458 -750
rect 457 -758 458 -756
rect 464 -752 465 -750
rect 464 -758 465 -756
rect 471 -752 472 -750
rect 471 -758 472 -756
rect 478 -752 479 -750
rect 478 -758 479 -756
rect 485 -752 486 -750
rect 492 -752 493 -750
rect 492 -758 493 -756
rect 495 -758 496 -756
rect 499 -752 500 -750
rect 499 -758 500 -756
rect 506 -752 507 -750
rect 506 -758 507 -756
rect 513 -752 514 -750
rect 513 -758 514 -756
rect 520 -752 521 -750
rect 520 -758 521 -756
rect 527 -758 528 -756
rect 530 -758 531 -756
rect 534 -752 535 -750
rect 534 -758 535 -756
rect 541 -758 542 -756
rect 544 -758 545 -756
rect 548 -752 549 -750
rect 548 -758 549 -756
rect 555 -752 556 -750
rect 555 -758 556 -756
rect 562 -752 563 -750
rect 565 -752 566 -750
rect 562 -758 563 -756
rect 569 -752 570 -750
rect 569 -758 570 -756
rect 576 -752 577 -750
rect 576 -758 577 -756
rect 583 -752 584 -750
rect 583 -758 584 -756
rect 586 -758 587 -756
rect 590 -752 591 -750
rect 590 -758 591 -756
rect 597 -752 598 -750
rect 597 -758 598 -756
rect 604 -752 605 -750
rect 604 -758 605 -756
rect 611 -752 612 -750
rect 611 -758 612 -756
rect 618 -752 619 -750
rect 618 -758 619 -756
rect 625 -752 626 -750
rect 625 -758 626 -756
rect 632 -752 633 -750
rect 632 -758 633 -756
rect 639 -752 640 -750
rect 639 -758 640 -756
rect 646 -752 647 -750
rect 646 -758 647 -756
rect 653 -752 654 -750
rect 653 -758 654 -756
rect 660 -752 661 -750
rect 660 -758 661 -756
rect 667 -752 668 -750
rect 667 -758 668 -756
rect 674 -752 675 -750
rect 674 -758 675 -756
rect 681 -752 682 -750
rect 681 -758 682 -756
rect 688 -752 689 -750
rect 688 -758 689 -756
rect 695 -752 696 -750
rect 695 -758 696 -756
rect 702 -752 703 -750
rect 702 -758 703 -756
rect 712 -758 713 -756
rect 716 -752 717 -750
rect 716 -758 717 -756
rect 723 -752 724 -750
rect 723 -758 724 -756
rect 733 -752 734 -750
rect 733 -758 734 -756
rect 737 -752 738 -750
rect 737 -758 738 -756
rect 744 -752 745 -750
rect 744 -758 745 -756
rect 754 -752 755 -750
rect 754 -758 755 -756
rect 800 -752 801 -750
rect 807 -752 808 -750
rect 807 -758 808 -756
rect 2 -829 3 -827
rect 2 -835 3 -833
rect 9 -829 10 -827
rect 9 -835 10 -833
rect 16 -829 17 -827
rect 16 -835 17 -833
rect 23 -829 24 -827
rect 30 -829 31 -827
rect 37 -829 38 -827
rect 37 -835 38 -833
rect 44 -829 45 -827
rect 44 -835 45 -833
rect 54 -829 55 -827
rect 54 -835 55 -833
rect 58 -829 59 -827
rect 58 -835 59 -833
rect 65 -829 66 -827
rect 65 -835 66 -833
rect 72 -829 73 -827
rect 72 -835 73 -833
rect 79 -829 80 -827
rect 82 -829 83 -827
rect 79 -835 80 -833
rect 82 -835 83 -833
rect 86 -829 87 -827
rect 89 -829 90 -827
rect 93 -829 94 -827
rect 93 -835 94 -833
rect 100 -829 101 -827
rect 100 -835 101 -833
rect 107 -829 108 -827
rect 110 -829 111 -827
rect 114 -829 115 -827
rect 114 -835 115 -833
rect 121 -829 122 -827
rect 124 -829 125 -827
rect 121 -835 122 -833
rect 128 -829 129 -827
rect 128 -835 129 -833
rect 135 -829 136 -827
rect 138 -829 139 -827
rect 138 -835 139 -833
rect 142 -835 143 -833
rect 145 -835 146 -833
rect 149 -829 150 -827
rect 149 -835 150 -833
rect 156 -829 157 -827
rect 156 -835 157 -833
rect 163 -829 164 -827
rect 166 -835 167 -833
rect 170 -829 171 -827
rect 170 -835 171 -833
rect 177 -829 178 -827
rect 177 -835 178 -833
rect 184 -829 185 -827
rect 184 -835 185 -833
rect 191 -829 192 -827
rect 198 -829 199 -827
rect 201 -829 202 -827
rect 201 -835 202 -833
rect 205 -829 206 -827
rect 205 -835 206 -833
rect 212 -829 213 -827
rect 215 -829 216 -827
rect 212 -835 213 -833
rect 215 -835 216 -833
rect 219 -829 220 -827
rect 222 -829 223 -827
rect 219 -835 220 -833
rect 226 -829 227 -827
rect 226 -835 227 -833
rect 233 -829 234 -827
rect 233 -835 234 -833
rect 240 -829 241 -827
rect 243 -829 244 -827
rect 240 -835 241 -833
rect 247 -829 248 -827
rect 247 -835 248 -833
rect 254 -829 255 -827
rect 254 -835 255 -833
rect 264 -829 265 -827
rect 268 -829 269 -827
rect 268 -835 269 -833
rect 275 -829 276 -827
rect 275 -835 276 -833
rect 285 -829 286 -827
rect 282 -835 283 -833
rect 289 -829 290 -827
rect 292 -829 293 -827
rect 292 -835 293 -833
rect 296 -829 297 -827
rect 299 -829 300 -827
rect 296 -835 297 -833
rect 299 -835 300 -833
rect 303 -829 304 -827
rect 303 -835 304 -833
rect 310 -829 311 -827
rect 310 -835 311 -833
rect 317 -829 318 -827
rect 317 -835 318 -833
rect 324 -829 325 -827
rect 324 -835 325 -833
rect 331 -829 332 -827
rect 334 -829 335 -827
rect 331 -835 332 -833
rect 334 -835 335 -833
rect 338 -829 339 -827
rect 338 -835 339 -833
rect 345 -829 346 -827
rect 345 -835 346 -833
rect 352 -829 353 -827
rect 352 -835 353 -833
rect 359 -829 360 -827
rect 359 -835 360 -833
rect 366 -829 367 -827
rect 366 -835 367 -833
rect 373 -829 374 -827
rect 373 -835 374 -833
rect 380 -829 381 -827
rect 383 -829 384 -827
rect 380 -835 381 -833
rect 387 -829 388 -827
rect 390 -829 391 -827
rect 390 -835 391 -833
rect 394 -829 395 -827
rect 394 -835 395 -833
rect 404 -829 405 -827
rect 401 -835 402 -833
rect 404 -835 405 -833
rect 408 -829 409 -827
rect 408 -835 409 -833
rect 418 -829 419 -827
rect 418 -835 419 -833
rect 422 -829 423 -827
rect 422 -835 423 -833
rect 429 -829 430 -827
rect 429 -835 430 -833
rect 436 -829 437 -827
rect 439 -829 440 -827
rect 436 -835 437 -833
rect 439 -835 440 -833
rect 443 -829 444 -827
rect 443 -835 444 -833
rect 450 -829 451 -827
rect 450 -835 451 -833
rect 457 -829 458 -827
rect 460 -829 461 -827
rect 460 -835 461 -833
rect 464 -829 465 -827
rect 464 -835 465 -833
rect 471 -829 472 -827
rect 471 -835 472 -833
rect 478 -829 479 -827
rect 478 -835 479 -833
rect 488 -829 489 -827
rect 485 -835 486 -833
rect 488 -835 489 -833
rect 495 -829 496 -827
rect 495 -835 496 -833
rect 499 -829 500 -827
rect 499 -835 500 -833
rect 506 -829 507 -827
rect 506 -835 507 -833
rect 513 -829 514 -827
rect 513 -835 514 -833
rect 520 -829 521 -827
rect 523 -829 524 -827
rect 523 -835 524 -833
rect 527 -835 528 -833
rect 530 -835 531 -833
rect 534 -829 535 -827
rect 534 -835 535 -833
rect 541 -829 542 -827
rect 541 -835 542 -833
rect 548 -829 549 -827
rect 548 -835 549 -833
rect 555 -829 556 -827
rect 555 -835 556 -833
rect 562 -829 563 -827
rect 562 -835 563 -833
rect 569 -829 570 -827
rect 569 -835 570 -833
rect 576 -829 577 -827
rect 576 -835 577 -833
rect 583 -829 584 -827
rect 583 -835 584 -833
rect 590 -829 591 -827
rect 590 -835 591 -833
rect 597 -829 598 -827
rect 597 -835 598 -833
rect 604 -829 605 -827
rect 604 -835 605 -833
rect 611 -829 612 -827
rect 611 -835 612 -833
rect 618 -829 619 -827
rect 618 -835 619 -833
rect 625 -829 626 -827
rect 625 -835 626 -833
rect 632 -829 633 -827
rect 632 -835 633 -833
rect 639 -829 640 -827
rect 639 -835 640 -833
rect 646 -829 647 -827
rect 646 -835 647 -833
rect 653 -829 654 -827
rect 653 -835 654 -833
rect 660 -829 661 -827
rect 660 -835 661 -833
rect 667 -829 668 -827
rect 667 -835 668 -833
rect 674 -829 675 -827
rect 674 -835 675 -833
rect 681 -829 682 -827
rect 681 -835 682 -833
rect 688 -829 689 -827
rect 688 -835 689 -833
rect 695 -829 696 -827
rect 695 -835 696 -833
rect 702 -829 703 -827
rect 702 -835 703 -833
rect 709 -829 710 -827
rect 709 -835 710 -833
rect 716 -829 717 -827
rect 716 -835 717 -833
rect 723 -829 724 -827
rect 723 -835 724 -833
rect 730 -829 731 -827
rect 730 -835 731 -833
rect 737 -829 738 -827
rect 737 -835 738 -833
rect 744 -829 745 -827
rect 744 -835 745 -833
rect 751 -829 752 -827
rect 751 -835 752 -833
rect 758 -829 759 -827
rect 758 -835 759 -833
rect 765 -829 766 -827
rect 765 -835 766 -833
rect 772 -829 773 -827
rect 772 -835 773 -833
rect 779 -829 780 -827
rect 779 -835 780 -833
rect 786 -829 787 -827
rect 786 -835 787 -833
rect 793 -829 794 -827
rect 793 -835 794 -833
rect 803 -829 804 -827
rect 803 -835 804 -833
rect 807 -829 808 -827
rect 807 -835 808 -833
rect 9 -916 10 -914
rect 9 -922 10 -920
rect 16 -916 17 -914
rect 16 -922 17 -920
rect 23 -916 24 -914
rect 23 -922 24 -920
rect 30 -916 31 -914
rect 30 -922 31 -920
rect 37 -916 38 -914
rect 37 -922 38 -920
rect 44 -916 45 -914
rect 44 -922 45 -920
rect 51 -916 52 -914
rect 51 -922 52 -920
rect 58 -916 59 -914
rect 58 -922 59 -920
rect 65 -916 66 -914
rect 72 -916 73 -914
rect 79 -916 80 -914
rect 79 -922 80 -920
rect 86 -916 87 -914
rect 86 -922 87 -920
rect 89 -922 90 -920
rect 93 -916 94 -914
rect 93 -922 94 -920
rect 100 -916 101 -914
rect 100 -922 101 -920
rect 107 -916 108 -914
rect 107 -922 108 -920
rect 114 -916 115 -914
rect 114 -922 115 -920
rect 121 -916 122 -914
rect 121 -922 122 -920
rect 128 -916 129 -914
rect 135 -916 136 -914
rect 135 -922 136 -920
rect 142 -916 143 -914
rect 142 -922 143 -920
rect 149 -916 150 -914
rect 152 -916 153 -914
rect 149 -922 150 -920
rect 152 -922 153 -920
rect 156 -916 157 -914
rect 159 -916 160 -914
rect 163 -916 164 -914
rect 163 -922 164 -920
rect 170 -916 171 -914
rect 173 -916 174 -914
rect 177 -916 178 -914
rect 180 -916 181 -914
rect 180 -922 181 -920
rect 184 -916 185 -914
rect 184 -922 185 -920
rect 191 -916 192 -914
rect 191 -922 192 -920
rect 201 -916 202 -914
rect 198 -922 199 -920
rect 201 -922 202 -920
rect 205 -916 206 -914
rect 205 -922 206 -920
rect 212 -916 213 -914
rect 212 -922 213 -920
rect 219 -916 220 -914
rect 219 -922 220 -920
rect 222 -922 223 -920
rect 226 -916 227 -914
rect 229 -916 230 -914
rect 226 -922 227 -920
rect 229 -922 230 -920
rect 233 -916 234 -914
rect 236 -916 237 -914
rect 233 -922 234 -920
rect 236 -922 237 -920
rect 240 -916 241 -914
rect 243 -916 244 -914
rect 243 -922 244 -920
rect 247 -916 248 -914
rect 247 -922 248 -920
rect 254 -916 255 -914
rect 254 -922 255 -920
rect 261 -916 262 -914
rect 261 -922 262 -920
rect 268 -916 269 -914
rect 268 -922 269 -920
rect 275 -916 276 -914
rect 278 -916 279 -914
rect 275 -922 276 -920
rect 278 -922 279 -920
rect 282 -916 283 -914
rect 285 -922 286 -920
rect 289 -916 290 -914
rect 289 -922 290 -920
rect 296 -916 297 -914
rect 296 -922 297 -920
rect 303 -916 304 -914
rect 303 -922 304 -920
rect 310 -916 311 -914
rect 310 -922 311 -920
rect 317 -916 318 -914
rect 317 -922 318 -920
rect 324 -916 325 -914
rect 324 -922 325 -920
rect 331 -916 332 -914
rect 331 -922 332 -920
rect 338 -916 339 -914
rect 338 -922 339 -920
rect 348 -916 349 -914
rect 345 -922 346 -920
rect 348 -922 349 -920
rect 352 -916 353 -914
rect 352 -922 353 -920
rect 359 -916 360 -914
rect 359 -922 360 -920
rect 366 -916 367 -914
rect 366 -922 367 -920
rect 373 -916 374 -914
rect 373 -922 374 -920
rect 383 -916 384 -914
rect 380 -922 381 -920
rect 387 -916 388 -914
rect 387 -922 388 -920
rect 394 -916 395 -914
rect 397 -916 398 -914
rect 394 -922 395 -920
rect 397 -922 398 -920
rect 401 -916 402 -914
rect 401 -922 402 -920
rect 408 -916 409 -914
rect 411 -916 412 -914
rect 408 -922 409 -920
rect 411 -922 412 -920
rect 415 -916 416 -914
rect 415 -922 416 -920
rect 418 -922 419 -920
rect 422 -916 423 -914
rect 422 -922 423 -920
rect 429 -916 430 -914
rect 429 -922 430 -920
rect 436 -916 437 -914
rect 436 -922 437 -920
rect 443 -916 444 -914
rect 443 -922 444 -920
rect 450 -916 451 -914
rect 450 -922 451 -920
rect 457 -916 458 -914
rect 460 -916 461 -914
rect 457 -922 458 -920
rect 460 -922 461 -920
rect 464 -916 465 -914
rect 467 -916 468 -914
rect 467 -922 468 -920
rect 471 -916 472 -914
rect 471 -922 472 -920
rect 478 -916 479 -914
rect 478 -922 479 -920
rect 488 -916 489 -914
rect 488 -922 489 -920
rect 492 -916 493 -914
rect 492 -922 493 -920
rect 499 -916 500 -914
rect 499 -922 500 -920
rect 502 -922 503 -920
rect 506 -916 507 -914
rect 506 -922 507 -920
rect 513 -916 514 -914
rect 513 -922 514 -920
rect 520 -916 521 -914
rect 520 -922 521 -920
rect 527 -916 528 -914
rect 527 -922 528 -920
rect 534 -916 535 -914
rect 534 -922 535 -920
rect 541 -916 542 -914
rect 541 -922 542 -920
rect 548 -916 549 -914
rect 548 -922 549 -920
rect 555 -916 556 -914
rect 555 -922 556 -920
rect 562 -916 563 -914
rect 562 -922 563 -920
rect 569 -916 570 -914
rect 569 -922 570 -920
rect 576 -922 577 -920
rect 579 -922 580 -920
rect 583 -916 584 -914
rect 583 -922 584 -920
rect 590 -916 591 -914
rect 590 -922 591 -920
rect 597 -916 598 -914
rect 597 -922 598 -920
rect 604 -916 605 -914
rect 604 -922 605 -920
rect 611 -916 612 -914
rect 611 -922 612 -920
rect 618 -916 619 -914
rect 618 -922 619 -920
rect 625 -916 626 -914
rect 625 -922 626 -920
rect 632 -916 633 -914
rect 632 -922 633 -920
rect 639 -916 640 -914
rect 639 -922 640 -920
rect 646 -916 647 -914
rect 646 -922 647 -920
rect 653 -916 654 -914
rect 653 -922 654 -920
rect 660 -916 661 -914
rect 660 -922 661 -920
rect 667 -916 668 -914
rect 667 -922 668 -920
rect 674 -916 675 -914
rect 674 -922 675 -920
rect 681 -916 682 -914
rect 681 -922 682 -920
rect 688 -916 689 -914
rect 688 -922 689 -920
rect 695 -916 696 -914
rect 695 -922 696 -920
rect 702 -916 703 -914
rect 702 -922 703 -920
rect 709 -916 710 -914
rect 709 -922 710 -920
rect 716 -916 717 -914
rect 716 -922 717 -920
rect 723 -916 724 -914
rect 723 -922 724 -920
rect 730 -916 731 -914
rect 730 -922 731 -920
rect 737 -916 738 -914
rect 737 -922 738 -920
rect 744 -916 745 -914
rect 744 -922 745 -920
rect 751 -916 752 -914
rect 751 -922 752 -920
rect 758 -916 759 -914
rect 758 -922 759 -920
rect 765 -916 766 -914
rect 765 -922 766 -920
rect 772 -916 773 -914
rect 775 -916 776 -914
rect 772 -922 773 -920
rect 775 -922 776 -920
rect 782 -916 783 -914
rect 779 -922 780 -920
rect 786 -916 787 -914
rect 786 -922 787 -920
rect 796 -916 797 -914
rect 9 -993 10 -991
rect 9 -999 10 -997
rect 16 -993 17 -991
rect 16 -999 17 -997
rect 23 -993 24 -991
rect 23 -999 24 -997
rect 30 -993 31 -991
rect 30 -999 31 -997
rect 37 -993 38 -991
rect 37 -999 38 -997
rect 44 -993 45 -991
rect 44 -999 45 -997
rect 51 -993 52 -991
rect 51 -999 52 -997
rect 58 -993 59 -991
rect 58 -999 59 -997
rect 65 -993 66 -991
rect 65 -999 66 -997
rect 75 -993 76 -991
rect 72 -999 73 -997
rect 79 -993 80 -991
rect 82 -993 83 -991
rect 79 -999 80 -997
rect 86 -993 87 -991
rect 86 -999 87 -997
rect 96 -993 97 -991
rect 96 -999 97 -997
rect 100 -993 101 -991
rect 103 -993 104 -991
rect 107 -993 108 -991
rect 107 -999 108 -997
rect 114 -993 115 -991
rect 117 -993 118 -991
rect 114 -999 115 -997
rect 117 -999 118 -997
rect 121 -993 122 -991
rect 121 -999 122 -997
rect 128 -993 129 -991
rect 128 -999 129 -997
rect 135 -993 136 -991
rect 135 -999 136 -997
rect 142 -993 143 -991
rect 142 -999 143 -997
rect 149 -993 150 -991
rect 149 -999 150 -997
rect 159 -993 160 -991
rect 156 -999 157 -997
rect 159 -999 160 -997
rect 163 -993 164 -991
rect 163 -999 164 -997
rect 170 -993 171 -991
rect 170 -999 171 -997
rect 177 -993 178 -991
rect 177 -999 178 -997
rect 184 -993 185 -991
rect 184 -999 185 -997
rect 191 -993 192 -991
rect 191 -999 192 -997
rect 198 -993 199 -991
rect 198 -999 199 -997
rect 205 -993 206 -991
rect 205 -999 206 -997
rect 212 -993 213 -991
rect 212 -999 213 -997
rect 219 -993 220 -991
rect 219 -999 220 -997
rect 222 -999 223 -997
rect 226 -993 227 -991
rect 226 -999 227 -997
rect 233 -993 234 -991
rect 236 -993 237 -991
rect 233 -999 234 -997
rect 240 -993 241 -991
rect 243 -993 244 -991
rect 240 -999 241 -997
rect 243 -999 244 -997
rect 247 -993 248 -991
rect 247 -999 248 -997
rect 254 -993 255 -991
rect 257 -993 258 -991
rect 254 -999 255 -997
rect 261 -993 262 -991
rect 261 -999 262 -997
rect 268 -993 269 -991
rect 268 -999 269 -997
rect 275 -993 276 -991
rect 275 -999 276 -997
rect 285 -993 286 -991
rect 282 -999 283 -997
rect 289 -993 290 -991
rect 289 -999 290 -997
rect 296 -993 297 -991
rect 296 -999 297 -997
rect 303 -993 304 -991
rect 303 -999 304 -997
rect 310 -993 311 -991
rect 313 -993 314 -991
rect 310 -999 311 -997
rect 313 -999 314 -997
rect 317 -993 318 -991
rect 317 -999 318 -997
rect 324 -993 325 -991
rect 324 -999 325 -997
rect 331 -993 332 -991
rect 331 -999 332 -997
rect 338 -993 339 -991
rect 338 -999 339 -997
rect 348 -993 349 -991
rect 345 -999 346 -997
rect 348 -999 349 -997
rect 352 -999 353 -997
rect 355 -999 356 -997
rect 362 -993 363 -991
rect 362 -999 363 -997
rect 369 -999 370 -997
rect 376 -993 377 -991
rect 373 -999 374 -997
rect 376 -999 377 -997
rect 380 -993 381 -991
rect 380 -999 381 -997
rect 390 -993 391 -991
rect 397 -993 398 -991
rect 397 -999 398 -997
rect 401 -993 402 -991
rect 401 -999 402 -997
rect 408 -993 409 -991
rect 408 -999 409 -997
rect 418 -993 419 -991
rect 415 -999 416 -997
rect 425 -993 426 -991
rect 425 -999 426 -997
rect 429 -993 430 -991
rect 432 -993 433 -991
rect 432 -999 433 -997
rect 436 -993 437 -991
rect 436 -999 437 -997
rect 443 -993 444 -991
rect 446 -993 447 -991
rect 443 -999 444 -997
rect 446 -999 447 -997
rect 450 -993 451 -991
rect 453 -999 454 -997
rect 457 -993 458 -991
rect 457 -999 458 -997
rect 464 -993 465 -991
rect 467 -999 468 -997
rect 471 -993 472 -991
rect 474 -993 475 -991
rect 471 -999 472 -997
rect 478 -993 479 -991
rect 478 -999 479 -997
rect 485 -993 486 -991
rect 485 -999 486 -997
rect 492 -993 493 -991
rect 492 -999 493 -997
rect 499 -993 500 -991
rect 499 -999 500 -997
rect 506 -993 507 -991
rect 506 -999 507 -997
rect 513 -993 514 -991
rect 513 -999 514 -997
rect 520 -993 521 -991
rect 520 -999 521 -997
rect 527 -993 528 -991
rect 527 -999 528 -997
rect 534 -993 535 -991
rect 534 -999 535 -997
rect 541 -993 542 -991
rect 541 -999 542 -997
rect 548 -993 549 -991
rect 548 -999 549 -997
rect 555 -993 556 -991
rect 555 -999 556 -997
rect 562 -993 563 -991
rect 562 -999 563 -997
rect 569 -993 570 -991
rect 569 -999 570 -997
rect 576 -993 577 -991
rect 576 -999 577 -997
rect 583 -993 584 -991
rect 583 -999 584 -997
rect 590 -993 591 -991
rect 590 -999 591 -997
rect 597 -993 598 -991
rect 597 -999 598 -997
rect 604 -993 605 -991
rect 604 -999 605 -997
rect 611 -993 612 -991
rect 611 -999 612 -997
rect 618 -993 619 -991
rect 618 -999 619 -997
rect 625 -993 626 -991
rect 625 -999 626 -997
rect 632 -993 633 -991
rect 632 -999 633 -997
rect 639 -993 640 -991
rect 639 -999 640 -997
rect 646 -993 647 -991
rect 646 -999 647 -997
rect 653 -993 654 -991
rect 653 -999 654 -997
rect 660 -993 661 -991
rect 660 -999 661 -997
rect 667 -993 668 -991
rect 667 -999 668 -997
rect 674 -993 675 -991
rect 674 -999 675 -997
rect 681 -993 682 -991
rect 681 -999 682 -997
rect 688 -993 689 -991
rect 688 -999 689 -997
rect 695 -993 696 -991
rect 695 -999 696 -997
rect 702 -993 703 -991
rect 702 -999 703 -997
rect 709 -993 710 -991
rect 709 -999 710 -997
rect 716 -993 717 -991
rect 716 -999 717 -997
rect 723 -993 724 -991
rect 723 -999 724 -997
rect 730 -993 731 -991
rect 730 -999 731 -997
rect 737 -993 738 -991
rect 740 -993 741 -991
rect 737 -999 738 -997
rect 740 -999 741 -997
rect 744 -999 745 -997
rect 754 -993 755 -991
rect 754 -999 755 -997
rect 758 -993 759 -991
rect 758 -999 759 -997
rect 23 -1068 24 -1066
rect 23 -1074 24 -1072
rect 33 -1068 34 -1066
rect 37 -1068 38 -1066
rect 37 -1074 38 -1072
rect 44 -1068 45 -1066
rect 44 -1074 45 -1072
rect 51 -1068 52 -1066
rect 51 -1074 52 -1072
rect 61 -1068 62 -1066
rect 65 -1068 66 -1066
rect 65 -1074 66 -1072
rect 75 -1068 76 -1066
rect 79 -1068 80 -1066
rect 79 -1074 80 -1072
rect 86 -1068 87 -1066
rect 93 -1068 94 -1066
rect 93 -1074 94 -1072
rect 103 -1068 104 -1066
rect 107 -1068 108 -1066
rect 114 -1068 115 -1066
rect 114 -1074 115 -1072
rect 121 -1068 122 -1066
rect 121 -1074 122 -1072
rect 128 -1068 129 -1066
rect 128 -1074 129 -1072
rect 135 -1068 136 -1066
rect 135 -1074 136 -1072
rect 142 -1068 143 -1066
rect 142 -1074 143 -1072
rect 149 -1068 150 -1066
rect 152 -1068 153 -1066
rect 149 -1074 150 -1072
rect 156 -1068 157 -1066
rect 156 -1074 157 -1072
rect 163 -1068 164 -1066
rect 166 -1068 167 -1066
rect 166 -1074 167 -1072
rect 170 -1068 171 -1066
rect 170 -1074 171 -1072
rect 177 -1068 178 -1066
rect 180 -1068 181 -1066
rect 177 -1074 178 -1072
rect 184 -1068 185 -1066
rect 184 -1074 185 -1072
rect 191 -1068 192 -1066
rect 194 -1068 195 -1066
rect 194 -1074 195 -1072
rect 198 -1074 199 -1072
rect 201 -1074 202 -1072
rect 205 -1068 206 -1066
rect 205 -1074 206 -1072
rect 212 -1068 213 -1066
rect 212 -1074 213 -1072
rect 219 -1068 220 -1066
rect 219 -1074 220 -1072
rect 226 -1068 227 -1066
rect 226 -1074 227 -1072
rect 233 -1068 234 -1066
rect 233 -1074 234 -1072
rect 243 -1068 244 -1066
rect 243 -1074 244 -1072
rect 250 -1068 251 -1066
rect 254 -1068 255 -1066
rect 254 -1074 255 -1072
rect 261 -1068 262 -1066
rect 261 -1074 262 -1072
rect 268 -1068 269 -1066
rect 268 -1074 269 -1072
rect 278 -1068 279 -1066
rect 278 -1074 279 -1072
rect 282 -1068 283 -1066
rect 282 -1074 283 -1072
rect 289 -1068 290 -1066
rect 289 -1074 290 -1072
rect 296 -1068 297 -1066
rect 296 -1074 297 -1072
rect 303 -1068 304 -1066
rect 303 -1074 304 -1072
rect 310 -1068 311 -1066
rect 313 -1068 314 -1066
rect 310 -1074 311 -1072
rect 317 -1068 318 -1066
rect 317 -1074 318 -1072
rect 324 -1068 325 -1066
rect 324 -1074 325 -1072
rect 334 -1068 335 -1066
rect 331 -1074 332 -1072
rect 334 -1074 335 -1072
rect 338 -1068 339 -1066
rect 338 -1074 339 -1072
rect 345 -1068 346 -1066
rect 345 -1074 346 -1072
rect 352 -1068 353 -1066
rect 352 -1074 353 -1072
rect 359 -1068 360 -1066
rect 359 -1074 360 -1072
rect 366 -1068 367 -1066
rect 366 -1074 367 -1072
rect 373 -1068 374 -1066
rect 373 -1074 374 -1072
rect 380 -1068 381 -1066
rect 380 -1074 381 -1072
rect 387 -1068 388 -1066
rect 387 -1074 388 -1072
rect 394 -1068 395 -1066
rect 394 -1074 395 -1072
rect 401 -1068 402 -1066
rect 404 -1068 405 -1066
rect 401 -1074 402 -1072
rect 408 -1068 409 -1066
rect 411 -1068 412 -1066
rect 411 -1074 412 -1072
rect 418 -1068 419 -1066
rect 415 -1074 416 -1072
rect 418 -1074 419 -1072
rect 425 -1068 426 -1066
rect 422 -1074 423 -1072
rect 425 -1074 426 -1072
rect 429 -1068 430 -1066
rect 429 -1074 430 -1072
rect 439 -1068 440 -1066
rect 439 -1074 440 -1072
rect 443 -1068 444 -1066
rect 443 -1074 444 -1072
rect 450 -1068 451 -1066
rect 450 -1074 451 -1072
rect 453 -1074 454 -1072
rect 457 -1068 458 -1066
rect 457 -1074 458 -1072
rect 464 -1068 465 -1066
rect 464 -1074 465 -1072
rect 474 -1074 475 -1072
rect 478 -1068 479 -1066
rect 478 -1074 479 -1072
rect 481 -1074 482 -1072
rect 485 -1068 486 -1066
rect 485 -1074 486 -1072
rect 492 -1068 493 -1066
rect 495 -1068 496 -1066
rect 492 -1074 493 -1072
rect 495 -1074 496 -1072
rect 499 -1068 500 -1066
rect 499 -1074 500 -1072
rect 506 -1074 507 -1072
rect 513 -1068 514 -1066
rect 513 -1074 514 -1072
rect 520 -1068 521 -1066
rect 523 -1074 524 -1072
rect 527 -1068 528 -1066
rect 527 -1074 528 -1072
rect 534 -1074 535 -1072
rect 537 -1074 538 -1072
rect 541 -1068 542 -1066
rect 541 -1074 542 -1072
rect 548 -1068 549 -1066
rect 548 -1074 549 -1072
rect 555 -1068 556 -1066
rect 555 -1074 556 -1072
rect 562 -1074 563 -1072
rect 565 -1074 566 -1072
rect 569 -1068 570 -1066
rect 569 -1074 570 -1072
rect 576 -1068 577 -1066
rect 576 -1074 577 -1072
rect 583 -1068 584 -1066
rect 583 -1074 584 -1072
rect 590 -1068 591 -1066
rect 590 -1074 591 -1072
rect 597 -1068 598 -1066
rect 597 -1074 598 -1072
rect 604 -1068 605 -1066
rect 604 -1074 605 -1072
rect 611 -1068 612 -1066
rect 611 -1074 612 -1072
rect 618 -1068 619 -1066
rect 618 -1074 619 -1072
rect 625 -1068 626 -1066
rect 625 -1074 626 -1072
rect 632 -1068 633 -1066
rect 632 -1074 633 -1072
rect 639 -1068 640 -1066
rect 639 -1074 640 -1072
rect 646 -1068 647 -1066
rect 646 -1074 647 -1072
rect 653 -1068 654 -1066
rect 653 -1074 654 -1072
rect 660 -1068 661 -1066
rect 660 -1074 661 -1072
rect 667 -1068 668 -1066
rect 667 -1074 668 -1072
rect 674 -1068 675 -1066
rect 674 -1074 675 -1072
rect 681 -1068 682 -1066
rect 681 -1074 682 -1072
rect 688 -1068 689 -1066
rect 691 -1068 692 -1066
rect 691 -1074 692 -1072
rect 695 -1068 696 -1066
rect 695 -1074 696 -1072
rect 702 -1068 703 -1066
rect 702 -1074 703 -1072
rect 709 -1068 710 -1066
rect 709 -1074 710 -1072
rect 716 -1068 717 -1066
rect 719 -1068 720 -1066
rect 716 -1074 717 -1072
rect 723 -1068 724 -1066
rect 723 -1074 724 -1072
rect 730 -1068 731 -1066
rect 730 -1074 731 -1072
rect 737 -1068 738 -1066
rect 737 -1074 738 -1072
rect 9 -1129 10 -1127
rect 9 -1135 10 -1133
rect 16 -1129 17 -1127
rect 16 -1135 17 -1133
rect 23 -1129 24 -1127
rect 23 -1135 24 -1133
rect 30 -1129 31 -1127
rect 37 -1129 38 -1127
rect 37 -1135 38 -1133
rect 44 -1135 45 -1133
rect 47 -1135 48 -1133
rect 51 -1129 52 -1127
rect 51 -1135 52 -1133
rect 58 -1129 59 -1127
rect 58 -1135 59 -1133
rect 65 -1129 66 -1127
rect 68 -1129 69 -1127
rect 72 -1129 73 -1127
rect 72 -1135 73 -1133
rect 82 -1129 83 -1127
rect 82 -1135 83 -1133
rect 86 -1129 87 -1127
rect 86 -1135 87 -1133
rect 93 -1129 94 -1127
rect 93 -1135 94 -1133
rect 100 -1129 101 -1127
rect 100 -1135 101 -1133
rect 107 -1129 108 -1127
rect 107 -1135 108 -1133
rect 114 -1129 115 -1127
rect 114 -1135 115 -1133
rect 124 -1129 125 -1127
rect 121 -1135 122 -1133
rect 128 -1129 129 -1127
rect 128 -1135 129 -1133
rect 135 -1129 136 -1127
rect 135 -1135 136 -1133
rect 142 -1129 143 -1127
rect 145 -1129 146 -1127
rect 142 -1135 143 -1133
rect 145 -1135 146 -1133
rect 149 -1129 150 -1127
rect 149 -1135 150 -1133
rect 159 -1129 160 -1127
rect 156 -1135 157 -1133
rect 163 -1135 164 -1133
rect 166 -1135 167 -1133
rect 170 -1135 171 -1133
rect 173 -1135 174 -1133
rect 177 -1129 178 -1127
rect 180 -1129 181 -1127
rect 180 -1135 181 -1133
rect 184 -1129 185 -1127
rect 187 -1129 188 -1127
rect 184 -1135 185 -1133
rect 191 -1135 192 -1133
rect 194 -1135 195 -1133
rect 198 -1129 199 -1127
rect 198 -1135 199 -1133
rect 205 -1129 206 -1127
rect 205 -1135 206 -1133
rect 215 -1129 216 -1127
rect 215 -1135 216 -1133
rect 219 -1129 220 -1127
rect 219 -1135 220 -1133
rect 226 -1129 227 -1127
rect 226 -1135 227 -1133
rect 233 -1129 234 -1127
rect 233 -1135 234 -1133
rect 240 -1129 241 -1127
rect 247 -1129 248 -1127
rect 247 -1135 248 -1133
rect 250 -1135 251 -1133
rect 254 -1129 255 -1127
rect 254 -1135 255 -1133
rect 261 -1129 262 -1127
rect 261 -1135 262 -1133
rect 268 -1129 269 -1127
rect 268 -1135 269 -1133
rect 275 -1129 276 -1127
rect 278 -1129 279 -1127
rect 275 -1135 276 -1133
rect 278 -1135 279 -1133
rect 282 -1129 283 -1127
rect 282 -1135 283 -1133
rect 289 -1129 290 -1127
rect 289 -1135 290 -1133
rect 296 -1129 297 -1127
rect 296 -1135 297 -1133
rect 303 -1129 304 -1127
rect 303 -1135 304 -1133
rect 310 -1129 311 -1127
rect 313 -1129 314 -1127
rect 310 -1135 311 -1133
rect 317 -1129 318 -1127
rect 317 -1135 318 -1133
rect 324 -1129 325 -1127
rect 324 -1135 325 -1133
rect 331 -1135 332 -1133
rect 334 -1135 335 -1133
rect 338 -1129 339 -1127
rect 338 -1135 339 -1133
rect 348 -1129 349 -1127
rect 345 -1135 346 -1133
rect 348 -1135 349 -1133
rect 352 -1129 353 -1127
rect 352 -1135 353 -1133
rect 362 -1129 363 -1127
rect 362 -1135 363 -1133
rect 366 -1135 367 -1133
rect 369 -1135 370 -1133
rect 376 -1129 377 -1127
rect 373 -1135 374 -1133
rect 380 -1129 381 -1127
rect 383 -1129 384 -1127
rect 387 -1129 388 -1127
rect 387 -1135 388 -1133
rect 390 -1135 391 -1133
rect 397 -1129 398 -1127
rect 394 -1135 395 -1133
rect 397 -1135 398 -1133
rect 401 -1129 402 -1127
rect 401 -1135 402 -1133
rect 408 -1129 409 -1127
rect 408 -1135 409 -1133
rect 415 -1129 416 -1127
rect 415 -1135 416 -1133
rect 422 -1129 423 -1127
rect 425 -1129 426 -1127
rect 422 -1135 423 -1133
rect 429 -1129 430 -1127
rect 429 -1135 430 -1133
rect 432 -1135 433 -1133
rect 436 -1129 437 -1127
rect 436 -1135 437 -1133
rect 443 -1129 444 -1127
rect 443 -1135 444 -1133
rect 450 -1129 451 -1127
rect 450 -1135 451 -1133
rect 457 -1129 458 -1127
rect 457 -1135 458 -1133
rect 464 -1129 465 -1127
rect 464 -1135 465 -1133
rect 471 -1129 472 -1127
rect 471 -1135 472 -1133
rect 478 -1129 479 -1127
rect 478 -1135 479 -1133
rect 485 -1129 486 -1127
rect 485 -1135 486 -1133
rect 492 -1129 493 -1127
rect 492 -1135 493 -1133
rect 499 -1129 500 -1127
rect 499 -1135 500 -1133
rect 506 -1129 507 -1127
rect 506 -1135 507 -1133
rect 513 -1129 514 -1127
rect 513 -1135 514 -1133
rect 523 -1129 524 -1127
rect 523 -1135 524 -1133
rect 527 -1129 528 -1127
rect 527 -1135 528 -1133
rect 534 -1129 535 -1127
rect 534 -1135 535 -1133
rect 541 -1129 542 -1127
rect 541 -1135 542 -1133
rect 548 -1129 549 -1127
rect 548 -1135 549 -1133
rect 555 -1129 556 -1127
rect 555 -1135 556 -1133
rect 562 -1129 563 -1127
rect 562 -1135 563 -1133
rect 569 -1129 570 -1127
rect 569 -1135 570 -1133
rect 576 -1129 577 -1127
rect 576 -1135 577 -1133
rect 583 -1129 584 -1127
rect 583 -1135 584 -1133
rect 590 -1129 591 -1127
rect 590 -1135 591 -1133
rect 597 -1129 598 -1127
rect 597 -1135 598 -1133
rect 604 -1129 605 -1127
rect 604 -1135 605 -1133
rect 611 -1129 612 -1127
rect 611 -1135 612 -1133
rect 618 -1129 619 -1127
rect 618 -1135 619 -1133
rect 625 -1129 626 -1127
rect 625 -1135 626 -1133
rect 632 -1129 633 -1127
rect 632 -1135 633 -1133
rect 639 -1129 640 -1127
rect 639 -1135 640 -1133
rect 646 -1129 647 -1127
rect 646 -1135 647 -1133
rect 653 -1129 654 -1127
rect 653 -1135 654 -1133
rect 660 -1129 661 -1127
rect 660 -1135 661 -1133
rect 667 -1129 668 -1127
rect 667 -1135 668 -1133
rect 674 -1129 675 -1127
rect 677 -1129 678 -1127
rect 674 -1135 675 -1133
rect 677 -1135 678 -1133
rect 681 -1129 682 -1127
rect 684 -1129 685 -1127
rect 688 -1129 689 -1127
rect 688 -1135 689 -1133
rect 695 -1129 696 -1127
rect 695 -1135 696 -1133
rect 702 -1129 703 -1127
rect 702 -1135 703 -1133
rect 709 -1129 710 -1127
rect 709 -1135 710 -1133
rect 2 -1186 3 -1184
rect 2 -1192 3 -1190
rect 9 -1186 10 -1184
rect 9 -1192 10 -1190
rect 19 -1186 20 -1184
rect 23 -1192 24 -1190
rect 30 -1186 31 -1184
rect 30 -1192 31 -1190
rect 37 -1186 38 -1184
rect 37 -1192 38 -1190
rect 44 -1186 45 -1184
rect 44 -1192 45 -1190
rect 51 -1186 52 -1184
rect 51 -1192 52 -1190
rect 58 -1186 59 -1184
rect 58 -1192 59 -1190
rect 65 -1186 66 -1184
rect 75 -1186 76 -1184
rect 72 -1192 73 -1190
rect 75 -1192 76 -1190
rect 79 -1186 80 -1184
rect 79 -1192 80 -1190
rect 86 -1186 87 -1184
rect 89 -1192 90 -1190
rect 93 -1186 94 -1184
rect 93 -1192 94 -1190
rect 100 -1192 101 -1190
rect 107 -1186 108 -1184
rect 110 -1186 111 -1184
rect 107 -1192 108 -1190
rect 114 -1186 115 -1184
rect 117 -1192 118 -1190
rect 121 -1186 122 -1184
rect 121 -1192 122 -1190
rect 128 -1186 129 -1184
rect 128 -1192 129 -1190
rect 135 -1186 136 -1184
rect 135 -1192 136 -1190
rect 142 -1186 143 -1184
rect 145 -1186 146 -1184
rect 145 -1192 146 -1190
rect 149 -1186 150 -1184
rect 152 -1186 153 -1184
rect 149 -1192 150 -1190
rect 152 -1192 153 -1190
rect 156 -1186 157 -1184
rect 159 -1186 160 -1184
rect 163 -1186 164 -1184
rect 163 -1192 164 -1190
rect 170 -1186 171 -1184
rect 170 -1192 171 -1190
rect 173 -1192 174 -1190
rect 177 -1186 178 -1184
rect 177 -1192 178 -1190
rect 184 -1186 185 -1184
rect 184 -1192 185 -1190
rect 194 -1186 195 -1184
rect 191 -1192 192 -1190
rect 198 -1186 199 -1184
rect 198 -1192 199 -1190
rect 205 -1186 206 -1184
rect 208 -1186 209 -1184
rect 215 -1192 216 -1190
rect 219 -1186 220 -1184
rect 219 -1192 220 -1190
rect 226 -1186 227 -1184
rect 226 -1192 227 -1190
rect 233 -1186 234 -1184
rect 236 -1186 237 -1184
rect 240 -1186 241 -1184
rect 240 -1192 241 -1190
rect 247 -1186 248 -1184
rect 247 -1192 248 -1190
rect 254 -1186 255 -1184
rect 254 -1192 255 -1190
rect 261 -1186 262 -1184
rect 261 -1192 262 -1190
rect 268 -1186 269 -1184
rect 268 -1192 269 -1190
rect 275 -1192 276 -1190
rect 282 -1186 283 -1184
rect 282 -1192 283 -1190
rect 289 -1186 290 -1184
rect 289 -1192 290 -1190
rect 296 -1186 297 -1184
rect 296 -1192 297 -1190
rect 303 -1186 304 -1184
rect 303 -1192 304 -1190
rect 306 -1192 307 -1190
rect 310 -1186 311 -1184
rect 310 -1192 311 -1190
rect 317 -1186 318 -1184
rect 320 -1186 321 -1184
rect 320 -1192 321 -1190
rect 324 -1186 325 -1184
rect 327 -1192 328 -1190
rect 331 -1186 332 -1184
rect 334 -1192 335 -1190
rect 338 -1186 339 -1184
rect 341 -1192 342 -1190
rect 348 -1186 349 -1184
rect 345 -1192 346 -1190
rect 348 -1192 349 -1190
rect 352 -1186 353 -1184
rect 352 -1192 353 -1190
rect 359 -1186 360 -1184
rect 359 -1192 360 -1190
rect 366 -1186 367 -1184
rect 366 -1192 367 -1190
rect 373 -1186 374 -1184
rect 373 -1192 374 -1190
rect 380 -1186 381 -1184
rect 380 -1192 381 -1190
rect 387 -1186 388 -1184
rect 390 -1186 391 -1184
rect 387 -1192 388 -1190
rect 390 -1192 391 -1190
rect 394 -1186 395 -1184
rect 394 -1192 395 -1190
rect 401 -1186 402 -1184
rect 401 -1192 402 -1190
rect 408 -1186 409 -1184
rect 408 -1192 409 -1190
rect 415 -1186 416 -1184
rect 415 -1192 416 -1190
rect 422 -1186 423 -1184
rect 422 -1192 423 -1190
rect 429 -1186 430 -1184
rect 429 -1192 430 -1190
rect 436 -1192 437 -1190
rect 443 -1186 444 -1184
rect 446 -1186 447 -1184
rect 443 -1192 444 -1190
rect 446 -1192 447 -1190
rect 450 -1186 451 -1184
rect 450 -1192 451 -1190
rect 453 -1192 454 -1190
rect 457 -1186 458 -1184
rect 457 -1192 458 -1190
rect 464 -1186 465 -1184
rect 467 -1192 468 -1190
rect 471 -1186 472 -1184
rect 471 -1192 472 -1190
rect 478 -1186 479 -1184
rect 478 -1192 479 -1190
rect 485 -1186 486 -1184
rect 485 -1192 486 -1190
rect 492 -1186 493 -1184
rect 492 -1192 493 -1190
rect 499 -1186 500 -1184
rect 499 -1192 500 -1190
rect 506 -1186 507 -1184
rect 506 -1192 507 -1190
rect 513 -1186 514 -1184
rect 513 -1192 514 -1190
rect 520 -1186 521 -1184
rect 520 -1192 521 -1190
rect 530 -1186 531 -1184
rect 530 -1192 531 -1190
rect 534 -1186 535 -1184
rect 534 -1192 535 -1190
rect 544 -1186 545 -1184
rect 541 -1192 542 -1190
rect 548 -1186 549 -1184
rect 548 -1192 549 -1190
rect 555 -1186 556 -1184
rect 555 -1192 556 -1190
rect 562 -1186 563 -1184
rect 562 -1192 563 -1190
rect 569 -1186 570 -1184
rect 569 -1192 570 -1190
rect 576 -1186 577 -1184
rect 576 -1192 577 -1190
rect 583 -1186 584 -1184
rect 583 -1192 584 -1190
rect 590 -1186 591 -1184
rect 590 -1192 591 -1190
rect 597 -1186 598 -1184
rect 597 -1192 598 -1190
rect 604 -1186 605 -1184
rect 604 -1192 605 -1190
rect 611 -1186 612 -1184
rect 611 -1192 612 -1190
rect 618 -1186 619 -1184
rect 618 -1192 619 -1190
rect 625 -1186 626 -1184
rect 625 -1192 626 -1190
rect 632 -1186 633 -1184
rect 632 -1192 633 -1190
rect 639 -1186 640 -1184
rect 639 -1192 640 -1190
rect 646 -1186 647 -1184
rect 646 -1192 647 -1190
rect 656 -1186 657 -1184
rect 660 -1186 661 -1184
rect 660 -1192 661 -1190
rect 667 -1186 668 -1184
rect 674 -1186 675 -1184
rect 677 -1186 678 -1184
rect 674 -1192 675 -1190
rect 681 -1186 682 -1184
rect 681 -1192 682 -1190
rect 688 -1186 689 -1184
rect 688 -1192 689 -1190
rect 702 -1186 703 -1184
rect 702 -1192 703 -1190
rect 709 -1186 710 -1184
rect 709 -1192 710 -1190
rect 2 -1257 3 -1255
rect 2 -1263 3 -1261
rect 9 -1257 10 -1255
rect 9 -1263 10 -1261
rect 16 -1257 17 -1255
rect 16 -1263 17 -1261
rect 23 -1257 24 -1255
rect 23 -1263 24 -1261
rect 30 -1257 31 -1255
rect 30 -1263 31 -1261
rect 37 -1257 38 -1255
rect 37 -1263 38 -1261
rect 44 -1263 45 -1261
rect 47 -1263 48 -1261
rect 54 -1257 55 -1255
rect 58 -1257 59 -1255
rect 61 -1263 62 -1261
rect 65 -1257 66 -1255
rect 65 -1263 66 -1261
rect 75 -1257 76 -1255
rect 72 -1263 73 -1261
rect 79 -1257 80 -1255
rect 79 -1263 80 -1261
rect 86 -1257 87 -1255
rect 86 -1263 87 -1261
rect 93 -1257 94 -1255
rect 93 -1263 94 -1261
rect 100 -1257 101 -1255
rect 103 -1263 104 -1261
rect 107 -1257 108 -1255
rect 110 -1257 111 -1255
rect 114 -1257 115 -1255
rect 114 -1263 115 -1261
rect 124 -1257 125 -1255
rect 121 -1263 122 -1261
rect 128 -1257 129 -1255
rect 128 -1263 129 -1261
rect 135 -1257 136 -1255
rect 135 -1263 136 -1261
rect 142 -1257 143 -1255
rect 145 -1263 146 -1261
rect 149 -1257 150 -1255
rect 149 -1263 150 -1261
rect 156 -1257 157 -1255
rect 156 -1263 157 -1261
rect 166 -1257 167 -1255
rect 163 -1263 164 -1261
rect 170 -1257 171 -1255
rect 170 -1263 171 -1261
rect 177 -1257 178 -1255
rect 177 -1263 178 -1261
rect 180 -1263 181 -1261
rect 187 -1257 188 -1255
rect 184 -1263 185 -1261
rect 187 -1263 188 -1261
rect 194 -1257 195 -1255
rect 191 -1263 192 -1261
rect 194 -1263 195 -1261
rect 201 -1257 202 -1255
rect 205 -1257 206 -1255
rect 205 -1263 206 -1261
rect 212 -1257 213 -1255
rect 212 -1263 213 -1261
rect 215 -1263 216 -1261
rect 219 -1263 220 -1261
rect 222 -1263 223 -1261
rect 226 -1257 227 -1255
rect 229 -1257 230 -1255
rect 233 -1257 234 -1255
rect 233 -1263 234 -1261
rect 236 -1263 237 -1261
rect 240 -1257 241 -1255
rect 240 -1263 241 -1261
rect 247 -1257 248 -1255
rect 250 -1257 251 -1255
rect 247 -1263 248 -1261
rect 250 -1263 251 -1261
rect 254 -1257 255 -1255
rect 257 -1257 258 -1255
rect 254 -1263 255 -1261
rect 257 -1263 258 -1261
rect 261 -1257 262 -1255
rect 261 -1263 262 -1261
rect 268 -1257 269 -1255
rect 268 -1263 269 -1261
rect 271 -1263 272 -1261
rect 275 -1257 276 -1255
rect 275 -1263 276 -1261
rect 282 -1257 283 -1255
rect 282 -1263 283 -1261
rect 289 -1257 290 -1255
rect 289 -1263 290 -1261
rect 296 -1257 297 -1255
rect 296 -1263 297 -1261
rect 306 -1257 307 -1255
rect 303 -1263 304 -1261
rect 306 -1263 307 -1261
rect 310 -1257 311 -1255
rect 313 -1263 314 -1261
rect 317 -1257 318 -1255
rect 317 -1263 318 -1261
rect 324 -1257 325 -1255
rect 327 -1257 328 -1255
rect 324 -1263 325 -1261
rect 327 -1263 328 -1261
rect 331 -1257 332 -1255
rect 331 -1263 332 -1261
rect 338 -1257 339 -1255
rect 338 -1263 339 -1261
rect 345 -1257 346 -1255
rect 345 -1263 346 -1261
rect 352 -1257 353 -1255
rect 359 -1257 360 -1255
rect 359 -1263 360 -1261
rect 366 -1257 367 -1255
rect 366 -1263 367 -1261
rect 373 -1257 374 -1255
rect 373 -1263 374 -1261
rect 380 -1257 381 -1255
rect 383 -1257 384 -1255
rect 380 -1263 381 -1261
rect 383 -1263 384 -1261
rect 387 -1257 388 -1255
rect 387 -1263 388 -1261
rect 394 -1257 395 -1255
rect 397 -1257 398 -1255
rect 397 -1263 398 -1261
rect 401 -1257 402 -1255
rect 401 -1263 402 -1261
rect 408 -1257 409 -1255
rect 408 -1263 409 -1261
rect 415 -1257 416 -1255
rect 415 -1263 416 -1261
rect 422 -1257 423 -1255
rect 422 -1263 423 -1261
rect 429 -1257 430 -1255
rect 432 -1257 433 -1255
rect 432 -1263 433 -1261
rect 436 -1257 437 -1255
rect 436 -1263 437 -1261
rect 443 -1257 444 -1255
rect 443 -1263 444 -1261
rect 450 -1257 451 -1255
rect 453 -1257 454 -1255
rect 453 -1263 454 -1261
rect 457 -1257 458 -1255
rect 460 -1257 461 -1255
rect 460 -1263 461 -1261
rect 464 -1257 465 -1255
rect 464 -1263 465 -1261
rect 471 -1257 472 -1255
rect 471 -1263 472 -1261
rect 478 -1257 479 -1255
rect 478 -1263 479 -1261
rect 485 -1257 486 -1255
rect 485 -1263 486 -1261
rect 492 -1257 493 -1255
rect 495 -1263 496 -1261
rect 499 -1257 500 -1255
rect 499 -1263 500 -1261
rect 506 -1257 507 -1255
rect 506 -1263 507 -1261
rect 513 -1257 514 -1255
rect 513 -1263 514 -1261
rect 520 -1257 521 -1255
rect 520 -1263 521 -1261
rect 527 -1257 528 -1255
rect 527 -1263 528 -1261
rect 534 -1257 535 -1255
rect 534 -1263 535 -1261
rect 541 -1257 542 -1255
rect 541 -1263 542 -1261
rect 548 -1257 549 -1255
rect 548 -1263 549 -1261
rect 555 -1257 556 -1255
rect 555 -1263 556 -1261
rect 562 -1257 563 -1255
rect 562 -1263 563 -1261
rect 569 -1257 570 -1255
rect 569 -1263 570 -1261
rect 576 -1257 577 -1255
rect 576 -1263 577 -1261
rect 583 -1257 584 -1255
rect 583 -1263 584 -1261
rect 590 -1257 591 -1255
rect 590 -1263 591 -1261
rect 597 -1257 598 -1255
rect 597 -1263 598 -1261
rect 604 -1257 605 -1255
rect 604 -1263 605 -1261
rect 611 -1257 612 -1255
rect 611 -1263 612 -1261
rect 618 -1257 619 -1255
rect 618 -1263 619 -1261
rect 625 -1257 626 -1255
rect 625 -1263 626 -1261
rect 632 -1257 633 -1255
rect 632 -1263 633 -1261
rect 639 -1257 640 -1255
rect 639 -1263 640 -1261
rect 646 -1257 647 -1255
rect 646 -1263 647 -1261
rect 653 -1257 654 -1255
rect 653 -1263 654 -1261
rect 660 -1257 661 -1255
rect 660 -1263 661 -1261
rect 667 -1257 668 -1255
rect 667 -1263 668 -1261
rect 674 -1257 675 -1255
rect 674 -1263 675 -1261
rect 681 -1257 682 -1255
rect 681 -1263 682 -1261
rect 688 -1257 689 -1255
rect 688 -1263 689 -1261
rect 695 -1257 696 -1255
rect 695 -1263 696 -1261
rect 702 -1257 703 -1255
rect 705 -1257 706 -1255
rect 702 -1263 703 -1261
rect 705 -1263 706 -1261
rect 712 -1257 713 -1255
rect 712 -1263 713 -1261
rect 716 -1257 717 -1255
rect 716 -1263 717 -1261
rect 2 -1328 3 -1326
rect 2 -1334 3 -1332
rect 9 -1328 10 -1326
rect 9 -1334 10 -1332
rect 19 -1334 20 -1332
rect 23 -1328 24 -1326
rect 23 -1334 24 -1332
rect 33 -1334 34 -1332
rect 40 -1328 41 -1326
rect 44 -1328 45 -1326
rect 44 -1334 45 -1332
rect 51 -1328 52 -1326
rect 51 -1334 52 -1332
rect 58 -1328 59 -1326
rect 58 -1334 59 -1332
rect 65 -1328 66 -1326
rect 65 -1334 66 -1332
rect 72 -1328 73 -1326
rect 75 -1334 76 -1332
rect 82 -1328 83 -1326
rect 82 -1334 83 -1332
rect 86 -1328 87 -1326
rect 86 -1334 87 -1332
rect 93 -1328 94 -1326
rect 93 -1334 94 -1332
rect 100 -1328 101 -1326
rect 100 -1334 101 -1332
rect 107 -1328 108 -1326
rect 107 -1334 108 -1332
rect 114 -1328 115 -1326
rect 114 -1334 115 -1332
rect 121 -1328 122 -1326
rect 121 -1334 122 -1332
rect 131 -1328 132 -1326
rect 131 -1334 132 -1332
rect 135 -1328 136 -1326
rect 138 -1328 139 -1326
rect 138 -1334 139 -1332
rect 142 -1328 143 -1326
rect 142 -1334 143 -1332
rect 152 -1334 153 -1332
rect 156 -1328 157 -1326
rect 156 -1334 157 -1332
rect 163 -1328 164 -1326
rect 163 -1334 164 -1332
rect 170 -1334 171 -1332
rect 173 -1334 174 -1332
rect 177 -1328 178 -1326
rect 180 -1328 181 -1326
rect 177 -1334 178 -1332
rect 184 -1328 185 -1326
rect 184 -1334 185 -1332
rect 191 -1328 192 -1326
rect 191 -1334 192 -1332
rect 198 -1328 199 -1326
rect 198 -1334 199 -1332
rect 205 -1328 206 -1326
rect 208 -1328 209 -1326
rect 212 -1328 213 -1326
rect 212 -1334 213 -1332
rect 219 -1328 220 -1326
rect 219 -1334 220 -1332
rect 226 -1328 227 -1326
rect 226 -1334 227 -1332
rect 233 -1328 234 -1326
rect 236 -1328 237 -1326
rect 233 -1334 234 -1332
rect 240 -1328 241 -1326
rect 240 -1334 241 -1332
rect 247 -1328 248 -1326
rect 247 -1334 248 -1332
rect 254 -1328 255 -1326
rect 254 -1334 255 -1332
rect 261 -1328 262 -1326
rect 261 -1334 262 -1332
rect 268 -1328 269 -1326
rect 268 -1334 269 -1332
rect 275 -1328 276 -1326
rect 275 -1334 276 -1332
rect 282 -1328 283 -1326
rect 285 -1328 286 -1326
rect 282 -1334 283 -1332
rect 285 -1334 286 -1332
rect 289 -1328 290 -1326
rect 289 -1334 290 -1332
rect 296 -1328 297 -1326
rect 296 -1334 297 -1332
rect 299 -1334 300 -1332
rect 303 -1328 304 -1326
rect 306 -1328 307 -1326
rect 310 -1328 311 -1326
rect 310 -1334 311 -1332
rect 317 -1328 318 -1326
rect 317 -1334 318 -1332
rect 324 -1328 325 -1326
rect 324 -1334 325 -1332
rect 327 -1334 328 -1332
rect 331 -1328 332 -1326
rect 331 -1334 332 -1332
rect 338 -1334 339 -1332
rect 341 -1334 342 -1332
rect 345 -1328 346 -1326
rect 345 -1334 346 -1332
rect 352 -1328 353 -1326
rect 355 -1328 356 -1326
rect 352 -1334 353 -1332
rect 362 -1328 363 -1326
rect 362 -1334 363 -1332
rect 366 -1328 367 -1326
rect 369 -1328 370 -1326
rect 366 -1334 367 -1332
rect 369 -1334 370 -1332
rect 373 -1328 374 -1326
rect 380 -1328 381 -1326
rect 380 -1334 381 -1332
rect 383 -1334 384 -1332
rect 390 -1328 391 -1326
rect 387 -1334 388 -1332
rect 390 -1334 391 -1332
rect 394 -1328 395 -1326
rect 397 -1328 398 -1326
rect 397 -1334 398 -1332
rect 401 -1328 402 -1326
rect 401 -1334 402 -1332
rect 408 -1328 409 -1326
rect 408 -1334 409 -1332
rect 415 -1328 416 -1326
rect 415 -1334 416 -1332
rect 422 -1328 423 -1326
rect 422 -1334 423 -1332
rect 425 -1334 426 -1332
rect 429 -1328 430 -1326
rect 429 -1334 430 -1332
rect 436 -1328 437 -1326
rect 436 -1334 437 -1332
rect 443 -1328 444 -1326
rect 443 -1334 444 -1332
rect 450 -1328 451 -1326
rect 457 -1328 458 -1326
rect 457 -1334 458 -1332
rect 464 -1328 465 -1326
rect 474 -1328 475 -1326
rect 471 -1334 472 -1332
rect 474 -1334 475 -1332
rect 478 -1328 479 -1326
rect 481 -1334 482 -1332
rect 485 -1328 486 -1326
rect 485 -1334 486 -1332
rect 492 -1328 493 -1326
rect 492 -1334 493 -1332
rect 499 -1328 500 -1326
rect 502 -1328 503 -1326
rect 499 -1334 500 -1332
rect 506 -1328 507 -1326
rect 506 -1334 507 -1332
rect 513 -1328 514 -1326
rect 513 -1334 514 -1332
rect 520 -1328 521 -1326
rect 520 -1334 521 -1332
rect 527 -1328 528 -1326
rect 527 -1334 528 -1332
rect 534 -1328 535 -1326
rect 534 -1334 535 -1332
rect 541 -1328 542 -1326
rect 541 -1334 542 -1332
rect 548 -1328 549 -1326
rect 548 -1334 549 -1332
rect 555 -1328 556 -1326
rect 555 -1334 556 -1332
rect 562 -1328 563 -1326
rect 562 -1334 563 -1332
rect 569 -1328 570 -1326
rect 569 -1334 570 -1332
rect 576 -1328 577 -1326
rect 576 -1334 577 -1332
rect 583 -1328 584 -1326
rect 583 -1334 584 -1332
rect 590 -1328 591 -1326
rect 590 -1334 591 -1332
rect 597 -1328 598 -1326
rect 597 -1334 598 -1332
rect 604 -1328 605 -1326
rect 604 -1334 605 -1332
rect 611 -1328 612 -1326
rect 611 -1334 612 -1332
rect 618 -1328 619 -1326
rect 618 -1334 619 -1332
rect 625 -1328 626 -1326
rect 625 -1334 626 -1332
rect 632 -1328 633 -1326
rect 632 -1334 633 -1332
rect 639 -1328 640 -1326
rect 639 -1334 640 -1332
rect 646 -1334 647 -1332
rect 653 -1328 654 -1326
rect 653 -1334 654 -1332
rect 660 -1328 661 -1326
rect 667 -1328 668 -1326
rect 670 -1328 671 -1326
rect 670 -1334 671 -1332
rect 674 -1328 675 -1326
rect 674 -1334 675 -1332
rect 681 -1328 682 -1326
rect 681 -1334 682 -1332
rect 702 -1328 703 -1326
rect 702 -1334 703 -1332
rect 33 -1393 34 -1391
rect 37 -1387 38 -1385
rect 37 -1393 38 -1391
rect 44 -1387 45 -1385
rect 44 -1393 45 -1391
rect 51 -1387 52 -1385
rect 51 -1393 52 -1391
rect 58 -1387 59 -1385
rect 58 -1393 59 -1391
rect 65 -1387 66 -1385
rect 65 -1393 66 -1391
rect 72 -1387 73 -1385
rect 72 -1393 73 -1391
rect 79 -1387 80 -1385
rect 79 -1393 80 -1391
rect 86 -1387 87 -1385
rect 86 -1393 87 -1391
rect 93 -1387 94 -1385
rect 93 -1393 94 -1391
rect 100 -1387 101 -1385
rect 103 -1393 104 -1391
rect 107 -1387 108 -1385
rect 107 -1393 108 -1391
rect 114 -1387 115 -1385
rect 114 -1393 115 -1391
rect 121 -1387 122 -1385
rect 124 -1387 125 -1385
rect 128 -1387 129 -1385
rect 128 -1393 129 -1391
rect 135 -1387 136 -1385
rect 138 -1387 139 -1385
rect 138 -1393 139 -1391
rect 145 -1387 146 -1385
rect 145 -1393 146 -1391
rect 149 -1387 150 -1385
rect 149 -1393 150 -1391
rect 159 -1387 160 -1385
rect 156 -1393 157 -1391
rect 163 -1387 164 -1385
rect 163 -1393 164 -1391
rect 170 -1387 171 -1385
rect 170 -1393 171 -1391
rect 177 -1387 178 -1385
rect 177 -1393 178 -1391
rect 184 -1387 185 -1385
rect 184 -1393 185 -1391
rect 187 -1393 188 -1391
rect 191 -1387 192 -1385
rect 191 -1393 192 -1391
rect 198 -1387 199 -1385
rect 201 -1387 202 -1385
rect 201 -1393 202 -1391
rect 205 -1387 206 -1385
rect 208 -1387 209 -1385
rect 205 -1393 206 -1391
rect 212 -1387 213 -1385
rect 212 -1393 213 -1391
rect 219 -1387 220 -1385
rect 222 -1387 223 -1385
rect 219 -1393 220 -1391
rect 226 -1387 227 -1385
rect 226 -1393 227 -1391
rect 233 -1393 234 -1391
rect 236 -1393 237 -1391
rect 240 -1387 241 -1385
rect 243 -1387 244 -1385
rect 243 -1393 244 -1391
rect 247 -1387 248 -1385
rect 250 -1387 251 -1385
rect 247 -1393 248 -1391
rect 254 -1387 255 -1385
rect 254 -1393 255 -1391
rect 261 -1387 262 -1385
rect 261 -1393 262 -1391
rect 268 -1387 269 -1385
rect 268 -1393 269 -1391
rect 275 -1387 276 -1385
rect 275 -1393 276 -1391
rect 282 -1387 283 -1385
rect 285 -1387 286 -1385
rect 282 -1393 283 -1391
rect 285 -1393 286 -1391
rect 289 -1387 290 -1385
rect 289 -1393 290 -1391
rect 296 -1387 297 -1385
rect 296 -1393 297 -1391
rect 303 -1387 304 -1385
rect 303 -1393 304 -1391
rect 310 -1387 311 -1385
rect 310 -1393 311 -1391
rect 317 -1387 318 -1385
rect 317 -1393 318 -1391
rect 324 -1387 325 -1385
rect 324 -1393 325 -1391
rect 331 -1387 332 -1385
rect 331 -1393 332 -1391
rect 338 -1387 339 -1385
rect 338 -1393 339 -1391
rect 345 -1387 346 -1385
rect 348 -1387 349 -1385
rect 352 -1387 353 -1385
rect 352 -1393 353 -1391
rect 359 -1387 360 -1385
rect 362 -1387 363 -1385
rect 366 -1387 367 -1385
rect 369 -1387 370 -1385
rect 366 -1393 367 -1391
rect 369 -1393 370 -1391
rect 373 -1387 374 -1385
rect 373 -1393 374 -1391
rect 383 -1387 384 -1385
rect 380 -1393 381 -1391
rect 383 -1393 384 -1391
rect 390 -1387 391 -1385
rect 387 -1393 388 -1391
rect 394 -1387 395 -1385
rect 394 -1393 395 -1391
rect 404 -1387 405 -1385
rect 401 -1393 402 -1391
rect 404 -1393 405 -1391
rect 408 -1387 409 -1385
rect 408 -1393 409 -1391
rect 418 -1387 419 -1385
rect 418 -1393 419 -1391
rect 425 -1387 426 -1385
rect 425 -1393 426 -1391
rect 429 -1393 430 -1391
rect 432 -1393 433 -1391
rect 436 -1387 437 -1385
rect 436 -1393 437 -1391
rect 443 -1387 444 -1385
rect 443 -1393 444 -1391
rect 450 -1387 451 -1385
rect 450 -1393 451 -1391
rect 460 -1387 461 -1385
rect 460 -1393 461 -1391
rect 464 -1387 465 -1385
rect 464 -1393 465 -1391
rect 471 -1387 472 -1385
rect 471 -1393 472 -1391
rect 478 -1387 479 -1385
rect 481 -1387 482 -1385
rect 485 -1387 486 -1385
rect 485 -1393 486 -1391
rect 492 -1387 493 -1385
rect 492 -1393 493 -1391
rect 499 -1387 500 -1385
rect 499 -1393 500 -1391
rect 506 -1387 507 -1385
rect 506 -1393 507 -1391
rect 513 -1387 514 -1385
rect 513 -1393 514 -1391
rect 520 -1387 521 -1385
rect 520 -1393 521 -1391
rect 527 -1387 528 -1385
rect 527 -1393 528 -1391
rect 534 -1387 535 -1385
rect 534 -1393 535 -1391
rect 541 -1387 542 -1385
rect 541 -1393 542 -1391
rect 548 -1387 549 -1385
rect 548 -1393 549 -1391
rect 555 -1387 556 -1385
rect 555 -1393 556 -1391
rect 562 -1387 563 -1385
rect 562 -1393 563 -1391
rect 569 -1387 570 -1385
rect 569 -1393 570 -1391
rect 576 -1387 577 -1385
rect 576 -1393 577 -1391
rect 583 -1387 584 -1385
rect 583 -1393 584 -1391
rect 590 -1387 591 -1385
rect 590 -1393 591 -1391
rect 600 -1387 601 -1385
rect 600 -1393 601 -1391
rect 604 -1387 605 -1385
rect 604 -1393 605 -1391
rect 611 -1387 612 -1385
rect 611 -1393 612 -1391
rect 621 -1387 622 -1385
rect 621 -1393 622 -1391
rect 625 -1387 626 -1385
rect 625 -1393 626 -1391
rect 635 -1393 636 -1391
rect 639 -1387 640 -1385
rect 639 -1393 640 -1391
rect 646 -1387 647 -1385
rect 646 -1393 647 -1391
rect 653 -1387 654 -1385
rect 656 -1387 657 -1385
rect 660 -1387 661 -1385
rect 660 -1393 661 -1391
rect 667 -1387 668 -1385
rect 667 -1393 668 -1391
rect 702 -1387 703 -1385
rect 705 -1393 706 -1391
rect 37 -1446 38 -1444
rect 37 -1452 38 -1450
rect 44 -1446 45 -1444
rect 44 -1452 45 -1450
rect 51 -1446 52 -1444
rect 51 -1452 52 -1450
rect 58 -1446 59 -1444
rect 58 -1452 59 -1450
rect 65 -1446 66 -1444
rect 65 -1452 66 -1450
rect 72 -1446 73 -1444
rect 72 -1452 73 -1450
rect 79 -1446 80 -1444
rect 79 -1452 80 -1450
rect 86 -1446 87 -1444
rect 86 -1452 87 -1450
rect 93 -1446 94 -1444
rect 93 -1452 94 -1450
rect 103 -1446 104 -1444
rect 107 -1446 108 -1444
rect 107 -1452 108 -1450
rect 117 -1446 118 -1444
rect 117 -1452 118 -1450
rect 121 -1446 122 -1444
rect 124 -1446 125 -1444
rect 128 -1446 129 -1444
rect 128 -1452 129 -1450
rect 135 -1446 136 -1444
rect 138 -1446 139 -1444
rect 135 -1452 136 -1450
rect 145 -1446 146 -1444
rect 142 -1452 143 -1450
rect 149 -1446 150 -1444
rect 149 -1452 150 -1450
rect 156 -1452 157 -1450
rect 159 -1452 160 -1450
rect 163 -1446 164 -1444
rect 163 -1452 164 -1450
rect 170 -1446 171 -1444
rect 170 -1452 171 -1450
rect 177 -1446 178 -1444
rect 177 -1452 178 -1450
rect 184 -1452 185 -1450
rect 191 -1446 192 -1444
rect 191 -1452 192 -1450
rect 198 -1452 199 -1450
rect 205 -1446 206 -1444
rect 205 -1452 206 -1450
rect 212 -1446 213 -1444
rect 215 -1446 216 -1444
rect 215 -1452 216 -1450
rect 219 -1446 220 -1444
rect 219 -1452 220 -1450
rect 226 -1446 227 -1444
rect 229 -1452 230 -1450
rect 233 -1446 234 -1444
rect 233 -1452 234 -1450
rect 240 -1446 241 -1444
rect 240 -1452 241 -1450
rect 243 -1452 244 -1450
rect 247 -1446 248 -1444
rect 247 -1452 248 -1450
rect 254 -1446 255 -1444
rect 254 -1452 255 -1450
rect 261 -1446 262 -1444
rect 261 -1452 262 -1450
rect 268 -1446 269 -1444
rect 271 -1446 272 -1444
rect 271 -1452 272 -1450
rect 275 -1446 276 -1444
rect 275 -1452 276 -1450
rect 282 -1446 283 -1444
rect 282 -1452 283 -1450
rect 289 -1446 290 -1444
rect 289 -1452 290 -1450
rect 296 -1446 297 -1444
rect 296 -1452 297 -1450
rect 303 -1446 304 -1444
rect 303 -1452 304 -1450
rect 310 -1446 311 -1444
rect 310 -1452 311 -1450
rect 317 -1446 318 -1444
rect 317 -1452 318 -1450
rect 327 -1446 328 -1444
rect 324 -1452 325 -1450
rect 327 -1452 328 -1450
rect 331 -1446 332 -1444
rect 331 -1452 332 -1450
rect 338 -1446 339 -1444
rect 338 -1452 339 -1450
rect 345 -1446 346 -1444
rect 345 -1452 346 -1450
rect 355 -1446 356 -1444
rect 359 -1446 360 -1444
rect 359 -1452 360 -1450
rect 366 -1446 367 -1444
rect 369 -1446 370 -1444
rect 373 -1446 374 -1444
rect 376 -1446 377 -1444
rect 380 -1446 381 -1444
rect 380 -1452 381 -1450
rect 387 -1446 388 -1444
rect 390 -1446 391 -1444
rect 387 -1452 388 -1450
rect 390 -1452 391 -1450
rect 394 -1446 395 -1444
rect 397 -1446 398 -1444
rect 401 -1446 402 -1444
rect 401 -1452 402 -1450
rect 408 -1446 409 -1444
rect 408 -1452 409 -1450
rect 415 -1446 416 -1444
rect 415 -1452 416 -1450
rect 422 -1446 423 -1444
rect 422 -1452 423 -1450
rect 429 -1446 430 -1444
rect 429 -1452 430 -1450
rect 436 -1446 437 -1444
rect 439 -1446 440 -1444
rect 439 -1452 440 -1450
rect 443 -1446 444 -1444
rect 446 -1446 447 -1444
rect 443 -1452 444 -1450
rect 446 -1452 447 -1450
rect 450 -1446 451 -1444
rect 453 -1446 454 -1444
rect 457 -1446 458 -1444
rect 457 -1452 458 -1450
rect 464 -1446 465 -1444
rect 464 -1452 465 -1450
rect 471 -1446 472 -1444
rect 471 -1452 472 -1450
rect 478 -1452 479 -1450
rect 485 -1446 486 -1444
rect 485 -1452 486 -1450
rect 492 -1446 493 -1444
rect 492 -1452 493 -1450
rect 499 -1446 500 -1444
rect 499 -1452 500 -1450
rect 506 -1446 507 -1444
rect 506 -1452 507 -1450
rect 513 -1446 514 -1444
rect 513 -1452 514 -1450
rect 520 -1446 521 -1444
rect 520 -1452 521 -1450
rect 527 -1446 528 -1444
rect 527 -1452 528 -1450
rect 534 -1446 535 -1444
rect 534 -1452 535 -1450
rect 541 -1446 542 -1444
rect 541 -1452 542 -1450
rect 548 -1446 549 -1444
rect 551 -1446 552 -1444
rect 555 -1446 556 -1444
rect 555 -1452 556 -1450
rect 565 -1446 566 -1444
rect 562 -1452 563 -1450
rect 565 -1452 566 -1450
rect 569 -1452 570 -1450
rect 572 -1452 573 -1450
rect 576 -1446 577 -1444
rect 576 -1452 577 -1450
rect 583 -1446 584 -1444
rect 583 -1452 584 -1450
rect 590 -1446 591 -1444
rect 590 -1452 591 -1450
rect 597 -1446 598 -1444
rect 597 -1452 598 -1450
rect 604 -1446 605 -1444
rect 604 -1452 605 -1450
rect 646 -1446 647 -1444
rect 705 -1446 706 -1444
rect 702 -1452 703 -1450
rect 712 -1452 713 -1450
rect 16 -1499 17 -1497
rect 16 -1505 17 -1503
rect 23 -1505 24 -1503
rect 30 -1499 31 -1497
rect 30 -1505 31 -1503
rect 37 -1499 38 -1497
rect 37 -1505 38 -1503
rect 44 -1499 45 -1497
rect 51 -1499 52 -1497
rect 51 -1505 52 -1503
rect 54 -1505 55 -1503
rect 58 -1499 59 -1497
rect 58 -1505 59 -1503
rect 65 -1499 66 -1497
rect 65 -1505 66 -1503
rect 72 -1499 73 -1497
rect 72 -1505 73 -1503
rect 79 -1499 80 -1497
rect 79 -1505 80 -1503
rect 86 -1499 87 -1497
rect 89 -1505 90 -1503
rect 93 -1499 94 -1497
rect 93 -1505 94 -1503
rect 100 -1499 101 -1497
rect 100 -1505 101 -1503
rect 107 -1499 108 -1497
rect 110 -1499 111 -1497
rect 114 -1499 115 -1497
rect 114 -1505 115 -1503
rect 124 -1499 125 -1497
rect 121 -1505 122 -1503
rect 128 -1499 129 -1497
rect 128 -1505 129 -1503
rect 135 -1499 136 -1497
rect 135 -1505 136 -1503
rect 142 -1499 143 -1497
rect 142 -1505 143 -1503
rect 149 -1505 150 -1503
rect 152 -1505 153 -1503
rect 156 -1499 157 -1497
rect 156 -1505 157 -1503
rect 163 -1499 164 -1497
rect 166 -1499 167 -1497
rect 170 -1505 171 -1503
rect 173 -1505 174 -1503
rect 177 -1499 178 -1497
rect 180 -1499 181 -1497
rect 180 -1505 181 -1503
rect 184 -1505 185 -1503
rect 187 -1505 188 -1503
rect 191 -1499 192 -1497
rect 191 -1505 192 -1503
rect 198 -1499 199 -1497
rect 198 -1505 199 -1503
rect 205 -1505 206 -1503
rect 208 -1505 209 -1503
rect 212 -1499 213 -1497
rect 212 -1505 213 -1503
rect 219 -1499 220 -1497
rect 219 -1505 220 -1503
rect 226 -1499 227 -1497
rect 229 -1505 230 -1503
rect 233 -1499 234 -1497
rect 236 -1505 237 -1503
rect 240 -1499 241 -1497
rect 240 -1505 241 -1503
rect 250 -1499 251 -1497
rect 247 -1505 248 -1503
rect 254 -1499 255 -1497
rect 254 -1505 255 -1503
rect 261 -1499 262 -1497
rect 261 -1505 262 -1503
rect 268 -1499 269 -1497
rect 271 -1499 272 -1497
rect 275 -1499 276 -1497
rect 275 -1505 276 -1503
rect 282 -1499 283 -1497
rect 282 -1505 283 -1503
rect 289 -1499 290 -1497
rect 292 -1499 293 -1497
rect 289 -1505 290 -1503
rect 292 -1505 293 -1503
rect 296 -1499 297 -1497
rect 296 -1505 297 -1503
rect 306 -1499 307 -1497
rect 303 -1505 304 -1503
rect 310 -1499 311 -1497
rect 310 -1505 311 -1503
rect 313 -1505 314 -1503
rect 317 -1505 318 -1503
rect 320 -1505 321 -1503
rect 324 -1499 325 -1497
rect 331 -1499 332 -1497
rect 331 -1505 332 -1503
rect 338 -1499 339 -1497
rect 338 -1505 339 -1503
rect 345 -1499 346 -1497
rect 345 -1505 346 -1503
rect 352 -1499 353 -1497
rect 352 -1505 353 -1503
rect 359 -1499 360 -1497
rect 359 -1505 360 -1503
rect 366 -1499 367 -1497
rect 369 -1499 370 -1497
rect 373 -1499 374 -1497
rect 373 -1505 374 -1503
rect 380 -1499 381 -1497
rect 380 -1505 381 -1503
rect 387 -1499 388 -1497
rect 387 -1505 388 -1503
rect 394 -1499 395 -1497
rect 394 -1505 395 -1503
rect 401 -1499 402 -1497
rect 401 -1505 402 -1503
rect 408 -1499 409 -1497
rect 408 -1505 409 -1503
rect 415 -1499 416 -1497
rect 415 -1505 416 -1503
rect 425 -1499 426 -1497
rect 422 -1505 423 -1503
rect 429 -1499 430 -1497
rect 432 -1499 433 -1497
rect 429 -1505 430 -1503
rect 436 -1499 437 -1497
rect 436 -1505 437 -1503
rect 443 -1499 444 -1497
rect 443 -1505 444 -1503
rect 450 -1499 451 -1497
rect 450 -1505 451 -1503
rect 457 -1499 458 -1497
rect 457 -1505 458 -1503
rect 464 -1499 465 -1497
rect 464 -1505 465 -1503
rect 471 -1499 472 -1497
rect 471 -1505 472 -1503
rect 478 -1499 479 -1497
rect 485 -1499 486 -1497
rect 485 -1505 486 -1503
rect 492 -1499 493 -1497
rect 492 -1505 493 -1503
rect 499 -1499 500 -1497
rect 499 -1505 500 -1503
rect 506 -1499 507 -1497
rect 506 -1505 507 -1503
rect 513 -1499 514 -1497
rect 513 -1505 514 -1503
rect 520 -1499 521 -1497
rect 520 -1505 521 -1503
rect 527 -1499 528 -1497
rect 527 -1505 528 -1503
rect 534 -1499 535 -1497
rect 534 -1505 535 -1503
rect 541 -1499 542 -1497
rect 541 -1505 542 -1503
rect 548 -1499 549 -1497
rect 548 -1505 549 -1503
rect 555 -1499 556 -1497
rect 555 -1505 556 -1503
rect 562 -1499 563 -1497
rect 565 -1499 566 -1497
rect 562 -1505 563 -1503
rect 565 -1505 566 -1503
rect 569 -1499 570 -1497
rect 569 -1505 570 -1503
rect 576 -1499 577 -1497
rect 576 -1505 577 -1503
rect 579 -1505 580 -1503
rect 583 -1499 584 -1497
rect 583 -1505 584 -1503
rect 590 -1499 591 -1497
rect 590 -1505 591 -1503
rect 51 -1548 52 -1546
rect 51 -1554 52 -1552
rect 58 -1548 59 -1546
rect 65 -1548 66 -1546
rect 65 -1554 66 -1552
rect 72 -1554 73 -1552
rect 75 -1554 76 -1552
rect 79 -1548 80 -1546
rect 79 -1554 80 -1552
rect 86 -1548 87 -1546
rect 86 -1554 87 -1552
rect 96 -1548 97 -1546
rect 96 -1554 97 -1552
rect 103 -1554 104 -1552
rect 110 -1548 111 -1546
rect 107 -1554 108 -1552
rect 114 -1548 115 -1546
rect 114 -1554 115 -1552
rect 121 -1548 122 -1546
rect 121 -1554 122 -1552
rect 128 -1548 129 -1546
rect 128 -1554 129 -1552
rect 135 -1548 136 -1546
rect 135 -1554 136 -1552
rect 142 -1548 143 -1546
rect 142 -1554 143 -1552
rect 152 -1548 153 -1546
rect 149 -1554 150 -1552
rect 152 -1554 153 -1552
rect 156 -1548 157 -1546
rect 156 -1554 157 -1552
rect 159 -1554 160 -1552
rect 163 -1548 164 -1546
rect 163 -1554 164 -1552
rect 170 -1548 171 -1546
rect 173 -1554 174 -1552
rect 177 -1548 178 -1546
rect 177 -1554 178 -1552
rect 184 -1548 185 -1546
rect 184 -1554 185 -1552
rect 191 -1554 192 -1552
rect 194 -1554 195 -1552
rect 198 -1548 199 -1546
rect 201 -1548 202 -1546
rect 205 -1548 206 -1546
rect 205 -1554 206 -1552
rect 212 -1548 213 -1546
rect 212 -1554 213 -1552
rect 222 -1554 223 -1552
rect 229 -1548 230 -1546
rect 236 -1548 237 -1546
rect 236 -1554 237 -1552
rect 240 -1548 241 -1546
rect 240 -1554 241 -1552
rect 243 -1554 244 -1552
rect 247 -1548 248 -1546
rect 247 -1554 248 -1552
rect 254 -1548 255 -1546
rect 254 -1554 255 -1552
rect 261 -1548 262 -1546
rect 261 -1554 262 -1552
rect 268 -1548 269 -1546
rect 268 -1554 269 -1552
rect 275 -1548 276 -1546
rect 275 -1554 276 -1552
rect 282 -1548 283 -1546
rect 285 -1554 286 -1552
rect 292 -1554 293 -1552
rect 296 -1548 297 -1546
rect 296 -1554 297 -1552
rect 303 -1548 304 -1546
rect 303 -1554 304 -1552
rect 310 -1548 311 -1546
rect 310 -1554 311 -1552
rect 317 -1548 318 -1546
rect 317 -1554 318 -1552
rect 327 -1548 328 -1546
rect 327 -1554 328 -1552
rect 331 -1548 332 -1546
rect 331 -1554 332 -1552
rect 338 -1548 339 -1546
rect 338 -1554 339 -1552
rect 345 -1548 346 -1546
rect 345 -1554 346 -1552
rect 352 -1548 353 -1546
rect 352 -1554 353 -1552
rect 359 -1548 360 -1546
rect 359 -1554 360 -1552
rect 369 -1548 370 -1546
rect 366 -1554 367 -1552
rect 369 -1554 370 -1552
rect 373 -1548 374 -1546
rect 373 -1554 374 -1552
rect 380 -1548 381 -1546
rect 383 -1548 384 -1546
rect 380 -1554 381 -1552
rect 387 -1548 388 -1546
rect 387 -1554 388 -1552
rect 394 -1548 395 -1546
rect 394 -1554 395 -1552
rect 401 -1548 402 -1546
rect 401 -1554 402 -1552
rect 408 -1548 409 -1546
rect 408 -1554 409 -1552
rect 415 -1554 416 -1552
rect 425 -1548 426 -1546
rect 422 -1554 423 -1552
rect 429 -1548 430 -1546
rect 429 -1554 430 -1552
rect 436 -1548 437 -1546
rect 436 -1554 437 -1552
rect 443 -1548 444 -1546
rect 443 -1554 444 -1552
rect 450 -1548 451 -1546
rect 450 -1554 451 -1552
rect 457 -1548 458 -1546
rect 457 -1554 458 -1552
rect 464 -1548 465 -1546
rect 464 -1554 465 -1552
rect 474 -1548 475 -1546
rect 478 -1548 479 -1546
rect 478 -1554 479 -1552
rect 488 -1548 489 -1546
rect 492 -1548 493 -1546
rect 492 -1554 493 -1552
rect 499 -1548 500 -1546
rect 499 -1554 500 -1552
rect 502 -1554 503 -1552
rect 506 -1548 507 -1546
rect 506 -1554 507 -1552
rect 513 -1548 514 -1546
rect 513 -1554 514 -1552
rect 520 -1548 521 -1546
rect 520 -1554 521 -1552
rect 527 -1548 528 -1546
rect 527 -1554 528 -1552
rect 586 -1554 587 -1552
rect 590 -1548 591 -1546
rect 590 -1554 591 -1552
rect 75 -1591 76 -1589
rect 79 -1585 80 -1583
rect 79 -1591 80 -1589
rect 128 -1585 129 -1583
rect 128 -1591 129 -1589
rect 135 -1585 136 -1583
rect 135 -1591 136 -1589
rect 142 -1585 143 -1583
rect 145 -1591 146 -1589
rect 152 -1585 153 -1583
rect 152 -1591 153 -1589
rect 159 -1585 160 -1583
rect 156 -1591 157 -1589
rect 163 -1585 164 -1583
rect 163 -1591 164 -1589
rect 170 -1585 171 -1583
rect 170 -1591 171 -1589
rect 177 -1585 178 -1583
rect 177 -1591 178 -1589
rect 184 -1585 185 -1583
rect 184 -1591 185 -1589
rect 191 -1585 192 -1583
rect 194 -1585 195 -1583
rect 191 -1591 192 -1589
rect 194 -1591 195 -1589
rect 198 -1585 199 -1583
rect 201 -1585 202 -1583
rect 205 -1591 206 -1589
rect 208 -1591 209 -1589
rect 212 -1585 213 -1583
rect 212 -1591 213 -1589
rect 219 -1585 220 -1583
rect 222 -1585 223 -1583
rect 226 -1585 227 -1583
rect 229 -1585 230 -1583
rect 226 -1591 227 -1589
rect 233 -1585 234 -1583
rect 233 -1591 234 -1589
rect 240 -1591 241 -1589
rect 243 -1591 244 -1589
rect 247 -1585 248 -1583
rect 247 -1591 248 -1589
rect 254 -1585 255 -1583
rect 254 -1591 255 -1589
rect 261 -1585 262 -1583
rect 261 -1591 262 -1589
rect 271 -1585 272 -1583
rect 268 -1591 269 -1589
rect 275 -1585 276 -1583
rect 275 -1591 276 -1589
rect 282 -1585 283 -1583
rect 282 -1591 283 -1589
rect 289 -1585 290 -1583
rect 289 -1591 290 -1589
rect 296 -1585 297 -1583
rect 296 -1591 297 -1589
rect 303 -1585 304 -1583
rect 303 -1591 304 -1589
rect 313 -1585 314 -1583
rect 310 -1591 311 -1589
rect 317 -1585 318 -1583
rect 317 -1591 318 -1589
rect 320 -1591 321 -1589
rect 324 -1585 325 -1583
rect 324 -1591 325 -1589
rect 331 -1585 332 -1583
rect 331 -1591 332 -1589
rect 338 -1591 339 -1589
rect 345 -1591 346 -1589
rect 352 -1585 353 -1583
rect 352 -1591 353 -1589
rect 359 -1585 360 -1583
rect 359 -1591 360 -1589
rect 366 -1585 367 -1583
rect 369 -1585 370 -1583
rect 369 -1591 370 -1589
rect 373 -1585 374 -1583
rect 373 -1591 374 -1589
rect 380 -1585 381 -1583
rect 390 -1585 391 -1583
rect 387 -1591 388 -1589
rect 394 -1585 395 -1583
rect 394 -1591 395 -1589
rect 401 -1585 402 -1583
rect 401 -1591 402 -1589
rect 422 -1591 423 -1589
rect 429 -1585 430 -1583
rect 429 -1591 430 -1589
rect 436 -1585 437 -1583
rect 436 -1591 437 -1589
rect 464 -1585 465 -1583
rect 464 -1591 465 -1589
rect 471 -1585 472 -1583
rect 471 -1591 472 -1589
rect 485 -1585 486 -1583
rect 485 -1591 486 -1589
rect 492 -1585 493 -1583
rect 492 -1591 493 -1589
rect 506 -1591 507 -1589
rect 513 -1585 514 -1583
rect 513 -1591 514 -1589
rect 33 -1624 34 -1622
rect 72 -1618 73 -1616
rect 72 -1624 73 -1622
rect 82 -1618 83 -1616
rect 89 -1618 90 -1616
rect 86 -1624 87 -1622
rect 89 -1624 90 -1622
rect 93 -1618 94 -1616
rect 93 -1624 94 -1622
rect 100 -1624 101 -1622
rect 114 -1618 115 -1616
rect 114 -1624 115 -1622
rect 121 -1624 122 -1622
rect 124 -1624 125 -1622
rect 131 -1618 132 -1616
rect 135 -1618 136 -1616
rect 135 -1624 136 -1622
rect 142 -1618 143 -1616
rect 142 -1624 143 -1622
rect 152 -1618 153 -1616
rect 149 -1624 150 -1622
rect 156 -1618 157 -1616
rect 156 -1624 157 -1622
rect 163 -1618 164 -1616
rect 163 -1624 164 -1622
rect 170 -1618 171 -1616
rect 170 -1624 171 -1622
rect 177 -1624 178 -1622
rect 180 -1624 181 -1622
rect 191 -1618 192 -1616
rect 201 -1618 202 -1616
rect 198 -1624 199 -1622
rect 205 -1618 206 -1616
rect 205 -1624 206 -1622
rect 215 -1618 216 -1616
rect 212 -1624 213 -1622
rect 215 -1624 216 -1622
rect 219 -1618 220 -1616
rect 219 -1624 220 -1622
rect 226 -1618 227 -1616
rect 226 -1624 227 -1622
rect 236 -1618 237 -1616
rect 236 -1624 237 -1622
rect 240 -1618 241 -1616
rect 243 -1618 244 -1616
rect 240 -1624 241 -1622
rect 250 -1618 251 -1616
rect 254 -1618 255 -1616
rect 254 -1624 255 -1622
rect 261 -1618 262 -1616
rect 264 -1624 265 -1622
rect 268 -1618 269 -1616
rect 275 -1618 276 -1616
rect 278 -1618 279 -1616
rect 275 -1624 276 -1622
rect 278 -1624 279 -1622
rect 282 -1618 283 -1616
rect 289 -1618 290 -1616
rect 289 -1624 290 -1622
rect 296 -1618 297 -1616
rect 299 -1618 300 -1616
rect 296 -1624 297 -1622
rect 303 -1618 304 -1616
rect 303 -1624 304 -1622
rect 310 -1618 311 -1616
rect 310 -1624 311 -1622
rect 317 -1618 318 -1616
rect 317 -1624 318 -1622
rect 324 -1618 325 -1616
rect 324 -1624 325 -1622
rect 334 -1618 335 -1616
rect 334 -1624 335 -1622
rect 338 -1618 339 -1616
rect 341 -1618 342 -1616
rect 345 -1618 346 -1616
rect 345 -1624 346 -1622
rect 352 -1618 353 -1616
rect 352 -1624 353 -1622
rect 359 -1618 360 -1616
rect 359 -1624 360 -1622
rect 366 -1618 367 -1616
rect 366 -1624 367 -1622
rect 380 -1618 381 -1616
rect 383 -1618 384 -1616
rect 387 -1618 388 -1616
rect 387 -1624 388 -1622
rect 394 -1618 395 -1616
rect 394 -1624 395 -1622
rect 443 -1618 444 -1616
rect 443 -1624 444 -1622
rect 467 -1624 468 -1622
rect 471 -1618 472 -1616
rect 471 -1624 472 -1622
rect 485 -1618 486 -1616
rect 488 -1624 489 -1622
rect 492 -1618 493 -1616
rect 492 -1624 493 -1622
rect 30 -1647 31 -1645
rect 37 -1647 38 -1645
rect 37 -1653 38 -1651
rect 44 -1647 45 -1645
rect 44 -1653 45 -1651
rect 51 -1647 52 -1645
rect 51 -1653 52 -1651
rect 58 -1647 59 -1645
rect 65 -1647 66 -1645
rect 65 -1653 66 -1651
rect 72 -1647 73 -1645
rect 72 -1653 73 -1651
rect 79 -1647 80 -1645
rect 79 -1653 80 -1651
rect 86 -1647 87 -1645
rect 86 -1653 87 -1651
rect 93 -1653 94 -1651
rect 96 -1653 97 -1651
rect 100 -1647 101 -1645
rect 100 -1653 101 -1651
rect 107 -1647 108 -1645
rect 110 -1647 111 -1645
rect 114 -1647 115 -1645
rect 114 -1653 115 -1651
rect 117 -1653 118 -1651
rect 124 -1647 125 -1645
rect 121 -1653 122 -1651
rect 124 -1653 125 -1651
rect 131 -1647 132 -1645
rect 128 -1653 129 -1651
rect 135 -1647 136 -1645
rect 138 -1647 139 -1645
rect 138 -1653 139 -1651
rect 145 -1647 146 -1645
rect 145 -1653 146 -1651
rect 149 -1647 150 -1645
rect 149 -1653 150 -1651
rect 156 -1647 157 -1645
rect 156 -1653 157 -1651
rect 163 -1647 164 -1645
rect 163 -1653 164 -1651
rect 170 -1647 171 -1645
rect 170 -1653 171 -1651
rect 177 -1647 178 -1645
rect 177 -1653 178 -1651
rect 184 -1653 185 -1651
rect 191 -1647 192 -1645
rect 191 -1653 192 -1651
rect 198 -1647 199 -1645
rect 201 -1647 202 -1645
rect 205 -1647 206 -1645
rect 205 -1653 206 -1651
rect 208 -1653 209 -1651
rect 212 -1653 213 -1651
rect 215 -1653 216 -1651
rect 219 -1647 220 -1645
rect 222 -1647 223 -1645
rect 219 -1653 220 -1651
rect 222 -1653 223 -1651
rect 226 -1647 227 -1645
rect 229 -1647 230 -1645
rect 226 -1653 227 -1651
rect 233 -1647 234 -1645
rect 236 -1653 237 -1651
rect 240 -1647 241 -1645
rect 240 -1653 241 -1651
rect 243 -1653 244 -1651
rect 247 -1647 248 -1645
rect 247 -1653 248 -1651
rect 254 -1647 255 -1645
rect 254 -1653 255 -1651
rect 261 -1647 262 -1645
rect 261 -1653 262 -1651
rect 271 -1647 272 -1645
rect 268 -1653 269 -1651
rect 271 -1653 272 -1651
rect 275 -1647 276 -1645
rect 275 -1653 276 -1651
rect 282 -1647 283 -1645
rect 282 -1653 283 -1651
rect 289 -1647 290 -1645
rect 289 -1653 290 -1651
rect 296 -1647 297 -1645
rect 296 -1653 297 -1651
rect 303 -1647 304 -1645
rect 310 -1647 311 -1645
rect 310 -1653 311 -1651
rect 317 -1647 318 -1645
rect 317 -1653 318 -1651
rect 327 -1647 328 -1645
rect 324 -1653 325 -1651
rect 331 -1647 332 -1645
rect 331 -1653 332 -1651
rect 338 -1647 339 -1645
rect 338 -1653 339 -1651
rect 345 -1647 346 -1645
rect 345 -1653 346 -1651
rect 352 -1647 353 -1645
rect 352 -1653 353 -1651
rect 359 -1647 360 -1645
rect 359 -1653 360 -1651
rect 366 -1647 367 -1645
rect 366 -1653 367 -1651
rect 373 -1647 374 -1645
rect 373 -1653 374 -1651
rect 380 -1647 381 -1645
rect 380 -1653 381 -1651
rect 387 -1647 388 -1645
rect 387 -1653 388 -1651
rect 394 -1647 395 -1645
rect 394 -1653 395 -1651
rect 401 -1647 402 -1645
rect 404 -1647 405 -1645
rect 2 -1688 3 -1686
rect 19 -1682 20 -1680
rect 23 -1682 24 -1680
rect 23 -1688 24 -1686
rect 33 -1688 34 -1686
rect 79 -1688 80 -1686
rect 103 -1682 104 -1680
rect 107 -1682 108 -1680
rect 107 -1688 108 -1686
rect 114 -1688 115 -1686
rect 121 -1682 122 -1680
rect 121 -1688 122 -1686
rect 131 -1688 132 -1686
rect 135 -1682 136 -1680
rect 135 -1688 136 -1686
rect 145 -1682 146 -1680
rect 149 -1682 150 -1680
rect 149 -1688 150 -1686
rect 156 -1682 157 -1680
rect 156 -1688 157 -1686
rect 163 -1682 164 -1680
rect 163 -1688 164 -1686
rect 170 -1688 171 -1686
rect 173 -1688 174 -1686
rect 177 -1688 178 -1686
rect 184 -1688 185 -1686
rect 191 -1682 192 -1680
rect 191 -1688 192 -1686
rect 198 -1682 199 -1680
rect 198 -1688 199 -1686
rect 205 -1682 206 -1680
rect 205 -1688 206 -1686
rect 212 -1682 213 -1680
rect 212 -1688 213 -1686
rect 222 -1682 223 -1680
rect 219 -1688 220 -1686
rect 226 -1682 227 -1680
rect 229 -1682 230 -1680
rect 226 -1688 227 -1686
rect 229 -1688 230 -1686
rect 233 -1682 234 -1680
rect 233 -1688 234 -1686
rect 240 -1682 241 -1680
rect 243 -1688 244 -1686
rect 247 -1682 248 -1680
rect 247 -1688 248 -1686
rect 254 -1688 255 -1686
rect 261 -1682 262 -1680
rect 264 -1688 265 -1686
rect 268 -1682 269 -1680
rect 268 -1688 269 -1686
rect 275 -1688 276 -1686
rect 285 -1682 286 -1680
rect 285 -1688 286 -1686
rect 289 -1688 290 -1686
rect 296 -1682 297 -1680
rect 296 -1688 297 -1686
rect 303 -1682 304 -1680
rect 303 -1688 304 -1686
rect 310 -1682 311 -1680
rect 310 -1688 311 -1686
rect 320 -1682 321 -1680
rect 317 -1688 318 -1686
rect 324 -1682 325 -1680
rect 324 -1688 325 -1686
rect 331 -1682 332 -1680
rect 331 -1688 332 -1686
rect 338 -1682 339 -1680
rect 338 -1688 339 -1686
rect 348 -1682 349 -1680
rect 352 -1682 353 -1680
rect 352 -1688 353 -1686
rect 359 -1688 360 -1686
rect 366 -1682 367 -1680
rect 373 -1682 374 -1680
rect 373 -1688 374 -1686
rect 380 -1682 381 -1680
rect 380 -1688 381 -1686
rect 390 -1682 391 -1680
rect 394 -1682 395 -1680
rect 394 -1688 395 -1686
rect 401 -1682 402 -1680
rect 401 -1688 402 -1686
rect 5 -1711 6 -1709
rect 9 -1705 10 -1703
rect 9 -1711 10 -1709
rect 16 -1705 17 -1703
rect 30 -1705 31 -1703
rect 79 -1705 80 -1703
rect 89 -1705 90 -1703
rect 96 -1705 97 -1703
rect 100 -1705 101 -1703
rect 117 -1705 118 -1703
rect 121 -1705 122 -1703
rect 128 -1705 129 -1703
rect 131 -1705 132 -1703
rect 128 -1711 129 -1709
rect 135 -1705 136 -1703
rect 135 -1711 136 -1709
rect 142 -1711 143 -1709
rect 152 -1711 153 -1709
rect 156 -1705 157 -1703
rect 156 -1711 157 -1709
rect 163 -1705 164 -1703
rect 163 -1711 164 -1709
rect 170 -1705 171 -1703
rect 170 -1711 171 -1709
rect 177 -1705 178 -1703
rect 177 -1711 178 -1709
rect 187 -1711 188 -1709
rect 194 -1705 195 -1703
rect 201 -1705 202 -1703
rect 201 -1711 202 -1709
rect 205 -1705 206 -1703
rect 205 -1711 206 -1709
rect 212 -1705 213 -1703
rect 212 -1711 213 -1709
rect 222 -1705 223 -1703
rect 219 -1711 220 -1709
rect 226 -1705 227 -1703
rect 226 -1711 227 -1709
rect 233 -1705 234 -1703
rect 233 -1711 234 -1709
rect 243 -1711 244 -1709
rect 257 -1705 258 -1703
rect 278 -1705 279 -1703
rect 285 -1705 286 -1703
rect 292 -1705 293 -1703
rect 296 -1705 297 -1703
rect 303 -1711 304 -1709
rect 310 -1705 311 -1703
rect 310 -1711 311 -1709
rect 317 -1711 318 -1709
rect 324 -1705 325 -1703
rect 324 -1711 325 -1709
rect 352 -1705 353 -1703
<< metal1 >>
rect 177 0 188 1
rect 198 0 206 1
rect 208 0 223 1
rect 240 0 248 1
rect 275 0 283 1
rect 289 0 300 1
rect 215 -2 234 -1
rect 243 -2 255 -1
rect 107 -13 111 -12
rect 142 -13 171 -12
rect 177 -13 195 -12
rect 219 -13 234 -12
rect 254 -13 269 -12
rect 289 -13 304 -12
rect 149 -15 160 -14
rect 163 -15 195 -14
rect 208 -15 220 -14
rect 226 -15 248 -14
rect 264 -15 276 -14
rect 282 -15 290 -14
rect 292 -15 311 -14
rect 184 -17 209 -16
rect 240 -17 248 -16
rect 296 -17 300 -16
rect 191 -19 199 -18
rect 198 -21 216 -20
rect 135 -32 146 -31
rect 152 -32 157 -31
rect 177 -32 227 -31
rect 233 -32 244 -31
rect 247 -32 262 -31
rect 282 -32 293 -31
rect 296 -32 304 -31
rect 310 -32 325 -31
rect 478 -32 486 -31
rect 579 -32 584 -31
rect 142 -34 181 -33
rect 191 -34 199 -33
rect 212 -34 220 -33
rect 240 -34 255 -33
rect 257 -34 269 -33
rect 285 -34 290 -33
rect 296 -34 304 -33
rect 317 -34 321 -33
rect 79 -45 83 -44
rect 135 -45 153 -44
rect 170 -45 174 -44
rect 184 -45 195 -44
rect 212 -45 216 -44
rect 219 -45 234 -44
rect 240 -45 283 -44
rect 289 -45 321 -44
rect 338 -45 346 -44
rect 352 -45 363 -44
rect 467 -45 472 -44
rect 478 -45 486 -44
rect 576 -45 584 -44
rect 177 -47 195 -46
rect 212 -47 244 -46
rect 247 -47 269 -46
rect 292 -47 318 -46
rect 184 -49 206 -48
rect 222 -49 227 -48
rect 233 -49 262 -48
rect 310 -49 325 -48
rect 229 -51 262 -50
rect 317 -51 342 -50
rect 247 -53 269 -52
rect 324 -53 335 -52
rect 250 -55 276 -54
rect 275 -57 283 -56
rect 142 -68 150 -67
rect 205 -68 213 -67
rect 219 -68 244 -67
rect 247 -68 262 -67
rect 268 -68 283 -67
rect 338 -68 346 -67
rect 474 -68 486 -67
rect 138 -70 220 -69
rect 226 -70 234 -69
rect 240 -70 290 -69
rect 345 -70 353 -69
rect 142 -72 164 -71
rect 166 -72 206 -71
rect 226 -72 276 -71
rect 278 -72 297 -71
rect 320 -72 353 -71
rect 149 -74 157 -73
rect 236 -74 290 -73
rect 296 -74 304 -73
rect 247 -76 255 -75
rect 261 -76 311 -75
rect 240 -78 255 -77
rect 268 -78 307 -77
rect 275 -80 318 -79
rect 128 -91 136 -90
rect 142 -91 146 -90
rect 149 -91 160 -90
rect 163 -91 227 -90
rect 233 -91 269 -90
rect 271 -91 360 -90
rect 397 -91 423 -90
rect 481 -91 486 -90
rect 576 -91 584 -90
rect 107 -93 143 -92
rect 152 -93 157 -92
rect 166 -93 171 -92
rect 177 -93 185 -92
rect 187 -93 199 -92
rect 205 -93 244 -92
rect 257 -93 262 -92
rect 289 -93 325 -92
rect 338 -93 349 -92
rect 352 -93 381 -92
rect 478 -93 486 -92
rect 576 -93 591 -92
rect 191 -95 202 -94
rect 219 -95 304 -94
rect 310 -95 367 -94
rect 478 -95 493 -94
rect 194 -97 227 -96
rect 240 -97 318 -96
rect 341 -97 346 -96
rect 212 -99 220 -98
rect 222 -99 353 -98
rect 212 -101 234 -100
rect 243 -101 248 -100
rect 250 -101 325 -100
rect 338 -101 346 -100
rect 254 -103 262 -102
rect 275 -103 311 -102
rect 317 -103 374 -102
rect 254 -105 321 -104
rect 296 -107 332 -106
rect 282 -109 297 -108
rect 180 -111 283 -110
rect 65 -122 108 -121
rect 131 -122 136 -121
rect 145 -122 171 -121
rect 173 -122 185 -121
rect 191 -122 206 -121
rect 208 -122 255 -121
rect 264 -122 279 -121
rect 289 -122 318 -121
rect 324 -122 339 -121
rect 359 -122 416 -121
rect 422 -122 444 -121
rect 478 -122 486 -121
rect 492 -122 500 -121
rect 576 -122 584 -121
rect 72 -124 101 -123
rect 107 -124 115 -123
rect 128 -124 136 -123
rect 149 -124 157 -123
rect 163 -124 237 -123
rect 243 -124 311 -123
rect 331 -124 423 -123
rect 86 -126 125 -125
rect 170 -126 209 -125
rect 219 -126 367 -125
rect 380 -126 430 -125
rect 93 -128 244 -127
rect 275 -128 374 -127
rect 387 -128 437 -127
rect 156 -130 220 -129
rect 222 -130 234 -129
rect 282 -130 311 -129
rect 334 -130 367 -129
rect 394 -130 402 -129
rect 177 -132 286 -131
rect 299 -132 360 -131
rect 184 -134 234 -133
rect 303 -134 374 -133
rect 191 -136 227 -135
rect 229 -136 290 -135
rect 352 -136 381 -135
rect 198 -138 213 -137
rect 222 -138 325 -137
rect 352 -138 395 -137
rect 198 -140 262 -139
rect 205 -142 248 -141
rect 261 -142 297 -141
rect 226 -144 269 -143
rect 240 -146 304 -145
rect 240 -148 276 -147
rect 257 -150 269 -149
rect 19 -161 27 -160
rect 65 -161 115 -160
rect 131 -161 160 -160
rect 163 -161 248 -160
rect 264 -161 311 -160
rect 317 -161 332 -160
rect 352 -161 430 -160
rect 499 -161 507 -160
rect 72 -163 122 -162
rect 149 -163 181 -162
rect 208 -163 416 -162
rect 79 -165 129 -164
rect 149 -165 157 -164
rect 219 -165 311 -164
rect 320 -165 437 -164
rect 79 -167 125 -166
rect 128 -167 185 -166
rect 226 -167 248 -166
rect 268 -167 437 -166
rect 86 -169 167 -168
rect 226 -169 332 -168
rect 345 -169 430 -168
rect 93 -171 146 -170
rect 236 -171 269 -170
rect 278 -171 461 -170
rect 100 -173 178 -172
rect 243 -173 339 -172
rect 352 -173 388 -172
rect 103 -175 143 -174
rect 177 -175 206 -174
rect 212 -175 339 -174
rect 359 -175 416 -174
rect 86 -177 143 -176
rect 212 -177 297 -176
rect 299 -177 423 -176
rect 107 -179 164 -178
rect 282 -179 318 -178
rect 324 -179 346 -178
rect 373 -179 465 -178
rect 107 -181 199 -180
rect 254 -181 325 -180
rect 373 -181 409 -180
rect 422 -181 444 -180
rect 114 -183 171 -182
rect 191 -183 255 -182
rect 299 -183 388 -182
rect 401 -183 409 -182
rect 93 -185 171 -184
rect 243 -185 444 -184
rect 121 -187 157 -186
rect 303 -187 360 -186
rect 394 -187 402 -186
rect 191 -189 304 -188
rect 380 -189 395 -188
rect 261 -191 381 -190
rect 240 -193 262 -192
rect 240 -195 276 -194
rect 275 -197 290 -196
rect 233 -199 290 -198
rect 79 -210 223 -209
rect 243 -210 325 -209
rect 348 -210 416 -209
rect 443 -210 454 -209
rect 506 -210 510 -209
rect 562 -210 573 -209
rect 86 -212 216 -211
rect 219 -212 339 -211
rect 380 -212 423 -211
rect 450 -212 461 -211
rect 100 -214 241 -213
rect 278 -214 437 -213
rect 107 -216 237 -215
rect 240 -216 255 -215
rect 296 -216 374 -215
rect 383 -216 395 -215
rect 114 -218 192 -217
rect 222 -218 465 -217
rect 114 -220 202 -219
rect 236 -220 283 -219
rect 317 -220 353 -219
rect 359 -220 374 -219
rect 128 -222 199 -221
rect 212 -222 318 -221
rect 320 -222 416 -221
rect 135 -224 146 -223
rect 156 -224 227 -223
rect 243 -224 437 -223
rect 128 -226 157 -225
rect 163 -226 276 -225
rect 282 -226 304 -225
rect 324 -226 346 -225
rect 135 -228 167 -227
rect 173 -228 265 -227
rect 289 -228 304 -227
rect 331 -228 444 -227
rect 142 -230 185 -229
rect 191 -230 248 -229
rect 254 -230 262 -229
rect 292 -230 332 -229
rect 338 -230 367 -229
rect 177 -232 216 -231
rect 226 -232 248 -231
rect 261 -232 395 -231
rect 184 -234 206 -233
rect 212 -234 293 -233
rect 296 -234 360 -233
rect 198 -236 311 -235
rect 345 -236 430 -235
rect 278 -238 311 -237
rect 352 -238 367 -237
rect 387 -238 430 -237
rect 275 -240 388 -239
rect 65 -251 94 -250
rect 107 -251 122 -250
rect 124 -251 160 -250
rect 177 -251 195 -250
rect 198 -251 262 -250
rect 292 -251 346 -250
rect 366 -251 402 -250
rect 415 -251 493 -250
rect 502 -251 521 -250
rect 590 -251 598 -250
rect 600 -251 612 -250
rect 79 -253 318 -252
rect 320 -253 339 -252
rect 422 -253 458 -252
rect 471 -253 500 -252
rect 506 -253 528 -252
rect 86 -255 129 -254
rect 135 -255 290 -254
rect 303 -255 402 -254
rect 429 -255 479 -254
rect 114 -257 328 -256
rect 338 -257 416 -256
rect 450 -257 486 -256
rect 114 -259 129 -258
rect 135 -259 171 -258
rect 173 -259 178 -258
rect 184 -259 230 -258
rect 254 -259 279 -258
rect 320 -259 409 -258
rect 464 -259 507 -258
rect 142 -261 237 -260
rect 257 -261 325 -260
rect 348 -261 423 -260
rect 436 -261 465 -260
rect 142 -263 185 -262
rect 187 -263 241 -262
rect 324 -263 360 -262
rect 373 -263 430 -262
rect 149 -265 157 -264
rect 163 -265 171 -264
rect 191 -265 244 -264
rect 303 -265 360 -264
rect 380 -265 409 -264
rect 149 -267 206 -266
rect 208 -267 234 -266
rect 236 -267 314 -266
rect 352 -267 374 -266
rect 387 -267 437 -266
rect 156 -269 220 -268
rect 222 -269 311 -268
rect 317 -269 353 -268
rect 394 -269 451 -268
rect 163 -271 244 -270
rect 331 -271 388 -270
rect 201 -273 276 -272
rect 299 -273 332 -272
rect 208 -275 367 -274
rect 219 -277 384 -276
rect 226 -279 283 -278
rect 275 -281 297 -280
rect 75 -292 255 -291
rect 257 -292 318 -291
rect 324 -292 479 -291
rect 516 -292 549 -291
rect 604 -292 612 -291
rect 646 -292 654 -291
rect 674 -292 682 -291
rect 79 -294 213 -293
rect 219 -294 297 -293
rect 303 -294 402 -293
rect 425 -294 458 -293
rect 464 -294 479 -293
rect 520 -294 542 -293
rect 649 -294 661 -293
rect 79 -296 108 -295
rect 114 -296 157 -295
rect 170 -296 178 -295
rect 187 -296 195 -295
rect 205 -296 283 -295
rect 289 -296 472 -295
rect 527 -296 545 -295
rect 86 -298 153 -297
rect 212 -298 234 -297
rect 236 -298 370 -297
rect 390 -298 493 -297
rect 506 -298 528 -297
rect 86 -300 143 -299
rect 219 -300 465 -299
rect 485 -300 507 -299
rect 93 -302 174 -301
rect 247 -302 321 -301
rect 324 -302 430 -301
rect 436 -302 535 -301
rect 93 -304 150 -303
rect 247 -304 346 -303
rect 348 -304 388 -303
rect 394 -304 430 -303
rect 100 -306 118 -305
rect 128 -306 143 -305
rect 254 -306 269 -305
rect 282 -306 486 -305
rect 103 -308 122 -307
rect 135 -308 199 -307
rect 261 -308 265 -307
rect 289 -308 339 -307
rect 341 -308 444 -307
rect 107 -310 164 -309
rect 198 -310 227 -309
rect 303 -310 423 -309
rect 443 -310 556 -309
rect 128 -312 136 -311
rect 163 -312 178 -311
rect 191 -312 227 -311
rect 313 -312 472 -311
rect 345 -314 451 -313
rect 352 -316 402 -315
rect 408 -316 451 -315
rect 331 -318 353 -317
rect 366 -318 381 -317
rect 408 -318 458 -317
rect 331 -320 388 -319
rect 415 -320 493 -319
rect 240 -322 416 -321
rect 422 -322 500 -321
rect 229 -324 241 -323
rect 366 -324 437 -323
rect 373 -326 395 -325
rect 359 -328 374 -327
rect 359 -330 521 -329
rect 44 -341 335 -340
rect 338 -341 528 -340
rect 541 -341 570 -340
rect 583 -341 605 -340
rect 642 -341 689 -340
rect 51 -343 115 -342
rect 128 -343 143 -342
rect 166 -343 237 -342
rect 243 -343 262 -342
rect 264 -343 626 -342
rect 649 -343 654 -342
rect 660 -343 682 -342
rect 58 -345 290 -344
rect 296 -345 314 -344
rect 341 -345 430 -344
rect 471 -345 514 -344
rect 523 -345 598 -344
rect 667 -345 675 -344
rect 79 -347 220 -346
rect 233 -347 346 -346
rect 359 -347 612 -346
rect 79 -349 171 -348
rect 177 -349 227 -348
rect 233 -349 353 -348
rect 362 -349 535 -348
rect 544 -349 640 -348
rect 86 -351 164 -350
rect 177 -351 216 -350
rect 222 -351 363 -350
rect 366 -351 619 -350
rect 86 -353 248 -352
rect 254 -353 269 -352
rect 275 -353 297 -352
rect 341 -353 528 -352
rect 548 -353 647 -352
rect 93 -355 157 -354
rect 159 -355 255 -354
rect 292 -355 367 -354
rect 380 -355 391 -354
rect 411 -355 437 -354
rect 460 -355 535 -354
rect 558 -355 563 -354
rect 72 -357 157 -356
rect 205 -357 286 -356
rect 327 -357 549 -356
rect 562 -357 654 -356
rect 72 -359 213 -358
rect 236 -359 272 -358
rect 327 -359 409 -358
rect 415 -359 437 -358
rect 471 -359 661 -358
rect 93 -361 101 -360
rect 114 -361 402 -360
rect 415 -361 426 -360
rect 478 -361 542 -360
rect 100 -363 122 -362
rect 128 -363 136 -362
rect 142 -363 230 -362
rect 373 -363 479 -362
rect 485 -363 591 -362
rect 68 -365 136 -364
rect 152 -365 220 -364
rect 380 -365 388 -364
rect 394 -365 402 -364
rect 422 -365 577 -364
rect 107 -367 153 -366
rect 205 -367 241 -366
rect 317 -367 395 -366
rect 422 -367 521 -366
rect 107 -369 248 -368
rect 317 -369 458 -368
rect 492 -369 605 -368
rect 110 -371 374 -370
rect 443 -371 486 -370
rect 499 -371 556 -370
rect 121 -373 192 -372
rect 303 -373 444 -372
rect 450 -373 493 -372
rect 506 -373 633 -372
rect 170 -375 241 -374
rect 303 -375 325 -374
rect 348 -375 500 -374
rect 184 -377 192 -376
rect 310 -377 325 -376
rect 429 -377 451 -376
rect 464 -377 507 -376
rect 184 -379 199 -378
rect 331 -379 465 -378
rect 138 -381 199 -380
rect 282 -381 332 -380
rect 2 -392 181 -391
rect 205 -392 227 -391
rect 233 -392 311 -391
rect 317 -392 353 -391
rect 359 -392 612 -391
rect 628 -392 640 -391
rect 649 -392 682 -391
rect 16 -394 293 -393
rect 303 -394 353 -393
rect 355 -394 360 -393
rect 373 -394 563 -393
rect 597 -394 612 -393
rect 667 -394 675 -393
rect 30 -396 38 -395
rect 44 -396 223 -395
rect 240 -396 465 -395
rect 597 -396 626 -395
rect 667 -396 689 -395
rect 44 -398 398 -397
rect 401 -398 423 -397
rect 436 -398 447 -397
rect 450 -398 647 -397
rect 51 -400 139 -399
rect 149 -400 192 -399
rect 215 -400 395 -399
rect 401 -400 633 -399
rect 51 -402 153 -401
rect 163 -402 185 -401
rect 219 -402 405 -401
rect 436 -402 535 -401
rect 576 -402 633 -401
rect 58 -404 342 -403
rect 373 -404 451 -403
rect 460 -404 549 -403
rect 558 -404 577 -403
rect 583 -404 626 -403
rect 58 -406 213 -405
rect 268 -406 290 -405
rect 317 -406 367 -405
rect 376 -406 416 -405
rect 439 -406 605 -405
rect 65 -408 304 -407
rect 334 -408 591 -407
rect 604 -408 654 -407
rect 72 -410 328 -409
rect 341 -410 479 -409
rect 492 -410 535 -409
rect 569 -410 584 -409
rect 653 -410 664 -409
rect 72 -412 188 -411
rect 254 -412 269 -411
rect 285 -412 297 -411
rect 369 -412 479 -411
rect 541 -412 570 -411
rect 79 -414 241 -413
rect 247 -414 297 -413
rect 387 -414 619 -413
rect 79 -416 216 -415
rect 247 -416 262 -415
rect 289 -416 332 -415
rect 387 -416 444 -415
rect 467 -416 591 -415
rect 86 -418 325 -417
rect 345 -418 444 -417
rect 471 -418 493 -417
rect 499 -418 542 -417
rect 555 -418 619 -417
rect 100 -420 160 -419
rect 184 -420 192 -419
rect 236 -420 346 -419
rect 408 -420 500 -419
rect 100 -422 146 -421
rect 159 -422 521 -421
rect 107 -424 199 -423
rect 236 -424 279 -423
rect 324 -424 507 -423
rect 114 -426 276 -425
rect 408 -426 458 -425
rect 114 -428 129 -427
rect 135 -428 167 -427
rect 198 -428 549 -427
rect 121 -430 311 -429
rect 415 -430 430 -429
rect 446 -430 472 -429
rect 86 -432 122 -431
rect 128 -432 171 -431
rect 261 -432 283 -431
rect 338 -432 430 -431
rect 142 -434 255 -433
rect 170 -436 178 -435
rect 205 -436 283 -435
rect 23 -438 178 -437
rect 9 -449 111 -448
rect 131 -449 521 -448
rect 541 -449 556 -448
rect 558 -449 584 -448
rect 611 -449 615 -448
rect 635 -449 654 -448
rect 660 -449 668 -448
rect 9 -451 356 -450
rect 369 -451 535 -450
rect 583 -451 605 -450
rect 653 -451 664 -450
rect 16 -453 237 -452
rect 247 -453 286 -452
rect 292 -453 416 -452
rect 418 -453 535 -452
rect 16 -455 115 -454
rect 142 -455 171 -454
rect 208 -455 332 -454
rect 373 -455 500 -454
rect 520 -455 563 -454
rect 23 -457 181 -456
rect 215 -457 262 -456
rect 275 -457 339 -456
rect 376 -457 514 -456
rect 23 -459 87 -458
rect 107 -459 171 -458
rect 177 -459 374 -458
rect 397 -459 493 -458
rect 499 -459 510 -458
rect 513 -459 528 -458
rect 30 -461 139 -460
rect 142 -461 297 -460
rect 324 -461 416 -460
rect 436 -461 542 -460
rect 33 -463 38 -462
rect 44 -463 157 -462
rect 159 -463 360 -462
rect 408 -463 423 -462
rect 436 -463 619 -462
rect 37 -465 108 -464
rect 121 -465 139 -464
rect 163 -465 188 -464
rect 233 -465 304 -464
rect 359 -465 388 -464
rect 457 -465 510 -464
rect 576 -465 619 -464
rect 44 -467 150 -466
rect 163 -467 346 -466
rect 387 -467 472 -466
rect 478 -467 563 -466
rect 576 -467 598 -466
rect 51 -469 185 -468
rect 219 -469 234 -468
rect 243 -469 493 -468
rect 597 -469 626 -468
rect 2 -471 244 -470
rect 247 -471 465 -470
rect 485 -471 528 -470
rect 51 -473 101 -472
rect 121 -473 265 -472
rect 275 -473 353 -472
rect 397 -473 486 -472
rect 58 -475 146 -474
rect 166 -475 185 -474
rect 205 -475 220 -474
rect 254 -475 290 -474
rect 296 -475 633 -474
rect 58 -477 402 -476
rect 429 -477 458 -476
rect 632 -477 640 -476
rect 65 -479 367 -478
rect 429 -479 444 -478
rect 450 -479 472 -478
rect 590 -479 640 -478
rect 65 -481 549 -480
rect 72 -483 202 -482
rect 212 -483 255 -482
rect 268 -483 290 -482
rect 345 -483 405 -482
rect 548 -483 570 -482
rect 72 -485 129 -484
rect 177 -485 192 -484
rect 215 -485 367 -484
rect 390 -485 444 -484
rect 79 -487 423 -486
rect 79 -489 94 -488
rect 100 -489 199 -488
rect 282 -489 465 -488
rect 86 -491 115 -490
rect 128 -491 192 -490
rect 282 -491 311 -490
rect 352 -491 451 -490
rect 310 -493 381 -492
rect 380 -495 570 -494
rect 5 -506 164 -505
rect 198 -506 363 -505
rect 366 -506 612 -505
rect 618 -506 629 -505
rect 653 -506 671 -505
rect 681 -506 689 -505
rect 9 -508 118 -507
rect 121 -508 125 -507
rect 152 -508 276 -507
rect 285 -508 570 -507
rect 583 -508 612 -507
rect 628 -508 647 -507
rect 667 -508 675 -507
rect 9 -510 62 -509
rect 65 -510 87 -509
rect 93 -510 101 -509
rect 121 -510 248 -509
rect 268 -510 297 -509
rect 310 -510 377 -509
rect 383 -510 493 -509
rect 499 -510 591 -509
rect 604 -510 615 -509
rect 618 -510 647 -509
rect 23 -512 59 -511
rect 68 -512 213 -511
rect 219 -512 276 -511
rect 289 -512 311 -511
rect 338 -512 349 -511
rect 369 -512 605 -511
rect 639 -512 654 -511
rect 23 -514 241 -513
rect 243 -514 563 -513
rect 576 -514 591 -513
rect 30 -516 209 -515
rect 212 -516 227 -515
rect 243 -516 388 -515
rect 390 -516 542 -515
rect 555 -516 563 -515
rect 30 -518 181 -517
rect 278 -518 556 -517
rect 37 -520 157 -519
rect 163 -520 437 -519
rect 450 -520 493 -519
rect 502 -520 514 -519
rect 37 -522 143 -521
rect 149 -522 220 -521
rect 292 -522 437 -521
rect 478 -522 570 -521
rect 16 -524 150 -523
rect 156 -524 234 -523
rect 296 -524 304 -523
rect 331 -524 542 -523
rect 16 -526 83 -525
rect 86 -526 101 -525
rect 114 -526 577 -525
rect 44 -528 216 -527
rect 303 -528 325 -527
rect 341 -528 451 -527
rect 457 -528 479 -527
rect 485 -528 584 -527
rect 44 -530 241 -529
rect 324 -530 346 -529
rect 373 -530 395 -529
rect 397 -530 598 -529
rect 72 -532 136 -531
rect 170 -532 227 -531
rect 345 -532 381 -531
rect 415 -532 528 -531
rect 548 -532 598 -531
rect 51 -534 73 -533
rect 93 -534 192 -533
rect 205 -534 234 -533
rect 359 -534 395 -533
rect 415 -534 430 -533
rect 471 -534 486 -533
rect 499 -534 528 -533
rect 534 -534 549 -533
rect 51 -536 80 -535
rect 107 -536 136 -535
rect 170 -536 283 -535
rect 401 -536 472 -535
rect 506 -536 521 -535
rect 107 -538 185 -537
rect 208 -538 430 -537
rect 464 -538 535 -537
rect 124 -540 248 -539
rect 261 -540 402 -539
rect 422 -540 640 -539
rect 128 -542 332 -541
rect 355 -542 465 -541
rect 513 -542 626 -541
rect 131 -544 206 -543
rect 313 -544 521 -543
rect 159 -546 185 -545
rect 355 -546 409 -545
rect 177 -548 199 -547
rect 408 -548 444 -547
rect 317 -550 444 -549
rect 271 -552 318 -551
rect 2 -563 269 -562
rect 275 -563 321 -562
rect 345 -563 423 -562
rect 436 -563 619 -562
rect 646 -563 668 -562
rect 670 -563 685 -562
rect 19 -565 307 -564
rect 310 -565 395 -564
rect 401 -565 633 -564
rect 653 -565 657 -564
rect 674 -565 678 -564
rect 23 -567 97 -566
rect 107 -567 293 -566
rect 296 -567 370 -566
rect 380 -567 402 -566
rect 404 -567 598 -566
rect 618 -567 626 -566
rect 653 -567 661 -566
rect 23 -569 122 -568
rect 128 -569 220 -568
rect 233 -569 269 -568
rect 278 -569 542 -568
rect 590 -569 647 -568
rect 9 -571 129 -570
rect 131 -571 605 -570
rect 9 -573 178 -572
rect 180 -573 472 -572
rect 478 -573 591 -572
rect 604 -573 626 -572
rect 30 -575 101 -574
rect 107 -575 171 -574
rect 243 -575 640 -574
rect 30 -577 234 -576
rect 247 -577 381 -576
rect 383 -577 479 -576
rect 499 -577 514 -576
rect 534 -577 542 -576
rect 562 -577 640 -576
rect 37 -579 342 -578
rect 345 -579 353 -578
rect 355 -579 444 -578
rect 457 -579 493 -578
rect 40 -581 181 -580
rect 184 -581 248 -580
rect 254 -581 475 -580
rect 485 -581 514 -580
rect 44 -583 143 -582
rect 163 -583 220 -582
rect 285 -583 339 -582
rect 366 -583 377 -582
rect 387 -583 598 -582
rect 51 -585 55 -584
rect 65 -585 83 -584
rect 93 -585 297 -584
rect 317 -585 570 -584
rect 16 -587 94 -586
rect 100 -587 118 -586
rect 121 -587 178 -586
rect 212 -587 255 -586
rect 289 -587 535 -586
rect 548 -587 570 -586
rect 51 -589 87 -588
rect 114 -589 157 -588
rect 163 -589 227 -588
rect 236 -589 318 -588
rect 366 -589 633 -588
rect 58 -591 115 -590
rect 131 -591 283 -590
rect 289 -591 468 -590
rect 471 -591 612 -590
rect 656 -591 661 -590
rect 65 -593 104 -592
rect 135 -593 195 -592
rect 198 -593 227 -592
rect 282 -593 304 -592
rect 373 -593 444 -592
rect 485 -593 521 -592
rect 583 -593 612 -592
rect 75 -595 311 -594
rect 359 -595 584 -594
rect 79 -597 185 -596
rect 198 -597 244 -596
rect 303 -597 556 -596
rect 135 -599 262 -598
rect 359 -599 426 -598
rect 429 -599 458 -598
rect 460 -599 521 -598
rect 527 -599 556 -598
rect 142 -601 188 -600
rect 205 -601 430 -600
rect 450 -601 528 -600
rect 170 -603 192 -602
rect 205 -603 314 -602
rect 373 -603 398 -602
rect 450 -603 465 -602
rect 506 -603 549 -602
rect 212 -605 265 -604
rect 331 -605 507 -604
rect 324 -607 332 -606
rect 387 -607 437 -606
rect 464 -607 563 -606
rect 72 -609 325 -608
rect 2 -620 395 -619
rect 411 -620 591 -619
rect 632 -620 703 -619
rect 716 -620 731 -619
rect 2 -622 45 -621
rect 51 -622 115 -621
rect 159 -622 248 -621
rect 285 -622 472 -621
rect 492 -622 640 -621
rect 653 -622 661 -621
rect 681 -622 689 -621
rect 695 -622 720 -621
rect 9 -624 188 -623
rect 194 -624 290 -623
rect 296 -624 349 -623
rect 355 -624 360 -623
rect 376 -624 521 -623
rect 527 -624 605 -623
rect 618 -624 661 -623
rect 9 -626 87 -625
rect 93 -626 101 -625
rect 107 -626 353 -625
rect 380 -626 654 -625
rect 23 -628 97 -627
rect 107 -628 150 -627
rect 166 -628 171 -627
rect 177 -628 388 -627
rect 390 -628 577 -627
rect 583 -628 619 -627
rect 23 -630 174 -629
rect 177 -630 213 -629
rect 226 -630 262 -629
rect 289 -630 374 -629
rect 383 -630 570 -629
rect 30 -632 370 -631
rect 394 -632 409 -631
rect 425 -632 549 -631
rect 562 -632 591 -631
rect 30 -634 164 -633
rect 184 -634 279 -633
rect 345 -634 381 -633
rect 453 -634 668 -633
rect 16 -636 279 -635
rect 345 -636 493 -635
rect 495 -636 549 -635
rect 37 -638 62 -637
rect 72 -638 122 -637
rect 128 -638 164 -637
rect 212 -638 220 -637
rect 240 -638 255 -637
rect 366 -638 570 -637
rect 44 -640 90 -639
rect 93 -640 521 -639
rect 541 -640 563 -639
rect 54 -642 255 -641
rect 303 -642 367 -641
rect 369 -642 556 -641
rect 58 -644 76 -643
rect 114 -644 157 -643
rect 240 -644 269 -643
rect 324 -644 556 -643
rect 117 -646 167 -645
rect 229 -646 269 -645
rect 324 -646 402 -645
rect 453 -646 633 -645
rect 121 -648 146 -647
rect 149 -648 206 -647
rect 243 -648 283 -647
rect 310 -648 402 -647
rect 464 -648 612 -647
rect 79 -650 311 -649
rect 387 -650 465 -649
rect 474 -650 640 -649
rect 79 -652 129 -651
rect 135 -652 220 -651
rect 282 -652 584 -651
rect 142 -654 248 -653
rect 506 -654 528 -653
rect 534 -654 612 -653
rect 142 -656 486 -655
rect 499 -656 535 -655
rect 156 -658 234 -657
rect 243 -658 507 -657
rect 513 -658 542 -657
rect 198 -660 206 -659
rect 338 -660 486 -659
rect 135 -662 199 -661
rect 457 -662 500 -661
rect 191 -664 339 -663
rect 457 -664 647 -663
rect 191 -666 678 -665
rect 478 -668 514 -667
rect 625 -668 647 -667
rect 443 -670 479 -669
rect 597 -670 626 -669
rect 299 -672 598 -671
rect 429 -674 444 -673
rect 415 -676 430 -675
rect 415 -678 437 -677
rect 422 -680 437 -679
rect 422 -682 577 -681
rect 2 -693 80 -692
rect 82 -693 437 -692
rect 450 -693 542 -692
rect 632 -693 724 -692
rect 730 -693 755 -692
rect 800 -693 808 -692
rect 9 -695 139 -694
rect 215 -695 311 -694
rect 341 -695 472 -694
rect 534 -695 717 -694
rect 16 -697 325 -696
rect 345 -697 528 -696
rect 674 -697 696 -696
rect 702 -697 745 -696
rect 19 -699 104 -698
rect 121 -699 164 -698
rect 226 -699 262 -698
rect 278 -699 584 -698
rect 653 -699 696 -698
rect 9 -701 227 -700
rect 236 -701 461 -700
rect 464 -701 612 -700
rect 646 -701 654 -700
rect 23 -703 188 -702
rect 254 -703 412 -702
rect 422 -703 689 -702
rect 23 -705 167 -704
rect 201 -705 423 -704
rect 429 -705 465 -704
rect 499 -705 535 -704
rect 569 -705 689 -704
rect 30 -707 241 -706
rect 254 -707 290 -706
rect 296 -707 402 -706
rect 408 -707 633 -706
rect 30 -709 94 -708
rect 100 -709 388 -708
rect 401 -709 458 -708
rect 467 -709 570 -708
rect 576 -709 612 -708
rect 37 -711 90 -710
rect 93 -711 157 -710
rect 240 -711 430 -710
rect 432 -711 626 -710
rect 2 -713 90 -712
rect 100 -713 738 -712
rect 40 -715 304 -714
rect 310 -715 332 -714
rect 352 -715 363 -714
rect 366 -715 619 -714
rect 44 -717 192 -716
rect 233 -717 353 -716
rect 359 -717 675 -716
rect 44 -719 125 -718
rect 135 -719 213 -718
rect 247 -719 363 -718
rect 373 -719 384 -718
rect 408 -719 605 -718
rect 58 -721 66 -720
rect 142 -721 304 -720
rect 317 -721 346 -720
rect 373 -721 454 -720
rect 548 -721 577 -720
rect 583 -721 682 -720
rect 65 -723 395 -722
rect 415 -723 500 -722
rect 562 -723 626 -722
rect 142 -725 283 -724
rect 296 -725 370 -724
rect 436 -725 521 -724
rect 565 -725 605 -724
rect 149 -727 213 -726
rect 247 -727 668 -726
rect 114 -729 150 -728
rect 156 -729 388 -728
rect 443 -729 458 -728
rect 492 -729 549 -728
rect 590 -729 647 -728
rect 114 -731 206 -730
rect 261 -731 734 -730
rect 184 -733 206 -732
rect 278 -733 325 -732
rect 331 -733 381 -732
rect 450 -733 472 -732
rect 492 -733 591 -732
rect 597 -733 619 -732
rect 639 -733 668 -732
rect 170 -735 185 -734
rect 191 -735 269 -734
rect 299 -735 339 -734
rect 348 -735 416 -734
rect 453 -735 661 -734
rect 107 -737 269 -736
rect 317 -737 328 -736
rect 366 -737 563 -736
rect 107 -739 178 -738
rect 243 -739 640 -738
rect 170 -741 199 -740
rect 376 -741 444 -740
rect 506 -741 521 -740
rect 555 -741 598 -740
rect 51 -743 199 -742
rect 380 -743 703 -742
rect 177 -745 293 -744
rect 383 -745 661 -744
rect 485 -747 507 -746
rect 513 -747 556 -746
rect 485 -749 514 -748
rect 30 -760 409 -759
rect 429 -760 752 -759
rect 30 -762 83 -761
rect 89 -762 150 -761
rect 177 -762 230 -761
rect 243 -762 276 -761
rect 289 -762 311 -761
rect 327 -762 640 -761
rect 674 -762 731 -761
rect 733 -762 745 -761
rect 2 -764 90 -763
rect 107 -764 202 -763
rect 226 -764 346 -763
rect 387 -764 717 -763
rect 723 -764 738 -763
rect 23 -766 388 -765
rect 390 -766 591 -765
rect 604 -766 766 -765
rect 23 -768 55 -767
rect 58 -768 87 -767
rect 100 -768 108 -767
rect 121 -768 139 -767
rect 142 -768 286 -767
rect 299 -768 409 -767
rect 422 -768 738 -767
rect 37 -770 94 -769
rect 100 -770 255 -769
rect 261 -770 325 -769
rect 334 -770 514 -769
rect 527 -770 626 -769
rect 632 -770 745 -769
rect 51 -772 675 -771
rect 702 -772 759 -771
rect 58 -774 192 -773
rect 247 -774 255 -773
rect 341 -774 444 -773
rect 495 -774 647 -773
rect 712 -774 787 -773
rect 65 -776 384 -775
rect 390 -776 423 -775
rect 436 -776 724 -775
rect 65 -778 87 -777
rect 93 -778 251 -777
rect 345 -778 353 -777
rect 373 -778 514 -777
rect 541 -778 654 -777
rect 72 -780 80 -779
rect 121 -780 717 -779
rect 72 -782 192 -781
rect 247 -782 318 -781
rect 352 -782 419 -781
rect 439 -782 640 -781
rect 79 -784 265 -783
rect 303 -784 654 -783
rect 124 -786 164 -785
rect 170 -786 311 -785
rect 373 -786 381 -785
rect 383 -786 773 -785
rect 2 -788 164 -787
rect 170 -788 293 -787
rect 303 -788 332 -787
rect 380 -788 605 -787
rect 611 -788 626 -787
rect 632 -788 668 -787
rect 9 -790 125 -789
rect 149 -790 241 -789
rect 394 -790 461 -789
rect 464 -790 542 -789
rect 544 -790 710 -789
rect 9 -792 129 -791
rect 156 -792 227 -791
rect 240 -792 794 -791
rect 16 -794 332 -793
rect 362 -794 465 -793
rect 488 -794 647 -793
rect 16 -796 136 -795
rect 156 -796 216 -795
rect 397 -796 451 -795
rect 453 -796 668 -795
rect 44 -798 136 -797
rect 177 -798 199 -797
rect 212 -798 318 -797
rect 366 -798 451 -797
rect 548 -798 584 -797
rect 586 -798 689 -797
rect 44 -800 339 -799
rect 404 -800 584 -799
rect 590 -800 598 -799
rect 618 -800 703 -799
rect 128 -802 220 -801
rect 222 -802 339 -801
rect 411 -802 444 -801
rect 534 -802 619 -801
rect 681 -802 689 -801
rect 103 -804 535 -803
rect 555 -804 682 -803
rect 184 -806 213 -805
rect 219 -806 269 -805
rect 415 -806 496 -805
rect 520 -806 556 -805
rect 562 -806 696 -805
rect 114 -808 185 -807
rect 198 -808 661 -807
rect 695 -808 755 -807
rect 110 -810 115 -809
rect 233 -810 367 -809
rect 436 -810 598 -809
rect 205 -812 234 -811
rect 268 -812 402 -811
rect 499 -812 563 -811
rect 569 -812 780 -811
rect 205 -814 237 -813
rect 359 -814 570 -813
rect 576 -814 612 -813
rect 296 -816 360 -815
rect 499 -816 507 -815
rect 520 -816 804 -815
rect 296 -818 549 -817
rect 471 -820 507 -819
rect 523 -820 577 -819
rect 457 -822 472 -821
rect 530 -822 661 -821
rect 457 -824 479 -823
rect 478 -826 493 -825
rect 9 -837 241 -836
rect 278 -837 794 -836
rect 803 -837 808 -836
rect 9 -839 150 -838
rect 159 -839 458 -838
rect 460 -839 766 -838
rect 16 -841 174 -840
rect 184 -841 297 -840
rect 366 -841 437 -840
rect 439 -841 780 -840
rect 16 -843 181 -842
rect 184 -843 353 -842
rect 359 -843 437 -842
rect 460 -843 738 -842
rect 751 -843 776 -842
rect 23 -845 146 -844
rect 149 -845 402 -844
rect 404 -845 563 -844
rect 730 -845 738 -844
rect 751 -845 783 -844
rect 30 -847 237 -846
rect 240 -847 248 -846
rect 268 -847 353 -846
rect 366 -847 388 -846
rect 390 -847 787 -846
rect 37 -849 87 -848
rect 107 -849 157 -848
rect 166 -849 213 -848
rect 215 -849 675 -848
rect 716 -849 731 -848
rect 786 -849 797 -848
rect 44 -851 139 -850
rect 156 -851 535 -850
rect 667 -851 675 -850
rect 54 -853 773 -852
rect 58 -855 300 -854
rect 338 -855 668 -854
rect 72 -857 248 -856
rect 268 -857 318 -856
rect 373 -857 535 -856
rect 646 -857 773 -856
rect 51 -859 73 -858
rect 82 -859 640 -858
rect 128 -861 213 -860
rect 219 -861 244 -860
rect 275 -861 339 -860
rect 383 -861 766 -860
rect 2 -863 276 -862
rect 282 -863 318 -862
rect 397 -863 605 -862
rect 44 -865 129 -864
rect 135 -865 430 -864
rect 467 -865 682 -864
rect 170 -867 188 -866
rect 201 -867 360 -866
rect 401 -867 416 -866
rect 418 -867 619 -866
rect 93 -869 202 -868
rect 226 -869 290 -868
rect 292 -869 717 -868
rect 58 -871 227 -870
rect 229 -871 661 -870
rect 93 -873 115 -872
rect 170 -873 255 -872
rect 282 -873 374 -872
rect 411 -873 661 -872
rect 114 -875 122 -874
rect 177 -875 220 -874
rect 233 -875 262 -874
rect 296 -875 311 -874
rect 334 -875 430 -874
rect 488 -875 710 -874
rect 37 -877 234 -876
rect 303 -877 311 -876
rect 348 -877 710 -876
rect 65 -879 122 -878
rect 177 -879 654 -878
rect 65 -881 164 -880
rect 187 -881 255 -880
rect 303 -881 395 -880
rect 422 -881 493 -880
rect 506 -881 521 -880
rect 523 -881 745 -880
rect 324 -883 423 -882
rect 488 -883 724 -882
rect 191 -885 325 -884
rect 394 -885 542 -884
rect 569 -885 647 -884
rect 653 -885 696 -884
rect 450 -887 542 -886
rect 576 -887 605 -886
rect 611 -887 682 -886
rect 695 -887 703 -886
rect 450 -889 759 -888
rect 464 -891 612 -890
rect 618 -891 633 -890
rect 152 -893 633 -892
rect 464 -895 570 -894
rect 583 -895 759 -894
rect 495 -897 703 -896
rect 499 -899 507 -898
rect 513 -899 563 -898
rect 583 -899 591 -898
rect 478 -901 514 -900
rect 527 -901 745 -900
rect 100 -903 479 -902
rect 499 -903 640 -902
rect 79 -905 101 -904
rect 443 -905 528 -904
rect 530 -905 549 -904
rect 590 -905 598 -904
rect 79 -907 346 -906
rect 485 -907 549 -906
rect 555 -907 598 -906
rect 331 -909 444 -908
rect 471 -909 556 -908
rect 331 -911 381 -910
rect 408 -911 472 -910
rect 408 -913 724 -912
rect 9 -924 223 -923
rect 229 -924 339 -923
rect 348 -924 612 -923
rect 723 -924 755 -923
rect 779 -924 787 -923
rect 9 -926 353 -925
rect 366 -926 444 -925
rect 446 -926 731 -925
rect 751 -926 776 -925
rect 16 -928 118 -927
rect 121 -928 129 -927
rect 142 -928 153 -927
rect 159 -928 426 -927
rect 432 -928 514 -927
rect 576 -928 731 -927
rect 16 -930 101 -929
rect 107 -930 143 -929
rect 149 -930 374 -929
rect 408 -930 535 -929
rect 576 -930 647 -929
rect 723 -930 741 -929
rect 23 -932 234 -931
rect 236 -932 654 -931
rect 23 -934 104 -933
rect 107 -934 276 -933
rect 285 -934 423 -933
rect 460 -934 738 -933
rect 30 -936 412 -935
rect 415 -936 486 -935
rect 499 -936 696 -935
rect 30 -938 185 -937
rect 191 -938 199 -937
rect 201 -938 503 -937
rect 513 -938 556 -937
rect 579 -938 605 -937
rect 681 -938 738 -937
rect 37 -940 83 -939
rect 86 -940 258 -939
rect 275 -940 304 -939
rect 310 -940 314 -939
rect 317 -940 381 -939
rect 418 -940 598 -939
rect 604 -940 626 -939
rect 674 -940 682 -939
rect 37 -942 76 -941
rect 86 -942 97 -941
rect 114 -942 122 -941
rect 135 -942 234 -941
rect 243 -942 262 -941
rect 296 -942 304 -941
rect 348 -942 402 -941
rect 418 -942 500 -941
rect 527 -942 626 -941
rect 44 -944 398 -943
rect 464 -944 766 -943
rect 51 -946 101 -945
rect 114 -946 654 -945
rect 51 -948 94 -947
rect 149 -948 286 -947
rect 359 -948 402 -947
rect 467 -948 745 -947
rect 65 -950 290 -949
rect 397 -950 437 -949
rect 471 -950 612 -949
rect 618 -950 675 -949
rect 79 -952 136 -951
rect 163 -952 409 -951
rect 488 -952 696 -951
rect 44 -954 80 -953
rect 89 -954 563 -953
rect 590 -954 647 -953
rect 163 -956 213 -955
rect 226 -956 339 -955
rect 429 -956 591 -955
rect 597 -956 661 -955
rect 58 -958 430 -957
rect 506 -958 563 -957
rect 618 -958 773 -957
rect 58 -960 475 -959
rect 478 -960 507 -959
rect 520 -960 528 -959
rect 534 -960 759 -959
rect 170 -962 444 -961
rect 457 -962 479 -961
rect 555 -962 570 -961
rect 632 -962 661 -961
rect 177 -964 377 -963
rect 390 -964 570 -963
rect 583 -964 633 -963
rect 180 -966 381 -965
rect 457 -966 493 -965
rect 583 -966 640 -965
rect 184 -968 269 -967
rect 278 -968 759 -967
rect 191 -970 206 -969
rect 212 -970 220 -969
rect 226 -970 318 -969
rect 471 -970 521 -969
rect 639 -970 668 -969
rect 205 -972 241 -971
rect 243 -972 332 -971
rect 492 -972 542 -971
rect 667 -972 703 -971
rect 198 -974 332 -973
rect 702 -974 710 -973
rect 219 -976 262 -975
rect 268 -976 325 -975
rect 709 -976 717 -975
rect 247 -978 346 -977
rect 394 -978 717 -977
rect 236 -980 248 -979
rect 254 -980 363 -979
rect 254 -982 542 -981
rect 289 -984 451 -983
rect 296 -986 451 -985
rect 310 -988 437 -987
rect 324 -990 388 -989
rect 9 -1001 318 -1000
rect 334 -1001 409 -1000
rect 411 -1001 514 -1000
rect 737 -1001 745 -1000
rect 16 -1003 195 -1002
rect 198 -1003 370 -1002
rect 373 -1003 384 -1002
rect 394 -1003 405 -1002
rect 408 -1003 465 -1002
rect 471 -1003 675 -1002
rect 740 -1003 759 -1002
rect 23 -1005 241 -1004
rect 243 -1005 360 -1004
rect 362 -1005 577 -1004
rect 23 -1007 150 -1006
rect 166 -1007 223 -1006
rect 233 -1007 332 -1006
rect 338 -1007 367 -1006
rect 373 -1007 556 -1006
rect 576 -1007 692 -1006
rect 30 -1009 244 -1008
rect 250 -1009 262 -1008
rect 268 -1009 318 -1008
rect 338 -1009 500 -1008
rect 33 -1011 181 -1010
rect 191 -1011 220 -1010
rect 247 -1011 262 -1010
rect 282 -1011 640 -1010
rect 37 -1013 80 -1012
rect 107 -1013 311 -1012
rect 345 -1013 731 -1012
rect 37 -1015 108 -1014
rect 114 -1015 755 -1014
rect 44 -1017 62 -1016
rect 65 -1017 94 -1016
rect 114 -1017 122 -1016
rect 142 -1017 153 -1016
rect 170 -1017 220 -1016
rect 296 -1017 346 -1016
rect 348 -1017 440 -1016
rect 443 -1017 549 -1016
rect 562 -1017 731 -1016
rect 51 -1019 118 -1018
rect 121 -1019 185 -1018
rect 205 -1019 255 -1018
rect 275 -1019 297 -1018
rect 352 -1019 619 -1018
rect 51 -1021 104 -1020
rect 135 -1021 143 -1020
rect 149 -1021 234 -1020
rect 352 -1021 356 -1020
rect 376 -1021 507 -1020
rect 590 -1021 619 -1020
rect 58 -1023 185 -1022
rect 191 -1023 206 -1022
rect 212 -1023 283 -1022
rect 380 -1023 388 -1022
rect 415 -1023 661 -1022
rect 65 -1025 97 -1024
rect 135 -1025 160 -1024
rect 163 -1025 255 -1024
rect 380 -1025 584 -1024
rect 590 -1025 598 -1024
rect 72 -1027 87 -1026
rect 170 -1027 227 -1026
rect 383 -1027 556 -1026
rect 597 -1027 654 -1026
rect 44 -1029 87 -1028
rect 156 -1029 227 -1028
rect 310 -1029 654 -1028
rect 75 -1031 164 -1030
rect 397 -1031 584 -1030
rect 79 -1033 129 -1032
rect 156 -1033 178 -1032
rect 418 -1033 458 -1032
rect 478 -1033 549 -1032
rect 128 -1035 290 -1034
rect 401 -1035 458 -1034
rect 478 -1035 710 -1034
rect 177 -1037 269 -1036
rect 289 -1037 325 -1036
rect 401 -1037 626 -1036
rect 646 -1037 710 -1036
rect 324 -1039 521 -1038
rect 625 -1039 696 -1038
rect 313 -1041 696 -1040
rect 212 -1043 314 -1042
rect 425 -1043 661 -1042
rect 432 -1045 675 -1044
rect 436 -1047 444 -1046
rect 446 -1047 493 -1046
rect 495 -1047 514 -1046
rect 520 -1047 535 -1046
rect 646 -1047 703 -1046
rect 450 -1049 612 -1048
rect 702 -1049 724 -1048
rect 453 -1051 668 -1050
rect 467 -1053 612 -1052
rect 667 -1053 717 -1052
rect 485 -1055 640 -1054
rect 716 -1055 738 -1054
rect 278 -1057 486 -1056
rect 492 -1057 570 -1056
rect 499 -1059 528 -1058
rect 541 -1059 724 -1058
rect 425 -1061 528 -1060
rect 569 -1061 633 -1060
rect 429 -1063 542 -1062
rect 632 -1063 682 -1062
rect 681 -1065 720 -1064
rect 9 -1076 122 -1075
rect 128 -1076 216 -1075
rect 243 -1076 363 -1075
rect 387 -1076 416 -1075
rect 418 -1076 661 -1075
rect 677 -1076 689 -1075
rect 16 -1078 31 -1077
rect 37 -1078 181 -1077
rect 187 -1078 262 -1077
rect 278 -1078 304 -1077
rect 313 -1078 409 -1077
rect 415 -1078 458 -1077
rect 478 -1078 692 -1077
rect 44 -1080 125 -1079
rect 128 -1080 213 -1079
rect 254 -1080 311 -1079
rect 324 -1080 388 -1079
rect 394 -1080 437 -1079
rect 485 -1080 717 -1079
rect 51 -1082 150 -1081
rect 166 -1082 202 -1081
rect 282 -1082 304 -1081
rect 310 -1082 682 -1081
rect 51 -1084 83 -1083
rect 86 -1084 241 -1083
rect 282 -1084 367 -1083
rect 401 -1084 479 -1083
rect 495 -1084 633 -1083
rect 65 -1086 178 -1085
rect 194 -1086 318 -1085
rect 324 -1086 349 -1085
rect 359 -1086 458 -1085
rect 464 -1086 486 -1085
rect 499 -1086 507 -1085
rect 534 -1086 591 -1085
rect 611 -1086 682 -1085
rect 58 -1088 66 -1087
rect 72 -1088 157 -1087
rect 177 -1088 262 -1087
rect 289 -1088 318 -1087
rect 334 -1088 619 -1087
rect 632 -1088 675 -1087
rect 79 -1090 160 -1089
rect 198 -1090 339 -1089
rect 345 -1090 402 -1089
rect 422 -1090 731 -1089
rect 23 -1092 199 -1091
rect 289 -1092 430 -1091
rect 439 -1092 500 -1091
rect 506 -1092 570 -1091
rect 583 -1092 591 -1091
rect 611 -1092 668 -1091
rect 93 -1094 384 -1093
rect 422 -1094 472 -1093
rect 513 -1094 535 -1093
rect 537 -1094 675 -1093
rect 37 -1096 94 -1095
rect 100 -1096 143 -1095
rect 145 -1096 255 -1095
rect 268 -1096 430 -1095
rect 453 -1096 668 -1095
rect 107 -1098 171 -1097
rect 268 -1098 482 -1097
rect 513 -1098 577 -1097
rect 583 -1098 598 -1097
rect 618 -1098 696 -1097
rect 135 -1100 279 -1099
rect 296 -1100 398 -1099
rect 523 -1100 570 -1099
rect 576 -1100 724 -1099
rect 135 -1102 227 -1101
rect 296 -1102 563 -1101
rect 565 -1102 605 -1101
rect 684 -1102 696 -1101
rect 142 -1104 381 -1103
rect 523 -1104 661 -1103
rect 149 -1106 234 -1105
rect 275 -1106 605 -1105
rect 184 -1108 227 -1107
rect 338 -1108 493 -1107
rect 541 -1108 647 -1107
rect 23 -1110 185 -1109
rect 219 -1110 234 -1109
rect 247 -1110 493 -1109
rect 555 -1110 563 -1109
rect 597 -1110 654 -1109
rect 68 -1112 647 -1111
rect 205 -1114 220 -1113
rect 373 -1114 465 -1113
rect 548 -1114 556 -1113
rect 205 -1116 332 -1115
rect 380 -1116 640 -1115
rect 376 -1118 640 -1117
rect 425 -1120 542 -1119
rect 548 -1120 626 -1119
rect 425 -1122 710 -1121
rect 450 -1124 654 -1123
rect 709 -1124 738 -1123
rect 411 -1126 451 -1125
rect 474 -1126 626 -1125
rect 2 -1137 129 -1136
rect 145 -1137 153 -1136
rect 159 -1137 269 -1136
rect 275 -1137 297 -1136
rect 303 -1137 311 -1136
rect 317 -1137 360 -1136
rect 369 -1137 640 -1136
rect 646 -1137 675 -1136
rect 677 -1137 710 -1136
rect 9 -1139 164 -1138
rect 170 -1139 563 -1138
rect 646 -1139 654 -1138
rect 677 -1139 682 -1138
rect 695 -1139 710 -1138
rect 9 -1141 248 -1140
rect 250 -1141 458 -1140
rect 506 -1141 521 -1140
rect 523 -1141 528 -1140
rect 530 -1141 535 -1140
rect 544 -1141 640 -1140
rect 16 -1143 45 -1142
rect 47 -1143 59 -1142
rect 72 -1143 195 -1142
rect 219 -1143 248 -1142
rect 261 -1143 374 -1142
rect 380 -1143 402 -1142
rect 429 -1143 556 -1142
rect 562 -1143 619 -1142
rect 37 -1145 66 -1144
rect 79 -1145 332 -1144
rect 334 -1145 444 -1144
rect 478 -1145 507 -1144
rect 590 -1145 619 -1144
rect 37 -1147 321 -1146
rect 331 -1147 493 -1146
rect 583 -1147 591 -1146
rect 44 -1149 216 -1148
rect 226 -1149 262 -1148
rect 278 -1149 626 -1148
rect 51 -1151 76 -1150
rect 93 -1151 181 -1150
rect 184 -1151 255 -1150
rect 282 -1151 423 -1150
rect 429 -1151 437 -1150
rect 471 -1151 479 -1150
rect 492 -1151 514 -1150
rect 541 -1151 584 -1150
rect 604 -1151 626 -1150
rect 51 -1153 150 -1152
rect 156 -1153 255 -1152
rect 310 -1153 325 -1152
rect 345 -1153 500 -1152
rect 19 -1155 325 -1154
rect 348 -1155 570 -1154
rect 58 -1157 206 -1156
rect 226 -1157 304 -1156
rect 317 -1157 668 -1156
rect 82 -1159 94 -1158
rect 100 -1159 195 -1158
rect 205 -1159 220 -1158
rect 233 -1159 269 -1158
rect 348 -1159 353 -1158
rect 373 -1159 409 -1158
rect 415 -1159 423 -1158
rect 432 -1159 535 -1158
rect 569 -1159 633 -1158
rect 660 -1159 668 -1158
rect 86 -1161 283 -1160
rect 387 -1161 409 -1160
rect 443 -1161 605 -1160
rect 632 -1161 657 -1160
rect 30 -1163 87 -1162
rect 107 -1163 209 -1162
rect 236 -1163 297 -1162
rect 394 -1163 402 -1162
rect 450 -1163 472 -1162
rect 485 -1163 500 -1162
rect 107 -1165 115 -1164
rect 121 -1165 234 -1164
rect 362 -1165 395 -1164
rect 397 -1165 577 -1164
rect 23 -1167 115 -1166
rect 121 -1167 339 -1166
rect 387 -1167 577 -1166
rect 110 -1169 129 -1168
rect 135 -1169 353 -1168
rect 450 -1169 549 -1168
rect 135 -1171 150 -1170
rect 156 -1171 178 -1170
rect 184 -1171 199 -1170
rect 338 -1171 514 -1170
rect 548 -1171 598 -1170
rect 142 -1173 661 -1172
rect 142 -1175 458 -1174
rect 485 -1175 675 -1174
rect 145 -1177 367 -1176
rect 597 -1177 612 -1176
rect 163 -1179 171 -1178
rect 173 -1179 241 -1178
rect 366 -1179 391 -1178
rect 446 -1179 612 -1178
rect 166 -1181 556 -1180
rect 191 -1183 199 -1182
rect 390 -1183 416 -1182
rect 2 -1194 153 -1193
rect 156 -1194 164 -1193
rect 166 -1194 192 -1193
rect 201 -1194 258 -1193
rect 275 -1194 297 -1193
rect 303 -1194 430 -1193
rect 436 -1194 577 -1193
rect 667 -1194 682 -1193
rect 702 -1194 706 -1193
rect 709 -1194 717 -1193
rect 2 -1196 108 -1195
rect 110 -1196 188 -1195
rect 215 -1196 248 -1195
rect 296 -1196 507 -1195
rect 530 -1196 633 -1195
rect 674 -1196 689 -1195
rect 9 -1198 24 -1197
rect 30 -1198 276 -1197
rect 306 -1198 353 -1197
rect 383 -1198 465 -1197
rect 541 -1198 591 -1197
rect 597 -1198 675 -1197
rect 9 -1200 45 -1199
rect 54 -1200 213 -1199
rect 229 -1200 283 -1199
rect 289 -1200 307 -1199
rect 310 -1200 318 -1199
rect 320 -1200 633 -1199
rect 16 -1202 76 -1201
rect 89 -1202 521 -1201
rect 562 -1202 654 -1201
rect 23 -1204 150 -1203
rect 198 -1204 290 -1203
rect 310 -1204 689 -1203
rect 30 -1206 108 -1205
rect 117 -1206 409 -1205
rect 436 -1206 472 -1205
rect 478 -1206 542 -1205
rect 562 -1206 703 -1205
rect 37 -1208 125 -1207
rect 142 -1208 507 -1207
rect 569 -1208 682 -1207
rect 37 -1210 185 -1209
rect 219 -1210 283 -1209
rect 324 -1210 374 -1209
rect 387 -1210 423 -1209
rect 443 -1210 556 -1209
rect 597 -1210 612 -1209
rect 58 -1212 174 -1211
rect 233 -1212 661 -1211
rect 58 -1214 87 -1213
rect 100 -1214 458 -1213
rect 460 -1214 577 -1213
rect 65 -1216 76 -1215
rect 100 -1216 115 -1215
rect 121 -1216 206 -1215
rect 240 -1216 339 -1215
rect 341 -1216 381 -1215
rect 387 -1216 454 -1215
rect 499 -1216 521 -1215
rect 548 -1216 556 -1215
rect 72 -1218 171 -1217
rect 194 -1218 241 -1217
rect 247 -1218 626 -1217
rect 145 -1220 251 -1219
rect 327 -1220 486 -1219
rect 513 -1220 570 -1219
rect 149 -1222 178 -1221
rect 254 -1222 486 -1221
rect 513 -1222 661 -1221
rect 51 -1224 178 -1223
rect 327 -1224 605 -1223
rect 334 -1226 479 -1225
rect 604 -1226 640 -1225
rect 348 -1228 626 -1227
rect 352 -1230 472 -1229
rect 583 -1230 640 -1229
rect 366 -1232 409 -1231
rect 429 -1232 549 -1231
rect 135 -1234 367 -1233
rect 373 -1234 398 -1233
rect 401 -1234 423 -1233
rect 432 -1234 444 -1233
rect 446 -1234 591 -1233
rect 79 -1236 136 -1235
rect 380 -1236 619 -1235
rect 79 -1238 129 -1237
rect 331 -1238 619 -1237
rect 128 -1240 227 -1239
rect 394 -1240 612 -1239
rect 226 -1242 262 -1241
rect 401 -1242 468 -1241
rect 534 -1242 584 -1241
rect 254 -1244 395 -1243
rect 450 -1244 647 -1243
rect 261 -1246 269 -1245
rect 415 -1246 647 -1245
rect 170 -1248 269 -1247
rect 345 -1248 416 -1247
rect 450 -1248 696 -1247
rect 345 -1250 391 -1249
rect 453 -1250 493 -1249
rect 534 -1250 713 -1249
rect 457 -1252 500 -1251
rect 492 -1254 528 -1253
rect 16 -1265 62 -1264
rect 72 -1265 689 -1264
rect 712 -1265 717 -1264
rect 2 -1267 73 -1266
rect 93 -1267 104 -1266
rect 107 -1267 314 -1266
rect 317 -1267 384 -1266
rect 394 -1267 682 -1266
rect 2 -1269 136 -1268
rect 142 -1269 157 -1268
rect 177 -1269 251 -1268
rect 254 -1269 262 -1268
rect 271 -1269 528 -1268
rect 667 -1269 671 -1268
rect 9 -1271 136 -1270
rect 145 -1271 290 -1270
rect 303 -1271 703 -1270
rect 9 -1273 188 -1272
rect 194 -1273 367 -1272
rect 397 -1273 612 -1272
rect 667 -1273 696 -1272
rect 702 -1273 706 -1272
rect 23 -1275 192 -1274
rect 208 -1275 220 -1274
rect 222 -1275 255 -1274
rect 257 -1275 290 -1274
rect 303 -1275 444 -1274
rect 460 -1275 528 -1274
rect 23 -1277 80 -1276
rect 86 -1277 94 -1276
rect 100 -1277 115 -1276
rect 128 -1277 199 -1276
rect 215 -1277 339 -1276
rect 352 -1277 598 -1276
rect 30 -1279 87 -1278
rect 114 -1279 234 -1278
rect 236 -1279 318 -1278
rect 324 -1279 409 -1278
rect 429 -1279 535 -1278
rect 576 -1279 598 -1278
rect 37 -1281 332 -1280
rect 362 -1281 521 -1280
rect 534 -1281 556 -1280
rect 569 -1281 577 -1280
rect 40 -1283 66 -1282
rect 131 -1283 237 -1282
rect 285 -1283 626 -1282
rect 44 -1285 83 -1284
rect 149 -1285 157 -1284
rect 177 -1285 647 -1284
rect 44 -1287 206 -1286
rect 219 -1287 475 -1286
rect 495 -1287 626 -1286
rect 47 -1289 479 -1288
rect 506 -1289 682 -1288
rect 51 -1291 164 -1290
rect 180 -1291 192 -1290
rect 226 -1291 248 -1290
rect 310 -1291 356 -1290
rect 366 -1291 570 -1290
rect 58 -1293 122 -1292
rect 163 -1293 276 -1292
rect 327 -1293 332 -1292
rect 380 -1293 612 -1292
rect 65 -1295 206 -1294
rect 233 -1295 454 -1294
rect 478 -1295 493 -1294
rect 513 -1295 640 -1294
rect 121 -1297 139 -1296
rect 184 -1297 297 -1296
rect 380 -1297 416 -1296
rect 422 -1297 556 -1296
rect 639 -1297 661 -1296
rect 170 -1299 185 -1298
rect 247 -1299 307 -1298
rect 373 -1299 416 -1298
rect 432 -1299 437 -1298
rect 443 -1299 503 -1298
rect 520 -1299 563 -1298
rect 632 -1299 661 -1298
rect 268 -1301 423 -1300
rect 436 -1301 486 -1300
rect 562 -1301 605 -1300
rect 268 -1303 283 -1302
rect 296 -1303 388 -1302
rect 397 -1303 458 -1302
rect 464 -1303 605 -1302
rect 261 -1305 283 -1304
rect 306 -1305 360 -1304
rect 373 -1305 514 -1304
rect 590 -1305 633 -1304
rect 275 -1307 370 -1306
rect 401 -1307 507 -1306
rect 324 -1309 591 -1308
rect 390 -1311 402 -1310
rect 408 -1311 472 -1310
rect 485 -1311 549 -1310
rect 464 -1313 619 -1312
rect 548 -1315 584 -1314
rect 618 -1315 654 -1314
rect 180 -1317 584 -1316
rect 499 -1319 654 -1318
rect 499 -1321 675 -1320
rect 541 -1323 675 -1322
rect 450 -1325 542 -1324
rect 2 -1336 178 -1335
rect 208 -1336 269 -1335
rect 303 -1336 398 -1335
rect 404 -1336 458 -1335
rect 460 -1336 605 -1335
rect 653 -1336 671 -1335
rect 9 -1338 202 -1337
rect 212 -1338 283 -1337
rect 338 -1338 591 -1337
rect 646 -1338 654 -1337
rect 667 -1338 682 -1337
rect 19 -1340 115 -1339
rect 135 -1340 234 -1339
rect 254 -1340 360 -1339
rect 366 -1340 598 -1339
rect 646 -1340 657 -1339
rect 33 -1342 132 -1341
rect 138 -1342 300 -1341
rect 338 -1342 416 -1341
rect 422 -1342 577 -1341
rect 590 -1342 640 -1341
rect 44 -1344 370 -1343
rect 373 -1344 514 -1343
rect 576 -1344 633 -1343
rect 51 -1346 244 -1345
rect 261 -1346 269 -1345
rect 275 -1346 283 -1345
rect 352 -1346 622 -1345
rect 58 -1348 83 -1347
rect 100 -1348 146 -1347
rect 149 -1348 157 -1347
rect 159 -1348 342 -1347
rect 366 -1348 556 -1347
rect 58 -1350 164 -1349
rect 177 -1350 185 -1349
rect 219 -1350 325 -1349
rect 380 -1350 395 -1349
rect 408 -1350 661 -1349
rect 37 -1352 185 -1351
rect 222 -1352 426 -1351
rect 450 -1352 542 -1351
rect 51 -1354 220 -1353
rect 226 -1354 255 -1353
rect 261 -1354 346 -1353
rect 348 -1354 409 -1353
rect 425 -1354 612 -1353
rect 65 -1356 328 -1355
rect 383 -1356 528 -1355
rect 541 -1356 675 -1355
rect 65 -1358 139 -1357
rect 163 -1358 199 -1357
rect 226 -1358 251 -1357
rect 285 -1358 346 -1357
rect 383 -1358 391 -1357
rect 474 -1358 619 -1357
rect 72 -1360 153 -1359
rect 240 -1360 276 -1359
rect 289 -1360 353 -1359
rect 387 -1360 437 -1359
rect 478 -1360 570 -1359
rect 583 -1360 612 -1359
rect 44 -1362 241 -1361
rect 285 -1362 290 -1361
rect 436 -1362 444 -1361
rect 481 -1362 626 -1361
rect 75 -1364 94 -1363
rect 100 -1364 171 -1363
rect 401 -1364 444 -1363
rect 481 -1364 605 -1363
rect 79 -1366 248 -1365
rect 492 -1366 528 -1365
rect 548 -1366 570 -1365
rect 600 -1366 626 -1365
rect 93 -1368 122 -1367
rect 124 -1368 325 -1367
rect 429 -1368 549 -1367
rect 562 -1368 584 -1367
rect 107 -1370 174 -1369
rect 212 -1370 248 -1369
rect 310 -1370 563 -1369
rect 107 -1372 206 -1371
rect 310 -1372 363 -1371
rect 492 -1372 507 -1371
rect 513 -1372 535 -1371
rect 114 -1374 143 -1373
rect 170 -1374 192 -1373
rect 362 -1374 556 -1373
rect 23 -1376 192 -1375
rect 471 -1376 535 -1375
rect 121 -1378 318 -1377
rect 331 -1378 472 -1377
rect 499 -1378 640 -1377
rect 128 -1380 199 -1379
rect 296 -1380 332 -1379
rect 369 -1380 500 -1379
rect 506 -1380 521 -1379
rect 296 -1382 419 -1381
rect 464 -1382 521 -1381
rect 317 -1384 391 -1383
rect 33 -1395 220 -1394
rect 233 -1395 297 -1394
rect 317 -1395 356 -1394
rect 366 -1395 451 -1394
rect 453 -1395 570 -1394
rect 600 -1395 668 -1394
rect 37 -1397 206 -1396
rect 233 -1397 521 -1396
rect 551 -1397 591 -1396
rect 621 -1397 640 -1396
rect 37 -1399 311 -1398
rect 317 -1399 328 -1398
rect 373 -1399 388 -1398
rect 390 -1399 444 -1398
rect 460 -1399 598 -1398
rect 635 -1399 661 -1398
rect 44 -1401 370 -1400
rect 380 -1401 486 -1400
rect 499 -1401 591 -1400
rect 44 -1403 139 -1402
rect 184 -1403 353 -1402
rect 369 -1403 563 -1402
rect 51 -1405 272 -1404
rect 275 -1405 286 -1404
rect 296 -1405 325 -1404
rect 331 -1405 381 -1404
rect 387 -1405 430 -1404
rect 432 -1405 535 -1404
rect 51 -1407 115 -1406
rect 124 -1407 136 -1406
rect 201 -1407 402 -1406
rect 404 -1407 430 -1406
rect 436 -1407 458 -1406
rect 464 -1407 507 -1406
rect 513 -1407 535 -1406
rect 58 -1409 157 -1408
rect 247 -1409 549 -1408
rect 58 -1411 164 -1410
rect 247 -1411 451 -1410
rect 464 -1411 584 -1410
rect 72 -1413 237 -1412
rect 261 -1413 377 -1412
rect 394 -1413 416 -1412
rect 418 -1413 528 -1412
rect 583 -1413 626 -1412
rect 72 -1415 150 -1414
rect 163 -1415 178 -1414
rect 187 -1415 395 -1414
rect 401 -1415 444 -1414
rect 485 -1415 542 -1414
rect 86 -1417 104 -1416
rect 107 -1417 346 -1416
rect 397 -1417 542 -1416
rect 79 -1419 87 -1418
rect 103 -1419 290 -1418
rect 310 -1419 374 -1418
rect 422 -1419 566 -1418
rect 79 -1421 227 -1420
rect 243 -1421 528 -1420
rect 107 -1423 122 -1422
rect 138 -1423 150 -1422
rect 177 -1423 360 -1422
rect 425 -1423 521 -1422
rect 205 -1425 227 -1424
rect 254 -1425 262 -1424
rect 268 -1425 367 -1424
rect 436 -1425 577 -1424
rect 219 -1427 269 -1426
rect 275 -1427 384 -1426
rect 492 -1427 507 -1426
rect 513 -1427 556 -1426
rect 576 -1427 612 -1426
rect 191 -1429 556 -1428
rect 191 -1431 213 -1430
rect 240 -1431 255 -1430
rect 282 -1431 500 -1430
rect 65 -1433 213 -1432
rect 215 -1433 283 -1432
rect 289 -1433 304 -1432
rect 331 -1433 339 -1432
rect 471 -1433 493 -1432
rect 65 -1435 171 -1434
rect 338 -1435 447 -1434
rect 128 -1437 304 -1436
rect 439 -1437 472 -1436
rect 117 -1439 129 -1438
rect 145 -1439 171 -1438
rect 145 -1441 409 -1440
rect 408 -1443 549 -1442
rect 16 -1454 178 -1453
rect 215 -1454 388 -1453
rect 429 -1454 570 -1453
rect 702 -1454 713 -1453
rect 44 -1456 118 -1455
rect 163 -1456 199 -1455
rect 254 -1456 307 -1455
rect 310 -1456 440 -1455
rect 443 -1456 535 -1455
rect 548 -1456 591 -1455
rect 51 -1458 181 -1457
rect 254 -1458 311 -1457
rect 327 -1458 332 -1457
rect 359 -1458 416 -1457
rect 422 -1458 444 -1457
rect 450 -1458 493 -1457
rect 562 -1458 605 -1457
rect 65 -1460 244 -1459
rect 268 -1460 395 -1459
rect 432 -1460 486 -1459
rect 492 -1460 528 -1459
rect 565 -1460 598 -1459
rect 51 -1462 66 -1461
rect 72 -1462 234 -1461
rect 271 -1462 409 -1461
rect 436 -1462 507 -1461
rect 534 -1462 566 -1461
rect 569 -1462 584 -1461
rect 72 -1464 192 -1463
rect 212 -1464 234 -1463
rect 240 -1464 409 -1463
rect 478 -1464 521 -1463
rect 572 -1464 584 -1463
rect 58 -1466 241 -1465
rect 271 -1466 304 -1465
rect 331 -1466 458 -1465
rect 478 -1466 542 -1465
rect 58 -1468 248 -1467
rect 282 -1468 367 -1467
rect 401 -1468 486 -1467
rect 506 -1468 563 -1467
rect 79 -1470 185 -1469
rect 250 -1470 402 -1469
rect 457 -1470 500 -1469
rect 520 -1470 577 -1469
rect 79 -1472 220 -1471
rect 261 -1472 283 -1471
rect 289 -1472 388 -1471
rect 429 -1472 500 -1471
rect 541 -1472 556 -1471
rect 576 -1472 591 -1471
rect 37 -1474 290 -1473
rect 292 -1474 374 -1473
rect 37 -1476 45 -1475
rect 86 -1476 157 -1475
rect 163 -1476 227 -1475
rect 261 -1476 339 -1475
rect 345 -1476 416 -1475
rect 30 -1478 87 -1477
rect 93 -1478 136 -1477
rect 142 -1478 199 -1477
rect 205 -1478 220 -1477
rect 296 -1478 346 -1477
rect 359 -1478 381 -1477
rect 93 -1480 108 -1479
rect 110 -1480 143 -1479
rect 149 -1480 192 -1479
rect 296 -1480 465 -1479
rect 100 -1482 426 -1481
rect 107 -1484 167 -1483
rect 170 -1484 230 -1483
rect 338 -1484 472 -1483
rect 114 -1486 129 -1485
rect 135 -1486 276 -1485
rect 369 -1486 556 -1485
rect 128 -1488 160 -1487
rect 177 -1488 353 -1487
rect 380 -1488 447 -1487
rect 471 -1488 514 -1487
rect 124 -1490 514 -1489
rect 156 -1492 528 -1491
rect 275 -1494 325 -1493
rect 390 -1494 465 -1493
rect 317 -1496 325 -1495
rect 16 -1507 171 -1506
rect 173 -1507 199 -1506
rect 205 -1507 276 -1506
rect 292 -1507 444 -1506
rect 464 -1507 475 -1506
rect 478 -1507 514 -1506
rect 565 -1507 570 -1506
rect 579 -1507 584 -1506
rect 23 -1509 55 -1508
rect 58 -1509 122 -1508
rect 142 -1509 178 -1508
rect 184 -1509 360 -1508
rect 369 -1509 437 -1508
rect 443 -1509 451 -1508
rect 488 -1509 556 -1508
rect 30 -1511 59 -1510
rect 72 -1511 150 -1510
rect 152 -1511 171 -1510
rect 184 -1511 290 -1510
rect 313 -1511 416 -1510
rect 422 -1511 521 -1510
rect 37 -1513 52 -1512
rect 79 -1513 122 -1512
rect 152 -1513 202 -1512
rect 240 -1513 542 -1512
rect 51 -1515 94 -1514
rect 100 -1515 143 -1514
rect 163 -1515 241 -1514
rect 247 -1515 304 -1514
rect 320 -1515 493 -1514
rect 513 -1515 549 -1514
rect 65 -1517 80 -1516
rect 86 -1517 255 -1516
rect 268 -1517 283 -1516
rect 303 -1517 346 -1516
rect 401 -1517 426 -1516
rect 429 -1517 465 -1516
rect 492 -1517 528 -1516
rect 65 -1519 209 -1518
rect 275 -1519 374 -1518
rect 387 -1519 528 -1518
rect 89 -1521 181 -1520
rect 187 -1521 255 -1520
rect 282 -1521 311 -1520
rect 327 -1521 486 -1520
rect 520 -1521 563 -1520
rect 110 -1523 129 -1522
rect 135 -1523 248 -1522
rect 261 -1523 311 -1522
rect 331 -1523 360 -1522
rect 373 -1523 381 -1522
rect 383 -1523 388 -1522
rect 436 -1523 458 -1522
rect 114 -1525 157 -1524
rect 191 -1525 206 -1524
rect 229 -1525 262 -1524
rect 380 -1525 402 -1524
rect 450 -1525 472 -1524
rect 96 -1527 115 -1526
rect 128 -1527 220 -1526
rect 236 -1527 332 -1526
rect 457 -1527 500 -1526
rect 135 -1529 297 -1528
rect 499 -1529 535 -1528
rect 156 -1531 430 -1530
rect 198 -1533 213 -1532
rect 236 -1533 346 -1532
rect 212 -1535 230 -1534
rect 296 -1535 318 -1534
rect 317 -1537 409 -1536
rect 352 -1539 409 -1538
rect 352 -1541 395 -1540
rect 338 -1543 395 -1542
rect 338 -1545 577 -1544
rect 51 -1556 108 -1555
rect 121 -1556 244 -1555
rect 261 -1556 286 -1555
rect 289 -1556 346 -1555
rect 359 -1556 388 -1555
rect 415 -1556 437 -1555
rect 450 -1556 472 -1555
rect 485 -1556 521 -1555
rect 586 -1556 591 -1555
rect 72 -1558 80 -1557
rect 86 -1558 223 -1557
rect 226 -1558 234 -1557
rect 236 -1558 248 -1557
rect 261 -1558 269 -1557
rect 271 -1558 360 -1557
rect 380 -1558 493 -1557
rect 75 -1560 80 -1559
rect 96 -1560 367 -1559
rect 422 -1560 503 -1559
rect 103 -1562 115 -1561
rect 128 -1562 328 -1561
rect 429 -1562 500 -1561
rect 149 -1564 178 -1563
rect 194 -1564 297 -1563
rect 310 -1564 370 -1563
rect 429 -1564 465 -1563
rect 492 -1564 507 -1563
rect 142 -1566 195 -1565
rect 198 -1566 223 -1565
rect 240 -1566 339 -1565
rect 369 -1566 395 -1565
rect 436 -1566 444 -1565
rect 457 -1566 465 -1565
rect 142 -1568 192 -1567
rect 205 -1568 230 -1567
rect 247 -1568 314 -1567
rect 317 -1568 391 -1567
rect 128 -1570 192 -1569
rect 219 -1570 255 -1569
rect 275 -1570 297 -1569
rect 317 -1570 479 -1569
rect 159 -1572 213 -1571
rect 254 -1572 283 -1571
rect 292 -1572 528 -1571
rect 65 -1574 160 -1573
rect 163 -1574 171 -1573
rect 173 -1574 202 -1573
rect 275 -1574 367 -1573
rect 373 -1574 395 -1573
rect 135 -1576 213 -1575
rect 324 -1576 381 -1575
rect 135 -1578 153 -1577
rect 163 -1578 185 -1577
rect 373 -1578 409 -1577
rect 152 -1580 178 -1579
rect 156 -1582 185 -1581
rect 72 -1593 83 -1592
rect 89 -1593 94 -1592
rect 128 -1593 157 -1592
rect 163 -1593 206 -1592
rect 219 -1593 241 -1592
rect 243 -1593 262 -1592
rect 282 -1593 290 -1592
rect 296 -1593 311 -1592
rect 320 -1593 339 -1592
rect 345 -1593 353 -1592
rect 366 -1593 374 -1592
rect 383 -1593 430 -1592
rect 471 -1593 486 -1592
rect 506 -1593 514 -1592
rect 75 -1595 80 -1594
rect 135 -1595 153 -1594
rect 163 -1595 195 -1594
rect 205 -1595 248 -1594
rect 254 -1595 370 -1594
rect 422 -1595 437 -1594
rect 443 -1595 486 -1594
rect 114 -1597 153 -1596
rect 177 -1597 269 -1596
rect 275 -1597 290 -1596
rect 317 -1597 346 -1596
rect 352 -1597 381 -1596
rect 464 -1597 472 -1596
rect 131 -1599 136 -1598
rect 142 -1599 146 -1598
rect 156 -1599 276 -1598
rect 282 -1599 311 -1598
rect 317 -1599 360 -1598
rect 184 -1601 216 -1600
rect 226 -1601 325 -1600
rect 331 -1601 335 -1600
rect 338 -1601 402 -1600
rect 191 -1603 202 -1602
rect 212 -1603 297 -1602
rect 299 -1603 360 -1602
rect 191 -1605 209 -1604
rect 226 -1605 342 -1604
rect 233 -1607 255 -1606
rect 261 -1607 304 -1606
rect 236 -1609 279 -1608
rect 240 -1611 269 -1610
rect 243 -1613 325 -1612
rect 250 -1615 304 -1614
rect 30 -1626 34 -1625
rect 37 -1626 181 -1625
rect 198 -1626 216 -1625
rect 233 -1626 237 -1625
rect 240 -1626 272 -1625
rect 275 -1626 318 -1625
rect 334 -1626 367 -1625
rect 401 -1626 444 -1625
rect 467 -1626 472 -1625
rect 488 -1626 493 -1625
rect 44 -1628 157 -1627
rect 177 -1628 220 -1627
rect 254 -1628 258 -1627
rect 261 -1628 353 -1627
rect 359 -1628 381 -1627
rect 51 -1630 87 -1629
rect 93 -1630 101 -1629
rect 121 -1630 143 -1629
rect 149 -1630 164 -1629
rect 177 -1630 202 -1629
rect 212 -1630 248 -1629
rect 254 -1630 290 -1629
rect 296 -1630 325 -1629
rect 327 -1630 353 -1629
rect 65 -1632 111 -1631
rect 124 -1632 136 -1631
rect 138 -1632 171 -1631
rect 191 -1632 241 -1631
rect 257 -1632 290 -1631
rect 303 -1632 360 -1631
rect 72 -1634 90 -1633
rect 100 -1634 125 -1633
rect 135 -1634 157 -1633
rect 163 -1634 227 -1633
rect 264 -1634 318 -1633
rect 345 -1634 367 -1633
rect 72 -1636 132 -1635
rect 170 -1636 230 -1635
rect 275 -1636 339 -1635
rect 345 -1636 405 -1635
rect 79 -1638 115 -1637
rect 198 -1638 223 -1637
rect 226 -1638 297 -1637
rect 303 -1638 311 -1637
rect 58 -1640 115 -1639
rect 219 -1640 332 -1639
rect 86 -1642 146 -1641
rect 278 -1642 374 -1641
rect 107 -1644 150 -1643
rect 282 -1644 311 -1643
rect 19 -1655 24 -1654
rect 37 -1655 223 -1654
rect 226 -1655 367 -1654
rect 387 -1655 391 -1654
rect 44 -1657 129 -1656
rect 149 -1657 216 -1656
rect 219 -1657 241 -1656
rect 243 -1657 262 -1656
rect 268 -1657 311 -1656
rect 317 -1657 402 -1656
rect 51 -1659 139 -1658
rect 163 -1659 185 -1658
rect 191 -1659 199 -1658
rect 212 -1659 290 -1658
rect 296 -1659 311 -1658
rect 324 -1659 374 -1658
rect 65 -1661 94 -1660
rect 100 -1661 136 -1660
rect 156 -1661 164 -1660
rect 212 -1661 297 -1660
rect 331 -1661 374 -1660
rect 72 -1663 97 -1662
rect 103 -1663 108 -1662
rect 117 -1663 192 -1662
rect 226 -1663 325 -1662
rect 331 -1663 346 -1662
rect 366 -1663 381 -1662
rect 79 -1665 125 -1664
rect 156 -1665 171 -1664
rect 222 -1665 381 -1664
rect 86 -1667 115 -1666
rect 121 -1667 146 -1666
rect 229 -1667 321 -1666
rect 338 -1667 395 -1666
rect 121 -1669 178 -1668
rect 205 -1669 395 -1668
rect 145 -1671 150 -1670
rect 205 -1671 272 -1670
rect 282 -1671 353 -1670
rect 233 -1673 248 -1672
rect 254 -1673 269 -1672
rect 285 -1673 339 -1672
rect 348 -1673 353 -1672
rect 208 -1675 248 -1674
rect 261 -1675 304 -1674
rect 236 -1677 360 -1676
rect 240 -1679 276 -1678
rect 2 -1690 10 -1689
rect 16 -1690 24 -1689
rect 30 -1690 34 -1689
rect 89 -1690 97 -1689
rect 100 -1690 108 -1689
rect 114 -1690 206 -1689
rect 222 -1690 244 -1689
rect 254 -1690 402 -1689
rect 121 -1692 213 -1691
rect 226 -1692 234 -1691
rect 257 -1692 297 -1691
rect 317 -1692 332 -1691
rect 359 -1692 374 -1691
rect 121 -1694 129 -1693
rect 156 -1694 185 -1693
rect 191 -1694 248 -1693
rect 264 -1694 311 -1693
rect 135 -1696 157 -1695
rect 163 -1696 171 -1695
rect 194 -1696 206 -1695
rect 226 -1696 325 -1695
rect 131 -1698 136 -1697
rect 149 -1698 164 -1697
rect 170 -1698 178 -1697
rect 198 -1698 220 -1697
rect 229 -1698 234 -1697
rect 268 -1698 286 -1697
rect 292 -1698 381 -1697
rect 117 -1700 132 -1699
rect 173 -1700 178 -1699
rect 201 -1700 213 -1699
rect 275 -1700 279 -1699
rect 285 -1700 290 -1699
rect 296 -1700 395 -1699
rect 303 -1702 311 -1701
rect 324 -1702 339 -1701
rect 5 -1713 10 -1712
rect 128 -1713 136 -1712
rect 142 -1713 164 -1712
rect 170 -1713 202 -1712
rect 212 -1713 220 -1712
rect 233 -1713 244 -1712
rect 303 -1713 311 -1712
rect 317 -1713 325 -1712
rect 152 -1715 157 -1714
rect 177 -1715 227 -1714
rect 187 -1717 206 -1716
<< m2contact >>
rect 177 0 178 1
rect 187 0 188 1
rect 198 0 199 1
rect 205 0 206 1
rect 208 0 209 1
rect 222 0 223 1
rect 240 0 241 1
rect 247 0 248 1
rect 275 0 276 1
rect 282 0 283 1
rect 289 0 290 1
rect 299 0 300 1
rect 215 -2 216 -1
rect 233 -2 234 -1
rect 243 -2 244 -1
rect 254 -2 255 -1
rect 107 -13 108 -12
rect 110 -13 111 -12
rect 142 -13 143 -12
rect 170 -13 171 -12
rect 177 -13 178 -12
rect 194 -13 195 -12
rect 219 -13 220 -12
rect 233 -13 234 -12
rect 254 -13 255 -12
rect 268 -13 269 -12
rect 289 -13 290 -12
rect 303 -13 304 -12
rect 149 -15 150 -14
rect 159 -15 160 -14
rect 163 -15 164 -14
rect 194 -15 195 -14
rect 208 -15 209 -14
rect 219 -15 220 -14
rect 226 -15 227 -14
rect 247 -15 248 -14
rect 264 -15 265 -14
rect 275 -15 276 -14
rect 282 -15 283 -14
rect 289 -15 290 -14
rect 292 -15 293 -14
rect 310 -15 311 -14
rect 184 -17 185 -16
rect 208 -17 209 -16
rect 240 -17 241 -16
rect 247 -17 248 -16
rect 296 -17 297 -16
rect 299 -17 300 -16
rect 191 -19 192 -18
rect 198 -19 199 -18
rect 198 -21 199 -20
rect 215 -21 216 -20
rect 135 -32 136 -31
rect 145 -32 146 -31
rect 152 -32 153 -31
rect 156 -32 157 -31
rect 177 -32 178 -31
rect 226 -32 227 -31
rect 233 -32 234 -31
rect 243 -32 244 -31
rect 247 -32 248 -31
rect 261 -32 262 -31
rect 282 -32 283 -31
rect 292 -32 293 -31
rect 296 -32 297 -31
rect 303 -32 304 -31
rect 310 -32 311 -31
rect 324 -32 325 -31
rect 478 -32 479 -31
rect 485 -32 486 -31
rect 579 -32 580 -31
rect 583 -32 584 -31
rect 142 -34 143 -33
rect 180 -34 181 -33
rect 191 -34 192 -33
rect 198 -34 199 -33
rect 212 -34 213 -33
rect 219 -34 220 -33
rect 240 -34 241 -33
rect 254 -34 255 -33
rect 257 -34 258 -33
rect 268 -34 269 -33
rect 285 -34 286 -33
rect 289 -34 290 -33
rect 296 -34 297 -33
rect 303 -34 304 -33
rect 317 -34 318 -33
rect 320 -34 321 -33
rect 79 -45 80 -44
rect 82 -45 83 -44
rect 135 -45 136 -44
rect 152 -45 153 -44
rect 170 -45 171 -44
rect 173 -45 174 -44
rect 184 -45 185 -44
rect 194 -45 195 -44
rect 212 -45 213 -44
rect 215 -45 216 -44
rect 219 -45 220 -44
rect 233 -45 234 -44
rect 240 -45 241 -44
rect 282 -45 283 -44
rect 289 -45 290 -44
rect 320 -45 321 -44
rect 338 -45 339 -44
rect 345 -45 346 -44
rect 352 -45 353 -44
rect 362 -45 363 -44
rect 467 -45 468 -44
rect 471 -45 472 -44
rect 478 -45 479 -44
rect 485 -45 486 -44
rect 576 -45 577 -44
rect 583 -45 584 -44
rect 177 -47 178 -46
rect 194 -47 195 -46
rect 212 -47 213 -46
rect 243 -47 244 -46
rect 247 -47 248 -46
rect 268 -47 269 -46
rect 292 -47 293 -46
rect 317 -47 318 -46
rect 184 -49 185 -48
rect 205 -49 206 -48
rect 222 -49 223 -48
rect 226 -49 227 -48
rect 233 -49 234 -48
rect 261 -49 262 -48
rect 310 -49 311 -48
rect 324 -49 325 -48
rect 229 -51 230 -50
rect 261 -51 262 -50
rect 317 -51 318 -50
rect 341 -51 342 -50
rect 247 -53 248 -52
rect 268 -53 269 -52
rect 324 -53 325 -52
rect 334 -53 335 -52
rect 250 -55 251 -54
rect 275 -55 276 -54
rect 275 -57 276 -56
rect 282 -57 283 -56
rect 142 -68 143 -67
rect 149 -68 150 -67
rect 205 -68 206 -67
rect 212 -68 213 -67
rect 219 -68 220 -67
rect 243 -68 244 -67
rect 247 -68 248 -67
rect 261 -68 262 -67
rect 268 -68 269 -67
rect 282 -68 283 -67
rect 338 -68 339 -67
rect 345 -68 346 -67
rect 474 -68 475 -67
rect 485 -68 486 -67
rect 138 -70 139 -69
rect 219 -70 220 -69
rect 226 -70 227 -69
rect 233 -70 234 -69
rect 240 -70 241 -69
rect 289 -70 290 -69
rect 345 -70 346 -69
rect 352 -70 353 -69
rect 142 -72 143 -71
rect 163 -72 164 -71
rect 166 -72 167 -71
rect 205 -72 206 -71
rect 226 -72 227 -71
rect 275 -72 276 -71
rect 278 -72 279 -71
rect 296 -72 297 -71
rect 320 -72 321 -71
rect 352 -72 353 -71
rect 149 -74 150 -73
rect 156 -74 157 -73
rect 236 -74 237 -73
rect 289 -74 290 -73
rect 296 -74 297 -73
rect 303 -74 304 -73
rect 247 -76 248 -75
rect 254 -76 255 -75
rect 261 -76 262 -75
rect 310 -76 311 -75
rect 240 -78 241 -77
rect 254 -78 255 -77
rect 268 -78 269 -77
rect 306 -78 307 -77
rect 275 -80 276 -79
rect 317 -80 318 -79
rect 128 -91 129 -90
rect 135 -91 136 -90
rect 142 -91 143 -90
rect 145 -91 146 -90
rect 149 -91 150 -90
rect 159 -91 160 -90
rect 163 -91 164 -90
rect 226 -91 227 -90
rect 233 -91 234 -90
rect 268 -91 269 -90
rect 271 -91 272 -90
rect 359 -91 360 -90
rect 397 -91 398 -90
rect 422 -91 423 -90
rect 481 -91 482 -90
rect 485 -91 486 -90
rect 576 -91 577 -90
rect 583 -91 584 -90
rect 107 -93 108 -92
rect 142 -93 143 -92
rect 152 -93 153 -92
rect 156 -93 157 -92
rect 166 -93 167 -92
rect 170 -93 171 -92
rect 177 -93 178 -92
rect 184 -93 185 -92
rect 187 -93 188 -92
rect 198 -93 199 -92
rect 205 -93 206 -92
rect 243 -93 244 -92
rect 257 -93 258 -92
rect 261 -93 262 -92
rect 289 -93 290 -92
rect 324 -93 325 -92
rect 338 -93 339 -92
rect 348 -93 349 -92
rect 352 -93 353 -92
rect 380 -93 381 -92
rect 478 -93 479 -92
rect 485 -93 486 -92
rect 576 -93 577 -92
rect 590 -93 591 -92
rect 191 -95 192 -94
rect 201 -95 202 -94
rect 219 -95 220 -94
rect 303 -95 304 -94
rect 310 -95 311 -94
rect 366 -95 367 -94
rect 478 -95 479 -94
rect 492 -95 493 -94
rect 194 -97 195 -96
rect 226 -97 227 -96
rect 240 -97 241 -96
rect 317 -97 318 -96
rect 341 -97 342 -96
rect 345 -97 346 -96
rect 212 -99 213 -98
rect 219 -99 220 -98
rect 222 -99 223 -98
rect 352 -99 353 -98
rect 212 -101 213 -100
rect 233 -101 234 -100
rect 243 -101 244 -100
rect 247 -101 248 -100
rect 250 -101 251 -100
rect 324 -101 325 -100
rect 338 -101 339 -100
rect 345 -101 346 -100
rect 254 -103 255 -102
rect 261 -103 262 -102
rect 275 -103 276 -102
rect 310 -103 311 -102
rect 317 -103 318 -102
rect 373 -103 374 -102
rect 254 -105 255 -104
rect 320 -105 321 -104
rect 296 -107 297 -106
rect 331 -107 332 -106
rect 282 -109 283 -108
rect 296 -109 297 -108
rect 180 -111 181 -110
rect 282 -111 283 -110
rect 65 -122 66 -121
rect 107 -122 108 -121
rect 131 -122 132 -121
rect 135 -122 136 -121
rect 145 -122 146 -121
rect 170 -122 171 -121
rect 173 -122 174 -121
rect 184 -122 185 -121
rect 191 -122 192 -121
rect 205 -122 206 -121
rect 208 -122 209 -121
rect 254 -122 255 -121
rect 264 -122 265 -121
rect 278 -122 279 -121
rect 289 -122 290 -121
rect 317 -122 318 -121
rect 324 -122 325 -121
rect 338 -122 339 -121
rect 359 -122 360 -121
rect 415 -122 416 -121
rect 422 -122 423 -121
rect 443 -122 444 -121
rect 478 -122 479 -121
rect 485 -122 486 -121
rect 492 -122 493 -121
rect 499 -122 500 -121
rect 576 -122 577 -121
rect 583 -122 584 -121
rect 72 -124 73 -123
rect 100 -124 101 -123
rect 107 -124 108 -123
rect 114 -124 115 -123
rect 128 -124 129 -123
rect 135 -124 136 -123
rect 149 -124 150 -123
rect 156 -124 157 -123
rect 163 -124 164 -123
rect 236 -124 237 -123
rect 243 -124 244 -123
rect 310 -124 311 -123
rect 331 -124 332 -123
rect 422 -124 423 -123
rect 86 -126 87 -125
rect 124 -126 125 -125
rect 170 -126 171 -125
rect 208 -126 209 -125
rect 219 -126 220 -125
rect 366 -126 367 -125
rect 380 -126 381 -125
rect 429 -126 430 -125
rect 93 -128 94 -127
rect 243 -128 244 -127
rect 275 -128 276 -127
rect 373 -128 374 -127
rect 387 -128 388 -127
rect 436 -128 437 -127
rect 156 -130 157 -129
rect 219 -130 220 -129
rect 222 -130 223 -129
rect 233 -130 234 -129
rect 282 -130 283 -129
rect 310 -130 311 -129
rect 334 -130 335 -129
rect 366 -130 367 -129
rect 394 -130 395 -129
rect 401 -130 402 -129
rect 177 -132 178 -131
rect 285 -132 286 -131
rect 299 -132 300 -131
rect 359 -132 360 -131
rect 184 -134 185 -133
rect 233 -134 234 -133
rect 303 -134 304 -133
rect 373 -134 374 -133
rect 191 -136 192 -135
rect 226 -136 227 -135
rect 229 -136 230 -135
rect 289 -136 290 -135
rect 352 -136 353 -135
rect 380 -136 381 -135
rect 198 -138 199 -137
rect 212 -138 213 -137
rect 222 -138 223 -137
rect 324 -138 325 -137
rect 352 -138 353 -137
rect 394 -138 395 -137
rect 198 -140 199 -139
rect 261 -140 262 -139
rect 205 -142 206 -141
rect 247 -142 248 -141
rect 261 -142 262 -141
rect 296 -142 297 -141
rect 226 -144 227 -143
rect 268 -144 269 -143
rect 240 -146 241 -145
rect 303 -146 304 -145
rect 240 -148 241 -147
rect 275 -148 276 -147
rect 257 -150 258 -149
rect 268 -150 269 -149
rect 19 -161 20 -160
rect 26 -161 27 -160
rect 65 -161 66 -160
rect 114 -161 115 -160
rect 131 -161 132 -160
rect 159 -161 160 -160
rect 163 -161 164 -160
rect 247 -161 248 -160
rect 264 -161 265 -160
rect 310 -161 311 -160
rect 317 -161 318 -160
rect 331 -161 332 -160
rect 352 -161 353 -160
rect 429 -161 430 -160
rect 499 -161 500 -160
rect 506 -161 507 -160
rect 72 -163 73 -162
rect 121 -163 122 -162
rect 149 -163 150 -162
rect 180 -163 181 -162
rect 208 -163 209 -162
rect 415 -163 416 -162
rect 79 -165 80 -164
rect 128 -165 129 -164
rect 149 -165 150 -164
rect 156 -165 157 -164
rect 219 -165 220 -164
rect 310 -165 311 -164
rect 320 -165 321 -164
rect 436 -165 437 -164
rect 79 -167 80 -166
rect 124 -167 125 -166
rect 128 -167 129 -166
rect 184 -167 185 -166
rect 226 -167 227 -166
rect 247 -167 248 -166
rect 268 -167 269 -166
rect 436 -167 437 -166
rect 86 -169 87 -168
rect 166 -169 167 -168
rect 226 -169 227 -168
rect 331 -169 332 -168
rect 345 -169 346 -168
rect 429 -169 430 -168
rect 93 -171 94 -170
rect 145 -171 146 -170
rect 236 -171 237 -170
rect 268 -171 269 -170
rect 278 -171 279 -170
rect 460 -171 461 -170
rect 100 -173 101 -172
rect 177 -173 178 -172
rect 243 -173 244 -172
rect 338 -173 339 -172
rect 352 -173 353 -172
rect 387 -173 388 -172
rect 103 -175 104 -174
rect 142 -175 143 -174
rect 177 -175 178 -174
rect 205 -175 206 -174
rect 212 -175 213 -174
rect 338 -175 339 -174
rect 359 -175 360 -174
rect 415 -175 416 -174
rect 86 -177 87 -176
rect 142 -177 143 -176
rect 212 -177 213 -176
rect 296 -177 297 -176
rect 299 -177 300 -176
rect 422 -177 423 -176
rect 107 -179 108 -178
rect 163 -179 164 -178
rect 282 -179 283 -178
rect 317 -179 318 -178
rect 324 -179 325 -178
rect 345 -179 346 -178
rect 373 -179 374 -178
rect 464 -179 465 -178
rect 107 -181 108 -180
rect 198 -181 199 -180
rect 254 -181 255 -180
rect 324 -181 325 -180
rect 373 -181 374 -180
rect 408 -181 409 -180
rect 422 -181 423 -180
rect 443 -181 444 -180
rect 114 -183 115 -182
rect 170 -183 171 -182
rect 191 -183 192 -182
rect 254 -183 255 -182
rect 299 -183 300 -182
rect 387 -183 388 -182
rect 401 -183 402 -182
rect 408 -183 409 -182
rect 93 -185 94 -184
rect 170 -185 171 -184
rect 243 -185 244 -184
rect 443 -185 444 -184
rect 121 -187 122 -186
rect 156 -187 157 -186
rect 303 -187 304 -186
rect 359 -187 360 -186
rect 394 -187 395 -186
rect 401 -187 402 -186
rect 191 -189 192 -188
rect 303 -189 304 -188
rect 380 -189 381 -188
rect 394 -189 395 -188
rect 261 -191 262 -190
rect 380 -191 381 -190
rect 240 -193 241 -192
rect 261 -193 262 -192
rect 240 -195 241 -194
rect 275 -195 276 -194
rect 275 -197 276 -196
rect 289 -197 290 -196
rect 233 -199 234 -198
rect 289 -199 290 -198
rect 79 -210 80 -209
rect 222 -210 223 -209
rect 243 -210 244 -209
rect 324 -210 325 -209
rect 348 -210 349 -209
rect 415 -210 416 -209
rect 443 -210 444 -209
rect 453 -210 454 -209
rect 506 -210 507 -209
rect 509 -210 510 -209
rect 562 -210 563 -209
rect 572 -210 573 -209
rect 86 -212 87 -211
rect 215 -212 216 -211
rect 219 -212 220 -211
rect 338 -212 339 -211
rect 380 -212 381 -211
rect 422 -212 423 -211
rect 450 -212 451 -211
rect 460 -212 461 -211
rect 100 -214 101 -213
rect 240 -214 241 -213
rect 278 -214 279 -213
rect 436 -214 437 -213
rect 107 -216 108 -215
rect 236 -216 237 -215
rect 240 -216 241 -215
rect 254 -216 255 -215
rect 296 -216 297 -215
rect 373 -216 374 -215
rect 383 -216 384 -215
rect 394 -216 395 -215
rect 114 -218 115 -217
rect 191 -218 192 -217
rect 222 -218 223 -217
rect 464 -218 465 -217
rect 114 -220 115 -219
rect 201 -220 202 -219
rect 236 -220 237 -219
rect 282 -220 283 -219
rect 317 -220 318 -219
rect 352 -220 353 -219
rect 359 -220 360 -219
rect 373 -220 374 -219
rect 128 -222 129 -221
rect 198 -222 199 -221
rect 212 -222 213 -221
rect 317 -222 318 -221
rect 320 -222 321 -221
rect 415 -222 416 -221
rect 135 -224 136 -223
rect 145 -224 146 -223
rect 156 -224 157 -223
rect 226 -224 227 -223
rect 243 -224 244 -223
rect 436 -224 437 -223
rect 128 -226 129 -225
rect 156 -226 157 -225
rect 163 -226 164 -225
rect 275 -226 276 -225
rect 282 -226 283 -225
rect 303 -226 304 -225
rect 324 -226 325 -225
rect 345 -226 346 -225
rect 135 -228 136 -227
rect 166 -228 167 -227
rect 173 -228 174 -227
rect 264 -228 265 -227
rect 289 -228 290 -227
rect 303 -228 304 -227
rect 331 -228 332 -227
rect 443 -228 444 -227
rect 142 -230 143 -229
rect 184 -230 185 -229
rect 191 -230 192 -229
rect 247 -230 248 -229
rect 254 -230 255 -229
rect 261 -230 262 -229
rect 292 -230 293 -229
rect 331 -230 332 -229
rect 338 -230 339 -229
rect 366 -230 367 -229
rect 177 -232 178 -231
rect 215 -232 216 -231
rect 226 -232 227 -231
rect 247 -232 248 -231
rect 261 -232 262 -231
rect 394 -232 395 -231
rect 184 -234 185 -233
rect 205 -234 206 -233
rect 212 -234 213 -233
rect 292 -234 293 -233
rect 296 -234 297 -233
rect 359 -234 360 -233
rect 198 -236 199 -235
rect 310 -236 311 -235
rect 345 -236 346 -235
rect 429 -236 430 -235
rect 278 -238 279 -237
rect 310 -238 311 -237
rect 352 -238 353 -237
rect 366 -238 367 -237
rect 387 -238 388 -237
rect 429 -238 430 -237
rect 275 -240 276 -239
rect 387 -240 388 -239
rect 65 -251 66 -250
rect 93 -251 94 -250
rect 107 -251 108 -250
rect 121 -251 122 -250
rect 124 -251 125 -250
rect 159 -251 160 -250
rect 177 -251 178 -250
rect 194 -251 195 -250
rect 198 -251 199 -250
rect 261 -251 262 -250
rect 292 -251 293 -250
rect 345 -251 346 -250
rect 366 -251 367 -250
rect 401 -251 402 -250
rect 415 -251 416 -250
rect 492 -251 493 -250
rect 502 -251 503 -250
rect 520 -251 521 -250
rect 590 -251 591 -250
rect 597 -251 598 -250
rect 600 -251 601 -250
rect 611 -251 612 -250
rect 79 -253 80 -252
rect 317 -253 318 -252
rect 320 -253 321 -252
rect 338 -253 339 -252
rect 422 -253 423 -252
rect 457 -253 458 -252
rect 471 -253 472 -252
rect 499 -253 500 -252
rect 506 -253 507 -252
rect 527 -253 528 -252
rect 86 -255 87 -254
rect 128 -255 129 -254
rect 135 -255 136 -254
rect 289 -255 290 -254
rect 303 -255 304 -254
rect 401 -255 402 -254
rect 429 -255 430 -254
rect 478 -255 479 -254
rect 114 -257 115 -256
rect 327 -257 328 -256
rect 338 -257 339 -256
rect 415 -257 416 -256
rect 450 -257 451 -256
rect 485 -257 486 -256
rect 114 -259 115 -258
rect 128 -259 129 -258
rect 135 -259 136 -258
rect 170 -259 171 -258
rect 173 -259 174 -258
rect 177 -259 178 -258
rect 184 -259 185 -258
rect 229 -259 230 -258
rect 254 -259 255 -258
rect 278 -259 279 -258
rect 320 -259 321 -258
rect 408 -259 409 -258
rect 464 -259 465 -258
rect 506 -259 507 -258
rect 142 -261 143 -260
rect 236 -261 237 -260
rect 257 -261 258 -260
rect 324 -261 325 -260
rect 348 -261 349 -260
rect 422 -261 423 -260
rect 436 -261 437 -260
rect 464 -261 465 -260
rect 142 -263 143 -262
rect 184 -263 185 -262
rect 187 -263 188 -262
rect 240 -263 241 -262
rect 324 -263 325 -262
rect 359 -263 360 -262
rect 373 -263 374 -262
rect 429 -263 430 -262
rect 149 -265 150 -264
rect 156 -265 157 -264
rect 163 -265 164 -264
rect 170 -265 171 -264
rect 191 -265 192 -264
rect 243 -265 244 -264
rect 303 -265 304 -264
rect 359 -265 360 -264
rect 380 -265 381 -264
rect 408 -265 409 -264
rect 149 -267 150 -266
rect 205 -267 206 -266
rect 208 -267 209 -266
rect 233 -267 234 -266
rect 236 -267 237 -266
rect 313 -267 314 -266
rect 352 -267 353 -266
rect 373 -267 374 -266
rect 387 -267 388 -266
rect 436 -267 437 -266
rect 156 -269 157 -268
rect 219 -269 220 -268
rect 222 -269 223 -268
rect 310 -269 311 -268
rect 317 -269 318 -268
rect 352 -269 353 -268
rect 394 -269 395 -268
rect 450 -269 451 -268
rect 163 -271 164 -270
rect 243 -271 244 -270
rect 331 -271 332 -270
rect 387 -271 388 -270
rect 201 -273 202 -272
rect 275 -273 276 -272
rect 299 -273 300 -272
rect 331 -273 332 -272
rect 208 -275 209 -274
rect 366 -275 367 -274
rect 219 -277 220 -276
rect 383 -277 384 -276
rect 226 -279 227 -278
rect 282 -279 283 -278
rect 275 -281 276 -280
rect 296 -281 297 -280
rect 75 -292 76 -291
rect 254 -292 255 -291
rect 257 -292 258 -291
rect 317 -292 318 -291
rect 324 -292 325 -291
rect 478 -292 479 -291
rect 516 -292 517 -291
rect 548 -292 549 -291
rect 604 -292 605 -291
rect 611 -292 612 -291
rect 646 -292 647 -291
rect 653 -292 654 -291
rect 674 -292 675 -291
rect 681 -292 682 -291
rect 79 -294 80 -293
rect 212 -294 213 -293
rect 219 -294 220 -293
rect 296 -294 297 -293
rect 303 -294 304 -293
rect 401 -294 402 -293
rect 425 -294 426 -293
rect 457 -294 458 -293
rect 464 -294 465 -293
rect 478 -294 479 -293
rect 520 -294 521 -293
rect 541 -294 542 -293
rect 649 -294 650 -293
rect 660 -294 661 -293
rect 79 -296 80 -295
rect 107 -296 108 -295
rect 114 -296 115 -295
rect 156 -296 157 -295
rect 170 -296 171 -295
rect 177 -296 178 -295
rect 187 -296 188 -295
rect 194 -296 195 -295
rect 205 -296 206 -295
rect 282 -296 283 -295
rect 289 -296 290 -295
rect 471 -296 472 -295
rect 527 -296 528 -295
rect 544 -296 545 -295
rect 86 -298 87 -297
rect 152 -298 153 -297
rect 212 -298 213 -297
rect 233 -298 234 -297
rect 236 -298 237 -297
rect 369 -298 370 -297
rect 390 -298 391 -297
rect 492 -298 493 -297
rect 506 -298 507 -297
rect 527 -298 528 -297
rect 86 -300 87 -299
rect 142 -300 143 -299
rect 219 -300 220 -299
rect 464 -300 465 -299
rect 485 -300 486 -299
rect 506 -300 507 -299
rect 93 -302 94 -301
rect 173 -302 174 -301
rect 247 -302 248 -301
rect 320 -302 321 -301
rect 324 -302 325 -301
rect 429 -302 430 -301
rect 436 -302 437 -301
rect 534 -302 535 -301
rect 93 -304 94 -303
rect 149 -304 150 -303
rect 247 -304 248 -303
rect 345 -304 346 -303
rect 348 -304 349 -303
rect 387 -304 388 -303
rect 394 -304 395 -303
rect 429 -304 430 -303
rect 100 -306 101 -305
rect 117 -306 118 -305
rect 128 -306 129 -305
rect 142 -306 143 -305
rect 254 -306 255 -305
rect 268 -306 269 -305
rect 282 -306 283 -305
rect 485 -306 486 -305
rect 103 -308 104 -307
rect 121 -308 122 -307
rect 135 -308 136 -307
rect 198 -308 199 -307
rect 261 -308 262 -307
rect 264 -308 265 -307
rect 289 -308 290 -307
rect 338 -308 339 -307
rect 341 -308 342 -307
rect 443 -308 444 -307
rect 107 -310 108 -309
rect 163 -310 164 -309
rect 198 -310 199 -309
rect 226 -310 227 -309
rect 303 -310 304 -309
rect 422 -310 423 -309
rect 443 -310 444 -309
rect 555 -310 556 -309
rect 128 -312 129 -311
rect 135 -312 136 -311
rect 163 -312 164 -311
rect 177 -312 178 -311
rect 191 -312 192 -311
rect 226 -312 227 -311
rect 313 -312 314 -311
rect 471 -312 472 -311
rect 345 -314 346 -313
rect 450 -314 451 -313
rect 352 -316 353 -315
rect 401 -316 402 -315
rect 408 -316 409 -315
rect 450 -316 451 -315
rect 331 -318 332 -317
rect 352 -318 353 -317
rect 366 -318 367 -317
rect 380 -318 381 -317
rect 408 -318 409 -317
rect 457 -318 458 -317
rect 331 -320 332 -319
rect 387 -320 388 -319
rect 415 -320 416 -319
rect 492 -320 493 -319
rect 240 -322 241 -321
rect 415 -322 416 -321
rect 422 -322 423 -321
rect 499 -322 500 -321
rect 229 -324 230 -323
rect 240 -324 241 -323
rect 366 -324 367 -323
rect 436 -324 437 -323
rect 373 -326 374 -325
rect 394 -326 395 -325
rect 359 -328 360 -327
rect 373 -328 374 -327
rect 359 -330 360 -329
rect 520 -330 521 -329
rect 44 -341 45 -340
rect 334 -341 335 -340
rect 338 -341 339 -340
rect 527 -341 528 -340
rect 541 -341 542 -340
rect 569 -341 570 -340
rect 583 -341 584 -340
rect 604 -341 605 -340
rect 642 -341 643 -340
rect 688 -341 689 -340
rect 51 -343 52 -342
rect 114 -343 115 -342
rect 128 -343 129 -342
rect 142 -343 143 -342
rect 166 -343 167 -342
rect 236 -343 237 -342
rect 243 -343 244 -342
rect 261 -343 262 -342
rect 264 -343 265 -342
rect 625 -343 626 -342
rect 649 -343 650 -342
rect 653 -343 654 -342
rect 660 -343 661 -342
rect 681 -343 682 -342
rect 58 -345 59 -344
rect 289 -345 290 -344
rect 296 -345 297 -344
rect 313 -345 314 -344
rect 341 -345 342 -344
rect 429 -345 430 -344
rect 471 -345 472 -344
rect 513 -345 514 -344
rect 523 -345 524 -344
rect 597 -345 598 -344
rect 667 -345 668 -344
rect 674 -345 675 -344
rect 79 -347 80 -346
rect 219 -347 220 -346
rect 233 -347 234 -346
rect 345 -347 346 -346
rect 359 -347 360 -346
rect 611 -347 612 -346
rect 79 -349 80 -348
rect 170 -349 171 -348
rect 177 -349 178 -348
rect 226 -349 227 -348
rect 233 -349 234 -348
rect 352 -349 353 -348
rect 362 -349 363 -348
rect 534 -349 535 -348
rect 544 -349 545 -348
rect 639 -349 640 -348
rect 86 -351 87 -350
rect 163 -351 164 -350
rect 177 -351 178 -350
rect 215 -351 216 -350
rect 222 -351 223 -350
rect 362 -351 363 -350
rect 366 -351 367 -350
rect 618 -351 619 -350
rect 86 -353 87 -352
rect 247 -353 248 -352
rect 254 -353 255 -352
rect 268 -353 269 -352
rect 275 -353 276 -352
rect 296 -353 297 -352
rect 341 -353 342 -352
rect 527 -353 528 -352
rect 548 -353 549 -352
rect 646 -353 647 -352
rect 93 -355 94 -354
rect 156 -355 157 -354
rect 159 -355 160 -354
rect 254 -355 255 -354
rect 292 -355 293 -354
rect 366 -355 367 -354
rect 380 -355 381 -354
rect 390 -355 391 -354
rect 411 -355 412 -354
rect 436 -355 437 -354
rect 460 -355 461 -354
rect 534 -355 535 -354
rect 558 -355 559 -354
rect 562 -355 563 -354
rect 72 -357 73 -356
rect 156 -357 157 -356
rect 205 -357 206 -356
rect 285 -357 286 -356
rect 327 -357 328 -356
rect 548 -357 549 -356
rect 562 -357 563 -356
rect 653 -357 654 -356
rect 72 -359 73 -358
rect 212 -359 213 -358
rect 236 -359 237 -358
rect 271 -359 272 -358
rect 327 -359 328 -358
rect 408 -359 409 -358
rect 415 -359 416 -358
rect 436 -359 437 -358
rect 471 -359 472 -358
rect 660 -359 661 -358
rect 93 -361 94 -360
rect 100 -361 101 -360
rect 114 -361 115 -360
rect 401 -361 402 -360
rect 415 -361 416 -360
rect 425 -361 426 -360
rect 478 -361 479 -360
rect 541 -361 542 -360
rect 100 -363 101 -362
rect 121 -363 122 -362
rect 128 -363 129 -362
rect 135 -363 136 -362
rect 142 -363 143 -362
rect 229 -363 230 -362
rect 373 -363 374 -362
rect 478 -363 479 -362
rect 485 -363 486 -362
rect 590 -363 591 -362
rect 68 -365 69 -364
rect 135 -365 136 -364
rect 152 -365 153 -364
rect 219 -365 220 -364
rect 380 -365 381 -364
rect 387 -365 388 -364
rect 394 -365 395 -364
rect 401 -365 402 -364
rect 422 -365 423 -364
rect 576 -365 577 -364
rect 107 -367 108 -366
rect 152 -367 153 -366
rect 205 -367 206 -366
rect 240 -367 241 -366
rect 317 -367 318 -366
rect 394 -367 395 -366
rect 422 -367 423 -366
rect 520 -367 521 -366
rect 107 -369 108 -368
rect 247 -369 248 -368
rect 317 -369 318 -368
rect 457 -369 458 -368
rect 492 -369 493 -368
rect 604 -369 605 -368
rect 110 -371 111 -370
rect 373 -371 374 -370
rect 443 -371 444 -370
rect 485 -371 486 -370
rect 499 -371 500 -370
rect 555 -371 556 -370
rect 121 -373 122 -372
rect 191 -373 192 -372
rect 303 -373 304 -372
rect 443 -373 444 -372
rect 450 -373 451 -372
rect 492 -373 493 -372
rect 506 -373 507 -372
rect 632 -373 633 -372
rect 170 -375 171 -374
rect 240 -375 241 -374
rect 303 -375 304 -374
rect 324 -375 325 -374
rect 348 -375 349 -374
rect 499 -375 500 -374
rect 184 -377 185 -376
rect 191 -377 192 -376
rect 310 -377 311 -376
rect 324 -377 325 -376
rect 429 -377 430 -376
rect 450 -377 451 -376
rect 464 -377 465 -376
rect 506 -377 507 -376
rect 184 -379 185 -378
rect 198 -379 199 -378
rect 331 -379 332 -378
rect 464 -379 465 -378
rect 138 -381 139 -380
rect 198 -381 199 -380
rect 282 -381 283 -380
rect 331 -381 332 -380
rect 2 -392 3 -391
rect 180 -392 181 -391
rect 205 -392 206 -391
rect 226 -392 227 -391
rect 233 -392 234 -391
rect 310 -392 311 -391
rect 317 -392 318 -391
rect 352 -392 353 -391
rect 359 -392 360 -391
rect 611 -392 612 -391
rect 628 -392 629 -391
rect 639 -392 640 -391
rect 649 -392 650 -391
rect 681 -392 682 -391
rect 16 -394 17 -393
rect 292 -394 293 -393
rect 303 -394 304 -393
rect 352 -394 353 -393
rect 355 -394 356 -393
rect 359 -394 360 -393
rect 373 -394 374 -393
rect 562 -394 563 -393
rect 597 -394 598 -393
rect 611 -394 612 -393
rect 667 -394 668 -393
rect 674 -394 675 -393
rect 30 -396 31 -395
rect 37 -396 38 -395
rect 44 -396 45 -395
rect 222 -396 223 -395
rect 240 -396 241 -395
rect 464 -396 465 -395
rect 597 -396 598 -395
rect 625 -396 626 -395
rect 667 -396 668 -395
rect 688 -396 689 -395
rect 44 -398 45 -397
rect 397 -398 398 -397
rect 401 -398 402 -397
rect 422 -398 423 -397
rect 436 -398 437 -397
rect 446 -398 447 -397
rect 450 -398 451 -397
rect 646 -398 647 -397
rect 51 -400 52 -399
rect 138 -400 139 -399
rect 149 -400 150 -399
rect 191 -400 192 -399
rect 215 -400 216 -399
rect 394 -400 395 -399
rect 401 -400 402 -399
rect 632 -400 633 -399
rect 51 -402 52 -401
rect 152 -402 153 -401
rect 163 -402 164 -401
rect 184 -402 185 -401
rect 219 -402 220 -401
rect 404 -402 405 -401
rect 436 -402 437 -401
rect 534 -402 535 -401
rect 576 -402 577 -401
rect 632 -402 633 -401
rect 58 -404 59 -403
rect 341 -404 342 -403
rect 373 -404 374 -403
rect 450 -404 451 -403
rect 460 -404 461 -403
rect 548 -404 549 -403
rect 558 -404 559 -403
rect 576 -404 577 -403
rect 583 -404 584 -403
rect 625 -404 626 -403
rect 58 -406 59 -405
rect 212 -406 213 -405
rect 268 -406 269 -405
rect 289 -406 290 -405
rect 317 -406 318 -405
rect 366 -406 367 -405
rect 376 -406 377 -405
rect 415 -406 416 -405
rect 439 -406 440 -405
rect 604 -406 605 -405
rect 65 -408 66 -407
rect 303 -408 304 -407
rect 334 -408 335 -407
rect 590 -408 591 -407
rect 604 -408 605 -407
rect 653 -408 654 -407
rect 72 -410 73 -409
rect 327 -410 328 -409
rect 341 -410 342 -409
rect 478 -410 479 -409
rect 492 -410 493 -409
rect 534 -410 535 -409
rect 569 -410 570 -409
rect 583 -410 584 -409
rect 653 -410 654 -409
rect 663 -410 664 -409
rect 72 -412 73 -411
rect 187 -412 188 -411
rect 254 -412 255 -411
rect 268 -412 269 -411
rect 285 -412 286 -411
rect 296 -412 297 -411
rect 369 -412 370 -411
rect 478 -412 479 -411
rect 541 -412 542 -411
rect 569 -412 570 -411
rect 79 -414 80 -413
rect 240 -414 241 -413
rect 247 -414 248 -413
rect 296 -414 297 -413
rect 387 -414 388 -413
rect 618 -414 619 -413
rect 79 -416 80 -415
rect 215 -416 216 -415
rect 247 -416 248 -415
rect 261 -416 262 -415
rect 289 -416 290 -415
rect 331 -416 332 -415
rect 387 -416 388 -415
rect 443 -416 444 -415
rect 467 -416 468 -415
rect 590 -416 591 -415
rect 86 -418 87 -417
rect 324 -418 325 -417
rect 345 -418 346 -417
rect 443 -418 444 -417
rect 471 -418 472 -417
rect 492 -418 493 -417
rect 499 -418 500 -417
rect 541 -418 542 -417
rect 555 -418 556 -417
rect 618 -418 619 -417
rect 100 -420 101 -419
rect 159 -420 160 -419
rect 184 -420 185 -419
rect 191 -420 192 -419
rect 236 -420 237 -419
rect 345 -420 346 -419
rect 408 -420 409 -419
rect 499 -420 500 -419
rect 100 -422 101 -421
rect 145 -422 146 -421
rect 159 -422 160 -421
rect 520 -422 521 -421
rect 107 -424 108 -423
rect 198 -424 199 -423
rect 236 -424 237 -423
rect 278 -424 279 -423
rect 324 -424 325 -423
rect 506 -424 507 -423
rect 114 -426 115 -425
rect 275 -426 276 -425
rect 408 -426 409 -425
rect 457 -426 458 -425
rect 114 -428 115 -427
rect 128 -428 129 -427
rect 135 -428 136 -427
rect 166 -428 167 -427
rect 198 -428 199 -427
rect 548 -428 549 -427
rect 121 -430 122 -429
rect 310 -430 311 -429
rect 415 -430 416 -429
rect 429 -430 430 -429
rect 446 -430 447 -429
rect 471 -430 472 -429
rect 86 -432 87 -431
rect 121 -432 122 -431
rect 128 -432 129 -431
rect 170 -432 171 -431
rect 261 -432 262 -431
rect 282 -432 283 -431
rect 338 -432 339 -431
rect 429 -432 430 -431
rect 142 -434 143 -433
rect 254 -434 255 -433
rect 170 -436 171 -435
rect 177 -436 178 -435
rect 205 -436 206 -435
rect 282 -436 283 -435
rect 23 -438 24 -437
rect 177 -438 178 -437
rect 9 -449 10 -448
rect 110 -449 111 -448
rect 131 -449 132 -448
rect 520 -449 521 -448
rect 541 -449 542 -448
rect 555 -449 556 -448
rect 558 -449 559 -448
rect 583 -449 584 -448
rect 611 -449 612 -448
rect 614 -449 615 -448
rect 635 -449 636 -448
rect 653 -449 654 -448
rect 660 -449 661 -448
rect 667 -449 668 -448
rect 9 -451 10 -450
rect 355 -451 356 -450
rect 369 -451 370 -450
rect 534 -451 535 -450
rect 583 -451 584 -450
rect 604 -451 605 -450
rect 653 -451 654 -450
rect 663 -451 664 -450
rect 16 -453 17 -452
rect 236 -453 237 -452
rect 247 -453 248 -452
rect 285 -453 286 -452
rect 292 -453 293 -452
rect 415 -453 416 -452
rect 418 -453 419 -452
rect 534 -453 535 -452
rect 16 -455 17 -454
rect 114 -455 115 -454
rect 142 -455 143 -454
rect 170 -455 171 -454
rect 208 -455 209 -454
rect 331 -455 332 -454
rect 373 -455 374 -454
rect 499 -455 500 -454
rect 520 -455 521 -454
rect 562 -455 563 -454
rect 23 -457 24 -456
rect 180 -457 181 -456
rect 215 -457 216 -456
rect 261 -457 262 -456
rect 275 -457 276 -456
rect 338 -457 339 -456
rect 376 -457 377 -456
rect 513 -457 514 -456
rect 23 -459 24 -458
rect 86 -459 87 -458
rect 107 -459 108 -458
rect 170 -459 171 -458
rect 177 -459 178 -458
rect 373 -459 374 -458
rect 397 -459 398 -458
rect 492 -459 493 -458
rect 499 -459 500 -458
rect 509 -459 510 -458
rect 513 -459 514 -458
rect 527 -459 528 -458
rect 30 -461 31 -460
rect 138 -461 139 -460
rect 142 -461 143 -460
rect 296 -461 297 -460
rect 324 -461 325 -460
rect 415 -461 416 -460
rect 436 -461 437 -460
rect 541 -461 542 -460
rect 33 -463 34 -462
rect 37 -463 38 -462
rect 44 -463 45 -462
rect 156 -463 157 -462
rect 159 -463 160 -462
rect 359 -463 360 -462
rect 408 -463 409 -462
rect 422 -463 423 -462
rect 436 -463 437 -462
rect 618 -463 619 -462
rect 37 -465 38 -464
rect 107 -465 108 -464
rect 121 -465 122 -464
rect 138 -465 139 -464
rect 163 -465 164 -464
rect 187 -465 188 -464
rect 233 -465 234 -464
rect 303 -465 304 -464
rect 359 -465 360 -464
rect 387 -465 388 -464
rect 457 -465 458 -464
rect 509 -465 510 -464
rect 576 -465 577 -464
rect 618 -465 619 -464
rect 44 -467 45 -466
rect 149 -467 150 -466
rect 163 -467 164 -466
rect 345 -467 346 -466
rect 387 -467 388 -466
rect 471 -467 472 -466
rect 478 -467 479 -466
rect 562 -467 563 -466
rect 576 -467 577 -466
rect 597 -467 598 -466
rect 51 -469 52 -468
rect 184 -469 185 -468
rect 219 -469 220 -468
rect 233 -469 234 -468
rect 243 -469 244 -468
rect 492 -469 493 -468
rect 597 -469 598 -468
rect 625 -469 626 -468
rect 2 -471 3 -470
rect 243 -471 244 -470
rect 247 -471 248 -470
rect 464 -471 465 -470
rect 485 -471 486 -470
rect 527 -471 528 -470
rect 51 -473 52 -472
rect 100 -473 101 -472
rect 121 -473 122 -472
rect 264 -473 265 -472
rect 275 -473 276 -472
rect 352 -473 353 -472
rect 397 -473 398 -472
rect 485 -473 486 -472
rect 58 -475 59 -474
rect 145 -475 146 -474
rect 166 -475 167 -474
rect 184 -475 185 -474
rect 205 -475 206 -474
rect 219 -475 220 -474
rect 254 -475 255 -474
rect 289 -475 290 -474
rect 296 -475 297 -474
rect 632 -475 633 -474
rect 58 -477 59 -476
rect 401 -477 402 -476
rect 429 -477 430 -476
rect 457 -477 458 -476
rect 632 -477 633 -476
rect 639 -477 640 -476
rect 65 -479 66 -478
rect 366 -479 367 -478
rect 429 -479 430 -478
rect 443 -479 444 -478
rect 450 -479 451 -478
rect 471 -479 472 -478
rect 590 -479 591 -478
rect 639 -479 640 -478
rect 65 -481 66 -480
rect 548 -481 549 -480
rect 72 -483 73 -482
rect 201 -483 202 -482
rect 212 -483 213 -482
rect 254 -483 255 -482
rect 268 -483 269 -482
rect 289 -483 290 -482
rect 345 -483 346 -482
rect 404 -483 405 -482
rect 548 -483 549 -482
rect 569 -483 570 -482
rect 72 -485 73 -484
rect 128 -485 129 -484
rect 177 -485 178 -484
rect 191 -485 192 -484
rect 215 -485 216 -484
rect 366 -485 367 -484
rect 390 -485 391 -484
rect 443 -485 444 -484
rect 79 -487 80 -486
rect 422 -487 423 -486
rect 79 -489 80 -488
rect 93 -489 94 -488
rect 100 -489 101 -488
rect 198 -489 199 -488
rect 282 -489 283 -488
rect 464 -489 465 -488
rect 86 -491 87 -490
rect 114 -491 115 -490
rect 128 -491 129 -490
rect 191 -491 192 -490
rect 282 -491 283 -490
rect 310 -491 311 -490
rect 352 -491 353 -490
rect 450 -491 451 -490
rect 310 -493 311 -492
rect 380 -493 381 -492
rect 380 -495 381 -494
rect 569 -495 570 -494
rect 5 -506 6 -505
rect 163 -506 164 -505
rect 198 -506 199 -505
rect 362 -506 363 -505
rect 366 -506 367 -505
rect 611 -506 612 -505
rect 618 -506 619 -505
rect 628 -506 629 -505
rect 653 -506 654 -505
rect 670 -506 671 -505
rect 681 -506 682 -505
rect 688 -506 689 -505
rect 9 -508 10 -507
rect 117 -508 118 -507
rect 121 -508 122 -507
rect 124 -508 125 -507
rect 152 -508 153 -507
rect 275 -508 276 -507
rect 285 -508 286 -507
rect 569 -508 570 -507
rect 583 -508 584 -507
rect 611 -508 612 -507
rect 628 -508 629 -507
rect 646 -508 647 -507
rect 667 -508 668 -507
rect 674 -508 675 -507
rect 9 -510 10 -509
rect 61 -510 62 -509
rect 65 -510 66 -509
rect 86 -510 87 -509
rect 93 -510 94 -509
rect 100 -510 101 -509
rect 121 -510 122 -509
rect 247 -510 248 -509
rect 268 -510 269 -509
rect 296 -510 297 -509
rect 310 -510 311 -509
rect 376 -510 377 -509
rect 383 -510 384 -509
rect 492 -510 493 -509
rect 499 -510 500 -509
rect 590 -510 591 -509
rect 604 -510 605 -509
rect 614 -510 615 -509
rect 618 -510 619 -509
rect 646 -510 647 -509
rect 23 -512 24 -511
rect 58 -512 59 -511
rect 68 -512 69 -511
rect 212 -512 213 -511
rect 219 -512 220 -511
rect 275 -512 276 -511
rect 289 -512 290 -511
rect 310 -512 311 -511
rect 338 -512 339 -511
rect 348 -512 349 -511
rect 369 -512 370 -511
rect 604 -512 605 -511
rect 639 -512 640 -511
rect 653 -512 654 -511
rect 23 -514 24 -513
rect 240 -514 241 -513
rect 243 -514 244 -513
rect 562 -514 563 -513
rect 576 -514 577 -513
rect 590 -514 591 -513
rect 30 -516 31 -515
rect 208 -516 209 -515
rect 212 -516 213 -515
rect 226 -516 227 -515
rect 243 -516 244 -515
rect 387 -516 388 -515
rect 390 -516 391 -515
rect 541 -516 542 -515
rect 555 -516 556 -515
rect 562 -516 563 -515
rect 30 -518 31 -517
rect 180 -518 181 -517
rect 278 -518 279 -517
rect 555 -518 556 -517
rect 37 -520 38 -519
rect 156 -520 157 -519
rect 163 -520 164 -519
rect 436 -520 437 -519
rect 450 -520 451 -519
rect 492 -520 493 -519
rect 502 -520 503 -519
rect 513 -520 514 -519
rect 37 -522 38 -521
rect 142 -522 143 -521
rect 149 -522 150 -521
rect 219 -522 220 -521
rect 292 -522 293 -521
rect 436 -522 437 -521
rect 478 -522 479 -521
rect 569 -522 570 -521
rect 16 -524 17 -523
rect 149 -524 150 -523
rect 156 -524 157 -523
rect 233 -524 234 -523
rect 296 -524 297 -523
rect 303 -524 304 -523
rect 331 -524 332 -523
rect 541 -524 542 -523
rect 16 -526 17 -525
rect 82 -526 83 -525
rect 86 -526 87 -525
rect 100 -526 101 -525
rect 114 -526 115 -525
rect 576 -526 577 -525
rect 44 -528 45 -527
rect 215 -528 216 -527
rect 303 -528 304 -527
rect 324 -528 325 -527
rect 341 -528 342 -527
rect 450 -528 451 -527
rect 457 -528 458 -527
rect 478 -528 479 -527
rect 485 -528 486 -527
rect 583 -528 584 -527
rect 44 -530 45 -529
rect 240 -530 241 -529
rect 324 -530 325 -529
rect 345 -530 346 -529
rect 373 -530 374 -529
rect 394 -530 395 -529
rect 397 -530 398 -529
rect 597 -530 598 -529
rect 72 -532 73 -531
rect 135 -532 136 -531
rect 170 -532 171 -531
rect 226 -532 227 -531
rect 345 -532 346 -531
rect 380 -532 381 -531
rect 415 -532 416 -531
rect 527 -532 528 -531
rect 548 -532 549 -531
rect 597 -532 598 -531
rect 51 -534 52 -533
rect 72 -534 73 -533
rect 93 -534 94 -533
rect 191 -534 192 -533
rect 205 -534 206 -533
rect 233 -534 234 -533
rect 359 -534 360 -533
rect 394 -534 395 -533
rect 415 -534 416 -533
rect 429 -534 430 -533
rect 471 -534 472 -533
rect 485 -534 486 -533
rect 499 -534 500 -533
rect 527 -534 528 -533
rect 534 -534 535 -533
rect 548 -534 549 -533
rect 51 -536 52 -535
rect 79 -536 80 -535
rect 107 -536 108 -535
rect 135 -536 136 -535
rect 170 -536 171 -535
rect 282 -536 283 -535
rect 401 -536 402 -535
rect 471 -536 472 -535
rect 506 -536 507 -535
rect 520 -536 521 -535
rect 107 -538 108 -537
rect 184 -538 185 -537
rect 208 -538 209 -537
rect 429 -538 430 -537
rect 464 -538 465 -537
rect 534 -538 535 -537
rect 124 -540 125 -539
rect 247 -540 248 -539
rect 261 -540 262 -539
rect 401 -540 402 -539
rect 422 -540 423 -539
rect 639 -540 640 -539
rect 128 -542 129 -541
rect 331 -542 332 -541
rect 355 -542 356 -541
rect 464 -542 465 -541
rect 513 -542 514 -541
rect 625 -542 626 -541
rect 131 -544 132 -543
rect 205 -544 206 -543
rect 313 -544 314 -543
rect 520 -544 521 -543
rect 159 -546 160 -545
rect 184 -546 185 -545
rect 355 -546 356 -545
rect 408 -546 409 -545
rect 177 -548 178 -547
rect 198 -548 199 -547
rect 408 -548 409 -547
rect 443 -548 444 -547
rect 317 -550 318 -549
rect 443 -550 444 -549
rect 271 -552 272 -551
rect 317 -552 318 -551
rect 2 -563 3 -562
rect 268 -563 269 -562
rect 275 -563 276 -562
rect 320 -563 321 -562
rect 345 -563 346 -562
rect 422 -563 423 -562
rect 436 -563 437 -562
rect 618 -563 619 -562
rect 646 -563 647 -562
rect 667 -563 668 -562
rect 670 -563 671 -562
rect 684 -563 685 -562
rect 19 -565 20 -564
rect 306 -565 307 -564
rect 310 -565 311 -564
rect 394 -565 395 -564
rect 401 -565 402 -564
rect 632 -565 633 -564
rect 653 -565 654 -564
rect 656 -565 657 -564
rect 674 -565 675 -564
rect 677 -565 678 -564
rect 23 -567 24 -566
rect 96 -567 97 -566
rect 107 -567 108 -566
rect 292 -567 293 -566
rect 296 -567 297 -566
rect 369 -567 370 -566
rect 380 -567 381 -566
rect 401 -567 402 -566
rect 404 -567 405 -566
rect 597 -567 598 -566
rect 618 -567 619 -566
rect 625 -567 626 -566
rect 653 -567 654 -566
rect 660 -567 661 -566
rect 23 -569 24 -568
rect 121 -569 122 -568
rect 128 -569 129 -568
rect 219 -569 220 -568
rect 233 -569 234 -568
rect 268 -569 269 -568
rect 278 -569 279 -568
rect 541 -569 542 -568
rect 590 -569 591 -568
rect 646 -569 647 -568
rect 9 -571 10 -570
rect 128 -571 129 -570
rect 131 -571 132 -570
rect 604 -571 605 -570
rect 9 -573 10 -572
rect 177 -573 178 -572
rect 180 -573 181 -572
rect 471 -573 472 -572
rect 478 -573 479 -572
rect 590 -573 591 -572
rect 604 -573 605 -572
rect 625 -573 626 -572
rect 30 -575 31 -574
rect 100 -575 101 -574
rect 107 -575 108 -574
rect 170 -575 171 -574
rect 243 -575 244 -574
rect 639 -575 640 -574
rect 30 -577 31 -576
rect 233 -577 234 -576
rect 247 -577 248 -576
rect 380 -577 381 -576
rect 383 -577 384 -576
rect 478 -577 479 -576
rect 499 -577 500 -576
rect 513 -577 514 -576
rect 534 -577 535 -576
rect 541 -577 542 -576
rect 562 -577 563 -576
rect 639 -577 640 -576
rect 37 -579 38 -578
rect 341 -579 342 -578
rect 345 -579 346 -578
rect 352 -579 353 -578
rect 355 -579 356 -578
rect 443 -579 444 -578
rect 457 -579 458 -578
rect 492 -579 493 -578
rect 40 -581 41 -580
rect 180 -581 181 -580
rect 184 -581 185 -580
rect 247 -581 248 -580
rect 254 -581 255 -580
rect 474 -581 475 -580
rect 485 -581 486 -580
rect 513 -581 514 -580
rect 44 -583 45 -582
rect 142 -583 143 -582
rect 163 -583 164 -582
rect 219 -583 220 -582
rect 285 -583 286 -582
rect 338 -583 339 -582
rect 366 -583 367 -582
rect 376 -583 377 -582
rect 387 -583 388 -582
rect 597 -583 598 -582
rect 51 -585 52 -584
rect 54 -585 55 -584
rect 65 -585 66 -584
rect 82 -585 83 -584
rect 93 -585 94 -584
rect 296 -585 297 -584
rect 317 -585 318 -584
rect 569 -585 570 -584
rect 16 -587 17 -586
rect 93 -587 94 -586
rect 100 -587 101 -586
rect 117 -587 118 -586
rect 121 -587 122 -586
rect 177 -587 178 -586
rect 212 -587 213 -586
rect 254 -587 255 -586
rect 289 -587 290 -586
rect 534 -587 535 -586
rect 548 -587 549 -586
rect 569 -587 570 -586
rect 51 -589 52 -588
rect 86 -589 87 -588
rect 114 -589 115 -588
rect 156 -589 157 -588
rect 163 -589 164 -588
rect 226 -589 227 -588
rect 236 -589 237 -588
rect 317 -589 318 -588
rect 366 -589 367 -588
rect 632 -589 633 -588
rect 58 -591 59 -590
rect 114 -591 115 -590
rect 131 -591 132 -590
rect 282 -591 283 -590
rect 289 -591 290 -590
rect 467 -591 468 -590
rect 471 -591 472 -590
rect 611 -591 612 -590
rect 656 -591 657 -590
rect 660 -591 661 -590
rect 65 -593 66 -592
rect 103 -593 104 -592
rect 135 -593 136 -592
rect 194 -593 195 -592
rect 198 -593 199 -592
rect 226 -593 227 -592
rect 282 -593 283 -592
rect 303 -593 304 -592
rect 373 -593 374 -592
rect 443 -593 444 -592
rect 485 -593 486 -592
rect 520 -593 521 -592
rect 583 -593 584 -592
rect 611 -593 612 -592
rect 75 -595 76 -594
rect 310 -595 311 -594
rect 359 -595 360 -594
rect 583 -595 584 -594
rect 79 -597 80 -596
rect 184 -597 185 -596
rect 198 -597 199 -596
rect 243 -597 244 -596
rect 303 -597 304 -596
rect 555 -597 556 -596
rect 135 -599 136 -598
rect 261 -599 262 -598
rect 359 -599 360 -598
rect 425 -599 426 -598
rect 429 -599 430 -598
rect 457 -599 458 -598
rect 460 -599 461 -598
rect 520 -599 521 -598
rect 527 -599 528 -598
rect 555 -599 556 -598
rect 142 -601 143 -600
rect 187 -601 188 -600
rect 205 -601 206 -600
rect 429 -601 430 -600
rect 450 -601 451 -600
rect 527 -601 528 -600
rect 170 -603 171 -602
rect 191 -603 192 -602
rect 205 -603 206 -602
rect 313 -603 314 -602
rect 373 -603 374 -602
rect 397 -603 398 -602
rect 450 -603 451 -602
rect 464 -603 465 -602
rect 506 -603 507 -602
rect 548 -603 549 -602
rect 212 -605 213 -604
rect 264 -605 265 -604
rect 331 -605 332 -604
rect 506 -605 507 -604
rect 324 -607 325 -606
rect 331 -607 332 -606
rect 387 -607 388 -606
rect 436 -607 437 -606
rect 464 -607 465 -606
rect 562 -607 563 -606
rect 72 -609 73 -608
rect 324 -609 325 -608
rect 2 -620 3 -619
rect 394 -620 395 -619
rect 411 -620 412 -619
rect 590 -620 591 -619
rect 632 -620 633 -619
rect 702 -620 703 -619
rect 716 -620 717 -619
rect 730 -620 731 -619
rect 2 -622 3 -621
rect 44 -622 45 -621
rect 51 -622 52 -621
rect 114 -622 115 -621
rect 159 -622 160 -621
rect 247 -622 248 -621
rect 285 -622 286 -621
rect 471 -622 472 -621
rect 492 -622 493 -621
rect 639 -622 640 -621
rect 653 -622 654 -621
rect 660 -622 661 -621
rect 681 -622 682 -621
rect 688 -622 689 -621
rect 695 -622 696 -621
rect 719 -622 720 -621
rect 9 -624 10 -623
rect 187 -624 188 -623
rect 194 -624 195 -623
rect 289 -624 290 -623
rect 296 -624 297 -623
rect 348 -624 349 -623
rect 355 -624 356 -623
rect 359 -624 360 -623
rect 376 -624 377 -623
rect 520 -624 521 -623
rect 527 -624 528 -623
rect 604 -624 605 -623
rect 618 -624 619 -623
rect 660 -624 661 -623
rect 9 -626 10 -625
rect 86 -626 87 -625
rect 93 -626 94 -625
rect 100 -626 101 -625
rect 107 -626 108 -625
rect 352 -626 353 -625
rect 380 -626 381 -625
rect 653 -626 654 -625
rect 23 -628 24 -627
rect 96 -628 97 -627
rect 107 -628 108 -627
rect 149 -628 150 -627
rect 166 -628 167 -627
rect 170 -628 171 -627
rect 177 -628 178 -627
rect 387 -628 388 -627
rect 390 -628 391 -627
rect 576 -628 577 -627
rect 583 -628 584 -627
rect 618 -628 619 -627
rect 23 -630 24 -629
rect 173 -630 174 -629
rect 177 -630 178 -629
rect 212 -630 213 -629
rect 226 -630 227 -629
rect 261 -630 262 -629
rect 289 -630 290 -629
rect 373 -630 374 -629
rect 383 -630 384 -629
rect 569 -630 570 -629
rect 30 -632 31 -631
rect 369 -632 370 -631
rect 394 -632 395 -631
rect 408 -632 409 -631
rect 425 -632 426 -631
rect 548 -632 549 -631
rect 562 -632 563 -631
rect 590 -632 591 -631
rect 30 -634 31 -633
rect 163 -634 164 -633
rect 184 -634 185 -633
rect 278 -634 279 -633
rect 345 -634 346 -633
rect 380 -634 381 -633
rect 453 -634 454 -633
rect 667 -634 668 -633
rect 16 -636 17 -635
rect 278 -636 279 -635
rect 345 -636 346 -635
rect 492 -636 493 -635
rect 495 -636 496 -635
rect 548 -636 549 -635
rect 37 -638 38 -637
rect 61 -638 62 -637
rect 72 -638 73 -637
rect 121 -638 122 -637
rect 128 -638 129 -637
rect 163 -638 164 -637
rect 212 -638 213 -637
rect 219 -638 220 -637
rect 240 -638 241 -637
rect 254 -638 255 -637
rect 366 -638 367 -637
rect 569 -638 570 -637
rect 44 -640 45 -639
rect 89 -640 90 -639
rect 93 -640 94 -639
rect 520 -640 521 -639
rect 541 -640 542 -639
rect 562 -640 563 -639
rect 54 -642 55 -641
rect 254 -642 255 -641
rect 303 -642 304 -641
rect 366 -642 367 -641
rect 369 -642 370 -641
rect 555 -642 556 -641
rect 58 -644 59 -643
rect 75 -644 76 -643
rect 114 -644 115 -643
rect 156 -644 157 -643
rect 240 -644 241 -643
rect 268 -644 269 -643
rect 324 -644 325 -643
rect 555 -644 556 -643
rect 117 -646 118 -645
rect 166 -646 167 -645
rect 229 -646 230 -645
rect 268 -646 269 -645
rect 324 -646 325 -645
rect 401 -646 402 -645
rect 453 -646 454 -645
rect 632 -646 633 -645
rect 121 -648 122 -647
rect 145 -648 146 -647
rect 149 -648 150 -647
rect 205 -648 206 -647
rect 243 -648 244 -647
rect 282 -648 283 -647
rect 310 -648 311 -647
rect 401 -648 402 -647
rect 464 -648 465 -647
rect 611 -648 612 -647
rect 79 -650 80 -649
rect 310 -650 311 -649
rect 387 -650 388 -649
rect 464 -650 465 -649
rect 474 -650 475 -649
rect 639 -650 640 -649
rect 79 -652 80 -651
rect 128 -652 129 -651
rect 135 -652 136 -651
rect 219 -652 220 -651
rect 282 -652 283 -651
rect 583 -652 584 -651
rect 142 -654 143 -653
rect 247 -654 248 -653
rect 506 -654 507 -653
rect 527 -654 528 -653
rect 534 -654 535 -653
rect 611 -654 612 -653
rect 142 -656 143 -655
rect 485 -656 486 -655
rect 499 -656 500 -655
rect 534 -656 535 -655
rect 156 -658 157 -657
rect 233 -658 234 -657
rect 243 -658 244 -657
rect 506 -658 507 -657
rect 513 -658 514 -657
rect 541 -658 542 -657
rect 198 -660 199 -659
rect 205 -660 206 -659
rect 338 -660 339 -659
rect 485 -660 486 -659
rect 135 -662 136 -661
rect 198 -662 199 -661
rect 457 -662 458 -661
rect 499 -662 500 -661
rect 191 -664 192 -663
rect 338 -664 339 -663
rect 457 -664 458 -663
rect 646 -664 647 -663
rect 191 -666 192 -665
rect 677 -666 678 -665
rect 478 -668 479 -667
rect 513 -668 514 -667
rect 625 -668 626 -667
rect 646 -668 647 -667
rect 443 -670 444 -669
rect 478 -670 479 -669
rect 597 -670 598 -669
rect 625 -670 626 -669
rect 299 -672 300 -671
rect 597 -672 598 -671
rect 429 -674 430 -673
rect 443 -674 444 -673
rect 415 -676 416 -675
rect 429 -676 430 -675
rect 415 -678 416 -677
rect 436 -678 437 -677
rect 422 -680 423 -679
rect 436 -680 437 -679
rect 422 -682 423 -681
rect 576 -682 577 -681
rect 2 -693 3 -692
rect 79 -693 80 -692
rect 82 -693 83 -692
rect 436 -693 437 -692
rect 450 -693 451 -692
rect 541 -693 542 -692
rect 632 -693 633 -692
rect 723 -693 724 -692
rect 730 -693 731 -692
rect 754 -693 755 -692
rect 800 -693 801 -692
rect 807 -693 808 -692
rect 9 -695 10 -694
rect 138 -695 139 -694
rect 215 -695 216 -694
rect 310 -695 311 -694
rect 341 -695 342 -694
rect 471 -695 472 -694
rect 534 -695 535 -694
rect 716 -695 717 -694
rect 16 -697 17 -696
rect 324 -697 325 -696
rect 345 -697 346 -696
rect 527 -697 528 -696
rect 674 -697 675 -696
rect 695 -697 696 -696
rect 702 -697 703 -696
rect 744 -697 745 -696
rect 19 -699 20 -698
rect 103 -699 104 -698
rect 121 -699 122 -698
rect 163 -699 164 -698
rect 226 -699 227 -698
rect 261 -699 262 -698
rect 278 -699 279 -698
rect 583 -699 584 -698
rect 653 -699 654 -698
rect 695 -699 696 -698
rect 9 -701 10 -700
rect 226 -701 227 -700
rect 236 -701 237 -700
rect 460 -701 461 -700
rect 464 -701 465 -700
rect 611 -701 612 -700
rect 646 -701 647 -700
rect 653 -701 654 -700
rect 23 -703 24 -702
rect 187 -703 188 -702
rect 254 -703 255 -702
rect 411 -703 412 -702
rect 422 -703 423 -702
rect 688 -703 689 -702
rect 23 -705 24 -704
rect 166 -705 167 -704
rect 201 -705 202 -704
rect 422 -705 423 -704
rect 429 -705 430 -704
rect 464 -705 465 -704
rect 499 -705 500 -704
rect 534 -705 535 -704
rect 569 -705 570 -704
rect 688 -705 689 -704
rect 30 -707 31 -706
rect 240 -707 241 -706
rect 254 -707 255 -706
rect 289 -707 290 -706
rect 296 -707 297 -706
rect 401 -707 402 -706
rect 408 -707 409 -706
rect 632 -707 633 -706
rect 30 -709 31 -708
rect 93 -709 94 -708
rect 100 -709 101 -708
rect 387 -709 388 -708
rect 401 -709 402 -708
rect 457 -709 458 -708
rect 467 -709 468 -708
rect 569 -709 570 -708
rect 576 -709 577 -708
rect 611 -709 612 -708
rect 37 -711 38 -710
rect 89 -711 90 -710
rect 93 -711 94 -710
rect 156 -711 157 -710
rect 240 -711 241 -710
rect 429 -711 430 -710
rect 432 -711 433 -710
rect 625 -711 626 -710
rect 2 -713 3 -712
rect 89 -713 90 -712
rect 100 -713 101 -712
rect 737 -713 738 -712
rect 40 -715 41 -714
rect 303 -715 304 -714
rect 310 -715 311 -714
rect 331 -715 332 -714
rect 352 -715 353 -714
rect 362 -715 363 -714
rect 366 -715 367 -714
rect 618 -715 619 -714
rect 44 -717 45 -716
rect 191 -717 192 -716
rect 233 -717 234 -716
rect 352 -717 353 -716
rect 359 -717 360 -716
rect 674 -717 675 -716
rect 44 -719 45 -718
rect 124 -719 125 -718
rect 135 -719 136 -718
rect 212 -719 213 -718
rect 247 -719 248 -718
rect 362 -719 363 -718
rect 373 -719 374 -718
rect 383 -719 384 -718
rect 408 -719 409 -718
rect 604 -719 605 -718
rect 58 -721 59 -720
rect 65 -721 66 -720
rect 142 -721 143 -720
rect 303 -721 304 -720
rect 317 -721 318 -720
rect 345 -721 346 -720
rect 373 -721 374 -720
rect 453 -721 454 -720
rect 548 -721 549 -720
rect 576 -721 577 -720
rect 583 -721 584 -720
rect 681 -721 682 -720
rect 65 -723 66 -722
rect 394 -723 395 -722
rect 415 -723 416 -722
rect 499 -723 500 -722
rect 562 -723 563 -722
rect 625 -723 626 -722
rect 142 -725 143 -724
rect 282 -725 283 -724
rect 296 -725 297 -724
rect 369 -725 370 -724
rect 436 -725 437 -724
rect 520 -725 521 -724
rect 565 -725 566 -724
rect 604 -725 605 -724
rect 149 -727 150 -726
rect 212 -727 213 -726
rect 247 -727 248 -726
rect 667 -727 668 -726
rect 114 -729 115 -728
rect 149 -729 150 -728
rect 156 -729 157 -728
rect 387 -729 388 -728
rect 443 -729 444 -728
rect 457 -729 458 -728
rect 492 -729 493 -728
rect 548 -729 549 -728
rect 590 -729 591 -728
rect 646 -729 647 -728
rect 114 -731 115 -730
rect 205 -731 206 -730
rect 261 -731 262 -730
rect 733 -731 734 -730
rect 184 -733 185 -732
rect 205 -733 206 -732
rect 278 -733 279 -732
rect 324 -733 325 -732
rect 331 -733 332 -732
rect 380 -733 381 -732
rect 450 -733 451 -732
rect 471 -733 472 -732
rect 492 -733 493 -732
rect 590 -733 591 -732
rect 597 -733 598 -732
rect 618 -733 619 -732
rect 639 -733 640 -732
rect 667 -733 668 -732
rect 170 -735 171 -734
rect 184 -735 185 -734
rect 191 -735 192 -734
rect 268 -735 269 -734
rect 299 -735 300 -734
rect 338 -735 339 -734
rect 348 -735 349 -734
rect 415 -735 416 -734
rect 453 -735 454 -734
rect 660 -735 661 -734
rect 107 -737 108 -736
rect 268 -737 269 -736
rect 317 -737 318 -736
rect 327 -737 328 -736
rect 366 -737 367 -736
rect 562 -737 563 -736
rect 107 -739 108 -738
rect 177 -739 178 -738
rect 243 -739 244 -738
rect 639 -739 640 -738
rect 170 -741 171 -740
rect 198 -741 199 -740
rect 376 -741 377 -740
rect 443 -741 444 -740
rect 506 -741 507 -740
rect 520 -741 521 -740
rect 555 -741 556 -740
rect 597 -741 598 -740
rect 51 -743 52 -742
rect 198 -743 199 -742
rect 380 -743 381 -742
rect 702 -743 703 -742
rect 177 -745 178 -744
rect 292 -745 293 -744
rect 383 -745 384 -744
rect 660 -745 661 -744
rect 485 -747 486 -746
rect 506 -747 507 -746
rect 513 -747 514 -746
rect 555 -747 556 -746
rect 485 -749 486 -748
rect 513 -749 514 -748
rect 30 -760 31 -759
rect 408 -760 409 -759
rect 429 -760 430 -759
rect 751 -760 752 -759
rect 30 -762 31 -761
rect 82 -762 83 -761
rect 89 -762 90 -761
rect 149 -762 150 -761
rect 177 -762 178 -761
rect 229 -762 230 -761
rect 243 -762 244 -761
rect 275 -762 276 -761
rect 289 -762 290 -761
rect 310 -762 311 -761
rect 327 -762 328 -761
rect 639 -762 640 -761
rect 674 -762 675 -761
rect 730 -762 731 -761
rect 733 -762 734 -761
rect 744 -762 745 -761
rect 2 -764 3 -763
rect 89 -764 90 -763
rect 107 -764 108 -763
rect 201 -764 202 -763
rect 226 -764 227 -763
rect 345 -764 346 -763
rect 387 -764 388 -763
rect 716 -764 717 -763
rect 723 -764 724 -763
rect 737 -764 738 -763
rect 23 -766 24 -765
rect 387 -766 388 -765
rect 390 -766 391 -765
rect 590 -766 591 -765
rect 604 -766 605 -765
rect 765 -766 766 -765
rect 23 -768 24 -767
rect 54 -768 55 -767
rect 58 -768 59 -767
rect 86 -768 87 -767
rect 100 -768 101 -767
rect 107 -768 108 -767
rect 121 -768 122 -767
rect 138 -768 139 -767
rect 142 -768 143 -767
rect 285 -768 286 -767
rect 299 -768 300 -767
rect 408 -768 409 -767
rect 422 -768 423 -767
rect 737 -768 738 -767
rect 37 -770 38 -769
rect 93 -770 94 -769
rect 100 -770 101 -769
rect 254 -770 255 -769
rect 261 -770 262 -769
rect 324 -770 325 -769
rect 334 -770 335 -769
rect 513 -770 514 -769
rect 527 -770 528 -769
rect 625 -770 626 -769
rect 632 -770 633 -769
rect 744 -770 745 -769
rect 51 -772 52 -771
rect 674 -772 675 -771
rect 702 -772 703 -771
rect 758 -772 759 -771
rect 58 -774 59 -773
rect 191 -774 192 -773
rect 247 -774 248 -773
rect 254 -774 255 -773
rect 341 -774 342 -773
rect 443 -774 444 -773
rect 495 -774 496 -773
rect 646 -774 647 -773
rect 712 -774 713 -773
rect 786 -774 787 -773
rect 65 -776 66 -775
rect 383 -776 384 -775
rect 390 -776 391 -775
rect 422 -776 423 -775
rect 436 -776 437 -775
rect 723 -776 724 -775
rect 65 -778 66 -777
rect 86 -778 87 -777
rect 93 -778 94 -777
rect 250 -778 251 -777
rect 345 -778 346 -777
rect 352 -778 353 -777
rect 373 -778 374 -777
rect 513 -778 514 -777
rect 541 -778 542 -777
rect 653 -778 654 -777
rect 72 -780 73 -779
rect 79 -780 80 -779
rect 121 -780 122 -779
rect 716 -780 717 -779
rect 72 -782 73 -781
rect 191 -782 192 -781
rect 247 -782 248 -781
rect 317 -782 318 -781
rect 352 -782 353 -781
rect 418 -782 419 -781
rect 439 -782 440 -781
rect 639 -782 640 -781
rect 79 -784 80 -783
rect 264 -784 265 -783
rect 303 -784 304 -783
rect 653 -784 654 -783
rect 124 -786 125 -785
rect 163 -786 164 -785
rect 170 -786 171 -785
rect 310 -786 311 -785
rect 373 -786 374 -785
rect 380 -786 381 -785
rect 383 -786 384 -785
rect 772 -786 773 -785
rect 2 -788 3 -787
rect 163 -788 164 -787
rect 170 -788 171 -787
rect 292 -788 293 -787
rect 303 -788 304 -787
rect 331 -788 332 -787
rect 380 -788 381 -787
rect 604 -788 605 -787
rect 611 -788 612 -787
rect 625 -788 626 -787
rect 632 -788 633 -787
rect 667 -788 668 -787
rect 9 -790 10 -789
rect 124 -790 125 -789
rect 149 -790 150 -789
rect 240 -790 241 -789
rect 394 -790 395 -789
rect 460 -790 461 -789
rect 464 -790 465 -789
rect 541 -790 542 -789
rect 544 -790 545 -789
rect 709 -790 710 -789
rect 9 -792 10 -791
rect 128 -792 129 -791
rect 156 -792 157 -791
rect 226 -792 227 -791
rect 240 -792 241 -791
rect 793 -792 794 -791
rect 16 -794 17 -793
rect 331 -794 332 -793
rect 362 -794 363 -793
rect 464 -794 465 -793
rect 488 -794 489 -793
rect 646 -794 647 -793
rect 16 -796 17 -795
rect 135 -796 136 -795
rect 156 -796 157 -795
rect 215 -796 216 -795
rect 397 -796 398 -795
rect 450 -796 451 -795
rect 453 -796 454 -795
rect 667 -796 668 -795
rect 44 -798 45 -797
rect 135 -798 136 -797
rect 177 -798 178 -797
rect 198 -798 199 -797
rect 212 -798 213 -797
rect 317 -798 318 -797
rect 366 -798 367 -797
rect 450 -798 451 -797
rect 548 -798 549 -797
rect 583 -798 584 -797
rect 586 -798 587 -797
rect 688 -798 689 -797
rect 44 -800 45 -799
rect 338 -800 339 -799
rect 404 -800 405 -799
rect 583 -800 584 -799
rect 590 -800 591 -799
rect 597 -800 598 -799
rect 618 -800 619 -799
rect 702 -800 703 -799
rect 128 -802 129 -801
rect 219 -802 220 -801
rect 222 -802 223 -801
rect 338 -802 339 -801
rect 411 -802 412 -801
rect 443 -802 444 -801
rect 534 -802 535 -801
rect 618 -802 619 -801
rect 681 -802 682 -801
rect 688 -802 689 -801
rect 103 -804 104 -803
rect 534 -804 535 -803
rect 555 -804 556 -803
rect 681 -804 682 -803
rect 184 -806 185 -805
rect 212 -806 213 -805
rect 219 -806 220 -805
rect 268 -806 269 -805
rect 415 -806 416 -805
rect 495 -806 496 -805
rect 520 -806 521 -805
rect 555 -806 556 -805
rect 562 -806 563 -805
rect 695 -806 696 -805
rect 114 -808 115 -807
rect 184 -808 185 -807
rect 198 -808 199 -807
rect 660 -808 661 -807
rect 695 -808 696 -807
rect 754 -808 755 -807
rect 110 -810 111 -809
rect 114 -810 115 -809
rect 233 -810 234 -809
rect 366 -810 367 -809
rect 436 -810 437 -809
rect 597 -810 598 -809
rect 205 -812 206 -811
rect 233 -812 234 -811
rect 268 -812 269 -811
rect 401 -812 402 -811
rect 499 -812 500 -811
rect 562 -812 563 -811
rect 569 -812 570 -811
rect 779 -812 780 -811
rect 205 -814 206 -813
rect 236 -814 237 -813
rect 359 -814 360 -813
rect 569 -814 570 -813
rect 576 -814 577 -813
rect 611 -814 612 -813
rect 296 -816 297 -815
rect 359 -816 360 -815
rect 499 -816 500 -815
rect 506 -816 507 -815
rect 520 -816 521 -815
rect 803 -816 804 -815
rect 296 -818 297 -817
rect 548 -818 549 -817
rect 471 -820 472 -819
rect 506 -820 507 -819
rect 523 -820 524 -819
rect 576 -820 577 -819
rect 457 -822 458 -821
rect 471 -822 472 -821
rect 530 -822 531 -821
rect 660 -822 661 -821
rect 457 -824 458 -823
rect 478 -824 479 -823
rect 478 -826 479 -825
rect 492 -826 493 -825
rect 9 -837 10 -836
rect 240 -837 241 -836
rect 278 -837 279 -836
rect 793 -837 794 -836
rect 803 -837 804 -836
rect 807 -837 808 -836
rect 9 -839 10 -838
rect 149 -839 150 -838
rect 159 -839 160 -838
rect 457 -839 458 -838
rect 460 -839 461 -838
rect 765 -839 766 -838
rect 16 -841 17 -840
rect 173 -841 174 -840
rect 184 -841 185 -840
rect 296 -841 297 -840
rect 366 -841 367 -840
rect 436 -841 437 -840
rect 439 -841 440 -840
rect 779 -841 780 -840
rect 16 -843 17 -842
rect 180 -843 181 -842
rect 184 -843 185 -842
rect 352 -843 353 -842
rect 359 -843 360 -842
rect 436 -843 437 -842
rect 460 -843 461 -842
rect 737 -843 738 -842
rect 751 -843 752 -842
rect 775 -843 776 -842
rect 23 -845 24 -844
rect 145 -845 146 -844
rect 149 -845 150 -844
rect 401 -845 402 -844
rect 404 -845 405 -844
rect 562 -845 563 -844
rect 730 -845 731 -844
rect 737 -845 738 -844
rect 751 -845 752 -844
rect 782 -845 783 -844
rect 30 -847 31 -846
rect 236 -847 237 -846
rect 240 -847 241 -846
rect 247 -847 248 -846
rect 268 -847 269 -846
rect 352 -847 353 -846
rect 366 -847 367 -846
rect 387 -847 388 -846
rect 390 -847 391 -846
rect 786 -847 787 -846
rect 37 -849 38 -848
rect 86 -849 87 -848
rect 107 -849 108 -848
rect 156 -849 157 -848
rect 166 -849 167 -848
rect 212 -849 213 -848
rect 215 -849 216 -848
rect 674 -849 675 -848
rect 716 -849 717 -848
rect 730 -849 731 -848
rect 786 -849 787 -848
rect 796 -849 797 -848
rect 44 -851 45 -850
rect 138 -851 139 -850
rect 156 -851 157 -850
rect 534 -851 535 -850
rect 667 -851 668 -850
rect 674 -851 675 -850
rect 54 -853 55 -852
rect 772 -853 773 -852
rect 58 -855 59 -854
rect 299 -855 300 -854
rect 338 -855 339 -854
rect 667 -855 668 -854
rect 72 -857 73 -856
rect 247 -857 248 -856
rect 268 -857 269 -856
rect 317 -857 318 -856
rect 373 -857 374 -856
rect 534 -857 535 -856
rect 646 -857 647 -856
rect 772 -857 773 -856
rect 51 -859 52 -858
rect 72 -859 73 -858
rect 82 -859 83 -858
rect 639 -859 640 -858
rect 128 -861 129 -860
rect 212 -861 213 -860
rect 219 -861 220 -860
rect 243 -861 244 -860
rect 275 -861 276 -860
rect 338 -861 339 -860
rect 383 -861 384 -860
rect 765 -861 766 -860
rect 2 -863 3 -862
rect 275 -863 276 -862
rect 282 -863 283 -862
rect 317 -863 318 -862
rect 397 -863 398 -862
rect 604 -863 605 -862
rect 44 -865 45 -864
rect 128 -865 129 -864
rect 135 -865 136 -864
rect 429 -865 430 -864
rect 467 -865 468 -864
rect 681 -865 682 -864
rect 170 -867 171 -866
rect 187 -867 188 -866
rect 201 -867 202 -866
rect 359 -867 360 -866
rect 401 -867 402 -866
rect 415 -867 416 -866
rect 418 -867 419 -866
rect 618 -867 619 -866
rect 93 -869 94 -868
rect 201 -869 202 -868
rect 226 -869 227 -868
rect 289 -869 290 -868
rect 292 -869 293 -868
rect 716 -869 717 -868
rect 58 -871 59 -870
rect 226 -871 227 -870
rect 229 -871 230 -870
rect 660 -871 661 -870
rect 93 -873 94 -872
rect 114 -873 115 -872
rect 170 -873 171 -872
rect 254 -873 255 -872
rect 282 -873 283 -872
rect 373 -873 374 -872
rect 411 -873 412 -872
rect 660 -873 661 -872
rect 114 -875 115 -874
rect 121 -875 122 -874
rect 177 -875 178 -874
rect 219 -875 220 -874
rect 233 -875 234 -874
rect 261 -875 262 -874
rect 296 -875 297 -874
rect 310 -875 311 -874
rect 334 -875 335 -874
rect 429 -875 430 -874
rect 488 -875 489 -874
rect 709 -875 710 -874
rect 37 -877 38 -876
rect 233 -877 234 -876
rect 303 -877 304 -876
rect 310 -877 311 -876
rect 348 -877 349 -876
rect 709 -877 710 -876
rect 65 -879 66 -878
rect 121 -879 122 -878
rect 177 -879 178 -878
rect 653 -879 654 -878
rect 65 -881 66 -880
rect 163 -881 164 -880
rect 187 -881 188 -880
rect 254 -881 255 -880
rect 303 -881 304 -880
rect 394 -881 395 -880
rect 422 -881 423 -880
rect 492 -881 493 -880
rect 506 -881 507 -880
rect 520 -881 521 -880
rect 523 -881 524 -880
rect 744 -881 745 -880
rect 324 -883 325 -882
rect 422 -883 423 -882
rect 488 -883 489 -882
rect 723 -883 724 -882
rect 191 -885 192 -884
rect 324 -885 325 -884
rect 394 -885 395 -884
rect 541 -885 542 -884
rect 569 -885 570 -884
rect 646 -885 647 -884
rect 653 -885 654 -884
rect 695 -885 696 -884
rect 450 -887 451 -886
rect 541 -887 542 -886
rect 576 -887 577 -886
rect 604 -887 605 -886
rect 611 -887 612 -886
rect 681 -887 682 -886
rect 695 -887 696 -886
rect 702 -887 703 -886
rect 450 -889 451 -888
rect 758 -889 759 -888
rect 464 -891 465 -890
rect 611 -891 612 -890
rect 618 -891 619 -890
rect 632 -891 633 -890
rect 152 -893 153 -892
rect 632 -893 633 -892
rect 464 -895 465 -894
rect 569 -895 570 -894
rect 583 -895 584 -894
rect 758 -895 759 -894
rect 495 -897 496 -896
rect 702 -897 703 -896
rect 499 -899 500 -898
rect 506 -899 507 -898
rect 513 -899 514 -898
rect 562 -899 563 -898
rect 583 -899 584 -898
rect 590 -899 591 -898
rect 478 -901 479 -900
rect 513 -901 514 -900
rect 527 -901 528 -900
rect 744 -901 745 -900
rect 100 -903 101 -902
rect 478 -903 479 -902
rect 499 -903 500 -902
rect 639 -903 640 -902
rect 79 -905 80 -904
rect 100 -905 101 -904
rect 443 -905 444 -904
rect 527 -905 528 -904
rect 530 -905 531 -904
rect 548 -905 549 -904
rect 590 -905 591 -904
rect 597 -905 598 -904
rect 79 -907 80 -906
rect 345 -907 346 -906
rect 485 -907 486 -906
rect 548 -907 549 -906
rect 555 -907 556 -906
rect 597 -907 598 -906
rect 331 -909 332 -908
rect 443 -909 444 -908
rect 471 -909 472 -908
rect 555 -909 556 -908
rect 331 -911 332 -910
rect 380 -911 381 -910
rect 408 -911 409 -910
rect 471 -911 472 -910
rect 408 -913 409 -912
rect 723 -913 724 -912
rect 9 -924 10 -923
rect 222 -924 223 -923
rect 229 -924 230 -923
rect 338 -924 339 -923
rect 348 -924 349 -923
rect 611 -924 612 -923
rect 723 -924 724 -923
rect 754 -924 755 -923
rect 779 -924 780 -923
rect 786 -924 787 -923
rect 9 -926 10 -925
rect 352 -926 353 -925
rect 366 -926 367 -925
rect 443 -926 444 -925
rect 446 -926 447 -925
rect 730 -926 731 -925
rect 751 -926 752 -925
rect 775 -926 776 -925
rect 16 -928 17 -927
rect 117 -928 118 -927
rect 121 -928 122 -927
rect 128 -928 129 -927
rect 142 -928 143 -927
rect 152 -928 153 -927
rect 159 -928 160 -927
rect 425 -928 426 -927
rect 432 -928 433 -927
rect 513 -928 514 -927
rect 576 -928 577 -927
rect 730 -928 731 -927
rect 16 -930 17 -929
rect 100 -930 101 -929
rect 107 -930 108 -929
rect 142 -930 143 -929
rect 149 -930 150 -929
rect 373 -930 374 -929
rect 408 -930 409 -929
rect 534 -930 535 -929
rect 576 -930 577 -929
rect 646 -930 647 -929
rect 723 -930 724 -929
rect 740 -930 741 -929
rect 23 -932 24 -931
rect 233 -932 234 -931
rect 236 -932 237 -931
rect 653 -932 654 -931
rect 23 -934 24 -933
rect 103 -934 104 -933
rect 107 -934 108 -933
rect 275 -934 276 -933
rect 285 -934 286 -933
rect 422 -934 423 -933
rect 460 -934 461 -933
rect 737 -934 738 -933
rect 30 -936 31 -935
rect 411 -936 412 -935
rect 415 -936 416 -935
rect 485 -936 486 -935
rect 499 -936 500 -935
rect 695 -936 696 -935
rect 30 -938 31 -937
rect 184 -938 185 -937
rect 191 -938 192 -937
rect 198 -938 199 -937
rect 201 -938 202 -937
rect 502 -938 503 -937
rect 513 -938 514 -937
rect 555 -938 556 -937
rect 579 -938 580 -937
rect 604 -938 605 -937
rect 681 -938 682 -937
rect 737 -938 738 -937
rect 37 -940 38 -939
rect 82 -940 83 -939
rect 86 -940 87 -939
rect 257 -940 258 -939
rect 275 -940 276 -939
rect 303 -940 304 -939
rect 310 -940 311 -939
rect 313 -940 314 -939
rect 317 -940 318 -939
rect 380 -940 381 -939
rect 418 -940 419 -939
rect 597 -940 598 -939
rect 604 -940 605 -939
rect 625 -940 626 -939
rect 674 -940 675 -939
rect 681 -940 682 -939
rect 37 -942 38 -941
rect 75 -942 76 -941
rect 86 -942 87 -941
rect 96 -942 97 -941
rect 114 -942 115 -941
rect 121 -942 122 -941
rect 135 -942 136 -941
rect 233 -942 234 -941
rect 243 -942 244 -941
rect 261 -942 262 -941
rect 296 -942 297 -941
rect 303 -942 304 -941
rect 348 -942 349 -941
rect 401 -942 402 -941
rect 418 -942 419 -941
rect 499 -942 500 -941
rect 527 -942 528 -941
rect 625 -942 626 -941
rect 44 -944 45 -943
rect 397 -944 398 -943
rect 464 -944 465 -943
rect 765 -944 766 -943
rect 51 -946 52 -945
rect 100 -946 101 -945
rect 114 -946 115 -945
rect 653 -946 654 -945
rect 51 -948 52 -947
rect 93 -948 94 -947
rect 149 -948 150 -947
rect 285 -948 286 -947
rect 359 -948 360 -947
rect 401 -948 402 -947
rect 467 -948 468 -947
rect 744 -948 745 -947
rect 65 -950 66 -949
rect 289 -950 290 -949
rect 397 -950 398 -949
rect 436 -950 437 -949
rect 471 -950 472 -949
rect 611 -950 612 -949
rect 618 -950 619 -949
rect 674 -950 675 -949
rect 79 -952 80 -951
rect 135 -952 136 -951
rect 163 -952 164 -951
rect 408 -952 409 -951
rect 488 -952 489 -951
rect 695 -952 696 -951
rect 44 -954 45 -953
rect 79 -954 80 -953
rect 89 -954 90 -953
rect 562 -954 563 -953
rect 590 -954 591 -953
rect 646 -954 647 -953
rect 163 -956 164 -955
rect 212 -956 213 -955
rect 226 -956 227 -955
rect 338 -956 339 -955
rect 429 -956 430 -955
rect 590 -956 591 -955
rect 597 -956 598 -955
rect 660 -956 661 -955
rect 58 -958 59 -957
rect 429 -958 430 -957
rect 506 -958 507 -957
rect 562 -958 563 -957
rect 618 -958 619 -957
rect 772 -958 773 -957
rect 58 -960 59 -959
rect 474 -960 475 -959
rect 478 -960 479 -959
rect 506 -960 507 -959
rect 520 -960 521 -959
rect 527 -960 528 -959
rect 534 -960 535 -959
rect 758 -960 759 -959
rect 170 -962 171 -961
rect 443 -962 444 -961
rect 457 -962 458 -961
rect 478 -962 479 -961
rect 555 -962 556 -961
rect 569 -962 570 -961
rect 632 -962 633 -961
rect 660 -962 661 -961
rect 177 -964 178 -963
rect 376 -964 377 -963
rect 390 -964 391 -963
rect 569 -964 570 -963
rect 583 -964 584 -963
rect 632 -964 633 -963
rect 180 -966 181 -965
rect 380 -966 381 -965
rect 457 -966 458 -965
rect 492 -966 493 -965
rect 583 -966 584 -965
rect 639 -966 640 -965
rect 184 -968 185 -967
rect 268 -968 269 -967
rect 278 -968 279 -967
rect 758 -968 759 -967
rect 191 -970 192 -969
rect 205 -970 206 -969
rect 212 -970 213 -969
rect 219 -970 220 -969
rect 226 -970 227 -969
rect 317 -970 318 -969
rect 471 -970 472 -969
rect 520 -970 521 -969
rect 639 -970 640 -969
rect 667 -970 668 -969
rect 205 -972 206 -971
rect 240 -972 241 -971
rect 243 -972 244 -971
rect 331 -972 332 -971
rect 492 -972 493 -971
rect 541 -972 542 -971
rect 667 -972 668 -971
rect 702 -972 703 -971
rect 198 -974 199 -973
rect 331 -974 332 -973
rect 702 -974 703 -973
rect 709 -974 710 -973
rect 219 -976 220 -975
rect 261 -976 262 -975
rect 268 -976 269 -975
rect 324 -976 325 -975
rect 709 -976 710 -975
rect 716 -976 717 -975
rect 247 -978 248 -977
rect 345 -978 346 -977
rect 394 -978 395 -977
rect 716 -978 717 -977
rect 236 -980 237 -979
rect 247 -980 248 -979
rect 254 -980 255 -979
rect 362 -980 363 -979
rect 254 -982 255 -981
rect 541 -982 542 -981
rect 289 -984 290 -983
rect 450 -984 451 -983
rect 296 -986 297 -985
rect 450 -986 451 -985
rect 310 -988 311 -987
rect 436 -988 437 -987
rect 324 -990 325 -989
rect 387 -990 388 -989
rect 9 -1001 10 -1000
rect 317 -1001 318 -1000
rect 334 -1001 335 -1000
rect 408 -1001 409 -1000
rect 411 -1001 412 -1000
rect 513 -1001 514 -1000
rect 737 -1001 738 -1000
rect 744 -1001 745 -1000
rect 16 -1003 17 -1002
rect 194 -1003 195 -1002
rect 198 -1003 199 -1002
rect 369 -1003 370 -1002
rect 373 -1003 374 -1002
rect 383 -1003 384 -1002
rect 394 -1003 395 -1002
rect 404 -1003 405 -1002
rect 408 -1003 409 -1002
rect 464 -1003 465 -1002
rect 471 -1003 472 -1002
rect 674 -1003 675 -1002
rect 740 -1003 741 -1002
rect 758 -1003 759 -1002
rect 23 -1005 24 -1004
rect 240 -1005 241 -1004
rect 243 -1005 244 -1004
rect 359 -1005 360 -1004
rect 362 -1005 363 -1004
rect 576 -1005 577 -1004
rect 23 -1007 24 -1006
rect 149 -1007 150 -1006
rect 166 -1007 167 -1006
rect 222 -1007 223 -1006
rect 233 -1007 234 -1006
rect 331 -1007 332 -1006
rect 338 -1007 339 -1006
rect 366 -1007 367 -1006
rect 373 -1007 374 -1006
rect 555 -1007 556 -1006
rect 576 -1007 577 -1006
rect 691 -1007 692 -1006
rect 30 -1009 31 -1008
rect 243 -1009 244 -1008
rect 250 -1009 251 -1008
rect 261 -1009 262 -1008
rect 268 -1009 269 -1008
rect 317 -1009 318 -1008
rect 338 -1009 339 -1008
rect 499 -1009 500 -1008
rect 33 -1011 34 -1010
rect 180 -1011 181 -1010
rect 191 -1011 192 -1010
rect 219 -1011 220 -1010
rect 247 -1011 248 -1010
rect 261 -1011 262 -1010
rect 282 -1011 283 -1010
rect 639 -1011 640 -1010
rect 37 -1013 38 -1012
rect 79 -1013 80 -1012
rect 107 -1013 108 -1012
rect 310 -1013 311 -1012
rect 345 -1013 346 -1012
rect 730 -1013 731 -1012
rect 37 -1015 38 -1014
rect 107 -1015 108 -1014
rect 114 -1015 115 -1014
rect 754 -1015 755 -1014
rect 44 -1017 45 -1016
rect 61 -1017 62 -1016
rect 65 -1017 66 -1016
rect 93 -1017 94 -1016
rect 114 -1017 115 -1016
rect 121 -1017 122 -1016
rect 142 -1017 143 -1016
rect 152 -1017 153 -1016
rect 170 -1017 171 -1016
rect 219 -1017 220 -1016
rect 296 -1017 297 -1016
rect 345 -1017 346 -1016
rect 348 -1017 349 -1016
rect 439 -1017 440 -1016
rect 443 -1017 444 -1016
rect 548 -1017 549 -1016
rect 562 -1017 563 -1016
rect 730 -1017 731 -1016
rect 51 -1019 52 -1018
rect 117 -1019 118 -1018
rect 121 -1019 122 -1018
rect 184 -1019 185 -1018
rect 205 -1019 206 -1018
rect 254 -1019 255 -1018
rect 275 -1019 276 -1018
rect 296 -1019 297 -1018
rect 352 -1019 353 -1018
rect 618 -1019 619 -1018
rect 51 -1021 52 -1020
rect 103 -1021 104 -1020
rect 135 -1021 136 -1020
rect 142 -1021 143 -1020
rect 149 -1021 150 -1020
rect 233 -1021 234 -1020
rect 352 -1021 353 -1020
rect 355 -1021 356 -1020
rect 376 -1021 377 -1020
rect 506 -1021 507 -1020
rect 590 -1021 591 -1020
rect 618 -1021 619 -1020
rect 58 -1023 59 -1022
rect 184 -1023 185 -1022
rect 191 -1023 192 -1022
rect 205 -1023 206 -1022
rect 212 -1023 213 -1022
rect 282 -1023 283 -1022
rect 380 -1023 381 -1022
rect 387 -1023 388 -1022
rect 415 -1023 416 -1022
rect 660 -1023 661 -1022
rect 65 -1025 66 -1024
rect 96 -1025 97 -1024
rect 135 -1025 136 -1024
rect 159 -1025 160 -1024
rect 163 -1025 164 -1024
rect 254 -1025 255 -1024
rect 380 -1025 381 -1024
rect 583 -1025 584 -1024
rect 590 -1025 591 -1024
rect 597 -1025 598 -1024
rect 72 -1027 73 -1026
rect 86 -1027 87 -1026
rect 170 -1027 171 -1026
rect 226 -1027 227 -1026
rect 383 -1027 384 -1026
rect 555 -1027 556 -1026
rect 597 -1027 598 -1026
rect 653 -1027 654 -1026
rect 44 -1029 45 -1028
rect 86 -1029 87 -1028
rect 156 -1029 157 -1028
rect 226 -1029 227 -1028
rect 310 -1029 311 -1028
rect 653 -1029 654 -1028
rect 75 -1031 76 -1030
rect 163 -1031 164 -1030
rect 397 -1031 398 -1030
rect 583 -1031 584 -1030
rect 79 -1033 80 -1032
rect 128 -1033 129 -1032
rect 156 -1033 157 -1032
rect 177 -1033 178 -1032
rect 418 -1033 419 -1032
rect 457 -1033 458 -1032
rect 478 -1033 479 -1032
rect 548 -1033 549 -1032
rect 128 -1035 129 -1034
rect 289 -1035 290 -1034
rect 401 -1035 402 -1034
rect 457 -1035 458 -1034
rect 478 -1035 479 -1034
rect 709 -1035 710 -1034
rect 177 -1037 178 -1036
rect 268 -1037 269 -1036
rect 289 -1037 290 -1036
rect 324 -1037 325 -1036
rect 401 -1037 402 -1036
rect 625 -1037 626 -1036
rect 646 -1037 647 -1036
rect 709 -1037 710 -1036
rect 324 -1039 325 -1038
rect 520 -1039 521 -1038
rect 625 -1039 626 -1038
rect 695 -1039 696 -1038
rect 313 -1041 314 -1040
rect 695 -1041 696 -1040
rect 212 -1043 213 -1042
rect 313 -1043 314 -1042
rect 425 -1043 426 -1042
rect 660 -1043 661 -1042
rect 432 -1045 433 -1044
rect 674 -1045 675 -1044
rect 436 -1047 437 -1046
rect 443 -1047 444 -1046
rect 446 -1047 447 -1046
rect 492 -1047 493 -1046
rect 495 -1047 496 -1046
rect 513 -1047 514 -1046
rect 520 -1047 521 -1046
rect 534 -1047 535 -1046
rect 646 -1047 647 -1046
rect 702 -1047 703 -1046
rect 450 -1049 451 -1048
rect 611 -1049 612 -1048
rect 702 -1049 703 -1048
rect 723 -1049 724 -1048
rect 453 -1051 454 -1050
rect 667 -1051 668 -1050
rect 467 -1053 468 -1052
rect 611 -1053 612 -1052
rect 667 -1053 668 -1052
rect 716 -1053 717 -1052
rect 485 -1055 486 -1054
rect 639 -1055 640 -1054
rect 716 -1055 717 -1054
rect 737 -1055 738 -1054
rect 278 -1057 279 -1056
rect 485 -1057 486 -1056
rect 492 -1057 493 -1056
rect 569 -1057 570 -1056
rect 499 -1059 500 -1058
rect 527 -1059 528 -1058
rect 541 -1059 542 -1058
rect 723 -1059 724 -1058
rect 425 -1061 426 -1060
rect 527 -1061 528 -1060
rect 569 -1061 570 -1060
rect 632 -1061 633 -1060
rect 429 -1063 430 -1062
rect 541 -1063 542 -1062
rect 632 -1063 633 -1062
rect 681 -1063 682 -1062
rect 681 -1065 682 -1064
rect 719 -1065 720 -1064
rect 9 -1076 10 -1075
rect 121 -1076 122 -1075
rect 128 -1076 129 -1075
rect 215 -1076 216 -1075
rect 243 -1076 244 -1075
rect 362 -1076 363 -1075
rect 387 -1076 388 -1075
rect 415 -1076 416 -1075
rect 418 -1076 419 -1075
rect 660 -1076 661 -1075
rect 677 -1076 678 -1075
rect 688 -1076 689 -1075
rect 16 -1078 17 -1077
rect 30 -1078 31 -1077
rect 37 -1078 38 -1077
rect 180 -1078 181 -1077
rect 187 -1078 188 -1077
rect 261 -1078 262 -1077
rect 278 -1078 279 -1077
rect 303 -1078 304 -1077
rect 313 -1078 314 -1077
rect 408 -1078 409 -1077
rect 415 -1078 416 -1077
rect 457 -1078 458 -1077
rect 478 -1078 479 -1077
rect 691 -1078 692 -1077
rect 44 -1080 45 -1079
rect 124 -1080 125 -1079
rect 128 -1080 129 -1079
rect 212 -1080 213 -1079
rect 254 -1080 255 -1079
rect 310 -1080 311 -1079
rect 324 -1080 325 -1079
rect 387 -1080 388 -1079
rect 394 -1080 395 -1079
rect 436 -1080 437 -1079
rect 485 -1080 486 -1079
rect 716 -1080 717 -1079
rect 51 -1082 52 -1081
rect 149 -1082 150 -1081
rect 166 -1082 167 -1081
rect 201 -1082 202 -1081
rect 282 -1082 283 -1081
rect 303 -1082 304 -1081
rect 310 -1082 311 -1081
rect 681 -1082 682 -1081
rect 51 -1084 52 -1083
rect 82 -1084 83 -1083
rect 86 -1084 87 -1083
rect 240 -1084 241 -1083
rect 282 -1084 283 -1083
rect 366 -1084 367 -1083
rect 401 -1084 402 -1083
rect 478 -1084 479 -1083
rect 495 -1084 496 -1083
rect 632 -1084 633 -1083
rect 65 -1086 66 -1085
rect 177 -1086 178 -1085
rect 194 -1086 195 -1085
rect 317 -1086 318 -1085
rect 324 -1086 325 -1085
rect 348 -1086 349 -1085
rect 359 -1086 360 -1085
rect 457 -1086 458 -1085
rect 464 -1086 465 -1085
rect 485 -1086 486 -1085
rect 499 -1086 500 -1085
rect 506 -1086 507 -1085
rect 534 -1086 535 -1085
rect 590 -1086 591 -1085
rect 611 -1086 612 -1085
rect 681 -1086 682 -1085
rect 58 -1088 59 -1087
rect 65 -1088 66 -1087
rect 72 -1088 73 -1087
rect 156 -1088 157 -1087
rect 177 -1088 178 -1087
rect 261 -1088 262 -1087
rect 289 -1088 290 -1087
rect 317 -1088 318 -1087
rect 334 -1088 335 -1087
rect 618 -1088 619 -1087
rect 632 -1088 633 -1087
rect 674 -1088 675 -1087
rect 79 -1090 80 -1089
rect 159 -1090 160 -1089
rect 198 -1090 199 -1089
rect 338 -1090 339 -1089
rect 345 -1090 346 -1089
rect 401 -1090 402 -1089
rect 422 -1090 423 -1089
rect 730 -1090 731 -1089
rect 23 -1092 24 -1091
rect 198 -1092 199 -1091
rect 289 -1092 290 -1091
rect 429 -1092 430 -1091
rect 439 -1092 440 -1091
rect 499 -1092 500 -1091
rect 506 -1092 507 -1091
rect 569 -1092 570 -1091
rect 583 -1092 584 -1091
rect 590 -1092 591 -1091
rect 611 -1092 612 -1091
rect 667 -1092 668 -1091
rect 93 -1094 94 -1093
rect 383 -1094 384 -1093
rect 422 -1094 423 -1093
rect 471 -1094 472 -1093
rect 513 -1094 514 -1093
rect 534 -1094 535 -1093
rect 537 -1094 538 -1093
rect 674 -1094 675 -1093
rect 37 -1096 38 -1095
rect 93 -1096 94 -1095
rect 100 -1096 101 -1095
rect 142 -1096 143 -1095
rect 145 -1096 146 -1095
rect 254 -1096 255 -1095
rect 268 -1096 269 -1095
rect 429 -1096 430 -1095
rect 453 -1096 454 -1095
rect 667 -1096 668 -1095
rect 107 -1098 108 -1097
rect 170 -1098 171 -1097
rect 268 -1098 269 -1097
rect 481 -1098 482 -1097
rect 513 -1098 514 -1097
rect 576 -1098 577 -1097
rect 583 -1098 584 -1097
rect 597 -1098 598 -1097
rect 618 -1098 619 -1097
rect 695 -1098 696 -1097
rect 135 -1100 136 -1099
rect 278 -1100 279 -1099
rect 296 -1100 297 -1099
rect 397 -1100 398 -1099
rect 523 -1100 524 -1099
rect 569 -1100 570 -1099
rect 576 -1100 577 -1099
rect 723 -1100 724 -1099
rect 135 -1102 136 -1101
rect 226 -1102 227 -1101
rect 296 -1102 297 -1101
rect 562 -1102 563 -1101
rect 565 -1102 566 -1101
rect 604 -1102 605 -1101
rect 684 -1102 685 -1101
rect 695 -1102 696 -1101
rect 142 -1104 143 -1103
rect 380 -1104 381 -1103
rect 523 -1104 524 -1103
rect 660 -1104 661 -1103
rect 149 -1106 150 -1105
rect 233 -1106 234 -1105
rect 275 -1106 276 -1105
rect 604 -1106 605 -1105
rect 184 -1108 185 -1107
rect 226 -1108 227 -1107
rect 338 -1108 339 -1107
rect 492 -1108 493 -1107
rect 541 -1108 542 -1107
rect 646 -1108 647 -1107
rect 23 -1110 24 -1109
rect 184 -1110 185 -1109
rect 219 -1110 220 -1109
rect 233 -1110 234 -1109
rect 247 -1110 248 -1109
rect 492 -1110 493 -1109
rect 555 -1110 556 -1109
rect 562 -1110 563 -1109
rect 597 -1110 598 -1109
rect 653 -1110 654 -1109
rect 68 -1112 69 -1111
rect 646 -1112 647 -1111
rect 205 -1114 206 -1113
rect 219 -1114 220 -1113
rect 373 -1114 374 -1113
rect 464 -1114 465 -1113
rect 548 -1114 549 -1113
rect 555 -1114 556 -1113
rect 205 -1116 206 -1115
rect 331 -1116 332 -1115
rect 380 -1116 381 -1115
rect 639 -1116 640 -1115
rect 376 -1118 377 -1117
rect 639 -1118 640 -1117
rect 425 -1120 426 -1119
rect 541 -1120 542 -1119
rect 548 -1120 549 -1119
rect 625 -1120 626 -1119
rect 425 -1122 426 -1121
rect 709 -1122 710 -1121
rect 450 -1124 451 -1123
rect 653 -1124 654 -1123
rect 709 -1124 710 -1123
rect 737 -1124 738 -1123
rect 411 -1126 412 -1125
rect 450 -1126 451 -1125
rect 474 -1126 475 -1125
rect 625 -1126 626 -1125
rect 2 -1137 3 -1136
rect 128 -1137 129 -1136
rect 145 -1137 146 -1136
rect 152 -1137 153 -1136
rect 159 -1137 160 -1136
rect 268 -1137 269 -1136
rect 275 -1137 276 -1136
rect 296 -1137 297 -1136
rect 303 -1137 304 -1136
rect 310 -1137 311 -1136
rect 317 -1137 318 -1136
rect 359 -1137 360 -1136
rect 369 -1137 370 -1136
rect 639 -1137 640 -1136
rect 646 -1137 647 -1136
rect 674 -1137 675 -1136
rect 677 -1137 678 -1136
rect 709 -1137 710 -1136
rect 9 -1139 10 -1138
rect 163 -1139 164 -1138
rect 170 -1139 171 -1138
rect 562 -1139 563 -1138
rect 646 -1139 647 -1138
rect 653 -1139 654 -1138
rect 677 -1139 678 -1138
rect 681 -1139 682 -1138
rect 695 -1139 696 -1138
rect 709 -1139 710 -1138
rect 9 -1141 10 -1140
rect 247 -1141 248 -1140
rect 250 -1141 251 -1140
rect 457 -1141 458 -1140
rect 506 -1141 507 -1140
rect 520 -1141 521 -1140
rect 523 -1141 524 -1140
rect 527 -1141 528 -1140
rect 530 -1141 531 -1140
rect 534 -1141 535 -1140
rect 544 -1141 545 -1140
rect 639 -1141 640 -1140
rect 16 -1143 17 -1142
rect 44 -1143 45 -1142
rect 47 -1143 48 -1142
rect 58 -1143 59 -1142
rect 72 -1143 73 -1142
rect 194 -1143 195 -1142
rect 219 -1143 220 -1142
rect 247 -1143 248 -1142
rect 261 -1143 262 -1142
rect 373 -1143 374 -1142
rect 380 -1143 381 -1142
rect 401 -1143 402 -1142
rect 429 -1143 430 -1142
rect 555 -1143 556 -1142
rect 562 -1143 563 -1142
rect 618 -1143 619 -1142
rect 37 -1145 38 -1144
rect 65 -1145 66 -1144
rect 79 -1145 80 -1144
rect 331 -1145 332 -1144
rect 334 -1145 335 -1144
rect 443 -1145 444 -1144
rect 478 -1145 479 -1144
rect 506 -1145 507 -1144
rect 590 -1145 591 -1144
rect 618 -1145 619 -1144
rect 37 -1147 38 -1146
rect 320 -1147 321 -1146
rect 331 -1147 332 -1146
rect 492 -1147 493 -1146
rect 583 -1147 584 -1146
rect 590 -1147 591 -1146
rect 44 -1149 45 -1148
rect 215 -1149 216 -1148
rect 226 -1149 227 -1148
rect 261 -1149 262 -1148
rect 278 -1149 279 -1148
rect 625 -1149 626 -1148
rect 51 -1151 52 -1150
rect 75 -1151 76 -1150
rect 93 -1151 94 -1150
rect 180 -1151 181 -1150
rect 184 -1151 185 -1150
rect 254 -1151 255 -1150
rect 282 -1151 283 -1150
rect 422 -1151 423 -1150
rect 429 -1151 430 -1150
rect 436 -1151 437 -1150
rect 471 -1151 472 -1150
rect 478 -1151 479 -1150
rect 492 -1151 493 -1150
rect 513 -1151 514 -1150
rect 541 -1151 542 -1150
rect 583 -1151 584 -1150
rect 604 -1151 605 -1150
rect 625 -1151 626 -1150
rect 51 -1153 52 -1152
rect 149 -1153 150 -1152
rect 156 -1153 157 -1152
rect 254 -1153 255 -1152
rect 310 -1153 311 -1152
rect 324 -1153 325 -1152
rect 345 -1153 346 -1152
rect 499 -1153 500 -1152
rect 19 -1155 20 -1154
rect 324 -1155 325 -1154
rect 348 -1155 349 -1154
rect 569 -1155 570 -1154
rect 58 -1157 59 -1156
rect 205 -1157 206 -1156
rect 226 -1157 227 -1156
rect 303 -1157 304 -1156
rect 317 -1157 318 -1156
rect 667 -1157 668 -1156
rect 82 -1159 83 -1158
rect 93 -1159 94 -1158
rect 100 -1159 101 -1158
rect 194 -1159 195 -1158
rect 205 -1159 206 -1158
rect 219 -1159 220 -1158
rect 233 -1159 234 -1158
rect 268 -1159 269 -1158
rect 348 -1159 349 -1158
rect 352 -1159 353 -1158
rect 373 -1159 374 -1158
rect 408 -1159 409 -1158
rect 415 -1159 416 -1158
rect 422 -1159 423 -1158
rect 432 -1159 433 -1158
rect 534 -1159 535 -1158
rect 569 -1159 570 -1158
rect 632 -1159 633 -1158
rect 660 -1159 661 -1158
rect 667 -1159 668 -1158
rect 86 -1161 87 -1160
rect 282 -1161 283 -1160
rect 387 -1161 388 -1160
rect 408 -1161 409 -1160
rect 443 -1161 444 -1160
rect 604 -1161 605 -1160
rect 632 -1161 633 -1160
rect 656 -1161 657 -1160
rect 30 -1163 31 -1162
rect 86 -1163 87 -1162
rect 107 -1163 108 -1162
rect 208 -1163 209 -1162
rect 236 -1163 237 -1162
rect 296 -1163 297 -1162
rect 394 -1163 395 -1162
rect 401 -1163 402 -1162
rect 450 -1163 451 -1162
rect 471 -1163 472 -1162
rect 485 -1163 486 -1162
rect 499 -1163 500 -1162
rect 107 -1165 108 -1164
rect 114 -1165 115 -1164
rect 121 -1165 122 -1164
rect 233 -1165 234 -1164
rect 362 -1165 363 -1164
rect 394 -1165 395 -1164
rect 397 -1165 398 -1164
rect 576 -1165 577 -1164
rect 23 -1167 24 -1166
rect 114 -1167 115 -1166
rect 121 -1167 122 -1166
rect 338 -1167 339 -1166
rect 387 -1167 388 -1166
rect 576 -1167 577 -1166
rect 110 -1169 111 -1168
rect 128 -1169 129 -1168
rect 135 -1169 136 -1168
rect 352 -1169 353 -1168
rect 450 -1169 451 -1168
rect 548 -1169 549 -1168
rect 135 -1171 136 -1170
rect 149 -1171 150 -1170
rect 156 -1171 157 -1170
rect 177 -1171 178 -1170
rect 184 -1171 185 -1170
rect 198 -1171 199 -1170
rect 338 -1171 339 -1170
rect 513 -1171 514 -1170
rect 548 -1171 549 -1170
rect 597 -1171 598 -1170
rect 142 -1173 143 -1172
rect 660 -1173 661 -1172
rect 142 -1175 143 -1174
rect 457 -1175 458 -1174
rect 485 -1175 486 -1174
rect 674 -1175 675 -1174
rect 145 -1177 146 -1176
rect 366 -1177 367 -1176
rect 597 -1177 598 -1176
rect 611 -1177 612 -1176
rect 163 -1179 164 -1178
rect 170 -1179 171 -1178
rect 173 -1179 174 -1178
rect 240 -1179 241 -1178
rect 366 -1179 367 -1178
rect 390 -1179 391 -1178
rect 446 -1179 447 -1178
rect 611 -1179 612 -1178
rect 166 -1181 167 -1180
rect 555 -1181 556 -1180
rect 191 -1183 192 -1182
rect 198 -1183 199 -1182
rect 390 -1183 391 -1182
rect 415 -1183 416 -1182
rect 2 -1194 3 -1193
rect 152 -1194 153 -1193
rect 156 -1194 157 -1193
rect 163 -1194 164 -1193
rect 166 -1194 167 -1193
rect 191 -1194 192 -1193
rect 201 -1194 202 -1193
rect 257 -1194 258 -1193
rect 275 -1194 276 -1193
rect 296 -1194 297 -1193
rect 303 -1194 304 -1193
rect 429 -1194 430 -1193
rect 436 -1194 437 -1193
rect 576 -1194 577 -1193
rect 667 -1194 668 -1193
rect 681 -1194 682 -1193
rect 702 -1194 703 -1193
rect 705 -1194 706 -1193
rect 709 -1194 710 -1193
rect 716 -1194 717 -1193
rect 2 -1196 3 -1195
rect 107 -1196 108 -1195
rect 110 -1196 111 -1195
rect 187 -1196 188 -1195
rect 215 -1196 216 -1195
rect 247 -1196 248 -1195
rect 296 -1196 297 -1195
rect 506 -1196 507 -1195
rect 530 -1196 531 -1195
rect 632 -1196 633 -1195
rect 674 -1196 675 -1195
rect 688 -1196 689 -1195
rect 9 -1198 10 -1197
rect 23 -1198 24 -1197
rect 30 -1198 31 -1197
rect 275 -1198 276 -1197
rect 306 -1198 307 -1197
rect 352 -1198 353 -1197
rect 383 -1198 384 -1197
rect 464 -1198 465 -1197
rect 541 -1198 542 -1197
rect 590 -1198 591 -1197
rect 597 -1198 598 -1197
rect 674 -1198 675 -1197
rect 9 -1200 10 -1199
rect 44 -1200 45 -1199
rect 54 -1200 55 -1199
rect 212 -1200 213 -1199
rect 229 -1200 230 -1199
rect 282 -1200 283 -1199
rect 289 -1200 290 -1199
rect 306 -1200 307 -1199
rect 310 -1200 311 -1199
rect 317 -1200 318 -1199
rect 320 -1200 321 -1199
rect 632 -1200 633 -1199
rect 16 -1202 17 -1201
rect 75 -1202 76 -1201
rect 89 -1202 90 -1201
rect 520 -1202 521 -1201
rect 562 -1202 563 -1201
rect 653 -1202 654 -1201
rect 23 -1204 24 -1203
rect 149 -1204 150 -1203
rect 198 -1204 199 -1203
rect 289 -1204 290 -1203
rect 310 -1204 311 -1203
rect 688 -1204 689 -1203
rect 30 -1206 31 -1205
rect 107 -1206 108 -1205
rect 117 -1206 118 -1205
rect 408 -1206 409 -1205
rect 436 -1206 437 -1205
rect 471 -1206 472 -1205
rect 478 -1206 479 -1205
rect 541 -1206 542 -1205
rect 562 -1206 563 -1205
rect 702 -1206 703 -1205
rect 37 -1208 38 -1207
rect 124 -1208 125 -1207
rect 142 -1208 143 -1207
rect 506 -1208 507 -1207
rect 569 -1208 570 -1207
rect 681 -1208 682 -1207
rect 37 -1210 38 -1209
rect 184 -1210 185 -1209
rect 219 -1210 220 -1209
rect 282 -1210 283 -1209
rect 324 -1210 325 -1209
rect 373 -1210 374 -1209
rect 387 -1210 388 -1209
rect 422 -1210 423 -1209
rect 443 -1210 444 -1209
rect 555 -1210 556 -1209
rect 597 -1210 598 -1209
rect 611 -1210 612 -1209
rect 58 -1212 59 -1211
rect 173 -1212 174 -1211
rect 233 -1212 234 -1211
rect 660 -1212 661 -1211
rect 58 -1214 59 -1213
rect 86 -1214 87 -1213
rect 100 -1214 101 -1213
rect 457 -1214 458 -1213
rect 460 -1214 461 -1213
rect 576 -1214 577 -1213
rect 65 -1216 66 -1215
rect 75 -1216 76 -1215
rect 100 -1216 101 -1215
rect 114 -1216 115 -1215
rect 121 -1216 122 -1215
rect 205 -1216 206 -1215
rect 240 -1216 241 -1215
rect 338 -1216 339 -1215
rect 341 -1216 342 -1215
rect 380 -1216 381 -1215
rect 387 -1216 388 -1215
rect 453 -1216 454 -1215
rect 499 -1216 500 -1215
rect 520 -1216 521 -1215
rect 548 -1216 549 -1215
rect 555 -1216 556 -1215
rect 72 -1218 73 -1217
rect 170 -1218 171 -1217
rect 194 -1218 195 -1217
rect 240 -1218 241 -1217
rect 247 -1218 248 -1217
rect 625 -1218 626 -1217
rect 145 -1220 146 -1219
rect 250 -1220 251 -1219
rect 327 -1220 328 -1219
rect 485 -1220 486 -1219
rect 513 -1220 514 -1219
rect 569 -1220 570 -1219
rect 149 -1222 150 -1221
rect 177 -1222 178 -1221
rect 254 -1222 255 -1221
rect 485 -1222 486 -1221
rect 513 -1222 514 -1221
rect 660 -1222 661 -1221
rect 51 -1224 52 -1223
rect 177 -1224 178 -1223
rect 327 -1224 328 -1223
rect 604 -1224 605 -1223
rect 334 -1226 335 -1225
rect 478 -1226 479 -1225
rect 604 -1226 605 -1225
rect 639 -1226 640 -1225
rect 348 -1228 349 -1227
rect 625 -1228 626 -1227
rect 352 -1230 353 -1229
rect 471 -1230 472 -1229
rect 583 -1230 584 -1229
rect 639 -1230 640 -1229
rect 366 -1232 367 -1231
rect 408 -1232 409 -1231
rect 429 -1232 430 -1231
rect 548 -1232 549 -1231
rect 135 -1234 136 -1233
rect 366 -1234 367 -1233
rect 373 -1234 374 -1233
rect 397 -1234 398 -1233
rect 401 -1234 402 -1233
rect 422 -1234 423 -1233
rect 432 -1234 433 -1233
rect 443 -1234 444 -1233
rect 446 -1234 447 -1233
rect 590 -1234 591 -1233
rect 79 -1236 80 -1235
rect 135 -1236 136 -1235
rect 380 -1236 381 -1235
rect 618 -1236 619 -1235
rect 79 -1238 80 -1237
rect 128 -1238 129 -1237
rect 331 -1238 332 -1237
rect 618 -1238 619 -1237
rect 128 -1240 129 -1239
rect 226 -1240 227 -1239
rect 394 -1240 395 -1239
rect 611 -1240 612 -1239
rect 226 -1242 227 -1241
rect 261 -1242 262 -1241
rect 401 -1242 402 -1241
rect 467 -1242 468 -1241
rect 534 -1242 535 -1241
rect 583 -1242 584 -1241
rect 254 -1244 255 -1243
rect 394 -1244 395 -1243
rect 450 -1244 451 -1243
rect 646 -1244 647 -1243
rect 261 -1246 262 -1245
rect 268 -1246 269 -1245
rect 415 -1246 416 -1245
rect 646 -1246 647 -1245
rect 170 -1248 171 -1247
rect 268 -1248 269 -1247
rect 345 -1248 346 -1247
rect 415 -1248 416 -1247
rect 450 -1248 451 -1247
rect 695 -1248 696 -1247
rect 345 -1250 346 -1249
rect 390 -1250 391 -1249
rect 453 -1250 454 -1249
rect 492 -1250 493 -1249
rect 534 -1250 535 -1249
rect 712 -1250 713 -1249
rect 457 -1252 458 -1251
rect 499 -1252 500 -1251
rect 492 -1254 493 -1253
rect 527 -1254 528 -1253
rect 16 -1265 17 -1264
rect 61 -1265 62 -1264
rect 72 -1265 73 -1264
rect 688 -1265 689 -1264
rect 712 -1265 713 -1264
rect 716 -1265 717 -1264
rect 2 -1267 3 -1266
rect 72 -1267 73 -1266
rect 93 -1267 94 -1266
rect 103 -1267 104 -1266
rect 107 -1267 108 -1266
rect 313 -1267 314 -1266
rect 317 -1267 318 -1266
rect 383 -1267 384 -1266
rect 394 -1267 395 -1266
rect 681 -1267 682 -1266
rect 2 -1269 3 -1268
rect 135 -1269 136 -1268
rect 142 -1269 143 -1268
rect 156 -1269 157 -1268
rect 177 -1269 178 -1268
rect 250 -1269 251 -1268
rect 254 -1269 255 -1268
rect 261 -1269 262 -1268
rect 271 -1269 272 -1268
rect 527 -1269 528 -1268
rect 667 -1269 668 -1268
rect 670 -1269 671 -1268
rect 9 -1271 10 -1270
rect 135 -1271 136 -1270
rect 145 -1271 146 -1270
rect 289 -1271 290 -1270
rect 303 -1271 304 -1270
rect 702 -1271 703 -1270
rect 9 -1273 10 -1272
rect 187 -1273 188 -1272
rect 194 -1273 195 -1272
rect 366 -1273 367 -1272
rect 397 -1273 398 -1272
rect 611 -1273 612 -1272
rect 667 -1273 668 -1272
rect 695 -1273 696 -1272
rect 702 -1273 703 -1272
rect 705 -1273 706 -1272
rect 23 -1275 24 -1274
rect 191 -1275 192 -1274
rect 208 -1275 209 -1274
rect 219 -1275 220 -1274
rect 222 -1275 223 -1274
rect 254 -1275 255 -1274
rect 257 -1275 258 -1274
rect 289 -1275 290 -1274
rect 303 -1275 304 -1274
rect 443 -1275 444 -1274
rect 460 -1275 461 -1274
rect 527 -1275 528 -1274
rect 23 -1277 24 -1276
rect 79 -1277 80 -1276
rect 86 -1277 87 -1276
rect 93 -1277 94 -1276
rect 100 -1277 101 -1276
rect 114 -1277 115 -1276
rect 128 -1277 129 -1276
rect 198 -1277 199 -1276
rect 215 -1277 216 -1276
rect 338 -1277 339 -1276
rect 352 -1277 353 -1276
rect 597 -1277 598 -1276
rect 30 -1279 31 -1278
rect 86 -1279 87 -1278
rect 114 -1279 115 -1278
rect 233 -1279 234 -1278
rect 236 -1279 237 -1278
rect 317 -1279 318 -1278
rect 324 -1279 325 -1278
rect 408 -1279 409 -1278
rect 429 -1279 430 -1278
rect 534 -1279 535 -1278
rect 576 -1279 577 -1278
rect 597 -1279 598 -1278
rect 37 -1281 38 -1280
rect 331 -1281 332 -1280
rect 362 -1281 363 -1280
rect 520 -1281 521 -1280
rect 534 -1281 535 -1280
rect 555 -1281 556 -1280
rect 569 -1281 570 -1280
rect 576 -1281 577 -1280
rect 40 -1283 41 -1282
rect 65 -1283 66 -1282
rect 131 -1283 132 -1282
rect 236 -1283 237 -1282
rect 285 -1283 286 -1282
rect 625 -1283 626 -1282
rect 44 -1285 45 -1284
rect 82 -1285 83 -1284
rect 149 -1285 150 -1284
rect 156 -1285 157 -1284
rect 177 -1285 178 -1284
rect 646 -1285 647 -1284
rect 44 -1287 45 -1286
rect 205 -1287 206 -1286
rect 219 -1287 220 -1286
rect 474 -1287 475 -1286
rect 495 -1287 496 -1286
rect 625 -1287 626 -1286
rect 47 -1289 48 -1288
rect 478 -1289 479 -1288
rect 506 -1289 507 -1288
rect 681 -1289 682 -1288
rect 51 -1291 52 -1290
rect 163 -1291 164 -1290
rect 180 -1291 181 -1290
rect 191 -1291 192 -1290
rect 226 -1291 227 -1290
rect 247 -1291 248 -1290
rect 310 -1291 311 -1290
rect 355 -1291 356 -1290
rect 366 -1291 367 -1290
rect 569 -1291 570 -1290
rect 58 -1293 59 -1292
rect 121 -1293 122 -1292
rect 163 -1293 164 -1292
rect 275 -1293 276 -1292
rect 327 -1293 328 -1292
rect 331 -1293 332 -1292
rect 380 -1293 381 -1292
rect 611 -1293 612 -1292
rect 65 -1295 66 -1294
rect 205 -1295 206 -1294
rect 233 -1295 234 -1294
rect 453 -1295 454 -1294
rect 478 -1295 479 -1294
rect 492 -1295 493 -1294
rect 513 -1295 514 -1294
rect 639 -1295 640 -1294
rect 121 -1297 122 -1296
rect 138 -1297 139 -1296
rect 184 -1297 185 -1296
rect 296 -1297 297 -1296
rect 380 -1297 381 -1296
rect 415 -1297 416 -1296
rect 422 -1297 423 -1296
rect 555 -1297 556 -1296
rect 639 -1297 640 -1296
rect 660 -1297 661 -1296
rect 170 -1299 171 -1298
rect 184 -1299 185 -1298
rect 247 -1299 248 -1298
rect 306 -1299 307 -1298
rect 373 -1299 374 -1298
rect 415 -1299 416 -1298
rect 432 -1299 433 -1298
rect 436 -1299 437 -1298
rect 443 -1299 444 -1298
rect 502 -1299 503 -1298
rect 520 -1299 521 -1298
rect 562 -1299 563 -1298
rect 632 -1299 633 -1298
rect 660 -1299 661 -1298
rect 268 -1301 269 -1300
rect 422 -1301 423 -1300
rect 436 -1301 437 -1300
rect 485 -1301 486 -1300
rect 562 -1301 563 -1300
rect 604 -1301 605 -1300
rect 268 -1303 269 -1302
rect 282 -1303 283 -1302
rect 296 -1303 297 -1302
rect 387 -1303 388 -1302
rect 397 -1303 398 -1302
rect 457 -1303 458 -1302
rect 464 -1303 465 -1302
rect 604 -1303 605 -1302
rect 261 -1305 262 -1304
rect 282 -1305 283 -1304
rect 306 -1305 307 -1304
rect 359 -1305 360 -1304
rect 373 -1305 374 -1304
rect 513 -1305 514 -1304
rect 590 -1305 591 -1304
rect 632 -1305 633 -1304
rect 275 -1307 276 -1306
rect 369 -1307 370 -1306
rect 401 -1307 402 -1306
rect 506 -1307 507 -1306
rect 324 -1309 325 -1308
rect 590 -1309 591 -1308
rect 390 -1311 391 -1310
rect 401 -1311 402 -1310
rect 408 -1311 409 -1310
rect 471 -1311 472 -1310
rect 485 -1311 486 -1310
rect 548 -1311 549 -1310
rect 464 -1313 465 -1312
rect 618 -1313 619 -1312
rect 548 -1315 549 -1314
rect 583 -1315 584 -1314
rect 618 -1315 619 -1314
rect 653 -1315 654 -1314
rect 180 -1317 181 -1316
rect 583 -1317 584 -1316
rect 499 -1319 500 -1318
rect 653 -1319 654 -1318
rect 499 -1321 500 -1320
rect 674 -1321 675 -1320
rect 541 -1323 542 -1322
rect 674 -1323 675 -1322
rect 450 -1325 451 -1324
rect 541 -1325 542 -1324
rect 2 -1336 3 -1335
rect 177 -1336 178 -1335
rect 208 -1336 209 -1335
rect 268 -1336 269 -1335
rect 303 -1336 304 -1335
rect 397 -1336 398 -1335
rect 404 -1336 405 -1335
rect 457 -1336 458 -1335
rect 460 -1336 461 -1335
rect 604 -1336 605 -1335
rect 653 -1336 654 -1335
rect 670 -1336 671 -1335
rect 9 -1338 10 -1337
rect 201 -1338 202 -1337
rect 212 -1338 213 -1337
rect 282 -1338 283 -1337
rect 338 -1338 339 -1337
rect 590 -1338 591 -1337
rect 646 -1338 647 -1337
rect 653 -1338 654 -1337
rect 667 -1338 668 -1337
rect 681 -1338 682 -1337
rect 19 -1340 20 -1339
rect 114 -1340 115 -1339
rect 135 -1340 136 -1339
rect 233 -1340 234 -1339
rect 254 -1340 255 -1339
rect 359 -1340 360 -1339
rect 366 -1340 367 -1339
rect 597 -1340 598 -1339
rect 646 -1340 647 -1339
rect 656 -1340 657 -1339
rect 33 -1342 34 -1341
rect 131 -1342 132 -1341
rect 138 -1342 139 -1341
rect 299 -1342 300 -1341
rect 338 -1342 339 -1341
rect 415 -1342 416 -1341
rect 422 -1342 423 -1341
rect 576 -1342 577 -1341
rect 590 -1342 591 -1341
rect 639 -1342 640 -1341
rect 44 -1344 45 -1343
rect 369 -1344 370 -1343
rect 373 -1344 374 -1343
rect 513 -1344 514 -1343
rect 576 -1344 577 -1343
rect 632 -1344 633 -1343
rect 51 -1346 52 -1345
rect 243 -1346 244 -1345
rect 261 -1346 262 -1345
rect 268 -1346 269 -1345
rect 275 -1346 276 -1345
rect 282 -1346 283 -1345
rect 352 -1346 353 -1345
rect 621 -1346 622 -1345
rect 58 -1348 59 -1347
rect 82 -1348 83 -1347
rect 100 -1348 101 -1347
rect 145 -1348 146 -1347
rect 149 -1348 150 -1347
rect 156 -1348 157 -1347
rect 159 -1348 160 -1347
rect 341 -1348 342 -1347
rect 366 -1348 367 -1347
rect 555 -1348 556 -1347
rect 58 -1350 59 -1349
rect 163 -1350 164 -1349
rect 177 -1350 178 -1349
rect 184 -1350 185 -1349
rect 219 -1350 220 -1349
rect 324 -1350 325 -1349
rect 380 -1350 381 -1349
rect 394 -1350 395 -1349
rect 408 -1350 409 -1349
rect 660 -1350 661 -1349
rect 37 -1352 38 -1351
rect 184 -1352 185 -1351
rect 222 -1352 223 -1351
rect 425 -1352 426 -1351
rect 450 -1352 451 -1351
rect 541 -1352 542 -1351
rect 51 -1354 52 -1353
rect 219 -1354 220 -1353
rect 226 -1354 227 -1353
rect 254 -1354 255 -1353
rect 261 -1354 262 -1353
rect 345 -1354 346 -1353
rect 348 -1354 349 -1353
rect 408 -1354 409 -1353
rect 425 -1354 426 -1353
rect 611 -1354 612 -1353
rect 65 -1356 66 -1355
rect 327 -1356 328 -1355
rect 383 -1356 384 -1355
rect 527 -1356 528 -1355
rect 541 -1356 542 -1355
rect 674 -1356 675 -1355
rect 65 -1358 66 -1357
rect 138 -1358 139 -1357
rect 163 -1358 164 -1357
rect 198 -1358 199 -1357
rect 226 -1358 227 -1357
rect 250 -1358 251 -1357
rect 285 -1358 286 -1357
rect 345 -1358 346 -1357
rect 383 -1358 384 -1357
rect 390 -1358 391 -1357
rect 474 -1358 475 -1357
rect 618 -1358 619 -1357
rect 72 -1360 73 -1359
rect 152 -1360 153 -1359
rect 240 -1360 241 -1359
rect 275 -1360 276 -1359
rect 289 -1360 290 -1359
rect 352 -1360 353 -1359
rect 387 -1360 388 -1359
rect 436 -1360 437 -1359
rect 478 -1360 479 -1359
rect 569 -1360 570 -1359
rect 583 -1360 584 -1359
rect 611 -1360 612 -1359
rect 44 -1362 45 -1361
rect 240 -1362 241 -1361
rect 285 -1362 286 -1361
rect 289 -1362 290 -1361
rect 436 -1362 437 -1361
rect 443 -1362 444 -1361
rect 481 -1362 482 -1361
rect 625 -1362 626 -1361
rect 75 -1364 76 -1363
rect 93 -1364 94 -1363
rect 100 -1364 101 -1363
rect 170 -1364 171 -1363
rect 401 -1364 402 -1363
rect 443 -1364 444 -1363
rect 481 -1364 482 -1363
rect 604 -1364 605 -1363
rect 79 -1366 80 -1365
rect 247 -1366 248 -1365
rect 492 -1366 493 -1365
rect 527 -1366 528 -1365
rect 548 -1366 549 -1365
rect 569 -1366 570 -1365
rect 600 -1366 601 -1365
rect 625 -1366 626 -1365
rect 93 -1368 94 -1367
rect 121 -1368 122 -1367
rect 124 -1368 125 -1367
rect 324 -1368 325 -1367
rect 429 -1368 430 -1367
rect 548 -1368 549 -1367
rect 562 -1368 563 -1367
rect 583 -1368 584 -1367
rect 107 -1370 108 -1369
rect 173 -1370 174 -1369
rect 212 -1370 213 -1369
rect 247 -1370 248 -1369
rect 310 -1370 311 -1369
rect 562 -1370 563 -1369
rect 107 -1372 108 -1371
rect 205 -1372 206 -1371
rect 310 -1372 311 -1371
rect 362 -1372 363 -1371
rect 492 -1372 493 -1371
rect 506 -1372 507 -1371
rect 513 -1372 514 -1371
rect 534 -1372 535 -1371
rect 114 -1374 115 -1373
rect 142 -1374 143 -1373
rect 170 -1374 171 -1373
rect 191 -1374 192 -1373
rect 362 -1374 363 -1373
rect 555 -1374 556 -1373
rect 23 -1376 24 -1375
rect 191 -1376 192 -1375
rect 471 -1376 472 -1375
rect 534 -1376 535 -1375
rect 121 -1378 122 -1377
rect 317 -1378 318 -1377
rect 331 -1378 332 -1377
rect 471 -1378 472 -1377
rect 499 -1378 500 -1377
rect 639 -1378 640 -1377
rect 128 -1380 129 -1379
rect 198 -1380 199 -1379
rect 296 -1380 297 -1379
rect 331 -1380 332 -1379
rect 369 -1380 370 -1379
rect 499 -1380 500 -1379
rect 506 -1380 507 -1379
rect 520 -1380 521 -1379
rect 296 -1382 297 -1381
rect 418 -1382 419 -1381
rect 464 -1382 465 -1381
rect 520 -1382 521 -1381
rect 317 -1384 318 -1383
rect 390 -1384 391 -1383
rect 33 -1395 34 -1394
rect 219 -1395 220 -1394
rect 233 -1395 234 -1394
rect 296 -1395 297 -1394
rect 317 -1395 318 -1394
rect 355 -1395 356 -1394
rect 366 -1395 367 -1394
rect 450 -1395 451 -1394
rect 453 -1395 454 -1394
rect 569 -1395 570 -1394
rect 600 -1395 601 -1394
rect 667 -1395 668 -1394
rect 37 -1397 38 -1396
rect 205 -1397 206 -1396
rect 233 -1397 234 -1396
rect 520 -1397 521 -1396
rect 551 -1397 552 -1396
rect 590 -1397 591 -1396
rect 621 -1397 622 -1396
rect 639 -1397 640 -1396
rect 37 -1399 38 -1398
rect 310 -1399 311 -1398
rect 317 -1399 318 -1398
rect 327 -1399 328 -1398
rect 373 -1399 374 -1398
rect 387 -1399 388 -1398
rect 390 -1399 391 -1398
rect 443 -1399 444 -1398
rect 460 -1399 461 -1398
rect 597 -1399 598 -1398
rect 635 -1399 636 -1398
rect 660 -1399 661 -1398
rect 44 -1401 45 -1400
rect 369 -1401 370 -1400
rect 380 -1401 381 -1400
rect 485 -1401 486 -1400
rect 499 -1401 500 -1400
rect 590 -1401 591 -1400
rect 44 -1403 45 -1402
rect 138 -1403 139 -1402
rect 184 -1403 185 -1402
rect 352 -1403 353 -1402
rect 369 -1403 370 -1402
rect 562 -1403 563 -1402
rect 51 -1405 52 -1404
rect 271 -1405 272 -1404
rect 275 -1405 276 -1404
rect 285 -1405 286 -1404
rect 296 -1405 297 -1404
rect 324 -1405 325 -1404
rect 331 -1405 332 -1404
rect 380 -1405 381 -1404
rect 387 -1405 388 -1404
rect 429 -1405 430 -1404
rect 432 -1405 433 -1404
rect 534 -1405 535 -1404
rect 51 -1407 52 -1406
rect 114 -1407 115 -1406
rect 124 -1407 125 -1406
rect 135 -1407 136 -1406
rect 201 -1407 202 -1406
rect 401 -1407 402 -1406
rect 404 -1407 405 -1406
rect 429 -1407 430 -1406
rect 436 -1407 437 -1406
rect 457 -1407 458 -1406
rect 464 -1407 465 -1406
rect 506 -1407 507 -1406
rect 513 -1407 514 -1406
rect 534 -1407 535 -1406
rect 58 -1409 59 -1408
rect 156 -1409 157 -1408
rect 247 -1409 248 -1408
rect 548 -1409 549 -1408
rect 58 -1411 59 -1410
rect 163 -1411 164 -1410
rect 247 -1411 248 -1410
rect 450 -1411 451 -1410
rect 464 -1411 465 -1410
rect 583 -1411 584 -1410
rect 72 -1413 73 -1412
rect 236 -1413 237 -1412
rect 261 -1413 262 -1412
rect 376 -1413 377 -1412
rect 394 -1413 395 -1412
rect 415 -1413 416 -1412
rect 418 -1413 419 -1412
rect 527 -1413 528 -1412
rect 583 -1413 584 -1412
rect 625 -1413 626 -1412
rect 72 -1415 73 -1414
rect 149 -1415 150 -1414
rect 163 -1415 164 -1414
rect 177 -1415 178 -1414
rect 187 -1415 188 -1414
rect 394 -1415 395 -1414
rect 401 -1415 402 -1414
rect 443 -1415 444 -1414
rect 485 -1415 486 -1414
rect 541 -1415 542 -1414
rect 86 -1417 87 -1416
rect 103 -1417 104 -1416
rect 107 -1417 108 -1416
rect 345 -1417 346 -1416
rect 397 -1417 398 -1416
rect 541 -1417 542 -1416
rect 79 -1419 80 -1418
rect 86 -1419 87 -1418
rect 103 -1419 104 -1418
rect 289 -1419 290 -1418
rect 310 -1419 311 -1418
rect 373 -1419 374 -1418
rect 422 -1419 423 -1418
rect 565 -1419 566 -1418
rect 79 -1421 80 -1420
rect 226 -1421 227 -1420
rect 243 -1421 244 -1420
rect 527 -1421 528 -1420
rect 107 -1423 108 -1422
rect 121 -1423 122 -1422
rect 138 -1423 139 -1422
rect 149 -1423 150 -1422
rect 177 -1423 178 -1422
rect 359 -1423 360 -1422
rect 425 -1423 426 -1422
rect 520 -1423 521 -1422
rect 205 -1425 206 -1424
rect 226 -1425 227 -1424
rect 254 -1425 255 -1424
rect 261 -1425 262 -1424
rect 268 -1425 269 -1424
rect 366 -1425 367 -1424
rect 436 -1425 437 -1424
rect 576 -1425 577 -1424
rect 219 -1427 220 -1426
rect 268 -1427 269 -1426
rect 275 -1427 276 -1426
rect 383 -1427 384 -1426
rect 492 -1427 493 -1426
rect 506 -1427 507 -1426
rect 513 -1427 514 -1426
rect 555 -1427 556 -1426
rect 576 -1427 577 -1426
rect 611 -1427 612 -1426
rect 191 -1429 192 -1428
rect 555 -1429 556 -1428
rect 191 -1431 192 -1430
rect 212 -1431 213 -1430
rect 240 -1431 241 -1430
rect 254 -1431 255 -1430
rect 282 -1431 283 -1430
rect 499 -1431 500 -1430
rect 65 -1433 66 -1432
rect 212 -1433 213 -1432
rect 215 -1433 216 -1432
rect 282 -1433 283 -1432
rect 289 -1433 290 -1432
rect 303 -1433 304 -1432
rect 331 -1433 332 -1432
rect 338 -1433 339 -1432
rect 471 -1433 472 -1432
rect 492 -1433 493 -1432
rect 65 -1435 66 -1434
rect 170 -1435 171 -1434
rect 338 -1435 339 -1434
rect 446 -1435 447 -1434
rect 128 -1437 129 -1436
rect 303 -1437 304 -1436
rect 439 -1437 440 -1436
rect 471 -1437 472 -1436
rect 117 -1439 118 -1438
rect 128 -1439 129 -1438
rect 145 -1439 146 -1438
rect 170 -1439 171 -1438
rect 145 -1441 146 -1440
rect 408 -1441 409 -1440
rect 408 -1443 409 -1442
rect 548 -1443 549 -1442
rect 16 -1454 17 -1453
rect 177 -1454 178 -1453
rect 215 -1454 216 -1453
rect 387 -1454 388 -1453
rect 429 -1454 430 -1453
rect 569 -1454 570 -1453
rect 702 -1454 703 -1453
rect 712 -1454 713 -1453
rect 44 -1456 45 -1455
rect 117 -1456 118 -1455
rect 163 -1456 164 -1455
rect 198 -1456 199 -1455
rect 254 -1456 255 -1455
rect 306 -1456 307 -1455
rect 310 -1456 311 -1455
rect 439 -1456 440 -1455
rect 443 -1456 444 -1455
rect 534 -1456 535 -1455
rect 548 -1456 549 -1455
rect 590 -1456 591 -1455
rect 51 -1458 52 -1457
rect 180 -1458 181 -1457
rect 254 -1458 255 -1457
rect 310 -1458 311 -1457
rect 327 -1458 328 -1457
rect 331 -1458 332 -1457
rect 359 -1458 360 -1457
rect 415 -1458 416 -1457
rect 422 -1458 423 -1457
rect 443 -1458 444 -1457
rect 450 -1458 451 -1457
rect 492 -1458 493 -1457
rect 562 -1458 563 -1457
rect 604 -1458 605 -1457
rect 65 -1460 66 -1459
rect 243 -1460 244 -1459
rect 268 -1460 269 -1459
rect 394 -1460 395 -1459
rect 432 -1460 433 -1459
rect 485 -1460 486 -1459
rect 492 -1460 493 -1459
rect 527 -1460 528 -1459
rect 565 -1460 566 -1459
rect 597 -1460 598 -1459
rect 51 -1462 52 -1461
rect 65 -1462 66 -1461
rect 72 -1462 73 -1461
rect 233 -1462 234 -1461
rect 271 -1462 272 -1461
rect 408 -1462 409 -1461
rect 436 -1462 437 -1461
rect 506 -1462 507 -1461
rect 534 -1462 535 -1461
rect 565 -1462 566 -1461
rect 569 -1462 570 -1461
rect 583 -1462 584 -1461
rect 72 -1464 73 -1463
rect 191 -1464 192 -1463
rect 212 -1464 213 -1463
rect 233 -1464 234 -1463
rect 240 -1464 241 -1463
rect 408 -1464 409 -1463
rect 478 -1464 479 -1463
rect 520 -1464 521 -1463
rect 572 -1464 573 -1463
rect 583 -1464 584 -1463
rect 58 -1466 59 -1465
rect 240 -1466 241 -1465
rect 271 -1466 272 -1465
rect 303 -1466 304 -1465
rect 331 -1466 332 -1465
rect 457 -1466 458 -1465
rect 478 -1466 479 -1465
rect 541 -1466 542 -1465
rect 58 -1468 59 -1467
rect 247 -1468 248 -1467
rect 282 -1468 283 -1467
rect 366 -1468 367 -1467
rect 401 -1468 402 -1467
rect 485 -1468 486 -1467
rect 506 -1468 507 -1467
rect 562 -1468 563 -1467
rect 79 -1470 80 -1469
rect 184 -1470 185 -1469
rect 250 -1470 251 -1469
rect 401 -1470 402 -1469
rect 457 -1470 458 -1469
rect 499 -1470 500 -1469
rect 520 -1470 521 -1469
rect 576 -1470 577 -1469
rect 79 -1472 80 -1471
rect 219 -1472 220 -1471
rect 261 -1472 262 -1471
rect 282 -1472 283 -1471
rect 289 -1472 290 -1471
rect 387 -1472 388 -1471
rect 429 -1472 430 -1471
rect 499 -1472 500 -1471
rect 541 -1472 542 -1471
rect 555 -1472 556 -1471
rect 576 -1472 577 -1471
rect 590 -1472 591 -1471
rect 37 -1474 38 -1473
rect 289 -1474 290 -1473
rect 292 -1474 293 -1473
rect 373 -1474 374 -1473
rect 37 -1476 38 -1475
rect 44 -1476 45 -1475
rect 86 -1476 87 -1475
rect 156 -1476 157 -1475
rect 163 -1476 164 -1475
rect 226 -1476 227 -1475
rect 261 -1476 262 -1475
rect 338 -1476 339 -1475
rect 345 -1476 346 -1475
rect 415 -1476 416 -1475
rect 30 -1478 31 -1477
rect 86 -1478 87 -1477
rect 93 -1478 94 -1477
rect 135 -1478 136 -1477
rect 142 -1478 143 -1477
rect 198 -1478 199 -1477
rect 205 -1478 206 -1477
rect 219 -1478 220 -1477
rect 296 -1478 297 -1477
rect 345 -1478 346 -1477
rect 359 -1478 360 -1477
rect 380 -1478 381 -1477
rect 93 -1480 94 -1479
rect 107 -1480 108 -1479
rect 110 -1480 111 -1479
rect 142 -1480 143 -1479
rect 149 -1480 150 -1479
rect 191 -1480 192 -1479
rect 296 -1480 297 -1479
rect 464 -1480 465 -1479
rect 100 -1482 101 -1481
rect 425 -1482 426 -1481
rect 107 -1484 108 -1483
rect 166 -1484 167 -1483
rect 170 -1484 171 -1483
rect 229 -1484 230 -1483
rect 338 -1484 339 -1483
rect 471 -1484 472 -1483
rect 114 -1486 115 -1485
rect 128 -1486 129 -1485
rect 135 -1486 136 -1485
rect 275 -1486 276 -1485
rect 369 -1486 370 -1485
rect 555 -1486 556 -1485
rect 128 -1488 129 -1487
rect 159 -1488 160 -1487
rect 177 -1488 178 -1487
rect 352 -1488 353 -1487
rect 380 -1488 381 -1487
rect 446 -1488 447 -1487
rect 471 -1488 472 -1487
rect 513 -1488 514 -1487
rect 124 -1490 125 -1489
rect 513 -1490 514 -1489
rect 156 -1492 157 -1491
rect 527 -1492 528 -1491
rect 275 -1494 276 -1493
rect 324 -1494 325 -1493
rect 390 -1494 391 -1493
rect 464 -1494 465 -1493
rect 317 -1496 318 -1495
rect 324 -1496 325 -1495
rect 16 -1507 17 -1506
rect 170 -1507 171 -1506
rect 173 -1507 174 -1506
rect 198 -1507 199 -1506
rect 205 -1507 206 -1506
rect 275 -1507 276 -1506
rect 292 -1507 293 -1506
rect 443 -1507 444 -1506
rect 464 -1507 465 -1506
rect 474 -1507 475 -1506
rect 478 -1507 479 -1506
rect 513 -1507 514 -1506
rect 565 -1507 566 -1506
rect 569 -1507 570 -1506
rect 579 -1507 580 -1506
rect 583 -1507 584 -1506
rect 23 -1509 24 -1508
rect 54 -1509 55 -1508
rect 58 -1509 59 -1508
rect 121 -1509 122 -1508
rect 142 -1509 143 -1508
rect 177 -1509 178 -1508
rect 184 -1509 185 -1508
rect 359 -1509 360 -1508
rect 369 -1509 370 -1508
rect 436 -1509 437 -1508
rect 443 -1509 444 -1508
rect 450 -1509 451 -1508
rect 488 -1509 489 -1508
rect 555 -1509 556 -1508
rect 30 -1511 31 -1510
rect 58 -1511 59 -1510
rect 72 -1511 73 -1510
rect 149 -1511 150 -1510
rect 152 -1511 153 -1510
rect 170 -1511 171 -1510
rect 184 -1511 185 -1510
rect 289 -1511 290 -1510
rect 313 -1511 314 -1510
rect 415 -1511 416 -1510
rect 422 -1511 423 -1510
rect 520 -1511 521 -1510
rect 37 -1513 38 -1512
rect 51 -1513 52 -1512
rect 79 -1513 80 -1512
rect 121 -1513 122 -1512
rect 152 -1513 153 -1512
rect 201 -1513 202 -1512
rect 240 -1513 241 -1512
rect 541 -1513 542 -1512
rect 51 -1515 52 -1514
rect 93 -1515 94 -1514
rect 100 -1515 101 -1514
rect 142 -1515 143 -1514
rect 163 -1515 164 -1514
rect 240 -1515 241 -1514
rect 247 -1515 248 -1514
rect 303 -1515 304 -1514
rect 320 -1515 321 -1514
rect 492 -1515 493 -1514
rect 513 -1515 514 -1514
rect 548 -1515 549 -1514
rect 65 -1517 66 -1516
rect 79 -1517 80 -1516
rect 86 -1517 87 -1516
rect 254 -1517 255 -1516
rect 268 -1517 269 -1516
rect 282 -1517 283 -1516
rect 303 -1517 304 -1516
rect 345 -1517 346 -1516
rect 401 -1517 402 -1516
rect 425 -1517 426 -1516
rect 429 -1517 430 -1516
rect 464 -1517 465 -1516
rect 492 -1517 493 -1516
rect 527 -1517 528 -1516
rect 65 -1519 66 -1518
rect 208 -1519 209 -1518
rect 275 -1519 276 -1518
rect 373 -1519 374 -1518
rect 387 -1519 388 -1518
rect 527 -1519 528 -1518
rect 89 -1521 90 -1520
rect 180 -1521 181 -1520
rect 187 -1521 188 -1520
rect 254 -1521 255 -1520
rect 282 -1521 283 -1520
rect 310 -1521 311 -1520
rect 327 -1521 328 -1520
rect 485 -1521 486 -1520
rect 520 -1521 521 -1520
rect 562 -1521 563 -1520
rect 110 -1523 111 -1522
rect 128 -1523 129 -1522
rect 135 -1523 136 -1522
rect 247 -1523 248 -1522
rect 261 -1523 262 -1522
rect 310 -1523 311 -1522
rect 331 -1523 332 -1522
rect 359 -1523 360 -1522
rect 373 -1523 374 -1522
rect 380 -1523 381 -1522
rect 383 -1523 384 -1522
rect 387 -1523 388 -1522
rect 436 -1523 437 -1522
rect 457 -1523 458 -1522
rect 114 -1525 115 -1524
rect 156 -1525 157 -1524
rect 191 -1525 192 -1524
rect 205 -1525 206 -1524
rect 229 -1525 230 -1524
rect 261 -1525 262 -1524
rect 380 -1525 381 -1524
rect 401 -1525 402 -1524
rect 450 -1525 451 -1524
rect 471 -1525 472 -1524
rect 96 -1527 97 -1526
rect 114 -1527 115 -1526
rect 128 -1527 129 -1526
rect 219 -1527 220 -1526
rect 236 -1527 237 -1526
rect 331 -1527 332 -1526
rect 457 -1527 458 -1526
rect 499 -1527 500 -1526
rect 135 -1529 136 -1528
rect 296 -1529 297 -1528
rect 499 -1529 500 -1528
rect 534 -1529 535 -1528
rect 156 -1531 157 -1530
rect 429 -1531 430 -1530
rect 198 -1533 199 -1532
rect 212 -1533 213 -1532
rect 236 -1533 237 -1532
rect 345 -1533 346 -1532
rect 212 -1535 213 -1534
rect 229 -1535 230 -1534
rect 296 -1535 297 -1534
rect 317 -1535 318 -1534
rect 317 -1537 318 -1536
rect 408 -1537 409 -1536
rect 352 -1539 353 -1538
rect 408 -1539 409 -1538
rect 352 -1541 353 -1540
rect 394 -1541 395 -1540
rect 338 -1543 339 -1542
rect 394 -1543 395 -1542
rect 338 -1545 339 -1544
rect 576 -1545 577 -1544
rect 51 -1556 52 -1555
rect 107 -1556 108 -1555
rect 121 -1556 122 -1555
rect 243 -1556 244 -1555
rect 261 -1556 262 -1555
rect 285 -1556 286 -1555
rect 289 -1556 290 -1555
rect 345 -1556 346 -1555
rect 359 -1556 360 -1555
rect 387 -1556 388 -1555
rect 415 -1556 416 -1555
rect 436 -1556 437 -1555
rect 450 -1556 451 -1555
rect 471 -1556 472 -1555
rect 485 -1556 486 -1555
rect 520 -1556 521 -1555
rect 586 -1556 587 -1555
rect 590 -1556 591 -1555
rect 72 -1558 73 -1557
rect 79 -1558 80 -1557
rect 86 -1558 87 -1557
rect 222 -1558 223 -1557
rect 226 -1558 227 -1557
rect 233 -1558 234 -1557
rect 236 -1558 237 -1557
rect 247 -1558 248 -1557
rect 261 -1558 262 -1557
rect 268 -1558 269 -1557
rect 271 -1558 272 -1557
rect 359 -1558 360 -1557
rect 380 -1558 381 -1557
rect 492 -1558 493 -1557
rect 75 -1560 76 -1559
rect 79 -1560 80 -1559
rect 96 -1560 97 -1559
rect 366 -1560 367 -1559
rect 422 -1560 423 -1559
rect 502 -1560 503 -1559
rect 103 -1562 104 -1561
rect 114 -1562 115 -1561
rect 128 -1562 129 -1561
rect 327 -1562 328 -1561
rect 429 -1562 430 -1561
rect 499 -1562 500 -1561
rect 149 -1564 150 -1563
rect 177 -1564 178 -1563
rect 194 -1564 195 -1563
rect 296 -1564 297 -1563
rect 310 -1564 311 -1563
rect 369 -1564 370 -1563
rect 429 -1564 430 -1563
rect 464 -1564 465 -1563
rect 492 -1564 493 -1563
rect 506 -1564 507 -1563
rect 142 -1566 143 -1565
rect 194 -1566 195 -1565
rect 198 -1566 199 -1565
rect 222 -1566 223 -1565
rect 240 -1566 241 -1565
rect 338 -1566 339 -1565
rect 369 -1566 370 -1565
rect 394 -1566 395 -1565
rect 436 -1566 437 -1565
rect 443 -1566 444 -1565
rect 457 -1566 458 -1565
rect 464 -1566 465 -1565
rect 142 -1568 143 -1567
rect 191 -1568 192 -1567
rect 205 -1568 206 -1567
rect 229 -1568 230 -1567
rect 247 -1568 248 -1567
rect 313 -1568 314 -1567
rect 317 -1568 318 -1567
rect 390 -1568 391 -1567
rect 128 -1570 129 -1569
rect 191 -1570 192 -1569
rect 219 -1570 220 -1569
rect 254 -1570 255 -1569
rect 275 -1570 276 -1569
rect 296 -1570 297 -1569
rect 317 -1570 318 -1569
rect 478 -1570 479 -1569
rect 159 -1572 160 -1571
rect 212 -1572 213 -1571
rect 254 -1572 255 -1571
rect 282 -1572 283 -1571
rect 292 -1572 293 -1571
rect 527 -1572 528 -1571
rect 65 -1574 66 -1573
rect 159 -1574 160 -1573
rect 163 -1574 164 -1573
rect 170 -1574 171 -1573
rect 173 -1574 174 -1573
rect 201 -1574 202 -1573
rect 275 -1574 276 -1573
rect 366 -1574 367 -1573
rect 373 -1574 374 -1573
rect 394 -1574 395 -1573
rect 135 -1576 136 -1575
rect 212 -1576 213 -1575
rect 324 -1576 325 -1575
rect 380 -1576 381 -1575
rect 135 -1578 136 -1577
rect 152 -1578 153 -1577
rect 163 -1578 164 -1577
rect 184 -1578 185 -1577
rect 373 -1578 374 -1577
rect 408 -1578 409 -1577
rect 152 -1580 153 -1579
rect 177 -1580 178 -1579
rect 156 -1582 157 -1581
rect 184 -1582 185 -1581
rect 72 -1593 73 -1592
rect 82 -1593 83 -1592
rect 89 -1593 90 -1592
rect 93 -1593 94 -1592
rect 128 -1593 129 -1592
rect 156 -1593 157 -1592
rect 163 -1593 164 -1592
rect 205 -1593 206 -1592
rect 219 -1593 220 -1592
rect 240 -1593 241 -1592
rect 243 -1593 244 -1592
rect 261 -1593 262 -1592
rect 282 -1593 283 -1592
rect 289 -1593 290 -1592
rect 296 -1593 297 -1592
rect 310 -1593 311 -1592
rect 320 -1593 321 -1592
rect 338 -1593 339 -1592
rect 345 -1593 346 -1592
rect 352 -1593 353 -1592
rect 366 -1593 367 -1592
rect 373 -1593 374 -1592
rect 383 -1593 384 -1592
rect 429 -1593 430 -1592
rect 471 -1593 472 -1592
rect 485 -1593 486 -1592
rect 506 -1593 507 -1592
rect 513 -1593 514 -1592
rect 75 -1595 76 -1594
rect 79 -1595 80 -1594
rect 135 -1595 136 -1594
rect 152 -1595 153 -1594
rect 163 -1595 164 -1594
rect 194 -1595 195 -1594
rect 205 -1595 206 -1594
rect 247 -1595 248 -1594
rect 254 -1595 255 -1594
rect 369 -1595 370 -1594
rect 422 -1595 423 -1594
rect 436 -1595 437 -1594
rect 443 -1595 444 -1594
rect 485 -1595 486 -1594
rect 114 -1597 115 -1596
rect 152 -1597 153 -1596
rect 177 -1597 178 -1596
rect 268 -1597 269 -1596
rect 275 -1597 276 -1596
rect 289 -1597 290 -1596
rect 317 -1597 318 -1596
rect 345 -1597 346 -1596
rect 352 -1597 353 -1596
rect 380 -1597 381 -1596
rect 464 -1597 465 -1596
rect 471 -1597 472 -1596
rect 131 -1599 132 -1598
rect 135 -1599 136 -1598
rect 142 -1599 143 -1598
rect 145 -1599 146 -1598
rect 156 -1599 157 -1598
rect 275 -1599 276 -1598
rect 282 -1599 283 -1598
rect 310 -1599 311 -1598
rect 317 -1599 318 -1598
rect 359 -1599 360 -1598
rect 184 -1601 185 -1600
rect 215 -1601 216 -1600
rect 226 -1601 227 -1600
rect 324 -1601 325 -1600
rect 331 -1601 332 -1600
rect 334 -1601 335 -1600
rect 338 -1601 339 -1600
rect 401 -1601 402 -1600
rect 191 -1603 192 -1602
rect 201 -1603 202 -1602
rect 212 -1603 213 -1602
rect 296 -1603 297 -1602
rect 299 -1603 300 -1602
rect 359 -1603 360 -1602
rect 191 -1605 192 -1604
rect 208 -1605 209 -1604
rect 226 -1605 227 -1604
rect 341 -1605 342 -1604
rect 233 -1607 234 -1606
rect 254 -1607 255 -1606
rect 261 -1607 262 -1606
rect 303 -1607 304 -1606
rect 236 -1609 237 -1608
rect 278 -1609 279 -1608
rect 240 -1611 241 -1610
rect 268 -1611 269 -1610
rect 243 -1613 244 -1612
rect 324 -1613 325 -1612
rect 250 -1615 251 -1614
rect 303 -1615 304 -1614
rect 30 -1626 31 -1625
rect 33 -1626 34 -1625
rect 37 -1626 38 -1625
rect 180 -1626 181 -1625
rect 198 -1626 199 -1625
rect 215 -1626 216 -1625
rect 233 -1626 234 -1625
rect 236 -1626 237 -1625
rect 240 -1626 241 -1625
rect 271 -1626 272 -1625
rect 275 -1626 276 -1625
rect 317 -1626 318 -1625
rect 334 -1626 335 -1625
rect 366 -1626 367 -1625
rect 401 -1626 402 -1625
rect 443 -1626 444 -1625
rect 467 -1626 468 -1625
rect 471 -1626 472 -1625
rect 488 -1626 489 -1625
rect 492 -1626 493 -1625
rect 44 -1628 45 -1627
rect 156 -1628 157 -1627
rect 177 -1628 178 -1627
rect 219 -1628 220 -1627
rect 254 -1628 255 -1627
rect 257 -1628 258 -1627
rect 261 -1628 262 -1627
rect 352 -1628 353 -1627
rect 359 -1628 360 -1627
rect 380 -1628 381 -1627
rect 51 -1630 52 -1629
rect 86 -1630 87 -1629
rect 93 -1630 94 -1629
rect 100 -1630 101 -1629
rect 121 -1630 122 -1629
rect 142 -1630 143 -1629
rect 149 -1630 150 -1629
rect 163 -1630 164 -1629
rect 177 -1630 178 -1629
rect 201 -1630 202 -1629
rect 212 -1630 213 -1629
rect 247 -1630 248 -1629
rect 254 -1630 255 -1629
rect 289 -1630 290 -1629
rect 296 -1630 297 -1629
rect 324 -1630 325 -1629
rect 327 -1630 328 -1629
rect 352 -1630 353 -1629
rect 65 -1632 66 -1631
rect 110 -1632 111 -1631
rect 124 -1632 125 -1631
rect 135 -1632 136 -1631
rect 138 -1632 139 -1631
rect 170 -1632 171 -1631
rect 191 -1632 192 -1631
rect 240 -1632 241 -1631
rect 257 -1632 258 -1631
rect 289 -1632 290 -1631
rect 303 -1632 304 -1631
rect 359 -1632 360 -1631
rect 72 -1634 73 -1633
rect 89 -1634 90 -1633
rect 100 -1634 101 -1633
rect 124 -1634 125 -1633
rect 135 -1634 136 -1633
rect 156 -1634 157 -1633
rect 163 -1634 164 -1633
rect 226 -1634 227 -1633
rect 264 -1634 265 -1633
rect 317 -1634 318 -1633
rect 345 -1634 346 -1633
rect 366 -1634 367 -1633
rect 72 -1636 73 -1635
rect 131 -1636 132 -1635
rect 170 -1636 171 -1635
rect 229 -1636 230 -1635
rect 275 -1636 276 -1635
rect 338 -1636 339 -1635
rect 345 -1636 346 -1635
rect 404 -1636 405 -1635
rect 79 -1638 80 -1637
rect 114 -1638 115 -1637
rect 198 -1638 199 -1637
rect 222 -1638 223 -1637
rect 226 -1638 227 -1637
rect 296 -1638 297 -1637
rect 303 -1638 304 -1637
rect 310 -1638 311 -1637
rect 58 -1640 59 -1639
rect 114 -1640 115 -1639
rect 219 -1640 220 -1639
rect 331 -1640 332 -1639
rect 86 -1642 87 -1641
rect 145 -1642 146 -1641
rect 278 -1642 279 -1641
rect 373 -1642 374 -1641
rect 107 -1644 108 -1643
rect 149 -1644 150 -1643
rect 282 -1644 283 -1643
rect 310 -1644 311 -1643
rect 19 -1655 20 -1654
rect 23 -1655 24 -1654
rect 37 -1655 38 -1654
rect 222 -1655 223 -1654
rect 226 -1655 227 -1654
rect 366 -1655 367 -1654
rect 387 -1655 388 -1654
rect 390 -1655 391 -1654
rect 44 -1657 45 -1656
rect 128 -1657 129 -1656
rect 149 -1657 150 -1656
rect 215 -1657 216 -1656
rect 219 -1657 220 -1656
rect 240 -1657 241 -1656
rect 243 -1657 244 -1656
rect 261 -1657 262 -1656
rect 268 -1657 269 -1656
rect 310 -1657 311 -1656
rect 317 -1657 318 -1656
rect 401 -1657 402 -1656
rect 51 -1659 52 -1658
rect 138 -1659 139 -1658
rect 163 -1659 164 -1658
rect 184 -1659 185 -1658
rect 191 -1659 192 -1658
rect 198 -1659 199 -1658
rect 212 -1659 213 -1658
rect 289 -1659 290 -1658
rect 296 -1659 297 -1658
rect 310 -1659 311 -1658
rect 324 -1659 325 -1658
rect 373 -1659 374 -1658
rect 65 -1661 66 -1660
rect 93 -1661 94 -1660
rect 100 -1661 101 -1660
rect 135 -1661 136 -1660
rect 156 -1661 157 -1660
rect 163 -1661 164 -1660
rect 212 -1661 213 -1660
rect 296 -1661 297 -1660
rect 331 -1661 332 -1660
rect 373 -1661 374 -1660
rect 72 -1663 73 -1662
rect 96 -1663 97 -1662
rect 103 -1663 104 -1662
rect 107 -1663 108 -1662
rect 117 -1663 118 -1662
rect 191 -1663 192 -1662
rect 226 -1663 227 -1662
rect 324 -1663 325 -1662
rect 331 -1663 332 -1662
rect 345 -1663 346 -1662
rect 366 -1663 367 -1662
rect 380 -1663 381 -1662
rect 79 -1665 80 -1664
rect 124 -1665 125 -1664
rect 156 -1665 157 -1664
rect 170 -1665 171 -1664
rect 222 -1665 223 -1664
rect 380 -1665 381 -1664
rect 86 -1667 87 -1666
rect 114 -1667 115 -1666
rect 121 -1667 122 -1666
rect 145 -1667 146 -1666
rect 229 -1667 230 -1666
rect 320 -1667 321 -1666
rect 338 -1667 339 -1666
rect 394 -1667 395 -1666
rect 121 -1669 122 -1668
rect 177 -1669 178 -1668
rect 205 -1669 206 -1668
rect 394 -1669 395 -1668
rect 145 -1671 146 -1670
rect 149 -1671 150 -1670
rect 205 -1671 206 -1670
rect 271 -1671 272 -1670
rect 282 -1671 283 -1670
rect 352 -1671 353 -1670
rect 233 -1673 234 -1672
rect 247 -1673 248 -1672
rect 254 -1673 255 -1672
rect 268 -1673 269 -1672
rect 285 -1673 286 -1672
rect 338 -1673 339 -1672
rect 348 -1673 349 -1672
rect 352 -1673 353 -1672
rect 208 -1675 209 -1674
rect 247 -1675 248 -1674
rect 261 -1675 262 -1674
rect 303 -1675 304 -1674
rect 236 -1677 237 -1676
rect 359 -1677 360 -1676
rect 240 -1679 241 -1678
rect 275 -1679 276 -1678
rect 2 -1690 3 -1689
rect 9 -1690 10 -1689
rect 16 -1690 17 -1689
rect 23 -1690 24 -1689
rect 30 -1690 31 -1689
rect 33 -1690 34 -1689
rect 89 -1690 90 -1689
rect 96 -1690 97 -1689
rect 100 -1690 101 -1689
rect 107 -1690 108 -1689
rect 114 -1690 115 -1689
rect 205 -1690 206 -1689
rect 222 -1690 223 -1689
rect 243 -1690 244 -1689
rect 254 -1690 255 -1689
rect 401 -1690 402 -1689
rect 121 -1692 122 -1691
rect 212 -1692 213 -1691
rect 226 -1692 227 -1691
rect 233 -1692 234 -1691
rect 257 -1692 258 -1691
rect 296 -1692 297 -1691
rect 317 -1692 318 -1691
rect 331 -1692 332 -1691
rect 359 -1692 360 -1691
rect 373 -1692 374 -1691
rect 121 -1694 122 -1693
rect 128 -1694 129 -1693
rect 156 -1694 157 -1693
rect 184 -1694 185 -1693
rect 191 -1694 192 -1693
rect 247 -1694 248 -1693
rect 264 -1694 265 -1693
rect 310 -1694 311 -1693
rect 135 -1696 136 -1695
rect 156 -1696 157 -1695
rect 163 -1696 164 -1695
rect 170 -1696 171 -1695
rect 194 -1696 195 -1695
rect 205 -1696 206 -1695
rect 226 -1696 227 -1695
rect 324 -1696 325 -1695
rect 131 -1698 132 -1697
rect 135 -1698 136 -1697
rect 149 -1698 150 -1697
rect 163 -1698 164 -1697
rect 170 -1698 171 -1697
rect 177 -1698 178 -1697
rect 198 -1698 199 -1697
rect 219 -1698 220 -1697
rect 229 -1698 230 -1697
rect 233 -1698 234 -1697
rect 268 -1698 269 -1697
rect 285 -1698 286 -1697
rect 292 -1698 293 -1697
rect 380 -1698 381 -1697
rect 117 -1700 118 -1699
rect 131 -1700 132 -1699
rect 173 -1700 174 -1699
rect 177 -1700 178 -1699
rect 201 -1700 202 -1699
rect 212 -1700 213 -1699
rect 275 -1700 276 -1699
rect 278 -1700 279 -1699
rect 285 -1700 286 -1699
rect 289 -1700 290 -1699
rect 296 -1700 297 -1699
rect 394 -1700 395 -1699
rect 303 -1702 304 -1701
rect 310 -1702 311 -1701
rect 324 -1702 325 -1701
rect 338 -1702 339 -1701
rect 5 -1713 6 -1712
rect 9 -1713 10 -1712
rect 128 -1713 129 -1712
rect 135 -1713 136 -1712
rect 142 -1713 143 -1712
rect 163 -1713 164 -1712
rect 170 -1713 171 -1712
rect 201 -1713 202 -1712
rect 212 -1713 213 -1712
rect 219 -1713 220 -1712
rect 233 -1713 234 -1712
rect 243 -1713 244 -1712
rect 303 -1713 304 -1712
rect 310 -1713 311 -1712
rect 317 -1713 318 -1712
rect 324 -1713 325 -1712
rect 152 -1715 153 -1714
rect 156 -1715 157 -1714
rect 177 -1715 178 -1714
rect 226 -1715 227 -1714
rect 187 -1717 188 -1716
rect 205 -1717 206 -1716
<< metal2 >>
rect 177 -3 178 1
rect 187 -3 188 1
rect 198 -3 199 1
rect 205 -3 206 1
rect 208 -3 209 1
rect 222 -3 223 1
rect 240 -3 241 1
rect 247 -3 248 1
rect 275 -3 276 1
rect 282 -3 283 1
rect 289 -3 290 1
rect 299 -3 300 1
rect 215 -3 216 -1
rect 233 -3 234 -1
rect 243 -3 244 -1
rect 254 -3 255 -1
rect 107 -13 108 -11
rect 110 -13 111 -11
rect 142 -22 143 -12
rect 170 -22 171 -12
rect 177 -13 178 -11
rect 194 -13 195 -11
rect 219 -13 220 -11
rect 233 -13 234 -11
rect 254 -13 255 -11
rect 268 -22 269 -12
rect 289 -13 290 -11
rect 303 -13 304 -11
rect 149 -22 150 -14
rect 159 -22 160 -14
rect 163 -22 164 -14
rect 194 -22 195 -14
rect 208 -15 209 -11
rect 219 -22 220 -14
rect 226 -15 227 -11
rect 247 -15 248 -11
rect 264 -22 265 -14
rect 275 -22 276 -14
rect 282 -15 283 -11
rect 289 -22 290 -14
rect 292 -22 293 -14
rect 310 -22 311 -14
rect 184 -22 185 -16
rect 208 -22 209 -16
rect 240 -22 241 -16
rect 247 -22 248 -16
rect 296 -22 297 -16
rect 299 -17 300 -11
rect 191 -19 192 -11
rect 198 -19 199 -11
rect 198 -22 199 -20
rect 215 -21 216 -11
rect 135 -35 136 -31
rect 145 -35 146 -31
rect 149 -32 150 -30
rect 149 -35 150 -31
rect 149 -32 150 -30
rect 149 -35 150 -31
rect 152 -35 153 -31
rect 156 -35 157 -31
rect 177 -32 178 -30
rect 226 -35 227 -31
rect 233 -35 234 -31
rect 243 -35 244 -31
rect 247 -35 248 -31
rect 261 -35 262 -31
rect 275 -32 276 -30
rect 275 -35 276 -31
rect 275 -32 276 -30
rect 275 -35 276 -31
rect 282 -35 283 -31
rect 292 -35 293 -31
rect 296 -32 297 -30
rect 303 -32 304 -30
rect 310 -32 311 -30
rect 324 -35 325 -31
rect 478 -35 479 -31
rect 485 -35 486 -31
rect 579 -35 580 -31
rect 583 -35 584 -31
rect 142 -34 143 -30
rect 180 -34 181 -30
rect 184 -34 185 -30
rect 184 -35 185 -33
rect 184 -34 185 -30
rect 184 -35 185 -33
rect 191 -34 192 -30
rect 198 -34 199 -30
rect 212 -34 213 -30
rect 219 -34 220 -30
rect 240 -34 241 -30
rect 254 -35 255 -33
rect 257 -34 258 -30
rect 268 -34 269 -30
rect 285 -34 286 -30
rect 289 -34 290 -30
rect 296 -35 297 -33
rect 303 -35 304 -33
rect 317 -35 318 -33
rect 320 -34 321 -30
rect 79 -58 80 -44
rect 82 -45 83 -43
rect 135 -45 136 -43
rect 152 -45 153 -43
rect 156 -45 157 -43
rect 156 -58 157 -44
rect 156 -45 157 -43
rect 156 -58 157 -44
rect 170 -58 171 -44
rect 173 -45 174 -43
rect 184 -45 185 -43
rect 194 -45 195 -43
rect 212 -45 213 -43
rect 215 -58 216 -44
rect 219 -58 220 -44
rect 233 -45 234 -43
rect 240 -58 241 -44
rect 282 -45 283 -43
rect 289 -58 290 -44
rect 320 -58 321 -44
rect 338 -58 339 -44
rect 345 -58 346 -44
rect 352 -58 353 -44
rect 362 -58 363 -44
rect 467 -58 468 -44
rect 471 -58 472 -44
rect 478 -58 479 -44
rect 485 -45 486 -43
rect 576 -58 577 -44
rect 583 -45 584 -43
rect 149 -47 150 -43
rect 149 -58 150 -46
rect 149 -47 150 -43
rect 149 -58 150 -46
rect 177 -58 178 -46
rect 194 -58 195 -46
rect 212 -58 213 -46
rect 243 -58 244 -46
rect 247 -47 248 -43
rect 268 -47 269 -43
rect 292 -47 293 -43
rect 317 -47 318 -43
rect 184 -58 185 -48
rect 205 -58 206 -48
rect 222 -49 223 -43
rect 226 -58 227 -48
rect 233 -58 234 -48
rect 261 -49 262 -43
rect 296 -49 297 -43
rect 296 -58 297 -48
rect 296 -49 297 -43
rect 296 -58 297 -48
rect 310 -49 311 -43
rect 324 -49 325 -43
rect 229 -51 230 -43
rect 261 -58 262 -50
rect 317 -58 318 -50
rect 341 -58 342 -50
rect 247 -58 248 -52
rect 268 -58 269 -52
rect 324 -58 325 -52
rect 334 -53 335 -43
rect 250 -55 251 -43
rect 275 -55 276 -43
rect 254 -57 255 -43
rect 254 -58 255 -56
rect 254 -57 255 -43
rect 254 -58 255 -56
rect 275 -58 276 -56
rect 282 -58 283 -56
rect 142 -68 143 -66
rect 149 -68 150 -66
rect 170 -68 171 -66
rect 170 -81 171 -67
rect 170 -68 171 -66
rect 170 -81 171 -67
rect 177 -68 178 -66
rect 177 -81 178 -67
rect 177 -68 178 -66
rect 177 -81 178 -67
rect 198 -68 199 -66
rect 198 -81 199 -67
rect 198 -68 199 -66
rect 198 -81 199 -67
rect 205 -68 206 -66
rect 212 -81 213 -67
rect 219 -68 220 -66
rect 243 -81 244 -67
rect 247 -68 248 -66
rect 261 -68 262 -66
rect 268 -68 269 -66
rect 282 -81 283 -67
rect 324 -68 325 -66
rect 324 -81 325 -67
rect 324 -68 325 -66
rect 324 -81 325 -67
rect 338 -81 339 -67
rect 345 -68 346 -66
rect 471 -68 472 -66
rect 471 -81 472 -67
rect 471 -68 472 -66
rect 471 -81 472 -67
rect 474 -81 475 -67
rect 485 -81 486 -67
rect 576 -68 577 -66
rect 576 -81 577 -67
rect 576 -68 577 -66
rect 576 -81 577 -67
rect 138 -81 139 -69
rect 219 -81 220 -69
rect 226 -70 227 -66
rect 233 -81 234 -69
rect 240 -70 241 -66
rect 289 -70 290 -66
rect 345 -81 346 -69
rect 352 -70 353 -66
rect 478 -70 479 -66
rect 478 -81 479 -69
rect 478 -70 479 -66
rect 478 -81 479 -69
rect 142 -81 143 -71
rect 163 -81 164 -71
rect 166 -81 167 -71
rect 205 -81 206 -71
rect 226 -81 227 -71
rect 275 -72 276 -66
rect 278 -81 279 -71
rect 296 -72 297 -66
rect 320 -72 321 -66
rect 352 -81 353 -71
rect 149 -81 150 -73
rect 156 -74 157 -66
rect 236 -74 237 -66
rect 289 -81 290 -73
rect 296 -81 297 -73
rect 303 -81 304 -73
rect 247 -81 248 -75
rect 254 -76 255 -66
rect 261 -81 262 -75
rect 310 -76 311 -66
rect 240 -81 241 -77
rect 254 -81 255 -77
rect 268 -81 269 -77
rect 306 -78 307 -66
rect 275 -81 276 -79
rect 317 -81 318 -79
rect 121 -91 122 -89
rect 121 -112 122 -90
rect 121 -91 122 -89
rect 121 -112 122 -90
rect 128 -112 129 -90
rect 135 -112 136 -90
rect 142 -91 143 -89
rect 145 -112 146 -90
rect 149 -91 150 -89
rect 159 -91 160 -89
rect 163 -112 164 -90
rect 226 -91 227 -89
rect 233 -91 234 -89
rect 268 -112 269 -90
rect 271 -91 272 -89
rect 359 -112 360 -90
rect 397 -112 398 -90
rect 422 -112 423 -90
rect 481 -112 482 -90
rect 485 -91 486 -89
rect 576 -91 577 -89
rect 583 -112 584 -90
rect 107 -112 108 -92
rect 142 -112 143 -92
rect 152 -112 153 -92
rect 156 -112 157 -92
rect 166 -93 167 -89
rect 170 -93 171 -89
rect 177 -93 178 -89
rect 184 -112 185 -92
rect 187 -93 188 -89
rect 198 -112 199 -92
rect 205 -93 206 -89
rect 243 -93 244 -89
rect 257 -112 258 -92
rect 261 -93 262 -89
rect 289 -112 290 -92
rect 324 -93 325 -89
rect 338 -93 339 -89
rect 348 -93 349 -89
rect 352 -93 353 -89
rect 380 -112 381 -92
rect 478 -93 479 -89
rect 485 -112 486 -92
rect 576 -112 577 -92
rect 590 -112 591 -92
rect 191 -112 192 -94
rect 201 -95 202 -89
rect 219 -95 220 -89
rect 303 -112 304 -94
rect 310 -95 311 -89
rect 366 -112 367 -94
rect 478 -112 479 -94
rect 492 -112 493 -94
rect 194 -97 195 -89
rect 226 -112 227 -96
rect 240 -97 241 -89
rect 317 -97 318 -89
rect 341 -112 342 -96
rect 345 -97 346 -89
rect 212 -99 213 -89
rect 219 -112 220 -98
rect 222 -112 223 -98
rect 352 -112 353 -98
rect 212 -112 213 -100
rect 233 -112 234 -100
rect 243 -112 244 -100
rect 247 -101 248 -89
rect 250 -112 251 -100
rect 324 -112 325 -100
rect 338 -112 339 -100
rect 345 -112 346 -100
rect 254 -103 255 -89
rect 261 -112 262 -102
rect 275 -112 276 -102
rect 310 -112 311 -102
rect 317 -112 318 -102
rect 373 -112 374 -102
rect 254 -112 255 -104
rect 320 -112 321 -104
rect 296 -107 297 -89
rect 331 -112 332 -106
rect 282 -109 283 -89
rect 296 -112 297 -108
rect 180 -112 181 -110
rect 282 -112 283 -110
rect 65 -151 66 -121
rect 107 -122 108 -120
rect 131 -151 132 -121
rect 135 -122 136 -120
rect 145 -122 146 -120
rect 170 -122 171 -120
rect 173 -122 174 -120
rect 184 -122 185 -120
rect 191 -122 192 -120
rect 205 -122 206 -120
rect 208 -122 209 -120
rect 254 -151 255 -121
rect 264 -151 265 -121
rect 278 -122 279 -120
rect 289 -122 290 -120
rect 317 -151 318 -121
rect 324 -122 325 -120
rect 338 -151 339 -121
rect 345 -122 346 -120
rect 345 -151 346 -121
rect 345 -122 346 -120
rect 345 -151 346 -121
rect 359 -122 360 -120
rect 415 -151 416 -121
rect 422 -122 423 -120
rect 443 -151 444 -121
rect 478 -122 479 -120
rect 485 -122 486 -120
rect 492 -122 493 -120
rect 499 -151 500 -121
rect 576 -122 577 -120
rect 583 -122 584 -120
rect 590 -122 591 -120
rect 590 -151 591 -121
rect 590 -122 591 -120
rect 590 -151 591 -121
rect 72 -151 73 -123
rect 100 -151 101 -123
rect 107 -151 108 -123
rect 114 -151 115 -123
rect 128 -151 129 -123
rect 135 -151 136 -123
rect 149 -151 150 -123
rect 156 -124 157 -120
rect 163 -124 164 -120
rect 236 -151 237 -123
rect 243 -124 244 -120
rect 310 -124 311 -120
rect 331 -124 332 -120
rect 422 -151 423 -123
rect 86 -151 87 -125
rect 124 -126 125 -120
rect 170 -151 171 -125
rect 208 -151 209 -125
rect 219 -126 220 -120
rect 366 -126 367 -120
rect 380 -126 381 -120
rect 429 -151 430 -125
rect 93 -151 94 -127
rect 243 -151 244 -127
rect 275 -128 276 -120
rect 373 -128 374 -120
rect 387 -151 388 -127
rect 436 -151 437 -127
rect 156 -151 157 -129
rect 219 -151 220 -129
rect 222 -130 223 -120
rect 233 -130 234 -120
rect 282 -130 283 -120
rect 310 -151 311 -129
rect 334 -151 335 -129
rect 366 -151 367 -129
rect 394 -130 395 -120
rect 401 -151 402 -129
rect 177 -151 178 -131
rect 285 -151 286 -131
rect 299 -151 300 -131
rect 359 -151 360 -131
rect 184 -151 185 -133
rect 233 -151 234 -133
rect 303 -134 304 -120
rect 373 -151 374 -133
rect 191 -151 192 -135
rect 226 -136 227 -120
rect 229 -151 230 -135
rect 289 -151 290 -135
rect 352 -136 353 -120
rect 380 -151 381 -135
rect 198 -138 199 -120
rect 212 -151 213 -137
rect 222 -151 223 -137
rect 324 -151 325 -137
rect 352 -151 353 -137
rect 394 -151 395 -137
rect 198 -151 199 -139
rect 261 -140 262 -120
rect 205 -151 206 -141
rect 247 -151 248 -141
rect 261 -151 262 -141
rect 296 -142 297 -120
rect 226 -151 227 -143
rect 268 -144 269 -120
rect 240 -146 241 -120
rect 303 -151 304 -145
rect 240 -151 241 -147
rect 275 -151 276 -147
rect 257 -150 258 -120
rect 268 -151 269 -149
rect 19 -200 20 -160
rect 26 -200 27 -160
rect 65 -161 66 -159
rect 114 -161 115 -159
rect 131 -161 132 -159
rect 159 -200 160 -160
rect 163 -161 164 -159
rect 247 -161 248 -159
rect 264 -161 265 -159
rect 310 -161 311 -159
rect 317 -161 318 -159
rect 331 -161 332 -159
rect 352 -161 353 -159
rect 429 -161 430 -159
rect 499 -161 500 -159
rect 506 -200 507 -160
rect 590 -161 591 -159
rect 590 -200 591 -160
rect 590 -161 591 -159
rect 590 -200 591 -160
rect 72 -163 73 -159
rect 121 -163 122 -159
rect 135 -163 136 -159
rect 135 -200 136 -162
rect 135 -163 136 -159
rect 135 -200 136 -162
rect 149 -163 150 -159
rect 180 -200 181 -162
rect 208 -163 209 -159
rect 415 -163 416 -159
rect 79 -165 80 -159
rect 128 -165 129 -159
rect 149 -200 150 -164
rect 156 -165 157 -159
rect 219 -200 220 -164
rect 310 -200 311 -164
rect 320 -200 321 -164
rect 436 -165 437 -159
rect 79 -200 80 -166
rect 124 -167 125 -159
rect 128 -200 129 -166
rect 184 -167 185 -159
rect 226 -167 227 -159
rect 247 -200 248 -166
rect 268 -167 269 -159
rect 436 -200 437 -166
rect 86 -169 87 -159
rect 166 -169 167 -159
rect 226 -200 227 -168
rect 331 -200 332 -168
rect 345 -169 346 -159
rect 429 -200 430 -168
rect 93 -171 94 -159
rect 145 -171 146 -159
rect 236 -200 237 -170
rect 268 -200 269 -170
rect 278 -200 279 -170
rect 460 -200 461 -170
rect 100 -200 101 -172
rect 177 -173 178 -159
rect 243 -173 244 -159
rect 338 -173 339 -159
rect 352 -200 353 -172
rect 387 -173 388 -159
rect 103 -175 104 -159
rect 142 -175 143 -159
rect 177 -200 178 -174
rect 205 -200 206 -174
rect 212 -175 213 -159
rect 338 -200 339 -174
rect 359 -175 360 -159
rect 415 -200 416 -174
rect 86 -200 87 -176
rect 142 -200 143 -176
rect 212 -200 213 -176
rect 296 -200 297 -176
rect 299 -177 300 -159
rect 422 -177 423 -159
rect 107 -179 108 -159
rect 163 -200 164 -178
rect 282 -200 283 -178
rect 317 -200 318 -178
rect 324 -179 325 -159
rect 345 -200 346 -178
rect 366 -179 367 -159
rect 366 -200 367 -178
rect 366 -179 367 -159
rect 366 -200 367 -178
rect 373 -179 374 -159
rect 464 -200 465 -178
rect 107 -200 108 -180
rect 198 -181 199 -159
rect 254 -181 255 -159
rect 324 -200 325 -180
rect 373 -200 374 -180
rect 408 -181 409 -159
rect 422 -200 423 -180
rect 443 -181 444 -159
rect 114 -200 115 -182
rect 170 -183 171 -159
rect 191 -183 192 -159
rect 254 -200 255 -182
rect 299 -200 300 -182
rect 387 -200 388 -182
rect 401 -183 402 -159
rect 408 -200 409 -182
rect 93 -200 94 -184
rect 170 -200 171 -184
rect 243 -200 244 -184
rect 443 -200 444 -184
rect 121 -200 122 -186
rect 156 -200 157 -186
rect 303 -187 304 -159
rect 359 -200 360 -186
rect 394 -187 395 -159
rect 401 -200 402 -186
rect 191 -200 192 -188
rect 303 -200 304 -188
rect 380 -189 381 -159
rect 394 -200 395 -188
rect 261 -191 262 -159
rect 380 -200 381 -190
rect 240 -193 241 -159
rect 261 -200 262 -192
rect 240 -200 241 -194
rect 275 -195 276 -159
rect 275 -200 276 -196
rect 289 -197 290 -159
rect 233 -199 234 -159
rect 289 -200 290 -198
rect 12 -210 13 -208
rect 12 -241 13 -209
rect 12 -210 13 -208
rect 12 -241 13 -209
rect 79 -210 80 -208
rect 222 -210 223 -208
rect 243 -210 244 -208
rect 324 -210 325 -208
rect 348 -241 349 -209
rect 415 -210 416 -208
rect 443 -210 444 -208
rect 453 -210 454 -208
rect 506 -210 507 -208
rect 509 -241 510 -209
rect 562 -241 563 -209
rect 572 -241 573 -209
rect 590 -210 591 -208
rect 590 -241 591 -209
rect 590 -210 591 -208
rect 590 -241 591 -209
rect 86 -212 87 -208
rect 215 -212 216 -208
rect 219 -212 220 -208
rect 338 -212 339 -208
rect 380 -212 381 -208
rect 422 -241 423 -211
rect 450 -241 451 -211
rect 460 -241 461 -211
rect 100 -214 101 -208
rect 240 -214 241 -208
rect 268 -214 269 -208
rect 268 -241 269 -213
rect 268 -214 269 -208
rect 268 -241 269 -213
rect 278 -214 279 -208
rect 436 -214 437 -208
rect 107 -216 108 -208
rect 236 -216 237 -208
rect 240 -241 241 -215
rect 254 -216 255 -208
rect 296 -216 297 -208
rect 373 -216 374 -208
rect 383 -241 384 -215
rect 394 -216 395 -208
rect 401 -216 402 -208
rect 401 -241 402 -215
rect 401 -216 402 -208
rect 401 -241 402 -215
rect 408 -216 409 -208
rect 408 -241 409 -215
rect 408 -216 409 -208
rect 408 -241 409 -215
rect 114 -218 115 -208
rect 191 -218 192 -208
rect 222 -241 223 -217
rect 464 -218 465 -208
rect 114 -241 115 -219
rect 201 -220 202 -208
rect 236 -241 237 -219
rect 282 -220 283 -208
rect 317 -220 318 -208
rect 352 -220 353 -208
rect 359 -220 360 -208
rect 373 -241 374 -219
rect 128 -222 129 -208
rect 198 -222 199 -208
rect 212 -222 213 -208
rect 317 -241 318 -221
rect 320 -241 321 -221
rect 415 -241 416 -221
rect 135 -224 136 -208
rect 145 -224 146 -208
rect 149 -224 150 -208
rect 149 -241 150 -223
rect 149 -224 150 -208
rect 149 -241 150 -223
rect 156 -224 157 -208
rect 226 -224 227 -208
rect 243 -241 244 -223
rect 436 -241 437 -223
rect 128 -241 129 -225
rect 156 -241 157 -225
rect 163 -241 164 -225
rect 275 -226 276 -208
rect 282 -241 283 -225
rect 303 -226 304 -208
rect 324 -241 325 -225
rect 345 -226 346 -208
rect 135 -241 136 -227
rect 166 -228 167 -208
rect 173 -228 174 -208
rect 264 -241 265 -227
rect 289 -241 290 -227
rect 303 -241 304 -227
rect 331 -228 332 -208
rect 443 -241 444 -227
rect 142 -241 143 -229
rect 184 -230 185 -208
rect 191 -241 192 -229
rect 247 -230 248 -208
rect 254 -241 255 -229
rect 261 -230 262 -208
rect 292 -230 293 -208
rect 331 -241 332 -229
rect 338 -241 339 -229
rect 366 -230 367 -208
rect 177 -241 178 -231
rect 215 -241 216 -231
rect 226 -241 227 -231
rect 247 -241 248 -231
rect 261 -241 262 -231
rect 394 -241 395 -231
rect 184 -241 185 -233
rect 205 -234 206 -208
rect 212 -241 213 -233
rect 292 -241 293 -233
rect 296 -241 297 -233
rect 359 -241 360 -233
rect 198 -241 199 -235
rect 310 -236 311 -208
rect 345 -241 346 -235
rect 429 -236 430 -208
rect 278 -241 279 -237
rect 310 -241 311 -237
rect 352 -241 353 -237
rect 366 -241 367 -237
rect 387 -238 388 -208
rect 429 -241 430 -237
rect 275 -241 276 -239
rect 387 -241 388 -239
rect 65 -282 66 -250
rect 93 -282 94 -250
rect 107 -282 108 -250
rect 121 -282 122 -250
rect 124 -251 125 -249
rect 159 -251 160 -249
rect 177 -251 178 -249
rect 194 -282 195 -250
rect 198 -251 199 -249
rect 261 -282 262 -250
rect 268 -251 269 -249
rect 268 -282 269 -250
rect 268 -251 269 -249
rect 268 -282 269 -250
rect 292 -282 293 -250
rect 345 -282 346 -250
rect 366 -251 367 -249
rect 401 -251 402 -249
rect 415 -251 416 -249
rect 492 -282 493 -250
rect 502 -282 503 -250
rect 520 -282 521 -250
rect 562 -251 563 -249
rect 562 -282 563 -250
rect 562 -251 563 -249
rect 562 -282 563 -250
rect 590 -251 591 -249
rect 597 -251 598 -249
rect 600 -251 601 -249
rect 611 -282 612 -250
rect 646 -251 647 -249
rect 646 -282 647 -250
rect 646 -251 647 -249
rect 646 -282 647 -250
rect 79 -282 80 -252
rect 317 -253 318 -249
rect 320 -253 321 -249
rect 338 -253 339 -249
rect 422 -253 423 -249
rect 457 -282 458 -252
rect 471 -282 472 -252
rect 499 -282 500 -252
rect 506 -253 507 -249
rect 527 -282 528 -252
rect 86 -282 87 -254
rect 128 -255 129 -249
rect 135 -255 136 -249
rect 289 -282 290 -254
rect 303 -255 304 -249
rect 401 -282 402 -254
rect 429 -255 430 -249
rect 478 -282 479 -254
rect 114 -257 115 -249
rect 327 -282 328 -256
rect 338 -282 339 -256
rect 415 -282 416 -256
rect 443 -257 444 -249
rect 443 -282 444 -256
rect 443 -257 444 -249
rect 443 -282 444 -256
rect 450 -257 451 -249
rect 485 -282 486 -256
rect 114 -282 115 -258
rect 128 -282 129 -258
rect 135 -282 136 -258
rect 170 -259 171 -249
rect 173 -282 174 -258
rect 177 -282 178 -258
rect 184 -259 185 -249
rect 229 -259 230 -249
rect 247 -259 248 -249
rect 247 -282 248 -258
rect 247 -259 248 -249
rect 247 -282 248 -258
rect 254 -259 255 -249
rect 278 -259 279 -249
rect 320 -282 321 -258
rect 408 -259 409 -249
rect 464 -259 465 -249
rect 506 -282 507 -258
rect 142 -261 143 -249
rect 236 -261 237 -249
rect 257 -282 258 -260
rect 324 -261 325 -249
rect 348 -261 349 -249
rect 422 -282 423 -260
rect 436 -261 437 -249
rect 464 -282 465 -260
rect 142 -282 143 -262
rect 184 -282 185 -262
rect 187 -282 188 -262
rect 240 -263 241 -249
rect 324 -282 325 -262
rect 359 -263 360 -249
rect 373 -263 374 -249
rect 429 -282 430 -262
rect 149 -265 150 -249
rect 156 -265 157 -249
rect 163 -265 164 -249
rect 170 -282 171 -264
rect 191 -265 192 -249
rect 243 -265 244 -249
rect 303 -282 304 -264
rect 359 -282 360 -264
rect 380 -265 381 -249
rect 408 -282 409 -264
rect 149 -282 150 -266
rect 205 -282 206 -266
rect 208 -267 209 -249
rect 233 -282 234 -266
rect 236 -282 237 -266
rect 313 -282 314 -266
rect 352 -267 353 -249
rect 373 -282 374 -266
rect 387 -267 388 -249
rect 436 -282 437 -266
rect 156 -282 157 -268
rect 219 -269 220 -249
rect 222 -269 223 -249
rect 310 -269 311 -249
rect 317 -282 318 -268
rect 352 -282 353 -268
rect 394 -269 395 -249
rect 450 -282 451 -268
rect 163 -282 164 -270
rect 243 -282 244 -270
rect 331 -271 332 -249
rect 387 -282 388 -270
rect 201 -282 202 -272
rect 275 -273 276 -249
rect 299 -282 300 -272
rect 331 -282 332 -272
rect 208 -282 209 -274
rect 366 -282 367 -274
rect 219 -282 220 -276
rect 383 -282 384 -276
rect 226 -282 227 -278
rect 282 -279 283 -249
rect 275 -282 276 -280
rect 296 -282 297 -280
rect 75 -292 76 -290
rect 254 -292 255 -290
rect 257 -292 258 -290
rect 317 -331 318 -291
rect 324 -292 325 -290
rect 478 -292 479 -290
rect 516 -331 517 -291
rect 548 -331 549 -291
rect 562 -292 563 -290
rect 562 -331 563 -291
rect 562 -292 563 -290
rect 562 -331 563 -291
rect 604 -331 605 -291
rect 611 -292 612 -290
rect 646 -292 647 -290
rect 653 -331 654 -291
rect 674 -331 675 -291
rect 681 -331 682 -291
rect 79 -294 80 -290
rect 212 -294 213 -290
rect 219 -294 220 -290
rect 296 -331 297 -293
rect 303 -294 304 -290
rect 401 -294 402 -290
rect 425 -331 426 -293
rect 457 -294 458 -290
rect 464 -294 465 -290
rect 478 -331 479 -293
rect 520 -294 521 -290
rect 541 -331 542 -293
rect 649 -331 650 -293
rect 660 -331 661 -293
rect 79 -331 80 -295
rect 107 -296 108 -290
rect 114 -331 115 -295
rect 156 -296 157 -290
rect 170 -331 171 -295
rect 177 -296 178 -290
rect 187 -296 188 -290
rect 194 -296 195 -290
rect 205 -331 206 -295
rect 282 -296 283 -290
rect 289 -296 290 -290
rect 471 -296 472 -290
rect 527 -296 528 -290
rect 544 -331 545 -295
rect 86 -298 87 -290
rect 152 -331 153 -297
rect 212 -331 213 -297
rect 233 -331 234 -297
rect 236 -298 237 -290
rect 369 -331 370 -297
rect 390 -331 391 -297
rect 492 -298 493 -290
rect 506 -298 507 -290
rect 527 -331 528 -297
rect 86 -331 87 -299
rect 142 -300 143 -290
rect 219 -331 220 -299
rect 464 -331 465 -299
rect 485 -300 486 -290
rect 506 -331 507 -299
rect 93 -302 94 -290
rect 173 -302 174 -290
rect 247 -302 248 -290
rect 320 -302 321 -290
rect 324 -331 325 -301
rect 429 -302 430 -290
rect 436 -302 437 -290
rect 534 -331 535 -301
rect 93 -331 94 -303
rect 149 -304 150 -290
rect 247 -331 248 -303
rect 345 -304 346 -290
rect 348 -331 349 -303
rect 387 -304 388 -290
rect 394 -304 395 -290
rect 429 -331 430 -303
rect 100 -331 101 -305
rect 117 -306 118 -290
rect 128 -306 129 -290
rect 142 -331 143 -305
rect 254 -331 255 -305
rect 268 -306 269 -290
rect 275 -306 276 -290
rect 275 -331 276 -305
rect 275 -306 276 -290
rect 275 -331 276 -305
rect 282 -331 283 -305
rect 485 -331 486 -305
rect 103 -308 104 -290
rect 121 -331 122 -307
rect 135 -308 136 -290
rect 198 -308 199 -290
rect 261 -308 262 -290
rect 264 -331 265 -307
rect 289 -331 290 -307
rect 338 -331 339 -307
rect 341 -308 342 -290
rect 443 -308 444 -290
rect 107 -331 108 -309
rect 163 -310 164 -290
rect 198 -331 199 -309
rect 226 -310 227 -290
rect 303 -331 304 -309
rect 422 -310 423 -290
rect 443 -331 444 -309
rect 555 -331 556 -309
rect 128 -331 129 -311
rect 135 -331 136 -311
rect 163 -331 164 -311
rect 177 -331 178 -311
rect 191 -331 192 -311
rect 226 -331 227 -311
rect 313 -331 314 -311
rect 471 -331 472 -311
rect 345 -331 346 -313
rect 450 -314 451 -290
rect 352 -316 353 -290
rect 401 -331 402 -315
rect 408 -316 409 -290
rect 450 -331 451 -315
rect 331 -318 332 -290
rect 352 -331 353 -317
rect 366 -318 367 -290
rect 380 -331 381 -317
rect 408 -331 409 -317
rect 457 -331 458 -317
rect 331 -331 332 -319
rect 387 -331 388 -319
rect 415 -320 416 -290
rect 492 -331 493 -319
rect 240 -322 241 -290
rect 415 -331 416 -321
rect 422 -331 423 -321
rect 499 -331 500 -321
rect 229 -331 230 -323
rect 240 -331 241 -323
rect 366 -331 367 -323
rect 436 -331 437 -323
rect 373 -326 374 -290
rect 394 -331 395 -325
rect 359 -328 360 -290
rect 373 -331 374 -327
rect 359 -331 360 -329
rect 520 -331 521 -329
rect 44 -382 45 -340
rect 334 -382 335 -340
rect 338 -382 339 -340
rect 527 -341 528 -339
rect 541 -341 542 -339
rect 569 -382 570 -340
rect 583 -382 584 -340
rect 604 -341 605 -339
rect 642 -382 643 -340
rect 688 -382 689 -340
rect 51 -382 52 -342
rect 114 -343 115 -339
rect 128 -343 129 -339
rect 142 -343 143 -339
rect 166 -382 167 -342
rect 236 -343 237 -339
rect 243 -382 244 -342
rect 261 -382 262 -342
rect 264 -343 265 -339
rect 625 -382 626 -342
rect 649 -343 650 -339
rect 653 -343 654 -339
rect 660 -343 661 -339
rect 681 -382 682 -342
rect 58 -382 59 -344
rect 289 -345 290 -339
rect 296 -345 297 -339
rect 313 -345 314 -339
rect 341 -345 342 -339
rect 429 -345 430 -339
rect 471 -345 472 -339
rect 513 -382 514 -344
rect 523 -382 524 -344
rect 597 -382 598 -344
rect 667 -382 668 -344
rect 674 -345 675 -339
rect 79 -347 80 -339
rect 219 -347 220 -339
rect 233 -347 234 -339
rect 345 -382 346 -346
rect 359 -347 360 -339
rect 611 -382 612 -346
rect 79 -382 80 -348
rect 170 -349 171 -339
rect 177 -349 178 -339
rect 226 -349 227 -339
rect 233 -382 234 -348
rect 352 -349 353 -339
rect 362 -349 363 -339
rect 534 -349 535 -339
rect 544 -349 545 -339
rect 639 -382 640 -348
rect 86 -351 87 -339
rect 163 -351 164 -339
rect 177 -382 178 -350
rect 215 -382 216 -350
rect 222 -382 223 -350
rect 362 -382 363 -350
rect 366 -351 367 -339
rect 618 -382 619 -350
rect 86 -382 87 -352
rect 247 -353 248 -339
rect 254 -353 255 -339
rect 268 -382 269 -352
rect 275 -353 276 -339
rect 296 -382 297 -352
rect 341 -382 342 -352
rect 527 -382 528 -352
rect 548 -353 549 -339
rect 646 -382 647 -352
rect 93 -355 94 -339
rect 156 -355 157 -339
rect 159 -382 160 -354
rect 254 -382 255 -354
rect 292 -382 293 -354
rect 366 -382 367 -354
rect 380 -355 381 -339
rect 390 -382 391 -354
rect 411 -355 412 -339
rect 436 -355 437 -339
rect 460 -382 461 -354
rect 534 -382 535 -354
rect 558 -355 559 -339
rect 562 -355 563 -339
rect 72 -357 73 -339
rect 156 -382 157 -356
rect 205 -357 206 -339
rect 285 -357 286 -339
rect 327 -357 328 -339
rect 548 -382 549 -356
rect 562 -382 563 -356
rect 653 -382 654 -356
rect 72 -382 73 -358
rect 212 -359 213 -339
rect 236 -382 237 -358
rect 271 -359 272 -339
rect 327 -382 328 -358
rect 408 -382 409 -358
rect 415 -359 416 -339
rect 436 -382 437 -358
rect 471 -382 472 -358
rect 660 -382 661 -358
rect 93 -382 94 -360
rect 100 -361 101 -339
rect 114 -382 115 -360
rect 401 -361 402 -339
rect 415 -382 416 -360
rect 425 -382 426 -360
rect 478 -361 479 -339
rect 541 -382 542 -360
rect 100 -382 101 -362
rect 121 -363 122 -339
rect 128 -382 129 -362
rect 135 -363 136 -339
rect 142 -382 143 -362
rect 229 -382 230 -362
rect 373 -363 374 -339
rect 478 -382 479 -362
rect 485 -363 486 -339
rect 590 -382 591 -362
rect 68 -382 69 -364
rect 135 -382 136 -364
rect 152 -365 153 -339
rect 219 -382 220 -364
rect 380 -382 381 -364
rect 387 -382 388 -364
rect 394 -365 395 -339
rect 401 -382 402 -364
rect 422 -365 423 -339
rect 576 -382 577 -364
rect 107 -367 108 -339
rect 152 -382 153 -366
rect 205 -382 206 -366
rect 240 -367 241 -339
rect 317 -367 318 -339
rect 394 -382 395 -366
rect 422 -382 423 -366
rect 520 -367 521 -339
rect 107 -382 108 -368
rect 247 -382 248 -368
rect 317 -382 318 -368
rect 457 -369 458 -339
rect 492 -369 493 -339
rect 604 -382 605 -368
rect 110 -382 111 -370
rect 373 -382 374 -370
rect 443 -371 444 -339
rect 485 -382 486 -370
rect 499 -371 500 -339
rect 555 -382 556 -370
rect 121 -382 122 -372
rect 191 -373 192 -339
rect 303 -373 304 -339
rect 443 -382 444 -372
rect 450 -373 451 -339
rect 492 -382 493 -372
rect 506 -373 507 -339
rect 632 -382 633 -372
rect 170 -382 171 -374
rect 240 -382 241 -374
rect 303 -382 304 -374
rect 324 -375 325 -339
rect 348 -375 349 -339
rect 499 -382 500 -374
rect 184 -377 185 -339
rect 191 -382 192 -376
rect 310 -382 311 -376
rect 324 -382 325 -376
rect 429 -382 430 -376
rect 450 -382 451 -376
rect 464 -377 465 -339
rect 506 -382 507 -376
rect 184 -382 185 -378
rect 198 -379 199 -339
rect 331 -379 332 -339
rect 464 -382 465 -378
rect 138 -382 139 -380
rect 198 -382 199 -380
rect 282 -382 283 -380
rect 331 -382 332 -380
rect 2 -439 3 -391
rect 180 -439 181 -391
rect 205 -392 206 -390
rect 226 -439 227 -391
rect 233 -439 234 -391
rect 310 -392 311 -390
rect 317 -392 318 -390
rect 352 -392 353 -390
rect 359 -392 360 -390
rect 611 -392 612 -390
rect 628 -439 629 -391
rect 639 -439 640 -391
rect 649 -439 650 -391
rect 681 -392 682 -390
rect 16 -439 17 -393
rect 292 -394 293 -390
rect 303 -394 304 -390
rect 352 -439 353 -393
rect 355 -394 356 -390
rect 359 -439 360 -393
rect 373 -394 374 -390
rect 562 -439 563 -393
rect 597 -394 598 -390
rect 611 -439 612 -393
rect 667 -394 668 -390
rect 674 -394 675 -390
rect 30 -396 31 -390
rect 37 -439 38 -395
rect 44 -396 45 -390
rect 222 -396 223 -390
rect 240 -396 241 -390
rect 464 -396 465 -390
rect 485 -396 486 -390
rect 485 -439 486 -395
rect 485 -396 486 -390
rect 485 -439 486 -395
rect 513 -396 514 -390
rect 513 -439 514 -395
rect 513 -396 514 -390
rect 513 -439 514 -395
rect 527 -396 528 -390
rect 527 -439 528 -395
rect 527 -396 528 -390
rect 527 -439 528 -395
rect 597 -439 598 -395
rect 625 -396 626 -390
rect 667 -439 668 -395
rect 688 -396 689 -390
rect 44 -439 45 -397
rect 397 -439 398 -397
rect 401 -398 402 -390
rect 422 -439 423 -397
rect 436 -398 437 -390
rect 446 -430 447 -397
rect 450 -398 451 -390
rect 646 -398 647 -390
rect 51 -400 52 -390
rect 138 -400 139 -390
rect 149 -439 150 -399
rect 191 -400 192 -390
rect 215 -400 216 -390
rect 394 -400 395 -390
rect 401 -439 402 -399
rect 632 -400 633 -390
rect 51 -439 52 -401
rect 152 -402 153 -390
rect 163 -439 164 -401
rect 184 -402 185 -390
rect 219 -439 220 -401
rect 404 -439 405 -401
rect 436 -439 437 -401
rect 534 -402 535 -390
rect 576 -402 577 -390
rect 632 -439 633 -401
rect 58 -404 59 -390
rect 341 -404 342 -390
rect 373 -439 374 -403
rect 450 -439 451 -403
rect 460 -404 461 -390
rect 548 -404 549 -390
rect 558 -439 559 -403
rect 576 -439 577 -403
rect 583 -404 584 -390
rect 625 -439 626 -403
rect 58 -439 59 -405
rect 212 -406 213 -390
rect 268 -406 269 -390
rect 289 -406 290 -390
rect 317 -439 318 -405
rect 366 -406 367 -390
rect 376 -439 377 -405
rect 415 -406 416 -390
rect 439 -439 440 -405
rect 604 -406 605 -390
rect 65 -439 66 -407
rect 303 -439 304 -407
rect 334 -408 335 -390
rect 590 -408 591 -390
rect 604 -439 605 -407
rect 653 -408 654 -390
rect 72 -410 73 -390
rect 327 -439 328 -409
rect 341 -439 342 -409
rect 478 -410 479 -390
rect 492 -410 493 -390
rect 534 -439 535 -409
rect 569 -410 570 -390
rect 583 -439 584 -409
rect 653 -439 654 -409
rect 663 -439 664 -409
rect 72 -439 73 -411
rect 187 -439 188 -411
rect 254 -412 255 -390
rect 268 -439 269 -411
rect 285 -439 286 -411
rect 296 -412 297 -390
rect 369 -439 370 -411
rect 478 -439 479 -411
rect 541 -412 542 -390
rect 569 -439 570 -411
rect 79 -414 80 -390
rect 240 -439 241 -413
rect 247 -414 248 -390
rect 296 -439 297 -413
rect 380 -414 381 -390
rect 380 -439 381 -413
rect 380 -414 381 -390
rect 380 -439 381 -413
rect 387 -414 388 -390
rect 618 -414 619 -390
rect 79 -439 80 -415
rect 215 -439 216 -415
rect 247 -439 248 -415
rect 261 -416 262 -390
rect 289 -439 290 -415
rect 331 -439 332 -415
rect 387 -439 388 -415
rect 443 -416 444 -390
rect 467 -439 468 -415
rect 590 -439 591 -415
rect 86 -418 87 -390
rect 324 -418 325 -390
rect 345 -418 346 -390
rect 443 -439 444 -417
rect 471 -418 472 -390
rect 492 -439 493 -417
rect 499 -418 500 -390
rect 541 -439 542 -417
rect 555 -418 556 -390
rect 618 -439 619 -417
rect 93 -420 94 -390
rect 93 -439 94 -419
rect 93 -420 94 -390
rect 93 -439 94 -419
rect 100 -420 101 -390
rect 159 -420 160 -390
rect 184 -439 185 -419
rect 191 -439 192 -419
rect 236 -420 237 -390
rect 345 -439 346 -419
rect 408 -420 409 -390
rect 499 -439 500 -419
rect 100 -439 101 -421
rect 145 -439 146 -421
rect 159 -439 160 -421
rect 520 -439 521 -421
rect 107 -439 108 -423
rect 198 -424 199 -390
rect 236 -439 237 -423
rect 278 -424 279 -390
rect 324 -439 325 -423
rect 506 -424 507 -390
rect 114 -426 115 -390
rect 275 -439 276 -425
rect 408 -439 409 -425
rect 457 -439 458 -425
rect 114 -439 115 -427
rect 128 -428 129 -390
rect 135 -439 136 -427
rect 166 -428 167 -390
rect 198 -439 199 -427
rect 548 -439 549 -427
rect 121 -430 122 -390
rect 310 -439 311 -429
rect 415 -439 416 -429
rect 429 -430 430 -390
rect 471 -439 472 -429
rect 86 -439 87 -431
rect 121 -439 122 -431
rect 128 -439 129 -431
rect 170 -432 171 -390
rect 261 -439 262 -431
rect 282 -432 283 -390
rect 338 -439 339 -431
rect 429 -439 430 -431
rect 142 -434 143 -390
rect 254 -439 255 -433
rect 170 -439 171 -435
rect 177 -436 178 -390
rect 205 -439 206 -435
rect 282 -439 283 -435
rect 23 -439 24 -437
rect 177 -439 178 -437
rect 9 -449 10 -447
rect 110 -496 111 -448
rect 131 -496 132 -448
rect 520 -449 521 -447
rect 541 -449 542 -447
rect 555 -496 556 -448
rect 558 -449 559 -447
rect 583 -449 584 -447
rect 611 -449 612 -447
rect 614 -496 615 -448
rect 635 -449 636 -447
rect 653 -449 654 -447
rect 660 -496 661 -448
rect 667 -449 668 -447
rect 9 -496 10 -450
rect 355 -496 356 -450
rect 369 -451 370 -447
rect 534 -451 535 -447
rect 583 -496 584 -450
rect 604 -451 605 -447
rect 646 -451 647 -447
rect 646 -496 647 -450
rect 646 -451 647 -447
rect 646 -496 647 -450
rect 653 -496 654 -450
rect 663 -451 664 -447
rect 16 -453 17 -447
rect 236 -453 237 -447
rect 247 -453 248 -447
rect 285 -453 286 -447
rect 292 -453 293 -447
rect 415 -453 416 -447
rect 418 -496 419 -452
rect 534 -496 535 -452
rect 16 -496 17 -454
rect 114 -455 115 -447
rect 142 -455 143 -447
rect 170 -455 171 -447
rect 208 -496 209 -454
rect 331 -455 332 -447
rect 373 -455 374 -447
rect 499 -455 500 -447
rect 520 -496 521 -454
rect 562 -455 563 -447
rect 23 -457 24 -447
rect 180 -457 181 -447
rect 215 -457 216 -447
rect 261 -457 262 -447
rect 275 -457 276 -447
rect 338 -496 339 -456
rect 376 -457 377 -447
rect 513 -457 514 -447
rect 23 -496 24 -458
rect 86 -459 87 -447
rect 107 -459 108 -447
rect 170 -496 171 -458
rect 177 -459 178 -447
rect 373 -496 374 -458
rect 397 -459 398 -447
rect 492 -459 493 -447
rect 499 -496 500 -458
rect 509 -459 510 -447
rect 513 -496 514 -458
rect 527 -459 528 -447
rect 30 -496 31 -460
rect 138 -461 139 -447
rect 142 -496 143 -460
rect 296 -461 297 -447
rect 317 -461 318 -447
rect 317 -496 318 -460
rect 317 -461 318 -447
rect 317 -496 318 -460
rect 324 -496 325 -460
rect 415 -496 416 -460
rect 436 -461 437 -447
rect 541 -496 542 -460
rect 33 -463 34 -447
rect 37 -463 38 -447
rect 44 -463 45 -447
rect 156 -496 157 -462
rect 159 -463 160 -447
rect 359 -463 360 -447
rect 408 -496 409 -462
rect 422 -463 423 -447
rect 436 -496 437 -462
rect 618 -463 619 -447
rect 37 -496 38 -464
rect 107 -496 108 -464
rect 121 -465 122 -447
rect 138 -496 139 -464
rect 163 -465 164 -447
rect 187 -465 188 -447
rect 226 -465 227 -447
rect 226 -496 227 -464
rect 226 -465 227 -447
rect 226 -496 227 -464
rect 233 -465 234 -447
rect 303 -496 304 -464
rect 359 -496 360 -464
rect 387 -465 388 -447
rect 457 -465 458 -447
rect 509 -496 510 -464
rect 576 -465 577 -447
rect 618 -496 619 -464
rect 44 -496 45 -466
rect 149 -467 150 -447
rect 163 -496 164 -466
rect 345 -467 346 -447
rect 387 -496 388 -466
rect 471 -467 472 -447
rect 478 -467 479 -447
rect 562 -496 563 -466
rect 576 -496 577 -466
rect 597 -467 598 -447
rect 51 -469 52 -447
rect 184 -469 185 -447
rect 219 -469 220 -447
rect 233 -496 234 -468
rect 243 -469 244 -447
rect 492 -496 493 -468
rect 597 -496 598 -468
rect 625 -469 626 -447
rect 2 -471 3 -447
rect 243 -496 244 -470
rect 247 -496 248 -470
rect 464 -471 465 -447
rect 485 -471 486 -447
rect 527 -496 528 -470
rect 51 -496 52 -472
rect 100 -473 101 -447
rect 121 -496 122 -472
rect 264 -496 265 -472
rect 275 -496 276 -472
rect 352 -473 353 -447
rect 397 -496 398 -472
rect 485 -496 486 -472
rect 58 -475 59 -447
rect 145 -475 146 -447
rect 166 -496 167 -474
rect 184 -496 185 -474
rect 205 -475 206 -447
rect 219 -496 220 -474
rect 254 -475 255 -447
rect 289 -475 290 -447
rect 296 -496 297 -474
rect 632 -475 633 -447
rect 58 -496 59 -476
rect 401 -496 402 -476
rect 429 -477 430 -447
rect 457 -496 458 -476
rect 632 -496 633 -476
rect 639 -477 640 -447
rect 65 -479 66 -447
rect 366 -479 367 -447
rect 429 -496 430 -478
rect 443 -479 444 -447
rect 450 -479 451 -447
rect 471 -496 472 -478
rect 590 -479 591 -447
rect 639 -496 640 -478
rect 65 -496 66 -480
rect 548 -481 549 -447
rect 72 -483 73 -447
rect 201 -496 202 -482
rect 212 -496 213 -482
rect 254 -496 255 -482
rect 268 -483 269 -447
rect 289 -496 290 -482
rect 345 -496 346 -482
rect 404 -483 405 -447
rect 548 -496 549 -482
rect 569 -483 570 -447
rect 72 -496 73 -484
rect 128 -485 129 -447
rect 177 -496 178 -484
rect 191 -485 192 -447
rect 215 -496 216 -484
rect 366 -496 367 -484
rect 390 -496 391 -484
rect 443 -496 444 -484
rect 79 -487 80 -447
rect 422 -496 423 -486
rect 79 -496 80 -488
rect 93 -489 94 -447
rect 100 -496 101 -488
rect 198 -489 199 -447
rect 282 -489 283 -447
rect 464 -496 465 -488
rect 86 -496 87 -490
rect 114 -496 115 -490
rect 128 -496 129 -490
rect 191 -496 192 -490
rect 282 -496 283 -490
rect 310 -491 311 -447
rect 352 -496 353 -490
rect 450 -496 451 -490
rect 310 -496 311 -492
rect 380 -493 381 -447
rect 380 -496 381 -494
rect 569 -496 570 -494
rect 5 -553 6 -505
rect 163 -506 164 -504
rect 198 -506 199 -504
rect 362 -553 363 -505
rect 366 -553 367 -505
rect 611 -506 612 -504
rect 618 -506 619 -504
rect 628 -506 629 -504
rect 632 -506 633 -504
rect 632 -553 633 -505
rect 632 -506 633 -504
rect 632 -553 633 -505
rect 653 -506 654 -504
rect 670 -506 671 -504
rect 681 -553 682 -505
rect 688 -553 689 -505
rect 9 -508 10 -504
rect 117 -553 118 -507
rect 121 -508 122 -504
rect 124 -540 125 -507
rect 152 -508 153 -504
rect 275 -508 276 -504
rect 285 -553 286 -507
rect 569 -508 570 -504
rect 583 -508 584 -504
rect 611 -553 612 -507
rect 628 -553 629 -507
rect 646 -508 647 -504
rect 660 -508 661 -504
rect 660 -553 661 -507
rect 660 -508 661 -504
rect 660 -553 661 -507
rect 667 -553 668 -507
rect 674 -553 675 -507
rect 9 -553 10 -509
rect 61 -553 62 -509
rect 65 -553 66 -509
rect 86 -510 87 -504
rect 93 -510 94 -504
rect 100 -510 101 -504
rect 121 -553 122 -509
rect 247 -510 248 -504
rect 254 -510 255 -504
rect 254 -553 255 -509
rect 254 -510 255 -504
rect 254 -553 255 -509
rect 268 -553 269 -509
rect 296 -510 297 -504
rect 310 -510 311 -504
rect 376 -553 377 -509
rect 383 -510 384 -504
rect 492 -510 493 -504
rect 499 -510 500 -504
rect 590 -510 591 -504
rect 604 -510 605 -504
rect 614 -510 615 -504
rect 618 -553 619 -509
rect 646 -553 647 -509
rect 23 -512 24 -504
rect 58 -553 59 -511
rect 68 -512 69 -504
rect 212 -512 213 -504
rect 219 -512 220 -504
rect 275 -553 276 -511
rect 289 -512 290 -504
rect 310 -553 311 -511
rect 338 -512 339 -504
rect 348 -553 349 -511
rect 369 -512 370 -504
rect 604 -553 605 -511
rect 639 -512 640 -504
rect 653 -553 654 -511
rect 23 -553 24 -513
rect 240 -514 241 -504
rect 243 -514 244 -504
rect 562 -514 563 -504
rect 576 -514 577 -504
rect 590 -553 591 -513
rect 30 -516 31 -504
rect 208 -516 209 -504
rect 212 -553 213 -515
rect 226 -516 227 -504
rect 243 -553 244 -515
rect 387 -553 388 -515
rect 390 -516 391 -504
rect 541 -516 542 -504
rect 555 -516 556 -504
rect 562 -553 563 -515
rect 30 -553 31 -517
rect 180 -553 181 -517
rect 278 -553 279 -517
rect 555 -553 556 -517
rect 37 -520 38 -504
rect 156 -520 157 -504
rect 163 -553 164 -519
rect 436 -520 437 -504
rect 450 -520 451 -504
rect 492 -553 493 -519
rect 502 -553 503 -519
rect 513 -520 514 -504
rect 37 -553 38 -521
rect 142 -522 143 -504
rect 149 -522 150 -504
rect 219 -553 220 -521
rect 292 -553 293 -521
rect 436 -553 437 -521
rect 478 -522 479 -504
rect 569 -553 570 -521
rect 16 -524 17 -504
rect 149 -553 150 -523
rect 156 -553 157 -523
rect 233 -524 234 -504
rect 296 -553 297 -523
rect 303 -524 304 -504
rect 331 -524 332 -504
rect 541 -553 542 -523
rect 16 -553 17 -525
rect 82 -553 83 -525
rect 86 -553 87 -525
rect 100 -553 101 -525
rect 114 -553 115 -525
rect 576 -553 577 -525
rect 44 -528 45 -504
rect 215 -528 216 -504
rect 303 -553 304 -527
rect 324 -528 325 -504
rect 341 -553 342 -527
rect 450 -553 451 -527
rect 457 -528 458 -504
rect 478 -553 479 -527
rect 485 -528 486 -504
rect 583 -553 584 -527
rect 44 -553 45 -529
rect 240 -553 241 -529
rect 324 -553 325 -529
rect 345 -530 346 -504
rect 373 -530 374 -504
rect 394 -530 395 -504
rect 397 -530 398 -504
rect 597 -530 598 -504
rect 72 -532 73 -504
rect 135 -532 136 -504
rect 170 -532 171 -504
rect 226 -553 227 -531
rect 345 -553 346 -531
rect 380 -553 381 -531
rect 415 -532 416 -504
rect 527 -532 528 -504
rect 548 -532 549 -504
rect 597 -553 598 -531
rect 51 -534 52 -504
rect 72 -553 73 -533
rect 93 -553 94 -533
rect 191 -534 192 -504
rect 205 -534 206 -504
rect 233 -553 234 -533
rect 359 -534 360 -504
rect 394 -553 395 -533
rect 415 -553 416 -533
rect 429 -534 430 -504
rect 471 -534 472 -504
rect 485 -553 486 -533
rect 499 -553 500 -533
rect 527 -553 528 -533
rect 534 -534 535 -504
rect 548 -553 549 -533
rect 51 -553 52 -535
rect 79 -536 80 -504
rect 107 -536 108 -504
rect 135 -553 136 -535
rect 170 -553 171 -535
rect 282 -536 283 -504
rect 401 -536 402 -504
rect 471 -553 472 -535
rect 506 -553 507 -535
rect 520 -536 521 -504
rect 107 -553 108 -537
rect 184 -538 185 -504
rect 208 -553 209 -537
rect 429 -553 430 -537
rect 464 -538 465 -504
rect 534 -553 535 -537
rect 247 -553 248 -539
rect 261 -553 262 -539
rect 401 -553 402 -539
rect 422 -540 423 -504
rect 639 -553 640 -539
rect 128 -553 129 -541
rect 331 -553 332 -541
rect 355 -542 356 -504
rect 464 -553 465 -541
rect 513 -553 514 -541
rect 625 -542 626 -504
rect 131 -553 132 -543
rect 205 -553 206 -543
rect 313 -553 314 -543
rect 520 -553 521 -543
rect 159 -546 160 -504
rect 184 -553 185 -545
rect 355 -553 356 -545
rect 408 -546 409 -504
rect 177 -548 178 -504
rect 198 -553 199 -547
rect 408 -553 409 -547
rect 443 -548 444 -504
rect 317 -550 318 -504
rect 443 -553 444 -549
rect 271 -552 272 -504
rect 317 -553 318 -551
rect 2 -610 3 -562
rect 268 -563 269 -561
rect 275 -610 276 -562
rect 320 -563 321 -561
rect 345 -563 346 -561
rect 422 -610 423 -562
rect 436 -563 437 -561
rect 618 -563 619 -561
rect 646 -563 647 -561
rect 667 -563 668 -561
rect 670 -563 671 -561
rect 684 -563 685 -561
rect 688 -563 689 -561
rect 688 -610 689 -562
rect 688 -563 689 -561
rect 688 -610 689 -562
rect 19 -610 20 -564
rect 306 -610 307 -564
rect 310 -565 311 -561
rect 394 -565 395 -561
rect 401 -565 402 -561
rect 632 -565 633 -561
rect 653 -565 654 -561
rect 656 -565 657 -561
rect 674 -565 675 -561
rect 677 -610 678 -564
rect 23 -567 24 -561
rect 96 -610 97 -566
rect 107 -567 108 -561
rect 292 -567 293 -561
rect 296 -567 297 -561
rect 369 -610 370 -566
rect 380 -567 381 -561
rect 401 -610 402 -566
rect 404 -567 405 -561
rect 597 -567 598 -561
rect 618 -610 619 -566
rect 625 -567 626 -561
rect 653 -610 654 -566
rect 660 -567 661 -561
rect 23 -610 24 -568
rect 121 -569 122 -561
rect 128 -569 129 -561
rect 219 -569 220 -561
rect 233 -569 234 -561
rect 268 -610 269 -568
rect 278 -569 279 -561
rect 541 -569 542 -561
rect 576 -569 577 -561
rect 576 -610 577 -568
rect 576 -569 577 -561
rect 576 -610 577 -568
rect 590 -569 591 -561
rect 646 -610 647 -568
rect 9 -571 10 -561
rect 128 -610 129 -570
rect 131 -571 132 -561
rect 604 -571 605 -561
rect 9 -610 10 -572
rect 177 -573 178 -561
rect 180 -573 181 -561
rect 471 -573 472 -561
rect 478 -573 479 -561
rect 590 -610 591 -572
rect 604 -610 605 -572
rect 625 -610 626 -572
rect 30 -575 31 -561
rect 100 -575 101 -561
rect 107 -610 108 -574
rect 170 -575 171 -561
rect 243 -575 244 -561
rect 639 -575 640 -561
rect 30 -610 31 -576
rect 233 -610 234 -576
rect 247 -577 248 -561
rect 380 -610 381 -576
rect 383 -610 384 -576
rect 478 -610 479 -576
rect 499 -610 500 -576
rect 513 -577 514 -561
rect 534 -577 535 -561
rect 541 -610 542 -576
rect 562 -577 563 -561
rect 639 -610 640 -576
rect 37 -579 38 -561
rect 341 -579 342 -561
rect 345 -610 346 -578
rect 352 -579 353 -561
rect 355 -579 356 -561
rect 443 -579 444 -561
rect 457 -579 458 -561
rect 492 -579 493 -561
rect 40 -610 41 -580
rect 180 -610 181 -580
rect 184 -581 185 -561
rect 247 -610 248 -580
rect 254 -581 255 -561
rect 474 -610 475 -580
rect 485 -581 486 -561
rect 513 -610 514 -580
rect 44 -583 45 -561
rect 142 -583 143 -561
rect 149 -583 150 -561
rect 149 -610 150 -582
rect 149 -583 150 -561
rect 149 -610 150 -582
rect 163 -583 164 -561
rect 219 -610 220 -582
rect 285 -583 286 -561
rect 338 -610 339 -582
rect 366 -583 367 -561
rect 376 -583 377 -561
rect 387 -583 388 -561
rect 597 -610 598 -582
rect 51 -585 52 -561
rect 54 -591 55 -584
rect 65 -585 66 -561
rect 82 -585 83 -561
rect 93 -585 94 -561
rect 296 -610 297 -584
rect 317 -585 318 -561
rect 569 -585 570 -561
rect 16 -587 17 -561
rect 93 -610 94 -586
rect 100 -610 101 -586
rect 117 -587 118 -561
rect 121 -610 122 -586
rect 177 -610 178 -586
rect 212 -587 213 -561
rect 254 -610 255 -586
rect 289 -587 290 -561
rect 534 -610 535 -586
rect 548 -587 549 -561
rect 569 -610 570 -586
rect 51 -610 52 -588
rect 114 -589 115 -561
rect 156 -589 157 -561
rect 163 -610 164 -588
rect 226 -589 227 -561
rect 236 -610 237 -588
rect 317 -610 318 -588
rect 366 -610 367 -588
rect 632 -610 633 -588
rect 58 -610 59 -590
rect 114 -610 115 -590
rect 131 -610 132 -590
rect 282 -591 283 -561
rect 289 -610 290 -590
rect 467 -610 468 -590
rect 471 -610 472 -590
rect 611 -591 612 -561
rect 656 -610 657 -590
rect 660 -610 661 -590
rect 65 -610 66 -592
rect 103 -610 104 -592
rect 135 -593 136 -561
rect 194 -593 195 -561
rect 198 -593 199 -561
rect 226 -610 227 -592
rect 282 -610 283 -592
rect 303 -593 304 -561
rect 373 -593 374 -561
rect 443 -610 444 -592
rect 485 -610 486 -592
rect 520 -593 521 -561
rect 583 -593 584 -561
rect 611 -610 612 -592
rect 75 -595 76 -561
rect 310 -610 311 -594
rect 359 -595 360 -561
rect 583 -610 584 -594
rect 79 -610 80 -596
rect 184 -610 185 -596
rect 198 -610 199 -596
rect 243 -610 244 -596
rect 303 -610 304 -596
rect 555 -597 556 -561
rect 135 -610 136 -598
rect 261 -599 262 -561
rect 359 -610 360 -598
rect 425 -599 426 -561
rect 429 -599 430 -561
rect 457 -610 458 -598
rect 460 -599 461 -561
rect 520 -610 521 -598
rect 527 -599 528 -561
rect 555 -610 556 -598
rect 142 -610 143 -600
rect 187 -610 188 -600
rect 205 -601 206 -561
rect 429 -610 430 -600
rect 450 -601 451 -561
rect 527 -610 528 -600
rect 170 -610 171 -602
rect 191 -610 192 -602
rect 205 -610 206 -602
rect 313 -603 314 -561
rect 373 -610 374 -602
rect 397 -610 398 -602
rect 408 -603 409 -561
rect 408 -610 409 -602
rect 408 -603 409 -561
rect 408 -610 409 -602
rect 415 -603 416 -561
rect 415 -610 416 -602
rect 415 -603 416 -561
rect 415 -610 416 -602
rect 450 -610 451 -602
rect 464 -603 465 -561
rect 506 -603 507 -561
rect 548 -610 549 -602
rect 212 -610 213 -604
rect 264 -610 265 -604
rect 331 -605 332 -561
rect 506 -610 507 -604
rect 324 -607 325 -561
rect 331 -610 332 -606
rect 387 -610 388 -606
rect 436 -610 437 -606
rect 464 -610 465 -606
rect 562 -610 563 -606
rect 72 -609 73 -561
rect 324 -610 325 -608
rect 2 -620 3 -618
rect 394 -620 395 -618
rect 411 -683 412 -619
rect 590 -620 591 -618
rect 632 -620 633 -618
rect 702 -683 703 -619
rect 716 -683 717 -619
rect 730 -683 731 -619
rect 2 -683 3 -621
rect 44 -622 45 -618
rect 51 -622 52 -618
rect 114 -622 115 -618
rect 159 -622 160 -618
rect 247 -622 248 -618
rect 285 -683 286 -621
rect 471 -683 472 -621
rect 492 -622 493 -618
rect 639 -622 640 -618
rect 653 -622 654 -618
rect 660 -622 661 -618
rect 681 -683 682 -621
rect 688 -683 689 -621
rect 695 -683 696 -621
rect 719 -683 720 -621
rect 9 -624 10 -618
rect 187 -624 188 -618
rect 194 -683 195 -623
rect 289 -624 290 -618
rect 296 -624 297 -618
rect 348 -683 349 -623
rect 355 -624 356 -618
rect 359 -624 360 -618
rect 376 -683 377 -623
rect 520 -624 521 -618
rect 527 -624 528 -618
rect 604 -683 605 -623
rect 618 -624 619 -618
rect 660 -683 661 -623
rect 9 -683 10 -625
rect 86 -626 87 -618
rect 93 -626 94 -618
rect 100 -626 101 -618
rect 107 -626 108 -618
rect 352 -683 353 -625
rect 380 -626 381 -618
rect 653 -683 654 -625
rect 23 -628 24 -618
rect 96 -683 97 -627
rect 107 -683 108 -627
rect 149 -628 150 -618
rect 166 -628 167 -618
rect 170 -683 171 -627
rect 177 -628 178 -618
rect 387 -628 388 -618
rect 390 -628 391 -618
rect 576 -628 577 -618
rect 583 -628 584 -618
rect 618 -683 619 -627
rect 23 -683 24 -629
rect 173 -630 174 -618
rect 177 -683 178 -629
rect 212 -630 213 -618
rect 226 -630 227 -618
rect 261 -683 262 -629
rect 289 -683 290 -629
rect 373 -630 374 -618
rect 383 -630 384 -618
rect 569 -630 570 -618
rect 30 -632 31 -618
rect 369 -632 370 -618
rect 394 -683 395 -631
rect 408 -632 409 -618
rect 425 -683 426 -631
rect 548 -632 549 -618
rect 562 -632 563 -618
rect 590 -683 591 -631
rect 30 -683 31 -633
rect 163 -634 164 -618
rect 184 -683 185 -633
rect 278 -634 279 -618
rect 317 -634 318 -618
rect 317 -683 318 -633
rect 317 -634 318 -618
rect 317 -683 318 -633
rect 331 -634 332 -618
rect 331 -683 332 -633
rect 331 -634 332 -618
rect 331 -683 332 -633
rect 345 -634 346 -618
rect 380 -683 381 -633
rect 453 -634 454 -618
rect 667 -683 668 -633
rect 16 -683 17 -635
rect 278 -683 279 -635
rect 345 -683 346 -635
rect 492 -683 493 -635
rect 495 -636 496 -618
rect 548 -683 549 -635
rect 37 -683 38 -637
rect 61 -683 62 -637
rect 65 -638 66 -618
rect 65 -683 66 -637
rect 65 -638 66 -618
rect 65 -683 66 -637
rect 72 -683 73 -637
rect 121 -638 122 -618
rect 128 -638 129 -618
rect 163 -683 164 -637
rect 212 -683 213 -637
rect 219 -638 220 -618
rect 240 -638 241 -618
rect 254 -638 255 -618
rect 366 -638 367 -618
rect 569 -683 570 -637
rect 44 -683 45 -639
rect 89 -683 90 -639
rect 93 -683 94 -639
rect 520 -683 521 -639
rect 541 -640 542 -618
rect 562 -683 563 -639
rect 54 -683 55 -641
rect 254 -683 255 -641
rect 303 -683 304 -641
rect 366 -683 367 -641
rect 369 -683 370 -641
rect 555 -642 556 -618
rect 58 -644 59 -618
rect 75 -644 76 -618
rect 114 -683 115 -643
rect 156 -644 157 -618
rect 240 -683 241 -643
rect 268 -644 269 -618
rect 324 -644 325 -618
rect 555 -683 556 -643
rect 117 -646 118 -618
rect 166 -683 167 -645
rect 229 -683 230 -645
rect 268 -683 269 -645
rect 324 -683 325 -645
rect 401 -646 402 -618
rect 453 -683 454 -645
rect 632 -683 633 -645
rect 121 -683 122 -647
rect 145 -683 146 -647
rect 149 -683 150 -647
rect 205 -648 206 -618
rect 243 -648 244 -618
rect 282 -648 283 -618
rect 310 -648 311 -618
rect 401 -683 402 -647
rect 464 -648 465 -618
rect 611 -648 612 -618
rect 79 -650 80 -618
rect 310 -683 311 -649
rect 387 -683 388 -649
rect 464 -683 465 -649
rect 474 -650 475 -618
rect 639 -683 640 -649
rect 79 -683 80 -651
rect 128 -683 129 -651
rect 135 -652 136 -618
rect 219 -683 220 -651
rect 282 -683 283 -651
rect 583 -683 584 -651
rect 142 -654 143 -618
rect 247 -683 248 -653
rect 506 -654 507 -618
rect 527 -683 528 -653
rect 534 -654 535 -618
rect 611 -683 612 -653
rect 142 -683 143 -655
rect 485 -656 486 -618
rect 499 -656 500 -618
rect 534 -683 535 -655
rect 156 -683 157 -657
rect 233 -683 234 -657
rect 243 -683 244 -657
rect 506 -683 507 -657
rect 513 -658 514 -618
rect 541 -683 542 -657
rect 198 -660 199 -618
rect 205 -683 206 -659
rect 338 -660 339 -618
rect 485 -683 486 -659
rect 135 -683 136 -661
rect 198 -683 199 -661
rect 457 -662 458 -618
rect 499 -683 500 -661
rect 191 -664 192 -618
rect 338 -683 339 -663
rect 457 -683 458 -663
rect 646 -664 647 -618
rect 191 -683 192 -665
rect 677 -683 678 -665
rect 478 -668 479 -618
rect 513 -683 514 -667
rect 625 -668 626 -618
rect 646 -683 647 -667
rect 443 -670 444 -618
rect 478 -683 479 -669
rect 597 -670 598 -618
rect 625 -683 626 -669
rect 299 -683 300 -671
rect 597 -683 598 -671
rect 429 -674 430 -618
rect 443 -683 444 -673
rect 415 -676 416 -618
rect 429 -683 430 -675
rect 415 -683 416 -677
rect 436 -678 437 -618
rect 422 -680 423 -618
rect 436 -683 437 -679
rect 422 -683 423 -681
rect 576 -683 577 -681
rect 2 -693 3 -691
rect 79 -750 80 -692
rect 82 -693 83 -691
rect 436 -693 437 -691
rect 450 -693 451 -691
rect 541 -693 542 -691
rect 632 -693 633 -691
rect 723 -750 724 -692
rect 730 -693 731 -691
rect 754 -750 755 -692
rect 800 -750 801 -692
rect 807 -750 808 -692
rect 9 -695 10 -691
rect 138 -695 139 -691
rect 215 -695 216 -691
rect 310 -695 311 -691
rect 341 -750 342 -694
rect 471 -695 472 -691
rect 478 -695 479 -691
rect 478 -750 479 -694
rect 478 -695 479 -691
rect 478 -750 479 -694
rect 534 -695 535 -691
rect 716 -750 717 -694
rect 16 -750 17 -696
rect 324 -697 325 -691
rect 345 -697 346 -691
rect 527 -697 528 -691
rect 674 -697 675 -691
rect 695 -697 696 -691
rect 702 -697 703 -691
rect 744 -750 745 -696
rect 19 -699 20 -691
rect 103 -699 104 -691
rect 121 -699 122 -691
rect 163 -750 164 -698
rect 219 -699 220 -691
rect 219 -750 220 -698
rect 219 -699 220 -691
rect 219 -750 220 -698
rect 226 -699 227 -691
rect 261 -699 262 -691
rect 278 -699 279 -691
rect 583 -699 584 -691
rect 653 -699 654 -691
rect 695 -750 696 -698
rect 9 -750 10 -700
rect 226 -750 227 -700
rect 236 -701 237 -691
rect 460 -701 461 -691
rect 464 -701 465 -691
rect 611 -701 612 -691
rect 646 -701 647 -691
rect 653 -750 654 -700
rect 23 -703 24 -691
rect 187 -703 188 -691
rect 254 -703 255 -691
rect 411 -703 412 -691
rect 422 -703 423 -691
rect 688 -703 689 -691
rect 23 -750 24 -704
rect 166 -705 167 -691
rect 201 -750 202 -704
rect 422 -750 423 -704
rect 429 -705 430 -691
rect 464 -750 465 -704
rect 499 -705 500 -691
rect 534 -750 535 -704
rect 569 -705 570 -691
rect 688 -750 689 -704
rect 30 -707 31 -691
rect 240 -707 241 -691
rect 254 -750 255 -706
rect 289 -707 290 -691
rect 296 -707 297 -691
rect 401 -707 402 -691
rect 408 -707 409 -691
rect 632 -750 633 -706
rect 30 -750 31 -708
rect 93 -709 94 -691
rect 100 -709 101 -691
rect 387 -709 388 -691
rect 401 -750 402 -708
rect 457 -709 458 -691
rect 467 -709 468 -691
rect 569 -750 570 -708
rect 576 -709 577 -691
rect 611 -750 612 -708
rect 37 -711 38 -691
rect 89 -711 90 -691
rect 93 -750 94 -710
rect 156 -711 157 -691
rect 240 -750 241 -710
rect 429 -750 430 -710
rect 432 -750 433 -710
rect 625 -711 626 -691
rect 2 -750 3 -712
rect 89 -750 90 -712
rect 100 -750 101 -712
rect 737 -750 738 -712
rect 40 -750 41 -714
rect 303 -715 304 -691
rect 310 -750 311 -714
rect 331 -715 332 -691
rect 352 -715 353 -691
rect 362 -715 363 -691
rect 366 -715 367 -691
rect 618 -715 619 -691
rect 44 -717 45 -691
rect 191 -717 192 -691
rect 233 -717 234 -691
rect 352 -750 353 -716
rect 359 -717 360 -691
rect 674 -750 675 -716
rect 44 -750 45 -718
rect 124 -750 125 -718
rect 128 -719 129 -691
rect 128 -750 129 -718
rect 128 -719 129 -691
rect 128 -750 129 -718
rect 135 -750 136 -718
rect 212 -719 213 -691
rect 247 -719 248 -691
rect 362 -750 363 -718
rect 373 -719 374 -691
rect 383 -745 384 -718
rect 408 -750 409 -718
rect 604 -719 605 -691
rect 58 -750 59 -720
rect 65 -721 66 -691
rect 72 -721 73 -691
rect 72 -750 73 -720
rect 72 -721 73 -691
rect 72 -750 73 -720
rect 142 -721 143 -691
rect 303 -750 304 -720
rect 317 -721 318 -691
rect 345 -750 346 -720
rect 373 -750 374 -720
rect 453 -721 454 -691
rect 548 -721 549 -691
rect 576 -750 577 -720
rect 583 -750 584 -720
rect 681 -750 682 -720
rect 65 -750 66 -722
rect 394 -723 395 -691
rect 415 -723 416 -691
rect 499 -750 500 -722
rect 562 -723 563 -691
rect 625 -750 626 -722
rect 142 -750 143 -724
rect 282 -750 283 -724
rect 296 -750 297 -724
rect 369 -725 370 -691
rect 436 -750 437 -724
rect 520 -725 521 -691
rect 565 -750 566 -724
rect 604 -750 605 -724
rect 149 -727 150 -691
rect 212 -750 213 -726
rect 247 -750 248 -726
rect 667 -727 668 -691
rect 114 -729 115 -691
rect 149 -750 150 -728
rect 156 -750 157 -728
rect 387 -750 388 -728
rect 443 -729 444 -691
rect 457 -750 458 -728
rect 492 -729 493 -691
rect 548 -750 549 -728
rect 590 -729 591 -691
rect 646 -750 647 -728
rect 114 -750 115 -730
rect 205 -731 206 -691
rect 261 -750 262 -730
rect 733 -750 734 -730
rect 184 -733 185 -691
rect 205 -750 206 -732
rect 278 -750 279 -732
rect 324 -750 325 -732
rect 331 -750 332 -732
rect 380 -733 381 -691
rect 450 -750 451 -732
rect 471 -750 472 -732
rect 492 -750 493 -732
rect 590 -750 591 -732
rect 597 -733 598 -691
rect 618 -750 619 -732
rect 639 -733 640 -691
rect 667 -750 668 -732
rect 170 -735 171 -691
rect 184 -750 185 -734
rect 191 -750 192 -734
rect 268 -735 269 -691
rect 299 -735 300 -691
rect 338 -735 339 -691
rect 348 -735 349 -691
rect 415 -750 416 -734
rect 453 -750 454 -734
rect 660 -735 661 -691
rect 107 -737 108 -691
rect 268 -750 269 -736
rect 317 -750 318 -736
rect 327 -750 328 -736
rect 366 -750 367 -736
rect 562 -750 563 -736
rect 107 -750 108 -738
rect 177 -739 178 -691
rect 243 -739 244 -691
rect 639 -750 640 -738
rect 170 -750 171 -740
rect 198 -741 199 -691
rect 376 -741 377 -691
rect 443 -750 444 -740
rect 506 -741 507 -691
rect 520 -750 521 -740
rect 555 -741 556 -691
rect 597 -750 598 -740
rect 51 -750 52 -742
rect 198 -750 199 -742
rect 380 -750 381 -742
rect 702 -750 703 -742
rect 177 -750 178 -744
rect 292 -750 293 -744
rect 660 -750 661 -744
rect 485 -747 486 -691
rect 506 -750 507 -746
rect 513 -747 514 -691
rect 555 -750 556 -746
rect 485 -750 486 -748
rect 513 -750 514 -748
rect 30 -760 31 -758
rect 408 -760 409 -758
rect 429 -827 430 -759
rect 751 -827 752 -759
rect 807 -760 808 -758
rect 807 -827 808 -759
rect 807 -760 808 -758
rect 807 -827 808 -759
rect 30 -827 31 -761
rect 82 -827 83 -761
rect 89 -762 90 -758
rect 149 -762 150 -758
rect 177 -762 178 -758
rect 229 -762 230 -758
rect 243 -827 244 -761
rect 275 -827 276 -761
rect 289 -827 290 -761
rect 310 -762 311 -758
rect 327 -762 328 -758
rect 639 -762 640 -758
rect 674 -762 675 -758
rect 730 -827 731 -761
rect 733 -762 734 -758
rect 744 -762 745 -758
rect 2 -764 3 -758
rect 89 -827 90 -763
rect 107 -764 108 -758
rect 201 -827 202 -763
rect 226 -764 227 -758
rect 345 -764 346 -758
rect 387 -764 388 -758
rect 716 -764 717 -758
rect 723 -764 724 -758
rect 737 -764 738 -758
rect 23 -766 24 -758
rect 387 -827 388 -765
rect 390 -766 391 -758
rect 590 -766 591 -758
rect 604 -766 605 -758
rect 765 -827 766 -765
rect 23 -827 24 -767
rect 54 -827 55 -767
rect 58 -768 59 -758
rect 86 -768 87 -758
rect 100 -768 101 -758
rect 107 -827 108 -767
rect 121 -768 122 -758
rect 138 -827 139 -767
rect 142 -768 143 -758
rect 285 -827 286 -767
rect 299 -827 300 -767
rect 408 -827 409 -767
rect 422 -768 423 -758
rect 737 -827 738 -767
rect 37 -827 38 -769
rect 93 -770 94 -758
rect 100 -827 101 -769
rect 254 -770 255 -758
rect 261 -770 262 -758
rect 324 -827 325 -769
rect 334 -827 335 -769
rect 513 -770 514 -758
rect 527 -770 528 -758
rect 625 -770 626 -758
rect 632 -770 633 -758
rect 744 -827 745 -769
rect 51 -772 52 -758
rect 674 -827 675 -771
rect 702 -772 703 -758
rect 758 -827 759 -771
rect 58 -827 59 -773
rect 191 -774 192 -758
rect 247 -774 248 -758
rect 254 -827 255 -773
rect 341 -774 342 -758
rect 443 -774 444 -758
rect 495 -774 496 -758
rect 646 -774 647 -758
rect 712 -774 713 -758
rect 786 -827 787 -773
rect 65 -776 66 -758
rect 383 -776 384 -758
rect 390 -827 391 -775
rect 422 -827 423 -775
rect 436 -776 437 -758
rect 723 -827 724 -775
rect 65 -827 66 -777
rect 86 -827 87 -777
rect 93 -827 94 -777
rect 250 -778 251 -758
rect 345 -827 346 -777
rect 352 -778 353 -758
rect 373 -778 374 -758
rect 513 -827 514 -777
rect 541 -778 542 -758
rect 653 -778 654 -758
rect 72 -780 73 -758
rect 79 -780 80 -758
rect 121 -827 122 -779
rect 716 -827 717 -779
rect 72 -827 73 -781
rect 191 -827 192 -781
rect 247 -827 248 -781
rect 317 -782 318 -758
rect 352 -827 353 -781
rect 418 -827 419 -781
rect 439 -827 440 -781
rect 639 -827 640 -781
rect 79 -827 80 -783
rect 264 -827 265 -783
rect 303 -784 304 -758
rect 653 -827 654 -783
rect 124 -786 125 -758
rect 163 -786 164 -758
rect 170 -786 171 -758
rect 310 -827 311 -785
rect 373 -827 374 -785
rect 380 -786 381 -758
rect 383 -827 384 -785
rect 772 -827 773 -785
rect 2 -827 3 -787
rect 163 -827 164 -787
rect 170 -827 171 -787
rect 292 -827 293 -787
rect 303 -827 304 -787
rect 331 -788 332 -758
rect 380 -827 381 -787
rect 604 -827 605 -787
rect 611 -788 612 -758
rect 625 -827 626 -787
rect 632 -827 633 -787
rect 667 -788 668 -758
rect 9 -790 10 -758
rect 124 -827 125 -789
rect 149 -827 150 -789
rect 240 -790 241 -758
rect 394 -827 395 -789
rect 460 -827 461 -789
rect 464 -790 465 -758
rect 541 -827 542 -789
rect 544 -790 545 -758
rect 709 -827 710 -789
rect 9 -827 10 -791
rect 128 -792 129 -758
rect 156 -792 157 -758
rect 226 -827 227 -791
rect 240 -827 241 -791
rect 793 -827 794 -791
rect 16 -794 17 -758
rect 331 -827 332 -793
rect 362 -794 363 -758
rect 464 -827 465 -793
rect 488 -827 489 -793
rect 646 -827 647 -793
rect 16 -827 17 -795
rect 135 -796 136 -758
rect 156 -827 157 -795
rect 215 -827 216 -795
rect 397 -796 398 -758
rect 450 -796 451 -758
rect 453 -796 454 -758
rect 667 -827 668 -795
rect 44 -798 45 -758
rect 135 -827 136 -797
rect 177 -827 178 -797
rect 198 -798 199 -758
rect 212 -798 213 -758
rect 317 -827 318 -797
rect 366 -798 367 -758
rect 450 -827 451 -797
rect 548 -798 549 -758
rect 583 -798 584 -758
rect 586 -798 587 -758
rect 688 -798 689 -758
rect 44 -827 45 -799
rect 338 -800 339 -758
rect 404 -827 405 -799
rect 583 -827 584 -799
rect 590 -827 591 -799
rect 597 -800 598 -758
rect 618 -800 619 -758
rect 702 -827 703 -799
rect 128 -827 129 -801
rect 219 -802 220 -758
rect 222 -827 223 -801
rect 338 -827 339 -801
rect 411 -802 412 -758
rect 443 -827 444 -801
rect 534 -802 535 -758
rect 618 -827 619 -801
rect 681 -802 682 -758
rect 688 -827 689 -801
rect 103 -804 104 -758
rect 534 -827 535 -803
rect 555 -804 556 -758
rect 681 -827 682 -803
rect 184 -806 185 -758
rect 212 -827 213 -805
rect 219 -827 220 -805
rect 268 -806 269 -758
rect 415 -806 416 -758
rect 495 -827 496 -805
rect 520 -806 521 -758
rect 555 -827 556 -805
rect 562 -806 563 -758
rect 695 -806 696 -758
rect 114 -808 115 -758
rect 184 -827 185 -807
rect 198 -827 199 -807
rect 660 -808 661 -758
rect 695 -827 696 -807
rect 754 -808 755 -758
rect 110 -827 111 -809
rect 114 -827 115 -809
rect 233 -810 234 -758
rect 366 -827 367 -809
rect 436 -827 437 -809
rect 597 -827 598 -809
rect 205 -812 206 -758
rect 233 -827 234 -811
rect 268 -827 269 -811
rect 401 -812 402 -758
rect 499 -812 500 -758
rect 562 -827 563 -811
rect 569 -812 570 -758
rect 779 -827 780 -811
rect 205 -827 206 -813
rect 236 -814 237 -758
rect 359 -814 360 -758
rect 569 -827 570 -813
rect 576 -814 577 -758
rect 611 -827 612 -813
rect 296 -816 297 -758
rect 359 -827 360 -815
rect 499 -827 500 -815
rect 506 -816 507 -758
rect 520 -827 521 -815
rect 803 -827 804 -815
rect 296 -827 297 -817
rect 548 -827 549 -817
rect 471 -820 472 -758
rect 506 -827 507 -819
rect 523 -827 524 -819
rect 576 -827 577 -819
rect 457 -822 458 -758
rect 471 -827 472 -821
rect 530 -822 531 -758
rect 660 -827 661 -821
rect 457 -827 458 -823
rect 478 -824 479 -758
rect 478 -827 479 -825
rect 492 -826 493 -758
rect 9 -837 10 -835
rect 240 -837 241 -835
rect 278 -914 279 -836
rect 793 -837 794 -835
rect 803 -837 804 -835
rect 807 -837 808 -835
rect 9 -914 10 -838
rect 149 -839 150 -835
rect 159 -914 160 -838
rect 457 -914 458 -838
rect 460 -839 461 -835
rect 765 -839 766 -835
rect 16 -841 17 -835
rect 173 -914 174 -840
rect 184 -841 185 -835
rect 296 -841 297 -835
rect 366 -841 367 -835
rect 436 -841 437 -835
rect 439 -841 440 -835
rect 779 -841 780 -835
rect 16 -914 17 -842
rect 180 -914 181 -842
rect 184 -914 185 -842
rect 352 -843 353 -835
rect 359 -843 360 -835
rect 436 -914 437 -842
rect 460 -914 461 -842
rect 737 -843 738 -835
rect 751 -843 752 -835
rect 775 -914 776 -842
rect 23 -914 24 -844
rect 145 -845 146 -835
rect 149 -914 150 -844
rect 401 -845 402 -835
rect 404 -845 405 -835
rect 562 -845 563 -835
rect 625 -845 626 -835
rect 625 -914 626 -844
rect 625 -845 626 -835
rect 625 -914 626 -844
rect 688 -845 689 -835
rect 688 -914 689 -844
rect 688 -845 689 -835
rect 688 -914 689 -844
rect 730 -845 731 -835
rect 737 -914 738 -844
rect 751 -914 752 -844
rect 782 -914 783 -844
rect 30 -914 31 -846
rect 236 -914 237 -846
rect 240 -914 241 -846
rect 247 -847 248 -835
rect 268 -847 269 -835
rect 352 -914 353 -846
rect 366 -914 367 -846
rect 387 -914 388 -846
rect 390 -847 391 -835
rect 786 -847 787 -835
rect 37 -849 38 -835
rect 86 -914 87 -848
rect 107 -914 108 -848
rect 156 -849 157 -835
rect 166 -849 167 -835
rect 212 -849 213 -835
rect 215 -849 216 -835
rect 674 -849 675 -835
rect 716 -849 717 -835
rect 730 -914 731 -848
rect 786 -914 787 -848
rect 796 -914 797 -848
rect 44 -851 45 -835
rect 138 -851 139 -835
rect 142 -851 143 -835
rect 142 -914 143 -850
rect 142 -851 143 -835
rect 142 -914 143 -850
rect 156 -914 157 -850
rect 534 -851 535 -835
rect 667 -851 668 -835
rect 674 -914 675 -850
rect 54 -853 55 -835
rect 772 -853 773 -835
rect 58 -855 59 -835
rect 299 -855 300 -835
rect 338 -855 339 -835
rect 667 -914 668 -854
rect 72 -857 73 -835
rect 247 -914 248 -856
rect 268 -914 269 -856
rect 317 -857 318 -835
rect 373 -857 374 -835
rect 534 -914 535 -856
rect 646 -857 647 -835
rect 772 -914 773 -856
rect 51 -914 52 -858
rect 72 -914 73 -858
rect 82 -859 83 -835
rect 639 -859 640 -835
rect 128 -861 129 -835
rect 212 -914 213 -860
rect 219 -861 220 -835
rect 243 -914 244 -860
rect 275 -861 276 -835
rect 338 -914 339 -860
rect 383 -914 384 -860
rect 765 -914 766 -860
rect 2 -863 3 -835
rect 275 -914 276 -862
rect 282 -863 283 -835
rect 317 -914 318 -862
rect 397 -914 398 -862
rect 604 -863 605 -835
rect 44 -914 45 -864
rect 128 -914 129 -864
rect 135 -914 136 -864
rect 429 -865 430 -835
rect 467 -914 468 -864
rect 681 -865 682 -835
rect 170 -867 171 -835
rect 187 -881 188 -866
rect 201 -867 202 -835
rect 359 -914 360 -866
rect 401 -914 402 -866
rect 415 -914 416 -866
rect 418 -867 419 -835
rect 618 -867 619 -835
rect 93 -869 94 -835
rect 201 -914 202 -868
rect 205 -869 206 -835
rect 205 -914 206 -868
rect 205 -869 206 -835
rect 205 -914 206 -868
rect 226 -869 227 -835
rect 289 -914 290 -868
rect 292 -869 293 -835
rect 716 -914 717 -868
rect 58 -914 59 -870
rect 226 -914 227 -870
rect 229 -914 230 -870
rect 660 -871 661 -835
rect 93 -914 94 -872
rect 114 -873 115 -835
rect 170 -914 171 -872
rect 254 -873 255 -835
rect 282 -914 283 -872
rect 373 -914 374 -872
rect 411 -914 412 -872
rect 660 -914 661 -872
rect 114 -914 115 -874
rect 121 -875 122 -835
rect 177 -875 178 -835
rect 219 -914 220 -874
rect 233 -875 234 -835
rect 261 -914 262 -874
rect 296 -914 297 -874
rect 310 -875 311 -835
rect 334 -875 335 -835
rect 429 -914 430 -874
rect 488 -875 489 -835
rect 709 -875 710 -835
rect 37 -914 38 -876
rect 233 -914 234 -876
rect 303 -877 304 -835
rect 310 -914 311 -876
rect 348 -914 349 -876
rect 709 -914 710 -876
rect 65 -879 66 -835
rect 121 -914 122 -878
rect 177 -914 178 -878
rect 653 -879 654 -835
rect 65 -914 66 -880
rect 163 -914 164 -880
rect 254 -914 255 -880
rect 303 -914 304 -880
rect 394 -881 395 -835
rect 422 -881 423 -835
rect 492 -914 493 -880
rect 506 -881 507 -835
rect 520 -914 521 -880
rect 523 -881 524 -835
rect 744 -881 745 -835
rect 324 -883 325 -835
rect 422 -914 423 -882
rect 488 -914 489 -882
rect 723 -883 724 -835
rect 191 -914 192 -884
rect 324 -914 325 -884
rect 394 -914 395 -884
rect 541 -885 542 -835
rect 569 -885 570 -835
rect 646 -914 647 -884
rect 653 -914 654 -884
rect 695 -885 696 -835
rect 450 -887 451 -835
rect 541 -914 542 -886
rect 576 -887 577 -835
rect 604 -914 605 -886
rect 611 -887 612 -835
rect 681 -914 682 -886
rect 695 -914 696 -886
rect 702 -887 703 -835
rect 450 -914 451 -888
rect 758 -889 759 -835
rect 464 -891 465 -835
rect 611 -914 612 -890
rect 618 -914 619 -890
rect 632 -891 633 -835
rect 152 -914 153 -892
rect 632 -914 633 -892
rect 464 -914 465 -894
rect 569 -914 570 -894
rect 583 -895 584 -835
rect 758 -914 759 -894
rect 495 -897 496 -835
rect 702 -914 703 -896
rect 499 -899 500 -835
rect 506 -914 507 -898
rect 513 -899 514 -835
rect 562 -914 563 -898
rect 583 -914 584 -898
rect 590 -899 591 -835
rect 478 -901 479 -835
rect 513 -914 514 -900
rect 527 -901 528 -835
rect 744 -914 745 -900
rect 100 -903 101 -835
rect 478 -914 479 -902
rect 499 -914 500 -902
rect 639 -914 640 -902
rect 79 -905 80 -835
rect 100 -914 101 -904
rect 443 -905 444 -835
rect 527 -914 528 -904
rect 530 -905 531 -835
rect 548 -905 549 -835
rect 590 -914 591 -904
rect 597 -905 598 -835
rect 79 -914 80 -906
rect 345 -907 346 -835
rect 485 -907 486 -835
rect 548 -914 549 -906
rect 555 -907 556 -835
rect 597 -914 598 -906
rect 331 -909 332 -835
rect 443 -914 444 -908
rect 471 -909 472 -835
rect 555 -914 556 -908
rect 331 -914 332 -910
rect 380 -911 381 -835
rect 408 -911 409 -835
rect 471 -914 472 -910
rect 408 -914 409 -912
rect 723 -914 724 -912
rect 9 -924 10 -922
rect 222 -924 223 -922
rect 229 -924 230 -922
rect 338 -924 339 -922
rect 348 -924 349 -922
rect 611 -924 612 -922
rect 688 -924 689 -922
rect 688 -991 689 -923
rect 688 -924 689 -922
rect 688 -991 689 -923
rect 723 -924 724 -922
rect 754 -991 755 -923
rect 779 -924 780 -922
rect 786 -924 787 -922
rect 9 -991 10 -925
rect 352 -926 353 -922
rect 366 -926 367 -922
rect 443 -926 444 -922
rect 446 -991 447 -925
rect 730 -926 731 -922
rect 751 -926 752 -922
rect 775 -926 776 -922
rect 16 -928 17 -922
rect 117 -991 118 -927
rect 121 -928 122 -922
rect 128 -991 129 -927
rect 142 -928 143 -922
rect 152 -928 153 -922
rect 159 -991 160 -927
rect 425 -991 426 -927
rect 432 -991 433 -927
rect 513 -928 514 -922
rect 548 -928 549 -922
rect 548 -991 549 -927
rect 548 -928 549 -922
rect 548 -991 549 -927
rect 576 -928 577 -922
rect 730 -991 731 -927
rect 16 -991 17 -929
rect 100 -930 101 -922
rect 107 -930 108 -922
rect 142 -991 143 -929
rect 149 -930 150 -922
rect 373 -930 374 -922
rect 408 -930 409 -922
rect 534 -930 535 -922
rect 576 -991 577 -929
rect 646 -930 647 -922
rect 723 -991 724 -929
rect 740 -991 741 -929
rect 23 -932 24 -922
rect 233 -932 234 -922
rect 236 -932 237 -922
rect 653 -932 654 -922
rect 23 -991 24 -933
rect 103 -991 104 -933
rect 107 -991 108 -933
rect 275 -934 276 -922
rect 285 -934 286 -922
rect 422 -934 423 -922
rect 460 -934 461 -922
rect 737 -934 738 -922
rect 30 -936 31 -922
rect 411 -936 412 -922
rect 415 -936 416 -922
rect 485 -991 486 -935
rect 499 -936 500 -922
rect 695 -936 696 -922
rect 30 -991 31 -937
rect 184 -938 185 -922
rect 191 -938 192 -922
rect 198 -938 199 -922
rect 201 -938 202 -922
rect 502 -938 503 -922
rect 513 -991 514 -937
rect 555 -938 556 -922
rect 579 -938 580 -922
rect 604 -938 605 -922
rect 681 -938 682 -922
rect 737 -991 738 -937
rect 37 -940 38 -922
rect 82 -991 83 -939
rect 86 -940 87 -922
rect 257 -991 258 -939
rect 275 -991 276 -939
rect 303 -940 304 -922
rect 310 -940 311 -922
rect 313 -991 314 -939
rect 317 -940 318 -922
rect 380 -940 381 -922
rect 418 -940 419 -922
rect 597 -940 598 -922
rect 604 -991 605 -939
rect 625 -940 626 -922
rect 674 -940 675 -922
rect 681 -991 682 -939
rect 37 -991 38 -941
rect 75 -991 76 -941
rect 86 -991 87 -941
rect 96 -991 97 -941
rect 114 -942 115 -922
rect 121 -991 122 -941
rect 135 -942 136 -922
rect 233 -991 234 -941
rect 243 -942 244 -922
rect 261 -942 262 -922
rect 296 -942 297 -922
rect 303 -991 304 -941
rect 348 -991 349 -941
rect 401 -942 402 -922
rect 418 -991 419 -941
rect 499 -991 500 -941
rect 527 -942 528 -922
rect 625 -991 626 -941
rect 44 -944 45 -922
rect 397 -944 398 -922
rect 464 -991 465 -943
rect 765 -944 766 -922
rect 51 -946 52 -922
rect 100 -991 101 -945
rect 114 -991 115 -945
rect 653 -991 654 -945
rect 51 -991 52 -947
rect 93 -948 94 -922
rect 149 -991 150 -947
rect 285 -991 286 -947
rect 359 -948 360 -922
rect 401 -991 402 -947
rect 467 -948 468 -922
rect 744 -948 745 -922
rect 65 -991 66 -949
rect 289 -950 290 -922
rect 397 -991 398 -949
rect 436 -950 437 -922
rect 471 -950 472 -922
rect 611 -991 612 -949
rect 618 -950 619 -922
rect 674 -991 675 -949
rect 79 -952 80 -922
rect 135 -991 136 -951
rect 163 -952 164 -922
rect 408 -991 409 -951
rect 488 -952 489 -922
rect 695 -991 696 -951
rect 44 -991 45 -953
rect 79 -991 80 -953
rect 89 -954 90 -922
rect 562 -954 563 -922
rect 590 -954 591 -922
rect 646 -991 647 -953
rect 163 -991 164 -955
rect 212 -956 213 -922
rect 226 -956 227 -922
rect 338 -991 339 -955
rect 429 -956 430 -922
rect 590 -991 591 -955
rect 597 -991 598 -955
rect 660 -956 661 -922
rect 58 -958 59 -922
rect 429 -991 430 -957
rect 506 -958 507 -922
rect 562 -991 563 -957
rect 618 -991 619 -957
rect 772 -958 773 -922
rect 58 -991 59 -959
rect 474 -991 475 -959
rect 478 -960 479 -922
rect 506 -991 507 -959
rect 520 -960 521 -922
rect 527 -991 528 -959
rect 534 -991 535 -959
rect 758 -960 759 -922
rect 170 -991 171 -961
rect 443 -991 444 -961
rect 457 -962 458 -922
rect 478 -991 479 -961
rect 555 -991 556 -961
rect 569 -962 570 -922
rect 632 -962 633 -922
rect 660 -991 661 -961
rect 177 -991 178 -963
rect 376 -991 377 -963
rect 390 -991 391 -963
rect 569 -991 570 -963
rect 583 -964 584 -922
rect 632 -991 633 -963
rect 180 -966 181 -922
rect 380 -991 381 -965
rect 457 -991 458 -965
rect 492 -966 493 -922
rect 583 -991 584 -965
rect 639 -966 640 -922
rect 184 -991 185 -967
rect 268 -968 269 -922
rect 278 -968 279 -922
rect 758 -991 759 -967
rect 191 -991 192 -969
rect 205 -970 206 -922
rect 212 -991 213 -969
rect 219 -970 220 -922
rect 226 -991 227 -969
rect 317 -991 318 -969
rect 471 -991 472 -969
rect 520 -991 521 -969
rect 639 -991 640 -969
rect 667 -970 668 -922
rect 205 -991 206 -971
rect 240 -991 241 -971
rect 243 -991 244 -971
rect 331 -972 332 -922
rect 492 -991 493 -971
rect 541 -972 542 -922
rect 667 -991 668 -971
rect 702 -972 703 -922
rect 198 -991 199 -973
rect 331 -991 332 -973
rect 702 -991 703 -973
rect 709 -974 710 -922
rect 219 -991 220 -975
rect 261 -991 262 -975
rect 268 -991 269 -975
rect 324 -976 325 -922
rect 709 -991 710 -975
rect 716 -976 717 -922
rect 247 -978 248 -922
rect 345 -978 346 -922
rect 394 -978 395 -922
rect 716 -991 717 -977
rect 236 -991 237 -979
rect 247 -991 248 -979
rect 254 -980 255 -922
rect 362 -991 363 -979
rect 254 -991 255 -981
rect 541 -991 542 -981
rect 289 -991 290 -983
rect 450 -984 451 -922
rect 296 -991 297 -985
rect 450 -991 451 -985
rect 310 -991 311 -987
rect 436 -991 437 -987
rect 324 -991 325 -989
rect 387 -990 388 -922
rect 9 -1001 10 -999
rect 317 -1001 318 -999
rect 334 -1066 335 -1000
rect 408 -1001 409 -999
rect 411 -1066 412 -1000
rect 513 -1001 514 -999
rect 604 -1001 605 -999
rect 604 -1066 605 -1000
rect 604 -1001 605 -999
rect 604 -1066 605 -1000
rect 688 -1001 689 -999
rect 688 -1066 689 -1000
rect 688 -1001 689 -999
rect 688 -1066 689 -1000
rect 737 -1001 738 -999
rect 744 -1001 745 -999
rect 16 -1003 17 -999
rect 194 -1066 195 -1002
rect 198 -1003 199 -999
rect 369 -1003 370 -999
rect 373 -1003 374 -999
rect 383 -1027 384 -1002
rect 394 -1066 395 -1002
rect 404 -1066 405 -1002
rect 408 -1066 409 -1002
rect 464 -1066 465 -1002
rect 471 -1003 472 -999
rect 674 -1003 675 -999
rect 740 -1003 741 -999
rect 758 -1003 759 -999
rect 23 -1005 24 -999
rect 240 -1005 241 -999
rect 243 -1005 244 -999
rect 359 -1066 360 -1004
rect 362 -1005 363 -999
rect 576 -1005 577 -999
rect 23 -1066 24 -1006
rect 149 -1007 150 -999
rect 166 -1066 167 -1006
rect 222 -1007 223 -999
rect 233 -1007 234 -999
rect 331 -1007 332 -999
rect 338 -1007 339 -999
rect 366 -1066 367 -1006
rect 373 -1066 374 -1006
rect 555 -1007 556 -999
rect 576 -1066 577 -1006
rect 691 -1066 692 -1006
rect 30 -1009 31 -999
rect 243 -1066 244 -1008
rect 250 -1066 251 -1008
rect 261 -1009 262 -999
rect 268 -1009 269 -999
rect 317 -1066 318 -1008
rect 338 -1066 339 -1008
rect 499 -1009 500 -999
rect 33 -1066 34 -1010
rect 180 -1066 181 -1010
rect 191 -1011 192 -999
rect 219 -1011 220 -999
rect 247 -1011 248 -999
rect 261 -1066 262 -1010
rect 282 -1011 283 -999
rect 639 -1011 640 -999
rect 37 -1013 38 -999
rect 79 -1013 80 -999
rect 107 -1013 108 -999
rect 310 -1013 311 -999
rect 345 -1013 346 -999
rect 730 -1013 731 -999
rect 37 -1066 38 -1014
rect 107 -1066 108 -1014
rect 114 -1015 115 -999
rect 754 -1015 755 -999
rect 44 -1017 45 -999
rect 61 -1066 62 -1016
rect 65 -1017 66 -999
rect 93 -1066 94 -1016
rect 114 -1066 115 -1016
rect 121 -1017 122 -999
rect 142 -1017 143 -999
rect 152 -1066 153 -1016
rect 170 -1017 171 -999
rect 219 -1066 220 -1016
rect 296 -1017 297 -999
rect 345 -1066 346 -1016
rect 348 -1017 349 -999
rect 439 -1066 440 -1016
rect 443 -1017 444 -999
rect 548 -1017 549 -999
rect 562 -1017 563 -999
rect 730 -1066 731 -1016
rect 51 -1019 52 -999
rect 117 -1019 118 -999
rect 121 -1066 122 -1018
rect 184 -1019 185 -999
rect 205 -1019 206 -999
rect 254 -1019 255 -999
rect 275 -1019 276 -999
rect 296 -1066 297 -1018
rect 303 -1019 304 -999
rect 303 -1066 304 -1018
rect 303 -1019 304 -999
rect 303 -1066 304 -1018
rect 352 -1019 353 -999
rect 618 -1019 619 -999
rect 51 -1066 52 -1020
rect 103 -1066 104 -1020
rect 135 -1021 136 -999
rect 142 -1066 143 -1020
rect 149 -1066 150 -1020
rect 233 -1066 234 -1020
rect 352 -1066 353 -1020
rect 355 -1021 356 -999
rect 376 -1021 377 -999
rect 506 -1021 507 -999
rect 590 -1021 591 -999
rect 618 -1066 619 -1020
rect 58 -1023 59 -999
rect 184 -1066 185 -1022
rect 191 -1066 192 -1022
rect 205 -1066 206 -1022
rect 212 -1023 213 -999
rect 282 -1066 283 -1022
rect 380 -1023 381 -999
rect 387 -1066 388 -1022
rect 415 -1023 416 -999
rect 660 -1023 661 -999
rect 65 -1066 66 -1024
rect 96 -1025 97 -999
rect 135 -1066 136 -1024
rect 159 -1025 160 -999
rect 163 -1025 164 -999
rect 254 -1066 255 -1024
rect 380 -1066 381 -1024
rect 583 -1025 584 -999
rect 590 -1066 591 -1024
rect 597 -1025 598 -999
rect 72 -1027 73 -999
rect 86 -1027 87 -999
rect 170 -1066 171 -1026
rect 226 -1027 227 -999
rect 555 -1066 556 -1026
rect 597 -1066 598 -1026
rect 653 -1027 654 -999
rect 44 -1066 45 -1028
rect 86 -1066 87 -1028
rect 156 -1029 157 -999
rect 226 -1066 227 -1028
rect 310 -1066 311 -1028
rect 653 -1066 654 -1028
rect 75 -1066 76 -1030
rect 163 -1066 164 -1030
rect 397 -1031 398 -999
rect 583 -1066 584 -1030
rect 79 -1066 80 -1032
rect 128 -1033 129 -999
rect 156 -1066 157 -1032
rect 177 -1033 178 -999
rect 418 -1066 419 -1032
rect 457 -1033 458 -999
rect 478 -1033 479 -999
rect 548 -1066 549 -1032
rect 128 -1066 129 -1034
rect 289 -1035 290 -999
rect 401 -1035 402 -999
rect 457 -1066 458 -1034
rect 478 -1066 479 -1034
rect 709 -1035 710 -999
rect 177 -1066 178 -1036
rect 268 -1066 269 -1036
rect 289 -1066 290 -1036
rect 324 -1037 325 -999
rect 401 -1066 402 -1036
rect 625 -1037 626 -999
rect 646 -1037 647 -999
rect 709 -1066 710 -1036
rect 324 -1066 325 -1038
rect 520 -1039 521 -999
rect 625 -1066 626 -1038
rect 695 -1039 696 -999
rect 313 -1041 314 -999
rect 695 -1066 696 -1040
rect 212 -1066 213 -1042
rect 313 -1066 314 -1042
rect 425 -1043 426 -999
rect 660 -1066 661 -1042
rect 432 -1045 433 -999
rect 674 -1066 675 -1044
rect 436 -1047 437 -999
rect 443 -1066 444 -1046
rect 446 -1047 447 -999
rect 492 -1047 493 -999
rect 495 -1066 496 -1046
rect 513 -1066 514 -1046
rect 520 -1066 521 -1046
rect 534 -1047 535 -999
rect 646 -1066 647 -1046
rect 702 -1047 703 -999
rect 450 -1066 451 -1048
rect 611 -1049 612 -999
rect 702 -1066 703 -1048
rect 723 -1049 724 -999
rect 453 -1051 454 -999
rect 667 -1051 668 -999
rect 467 -1053 468 -999
rect 611 -1066 612 -1052
rect 667 -1066 668 -1052
rect 716 -1053 717 -999
rect 485 -1055 486 -999
rect 639 -1066 640 -1054
rect 716 -1066 717 -1054
rect 737 -1066 738 -1054
rect 278 -1066 279 -1056
rect 485 -1066 486 -1056
rect 492 -1066 493 -1056
rect 569 -1057 570 -999
rect 499 -1066 500 -1058
rect 527 -1059 528 -999
rect 541 -1059 542 -999
rect 723 -1066 724 -1058
rect 425 -1066 426 -1060
rect 527 -1066 528 -1060
rect 569 -1066 570 -1060
rect 632 -1061 633 -999
rect 429 -1066 430 -1062
rect 541 -1066 542 -1062
rect 632 -1066 633 -1062
rect 681 -1063 682 -999
rect 681 -1066 682 -1064
rect 719 -1066 720 -1064
rect 9 -1127 10 -1075
rect 121 -1076 122 -1074
rect 128 -1076 129 -1074
rect 215 -1127 216 -1075
rect 243 -1076 244 -1074
rect 362 -1127 363 -1075
rect 387 -1076 388 -1074
rect 415 -1076 416 -1074
rect 418 -1076 419 -1074
rect 660 -1076 661 -1074
rect 677 -1127 678 -1075
rect 688 -1127 689 -1075
rect 702 -1076 703 -1074
rect 702 -1127 703 -1075
rect 702 -1076 703 -1074
rect 702 -1127 703 -1075
rect 16 -1127 17 -1077
rect 30 -1127 31 -1077
rect 37 -1078 38 -1074
rect 180 -1127 181 -1077
rect 187 -1127 188 -1077
rect 261 -1078 262 -1074
rect 278 -1078 279 -1074
rect 303 -1078 304 -1074
rect 313 -1127 314 -1077
rect 408 -1127 409 -1077
rect 415 -1127 416 -1077
rect 457 -1078 458 -1074
rect 478 -1078 479 -1074
rect 691 -1078 692 -1074
rect 44 -1080 45 -1074
rect 124 -1127 125 -1079
rect 128 -1127 129 -1079
rect 212 -1080 213 -1074
rect 254 -1080 255 -1074
rect 310 -1080 311 -1074
rect 324 -1080 325 -1074
rect 387 -1127 388 -1079
rect 394 -1080 395 -1074
rect 436 -1127 437 -1079
rect 443 -1080 444 -1074
rect 443 -1127 444 -1079
rect 443 -1080 444 -1074
rect 443 -1127 444 -1079
rect 485 -1080 486 -1074
rect 716 -1080 717 -1074
rect 51 -1082 52 -1074
rect 149 -1082 150 -1074
rect 166 -1082 167 -1074
rect 201 -1082 202 -1074
rect 282 -1082 283 -1074
rect 303 -1127 304 -1081
rect 310 -1127 311 -1081
rect 681 -1082 682 -1074
rect 51 -1127 52 -1083
rect 82 -1127 83 -1083
rect 86 -1127 87 -1083
rect 240 -1127 241 -1083
rect 282 -1127 283 -1083
rect 366 -1084 367 -1074
rect 401 -1084 402 -1074
rect 478 -1127 479 -1083
rect 495 -1084 496 -1074
rect 632 -1084 633 -1074
rect 65 -1086 66 -1074
rect 177 -1086 178 -1074
rect 194 -1086 195 -1074
rect 317 -1086 318 -1074
rect 324 -1127 325 -1085
rect 348 -1127 349 -1085
rect 352 -1086 353 -1074
rect 352 -1127 353 -1085
rect 352 -1086 353 -1074
rect 352 -1127 353 -1085
rect 359 -1086 360 -1074
rect 457 -1127 458 -1085
rect 464 -1086 465 -1074
rect 485 -1127 486 -1085
rect 499 -1086 500 -1074
rect 506 -1086 507 -1074
rect 527 -1086 528 -1074
rect 527 -1127 528 -1085
rect 527 -1086 528 -1074
rect 527 -1127 528 -1085
rect 534 -1086 535 -1074
rect 590 -1086 591 -1074
rect 611 -1086 612 -1074
rect 681 -1127 682 -1085
rect 58 -1127 59 -1087
rect 65 -1127 66 -1087
rect 72 -1127 73 -1087
rect 156 -1088 157 -1074
rect 177 -1127 178 -1087
rect 261 -1127 262 -1087
rect 289 -1088 290 -1074
rect 317 -1127 318 -1087
rect 334 -1088 335 -1074
rect 618 -1088 619 -1074
rect 632 -1127 633 -1087
rect 674 -1088 675 -1074
rect 79 -1090 80 -1074
rect 159 -1127 160 -1089
rect 198 -1090 199 -1074
rect 338 -1090 339 -1074
rect 345 -1090 346 -1074
rect 401 -1127 402 -1089
rect 422 -1090 423 -1074
rect 730 -1090 731 -1074
rect 23 -1092 24 -1074
rect 198 -1127 199 -1091
rect 289 -1127 290 -1091
rect 429 -1092 430 -1074
rect 439 -1092 440 -1074
rect 499 -1127 500 -1091
rect 506 -1127 507 -1091
rect 569 -1092 570 -1074
rect 583 -1092 584 -1074
rect 590 -1127 591 -1091
rect 611 -1127 612 -1091
rect 667 -1092 668 -1074
rect 93 -1094 94 -1074
rect 383 -1127 384 -1093
rect 422 -1127 423 -1093
rect 471 -1127 472 -1093
rect 513 -1094 514 -1074
rect 534 -1127 535 -1093
rect 537 -1094 538 -1074
rect 674 -1127 675 -1093
rect 37 -1127 38 -1095
rect 93 -1127 94 -1095
rect 100 -1127 101 -1095
rect 142 -1096 143 -1074
rect 145 -1127 146 -1095
rect 254 -1127 255 -1095
rect 268 -1096 269 -1074
rect 429 -1127 430 -1095
rect 453 -1096 454 -1074
rect 667 -1127 668 -1095
rect 107 -1127 108 -1097
rect 170 -1098 171 -1074
rect 268 -1127 269 -1097
rect 481 -1098 482 -1074
rect 513 -1127 514 -1097
rect 576 -1098 577 -1074
rect 583 -1127 584 -1097
rect 597 -1098 598 -1074
rect 618 -1127 619 -1097
rect 695 -1098 696 -1074
rect 114 -1100 115 -1074
rect 114 -1127 115 -1099
rect 114 -1100 115 -1074
rect 114 -1127 115 -1099
rect 135 -1100 136 -1074
rect 278 -1127 279 -1099
rect 296 -1100 297 -1074
rect 397 -1127 398 -1099
rect 523 -1100 524 -1074
rect 569 -1127 570 -1099
rect 576 -1127 577 -1099
rect 723 -1100 724 -1074
rect 135 -1127 136 -1101
rect 226 -1102 227 -1074
rect 296 -1127 297 -1101
rect 562 -1102 563 -1074
rect 565 -1102 566 -1074
rect 604 -1102 605 -1074
rect 684 -1127 685 -1101
rect 695 -1127 696 -1101
rect 142 -1127 143 -1103
rect 380 -1104 381 -1074
rect 523 -1127 524 -1103
rect 660 -1127 661 -1103
rect 149 -1127 150 -1105
rect 233 -1106 234 -1074
rect 275 -1127 276 -1105
rect 604 -1127 605 -1105
rect 184 -1108 185 -1074
rect 226 -1127 227 -1107
rect 338 -1127 339 -1107
rect 492 -1108 493 -1074
rect 541 -1108 542 -1074
rect 646 -1108 647 -1074
rect 23 -1127 24 -1109
rect 184 -1127 185 -1109
rect 219 -1110 220 -1074
rect 233 -1127 234 -1109
rect 247 -1127 248 -1109
rect 492 -1127 493 -1109
rect 555 -1110 556 -1074
rect 562 -1127 563 -1109
rect 597 -1127 598 -1109
rect 653 -1110 654 -1074
rect 68 -1127 69 -1111
rect 646 -1127 647 -1111
rect 205 -1114 206 -1074
rect 219 -1127 220 -1113
rect 373 -1114 374 -1074
rect 464 -1127 465 -1113
rect 548 -1114 549 -1074
rect 555 -1127 556 -1113
rect 205 -1127 206 -1115
rect 331 -1116 332 -1074
rect 380 -1127 381 -1115
rect 639 -1116 640 -1074
rect 376 -1127 377 -1117
rect 639 -1127 640 -1117
rect 425 -1120 426 -1074
rect 541 -1127 542 -1119
rect 548 -1127 549 -1119
rect 625 -1120 626 -1074
rect 425 -1127 426 -1121
rect 709 -1122 710 -1074
rect 450 -1124 451 -1074
rect 653 -1127 654 -1123
rect 709 -1127 710 -1123
rect 737 -1124 738 -1074
rect 411 -1126 412 -1074
rect 450 -1127 451 -1125
rect 474 -1126 475 -1074
rect 625 -1127 626 -1125
rect 2 -1184 3 -1136
rect 128 -1137 129 -1135
rect 145 -1137 146 -1135
rect 152 -1184 153 -1136
rect 159 -1184 160 -1136
rect 268 -1137 269 -1135
rect 275 -1137 276 -1135
rect 296 -1137 297 -1135
rect 303 -1137 304 -1135
rect 310 -1137 311 -1135
rect 317 -1137 318 -1135
rect 359 -1184 360 -1136
rect 369 -1137 370 -1135
rect 639 -1137 640 -1135
rect 646 -1137 647 -1135
rect 674 -1137 675 -1135
rect 677 -1137 678 -1135
rect 709 -1137 710 -1135
rect 9 -1139 10 -1135
rect 163 -1139 164 -1135
rect 170 -1139 171 -1135
rect 562 -1139 563 -1135
rect 646 -1184 647 -1138
rect 653 -1139 654 -1135
rect 677 -1184 678 -1138
rect 681 -1184 682 -1138
rect 688 -1139 689 -1135
rect 688 -1184 689 -1138
rect 688 -1139 689 -1135
rect 688 -1184 689 -1138
rect 695 -1139 696 -1135
rect 709 -1184 710 -1138
rect 9 -1184 10 -1140
rect 247 -1141 248 -1135
rect 250 -1141 251 -1135
rect 457 -1141 458 -1135
rect 464 -1141 465 -1135
rect 464 -1184 465 -1140
rect 464 -1141 465 -1135
rect 464 -1184 465 -1140
rect 506 -1141 507 -1135
rect 520 -1184 521 -1140
rect 523 -1141 524 -1135
rect 527 -1141 528 -1135
rect 530 -1184 531 -1140
rect 534 -1141 535 -1135
rect 544 -1184 545 -1140
rect 639 -1184 640 -1140
rect 702 -1141 703 -1135
rect 702 -1184 703 -1140
rect 702 -1141 703 -1135
rect 702 -1184 703 -1140
rect 16 -1143 17 -1135
rect 44 -1143 45 -1135
rect 47 -1143 48 -1135
rect 58 -1143 59 -1135
rect 72 -1143 73 -1135
rect 194 -1143 195 -1135
rect 219 -1143 220 -1135
rect 247 -1184 248 -1142
rect 261 -1143 262 -1135
rect 373 -1143 374 -1135
rect 380 -1184 381 -1142
rect 401 -1143 402 -1135
rect 429 -1143 430 -1135
rect 555 -1143 556 -1135
rect 562 -1184 563 -1142
rect 618 -1143 619 -1135
rect 37 -1145 38 -1135
rect 65 -1184 66 -1144
rect 79 -1184 80 -1144
rect 331 -1145 332 -1135
rect 334 -1145 335 -1135
rect 443 -1145 444 -1135
rect 478 -1145 479 -1135
rect 506 -1184 507 -1144
rect 590 -1145 591 -1135
rect 618 -1184 619 -1144
rect 37 -1184 38 -1146
rect 320 -1184 321 -1146
rect 331 -1184 332 -1146
rect 492 -1147 493 -1135
rect 583 -1147 584 -1135
rect 590 -1184 591 -1146
rect 44 -1184 45 -1148
rect 215 -1149 216 -1135
rect 226 -1149 227 -1135
rect 261 -1184 262 -1148
rect 278 -1149 279 -1135
rect 625 -1149 626 -1135
rect 51 -1151 52 -1135
rect 75 -1184 76 -1150
rect 93 -1151 94 -1135
rect 180 -1151 181 -1135
rect 184 -1151 185 -1135
rect 254 -1151 255 -1135
rect 282 -1151 283 -1135
rect 422 -1151 423 -1135
rect 429 -1184 430 -1150
rect 436 -1151 437 -1135
rect 471 -1151 472 -1135
rect 478 -1184 479 -1150
rect 492 -1184 493 -1150
rect 513 -1151 514 -1135
rect 541 -1151 542 -1135
rect 583 -1184 584 -1150
rect 604 -1151 605 -1135
rect 625 -1184 626 -1150
rect 51 -1184 52 -1152
rect 149 -1153 150 -1135
rect 156 -1153 157 -1135
rect 254 -1184 255 -1152
rect 289 -1153 290 -1135
rect 289 -1184 290 -1152
rect 289 -1153 290 -1135
rect 289 -1184 290 -1152
rect 310 -1184 311 -1152
rect 324 -1153 325 -1135
rect 345 -1153 346 -1135
rect 499 -1153 500 -1135
rect 19 -1184 20 -1154
rect 324 -1184 325 -1154
rect 348 -1155 349 -1135
rect 569 -1155 570 -1135
rect 58 -1184 59 -1156
rect 205 -1157 206 -1135
rect 226 -1184 227 -1156
rect 303 -1184 304 -1156
rect 317 -1184 318 -1156
rect 667 -1157 668 -1135
rect 82 -1159 83 -1135
rect 93 -1184 94 -1158
rect 100 -1159 101 -1135
rect 194 -1184 195 -1158
rect 205 -1184 206 -1158
rect 219 -1184 220 -1158
rect 233 -1159 234 -1135
rect 268 -1184 269 -1158
rect 348 -1184 349 -1158
rect 352 -1159 353 -1135
rect 373 -1184 374 -1158
rect 408 -1159 409 -1135
rect 415 -1159 416 -1135
rect 422 -1184 423 -1158
rect 432 -1159 433 -1135
rect 534 -1184 535 -1158
rect 569 -1184 570 -1158
rect 632 -1159 633 -1135
rect 660 -1159 661 -1135
rect 667 -1184 668 -1158
rect 86 -1161 87 -1135
rect 282 -1184 283 -1160
rect 387 -1161 388 -1135
rect 408 -1184 409 -1160
rect 443 -1184 444 -1160
rect 604 -1184 605 -1160
rect 632 -1184 633 -1160
rect 656 -1184 657 -1160
rect 30 -1184 31 -1162
rect 86 -1184 87 -1162
rect 107 -1163 108 -1135
rect 208 -1184 209 -1162
rect 236 -1184 237 -1162
rect 296 -1184 297 -1162
rect 394 -1163 395 -1135
rect 401 -1184 402 -1162
rect 450 -1163 451 -1135
rect 471 -1184 472 -1162
rect 485 -1163 486 -1135
rect 499 -1184 500 -1162
rect 107 -1184 108 -1164
rect 114 -1165 115 -1135
rect 121 -1165 122 -1135
rect 233 -1184 234 -1164
rect 362 -1165 363 -1135
rect 394 -1184 395 -1164
rect 397 -1165 398 -1135
rect 576 -1165 577 -1135
rect 23 -1167 24 -1135
rect 114 -1184 115 -1166
rect 121 -1184 122 -1166
rect 338 -1167 339 -1135
rect 387 -1184 388 -1166
rect 576 -1184 577 -1166
rect 110 -1184 111 -1168
rect 128 -1184 129 -1168
rect 135 -1169 136 -1135
rect 352 -1184 353 -1168
rect 450 -1184 451 -1168
rect 548 -1169 549 -1135
rect 135 -1184 136 -1170
rect 149 -1184 150 -1170
rect 156 -1184 157 -1170
rect 177 -1184 178 -1170
rect 184 -1184 185 -1170
rect 198 -1171 199 -1135
rect 338 -1184 339 -1170
rect 513 -1184 514 -1170
rect 548 -1184 549 -1170
rect 597 -1171 598 -1135
rect 142 -1173 143 -1135
rect 660 -1184 661 -1172
rect 142 -1184 143 -1174
rect 457 -1184 458 -1174
rect 485 -1184 486 -1174
rect 674 -1184 675 -1174
rect 145 -1184 146 -1176
rect 366 -1177 367 -1135
rect 597 -1184 598 -1176
rect 611 -1177 612 -1135
rect 163 -1184 164 -1178
rect 170 -1184 171 -1178
rect 173 -1179 174 -1135
rect 240 -1184 241 -1178
rect 366 -1184 367 -1178
rect 390 -1179 391 -1135
rect 446 -1184 447 -1178
rect 611 -1184 612 -1178
rect 166 -1181 167 -1135
rect 555 -1184 556 -1180
rect 191 -1183 192 -1135
rect 198 -1184 199 -1182
rect 390 -1184 391 -1182
rect 415 -1184 416 -1182
rect 2 -1194 3 -1192
rect 152 -1194 153 -1192
rect 156 -1255 157 -1193
rect 163 -1194 164 -1192
rect 166 -1255 167 -1193
rect 191 -1194 192 -1192
rect 201 -1255 202 -1193
rect 257 -1255 258 -1193
rect 275 -1194 276 -1192
rect 296 -1194 297 -1192
rect 303 -1194 304 -1192
rect 429 -1194 430 -1192
rect 436 -1194 437 -1192
rect 576 -1194 577 -1192
rect 667 -1255 668 -1193
rect 681 -1194 682 -1192
rect 702 -1194 703 -1192
rect 705 -1255 706 -1193
rect 709 -1194 710 -1192
rect 716 -1255 717 -1193
rect 2 -1255 3 -1195
rect 107 -1196 108 -1192
rect 110 -1255 111 -1195
rect 187 -1255 188 -1195
rect 215 -1196 216 -1192
rect 247 -1196 248 -1192
rect 296 -1255 297 -1195
rect 506 -1196 507 -1192
rect 530 -1196 531 -1192
rect 632 -1196 633 -1192
rect 674 -1196 675 -1192
rect 688 -1196 689 -1192
rect 9 -1198 10 -1192
rect 23 -1198 24 -1192
rect 30 -1198 31 -1192
rect 275 -1255 276 -1197
rect 306 -1198 307 -1192
rect 352 -1198 353 -1192
rect 359 -1198 360 -1192
rect 359 -1255 360 -1197
rect 359 -1198 360 -1192
rect 359 -1255 360 -1197
rect 383 -1255 384 -1197
rect 464 -1255 465 -1197
rect 541 -1198 542 -1192
rect 590 -1198 591 -1192
rect 597 -1198 598 -1192
rect 674 -1255 675 -1197
rect 9 -1255 10 -1199
rect 44 -1200 45 -1192
rect 54 -1255 55 -1199
rect 212 -1255 213 -1199
rect 229 -1255 230 -1199
rect 282 -1200 283 -1192
rect 289 -1200 290 -1192
rect 306 -1255 307 -1199
rect 310 -1200 311 -1192
rect 317 -1255 318 -1199
rect 320 -1200 321 -1192
rect 632 -1255 633 -1199
rect 16 -1255 17 -1201
rect 75 -1202 76 -1192
rect 89 -1202 90 -1192
rect 520 -1202 521 -1192
rect 562 -1202 563 -1192
rect 653 -1255 654 -1201
rect 23 -1255 24 -1203
rect 149 -1204 150 -1192
rect 198 -1204 199 -1192
rect 289 -1255 290 -1203
rect 310 -1255 311 -1203
rect 688 -1255 689 -1203
rect 30 -1255 31 -1205
rect 107 -1255 108 -1205
rect 117 -1206 118 -1192
rect 408 -1206 409 -1192
rect 436 -1255 437 -1205
rect 471 -1206 472 -1192
rect 478 -1206 479 -1192
rect 541 -1255 542 -1205
rect 562 -1255 563 -1205
rect 702 -1255 703 -1205
rect 37 -1208 38 -1192
rect 124 -1255 125 -1207
rect 142 -1255 143 -1207
rect 506 -1255 507 -1207
rect 569 -1208 570 -1192
rect 681 -1255 682 -1207
rect 37 -1255 38 -1209
rect 184 -1210 185 -1192
rect 219 -1210 220 -1192
rect 282 -1255 283 -1209
rect 324 -1255 325 -1209
rect 373 -1210 374 -1192
rect 387 -1210 388 -1192
rect 422 -1210 423 -1192
rect 443 -1210 444 -1192
rect 555 -1210 556 -1192
rect 597 -1255 598 -1209
rect 611 -1210 612 -1192
rect 58 -1212 59 -1192
rect 173 -1212 174 -1192
rect 233 -1255 234 -1211
rect 660 -1212 661 -1192
rect 58 -1255 59 -1213
rect 86 -1255 87 -1213
rect 93 -1214 94 -1192
rect 93 -1255 94 -1213
rect 93 -1214 94 -1192
rect 93 -1255 94 -1213
rect 100 -1214 101 -1192
rect 457 -1214 458 -1192
rect 460 -1255 461 -1213
rect 576 -1255 577 -1213
rect 65 -1255 66 -1215
rect 75 -1255 76 -1215
rect 100 -1255 101 -1215
rect 114 -1255 115 -1215
rect 121 -1216 122 -1192
rect 205 -1255 206 -1215
rect 240 -1216 241 -1192
rect 338 -1255 339 -1215
rect 341 -1216 342 -1192
rect 380 -1216 381 -1192
rect 387 -1255 388 -1215
rect 453 -1216 454 -1192
rect 499 -1216 500 -1192
rect 520 -1255 521 -1215
rect 548 -1216 549 -1192
rect 555 -1255 556 -1215
rect 72 -1218 73 -1192
rect 170 -1218 171 -1192
rect 194 -1255 195 -1217
rect 240 -1255 241 -1217
rect 247 -1255 248 -1217
rect 625 -1218 626 -1192
rect 145 -1220 146 -1192
rect 250 -1255 251 -1219
rect 327 -1220 328 -1192
rect 485 -1220 486 -1192
rect 513 -1220 514 -1192
rect 569 -1255 570 -1219
rect 149 -1255 150 -1221
rect 177 -1222 178 -1192
rect 254 -1222 255 -1192
rect 485 -1255 486 -1221
rect 513 -1255 514 -1221
rect 660 -1255 661 -1221
rect 51 -1224 52 -1192
rect 177 -1255 178 -1223
rect 327 -1255 328 -1223
rect 604 -1224 605 -1192
rect 334 -1226 335 -1192
rect 478 -1255 479 -1225
rect 604 -1255 605 -1225
rect 639 -1226 640 -1192
rect 348 -1228 349 -1192
rect 625 -1255 626 -1227
rect 352 -1255 353 -1229
rect 471 -1255 472 -1229
rect 583 -1230 584 -1192
rect 639 -1255 640 -1229
rect 366 -1232 367 -1192
rect 408 -1255 409 -1231
rect 429 -1255 430 -1231
rect 548 -1255 549 -1231
rect 135 -1234 136 -1192
rect 366 -1255 367 -1233
rect 373 -1255 374 -1233
rect 397 -1255 398 -1233
rect 401 -1234 402 -1192
rect 422 -1255 423 -1233
rect 432 -1255 433 -1233
rect 443 -1255 444 -1233
rect 446 -1234 447 -1192
rect 590 -1255 591 -1233
rect 79 -1236 80 -1192
rect 135 -1255 136 -1235
rect 380 -1255 381 -1235
rect 618 -1236 619 -1192
rect 79 -1255 80 -1237
rect 128 -1238 129 -1192
rect 331 -1255 332 -1237
rect 618 -1255 619 -1237
rect 128 -1255 129 -1239
rect 226 -1240 227 -1192
rect 394 -1240 395 -1192
rect 611 -1255 612 -1239
rect 226 -1255 227 -1241
rect 261 -1242 262 -1192
rect 401 -1255 402 -1241
rect 467 -1242 468 -1192
rect 534 -1242 535 -1192
rect 583 -1255 584 -1241
rect 254 -1255 255 -1243
rect 394 -1255 395 -1243
rect 450 -1244 451 -1192
rect 646 -1244 647 -1192
rect 261 -1255 262 -1245
rect 268 -1246 269 -1192
rect 415 -1246 416 -1192
rect 646 -1255 647 -1245
rect 170 -1255 171 -1247
rect 268 -1255 269 -1247
rect 345 -1248 346 -1192
rect 415 -1255 416 -1247
rect 450 -1255 451 -1247
rect 695 -1255 696 -1247
rect 345 -1255 346 -1249
rect 390 -1250 391 -1192
rect 453 -1255 454 -1249
rect 492 -1250 493 -1192
rect 534 -1255 535 -1249
rect 712 -1255 713 -1249
rect 457 -1255 458 -1251
rect 499 -1255 500 -1251
rect 492 -1255 493 -1253
rect 527 -1255 528 -1253
rect 16 -1265 17 -1263
rect 61 -1265 62 -1263
rect 72 -1265 73 -1263
rect 688 -1265 689 -1263
rect 712 -1265 713 -1263
rect 716 -1265 717 -1263
rect 2 -1267 3 -1263
rect 72 -1326 73 -1266
rect 93 -1267 94 -1263
rect 103 -1267 104 -1263
rect 107 -1326 108 -1266
rect 313 -1267 314 -1263
rect 317 -1267 318 -1263
rect 383 -1267 384 -1263
rect 394 -1326 395 -1266
rect 681 -1267 682 -1263
rect 2 -1326 3 -1268
rect 135 -1269 136 -1263
rect 142 -1326 143 -1268
rect 156 -1269 157 -1263
rect 177 -1269 178 -1263
rect 250 -1269 251 -1263
rect 254 -1269 255 -1263
rect 261 -1269 262 -1263
rect 271 -1269 272 -1263
rect 527 -1269 528 -1263
rect 667 -1269 668 -1263
rect 670 -1326 671 -1268
rect 9 -1271 10 -1263
rect 135 -1326 136 -1270
rect 145 -1271 146 -1263
rect 289 -1271 290 -1263
rect 303 -1271 304 -1263
rect 702 -1271 703 -1263
rect 9 -1326 10 -1272
rect 187 -1273 188 -1263
rect 194 -1273 195 -1263
rect 366 -1273 367 -1263
rect 397 -1273 398 -1263
rect 611 -1273 612 -1263
rect 667 -1326 668 -1272
rect 695 -1273 696 -1263
rect 702 -1326 703 -1272
rect 705 -1273 706 -1263
rect 23 -1275 24 -1263
rect 191 -1275 192 -1263
rect 208 -1326 209 -1274
rect 219 -1275 220 -1263
rect 222 -1275 223 -1263
rect 254 -1326 255 -1274
rect 257 -1275 258 -1263
rect 289 -1326 290 -1274
rect 303 -1326 304 -1274
rect 443 -1275 444 -1263
rect 460 -1275 461 -1263
rect 527 -1326 528 -1274
rect 23 -1326 24 -1276
rect 79 -1277 80 -1263
rect 86 -1277 87 -1263
rect 93 -1326 94 -1276
rect 100 -1326 101 -1276
rect 114 -1277 115 -1263
rect 128 -1277 129 -1263
rect 198 -1326 199 -1276
rect 212 -1277 213 -1263
rect 212 -1326 213 -1276
rect 212 -1277 213 -1263
rect 212 -1326 213 -1276
rect 215 -1277 216 -1263
rect 338 -1277 339 -1263
rect 345 -1277 346 -1263
rect 345 -1326 346 -1276
rect 345 -1277 346 -1263
rect 345 -1326 346 -1276
rect 352 -1326 353 -1276
rect 597 -1277 598 -1263
rect 30 -1279 31 -1263
rect 86 -1326 87 -1278
rect 114 -1326 115 -1278
rect 233 -1279 234 -1263
rect 236 -1279 237 -1263
rect 317 -1326 318 -1278
rect 324 -1279 325 -1263
rect 408 -1279 409 -1263
rect 429 -1326 430 -1278
rect 534 -1279 535 -1263
rect 576 -1279 577 -1263
rect 597 -1326 598 -1278
rect 37 -1281 38 -1263
rect 331 -1281 332 -1263
rect 362 -1326 363 -1280
rect 520 -1281 521 -1263
rect 534 -1326 535 -1280
rect 555 -1281 556 -1263
rect 569 -1281 570 -1263
rect 576 -1326 577 -1280
rect 40 -1326 41 -1282
rect 65 -1283 66 -1263
rect 131 -1326 132 -1282
rect 236 -1326 237 -1282
rect 240 -1283 241 -1263
rect 240 -1326 241 -1282
rect 240 -1283 241 -1263
rect 240 -1326 241 -1282
rect 285 -1326 286 -1282
rect 625 -1283 626 -1263
rect 44 -1285 45 -1263
rect 82 -1326 83 -1284
rect 149 -1285 150 -1263
rect 156 -1326 157 -1284
rect 177 -1326 178 -1284
rect 646 -1285 647 -1263
rect 44 -1326 45 -1286
rect 205 -1287 206 -1263
rect 219 -1326 220 -1286
rect 474 -1326 475 -1286
rect 495 -1287 496 -1263
rect 625 -1326 626 -1286
rect 47 -1289 48 -1263
rect 478 -1289 479 -1263
rect 506 -1289 507 -1263
rect 681 -1326 682 -1288
rect 51 -1326 52 -1290
rect 163 -1291 164 -1263
rect 180 -1291 181 -1263
rect 191 -1326 192 -1290
rect 226 -1326 227 -1290
rect 247 -1291 248 -1263
rect 310 -1326 311 -1290
rect 355 -1326 356 -1290
rect 366 -1326 367 -1290
rect 569 -1326 570 -1290
rect 58 -1326 59 -1292
rect 121 -1293 122 -1263
rect 163 -1326 164 -1292
rect 275 -1293 276 -1263
rect 327 -1293 328 -1263
rect 331 -1326 332 -1292
rect 380 -1293 381 -1263
rect 611 -1326 612 -1292
rect 65 -1326 66 -1294
rect 205 -1326 206 -1294
rect 233 -1326 234 -1294
rect 453 -1295 454 -1263
rect 478 -1326 479 -1294
rect 492 -1326 493 -1294
rect 513 -1295 514 -1263
rect 639 -1295 640 -1263
rect 121 -1326 122 -1296
rect 138 -1326 139 -1296
rect 184 -1297 185 -1263
rect 296 -1297 297 -1263
rect 380 -1326 381 -1296
rect 415 -1297 416 -1263
rect 422 -1297 423 -1263
rect 555 -1326 556 -1296
rect 639 -1326 640 -1296
rect 660 -1297 661 -1263
rect 170 -1299 171 -1263
rect 184 -1326 185 -1298
rect 247 -1326 248 -1298
rect 306 -1299 307 -1263
rect 373 -1299 374 -1263
rect 415 -1326 416 -1298
rect 432 -1299 433 -1263
rect 436 -1299 437 -1263
rect 443 -1326 444 -1298
rect 502 -1326 503 -1298
rect 520 -1326 521 -1298
rect 562 -1299 563 -1263
rect 632 -1299 633 -1263
rect 660 -1326 661 -1298
rect 268 -1301 269 -1263
rect 422 -1326 423 -1300
rect 436 -1326 437 -1300
rect 485 -1301 486 -1263
rect 562 -1326 563 -1300
rect 604 -1301 605 -1263
rect 268 -1326 269 -1302
rect 282 -1303 283 -1263
rect 296 -1326 297 -1302
rect 387 -1303 388 -1263
rect 397 -1326 398 -1302
rect 457 -1326 458 -1302
rect 464 -1303 465 -1263
rect 604 -1326 605 -1302
rect 261 -1326 262 -1304
rect 282 -1326 283 -1304
rect 306 -1326 307 -1304
rect 359 -1305 360 -1263
rect 373 -1326 374 -1304
rect 513 -1326 514 -1304
rect 590 -1305 591 -1263
rect 632 -1326 633 -1304
rect 275 -1326 276 -1306
rect 369 -1326 370 -1306
rect 401 -1307 402 -1263
rect 506 -1326 507 -1306
rect 324 -1326 325 -1308
rect 590 -1326 591 -1308
rect 390 -1326 391 -1310
rect 401 -1326 402 -1310
rect 408 -1326 409 -1310
rect 471 -1311 472 -1263
rect 485 -1326 486 -1310
rect 548 -1311 549 -1263
rect 464 -1326 465 -1312
rect 618 -1313 619 -1263
rect 548 -1326 549 -1314
rect 583 -1315 584 -1263
rect 618 -1326 619 -1314
rect 653 -1315 654 -1263
rect 180 -1326 181 -1316
rect 583 -1326 584 -1316
rect 499 -1319 500 -1263
rect 653 -1326 654 -1318
rect 499 -1326 500 -1320
rect 674 -1321 675 -1263
rect 541 -1323 542 -1263
rect 674 -1326 675 -1322
rect 450 -1326 451 -1324
rect 541 -1326 542 -1324
rect 2 -1336 3 -1334
rect 177 -1336 178 -1334
rect 208 -1385 209 -1335
rect 268 -1336 269 -1334
rect 303 -1385 304 -1335
rect 397 -1336 398 -1334
rect 404 -1385 405 -1335
rect 457 -1336 458 -1334
rect 460 -1385 461 -1335
rect 604 -1336 605 -1334
rect 653 -1336 654 -1334
rect 670 -1336 671 -1334
rect 702 -1336 703 -1334
rect 702 -1385 703 -1335
rect 702 -1336 703 -1334
rect 702 -1385 703 -1335
rect 9 -1338 10 -1334
rect 201 -1385 202 -1337
rect 212 -1338 213 -1334
rect 282 -1338 283 -1334
rect 338 -1338 339 -1334
rect 590 -1338 591 -1334
rect 646 -1338 647 -1334
rect 653 -1385 654 -1337
rect 667 -1385 668 -1337
rect 681 -1338 682 -1334
rect 19 -1340 20 -1334
rect 114 -1340 115 -1334
rect 135 -1385 136 -1339
rect 233 -1340 234 -1334
rect 254 -1340 255 -1334
rect 359 -1385 360 -1339
rect 366 -1340 367 -1334
rect 597 -1340 598 -1334
rect 646 -1385 647 -1339
rect 656 -1385 657 -1339
rect 33 -1342 34 -1334
rect 131 -1342 132 -1334
rect 138 -1342 139 -1334
rect 299 -1342 300 -1334
rect 338 -1385 339 -1341
rect 415 -1342 416 -1334
rect 422 -1342 423 -1334
rect 576 -1342 577 -1334
rect 590 -1385 591 -1341
rect 639 -1342 640 -1334
rect 44 -1344 45 -1334
rect 369 -1344 370 -1334
rect 373 -1385 374 -1343
rect 513 -1344 514 -1334
rect 576 -1385 577 -1343
rect 632 -1344 633 -1334
rect 51 -1346 52 -1334
rect 243 -1385 244 -1345
rect 261 -1346 262 -1334
rect 268 -1385 269 -1345
rect 275 -1346 276 -1334
rect 282 -1385 283 -1345
rect 352 -1346 353 -1334
rect 621 -1385 622 -1345
rect 58 -1348 59 -1334
rect 82 -1348 83 -1334
rect 86 -1348 87 -1334
rect 86 -1385 87 -1347
rect 86 -1348 87 -1334
rect 86 -1385 87 -1347
rect 100 -1348 101 -1334
rect 145 -1385 146 -1347
rect 149 -1385 150 -1347
rect 156 -1348 157 -1334
rect 159 -1385 160 -1347
rect 341 -1348 342 -1334
rect 366 -1385 367 -1347
rect 555 -1348 556 -1334
rect 58 -1385 59 -1349
rect 163 -1350 164 -1334
rect 177 -1385 178 -1349
rect 184 -1350 185 -1334
rect 219 -1350 220 -1334
rect 324 -1350 325 -1334
rect 380 -1350 381 -1334
rect 394 -1385 395 -1349
rect 408 -1350 409 -1334
rect 660 -1385 661 -1349
rect 37 -1385 38 -1351
rect 184 -1385 185 -1351
rect 222 -1385 223 -1351
rect 425 -1352 426 -1334
rect 450 -1385 451 -1351
rect 541 -1352 542 -1334
rect 51 -1385 52 -1353
rect 219 -1385 220 -1353
rect 226 -1354 227 -1334
rect 254 -1385 255 -1353
rect 261 -1385 262 -1353
rect 345 -1354 346 -1334
rect 348 -1385 349 -1353
rect 408 -1385 409 -1353
rect 425 -1385 426 -1353
rect 611 -1354 612 -1334
rect 65 -1356 66 -1334
rect 327 -1356 328 -1334
rect 383 -1356 384 -1334
rect 527 -1356 528 -1334
rect 541 -1385 542 -1355
rect 674 -1356 675 -1334
rect 65 -1385 66 -1357
rect 138 -1385 139 -1357
rect 163 -1385 164 -1357
rect 198 -1358 199 -1334
rect 226 -1385 227 -1357
rect 250 -1385 251 -1357
rect 285 -1358 286 -1334
rect 345 -1385 346 -1357
rect 383 -1385 384 -1357
rect 390 -1358 391 -1334
rect 474 -1358 475 -1334
rect 618 -1358 619 -1334
rect 72 -1385 73 -1359
rect 152 -1360 153 -1334
rect 240 -1360 241 -1334
rect 275 -1385 276 -1359
rect 289 -1360 290 -1334
rect 352 -1385 353 -1359
rect 387 -1360 388 -1334
rect 436 -1360 437 -1334
rect 478 -1385 479 -1359
rect 569 -1360 570 -1334
rect 583 -1360 584 -1334
rect 611 -1385 612 -1359
rect 44 -1385 45 -1361
rect 240 -1385 241 -1361
rect 285 -1385 286 -1361
rect 289 -1385 290 -1361
rect 436 -1385 437 -1361
rect 443 -1362 444 -1334
rect 481 -1362 482 -1334
rect 625 -1362 626 -1334
rect 75 -1364 76 -1334
rect 93 -1364 94 -1334
rect 100 -1385 101 -1363
rect 170 -1364 171 -1334
rect 401 -1364 402 -1334
rect 443 -1385 444 -1363
rect 481 -1385 482 -1363
rect 604 -1385 605 -1363
rect 79 -1385 80 -1365
rect 247 -1366 248 -1334
rect 485 -1366 486 -1334
rect 485 -1385 486 -1365
rect 485 -1366 486 -1334
rect 485 -1385 486 -1365
rect 492 -1366 493 -1334
rect 527 -1385 528 -1365
rect 548 -1366 549 -1334
rect 569 -1385 570 -1365
rect 600 -1385 601 -1365
rect 625 -1385 626 -1365
rect 93 -1385 94 -1367
rect 121 -1368 122 -1334
rect 124 -1385 125 -1367
rect 324 -1385 325 -1367
rect 429 -1368 430 -1334
rect 548 -1385 549 -1367
rect 562 -1368 563 -1334
rect 583 -1385 584 -1367
rect 107 -1370 108 -1334
rect 173 -1370 174 -1334
rect 212 -1385 213 -1369
rect 247 -1385 248 -1369
rect 310 -1370 311 -1334
rect 562 -1385 563 -1369
rect 107 -1385 108 -1371
rect 205 -1385 206 -1371
rect 310 -1385 311 -1371
rect 362 -1372 363 -1334
rect 492 -1385 493 -1371
rect 506 -1372 507 -1334
rect 513 -1385 514 -1371
rect 534 -1372 535 -1334
rect 114 -1385 115 -1373
rect 142 -1374 143 -1334
rect 170 -1385 171 -1373
rect 191 -1374 192 -1334
rect 362 -1385 363 -1373
rect 555 -1385 556 -1373
rect 23 -1376 24 -1334
rect 191 -1385 192 -1375
rect 471 -1376 472 -1334
rect 534 -1385 535 -1375
rect 121 -1385 122 -1377
rect 317 -1378 318 -1334
rect 331 -1378 332 -1334
rect 471 -1385 472 -1377
rect 499 -1378 500 -1334
rect 639 -1385 640 -1377
rect 128 -1385 129 -1379
rect 198 -1385 199 -1379
rect 296 -1380 297 -1334
rect 331 -1385 332 -1379
rect 369 -1385 370 -1379
rect 499 -1385 500 -1379
rect 506 -1385 507 -1379
rect 520 -1380 521 -1334
rect 296 -1385 297 -1381
rect 418 -1385 419 -1381
rect 464 -1385 465 -1381
rect 520 -1385 521 -1381
rect 317 -1385 318 -1383
rect 390 -1385 391 -1383
rect 33 -1395 34 -1393
rect 219 -1395 220 -1393
rect 233 -1395 234 -1393
rect 296 -1395 297 -1393
rect 317 -1395 318 -1393
rect 355 -1444 356 -1394
rect 366 -1395 367 -1393
rect 450 -1395 451 -1393
rect 453 -1444 454 -1394
rect 569 -1395 570 -1393
rect 600 -1395 601 -1393
rect 667 -1395 668 -1393
rect 705 -1395 706 -1393
rect 705 -1444 706 -1394
rect 705 -1395 706 -1393
rect 705 -1444 706 -1394
rect 37 -1397 38 -1393
rect 205 -1397 206 -1393
rect 233 -1444 234 -1396
rect 520 -1397 521 -1393
rect 551 -1444 552 -1396
rect 590 -1397 591 -1393
rect 604 -1397 605 -1393
rect 604 -1444 605 -1396
rect 604 -1397 605 -1393
rect 604 -1444 605 -1396
rect 621 -1397 622 -1393
rect 639 -1397 640 -1393
rect 646 -1397 647 -1393
rect 646 -1444 647 -1396
rect 646 -1397 647 -1393
rect 646 -1444 647 -1396
rect 37 -1444 38 -1398
rect 310 -1399 311 -1393
rect 317 -1444 318 -1398
rect 327 -1444 328 -1398
rect 373 -1399 374 -1393
rect 387 -1399 388 -1393
rect 390 -1444 391 -1398
rect 443 -1399 444 -1393
rect 460 -1399 461 -1393
rect 597 -1444 598 -1398
rect 635 -1399 636 -1393
rect 660 -1399 661 -1393
rect 44 -1401 45 -1393
rect 369 -1401 370 -1393
rect 380 -1401 381 -1393
rect 485 -1401 486 -1393
rect 499 -1401 500 -1393
rect 590 -1444 591 -1400
rect 44 -1444 45 -1402
rect 138 -1403 139 -1393
rect 184 -1403 185 -1393
rect 352 -1403 353 -1393
rect 369 -1444 370 -1402
rect 562 -1403 563 -1393
rect 51 -1405 52 -1393
rect 271 -1444 272 -1404
rect 275 -1405 276 -1393
rect 285 -1405 286 -1393
rect 296 -1444 297 -1404
rect 324 -1405 325 -1393
rect 331 -1405 332 -1393
rect 380 -1444 381 -1404
rect 387 -1444 388 -1404
rect 429 -1405 430 -1393
rect 432 -1405 433 -1393
rect 534 -1405 535 -1393
rect 51 -1444 52 -1406
rect 114 -1407 115 -1393
rect 124 -1444 125 -1406
rect 135 -1444 136 -1406
rect 201 -1407 202 -1393
rect 401 -1407 402 -1393
rect 404 -1407 405 -1393
rect 429 -1444 430 -1406
rect 436 -1407 437 -1393
rect 457 -1444 458 -1406
rect 464 -1407 465 -1393
rect 506 -1407 507 -1393
rect 513 -1407 514 -1393
rect 534 -1444 535 -1406
rect 58 -1409 59 -1393
rect 156 -1409 157 -1393
rect 247 -1409 248 -1393
rect 548 -1409 549 -1393
rect 58 -1444 59 -1410
rect 163 -1411 164 -1393
rect 247 -1444 248 -1410
rect 450 -1444 451 -1410
rect 464 -1444 465 -1410
rect 583 -1411 584 -1393
rect 72 -1413 73 -1393
rect 236 -1413 237 -1393
rect 261 -1413 262 -1393
rect 376 -1444 377 -1412
rect 394 -1413 395 -1393
rect 415 -1444 416 -1412
rect 418 -1413 419 -1393
rect 527 -1413 528 -1393
rect 583 -1444 584 -1412
rect 625 -1413 626 -1393
rect 72 -1444 73 -1414
rect 149 -1415 150 -1393
rect 163 -1444 164 -1414
rect 177 -1415 178 -1393
rect 187 -1415 188 -1393
rect 394 -1444 395 -1414
rect 401 -1444 402 -1414
rect 443 -1444 444 -1414
rect 485 -1444 486 -1414
rect 541 -1415 542 -1393
rect 86 -1417 87 -1393
rect 103 -1417 104 -1393
rect 107 -1417 108 -1393
rect 345 -1444 346 -1416
rect 397 -1444 398 -1416
rect 541 -1444 542 -1416
rect 79 -1419 80 -1393
rect 86 -1444 87 -1418
rect 93 -1419 94 -1393
rect 93 -1444 94 -1418
rect 93 -1419 94 -1393
rect 93 -1444 94 -1418
rect 103 -1444 104 -1418
rect 289 -1419 290 -1393
rect 310 -1444 311 -1418
rect 373 -1444 374 -1418
rect 422 -1444 423 -1418
rect 565 -1444 566 -1418
rect 79 -1444 80 -1420
rect 226 -1421 227 -1393
rect 243 -1421 244 -1393
rect 527 -1444 528 -1420
rect 107 -1444 108 -1422
rect 121 -1444 122 -1422
rect 138 -1444 139 -1422
rect 149 -1444 150 -1422
rect 177 -1444 178 -1422
rect 359 -1444 360 -1422
rect 425 -1423 426 -1393
rect 520 -1444 521 -1422
rect 205 -1444 206 -1424
rect 226 -1444 227 -1424
rect 254 -1425 255 -1393
rect 261 -1444 262 -1424
rect 268 -1425 269 -1393
rect 366 -1444 367 -1424
rect 436 -1444 437 -1424
rect 576 -1425 577 -1393
rect 219 -1444 220 -1426
rect 268 -1444 269 -1426
rect 275 -1444 276 -1426
rect 383 -1427 384 -1393
rect 492 -1427 493 -1393
rect 506 -1444 507 -1426
rect 513 -1444 514 -1426
rect 555 -1427 556 -1393
rect 576 -1444 577 -1426
rect 611 -1427 612 -1393
rect 191 -1429 192 -1393
rect 555 -1444 556 -1428
rect 191 -1444 192 -1430
rect 212 -1431 213 -1393
rect 240 -1444 241 -1430
rect 254 -1444 255 -1430
rect 282 -1431 283 -1393
rect 499 -1444 500 -1430
rect 65 -1433 66 -1393
rect 212 -1444 213 -1432
rect 215 -1444 216 -1432
rect 282 -1444 283 -1432
rect 289 -1444 290 -1432
rect 303 -1433 304 -1393
rect 331 -1444 332 -1432
rect 338 -1433 339 -1393
rect 471 -1433 472 -1393
rect 492 -1444 493 -1432
rect 65 -1444 66 -1434
rect 170 -1435 171 -1393
rect 338 -1444 339 -1434
rect 446 -1444 447 -1434
rect 128 -1437 129 -1393
rect 303 -1444 304 -1436
rect 439 -1444 440 -1436
rect 471 -1444 472 -1436
rect 117 -1444 118 -1438
rect 128 -1444 129 -1438
rect 145 -1439 146 -1393
rect 170 -1444 171 -1438
rect 145 -1444 146 -1440
rect 408 -1441 409 -1393
rect 408 -1444 409 -1442
rect 548 -1444 549 -1442
rect 16 -1497 17 -1453
rect 177 -1454 178 -1452
rect 215 -1454 216 -1452
rect 387 -1454 388 -1452
rect 429 -1454 430 -1452
rect 569 -1454 570 -1452
rect 702 -1454 703 -1452
rect 712 -1454 713 -1452
rect 44 -1456 45 -1452
rect 117 -1456 118 -1452
rect 163 -1456 164 -1452
rect 198 -1456 199 -1452
rect 254 -1456 255 -1452
rect 306 -1497 307 -1455
rect 310 -1456 311 -1452
rect 439 -1456 440 -1452
rect 443 -1456 444 -1452
rect 534 -1456 535 -1452
rect 548 -1497 549 -1455
rect 590 -1456 591 -1452
rect 51 -1458 52 -1452
rect 180 -1497 181 -1457
rect 254 -1497 255 -1457
rect 310 -1497 311 -1457
rect 327 -1458 328 -1452
rect 331 -1458 332 -1452
rect 359 -1458 360 -1452
rect 415 -1458 416 -1452
rect 422 -1458 423 -1452
rect 443 -1497 444 -1457
rect 450 -1497 451 -1457
rect 492 -1458 493 -1452
rect 562 -1458 563 -1452
rect 604 -1458 605 -1452
rect 65 -1460 66 -1452
rect 243 -1460 244 -1452
rect 268 -1497 269 -1459
rect 394 -1497 395 -1459
rect 432 -1497 433 -1459
rect 485 -1460 486 -1452
rect 492 -1497 493 -1459
rect 527 -1460 528 -1452
rect 565 -1460 566 -1452
rect 597 -1460 598 -1452
rect 51 -1497 52 -1461
rect 65 -1497 66 -1461
rect 72 -1462 73 -1452
rect 233 -1462 234 -1452
rect 271 -1462 272 -1452
rect 408 -1462 409 -1452
rect 436 -1497 437 -1461
rect 506 -1462 507 -1452
rect 534 -1497 535 -1461
rect 565 -1497 566 -1461
rect 569 -1497 570 -1461
rect 583 -1462 584 -1452
rect 72 -1497 73 -1463
rect 191 -1464 192 -1452
rect 212 -1497 213 -1463
rect 233 -1497 234 -1463
rect 240 -1464 241 -1452
rect 408 -1497 409 -1463
rect 478 -1464 479 -1452
rect 520 -1464 521 -1452
rect 572 -1464 573 -1452
rect 583 -1497 584 -1463
rect 58 -1466 59 -1452
rect 240 -1497 241 -1465
rect 271 -1497 272 -1465
rect 303 -1466 304 -1452
rect 331 -1497 332 -1465
rect 457 -1466 458 -1452
rect 478 -1497 479 -1465
rect 541 -1466 542 -1452
rect 58 -1497 59 -1467
rect 247 -1468 248 -1452
rect 282 -1468 283 -1452
rect 366 -1497 367 -1467
rect 401 -1468 402 -1452
rect 485 -1497 486 -1467
rect 506 -1497 507 -1467
rect 562 -1497 563 -1467
rect 79 -1470 80 -1452
rect 184 -1470 185 -1452
rect 250 -1497 251 -1469
rect 401 -1497 402 -1469
rect 457 -1497 458 -1469
rect 499 -1470 500 -1452
rect 520 -1497 521 -1469
rect 576 -1470 577 -1452
rect 79 -1497 80 -1471
rect 219 -1472 220 -1452
rect 261 -1472 262 -1452
rect 282 -1497 283 -1471
rect 289 -1472 290 -1452
rect 387 -1497 388 -1471
rect 429 -1497 430 -1471
rect 499 -1497 500 -1471
rect 541 -1497 542 -1471
rect 555 -1472 556 -1452
rect 576 -1497 577 -1471
rect 590 -1497 591 -1471
rect 37 -1474 38 -1452
rect 289 -1497 290 -1473
rect 292 -1497 293 -1473
rect 373 -1497 374 -1473
rect 37 -1497 38 -1475
rect 44 -1497 45 -1475
rect 86 -1476 87 -1452
rect 156 -1476 157 -1452
rect 163 -1497 164 -1475
rect 226 -1497 227 -1475
rect 261 -1497 262 -1475
rect 338 -1476 339 -1452
rect 345 -1476 346 -1452
rect 415 -1497 416 -1475
rect 30 -1497 31 -1477
rect 86 -1497 87 -1477
rect 93 -1478 94 -1452
rect 135 -1478 136 -1452
rect 142 -1478 143 -1452
rect 198 -1497 199 -1477
rect 205 -1478 206 -1452
rect 219 -1497 220 -1477
rect 296 -1478 297 -1452
rect 345 -1497 346 -1477
rect 359 -1497 360 -1477
rect 380 -1478 381 -1452
rect 93 -1497 94 -1479
rect 107 -1480 108 -1452
rect 110 -1497 111 -1479
rect 142 -1497 143 -1479
rect 149 -1480 150 -1452
rect 191 -1497 192 -1479
rect 296 -1497 297 -1479
rect 464 -1480 465 -1452
rect 100 -1497 101 -1481
rect 425 -1497 426 -1481
rect 107 -1497 108 -1483
rect 166 -1497 167 -1483
rect 170 -1484 171 -1452
rect 229 -1484 230 -1452
rect 338 -1497 339 -1483
rect 471 -1484 472 -1452
rect 114 -1497 115 -1485
rect 128 -1486 129 -1452
rect 135 -1497 136 -1485
rect 275 -1486 276 -1452
rect 369 -1497 370 -1485
rect 555 -1497 556 -1485
rect 128 -1497 129 -1487
rect 159 -1488 160 -1452
rect 177 -1497 178 -1487
rect 352 -1497 353 -1487
rect 380 -1497 381 -1487
rect 446 -1488 447 -1452
rect 471 -1497 472 -1487
rect 513 -1488 514 -1452
rect 124 -1497 125 -1489
rect 513 -1497 514 -1489
rect 156 -1497 157 -1491
rect 527 -1497 528 -1491
rect 275 -1497 276 -1493
rect 324 -1494 325 -1452
rect 390 -1494 391 -1452
rect 464 -1497 465 -1493
rect 317 -1496 318 -1452
rect 324 -1497 325 -1495
rect 16 -1507 17 -1505
rect 170 -1507 171 -1505
rect 173 -1507 174 -1505
rect 198 -1507 199 -1505
rect 205 -1507 206 -1505
rect 275 -1507 276 -1505
rect 292 -1507 293 -1505
rect 443 -1507 444 -1505
rect 464 -1507 465 -1505
rect 474 -1546 475 -1506
rect 478 -1546 479 -1506
rect 513 -1507 514 -1505
rect 565 -1507 566 -1505
rect 569 -1507 570 -1505
rect 579 -1507 580 -1505
rect 583 -1507 584 -1505
rect 590 -1507 591 -1505
rect 590 -1546 591 -1506
rect 590 -1507 591 -1505
rect 590 -1546 591 -1506
rect 23 -1509 24 -1505
rect 54 -1509 55 -1505
rect 58 -1509 59 -1505
rect 121 -1509 122 -1505
rect 142 -1509 143 -1505
rect 177 -1546 178 -1508
rect 184 -1509 185 -1505
rect 359 -1509 360 -1505
rect 369 -1546 370 -1508
rect 436 -1509 437 -1505
rect 443 -1546 444 -1508
rect 450 -1509 451 -1505
rect 488 -1546 489 -1508
rect 555 -1509 556 -1505
rect 30 -1511 31 -1505
rect 58 -1546 59 -1510
rect 72 -1511 73 -1505
rect 149 -1511 150 -1505
rect 152 -1511 153 -1505
rect 170 -1546 171 -1510
rect 184 -1546 185 -1510
rect 289 -1511 290 -1505
rect 313 -1511 314 -1505
rect 415 -1511 416 -1505
rect 422 -1511 423 -1505
rect 520 -1511 521 -1505
rect 37 -1513 38 -1505
rect 51 -1513 52 -1505
rect 79 -1513 80 -1505
rect 121 -1546 122 -1512
rect 152 -1546 153 -1512
rect 201 -1546 202 -1512
rect 240 -1513 241 -1505
rect 541 -1513 542 -1505
rect 51 -1546 52 -1514
rect 93 -1515 94 -1505
rect 100 -1515 101 -1505
rect 142 -1546 143 -1514
rect 163 -1546 164 -1514
rect 240 -1546 241 -1514
rect 247 -1515 248 -1505
rect 303 -1515 304 -1505
rect 320 -1515 321 -1505
rect 492 -1515 493 -1505
rect 506 -1515 507 -1505
rect 506 -1546 507 -1514
rect 506 -1515 507 -1505
rect 506 -1546 507 -1514
rect 513 -1546 514 -1514
rect 548 -1515 549 -1505
rect 65 -1517 66 -1505
rect 79 -1546 80 -1516
rect 86 -1546 87 -1516
rect 254 -1517 255 -1505
rect 268 -1546 269 -1516
rect 282 -1517 283 -1505
rect 303 -1546 304 -1516
rect 345 -1517 346 -1505
rect 401 -1517 402 -1505
rect 425 -1546 426 -1516
rect 429 -1517 430 -1505
rect 464 -1546 465 -1516
rect 492 -1546 493 -1516
rect 527 -1517 528 -1505
rect 65 -1546 66 -1518
rect 208 -1519 209 -1505
rect 275 -1546 276 -1518
rect 373 -1519 374 -1505
rect 387 -1519 388 -1505
rect 527 -1546 528 -1518
rect 89 -1521 90 -1505
rect 180 -1521 181 -1505
rect 187 -1521 188 -1505
rect 254 -1546 255 -1520
rect 282 -1546 283 -1520
rect 310 -1521 311 -1505
rect 327 -1546 328 -1520
rect 485 -1521 486 -1505
rect 520 -1546 521 -1520
rect 562 -1521 563 -1505
rect 110 -1546 111 -1522
rect 128 -1523 129 -1505
rect 135 -1523 136 -1505
rect 247 -1546 248 -1522
rect 261 -1523 262 -1505
rect 310 -1546 311 -1522
rect 331 -1523 332 -1505
rect 359 -1546 360 -1522
rect 373 -1546 374 -1522
rect 380 -1523 381 -1505
rect 383 -1546 384 -1522
rect 387 -1546 388 -1522
rect 436 -1546 437 -1522
rect 457 -1523 458 -1505
rect 114 -1525 115 -1505
rect 156 -1525 157 -1505
rect 191 -1525 192 -1505
rect 205 -1546 206 -1524
rect 229 -1525 230 -1505
rect 261 -1546 262 -1524
rect 380 -1546 381 -1524
rect 401 -1546 402 -1524
rect 450 -1546 451 -1524
rect 471 -1525 472 -1505
rect 96 -1546 97 -1526
rect 114 -1546 115 -1526
rect 128 -1546 129 -1526
rect 219 -1527 220 -1505
rect 236 -1527 237 -1505
rect 331 -1546 332 -1526
rect 457 -1546 458 -1526
rect 499 -1527 500 -1505
rect 135 -1546 136 -1528
rect 296 -1529 297 -1505
rect 499 -1546 500 -1528
rect 534 -1529 535 -1505
rect 156 -1546 157 -1530
rect 429 -1546 430 -1530
rect 198 -1546 199 -1532
rect 212 -1533 213 -1505
rect 236 -1546 237 -1532
rect 345 -1546 346 -1532
rect 212 -1546 213 -1534
rect 229 -1546 230 -1534
rect 296 -1546 297 -1534
rect 317 -1535 318 -1505
rect 317 -1546 318 -1536
rect 408 -1537 409 -1505
rect 352 -1539 353 -1505
rect 408 -1546 409 -1538
rect 352 -1546 353 -1540
rect 394 -1541 395 -1505
rect 338 -1543 339 -1505
rect 394 -1546 395 -1542
rect 338 -1546 339 -1544
rect 576 -1545 577 -1505
rect 51 -1556 52 -1554
rect 107 -1556 108 -1554
rect 121 -1556 122 -1554
rect 243 -1556 244 -1554
rect 261 -1556 262 -1554
rect 285 -1556 286 -1554
rect 289 -1583 290 -1555
rect 345 -1556 346 -1554
rect 352 -1556 353 -1554
rect 352 -1583 353 -1555
rect 352 -1556 353 -1554
rect 352 -1583 353 -1555
rect 359 -1556 360 -1554
rect 387 -1556 388 -1554
rect 401 -1556 402 -1554
rect 401 -1583 402 -1555
rect 401 -1556 402 -1554
rect 401 -1583 402 -1555
rect 415 -1556 416 -1554
rect 436 -1556 437 -1554
rect 450 -1556 451 -1554
rect 471 -1583 472 -1555
rect 485 -1583 486 -1555
rect 520 -1556 521 -1554
rect 586 -1556 587 -1554
rect 590 -1556 591 -1554
rect 72 -1558 73 -1554
rect 79 -1558 80 -1554
rect 86 -1558 87 -1554
rect 222 -1558 223 -1554
rect 226 -1583 227 -1557
rect 233 -1583 234 -1557
rect 236 -1558 237 -1554
rect 247 -1558 248 -1554
rect 261 -1583 262 -1557
rect 268 -1558 269 -1554
rect 271 -1583 272 -1557
rect 359 -1583 360 -1557
rect 380 -1558 381 -1554
rect 492 -1558 493 -1554
rect 513 -1558 514 -1554
rect 513 -1583 514 -1557
rect 513 -1558 514 -1554
rect 513 -1583 514 -1557
rect 75 -1560 76 -1554
rect 79 -1583 80 -1559
rect 96 -1560 97 -1554
rect 366 -1560 367 -1554
rect 422 -1560 423 -1554
rect 502 -1560 503 -1554
rect 103 -1562 104 -1554
rect 114 -1562 115 -1554
rect 128 -1562 129 -1554
rect 327 -1562 328 -1554
rect 331 -1562 332 -1554
rect 331 -1583 332 -1561
rect 331 -1562 332 -1554
rect 331 -1583 332 -1561
rect 429 -1562 430 -1554
rect 499 -1562 500 -1554
rect 149 -1564 150 -1554
rect 177 -1564 178 -1554
rect 194 -1564 195 -1554
rect 296 -1564 297 -1554
rect 303 -1564 304 -1554
rect 303 -1583 304 -1563
rect 303 -1564 304 -1554
rect 303 -1583 304 -1563
rect 310 -1564 311 -1554
rect 369 -1564 370 -1554
rect 429 -1583 430 -1563
rect 464 -1564 465 -1554
rect 492 -1583 493 -1563
rect 506 -1564 507 -1554
rect 142 -1566 143 -1554
rect 194 -1583 195 -1565
rect 198 -1583 199 -1565
rect 222 -1583 223 -1565
rect 240 -1566 241 -1554
rect 338 -1566 339 -1554
rect 369 -1583 370 -1565
rect 394 -1566 395 -1554
rect 436 -1583 437 -1565
rect 443 -1566 444 -1554
rect 457 -1566 458 -1554
rect 464 -1583 465 -1565
rect 142 -1583 143 -1567
rect 191 -1568 192 -1554
rect 205 -1568 206 -1554
rect 229 -1583 230 -1567
rect 247 -1583 248 -1567
rect 313 -1583 314 -1567
rect 317 -1568 318 -1554
rect 390 -1583 391 -1567
rect 128 -1583 129 -1569
rect 191 -1583 192 -1569
rect 219 -1583 220 -1569
rect 254 -1570 255 -1554
rect 275 -1570 276 -1554
rect 296 -1583 297 -1569
rect 317 -1583 318 -1569
rect 478 -1570 479 -1554
rect 159 -1572 160 -1554
rect 212 -1572 213 -1554
rect 254 -1583 255 -1571
rect 282 -1583 283 -1571
rect 292 -1572 293 -1554
rect 527 -1572 528 -1554
rect 65 -1574 66 -1554
rect 159 -1583 160 -1573
rect 163 -1574 164 -1554
rect 170 -1583 171 -1573
rect 173 -1574 174 -1554
rect 201 -1583 202 -1573
rect 275 -1583 276 -1573
rect 366 -1583 367 -1573
rect 373 -1574 374 -1554
rect 394 -1583 395 -1573
rect 135 -1576 136 -1554
rect 212 -1583 213 -1575
rect 324 -1583 325 -1575
rect 380 -1583 381 -1575
rect 135 -1583 136 -1577
rect 152 -1578 153 -1554
rect 163 -1583 164 -1577
rect 184 -1578 185 -1554
rect 373 -1583 374 -1577
rect 408 -1578 409 -1554
rect 152 -1583 153 -1579
rect 177 -1583 178 -1579
rect 156 -1582 157 -1554
rect 184 -1583 185 -1581
rect 72 -1616 73 -1592
rect 82 -1616 83 -1592
rect 89 -1616 90 -1592
rect 93 -1616 94 -1592
rect 128 -1593 129 -1591
rect 156 -1593 157 -1591
rect 163 -1593 164 -1591
rect 205 -1593 206 -1591
rect 219 -1616 220 -1592
rect 240 -1593 241 -1591
rect 243 -1593 244 -1591
rect 261 -1593 262 -1591
rect 282 -1593 283 -1591
rect 289 -1593 290 -1591
rect 296 -1593 297 -1591
rect 310 -1593 311 -1591
rect 320 -1593 321 -1591
rect 338 -1593 339 -1591
rect 345 -1593 346 -1591
rect 352 -1593 353 -1591
rect 366 -1616 367 -1592
rect 373 -1593 374 -1591
rect 383 -1616 384 -1592
rect 429 -1593 430 -1591
rect 471 -1593 472 -1591
rect 485 -1593 486 -1591
rect 492 -1593 493 -1591
rect 492 -1616 493 -1592
rect 492 -1593 493 -1591
rect 492 -1616 493 -1592
rect 506 -1593 507 -1591
rect 513 -1593 514 -1591
rect 75 -1595 76 -1591
rect 79 -1595 80 -1591
rect 135 -1595 136 -1591
rect 152 -1595 153 -1591
rect 163 -1616 164 -1594
rect 194 -1595 195 -1591
rect 205 -1616 206 -1594
rect 247 -1595 248 -1591
rect 254 -1595 255 -1591
rect 369 -1595 370 -1591
rect 387 -1595 388 -1591
rect 387 -1616 388 -1594
rect 387 -1595 388 -1591
rect 387 -1616 388 -1594
rect 394 -1595 395 -1591
rect 394 -1616 395 -1594
rect 394 -1595 395 -1591
rect 394 -1616 395 -1594
rect 422 -1595 423 -1591
rect 436 -1595 437 -1591
rect 443 -1616 444 -1594
rect 485 -1616 486 -1594
rect 114 -1616 115 -1596
rect 152 -1616 153 -1596
rect 170 -1597 171 -1591
rect 170 -1616 171 -1596
rect 170 -1597 171 -1591
rect 170 -1616 171 -1596
rect 177 -1597 178 -1591
rect 268 -1597 269 -1591
rect 275 -1597 276 -1591
rect 289 -1616 290 -1596
rect 317 -1597 318 -1591
rect 345 -1616 346 -1596
rect 352 -1616 353 -1596
rect 380 -1616 381 -1596
rect 464 -1597 465 -1591
rect 471 -1616 472 -1596
rect 131 -1616 132 -1598
rect 135 -1616 136 -1598
rect 142 -1616 143 -1598
rect 145 -1599 146 -1591
rect 156 -1616 157 -1598
rect 275 -1616 276 -1598
rect 282 -1616 283 -1598
rect 310 -1616 311 -1598
rect 317 -1616 318 -1598
rect 359 -1599 360 -1591
rect 184 -1601 185 -1591
rect 215 -1616 216 -1600
rect 226 -1601 227 -1591
rect 324 -1601 325 -1591
rect 331 -1601 332 -1591
rect 334 -1616 335 -1600
rect 338 -1616 339 -1600
rect 401 -1601 402 -1591
rect 191 -1603 192 -1591
rect 201 -1616 202 -1602
rect 212 -1603 213 -1591
rect 296 -1616 297 -1602
rect 299 -1616 300 -1602
rect 359 -1616 360 -1602
rect 191 -1616 192 -1604
rect 208 -1605 209 -1591
rect 226 -1616 227 -1604
rect 341 -1616 342 -1604
rect 233 -1607 234 -1591
rect 254 -1616 255 -1606
rect 261 -1616 262 -1606
rect 303 -1607 304 -1591
rect 236 -1616 237 -1608
rect 278 -1616 279 -1608
rect 240 -1616 241 -1610
rect 268 -1616 269 -1610
rect 243 -1616 244 -1612
rect 324 -1616 325 -1612
rect 250 -1616 251 -1614
rect 303 -1616 304 -1614
rect 30 -1645 31 -1625
rect 33 -1626 34 -1624
rect 37 -1645 38 -1625
rect 180 -1626 181 -1624
rect 198 -1626 199 -1624
rect 215 -1626 216 -1624
rect 233 -1645 234 -1625
rect 236 -1626 237 -1624
rect 240 -1626 241 -1624
rect 271 -1645 272 -1625
rect 275 -1626 276 -1624
rect 317 -1626 318 -1624
rect 334 -1626 335 -1624
rect 366 -1626 367 -1624
rect 387 -1626 388 -1624
rect 387 -1645 388 -1625
rect 387 -1626 388 -1624
rect 387 -1645 388 -1625
rect 394 -1626 395 -1624
rect 394 -1645 395 -1625
rect 394 -1626 395 -1624
rect 394 -1645 395 -1625
rect 401 -1645 402 -1625
rect 443 -1626 444 -1624
rect 467 -1626 468 -1624
rect 471 -1626 472 -1624
rect 488 -1626 489 -1624
rect 492 -1626 493 -1624
rect 44 -1645 45 -1627
rect 156 -1628 157 -1624
rect 177 -1628 178 -1624
rect 219 -1628 220 -1624
rect 254 -1628 255 -1624
rect 257 -1632 258 -1627
rect 261 -1645 262 -1627
rect 352 -1628 353 -1624
rect 359 -1628 360 -1624
rect 380 -1645 381 -1627
rect 51 -1645 52 -1629
rect 86 -1630 87 -1624
rect 93 -1630 94 -1624
rect 100 -1630 101 -1624
rect 121 -1630 122 -1624
rect 142 -1630 143 -1624
rect 149 -1630 150 -1624
rect 163 -1630 164 -1624
rect 177 -1645 178 -1629
rect 201 -1645 202 -1629
rect 205 -1630 206 -1624
rect 205 -1645 206 -1629
rect 205 -1630 206 -1624
rect 205 -1645 206 -1629
rect 212 -1630 213 -1624
rect 247 -1645 248 -1629
rect 254 -1645 255 -1629
rect 289 -1630 290 -1624
rect 296 -1630 297 -1624
rect 324 -1630 325 -1624
rect 327 -1645 328 -1629
rect 352 -1645 353 -1629
rect 65 -1645 66 -1631
rect 110 -1645 111 -1631
rect 124 -1632 125 -1624
rect 135 -1632 136 -1624
rect 138 -1645 139 -1631
rect 170 -1632 171 -1624
rect 191 -1645 192 -1631
rect 240 -1645 241 -1631
rect 289 -1645 290 -1631
rect 303 -1632 304 -1624
rect 359 -1645 360 -1631
rect 72 -1634 73 -1624
rect 89 -1634 90 -1624
rect 100 -1645 101 -1633
rect 124 -1645 125 -1633
rect 135 -1645 136 -1633
rect 156 -1645 157 -1633
rect 163 -1645 164 -1633
rect 226 -1634 227 -1624
rect 264 -1634 265 -1624
rect 317 -1645 318 -1633
rect 345 -1634 346 -1624
rect 366 -1645 367 -1633
rect 72 -1645 73 -1635
rect 131 -1645 132 -1635
rect 170 -1645 171 -1635
rect 229 -1645 230 -1635
rect 275 -1645 276 -1635
rect 338 -1645 339 -1635
rect 345 -1645 346 -1635
rect 404 -1645 405 -1635
rect 79 -1645 80 -1637
rect 114 -1638 115 -1624
rect 198 -1645 199 -1637
rect 222 -1645 223 -1637
rect 226 -1645 227 -1637
rect 296 -1645 297 -1637
rect 303 -1645 304 -1637
rect 310 -1638 311 -1624
rect 58 -1645 59 -1639
rect 114 -1645 115 -1639
rect 219 -1645 220 -1639
rect 331 -1645 332 -1639
rect 86 -1645 87 -1641
rect 145 -1645 146 -1641
rect 278 -1642 279 -1624
rect 373 -1645 374 -1641
rect 107 -1645 108 -1643
rect 149 -1645 150 -1643
rect 282 -1645 283 -1643
rect 310 -1645 311 -1643
rect 19 -1680 20 -1654
rect 23 -1680 24 -1654
rect 37 -1655 38 -1653
rect 222 -1655 223 -1653
rect 226 -1655 227 -1653
rect 366 -1655 367 -1653
rect 387 -1655 388 -1653
rect 390 -1680 391 -1654
rect 44 -1657 45 -1653
rect 128 -1657 129 -1653
rect 149 -1657 150 -1653
rect 215 -1657 216 -1653
rect 219 -1657 220 -1653
rect 240 -1657 241 -1653
rect 243 -1657 244 -1653
rect 261 -1657 262 -1653
rect 268 -1657 269 -1653
rect 310 -1657 311 -1653
rect 317 -1657 318 -1653
rect 401 -1680 402 -1656
rect 51 -1659 52 -1653
rect 138 -1659 139 -1653
rect 163 -1659 164 -1653
rect 184 -1659 185 -1653
rect 191 -1659 192 -1653
rect 198 -1680 199 -1658
rect 212 -1659 213 -1653
rect 289 -1659 290 -1653
rect 296 -1659 297 -1653
rect 310 -1680 311 -1658
rect 324 -1659 325 -1653
rect 373 -1659 374 -1653
rect 65 -1661 66 -1653
rect 93 -1661 94 -1653
rect 100 -1661 101 -1653
rect 135 -1680 136 -1660
rect 156 -1661 157 -1653
rect 163 -1680 164 -1660
rect 212 -1680 213 -1660
rect 296 -1680 297 -1660
rect 331 -1661 332 -1653
rect 373 -1680 374 -1660
rect 72 -1663 73 -1653
rect 96 -1663 97 -1653
rect 103 -1680 104 -1662
rect 107 -1680 108 -1662
rect 117 -1663 118 -1653
rect 191 -1680 192 -1662
rect 226 -1680 227 -1662
rect 324 -1680 325 -1662
rect 331 -1680 332 -1662
rect 345 -1663 346 -1653
rect 366 -1680 367 -1662
rect 380 -1663 381 -1653
rect 79 -1665 80 -1653
rect 124 -1665 125 -1653
rect 156 -1680 157 -1664
rect 170 -1665 171 -1653
rect 222 -1680 223 -1664
rect 380 -1680 381 -1664
rect 86 -1667 87 -1653
rect 114 -1667 115 -1653
rect 121 -1667 122 -1653
rect 145 -1667 146 -1653
rect 229 -1680 230 -1666
rect 320 -1680 321 -1666
rect 338 -1667 339 -1653
rect 394 -1667 395 -1653
rect 121 -1680 122 -1668
rect 177 -1669 178 -1653
rect 205 -1669 206 -1653
rect 394 -1680 395 -1668
rect 145 -1680 146 -1670
rect 149 -1680 150 -1670
rect 205 -1680 206 -1670
rect 271 -1671 272 -1653
rect 282 -1671 283 -1653
rect 352 -1671 353 -1653
rect 233 -1680 234 -1672
rect 247 -1673 248 -1653
rect 254 -1673 255 -1653
rect 268 -1680 269 -1672
rect 285 -1680 286 -1672
rect 338 -1680 339 -1672
rect 348 -1680 349 -1672
rect 352 -1680 353 -1672
rect 208 -1675 209 -1653
rect 247 -1680 248 -1674
rect 261 -1680 262 -1674
rect 303 -1680 304 -1674
rect 236 -1677 237 -1653
rect 359 -1677 360 -1653
rect 240 -1680 241 -1678
rect 275 -1679 276 -1653
rect 2 -1690 3 -1688
rect 9 -1703 10 -1689
rect 16 -1703 17 -1689
rect 23 -1690 24 -1688
rect 30 -1703 31 -1689
rect 33 -1690 34 -1688
rect 79 -1690 80 -1688
rect 79 -1703 80 -1689
rect 79 -1690 80 -1688
rect 79 -1703 80 -1689
rect 89 -1703 90 -1689
rect 96 -1703 97 -1689
rect 100 -1703 101 -1689
rect 107 -1690 108 -1688
rect 114 -1690 115 -1688
rect 205 -1690 206 -1688
rect 222 -1703 223 -1689
rect 243 -1690 244 -1688
rect 254 -1690 255 -1688
rect 401 -1690 402 -1688
rect 121 -1692 122 -1688
rect 212 -1692 213 -1688
rect 226 -1692 227 -1688
rect 233 -1692 234 -1688
rect 257 -1703 258 -1691
rect 296 -1692 297 -1688
rect 317 -1692 318 -1688
rect 331 -1692 332 -1688
rect 352 -1692 353 -1688
rect 352 -1703 353 -1691
rect 352 -1692 353 -1688
rect 352 -1703 353 -1691
rect 359 -1692 360 -1688
rect 373 -1692 374 -1688
rect 121 -1703 122 -1693
rect 128 -1703 129 -1693
rect 156 -1694 157 -1688
rect 184 -1694 185 -1688
rect 191 -1694 192 -1688
rect 247 -1694 248 -1688
rect 264 -1694 265 -1688
rect 310 -1694 311 -1688
rect 135 -1696 136 -1688
rect 156 -1703 157 -1695
rect 163 -1696 164 -1688
rect 170 -1696 171 -1688
rect 194 -1703 195 -1695
rect 205 -1703 206 -1695
rect 226 -1703 227 -1695
rect 324 -1696 325 -1688
rect 131 -1698 132 -1688
rect 135 -1703 136 -1697
rect 149 -1698 150 -1688
rect 163 -1703 164 -1697
rect 170 -1703 171 -1697
rect 177 -1698 178 -1688
rect 198 -1698 199 -1688
rect 219 -1698 220 -1688
rect 229 -1698 230 -1688
rect 233 -1703 234 -1697
rect 268 -1698 269 -1688
rect 285 -1698 286 -1688
rect 292 -1703 293 -1697
rect 380 -1698 381 -1688
rect 117 -1703 118 -1699
rect 131 -1703 132 -1699
rect 173 -1700 174 -1688
rect 177 -1703 178 -1699
rect 201 -1703 202 -1699
rect 212 -1703 213 -1699
rect 275 -1700 276 -1688
rect 278 -1703 279 -1699
rect 285 -1703 286 -1699
rect 289 -1700 290 -1688
rect 296 -1703 297 -1699
rect 394 -1700 395 -1688
rect 303 -1702 304 -1688
rect 310 -1703 311 -1701
rect 324 -1703 325 -1701
rect 338 -1702 339 -1688
rect 5 -1713 6 -1711
rect 9 -1713 10 -1711
rect 128 -1713 129 -1711
rect 135 -1713 136 -1711
rect 142 -1713 143 -1711
rect 163 -1713 164 -1711
rect 170 -1713 171 -1711
rect 201 -1713 202 -1711
rect 212 -1713 213 -1711
rect 219 -1713 220 -1711
rect 233 -1713 234 -1711
rect 243 -1713 244 -1711
rect 303 -1713 304 -1711
rect 310 -1713 311 -1711
rect 317 -1713 318 -1711
rect 324 -1713 325 -1711
rect 152 -1715 153 -1711
rect 156 -1715 157 -1711
rect 177 -1715 178 -1711
rect 226 -1715 227 -1711
rect 187 -1717 188 -1711
rect 205 -1717 206 -1711
<< labels >>
rlabel pdiffusion 3 -8 3 -8 0 cellNo=8
rlabel pdiffusion 10 -8 10 -8 0 cellNo=988
rlabel pdiffusion 17 -8 17 -8 0 cellNo=55
rlabel pdiffusion 24 -8 24 -8 0 cellNo=725
rlabel pdiffusion 31 -8 31 -8 0 cellNo=438
rlabel pdiffusion 38 -8 38 -8 0 cellNo=245
rlabel pdiffusion 45 -8 45 -8 0 cellNo=394
rlabel pdiffusion 52 -8 52 -8 0 cellNo=464
rlabel pdiffusion 59 -8 59 -8 0 cellNo=603
rlabel pdiffusion 66 -8 66 -8 0 cellNo=807
rlabel pdiffusion 108 -8 108 -8 0 cellNo=16
rlabel pdiffusion 178 -8 178 -8 0 feedthrough
rlabel pdiffusion 185 -8 185 -8 0 cellNo=965
rlabel pdiffusion 192 -8 192 -8 0 cellNo=393
rlabel pdiffusion 199 -8 199 -8 0 feedthrough
rlabel pdiffusion 206 -8 206 -8 0 cellNo=382
rlabel pdiffusion 213 -8 213 -8 0 cellNo=252
rlabel pdiffusion 220 -8 220 -8 0 cellNo=545
rlabel pdiffusion 227 -8 227 -8 0 cellNo=682
rlabel pdiffusion 234 -8 234 -8 0 feedthrough
rlabel pdiffusion 241 -8 241 -8 0 cellNo=125
rlabel pdiffusion 248 -8 248 -8 0 feedthrough
rlabel pdiffusion 255 -8 255 -8 0 feedthrough
rlabel pdiffusion 276 -8 276 -8 0 cellNo=449
rlabel pdiffusion 283 -8 283 -8 0 feedthrough
rlabel pdiffusion 290 -8 290 -8 0 feedthrough
rlabel pdiffusion 297 -8 297 -8 0 cellNo=343
rlabel pdiffusion 304 -8 304 -8 0 cellNo=466
rlabel pdiffusion 3 -27 3 -27 0 cellNo=68
rlabel pdiffusion 10 -27 10 -27 0 cellNo=467
rlabel pdiffusion 17 -27 17 -27 0 cellNo=539
rlabel pdiffusion 24 -27 24 -27 0 cellNo=101
rlabel pdiffusion 31 -27 31 -27 0 cellNo=180
rlabel pdiffusion 38 -27 38 -27 0 cellNo=351
rlabel pdiffusion 45 -27 45 -27 0 cellNo=531
rlabel pdiffusion 52 -27 52 -27 0 cellNo=951
rlabel pdiffusion 143 -27 143 -27 0 feedthrough
rlabel pdiffusion 150 -27 150 -27 0 feedthrough
rlabel pdiffusion 157 -27 157 -27 0 cellNo=229
rlabel pdiffusion 164 -27 164 -27 0 cellNo=379
rlabel pdiffusion 171 -27 171 -27 0 cellNo=703
rlabel pdiffusion 178 -27 178 -27 0 cellNo=513
rlabel pdiffusion 185 -27 185 -27 0 feedthrough
rlabel pdiffusion 192 -27 192 -27 0 cellNo=317
rlabel pdiffusion 199 -27 199 -27 0 feedthrough
rlabel pdiffusion 206 -27 206 -27 0 cellNo=399
rlabel pdiffusion 213 -27 213 -27 0 cellNo=310
rlabel pdiffusion 220 -27 220 -27 0 feedthrough
rlabel pdiffusion 241 -27 241 -27 0 feedthrough
rlabel pdiffusion 248 -27 248 -27 0 cellNo=200
rlabel pdiffusion 255 -27 255 -27 0 cellNo=573
rlabel pdiffusion 262 -27 262 -27 0 cellNo=171
rlabel pdiffusion 269 -27 269 -27 0 feedthrough
rlabel pdiffusion 276 -27 276 -27 0 feedthrough
rlabel pdiffusion 283 -27 283 -27 0 cellNo=177
rlabel pdiffusion 290 -27 290 -27 0 cellNo=836
rlabel pdiffusion 297 -27 297 -27 0 feedthrough
rlabel pdiffusion 304 -27 304 -27 0 cellNo=790
rlabel pdiffusion 311 -27 311 -27 0 feedthrough
rlabel pdiffusion 318 -27 318 -27 0 cellNo=287
rlabel pdiffusion 3 -40 3 -40 0 cellNo=100
rlabel pdiffusion 10 -40 10 -40 0 cellNo=582
rlabel pdiffusion 17 -40 17 -40 0 cellNo=761
rlabel pdiffusion 24 -40 24 -40 0 cellNo=213
rlabel pdiffusion 31 -40 31 -40 0 cellNo=339
rlabel pdiffusion 38 -40 38 -40 0 cellNo=418
rlabel pdiffusion 45 -40 45 -40 0 cellNo=631
rlabel pdiffusion 52 -40 52 -40 0 cellNo=731
rlabel pdiffusion 80 -40 80 -40 0 cellNo=254
rlabel pdiffusion 136 -40 136 -40 0 feedthrough
rlabel pdiffusion 143 -40 143 -40 0 cellNo=510
rlabel pdiffusion 150 -40 150 -40 0 cellNo=400
rlabel pdiffusion 157 -40 157 -40 0 feedthrough
rlabel pdiffusion 171 -40 171 -40 0 cellNo=210
rlabel pdiffusion 185 -40 185 -40 0 feedthrough
rlabel pdiffusion 192 -40 192 -40 0 cellNo=330
rlabel pdiffusion 213 -40 213 -40 0 cellNo=969
rlabel pdiffusion 220 -40 220 -40 0 cellNo=888
rlabel pdiffusion 227 -40 227 -40 0 cellNo=137
rlabel pdiffusion 234 -40 234 -40 0 feedthrough
rlabel pdiffusion 241 -40 241 -40 0 cellNo=302
rlabel pdiffusion 248 -40 248 -40 0 cellNo=537
rlabel pdiffusion 255 -40 255 -40 0 feedthrough
rlabel pdiffusion 262 -40 262 -40 0 feedthrough
rlabel pdiffusion 269 -40 269 -40 0 cellNo=110
rlabel pdiffusion 276 -40 276 -40 0 feedthrough
rlabel pdiffusion 283 -40 283 -40 0 feedthrough
rlabel pdiffusion 290 -40 290 -40 0 cellNo=163
rlabel pdiffusion 297 -40 297 -40 0 feedthrough
rlabel pdiffusion 304 -40 304 -40 0 cellNo=957
rlabel pdiffusion 311 -40 311 -40 0 cellNo=59
rlabel pdiffusion 318 -40 318 -40 0 feedthrough
rlabel pdiffusion 325 -40 325 -40 0 feedthrough
rlabel pdiffusion 332 -40 332 -40 0 cellNo=598
rlabel pdiffusion 479 -40 479 -40 0 cellNo=41
rlabel pdiffusion 486 -40 486 -40 0 feedthrough
rlabel pdiffusion 577 -40 577 -40 0 cellNo=300
rlabel pdiffusion 584 -40 584 -40 0 feedthrough
rlabel pdiffusion 3 -63 3 -63 0 cellNo=95
rlabel pdiffusion 10 -63 10 -63 0 cellNo=855
rlabel pdiffusion 17 -63 17 -63 0 cellNo=161
rlabel pdiffusion 24 -63 24 -63 0 cellNo=315
rlabel pdiffusion 31 -63 31 -63 0 cellNo=388
rlabel pdiffusion 38 -63 38 -63 0 cellNo=697
rlabel pdiffusion 45 -63 45 -63 0 cellNo=496
rlabel pdiffusion 52 -63 52 -63 0 cellNo=704
rlabel pdiffusion 80 -63 80 -63 0 cellNo=117
rlabel pdiffusion 143 -63 143 -63 0 cellNo=165
rlabel pdiffusion 150 -63 150 -63 0 feedthrough
rlabel pdiffusion 157 -63 157 -63 0 feedthrough
rlabel pdiffusion 171 -63 171 -63 0 feedthrough
rlabel pdiffusion 178 -63 178 -63 0 cellNo=712
rlabel pdiffusion 185 -63 185 -63 0 cellNo=234
rlabel pdiffusion 192 -63 192 -63 0 cellNo=518
rlabel pdiffusion 199 -63 199 -63 0 cellNo=204
rlabel pdiffusion 206 -63 206 -63 0 feedthrough
rlabel pdiffusion 213 -63 213 -63 0 cellNo=187
rlabel pdiffusion 220 -63 220 -63 0 feedthrough
rlabel pdiffusion 227 -63 227 -63 0 feedthrough
rlabel pdiffusion 234 -63 234 -63 0 cellNo=591
rlabel pdiffusion 241 -63 241 -63 0 cellNo=755
rlabel pdiffusion 248 -63 248 -63 0 cellNo=160
rlabel pdiffusion 255 -63 255 -63 0 feedthrough
rlabel pdiffusion 262 -63 262 -63 0 feedthrough
rlabel pdiffusion 269 -63 269 -63 0 feedthrough
rlabel pdiffusion 276 -63 276 -63 0 feedthrough
rlabel pdiffusion 283 -63 283 -63 0 cellNo=235
rlabel pdiffusion 290 -63 290 -63 0 feedthrough
rlabel pdiffusion 297 -63 297 -63 0 feedthrough
rlabel pdiffusion 304 -63 304 -63 0 cellNo=195
rlabel pdiffusion 311 -63 311 -63 0 cellNo=186
rlabel pdiffusion 318 -63 318 -63 0 cellNo=558
rlabel pdiffusion 325 -63 325 -63 0 feedthrough
rlabel pdiffusion 339 -63 339 -63 0 cellNo=520
rlabel pdiffusion 346 -63 346 -63 0 feedthrough
rlabel pdiffusion 353 -63 353 -63 0 feedthrough
rlabel pdiffusion 360 -63 360 -63 0 cellNo=584
rlabel pdiffusion 465 -63 465 -63 0 cellNo=2
rlabel pdiffusion 472 -63 472 -63 0 feedthrough
rlabel pdiffusion 479 -63 479 -63 0 feedthrough
rlabel pdiffusion 577 -63 577 -63 0 feedthrough
rlabel pdiffusion 3 -86 3 -86 0 cellNo=151
rlabel pdiffusion 10 -86 10 -86 0 cellNo=498
rlabel pdiffusion 17 -86 17 -86 0 cellNo=301
rlabel pdiffusion 24 -86 24 -86 0 cellNo=741
rlabel pdiffusion 31 -86 31 -86 0 cellNo=458
rlabel pdiffusion 38 -86 38 -86 0 cellNo=506
rlabel pdiffusion 45 -86 45 -86 0 cellNo=670
rlabel pdiffusion 122 -86 122 -86 0 cellNo=497
rlabel pdiffusion 136 -86 136 -86 0 cellNo=843
rlabel pdiffusion 143 -86 143 -86 0 feedthrough
rlabel pdiffusion 150 -86 150 -86 0 feedthrough
rlabel pdiffusion 157 -86 157 -86 0 cellNo=437
rlabel pdiffusion 164 -86 164 -86 0 cellNo=789
rlabel pdiffusion 171 -86 171 -86 0 feedthrough
rlabel pdiffusion 178 -86 178 -86 0 feedthrough
rlabel pdiffusion 185 -86 185 -86 0 cellNo=870
rlabel pdiffusion 192 -86 192 -86 0 cellNo=264
rlabel pdiffusion 199 -86 199 -86 0 cellNo=154
rlabel pdiffusion 206 -86 206 -86 0 cellNo=49
rlabel pdiffusion 213 -86 213 -86 0 feedthrough
rlabel pdiffusion 220 -86 220 -86 0 feedthrough
rlabel pdiffusion 227 -86 227 -86 0 feedthrough
rlabel pdiffusion 234 -86 234 -86 0 feedthrough
rlabel pdiffusion 241 -86 241 -86 0 cellNo=214
rlabel pdiffusion 248 -86 248 -86 0 feedthrough
rlabel pdiffusion 255 -86 255 -86 0 feedthrough
rlabel pdiffusion 262 -86 262 -86 0 feedthrough
rlabel pdiffusion 269 -86 269 -86 0 cellNo=875
rlabel pdiffusion 276 -86 276 -86 0 cellNo=175
rlabel pdiffusion 283 -86 283 -86 0 feedthrough
rlabel pdiffusion 290 -86 290 -86 0 cellNo=416
rlabel pdiffusion 297 -86 297 -86 0 feedthrough
rlabel pdiffusion 304 -86 304 -86 0 cellNo=48
rlabel pdiffusion 311 -86 311 -86 0 cellNo=367
rlabel pdiffusion 318 -86 318 -86 0 feedthrough
rlabel pdiffusion 325 -86 325 -86 0 cellNo=152
rlabel pdiffusion 339 -86 339 -86 0 feedthrough
rlabel pdiffusion 346 -86 346 -86 0 cellNo=206
rlabel pdiffusion 353 -86 353 -86 0 feedthrough
rlabel pdiffusion 472 -86 472 -86 0 cellNo=471
rlabel pdiffusion 479 -86 479 -86 0 feedthrough
rlabel pdiffusion 486 -86 486 -86 0 feedthrough
rlabel pdiffusion 577 -86 577 -86 0 feedthrough
rlabel pdiffusion 3 -117 3 -117 0 cellNo=109
rlabel pdiffusion 10 -117 10 -117 0 cellNo=294
rlabel pdiffusion 17 -117 17 -117 0 cellNo=377
rlabel pdiffusion 24 -117 24 -117 0 cellNo=456
rlabel pdiffusion 31 -117 31 -117 0 cellNo=485
rlabel pdiffusion 38 -117 38 -117 0 cellNo=650
rlabel pdiffusion 108 -117 108 -117 0 feedthrough
rlabel pdiffusion 122 -117 122 -117 0 cellNo=230
rlabel pdiffusion 129 -117 129 -117 0 cellNo=714
rlabel pdiffusion 136 -117 136 -117 0 feedthrough
rlabel pdiffusion 143 -117 143 -117 0 cellNo=326
rlabel pdiffusion 150 -117 150 -117 0 cellNo=261
rlabel pdiffusion 157 -117 157 -117 0 feedthrough
rlabel pdiffusion 164 -117 164 -117 0 feedthrough
rlabel pdiffusion 171 -117 171 -117 0 cellNo=547
rlabel pdiffusion 178 -117 178 -117 0 cellNo=107
rlabel pdiffusion 185 -117 185 -117 0 feedthrough
rlabel pdiffusion 192 -117 192 -117 0 feedthrough
rlabel pdiffusion 199 -117 199 -117 0 feedthrough
rlabel pdiffusion 206 -117 206 -117 0 cellNo=188
rlabel pdiffusion 213 -117 213 -117 0 cellNo=14
rlabel pdiffusion 220 -117 220 -117 0 cellNo=27
rlabel pdiffusion 227 -117 227 -117 0 feedthrough
rlabel pdiffusion 234 -117 234 -117 0 feedthrough
rlabel pdiffusion 241 -117 241 -117 0 cellNo=153
rlabel pdiffusion 248 -117 248 -117 0 cellNo=43
rlabel pdiffusion 255 -117 255 -117 0 cellNo=548
rlabel pdiffusion 262 -117 262 -117 0 feedthrough
rlabel pdiffusion 269 -117 269 -117 0 feedthrough
rlabel pdiffusion 276 -117 276 -117 0 cellNo=325
rlabel pdiffusion 283 -117 283 -117 0 feedthrough
rlabel pdiffusion 290 -117 290 -117 0 feedthrough
rlabel pdiffusion 297 -117 297 -117 0 feedthrough
rlabel pdiffusion 304 -117 304 -117 0 feedthrough
rlabel pdiffusion 311 -117 311 -117 0 feedthrough
rlabel pdiffusion 318 -117 318 -117 0 cellNo=845
rlabel pdiffusion 325 -117 325 -117 0 feedthrough
rlabel pdiffusion 332 -117 332 -117 0 feedthrough
rlabel pdiffusion 339 -117 339 -117 0 cellNo=236
rlabel pdiffusion 346 -117 346 -117 0 feedthrough
rlabel pdiffusion 353 -117 353 -117 0 feedthrough
rlabel pdiffusion 360 -117 360 -117 0 feedthrough
rlabel pdiffusion 367 -117 367 -117 0 feedthrough
rlabel pdiffusion 374 -117 374 -117 0 feedthrough
rlabel pdiffusion 381 -117 381 -117 0 feedthrough
rlabel pdiffusion 395 -117 395 -117 0 cellNo=964
rlabel pdiffusion 423 -117 423 -117 0 feedthrough
rlabel pdiffusion 479 -117 479 -117 0 cellNo=460
rlabel pdiffusion 486 -117 486 -117 0 feedthrough
rlabel pdiffusion 493 -117 493 -117 0 feedthrough
rlabel pdiffusion 577 -117 577 -117 0 cellNo=433
rlabel pdiffusion 584 -117 584 -117 0 feedthrough
rlabel pdiffusion 591 -117 591 -117 0 feedthrough
rlabel pdiffusion 3 -156 3 -156 0 cellNo=292
rlabel pdiffusion 10 -156 10 -156 0 cellNo=357
rlabel pdiffusion 17 -156 17 -156 0 cellNo=444
rlabel pdiffusion 24 -156 24 -156 0 cellNo=473
rlabel pdiffusion 31 -156 31 -156 0 cellNo=943
rlabel pdiffusion 66 -156 66 -156 0 feedthrough
rlabel pdiffusion 73 -156 73 -156 0 feedthrough
rlabel pdiffusion 80 -156 80 -156 0 cellNo=440
rlabel pdiffusion 87 -156 87 -156 0 feedthrough
rlabel pdiffusion 94 -156 94 -156 0 feedthrough
rlabel pdiffusion 101 -156 101 -156 0 cellNo=233
rlabel pdiffusion 108 -156 108 -156 0 feedthrough
rlabel pdiffusion 115 -156 115 -156 0 cellNo=493
rlabel pdiffusion 122 -156 122 -156 0 cellNo=740
rlabel pdiffusion 129 -156 129 -156 0 cellNo=465
rlabel pdiffusion 136 -156 136 -156 0 feedthrough
rlabel pdiffusion 143 -156 143 -156 0 cellNo=443
rlabel pdiffusion 150 -156 150 -156 0 feedthrough
rlabel pdiffusion 157 -156 157 -156 0 feedthrough
rlabel pdiffusion 164 -156 164 -156 0 cellNo=144
rlabel pdiffusion 171 -156 171 -156 0 feedthrough
rlabel pdiffusion 178 -156 178 -156 0 feedthrough
rlabel pdiffusion 185 -156 185 -156 0 feedthrough
rlabel pdiffusion 192 -156 192 -156 0 feedthrough
rlabel pdiffusion 199 -156 199 -156 0 feedthrough
rlabel pdiffusion 206 -156 206 -156 0 cellNo=765
rlabel pdiffusion 213 -156 213 -156 0 cellNo=472
rlabel pdiffusion 220 -156 220 -156 0 cellNo=962
rlabel pdiffusion 227 -156 227 -156 0 cellNo=24
rlabel pdiffusion 234 -156 234 -156 0 cellNo=639
rlabel pdiffusion 241 -156 241 -156 0 cellNo=174
rlabel pdiffusion 248 -156 248 -156 0 feedthrough
rlabel pdiffusion 255 -156 255 -156 0 feedthrough
rlabel pdiffusion 262 -156 262 -156 0 cellNo=239
rlabel pdiffusion 269 -156 269 -156 0 feedthrough
rlabel pdiffusion 276 -156 276 -156 0 feedthrough
rlabel pdiffusion 283 -156 283 -156 0 cellNo=52
rlabel pdiffusion 290 -156 290 -156 0 feedthrough
rlabel pdiffusion 297 -156 297 -156 0 cellNo=130
rlabel pdiffusion 304 -156 304 -156 0 feedthrough
rlabel pdiffusion 311 -156 311 -156 0 feedthrough
rlabel pdiffusion 318 -156 318 -156 0 feedthrough
rlabel pdiffusion 325 -156 325 -156 0 feedthrough
rlabel pdiffusion 332 -156 332 -156 0 cellNo=651
rlabel pdiffusion 339 -156 339 -156 0 feedthrough
rlabel pdiffusion 346 -156 346 -156 0 feedthrough
rlabel pdiffusion 353 -156 353 -156 0 cellNo=259
rlabel pdiffusion 360 -156 360 -156 0 feedthrough
rlabel pdiffusion 367 -156 367 -156 0 feedthrough
rlabel pdiffusion 374 -156 374 -156 0 feedthrough
rlabel pdiffusion 381 -156 381 -156 0 feedthrough
rlabel pdiffusion 388 -156 388 -156 0 cellNo=720
rlabel pdiffusion 395 -156 395 -156 0 feedthrough
rlabel pdiffusion 402 -156 402 -156 0 feedthrough
rlabel pdiffusion 409 -156 409 -156 0 cellNo=362
rlabel pdiffusion 416 -156 416 -156 0 feedthrough
rlabel pdiffusion 423 -156 423 -156 0 feedthrough
rlabel pdiffusion 430 -156 430 -156 0 feedthrough
rlabel pdiffusion 437 -156 437 -156 0 feedthrough
rlabel pdiffusion 444 -156 444 -156 0 feedthrough
rlabel pdiffusion 500 -156 500 -156 0 feedthrough
rlabel pdiffusion 591 -156 591 -156 0 feedthrough
rlabel pdiffusion 3 -205 3 -205 0 cellNo=758
rlabel pdiffusion 10 -205 10 -205 0 cellNo=247
rlabel pdiffusion 17 -205 17 -205 0 cellNo=511
rlabel pdiffusion 24 -205 24 -205 0 cellNo=250
rlabel pdiffusion 31 -205 31 -205 0 cellNo=947
rlabel pdiffusion 80 -205 80 -205 0 feedthrough
rlabel pdiffusion 87 -205 87 -205 0 feedthrough
rlabel pdiffusion 94 -205 94 -205 0 cellNo=328
rlabel pdiffusion 101 -205 101 -205 0 feedthrough
rlabel pdiffusion 108 -205 108 -205 0 feedthrough
rlabel pdiffusion 115 -205 115 -205 0 feedthrough
rlabel pdiffusion 122 -205 122 -205 0 cellNo=515
rlabel pdiffusion 129 -205 129 -205 0 feedthrough
rlabel pdiffusion 136 -205 136 -205 0 feedthrough
rlabel pdiffusion 143 -205 143 -205 0 cellNo=406
rlabel pdiffusion 150 -205 150 -205 0 feedthrough
rlabel pdiffusion 157 -205 157 -205 0 cellNo=322
rlabel pdiffusion 164 -205 164 -205 0 cellNo=348
rlabel pdiffusion 171 -205 171 -205 0 cellNo=607
rlabel pdiffusion 178 -205 178 -205 0 cellNo=342
rlabel pdiffusion 185 -205 185 -205 0 cellNo=283
rlabel pdiffusion 192 -205 192 -205 0 cellNo=792
rlabel pdiffusion 199 -205 199 -205 0 cellNo=483
rlabel pdiffusion 206 -205 206 -205 0 feedthrough
rlabel pdiffusion 213 -205 213 -205 0 cellNo=262
rlabel pdiffusion 220 -205 220 -205 0 cellNo=652
rlabel pdiffusion 227 -205 227 -205 0 cellNo=838
rlabel pdiffusion 234 -205 234 -205 0 cellNo=286
rlabel pdiffusion 241 -205 241 -205 0 cellNo=517
rlabel pdiffusion 248 -205 248 -205 0 feedthrough
rlabel pdiffusion 255 -205 255 -205 0 feedthrough
rlabel pdiffusion 262 -205 262 -205 0 feedthrough
rlabel pdiffusion 269 -205 269 -205 0 feedthrough
rlabel pdiffusion 276 -205 276 -205 0 cellNo=955
rlabel pdiffusion 283 -205 283 -205 0 feedthrough
rlabel pdiffusion 290 -205 290 -205 0 cellNo=612
rlabel pdiffusion 297 -205 297 -205 0 cellNo=69
rlabel pdiffusion 304 -205 304 -205 0 feedthrough
rlabel pdiffusion 311 -205 311 -205 0 feedthrough
rlabel pdiffusion 318 -205 318 -205 0 cellNo=904
rlabel pdiffusion 325 -205 325 -205 0 feedthrough
rlabel pdiffusion 332 -205 332 -205 0 feedthrough
rlabel pdiffusion 339 -205 339 -205 0 feedthrough
rlabel pdiffusion 346 -205 346 -205 0 feedthrough
rlabel pdiffusion 353 -205 353 -205 0 feedthrough
rlabel pdiffusion 360 -205 360 -205 0 feedthrough
rlabel pdiffusion 367 -205 367 -205 0 feedthrough
rlabel pdiffusion 374 -205 374 -205 0 feedthrough
rlabel pdiffusion 381 -205 381 -205 0 feedthrough
rlabel pdiffusion 388 -205 388 -205 0 feedthrough
rlabel pdiffusion 395 -205 395 -205 0 feedthrough
rlabel pdiffusion 402 -205 402 -205 0 feedthrough
rlabel pdiffusion 409 -205 409 -205 0 feedthrough
rlabel pdiffusion 416 -205 416 -205 0 feedthrough
rlabel pdiffusion 423 -205 423 -205 0 cellNo=653
rlabel pdiffusion 430 -205 430 -205 0 feedthrough
rlabel pdiffusion 437 -205 437 -205 0 feedthrough
rlabel pdiffusion 444 -205 444 -205 0 feedthrough
rlabel pdiffusion 451 -205 451 -205 0 cellNo=784
rlabel pdiffusion 458 -205 458 -205 0 cellNo=93
rlabel pdiffusion 465 -205 465 -205 0 feedthrough
rlabel pdiffusion 507 -205 507 -205 0 feedthrough
rlabel pdiffusion 591 -205 591 -205 0 feedthrough
rlabel pdiffusion 3 -246 3 -246 0 cellNo=407
rlabel pdiffusion 10 -246 10 -246 0 cellNo=694
rlabel pdiffusion 17 -246 17 -246 0 cellNo=643
rlabel pdiffusion 24 -246 24 -246 0 cellNo=934
rlabel pdiffusion 115 -246 115 -246 0 feedthrough
rlabel pdiffusion 122 -246 122 -246 0 cellNo=281
rlabel pdiffusion 129 -246 129 -246 0 feedthrough
rlabel pdiffusion 136 -246 136 -246 0 feedthrough
rlabel pdiffusion 143 -246 143 -246 0 feedthrough
rlabel pdiffusion 150 -246 150 -246 0 feedthrough
rlabel pdiffusion 157 -246 157 -246 0 cellNo=529
rlabel pdiffusion 164 -246 164 -246 0 feedthrough
rlabel pdiffusion 171 -246 171 -246 0 cellNo=899
rlabel pdiffusion 178 -246 178 -246 0 feedthrough
rlabel pdiffusion 185 -246 185 -246 0 feedthrough
rlabel pdiffusion 192 -246 192 -246 0 feedthrough
rlabel pdiffusion 199 -246 199 -246 0 feedthrough
rlabel pdiffusion 206 -246 206 -246 0 cellNo=750
rlabel pdiffusion 213 -246 213 -246 0 cellNo=291
rlabel pdiffusion 220 -246 220 -246 0 cellNo=887
rlabel pdiffusion 227 -246 227 -246 0 cellNo=54
rlabel pdiffusion 234 -246 234 -246 0 cellNo=402
rlabel pdiffusion 241 -246 241 -246 0 cellNo=563
rlabel pdiffusion 248 -246 248 -246 0 feedthrough
rlabel pdiffusion 255 -246 255 -246 0 feedthrough
rlabel pdiffusion 262 -246 262 -246 0 cellNo=97
rlabel pdiffusion 269 -246 269 -246 0 feedthrough
rlabel pdiffusion 276 -246 276 -246 0 cellNo=699
rlabel pdiffusion 283 -246 283 -246 0 feedthrough
rlabel pdiffusion 290 -246 290 -246 0 cellNo=689
rlabel pdiffusion 297 -246 297 -246 0 cellNo=953
rlabel pdiffusion 304 -246 304 -246 0 feedthrough
rlabel pdiffusion 311 -246 311 -246 0 feedthrough
rlabel pdiffusion 318 -246 318 -246 0 cellNo=861
rlabel pdiffusion 325 -246 325 -246 0 feedthrough
rlabel pdiffusion 332 -246 332 -246 0 feedthrough
rlabel pdiffusion 339 -246 339 -246 0 feedthrough
rlabel pdiffusion 346 -246 346 -246 0 cellNo=164
rlabel pdiffusion 353 -246 353 -246 0 feedthrough
rlabel pdiffusion 360 -246 360 -246 0 feedthrough
rlabel pdiffusion 367 -246 367 -246 0 cellNo=25
rlabel pdiffusion 374 -246 374 -246 0 feedthrough
rlabel pdiffusion 381 -246 381 -246 0 cellNo=884
rlabel pdiffusion 388 -246 388 -246 0 feedthrough
rlabel pdiffusion 395 -246 395 -246 0 feedthrough
rlabel pdiffusion 402 -246 402 -246 0 feedthrough
rlabel pdiffusion 409 -246 409 -246 0 feedthrough
rlabel pdiffusion 416 -246 416 -246 0 feedthrough
rlabel pdiffusion 423 -246 423 -246 0 feedthrough
rlabel pdiffusion 430 -246 430 -246 0 feedthrough
rlabel pdiffusion 437 -246 437 -246 0 feedthrough
rlabel pdiffusion 444 -246 444 -246 0 feedthrough
rlabel pdiffusion 451 -246 451 -246 0 feedthrough
rlabel pdiffusion 458 -246 458 -246 0 cellNo=70
rlabel pdiffusion 465 -246 465 -246 0 cellNo=524
rlabel pdiffusion 507 -246 507 -246 0 cellNo=4
rlabel pdiffusion 563 -246 563 -246 0 cellNo=157
rlabel pdiffusion 570 -246 570 -246 0 cellNo=775
rlabel pdiffusion 591 -246 591 -246 0 feedthrough
rlabel pdiffusion 598 -246 598 -246 0 cellNo=211
rlabel pdiffusion 647 -246 647 -246 0 cellNo=44
rlabel pdiffusion 3 -287 3 -287 0 cellNo=470
rlabel pdiffusion 10 -287 10 -287 0 cellNo=642
rlabel pdiffusion 17 -287 17 -287 0 cellNo=897
rlabel pdiffusion 66 -287 66 -287 0 cellNo=425
rlabel pdiffusion 73 -287 73 -287 0 cellNo=145
rlabel pdiffusion 80 -287 80 -287 0 feedthrough
rlabel pdiffusion 87 -287 87 -287 0 feedthrough
rlabel pdiffusion 94 -287 94 -287 0 feedthrough
rlabel pdiffusion 101 -287 101 -287 0 cellNo=238
rlabel pdiffusion 108 -287 108 -287 0 feedthrough
rlabel pdiffusion 115 -287 115 -287 0 cellNo=569
rlabel pdiffusion 122 -287 122 -287 0 cellNo=580
rlabel pdiffusion 129 -287 129 -287 0 feedthrough
rlabel pdiffusion 136 -287 136 -287 0 feedthrough
rlabel pdiffusion 143 -287 143 -287 0 feedthrough
rlabel pdiffusion 150 -287 150 -287 0 feedthrough
rlabel pdiffusion 157 -287 157 -287 0 feedthrough
rlabel pdiffusion 164 -287 164 -287 0 feedthrough
rlabel pdiffusion 171 -287 171 -287 0 cellNo=386
rlabel pdiffusion 178 -287 178 -287 0 feedthrough
rlabel pdiffusion 185 -287 185 -287 0 cellNo=141
rlabel pdiffusion 192 -287 192 -287 0 cellNo=159
rlabel pdiffusion 199 -287 199 -287 0 cellNo=649
rlabel pdiffusion 206 -287 206 -287 0 cellNo=488
rlabel pdiffusion 213 -287 213 -287 0 cellNo=306
rlabel pdiffusion 220 -287 220 -287 0 feedthrough
rlabel pdiffusion 227 -287 227 -287 0 feedthrough
rlabel pdiffusion 234 -287 234 -287 0 cellNo=29
rlabel pdiffusion 241 -287 241 -287 0 cellNo=533
rlabel pdiffusion 248 -287 248 -287 0 feedthrough
rlabel pdiffusion 255 -287 255 -287 0 cellNo=900
rlabel pdiffusion 262 -287 262 -287 0 feedthrough
rlabel pdiffusion 269 -287 269 -287 0 feedthrough
rlabel pdiffusion 276 -287 276 -287 0 feedthrough
rlabel pdiffusion 283 -287 283 -287 0 cellNo=577
rlabel pdiffusion 290 -287 290 -287 0 cellNo=430
rlabel pdiffusion 297 -287 297 -287 0 cellNo=596
rlabel pdiffusion 304 -287 304 -287 0 cellNo=940
rlabel pdiffusion 311 -287 311 -287 0 cellNo=237
rlabel pdiffusion 318 -287 318 -287 0 cellNo=104
rlabel pdiffusion 325 -287 325 -287 0 cellNo=732
rlabel pdiffusion 332 -287 332 -287 0 feedthrough
rlabel pdiffusion 339 -287 339 -287 0 cellNo=587
rlabel pdiffusion 346 -287 346 -287 0 feedthrough
rlabel pdiffusion 353 -287 353 -287 0 feedthrough
rlabel pdiffusion 360 -287 360 -287 0 feedthrough
rlabel pdiffusion 367 -287 367 -287 0 feedthrough
rlabel pdiffusion 374 -287 374 -287 0 feedthrough
rlabel pdiffusion 381 -287 381 -287 0 cellNo=82
rlabel pdiffusion 388 -287 388 -287 0 feedthrough
rlabel pdiffusion 395 -287 395 -287 0 cellNo=215
rlabel pdiffusion 402 -287 402 -287 0 feedthrough
rlabel pdiffusion 409 -287 409 -287 0 feedthrough
rlabel pdiffusion 416 -287 416 -287 0 feedthrough
rlabel pdiffusion 423 -287 423 -287 0 feedthrough
rlabel pdiffusion 430 -287 430 -287 0 feedthrough
rlabel pdiffusion 437 -287 437 -287 0 feedthrough
rlabel pdiffusion 444 -287 444 -287 0 feedthrough
rlabel pdiffusion 451 -287 451 -287 0 feedthrough
rlabel pdiffusion 458 -287 458 -287 0 feedthrough
rlabel pdiffusion 465 -287 465 -287 0 feedthrough
rlabel pdiffusion 472 -287 472 -287 0 feedthrough
rlabel pdiffusion 479 -287 479 -287 0 feedthrough
rlabel pdiffusion 486 -287 486 -287 0 feedthrough
rlabel pdiffusion 493 -287 493 -287 0 feedthrough
rlabel pdiffusion 500 -287 500 -287 0 cellNo=627
rlabel pdiffusion 507 -287 507 -287 0 feedthrough
rlabel pdiffusion 521 -287 521 -287 0 feedthrough
rlabel pdiffusion 528 -287 528 -287 0 feedthrough
rlabel pdiffusion 563 -287 563 -287 0 feedthrough
rlabel pdiffusion 612 -287 612 -287 0 feedthrough
rlabel pdiffusion 647 -287 647 -287 0 feedthrough
rlabel pdiffusion 3 -336 3 -336 0 cellNo=633
rlabel pdiffusion 10 -336 10 -336 0 cellNo=877
rlabel pdiffusion 73 -336 73 -336 0 cellNo=528
rlabel pdiffusion 80 -336 80 -336 0 feedthrough
rlabel pdiffusion 87 -336 87 -336 0 feedthrough
rlabel pdiffusion 94 -336 94 -336 0 feedthrough
rlabel pdiffusion 101 -336 101 -336 0 feedthrough
rlabel pdiffusion 108 -336 108 -336 0 feedthrough
rlabel pdiffusion 115 -336 115 -336 0 feedthrough
rlabel pdiffusion 122 -336 122 -336 0 feedthrough
rlabel pdiffusion 129 -336 129 -336 0 cellNo=804
rlabel pdiffusion 136 -336 136 -336 0 feedthrough
rlabel pdiffusion 143 -336 143 -336 0 feedthrough
rlabel pdiffusion 150 -336 150 -336 0 cellNo=111
rlabel pdiffusion 157 -336 157 -336 0 cellNo=932
rlabel pdiffusion 164 -336 164 -336 0 cellNo=277
rlabel pdiffusion 171 -336 171 -336 0 feedthrough
rlabel pdiffusion 178 -336 178 -336 0 feedthrough
rlabel pdiffusion 185 -336 185 -336 0 cellNo=759
rlabel pdiffusion 192 -336 192 -336 0 feedthrough
rlabel pdiffusion 199 -336 199 -336 0 feedthrough
rlabel pdiffusion 206 -336 206 -336 0 feedthrough
rlabel pdiffusion 213 -336 213 -336 0 feedthrough
rlabel pdiffusion 220 -336 220 -336 0 cellNo=805
rlabel pdiffusion 227 -336 227 -336 0 cellNo=681
rlabel pdiffusion 234 -336 234 -336 0 cellNo=98
rlabel pdiffusion 241 -336 241 -336 0 feedthrough
rlabel pdiffusion 248 -336 248 -336 0 feedthrough
rlabel pdiffusion 255 -336 255 -336 0 feedthrough
rlabel pdiffusion 262 -336 262 -336 0 cellNo=176
rlabel pdiffusion 269 -336 269 -336 0 cellNo=12
rlabel pdiffusion 276 -336 276 -336 0 feedthrough
rlabel pdiffusion 283 -336 283 -336 0 cellNo=398
rlabel pdiffusion 290 -336 290 -336 0 feedthrough
rlabel pdiffusion 297 -336 297 -336 0 feedthrough
rlabel pdiffusion 304 -336 304 -336 0 feedthrough
rlabel pdiffusion 311 -336 311 -336 0 cellNo=65
rlabel pdiffusion 318 -336 318 -336 0 feedthrough
rlabel pdiffusion 325 -336 325 -336 0 cellNo=190
rlabel pdiffusion 332 -336 332 -336 0 feedthrough
rlabel pdiffusion 339 -336 339 -336 0 cellNo=149
rlabel pdiffusion 346 -336 346 -336 0 cellNo=771
rlabel pdiffusion 353 -336 353 -336 0 feedthrough
rlabel pdiffusion 360 -336 360 -336 0 cellNo=37
rlabel pdiffusion 367 -336 367 -336 0 cellNo=655
rlabel pdiffusion 374 -336 374 -336 0 feedthrough
rlabel pdiffusion 381 -336 381 -336 0 feedthrough
rlabel pdiffusion 388 -336 388 -336 0 cellNo=30
rlabel pdiffusion 395 -336 395 -336 0 feedthrough
rlabel pdiffusion 402 -336 402 -336 0 feedthrough
rlabel pdiffusion 409 -336 409 -336 0 cellNo=106
rlabel pdiffusion 416 -336 416 -336 0 feedthrough
rlabel pdiffusion 423 -336 423 -336 0 cellNo=514
rlabel pdiffusion 430 -336 430 -336 0 feedthrough
rlabel pdiffusion 437 -336 437 -336 0 feedthrough
rlabel pdiffusion 444 -336 444 -336 0 feedthrough
rlabel pdiffusion 451 -336 451 -336 0 feedthrough
rlabel pdiffusion 458 -336 458 -336 0 feedthrough
rlabel pdiffusion 465 -336 465 -336 0 feedthrough
rlabel pdiffusion 472 -336 472 -336 0 feedthrough
rlabel pdiffusion 479 -336 479 -336 0 feedthrough
rlabel pdiffusion 486 -336 486 -336 0 feedthrough
rlabel pdiffusion 493 -336 493 -336 0 feedthrough
rlabel pdiffusion 500 -336 500 -336 0 feedthrough
rlabel pdiffusion 507 -336 507 -336 0 feedthrough
rlabel pdiffusion 514 -336 514 -336 0 cellNo=455
rlabel pdiffusion 521 -336 521 -336 0 feedthrough
rlabel pdiffusion 528 -336 528 -336 0 feedthrough
rlabel pdiffusion 535 -336 535 -336 0 feedthrough
rlabel pdiffusion 542 -336 542 -336 0 cellNo=595
rlabel pdiffusion 549 -336 549 -336 0 feedthrough
rlabel pdiffusion 556 -336 556 -336 0 cellNo=613
rlabel pdiffusion 563 -336 563 -336 0 feedthrough
rlabel pdiffusion 605 -336 605 -336 0 feedthrough
rlabel pdiffusion 647 -336 647 -336 0 cellNo=635
rlabel pdiffusion 654 -336 654 -336 0 feedthrough
rlabel pdiffusion 661 -336 661 -336 0 feedthrough
rlabel pdiffusion 675 -336 675 -336 0 feedthrough
rlabel pdiffusion 682 -336 682 -336 0 cellNo=892
rlabel pdiffusion 3 -387 3 -387 0 cellNo=860
rlabel pdiffusion 31 -387 31 -387 0 cellNo=168
rlabel pdiffusion 45 -387 45 -387 0 feedthrough
rlabel pdiffusion 52 -387 52 -387 0 feedthrough
rlabel pdiffusion 59 -387 59 -387 0 feedthrough
rlabel pdiffusion 66 -387 66 -387 0 cellNo=492
rlabel pdiffusion 73 -387 73 -387 0 feedthrough
rlabel pdiffusion 80 -387 80 -387 0 feedthrough
rlabel pdiffusion 87 -387 87 -387 0 feedthrough
rlabel pdiffusion 94 -387 94 -387 0 feedthrough
rlabel pdiffusion 101 -387 101 -387 0 feedthrough
rlabel pdiffusion 108 -387 108 -387 0 cellNo=479
rlabel pdiffusion 115 -387 115 -387 0 feedthrough
rlabel pdiffusion 122 -387 122 -387 0 feedthrough
rlabel pdiffusion 129 -387 129 -387 0 feedthrough
rlabel pdiffusion 136 -387 136 -387 0 cellNo=560
rlabel pdiffusion 143 -387 143 -387 0 feedthrough
rlabel pdiffusion 150 -387 150 -387 0 cellNo=199
rlabel pdiffusion 157 -387 157 -387 0 cellNo=244
rlabel pdiffusion 164 -387 164 -387 0 cellNo=984
rlabel pdiffusion 171 -387 171 -387 0 feedthrough
rlabel pdiffusion 178 -387 178 -387 0 feedthrough
rlabel pdiffusion 185 -387 185 -387 0 feedthrough
rlabel pdiffusion 192 -387 192 -387 0 feedthrough
rlabel pdiffusion 199 -387 199 -387 0 feedthrough
rlabel pdiffusion 206 -387 206 -387 0 feedthrough
rlabel pdiffusion 213 -387 213 -387 0 cellNo=436
rlabel pdiffusion 220 -387 220 -387 0 cellNo=45
rlabel pdiffusion 227 -387 227 -387 0 cellNo=924
rlabel pdiffusion 234 -387 234 -387 0 cellNo=656
rlabel pdiffusion 241 -387 241 -387 0 cellNo=366
rlabel pdiffusion 248 -387 248 -387 0 feedthrough
rlabel pdiffusion 255 -387 255 -387 0 feedthrough
rlabel pdiffusion 262 -387 262 -387 0 feedthrough
rlabel pdiffusion 269 -387 269 -387 0 feedthrough
rlabel pdiffusion 276 -387 276 -387 0 cellNo=489
rlabel pdiffusion 283 -387 283 -387 0 feedthrough
rlabel pdiffusion 290 -387 290 -387 0 cellNo=158
rlabel pdiffusion 297 -387 297 -387 0 feedthrough
rlabel pdiffusion 304 -387 304 -387 0 feedthrough
rlabel pdiffusion 311 -387 311 -387 0 feedthrough
rlabel pdiffusion 318 -387 318 -387 0 feedthrough
rlabel pdiffusion 325 -387 325 -387 0 cellNo=223
rlabel pdiffusion 332 -387 332 -387 0 cellNo=474
rlabel pdiffusion 339 -387 339 -387 0 cellNo=28
rlabel pdiffusion 346 -387 346 -387 0 feedthrough
rlabel pdiffusion 353 -387 353 -387 0 cellNo=354
rlabel pdiffusion 360 -387 360 -387 0 cellNo=617
rlabel pdiffusion 367 -387 367 -387 0 feedthrough
rlabel pdiffusion 374 -387 374 -387 0 feedthrough
rlabel pdiffusion 381 -387 381 -387 0 feedthrough
rlabel pdiffusion 388 -387 388 -387 0 cellNo=432
rlabel pdiffusion 395 -387 395 -387 0 feedthrough
rlabel pdiffusion 402 -387 402 -387 0 feedthrough
rlabel pdiffusion 409 -387 409 -387 0 feedthrough
rlabel pdiffusion 416 -387 416 -387 0 feedthrough
rlabel pdiffusion 423 -387 423 -387 0 cellNo=954
rlabel pdiffusion 430 -387 430 -387 0 feedthrough
rlabel pdiffusion 437 -387 437 -387 0 feedthrough
rlabel pdiffusion 444 -387 444 -387 0 feedthrough
rlabel pdiffusion 451 -387 451 -387 0 cellNo=92
rlabel pdiffusion 458 -387 458 -387 0 cellNo=781
rlabel pdiffusion 465 -387 465 -387 0 feedthrough
rlabel pdiffusion 472 -387 472 -387 0 feedthrough
rlabel pdiffusion 479 -387 479 -387 0 feedthrough
rlabel pdiffusion 486 -387 486 -387 0 feedthrough
rlabel pdiffusion 493 -387 493 -387 0 feedthrough
rlabel pdiffusion 500 -387 500 -387 0 feedthrough
rlabel pdiffusion 507 -387 507 -387 0 feedthrough
rlabel pdiffusion 514 -387 514 -387 0 feedthrough
rlabel pdiffusion 521 -387 521 -387 0 cellNo=535
rlabel pdiffusion 528 -387 528 -387 0 feedthrough
rlabel pdiffusion 535 -387 535 -387 0 feedthrough
rlabel pdiffusion 542 -387 542 -387 0 feedthrough
rlabel pdiffusion 549 -387 549 -387 0 feedthrough
rlabel pdiffusion 556 -387 556 -387 0 feedthrough
rlabel pdiffusion 563 -387 563 -387 0 cellNo=303
rlabel pdiffusion 570 -387 570 -387 0 feedthrough
rlabel pdiffusion 577 -387 577 -387 0 feedthrough
rlabel pdiffusion 584 -387 584 -387 0 feedthrough
rlabel pdiffusion 591 -387 591 -387 0 feedthrough
rlabel pdiffusion 598 -387 598 -387 0 feedthrough
rlabel pdiffusion 605 -387 605 -387 0 feedthrough
rlabel pdiffusion 612 -387 612 -387 0 feedthrough
rlabel pdiffusion 619 -387 619 -387 0 feedthrough
rlabel pdiffusion 626 -387 626 -387 0 feedthrough
rlabel pdiffusion 633 -387 633 -387 0 feedthrough
rlabel pdiffusion 640 -387 640 -387 0 cellNo=184
rlabel pdiffusion 647 -387 647 -387 0 feedthrough
rlabel pdiffusion 654 -387 654 -387 0 feedthrough
rlabel pdiffusion 661 -387 661 -387 0 cellNo=345
rlabel pdiffusion 668 -387 668 -387 0 feedthrough
rlabel pdiffusion 675 -387 675 -387 0 cellNo=424
rlabel pdiffusion 682 -387 682 -387 0 feedthrough
rlabel pdiffusion 689 -387 689 -387 0 feedthrough
rlabel pdiffusion 3 -444 3 -444 0 feedthrough
rlabel pdiffusion 10 -444 10 -444 0 cellNo=491
rlabel pdiffusion 17 -444 17 -444 0 feedthrough
rlabel pdiffusion 24 -444 24 -444 0 feedthrough
rlabel pdiffusion 31 -444 31 -444 0 cellNo=40
rlabel pdiffusion 38 -444 38 -444 0 feedthrough
rlabel pdiffusion 45 -444 45 -444 0 feedthrough
rlabel pdiffusion 52 -444 52 -444 0 feedthrough
rlabel pdiffusion 59 -444 59 -444 0 feedthrough
rlabel pdiffusion 66 -444 66 -444 0 feedthrough
rlabel pdiffusion 73 -444 73 -444 0 feedthrough
rlabel pdiffusion 80 -444 80 -444 0 feedthrough
rlabel pdiffusion 87 -444 87 -444 0 cellNo=241
rlabel pdiffusion 94 -444 94 -444 0 feedthrough
rlabel pdiffusion 101 -444 101 -444 0 feedthrough
rlabel pdiffusion 108 -444 108 -444 0 feedthrough
rlabel pdiffusion 115 -444 115 -444 0 cellNo=191
rlabel pdiffusion 122 -444 122 -444 0 feedthrough
rlabel pdiffusion 129 -444 129 -444 0 feedthrough
rlabel pdiffusion 136 -444 136 -444 0 cellNo=88
rlabel pdiffusion 143 -444 143 -444 0 cellNo=324
rlabel pdiffusion 150 -444 150 -444 0 feedthrough
rlabel pdiffusion 157 -444 157 -444 0 cellNo=618
rlabel pdiffusion 164 -444 164 -444 0 feedthrough
rlabel pdiffusion 171 -444 171 -444 0 feedthrough
rlabel pdiffusion 178 -444 178 -444 0 cellNo=21
rlabel pdiffusion 185 -444 185 -444 0 cellNo=601
rlabel pdiffusion 192 -444 192 -444 0 feedthrough
rlabel pdiffusion 199 -444 199 -444 0 cellNo=992
rlabel pdiffusion 206 -444 206 -444 0 feedthrough
rlabel pdiffusion 213 -444 213 -444 0 cellNo=743
rlabel pdiffusion 220 -444 220 -444 0 feedthrough
rlabel pdiffusion 227 -444 227 -444 0 feedthrough
rlabel pdiffusion 234 -444 234 -444 0 cellNo=258
rlabel pdiffusion 241 -444 241 -444 0 cellNo=429
rlabel pdiffusion 248 -444 248 -444 0 feedthrough
rlabel pdiffusion 255 -444 255 -444 0 feedthrough
rlabel pdiffusion 262 -444 262 -444 0 feedthrough
rlabel pdiffusion 269 -444 269 -444 0 feedthrough
rlabel pdiffusion 276 -444 276 -444 0 feedthrough
rlabel pdiffusion 283 -444 283 -444 0 cellNo=403
rlabel pdiffusion 290 -444 290 -444 0 cellNo=198
rlabel pdiffusion 297 -444 297 -444 0 feedthrough
rlabel pdiffusion 304 -444 304 -444 0 cellNo=288
rlabel pdiffusion 311 -444 311 -444 0 feedthrough
rlabel pdiffusion 318 -444 318 -444 0 feedthrough
rlabel pdiffusion 325 -444 325 -444 0 cellNo=89
rlabel pdiffusion 332 -444 332 -444 0 feedthrough
rlabel pdiffusion 339 -444 339 -444 0 cellNo=298
rlabel pdiffusion 346 -444 346 -444 0 feedthrough
rlabel pdiffusion 353 -444 353 -444 0 feedthrough
rlabel pdiffusion 360 -444 360 -444 0 feedthrough
rlabel pdiffusion 367 -444 367 -444 0 cellNo=512
rlabel pdiffusion 374 -444 374 -444 0 cellNo=396
rlabel pdiffusion 381 -444 381 -444 0 feedthrough
rlabel pdiffusion 388 -444 388 -444 0 feedthrough
rlabel pdiffusion 395 -444 395 -444 0 cellNo=777
rlabel pdiffusion 402 -444 402 -444 0 cellNo=994
rlabel pdiffusion 409 -444 409 -444 0 cellNo=581
rlabel pdiffusion 416 -444 416 -444 0 feedthrough
rlabel pdiffusion 423 -444 423 -444 0 feedthrough
rlabel pdiffusion 430 -444 430 -444 0 feedthrough
rlabel pdiffusion 437 -444 437 -444 0 cellNo=851
rlabel pdiffusion 444 -444 444 -444 0 feedthrough
rlabel pdiffusion 451 -444 451 -444 0 feedthrough
rlabel pdiffusion 458 -444 458 -444 0 feedthrough
rlabel pdiffusion 465 -444 465 -444 0 cellNo=62
rlabel pdiffusion 472 -444 472 -444 0 feedthrough
rlabel pdiffusion 479 -444 479 -444 0 feedthrough
rlabel pdiffusion 486 -444 486 -444 0 feedthrough
rlabel pdiffusion 493 -444 493 -444 0 feedthrough
rlabel pdiffusion 500 -444 500 -444 0 feedthrough
rlabel pdiffusion 507 -444 507 -444 0 cellNo=658
rlabel pdiffusion 514 -444 514 -444 0 feedthrough
rlabel pdiffusion 521 -444 521 -444 0 feedthrough
rlabel pdiffusion 528 -444 528 -444 0 feedthrough
rlabel pdiffusion 535 -444 535 -444 0 feedthrough
rlabel pdiffusion 542 -444 542 -444 0 feedthrough
rlabel pdiffusion 549 -444 549 -444 0 feedthrough
rlabel pdiffusion 556 -444 556 -444 0 cellNo=574
rlabel pdiffusion 563 -444 563 -444 0 feedthrough
rlabel pdiffusion 570 -444 570 -444 0 feedthrough
rlabel pdiffusion 577 -444 577 -444 0 feedthrough
rlabel pdiffusion 584 -444 584 -444 0 feedthrough
rlabel pdiffusion 591 -444 591 -444 0 feedthrough
rlabel pdiffusion 598 -444 598 -444 0 feedthrough
rlabel pdiffusion 605 -444 605 -444 0 feedthrough
rlabel pdiffusion 612 -444 612 -444 0 feedthrough
rlabel pdiffusion 619 -444 619 -444 0 feedthrough
rlabel pdiffusion 626 -444 626 -444 0 cellNo=53
rlabel pdiffusion 633 -444 633 -444 0 cellNo=821
rlabel pdiffusion 640 -444 640 -444 0 feedthrough
rlabel pdiffusion 647 -444 647 -444 0 cellNo=201
rlabel pdiffusion 654 -444 654 -444 0 feedthrough
rlabel pdiffusion 661 -444 661 -444 0 cellNo=203
rlabel pdiffusion 668 -444 668 -444 0 feedthrough
rlabel pdiffusion 10 -501 10 -501 0 feedthrough
rlabel pdiffusion 17 -501 17 -501 0 feedthrough
rlabel pdiffusion 24 -501 24 -501 0 feedthrough
rlabel pdiffusion 31 -501 31 -501 0 feedthrough
rlabel pdiffusion 38 -501 38 -501 0 feedthrough
rlabel pdiffusion 45 -501 45 -501 0 feedthrough
rlabel pdiffusion 52 -501 52 -501 0 feedthrough
rlabel pdiffusion 59 -501 59 -501 0 cellNo=918
rlabel pdiffusion 66 -501 66 -501 0 cellNo=378
rlabel pdiffusion 73 -501 73 -501 0 feedthrough
rlabel pdiffusion 80 -501 80 -501 0 feedthrough
rlabel pdiffusion 87 -501 87 -501 0 feedthrough
rlabel pdiffusion 94 -501 94 -501 0 cellNo=15
rlabel pdiffusion 101 -501 101 -501 0 feedthrough
rlabel pdiffusion 108 -501 108 -501 0 cellNo=78
rlabel pdiffusion 115 -501 115 -501 0 cellNo=634
rlabel pdiffusion 122 -501 122 -501 0 feedthrough
rlabel pdiffusion 129 -501 129 -501 0 cellNo=225
rlabel pdiffusion 136 -501 136 -501 0 cellNo=920
rlabel pdiffusion 143 -501 143 -501 0 feedthrough
rlabel pdiffusion 150 -501 150 -501 0 cellNo=793
rlabel pdiffusion 157 -501 157 -501 0 cellNo=34
rlabel pdiffusion 164 -501 164 -501 0 cellNo=419
rlabel pdiffusion 171 -501 171 -501 0 feedthrough
rlabel pdiffusion 178 -501 178 -501 0 feedthrough
rlabel pdiffusion 185 -501 185 -501 0 feedthrough
rlabel pdiffusion 192 -501 192 -501 0 feedthrough
rlabel pdiffusion 199 -501 199 -501 0 cellNo=249
rlabel pdiffusion 206 -501 206 -501 0 cellNo=509
rlabel pdiffusion 213 -501 213 -501 0 cellNo=975
rlabel pdiffusion 220 -501 220 -501 0 feedthrough
rlabel pdiffusion 227 -501 227 -501 0 feedthrough
rlabel pdiffusion 234 -501 234 -501 0 feedthrough
rlabel pdiffusion 241 -501 241 -501 0 cellNo=986
rlabel pdiffusion 248 -501 248 -501 0 feedthrough
rlabel pdiffusion 255 -501 255 -501 0 feedthrough
rlabel pdiffusion 262 -501 262 -501 0 cellNo=586
rlabel pdiffusion 269 -501 269 -501 0 cellNo=865
rlabel pdiffusion 276 -501 276 -501 0 feedthrough
rlabel pdiffusion 283 -501 283 -501 0 feedthrough
rlabel pdiffusion 290 -501 290 -501 0 feedthrough
rlabel pdiffusion 297 -501 297 -501 0 feedthrough
rlabel pdiffusion 304 -501 304 -501 0 feedthrough
rlabel pdiffusion 311 -501 311 -501 0 feedthrough
rlabel pdiffusion 318 -501 318 -501 0 feedthrough
rlabel pdiffusion 325 -501 325 -501 0 feedthrough
rlabel pdiffusion 332 -501 332 -501 0 cellNo=372
rlabel pdiffusion 339 -501 339 -501 0 feedthrough
rlabel pdiffusion 346 -501 346 -501 0 feedthrough
rlabel pdiffusion 353 -501 353 -501 0 cellNo=766
rlabel pdiffusion 360 -501 360 -501 0 feedthrough
rlabel pdiffusion 367 -501 367 -501 0 cellNo=729
rlabel pdiffusion 374 -501 374 -501 0 feedthrough
rlabel pdiffusion 381 -501 381 -501 0 cellNo=459
rlabel pdiffusion 388 -501 388 -501 0 cellNo=143
rlabel pdiffusion 395 -501 395 -501 0 cellNo=257
rlabel pdiffusion 402 -501 402 -501 0 feedthrough
rlabel pdiffusion 409 -501 409 -501 0 feedthrough
rlabel pdiffusion 416 -501 416 -501 0 cellNo=138
rlabel pdiffusion 423 -501 423 -501 0 feedthrough
rlabel pdiffusion 430 -501 430 -501 0 feedthrough
rlabel pdiffusion 437 -501 437 -501 0 cellNo=260
rlabel pdiffusion 444 -501 444 -501 0 feedthrough
rlabel pdiffusion 451 -501 451 -501 0 feedthrough
rlabel pdiffusion 458 -501 458 -501 0 feedthrough
rlabel pdiffusion 465 -501 465 -501 0 feedthrough
rlabel pdiffusion 472 -501 472 -501 0 feedthrough
rlabel pdiffusion 479 -501 479 -501 0 cellNo=131
rlabel pdiffusion 486 -501 486 -501 0 feedthrough
rlabel pdiffusion 493 -501 493 -501 0 feedthrough
rlabel pdiffusion 500 -501 500 -501 0 feedthrough
rlabel pdiffusion 507 -501 507 -501 0 cellNo=274
rlabel pdiffusion 514 -501 514 -501 0 feedthrough
rlabel pdiffusion 521 -501 521 -501 0 feedthrough
rlabel pdiffusion 528 -501 528 -501 0 feedthrough
rlabel pdiffusion 535 -501 535 -501 0 feedthrough
rlabel pdiffusion 542 -501 542 -501 0 feedthrough
rlabel pdiffusion 549 -501 549 -501 0 feedthrough
rlabel pdiffusion 556 -501 556 -501 0 feedthrough
rlabel pdiffusion 563 -501 563 -501 0 feedthrough
rlabel pdiffusion 570 -501 570 -501 0 feedthrough
rlabel pdiffusion 577 -501 577 -501 0 feedthrough
rlabel pdiffusion 584 -501 584 -501 0 feedthrough
rlabel pdiffusion 591 -501 591 -501 0 cellNo=487
rlabel pdiffusion 598 -501 598 -501 0 feedthrough
rlabel pdiffusion 605 -501 605 -501 0 cellNo=797
rlabel pdiffusion 612 -501 612 -501 0 cellNo=711
rlabel pdiffusion 619 -501 619 -501 0 feedthrough
rlabel pdiffusion 626 -501 626 -501 0 cellNo=993
rlabel pdiffusion 633 -501 633 -501 0 feedthrough
rlabel pdiffusion 640 -501 640 -501 0 feedthrough
rlabel pdiffusion 647 -501 647 -501 0 feedthrough
rlabel pdiffusion 654 -501 654 -501 0 feedthrough
rlabel pdiffusion 661 -501 661 -501 0 feedthrough
rlabel pdiffusion 668 -501 668 -501 0 cellNo=352
rlabel pdiffusion 3 -558 3 -558 0 cellNo=60
rlabel pdiffusion 10 -558 10 -558 0 feedthrough
rlabel pdiffusion 17 -558 17 -558 0 feedthrough
rlabel pdiffusion 24 -558 24 -558 0 feedthrough
rlabel pdiffusion 31 -558 31 -558 0 feedthrough
rlabel pdiffusion 38 -558 38 -558 0 feedthrough
rlabel pdiffusion 45 -558 45 -558 0 feedthrough
rlabel pdiffusion 52 -558 52 -558 0 feedthrough
rlabel pdiffusion 59 -558 59 -558 0 cellNo=397
rlabel pdiffusion 66 -558 66 -558 0 feedthrough
rlabel pdiffusion 73 -558 73 -558 0 cellNo=782
rlabel pdiffusion 80 -558 80 -558 0 cellNo=9
rlabel pdiffusion 87 -558 87 -558 0 feedthrough
rlabel pdiffusion 94 -558 94 -558 0 feedthrough
rlabel pdiffusion 101 -558 101 -558 0 cellNo=594
rlabel pdiffusion 108 -558 108 -558 0 feedthrough
rlabel pdiffusion 115 -558 115 -558 0 cellNo=977
rlabel pdiffusion 122 -558 122 -558 0 feedthrough
rlabel pdiffusion 129 -558 129 -558 0 cellNo=332
rlabel pdiffusion 136 -558 136 -558 0 feedthrough
rlabel pdiffusion 143 -558 143 -558 0 cellNo=723
rlabel pdiffusion 150 -558 150 -558 0 cellNo=380
rlabel pdiffusion 157 -558 157 -558 0 feedthrough
rlabel pdiffusion 164 -558 164 -558 0 feedthrough
rlabel pdiffusion 171 -558 171 -558 0 feedthrough
rlabel pdiffusion 178 -558 178 -558 0 cellNo=361
rlabel pdiffusion 185 -558 185 -558 0 feedthrough
rlabel pdiffusion 192 -558 192 -558 0 cellNo=486
rlabel pdiffusion 199 -558 199 -558 0 feedthrough
rlabel pdiffusion 206 -558 206 -558 0 cellNo=647
rlabel pdiffusion 213 -558 213 -558 0 feedthrough
rlabel pdiffusion 220 -558 220 -558 0 feedthrough
rlabel pdiffusion 227 -558 227 -558 0 feedthrough
rlabel pdiffusion 234 -558 234 -558 0 feedthrough
rlabel pdiffusion 241 -558 241 -558 0 cellNo=726
rlabel pdiffusion 248 -558 248 -558 0 feedthrough
rlabel pdiffusion 255 -558 255 -558 0 feedthrough
rlabel pdiffusion 262 -558 262 -558 0 feedthrough
rlabel pdiffusion 269 -558 269 -558 0 feedthrough
rlabel pdiffusion 276 -558 276 -558 0 cellNo=842
rlabel pdiffusion 283 -558 283 -558 0 cellNo=375
rlabel pdiffusion 290 -558 290 -558 0 cellNo=995
rlabel pdiffusion 297 -558 297 -558 0 feedthrough
rlabel pdiffusion 304 -558 304 -558 0 feedthrough
rlabel pdiffusion 311 -558 311 -558 0 cellNo=527
rlabel pdiffusion 318 -558 318 -558 0 cellNo=102
rlabel pdiffusion 325 -558 325 -558 0 feedthrough
rlabel pdiffusion 332 -558 332 -558 0 feedthrough
rlabel pdiffusion 339 -558 339 -558 0 cellNo=933
rlabel pdiffusion 346 -558 346 -558 0 cellNo=783
rlabel pdiffusion 353 -558 353 -558 0 cellNo=115
rlabel pdiffusion 360 -558 360 -558 0 cellNo=504
rlabel pdiffusion 367 -558 367 -558 0 feedthrough
rlabel pdiffusion 374 -558 374 -558 0 cellNo=481
rlabel pdiffusion 381 -558 381 -558 0 feedthrough
rlabel pdiffusion 388 -558 388 -558 0 feedthrough
rlabel pdiffusion 395 -558 395 -558 0 feedthrough
rlabel pdiffusion 402 -558 402 -558 0 cellNo=336
rlabel pdiffusion 409 -558 409 -558 0 feedthrough
rlabel pdiffusion 416 -558 416 -558 0 feedthrough
rlabel pdiffusion 423 -558 423 -558 0 cellNo=275
rlabel pdiffusion 430 -558 430 -558 0 feedthrough
rlabel pdiffusion 437 -558 437 -558 0 feedthrough
rlabel pdiffusion 444 -558 444 -558 0 feedthrough
rlabel pdiffusion 451 -558 451 -558 0 feedthrough
rlabel pdiffusion 458 -558 458 -558 0 cellNo=640
rlabel pdiffusion 465 -558 465 -558 0 feedthrough
rlabel pdiffusion 472 -558 472 -558 0 feedthrough
rlabel pdiffusion 479 -558 479 -558 0 cellNo=748
rlabel pdiffusion 486 -558 486 -558 0 feedthrough
rlabel pdiffusion 493 -558 493 -558 0 feedthrough
rlabel pdiffusion 500 -558 500 -558 0 cellNo=828
rlabel pdiffusion 507 -558 507 -558 0 feedthrough
rlabel pdiffusion 514 -558 514 -558 0 feedthrough
rlabel pdiffusion 521 -558 521 -558 0 feedthrough
rlabel pdiffusion 528 -558 528 -558 0 feedthrough
rlabel pdiffusion 535 -558 535 -558 0 feedthrough
rlabel pdiffusion 542 -558 542 -558 0 feedthrough
rlabel pdiffusion 549 -558 549 -558 0 feedthrough
rlabel pdiffusion 556 -558 556 -558 0 feedthrough
rlabel pdiffusion 563 -558 563 -558 0 feedthrough
rlabel pdiffusion 570 -558 570 -558 0 feedthrough
rlabel pdiffusion 577 -558 577 -558 0 feedthrough
rlabel pdiffusion 584 -558 584 -558 0 feedthrough
rlabel pdiffusion 591 -558 591 -558 0 feedthrough
rlabel pdiffusion 598 -558 598 -558 0 feedthrough
rlabel pdiffusion 605 -558 605 -558 0 feedthrough
rlabel pdiffusion 612 -558 612 -558 0 feedthrough
rlabel pdiffusion 619 -558 619 -558 0 cellNo=132
rlabel pdiffusion 626 -558 626 -558 0 cellNo=454
rlabel pdiffusion 633 -558 633 -558 0 feedthrough
rlabel pdiffusion 640 -558 640 -558 0 feedthrough
rlabel pdiffusion 647 -558 647 -558 0 feedthrough
rlabel pdiffusion 654 -558 654 -558 0 feedthrough
rlabel pdiffusion 661 -558 661 -558 0 feedthrough
rlabel pdiffusion 668 -558 668 -558 0 cellNo=212
rlabel pdiffusion 675 -558 675 -558 0 feedthrough
rlabel pdiffusion 682 -558 682 -558 0 cellNo=376
rlabel pdiffusion 689 -558 689 -558 0 feedthrough
rlabel pdiffusion 3 -615 3 -615 0 feedthrough
rlabel pdiffusion 10 -615 10 -615 0 feedthrough
rlabel pdiffusion 17 -615 17 -615 0 cellNo=500
rlabel pdiffusion 24 -615 24 -615 0 feedthrough
rlabel pdiffusion 31 -615 31 -615 0 feedthrough
rlabel pdiffusion 38 -615 38 -615 0 cellNo=702
rlabel pdiffusion 45 -615 45 -615 0 cellNo=605
rlabel pdiffusion 52 -615 52 -615 0 feedthrough
rlabel pdiffusion 59 -615 59 -615 0 feedthrough
rlabel pdiffusion 66 -615 66 -615 0 feedthrough
rlabel pdiffusion 73 -615 73 -615 0 cellNo=675
rlabel pdiffusion 80 -615 80 -615 0 feedthrough
rlabel pdiffusion 87 -615 87 -615 0 cellNo=263
rlabel pdiffusion 94 -615 94 -615 0 cellNo=847
rlabel pdiffusion 101 -615 101 -615 0 cellNo=632
rlabel pdiffusion 108 -615 108 -615 0 feedthrough
rlabel pdiffusion 115 -615 115 -615 0 cellNo=279
rlabel pdiffusion 122 -615 122 -615 0 feedthrough
rlabel pdiffusion 129 -615 129 -615 0 cellNo=126
rlabel pdiffusion 136 -615 136 -615 0 feedthrough
rlabel pdiffusion 143 -615 143 -615 0 feedthrough
rlabel pdiffusion 150 -615 150 -615 0 feedthrough
rlabel pdiffusion 157 -615 157 -615 0 cellNo=705
rlabel pdiffusion 164 -615 164 -615 0 cellNo=835
rlabel pdiffusion 171 -615 171 -615 0 cellNo=754
rlabel pdiffusion 178 -615 178 -615 0 cellNo=858
rlabel pdiffusion 185 -615 185 -615 0 cellNo=269
rlabel pdiffusion 192 -615 192 -615 0 feedthrough
rlabel pdiffusion 199 -615 199 -615 0 feedthrough
rlabel pdiffusion 206 -615 206 -615 0 feedthrough
rlabel pdiffusion 213 -615 213 -615 0 feedthrough
rlabel pdiffusion 220 -615 220 -615 0 feedthrough
rlabel pdiffusion 227 -615 227 -615 0 feedthrough
rlabel pdiffusion 234 -615 234 -615 0 cellNo=808
rlabel pdiffusion 241 -615 241 -615 0 cellNo=839
rlabel pdiffusion 248 -615 248 -615 0 feedthrough
rlabel pdiffusion 255 -615 255 -615 0 feedthrough
rlabel pdiffusion 262 -615 262 -615 0 cellNo=139
rlabel pdiffusion 269 -615 269 -615 0 feedthrough
rlabel pdiffusion 276 -615 276 -615 0 cellNo=96
rlabel pdiffusion 283 -615 283 -615 0 feedthrough
rlabel pdiffusion 290 -615 290 -615 0 feedthrough
rlabel pdiffusion 297 -615 297 -615 0 feedthrough
rlabel pdiffusion 304 -615 304 -615 0 cellNo=691
rlabel pdiffusion 311 -615 311 -615 0 feedthrough
rlabel pdiffusion 318 -615 318 -615 0 feedthrough
rlabel pdiffusion 325 -615 325 -615 0 feedthrough
rlabel pdiffusion 332 -615 332 -615 0 feedthrough
rlabel pdiffusion 339 -615 339 -615 0 feedthrough
rlabel pdiffusion 346 -615 346 -615 0 feedthrough
rlabel pdiffusion 353 -615 353 -615 0 cellNo=243
rlabel pdiffusion 360 -615 360 -615 0 feedthrough
rlabel pdiffusion 367 -615 367 -615 0 cellNo=309
rlabel pdiffusion 374 -615 374 -615 0 feedthrough
rlabel pdiffusion 381 -615 381 -615 0 cellNo=745
rlabel pdiffusion 388 -615 388 -615 0 cellNo=978
rlabel pdiffusion 395 -615 395 -615 0 cellNo=903
rlabel pdiffusion 402 -615 402 -615 0 feedthrough
rlabel pdiffusion 409 -615 409 -615 0 feedthrough
rlabel pdiffusion 416 -615 416 -615 0 feedthrough
rlabel pdiffusion 423 -615 423 -615 0 feedthrough
rlabel pdiffusion 430 -615 430 -615 0 feedthrough
rlabel pdiffusion 437 -615 437 -615 0 feedthrough
rlabel pdiffusion 444 -615 444 -615 0 feedthrough
rlabel pdiffusion 451 -615 451 -615 0 cellNo=22
rlabel pdiffusion 458 -615 458 -615 0 feedthrough
rlabel pdiffusion 465 -615 465 -615 0 cellNo=446
rlabel pdiffusion 472 -615 472 -615 0 cellNo=780
rlabel pdiffusion 479 -615 479 -615 0 feedthrough
rlabel pdiffusion 486 -615 486 -615 0 feedthrough
rlabel pdiffusion 493 -615 493 -615 0 cellNo=614
rlabel pdiffusion 500 -615 500 -615 0 feedthrough
rlabel pdiffusion 507 -615 507 -615 0 feedthrough
rlabel pdiffusion 514 -615 514 -615 0 feedthrough
rlabel pdiffusion 521 -615 521 -615 0 feedthrough
rlabel pdiffusion 528 -615 528 -615 0 feedthrough
rlabel pdiffusion 535 -615 535 -615 0 feedthrough
rlabel pdiffusion 542 -615 542 -615 0 feedthrough
rlabel pdiffusion 549 -615 549 -615 0 feedthrough
rlabel pdiffusion 556 -615 556 -615 0 feedthrough
rlabel pdiffusion 563 -615 563 -615 0 feedthrough
rlabel pdiffusion 570 -615 570 -615 0 feedthrough
rlabel pdiffusion 577 -615 577 -615 0 feedthrough
rlabel pdiffusion 584 -615 584 -615 0 feedthrough
rlabel pdiffusion 591 -615 591 -615 0 feedthrough
rlabel pdiffusion 598 -615 598 -615 0 feedthrough
rlabel pdiffusion 605 -615 605 -615 0 cellNo=216
rlabel pdiffusion 612 -615 612 -615 0 feedthrough
rlabel pdiffusion 619 -615 619 -615 0 feedthrough
rlabel pdiffusion 626 -615 626 -615 0 feedthrough
rlabel pdiffusion 633 -615 633 -615 0 feedthrough
rlabel pdiffusion 640 -615 640 -615 0 feedthrough
rlabel pdiffusion 647 -615 647 -615 0 feedthrough
rlabel pdiffusion 654 -615 654 -615 0 cellNo=304
rlabel pdiffusion 661 -615 661 -615 0 feedthrough
rlabel pdiffusion 675 -615 675 -615 0 cellNo=937
rlabel pdiffusion 689 -615 689 -615 0 cellNo=340
rlabel pdiffusion 3 -688 3 -688 0 feedthrough
rlabel pdiffusion 10 -688 10 -688 0 feedthrough
rlabel pdiffusion 17 -688 17 -688 0 cellNo=526
rlabel pdiffusion 24 -688 24 -688 0 feedthrough
rlabel pdiffusion 31 -688 31 -688 0 feedthrough
rlabel pdiffusion 38 -688 38 -688 0 feedthrough
rlabel pdiffusion 45 -688 45 -688 0 feedthrough
rlabel pdiffusion 52 -688 52 -688 0 cellNo=709
rlabel pdiffusion 59 -688 59 -688 0 cellNo=830
rlabel pdiffusion 66 -688 66 -688 0 feedthrough
rlabel pdiffusion 73 -688 73 -688 0 feedthrough
rlabel pdiffusion 80 -688 80 -688 0 cellNo=564
rlabel pdiffusion 87 -688 87 -688 0 cellNo=50
rlabel pdiffusion 94 -688 94 -688 0 cellNo=32
rlabel pdiffusion 101 -688 101 -688 0 cellNo=698
rlabel pdiffusion 108 -688 108 -688 0 feedthrough
rlabel pdiffusion 115 -688 115 -688 0 feedthrough
rlabel pdiffusion 122 -688 122 -688 0 feedthrough
rlabel pdiffusion 129 -688 129 -688 0 feedthrough
rlabel pdiffusion 136 -688 136 -688 0 cellNo=74
rlabel pdiffusion 143 -688 143 -688 0 cellNo=123
rlabel pdiffusion 150 -688 150 -688 0 feedthrough
rlabel pdiffusion 157 -688 157 -688 0 feedthrough
rlabel pdiffusion 164 -688 164 -688 0 cellNo=365
rlabel pdiffusion 171 -688 171 -688 0 feedthrough
rlabel pdiffusion 178 -688 178 -688 0 feedthrough
rlabel pdiffusion 185 -688 185 -688 0 cellNo=166
rlabel pdiffusion 192 -688 192 -688 0 cellNo=849
rlabel pdiffusion 199 -688 199 -688 0 feedthrough
rlabel pdiffusion 206 -688 206 -688 0 feedthrough
rlabel pdiffusion 213 -688 213 -688 0 cellNo=77
rlabel pdiffusion 220 -688 220 -688 0 feedthrough
rlabel pdiffusion 227 -688 227 -688 0 cellNo=823
rlabel pdiffusion 234 -688 234 -688 0 cellNo=767
rlabel pdiffusion 241 -688 241 -688 0 cellNo=297
rlabel pdiffusion 248 -688 248 -688 0 feedthrough
rlabel pdiffusion 255 -688 255 -688 0 feedthrough
rlabel pdiffusion 262 -688 262 -688 0 feedthrough
rlabel pdiffusion 269 -688 269 -688 0 feedthrough
rlabel pdiffusion 276 -688 276 -688 0 cellNo=358
rlabel pdiffusion 283 -688 283 -688 0 cellNo=802
rlabel pdiffusion 290 -688 290 -688 0 feedthrough
rlabel pdiffusion 297 -688 297 -688 0 cellNo=421
rlabel pdiffusion 304 -688 304 -688 0 feedthrough
rlabel pdiffusion 311 -688 311 -688 0 feedthrough
rlabel pdiffusion 318 -688 318 -688 0 feedthrough
rlabel pdiffusion 325 -688 325 -688 0 feedthrough
rlabel pdiffusion 332 -688 332 -688 0 feedthrough
rlabel pdiffusion 339 -688 339 -688 0 feedthrough
rlabel pdiffusion 346 -688 346 -688 0 cellNo=907
rlabel pdiffusion 353 -688 353 -688 0 feedthrough
rlabel pdiffusion 360 -688 360 -688 0 cellNo=461
rlabel pdiffusion 367 -688 367 -688 0 cellNo=307
rlabel pdiffusion 374 -688 374 -688 0 cellNo=240
rlabel pdiffusion 381 -688 381 -688 0 feedthrough
rlabel pdiffusion 388 -688 388 -688 0 feedthrough
rlabel pdiffusion 395 -688 395 -688 0 feedthrough
rlabel pdiffusion 402 -688 402 -688 0 feedthrough
rlabel pdiffusion 409 -688 409 -688 0 cellNo=341
rlabel pdiffusion 416 -688 416 -688 0 feedthrough
rlabel pdiffusion 423 -688 423 -688 0 cellNo=5
rlabel pdiffusion 430 -688 430 -688 0 feedthrough
rlabel pdiffusion 437 -688 437 -688 0 feedthrough
rlabel pdiffusion 444 -688 444 -688 0 feedthrough
rlabel pdiffusion 451 -688 451 -688 0 cellNo=542
rlabel pdiffusion 458 -688 458 -688 0 cellNo=67
rlabel pdiffusion 465 -688 465 -688 0 cellNo=228
rlabel pdiffusion 472 -688 472 -688 0 feedthrough
rlabel pdiffusion 479 -688 479 -688 0 feedthrough
rlabel pdiffusion 486 -688 486 -688 0 feedthrough
rlabel pdiffusion 493 -688 493 -688 0 feedthrough
rlabel pdiffusion 500 -688 500 -688 0 feedthrough
rlabel pdiffusion 507 -688 507 -688 0 feedthrough
rlabel pdiffusion 514 -688 514 -688 0 feedthrough
rlabel pdiffusion 521 -688 521 -688 0 feedthrough
rlabel pdiffusion 528 -688 528 -688 0 feedthrough
rlabel pdiffusion 535 -688 535 -688 0 feedthrough
rlabel pdiffusion 542 -688 542 -688 0 feedthrough
rlabel pdiffusion 549 -688 549 -688 0 feedthrough
rlabel pdiffusion 556 -688 556 -688 0 feedthrough
rlabel pdiffusion 563 -688 563 -688 0 feedthrough
rlabel pdiffusion 570 -688 570 -688 0 feedthrough
rlabel pdiffusion 577 -688 577 -688 0 feedthrough
rlabel pdiffusion 584 -688 584 -688 0 feedthrough
rlabel pdiffusion 591 -688 591 -688 0 feedthrough
rlabel pdiffusion 598 -688 598 -688 0 feedthrough
rlabel pdiffusion 605 -688 605 -688 0 feedthrough
rlabel pdiffusion 612 -688 612 -688 0 feedthrough
rlabel pdiffusion 619 -688 619 -688 0 feedthrough
rlabel pdiffusion 626 -688 626 -688 0 feedthrough
rlabel pdiffusion 633 -688 633 -688 0 feedthrough
rlabel pdiffusion 640 -688 640 -688 0 feedthrough
rlabel pdiffusion 647 -688 647 -688 0 feedthrough
rlabel pdiffusion 654 -688 654 -688 0 feedthrough
rlabel pdiffusion 661 -688 661 -688 0 feedthrough
rlabel pdiffusion 668 -688 668 -688 0 feedthrough
rlabel pdiffusion 675 -688 675 -688 0 cellNo=674
rlabel pdiffusion 682 -688 682 -688 0 cellNo=834
rlabel pdiffusion 689 -688 689 -688 0 feedthrough
rlabel pdiffusion 696 -688 696 -688 0 feedthrough
rlabel pdiffusion 703 -688 703 -688 0 feedthrough
rlabel pdiffusion 717 -688 717 -688 0 cellNo=791
rlabel pdiffusion 731 -688 731 -688 0 feedthrough
rlabel pdiffusion 3 -755 3 -755 0 feedthrough
rlabel pdiffusion 10 -755 10 -755 0 feedthrough
rlabel pdiffusion 17 -755 17 -755 0 feedthrough
rlabel pdiffusion 24 -755 24 -755 0 feedthrough
rlabel pdiffusion 31 -755 31 -755 0 feedthrough
rlabel pdiffusion 38 -755 38 -755 0 cellNo=289
rlabel pdiffusion 45 -755 45 -755 0 feedthrough
rlabel pdiffusion 52 -755 52 -755 0 feedthrough
rlabel pdiffusion 59 -755 59 -755 0 feedthrough
rlabel pdiffusion 66 -755 66 -755 0 feedthrough
rlabel pdiffusion 73 -755 73 -755 0 feedthrough
rlabel pdiffusion 80 -755 80 -755 0 cellNo=427
rlabel pdiffusion 87 -755 87 -755 0 cellNo=710
rlabel pdiffusion 94 -755 94 -755 0 feedthrough
rlabel pdiffusion 101 -755 101 -755 0 cellNo=863
rlabel pdiffusion 108 -755 108 -755 0 feedthrough
rlabel pdiffusion 115 -755 115 -755 0 feedthrough
rlabel pdiffusion 122 -755 122 -755 0 cellNo=795
rlabel pdiffusion 129 -755 129 -755 0 feedthrough
rlabel pdiffusion 136 -755 136 -755 0 feedthrough
rlabel pdiffusion 143 -755 143 -755 0 feedthrough
rlabel pdiffusion 150 -755 150 -755 0 feedthrough
rlabel pdiffusion 157 -755 157 -755 0 feedthrough
rlabel pdiffusion 164 -755 164 -755 0 feedthrough
rlabel pdiffusion 171 -755 171 -755 0 feedthrough
rlabel pdiffusion 178 -755 178 -755 0 feedthrough
rlabel pdiffusion 185 -755 185 -755 0 feedthrough
rlabel pdiffusion 192 -755 192 -755 0 feedthrough
rlabel pdiffusion 199 -755 199 -755 0 cellNo=606
rlabel pdiffusion 206 -755 206 -755 0 feedthrough
rlabel pdiffusion 213 -755 213 -755 0 feedthrough
rlabel pdiffusion 220 -755 220 -755 0 feedthrough
rlabel pdiffusion 227 -755 227 -755 0 cellNo=905
rlabel pdiffusion 234 -755 234 -755 0 cellNo=816
rlabel pdiffusion 241 -755 241 -755 0 feedthrough
rlabel pdiffusion 248 -755 248 -755 0 cellNo=588
rlabel pdiffusion 255 -755 255 -755 0 feedthrough
rlabel pdiffusion 262 -755 262 -755 0 feedthrough
rlabel pdiffusion 269 -755 269 -755 0 feedthrough
rlabel pdiffusion 276 -755 276 -755 0 cellNo=997
rlabel pdiffusion 283 -755 283 -755 0 cellNo=321
rlabel pdiffusion 290 -755 290 -755 0 cellNo=654
rlabel pdiffusion 297 -755 297 -755 0 feedthrough
rlabel pdiffusion 304 -755 304 -755 0 feedthrough
rlabel pdiffusion 311 -755 311 -755 0 feedthrough
rlabel pdiffusion 318 -755 318 -755 0 feedthrough
rlabel pdiffusion 325 -755 325 -755 0 cellNo=401
rlabel pdiffusion 332 -755 332 -755 0 feedthrough
rlabel pdiffusion 339 -755 339 -755 0 cellNo=549
rlabel pdiffusion 346 -755 346 -755 0 feedthrough
rlabel pdiffusion 353 -755 353 -755 0 feedthrough
rlabel pdiffusion 360 -755 360 -755 0 cellNo=815
rlabel pdiffusion 367 -755 367 -755 0 feedthrough
rlabel pdiffusion 374 -755 374 -755 0 feedthrough
rlabel pdiffusion 381 -755 381 -755 0 cellNo=475
rlabel pdiffusion 388 -755 388 -755 0 cellNo=553
rlabel pdiffusion 395 -755 395 -755 0 cellNo=451
rlabel pdiffusion 402 -755 402 -755 0 feedthrough
rlabel pdiffusion 409 -755 409 -755 0 cellNo=64
rlabel pdiffusion 416 -755 416 -755 0 feedthrough
rlabel pdiffusion 423 -755 423 -755 0 feedthrough
rlabel pdiffusion 430 -755 430 -755 0 cellNo=217
rlabel pdiffusion 437 -755 437 -755 0 feedthrough
rlabel pdiffusion 444 -755 444 -755 0 feedthrough
rlabel pdiffusion 451 -755 451 -755 0 cellNo=744
rlabel pdiffusion 458 -755 458 -755 0 feedthrough
rlabel pdiffusion 465 -755 465 -755 0 feedthrough
rlabel pdiffusion 472 -755 472 -755 0 feedthrough
rlabel pdiffusion 479 -755 479 -755 0 feedthrough
rlabel pdiffusion 486 -755 486 -755 0 cellNo=469
rlabel pdiffusion 493 -755 493 -755 0 cellNo=638
rlabel pdiffusion 500 -755 500 -755 0 feedthrough
rlabel pdiffusion 507 -755 507 -755 0 feedthrough
rlabel pdiffusion 514 -755 514 -755 0 feedthrough
rlabel pdiffusion 521 -755 521 -755 0 feedthrough
rlabel pdiffusion 528 -755 528 -755 0 cellNo=609
rlabel pdiffusion 535 -755 535 -755 0 feedthrough
rlabel pdiffusion 542 -755 542 -755 0 cellNo=757
rlabel pdiffusion 549 -755 549 -755 0 feedthrough
rlabel pdiffusion 556 -755 556 -755 0 feedthrough
rlabel pdiffusion 563 -755 563 -755 0 cellNo=876
rlabel pdiffusion 570 -755 570 -755 0 feedthrough
rlabel pdiffusion 577 -755 577 -755 0 feedthrough
rlabel pdiffusion 584 -755 584 -755 0 cellNo=611
rlabel pdiffusion 591 -755 591 -755 0 feedthrough
rlabel pdiffusion 598 -755 598 -755 0 feedthrough
rlabel pdiffusion 605 -755 605 -755 0 feedthrough
rlabel pdiffusion 612 -755 612 -755 0 feedthrough
rlabel pdiffusion 619 -755 619 -755 0 feedthrough
rlabel pdiffusion 626 -755 626 -755 0 feedthrough
rlabel pdiffusion 633 -755 633 -755 0 feedthrough
rlabel pdiffusion 640 -755 640 -755 0 feedthrough
rlabel pdiffusion 647 -755 647 -755 0 feedthrough
rlabel pdiffusion 654 -755 654 -755 0 feedthrough
rlabel pdiffusion 661 -755 661 -755 0 feedthrough
rlabel pdiffusion 668 -755 668 -755 0 feedthrough
rlabel pdiffusion 675 -755 675 -755 0 feedthrough
rlabel pdiffusion 682 -755 682 -755 0 feedthrough
rlabel pdiffusion 689 -755 689 -755 0 feedthrough
rlabel pdiffusion 696 -755 696 -755 0 feedthrough
rlabel pdiffusion 703 -755 703 -755 0 feedthrough
rlabel pdiffusion 710 -755 710 -755 0 cellNo=973
rlabel pdiffusion 717 -755 717 -755 0 feedthrough
rlabel pdiffusion 724 -755 724 -755 0 feedthrough
rlabel pdiffusion 731 -755 731 -755 0 cellNo=81
rlabel pdiffusion 738 -755 738 -755 0 cellNo=208
rlabel pdiffusion 745 -755 745 -755 0 feedthrough
rlabel pdiffusion 752 -755 752 -755 0 cellNo=624
rlabel pdiffusion 801 -755 801 -755 0 cellNo=256
rlabel pdiffusion 808 -755 808 -755 0 feedthrough
rlabel pdiffusion 3 -832 3 -832 0 feedthrough
rlabel pdiffusion 10 -832 10 -832 0 feedthrough
rlabel pdiffusion 17 -832 17 -832 0 feedthrough
rlabel pdiffusion 24 -832 24 -832 0 cellNo=415
rlabel pdiffusion 31 -832 31 -832 0 cellNo=90
rlabel pdiffusion 38 -832 38 -832 0 feedthrough
rlabel pdiffusion 45 -832 45 -832 0 feedthrough
rlabel pdiffusion 52 -832 52 -832 0 cellNo=121
rlabel pdiffusion 59 -832 59 -832 0 feedthrough
rlabel pdiffusion 66 -832 66 -832 0 feedthrough
rlabel pdiffusion 73 -832 73 -832 0 feedthrough
rlabel pdiffusion 80 -832 80 -832 0 cellNo=593
rlabel pdiffusion 87 -832 87 -832 0 cellNo=942
rlabel pdiffusion 94 -832 94 -832 0 feedthrough
rlabel pdiffusion 101 -832 101 -832 0 feedthrough
rlabel pdiffusion 108 -832 108 -832 0 cellNo=503
rlabel pdiffusion 115 -832 115 -832 0 feedthrough
rlabel pdiffusion 122 -832 122 -832 0 cellNo=752
rlabel pdiffusion 129 -832 129 -832 0 feedthrough
rlabel pdiffusion 136 -832 136 -832 0 cellNo=645
rlabel pdiffusion 143 -832 143 -832 0 cellNo=38
rlabel pdiffusion 150 -832 150 -832 0 feedthrough
rlabel pdiffusion 157 -832 157 -832 0 feedthrough
rlabel pdiffusion 164 -832 164 -832 0 cellNo=885
rlabel pdiffusion 171 -832 171 -832 0 feedthrough
rlabel pdiffusion 178 -832 178 -832 0 feedthrough
rlabel pdiffusion 185 -832 185 -832 0 feedthrough
rlabel pdiffusion 192 -832 192 -832 0 cellNo=788
rlabel pdiffusion 199 -832 199 -832 0 cellNo=173
rlabel pdiffusion 206 -832 206 -832 0 feedthrough
rlabel pdiffusion 213 -832 213 -832 0 cellNo=669
rlabel pdiffusion 220 -832 220 -832 0 cellNo=915
rlabel pdiffusion 227 -832 227 -832 0 feedthrough
rlabel pdiffusion 234 -832 234 -832 0 feedthrough
rlabel pdiffusion 241 -832 241 -832 0 cellNo=278
rlabel pdiffusion 248 -832 248 -832 0 feedthrough
rlabel pdiffusion 255 -832 255 -832 0 feedthrough
rlabel pdiffusion 262 -832 262 -832 0 cellNo=550
rlabel pdiffusion 269 -832 269 -832 0 feedthrough
rlabel pdiffusion 276 -832 276 -832 0 feedthrough
rlabel pdiffusion 283 -832 283 -832 0 cellNo=499
rlabel pdiffusion 290 -832 290 -832 0 cellNo=408
rlabel pdiffusion 297 -832 297 -832 0 cellNo=205
rlabel pdiffusion 304 -832 304 -832 0 feedthrough
rlabel pdiffusion 311 -832 311 -832 0 feedthrough
rlabel pdiffusion 318 -832 318 -832 0 feedthrough
rlabel pdiffusion 325 -832 325 -832 0 feedthrough
rlabel pdiffusion 332 -832 332 -832 0 cellNo=31
rlabel pdiffusion 339 -832 339 -832 0 feedthrough
rlabel pdiffusion 346 -832 346 -832 0 feedthrough
rlabel pdiffusion 353 -832 353 -832 0 feedthrough
rlabel pdiffusion 360 -832 360 -832 0 feedthrough
rlabel pdiffusion 367 -832 367 -832 0 feedthrough
rlabel pdiffusion 374 -832 374 -832 0 feedthrough
rlabel pdiffusion 381 -832 381 -832 0 cellNo=312
rlabel pdiffusion 388 -832 388 -832 0 cellNo=666
rlabel pdiffusion 395 -832 395 -832 0 feedthrough
rlabel pdiffusion 402 -832 402 -832 0 cellNo=135
rlabel pdiffusion 409 -832 409 -832 0 feedthrough
rlabel pdiffusion 416 -832 416 -832 0 cellNo=837
rlabel pdiffusion 423 -832 423 -832 0 feedthrough
rlabel pdiffusion 430 -832 430 -832 0 cellNo=349
rlabel pdiffusion 437 -832 437 -832 0 cellNo=246
rlabel pdiffusion 444 -832 444 -832 0 feedthrough
rlabel pdiffusion 451 -832 451 -832 0 feedthrough
rlabel pdiffusion 458 -832 458 -832 0 cellNo=169
rlabel pdiffusion 465 -832 465 -832 0 feedthrough
rlabel pdiffusion 472 -832 472 -832 0 feedthrough
rlabel pdiffusion 479 -832 479 -832 0 feedthrough
rlabel pdiffusion 486 -832 486 -832 0 cellNo=628
rlabel pdiffusion 493 -832 493 -832 0 cellNo=99
rlabel pdiffusion 500 -832 500 -832 0 feedthrough
rlabel pdiffusion 507 -832 507 -832 0 feedthrough
rlabel pdiffusion 514 -832 514 -832 0 feedthrough
rlabel pdiffusion 521 -832 521 -832 0 cellNo=833
rlabel pdiffusion 528 -832 528 -832 0 cellNo=73
rlabel pdiffusion 535 -832 535 -832 0 feedthrough
rlabel pdiffusion 542 -832 542 -832 0 feedthrough
rlabel pdiffusion 549 -832 549 -832 0 feedthrough
rlabel pdiffusion 556 -832 556 -832 0 feedthrough
rlabel pdiffusion 563 -832 563 -832 0 feedthrough
rlabel pdiffusion 570 -832 570 -832 0 feedthrough
rlabel pdiffusion 577 -832 577 -832 0 feedthrough
rlabel pdiffusion 584 -832 584 -832 0 feedthrough
rlabel pdiffusion 591 -832 591 -832 0 feedthrough
rlabel pdiffusion 598 -832 598 -832 0 feedthrough
rlabel pdiffusion 605 -832 605 -832 0 feedthrough
rlabel pdiffusion 612 -832 612 -832 0 feedthrough
rlabel pdiffusion 619 -832 619 -832 0 feedthrough
rlabel pdiffusion 626 -832 626 -832 0 feedthrough
rlabel pdiffusion 633 -832 633 -832 0 feedthrough
rlabel pdiffusion 640 -832 640 -832 0 feedthrough
rlabel pdiffusion 647 -832 647 -832 0 feedthrough
rlabel pdiffusion 654 -832 654 -832 0 feedthrough
rlabel pdiffusion 661 -832 661 -832 0 feedthrough
rlabel pdiffusion 668 -832 668 -832 0 feedthrough
rlabel pdiffusion 675 -832 675 -832 0 feedthrough
rlabel pdiffusion 682 -832 682 -832 0 feedthrough
rlabel pdiffusion 689 -832 689 -832 0 feedthrough
rlabel pdiffusion 696 -832 696 -832 0 feedthrough
rlabel pdiffusion 703 -832 703 -832 0 feedthrough
rlabel pdiffusion 710 -832 710 -832 0 feedthrough
rlabel pdiffusion 717 -832 717 -832 0 feedthrough
rlabel pdiffusion 724 -832 724 -832 0 feedthrough
rlabel pdiffusion 731 -832 731 -832 0 feedthrough
rlabel pdiffusion 738 -832 738 -832 0 feedthrough
rlabel pdiffusion 745 -832 745 -832 0 feedthrough
rlabel pdiffusion 752 -832 752 -832 0 feedthrough
rlabel pdiffusion 759 -832 759 -832 0 feedthrough
rlabel pdiffusion 766 -832 766 -832 0 feedthrough
rlabel pdiffusion 773 -832 773 -832 0 feedthrough
rlabel pdiffusion 780 -832 780 -832 0 feedthrough
rlabel pdiffusion 787 -832 787 -832 0 feedthrough
rlabel pdiffusion 794 -832 794 -832 0 feedthrough
rlabel pdiffusion 801 -832 801 -832 0 cellNo=266
rlabel pdiffusion 808 -832 808 -832 0 feedthrough
rlabel pdiffusion 10 -919 10 -919 0 feedthrough
rlabel pdiffusion 17 -919 17 -919 0 feedthrough
rlabel pdiffusion 24 -919 24 -919 0 feedthrough
rlabel pdiffusion 31 -919 31 -919 0 feedthrough
rlabel pdiffusion 38 -919 38 -919 0 feedthrough
rlabel pdiffusion 45 -919 45 -919 0 feedthrough
rlabel pdiffusion 52 -919 52 -919 0 feedthrough
rlabel pdiffusion 59 -919 59 -919 0 feedthrough
rlabel pdiffusion 66 -919 66 -919 0 cellNo=557
rlabel pdiffusion 73 -919 73 -919 0 cellNo=7
rlabel pdiffusion 80 -919 80 -919 0 feedthrough
rlabel pdiffusion 87 -919 87 -919 0 cellNo=119
rlabel pdiffusion 94 -919 94 -919 0 feedthrough
rlabel pdiffusion 101 -919 101 -919 0 feedthrough
rlabel pdiffusion 108 -919 108 -919 0 feedthrough
rlabel pdiffusion 115 -919 115 -919 0 feedthrough
rlabel pdiffusion 122 -919 122 -919 0 feedthrough
rlabel pdiffusion 129 -919 129 -919 0 cellNo=693
rlabel pdiffusion 136 -919 136 -919 0 feedthrough
rlabel pdiffusion 143 -919 143 -919 0 feedthrough
rlabel pdiffusion 150 -919 150 -919 0 cellNo=194
rlabel pdiffusion 157 -919 157 -919 0 cellNo=536
rlabel pdiffusion 164 -919 164 -919 0 feedthrough
rlabel pdiffusion 171 -919 171 -919 0 cellNo=604
rlabel pdiffusion 178 -919 178 -919 0 cellNo=185
rlabel pdiffusion 185 -919 185 -919 0 feedthrough
rlabel pdiffusion 192 -919 192 -919 0 cellNo=442
rlabel pdiffusion 199 -919 199 -919 0 cellNo=333
rlabel pdiffusion 206 -919 206 -919 0 feedthrough
rlabel pdiffusion 213 -919 213 -919 0 feedthrough
rlabel pdiffusion 220 -919 220 -919 0 cellNo=113
rlabel pdiffusion 227 -919 227 -919 0 cellNo=46
rlabel pdiffusion 234 -919 234 -919 0 cellNo=428
rlabel pdiffusion 241 -919 241 -919 0 cellNo=813
rlabel pdiffusion 248 -919 248 -919 0 feedthrough
rlabel pdiffusion 255 -919 255 -919 0 feedthrough
rlabel pdiffusion 262 -919 262 -919 0 feedthrough
rlabel pdiffusion 269 -919 269 -919 0 feedthrough
rlabel pdiffusion 276 -919 276 -919 0 cellNo=337
rlabel pdiffusion 283 -919 283 -919 0 cellNo=391
rlabel pdiffusion 290 -919 290 -919 0 feedthrough
rlabel pdiffusion 297 -919 297 -919 0 feedthrough
rlabel pdiffusion 304 -919 304 -919 0 feedthrough
rlabel pdiffusion 311 -919 311 -919 0 feedthrough
rlabel pdiffusion 318 -919 318 -919 0 feedthrough
rlabel pdiffusion 325 -919 325 -919 0 feedthrough
rlabel pdiffusion 332 -919 332 -919 0 feedthrough
rlabel pdiffusion 339 -919 339 -919 0 feedthrough
rlabel pdiffusion 346 -919 346 -919 0 cellNo=411
rlabel pdiffusion 353 -919 353 -919 0 feedthrough
rlabel pdiffusion 360 -919 360 -919 0 feedthrough
rlabel pdiffusion 367 -919 367 -919 0 cellNo=369
rlabel pdiffusion 374 -919 374 -919 0 feedthrough
rlabel pdiffusion 381 -919 381 -919 0 cellNo=910
rlabel pdiffusion 388 -919 388 -919 0 feedthrough
rlabel pdiffusion 395 -919 395 -919 0 cellNo=494
rlabel pdiffusion 402 -919 402 -919 0 feedthrough
rlabel pdiffusion 409 -919 409 -919 0 cellNo=559
rlabel pdiffusion 416 -919 416 -919 0 cellNo=255
rlabel pdiffusion 423 -919 423 -919 0 feedthrough
rlabel pdiffusion 430 -919 430 -919 0 feedthrough
rlabel pdiffusion 437 -919 437 -919 0 feedthrough
rlabel pdiffusion 444 -919 444 -919 0 feedthrough
rlabel pdiffusion 451 -919 451 -919 0 cellNo=36
rlabel pdiffusion 458 -919 458 -919 0 cellNo=155
rlabel pdiffusion 465 -919 465 -919 0 cellNo=773
rlabel pdiffusion 472 -919 472 -919 0 feedthrough
rlabel pdiffusion 479 -919 479 -919 0 feedthrough
rlabel pdiffusion 486 -919 486 -919 0 cellNo=314
rlabel pdiffusion 493 -919 493 -919 0 feedthrough
rlabel pdiffusion 500 -919 500 -919 0 cellNo=108
rlabel pdiffusion 507 -919 507 -919 0 feedthrough
rlabel pdiffusion 514 -919 514 -919 0 feedthrough
rlabel pdiffusion 521 -919 521 -919 0 feedthrough
rlabel pdiffusion 528 -919 528 -919 0 feedthrough
rlabel pdiffusion 535 -919 535 -919 0 feedthrough
rlabel pdiffusion 542 -919 542 -919 0 feedthrough
rlabel pdiffusion 549 -919 549 -919 0 feedthrough
rlabel pdiffusion 556 -919 556 -919 0 feedthrough
rlabel pdiffusion 563 -919 563 -919 0 feedthrough
rlabel pdiffusion 570 -919 570 -919 0 feedthrough
rlabel pdiffusion 577 -919 577 -919 0 cellNo=636
rlabel pdiffusion 584 -919 584 -919 0 feedthrough
rlabel pdiffusion 591 -919 591 -919 0 feedthrough
rlabel pdiffusion 598 -919 598 -919 0 feedthrough
rlabel pdiffusion 605 -919 605 -919 0 feedthrough
rlabel pdiffusion 612 -919 612 -919 0 feedthrough
rlabel pdiffusion 619 -919 619 -919 0 feedthrough
rlabel pdiffusion 626 -919 626 -919 0 feedthrough
rlabel pdiffusion 633 -919 633 -919 0 feedthrough
rlabel pdiffusion 640 -919 640 -919 0 feedthrough
rlabel pdiffusion 647 -919 647 -919 0 feedthrough
rlabel pdiffusion 654 -919 654 -919 0 feedthrough
rlabel pdiffusion 661 -919 661 -919 0 feedthrough
rlabel pdiffusion 668 -919 668 -919 0 feedthrough
rlabel pdiffusion 675 -919 675 -919 0 feedthrough
rlabel pdiffusion 682 -919 682 -919 0 feedthrough
rlabel pdiffusion 689 -919 689 -919 0 feedthrough
rlabel pdiffusion 696 -919 696 -919 0 feedthrough
rlabel pdiffusion 703 -919 703 -919 0 feedthrough
rlabel pdiffusion 710 -919 710 -919 0 feedthrough
rlabel pdiffusion 717 -919 717 -919 0 feedthrough
rlabel pdiffusion 724 -919 724 -919 0 feedthrough
rlabel pdiffusion 731 -919 731 -919 0 feedthrough
rlabel pdiffusion 738 -919 738 -919 0 feedthrough
rlabel pdiffusion 745 -919 745 -919 0 feedthrough
rlabel pdiffusion 752 -919 752 -919 0 feedthrough
rlabel pdiffusion 759 -919 759 -919 0 feedthrough
rlabel pdiffusion 766 -919 766 -919 0 feedthrough
rlabel pdiffusion 773 -919 773 -919 0 cellNo=453
rlabel pdiffusion 780 -919 780 -919 0 cellNo=916
rlabel pdiffusion 787 -919 787 -919 0 feedthrough
rlabel pdiffusion 794 -919 794 -919 0 cellNo=976
rlabel pdiffusion 10 -996 10 -996 0 feedthrough
rlabel pdiffusion 17 -996 17 -996 0 feedthrough
rlabel pdiffusion 24 -996 24 -996 0 feedthrough
rlabel pdiffusion 31 -996 31 -996 0 feedthrough
rlabel pdiffusion 38 -996 38 -996 0 feedthrough
rlabel pdiffusion 45 -996 45 -996 0 feedthrough
rlabel pdiffusion 52 -996 52 -996 0 feedthrough
rlabel pdiffusion 59 -996 59 -996 0 feedthrough
rlabel pdiffusion 66 -996 66 -996 0 feedthrough
rlabel pdiffusion 73 -996 73 -996 0 cellNo=124
rlabel pdiffusion 80 -996 80 -996 0 cellNo=521
rlabel pdiffusion 87 -996 87 -996 0 feedthrough
rlabel pdiffusion 94 -996 94 -996 0 cellNo=881
rlabel pdiffusion 101 -996 101 -996 0 cellNo=422
rlabel pdiffusion 108 -996 108 -996 0 feedthrough
rlabel pdiffusion 115 -996 115 -996 0 cellNo=51
rlabel pdiffusion 122 -996 122 -996 0 feedthrough
rlabel pdiffusion 129 -996 129 -996 0 feedthrough
rlabel pdiffusion 136 -996 136 -996 0 feedthrough
rlabel pdiffusion 143 -996 143 -996 0 feedthrough
rlabel pdiffusion 150 -996 150 -996 0 feedthrough
rlabel pdiffusion 157 -996 157 -996 0 cellNo=480
rlabel pdiffusion 164 -996 164 -996 0 feedthrough
rlabel pdiffusion 171 -996 171 -996 0 feedthrough
rlabel pdiffusion 178 -996 178 -996 0 feedthrough
rlabel pdiffusion 185 -996 185 -996 0 feedthrough
rlabel pdiffusion 192 -996 192 -996 0 feedthrough
rlabel pdiffusion 199 -996 199 -996 0 cellNo=360
rlabel pdiffusion 206 -996 206 -996 0 feedthrough
rlabel pdiffusion 213 -996 213 -996 0 feedthrough
rlabel pdiffusion 220 -996 220 -996 0 cellNo=116
rlabel pdiffusion 227 -996 227 -996 0 feedthrough
rlabel pdiffusion 234 -996 234 -996 0 cellNo=209
rlabel pdiffusion 241 -996 241 -996 0 cellNo=502
rlabel pdiffusion 248 -996 248 -996 0 feedthrough
rlabel pdiffusion 255 -996 255 -996 0 cellNo=371
rlabel pdiffusion 262 -996 262 -996 0 feedthrough
rlabel pdiffusion 269 -996 269 -996 0 feedthrough
rlabel pdiffusion 276 -996 276 -996 0 feedthrough
rlabel pdiffusion 283 -996 283 -996 0 cellNo=383
rlabel pdiffusion 290 -996 290 -996 0 feedthrough
rlabel pdiffusion 297 -996 297 -996 0 feedthrough
rlabel pdiffusion 304 -996 304 -996 0 feedthrough
rlabel pdiffusion 311 -996 311 -996 0 cellNo=146
rlabel pdiffusion 318 -996 318 -996 0 cellNo=134
rlabel pdiffusion 325 -996 325 -996 0 feedthrough
rlabel pdiffusion 332 -996 332 -996 0 feedthrough
rlabel pdiffusion 339 -996 339 -996 0 feedthrough
rlabel pdiffusion 346 -996 346 -996 0 cellNo=196
rlabel pdiffusion 353 -996 353 -996 0 cellNo=133
rlabel pdiffusion 360 -996 360 -996 0 cellNo=516
rlabel pdiffusion 367 -996 367 -996 0 cellNo=890
rlabel pdiffusion 374 -996 374 -996 0 cellNo=58
rlabel pdiffusion 381 -996 381 -996 0 feedthrough
rlabel pdiffusion 388 -996 388 -996 0 cellNo=737
rlabel pdiffusion 395 -996 395 -996 0 cellNo=329
rlabel pdiffusion 402 -996 402 -996 0 feedthrough
rlabel pdiffusion 409 -996 409 -996 0 feedthrough
rlabel pdiffusion 416 -996 416 -996 0 cellNo=271
rlabel pdiffusion 423 -996 423 -996 0 cellNo=859
rlabel pdiffusion 430 -996 430 -996 0 cellNo=958
rlabel pdiffusion 437 -996 437 -996 0 feedthrough
rlabel pdiffusion 444 -996 444 -996 0 cellNo=680
rlabel pdiffusion 451 -996 451 -996 0 cellNo=753
rlabel pdiffusion 458 -996 458 -996 0 feedthrough
rlabel pdiffusion 465 -996 465 -996 0 cellNo=91
rlabel pdiffusion 472 -996 472 -996 0 cellNo=83
rlabel pdiffusion 479 -996 479 -996 0 feedthrough
rlabel pdiffusion 486 -996 486 -996 0 feedthrough
rlabel pdiffusion 493 -996 493 -996 0 feedthrough
rlabel pdiffusion 500 -996 500 -996 0 feedthrough
rlabel pdiffusion 507 -996 507 -996 0 feedthrough
rlabel pdiffusion 514 -996 514 -996 0 feedthrough
rlabel pdiffusion 521 -996 521 -996 0 feedthrough
rlabel pdiffusion 528 -996 528 -996 0 feedthrough
rlabel pdiffusion 535 -996 535 -996 0 cellNo=114
rlabel pdiffusion 542 -996 542 -996 0 feedthrough
rlabel pdiffusion 549 -996 549 -996 0 feedthrough
rlabel pdiffusion 556 -996 556 -996 0 feedthrough
rlabel pdiffusion 563 -996 563 -996 0 feedthrough
rlabel pdiffusion 570 -996 570 -996 0 feedthrough
rlabel pdiffusion 577 -996 577 -996 0 feedthrough
rlabel pdiffusion 584 -996 584 -996 0 feedthrough
rlabel pdiffusion 591 -996 591 -996 0 feedthrough
rlabel pdiffusion 598 -996 598 -996 0 feedthrough
rlabel pdiffusion 605 -996 605 -996 0 feedthrough
rlabel pdiffusion 612 -996 612 -996 0 feedthrough
rlabel pdiffusion 619 -996 619 -996 0 feedthrough
rlabel pdiffusion 626 -996 626 -996 0 feedthrough
rlabel pdiffusion 633 -996 633 -996 0 feedthrough
rlabel pdiffusion 640 -996 640 -996 0 feedthrough
rlabel pdiffusion 647 -996 647 -996 0 feedthrough
rlabel pdiffusion 654 -996 654 -996 0 feedthrough
rlabel pdiffusion 661 -996 661 -996 0 feedthrough
rlabel pdiffusion 668 -996 668 -996 0 feedthrough
rlabel pdiffusion 675 -996 675 -996 0 feedthrough
rlabel pdiffusion 682 -996 682 -996 0 feedthrough
rlabel pdiffusion 689 -996 689 -996 0 feedthrough
rlabel pdiffusion 696 -996 696 -996 0 feedthrough
rlabel pdiffusion 703 -996 703 -996 0 feedthrough
rlabel pdiffusion 710 -996 710 -996 0 feedthrough
rlabel pdiffusion 717 -996 717 -996 0 feedthrough
rlabel pdiffusion 724 -996 724 -996 0 feedthrough
rlabel pdiffusion 731 -996 731 -996 0 feedthrough
rlabel pdiffusion 738 -996 738 -996 0 cellNo=447
rlabel pdiffusion 745 -996 745 -996 0 cellNo=972
rlabel pdiffusion 752 -996 752 -996 0 cellNo=912
rlabel pdiffusion 759 -996 759 -996 0 feedthrough
rlabel pdiffusion 24 -1071 24 -1071 0 feedthrough
rlabel pdiffusion 31 -1071 31 -1071 0 cellNo=75
rlabel pdiffusion 38 -1071 38 -1071 0 feedthrough
rlabel pdiffusion 45 -1071 45 -1071 0 feedthrough
rlabel pdiffusion 52 -1071 52 -1071 0 feedthrough
rlabel pdiffusion 59 -1071 59 -1071 0 cellNo=189
rlabel pdiffusion 66 -1071 66 -1071 0 feedthrough
rlabel pdiffusion 73 -1071 73 -1071 0 cellNo=268
rlabel pdiffusion 80 -1071 80 -1071 0 feedthrough
rlabel pdiffusion 87 -1071 87 -1071 0 cellNo=273
rlabel pdiffusion 94 -1071 94 -1071 0 feedthrough
rlabel pdiffusion 101 -1071 101 -1071 0 cellNo=305
rlabel pdiffusion 108 -1071 108 -1071 0 cellNo=320
rlabel pdiffusion 115 -1071 115 -1071 0 feedthrough
rlabel pdiffusion 122 -1071 122 -1071 0 feedthrough
rlabel pdiffusion 129 -1071 129 -1071 0 feedthrough
rlabel pdiffusion 136 -1071 136 -1071 0 feedthrough
rlabel pdiffusion 143 -1071 143 -1071 0 feedthrough
rlabel pdiffusion 150 -1071 150 -1071 0 cellNo=105
rlabel pdiffusion 157 -1071 157 -1071 0 feedthrough
rlabel pdiffusion 164 -1071 164 -1071 0 cellNo=695
rlabel pdiffusion 171 -1071 171 -1071 0 feedthrough
rlabel pdiffusion 178 -1071 178 -1071 0 cellNo=334
rlabel pdiffusion 185 -1071 185 -1071 0 feedthrough
rlabel pdiffusion 192 -1071 192 -1071 0 cellNo=346
rlabel pdiffusion 199 -1071 199 -1071 0 cellNo=534
rlabel pdiffusion 206 -1071 206 -1071 0 feedthrough
rlabel pdiffusion 213 -1071 213 -1071 0 feedthrough
rlabel pdiffusion 220 -1071 220 -1071 0 feedthrough
rlabel pdiffusion 227 -1071 227 -1071 0 feedthrough
rlabel pdiffusion 234 -1071 234 -1071 0 feedthrough
rlabel pdiffusion 241 -1071 241 -1071 0 cellNo=811
rlabel pdiffusion 248 -1071 248 -1071 0 cellNo=891
rlabel pdiffusion 255 -1071 255 -1071 0 feedthrough
rlabel pdiffusion 262 -1071 262 -1071 0 feedthrough
rlabel pdiffusion 269 -1071 269 -1071 0 feedthrough
rlabel pdiffusion 276 -1071 276 -1071 0 cellNo=679
rlabel pdiffusion 283 -1071 283 -1071 0 feedthrough
rlabel pdiffusion 290 -1071 290 -1071 0 feedthrough
rlabel pdiffusion 297 -1071 297 -1071 0 feedthrough
rlabel pdiffusion 304 -1071 304 -1071 0 feedthrough
rlabel pdiffusion 311 -1071 311 -1071 0 cellNo=914
rlabel pdiffusion 318 -1071 318 -1071 0 feedthrough
rlabel pdiffusion 325 -1071 325 -1071 0 feedthrough
rlabel pdiffusion 332 -1071 332 -1071 0 cellNo=79
rlabel pdiffusion 339 -1071 339 -1071 0 feedthrough
rlabel pdiffusion 346 -1071 346 -1071 0 feedthrough
rlabel pdiffusion 353 -1071 353 -1071 0 feedthrough
rlabel pdiffusion 360 -1071 360 -1071 0 feedthrough
rlabel pdiffusion 367 -1071 367 -1071 0 feedthrough
rlabel pdiffusion 374 -1071 374 -1071 0 feedthrough
rlabel pdiffusion 381 -1071 381 -1071 0 feedthrough
rlabel pdiffusion 388 -1071 388 -1071 0 feedthrough
rlabel pdiffusion 395 -1071 395 -1071 0 feedthrough
rlabel pdiffusion 402 -1071 402 -1071 0 cellNo=17
rlabel pdiffusion 409 -1071 409 -1071 0 cellNo=519
rlabel pdiffusion 416 -1071 416 -1071 0 cellNo=80
rlabel pdiffusion 423 -1071 423 -1071 0 cellNo=462
rlabel pdiffusion 430 -1071 430 -1071 0 feedthrough
rlabel pdiffusion 437 -1071 437 -1071 0 cellNo=323
rlabel pdiffusion 444 -1071 444 -1071 0 feedthrough
rlabel pdiffusion 451 -1071 451 -1071 0 cellNo=253
rlabel pdiffusion 458 -1071 458 -1071 0 feedthrough
rlabel pdiffusion 465 -1071 465 -1071 0 feedthrough
rlabel pdiffusion 472 -1071 472 -1071 0 cellNo=381
rlabel pdiffusion 479 -1071 479 -1071 0 cellNo=590
rlabel pdiffusion 486 -1071 486 -1071 0 feedthrough
rlabel pdiffusion 493 -1071 493 -1071 0 cellNo=822
rlabel pdiffusion 500 -1071 500 -1071 0 feedthrough
rlabel pdiffusion 507 -1071 507 -1071 0 cellNo=708
rlabel pdiffusion 514 -1071 514 -1071 0 feedthrough
rlabel pdiffusion 521 -1071 521 -1071 0 cellNo=979
rlabel pdiffusion 528 -1071 528 -1071 0 feedthrough
rlabel pdiffusion 535 -1071 535 -1071 0 cellNo=468
rlabel pdiffusion 542 -1071 542 -1071 0 cellNo=853
rlabel pdiffusion 549 -1071 549 -1071 0 feedthrough
rlabel pdiffusion 556 -1071 556 -1071 0 feedthrough
rlabel pdiffusion 563 -1071 563 -1071 0 cellNo=284
rlabel pdiffusion 570 -1071 570 -1071 0 feedthrough
rlabel pdiffusion 577 -1071 577 -1071 0 feedthrough
rlabel pdiffusion 584 -1071 584 -1071 0 feedthrough
rlabel pdiffusion 591 -1071 591 -1071 0 feedthrough
rlabel pdiffusion 598 -1071 598 -1071 0 feedthrough
rlabel pdiffusion 605 -1071 605 -1071 0 feedthrough
rlabel pdiffusion 612 -1071 612 -1071 0 feedthrough
rlabel pdiffusion 619 -1071 619 -1071 0 feedthrough
rlabel pdiffusion 626 -1071 626 -1071 0 feedthrough
rlabel pdiffusion 633 -1071 633 -1071 0 feedthrough
rlabel pdiffusion 640 -1071 640 -1071 0 feedthrough
rlabel pdiffusion 647 -1071 647 -1071 0 feedthrough
rlabel pdiffusion 654 -1071 654 -1071 0 feedthrough
rlabel pdiffusion 661 -1071 661 -1071 0 feedthrough
rlabel pdiffusion 668 -1071 668 -1071 0 feedthrough
rlabel pdiffusion 675 -1071 675 -1071 0 feedthrough
rlabel pdiffusion 682 -1071 682 -1071 0 feedthrough
rlabel pdiffusion 689 -1071 689 -1071 0 cellNo=589
rlabel pdiffusion 696 -1071 696 -1071 0 feedthrough
rlabel pdiffusion 703 -1071 703 -1071 0 feedthrough
rlabel pdiffusion 710 -1071 710 -1071 0 feedthrough
rlabel pdiffusion 717 -1071 717 -1071 0 cellNo=676
rlabel pdiffusion 724 -1071 724 -1071 0 feedthrough
rlabel pdiffusion 731 -1071 731 -1071 0 feedthrough
rlabel pdiffusion 738 -1071 738 -1071 0 feedthrough
rlabel pdiffusion 10 -1132 10 -1132 0 feedthrough
rlabel pdiffusion 17 -1132 17 -1132 0 feedthrough
rlabel pdiffusion 24 -1132 24 -1132 0 feedthrough
rlabel pdiffusion 31 -1132 31 -1132 0 cellNo=684
rlabel pdiffusion 38 -1132 38 -1132 0 feedthrough
rlabel pdiffusion 45 -1132 45 -1132 0 cellNo=970
rlabel pdiffusion 52 -1132 52 -1132 0 feedthrough
rlabel pdiffusion 59 -1132 59 -1132 0 feedthrough
rlabel pdiffusion 66 -1132 66 -1132 0 cellNo=353
rlabel pdiffusion 73 -1132 73 -1132 0 feedthrough
rlabel pdiffusion 80 -1132 80 -1132 0 cellNo=136
rlabel pdiffusion 87 -1132 87 -1132 0 feedthrough
rlabel pdiffusion 94 -1132 94 -1132 0 cellNo=505
rlabel pdiffusion 101 -1132 101 -1132 0 feedthrough
rlabel pdiffusion 108 -1132 108 -1132 0 feedthrough
rlabel pdiffusion 115 -1132 115 -1132 0 feedthrough
rlabel pdiffusion 122 -1132 122 -1132 0 cellNo=554
rlabel pdiffusion 129 -1132 129 -1132 0 feedthrough
rlabel pdiffusion 136 -1132 136 -1132 0 feedthrough
rlabel pdiffusion 143 -1132 143 -1132 0 cellNo=363
rlabel pdiffusion 150 -1132 150 -1132 0 feedthrough
rlabel pdiffusion 157 -1132 157 -1132 0 cellNo=928
rlabel pdiffusion 164 -1132 164 -1132 0 cellNo=344
rlabel pdiffusion 171 -1132 171 -1132 0 cellNo=61
rlabel pdiffusion 178 -1132 178 -1132 0 cellNo=850
rlabel pdiffusion 185 -1132 185 -1132 0 cellNo=525
rlabel pdiffusion 192 -1132 192 -1132 0 cellNo=944
rlabel pdiffusion 199 -1132 199 -1132 0 cellNo=854
rlabel pdiffusion 206 -1132 206 -1132 0 feedthrough
rlabel pdiffusion 213 -1132 213 -1132 0 cellNo=122
rlabel pdiffusion 220 -1132 220 -1132 0 feedthrough
rlabel pdiffusion 227 -1132 227 -1132 0 feedthrough
rlabel pdiffusion 234 -1132 234 -1132 0 feedthrough
rlabel pdiffusion 241 -1132 241 -1132 0 cellNo=94
rlabel pdiffusion 248 -1132 248 -1132 0 cellNo=896
rlabel pdiffusion 255 -1132 255 -1132 0 feedthrough
rlabel pdiffusion 262 -1132 262 -1132 0 feedthrough
rlabel pdiffusion 269 -1132 269 -1132 0 feedthrough
rlabel pdiffusion 276 -1132 276 -1132 0 cellNo=556
rlabel pdiffusion 283 -1132 283 -1132 0 feedthrough
rlabel pdiffusion 290 -1132 290 -1132 0 feedthrough
rlabel pdiffusion 297 -1132 297 -1132 0 feedthrough
rlabel pdiffusion 304 -1132 304 -1132 0 feedthrough
rlabel pdiffusion 311 -1132 311 -1132 0 cellNo=290
rlabel pdiffusion 318 -1132 318 -1132 0 feedthrough
rlabel pdiffusion 325 -1132 325 -1132 0 feedthrough
rlabel pdiffusion 332 -1132 332 -1132 0 cellNo=392
rlabel pdiffusion 339 -1132 339 -1132 0 feedthrough
rlabel pdiffusion 346 -1132 346 -1132 0 cellNo=319
rlabel pdiffusion 353 -1132 353 -1132 0 feedthrough
rlabel pdiffusion 360 -1132 360 -1132 0 cellNo=338
rlabel pdiffusion 367 -1132 367 -1132 0 cellNo=683
rlabel pdiffusion 374 -1132 374 -1132 0 cellNo=311
rlabel pdiffusion 381 -1132 381 -1132 0 cellNo=756
rlabel pdiffusion 388 -1132 388 -1132 0 cellNo=840
rlabel pdiffusion 395 -1132 395 -1132 0 cellNo=935
rlabel pdiffusion 402 -1132 402 -1132 0 feedthrough
rlabel pdiffusion 409 -1132 409 -1132 0 feedthrough
rlabel pdiffusion 416 -1132 416 -1132 0 feedthrough
rlabel pdiffusion 423 -1132 423 -1132 0 cellNo=251
rlabel pdiffusion 430 -1132 430 -1132 0 cellNo=368
rlabel pdiffusion 437 -1132 437 -1132 0 feedthrough
rlabel pdiffusion 444 -1132 444 -1132 0 feedthrough
rlabel pdiffusion 451 -1132 451 -1132 0 feedthrough
rlabel pdiffusion 458 -1132 458 -1132 0 feedthrough
rlabel pdiffusion 465 -1132 465 -1132 0 feedthrough
rlabel pdiffusion 472 -1132 472 -1132 0 feedthrough
rlabel pdiffusion 479 -1132 479 -1132 0 feedthrough
rlabel pdiffusion 486 -1132 486 -1132 0 feedthrough
rlabel pdiffusion 493 -1132 493 -1132 0 feedthrough
rlabel pdiffusion 500 -1132 500 -1132 0 feedthrough
rlabel pdiffusion 507 -1132 507 -1132 0 cellNo=10
rlabel pdiffusion 514 -1132 514 -1132 0 feedthrough
rlabel pdiffusion 521 -1132 521 -1132 0 cellNo=282
rlabel pdiffusion 528 -1132 528 -1132 0 feedthrough
rlabel pdiffusion 535 -1132 535 -1132 0 feedthrough
rlabel pdiffusion 542 -1132 542 -1132 0 feedthrough
rlabel pdiffusion 549 -1132 549 -1132 0 feedthrough
rlabel pdiffusion 556 -1132 556 -1132 0 feedthrough
rlabel pdiffusion 563 -1132 563 -1132 0 feedthrough
rlabel pdiffusion 570 -1132 570 -1132 0 feedthrough
rlabel pdiffusion 577 -1132 577 -1132 0 feedthrough
rlabel pdiffusion 584 -1132 584 -1132 0 feedthrough
rlabel pdiffusion 591 -1132 591 -1132 0 feedthrough
rlabel pdiffusion 598 -1132 598 -1132 0 feedthrough
rlabel pdiffusion 605 -1132 605 -1132 0 feedthrough
rlabel pdiffusion 612 -1132 612 -1132 0 feedthrough
rlabel pdiffusion 619 -1132 619 -1132 0 feedthrough
rlabel pdiffusion 626 -1132 626 -1132 0 feedthrough
rlabel pdiffusion 633 -1132 633 -1132 0 feedthrough
rlabel pdiffusion 640 -1132 640 -1132 0 feedthrough
rlabel pdiffusion 647 -1132 647 -1132 0 feedthrough
rlabel pdiffusion 654 -1132 654 -1132 0 feedthrough
rlabel pdiffusion 661 -1132 661 -1132 0 feedthrough
rlabel pdiffusion 668 -1132 668 -1132 0 feedthrough
rlabel pdiffusion 675 -1132 675 -1132 0 cellNo=989
rlabel pdiffusion 682 -1132 682 -1132 0 cellNo=478
rlabel pdiffusion 689 -1132 689 -1132 0 feedthrough
rlabel pdiffusion 696 -1132 696 -1132 0 feedthrough
rlabel pdiffusion 703 -1132 703 -1132 0 feedthrough
rlabel pdiffusion 710 -1132 710 -1132 0 feedthrough
rlabel pdiffusion 3 -1189 3 -1189 0 feedthrough
rlabel pdiffusion 10 -1189 10 -1189 0 feedthrough
rlabel pdiffusion 17 -1189 17 -1189 0 cellNo=242
rlabel pdiffusion 24 -1189 24 -1189 0 cellNo=221
rlabel pdiffusion 31 -1189 31 -1189 0 feedthrough
rlabel pdiffusion 38 -1189 38 -1189 0 feedthrough
rlabel pdiffusion 45 -1189 45 -1189 0 feedthrough
rlabel pdiffusion 52 -1189 52 -1189 0 feedthrough
rlabel pdiffusion 59 -1189 59 -1189 0 feedthrough
rlabel pdiffusion 66 -1189 66 -1189 0 cellNo=730
rlabel pdiffusion 73 -1189 73 -1189 0 cellNo=616
rlabel pdiffusion 80 -1189 80 -1189 0 feedthrough
rlabel pdiffusion 87 -1189 87 -1189 0 cellNo=224
rlabel pdiffusion 94 -1189 94 -1189 0 feedthrough
rlabel pdiffusion 101 -1189 101 -1189 0 cellNo=733
rlabel pdiffusion 108 -1189 108 -1189 0 cellNo=948
rlabel pdiffusion 115 -1189 115 -1189 0 cellNo=85
rlabel pdiffusion 122 -1189 122 -1189 0 feedthrough
rlabel pdiffusion 129 -1189 129 -1189 0 feedthrough
rlabel pdiffusion 136 -1189 136 -1189 0 feedthrough
rlabel pdiffusion 143 -1189 143 -1189 0 cellNo=814
rlabel pdiffusion 150 -1189 150 -1189 0 cellNo=405
rlabel pdiffusion 157 -1189 157 -1189 0 cellNo=760
rlabel pdiffusion 164 -1189 164 -1189 0 feedthrough
rlabel pdiffusion 171 -1189 171 -1189 0 cellNo=867
rlabel pdiffusion 178 -1189 178 -1189 0 feedthrough
rlabel pdiffusion 185 -1189 185 -1189 0 feedthrough
rlabel pdiffusion 192 -1189 192 -1189 0 cellNo=662
rlabel pdiffusion 199 -1189 199 -1189 0 feedthrough
rlabel pdiffusion 206 -1189 206 -1189 0 cellNo=717
rlabel pdiffusion 213 -1189 213 -1189 0 cellNo=659
rlabel pdiffusion 220 -1189 220 -1189 0 feedthrough
rlabel pdiffusion 227 -1189 227 -1189 0 feedthrough
rlabel pdiffusion 234 -1189 234 -1189 0 cellNo=597
rlabel pdiffusion 241 -1189 241 -1189 0 feedthrough
rlabel pdiffusion 248 -1189 248 -1189 0 feedthrough
rlabel pdiffusion 255 -1189 255 -1189 0 feedthrough
rlabel pdiffusion 262 -1189 262 -1189 0 feedthrough
rlabel pdiffusion 269 -1189 269 -1189 0 feedthrough
rlabel pdiffusion 276 -1189 276 -1189 0 cellNo=980
rlabel pdiffusion 283 -1189 283 -1189 0 feedthrough
rlabel pdiffusion 290 -1189 290 -1189 0 feedthrough
rlabel pdiffusion 297 -1189 297 -1189 0 feedthrough
rlabel pdiffusion 304 -1189 304 -1189 0 cellNo=11
rlabel pdiffusion 311 -1189 311 -1189 0 feedthrough
rlabel pdiffusion 318 -1189 318 -1189 0 cellNo=231
rlabel pdiffusion 325 -1189 325 -1189 0 cellNo=763
rlabel pdiffusion 332 -1189 332 -1189 0 cellNo=448
rlabel pdiffusion 339 -1189 339 -1189 0 cellNo=630
rlabel pdiffusion 346 -1189 346 -1189 0 cellNo=913
rlabel pdiffusion 353 -1189 353 -1189 0 feedthrough
rlabel pdiffusion 360 -1189 360 -1189 0 feedthrough
rlabel pdiffusion 367 -1189 367 -1189 0 feedthrough
rlabel pdiffusion 374 -1189 374 -1189 0 feedthrough
rlabel pdiffusion 381 -1189 381 -1189 0 feedthrough
rlabel pdiffusion 388 -1189 388 -1189 0 cellNo=939
rlabel pdiffusion 395 -1189 395 -1189 0 feedthrough
rlabel pdiffusion 402 -1189 402 -1189 0 feedthrough
rlabel pdiffusion 409 -1189 409 -1189 0 feedthrough
rlabel pdiffusion 416 -1189 416 -1189 0 feedthrough
rlabel pdiffusion 423 -1189 423 -1189 0 feedthrough
rlabel pdiffusion 430 -1189 430 -1189 0 feedthrough
rlabel pdiffusion 437 -1189 437 -1189 0 cellNo=735
rlabel pdiffusion 444 -1189 444 -1189 0 cellNo=170
rlabel pdiffusion 451 -1189 451 -1189 0 cellNo=945
rlabel pdiffusion 458 -1189 458 -1189 0 feedthrough
rlabel pdiffusion 465 -1189 465 -1189 0 cellNo=667
rlabel pdiffusion 472 -1189 472 -1189 0 feedthrough
rlabel pdiffusion 479 -1189 479 -1189 0 feedthrough
rlabel pdiffusion 486 -1189 486 -1189 0 feedthrough
rlabel pdiffusion 493 -1189 493 -1189 0 feedthrough
rlabel pdiffusion 500 -1189 500 -1189 0 feedthrough
rlabel pdiffusion 507 -1189 507 -1189 0 feedthrough
rlabel pdiffusion 514 -1189 514 -1189 0 feedthrough
rlabel pdiffusion 521 -1189 521 -1189 0 feedthrough
rlabel pdiffusion 528 -1189 528 -1189 0 cellNo=749
rlabel pdiffusion 535 -1189 535 -1189 0 feedthrough
rlabel pdiffusion 542 -1189 542 -1189 0 cellNo=227
rlabel pdiffusion 549 -1189 549 -1189 0 feedthrough
rlabel pdiffusion 556 -1189 556 -1189 0 feedthrough
rlabel pdiffusion 563 -1189 563 -1189 0 feedthrough
rlabel pdiffusion 570 -1189 570 -1189 0 feedthrough
rlabel pdiffusion 577 -1189 577 -1189 0 feedthrough
rlabel pdiffusion 584 -1189 584 -1189 0 feedthrough
rlabel pdiffusion 591 -1189 591 -1189 0 feedthrough
rlabel pdiffusion 598 -1189 598 -1189 0 feedthrough
rlabel pdiffusion 605 -1189 605 -1189 0 feedthrough
rlabel pdiffusion 612 -1189 612 -1189 0 feedthrough
rlabel pdiffusion 619 -1189 619 -1189 0 feedthrough
rlabel pdiffusion 626 -1189 626 -1189 0 feedthrough
rlabel pdiffusion 633 -1189 633 -1189 0 feedthrough
rlabel pdiffusion 640 -1189 640 -1189 0 feedthrough
rlabel pdiffusion 647 -1189 647 -1189 0 feedthrough
rlabel pdiffusion 654 -1189 654 -1189 0 cellNo=293
rlabel pdiffusion 661 -1189 661 -1189 0 feedthrough
rlabel pdiffusion 668 -1189 668 -1189 0 cellNo=724
rlabel pdiffusion 675 -1189 675 -1189 0 cellNo=501
rlabel pdiffusion 682 -1189 682 -1189 0 feedthrough
rlabel pdiffusion 689 -1189 689 -1189 0 feedthrough
rlabel pdiffusion 703 -1189 703 -1189 0 feedthrough
rlabel pdiffusion 710 -1189 710 -1189 0 feedthrough
rlabel pdiffusion 3 -1260 3 -1260 0 feedthrough
rlabel pdiffusion 10 -1260 10 -1260 0 feedthrough
rlabel pdiffusion 17 -1260 17 -1260 0 feedthrough
rlabel pdiffusion 24 -1260 24 -1260 0 feedthrough
rlabel pdiffusion 31 -1260 31 -1260 0 feedthrough
rlabel pdiffusion 38 -1260 38 -1260 0 feedthrough
rlabel pdiffusion 45 -1260 45 -1260 0 cellNo=356
rlabel pdiffusion 52 -1260 52 -1260 0 cellNo=817
rlabel pdiffusion 59 -1260 59 -1260 0 cellNo=248
rlabel pdiffusion 66 -1260 66 -1260 0 feedthrough
rlabel pdiffusion 73 -1260 73 -1260 0 cellNo=435
rlabel pdiffusion 80 -1260 80 -1260 0 feedthrough
rlabel pdiffusion 87 -1260 87 -1260 0 feedthrough
rlabel pdiffusion 94 -1260 94 -1260 0 feedthrough
rlabel pdiffusion 101 -1260 101 -1260 0 cellNo=6
rlabel pdiffusion 108 -1260 108 -1260 0 cellNo=571
rlabel pdiffusion 115 -1260 115 -1260 0 feedthrough
rlabel pdiffusion 122 -1260 122 -1260 0 cellNo=848
rlabel pdiffusion 129 -1260 129 -1260 0 feedthrough
rlabel pdiffusion 136 -1260 136 -1260 0 feedthrough
rlabel pdiffusion 143 -1260 143 -1260 0 cellNo=678
rlabel pdiffusion 150 -1260 150 -1260 0 feedthrough
rlabel pdiffusion 157 -1260 157 -1260 0 feedthrough
rlabel pdiffusion 164 -1260 164 -1260 0 cellNo=495
rlabel pdiffusion 171 -1260 171 -1260 0 feedthrough
rlabel pdiffusion 178 -1260 178 -1260 0 cellNo=272
rlabel pdiffusion 185 -1260 185 -1260 0 cellNo=764
rlabel pdiffusion 192 -1260 192 -1260 0 cellNo=908
rlabel pdiffusion 199 -1260 199 -1260 0 cellNo=869
rlabel pdiffusion 206 -1260 206 -1260 0 feedthrough
rlabel pdiffusion 213 -1260 213 -1260 0 cellNo=663
rlabel pdiffusion 220 -1260 220 -1260 0 cellNo=318
rlabel pdiffusion 227 -1260 227 -1260 0 cellNo=796
rlabel pdiffusion 234 -1260 234 -1260 0 cellNo=127
rlabel pdiffusion 241 -1260 241 -1260 0 feedthrough
rlabel pdiffusion 248 -1260 248 -1260 0 cellNo=162
rlabel pdiffusion 255 -1260 255 -1260 0 cellNo=578
rlabel pdiffusion 262 -1260 262 -1260 0 feedthrough
rlabel pdiffusion 269 -1260 269 -1260 0 cellNo=546
rlabel pdiffusion 276 -1260 276 -1260 0 feedthrough
rlabel pdiffusion 283 -1260 283 -1260 0 feedthrough
rlabel pdiffusion 290 -1260 290 -1260 0 feedthrough
rlabel pdiffusion 297 -1260 297 -1260 0 feedthrough
rlabel pdiffusion 304 -1260 304 -1260 0 cellNo=568
rlabel pdiffusion 311 -1260 311 -1260 0 cellNo=615
rlabel pdiffusion 318 -1260 318 -1260 0 feedthrough
rlabel pdiffusion 325 -1260 325 -1260 0 cellNo=779
rlabel pdiffusion 332 -1260 332 -1260 0 cellNo=671
rlabel pdiffusion 339 -1260 339 -1260 0 feedthrough
rlabel pdiffusion 346 -1260 346 -1260 0 feedthrough
rlabel pdiffusion 353 -1260 353 -1260 0 cellNo=182
rlabel pdiffusion 360 -1260 360 -1260 0 feedthrough
rlabel pdiffusion 367 -1260 367 -1260 0 feedthrough
rlabel pdiffusion 374 -1260 374 -1260 0 feedthrough
rlabel pdiffusion 381 -1260 381 -1260 0 cellNo=715
rlabel pdiffusion 388 -1260 388 -1260 0 feedthrough
rlabel pdiffusion 395 -1260 395 -1260 0 cellNo=47
rlabel pdiffusion 402 -1260 402 -1260 0 feedthrough
rlabel pdiffusion 409 -1260 409 -1260 0 feedthrough
rlabel pdiffusion 416 -1260 416 -1260 0 feedthrough
rlabel pdiffusion 423 -1260 423 -1260 0 feedthrough
rlabel pdiffusion 430 -1260 430 -1260 0 cellNo=197
rlabel pdiffusion 437 -1260 437 -1260 0 feedthrough
rlabel pdiffusion 444 -1260 444 -1260 0 feedthrough
rlabel pdiffusion 451 -1260 451 -1260 0 cellNo=103
rlabel pdiffusion 458 -1260 458 -1260 0 cellNo=960
rlabel pdiffusion 465 -1260 465 -1260 0 feedthrough
rlabel pdiffusion 472 -1260 472 -1260 0 feedthrough
rlabel pdiffusion 479 -1260 479 -1260 0 feedthrough
rlabel pdiffusion 486 -1260 486 -1260 0 feedthrough
rlabel pdiffusion 493 -1260 493 -1260 0 cellNo=718
rlabel pdiffusion 500 -1260 500 -1260 0 feedthrough
rlabel pdiffusion 507 -1260 507 -1260 0 feedthrough
rlabel pdiffusion 514 -1260 514 -1260 0 cellNo=463
rlabel pdiffusion 521 -1260 521 -1260 0 feedthrough
rlabel pdiffusion 528 -1260 528 -1260 0 feedthrough
rlabel pdiffusion 535 -1260 535 -1260 0 feedthrough
rlabel pdiffusion 542 -1260 542 -1260 0 feedthrough
rlabel pdiffusion 549 -1260 549 -1260 0 feedthrough
rlabel pdiffusion 556 -1260 556 -1260 0 feedthrough
rlabel pdiffusion 563 -1260 563 -1260 0 feedthrough
rlabel pdiffusion 570 -1260 570 -1260 0 feedthrough
rlabel pdiffusion 577 -1260 577 -1260 0 feedthrough
rlabel pdiffusion 584 -1260 584 -1260 0 feedthrough
rlabel pdiffusion 591 -1260 591 -1260 0 feedthrough
rlabel pdiffusion 598 -1260 598 -1260 0 feedthrough
rlabel pdiffusion 605 -1260 605 -1260 0 feedthrough
rlabel pdiffusion 612 -1260 612 -1260 0 feedthrough
rlabel pdiffusion 619 -1260 619 -1260 0 feedthrough
rlabel pdiffusion 626 -1260 626 -1260 0 feedthrough
rlabel pdiffusion 633 -1260 633 -1260 0 feedthrough
rlabel pdiffusion 640 -1260 640 -1260 0 feedthrough
rlabel pdiffusion 647 -1260 647 -1260 0 feedthrough
rlabel pdiffusion 654 -1260 654 -1260 0 feedthrough
rlabel pdiffusion 661 -1260 661 -1260 0 feedthrough
rlabel pdiffusion 668 -1260 668 -1260 0 feedthrough
rlabel pdiffusion 675 -1260 675 -1260 0 feedthrough
rlabel pdiffusion 682 -1260 682 -1260 0 feedthrough
rlabel pdiffusion 689 -1260 689 -1260 0 feedthrough
rlabel pdiffusion 696 -1260 696 -1260 0 feedthrough
rlabel pdiffusion 703 -1260 703 -1260 0 cellNo=819
rlabel pdiffusion 710 -1260 710 -1260 0 cellNo=579
rlabel pdiffusion 717 -1260 717 -1260 0 feedthrough
rlabel pdiffusion 3 -1331 3 -1331 0 feedthrough
rlabel pdiffusion 10 -1331 10 -1331 0 feedthrough
rlabel pdiffusion 17 -1331 17 -1331 0 cellNo=873
rlabel pdiffusion 24 -1331 24 -1331 0 feedthrough
rlabel pdiffusion 31 -1331 31 -1331 0 cellNo=445
rlabel pdiffusion 38 -1331 38 -1331 0 cellNo=803
rlabel pdiffusion 45 -1331 45 -1331 0 feedthrough
rlabel pdiffusion 52 -1331 52 -1331 0 feedthrough
rlabel pdiffusion 59 -1331 59 -1331 0 feedthrough
rlabel pdiffusion 66 -1331 66 -1331 0 feedthrough
rlabel pdiffusion 73 -1331 73 -1331 0 cellNo=608
rlabel pdiffusion 80 -1331 80 -1331 0 cellNo=672
rlabel pdiffusion 87 -1331 87 -1331 0 feedthrough
rlabel pdiffusion 94 -1331 94 -1331 0 feedthrough
rlabel pdiffusion 101 -1331 101 -1331 0 feedthrough
rlabel pdiffusion 108 -1331 108 -1331 0 feedthrough
rlabel pdiffusion 115 -1331 115 -1331 0 feedthrough
rlabel pdiffusion 122 -1331 122 -1331 0 feedthrough
rlabel pdiffusion 129 -1331 129 -1331 0 cellNo=412
rlabel pdiffusion 136 -1331 136 -1331 0 cellNo=622
rlabel pdiffusion 143 -1331 143 -1331 0 feedthrough
rlabel pdiffusion 150 -1331 150 -1331 0 cellNo=129
rlabel pdiffusion 157 -1331 157 -1331 0 feedthrough
rlabel pdiffusion 164 -1331 164 -1331 0 feedthrough
rlabel pdiffusion 171 -1331 171 -1331 0 cellNo=308
rlabel pdiffusion 178 -1331 178 -1331 0 cellNo=561
rlabel pdiffusion 185 -1331 185 -1331 0 feedthrough
rlabel pdiffusion 192 -1331 192 -1331 0 feedthrough
rlabel pdiffusion 199 -1331 199 -1331 0 feedthrough
rlabel pdiffusion 206 -1331 206 -1331 0 cellNo=477
rlabel pdiffusion 213 -1331 213 -1331 0 feedthrough
rlabel pdiffusion 220 -1331 220 -1331 0 feedthrough
rlabel pdiffusion 227 -1331 227 -1331 0 feedthrough
rlabel pdiffusion 234 -1331 234 -1331 0 cellNo=335
rlabel pdiffusion 241 -1331 241 -1331 0 feedthrough
rlabel pdiffusion 248 -1331 248 -1331 0 feedthrough
rlabel pdiffusion 255 -1331 255 -1331 0 feedthrough
rlabel pdiffusion 262 -1331 262 -1331 0 feedthrough
rlabel pdiffusion 269 -1331 269 -1331 0 feedthrough
rlabel pdiffusion 276 -1331 276 -1331 0 feedthrough
rlabel pdiffusion 283 -1331 283 -1331 0 cellNo=544
rlabel pdiffusion 290 -1331 290 -1331 0 feedthrough
rlabel pdiffusion 297 -1331 297 -1331 0 cellNo=71
rlabel pdiffusion 304 -1331 304 -1331 0 cellNo=736
rlabel pdiffusion 311 -1331 311 -1331 0 feedthrough
rlabel pdiffusion 318 -1331 318 -1331 0 feedthrough
rlabel pdiffusion 325 -1331 325 -1331 0 cellNo=373
rlabel pdiffusion 332 -1331 332 -1331 0 feedthrough
rlabel pdiffusion 339 -1331 339 -1331 0 cellNo=87
rlabel pdiffusion 346 -1331 346 -1331 0 feedthrough
rlabel pdiffusion 353 -1331 353 -1331 0 cellNo=868
rlabel pdiffusion 360 -1331 360 -1331 0 cellNo=420
rlabel pdiffusion 367 -1331 367 -1331 0 cellNo=84
rlabel pdiffusion 374 -1331 374 -1331 0 cellNo=118
rlabel pdiffusion 381 -1331 381 -1331 0 cellNo=35
rlabel pdiffusion 388 -1331 388 -1331 0 cellNo=952
rlabel pdiffusion 395 -1331 395 -1331 0 cellNo=968
rlabel pdiffusion 402 -1331 402 -1331 0 feedthrough
rlabel pdiffusion 409 -1331 409 -1331 0 cellNo=799
rlabel pdiffusion 416 -1331 416 -1331 0 feedthrough
rlabel pdiffusion 423 -1331 423 -1331 0 cellNo=540
rlabel pdiffusion 430 -1331 430 -1331 0 feedthrough
rlabel pdiffusion 437 -1331 437 -1331 0 feedthrough
rlabel pdiffusion 444 -1331 444 -1331 0 feedthrough
rlabel pdiffusion 451 -1331 451 -1331 0 cellNo=551
rlabel pdiffusion 458 -1331 458 -1331 0 feedthrough
rlabel pdiffusion 465 -1331 465 -1331 0 cellNo=575
rlabel pdiffusion 472 -1331 472 -1331 0 cellNo=76
rlabel pdiffusion 479 -1331 479 -1331 0 cellNo=769
rlabel pdiffusion 486 -1331 486 -1331 0 feedthrough
rlabel pdiffusion 493 -1331 493 -1331 0 feedthrough
rlabel pdiffusion 500 -1331 500 -1331 0 cellNo=987
rlabel pdiffusion 507 -1331 507 -1331 0 feedthrough
rlabel pdiffusion 514 -1331 514 -1331 0 feedthrough
rlabel pdiffusion 521 -1331 521 -1331 0 feedthrough
rlabel pdiffusion 528 -1331 528 -1331 0 feedthrough
rlabel pdiffusion 535 -1331 535 -1331 0 feedthrough
rlabel pdiffusion 542 -1331 542 -1331 0 feedthrough
rlabel pdiffusion 549 -1331 549 -1331 0 feedthrough
rlabel pdiffusion 556 -1331 556 -1331 0 feedthrough
rlabel pdiffusion 563 -1331 563 -1331 0 feedthrough
rlabel pdiffusion 570 -1331 570 -1331 0 feedthrough
rlabel pdiffusion 577 -1331 577 -1331 0 feedthrough
rlabel pdiffusion 584 -1331 584 -1331 0 feedthrough
rlabel pdiffusion 591 -1331 591 -1331 0 feedthrough
rlabel pdiffusion 598 -1331 598 -1331 0 feedthrough
rlabel pdiffusion 605 -1331 605 -1331 0 feedthrough
rlabel pdiffusion 612 -1331 612 -1331 0 feedthrough
rlabel pdiffusion 619 -1331 619 -1331 0 feedthrough
rlabel pdiffusion 626 -1331 626 -1331 0 feedthrough
rlabel pdiffusion 633 -1331 633 -1331 0 feedthrough
rlabel pdiffusion 640 -1331 640 -1331 0 feedthrough
rlabel pdiffusion 647 -1331 647 -1331 0 cellNo=930
rlabel pdiffusion 654 -1331 654 -1331 0 feedthrough
rlabel pdiffusion 661 -1331 661 -1331 0 cellNo=880
rlabel pdiffusion 668 -1331 668 -1331 0 cellNo=866
rlabel pdiffusion 675 -1331 675 -1331 0 feedthrough
rlabel pdiffusion 682 -1331 682 -1331 0 feedthrough
rlabel pdiffusion 703 -1331 703 -1331 0 feedthrough
rlabel pdiffusion 31 -1390 31 -1390 0 cellNo=232
rlabel pdiffusion 38 -1390 38 -1390 0 feedthrough
rlabel pdiffusion 45 -1390 45 -1390 0 feedthrough
rlabel pdiffusion 52 -1390 52 -1390 0 feedthrough
rlabel pdiffusion 59 -1390 59 -1390 0 feedthrough
rlabel pdiffusion 66 -1390 66 -1390 0 feedthrough
rlabel pdiffusion 73 -1390 73 -1390 0 feedthrough
rlabel pdiffusion 80 -1390 80 -1390 0 feedthrough
rlabel pdiffusion 87 -1390 87 -1390 0 feedthrough
rlabel pdiffusion 94 -1390 94 -1390 0 feedthrough
rlabel pdiffusion 101 -1390 101 -1390 0 cellNo=812
rlabel pdiffusion 108 -1390 108 -1390 0 feedthrough
rlabel pdiffusion 115 -1390 115 -1390 0 feedthrough
rlabel pdiffusion 122 -1390 122 -1390 0 cellNo=690
rlabel pdiffusion 129 -1390 129 -1390 0 feedthrough
rlabel pdiffusion 136 -1390 136 -1390 0 cellNo=414
rlabel pdiffusion 143 -1390 143 -1390 0 cellNo=181
rlabel pdiffusion 150 -1390 150 -1390 0 feedthrough
rlabel pdiffusion 157 -1390 157 -1390 0 cellNo=673
rlabel pdiffusion 164 -1390 164 -1390 0 feedthrough
rlabel pdiffusion 171 -1390 171 -1390 0 feedthrough
rlabel pdiffusion 178 -1390 178 -1390 0 feedthrough
rlabel pdiffusion 185 -1390 185 -1390 0 cellNo=911
rlabel pdiffusion 192 -1390 192 -1390 0 cellNo=18
rlabel pdiffusion 199 -1390 199 -1390 0 cellNo=841
rlabel pdiffusion 206 -1390 206 -1390 0 cellNo=620
rlabel pdiffusion 213 -1390 213 -1390 0 feedthrough
rlabel pdiffusion 220 -1390 220 -1390 0 cellNo=747
rlabel pdiffusion 227 -1390 227 -1390 0 feedthrough
rlabel pdiffusion 234 -1390 234 -1390 0 cellNo=936
rlabel pdiffusion 241 -1390 241 -1390 0 cellNo=707
rlabel pdiffusion 248 -1390 248 -1390 0 cellNo=172
rlabel pdiffusion 255 -1390 255 -1390 0 feedthrough
rlabel pdiffusion 262 -1390 262 -1390 0 feedthrough
rlabel pdiffusion 269 -1390 269 -1390 0 feedthrough
rlabel pdiffusion 276 -1390 276 -1390 0 feedthrough
rlabel pdiffusion 283 -1390 283 -1390 0 cellNo=801
rlabel pdiffusion 290 -1390 290 -1390 0 feedthrough
rlabel pdiffusion 297 -1390 297 -1390 0 feedthrough
rlabel pdiffusion 304 -1390 304 -1390 0 feedthrough
rlabel pdiffusion 311 -1390 311 -1390 0 feedthrough
rlabel pdiffusion 318 -1390 318 -1390 0 feedthrough
rlabel pdiffusion 325 -1390 325 -1390 0 feedthrough
rlabel pdiffusion 332 -1390 332 -1390 0 feedthrough
rlabel pdiffusion 339 -1390 339 -1390 0 feedthrough
rlabel pdiffusion 346 -1390 346 -1390 0 cellNo=265
rlabel pdiffusion 353 -1390 353 -1390 0 feedthrough
rlabel pdiffusion 360 -1390 360 -1390 0 cellNo=776
rlabel pdiffusion 367 -1390 367 -1390 0 cellNo=566
rlabel pdiffusion 374 -1390 374 -1390 0 feedthrough
rlabel pdiffusion 381 -1390 381 -1390 0 cellNo=599
rlabel pdiffusion 388 -1390 388 -1390 0 cellNo=871
rlabel pdiffusion 395 -1390 395 -1390 0 feedthrough
rlabel pdiffusion 402 -1390 402 -1390 0 cellNo=374
rlabel pdiffusion 409 -1390 409 -1390 0 feedthrough
rlabel pdiffusion 416 -1390 416 -1390 0 cellNo=434
rlabel pdiffusion 423 -1390 423 -1390 0 cellNo=770
rlabel pdiffusion 430 -1390 430 -1390 0 cellNo=832
rlabel pdiffusion 437 -1390 437 -1390 0 feedthrough
rlabel pdiffusion 444 -1390 444 -1390 0 feedthrough
rlabel pdiffusion 451 -1390 451 -1390 0 feedthrough
rlabel pdiffusion 458 -1390 458 -1390 0 cellNo=431
rlabel pdiffusion 465 -1390 465 -1390 0 cellNo=925
rlabel pdiffusion 472 -1390 472 -1390 0 feedthrough
rlabel pdiffusion 479 -1390 479 -1390 0 cellNo=33
rlabel pdiffusion 486 -1390 486 -1390 0 feedthrough
rlabel pdiffusion 493 -1390 493 -1390 0 feedthrough
rlabel pdiffusion 500 -1390 500 -1390 0 feedthrough
rlabel pdiffusion 507 -1390 507 -1390 0 feedthrough
rlabel pdiffusion 514 -1390 514 -1390 0 feedthrough
rlabel pdiffusion 521 -1390 521 -1390 0 feedthrough
rlabel pdiffusion 528 -1390 528 -1390 0 feedthrough
rlabel pdiffusion 535 -1390 535 -1390 0 feedthrough
rlabel pdiffusion 542 -1390 542 -1390 0 feedthrough
rlabel pdiffusion 549 -1390 549 -1390 0 feedthrough
rlabel pdiffusion 556 -1390 556 -1390 0 feedthrough
rlabel pdiffusion 563 -1390 563 -1390 0 feedthrough
rlabel pdiffusion 570 -1390 570 -1390 0 feedthrough
rlabel pdiffusion 577 -1390 577 -1390 0 feedthrough
rlabel pdiffusion 584 -1390 584 -1390 0 feedthrough
rlabel pdiffusion 591 -1390 591 -1390 0 feedthrough
rlabel pdiffusion 598 -1390 598 -1390 0 cellNo=778
rlabel pdiffusion 605 -1390 605 -1390 0 feedthrough
rlabel pdiffusion 612 -1390 612 -1390 0 feedthrough
rlabel pdiffusion 619 -1390 619 -1390 0 cellNo=592
rlabel pdiffusion 626 -1390 626 -1390 0 feedthrough
rlabel pdiffusion 633 -1390 633 -1390 0 cellNo=660
rlabel pdiffusion 640 -1390 640 -1390 0 feedthrough
rlabel pdiffusion 647 -1390 647 -1390 0 feedthrough
rlabel pdiffusion 654 -1390 654 -1390 0 cellNo=810
rlabel pdiffusion 661 -1390 661 -1390 0 feedthrough
rlabel pdiffusion 668 -1390 668 -1390 0 feedthrough
rlabel pdiffusion 703 -1390 703 -1390 0 cellNo=63
rlabel pdiffusion 38 -1449 38 -1449 0 feedthrough
rlabel pdiffusion 45 -1449 45 -1449 0 feedthrough
rlabel pdiffusion 52 -1449 52 -1449 0 feedthrough
rlabel pdiffusion 59 -1449 59 -1449 0 feedthrough
rlabel pdiffusion 66 -1449 66 -1449 0 feedthrough
rlabel pdiffusion 73 -1449 73 -1449 0 feedthrough
rlabel pdiffusion 80 -1449 80 -1449 0 feedthrough
rlabel pdiffusion 87 -1449 87 -1449 0 feedthrough
rlabel pdiffusion 94 -1449 94 -1449 0 feedthrough
rlabel pdiffusion 101 -1449 101 -1449 0 cellNo=734
rlabel pdiffusion 108 -1449 108 -1449 0 feedthrough
rlabel pdiffusion 115 -1449 115 -1449 0 cellNo=86
rlabel pdiffusion 122 -1449 122 -1449 0 cellNo=774
rlabel pdiffusion 129 -1449 129 -1449 0 feedthrough
rlabel pdiffusion 136 -1449 136 -1449 0 cellNo=700
rlabel pdiffusion 143 -1449 143 -1449 0 cellNo=820
rlabel pdiffusion 150 -1449 150 -1449 0 feedthrough
rlabel pdiffusion 157 -1449 157 -1449 0 cellNo=927
rlabel pdiffusion 164 -1449 164 -1449 0 feedthrough
rlabel pdiffusion 171 -1449 171 -1449 0 feedthrough
rlabel pdiffusion 178 -1449 178 -1449 0 feedthrough
rlabel pdiffusion 185 -1449 185 -1449 0 cellNo=20
rlabel pdiffusion 192 -1449 192 -1449 0 feedthrough
rlabel pdiffusion 199 -1449 199 -1449 0 cellNo=385
rlabel pdiffusion 206 -1449 206 -1449 0 feedthrough
rlabel pdiffusion 213 -1449 213 -1449 0 cellNo=327
rlabel pdiffusion 220 -1449 220 -1449 0 feedthrough
rlabel pdiffusion 227 -1449 227 -1449 0 cellNo=971
rlabel pdiffusion 234 -1449 234 -1449 0 cellNo=441
rlabel pdiffusion 241 -1449 241 -1449 0 cellNo=706
rlabel pdiffusion 248 -1449 248 -1449 0 feedthrough
rlabel pdiffusion 255 -1449 255 -1449 0 feedthrough
rlabel pdiffusion 262 -1449 262 -1449 0 feedthrough
rlabel pdiffusion 269 -1449 269 -1449 0 cellNo=57
rlabel pdiffusion 276 -1449 276 -1449 0 feedthrough
rlabel pdiffusion 283 -1449 283 -1449 0 feedthrough
rlabel pdiffusion 290 -1449 290 -1449 0 feedthrough
rlabel pdiffusion 297 -1449 297 -1449 0 feedthrough
rlabel pdiffusion 304 -1449 304 -1449 0 feedthrough
rlabel pdiffusion 311 -1449 311 -1449 0 feedthrough
rlabel pdiffusion 318 -1449 318 -1449 0 feedthrough
rlabel pdiffusion 325 -1449 325 -1449 0 cellNo=417
rlabel pdiffusion 332 -1449 332 -1449 0 feedthrough
rlabel pdiffusion 339 -1449 339 -1449 0 feedthrough
rlabel pdiffusion 346 -1449 346 -1449 0 feedthrough
rlabel pdiffusion 353 -1449 353 -1449 0 cellNo=629
rlabel pdiffusion 360 -1449 360 -1449 0 cellNo=476
rlabel pdiffusion 367 -1449 367 -1449 0 cellNo=389
rlabel pdiffusion 374 -1449 374 -1449 0 cellNo=178
rlabel pdiffusion 381 -1449 381 -1449 0 feedthrough
rlabel pdiffusion 388 -1449 388 -1449 0 cellNo=692
rlabel pdiffusion 395 -1449 395 -1449 0 cellNo=787
rlabel pdiffusion 402 -1449 402 -1449 0 feedthrough
rlabel pdiffusion 409 -1449 409 -1449 0 feedthrough
rlabel pdiffusion 416 -1449 416 -1449 0 feedthrough
rlabel pdiffusion 423 -1449 423 -1449 0 feedthrough
rlabel pdiffusion 430 -1449 430 -1449 0 feedthrough
rlabel pdiffusion 437 -1449 437 -1449 0 cellNo=583
rlabel pdiffusion 444 -1449 444 -1449 0 cellNo=192
rlabel pdiffusion 451 -1449 451 -1449 0 cellNo=898
rlabel pdiffusion 458 -1449 458 -1449 0 feedthrough
rlabel pdiffusion 465 -1449 465 -1449 0 cellNo=938
rlabel pdiffusion 472 -1449 472 -1449 0 feedthrough
rlabel pdiffusion 479 -1449 479 -1449 0 cellNo=450
rlabel pdiffusion 486 -1449 486 -1449 0 feedthrough
rlabel pdiffusion 493 -1449 493 -1449 0 feedthrough
rlabel pdiffusion 500 -1449 500 -1449 0 feedthrough
rlabel pdiffusion 507 -1449 507 -1449 0 feedthrough
rlabel pdiffusion 514 -1449 514 -1449 0 feedthrough
rlabel pdiffusion 521 -1449 521 -1449 0 feedthrough
rlabel pdiffusion 528 -1449 528 -1449 0 feedthrough
rlabel pdiffusion 535 -1449 535 -1449 0 feedthrough
rlabel pdiffusion 542 -1449 542 -1449 0 feedthrough
rlabel pdiffusion 549 -1449 549 -1449 0 cellNo=722
rlabel pdiffusion 556 -1449 556 -1449 0 feedthrough
rlabel pdiffusion 563 -1449 563 -1449 0 cellNo=42
rlabel pdiffusion 570 -1449 570 -1449 0 cellNo=800
rlabel pdiffusion 577 -1449 577 -1449 0 feedthrough
rlabel pdiffusion 584 -1449 584 -1449 0 feedthrough
rlabel pdiffusion 591 -1449 591 -1449 0 feedthrough
rlabel pdiffusion 598 -1449 598 -1449 0 feedthrough
rlabel pdiffusion 605 -1449 605 -1449 0 feedthrough
rlabel pdiffusion 647 -1449 647 -1449 0 cellNo=295
rlabel pdiffusion 703 -1449 703 -1449 0 cellNo=856
rlabel pdiffusion 710 -1449 710 -1449 0 cellNo=13
rlabel pdiffusion 17 -1502 17 -1502 0 feedthrough
rlabel pdiffusion 24 -1502 24 -1502 0 cellNo=457
rlabel pdiffusion 31 -1502 31 -1502 0 feedthrough
rlabel pdiffusion 38 -1502 38 -1502 0 feedthrough
rlabel pdiffusion 45 -1502 45 -1502 0 cellNo=364
rlabel pdiffusion 52 -1502 52 -1502 0 cellNo=404
rlabel pdiffusion 59 -1502 59 -1502 0 feedthrough
rlabel pdiffusion 66 -1502 66 -1502 0 feedthrough
rlabel pdiffusion 73 -1502 73 -1502 0 feedthrough
rlabel pdiffusion 80 -1502 80 -1502 0 feedthrough
rlabel pdiffusion 87 -1502 87 -1502 0 cellNo=3
rlabel pdiffusion 94 -1502 94 -1502 0 feedthrough
rlabel pdiffusion 101 -1502 101 -1502 0 feedthrough
rlabel pdiffusion 108 -1502 108 -1502 0 cellNo=276
rlabel pdiffusion 115 -1502 115 -1502 0 feedthrough
rlabel pdiffusion 122 -1502 122 -1502 0 cellNo=482
rlabel pdiffusion 129 -1502 129 -1502 0 feedthrough
rlabel pdiffusion 136 -1502 136 -1502 0 feedthrough
rlabel pdiffusion 143 -1502 143 -1502 0 feedthrough
rlabel pdiffusion 150 -1502 150 -1502 0 cellNo=981
rlabel pdiffusion 157 -1502 157 -1502 0 cellNo=452
rlabel pdiffusion 164 -1502 164 -1502 0 cellNo=552
rlabel pdiffusion 171 -1502 171 -1502 0 cellNo=852
rlabel pdiffusion 178 -1502 178 -1502 0 cellNo=532
rlabel pdiffusion 185 -1502 185 -1502 0 cellNo=19
rlabel pdiffusion 192 -1502 192 -1502 0 feedthrough
rlabel pdiffusion 199 -1502 199 -1502 0 feedthrough
rlabel pdiffusion 206 -1502 206 -1502 0 cellNo=576
rlabel pdiffusion 213 -1502 213 -1502 0 feedthrough
rlabel pdiffusion 220 -1502 220 -1502 0 feedthrough
rlabel pdiffusion 227 -1502 227 -1502 0 cellNo=413
rlabel pdiffusion 234 -1502 234 -1502 0 cellNo=567
rlabel pdiffusion 241 -1502 241 -1502 0 cellNo=878
rlabel pdiffusion 248 -1502 248 -1502 0 cellNo=1
rlabel pdiffusion 255 -1502 255 -1502 0 feedthrough
rlabel pdiffusion 262 -1502 262 -1502 0 feedthrough
rlabel pdiffusion 269 -1502 269 -1502 0 cellNo=219
rlabel pdiffusion 276 -1502 276 -1502 0 feedthrough
rlabel pdiffusion 283 -1502 283 -1502 0 feedthrough
rlabel pdiffusion 290 -1502 290 -1502 0 cellNo=150
rlabel pdiffusion 297 -1502 297 -1502 0 feedthrough
rlabel pdiffusion 304 -1502 304 -1502 0 cellNo=895
rlabel pdiffusion 311 -1502 311 -1502 0 cellNo=713
rlabel pdiffusion 318 -1502 318 -1502 0 cellNo=409
rlabel pdiffusion 325 -1502 325 -1502 0 cellNo=56
rlabel pdiffusion 332 -1502 332 -1502 0 feedthrough
rlabel pdiffusion 339 -1502 339 -1502 0 feedthrough
rlabel pdiffusion 346 -1502 346 -1502 0 feedthrough
rlabel pdiffusion 353 -1502 353 -1502 0 feedthrough
rlabel pdiffusion 360 -1502 360 -1502 0 feedthrough
rlabel pdiffusion 367 -1502 367 -1502 0 cellNo=543
rlabel pdiffusion 374 -1502 374 -1502 0 feedthrough
rlabel pdiffusion 381 -1502 381 -1502 0 feedthrough
rlabel pdiffusion 388 -1502 388 -1502 0 feedthrough
rlabel pdiffusion 395 -1502 395 -1502 0 feedthrough
rlabel pdiffusion 402 -1502 402 -1502 0 feedthrough
rlabel pdiffusion 409 -1502 409 -1502 0 feedthrough
rlabel pdiffusion 416 -1502 416 -1502 0 feedthrough
rlabel pdiffusion 423 -1502 423 -1502 0 cellNo=267
rlabel pdiffusion 430 -1502 430 -1502 0 cellNo=949
rlabel pdiffusion 437 -1502 437 -1502 0 feedthrough
rlabel pdiffusion 444 -1502 444 -1502 0 feedthrough
rlabel pdiffusion 451 -1502 451 -1502 0 feedthrough
rlabel pdiffusion 458 -1502 458 -1502 0 feedthrough
rlabel pdiffusion 465 -1502 465 -1502 0 feedthrough
rlabel pdiffusion 472 -1502 472 -1502 0 feedthrough
rlabel pdiffusion 479 -1502 479 -1502 0 cellNo=798
rlabel pdiffusion 486 -1502 486 -1502 0 feedthrough
rlabel pdiffusion 493 -1502 493 -1502 0 feedthrough
rlabel pdiffusion 500 -1502 500 -1502 0 feedthrough
rlabel pdiffusion 507 -1502 507 -1502 0 feedthrough
rlabel pdiffusion 514 -1502 514 -1502 0 feedthrough
rlabel pdiffusion 521 -1502 521 -1502 0 feedthrough
rlabel pdiffusion 528 -1502 528 -1502 0 feedthrough
rlabel pdiffusion 535 -1502 535 -1502 0 feedthrough
rlabel pdiffusion 542 -1502 542 -1502 0 feedthrough
rlabel pdiffusion 549 -1502 549 -1502 0 feedthrough
rlabel pdiffusion 556 -1502 556 -1502 0 feedthrough
rlabel pdiffusion 563 -1502 563 -1502 0 cellNo=824
rlabel pdiffusion 570 -1502 570 -1502 0 feedthrough
rlabel pdiffusion 577 -1502 577 -1502 0 cellNo=864
rlabel pdiffusion 584 -1502 584 -1502 0 feedthrough
rlabel pdiffusion 591 -1502 591 -1502 0 feedthrough
rlabel pdiffusion 52 -1551 52 -1551 0 feedthrough
rlabel pdiffusion 59 -1551 59 -1551 0 cellNo=423
rlabel pdiffusion 66 -1551 66 -1551 0 feedthrough
rlabel pdiffusion 73 -1551 73 -1551 0 cellNo=929
rlabel pdiffusion 80 -1551 80 -1551 0 feedthrough
rlabel pdiffusion 87 -1551 87 -1551 0 feedthrough
rlabel pdiffusion 94 -1551 94 -1551 0 cellNo=919
rlabel pdiffusion 101 -1551 101 -1551 0 cellNo=347
rlabel pdiffusion 108 -1551 108 -1551 0 cellNo=901
rlabel pdiffusion 115 -1551 115 -1551 0 feedthrough
rlabel pdiffusion 122 -1551 122 -1551 0 feedthrough
rlabel pdiffusion 129 -1551 129 -1551 0 feedthrough
rlabel pdiffusion 136 -1551 136 -1551 0 feedthrough
rlabel pdiffusion 143 -1551 143 -1551 0 feedthrough
rlabel pdiffusion 150 -1551 150 -1551 0 cellNo=183
rlabel pdiffusion 157 -1551 157 -1551 0 cellNo=350
rlabel pdiffusion 164 -1551 164 -1551 0 feedthrough
rlabel pdiffusion 171 -1551 171 -1551 0 cellNo=193
rlabel pdiffusion 178 -1551 178 -1551 0 feedthrough
rlabel pdiffusion 185 -1551 185 -1551 0 feedthrough
rlabel pdiffusion 192 -1551 192 -1551 0 cellNo=410
rlabel pdiffusion 199 -1551 199 -1551 0 cellNo=530
rlabel pdiffusion 206 -1551 206 -1551 0 feedthrough
rlabel pdiffusion 213 -1551 213 -1551 0 feedthrough
rlabel pdiffusion 220 -1551 220 -1551 0 cellNo=641
rlabel pdiffusion 227 -1551 227 -1551 0 cellNo=299
rlabel pdiffusion 234 -1551 234 -1551 0 cellNo=296
rlabel pdiffusion 241 -1551 241 -1551 0 cellNo=222
rlabel pdiffusion 248 -1551 248 -1551 0 feedthrough
rlabel pdiffusion 255 -1551 255 -1551 0 feedthrough
rlabel pdiffusion 262 -1551 262 -1551 0 feedthrough
rlabel pdiffusion 269 -1551 269 -1551 0 feedthrough
rlabel pdiffusion 276 -1551 276 -1551 0 feedthrough
rlabel pdiffusion 283 -1551 283 -1551 0 cellNo=220
rlabel pdiffusion 290 -1551 290 -1551 0 cellNo=738
rlabel pdiffusion 297 -1551 297 -1551 0 feedthrough
rlabel pdiffusion 304 -1551 304 -1551 0 feedthrough
rlabel pdiffusion 311 -1551 311 -1551 0 feedthrough
rlabel pdiffusion 318 -1551 318 -1551 0 feedthrough
rlabel pdiffusion 325 -1551 325 -1551 0 cellNo=961
rlabel pdiffusion 332 -1551 332 -1551 0 feedthrough
rlabel pdiffusion 339 -1551 339 -1551 0 feedthrough
rlabel pdiffusion 346 -1551 346 -1551 0 feedthrough
rlabel pdiffusion 353 -1551 353 -1551 0 feedthrough
rlabel pdiffusion 360 -1551 360 -1551 0 feedthrough
rlabel pdiffusion 367 -1551 367 -1551 0 cellNo=872
rlabel pdiffusion 374 -1551 374 -1551 0 feedthrough
rlabel pdiffusion 381 -1551 381 -1551 0 cellNo=39
rlabel pdiffusion 388 -1551 388 -1551 0 cellNo=883
rlabel pdiffusion 395 -1551 395 -1551 0 feedthrough
rlabel pdiffusion 402 -1551 402 -1551 0 feedthrough
rlabel pdiffusion 409 -1551 409 -1551 0 feedthrough
rlabel pdiffusion 416 -1551 416 -1551 0 cellNo=387
rlabel pdiffusion 423 -1551 423 -1551 0 cellNo=956
rlabel pdiffusion 430 -1551 430 -1551 0 feedthrough
rlabel pdiffusion 437 -1551 437 -1551 0 feedthrough
rlabel pdiffusion 444 -1551 444 -1551 0 feedthrough
rlabel pdiffusion 451 -1551 451 -1551 0 feedthrough
rlabel pdiffusion 458 -1551 458 -1551 0 feedthrough
rlabel pdiffusion 465 -1551 465 -1551 0 feedthrough
rlabel pdiffusion 472 -1551 472 -1551 0 cellNo=846
rlabel pdiffusion 479 -1551 479 -1551 0 feedthrough
rlabel pdiffusion 486 -1551 486 -1551 0 cellNo=991
rlabel pdiffusion 493 -1551 493 -1551 0 feedthrough
rlabel pdiffusion 500 -1551 500 -1551 0 cellNo=786
rlabel pdiffusion 507 -1551 507 -1551 0 feedthrough
rlabel pdiffusion 514 -1551 514 -1551 0 feedthrough
rlabel pdiffusion 521 -1551 521 -1551 0 feedthrough
rlabel pdiffusion 528 -1551 528 -1551 0 feedthrough
rlabel pdiffusion 584 -1551 584 -1551 0 cellNo=677
rlabel pdiffusion 591 -1551 591 -1551 0 feedthrough
rlabel pdiffusion 73 -1588 73 -1588 0 cellNo=688
rlabel pdiffusion 80 -1588 80 -1588 0 feedthrough
rlabel pdiffusion 129 -1588 129 -1588 0 feedthrough
rlabel pdiffusion 136 -1588 136 -1588 0 feedthrough
rlabel pdiffusion 143 -1588 143 -1588 0 cellNo=484
rlabel pdiffusion 150 -1588 150 -1588 0 cellNo=857
rlabel pdiffusion 157 -1588 157 -1588 0 cellNo=686
rlabel pdiffusion 164 -1588 164 -1588 0 feedthrough
rlabel pdiffusion 171 -1588 171 -1588 0 feedthrough
rlabel pdiffusion 178 -1588 178 -1588 0 cellNo=893
rlabel pdiffusion 185 -1588 185 -1588 0 cellNo=657
rlabel pdiffusion 192 -1588 192 -1588 0 cellNo=742
rlabel pdiffusion 199 -1588 199 -1588 0 cellNo=626
rlabel pdiffusion 206 -1588 206 -1588 0 cellNo=331
rlabel pdiffusion 213 -1588 213 -1588 0 feedthrough
rlabel pdiffusion 220 -1588 220 -1588 0 cellNo=889
rlabel pdiffusion 227 -1588 227 -1588 0 cellNo=555
rlabel pdiffusion 234 -1588 234 -1588 0 feedthrough
rlabel pdiffusion 241 -1588 241 -1588 0 cellNo=644
rlabel pdiffusion 248 -1588 248 -1588 0 feedthrough
rlabel pdiffusion 255 -1588 255 -1588 0 feedthrough
rlabel pdiffusion 262 -1588 262 -1588 0 feedthrough
rlabel pdiffusion 269 -1588 269 -1588 0 cellNo=270
rlabel pdiffusion 276 -1588 276 -1588 0 feedthrough
rlabel pdiffusion 283 -1588 283 -1588 0 cellNo=982
rlabel pdiffusion 290 -1588 290 -1588 0 feedthrough
rlabel pdiffusion 297 -1588 297 -1588 0 feedthrough
rlabel pdiffusion 304 -1588 304 -1588 0 feedthrough
rlabel pdiffusion 311 -1588 311 -1588 0 cellNo=66
rlabel pdiffusion 318 -1588 318 -1588 0 cellNo=879
rlabel pdiffusion 325 -1588 325 -1588 0 feedthrough
rlabel pdiffusion 332 -1588 332 -1588 0 feedthrough
rlabel pdiffusion 339 -1588 339 -1588 0 cellNo=941
rlabel pdiffusion 346 -1588 346 -1588 0 cellNo=794
rlabel pdiffusion 353 -1588 353 -1588 0 feedthrough
rlabel pdiffusion 360 -1588 360 -1588 0 feedthrough
rlabel pdiffusion 367 -1588 367 -1588 0 cellNo=751
rlabel pdiffusion 374 -1588 374 -1588 0 feedthrough
rlabel pdiffusion 381 -1588 381 -1588 0 cellNo=701
rlabel pdiffusion 388 -1588 388 -1588 0 cellNo=862
rlabel pdiffusion 395 -1588 395 -1588 0 feedthrough
rlabel pdiffusion 402 -1588 402 -1588 0 feedthrough
rlabel pdiffusion 423 -1588 423 -1588 0 cellNo=806
rlabel pdiffusion 430 -1588 430 -1588 0 feedthrough
rlabel pdiffusion 437 -1588 437 -1588 0 feedthrough
rlabel pdiffusion 465 -1588 465 -1588 0 feedthrough
rlabel pdiffusion 472 -1588 472 -1588 0 feedthrough
rlabel pdiffusion 486 -1588 486 -1588 0 cellNo=395
rlabel pdiffusion 493 -1588 493 -1588 0 feedthrough
rlabel pdiffusion 507 -1588 507 -1588 0 cellNo=226
rlabel pdiffusion 514 -1588 514 -1588 0 feedthrough
rlabel pdiffusion 31 -1621 31 -1621 0 cellNo=950
rlabel pdiffusion 73 -1621 73 -1621 0 feedthrough
rlabel pdiffusion 80 -1621 80 -1621 0 cellNo=600
rlabel pdiffusion 87 -1621 87 -1621 0 cellNo=572
rlabel pdiffusion 94 -1621 94 -1621 0 feedthrough
rlabel pdiffusion 101 -1621 101 -1621 0 cellNo=585
rlabel pdiffusion 115 -1621 115 -1621 0 feedthrough
rlabel pdiffusion 122 -1621 122 -1621 0 cellNo=384
rlabel pdiffusion 129 -1621 129 -1621 0 cellNo=785
rlabel pdiffusion 136 -1621 136 -1621 0 feedthrough
rlabel pdiffusion 143 -1621 143 -1621 0 feedthrough
rlabel pdiffusion 150 -1621 150 -1621 0 cellNo=565
rlabel pdiffusion 157 -1621 157 -1621 0 feedthrough
rlabel pdiffusion 164 -1621 164 -1621 0 feedthrough
rlabel pdiffusion 171 -1621 171 -1621 0 cellNo=716
rlabel pdiffusion 178 -1621 178 -1621 0 cellNo=923
rlabel pdiffusion 192 -1621 192 -1621 0 cellNo=207
rlabel pdiffusion 199 -1621 199 -1621 0 cellNo=637
rlabel pdiffusion 206 -1621 206 -1621 0 feedthrough
rlabel pdiffusion 213 -1621 213 -1621 0 cellNo=829
rlabel pdiffusion 220 -1621 220 -1621 0 feedthrough
rlabel pdiffusion 227 -1621 227 -1621 0 feedthrough
rlabel pdiffusion 234 -1621 234 -1621 0 cellNo=685
rlabel pdiffusion 241 -1621 241 -1621 0 cellNo=120
rlabel pdiffusion 248 -1621 248 -1621 0 cellNo=280
rlabel pdiffusion 255 -1621 255 -1621 0 feedthrough
rlabel pdiffusion 262 -1621 262 -1621 0 cellNo=922
rlabel pdiffusion 269 -1621 269 -1621 0 cellNo=902
rlabel pdiffusion 276 -1621 276 -1621 0 cellNo=967
rlabel pdiffusion 283 -1621 283 -1621 0 cellNo=728
rlabel pdiffusion 290 -1621 290 -1621 0 feedthrough
rlabel pdiffusion 297 -1621 297 -1621 0 cellNo=72
rlabel pdiffusion 304 -1621 304 -1621 0 feedthrough
rlabel pdiffusion 311 -1621 311 -1621 0 feedthrough
rlabel pdiffusion 318 -1621 318 -1621 0 feedthrough
rlabel pdiffusion 325 -1621 325 -1621 0 feedthrough
rlabel pdiffusion 332 -1621 332 -1621 0 cellNo=826
rlabel pdiffusion 339 -1621 339 -1621 0 cellNo=523
rlabel pdiffusion 346 -1621 346 -1621 0 feedthrough
rlabel pdiffusion 353 -1621 353 -1621 0 feedthrough
rlabel pdiffusion 360 -1621 360 -1621 0 feedthrough
rlabel pdiffusion 367 -1621 367 -1621 0 feedthrough
rlabel pdiffusion 381 -1621 381 -1621 0 cellNo=762
rlabel pdiffusion 388 -1621 388 -1621 0 feedthrough
rlabel pdiffusion 395 -1621 395 -1621 0 feedthrough
rlabel pdiffusion 444 -1621 444 -1621 0 feedthrough
rlabel pdiffusion 465 -1621 465 -1621 0 cellNo=355
rlabel pdiffusion 472 -1621 472 -1621 0 feedthrough
rlabel pdiffusion 486 -1621 486 -1621 0 cellNo=128
rlabel pdiffusion 493 -1621 493 -1621 0 feedthrough
rlabel pdiffusion 31 -1650 31 -1650 0 cellNo=721
rlabel pdiffusion 38 -1650 38 -1650 0 feedthrough
rlabel pdiffusion 45 -1650 45 -1650 0 feedthrough
rlabel pdiffusion 52 -1650 52 -1650 0 feedthrough
rlabel pdiffusion 59 -1650 59 -1650 0 cellNo=746
rlabel pdiffusion 66 -1650 66 -1650 0 feedthrough
rlabel pdiffusion 73 -1650 73 -1650 0 feedthrough
rlabel pdiffusion 80 -1650 80 -1650 0 feedthrough
rlabel pdiffusion 87 -1650 87 -1650 0 feedthrough
rlabel pdiffusion 94 -1650 94 -1650 0 cellNo=562
rlabel pdiffusion 101 -1650 101 -1650 0 feedthrough
rlabel pdiffusion 108 -1650 108 -1650 0 cellNo=906
rlabel pdiffusion 115 -1650 115 -1650 0 cellNo=844
rlabel pdiffusion 122 -1650 122 -1650 0 cellNo=541
rlabel pdiffusion 129 -1650 129 -1650 0 cellNo=507
rlabel pdiffusion 136 -1650 136 -1650 0 cellNo=959
rlabel pdiffusion 143 -1650 143 -1650 0 cellNo=426
rlabel pdiffusion 150 -1650 150 -1650 0 feedthrough
rlabel pdiffusion 157 -1650 157 -1650 0 feedthrough
rlabel pdiffusion 164 -1650 164 -1650 0 feedthrough
rlabel pdiffusion 171 -1650 171 -1650 0 feedthrough
rlabel pdiffusion 178 -1650 178 -1650 0 feedthrough
rlabel pdiffusion 185 -1650 185 -1650 0 cellNo=661
rlabel pdiffusion 192 -1650 192 -1650 0 feedthrough
rlabel pdiffusion 199 -1650 199 -1650 0 cellNo=963
rlabel pdiffusion 206 -1650 206 -1650 0 cellNo=148
rlabel pdiffusion 213 -1650 213 -1650 0 cellNo=739
rlabel pdiffusion 220 -1650 220 -1650 0 cellNo=602
rlabel pdiffusion 227 -1650 227 -1650 0 cellNo=719
rlabel pdiffusion 234 -1650 234 -1650 0 cellNo=179
rlabel pdiffusion 241 -1650 241 -1650 0 cellNo=825
rlabel pdiffusion 248 -1650 248 -1650 0 feedthrough
rlabel pdiffusion 255 -1650 255 -1650 0 feedthrough
rlabel pdiffusion 262 -1650 262 -1650 0 feedthrough
rlabel pdiffusion 269 -1650 269 -1650 0 cellNo=696
rlabel pdiffusion 276 -1650 276 -1650 0 cellNo=218
rlabel pdiffusion 283 -1650 283 -1650 0 cellNo=974
rlabel pdiffusion 290 -1650 290 -1650 0 feedthrough
rlabel pdiffusion 297 -1650 297 -1650 0 feedthrough
rlabel pdiffusion 304 -1650 304 -1650 0 cellNo=926
rlabel pdiffusion 311 -1650 311 -1650 0 feedthrough
rlabel pdiffusion 318 -1650 318 -1650 0 feedthrough
rlabel pdiffusion 325 -1650 325 -1650 0 cellNo=996
rlabel pdiffusion 332 -1650 332 -1650 0 feedthrough
rlabel pdiffusion 339 -1650 339 -1650 0 feedthrough
rlabel pdiffusion 346 -1650 346 -1650 0 feedthrough
rlabel pdiffusion 353 -1650 353 -1650 0 feedthrough
rlabel pdiffusion 360 -1650 360 -1650 0 feedthrough
rlabel pdiffusion 367 -1650 367 -1650 0 feedthrough
rlabel pdiffusion 374 -1650 374 -1650 0 feedthrough
rlabel pdiffusion 381 -1650 381 -1650 0 feedthrough
rlabel pdiffusion 388 -1650 388 -1650 0 feedthrough
rlabel pdiffusion 395 -1650 395 -1650 0 cellNo=894
rlabel pdiffusion 402 -1650 402 -1650 0 cellNo=142
rlabel pdiffusion 3 -1685 3 -1685 0 cellNo=921
rlabel pdiffusion 17 -1685 17 -1685 0 cellNo=809
rlabel pdiffusion 24 -1685 24 -1685 0 feedthrough
rlabel pdiffusion 31 -1685 31 -1685 0 cellNo=538
rlabel pdiffusion 80 -1685 80 -1685 0 cellNo=625
rlabel pdiffusion 101 -1685 101 -1685 0 cellNo=687
rlabel pdiffusion 108 -1685 108 -1685 0 feedthrough
rlabel pdiffusion 115 -1685 115 -1685 0 cellNo=874
rlabel pdiffusion 122 -1685 122 -1685 0 feedthrough
rlabel pdiffusion 129 -1685 129 -1685 0 cellNo=668
rlabel pdiffusion 136 -1685 136 -1685 0 feedthrough
rlabel pdiffusion 143 -1685 143 -1685 0 cellNo=665
rlabel pdiffusion 150 -1685 150 -1685 0 feedthrough
rlabel pdiffusion 157 -1685 157 -1685 0 feedthrough
rlabel pdiffusion 164 -1685 164 -1685 0 feedthrough
rlabel pdiffusion 171 -1685 171 -1685 0 cellNo=917
rlabel pdiffusion 178 -1685 178 -1685 0 cellNo=140
rlabel pdiffusion 185 -1685 185 -1685 0 cellNo=946
rlabel pdiffusion 192 -1685 192 -1685 0 cellNo=646
rlabel pdiffusion 199 -1685 199 -1685 0 feedthrough
rlabel pdiffusion 206 -1685 206 -1685 0 cellNo=623
rlabel pdiffusion 213 -1685 213 -1685 0 cellNo=390
rlabel pdiffusion 220 -1685 220 -1685 0 cellNo=648
rlabel pdiffusion 227 -1685 227 -1685 0 cellNo=167
rlabel pdiffusion 234 -1685 234 -1685 0 feedthrough
rlabel pdiffusion 241 -1685 241 -1685 0 cellNo=983
rlabel pdiffusion 248 -1685 248 -1685 0 feedthrough
rlabel pdiffusion 255 -1685 255 -1685 0 cellNo=882
rlabel pdiffusion 262 -1685 262 -1685 0 cellNo=490
rlabel pdiffusion 269 -1685 269 -1685 0 feedthrough
rlabel pdiffusion 276 -1685 276 -1685 0 cellNo=931
rlabel pdiffusion 283 -1685 283 -1685 0 cellNo=827
rlabel pdiffusion 290 -1685 290 -1685 0 cellNo=909
rlabel pdiffusion 297 -1685 297 -1685 0 feedthrough
rlabel pdiffusion 304 -1685 304 -1685 0 feedthrough
rlabel pdiffusion 311 -1685 311 -1685 0 feedthrough
rlabel pdiffusion 318 -1685 318 -1685 0 cellNo=570
rlabel pdiffusion 325 -1685 325 -1685 0 feedthrough
rlabel pdiffusion 332 -1685 332 -1685 0 feedthrough
rlabel pdiffusion 339 -1685 339 -1685 0 feedthrough
rlabel pdiffusion 346 -1685 346 -1685 0 cellNo=26
rlabel pdiffusion 353 -1685 353 -1685 0 feedthrough
rlabel pdiffusion 360 -1685 360 -1685 0 cellNo=610
rlabel pdiffusion 367 -1685 367 -1685 0 cellNo=370
rlabel pdiffusion 374 -1685 374 -1685 0 feedthrough
rlabel pdiffusion 381 -1685 381 -1685 0 feedthrough
rlabel pdiffusion 388 -1685 388 -1685 0 cellNo=998
rlabel pdiffusion 395 -1685 395 -1685 0 feedthrough
rlabel pdiffusion 402 -1685 402 -1685 0 feedthrough
rlabel pdiffusion 3 -1708 3 -1708 0 cellNo=316
rlabel pdiffusion 10 -1708 10 -1708 0 feedthrough
rlabel pdiffusion 17 -1708 17 -1708 0 cellNo=1000
rlabel pdiffusion 31 -1708 31 -1708 0 cellNo=985
rlabel pdiffusion 80 -1708 80 -1708 0 cellNo=439
rlabel pdiffusion 87 -1708 87 -1708 0 cellNo=359
rlabel pdiffusion 94 -1708 94 -1708 0 cellNo=886
rlabel pdiffusion 101 -1708 101 -1708 0 cellNo=112
rlabel pdiffusion 115 -1708 115 -1708 0 cellNo=966
rlabel pdiffusion 122 -1708 122 -1708 0 cellNo=619
rlabel pdiffusion 129 -1708 129 -1708 0 cellNo=508
rlabel pdiffusion 136 -1708 136 -1708 0 feedthrough
rlabel pdiffusion 143 -1708 143 -1708 0 cellNo=990
rlabel pdiffusion 150 -1708 150 -1708 0 cellNo=621
rlabel pdiffusion 157 -1708 157 -1708 0 feedthrough
rlabel pdiffusion 164 -1708 164 -1708 0 feedthrough
rlabel pdiffusion 171 -1708 171 -1708 0 feedthrough
rlabel pdiffusion 178 -1708 178 -1708 0 feedthrough
rlabel pdiffusion 185 -1708 185 -1708 0 cellNo=999
rlabel pdiffusion 192 -1708 192 -1708 0 cellNo=522
rlabel pdiffusion 199 -1708 199 -1708 0 cellNo=202
rlabel pdiffusion 206 -1708 206 -1708 0 feedthrough
rlabel pdiffusion 213 -1708 213 -1708 0 feedthrough
rlabel pdiffusion 220 -1708 220 -1708 0 cellNo=147
rlabel pdiffusion 227 -1708 227 -1708 0 cellNo=831
rlabel pdiffusion 234 -1708 234 -1708 0 feedthrough
rlabel pdiffusion 241 -1708 241 -1708 0 cellNo=156
rlabel pdiffusion 255 -1708 255 -1708 0 cellNo=772
rlabel pdiffusion 276 -1708 276 -1708 0 cellNo=23
rlabel pdiffusion 283 -1708 283 -1708 0 cellNo=285
rlabel pdiffusion 290 -1708 290 -1708 0 cellNo=313
rlabel pdiffusion 297 -1708 297 -1708 0 cellNo=768
rlabel pdiffusion 304 -1708 304 -1708 0 cellNo=727
rlabel pdiffusion 311 -1708 311 -1708 0 feedthrough
rlabel pdiffusion 318 -1708 318 -1708 0 cellNo=818
rlabel pdiffusion 325 -1708 325 -1708 0 feedthrough
rlabel pdiffusion 353 -1708 353 -1708 0 cellNo=664
rlabel polysilicon 107 -10 107 -10 0 3
rlabel polysilicon 110 -10 110 -10 0 4
rlabel polysilicon 177 -4 177 -4 0 1
rlabel polysilicon 177 -10 177 -10 0 3
rlabel polysilicon 187 -4 187 -4 0 2
rlabel polysilicon 191 -10 191 -10 0 3
rlabel polysilicon 194 -10 194 -10 0 4
rlabel polysilicon 198 -4 198 -4 0 1
rlabel polysilicon 198 -10 198 -10 0 3
rlabel polysilicon 205 -4 205 -4 0 1
rlabel polysilicon 208 -4 208 -4 0 2
rlabel polysilicon 208 -10 208 -10 0 4
rlabel polysilicon 215 -4 215 -4 0 2
rlabel polysilicon 215 -10 215 -10 0 4
rlabel polysilicon 222 -4 222 -4 0 2
rlabel polysilicon 219 -10 219 -10 0 3
rlabel polysilicon 226 -10 226 -10 0 3
rlabel polysilicon 233 -4 233 -4 0 1
rlabel polysilicon 233 -10 233 -10 0 3
rlabel polysilicon 240 -4 240 -4 0 1
rlabel polysilicon 243 -4 243 -4 0 2
rlabel polysilicon 247 -4 247 -4 0 1
rlabel polysilicon 247 -10 247 -10 0 3
rlabel polysilicon 254 -4 254 -4 0 1
rlabel polysilicon 254 -10 254 -10 0 3
rlabel polysilicon 275 -4 275 -4 0 1
rlabel polysilicon 282 -4 282 -4 0 1
rlabel polysilicon 282 -10 282 -10 0 3
rlabel polysilicon 289 -4 289 -4 0 1
rlabel polysilicon 289 -10 289 -10 0 3
rlabel polysilicon 299 -4 299 -4 0 2
rlabel polysilicon 299 -10 299 -10 0 4
rlabel polysilicon 303 -10 303 -10 0 3
rlabel polysilicon 142 -23 142 -23 0 1
rlabel polysilicon 142 -29 142 -29 0 3
rlabel polysilicon 149 -23 149 -23 0 1
rlabel polysilicon 149 -29 149 -29 0 3
rlabel polysilicon 159 -23 159 -23 0 2
rlabel polysilicon 163 -23 163 -23 0 1
rlabel polysilicon 170 -23 170 -23 0 1
rlabel polysilicon 177 -29 177 -29 0 3
rlabel polysilicon 180 -29 180 -29 0 4
rlabel polysilicon 184 -23 184 -23 0 1
rlabel polysilicon 184 -29 184 -29 0 3
rlabel polysilicon 194 -23 194 -23 0 2
rlabel polysilicon 191 -29 191 -29 0 3
rlabel polysilicon 198 -23 198 -23 0 1
rlabel polysilicon 198 -29 198 -29 0 3
rlabel polysilicon 208 -23 208 -23 0 2
rlabel polysilicon 212 -29 212 -29 0 3
rlabel polysilicon 219 -23 219 -23 0 1
rlabel polysilicon 219 -29 219 -29 0 3
rlabel polysilicon 240 -23 240 -23 0 1
rlabel polysilicon 240 -29 240 -29 0 3
rlabel polysilicon 247 -23 247 -23 0 1
rlabel polysilicon 257 -29 257 -29 0 4
rlabel polysilicon 264 -23 264 -23 0 2
rlabel polysilicon 268 -23 268 -23 0 1
rlabel polysilicon 268 -29 268 -29 0 3
rlabel polysilicon 275 -23 275 -23 0 1
rlabel polysilicon 275 -29 275 -29 0 3
rlabel polysilicon 285 -29 285 -29 0 4
rlabel polysilicon 289 -23 289 -23 0 1
rlabel polysilicon 292 -23 292 -23 0 2
rlabel polysilicon 289 -29 289 -29 0 3
rlabel polysilicon 296 -23 296 -23 0 1
rlabel polysilicon 296 -29 296 -29 0 3
rlabel polysilicon 303 -29 303 -29 0 3
rlabel polysilicon 310 -23 310 -23 0 1
rlabel polysilicon 310 -29 310 -29 0 3
rlabel polysilicon 320 -29 320 -29 0 4
rlabel polysilicon 82 -42 82 -42 0 4
rlabel polysilicon 135 -36 135 -36 0 1
rlabel polysilicon 135 -42 135 -42 0 3
rlabel polysilicon 145 -36 145 -36 0 2
rlabel polysilicon 149 -36 149 -36 0 1
rlabel polysilicon 152 -36 152 -36 0 2
rlabel polysilicon 149 -42 149 -42 0 3
rlabel polysilicon 152 -42 152 -42 0 4
rlabel polysilicon 156 -36 156 -36 0 1
rlabel polysilicon 156 -42 156 -42 0 3
rlabel polysilicon 173 -42 173 -42 0 4
rlabel polysilicon 184 -36 184 -36 0 1
rlabel polysilicon 184 -42 184 -42 0 3
rlabel polysilicon 194 -42 194 -42 0 4
rlabel polysilicon 212 -42 212 -42 0 3
rlabel polysilicon 222 -42 222 -42 0 4
rlabel polysilicon 226 -36 226 -36 0 1
rlabel polysilicon 229 -42 229 -42 0 4
rlabel polysilicon 233 -36 233 -36 0 1
rlabel polysilicon 233 -42 233 -42 0 3
rlabel polysilicon 243 -36 243 -36 0 2
rlabel polysilicon 247 -36 247 -36 0 1
rlabel polysilicon 247 -42 247 -42 0 3
rlabel polysilicon 250 -42 250 -42 0 4
rlabel polysilicon 254 -36 254 -36 0 1
rlabel polysilicon 254 -42 254 -42 0 3
rlabel polysilicon 261 -36 261 -36 0 1
rlabel polysilicon 261 -42 261 -42 0 3
rlabel polysilicon 268 -42 268 -42 0 3
rlabel polysilicon 275 -36 275 -36 0 1
rlabel polysilicon 275 -42 275 -42 0 3
rlabel polysilicon 282 -36 282 -36 0 1
rlabel polysilicon 282 -42 282 -42 0 3
rlabel polysilicon 292 -36 292 -36 0 2
rlabel polysilicon 292 -42 292 -42 0 4
rlabel polysilicon 296 -36 296 -36 0 1
rlabel polysilicon 296 -42 296 -42 0 3
rlabel polysilicon 303 -36 303 -36 0 1
rlabel polysilicon 310 -42 310 -42 0 3
rlabel polysilicon 317 -36 317 -36 0 1
rlabel polysilicon 317 -42 317 -42 0 3
rlabel polysilicon 324 -36 324 -36 0 1
rlabel polysilicon 324 -42 324 -42 0 3
rlabel polysilicon 334 -42 334 -42 0 4
rlabel polysilicon 478 -36 478 -36 0 1
rlabel polysilicon 485 -36 485 -36 0 1
rlabel polysilicon 485 -42 485 -42 0 3
rlabel polysilicon 579 -36 579 -36 0 2
rlabel polysilicon 583 -36 583 -36 0 1
rlabel polysilicon 583 -42 583 -42 0 3
rlabel polysilicon 79 -59 79 -59 0 1
rlabel polysilicon 142 -65 142 -65 0 3
rlabel polysilicon 149 -59 149 -59 0 1
rlabel polysilicon 149 -65 149 -65 0 3
rlabel polysilicon 156 -59 156 -59 0 1
rlabel polysilicon 156 -65 156 -65 0 3
rlabel polysilicon 170 -59 170 -59 0 1
rlabel polysilicon 170 -65 170 -65 0 3
rlabel polysilicon 177 -59 177 -59 0 1
rlabel polysilicon 177 -65 177 -65 0 3
rlabel polysilicon 184 -59 184 -59 0 1
rlabel polysilicon 194 -59 194 -59 0 2
rlabel polysilicon 198 -65 198 -65 0 3
rlabel polysilicon 205 -59 205 -59 0 1
rlabel polysilicon 205 -65 205 -65 0 3
rlabel polysilicon 212 -59 212 -59 0 1
rlabel polysilicon 215 -59 215 -59 0 2
rlabel polysilicon 219 -59 219 -59 0 1
rlabel polysilicon 219 -65 219 -65 0 3
rlabel polysilicon 226 -59 226 -59 0 1
rlabel polysilicon 226 -65 226 -65 0 3
rlabel polysilicon 233 -59 233 -59 0 1
rlabel polysilicon 236 -65 236 -65 0 4
rlabel polysilicon 240 -59 240 -59 0 1
rlabel polysilicon 243 -59 243 -59 0 2
rlabel polysilicon 240 -65 240 -65 0 3
rlabel polysilicon 247 -59 247 -59 0 1
rlabel polysilicon 247 -65 247 -65 0 3
rlabel polysilicon 254 -59 254 -59 0 1
rlabel polysilicon 254 -65 254 -65 0 3
rlabel polysilicon 261 -59 261 -59 0 1
rlabel polysilicon 261 -65 261 -65 0 3
rlabel polysilicon 268 -59 268 -59 0 1
rlabel polysilicon 268 -65 268 -65 0 3
rlabel polysilicon 275 -59 275 -59 0 1
rlabel polysilicon 275 -65 275 -65 0 3
rlabel polysilicon 282 -59 282 -59 0 1
rlabel polysilicon 289 -59 289 -59 0 1
rlabel polysilicon 289 -65 289 -65 0 3
rlabel polysilicon 296 -59 296 -59 0 1
rlabel polysilicon 296 -65 296 -65 0 3
rlabel polysilicon 306 -65 306 -65 0 4
rlabel polysilicon 310 -65 310 -65 0 3
rlabel polysilicon 317 -59 317 -59 0 1
rlabel polysilicon 320 -59 320 -59 0 2
rlabel polysilicon 320 -65 320 -65 0 4
rlabel polysilicon 324 -59 324 -59 0 1
rlabel polysilicon 324 -65 324 -65 0 3
rlabel polysilicon 338 -59 338 -59 0 1
rlabel polysilicon 341 -59 341 -59 0 2
rlabel polysilicon 345 -59 345 -59 0 1
rlabel polysilicon 345 -65 345 -65 0 3
rlabel polysilicon 352 -59 352 -59 0 1
rlabel polysilicon 352 -65 352 -65 0 3
rlabel polysilicon 362 -59 362 -59 0 2
rlabel polysilicon 467 -59 467 -59 0 2
rlabel polysilicon 471 -59 471 -59 0 1
rlabel polysilicon 471 -65 471 -65 0 3
rlabel polysilicon 478 -59 478 -59 0 1
rlabel polysilicon 478 -65 478 -65 0 3
rlabel polysilicon 576 -59 576 -59 0 1
rlabel polysilicon 576 -65 576 -65 0 3
rlabel polysilicon 121 -88 121 -88 0 3
rlabel polysilicon 138 -82 138 -82 0 2
rlabel polysilicon 142 -82 142 -82 0 1
rlabel polysilicon 142 -88 142 -88 0 3
rlabel polysilicon 149 -82 149 -82 0 1
rlabel polysilicon 149 -88 149 -88 0 3
rlabel polysilicon 159 -88 159 -88 0 4
rlabel polysilicon 163 -82 163 -82 0 1
rlabel polysilicon 166 -82 166 -82 0 2
rlabel polysilicon 166 -88 166 -88 0 4
rlabel polysilicon 170 -82 170 -82 0 1
rlabel polysilicon 170 -88 170 -88 0 3
rlabel polysilicon 177 -82 177 -82 0 1
rlabel polysilicon 177 -88 177 -88 0 3
rlabel polysilicon 187 -88 187 -88 0 4
rlabel polysilicon 194 -88 194 -88 0 4
rlabel polysilicon 198 -82 198 -82 0 1
rlabel polysilicon 201 -88 201 -88 0 4
rlabel polysilicon 205 -82 205 -82 0 1
rlabel polysilicon 205 -88 205 -88 0 3
rlabel polysilicon 212 -82 212 -82 0 1
rlabel polysilicon 212 -88 212 -88 0 3
rlabel polysilicon 219 -82 219 -82 0 1
rlabel polysilicon 219 -88 219 -88 0 3
rlabel polysilicon 226 -82 226 -82 0 1
rlabel polysilicon 226 -88 226 -88 0 3
rlabel polysilicon 233 -82 233 -82 0 1
rlabel polysilicon 233 -88 233 -88 0 3
rlabel polysilicon 240 -82 240 -82 0 1
rlabel polysilicon 243 -82 243 -82 0 2
rlabel polysilicon 240 -88 240 -88 0 3
rlabel polysilicon 243 -88 243 -88 0 4
rlabel polysilicon 247 -82 247 -82 0 1
rlabel polysilicon 247 -88 247 -88 0 3
rlabel polysilicon 254 -82 254 -82 0 1
rlabel polysilicon 254 -88 254 -88 0 3
rlabel polysilicon 261 -82 261 -82 0 1
rlabel polysilicon 261 -88 261 -88 0 3
rlabel polysilicon 268 -82 268 -82 0 1
rlabel polysilicon 271 -88 271 -88 0 4
rlabel polysilicon 275 -82 275 -82 0 1
rlabel polysilicon 278 -82 278 -82 0 2
rlabel polysilicon 282 -82 282 -82 0 1
rlabel polysilicon 282 -88 282 -88 0 3
rlabel polysilicon 289 -82 289 -82 0 1
rlabel polysilicon 296 -82 296 -82 0 1
rlabel polysilicon 296 -88 296 -88 0 3
rlabel polysilicon 303 -82 303 -82 0 1
rlabel polysilicon 310 -88 310 -88 0 3
rlabel polysilicon 317 -82 317 -82 0 1
rlabel polysilicon 317 -88 317 -88 0 3
rlabel polysilicon 324 -82 324 -82 0 1
rlabel polysilicon 324 -88 324 -88 0 3
rlabel polysilicon 338 -82 338 -82 0 1
rlabel polysilicon 338 -88 338 -88 0 3
rlabel polysilicon 345 -82 345 -82 0 1
rlabel polysilicon 345 -88 345 -88 0 3
rlabel polysilicon 348 -88 348 -88 0 4
rlabel polysilicon 352 -82 352 -82 0 1
rlabel polysilicon 352 -88 352 -88 0 3
rlabel polysilicon 471 -82 471 -82 0 1
rlabel polysilicon 474 -82 474 -82 0 2
rlabel polysilicon 478 -82 478 -82 0 1
rlabel polysilicon 478 -88 478 -88 0 3
rlabel polysilicon 485 -82 485 -82 0 1
rlabel polysilicon 485 -88 485 -88 0 3
rlabel polysilicon 576 -82 576 -82 0 1
rlabel polysilicon 576 -88 576 -88 0 3
rlabel polysilicon 107 -113 107 -113 0 1
rlabel polysilicon 107 -119 107 -119 0 3
rlabel polysilicon 121 -113 121 -113 0 1
rlabel polysilicon 124 -119 124 -119 0 4
rlabel polysilicon 128 -113 128 -113 0 1
rlabel polysilicon 135 -113 135 -113 0 1
rlabel polysilicon 135 -119 135 -119 0 3
rlabel polysilicon 142 -113 142 -113 0 1
rlabel polysilicon 145 -113 145 -113 0 2
rlabel polysilicon 145 -119 145 -119 0 4
rlabel polysilicon 152 -113 152 -113 0 2
rlabel polysilicon 156 -113 156 -113 0 1
rlabel polysilicon 156 -119 156 -119 0 3
rlabel polysilicon 163 -113 163 -113 0 1
rlabel polysilicon 163 -119 163 -119 0 3
rlabel polysilicon 170 -119 170 -119 0 3
rlabel polysilicon 173 -119 173 -119 0 4
rlabel polysilicon 180 -113 180 -113 0 2
rlabel polysilicon 184 -113 184 -113 0 1
rlabel polysilicon 184 -119 184 -119 0 3
rlabel polysilicon 191 -113 191 -113 0 1
rlabel polysilicon 191 -119 191 -119 0 3
rlabel polysilicon 198 -113 198 -113 0 1
rlabel polysilicon 198 -119 198 -119 0 3
rlabel polysilicon 205 -119 205 -119 0 3
rlabel polysilicon 208 -119 208 -119 0 4
rlabel polysilicon 212 -113 212 -113 0 1
rlabel polysilicon 219 -113 219 -113 0 1
rlabel polysilicon 222 -113 222 -113 0 2
rlabel polysilicon 219 -119 219 -119 0 3
rlabel polysilicon 222 -119 222 -119 0 4
rlabel polysilicon 226 -113 226 -113 0 1
rlabel polysilicon 226 -119 226 -119 0 3
rlabel polysilicon 233 -113 233 -113 0 1
rlabel polysilicon 233 -119 233 -119 0 3
rlabel polysilicon 243 -113 243 -113 0 2
rlabel polysilicon 240 -119 240 -119 0 3
rlabel polysilicon 243 -119 243 -119 0 4
rlabel polysilicon 250 -113 250 -113 0 2
rlabel polysilicon 254 -113 254 -113 0 1
rlabel polysilicon 257 -113 257 -113 0 2
rlabel polysilicon 257 -119 257 -119 0 4
rlabel polysilicon 261 -113 261 -113 0 1
rlabel polysilicon 261 -119 261 -119 0 3
rlabel polysilicon 268 -113 268 -113 0 1
rlabel polysilicon 268 -119 268 -119 0 3
rlabel polysilicon 275 -113 275 -113 0 1
rlabel polysilicon 275 -119 275 -119 0 3
rlabel polysilicon 278 -119 278 -119 0 4
rlabel polysilicon 282 -113 282 -113 0 1
rlabel polysilicon 282 -119 282 -119 0 3
rlabel polysilicon 289 -113 289 -113 0 1
rlabel polysilicon 289 -119 289 -119 0 3
rlabel polysilicon 296 -113 296 -113 0 1
rlabel polysilicon 296 -119 296 -119 0 3
rlabel polysilicon 303 -113 303 -113 0 1
rlabel polysilicon 303 -119 303 -119 0 3
rlabel polysilicon 310 -113 310 -113 0 1
rlabel polysilicon 310 -119 310 -119 0 3
rlabel polysilicon 317 -113 317 -113 0 1
rlabel polysilicon 320 -113 320 -113 0 2
rlabel polysilicon 324 -113 324 -113 0 1
rlabel polysilicon 324 -119 324 -119 0 3
rlabel polysilicon 331 -113 331 -113 0 1
rlabel polysilicon 331 -119 331 -119 0 3
rlabel polysilicon 338 -113 338 -113 0 1
rlabel polysilicon 341 -113 341 -113 0 2
rlabel polysilicon 345 -113 345 -113 0 1
rlabel polysilicon 345 -119 345 -119 0 3
rlabel polysilicon 352 -113 352 -113 0 1
rlabel polysilicon 352 -119 352 -119 0 3
rlabel polysilicon 359 -113 359 -113 0 1
rlabel polysilicon 359 -119 359 -119 0 3
rlabel polysilicon 366 -113 366 -113 0 1
rlabel polysilicon 366 -119 366 -119 0 3
rlabel polysilicon 373 -113 373 -113 0 1
rlabel polysilicon 373 -119 373 -119 0 3
rlabel polysilicon 380 -113 380 -113 0 1
rlabel polysilicon 380 -119 380 -119 0 3
rlabel polysilicon 397 -113 397 -113 0 2
rlabel polysilicon 394 -119 394 -119 0 3
rlabel polysilicon 422 -113 422 -113 0 1
rlabel polysilicon 422 -119 422 -119 0 3
rlabel polysilicon 478 -113 478 -113 0 1
rlabel polysilicon 481 -113 481 -113 0 2
rlabel polysilicon 478 -119 478 -119 0 3
rlabel polysilicon 485 -113 485 -113 0 1
rlabel polysilicon 485 -119 485 -119 0 3
rlabel polysilicon 492 -113 492 -113 0 1
rlabel polysilicon 492 -119 492 -119 0 3
rlabel polysilicon 576 -113 576 -113 0 1
rlabel polysilicon 576 -119 576 -119 0 3
rlabel polysilicon 583 -113 583 -113 0 1
rlabel polysilicon 583 -119 583 -119 0 3
rlabel polysilicon 590 -113 590 -113 0 1
rlabel polysilicon 590 -119 590 -119 0 3
rlabel polysilicon 65 -152 65 -152 0 1
rlabel polysilicon 65 -158 65 -158 0 3
rlabel polysilicon 72 -152 72 -152 0 1
rlabel polysilicon 72 -158 72 -158 0 3
rlabel polysilicon 79 -158 79 -158 0 3
rlabel polysilicon 86 -152 86 -152 0 1
rlabel polysilicon 86 -158 86 -158 0 3
rlabel polysilicon 93 -152 93 -152 0 1
rlabel polysilicon 93 -158 93 -158 0 3
rlabel polysilicon 100 -152 100 -152 0 1
rlabel polysilicon 103 -158 103 -158 0 4
rlabel polysilicon 107 -152 107 -152 0 1
rlabel polysilicon 107 -158 107 -158 0 3
rlabel polysilicon 114 -152 114 -152 0 1
rlabel polysilicon 114 -158 114 -158 0 3
rlabel polysilicon 121 -158 121 -158 0 3
rlabel polysilicon 124 -158 124 -158 0 4
rlabel polysilicon 128 -152 128 -152 0 1
rlabel polysilicon 131 -152 131 -152 0 2
rlabel polysilicon 128 -158 128 -158 0 3
rlabel polysilicon 131 -158 131 -158 0 4
rlabel polysilicon 135 -152 135 -152 0 1
rlabel polysilicon 135 -158 135 -158 0 3
rlabel polysilicon 142 -158 142 -158 0 3
rlabel polysilicon 145 -158 145 -158 0 4
rlabel polysilicon 149 -152 149 -152 0 1
rlabel polysilicon 149 -158 149 -158 0 3
rlabel polysilicon 156 -152 156 -152 0 1
rlabel polysilicon 156 -158 156 -158 0 3
rlabel polysilicon 163 -158 163 -158 0 3
rlabel polysilicon 166 -158 166 -158 0 4
rlabel polysilicon 170 -152 170 -152 0 1
rlabel polysilicon 170 -158 170 -158 0 3
rlabel polysilicon 177 -152 177 -152 0 1
rlabel polysilicon 177 -158 177 -158 0 3
rlabel polysilicon 184 -152 184 -152 0 1
rlabel polysilicon 184 -158 184 -158 0 3
rlabel polysilicon 191 -152 191 -152 0 1
rlabel polysilicon 191 -158 191 -158 0 3
rlabel polysilicon 198 -152 198 -152 0 1
rlabel polysilicon 198 -158 198 -158 0 3
rlabel polysilicon 205 -152 205 -152 0 1
rlabel polysilicon 208 -152 208 -152 0 2
rlabel polysilicon 208 -158 208 -158 0 4
rlabel polysilicon 212 -152 212 -152 0 1
rlabel polysilicon 212 -158 212 -158 0 3
rlabel polysilicon 219 -152 219 -152 0 1
rlabel polysilicon 222 -152 222 -152 0 2
rlabel polysilicon 226 -152 226 -152 0 1
rlabel polysilicon 229 -152 229 -152 0 2
rlabel polysilicon 226 -158 226 -158 0 3
rlabel polysilicon 233 -152 233 -152 0 1
rlabel polysilicon 236 -152 236 -152 0 2
rlabel polysilicon 233 -158 233 -158 0 3
rlabel polysilicon 240 -152 240 -152 0 1
rlabel polysilicon 243 -152 243 -152 0 2
rlabel polysilicon 240 -158 240 -158 0 3
rlabel polysilicon 243 -158 243 -158 0 4
rlabel polysilicon 247 -152 247 -152 0 1
rlabel polysilicon 247 -158 247 -158 0 3
rlabel polysilicon 254 -152 254 -152 0 1
rlabel polysilicon 254 -158 254 -158 0 3
rlabel polysilicon 261 -152 261 -152 0 1
rlabel polysilicon 264 -152 264 -152 0 2
rlabel polysilicon 261 -158 261 -158 0 3
rlabel polysilicon 264 -158 264 -158 0 4
rlabel polysilicon 268 -152 268 -152 0 1
rlabel polysilicon 268 -158 268 -158 0 3
rlabel polysilicon 275 -152 275 -152 0 1
rlabel polysilicon 275 -158 275 -158 0 3
rlabel polysilicon 285 -152 285 -152 0 2
rlabel polysilicon 289 -152 289 -152 0 1
rlabel polysilicon 289 -158 289 -158 0 3
rlabel polysilicon 299 -152 299 -152 0 2
rlabel polysilicon 299 -158 299 -158 0 4
rlabel polysilicon 303 -152 303 -152 0 1
rlabel polysilicon 303 -158 303 -158 0 3
rlabel polysilicon 310 -152 310 -152 0 1
rlabel polysilicon 310 -158 310 -158 0 3
rlabel polysilicon 317 -152 317 -152 0 1
rlabel polysilicon 317 -158 317 -158 0 3
rlabel polysilicon 324 -152 324 -152 0 1
rlabel polysilicon 324 -158 324 -158 0 3
rlabel polysilicon 334 -152 334 -152 0 2
rlabel polysilicon 331 -158 331 -158 0 3
rlabel polysilicon 338 -152 338 -152 0 1
rlabel polysilicon 338 -158 338 -158 0 3
rlabel polysilicon 345 -152 345 -152 0 1
rlabel polysilicon 345 -158 345 -158 0 3
rlabel polysilicon 352 -152 352 -152 0 1
rlabel polysilicon 352 -158 352 -158 0 3
rlabel polysilicon 359 -152 359 -152 0 1
rlabel polysilicon 359 -158 359 -158 0 3
rlabel polysilicon 366 -152 366 -152 0 1
rlabel polysilicon 366 -158 366 -158 0 3
rlabel polysilicon 373 -152 373 -152 0 1
rlabel polysilicon 373 -158 373 -158 0 3
rlabel polysilicon 380 -152 380 -152 0 1
rlabel polysilicon 380 -158 380 -158 0 3
rlabel polysilicon 387 -152 387 -152 0 1
rlabel polysilicon 387 -158 387 -158 0 3
rlabel polysilicon 394 -152 394 -152 0 1
rlabel polysilicon 394 -158 394 -158 0 3
rlabel polysilicon 401 -152 401 -152 0 1
rlabel polysilicon 401 -158 401 -158 0 3
rlabel polysilicon 408 -158 408 -158 0 3
rlabel polysilicon 415 -152 415 -152 0 1
rlabel polysilicon 415 -158 415 -158 0 3
rlabel polysilicon 422 -152 422 -152 0 1
rlabel polysilicon 422 -158 422 -158 0 3
rlabel polysilicon 429 -152 429 -152 0 1
rlabel polysilicon 429 -158 429 -158 0 3
rlabel polysilicon 436 -152 436 -152 0 1
rlabel polysilicon 436 -158 436 -158 0 3
rlabel polysilicon 443 -152 443 -152 0 1
rlabel polysilicon 443 -158 443 -158 0 3
rlabel polysilicon 499 -152 499 -152 0 1
rlabel polysilicon 499 -158 499 -158 0 3
rlabel polysilicon 590 -152 590 -152 0 1
rlabel polysilicon 590 -158 590 -158 0 3
rlabel polysilicon 12 -207 12 -207 0 4
rlabel polysilicon 19 -201 19 -201 0 2
rlabel polysilicon 26 -201 26 -201 0 2
rlabel polysilicon 79 -201 79 -201 0 1
rlabel polysilicon 79 -207 79 -207 0 3
rlabel polysilicon 86 -201 86 -201 0 1
rlabel polysilicon 86 -207 86 -207 0 3
rlabel polysilicon 93 -201 93 -201 0 1
rlabel polysilicon 100 -201 100 -201 0 1
rlabel polysilicon 100 -207 100 -207 0 3
rlabel polysilicon 107 -201 107 -201 0 1
rlabel polysilicon 107 -207 107 -207 0 3
rlabel polysilicon 114 -201 114 -201 0 1
rlabel polysilicon 114 -207 114 -207 0 3
rlabel polysilicon 121 -201 121 -201 0 1
rlabel polysilicon 128 -201 128 -201 0 1
rlabel polysilicon 128 -207 128 -207 0 3
rlabel polysilicon 135 -201 135 -201 0 1
rlabel polysilicon 135 -207 135 -207 0 3
rlabel polysilicon 142 -201 142 -201 0 1
rlabel polysilicon 145 -207 145 -207 0 4
rlabel polysilicon 149 -201 149 -201 0 1
rlabel polysilicon 149 -207 149 -207 0 3
rlabel polysilicon 156 -201 156 -201 0 1
rlabel polysilicon 159 -201 159 -201 0 2
rlabel polysilicon 156 -207 156 -207 0 3
rlabel polysilicon 163 -201 163 -201 0 1
rlabel polysilicon 166 -207 166 -207 0 4
rlabel polysilicon 170 -201 170 -201 0 1
rlabel polysilicon 173 -207 173 -207 0 4
rlabel polysilicon 177 -201 177 -201 0 1
rlabel polysilicon 180 -201 180 -201 0 2
rlabel polysilicon 184 -207 184 -207 0 3
rlabel polysilicon 191 -201 191 -201 0 1
rlabel polysilicon 191 -207 191 -207 0 3
rlabel polysilicon 198 -207 198 -207 0 3
rlabel polysilicon 201 -207 201 -207 0 4
rlabel polysilicon 205 -201 205 -201 0 1
rlabel polysilicon 205 -207 205 -207 0 3
rlabel polysilicon 212 -201 212 -201 0 1
rlabel polysilicon 212 -207 212 -207 0 3
rlabel polysilicon 215 -207 215 -207 0 4
rlabel polysilicon 219 -201 219 -201 0 1
rlabel polysilicon 219 -207 219 -207 0 3
rlabel polysilicon 222 -207 222 -207 0 4
rlabel polysilicon 226 -201 226 -201 0 1
rlabel polysilicon 226 -207 226 -207 0 3
rlabel polysilicon 236 -201 236 -201 0 2
rlabel polysilicon 236 -207 236 -207 0 4
rlabel polysilicon 240 -201 240 -201 0 1
rlabel polysilicon 243 -201 243 -201 0 2
rlabel polysilicon 240 -207 240 -207 0 3
rlabel polysilicon 243 -207 243 -207 0 4
rlabel polysilicon 247 -201 247 -201 0 1
rlabel polysilicon 247 -207 247 -207 0 3
rlabel polysilicon 254 -201 254 -201 0 1
rlabel polysilicon 254 -207 254 -207 0 3
rlabel polysilicon 261 -201 261 -201 0 1
rlabel polysilicon 261 -207 261 -207 0 3
rlabel polysilicon 268 -201 268 -201 0 1
rlabel polysilicon 268 -207 268 -207 0 3
rlabel polysilicon 275 -201 275 -201 0 1
rlabel polysilicon 278 -201 278 -201 0 2
rlabel polysilicon 275 -207 275 -207 0 3
rlabel polysilicon 278 -207 278 -207 0 4
rlabel polysilicon 282 -201 282 -201 0 1
rlabel polysilicon 282 -207 282 -207 0 3
rlabel polysilicon 289 -201 289 -201 0 1
rlabel polysilicon 292 -207 292 -207 0 4
rlabel polysilicon 296 -201 296 -201 0 1
rlabel polysilicon 299 -201 299 -201 0 2
rlabel polysilicon 296 -207 296 -207 0 3
rlabel polysilicon 303 -201 303 -201 0 1
rlabel polysilicon 303 -207 303 -207 0 3
rlabel polysilicon 310 -201 310 -201 0 1
rlabel polysilicon 310 -207 310 -207 0 3
rlabel polysilicon 317 -201 317 -201 0 1
rlabel polysilicon 320 -201 320 -201 0 2
rlabel polysilicon 317 -207 317 -207 0 3
rlabel polysilicon 324 -201 324 -201 0 1
rlabel polysilicon 324 -207 324 -207 0 3
rlabel polysilicon 331 -201 331 -201 0 1
rlabel polysilicon 331 -207 331 -207 0 3
rlabel polysilicon 338 -201 338 -201 0 1
rlabel polysilicon 338 -207 338 -207 0 3
rlabel polysilicon 345 -201 345 -201 0 1
rlabel polysilicon 345 -207 345 -207 0 3
rlabel polysilicon 352 -201 352 -201 0 1
rlabel polysilicon 352 -207 352 -207 0 3
rlabel polysilicon 359 -201 359 -201 0 1
rlabel polysilicon 359 -207 359 -207 0 3
rlabel polysilicon 366 -201 366 -201 0 1
rlabel polysilicon 366 -207 366 -207 0 3
rlabel polysilicon 373 -201 373 -201 0 1
rlabel polysilicon 373 -207 373 -207 0 3
rlabel polysilicon 380 -201 380 -201 0 1
rlabel polysilicon 380 -207 380 -207 0 3
rlabel polysilicon 387 -201 387 -201 0 1
rlabel polysilicon 387 -207 387 -207 0 3
rlabel polysilicon 394 -201 394 -201 0 1
rlabel polysilicon 394 -207 394 -207 0 3
rlabel polysilicon 401 -201 401 -201 0 1
rlabel polysilicon 401 -207 401 -207 0 3
rlabel polysilicon 408 -201 408 -201 0 1
rlabel polysilicon 408 -207 408 -207 0 3
rlabel polysilicon 415 -201 415 -201 0 1
rlabel polysilicon 415 -207 415 -207 0 3
rlabel polysilicon 422 -201 422 -201 0 1
rlabel polysilicon 429 -201 429 -201 0 1
rlabel polysilicon 429 -207 429 -207 0 3
rlabel polysilicon 436 -201 436 -201 0 1
rlabel polysilicon 436 -207 436 -207 0 3
rlabel polysilicon 443 -201 443 -201 0 1
rlabel polysilicon 443 -207 443 -207 0 3
rlabel polysilicon 453 -207 453 -207 0 4
rlabel polysilicon 460 -201 460 -201 0 2
rlabel polysilicon 464 -201 464 -201 0 1
rlabel polysilicon 464 -207 464 -207 0 3
rlabel polysilicon 506 -201 506 -201 0 1
rlabel polysilicon 506 -207 506 -207 0 3
rlabel polysilicon 590 -201 590 -201 0 1
rlabel polysilicon 590 -207 590 -207 0 3
rlabel polysilicon 12 -242 12 -242 0 2
rlabel polysilicon 114 -242 114 -242 0 1
rlabel polysilicon 114 -248 114 -248 0 3
rlabel polysilicon 124 -248 124 -248 0 4
rlabel polysilicon 128 -242 128 -242 0 1
rlabel polysilicon 128 -248 128 -248 0 3
rlabel polysilicon 135 -242 135 -242 0 1
rlabel polysilicon 135 -248 135 -248 0 3
rlabel polysilicon 142 -242 142 -242 0 1
rlabel polysilicon 142 -248 142 -248 0 3
rlabel polysilicon 149 -242 149 -242 0 1
rlabel polysilicon 149 -248 149 -248 0 3
rlabel polysilicon 156 -242 156 -242 0 1
rlabel polysilicon 156 -248 156 -248 0 3
rlabel polysilicon 159 -248 159 -248 0 4
rlabel polysilicon 163 -242 163 -242 0 1
rlabel polysilicon 163 -248 163 -248 0 3
rlabel polysilicon 170 -248 170 -248 0 3
rlabel polysilicon 177 -242 177 -242 0 1
rlabel polysilicon 177 -248 177 -248 0 3
rlabel polysilicon 184 -242 184 -242 0 1
rlabel polysilicon 184 -248 184 -248 0 3
rlabel polysilicon 191 -242 191 -242 0 1
rlabel polysilicon 191 -248 191 -248 0 3
rlabel polysilicon 198 -242 198 -242 0 1
rlabel polysilicon 198 -248 198 -248 0 3
rlabel polysilicon 208 -248 208 -248 0 4
rlabel polysilicon 212 -242 212 -242 0 1
rlabel polysilicon 215 -242 215 -242 0 2
rlabel polysilicon 222 -242 222 -242 0 2
rlabel polysilicon 219 -248 219 -248 0 3
rlabel polysilicon 222 -248 222 -248 0 4
rlabel polysilicon 226 -242 226 -242 0 1
rlabel polysilicon 229 -248 229 -248 0 4
rlabel polysilicon 236 -242 236 -242 0 2
rlabel polysilicon 236 -248 236 -248 0 4
rlabel polysilicon 240 -242 240 -242 0 1
rlabel polysilicon 243 -242 243 -242 0 2
rlabel polysilicon 240 -248 240 -248 0 3
rlabel polysilicon 243 -248 243 -248 0 4
rlabel polysilicon 247 -242 247 -242 0 1
rlabel polysilicon 247 -248 247 -248 0 3
rlabel polysilicon 254 -242 254 -242 0 1
rlabel polysilicon 254 -248 254 -248 0 3
rlabel polysilicon 261 -242 261 -242 0 1
rlabel polysilicon 264 -242 264 -242 0 2
rlabel polysilicon 268 -242 268 -242 0 1
rlabel polysilicon 268 -248 268 -248 0 3
rlabel polysilicon 275 -242 275 -242 0 1
rlabel polysilicon 278 -242 278 -242 0 2
rlabel polysilicon 275 -248 275 -248 0 3
rlabel polysilicon 278 -248 278 -248 0 4
rlabel polysilicon 282 -242 282 -242 0 1
rlabel polysilicon 282 -248 282 -248 0 3
rlabel polysilicon 289 -242 289 -242 0 1
rlabel polysilicon 292 -242 292 -242 0 2
rlabel polysilicon 296 -242 296 -242 0 1
rlabel polysilicon 303 -242 303 -242 0 1
rlabel polysilicon 303 -248 303 -248 0 3
rlabel polysilicon 310 -242 310 -242 0 1
rlabel polysilicon 310 -248 310 -248 0 3
rlabel polysilicon 317 -242 317 -242 0 1
rlabel polysilicon 320 -242 320 -242 0 2
rlabel polysilicon 317 -248 317 -248 0 3
rlabel polysilicon 320 -248 320 -248 0 4
rlabel polysilicon 324 -242 324 -242 0 1
rlabel polysilicon 324 -248 324 -248 0 3
rlabel polysilicon 331 -242 331 -242 0 1
rlabel polysilicon 331 -248 331 -248 0 3
rlabel polysilicon 338 -242 338 -242 0 1
rlabel polysilicon 338 -248 338 -248 0 3
rlabel polysilicon 345 -242 345 -242 0 1
rlabel polysilicon 348 -242 348 -242 0 2
rlabel polysilicon 348 -248 348 -248 0 4
rlabel polysilicon 352 -242 352 -242 0 1
rlabel polysilicon 352 -248 352 -248 0 3
rlabel polysilicon 359 -242 359 -242 0 1
rlabel polysilicon 359 -248 359 -248 0 3
rlabel polysilicon 366 -242 366 -242 0 1
rlabel polysilicon 366 -248 366 -248 0 3
rlabel polysilicon 373 -242 373 -242 0 1
rlabel polysilicon 373 -248 373 -248 0 3
rlabel polysilicon 383 -242 383 -242 0 2
rlabel polysilicon 380 -248 380 -248 0 3
rlabel polysilicon 387 -242 387 -242 0 1
rlabel polysilicon 387 -248 387 -248 0 3
rlabel polysilicon 394 -242 394 -242 0 1
rlabel polysilicon 394 -248 394 -248 0 3
rlabel polysilicon 401 -242 401 -242 0 1
rlabel polysilicon 401 -248 401 -248 0 3
rlabel polysilicon 408 -242 408 -242 0 1
rlabel polysilicon 408 -248 408 -248 0 3
rlabel polysilicon 415 -242 415 -242 0 1
rlabel polysilicon 415 -248 415 -248 0 3
rlabel polysilicon 422 -242 422 -242 0 1
rlabel polysilicon 422 -248 422 -248 0 3
rlabel polysilicon 429 -242 429 -242 0 1
rlabel polysilicon 429 -248 429 -248 0 3
rlabel polysilicon 436 -242 436 -242 0 1
rlabel polysilicon 436 -248 436 -248 0 3
rlabel polysilicon 443 -242 443 -242 0 1
rlabel polysilicon 443 -248 443 -248 0 3
rlabel polysilicon 450 -242 450 -242 0 1
rlabel polysilicon 450 -248 450 -248 0 3
rlabel polysilicon 460 -242 460 -242 0 2
rlabel polysilicon 464 -248 464 -248 0 3
rlabel polysilicon 509 -242 509 -242 0 2
rlabel polysilicon 506 -248 506 -248 0 3
rlabel polysilicon 562 -242 562 -242 0 1
rlabel polysilicon 562 -248 562 -248 0 3
rlabel polysilicon 572 -242 572 -242 0 2
rlabel polysilicon 590 -242 590 -242 0 1
rlabel polysilicon 590 -248 590 -248 0 3
rlabel polysilicon 597 -248 597 -248 0 3
rlabel polysilicon 600 -248 600 -248 0 4
rlabel polysilicon 646 -248 646 -248 0 3
rlabel polysilicon 65 -283 65 -283 0 1
rlabel polysilicon 75 -289 75 -289 0 4
rlabel polysilicon 79 -283 79 -283 0 1
rlabel polysilicon 79 -289 79 -289 0 3
rlabel polysilicon 86 -283 86 -283 0 1
rlabel polysilicon 86 -289 86 -289 0 3
rlabel polysilicon 93 -283 93 -283 0 1
rlabel polysilicon 93 -289 93 -289 0 3
rlabel polysilicon 103 -289 103 -289 0 4
rlabel polysilicon 107 -283 107 -283 0 1
rlabel polysilicon 107 -289 107 -289 0 3
rlabel polysilicon 114 -283 114 -283 0 1
rlabel polysilicon 117 -289 117 -289 0 4
rlabel polysilicon 121 -283 121 -283 0 1
rlabel polysilicon 128 -283 128 -283 0 1
rlabel polysilicon 128 -289 128 -289 0 3
rlabel polysilicon 135 -283 135 -283 0 1
rlabel polysilicon 135 -289 135 -289 0 3
rlabel polysilicon 142 -283 142 -283 0 1
rlabel polysilicon 142 -289 142 -289 0 3
rlabel polysilicon 149 -283 149 -283 0 1
rlabel polysilicon 149 -289 149 -289 0 3
rlabel polysilicon 156 -283 156 -283 0 1
rlabel polysilicon 156 -289 156 -289 0 3
rlabel polysilicon 163 -283 163 -283 0 1
rlabel polysilicon 163 -289 163 -289 0 3
rlabel polysilicon 170 -283 170 -283 0 1
rlabel polysilicon 173 -283 173 -283 0 2
rlabel polysilicon 173 -289 173 -289 0 4
rlabel polysilicon 177 -283 177 -283 0 1
rlabel polysilicon 177 -289 177 -289 0 3
rlabel polysilicon 184 -283 184 -283 0 1
rlabel polysilicon 187 -283 187 -283 0 2
rlabel polysilicon 187 -289 187 -289 0 4
rlabel polysilicon 194 -283 194 -283 0 2
rlabel polysilicon 194 -289 194 -289 0 4
rlabel polysilicon 201 -283 201 -283 0 2
rlabel polysilicon 198 -289 198 -289 0 3
rlabel polysilicon 205 -283 205 -283 0 1
rlabel polysilicon 208 -283 208 -283 0 2
rlabel polysilicon 212 -289 212 -289 0 3
rlabel polysilicon 219 -283 219 -283 0 1
rlabel polysilicon 219 -289 219 -289 0 3
rlabel polysilicon 226 -283 226 -283 0 1
rlabel polysilicon 226 -289 226 -289 0 3
rlabel polysilicon 233 -283 233 -283 0 1
rlabel polysilicon 236 -283 236 -283 0 2
rlabel polysilicon 236 -289 236 -289 0 4
rlabel polysilicon 243 -283 243 -283 0 2
rlabel polysilicon 240 -289 240 -289 0 3
rlabel polysilicon 247 -283 247 -283 0 1
rlabel polysilicon 247 -289 247 -289 0 3
rlabel polysilicon 257 -283 257 -283 0 2
rlabel polysilicon 254 -289 254 -289 0 3
rlabel polysilicon 257 -289 257 -289 0 4
rlabel polysilicon 261 -283 261 -283 0 1
rlabel polysilicon 261 -289 261 -289 0 3
rlabel polysilicon 268 -283 268 -283 0 1
rlabel polysilicon 268 -289 268 -289 0 3
rlabel polysilicon 275 -283 275 -283 0 1
rlabel polysilicon 275 -289 275 -289 0 3
rlabel polysilicon 282 -289 282 -289 0 3
rlabel polysilicon 289 -283 289 -283 0 1
rlabel polysilicon 292 -283 292 -283 0 2
rlabel polysilicon 289 -289 289 -289 0 3
rlabel polysilicon 296 -283 296 -283 0 1
rlabel polysilicon 299 -283 299 -283 0 2
rlabel polysilicon 303 -283 303 -283 0 1
rlabel polysilicon 303 -289 303 -289 0 3
rlabel polysilicon 313 -283 313 -283 0 2
rlabel polysilicon 317 -283 317 -283 0 1
rlabel polysilicon 320 -283 320 -283 0 2
rlabel polysilicon 320 -289 320 -289 0 4
rlabel polysilicon 324 -283 324 -283 0 1
rlabel polysilicon 327 -283 327 -283 0 2
rlabel polysilicon 324 -289 324 -289 0 3
rlabel polysilicon 331 -283 331 -283 0 1
rlabel polysilicon 331 -289 331 -289 0 3
rlabel polysilicon 338 -283 338 -283 0 1
rlabel polysilicon 341 -289 341 -289 0 4
rlabel polysilicon 345 -283 345 -283 0 1
rlabel polysilicon 345 -289 345 -289 0 3
rlabel polysilicon 352 -283 352 -283 0 1
rlabel polysilicon 352 -289 352 -289 0 3
rlabel polysilicon 359 -283 359 -283 0 1
rlabel polysilicon 359 -289 359 -289 0 3
rlabel polysilicon 366 -283 366 -283 0 1
rlabel polysilicon 366 -289 366 -289 0 3
rlabel polysilicon 373 -283 373 -283 0 1
rlabel polysilicon 373 -289 373 -289 0 3
rlabel polysilicon 383 -283 383 -283 0 2
rlabel polysilicon 387 -283 387 -283 0 1
rlabel polysilicon 387 -289 387 -289 0 3
rlabel polysilicon 394 -289 394 -289 0 3
rlabel polysilicon 401 -283 401 -283 0 1
rlabel polysilicon 401 -289 401 -289 0 3
rlabel polysilicon 408 -283 408 -283 0 1
rlabel polysilicon 408 -289 408 -289 0 3
rlabel polysilicon 415 -283 415 -283 0 1
rlabel polysilicon 415 -289 415 -289 0 3
rlabel polysilicon 422 -283 422 -283 0 1
rlabel polysilicon 422 -289 422 -289 0 3
rlabel polysilicon 429 -283 429 -283 0 1
rlabel polysilicon 429 -289 429 -289 0 3
rlabel polysilicon 436 -283 436 -283 0 1
rlabel polysilicon 436 -289 436 -289 0 3
rlabel polysilicon 443 -283 443 -283 0 1
rlabel polysilicon 443 -289 443 -289 0 3
rlabel polysilicon 450 -283 450 -283 0 1
rlabel polysilicon 450 -289 450 -289 0 3
rlabel polysilicon 457 -283 457 -283 0 1
rlabel polysilicon 457 -289 457 -289 0 3
rlabel polysilicon 464 -283 464 -283 0 1
rlabel polysilicon 464 -289 464 -289 0 3
rlabel polysilicon 471 -283 471 -283 0 1
rlabel polysilicon 471 -289 471 -289 0 3
rlabel polysilicon 478 -283 478 -283 0 1
rlabel polysilicon 478 -289 478 -289 0 3
rlabel polysilicon 485 -283 485 -283 0 1
rlabel polysilicon 485 -289 485 -289 0 3
rlabel polysilicon 492 -283 492 -283 0 1
rlabel polysilicon 492 -289 492 -289 0 3
rlabel polysilicon 499 -283 499 -283 0 1
rlabel polysilicon 502 -283 502 -283 0 2
rlabel polysilicon 506 -283 506 -283 0 1
rlabel polysilicon 506 -289 506 -289 0 3
rlabel polysilicon 520 -283 520 -283 0 1
rlabel polysilicon 520 -289 520 -289 0 3
rlabel polysilicon 527 -283 527 -283 0 1
rlabel polysilicon 527 -289 527 -289 0 3
rlabel polysilicon 562 -283 562 -283 0 1
rlabel polysilicon 562 -289 562 -289 0 3
rlabel polysilicon 611 -283 611 -283 0 1
rlabel polysilicon 611 -289 611 -289 0 3
rlabel polysilicon 646 -283 646 -283 0 1
rlabel polysilicon 646 -289 646 -289 0 3
rlabel polysilicon 72 -338 72 -338 0 3
rlabel polysilicon 79 -332 79 -332 0 1
rlabel polysilicon 79 -338 79 -338 0 3
rlabel polysilicon 86 -332 86 -332 0 1
rlabel polysilicon 86 -338 86 -338 0 3
rlabel polysilicon 93 -332 93 -332 0 1
rlabel polysilicon 93 -338 93 -338 0 3
rlabel polysilicon 100 -332 100 -332 0 1
rlabel polysilicon 100 -338 100 -338 0 3
rlabel polysilicon 107 -332 107 -332 0 1
rlabel polysilicon 107 -338 107 -338 0 3
rlabel polysilicon 114 -332 114 -332 0 1
rlabel polysilicon 114 -338 114 -338 0 3
rlabel polysilicon 121 -332 121 -332 0 1
rlabel polysilicon 121 -338 121 -338 0 3
rlabel polysilicon 128 -332 128 -332 0 1
rlabel polysilicon 128 -338 128 -338 0 3
rlabel polysilicon 135 -332 135 -332 0 1
rlabel polysilicon 135 -338 135 -338 0 3
rlabel polysilicon 142 -332 142 -332 0 1
rlabel polysilicon 142 -338 142 -338 0 3
rlabel polysilicon 152 -332 152 -332 0 2
rlabel polysilicon 152 -338 152 -338 0 4
rlabel polysilicon 156 -338 156 -338 0 3
rlabel polysilicon 163 -332 163 -332 0 1
rlabel polysilicon 163 -338 163 -338 0 3
rlabel polysilicon 170 -332 170 -332 0 1
rlabel polysilicon 170 -338 170 -338 0 3
rlabel polysilicon 177 -332 177 -332 0 1
rlabel polysilicon 177 -338 177 -338 0 3
rlabel polysilicon 184 -338 184 -338 0 3
rlabel polysilicon 191 -332 191 -332 0 1
rlabel polysilicon 191 -338 191 -338 0 3
rlabel polysilicon 198 -332 198 -332 0 1
rlabel polysilicon 198 -338 198 -338 0 3
rlabel polysilicon 205 -332 205 -332 0 1
rlabel polysilicon 205 -338 205 -338 0 3
rlabel polysilicon 212 -332 212 -332 0 1
rlabel polysilicon 212 -338 212 -338 0 3
rlabel polysilicon 219 -332 219 -332 0 1
rlabel polysilicon 219 -338 219 -338 0 3
rlabel polysilicon 226 -332 226 -332 0 1
rlabel polysilicon 229 -332 229 -332 0 2
rlabel polysilicon 226 -338 226 -338 0 3
rlabel polysilicon 233 -332 233 -332 0 1
rlabel polysilicon 233 -338 233 -338 0 3
rlabel polysilicon 236 -338 236 -338 0 4
rlabel polysilicon 240 -332 240 -332 0 1
rlabel polysilicon 240 -338 240 -338 0 3
rlabel polysilicon 247 -332 247 -332 0 1
rlabel polysilicon 247 -338 247 -338 0 3
rlabel polysilicon 254 -332 254 -332 0 1
rlabel polysilicon 254 -338 254 -338 0 3
rlabel polysilicon 264 -332 264 -332 0 2
rlabel polysilicon 264 -338 264 -338 0 4
rlabel polysilicon 271 -338 271 -338 0 4
rlabel polysilicon 275 -332 275 -332 0 1
rlabel polysilicon 275 -338 275 -338 0 3
rlabel polysilicon 282 -332 282 -332 0 1
rlabel polysilicon 285 -338 285 -338 0 4
rlabel polysilicon 289 -332 289 -332 0 1
rlabel polysilicon 289 -338 289 -338 0 3
rlabel polysilicon 296 -332 296 -332 0 1
rlabel polysilicon 296 -338 296 -338 0 3
rlabel polysilicon 303 -332 303 -332 0 1
rlabel polysilicon 303 -338 303 -338 0 3
rlabel polysilicon 313 -332 313 -332 0 2
rlabel polysilicon 313 -338 313 -338 0 4
rlabel polysilicon 317 -332 317 -332 0 1
rlabel polysilicon 317 -338 317 -338 0 3
rlabel polysilicon 324 -332 324 -332 0 1
rlabel polysilicon 324 -338 324 -338 0 3
rlabel polysilicon 327 -338 327 -338 0 4
rlabel polysilicon 331 -332 331 -332 0 1
rlabel polysilicon 331 -338 331 -338 0 3
rlabel polysilicon 338 -332 338 -332 0 1
rlabel polysilicon 341 -338 341 -338 0 4
rlabel polysilicon 345 -332 345 -332 0 1
rlabel polysilicon 348 -332 348 -332 0 2
rlabel polysilicon 348 -338 348 -338 0 4
rlabel polysilicon 352 -332 352 -332 0 1
rlabel polysilicon 352 -338 352 -338 0 3
rlabel polysilicon 359 -332 359 -332 0 1
rlabel polysilicon 359 -338 359 -338 0 3
rlabel polysilicon 362 -338 362 -338 0 4
rlabel polysilicon 366 -332 366 -332 0 1
rlabel polysilicon 369 -332 369 -332 0 2
rlabel polysilicon 366 -338 366 -338 0 3
rlabel polysilicon 373 -332 373 -332 0 1
rlabel polysilicon 373 -338 373 -338 0 3
rlabel polysilicon 380 -332 380 -332 0 1
rlabel polysilicon 380 -338 380 -338 0 3
rlabel polysilicon 387 -332 387 -332 0 1
rlabel polysilicon 390 -332 390 -332 0 2
rlabel polysilicon 394 -332 394 -332 0 1
rlabel polysilicon 394 -338 394 -338 0 3
rlabel polysilicon 401 -332 401 -332 0 1
rlabel polysilicon 401 -338 401 -338 0 3
rlabel polysilicon 408 -332 408 -332 0 1
rlabel polysilicon 411 -338 411 -338 0 4
rlabel polysilicon 415 -332 415 -332 0 1
rlabel polysilicon 415 -338 415 -338 0 3
rlabel polysilicon 422 -332 422 -332 0 1
rlabel polysilicon 425 -332 425 -332 0 2
rlabel polysilicon 422 -338 422 -338 0 3
rlabel polysilicon 429 -332 429 -332 0 1
rlabel polysilicon 429 -338 429 -338 0 3
rlabel polysilicon 436 -332 436 -332 0 1
rlabel polysilicon 436 -338 436 -338 0 3
rlabel polysilicon 443 -332 443 -332 0 1
rlabel polysilicon 443 -338 443 -338 0 3
rlabel polysilicon 450 -332 450 -332 0 1
rlabel polysilicon 450 -338 450 -338 0 3
rlabel polysilicon 457 -332 457 -332 0 1
rlabel polysilicon 457 -338 457 -338 0 3
rlabel polysilicon 464 -332 464 -332 0 1
rlabel polysilicon 464 -338 464 -338 0 3
rlabel polysilicon 471 -332 471 -332 0 1
rlabel polysilicon 471 -338 471 -338 0 3
rlabel polysilicon 478 -332 478 -332 0 1
rlabel polysilicon 478 -338 478 -338 0 3
rlabel polysilicon 485 -332 485 -332 0 1
rlabel polysilicon 485 -338 485 -338 0 3
rlabel polysilicon 492 -332 492 -332 0 1
rlabel polysilicon 492 -338 492 -338 0 3
rlabel polysilicon 499 -332 499 -332 0 1
rlabel polysilicon 499 -338 499 -338 0 3
rlabel polysilicon 506 -332 506 -332 0 1
rlabel polysilicon 506 -338 506 -338 0 3
rlabel polysilicon 516 -332 516 -332 0 2
rlabel polysilicon 520 -332 520 -332 0 1
rlabel polysilicon 520 -338 520 -338 0 3
rlabel polysilicon 527 -332 527 -332 0 1
rlabel polysilicon 527 -338 527 -338 0 3
rlabel polysilicon 534 -332 534 -332 0 1
rlabel polysilicon 534 -338 534 -338 0 3
rlabel polysilicon 541 -332 541 -332 0 1
rlabel polysilicon 544 -332 544 -332 0 2
rlabel polysilicon 541 -338 541 -338 0 3
rlabel polysilicon 544 -338 544 -338 0 4
rlabel polysilicon 548 -332 548 -332 0 1
rlabel polysilicon 548 -338 548 -338 0 3
rlabel polysilicon 555 -332 555 -332 0 1
rlabel polysilicon 558 -338 558 -338 0 4
rlabel polysilicon 562 -332 562 -332 0 1
rlabel polysilicon 562 -338 562 -338 0 3
rlabel polysilicon 604 -332 604 -332 0 1
rlabel polysilicon 604 -338 604 -338 0 3
rlabel polysilicon 649 -332 649 -332 0 2
rlabel polysilicon 649 -338 649 -338 0 4
rlabel polysilicon 653 -332 653 -332 0 1
rlabel polysilicon 653 -338 653 -338 0 3
rlabel polysilicon 660 -332 660 -332 0 1
rlabel polysilicon 660 -338 660 -338 0 3
rlabel polysilicon 674 -332 674 -332 0 1
rlabel polysilicon 674 -338 674 -338 0 3
rlabel polysilicon 681 -332 681 -332 0 1
rlabel polysilicon 30 -389 30 -389 0 3
rlabel polysilicon 44 -383 44 -383 0 1
rlabel polysilicon 44 -389 44 -389 0 3
rlabel polysilicon 51 -383 51 -383 0 1
rlabel polysilicon 51 -389 51 -389 0 3
rlabel polysilicon 58 -383 58 -383 0 1
rlabel polysilicon 58 -389 58 -389 0 3
rlabel polysilicon 68 -383 68 -383 0 2
rlabel polysilicon 72 -383 72 -383 0 1
rlabel polysilicon 72 -389 72 -389 0 3
rlabel polysilicon 79 -383 79 -383 0 1
rlabel polysilicon 79 -389 79 -389 0 3
rlabel polysilicon 86 -383 86 -383 0 1
rlabel polysilicon 86 -389 86 -389 0 3
rlabel polysilicon 93 -383 93 -383 0 1
rlabel polysilicon 93 -389 93 -389 0 3
rlabel polysilicon 100 -383 100 -383 0 1
rlabel polysilicon 100 -389 100 -389 0 3
rlabel polysilicon 107 -383 107 -383 0 1
rlabel polysilicon 110 -383 110 -383 0 2
rlabel polysilicon 114 -383 114 -383 0 1
rlabel polysilicon 114 -389 114 -389 0 3
rlabel polysilicon 121 -383 121 -383 0 1
rlabel polysilicon 121 -389 121 -389 0 3
rlabel polysilicon 128 -383 128 -383 0 1
rlabel polysilicon 128 -389 128 -389 0 3
rlabel polysilicon 135 -383 135 -383 0 1
rlabel polysilicon 138 -383 138 -383 0 2
rlabel polysilicon 138 -389 138 -389 0 4
rlabel polysilicon 142 -383 142 -383 0 1
rlabel polysilicon 142 -389 142 -389 0 3
rlabel polysilicon 152 -383 152 -383 0 2
rlabel polysilicon 152 -389 152 -389 0 4
rlabel polysilicon 156 -383 156 -383 0 1
rlabel polysilicon 159 -383 159 -383 0 2
rlabel polysilicon 159 -389 159 -389 0 4
rlabel polysilicon 166 -383 166 -383 0 2
rlabel polysilicon 166 -389 166 -389 0 4
rlabel polysilicon 170 -383 170 -383 0 1
rlabel polysilicon 170 -389 170 -389 0 3
rlabel polysilicon 177 -383 177 -383 0 1
rlabel polysilicon 177 -389 177 -389 0 3
rlabel polysilicon 184 -383 184 -383 0 1
rlabel polysilicon 184 -389 184 -389 0 3
rlabel polysilicon 191 -383 191 -383 0 1
rlabel polysilicon 191 -389 191 -389 0 3
rlabel polysilicon 198 -383 198 -383 0 1
rlabel polysilicon 198 -389 198 -389 0 3
rlabel polysilicon 205 -383 205 -383 0 1
rlabel polysilicon 205 -389 205 -389 0 3
rlabel polysilicon 215 -383 215 -383 0 2
rlabel polysilicon 212 -389 212 -389 0 3
rlabel polysilicon 215 -389 215 -389 0 4
rlabel polysilicon 219 -383 219 -383 0 1
rlabel polysilicon 222 -383 222 -383 0 2
rlabel polysilicon 222 -389 222 -389 0 4
rlabel polysilicon 229 -383 229 -383 0 2
rlabel polysilicon 233 -383 233 -383 0 1
rlabel polysilicon 236 -383 236 -383 0 2
rlabel polysilicon 236 -389 236 -389 0 4
rlabel polysilicon 240 -383 240 -383 0 1
rlabel polysilicon 243 -383 243 -383 0 2
rlabel polysilicon 240 -389 240 -389 0 3
rlabel polysilicon 247 -383 247 -383 0 1
rlabel polysilicon 247 -389 247 -389 0 3
rlabel polysilicon 254 -383 254 -383 0 1
rlabel polysilicon 254 -389 254 -389 0 3
rlabel polysilicon 261 -383 261 -383 0 1
rlabel polysilicon 261 -389 261 -389 0 3
rlabel polysilicon 268 -383 268 -383 0 1
rlabel polysilicon 268 -389 268 -389 0 3
rlabel polysilicon 278 -389 278 -389 0 4
rlabel polysilicon 282 -383 282 -383 0 1
rlabel polysilicon 282 -389 282 -389 0 3
rlabel polysilicon 292 -383 292 -383 0 2
rlabel polysilicon 289 -389 289 -389 0 3
rlabel polysilicon 292 -389 292 -389 0 4
rlabel polysilicon 296 -383 296 -383 0 1
rlabel polysilicon 296 -389 296 -389 0 3
rlabel polysilicon 303 -383 303 -383 0 1
rlabel polysilicon 303 -389 303 -389 0 3
rlabel polysilicon 310 -383 310 -383 0 1
rlabel polysilicon 310 -389 310 -389 0 3
rlabel polysilicon 317 -383 317 -383 0 1
rlabel polysilicon 317 -389 317 -389 0 3
rlabel polysilicon 324 -383 324 -383 0 1
rlabel polysilicon 327 -383 327 -383 0 2
rlabel polysilicon 324 -389 324 -389 0 3
rlabel polysilicon 331 -383 331 -383 0 1
rlabel polysilicon 334 -383 334 -383 0 2
rlabel polysilicon 334 -389 334 -389 0 4
rlabel polysilicon 338 -383 338 -383 0 1
rlabel polysilicon 341 -383 341 -383 0 2
rlabel polysilicon 341 -389 341 -389 0 4
rlabel polysilicon 345 -383 345 -383 0 1
rlabel polysilicon 345 -389 345 -389 0 3
rlabel polysilicon 352 -389 352 -389 0 3
rlabel polysilicon 355 -389 355 -389 0 4
rlabel polysilicon 362 -383 362 -383 0 2
rlabel polysilicon 359 -389 359 -389 0 3
rlabel polysilicon 366 -383 366 -383 0 1
rlabel polysilicon 366 -389 366 -389 0 3
rlabel polysilicon 373 -383 373 -383 0 1
rlabel polysilicon 373 -389 373 -389 0 3
rlabel polysilicon 380 -383 380 -383 0 1
rlabel polysilicon 380 -389 380 -389 0 3
rlabel polysilicon 387 -383 387 -383 0 1
rlabel polysilicon 390 -383 390 -383 0 2
rlabel polysilicon 387 -389 387 -389 0 3
rlabel polysilicon 394 -383 394 -383 0 1
rlabel polysilicon 394 -389 394 -389 0 3
rlabel polysilicon 401 -383 401 -383 0 1
rlabel polysilicon 401 -389 401 -389 0 3
rlabel polysilicon 408 -383 408 -383 0 1
rlabel polysilicon 408 -389 408 -389 0 3
rlabel polysilicon 415 -383 415 -383 0 1
rlabel polysilicon 415 -389 415 -389 0 3
rlabel polysilicon 422 -383 422 -383 0 1
rlabel polysilicon 425 -383 425 -383 0 2
rlabel polysilicon 429 -383 429 -383 0 1
rlabel polysilicon 429 -389 429 -389 0 3
rlabel polysilicon 436 -383 436 -383 0 1
rlabel polysilicon 436 -389 436 -389 0 3
rlabel polysilicon 443 -383 443 -383 0 1
rlabel polysilicon 443 -389 443 -389 0 3
rlabel polysilicon 450 -383 450 -383 0 1
rlabel polysilicon 450 -389 450 -389 0 3
rlabel polysilicon 460 -383 460 -383 0 2
rlabel polysilicon 460 -389 460 -389 0 4
rlabel polysilicon 464 -383 464 -383 0 1
rlabel polysilicon 464 -389 464 -389 0 3
rlabel polysilicon 471 -383 471 -383 0 1
rlabel polysilicon 471 -389 471 -389 0 3
rlabel polysilicon 478 -383 478 -383 0 1
rlabel polysilicon 478 -389 478 -389 0 3
rlabel polysilicon 485 -383 485 -383 0 1
rlabel polysilicon 485 -389 485 -389 0 3
rlabel polysilicon 492 -383 492 -383 0 1
rlabel polysilicon 492 -389 492 -389 0 3
rlabel polysilicon 499 -383 499 -383 0 1
rlabel polysilicon 499 -389 499 -389 0 3
rlabel polysilicon 506 -383 506 -383 0 1
rlabel polysilicon 506 -389 506 -389 0 3
rlabel polysilicon 513 -383 513 -383 0 1
rlabel polysilicon 513 -389 513 -389 0 3
rlabel polysilicon 523 -383 523 -383 0 2
rlabel polysilicon 527 -383 527 -383 0 1
rlabel polysilicon 527 -389 527 -389 0 3
rlabel polysilicon 534 -383 534 -383 0 1
rlabel polysilicon 534 -389 534 -389 0 3
rlabel polysilicon 541 -383 541 -383 0 1
rlabel polysilicon 541 -389 541 -389 0 3
rlabel polysilicon 548 -383 548 -383 0 1
rlabel polysilicon 548 -389 548 -389 0 3
rlabel polysilicon 555 -383 555 -383 0 1
rlabel polysilicon 555 -389 555 -389 0 3
rlabel polysilicon 562 -383 562 -383 0 1
rlabel polysilicon 569 -383 569 -383 0 1
rlabel polysilicon 569 -389 569 -389 0 3
rlabel polysilicon 576 -383 576 -383 0 1
rlabel polysilicon 576 -389 576 -389 0 3
rlabel polysilicon 583 -383 583 -383 0 1
rlabel polysilicon 583 -389 583 -389 0 3
rlabel polysilicon 590 -383 590 -383 0 1
rlabel polysilicon 590 -389 590 -389 0 3
rlabel polysilicon 597 -383 597 -383 0 1
rlabel polysilicon 597 -389 597 -389 0 3
rlabel polysilicon 604 -383 604 -383 0 1
rlabel polysilicon 604 -389 604 -389 0 3
rlabel polysilicon 611 -383 611 -383 0 1
rlabel polysilicon 611 -389 611 -389 0 3
rlabel polysilicon 618 -383 618 -383 0 1
rlabel polysilicon 618 -389 618 -389 0 3
rlabel polysilicon 625 -383 625 -383 0 1
rlabel polysilicon 625 -389 625 -389 0 3
rlabel polysilicon 632 -383 632 -383 0 1
rlabel polysilicon 632 -389 632 -389 0 3
rlabel polysilicon 639 -383 639 -383 0 1
rlabel polysilicon 642 -383 642 -383 0 2
rlabel polysilicon 646 -383 646 -383 0 1
rlabel polysilicon 646 -389 646 -389 0 3
rlabel polysilicon 653 -383 653 -383 0 1
rlabel polysilicon 653 -389 653 -389 0 3
rlabel polysilicon 660 -383 660 -383 0 1
rlabel polysilicon 667 -383 667 -383 0 1
rlabel polysilicon 667 -389 667 -389 0 3
rlabel polysilicon 674 -389 674 -389 0 3
rlabel polysilicon 681 -383 681 -383 0 1
rlabel polysilicon 681 -389 681 -389 0 3
rlabel polysilicon 688 -383 688 -383 0 1
rlabel polysilicon 688 -389 688 -389 0 3
rlabel polysilicon 2 -440 2 -440 0 1
rlabel polysilicon 2 -446 2 -446 0 3
rlabel polysilicon 9 -446 9 -446 0 3
rlabel polysilicon 16 -440 16 -440 0 1
rlabel polysilicon 16 -446 16 -446 0 3
rlabel polysilicon 23 -440 23 -440 0 1
rlabel polysilicon 23 -446 23 -446 0 3
rlabel polysilicon 33 -446 33 -446 0 4
rlabel polysilicon 37 -440 37 -440 0 1
rlabel polysilicon 37 -446 37 -446 0 3
rlabel polysilicon 44 -440 44 -440 0 1
rlabel polysilicon 44 -446 44 -446 0 3
rlabel polysilicon 51 -440 51 -440 0 1
rlabel polysilicon 51 -446 51 -446 0 3
rlabel polysilicon 58 -440 58 -440 0 1
rlabel polysilicon 58 -446 58 -446 0 3
rlabel polysilicon 65 -440 65 -440 0 1
rlabel polysilicon 65 -446 65 -446 0 3
rlabel polysilicon 72 -440 72 -440 0 1
rlabel polysilicon 72 -446 72 -446 0 3
rlabel polysilicon 79 -440 79 -440 0 1
rlabel polysilicon 79 -446 79 -446 0 3
rlabel polysilicon 86 -440 86 -440 0 1
rlabel polysilicon 86 -446 86 -446 0 3
rlabel polysilicon 93 -440 93 -440 0 1
rlabel polysilicon 93 -446 93 -446 0 3
rlabel polysilicon 100 -440 100 -440 0 1
rlabel polysilicon 100 -446 100 -446 0 3
rlabel polysilicon 107 -440 107 -440 0 1
rlabel polysilicon 107 -446 107 -446 0 3
rlabel polysilicon 114 -440 114 -440 0 1
rlabel polysilicon 114 -446 114 -446 0 3
rlabel polysilicon 121 -440 121 -440 0 1
rlabel polysilicon 121 -446 121 -446 0 3
rlabel polysilicon 128 -440 128 -440 0 1
rlabel polysilicon 128 -446 128 -446 0 3
rlabel polysilicon 135 -440 135 -440 0 1
rlabel polysilicon 138 -446 138 -446 0 4
rlabel polysilicon 145 -440 145 -440 0 2
rlabel polysilicon 142 -446 142 -446 0 3
rlabel polysilicon 145 -446 145 -446 0 4
rlabel polysilicon 149 -440 149 -440 0 1
rlabel polysilicon 149 -446 149 -446 0 3
rlabel polysilicon 159 -440 159 -440 0 2
rlabel polysilicon 159 -446 159 -446 0 4
rlabel polysilicon 163 -440 163 -440 0 1
rlabel polysilicon 163 -446 163 -446 0 3
rlabel polysilicon 170 -440 170 -440 0 1
rlabel polysilicon 170 -446 170 -446 0 3
rlabel polysilicon 177 -440 177 -440 0 1
rlabel polysilicon 180 -440 180 -440 0 2
rlabel polysilicon 177 -446 177 -446 0 3
rlabel polysilicon 180 -446 180 -446 0 4
rlabel polysilicon 184 -440 184 -440 0 1
rlabel polysilicon 187 -440 187 -440 0 2
rlabel polysilicon 184 -446 184 -446 0 3
rlabel polysilicon 187 -446 187 -446 0 4
rlabel polysilicon 191 -440 191 -440 0 1
rlabel polysilicon 191 -446 191 -446 0 3
rlabel polysilicon 198 -440 198 -440 0 1
rlabel polysilicon 198 -446 198 -446 0 3
rlabel polysilicon 205 -440 205 -440 0 1
rlabel polysilicon 205 -446 205 -446 0 3
rlabel polysilicon 215 -440 215 -440 0 2
rlabel polysilicon 215 -446 215 -446 0 4
rlabel polysilicon 219 -440 219 -440 0 1
rlabel polysilicon 219 -446 219 -446 0 3
rlabel polysilicon 226 -440 226 -440 0 1
rlabel polysilicon 226 -446 226 -446 0 3
rlabel polysilicon 233 -440 233 -440 0 1
rlabel polysilicon 236 -440 236 -440 0 2
rlabel polysilicon 233 -446 233 -446 0 3
rlabel polysilicon 236 -446 236 -446 0 4
rlabel polysilicon 240 -440 240 -440 0 1
rlabel polysilicon 243 -446 243 -446 0 4
rlabel polysilicon 247 -440 247 -440 0 1
rlabel polysilicon 247 -446 247 -446 0 3
rlabel polysilicon 254 -440 254 -440 0 1
rlabel polysilicon 254 -446 254 -446 0 3
rlabel polysilicon 261 -440 261 -440 0 1
rlabel polysilicon 261 -446 261 -446 0 3
rlabel polysilicon 268 -440 268 -440 0 1
rlabel polysilicon 268 -446 268 -446 0 3
rlabel polysilicon 275 -440 275 -440 0 1
rlabel polysilicon 275 -446 275 -446 0 3
rlabel polysilicon 282 -440 282 -440 0 1
rlabel polysilicon 285 -440 285 -440 0 2
rlabel polysilicon 282 -446 282 -446 0 3
rlabel polysilicon 285 -446 285 -446 0 4
rlabel polysilicon 289 -440 289 -440 0 1
rlabel polysilicon 289 -446 289 -446 0 3
rlabel polysilicon 292 -446 292 -446 0 4
rlabel polysilicon 296 -440 296 -440 0 1
rlabel polysilicon 296 -446 296 -446 0 3
rlabel polysilicon 303 -440 303 -440 0 1
rlabel polysilicon 310 -440 310 -440 0 1
rlabel polysilicon 310 -446 310 -446 0 3
rlabel polysilicon 317 -440 317 -440 0 1
rlabel polysilicon 317 -446 317 -446 0 3
rlabel polysilicon 324 -440 324 -440 0 1
rlabel polysilicon 327 -440 327 -440 0 2
rlabel polysilicon 331 -440 331 -440 0 1
rlabel polysilicon 331 -446 331 -446 0 3
rlabel polysilicon 338 -440 338 -440 0 1
rlabel polysilicon 341 -440 341 -440 0 2
rlabel polysilicon 345 -440 345 -440 0 1
rlabel polysilicon 345 -446 345 -446 0 3
rlabel polysilicon 352 -440 352 -440 0 1
rlabel polysilicon 352 -446 352 -446 0 3
rlabel polysilicon 359 -440 359 -440 0 1
rlabel polysilicon 359 -446 359 -446 0 3
rlabel polysilicon 369 -440 369 -440 0 2
rlabel polysilicon 366 -446 366 -446 0 3
rlabel polysilicon 369 -446 369 -446 0 4
rlabel polysilicon 373 -440 373 -440 0 1
rlabel polysilicon 376 -440 376 -440 0 2
rlabel polysilicon 373 -446 373 -446 0 3
rlabel polysilicon 376 -446 376 -446 0 4
rlabel polysilicon 380 -440 380 -440 0 1
rlabel polysilicon 380 -446 380 -446 0 3
rlabel polysilicon 387 -440 387 -440 0 1
rlabel polysilicon 387 -446 387 -446 0 3
rlabel polysilicon 397 -440 397 -440 0 2
rlabel polysilicon 397 -446 397 -446 0 4
rlabel polysilicon 401 -440 401 -440 0 1
rlabel polysilicon 404 -440 404 -440 0 2
rlabel polysilicon 404 -446 404 -446 0 4
rlabel polysilicon 408 -440 408 -440 0 1
rlabel polysilicon 415 -440 415 -440 0 1
rlabel polysilicon 415 -446 415 -446 0 3
rlabel polysilicon 422 -440 422 -440 0 1
rlabel polysilicon 422 -446 422 -446 0 3
rlabel polysilicon 429 -440 429 -440 0 1
rlabel polysilicon 429 -446 429 -446 0 3
rlabel polysilicon 436 -440 436 -440 0 1
rlabel polysilicon 439 -440 439 -440 0 2
rlabel polysilicon 436 -446 436 -446 0 3
rlabel polysilicon 443 -440 443 -440 0 1
rlabel polysilicon 443 -446 443 -446 0 3
rlabel polysilicon 450 -440 450 -440 0 1
rlabel polysilicon 450 -446 450 -446 0 3
rlabel polysilicon 457 -440 457 -440 0 1
rlabel polysilicon 457 -446 457 -446 0 3
rlabel polysilicon 467 -440 467 -440 0 2
rlabel polysilicon 464 -446 464 -446 0 3
rlabel polysilicon 471 -440 471 -440 0 1
rlabel polysilicon 471 -446 471 -446 0 3
rlabel polysilicon 478 -440 478 -440 0 1
rlabel polysilicon 478 -446 478 -446 0 3
rlabel polysilicon 485 -440 485 -440 0 1
rlabel polysilicon 485 -446 485 -446 0 3
rlabel polysilicon 492 -440 492 -440 0 1
rlabel polysilicon 492 -446 492 -446 0 3
rlabel polysilicon 499 -440 499 -440 0 1
rlabel polysilicon 499 -446 499 -446 0 3
rlabel polysilicon 509 -446 509 -446 0 4
rlabel polysilicon 513 -440 513 -440 0 1
rlabel polysilicon 513 -446 513 -446 0 3
rlabel polysilicon 520 -440 520 -440 0 1
rlabel polysilicon 520 -446 520 -446 0 3
rlabel polysilicon 527 -440 527 -440 0 1
rlabel polysilicon 527 -446 527 -446 0 3
rlabel polysilicon 534 -440 534 -440 0 1
rlabel polysilicon 534 -446 534 -446 0 3
rlabel polysilicon 541 -440 541 -440 0 1
rlabel polysilicon 541 -446 541 -446 0 3
rlabel polysilicon 548 -440 548 -440 0 1
rlabel polysilicon 548 -446 548 -446 0 3
rlabel polysilicon 558 -440 558 -440 0 2
rlabel polysilicon 558 -446 558 -446 0 4
rlabel polysilicon 562 -440 562 -440 0 1
rlabel polysilicon 562 -446 562 -446 0 3
rlabel polysilicon 569 -440 569 -440 0 1
rlabel polysilicon 569 -446 569 -446 0 3
rlabel polysilicon 576 -440 576 -440 0 1
rlabel polysilicon 576 -446 576 -446 0 3
rlabel polysilicon 583 -440 583 -440 0 1
rlabel polysilicon 583 -446 583 -446 0 3
rlabel polysilicon 590 -440 590 -440 0 1
rlabel polysilicon 590 -446 590 -446 0 3
rlabel polysilicon 597 -440 597 -440 0 1
rlabel polysilicon 597 -446 597 -446 0 3
rlabel polysilicon 604 -440 604 -440 0 1
rlabel polysilicon 604 -446 604 -446 0 3
rlabel polysilicon 611 -440 611 -440 0 1
rlabel polysilicon 611 -446 611 -446 0 3
rlabel polysilicon 618 -440 618 -440 0 1
rlabel polysilicon 618 -446 618 -446 0 3
rlabel polysilicon 625 -440 625 -440 0 1
rlabel polysilicon 628 -440 628 -440 0 2
rlabel polysilicon 625 -446 625 -446 0 3
rlabel polysilicon 632 -440 632 -440 0 1
rlabel polysilicon 632 -446 632 -446 0 3
rlabel polysilicon 635 -446 635 -446 0 4
rlabel polysilicon 639 -440 639 -440 0 1
rlabel polysilicon 639 -446 639 -446 0 3
rlabel polysilicon 649 -440 649 -440 0 2
rlabel polysilicon 646 -446 646 -446 0 3
rlabel polysilicon 653 -440 653 -440 0 1
rlabel polysilicon 653 -446 653 -446 0 3
rlabel polysilicon 663 -440 663 -440 0 2
rlabel polysilicon 663 -446 663 -446 0 4
rlabel polysilicon 667 -440 667 -440 0 1
rlabel polysilicon 667 -446 667 -446 0 3
rlabel polysilicon 9 -497 9 -497 0 1
rlabel polysilicon 9 -503 9 -503 0 3
rlabel polysilicon 16 -497 16 -497 0 1
rlabel polysilicon 16 -503 16 -503 0 3
rlabel polysilicon 23 -497 23 -497 0 1
rlabel polysilicon 23 -503 23 -503 0 3
rlabel polysilicon 30 -497 30 -497 0 1
rlabel polysilicon 30 -503 30 -503 0 3
rlabel polysilicon 37 -497 37 -497 0 1
rlabel polysilicon 37 -503 37 -503 0 3
rlabel polysilicon 44 -497 44 -497 0 1
rlabel polysilicon 44 -503 44 -503 0 3
rlabel polysilicon 51 -497 51 -497 0 1
rlabel polysilicon 51 -503 51 -503 0 3
rlabel polysilicon 58 -497 58 -497 0 1
rlabel polysilicon 65 -497 65 -497 0 1
rlabel polysilicon 68 -503 68 -503 0 4
rlabel polysilicon 72 -497 72 -497 0 1
rlabel polysilicon 72 -503 72 -503 0 3
rlabel polysilicon 79 -497 79 -497 0 1
rlabel polysilicon 79 -503 79 -503 0 3
rlabel polysilicon 86 -497 86 -497 0 1
rlabel polysilicon 86 -503 86 -503 0 3
rlabel polysilicon 93 -503 93 -503 0 3
rlabel polysilicon 100 -497 100 -497 0 1
rlabel polysilicon 100 -503 100 -503 0 3
rlabel polysilicon 107 -497 107 -497 0 1
rlabel polysilicon 110 -497 110 -497 0 2
rlabel polysilicon 107 -503 107 -503 0 3
rlabel polysilicon 114 -497 114 -497 0 1
rlabel polysilicon 121 -497 121 -497 0 1
rlabel polysilicon 121 -503 121 -503 0 3
rlabel polysilicon 128 -497 128 -497 0 1
rlabel polysilicon 131 -497 131 -497 0 2
rlabel polysilicon 138 -497 138 -497 0 2
rlabel polysilicon 135 -503 135 -503 0 3
rlabel polysilicon 142 -497 142 -497 0 1
rlabel polysilicon 142 -503 142 -503 0 3
rlabel polysilicon 149 -503 149 -503 0 3
rlabel polysilicon 152 -503 152 -503 0 4
rlabel polysilicon 156 -497 156 -497 0 1
rlabel polysilicon 156 -503 156 -503 0 3
rlabel polysilicon 159 -503 159 -503 0 4
rlabel polysilicon 163 -497 163 -497 0 1
rlabel polysilicon 166 -497 166 -497 0 2
rlabel polysilicon 163 -503 163 -503 0 3
rlabel polysilicon 170 -497 170 -497 0 1
rlabel polysilicon 170 -503 170 -503 0 3
rlabel polysilicon 177 -497 177 -497 0 1
rlabel polysilicon 177 -503 177 -503 0 3
rlabel polysilicon 184 -497 184 -497 0 1
rlabel polysilicon 184 -503 184 -503 0 3
rlabel polysilicon 191 -497 191 -497 0 1
rlabel polysilicon 191 -503 191 -503 0 3
rlabel polysilicon 201 -497 201 -497 0 2
rlabel polysilicon 198 -503 198 -503 0 3
rlabel polysilicon 208 -497 208 -497 0 2
rlabel polysilicon 205 -503 205 -503 0 3
rlabel polysilicon 208 -503 208 -503 0 4
rlabel polysilicon 212 -497 212 -497 0 1
rlabel polysilicon 215 -497 215 -497 0 2
rlabel polysilicon 212 -503 212 -503 0 3
rlabel polysilicon 215 -503 215 -503 0 4
rlabel polysilicon 219 -497 219 -497 0 1
rlabel polysilicon 219 -503 219 -503 0 3
rlabel polysilicon 226 -497 226 -497 0 1
rlabel polysilicon 226 -503 226 -503 0 3
rlabel polysilicon 233 -497 233 -497 0 1
rlabel polysilicon 233 -503 233 -503 0 3
rlabel polysilicon 243 -497 243 -497 0 2
rlabel polysilicon 240 -503 240 -503 0 3
rlabel polysilicon 243 -503 243 -503 0 4
rlabel polysilicon 247 -497 247 -497 0 1
rlabel polysilicon 247 -503 247 -503 0 3
rlabel polysilicon 254 -497 254 -497 0 1
rlabel polysilicon 254 -503 254 -503 0 3
rlabel polysilicon 264 -497 264 -497 0 2
rlabel polysilicon 271 -503 271 -503 0 4
rlabel polysilicon 275 -497 275 -497 0 1
rlabel polysilicon 275 -503 275 -503 0 3
rlabel polysilicon 282 -497 282 -497 0 1
rlabel polysilicon 282 -503 282 -503 0 3
rlabel polysilicon 289 -497 289 -497 0 1
rlabel polysilicon 289 -503 289 -503 0 3
rlabel polysilicon 296 -497 296 -497 0 1
rlabel polysilicon 296 -503 296 -503 0 3
rlabel polysilicon 303 -497 303 -497 0 1
rlabel polysilicon 303 -503 303 -503 0 3
rlabel polysilicon 310 -497 310 -497 0 1
rlabel polysilicon 310 -503 310 -503 0 3
rlabel polysilicon 317 -497 317 -497 0 1
rlabel polysilicon 317 -503 317 -503 0 3
rlabel polysilicon 324 -497 324 -497 0 1
rlabel polysilicon 324 -503 324 -503 0 3
rlabel polysilicon 331 -503 331 -503 0 3
rlabel polysilicon 338 -497 338 -497 0 1
rlabel polysilicon 338 -503 338 -503 0 3
rlabel polysilicon 345 -497 345 -497 0 1
rlabel polysilicon 345 -503 345 -503 0 3
rlabel polysilicon 352 -497 352 -497 0 1
rlabel polysilicon 355 -497 355 -497 0 2
rlabel polysilicon 355 -503 355 -503 0 4
rlabel polysilicon 359 -497 359 -497 0 1
rlabel polysilicon 359 -503 359 -503 0 3
rlabel polysilicon 366 -497 366 -497 0 1
rlabel polysilicon 369 -503 369 -503 0 4
rlabel polysilicon 373 -497 373 -497 0 1
rlabel polysilicon 373 -503 373 -503 0 3
rlabel polysilicon 380 -497 380 -497 0 1
rlabel polysilicon 383 -503 383 -503 0 4
rlabel polysilicon 387 -497 387 -497 0 1
rlabel polysilicon 390 -497 390 -497 0 2
rlabel polysilicon 390 -503 390 -503 0 4
rlabel polysilicon 397 -497 397 -497 0 2
rlabel polysilicon 394 -503 394 -503 0 3
rlabel polysilicon 397 -503 397 -503 0 4
rlabel polysilicon 401 -497 401 -497 0 1
rlabel polysilicon 401 -503 401 -503 0 3
rlabel polysilicon 408 -497 408 -497 0 1
rlabel polysilicon 408 -503 408 -503 0 3
rlabel polysilicon 415 -497 415 -497 0 1
rlabel polysilicon 418 -497 418 -497 0 2
rlabel polysilicon 415 -503 415 -503 0 3
rlabel polysilicon 422 -497 422 -497 0 1
rlabel polysilicon 422 -503 422 -503 0 3
rlabel polysilicon 429 -497 429 -497 0 1
rlabel polysilicon 429 -503 429 -503 0 3
rlabel polysilicon 436 -497 436 -497 0 1
rlabel polysilicon 436 -503 436 -503 0 3
rlabel polysilicon 443 -497 443 -497 0 1
rlabel polysilicon 443 -503 443 -503 0 3
rlabel polysilicon 450 -497 450 -497 0 1
rlabel polysilicon 450 -503 450 -503 0 3
rlabel polysilicon 457 -497 457 -497 0 1
rlabel polysilicon 457 -503 457 -503 0 3
rlabel polysilicon 464 -497 464 -497 0 1
rlabel polysilicon 464 -503 464 -503 0 3
rlabel polysilicon 471 -497 471 -497 0 1
rlabel polysilicon 471 -503 471 -503 0 3
rlabel polysilicon 478 -503 478 -503 0 3
rlabel polysilicon 485 -497 485 -497 0 1
rlabel polysilicon 485 -503 485 -503 0 3
rlabel polysilicon 492 -497 492 -497 0 1
rlabel polysilicon 492 -503 492 -503 0 3
rlabel polysilicon 499 -497 499 -497 0 1
rlabel polysilicon 499 -503 499 -503 0 3
rlabel polysilicon 509 -497 509 -497 0 2
rlabel polysilicon 513 -497 513 -497 0 1
rlabel polysilicon 513 -503 513 -503 0 3
rlabel polysilicon 520 -497 520 -497 0 1
rlabel polysilicon 520 -503 520 -503 0 3
rlabel polysilicon 527 -497 527 -497 0 1
rlabel polysilicon 527 -503 527 -503 0 3
rlabel polysilicon 534 -497 534 -497 0 1
rlabel polysilicon 534 -503 534 -503 0 3
rlabel polysilicon 541 -497 541 -497 0 1
rlabel polysilicon 541 -503 541 -503 0 3
rlabel polysilicon 548 -497 548 -497 0 1
rlabel polysilicon 548 -503 548 -503 0 3
rlabel polysilicon 555 -497 555 -497 0 1
rlabel polysilicon 555 -503 555 -503 0 3
rlabel polysilicon 562 -497 562 -497 0 1
rlabel polysilicon 562 -503 562 -503 0 3
rlabel polysilicon 569 -497 569 -497 0 1
rlabel polysilicon 569 -503 569 -503 0 3
rlabel polysilicon 576 -497 576 -497 0 1
rlabel polysilicon 576 -503 576 -503 0 3
rlabel polysilicon 583 -497 583 -497 0 1
rlabel polysilicon 583 -503 583 -503 0 3
rlabel polysilicon 590 -503 590 -503 0 3
rlabel polysilicon 597 -497 597 -497 0 1
rlabel polysilicon 597 -503 597 -503 0 3
rlabel polysilicon 604 -503 604 -503 0 3
rlabel polysilicon 614 -497 614 -497 0 2
rlabel polysilicon 611 -503 611 -503 0 3
rlabel polysilicon 614 -503 614 -503 0 4
rlabel polysilicon 618 -497 618 -497 0 1
rlabel polysilicon 618 -503 618 -503 0 3
rlabel polysilicon 625 -503 625 -503 0 3
rlabel polysilicon 628 -503 628 -503 0 4
rlabel polysilicon 632 -497 632 -497 0 1
rlabel polysilicon 632 -503 632 -503 0 3
rlabel polysilicon 639 -497 639 -497 0 1
rlabel polysilicon 639 -503 639 -503 0 3
rlabel polysilicon 646 -497 646 -497 0 1
rlabel polysilicon 646 -503 646 -503 0 3
rlabel polysilicon 653 -497 653 -497 0 1
rlabel polysilicon 653 -503 653 -503 0 3
rlabel polysilicon 660 -497 660 -497 0 1
rlabel polysilicon 660 -503 660 -503 0 3
rlabel polysilicon 670 -503 670 -503 0 4
rlabel polysilicon 5 -554 5 -554 0 2
rlabel polysilicon 9 -554 9 -554 0 1
rlabel polysilicon 9 -560 9 -560 0 3
rlabel polysilicon 16 -554 16 -554 0 1
rlabel polysilicon 16 -560 16 -560 0 3
rlabel polysilicon 23 -554 23 -554 0 1
rlabel polysilicon 23 -560 23 -560 0 3
rlabel polysilicon 30 -554 30 -554 0 1
rlabel polysilicon 30 -560 30 -560 0 3
rlabel polysilicon 37 -554 37 -554 0 1
rlabel polysilicon 37 -560 37 -560 0 3
rlabel polysilicon 44 -554 44 -554 0 1
rlabel polysilicon 44 -560 44 -560 0 3
rlabel polysilicon 51 -554 51 -554 0 1
rlabel polysilicon 51 -560 51 -560 0 3
rlabel polysilicon 58 -554 58 -554 0 1
rlabel polysilicon 61 -554 61 -554 0 2
rlabel polysilicon 65 -554 65 -554 0 1
rlabel polysilicon 65 -560 65 -560 0 3
rlabel polysilicon 72 -554 72 -554 0 1
rlabel polysilicon 72 -560 72 -560 0 3
rlabel polysilicon 75 -560 75 -560 0 4
rlabel polysilicon 82 -554 82 -554 0 2
rlabel polysilicon 82 -560 82 -560 0 4
rlabel polysilicon 86 -554 86 -554 0 1
rlabel polysilicon 93 -554 93 -554 0 1
rlabel polysilicon 93 -560 93 -560 0 3
rlabel polysilicon 100 -554 100 -554 0 1
rlabel polysilicon 100 -560 100 -560 0 3
rlabel polysilicon 107 -554 107 -554 0 1
rlabel polysilicon 107 -560 107 -560 0 3
rlabel polysilicon 114 -554 114 -554 0 1
rlabel polysilicon 117 -554 117 -554 0 2
rlabel polysilicon 114 -560 114 -560 0 3
rlabel polysilicon 117 -560 117 -560 0 4
rlabel polysilicon 121 -554 121 -554 0 1
rlabel polysilicon 121 -560 121 -560 0 3
rlabel polysilicon 128 -554 128 -554 0 1
rlabel polysilicon 131 -554 131 -554 0 2
rlabel polysilicon 128 -560 128 -560 0 3
rlabel polysilicon 131 -560 131 -560 0 4
rlabel polysilicon 135 -554 135 -554 0 1
rlabel polysilicon 135 -560 135 -560 0 3
rlabel polysilicon 142 -560 142 -560 0 3
rlabel polysilicon 149 -554 149 -554 0 1
rlabel polysilicon 149 -560 149 -560 0 3
rlabel polysilicon 156 -554 156 -554 0 1
rlabel polysilicon 156 -560 156 -560 0 3
rlabel polysilicon 163 -554 163 -554 0 1
rlabel polysilicon 163 -560 163 -560 0 3
rlabel polysilicon 170 -554 170 -554 0 1
rlabel polysilicon 170 -560 170 -560 0 3
rlabel polysilicon 180 -554 180 -554 0 2
rlabel polysilicon 177 -560 177 -560 0 3
rlabel polysilicon 180 -560 180 -560 0 4
rlabel polysilicon 184 -554 184 -554 0 1
rlabel polysilicon 184 -560 184 -560 0 3
rlabel polysilicon 194 -560 194 -560 0 4
rlabel polysilicon 198 -554 198 -554 0 1
rlabel polysilicon 198 -560 198 -560 0 3
rlabel polysilicon 205 -554 205 -554 0 1
rlabel polysilicon 208 -554 208 -554 0 2
rlabel polysilicon 205 -560 205 -560 0 3
rlabel polysilicon 212 -554 212 -554 0 1
rlabel polysilicon 212 -560 212 -560 0 3
rlabel polysilicon 219 -554 219 -554 0 1
rlabel polysilicon 219 -560 219 -560 0 3
rlabel polysilicon 226 -554 226 -554 0 1
rlabel polysilicon 226 -560 226 -560 0 3
rlabel polysilicon 233 -554 233 -554 0 1
rlabel polysilicon 233 -560 233 -560 0 3
rlabel polysilicon 240 -554 240 -554 0 1
rlabel polysilicon 243 -554 243 -554 0 2
rlabel polysilicon 243 -560 243 -560 0 4
rlabel polysilicon 247 -554 247 -554 0 1
rlabel polysilicon 247 -560 247 -560 0 3
rlabel polysilicon 254 -554 254 -554 0 1
rlabel polysilicon 254 -560 254 -560 0 3
rlabel polysilicon 261 -554 261 -554 0 1
rlabel polysilicon 261 -560 261 -560 0 3
rlabel polysilicon 268 -554 268 -554 0 1
rlabel polysilicon 268 -560 268 -560 0 3
rlabel polysilicon 275 -554 275 -554 0 1
rlabel polysilicon 278 -554 278 -554 0 2
rlabel polysilicon 278 -560 278 -560 0 4
rlabel polysilicon 285 -554 285 -554 0 2
rlabel polysilicon 282 -560 282 -560 0 3
rlabel polysilicon 285 -560 285 -560 0 4
rlabel polysilicon 292 -554 292 -554 0 2
rlabel polysilicon 289 -560 289 -560 0 3
rlabel polysilicon 292 -560 292 -560 0 4
rlabel polysilicon 296 -554 296 -554 0 1
rlabel polysilicon 296 -560 296 -560 0 3
rlabel polysilicon 303 -554 303 -554 0 1
rlabel polysilicon 303 -560 303 -560 0 3
rlabel polysilicon 310 -554 310 -554 0 1
rlabel polysilicon 313 -554 313 -554 0 2
rlabel polysilicon 310 -560 310 -560 0 3
rlabel polysilicon 313 -560 313 -560 0 4
rlabel polysilicon 317 -554 317 -554 0 1
rlabel polysilicon 317 -560 317 -560 0 3
rlabel polysilicon 320 -560 320 -560 0 4
rlabel polysilicon 324 -554 324 -554 0 1
rlabel polysilicon 324 -560 324 -560 0 3
rlabel polysilicon 331 -554 331 -554 0 1
rlabel polysilicon 331 -560 331 -560 0 3
rlabel polysilicon 341 -554 341 -554 0 2
rlabel polysilicon 341 -560 341 -560 0 4
rlabel polysilicon 345 -554 345 -554 0 1
rlabel polysilicon 348 -554 348 -554 0 2
rlabel polysilicon 345 -560 345 -560 0 3
rlabel polysilicon 355 -554 355 -554 0 2
rlabel polysilicon 352 -560 352 -560 0 3
rlabel polysilicon 355 -560 355 -560 0 4
rlabel polysilicon 362 -554 362 -554 0 2
rlabel polysilicon 359 -560 359 -560 0 3
rlabel polysilicon 366 -554 366 -554 0 1
rlabel polysilicon 366 -560 366 -560 0 3
rlabel polysilicon 376 -554 376 -554 0 2
rlabel polysilicon 373 -560 373 -560 0 3
rlabel polysilicon 376 -560 376 -560 0 4
rlabel polysilicon 380 -554 380 -554 0 1
rlabel polysilicon 380 -560 380 -560 0 3
rlabel polysilicon 387 -554 387 -554 0 1
rlabel polysilicon 387 -560 387 -560 0 3
rlabel polysilicon 394 -554 394 -554 0 1
rlabel polysilicon 394 -560 394 -560 0 3
rlabel polysilicon 401 -554 401 -554 0 1
rlabel polysilicon 401 -560 401 -560 0 3
rlabel polysilicon 404 -560 404 -560 0 4
rlabel polysilicon 408 -554 408 -554 0 1
rlabel polysilicon 408 -560 408 -560 0 3
rlabel polysilicon 415 -554 415 -554 0 1
rlabel polysilicon 415 -560 415 -560 0 3
rlabel polysilicon 425 -560 425 -560 0 4
rlabel polysilicon 429 -554 429 -554 0 1
rlabel polysilicon 429 -560 429 -560 0 3
rlabel polysilicon 436 -554 436 -554 0 1
rlabel polysilicon 436 -560 436 -560 0 3
rlabel polysilicon 443 -554 443 -554 0 1
rlabel polysilicon 443 -560 443 -560 0 3
rlabel polysilicon 450 -554 450 -554 0 1
rlabel polysilicon 450 -560 450 -560 0 3
rlabel polysilicon 457 -560 457 -560 0 3
rlabel polysilicon 460 -560 460 -560 0 4
rlabel polysilicon 464 -554 464 -554 0 1
rlabel polysilicon 464 -560 464 -560 0 3
rlabel polysilicon 471 -554 471 -554 0 1
rlabel polysilicon 471 -560 471 -560 0 3
rlabel polysilicon 478 -554 478 -554 0 1
rlabel polysilicon 478 -560 478 -560 0 3
rlabel polysilicon 485 -554 485 -554 0 1
rlabel polysilicon 485 -560 485 -560 0 3
rlabel polysilicon 492 -554 492 -554 0 1
rlabel polysilicon 492 -560 492 -560 0 3
rlabel polysilicon 499 -554 499 -554 0 1
rlabel polysilicon 502 -554 502 -554 0 2
rlabel polysilicon 506 -554 506 -554 0 1
rlabel polysilicon 506 -560 506 -560 0 3
rlabel polysilicon 513 -554 513 -554 0 1
rlabel polysilicon 513 -560 513 -560 0 3
rlabel polysilicon 520 -554 520 -554 0 1
rlabel polysilicon 520 -560 520 -560 0 3
rlabel polysilicon 527 -554 527 -554 0 1
rlabel polysilicon 527 -560 527 -560 0 3
rlabel polysilicon 534 -554 534 -554 0 1
rlabel polysilicon 534 -560 534 -560 0 3
rlabel polysilicon 541 -554 541 -554 0 1
rlabel polysilicon 541 -560 541 -560 0 3
rlabel polysilicon 548 -554 548 -554 0 1
rlabel polysilicon 548 -560 548 -560 0 3
rlabel polysilicon 555 -554 555 -554 0 1
rlabel polysilicon 555 -560 555 -560 0 3
rlabel polysilicon 562 -554 562 -554 0 1
rlabel polysilicon 562 -560 562 -560 0 3
rlabel polysilicon 569 -554 569 -554 0 1
rlabel polysilicon 569 -560 569 -560 0 3
rlabel polysilicon 576 -554 576 -554 0 1
rlabel polysilicon 576 -560 576 -560 0 3
rlabel polysilicon 583 -554 583 -554 0 1
rlabel polysilicon 583 -560 583 -560 0 3
rlabel polysilicon 590 -554 590 -554 0 1
rlabel polysilicon 590 -560 590 -560 0 3
rlabel polysilicon 597 -554 597 -554 0 1
rlabel polysilicon 597 -560 597 -560 0 3
rlabel polysilicon 604 -554 604 -554 0 1
rlabel polysilicon 604 -560 604 -560 0 3
rlabel polysilicon 611 -554 611 -554 0 1
rlabel polysilicon 611 -560 611 -560 0 3
rlabel polysilicon 618 -554 618 -554 0 1
rlabel polysilicon 618 -560 618 -560 0 3
rlabel polysilicon 628 -554 628 -554 0 2
rlabel polysilicon 625 -560 625 -560 0 3
rlabel polysilicon 632 -554 632 -554 0 1
rlabel polysilicon 632 -560 632 -560 0 3
rlabel polysilicon 639 -554 639 -554 0 1
rlabel polysilicon 639 -560 639 -560 0 3
rlabel polysilicon 646 -554 646 -554 0 1
rlabel polysilicon 646 -560 646 -560 0 3
rlabel polysilicon 653 -554 653 -554 0 1
rlabel polysilicon 653 -560 653 -560 0 3
rlabel polysilicon 656 -560 656 -560 0 4
rlabel polysilicon 660 -554 660 -554 0 1
rlabel polysilicon 660 -560 660 -560 0 3
rlabel polysilicon 667 -554 667 -554 0 1
rlabel polysilicon 667 -560 667 -560 0 3
rlabel polysilicon 670 -560 670 -560 0 4
rlabel polysilicon 674 -554 674 -554 0 1
rlabel polysilicon 674 -560 674 -560 0 3
rlabel polysilicon 681 -554 681 -554 0 1
rlabel polysilicon 684 -560 684 -560 0 4
rlabel polysilicon 688 -554 688 -554 0 1
rlabel polysilicon 688 -560 688 -560 0 3
rlabel polysilicon 2 -611 2 -611 0 1
rlabel polysilicon 2 -617 2 -617 0 3
rlabel polysilicon 9 -611 9 -611 0 1
rlabel polysilicon 9 -617 9 -617 0 3
rlabel polysilicon 19 -611 19 -611 0 2
rlabel polysilicon 23 -611 23 -611 0 1
rlabel polysilicon 23 -617 23 -617 0 3
rlabel polysilicon 30 -611 30 -611 0 1
rlabel polysilicon 30 -617 30 -617 0 3
rlabel polysilicon 40 -611 40 -611 0 2
rlabel polysilicon 44 -617 44 -617 0 3
rlabel polysilicon 51 -611 51 -611 0 1
rlabel polysilicon 51 -617 51 -617 0 3
rlabel polysilicon 58 -611 58 -611 0 1
rlabel polysilicon 58 -617 58 -617 0 3
rlabel polysilicon 65 -611 65 -611 0 1
rlabel polysilicon 65 -617 65 -617 0 3
rlabel polysilicon 75 -617 75 -617 0 4
rlabel polysilicon 79 -611 79 -611 0 1
rlabel polysilicon 79 -617 79 -617 0 3
rlabel polysilicon 86 -617 86 -617 0 3
rlabel polysilicon 93 -611 93 -611 0 1
rlabel polysilicon 96 -611 96 -611 0 2
rlabel polysilicon 93 -617 93 -617 0 3
rlabel polysilicon 100 -611 100 -611 0 1
rlabel polysilicon 103 -611 103 -611 0 2
rlabel polysilicon 100 -617 100 -617 0 3
rlabel polysilicon 107 -611 107 -611 0 1
rlabel polysilicon 107 -617 107 -617 0 3
rlabel polysilicon 114 -611 114 -611 0 1
rlabel polysilicon 114 -617 114 -617 0 3
rlabel polysilicon 117 -617 117 -617 0 4
rlabel polysilicon 121 -611 121 -611 0 1
rlabel polysilicon 121 -617 121 -617 0 3
rlabel polysilicon 128 -611 128 -611 0 1
rlabel polysilicon 131 -611 131 -611 0 2
rlabel polysilicon 128 -617 128 -617 0 3
rlabel polysilicon 135 -611 135 -611 0 1
rlabel polysilicon 135 -617 135 -617 0 3
rlabel polysilicon 142 -611 142 -611 0 1
rlabel polysilicon 142 -617 142 -617 0 3
rlabel polysilicon 149 -611 149 -611 0 1
rlabel polysilicon 149 -617 149 -617 0 3
rlabel polysilicon 156 -617 156 -617 0 3
rlabel polysilicon 159 -617 159 -617 0 4
rlabel polysilicon 163 -611 163 -611 0 1
rlabel polysilicon 163 -617 163 -617 0 3
rlabel polysilicon 166 -617 166 -617 0 4
rlabel polysilicon 170 -611 170 -611 0 1
rlabel polysilicon 173 -617 173 -617 0 4
rlabel polysilicon 177 -611 177 -611 0 1
rlabel polysilicon 180 -611 180 -611 0 2
rlabel polysilicon 177 -617 177 -617 0 3
rlabel polysilicon 184 -611 184 -611 0 1
rlabel polysilicon 187 -611 187 -611 0 2
rlabel polysilicon 187 -617 187 -617 0 4
rlabel polysilicon 191 -611 191 -611 0 1
rlabel polysilicon 191 -617 191 -617 0 3
rlabel polysilicon 198 -611 198 -611 0 1
rlabel polysilicon 198 -617 198 -617 0 3
rlabel polysilicon 205 -611 205 -611 0 1
rlabel polysilicon 205 -617 205 -617 0 3
rlabel polysilicon 212 -611 212 -611 0 1
rlabel polysilicon 212 -617 212 -617 0 3
rlabel polysilicon 219 -611 219 -611 0 1
rlabel polysilicon 219 -617 219 -617 0 3
rlabel polysilicon 226 -611 226 -611 0 1
rlabel polysilicon 226 -617 226 -617 0 3
rlabel polysilicon 233 -611 233 -611 0 1
rlabel polysilicon 236 -611 236 -611 0 2
rlabel polysilicon 243 -611 243 -611 0 2
rlabel polysilicon 240 -617 240 -617 0 3
rlabel polysilicon 243 -617 243 -617 0 4
rlabel polysilicon 247 -611 247 -611 0 1
rlabel polysilicon 247 -617 247 -617 0 3
rlabel polysilicon 254 -611 254 -611 0 1
rlabel polysilicon 254 -617 254 -617 0 3
rlabel polysilicon 264 -611 264 -611 0 2
rlabel polysilicon 268 -611 268 -611 0 1
rlabel polysilicon 268 -617 268 -617 0 3
rlabel polysilicon 275 -611 275 -611 0 1
rlabel polysilicon 278 -617 278 -617 0 4
rlabel polysilicon 282 -611 282 -611 0 1
rlabel polysilicon 282 -617 282 -617 0 3
rlabel polysilicon 289 -611 289 -611 0 1
rlabel polysilicon 289 -617 289 -617 0 3
rlabel polysilicon 296 -611 296 -611 0 1
rlabel polysilicon 296 -617 296 -617 0 3
rlabel polysilicon 303 -611 303 -611 0 1
rlabel polysilicon 306 -611 306 -611 0 2
rlabel polysilicon 310 -611 310 -611 0 1
rlabel polysilicon 310 -617 310 -617 0 3
rlabel polysilicon 317 -611 317 -611 0 1
rlabel polysilicon 317 -617 317 -617 0 3
rlabel polysilicon 324 -611 324 -611 0 1
rlabel polysilicon 324 -617 324 -617 0 3
rlabel polysilicon 331 -611 331 -611 0 1
rlabel polysilicon 331 -617 331 -617 0 3
rlabel polysilicon 338 -611 338 -611 0 1
rlabel polysilicon 338 -617 338 -617 0 3
rlabel polysilicon 345 -611 345 -611 0 1
rlabel polysilicon 345 -617 345 -617 0 3
rlabel polysilicon 355 -617 355 -617 0 4
rlabel polysilicon 359 -611 359 -611 0 1
rlabel polysilicon 359 -617 359 -617 0 3
rlabel polysilicon 366 -611 366 -611 0 1
rlabel polysilicon 369 -611 369 -611 0 2
rlabel polysilicon 366 -617 366 -617 0 3
rlabel polysilicon 369 -617 369 -617 0 4
rlabel polysilicon 373 -611 373 -611 0 1
rlabel polysilicon 373 -617 373 -617 0 3
rlabel polysilicon 380 -611 380 -611 0 1
rlabel polysilicon 383 -611 383 -611 0 2
rlabel polysilicon 380 -617 380 -617 0 3
rlabel polysilicon 383 -617 383 -617 0 4
rlabel polysilicon 387 -611 387 -611 0 1
rlabel polysilicon 387 -617 387 -617 0 3
rlabel polysilicon 390 -617 390 -617 0 4
rlabel polysilicon 397 -611 397 -611 0 2
rlabel polysilicon 394 -617 394 -617 0 3
rlabel polysilicon 401 -611 401 -611 0 1
rlabel polysilicon 401 -617 401 -617 0 3
rlabel polysilicon 408 -611 408 -611 0 1
rlabel polysilicon 408 -617 408 -617 0 3
rlabel polysilicon 415 -611 415 -611 0 1
rlabel polysilicon 415 -617 415 -617 0 3
rlabel polysilicon 422 -611 422 -611 0 1
rlabel polysilicon 422 -617 422 -617 0 3
rlabel polysilicon 429 -611 429 -611 0 1
rlabel polysilicon 429 -617 429 -617 0 3
rlabel polysilicon 436 -611 436 -611 0 1
rlabel polysilicon 436 -617 436 -617 0 3
rlabel polysilicon 443 -611 443 -611 0 1
rlabel polysilicon 443 -617 443 -617 0 3
rlabel polysilicon 450 -611 450 -611 0 1
rlabel polysilicon 453 -617 453 -617 0 4
rlabel polysilicon 457 -611 457 -611 0 1
rlabel polysilicon 457 -617 457 -617 0 3
rlabel polysilicon 464 -611 464 -611 0 1
rlabel polysilicon 467 -611 467 -611 0 2
rlabel polysilicon 464 -617 464 -617 0 3
rlabel polysilicon 471 -611 471 -611 0 1
rlabel polysilicon 474 -611 474 -611 0 2
rlabel polysilicon 474 -617 474 -617 0 4
rlabel polysilicon 478 -611 478 -611 0 1
rlabel polysilicon 478 -617 478 -617 0 3
rlabel polysilicon 485 -611 485 -611 0 1
rlabel polysilicon 485 -617 485 -617 0 3
rlabel polysilicon 492 -617 492 -617 0 3
rlabel polysilicon 495 -617 495 -617 0 4
rlabel polysilicon 499 -611 499 -611 0 1
rlabel polysilicon 499 -617 499 -617 0 3
rlabel polysilicon 506 -611 506 -611 0 1
rlabel polysilicon 506 -617 506 -617 0 3
rlabel polysilicon 513 -611 513 -611 0 1
rlabel polysilicon 513 -617 513 -617 0 3
rlabel polysilicon 520 -611 520 -611 0 1
rlabel polysilicon 520 -617 520 -617 0 3
rlabel polysilicon 527 -611 527 -611 0 1
rlabel polysilicon 527 -617 527 -617 0 3
rlabel polysilicon 534 -611 534 -611 0 1
rlabel polysilicon 534 -617 534 -617 0 3
rlabel polysilicon 541 -611 541 -611 0 1
rlabel polysilicon 541 -617 541 -617 0 3
rlabel polysilicon 548 -611 548 -611 0 1
rlabel polysilicon 548 -617 548 -617 0 3
rlabel polysilicon 555 -611 555 -611 0 1
rlabel polysilicon 555 -617 555 -617 0 3
rlabel polysilicon 562 -611 562 -611 0 1
rlabel polysilicon 562 -617 562 -617 0 3
rlabel polysilicon 569 -611 569 -611 0 1
rlabel polysilicon 569 -617 569 -617 0 3
rlabel polysilicon 576 -611 576 -611 0 1
rlabel polysilicon 576 -617 576 -617 0 3
rlabel polysilicon 583 -611 583 -611 0 1
rlabel polysilicon 583 -617 583 -617 0 3
rlabel polysilicon 590 -611 590 -611 0 1
rlabel polysilicon 590 -617 590 -617 0 3
rlabel polysilicon 597 -611 597 -611 0 1
rlabel polysilicon 597 -617 597 -617 0 3
rlabel polysilicon 604 -611 604 -611 0 1
rlabel polysilicon 611 -611 611 -611 0 1
rlabel polysilicon 611 -617 611 -617 0 3
rlabel polysilicon 618 -611 618 -611 0 1
rlabel polysilicon 618 -617 618 -617 0 3
rlabel polysilicon 625 -611 625 -611 0 1
rlabel polysilicon 625 -617 625 -617 0 3
rlabel polysilicon 632 -611 632 -611 0 1
rlabel polysilicon 632 -617 632 -617 0 3
rlabel polysilicon 639 -611 639 -611 0 1
rlabel polysilicon 639 -617 639 -617 0 3
rlabel polysilicon 646 -611 646 -611 0 1
rlabel polysilicon 646 -617 646 -617 0 3
rlabel polysilicon 653 -611 653 -611 0 1
rlabel polysilicon 656 -611 656 -611 0 2
rlabel polysilicon 653 -617 653 -617 0 3
rlabel polysilicon 660 -611 660 -611 0 1
rlabel polysilicon 660 -617 660 -617 0 3
rlabel polysilicon 677 -611 677 -611 0 2
rlabel polysilicon 688 -611 688 -611 0 1
rlabel polysilicon 2 -684 2 -684 0 1
rlabel polysilicon 2 -690 2 -690 0 3
rlabel polysilicon 9 -684 9 -684 0 1
rlabel polysilicon 9 -690 9 -690 0 3
rlabel polysilicon 16 -684 16 -684 0 1
rlabel polysilicon 19 -690 19 -690 0 4
rlabel polysilicon 23 -684 23 -684 0 1
rlabel polysilicon 23 -690 23 -690 0 3
rlabel polysilicon 30 -684 30 -684 0 1
rlabel polysilicon 30 -690 30 -690 0 3
rlabel polysilicon 37 -684 37 -684 0 1
rlabel polysilicon 37 -690 37 -690 0 3
rlabel polysilicon 44 -684 44 -684 0 1
rlabel polysilicon 44 -690 44 -690 0 3
rlabel polysilicon 54 -684 54 -684 0 2
rlabel polysilicon 61 -684 61 -684 0 2
rlabel polysilicon 65 -684 65 -684 0 1
rlabel polysilicon 65 -690 65 -690 0 3
rlabel polysilicon 72 -684 72 -684 0 1
rlabel polysilicon 72 -690 72 -690 0 3
rlabel polysilicon 79 -684 79 -684 0 1
rlabel polysilicon 82 -690 82 -690 0 4
rlabel polysilicon 89 -684 89 -684 0 2
rlabel polysilicon 89 -690 89 -690 0 4
rlabel polysilicon 93 -684 93 -684 0 1
rlabel polysilicon 96 -684 96 -684 0 2
rlabel polysilicon 93 -690 93 -690 0 3
rlabel polysilicon 100 -690 100 -690 0 3
rlabel polysilicon 103 -690 103 -690 0 4
rlabel polysilicon 107 -684 107 -684 0 1
rlabel polysilicon 107 -690 107 -690 0 3
rlabel polysilicon 114 -684 114 -684 0 1
rlabel polysilicon 114 -690 114 -690 0 3
rlabel polysilicon 121 -684 121 -684 0 1
rlabel polysilicon 121 -690 121 -690 0 3
rlabel polysilicon 128 -684 128 -684 0 1
rlabel polysilicon 128 -690 128 -690 0 3
rlabel polysilicon 135 -684 135 -684 0 1
rlabel polysilicon 138 -690 138 -690 0 4
rlabel polysilicon 142 -684 142 -684 0 1
rlabel polysilicon 145 -684 145 -684 0 2
rlabel polysilicon 142 -690 142 -690 0 3
rlabel polysilicon 149 -684 149 -684 0 1
rlabel polysilicon 149 -690 149 -690 0 3
rlabel polysilicon 156 -684 156 -684 0 1
rlabel polysilicon 156 -690 156 -690 0 3
rlabel polysilicon 163 -684 163 -684 0 1
rlabel polysilicon 166 -684 166 -684 0 2
rlabel polysilicon 166 -690 166 -690 0 4
rlabel polysilicon 170 -684 170 -684 0 1
rlabel polysilicon 170 -690 170 -690 0 3
rlabel polysilicon 177 -684 177 -684 0 1
rlabel polysilicon 177 -690 177 -690 0 3
rlabel polysilicon 184 -684 184 -684 0 1
rlabel polysilicon 184 -690 184 -690 0 3
rlabel polysilicon 187 -690 187 -690 0 4
rlabel polysilicon 191 -684 191 -684 0 1
rlabel polysilicon 194 -684 194 -684 0 2
rlabel polysilicon 191 -690 191 -690 0 3
rlabel polysilicon 198 -684 198 -684 0 1
rlabel polysilicon 198 -690 198 -690 0 3
rlabel polysilicon 205 -684 205 -684 0 1
rlabel polysilicon 205 -690 205 -690 0 3
rlabel polysilicon 212 -684 212 -684 0 1
rlabel polysilicon 212 -690 212 -690 0 3
rlabel polysilicon 215 -690 215 -690 0 4
rlabel polysilicon 219 -684 219 -684 0 1
rlabel polysilicon 219 -690 219 -690 0 3
rlabel polysilicon 229 -684 229 -684 0 2
rlabel polysilicon 226 -690 226 -690 0 3
rlabel polysilicon 233 -684 233 -684 0 1
rlabel polysilicon 233 -690 233 -690 0 3
rlabel polysilicon 236 -690 236 -690 0 4
rlabel polysilicon 240 -684 240 -684 0 1
rlabel polysilicon 243 -684 243 -684 0 2
rlabel polysilicon 240 -690 240 -690 0 3
rlabel polysilicon 243 -690 243 -690 0 4
rlabel polysilicon 247 -684 247 -684 0 1
rlabel polysilicon 247 -690 247 -690 0 3
rlabel polysilicon 254 -684 254 -684 0 1
rlabel polysilicon 254 -690 254 -690 0 3
rlabel polysilicon 261 -684 261 -684 0 1
rlabel polysilicon 261 -690 261 -690 0 3
rlabel polysilicon 268 -684 268 -684 0 1
rlabel polysilicon 268 -690 268 -690 0 3
rlabel polysilicon 278 -684 278 -684 0 2
rlabel polysilicon 278 -690 278 -690 0 4
rlabel polysilicon 282 -684 282 -684 0 1
rlabel polysilicon 285 -684 285 -684 0 2
rlabel polysilicon 289 -684 289 -684 0 1
rlabel polysilicon 289 -690 289 -690 0 3
rlabel polysilicon 299 -684 299 -684 0 2
rlabel polysilicon 296 -690 296 -690 0 3
rlabel polysilicon 299 -690 299 -690 0 4
rlabel polysilicon 303 -684 303 -684 0 1
rlabel polysilicon 303 -690 303 -690 0 3
rlabel polysilicon 310 -684 310 -684 0 1
rlabel polysilicon 310 -690 310 -690 0 3
rlabel polysilicon 317 -684 317 -684 0 1
rlabel polysilicon 317 -690 317 -690 0 3
rlabel polysilicon 324 -684 324 -684 0 1
rlabel polysilicon 324 -690 324 -690 0 3
rlabel polysilicon 331 -684 331 -684 0 1
rlabel polysilicon 331 -690 331 -690 0 3
rlabel polysilicon 338 -684 338 -684 0 1
rlabel polysilicon 338 -690 338 -690 0 3
rlabel polysilicon 345 -684 345 -684 0 1
rlabel polysilicon 348 -684 348 -684 0 2
rlabel polysilicon 345 -690 345 -690 0 3
rlabel polysilicon 348 -690 348 -690 0 4
rlabel polysilicon 352 -684 352 -684 0 1
rlabel polysilicon 352 -690 352 -690 0 3
rlabel polysilicon 359 -690 359 -690 0 3
rlabel polysilicon 362 -690 362 -690 0 4
rlabel polysilicon 366 -684 366 -684 0 1
rlabel polysilicon 369 -684 369 -684 0 2
rlabel polysilicon 366 -690 366 -690 0 3
rlabel polysilicon 369 -690 369 -690 0 4
rlabel polysilicon 376 -684 376 -684 0 2
rlabel polysilicon 373 -690 373 -690 0 3
rlabel polysilicon 376 -690 376 -690 0 4
rlabel polysilicon 380 -684 380 -684 0 1
rlabel polysilicon 380 -690 380 -690 0 3
rlabel polysilicon 387 -684 387 -684 0 1
rlabel polysilicon 387 -690 387 -690 0 3
rlabel polysilicon 394 -684 394 -684 0 1
rlabel polysilicon 394 -690 394 -690 0 3
rlabel polysilicon 401 -684 401 -684 0 1
rlabel polysilicon 401 -690 401 -690 0 3
rlabel polysilicon 411 -684 411 -684 0 2
rlabel polysilicon 408 -690 408 -690 0 3
rlabel polysilicon 411 -690 411 -690 0 4
rlabel polysilicon 415 -684 415 -684 0 1
rlabel polysilicon 415 -690 415 -690 0 3
rlabel polysilicon 422 -684 422 -684 0 1
rlabel polysilicon 425 -684 425 -684 0 2
rlabel polysilicon 422 -690 422 -690 0 3
rlabel polysilicon 429 -684 429 -684 0 1
rlabel polysilicon 429 -690 429 -690 0 3
rlabel polysilicon 436 -684 436 -684 0 1
rlabel polysilicon 436 -690 436 -690 0 3
rlabel polysilicon 443 -684 443 -684 0 1
rlabel polysilicon 443 -690 443 -690 0 3
rlabel polysilicon 453 -684 453 -684 0 2
rlabel polysilicon 450 -690 450 -690 0 3
rlabel polysilicon 453 -690 453 -690 0 4
rlabel polysilicon 457 -684 457 -684 0 1
rlabel polysilicon 457 -690 457 -690 0 3
rlabel polysilicon 460 -690 460 -690 0 4
rlabel polysilicon 464 -684 464 -684 0 1
rlabel polysilicon 464 -690 464 -690 0 3
rlabel polysilicon 467 -690 467 -690 0 4
rlabel polysilicon 471 -684 471 -684 0 1
rlabel polysilicon 471 -690 471 -690 0 3
rlabel polysilicon 478 -684 478 -684 0 1
rlabel polysilicon 478 -690 478 -690 0 3
rlabel polysilicon 485 -684 485 -684 0 1
rlabel polysilicon 485 -690 485 -690 0 3
rlabel polysilicon 492 -684 492 -684 0 1
rlabel polysilicon 492 -690 492 -690 0 3
rlabel polysilicon 499 -684 499 -684 0 1
rlabel polysilicon 499 -690 499 -690 0 3
rlabel polysilicon 506 -684 506 -684 0 1
rlabel polysilicon 506 -690 506 -690 0 3
rlabel polysilicon 513 -684 513 -684 0 1
rlabel polysilicon 513 -690 513 -690 0 3
rlabel polysilicon 520 -684 520 -684 0 1
rlabel polysilicon 520 -690 520 -690 0 3
rlabel polysilicon 527 -684 527 -684 0 1
rlabel polysilicon 527 -690 527 -690 0 3
rlabel polysilicon 534 -684 534 -684 0 1
rlabel polysilicon 534 -690 534 -690 0 3
rlabel polysilicon 541 -684 541 -684 0 1
rlabel polysilicon 541 -690 541 -690 0 3
rlabel polysilicon 548 -684 548 -684 0 1
rlabel polysilicon 548 -690 548 -690 0 3
rlabel polysilicon 555 -684 555 -684 0 1
rlabel polysilicon 555 -690 555 -690 0 3
rlabel polysilicon 562 -684 562 -684 0 1
rlabel polysilicon 562 -690 562 -690 0 3
rlabel polysilicon 569 -684 569 -684 0 1
rlabel polysilicon 569 -690 569 -690 0 3
rlabel polysilicon 576 -684 576 -684 0 1
rlabel polysilicon 576 -690 576 -690 0 3
rlabel polysilicon 583 -684 583 -684 0 1
rlabel polysilicon 583 -690 583 -690 0 3
rlabel polysilicon 590 -684 590 -684 0 1
rlabel polysilicon 590 -690 590 -690 0 3
rlabel polysilicon 597 -684 597 -684 0 1
rlabel polysilicon 597 -690 597 -690 0 3
rlabel polysilicon 604 -684 604 -684 0 1
rlabel polysilicon 604 -690 604 -690 0 3
rlabel polysilicon 611 -684 611 -684 0 1
rlabel polysilicon 611 -690 611 -690 0 3
rlabel polysilicon 618 -684 618 -684 0 1
rlabel polysilicon 618 -690 618 -690 0 3
rlabel polysilicon 625 -684 625 -684 0 1
rlabel polysilicon 625 -690 625 -690 0 3
rlabel polysilicon 632 -684 632 -684 0 1
rlabel polysilicon 632 -690 632 -690 0 3
rlabel polysilicon 639 -684 639 -684 0 1
rlabel polysilicon 639 -690 639 -690 0 3
rlabel polysilicon 646 -684 646 -684 0 1
rlabel polysilicon 646 -690 646 -690 0 3
rlabel polysilicon 653 -684 653 -684 0 1
rlabel polysilicon 653 -690 653 -690 0 3
rlabel polysilicon 660 -684 660 -684 0 1
rlabel polysilicon 660 -690 660 -690 0 3
rlabel polysilicon 667 -684 667 -684 0 1
rlabel polysilicon 667 -690 667 -690 0 3
rlabel polysilicon 677 -684 677 -684 0 2
rlabel polysilicon 674 -690 674 -690 0 3
rlabel polysilicon 681 -684 681 -684 0 1
rlabel polysilicon 688 -684 688 -684 0 1
rlabel polysilicon 688 -690 688 -690 0 3
rlabel polysilicon 695 -684 695 -684 0 1
rlabel polysilicon 695 -690 695 -690 0 3
rlabel polysilicon 702 -684 702 -684 0 1
rlabel polysilicon 702 -690 702 -690 0 3
rlabel polysilicon 716 -684 716 -684 0 1
rlabel polysilicon 719 -684 719 -684 0 2
rlabel polysilicon 730 -684 730 -684 0 1
rlabel polysilicon 730 -690 730 -690 0 3
rlabel polysilicon 2 -751 2 -751 0 1
rlabel polysilicon 2 -757 2 -757 0 3
rlabel polysilicon 9 -751 9 -751 0 1
rlabel polysilicon 9 -757 9 -757 0 3
rlabel polysilicon 16 -751 16 -751 0 1
rlabel polysilicon 16 -757 16 -757 0 3
rlabel polysilicon 23 -751 23 -751 0 1
rlabel polysilicon 23 -757 23 -757 0 3
rlabel polysilicon 30 -751 30 -751 0 1
rlabel polysilicon 30 -757 30 -757 0 3
rlabel polysilicon 40 -751 40 -751 0 2
rlabel polysilicon 44 -751 44 -751 0 1
rlabel polysilicon 44 -757 44 -757 0 3
rlabel polysilicon 51 -751 51 -751 0 1
rlabel polysilicon 51 -757 51 -757 0 3
rlabel polysilicon 58 -751 58 -751 0 1
rlabel polysilicon 58 -757 58 -757 0 3
rlabel polysilicon 65 -751 65 -751 0 1
rlabel polysilicon 65 -757 65 -757 0 3
rlabel polysilicon 72 -751 72 -751 0 1
rlabel polysilicon 72 -757 72 -757 0 3
rlabel polysilicon 79 -751 79 -751 0 1
rlabel polysilicon 79 -757 79 -757 0 3
rlabel polysilicon 89 -751 89 -751 0 2
rlabel polysilicon 86 -757 86 -757 0 3
rlabel polysilicon 89 -757 89 -757 0 4
rlabel polysilicon 93 -751 93 -751 0 1
rlabel polysilicon 93 -757 93 -757 0 3
rlabel polysilicon 100 -751 100 -751 0 1
rlabel polysilicon 100 -757 100 -757 0 3
rlabel polysilicon 103 -757 103 -757 0 4
rlabel polysilicon 107 -751 107 -751 0 1
rlabel polysilicon 107 -757 107 -757 0 3
rlabel polysilicon 114 -751 114 -751 0 1
rlabel polysilicon 114 -757 114 -757 0 3
rlabel polysilicon 124 -751 124 -751 0 2
rlabel polysilicon 121 -757 121 -757 0 3
rlabel polysilicon 124 -757 124 -757 0 4
rlabel polysilicon 128 -751 128 -751 0 1
rlabel polysilicon 128 -757 128 -757 0 3
rlabel polysilicon 135 -751 135 -751 0 1
rlabel polysilicon 135 -757 135 -757 0 3
rlabel polysilicon 142 -751 142 -751 0 1
rlabel polysilicon 142 -757 142 -757 0 3
rlabel polysilicon 149 -751 149 -751 0 1
rlabel polysilicon 149 -757 149 -757 0 3
rlabel polysilicon 156 -751 156 -751 0 1
rlabel polysilicon 156 -757 156 -757 0 3
rlabel polysilicon 163 -751 163 -751 0 1
rlabel polysilicon 163 -757 163 -757 0 3
rlabel polysilicon 170 -751 170 -751 0 1
rlabel polysilicon 170 -757 170 -757 0 3
rlabel polysilicon 177 -751 177 -751 0 1
rlabel polysilicon 177 -757 177 -757 0 3
rlabel polysilicon 184 -751 184 -751 0 1
rlabel polysilicon 184 -757 184 -757 0 3
rlabel polysilicon 191 -751 191 -751 0 1
rlabel polysilicon 191 -757 191 -757 0 3
rlabel polysilicon 198 -751 198 -751 0 1
rlabel polysilicon 201 -751 201 -751 0 2
rlabel polysilicon 198 -757 198 -757 0 3
rlabel polysilicon 205 -751 205 -751 0 1
rlabel polysilicon 205 -757 205 -757 0 3
rlabel polysilicon 212 -751 212 -751 0 1
rlabel polysilicon 212 -757 212 -757 0 3
rlabel polysilicon 219 -751 219 -751 0 1
rlabel polysilicon 219 -757 219 -757 0 3
rlabel polysilicon 226 -751 226 -751 0 1
rlabel polysilicon 226 -757 226 -757 0 3
rlabel polysilicon 229 -757 229 -757 0 4
rlabel polysilicon 233 -757 233 -757 0 3
rlabel polysilicon 236 -757 236 -757 0 4
rlabel polysilicon 240 -751 240 -751 0 1
rlabel polysilicon 240 -757 240 -757 0 3
rlabel polysilicon 247 -751 247 -751 0 1
rlabel polysilicon 247 -757 247 -757 0 3
rlabel polysilicon 250 -757 250 -757 0 4
rlabel polysilicon 254 -751 254 -751 0 1
rlabel polysilicon 254 -757 254 -757 0 3
rlabel polysilicon 261 -751 261 -751 0 1
rlabel polysilicon 261 -757 261 -757 0 3
rlabel polysilicon 268 -751 268 -751 0 1
rlabel polysilicon 268 -757 268 -757 0 3
rlabel polysilicon 278 -751 278 -751 0 2
rlabel polysilicon 282 -751 282 -751 0 1
rlabel polysilicon 292 -751 292 -751 0 2
rlabel polysilicon 296 -751 296 -751 0 1
rlabel polysilicon 296 -757 296 -757 0 3
rlabel polysilicon 303 -751 303 -751 0 1
rlabel polysilicon 303 -757 303 -757 0 3
rlabel polysilicon 310 -751 310 -751 0 1
rlabel polysilicon 310 -757 310 -757 0 3
rlabel polysilicon 317 -751 317 -751 0 1
rlabel polysilicon 317 -757 317 -757 0 3
rlabel polysilicon 324 -751 324 -751 0 1
rlabel polysilicon 327 -751 327 -751 0 2
rlabel polysilicon 327 -757 327 -757 0 4
rlabel polysilicon 331 -751 331 -751 0 1
rlabel polysilicon 331 -757 331 -757 0 3
rlabel polysilicon 341 -751 341 -751 0 2
rlabel polysilicon 338 -757 338 -757 0 3
rlabel polysilicon 341 -757 341 -757 0 4
rlabel polysilicon 345 -751 345 -751 0 1
rlabel polysilicon 345 -757 345 -757 0 3
rlabel polysilicon 352 -751 352 -751 0 1
rlabel polysilicon 352 -757 352 -757 0 3
rlabel polysilicon 362 -751 362 -751 0 2
rlabel polysilicon 359 -757 359 -757 0 3
rlabel polysilicon 362 -757 362 -757 0 4
rlabel polysilicon 366 -751 366 -751 0 1
rlabel polysilicon 366 -757 366 -757 0 3
rlabel polysilicon 373 -751 373 -751 0 1
rlabel polysilicon 373 -757 373 -757 0 3
rlabel polysilicon 380 -751 380 -751 0 1
rlabel polysilicon 380 -757 380 -757 0 3
rlabel polysilicon 383 -757 383 -757 0 4
rlabel polysilicon 387 -751 387 -751 0 1
rlabel polysilicon 387 -757 387 -757 0 3
rlabel polysilicon 390 -757 390 -757 0 4
rlabel polysilicon 397 -757 397 -757 0 4
rlabel polysilicon 401 -751 401 -751 0 1
rlabel polysilicon 401 -757 401 -757 0 3
rlabel polysilicon 408 -751 408 -751 0 1
rlabel polysilicon 408 -757 408 -757 0 3
rlabel polysilicon 411 -757 411 -757 0 4
rlabel polysilicon 415 -751 415 -751 0 1
rlabel polysilicon 415 -757 415 -757 0 3
rlabel polysilicon 422 -751 422 -751 0 1
rlabel polysilicon 422 -757 422 -757 0 3
rlabel polysilicon 429 -751 429 -751 0 1
rlabel polysilicon 432 -751 432 -751 0 2
rlabel polysilicon 436 -751 436 -751 0 1
rlabel polysilicon 436 -757 436 -757 0 3
rlabel polysilicon 443 -751 443 -751 0 1
rlabel polysilicon 443 -757 443 -757 0 3
rlabel polysilicon 450 -751 450 -751 0 1
rlabel polysilicon 453 -751 453 -751 0 2
rlabel polysilicon 450 -757 450 -757 0 3
rlabel polysilicon 453 -757 453 -757 0 4
rlabel polysilicon 457 -751 457 -751 0 1
rlabel polysilicon 457 -757 457 -757 0 3
rlabel polysilicon 464 -751 464 -751 0 1
rlabel polysilicon 464 -757 464 -757 0 3
rlabel polysilicon 471 -751 471 -751 0 1
rlabel polysilicon 471 -757 471 -757 0 3
rlabel polysilicon 478 -751 478 -751 0 1
rlabel polysilicon 478 -757 478 -757 0 3
rlabel polysilicon 485 -751 485 -751 0 1
rlabel polysilicon 492 -751 492 -751 0 1
rlabel polysilicon 492 -757 492 -757 0 3
rlabel polysilicon 495 -757 495 -757 0 4
rlabel polysilicon 499 -751 499 -751 0 1
rlabel polysilicon 499 -757 499 -757 0 3
rlabel polysilicon 506 -751 506 -751 0 1
rlabel polysilicon 506 -757 506 -757 0 3
rlabel polysilicon 513 -751 513 -751 0 1
rlabel polysilicon 513 -757 513 -757 0 3
rlabel polysilicon 520 -751 520 -751 0 1
rlabel polysilicon 520 -757 520 -757 0 3
rlabel polysilicon 527 -757 527 -757 0 3
rlabel polysilicon 530 -757 530 -757 0 4
rlabel polysilicon 534 -751 534 -751 0 1
rlabel polysilicon 534 -757 534 -757 0 3
rlabel polysilicon 541 -757 541 -757 0 3
rlabel polysilicon 544 -757 544 -757 0 4
rlabel polysilicon 548 -751 548 -751 0 1
rlabel polysilicon 548 -757 548 -757 0 3
rlabel polysilicon 555 -751 555 -751 0 1
rlabel polysilicon 555 -757 555 -757 0 3
rlabel polysilicon 562 -751 562 -751 0 1
rlabel polysilicon 565 -751 565 -751 0 2
rlabel polysilicon 562 -757 562 -757 0 3
rlabel polysilicon 569 -751 569 -751 0 1
rlabel polysilicon 569 -757 569 -757 0 3
rlabel polysilicon 576 -751 576 -751 0 1
rlabel polysilicon 576 -757 576 -757 0 3
rlabel polysilicon 583 -751 583 -751 0 1
rlabel polysilicon 583 -757 583 -757 0 3
rlabel polysilicon 586 -757 586 -757 0 4
rlabel polysilicon 590 -751 590 -751 0 1
rlabel polysilicon 590 -757 590 -757 0 3
rlabel polysilicon 597 -751 597 -751 0 1
rlabel polysilicon 597 -757 597 -757 0 3
rlabel polysilicon 604 -751 604 -751 0 1
rlabel polysilicon 604 -757 604 -757 0 3
rlabel polysilicon 611 -751 611 -751 0 1
rlabel polysilicon 611 -757 611 -757 0 3
rlabel polysilicon 618 -751 618 -751 0 1
rlabel polysilicon 618 -757 618 -757 0 3
rlabel polysilicon 625 -751 625 -751 0 1
rlabel polysilicon 625 -757 625 -757 0 3
rlabel polysilicon 632 -751 632 -751 0 1
rlabel polysilicon 632 -757 632 -757 0 3
rlabel polysilicon 639 -751 639 -751 0 1
rlabel polysilicon 639 -757 639 -757 0 3
rlabel polysilicon 646 -751 646 -751 0 1
rlabel polysilicon 646 -757 646 -757 0 3
rlabel polysilicon 653 -751 653 -751 0 1
rlabel polysilicon 653 -757 653 -757 0 3
rlabel polysilicon 660 -751 660 -751 0 1
rlabel polysilicon 660 -757 660 -757 0 3
rlabel polysilicon 667 -751 667 -751 0 1
rlabel polysilicon 667 -757 667 -757 0 3
rlabel polysilicon 674 -751 674 -751 0 1
rlabel polysilicon 674 -757 674 -757 0 3
rlabel polysilicon 681 -751 681 -751 0 1
rlabel polysilicon 681 -757 681 -757 0 3
rlabel polysilicon 688 -751 688 -751 0 1
rlabel polysilicon 688 -757 688 -757 0 3
rlabel polysilicon 695 -751 695 -751 0 1
rlabel polysilicon 695 -757 695 -757 0 3
rlabel polysilicon 702 -751 702 -751 0 1
rlabel polysilicon 702 -757 702 -757 0 3
rlabel polysilicon 712 -757 712 -757 0 4
rlabel polysilicon 716 -751 716 -751 0 1
rlabel polysilicon 716 -757 716 -757 0 3
rlabel polysilicon 723 -751 723 -751 0 1
rlabel polysilicon 723 -757 723 -757 0 3
rlabel polysilicon 733 -751 733 -751 0 2
rlabel polysilicon 733 -757 733 -757 0 4
rlabel polysilicon 737 -751 737 -751 0 1
rlabel polysilicon 737 -757 737 -757 0 3
rlabel polysilicon 744 -751 744 -751 0 1
rlabel polysilicon 744 -757 744 -757 0 3
rlabel polysilicon 754 -751 754 -751 0 2
rlabel polysilicon 754 -757 754 -757 0 4
rlabel polysilicon 800 -751 800 -751 0 1
rlabel polysilicon 807 -751 807 -751 0 1
rlabel polysilicon 807 -757 807 -757 0 3
rlabel polysilicon 2 -828 2 -828 0 1
rlabel polysilicon 2 -834 2 -834 0 3
rlabel polysilicon 9 -828 9 -828 0 1
rlabel polysilicon 9 -834 9 -834 0 3
rlabel polysilicon 16 -828 16 -828 0 1
rlabel polysilicon 16 -834 16 -834 0 3
rlabel polysilicon 23 -828 23 -828 0 1
rlabel polysilicon 30 -828 30 -828 0 1
rlabel polysilicon 37 -828 37 -828 0 1
rlabel polysilicon 37 -834 37 -834 0 3
rlabel polysilicon 44 -828 44 -828 0 1
rlabel polysilicon 44 -834 44 -834 0 3
rlabel polysilicon 54 -828 54 -828 0 2
rlabel polysilicon 54 -834 54 -834 0 4
rlabel polysilicon 58 -828 58 -828 0 1
rlabel polysilicon 58 -834 58 -834 0 3
rlabel polysilicon 65 -828 65 -828 0 1
rlabel polysilicon 65 -834 65 -834 0 3
rlabel polysilicon 72 -828 72 -828 0 1
rlabel polysilicon 72 -834 72 -834 0 3
rlabel polysilicon 79 -828 79 -828 0 1
rlabel polysilicon 82 -828 82 -828 0 2
rlabel polysilicon 79 -834 79 -834 0 3
rlabel polysilicon 82 -834 82 -834 0 4
rlabel polysilicon 86 -828 86 -828 0 1
rlabel polysilicon 89 -828 89 -828 0 2
rlabel polysilicon 93 -828 93 -828 0 1
rlabel polysilicon 93 -834 93 -834 0 3
rlabel polysilicon 100 -828 100 -828 0 1
rlabel polysilicon 100 -834 100 -834 0 3
rlabel polysilicon 107 -828 107 -828 0 1
rlabel polysilicon 110 -828 110 -828 0 2
rlabel polysilicon 114 -828 114 -828 0 1
rlabel polysilicon 114 -834 114 -834 0 3
rlabel polysilicon 121 -828 121 -828 0 1
rlabel polysilicon 124 -828 124 -828 0 2
rlabel polysilicon 121 -834 121 -834 0 3
rlabel polysilicon 128 -828 128 -828 0 1
rlabel polysilicon 128 -834 128 -834 0 3
rlabel polysilicon 135 -828 135 -828 0 1
rlabel polysilicon 138 -828 138 -828 0 2
rlabel polysilicon 138 -834 138 -834 0 4
rlabel polysilicon 142 -834 142 -834 0 3
rlabel polysilicon 145 -834 145 -834 0 4
rlabel polysilicon 149 -828 149 -828 0 1
rlabel polysilicon 149 -834 149 -834 0 3
rlabel polysilicon 156 -828 156 -828 0 1
rlabel polysilicon 156 -834 156 -834 0 3
rlabel polysilicon 163 -828 163 -828 0 1
rlabel polysilicon 166 -834 166 -834 0 4
rlabel polysilicon 170 -828 170 -828 0 1
rlabel polysilicon 170 -834 170 -834 0 3
rlabel polysilicon 177 -828 177 -828 0 1
rlabel polysilicon 177 -834 177 -834 0 3
rlabel polysilicon 184 -828 184 -828 0 1
rlabel polysilicon 184 -834 184 -834 0 3
rlabel polysilicon 191 -828 191 -828 0 1
rlabel polysilicon 198 -828 198 -828 0 1
rlabel polysilicon 201 -828 201 -828 0 2
rlabel polysilicon 201 -834 201 -834 0 4
rlabel polysilicon 205 -828 205 -828 0 1
rlabel polysilicon 205 -834 205 -834 0 3
rlabel polysilicon 212 -828 212 -828 0 1
rlabel polysilicon 215 -828 215 -828 0 2
rlabel polysilicon 212 -834 212 -834 0 3
rlabel polysilicon 215 -834 215 -834 0 4
rlabel polysilicon 219 -828 219 -828 0 1
rlabel polysilicon 222 -828 222 -828 0 2
rlabel polysilicon 219 -834 219 -834 0 3
rlabel polysilicon 226 -828 226 -828 0 1
rlabel polysilicon 226 -834 226 -834 0 3
rlabel polysilicon 233 -828 233 -828 0 1
rlabel polysilicon 233 -834 233 -834 0 3
rlabel polysilicon 240 -828 240 -828 0 1
rlabel polysilicon 243 -828 243 -828 0 2
rlabel polysilicon 240 -834 240 -834 0 3
rlabel polysilicon 247 -828 247 -828 0 1
rlabel polysilicon 247 -834 247 -834 0 3
rlabel polysilicon 254 -828 254 -828 0 1
rlabel polysilicon 254 -834 254 -834 0 3
rlabel polysilicon 264 -828 264 -828 0 2
rlabel polysilicon 268 -828 268 -828 0 1
rlabel polysilicon 268 -834 268 -834 0 3
rlabel polysilicon 275 -828 275 -828 0 1
rlabel polysilicon 275 -834 275 -834 0 3
rlabel polysilicon 285 -828 285 -828 0 2
rlabel polysilicon 282 -834 282 -834 0 3
rlabel polysilicon 289 -828 289 -828 0 1
rlabel polysilicon 292 -828 292 -828 0 2
rlabel polysilicon 292 -834 292 -834 0 4
rlabel polysilicon 296 -828 296 -828 0 1
rlabel polysilicon 299 -828 299 -828 0 2
rlabel polysilicon 296 -834 296 -834 0 3
rlabel polysilicon 299 -834 299 -834 0 4
rlabel polysilicon 303 -828 303 -828 0 1
rlabel polysilicon 303 -834 303 -834 0 3
rlabel polysilicon 310 -828 310 -828 0 1
rlabel polysilicon 310 -834 310 -834 0 3
rlabel polysilicon 317 -828 317 -828 0 1
rlabel polysilicon 317 -834 317 -834 0 3
rlabel polysilicon 324 -828 324 -828 0 1
rlabel polysilicon 324 -834 324 -834 0 3
rlabel polysilicon 331 -828 331 -828 0 1
rlabel polysilicon 334 -828 334 -828 0 2
rlabel polysilicon 331 -834 331 -834 0 3
rlabel polysilicon 334 -834 334 -834 0 4
rlabel polysilicon 338 -828 338 -828 0 1
rlabel polysilicon 338 -834 338 -834 0 3
rlabel polysilicon 345 -828 345 -828 0 1
rlabel polysilicon 345 -834 345 -834 0 3
rlabel polysilicon 352 -828 352 -828 0 1
rlabel polysilicon 352 -834 352 -834 0 3
rlabel polysilicon 359 -828 359 -828 0 1
rlabel polysilicon 359 -834 359 -834 0 3
rlabel polysilicon 366 -828 366 -828 0 1
rlabel polysilicon 366 -834 366 -834 0 3
rlabel polysilicon 373 -828 373 -828 0 1
rlabel polysilicon 373 -834 373 -834 0 3
rlabel polysilicon 380 -828 380 -828 0 1
rlabel polysilicon 383 -828 383 -828 0 2
rlabel polysilicon 380 -834 380 -834 0 3
rlabel polysilicon 387 -828 387 -828 0 1
rlabel polysilicon 390 -828 390 -828 0 2
rlabel polysilicon 390 -834 390 -834 0 4
rlabel polysilicon 394 -828 394 -828 0 1
rlabel polysilicon 394 -834 394 -834 0 3
rlabel polysilicon 404 -828 404 -828 0 2
rlabel polysilicon 401 -834 401 -834 0 3
rlabel polysilicon 404 -834 404 -834 0 4
rlabel polysilicon 408 -828 408 -828 0 1
rlabel polysilicon 408 -834 408 -834 0 3
rlabel polysilicon 418 -828 418 -828 0 2
rlabel polysilicon 418 -834 418 -834 0 4
rlabel polysilicon 422 -828 422 -828 0 1
rlabel polysilicon 422 -834 422 -834 0 3
rlabel polysilicon 429 -828 429 -828 0 1
rlabel polysilicon 429 -834 429 -834 0 3
rlabel polysilicon 436 -828 436 -828 0 1
rlabel polysilicon 439 -828 439 -828 0 2
rlabel polysilicon 436 -834 436 -834 0 3
rlabel polysilicon 439 -834 439 -834 0 4
rlabel polysilicon 443 -828 443 -828 0 1
rlabel polysilicon 443 -834 443 -834 0 3
rlabel polysilicon 450 -828 450 -828 0 1
rlabel polysilicon 450 -834 450 -834 0 3
rlabel polysilicon 457 -828 457 -828 0 1
rlabel polysilicon 460 -828 460 -828 0 2
rlabel polysilicon 460 -834 460 -834 0 4
rlabel polysilicon 464 -828 464 -828 0 1
rlabel polysilicon 464 -834 464 -834 0 3
rlabel polysilicon 471 -828 471 -828 0 1
rlabel polysilicon 471 -834 471 -834 0 3
rlabel polysilicon 478 -828 478 -828 0 1
rlabel polysilicon 478 -834 478 -834 0 3
rlabel polysilicon 488 -828 488 -828 0 2
rlabel polysilicon 485 -834 485 -834 0 3
rlabel polysilicon 488 -834 488 -834 0 4
rlabel polysilicon 495 -828 495 -828 0 2
rlabel polysilicon 495 -834 495 -834 0 4
rlabel polysilicon 499 -828 499 -828 0 1
rlabel polysilicon 499 -834 499 -834 0 3
rlabel polysilicon 506 -828 506 -828 0 1
rlabel polysilicon 506 -834 506 -834 0 3
rlabel polysilicon 513 -828 513 -828 0 1
rlabel polysilicon 513 -834 513 -834 0 3
rlabel polysilicon 520 -828 520 -828 0 1
rlabel polysilicon 523 -828 523 -828 0 2
rlabel polysilicon 523 -834 523 -834 0 4
rlabel polysilicon 527 -834 527 -834 0 3
rlabel polysilicon 530 -834 530 -834 0 4
rlabel polysilicon 534 -828 534 -828 0 1
rlabel polysilicon 534 -834 534 -834 0 3
rlabel polysilicon 541 -828 541 -828 0 1
rlabel polysilicon 541 -834 541 -834 0 3
rlabel polysilicon 548 -828 548 -828 0 1
rlabel polysilicon 548 -834 548 -834 0 3
rlabel polysilicon 555 -828 555 -828 0 1
rlabel polysilicon 555 -834 555 -834 0 3
rlabel polysilicon 562 -828 562 -828 0 1
rlabel polysilicon 562 -834 562 -834 0 3
rlabel polysilicon 569 -828 569 -828 0 1
rlabel polysilicon 569 -834 569 -834 0 3
rlabel polysilicon 576 -828 576 -828 0 1
rlabel polysilicon 576 -834 576 -834 0 3
rlabel polysilicon 583 -828 583 -828 0 1
rlabel polysilicon 583 -834 583 -834 0 3
rlabel polysilicon 590 -828 590 -828 0 1
rlabel polysilicon 590 -834 590 -834 0 3
rlabel polysilicon 597 -828 597 -828 0 1
rlabel polysilicon 597 -834 597 -834 0 3
rlabel polysilicon 604 -828 604 -828 0 1
rlabel polysilicon 604 -834 604 -834 0 3
rlabel polysilicon 611 -828 611 -828 0 1
rlabel polysilicon 611 -834 611 -834 0 3
rlabel polysilicon 618 -828 618 -828 0 1
rlabel polysilicon 618 -834 618 -834 0 3
rlabel polysilicon 625 -828 625 -828 0 1
rlabel polysilicon 625 -834 625 -834 0 3
rlabel polysilicon 632 -828 632 -828 0 1
rlabel polysilicon 632 -834 632 -834 0 3
rlabel polysilicon 639 -828 639 -828 0 1
rlabel polysilicon 639 -834 639 -834 0 3
rlabel polysilicon 646 -828 646 -828 0 1
rlabel polysilicon 646 -834 646 -834 0 3
rlabel polysilicon 653 -828 653 -828 0 1
rlabel polysilicon 653 -834 653 -834 0 3
rlabel polysilicon 660 -828 660 -828 0 1
rlabel polysilicon 660 -834 660 -834 0 3
rlabel polysilicon 667 -828 667 -828 0 1
rlabel polysilicon 667 -834 667 -834 0 3
rlabel polysilicon 674 -828 674 -828 0 1
rlabel polysilicon 674 -834 674 -834 0 3
rlabel polysilicon 681 -828 681 -828 0 1
rlabel polysilicon 681 -834 681 -834 0 3
rlabel polysilicon 688 -828 688 -828 0 1
rlabel polysilicon 688 -834 688 -834 0 3
rlabel polysilicon 695 -828 695 -828 0 1
rlabel polysilicon 695 -834 695 -834 0 3
rlabel polysilicon 702 -828 702 -828 0 1
rlabel polysilicon 702 -834 702 -834 0 3
rlabel polysilicon 709 -828 709 -828 0 1
rlabel polysilicon 709 -834 709 -834 0 3
rlabel polysilicon 716 -828 716 -828 0 1
rlabel polysilicon 716 -834 716 -834 0 3
rlabel polysilicon 723 -828 723 -828 0 1
rlabel polysilicon 723 -834 723 -834 0 3
rlabel polysilicon 730 -828 730 -828 0 1
rlabel polysilicon 730 -834 730 -834 0 3
rlabel polysilicon 737 -828 737 -828 0 1
rlabel polysilicon 737 -834 737 -834 0 3
rlabel polysilicon 744 -828 744 -828 0 1
rlabel polysilicon 744 -834 744 -834 0 3
rlabel polysilicon 751 -828 751 -828 0 1
rlabel polysilicon 751 -834 751 -834 0 3
rlabel polysilicon 758 -828 758 -828 0 1
rlabel polysilicon 758 -834 758 -834 0 3
rlabel polysilicon 765 -828 765 -828 0 1
rlabel polysilicon 765 -834 765 -834 0 3
rlabel polysilicon 772 -828 772 -828 0 1
rlabel polysilicon 772 -834 772 -834 0 3
rlabel polysilicon 779 -828 779 -828 0 1
rlabel polysilicon 779 -834 779 -834 0 3
rlabel polysilicon 786 -828 786 -828 0 1
rlabel polysilicon 786 -834 786 -834 0 3
rlabel polysilicon 793 -828 793 -828 0 1
rlabel polysilicon 793 -834 793 -834 0 3
rlabel polysilicon 803 -828 803 -828 0 2
rlabel polysilicon 803 -834 803 -834 0 4
rlabel polysilicon 807 -828 807 -828 0 1
rlabel polysilicon 807 -834 807 -834 0 3
rlabel polysilicon 9 -915 9 -915 0 1
rlabel polysilicon 9 -921 9 -921 0 3
rlabel polysilicon 16 -915 16 -915 0 1
rlabel polysilicon 16 -921 16 -921 0 3
rlabel polysilicon 23 -915 23 -915 0 1
rlabel polysilicon 23 -921 23 -921 0 3
rlabel polysilicon 30 -915 30 -915 0 1
rlabel polysilicon 30 -921 30 -921 0 3
rlabel polysilicon 37 -915 37 -915 0 1
rlabel polysilicon 37 -921 37 -921 0 3
rlabel polysilicon 44 -915 44 -915 0 1
rlabel polysilicon 44 -921 44 -921 0 3
rlabel polysilicon 51 -915 51 -915 0 1
rlabel polysilicon 51 -921 51 -921 0 3
rlabel polysilicon 58 -915 58 -915 0 1
rlabel polysilicon 58 -921 58 -921 0 3
rlabel polysilicon 65 -915 65 -915 0 1
rlabel polysilicon 72 -915 72 -915 0 1
rlabel polysilicon 79 -915 79 -915 0 1
rlabel polysilicon 79 -921 79 -921 0 3
rlabel polysilicon 86 -915 86 -915 0 1
rlabel polysilicon 86 -921 86 -921 0 3
rlabel polysilicon 89 -921 89 -921 0 4
rlabel polysilicon 93 -915 93 -915 0 1
rlabel polysilicon 93 -921 93 -921 0 3
rlabel polysilicon 100 -915 100 -915 0 1
rlabel polysilicon 100 -921 100 -921 0 3
rlabel polysilicon 107 -915 107 -915 0 1
rlabel polysilicon 107 -921 107 -921 0 3
rlabel polysilicon 114 -915 114 -915 0 1
rlabel polysilicon 114 -921 114 -921 0 3
rlabel polysilicon 121 -915 121 -915 0 1
rlabel polysilicon 121 -921 121 -921 0 3
rlabel polysilicon 128 -915 128 -915 0 1
rlabel polysilicon 135 -915 135 -915 0 1
rlabel polysilicon 135 -921 135 -921 0 3
rlabel polysilicon 142 -915 142 -915 0 1
rlabel polysilicon 142 -921 142 -921 0 3
rlabel polysilicon 149 -915 149 -915 0 1
rlabel polysilicon 152 -915 152 -915 0 2
rlabel polysilicon 149 -921 149 -921 0 3
rlabel polysilicon 152 -921 152 -921 0 4
rlabel polysilicon 156 -915 156 -915 0 1
rlabel polysilicon 159 -915 159 -915 0 2
rlabel polysilicon 163 -915 163 -915 0 1
rlabel polysilicon 163 -921 163 -921 0 3
rlabel polysilicon 170 -915 170 -915 0 1
rlabel polysilicon 173 -915 173 -915 0 2
rlabel polysilicon 177 -915 177 -915 0 1
rlabel polysilicon 180 -915 180 -915 0 2
rlabel polysilicon 180 -921 180 -921 0 4
rlabel polysilicon 184 -915 184 -915 0 1
rlabel polysilicon 184 -921 184 -921 0 3
rlabel polysilicon 191 -915 191 -915 0 1
rlabel polysilicon 191 -921 191 -921 0 3
rlabel polysilicon 201 -915 201 -915 0 2
rlabel polysilicon 198 -921 198 -921 0 3
rlabel polysilicon 201 -921 201 -921 0 4
rlabel polysilicon 205 -915 205 -915 0 1
rlabel polysilicon 205 -921 205 -921 0 3
rlabel polysilicon 212 -915 212 -915 0 1
rlabel polysilicon 212 -921 212 -921 0 3
rlabel polysilicon 219 -915 219 -915 0 1
rlabel polysilicon 219 -921 219 -921 0 3
rlabel polysilicon 222 -921 222 -921 0 4
rlabel polysilicon 226 -915 226 -915 0 1
rlabel polysilicon 229 -915 229 -915 0 2
rlabel polysilicon 226 -921 226 -921 0 3
rlabel polysilicon 229 -921 229 -921 0 4
rlabel polysilicon 233 -915 233 -915 0 1
rlabel polysilicon 236 -915 236 -915 0 2
rlabel polysilicon 233 -921 233 -921 0 3
rlabel polysilicon 236 -921 236 -921 0 4
rlabel polysilicon 240 -915 240 -915 0 1
rlabel polysilicon 243 -915 243 -915 0 2
rlabel polysilicon 243 -921 243 -921 0 4
rlabel polysilicon 247 -915 247 -915 0 1
rlabel polysilicon 247 -921 247 -921 0 3
rlabel polysilicon 254 -915 254 -915 0 1
rlabel polysilicon 254 -921 254 -921 0 3
rlabel polysilicon 261 -915 261 -915 0 1
rlabel polysilicon 261 -921 261 -921 0 3
rlabel polysilicon 268 -915 268 -915 0 1
rlabel polysilicon 268 -921 268 -921 0 3
rlabel polysilicon 275 -915 275 -915 0 1
rlabel polysilicon 278 -915 278 -915 0 2
rlabel polysilicon 275 -921 275 -921 0 3
rlabel polysilicon 278 -921 278 -921 0 4
rlabel polysilicon 282 -915 282 -915 0 1
rlabel polysilicon 285 -921 285 -921 0 4
rlabel polysilicon 289 -915 289 -915 0 1
rlabel polysilicon 289 -921 289 -921 0 3
rlabel polysilicon 296 -915 296 -915 0 1
rlabel polysilicon 296 -921 296 -921 0 3
rlabel polysilicon 303 -915 303 -915 0 1
rlabel polysilicon 303 -921 303 -921 0 3
rlabel polysilicon 310 -915 310 -915 0 1
rlabel polysilicon 310 -921 310 -921 0 3
rlabel polysilicon 317 -915 317 -915 0 1
rlabel polysilicon 317 -921 317 -921 0 3
rlabel polysilicon 324 -915 324 -915 0 1
rlabel polysilicon 324 -921 324 -921 0 3
rlabel polysilicon 331 -915 331 -915 0 1
rlabel polysilicon 331 -921 331 -921 0 3
rlabel polysilicon 338 -915 338 -915 0 1
rlabel polysilicon 338 -921 338 -921 0 3
rlabel polysilicon 348 -915 348 -915 0 2
rlabel polysilicon 345 -921 345 -921 0 3
rlabel polysilicon 348 -921 348 -921 0 4
rlabel polysilicon 352 -915 352 -915 0 1
rlabel polysilicon 352 -921 352 -921 0 3
rlabel polysilicon 359 -915 359 -915 0 1
rlabel polysilicon 359 -921 359 -921 0 3
rlabel polysilicon 366 -915 366 -915 0 1
rlabel polysilicon 366 -921 366 -921 0 3
rlabel polysilicon 373 -915 373 -915 0 1
rlabel polysilicon 373 -921 373 -921 0 3
rlabel polysilicon 383 -915 383 -915 0 2
rlabel polysilicon 380 -921 380 -921 0 3
rlabel polysilicon 387 -915 387 -915 0 1
rlabel polysilicon 387 -921 387 -921 0 3
rlabel polysilicon 394 -915 394 -915 0 1
rlabel polysilicon 397 -915 397 -915 0 2
rlabel polysilicon 394 -921 394 -921 0 3
rlabel polysilicon 397 -921 397 -921 0 4
rlabel polysilicon 401 -915 401 -915 0 1
rlabel polysilicon 401 -921 401 -921 0 3
rlabel polysilicon 408 -915 408 -915 0 1
rlabel polysilicon 411 -915 411 -915 0 2
rlabel polysilicon 408 -921 408 -921 0 3
rlabel polysilicon 411 -921 411 -921 0 4
rlabel polysilicon 415 -915 415 -915 0 1
rlabel polysilicon 415 -921 415 -921 0 3
rlabel polysilicon 418 -921 418 -921 0 4
rlabel polysilicon 422 -915 422 -915 0 1
rlabel polysilicon 422 -921 422 -921 0 3
rlabel polysilicon 429 -915 429 -915 0 1
rlabel polysilicon 429 -921 429 -921 0 3
rlabel polysilicon 436 -915 436 -915 0 1
rlabel polysilicon 436 -921 436 -921 0 3
rlabel polysilicon 443 -915 443 -915 0 1
rlabel polysilicon 443 -921 443 -921 0 3
rlabel polysilicon 450 -915 450 -915 0 1
rlabel polysilicon 450 -921 450 -921 0 3
rlabel polysilicon 457 -915 457 -915 0 1
rlabel polysilicon 460 -915 460 -915 0 2
rlabel polysilicon 457 -921 457 -921 0 3
rlabel polysilicon 460 -921 460 -921 0 4
rlabel polysilicon 464 -915 464 -915 0 1
rlabel polysilicon 467 -915 467 -915 0 2
rlabel polysilicon 467 -921 467 -921 0 4
rlabel polysilicon 471 -915 471 -915 0 1
rlabel polysilicon 471 -921 471 -921 0 3
rlabel polysilicon 478 -915 478 -915 0 1
rlabel polysilicon 478 -921 478 -921 0 3
rlabel polysilicon 488 -915 488 -915 0 2
rlabel polysilicon 488 -921 488 -921 0 4
rlabel polysilicon 492 -915 492 -915 0 1
rlabel polysilicon 492 -921 492 -921 0 3
rlabel polysilicon 499 -915 499 -915 0 1
rlabel polysilicon 499 -921 499 -921 0 3
rlabel polysilicon 502 -921 502 -921 0 4
rlabel polysilicon 506 -915 506 -915 0 1
rlabel polysilicon 506 -921 506 -921 0 3
rlabel polysilicon 513 -915 513 -915 0 1
rlabel polysilicon 513 -921 513 -921 0 3
rlabel polysilicon 520 -915 520 -915 0 1
rlabel polysilicon 520 -921 520 -921 0 3
rlabel polysilicon 527 -915 527 -915 0 1
rlabel polysilicon 527 -921 527 -921 0 3
rlabel polysilicon 534 -915 534 -915 0 1
rlabel polysilicon 534 -921 534 -921 0 3
rlabel polysilicon 541 -915 541 -915 0 1
rlabel polysilicon 541 -921 541 -921 0 3
rlabel polysilicon 548 -915 548 -915 0 1
rlabel polysilicon 548 -921 548 -921 0 3
rlabel polysilicon 555 -915 555 -915 0 1
rlabel polysilicon 555 -921 555 -921 0 3
rlabel polysilicon 562 -915 562 -915 0 1
rlabel polysilicon 562 -921 562 -921 0 3
rlabel polysilicon 569 -915 569 -915 0 1
rlabel polysilicon 569 -921 569 -921 0 3
rlabel polysilicon 576 -921 576 -921 0 3
rlabel polysilicon 579 -921 579 -921 0 4
rlabel polysilicon 583 -915 583 -915 0 1
rlabel polysilicon 583 -921 583 -921 0 3
rlabel polysilicon 590 -915 590 -915 0 1
rlabel polysilicon 590 -921 590 -921 0 3
rlabel polysilicon 597 -915 597 -915 0 1
rlabel polysilicon 597 -921 597 -921 0 3
rlabel polysilicon 604 -915 604 -915 0 1
rlabel polysilicon 604 -921 604 -921 0 3
rlabel polysilicon 611 -915 611 -915 0 1
rlabel polysilicon 611 -921 611 -921 0 3
rlabel polysilicon 618 -915 618 -915 0 1
rlabel polysilicon 618 -921 618 -921 0 3
rlabel polysilicon 625 -915 625 -915 0 1
rlabel polysilicon 625 -921 625 -921 0 3
rlabel polysilicon 632 -915 632 -915 0 1
rlabel polysilicon 632 -921 632 -921 0 3
rlabel polysilicon 639 -915 639 -915 0 1
rlabel polysilicon 639 -921 639 -921 0 3
rlabel polysilicon 646 -915 646 -915 0 1
rlabel polysilicon 646 -921 646 -921 0 3
rlabel polysilicon 653 -915 653 -915 0 1
rlabel polysilicon 653 -921 653 -921 0 3
rlabel polysilicon 660 -915 660 -915 0 1
rlabel polysilicon 660 -921 660 -921 0 3
rlabel polysilicon 667 -915 667 -915 0 1
rlabel polysilicon 667 -921 667 -921 0 3
rlabel polysilicon 674 -915 674 -915 0 1
rlabel polysilicon 674 -921 674 -921 0 3
rlabel polysilicon 681 -915 681 -915 0 1
rlabel polysilicon 681 -921 681 -921 0 3
rlabel polysilicon 688 -915 688 -915 0 1
rlabel polysilicon 688 -921 688 -921 0 3
rlabel polysilicon 695 -915 695 -915 0 1
rlabel polysilicon 695 -921 695 -921 0 3
rlabel polysilicon 702 -915 702 -915 0 1
rlabel polysilicon 702 -921 702 -921 0 3
rlabel polysilicon 709 -915 709 -915 0 1
rlabel polysilicon 709 -921 709 -921 0 3
rlabel polysilicon 716 -915 716 -915 0 1
rlabel polysilicon 716 -921 716 -921 0 3
rlabel polysilicon 723 -915 723 -915 0 1
rlabel polysilicon 723 -921 723 -921 0 3
rlabel polysilicon 730 -915 730 -915 0 1
rlabel polysilicon 730 -921 730 -921 0 3
rlabel polysilicon 737 -915 737 -915 0 1
rlabel polysilicon 737 -921 737 -921 0 3
rlabel polysilicon 744 -915 744 -915 0 1
rlabel polysilicon 744 -921 744 -921 0 3
rlabel polysilicon 751 -915 751 -915 0 1
rlabel polysilicon 751 -921 751 -921 0 3
rlabel polysilicon 758 -915 758 -915 0 1
rlabel polysilicon 758 -921 758 -921 0 3
rlabel polysilicon 765 -915 765 -915 0 1
rlabel polysilicon 765 -921 765 -921 0 3
rlabel polysilicon 772 -915 772 -915 0 1
rlabel polysilicon 775 -915 775 -915 0 2
rlabel polysilicon 772 -921 772 -921 0 3
rlabel polysilicon 775 -921 775 -921 0 4
rlabel polysilicon 782 -915 782 -915 0 2
rlabel polysilicon 779 -921 779 -921 0 3
rlabel polysilicon 786 -915 786 -915 0 1
rlabel polysilicon 786 -921 786 -921 0 3
rlabel polysilicon 796 -915 796 -915 0 2
rlabel polysilicon 9 -992 9 -992 0 1
rlabel polysilicon 9 -998 9 -998 0 3
rlabel polysilicon 16 -992 16 -992 0 1
rlabel polysilicon 16 -998 16 -998 0 3
rlabel polysilicon 23 -992 23 -992 0 1
rlabel polysilicon 23 -998 23 -998 0 3
rlabel polysilicon 30 -992 30 -992 0 1
rlabel polysilicon 30 -998 30 -998 0 3
rlabel polysilicon 37 -992 37 -992 0 1
rlabel polysilicon 37 -998 37 -998 0 3
rlabel polysilicon 44 -992 44 -992 0 1
rlabel polysilicon 44 -998 44 -998 0 3
rlabel polysilicon 51 -992 51 -992 0 1
rlabel polysilicon 51 -998 51 -998 0 3
rlabel polysilicon 58 -992 58 -992 0 1
rlabel polysilicon 58 -998 58 -998 0 3
rlabel polysilicon 65 -992 65 -992 0 1
rlabel polysilicon 65 -998 65 -998 0 3
rlabel polysilicon 75 -992 75 -992 0 2
rlabel polysilicon 72 -998 72 -998 0 3
rlabel polysilicon 79 -992 79 -992 0 1
rlabel polysilicon 82 -992 82 -992 0 2
rlabel polysilicon 79 -998 79 -998 0 3
rlabel polysilicon 86 -992 86 -992 0 1
rlabel polysilicon 86 -998 86 -998 0 3
rlabel polysilicon 96 -992 96 -992 0 2
rlabel polysilicon 96 -998 96 -998 0 4
rlabel polysilicon 100 -992 100 -992 0 1
rlabel polysilicon 103 -992 103 -992 0 2
rlabel polysilicon 107 -992 107 -992 0 1
rlabel polysilicon 107 -998 107 -998 0 3
rlabel polysilicon 114 -992 114 -992 0 1
rlabel polysilicon 117 -992 117 -992 0 2
rlabel polysilicon 114 -998 114 -998 0 3
rlabel polysilicon 117 -998 117 -998 0 4
rlabel polysilicon 121 -992 121 -992 0 1
rlabel polysilicon 121 -998 121 -998 0 3
rlabel polysilicon 128 -992 128 -992 0 1
rlabel polysilicon 128 -998 128 -998 0 3
rlabel polysilicon 135 -992 135 -992 0 1
rlabel polysilicon 135 -998 135 -998 0 3
rlabel polysilicon 142 -992 142 -992 0 1
rlabel polysilicon 142 -998 142 -998 0 3
rlabel polysilicon 149 -992 149 -992 0 1
rlabel polysilicon 149 -998 149 -998 0 3
rlabel polysilicon 159 -992 159 -992 0 2
rlabel polysilicon 156 -998 156 -998 0 3
rlabel polysilicon 159 -998 159 -998 0 4
rlabel polysilicon 163 -992 163 -992 0 1
rlabel polysilicon 163 -998 163 -998 0 3
rlabel polysilicon 170 -992 170 -992 0 1
rlabel polysilicon 170 -998 170 -998 0 3
rlabel polysilicon 177 -992 177 -992 0 1
rlabel polysilicon 177 -998 177 -998 0 3
rlabel polysilicon 184 -992 184 -992 0 1
rlabel polysilicon 184 -998 184 -998 0 3
rlabel polysilicon 191 -992 191 -992 0 1
rlabel polysilicon 191 -998 191 -998 0 3
rlabel polysilicon 198 -992 198 -992 0 1
rlabel polysilicon 198 -998 198 -998 0 3
rlabel polysilicon 205 -992 205 -992 0 1
rlabel polysilicon 205 -998 205 -998 0 3
rlabel polysilicon 212 -992 212 -992 0 1
rlabel polysilicon 212 -998 212 -998 0 3
rlabel polysilicon 219 -992 219 -992 0 1
rlabel polysilicon 219 -998 219 -998 0 3
rlabel polysilicon 222 -998 222 -998 0 4
rlabel polysilicon 226 -992 226 -992 0 1
rlabel polysilicon 226 -998 226 -998 0 3
rlabel polysilicon 233 -992 233 -992 0 1
rlabel polysilicon 236 -992 236 -992 0 2
rlabel polysilicon 233 -998 233 -998 0 3
rlabel polysilicon 240 -992 240 -992 0 1
rlabel polysilicon 243 -992 243 -992 0 2
rlabel polysilicon 240 -998 240 -998 0 3
rlabel polysilicon 243 -998 243 -998 0 4
rlabel polysilicon 247 -992 247 -992 0 1
rlabel polysilicon 247 -998 247 -998 0 3
rlabel polysilicon 254 -992 254 -992 0 1
rlabel polysilicon 257 -992 257 -992 0 2
rlabel polysilicon 254 -998 254 -998 0 3
rlabel polysilicon 261 -992 261 -992 0 1
rlabel polysilicon 261 -998 261 -998 0 3
rlabel polysilicon 268 -992 268 -992 0 1
rlabel polysilicon 268 -998 268 -998 0 3
rlabel polysilicon 275 -992 275 -992 0 1
rlabel polysilicon 275 -998 275 -998 0 3
rlabel polysilicon 285 -992 285 -992 0 2
rlabel polysilicon 282 -998 282 -998 0 3
rlabel polysilicon 289 -992 289 -992 0 1
rlabel polysilicon 289 -998 289 -998 0 3
rlabel polysilicon 296 -992 296 -992 0 1
rlabel polysilicon 296 -998 296 -998 0 3
rlabel polysilicon 303 -992 303 -992 0 1
rlabel polysilicon 303 -998 303 -998 0 3
rlabel polysilicon 310 -992 310 -992 0 1
rlabel polysilicon 313 -992 313 -992 0 2
rlabel polysilicon 310 -998 310 -998 0 3
rlabel polysilicon 313 -998 313 -998 0 4
rlabel polysilicon 317 -992 317 -992 0 1
rlabel polysilicon 317 -998 317 -998 0 3
rlabel polysilicon 324 -992 324 -992 0 1
rlabel polysilicon 324 -998 324 -998 0 3
rlabel polysilicon 331 -992 331 -992 0 1
rlabel polysilicon 331 -998 331 -998 0 3
rlabel polysilicon 338 -992 338 -992 0 1
rlabel polysilicon 338 -998 338 -998 0 3
rlabel polysilicon 348 -992 348 -992 0 2
rlabel polysilicon 345 -998 345 -998 0 3
rlabel polysilicon 348 -998 348 -998 0 4
rlabel polysilicon 352 -998 352 -998 0 3
rlabel polysilicon 355 -998 355 -998 0 4
rlabel polysilicon 362 -992 362 -992 0 2
rlabel polysilicon 362 -998 362 -998 0 4
rlabel polysilicon 369 -998 369 -998 0 4
rlabel polysilicon 376 -992 376 -992 0 2
rlabel polysilicon 373 -998 373 -998 0 3
rlabel polysilicon 376 -998 376 -998 0 4
rlabel polysilicon 380 -992 380 -992 0 1
rlabel polysilicon 380 -998 380 -998 0 3
rlabel polysilicon 390 -992 390 -992 0 2
rlabel polysilicon 397 -992 397 -992 0 2
rlabel polysilicon 397 -998 397 -998 0 4
rlabel polysilicon 401 -992 401 -992 0 1
rlabel polysilicon 401 -998 401 -998 0 3
rlabel polysilicon 408 -992 408 -992 0 1
rlabel polysilicon 408 -998 408 -998 0 3
rlabel polysilicon 418 -992 418 -992 0 2
rlabel polysilicon 415 -998 415 -998 0 3
rlabel polysilicon 425 -992 425 -992 0 2
rlabel polysilicon 425 -998 425 -998 0 4
rlabel polysilicon 429 -992 429 -992 0 1
rlabel polysilicon 432 -992 432 -992 0 2
rlabel polysilicon 432 -998 432 -998 0 4
rlabel polysilicon 436 -992 436 -992 0 1
rlabel polysilicon 436 -998 436 -998 0 3
rlabel polysilicon 443 -992 443 -992 0 1
rlabel polysilicon 446 -992 446 -992 0 2
rlabel polysilicon 443 -998 443 -998 0 3
rlabel polysilicon 446 -998 446 -998 0 4
rlabel polysilicon 450 -992 450 -992 0 1
rlabel polysilicon 453 -998 453 -998 0 4
rlabel polysilicon 457 -992 457 -992 0 1
rlabel polysilicon 457 -998 457 -998 0 3
rlabel polysilicon 464 -992 464 -992 0 1
rlabel polysilicon 467 -998 467 -998 0 4
rlabel polysilicon 471 -992 471 -992 0 1
rlabel polysilicon 474 -992 474 -992 0 2
rlabel polysilicon 471 -998 471 -998 0 3
rlabel polysilicon 478 -992 478 -992 0 1
rlabel polysilicon 478 -998 478 -998 0 3
rlabel polysilicon 485 -992 485 -992 0 1
rlabel polysilicon 485 -998 485 -998 0 3
rlabel polysilicon 492 -992 492 -992 0 1
rlabel polysilicon 492 -998 492 -998 0 3
rlabel polysilicon 499 -992 499 -992 0 1
rlabel polysilicon 499 -998 499 -998 0 3
rlabel polysilicon 506 -992 506 -992 0 1
rlabel polysilicon 506 -998 506 -998 0 3
rlabel polysilicon 513 -992 513 -992 0 1
rlabel polysilicon 513 -998 513 -998 0 3
rlabel polysilicon 520 -992 520 -992 0 1
rlabel polysilicon 520 -998 520 -998 0 3
rlabel polysilicon 527 -992 527 -992 0 1
rlabel polysilicon 527 -998 527 -998 0 3
rlabel polysilicon 534 -992 534 -992 0 1
rlabel polysilicon 534 -998 534 -998 0 3
rlabel polysilicon 541 -992 541 -992 0 1
rlabel polysilicon 541 -998 541 -998 0 3
rlabel polysilicon 548 -992 548 -992 0 1
rlabel polysilicon 548 -998 548 -998 0 3
rlabel polysilicon 555 -992 555 -992 0 1
rlabel polysilicon 555 -998 555 -998 0 3
rlabel polysilicon 562 -992 562 -992 0 1
rlabel polysilicon 562 -998 562 -998 0 3
rlabel polysilicon 569 -992 569 -992 0 1
rlabel polysilicon 569 -998 569 -998 0 3
rlabel polysilicon 576 -992 576 -992 0 1
rlabel polysilicon 576 -998 576 -998 0 3
rlabel polysilicon 583 -992 583 -992 0 1
rlabel polysilicon 583 -998 583 -998 0 3
rlabel polysilicon 590 -992 590 -992 0 1
rlabel polysilicon 590 -998 590 -998 0 3
rlabel polysilicon 597 -992 597 -992 0 1
rlabel polysilicon 597 -998 597 -998 0 3
rlabel polysilicon 604 -992 604 -992 0 1
rlabel polysilicon 604 -998 604 -998 0 3
rlabel polysilicon 611 -992 611 -992 0 1
rlabel polysilicon 611 -998 611 -998 0 3
rlabel polysilicon 618 -992 618 -992 0 1
rlabel polysilicon 618 -998 618 -998 0 3
rlabel polysilicon 625 -992 625 -992 0 1
rlabel polysilicon 625 -998 625 -998 0 3
rlabel polysilicon 632 -992 632 -992 0 1
rlabel polysilicon 632 -998 632 -998 0 3
rlabel polysilicon 639 -992 639 -992 0 1
rlabel polysilicon 639 -998 639 -998 0 3
rlabel polysilicon 646 -992 646 -992 0 1
rlabel polysilicon 646 -998 646 -998 0 3
rlabel polysilicon 653 -992 653 -992 0 1
rlabel polysilicon 653 -998 653 -998 0 3
rlabel polysilicon 660 -992 660 -992 0 1
rlabel polysilicon 660 -998 660 -998 0 3
rlabel polysilicon 667 -992 667 -992 0 1
rlabel polysilicon 667 -998 667 -998 0 3
rlabel polysilicon 674 -992 674 -992 0 1
rlabel polysilicon 674 -998 674 -998 0 3
rlabel polysilicon 681 -992 681 -992 0 1
rlabel polysilicon 681 -998 681 -998 0 3
rlabel polysilicon 688 -992 688 -992 0 1
rlabel polysilicon 688 -998 688 -998 0 3
rlabel polysilicon 695 -992 695 -992 0 1
rlabel polysilicon 695 -998 695 -998 0 3
rlabel polysilicon 702 -992 702 -992 0 1
rlabel polysilicon 702 -998 702 -998 0 3
rlabel polysilicon 709 -992 709 -992 0 1
rlabel polysilicon 709 -998 709 -998 0 3
rlabel polysilicon 716 -992 716 -992 0 1
rlabel polysilicon 716 -998 716 -998 0 3
rlabel polysilicon 723 -992 723 -992 0 1
rlabel polysilicon 723 -998 723 -998 0 3
rlabel polysilicon 730 -992 730 -992 0 1
rlabel polysilicon 730 -998 730 -998 0 3
rlabel polysilicon 737 -992 737 -992 0 1
rlabel polysilicon 740 -992 740 -992 0 2
rlabel polysilicon 737 -998 737 -998 0 3
rlabel polysilicon 740 -998 740 -998 0 4
rlabel polysilicon 744 -998 744 -998 0 3
rlabel polysilicon 754 -992 754 -992 0 2
rlabel polysilicon 754 -998 754 -998 0 4
rlabel polysilicon 758 -992 758 -992 0 1
rlabel polysilicon 758 -998 758 -998 0 3
rlabel polysilicon 23 -1067 23 -1067 0 1
rlabel polysilicon 23 -1073 23 -1073 0 3
rlabel polysilicon 33 -1067 33 -1067 0 2
rlabel polysilicon 37 -1067 37 -1067 0 1
rlabel polysilicon 37 -1073 37 -1073 0 3
rlabel polysilicon 44 -1067 44 -1067 0 1
rlabel polysilicon 44 -1073 44 -1073 0 3
rlabel polysilicon 51 -1067 51 -1067 0 1
rlabel polysilicon 51 -1073 51 -1073 0 3
rlabel polysilicon 61 -1067 61 -1067 0 2
rlabel polysilicon 65 -1067 65 -1067 0 1
rlabel polysilicon 65 -1073 65 -1073 0 3
rlabel polysilicon 75 -1067 75 -1067 0 2
rlabel polysilicon 79 -1067 79 -1067 0 1
rlabel polysilicon 79 -1073 79 -1073 0 3
rlabel polysilicon 86 -1067 86 -1067 0 1
rlabel polysilicon 93 -1067 93 -1067 0 1
rlabel polysilicon 93 -1073 93 -1073 0 3
rlabel polysilicon 103 -1067 103 -1067 0 2
rlabel polysilicon 107 -1067 107 -1067 0 1
rlabel polysilicon 114 -1067 114 -1067 0 1
rlabel polysilicon 114 -1073 114 -1073 0 3
rlabel polysilicon 121 -1067 121 -1067 0 1
rlabel polysilicon 121 -1073 121 -1073 0 3
rlabel polysilicon 128 -1067 128 -1067 0 1
rlabel polysilicon 128 -1073 128 -1073 0 3
rlabel polysilicon 135 -1067 135 -1067 0 1
rlabel polysilicon 135 -1073 135 -1073 0 3
rlabel polysilicon 142 -1067 142 -1067 0 1
rlabel polysilicon 142 -1073 142 -1073 0 3
rlabel polysilicon 149 -1067 149 -1067 0 1
rlabel polysilicon 152 -1067 152 -1067 0 2
rlabel polysilicon 149 -1073 149 -1073 0 3
rlabel polysilicon 156 -1067 156 -1067 0 1
rlabel polysilicon 156 -1073 156 -1073 0 3
rlabel polysilicon 163 -1067 163 -1067 0 1
rlabel polysilicon 166 -1067 166 -1067 0 2
rlabel polysilicon 166 -1073 166 -1073 0 4
rlabel polysilicon 170 -1067 170 -1067 0 1
rlabel polysilicon 170 -1073 170 -1073 0 3
rlabel polysilicon 177 -1067 177 -1067 0 1
rlabel polysilicon 180 -1067 180 -1067 0 2
rlabel polysilicon 177 -1073 177 -1073 0 3
rlabel polysilicon 184 -1067 184 -1067 0 1
rlabel polysilicon 184 -1073 184 -1073 0 3
rlabel polysilicon 191 -1067 191 -1067 0 1
rlabel polysilicon 194 -1067 194 -1067 0 2
rlabel polysilicon 194 -1073 194 -1073 0 4
rlabel polysilicon 198 -1073 198 -1073 0 3
rlabel polysilicon 201 -1073 201 -1073 0 4
rlabel polysilicon 205 -1067 205 -1067 0 1
rlabel polysilicon 205 -1073 205 -1073 0 3
rlabel polysilicon 212 -1067 212 -1067 0 1
rlabel polysilicon 212 -1073 212 -1073 0 3
rlabel polysilicon 219 -1067 219 -1067 0 1
rlabel polysilicon 219 -1073 219 -1073 0 3
rlabel polysilicon 226 -1067 226 -1067 0 1
rlabel polysilicon 226 -1073 226 -1073 0 3
rlabel polysilicon 233 -1067 233 -1067 0 1
rlabel polysilicon 233 -1073 233 -1073 0 3
rlabel polysilicon 243 -1067 243 -1067 0 2
rlabel polysilicon 243 -1073 243 -1073 0 4
rlabel polysilicon 250 -1067 250 -1067 0 2
rlabel polysilicon 254 -1067 254 -1067 0 1
rlabel polysilicon 254 -1073 254 -1073 0 3
rlabel polysilicon 261 -1067 261 -1067 0 1
rlabel polysilicon 261 -1073 261 -1073 0 3
rlabel polysilicon 268 -1067 268 -1067 0 1
rlabel polysilicon 268 -1073 268 -1073 0 3
rlabel polysilicon 278 -1067 278 -1067 0 2
rlabel polysilicon 278 -1073 278 -1073 0 4
rlabel polysilicon 282 -1067 282 -1067 0 1
rlabel polysilicon 282 -1073 282 -1073 0 3
rlabel polysilicon 289 -1067 289 -1067 0 1
rlabel polysilicon 289 -1073 289 -1073 0 3
rlabel polysilicon 296 -1067 296 -1067 0 1
rlabel polysilicon 296 -1073 296 -1073 0 3
rlabel polysilicon 303 -1067 303 -1067 0 1
rlabel polysilicon 303 -1073 303 -1073 0 3
rlabel polysilicon 310 -1067 310 -1067 0 1
rlabel polysilicon 313 -1067 313 -1067 0 2
rlabel polysilicon 310 -1073 310 -1073 0 3
rlabel polysilicon 317 -1067 317 -1067 0 1
rlabel polysilicon 317 -1073 317 -1073 0 3
rlabel polysilicon 324 -1067 324 -1067 0 1
rlabel polysilicon 324 -1073 324 -1073 0 3
rlabel polysilicon 334 -1067 334 -1067 0 2
rlabel polysilicon 331 -1073 331 -1073 0 3
rlabel polysilicon 334 -1073 334 -1073 0 4
rlabel polysilicon 338 -1067 338 -1067 0 1
rlabel polysilicon 338 -1073 338 -1073 0 3
rlabel polysilicon 345 -1067 345 -1067 0 1
rlabel polysilicon 345 -1073 345 -1073 0 3
rlabel polysilicon 352 -1067 352 -1067 0 1
rlabel polysilicon 352 -1073 352 -1073 0 3
rlabel polysilicon 359 -1067 359 -1067 0 1
rlabel polysilicon 359 -1073 359 -1073 0 3
rlabel polysilicon 366 -1067 366 -1067 0 1
rlabel polysilicon 366 -1073 366 -1073 0 3
rlabel polysilicon 373 -1067 373 -1067 0 1
rlabel polysilicon 373 -1073 373 -1073 0 3
rlabel polysilicon 380 -1067 380 -1067 0 1
rlabel polysilicon 380 -1073 380 -1073 0 3
rlabel polysilicon 387 -1067 387 -1067 0 1
rlabel polysilicon 387 -1073 387 -1073 0 3
rlabel polysilicon 394 -1067 394 -1067 0 1
rlabel polysilicon 394 -1073 394 -1073 0 3
rlabel polysilicon 401 -1067 401 -1067 0 1
rlabel polysilicon 404 -1067 404 -1067 0 2
rlabel polysilicon 401 -1073 401 -1073 0 3
rlabel polysilicon 408 -1067 408 -1067 0 1
rlabel polysilicon 411 -1067 411 -1067 0 2
rlabel polysilicon 411 -1073 411 -1073 0 4
rlabel polysilicon 418 -1067 418 -1067 0 2
rlabel polysilicon 415 -1073 415 -1073 0 3
rlabel polysilicon 418 -1073 418 -1073 0 4
rlabel polysilicon 425 -1067 425 -1067 0 2
rlabel polysilicon 422 -1073 422 -1073 0 3
rlabel polysilicon 425 -1073 425 -1073 0 4
rlabel polysilicon 429 -1067 429 -1067 0 1
rlabel polysilicon 429 -1073 429 -1073 0 3
rlabel polysilicon 439 -1067 439 -1067 0 2
rlabel polysilicon 439 -1073 439 -1073 0 4
rlabel polysilicon 443 -1067 443 -1067 0 1
rlabel polysilicon 443 -1073 443 -1073 0 3
rlabel polysilicon 450 -1067 450 -1067 0 1
rlabel polysilicon 450 -1073 450 -1073 0 3
rlabel polysilicon 453 -1073 453 -1073 0 4
rlabel polysilicon 457 -1067 457 -1067 0 1
rlabel polysilicon 457 -1073 457 -1073 0 3
rlabel polysilicon 464 -1067 464 -1067 0 1
rlabel polysilicon 464 -1073 464 -1073 0 3
rlabel polysilicon 474 -1073 474 -1073 0 4
rlabel polysilicon 478 -1067 478 -1067 0 1
rlabel polysilicon 478 -1073 478 -1073 0 3
rlabel polysilicon 481 -1073 481 -1073 0 4
rlabel polysilicon 485 -1067 485 -1067 0 1
rlabel polysilicon 485 -1073 485 -1073 0 3
rlabel polysilicon 492 -1067 492 -1067 0 1
rlabel polysilicon 495 -1067 495 -1067 0 2
rlabel polysilicon 492 -1073 492 -1073 0 3
rlabel polysilicon 495 -1073 495 -1073 0 4
rlabel polysilicon 499 -1067 499 -1067 0 1
rlabel polysilicon 499 -1073 499 -1073 0 3
rlabel polysilicon 506 -1073 506 -1073 0 3
rlabel polysilicon 513 -1067 513 -1067 0 1
rlabel polysilicon 513 -1073 513 -1073 0 3
rlabel polysilicon 520 -1067 520 -1067 0 1
rlabel polysilicon 523 -1073 523 -1073 0 4
rlabel polysilicon 527 -1067 527 -1067 0 1
rlabel polysilicon 527 -1073 527 -1073 0 3
rlabel polysilicon 534 -1073 534 -1073 0 3
rlabel polysilicon 537 -1073 537 -1073 0 4
rlabel polysilicon 541 -1067 541 -1067 0 1
rlabel polysilicon 541 -1073 541 -1073 0 3
rlabel polysilicon 548 -1067 548 -1067 0 1
rlabel polysilicon 548 -1073 548 -1073 0 3
rlabel polysilicon 555 -1067 555 -1067 0 1
rlabel polysilicon 555 -1073 555 -1073 0 3
rlabel polysilicon 562 -1073 562 -1073 0 3
rlabel polysilicon 565 -1073 565 -1073 0 4
rlabel polysilicon 569 -1067 569 -1067 0 1
rlabel polysilicon 569 -1073 569 -1073 0 3
rlabel polysilicon 576 -1067 576 -1067 0 1
rlabel polysilicon 576 -1073 576 -1073 0 3
rlabel polysilicon 583 -1067 583 -1067 0 1
rlabel polysilicon 583 -1073 583 -1073 0 3
rlabel polysilicon 590 -1067 590 -1067 0 1
rlabel polysilicon 590 -1073 590 -1073 0 3
rlabel polysilicon 597 -1067 597 -1067 0 1
rlabel polysilicon 597 -1073 597 -1073 0 3
rlabel polysilicon 604 -1067 604 -1067 0 1
rlabel polysilicon 604 -1073 604 -1073 0 3
rlabel polysilicon 611 -1067 611 -1067 0 1
rlabel polysilicon 611 -1073 611 -1073 0 3
rlabel polysilicon 618 -1067 618 -1067 0 1
rlabel polysilicon 618 -1073 618 -1073 0 3
rlabel polysilicon 625 -1067 625 -1067 0 1
rlabel polysilicon 625 -1073 625 -1073 0 3
rlabel polysilicon 632 -1067 632 -1067 0 1
rlabel polysilicon 632 -1073 632 -1073 0 3
rlabel polysilicon 639 -1067 639 -1067 0 1
rlabel polysilicon 639 -1073 639 -1073 0 3
rlabel polysilicon 646 -1067 646 -1067 0 1
rlabel polysilicon 646 -1073 646 -1073 0 3
rlabel polysilicon 653 -1067 653 -1067 0 1
rlabel polysilicon 653 -1073 653 -1073 0 3
rlabel polysilicon 660 -1067 660 -1067 0 1
rlabel polysilicon 660 -1073 660 -1073 0 3
rlabel polysilicon 667 -1067 667 -1067 0 1
rlabel polysilicon 667 -1073 667 -1073 0 3
rlabel polysilicon 674 -1067 674 -1067 0 1
rlabel polysilicon 674 -1073 674 -1073 0 3
rlabel polysilicon 681 -1067 681 -1067 0 1
rlabel polysilicon 681 -1073 681 -1073 0 3
rlabel polysilicon 688 -1067 688 -1067 0 1
rlabel polysilicon 691 -1067 691 -1067 0 2
rlabel polysilicon 691 -1073 691 -1073 0 4
rlabel polysilicon 695 -1067 695 -1067 0 1
rlabel polysilicon 695 -1073 695 -1073 0 3
rlabel polysilicon 702 -1067 702 -1067 0 1
rlabel polysilicon 702 -1073 702 -1073 0 3
rlabel polysilicon 709 -1067 709 -1067 0 1
rlabel polysilicon 709 -1073 709 -1073 0 3
rlabel polysilicon 716 -1067 716 -1067 0 1
rlabel polysilicon 719 -1067 719 -1067 0 2
rlabel polysilicon 716 -1073 716 -1073 0 3
rlabel polysilicon 723 -1067 723 -1067 0 1
rlabel polysilicon 723 -1073 723 -1073 0 3
rlabel polysilicon 730 -1067 730 -1067 0 1
rlabel polysilicon 730 -1073 730 -1073 0 3
rlabel polysilicon 737 -1067 737 -1067 0 1
rlabel polysilicon 737 -1073 737 -1073 0 3
rlabel polysilicon 9 -1128 9 -1128 0 1
rlabel polysilicon 9 -1134 9 -1134 0 3
rlabel polysilicon 16 -1128 16 -1128 0 1
rlabel polysilicon 16 -1134 16 -1134 0 3
rlabel polysilicon 23 -1128 23 -1128 0 1
rlabel polysilicon 23 -1134 23 -1134 0 3
rlabel polysilicon 30 -1128 30 -1128 0 1
rlabel polysilicon 37 -1128 37 -1128 0 1
rlabel polysilicon 37 -1134 37 -1134 0 3
rlabel polysilicon 44 -1134 44 -1134 0 3
rlabel polysilicon 47 -1134 47 -1134 0 4
rlabel polysilicon 51 -1128 51 -1128 0 1
rlabel polysilicon 51 -1134 51 -1134 0 3
rlabel polysilicon 58 -1128 58 -1128 0 1
rlabel polysilicon 58 -1134 58 -1134 0 3
rlabel polysilicon 65 -1128 65 -1128 0 1
rlabel polysilicon 68 -1128 68 -1128 0 2
rlabel polysilicon 72 -1128 72 -1128 0 1
rlabel polysilicon 72 -1134 72 -1134 0 3
rlabel polysilicon 82 -1128 82 -1128 0 2
rlabel polysilicon 82 -1134 82 -1134 0 4
rlabel polysilicon 86 -1128 86 -1128 0 1
rlabel polysilicon 86 -1134 86 -1134 0 3
rlabel polysilicon 93 -1128 93 -1128 0 1
rlabel polysilicon 93 -1134 93 -1134 0 3
rlabel polysilicon 100 -1128 100 -1128 0 1
rlabel polysilicon 100 -1134 100 -1134 0 3
rlabel polysilicon 107 -1128 107 -1128 0 1
rlabel polysilicon 107 -1134 107 -1134 0 3
rlabel polysilicon 114 -1128 114 -1128 0 1
rlabel polysilicon 114 -1134 114 -1134 0 3
rlabel polysilicon 124 -1128 124 -1128 0 2
rlabel polysilicon 121 -1134 121 -1134 0 3
rlabel polysilicon 128 -1128 128 -1128 0 1
rlabel polysilicon 128 -1134 128 -1134 0 3
rlabel polysilicon 135 -1128 135 -1128 0 1
rlabel polysilicon 135 -1134 135 -1134 0 3
rlabel polysilicon 142 -1128 142 -1128 0 1
rlabel polysilicon 145 -1128 145 -1128 0 2
rlabel polysilicon 142 -1134 142 -1134 0 3
rlabel polysilicon 145 -1134 145 -1134 0 4
rlabel polysilicon 149 -1128 149 -1128 0 1
rlabel polysilicon 149 -1134 149 -1134 0 3
rlabel polysilicon 159 -1128 159 -1128 0 2
rlabel polysilicon 156 -1134 156 -1134 0 3
rlabel polysilicon 163 -1134 163 -1134 0 3
rlabel polysilicon 166 -1134 166 -1134 0 4
rlabel polysilicon 170 -1134 170 -1134 0 3
rlabel polysilicon 173 -1134 173 -1134 0 4
rlabel polysilicon 177 -1128 177 -1128 0 1
rlabel polysilicon 180 -1128 180 -1128 0 2
rlabel polysilicon 180 -1134 180 -1134 0 4
rlabel polysilicon 184 -1128 184 -1128 0 1
rlabel polysilicon 187 -1128 187 -1128 0 2
rlabel polysilicon 184 -1134 184 -1134 0 3
rlabel polysilicon 191 -1134 191 -1134 0 3
rlabel polysilicon 194 -1134 194 -1134 0 4
rlabel polysilicon 198 -1128 198 -1128 0 1
rlabel polysilicon 198 -1134 198 -1134 0 3
rlabel polysilicon 205 -1128 205 -1128 0 1
rlabel polysilicon 205 -1134 205 -1134 0 3
rlabel polysilicon 215 -1128 215 -1128 0 2
rlabel polysilicon 215 -1134 215 -1134 0 4
rlabel polysilicon 219 -1128 219 -1128 0 1
rlabel polysilicon 219 -1134 219 -1134 0 3
rlabel polysilicon 226 -1128 226 -1128 0 1
rlabel polysilicon 226 -1134 226 -1134 0 3
rlabel polysilicon 233 -1128 233 -1128 0 1
rlabel polysilicon 233 -1134 233 -1134 0 3
rlabel polysilicon 240 -1128 240 -1128 0 1
rlabel polysilicon 247 -1128 247 -1128 0 1
rlabel polysilicon 247 -1134 247 -1134 0 3
rlabel polysilicon 250 -1134 250 -1134 0 4
rlabel polysilicon 254 -1128 254 -1128 0 1
rlabel polysilicon 254 -1134 254 -1134 0 3
rlabel polysilicon 261 -1128 261 -1128 0 1
rlabel polysilicon 261 -1134 261 -1134 0 3
rlabel polysilicon 268 -1128 268 -1128 0 1
rlabel polysilicon 268 -1134 268 -1134 0 3
rlabel polysilicon 275 -1128 275 -1128 0 1
rlabel polysilicon 278 -1128 278 -1128 0 2
rlabel polysilicon 275 -1134 275 -1134 0 3
rlabel polysilicon 278 -1134 278 -1134 0 4
rlabel polysilicon 282 -1128 282 -1128 0 1
rlabel polysilicon 282 -1134 282 -1134 0 3
rlabel polysilicon 289 -1128 289 -1128 0 1
rlabel polysilicon 289 -1134 289 -1134 0 3
rlabel polysilicon 296 -1128 296 -1128 0 1
rlabel polysilicon 296 -1134 296 -1134 0 3
rlabel polysilicon 303 -1128 303 -1128 0 1
rlabel polysilicon 303 -1134 303 -1134 0 3
rlabel polysilicon 310 -1128 310 -1128 0 1
rlabel polysilicon 313 -1128 313 -1128 0 2
rlabel polysilicon 310 -1134 310 -1134 0 3
rlabel polysilicon 317 -1128 317 -1128 0 1
rlabel polysilicon 317 -1134 317 -1134 0 3
rlabel polysilicon 324 -1128 324 -1128 0 1
rlabel polysilicon 324 -1134 324 -1134 0 3
rlabel polysilicon 331 -1134 331 -1134 0 3
rlabel polysilicon 334 -1134 334 -1134 0 4
rlabel polysilicon 338 -1128 338 -1128 0 1
rlabel polysilicon 338 -1134 338 -1134 0 3
rlabel polysilicon 348 -1128 348 -1128 0 2
rlabel polysilicon 345 -1134 345 -1134 0 3
rlabel polysilicon 348 -1134 348 -1134 0 4
rlabel polysilicon 352 -1128 352 -1128 0 1
rlabel polysilicon 352 -1134 352 -1134 0 3
rlabel polysilicon 362 -1128 362 -1128 0 2
rlabel polysilicon 362 -1134 362 -1134 0 4
rlabel polysilicon 366 -1134 366 -1134 0 3
rlabel polysilicon 369 -1134 369 -1134 0 4
rlabel polysilicon 376 -1128 376 -1128 0 2
rlabel polysilicon 373 -1134 373 -1134 0 3
rlabel polysilicon 380 -1128 380 -1128 0 1
rlabel polysilicon 383 -1128 383 -1128 0 2
rlabel polysilicon 387 -1128 387 -1128 0 1
rlabel polysilicon 387 -1134 387 -1134 0 3
rlabel polysilicon 390 -1134 390 -1134 0 4
rlabel polysilicon 397 -1128 397 -1128 0 2
rlabel polysilicon 394 -1134 394 -1134 0 3
rlabel polysilicon 397 -1134 397 -1134 0 4
rlabel polysilicon 401 -1128 401 -1128 0 1
rlabel polysilicon 401 -1134 401 -1134 0 3
rlabel polysilicon 408 -1128 408 -1128 0 1
rlabel polysilicon 408 -1134 408 -1134 0 3
rlabel polysilicon 415 -1128 415 -1128 0 1
rlabel polysilicon 415 -1134 415 -1134 0 3
rlabel polysilicon 422 -1128 422 -1128 0 1
rlabel polysilicon 425 -1128 425 -1128 0 2
rlabel polysilicon 422 -1134 422 -1134 0 3
rlabel polysilicon 429 -1128 429 -1128 0 1
rlabel polysilicon 429 -1134 429 -1134 0 3
rlabel polysilicon 432 -1134 432 -1134 0 4
rlabel polysilicon 436 -1128 436 -1128 0 1
rlabel polysilicon 436 -1134 436 -1134 0 3
rlabel polysilicon 443 -1128 443 -1128 0 1
rlabel polysilicon 443 -1134 443 -1134 0 3
rlabel polysilicon 450 -1128 450 -1128 0 1
rlabel polysilicon 450 -1134 450 -1134 0 3
rlabel polysilicon 457 -1128 457 -1128 0 1
rlabel polysilicon 457 -1134 457 -1134 0 3
rlabel polysilicon 464 -1128 464 -1128 0 1
rlabel polysilicon 464 -1134 464 -1134 0 3
rlabel polysilicon 471 -1128 471 -1128 0 1
rlabel polysilicon 471 -1134 471 -1134 0 3
rlabel polysilicon 478 -1128 478 -1128 0 1
rlabel polysilicon 478 -1134 478 -1134 0 3
rlabel polysilicon 485 -1128 485 -1128 0 1
rlabel polysilicon 485 -1134 485 -1134 0 3
rlabel polysilicon 492 -1128 492 -1128 0 1
rlabel polysilicon 492 -1134 492 -1134 0 3
rlabel polysilicon 499 -1128 499 -1128 0 1
rlabel polysilicon 499 -1134 499 -1134 0 3
rlabel polysilicon 506 -1128 506 -1128 0 1
rlabel polysilicon 506 -1134 506 -1134 0 3
rlabel polysilicon 513 -1128 513 -1128 0 1
rlabel polysilicon 513 -1134 513 -1134 0 3
rlabel polysilicon 523 -1128 523 -1128 0 2
rlabel polysilicon 523 -1134 523 -1134 0 4
rlabel polysilicon 527 -1128 527 -1128 0 1
rlabel polysilicon 527 -1134 527 -1134 0 3
rlabel polysilicon 534 -1128 534 -1128 0 1
rlabel polysilicon 534 -1134 534 -1134 0 3
rlabel polysilicon 541 -1128 541 -1128 0 1
rlabel polysilicon 541 -1134 541 -1134 0 3
rlabel polysilicon 548 -1128 548 -1128 0 1
rlabel polysilicon 548 -1134 548 -1134 0 3
rlabel polysilicon 555 -1128 555 -1128 0 1
rlabel polysilicon 555 -1134 555 -1134 0 3
rlabel polysilicon 562 -1128 562 -1128 0 1
rlabel polysilicon 562 -1134 562 -1134 0 3
rlabel polysilicon 569 -1128 569 -1128 0 1
rlabel polysilicon 569 -1134 569 -1134 0 3
rlabel polysilicon 576 -1128 576 -1128 0 1
rlabel polysilicon 576 -1134 576 -1134 0 3
rlabel polysilicon 583 -1128 583 -1128 0 1
rlabel polysilicon 583 -1134 583 -1134 0 3
rlabel polysilicon 590 -1128 590 -1128 0 1
rlabel polysilicon 590 -1134 590 -1134 0 3
rlabel polysilicon 597 -1128 597 -1128 0 1
rlabel polysilicon 597 -1134 597 -1134 0 3
rlabel polysilicon 604 -1128 604 -1128 0 1
rlabel polysilicon 604 -1134 604 -1134 0 3
rlabel polysilicon 611 -1128 611 -1128 0 1
rlabel polysilicon 611 -1134 611 -1134 0 3
rlabel polysilicon 618 -1128 618 -1128 0 1
rlabel polysilicon 618 -1134 618 -1134 0 3
rlabel polysilicon 625 -1128 625 -1128 0 1
rlabel polysilicon 625 -1134 625 -1134 0 3
rlabel polysilicon 632 -1128 632 -1128 0 1
rlabel polysilicon 632 -1134 632 -1134 0 3
rlabel polysilicon 639 -1128 639 -1128 0 1
rlabel polysilicon 639 -1134 639 -1134 0 3
rlabel polysilicon 646 -1128 646 -1128 0 1
rlabel polysilicon 646 -1134 646 -1134 0 3
rlabel polysilicon 653 -1128 653 -1128 0 1
rlabel polysilicon 653 -1134 653 -1134 0 3
rlabel polysilicon 660 -1128 660 -1128 0 1
rlabel polysilicon 660 -1134 660 -1134 0 3
rlabel polysilicon 667 -1128 667 -1128 0 1
rlabel polysilicon 667 -1134 667 -1134 0 3
rlabel polysilicon 674 -1128 674 -1128 0 1
rlabel polysilicon 677 -1128 677 -1128 0 2
rlabel polysilicon 674 -1134 674 -1134 0 3
rlabel polysilicon 677 -1134 677 -1134 0 4
rlabel polysilicon 681 -1128 681 -1128 0 1
rlabel polysilicon 684 -1128 684 -1128 0 2
rlabel polysilicon 688 -1128 688 -1128 0 1
rlabel polysilicon 688 -1134 688 -1134 0 3
rlabel polysilicon 695 -1128 695 -1128 0 1
rlabel polysilicon 695 -1134 695 -1134 0 3
rlabel polysilicon 702 -1128 702 -1128 0 1
rlabel polysilicon 702 -1134 702 -1134 0 3
rlabel polysilicon 709 -1128 709 -1128 0 1
rlabel polysilicon 709 -1134 709 -1134 0 3
rlabel polysilicon 2 -1185 2 -1185 0 1
rlabel polysilicon 2 -1191 2 -1191 0 3
rlabel polysilicon 9 -1185 9 -1185 0 1
rlabel polysilicon 9 -1191 9 -1191 0 3
rlabel polysilicon 19 -1185 19 -1185 0 2
rlabel polysilicon 23 -1191 23 -1191 0 3
rlabel polysilicon 30 -1185 30 -1185 0 1
rlabel polysilicon 30 -1191 30 -1191 0 3
rlabel polysilicon 37 -1185 37 -1185 0 1
rlabel polysilicon 37 -1191 37 -1191 0 3
rlabel polysilicon 44 -1185 44 -1185 0 1
rlabel polysilicon 44 -1191 44 -1191 0 3
rlabel polysilicon 51 -1185 51 -1185 0 1
rlabel polysilicon 51 -1191 51 -1191 0 3
rlabel polysilicon 58 -1185 58 -1185 0 1
rlabel polysilicon 58 -1191 58 -1191 0 3
rlabel polysilicon 65 -1185 65 -1185 0 1
rlabel polysilicon 75 -1185 75 -1185 0 2
rlabel polysilicon 72 -1191 72 -1191 0 3
rlabel polysilicon 75 -1191 75 -1191 0 4
rlabel polysilicon 79 -1185 79 -1185 0 1
rlabel polysilicon 79 -1191 79 -1191 0 3
rlabel polysilicon 86 -1185 86 -1185 0 1
rlabel polysilicon 89 -1191 89 -1191 0 4
rlabel polysilicon 93 -1185 93 -1185 0 1
rlabel polysilicon 93 -1191 93 -1191 0 3
rlabel polysilicon 100 -1191 100 -1191 0 3
rlabel polysilicon 107 -1185 107 -1185 0 1
rlabel polysilicon 110 -1185 110 -1185 0 2
rlabel polysilicon 107 -1191 107 -1191 0 3
rlabel polysilicon 114 -1185 114 -1185 0 1
rlabel polysilicon 117 -1191 117 -1191 0 4
rlabel polysilicon 121 -1185 121 -1185 0 1
rlabel polysilicon 121 -1191 121 -1191 0 3
rlabel polysilicon 128 -1185 128 -1185 0 1
rlabel polysilicon 128 -1191 128 -1191 0 3
rlabel polysilicon 135 -1185 135 -1185 0 1
rlabel polysilicon 135 -1191 135 -1191 0 3
rlabel polysilicon 142 -1185 142 -1185 0 1
rlabel polysilicon 145 -1185 145 -1185 0 2
rlabel polysilicon 145 -1191 145 -1191 0 4
rlabel polysilicon 149 -1185 149 -1185 0 1
rlabel polysilicon 152 -1185 152 -1185 0 2
rlabel polysilicon 149 -1191 149 -1191 0 3
rlabel polysilicon 152 -1191 152 -1191 0 4
rlabel polysilicon 156 -1185 156 -1185 0 1
rlabel polysilicon 159 -1185 159 -1185 0 2
rlabel polysilicon 163 -1185 163 -1185 0 1
rlabel polysilicon 163 -1191 163 -1191 0 3
rlabel polysilicon 170 -1185 170 -1185 0 1
rlabel polysilicon 170 -1191 170 -1191 0 3
rlabel polysilicon 173 -1191 173 -1191 0 4
rlabel polysilicon 177 -1185 177 -1185 0 1
rlabel polysilicon 177 -1191 177 -1191 0 3
rlabel polysilicon 184 -1185 184 -1185 0 1
rlabel polysilicon 184 -1191 184 -1191 0 3
rlabel polysilicon 194 -1185 194 -1185 0 2
rlabel polysilicon 191 -1191 191 -1191 0 3
rlabel polysilicon 198 -1185 198 -1185 0 1
rlabel polysilicon 198 -1191 198 -1191 0 3
rlabel polysilicon 205 -1185 205 -1185 0 1
rlabel polysilicon 208 -1185 208 -1185 0 2
rlabel polysilicon 215 -1191 215 -1191 0 4
rlabel polysilicon 219 -1185 219 -1185 0 1
rlabel polysilicon 219 -1191 219 -1191 0 3
rlabel polysilicon 226 -1185 226 -1185 0 1
rlabel polysilicon 226 -1191 226 -1191 0 3
rlabel polysilicon 233 -1185 233 -1185 0 1
rlabel polysilicon 236 -1185 236 -1185 0 2
rlabel polysilicon 240 -1185 240 -1185 0 1
rlabel polysilicon 240 -1191 240 -1191 0 3
rlabel polysilicon 247 -1185 247 -1185 0 1
rlabel polysilicon 247 -1191 247 -1191 0 3
rlabel polysilicon 254 -1185 254 -1185 0 1
rlabel polysilicon 254 -1191 254 -1191 0 3
rlabel polysilicon 261 -1185 261 -1185 0 1
rlabel polysilicon 261 -1191 261 -1191 0 3
rlabel polysilicon 268 -1185 268 -1185 0 1
rlabel polysilicon 268 -1191 268 -1191 0 3
rlabel polysilicon 275 -1191 275 -1191 0 3
rlabel polysilicon 282 -1185 282 -1185 0 1
rlabel polysilicon 282 -1191 282 -1191 0 3
rlabel polysilicon 289 -1185 289 -1185 0 1
rlabel polysilicon 289 -1191 289 -1191 0 3
rlabel polysilicon 296 -1185 296 -1185 0 1
rlabel polysilicon 296 -1191 296 -1191 0 3
rlabel polysilicon 303 -1185 303 -1185 0 1
rlabel polysilicon 303 -1191 303 -1191 0 3
rlabel polysilicon 306 -1191 306 -1191 0 4
rlabel polysilicon 310 -1185 310 -1185 0 1
rlabel polysilicon 310 -1191 310 -1191 0 3
rlabel polysilicon 317 -1185 317 -1185 0 1
rlabel polysilicon 320 -1185 320 -1185 0 2
rlabel polysilicon 320 -1191 320 -1191 0 4
rlabel polysilicon 324 -1185 324 -1185 0 1
rlabel polysilicon 327 -1191 327 -1191 0 4
rlabel polysilicon 331 -1185 331 -1185 0 1
rlabel polysilicon 334 -1191 334 -1191 0 4
rlabel polysilicon 338 -1185 338 -1185 0 1
rlabel polysilicon 341 -1191 341 -1191 0 4
rlabel polysilicon 348 -1185 348 -1185 0 2
rlabel polysilicon 345 -1191 345 -1191 0 3
rlabel polysilicon 348 -1191 348 -1191 0 4
rlabel polysilicon 352 -1185 352 -1185 0 1
rlabel polysilicon 352 -1191 352 -1191 0 3
rlabel polysilicon 359 -1185 359 -1185 0 1
rlabel polysilicon 359 -1191 359 -1191 0 3
rlabel polysilicon 366 -1185 366 -1185 0 1
rlabel polysilicon 366 -1191 366 -1191 0 3
rlabel polysilicon 373 -1185 373 -1185 0 1
rlabel polysilicon 373 -1191 373 -1191 0 3
rlabel polysilicon 380 -1185 380 -1185 0 1
rlabel polysilicon 380 -1191 380 -1191 0 3
rlabel polysilicon 387 -1185 387 -1185 0 1
rlabel polysilicon 390 -1185 390 -1185 0 2
rlabel polysilicon 387 -1191 387 -1191 0 3
rlabel polysilicon 390 -1191 390 -1191 0 4
rlabel polysilicon 394 -1185 394 -1185 0 1
rlabel polysilicon 394 -1191 394 -1191 0 3
rlabel polysilicon 401 -1185 401 -1185 0 1
rlabel polysilicon 401 -1191 401 -1191 0 3
rlabel polysilicon 408 -1185 408 -1185 0 1
rlabel polysilicon 408 -1191 408 -1191 0 3
rlabel polysilicon 415 -1185 415 -1185 0 1
rlabel polysilicon 415 -1191 415 -1191 0 3
rlabel polysilicon 422 -1185 422 -1185 0 1
rlabel polysilicon 422 -1191 422 -1191 0 3
rlabel polysilicon 429 -1185 429 -1185 0 1
rlabel polysilicon 429 -1191 429 -1191 0 3
rlabel polysilicon 436 -1191 436 -1191 0 3
rlabel polysilicon 443 -1185 443 -1185 0 1
rlabel polysilicon 446 -1185 446 -1185 0 2
rlabel polysilicon 443 -1191 443 -1191 0 3
rlabel polysilicon 446 -1191 446 -1191 0 4
rlabel polysilicon 450 -1185 450 -1185 0 1
rlabel polysilicon 450 -1191 450 -1191 0 3
rlabel polysilicon 453 -1191 453 -1191 0 4
rlabel polysilicon 457 -1185 457 -1185 0 1
rlabel polysilicon 457 -1191 457 -1191 0 3
rlabel polysilicon 464 -1185 464 -1185 0 1
rlabel polysilicon 467 -1191 467 -1191 0 4
rlabel polysilicon 471 -1185 471 -1185 0 1
rlabel polysilicon 471 -1191 471 -1191 0 3
rlabel polysilicon 478 -1185 478 -1185 0 1
rlabel polysilicon 478 -1191 478 -1191 0 3
rlabel polysilicon 485 -1185 485 -1185 0 1
rlabel polysilicon 485 -1191 485 -1191 0 3
rlabel polysilicon 492 -1185 492 -1185 0 1
rlabel polysilicon 492 -1191 492 -1191 0 3
rlabel polysilicon 499 -1185 499 -1185 0 1
rlabel polysilicon 499 -1191 499 -1191 0 3
rlabel polysilicon 506 -1185 506 -1185 0 1
rlabel polysilicon 506 -1191 506 -1191 0 3
rlabel polysilicon 513 -1185 513 -1185 0 1
rlabel polysilicon 513 -1191 513 -1191 0 3
rlabel polysilicon 520 -1185 520 -1185 0 1
rlabel polysilicon 520 -1191 520 -1191 0 3
rlabel polysilicon 530 -1185 530 -1185 0 2
rlabel polysilicon 530 -1191 530 -1191 0 4
rlabel polysilicon 534 -1185 534 -1185 0 1
rlabel polysilicon 534 -1191 534 -1191 0 3
rlabel polysilicon 544 -1185 544 -1185 0 2
rlabel polysilicon 541 -1191 541 -1191 0 3
rlabel polysilicon 548 -1185 548 -1185 0 1
rlabel polysilicon 548 -1191 548 -1191 0 3
rlabel polysilicon 555 -1185 555 -1185 0 1
rlabel polysilicon 555 -1191 555 -1191 0 3
rlabel polysilicon 562 -1185 562 -1185 0 1
rlabel polysilicon 562 -1191 562 -1191 0 3
rlabel polysilicon 569 -1185 569 -1185 0 1
rlabel polysilicon 569 -1191 569 -1191 0 3
rlabel polysilicon 576 -1185 576 -1185 0 1
rlabel polysilicon 576 -1191 576 -1191 0 3
rlabel polysilicon 583 -1185 583 -1185 0 1
rlabel polysilicon 583 -1191 583 -1191 0 3
rlabel polysilicon 590 -1185 590 -1185 0 1
rlabel polysilicon 590 -1191 590 -1191 0 3
rlabel polysilicon 597 -1185 597 -1185 0 1
rlabel polysilicon 597 -1191 597 -1191 0 3
rlabel polysilicon 604 -1185 604 -1185 0 1
rlabel polysilicon 604 -1191 604 -1191 0 3
rlabel polysilicon 611 -1185 611 -1185 0 1
rlabel polysilicon 611 -1191 611 -1191 0 3
rlabel polysilicon 618 -1185 618 -1185 0 1
rlabel polysilicon 618 -1191 618 -1191 0 3
rlabel polysilicon 625 -1185 625 -1185 0 1
rlabel polysilicon 625 -1191 625 -1191 0 3
rlabel polysilicon 632 -1185 632 -1185 0 1
rlabel polysilicon 632 -1191 632 -1191 0 3
rlabel polysilicon 639 -1185 639 -1185 0 1
rlabel polysilicon 639 -1191 639 -1191 0 3
rlabel polysilicon 646 -1185 646 -1185 0 1
rlabel polysilicon 646 -1191 646 -1191 0 3
rlabel polysilicon 656 -1185 656 -1185 0 2
rlabel polysilicon 660 -1185 660 -1185 0 1
rlabel polysilicon 660 -1191 660 -1191 0 3
rlabel polysilicon 667 -1185 667 -1185 0 1
rlabel polysilicon 674 -1185 674 -1185 0 1
rlabel polysilicon 677 -1185 677 -1185 0 2
rlabel polysilicon 674 -1191 674 -1191 0 3
rlabel polysilicon 681 -1185 681 -1185 0 1
rlabel polysilicon 681 -1191 681 -1191 0 3
rlabel polysilicon 688 -1185 688 -1185 0 1
rlabel polysilicon 688 -1191 688 -1191 0 3
rlabel polysilicon 702 -1185 702 -1185 0 1
rlabel polysilicon 702 -1191 702 -1191 0 3
rlabel polysilicon 709 -1185 709 -1185 0 1
rlabel polysilicon 709 -1191 709 -1191 0 3
rlabel polysilicon 2 -1256 2 -1256 0 1
rlabel polysilicon 2 -1262 2 -1262 0 3
rlabel polysilicon 9 -1256 9 -1256 0 1
rlabel polysilicon 9 -1262 9 -1262 0 3
rlabel polysilicon 16 -1256 16 -1256 0 1
rlabel polysilicon 16 -1262 16 -1262 0 3
rlabel polysilicon 23 -1256 23 -1256 0 1
rlabel polysilicon 23 -1262 23 -1262 0 3
rlabel polysilicon 30 -1256 30 -1256 0 1
rlabel polysilicon 30 -1262 30 -1262 0 3
rlabel polysilicon 37 -1256 37 -1256 0 1
rlabel polysilicon 37 -1262 37 -1262 0 3
rlabel polysilicon 44 -1262 44 -1262 0 3
rlabel polysilicon 47 -1262 47 -1262 0 4
rlabel polysilicon 54 -1256 54 -1256 0 2
rlabel polysilicon 58 -1256 58 -1256 0 1
rlabel polysilicon 61 -1262 61 -1262 0 4
rlabel polysilicon 65 -1256 65 -1256 0 1
rlabel polysilicon 65 -1262 65 -1262 0 3
rlabel polysilicon 75 -1256 75 -1256 0 2
rlabel polysilicon 72 -1262 72 -1262 0 3
rlabel polysilicon 79 -1256 79 -1256 0 1
rlabel polysilicon 79 -1262 79 -1262 0 3
rlabel polysilicon 86 -1256 86 -1256 0 1
rlabel polysilicon 86 -1262 86 -1262 0 3
rlabel polysilicon 93 -1256 93 -1256 0 1
rlabel polysilicon 93 -1262 93 -1262 0 3
rlabel polysilicon 100 -1256 100 -1256 0 1
rlabel polysilicon 103 -1262 103 -1262 0 4
rlabel polysilicon 107 -1256 107 -1256 0 1
rlabel polysilicon 110 -1256 110 -1256 0 2
rlabel polysilicon 114 -1256 114 -1256 0 1
rlabel polysilicon 114 -1262 114 -1262 0 3
rlabel polysilicon 124 -1256 124 -1256 0 2
rlabel polysilicon 121 -1262 121 -1262 0 3
rlabel polysilicon 128 -1256 128 -1256 0 1
rlabel polysilicon 128 -1262 128 -1262 0 3
rlabel polysilicon 135 -1256 135 -1256 0 1
rlabel polysilicon 135 -1262 135 -1262 0 3
rlabel polysilicon 142 -1256 142 -1256 0 1
rlabel polysilicon 145 -1262 145 -1262 0 4
rlabel polysilicon 149 -1256 149 -1256 0 1
rlabel polysilicon 149 -1262 149 -1262 0 3
rlabel polysilicon 156 -1256 156 -1256 0 1
rlabel polysilicon 156 -1262 156 -1262 0 3
rlabel polysilicon 166 -1256 166 -1256 0 2
rlabel polysilicon 163 -1262 163 -1262 0 3
rlabel polysilicon 170 -1256 170 -1256 0 1
rlabel polysilicon 170 -1262 170 -1262 0 3
rlabel polysilicon 177 -1256 177 -1256 0 1
rlabel polysilicon 177 -1262 177 -1262 0 3
rlabel polysilicon 180 -1262 180 -1262 0 4
rlabel polysilicon 187 -1256 187 -1256 0 2
rlabel polysilicon 184 -1262 184 -1262 0 3
rlabel polysilicon 187 -1262 187 -1262 0 4
rlabel polysilicon 194 -1256 194 -1256 0 2
rlabel polysilicon 191 -1262 191 -1262 0 3
rlabel polysilicon 194 -1262 194 -1262 0 4
rlabel polysilicon 201 -1256 201 -1256 0 2
rlabel polysilicon 205 -1256 205 -1256 0 1
rlabel polysilicon 205 -1262 205 -1262 0 3
rlabel polysilicon 212 -1256 212 -1256 0 1
rlabel polysilicon 212 -1262 212 -1262 0 3
rlabel polysilicon 215 -1262 215 -1262 0 4
rlabel polysilicon 219 -1262 219 -1262 0 3
rlabel polysilicon 222 -1262 222 -1262 0 4
rlabel polysilicon 226 -1256 226 -1256 0 1
rlabel polysilicon 229 -1256 229 -1256 0 2
rlabel polysilicon 233 -1256 233 -1256 0 1
rlabel polysilicon 233 -1262 233 -1262 0 3
rlabel polysilicon 236 -1262 236 -1262 0 4
rlabel polysilicon 240 -1256 240 -1256 0 1
rlabel polysilicon 240 -1262 240 -1262 0 3
rlabel polysilicon 247 -1256 247 -1256 0 1
rlabel polysilicon 250 -1256 250 -1256 0 2
rlabel polysilicon 247 -1262 247 -1262 0 3
rlabel polysilicon 250 -1262 250 -1262 0 4
rlabel polysilicon 254 -1256 254 -1256 0 1
rlabel polysilicon 257 -1256 257 -1256 0 2
rlabel polysilicon 254 -1262 254 -1262 0 3
rlabel polysilicon 257 -1262 257 -1262 0 4
rlabel polysilicon 261 -1256 261 -1256 0 1
rlabel polysilicon 261 -1262 261 -1262 0 3
rlabel polysilicon 268 -1256 268 -1256 0 1
rlabel polysilicon 268 -1262 268 -1262 0 3
rlabel polysilicon 271 -1262 271 -1262 0 4
rlabel polysilicon 275 -1256 275 -1256 0 1
rlabel polysilicon 275 -1262 275 -1262 0 3
rlabel polysilicon 282 -1256 282 -1256 0 1
rlabel polysilicon 282 -1262 282 -1262 0 3
rlabel polysilicon 289 -1256 289 -1256 0 1
rlabel polysilicon 289 -1262 289 -1262 0 3
rlabel polysilicon 296 -1256 296 -1256 0 1
rlabel polysilicon 296 -1262 296 -1262 0 3
rlabel polysilicon 306 -1256 306 -1256 0 2
rlabel polysilicon 303 -1262 303 -1262 0 3
rlabel polysilicon 306 -1262 306 -1262 0 4
rlabel polysilicon 310 -1256 310 -1256 0 1
rlabel polysilicon 313 -1262 313 -1262 0 4
rlabel polysilicon 317 -1256 317 -1256 0 1
rlabel polysilicon 317 -1262 317 -1262 0 3
rlabel polysilicon 324 -1256 324 -1256 0 1
rlabel polysilicon 327 -1256 327 -1256 0 2
rlabel polysilicon 324 -1262 324 -1262 0 3
rlabel polysilicon 327 -1262 327 -1262 0 4
rlabel polysilicon 331 -1256 331 -1256 0 1
rlabel polysilicon 331 -1262 331 -1262 0 3
rlabel polysilicon 338 -1256 338 -1256 0 1
rlabel polysilicon 338 -1262 338 -1262 0 3
rlabel polysilicon 345 -1256 345 -1256 0 1
rlabel polysilicon 345 -1262 345 -1262 0 3
rlabel polysilicon 352 -1256 352 -1256 0 1
rlabel polysilicon 359 -1256 359 -1256 0 1
rlabel polysilicon 359 -1262 359 -1262 0 3
rlabel polysilicon 366 -1256 366 -1256 0 1
rlabel polysilicon 366 -1262 366 -1262 0 3
rlabel polysilicon 373 -1256 373 -1256 0 1
rlabel polysilicon 373 -1262 373 -1262 0 3
rlabel polysilicon 380 -1256 380 -1256 0 1
rlabel polysilicon 383 -1256 383 -1256 0 2
rlabel polysilicon 380 -1262 380 -1262 0 3
rlabel polysilicon 383 -1262 383 -1262 0 4
rlabel polysilicon 387 -1256 387 -1256 0 1
rlabel polysilicon 387 -1262 387 -1262 0 3
rlabel polysilicon 394 -1256 394 -1256 0 1
rlabel polysilicon 397 -1256 397 -1256 0 2
rlabel polysilicon 397 -1262 397 -1262 0 4
rlabel polysilicon 401 -1256 401 -1256 0 1
rlabel polysilicon 401 -1262 401 -1262 0 3
rlabel polysilicon 408 -1256 408 -1256 0 1
rlabel polysilicon 408 -1262 408 -1262 0 3
rlabel polysilicon 415 -1256 415 -1256 0 1
rlabel polysilicon 415 -1262 415 -1262 0 3
rlabel polysilicon 422 -1256 422 -1256 0 1
rlabel polysilicon 422 -1262 422 -1262 0 3
rlabel polysilicon 429 -1256 429 -1256 0 1
rlabel polysilicon 432 -1256 432 -1256 0 2
rlabel polysilicon 432 -1262 432 -1262 0 4
rlabel polysilicon 436 -1256 436 -1256 0 1
rlabel polysilicon 436 -1262 436 -1262 0 3
rlabel polysilicon 443 -1256 443 -1256 0 1
rlabel polysilicon 443 -1262 443 -1262 0 3
rlabel polysilicon 450 -1256 450 -1256 0 1
rlabel polysilicon 453 -1256 453 -1256 0 2
rlabel polysilicon 453 -1262 453 -1262 0 4
rlabel polysilicon 457 -1256 457 -1256 0 1
rlabel polysilicon 460 -1256 460 -1256 0 2
rlabel polysilicon 460 -1262 460 -1262 0 4
rlabel polysilicon 464 -1256 464 -1256 0 1
rlabel polysilicon 464 -1262 464 -1262 0 3
rlabel polysilicon 471 -1256 471 -1256 0 1
rlabel polysilicon 471 -1262 471 -1262 0 3
rlabel polysilicon 478 -1256 478 -1256 0 1
rlabel polysilicon 478 -1262 478 -1262 0 3
rlabel polysilicon 485 -1256 485 -1256 0 1
rlabel polysilicon 485 -1262 485 -1262 0 3
rlabel polysilicon 492 -1256 492 -1256 0 1
rlabel polysilicon 495 -1262 495 -1262 0 4
rlabel polysilicon 499 -1256 499 -1256 0 1
rlabel polysilicon 499 -1262 499 -1262 0 3
rlabel polysilicon 506 -1256 506 -1256 0 1
rlabel polysilicon 506 -1262 506 -1262 0 3
rlabel polysilicon 513 -1256 513 -1256 0 1
rlabel polysilicon 513 -1262 513 -1262 0 3
rlabel polysilicon 520 -1256 520 -1256 0 1
rlabel polysilicon 520 -1262 520 -1262 0 3
rlabel polysilicon 527 -1256 527 -1256 0 1
rlabel polysilicon 527 -1262 527 -1262 0 3
rlabel polysilicon 534 -1256 534 -1256 0 1
rlabel polysilicon 534 -1262 534 -1262 0 3
rlabel polysilicon 541 -1256 541 -1256 0 1
rlabel polysilicon 541 -1262 541 -1262 0 3
rlabel polysilicon 548 -1256 548 -1256 0 1
rlabel polysilicon 548 -1262 548 -1262 0 3
rlabel polysilicon 555 -1256 555 -1256 0 1
rlabel polysilicon 555 -1262 555 -1262 0 3
rlabel polysilicon 562 -1256 562 -1256 0 1
rlabel polysilicon 562 -1262 562 -1262 0 3
rlabel polysilicon 569 -1256 569 -1256 0 1
rlabel polysilicon 569 -1262 569 -1262 0 3
rlabel polysilicon 576 -1256 576 -1256 0 1
rlabel polysilicon 576 -1262 576 -1262 0 3
rlabel polysilicon 583 -1256 583 -1256 0 1
rlabel polysilicon 583 -1262 583 -1262 0 3
rlabel polysilicon 590 -1256 590 -1256 0 1
rlabel polysilicon 590 -1262 590 -1262 0 3
rlabel polysilicon 597 -1256 597 -1256 0 1
rlabel polysilicon 597 -1262 597 -1262 0 3
rlabel polysilicon 604 -1256 604 -1256 0 1
rlabel polysilicon 604 -1262 604 -1262 0 3
rlabel polysilicon 611 -1256 611 -1256 0 1
rlabel polysilicon 611 -1262 611 -1262 0 3
rlabel polysilicon 618 -1256 618 -1256 0 1
rlabel polysilicon 618 -1262 618 -1262 0 3
rlabel polysilicon 625 -1256 625 -1256 0 1
rlabel polysilicon 625 -1262 625 -1262 0 3
rlabel polysilicon 632 -1256 632 -1256 0 1
rlabel polysilicon 632 -1262 632 -1262 0 3
rlabel polysilicon 639 -1256 639 -1256 0 1
rlabel polysilicon 639 -1262 639 -1262 0 3
rlabel polysilicon 646 -1256 646 -1256 0 1
rlabel polysilicon 646 -1262 646 -1262 0 3
rlabel polysilicon 653 -1256 653 -1256 0 1
rlabel polysilicon 653 -1262 653 -1262 0 3
rlabel polysilicon 660 -1256 660 -1256 0 1
rlabel polysilicon 660 -1262 660 -1262 0 3
rlabel polysilicon 667 -1256 667 -1256 0 1
rlabel polysilicon 667 -1262 667 -1262 0 3
rlabel polysilicon 674 -1256 674 -1256 0 1
rlabel polysilicon 674 -1262 674 -1262 0 3
rlabel polysilicon 681 -1256 681 -1256 0 1
rlabel polysilicon 681 -1262 681 -1262 0 3
rlabel polysilicon 688 -1256 688 -1256 0 1
rlabel polysilicon 688 -1262 688 -1262 0 3
rlabel polysilicon 695 -1256 695 -1256 0 1
rlabel polysilicon 695 -1262 695 -1262 0 3
rlabel polysilicon 702 -1256 702 -1256 0 1
rlabel polysilicon 705 -1256 705 -1256 0 2
rlabel polysilicon 702 -1262 702 -1262 0 3
rlabel polysilicon 705 -1262 705 -1262 0 4
rlabel polysilicon 712 -1256 712 -1256 0 2
rlabel polysilicon 712 -1262 712 -1262 0 4
rlabel polysilicon 716 -1256 716 -1256 0 1
rlabel polysilicon 716 -1262 716 -1262 0 3
rlabel polysilicon 2 -1327 2 -1327 0 1
rlabel polysilicon 2 -1333 2 -1333 0 3
rlabel polysilicon 9 -1327 9 -1327 0 1
rlabel polysilicon 9 -1333 9 -1333 0 3
rlabel polysilicon 19 -1333 19 -1333 0 4
rlabel polysilicon 23 -1327 23 -1327 0 1
rlabel polysilicon 23 -1333 23 -1333 0 3
rlabel polysilicon 33 -1333 33 -1333 0 4
rlabel polysilicon 40 -1327 40 -1327 0 2
rlabel polysilicon 44 -1327 44 -1327 0 1
rlabel polysilicon 44 -1333 44 -1333 0 3
rlabel polysilicon 51 -1327 51 -1327 0 1
rlabel polysilicon 51 -1333 51 -1333 0 3
rlabel polysilicon 58 -1327 58 -1327 0 1
rlabel polysilicon 58 -1333 58 -1333 0 3
rlabel polysilicon 65 -1327 65 -1327 0 1
rlabel polysilicon 65 -1333 65 -1333 0 3
rlabel polysilicon 72 -1327 72 -1327 0 1
rlabel polysilicon 75 -1333 75 -1333 0 4
rlabel polysilicon 82 -1327 82 -1327 0 2
rlabel polysilicon 82 -1333 82 -1333 0 4
rlabel polysilicon 86 -1327 86 -1327 0 1
rlabel polysilicon 86 -1333 86 -1333 0 3
rlabel polysilicon 93 -1327 93 -1327 0 1
rlabel polysilicon 93 -1333 93 -1333 0 3
rlabel polysilicon 100 -1327 100 -1327 0 1
rlabel polysilicon 100 -1333 100 -1333 0 3
rlabel polysilicon 107 -1327 107 -1327 0 1
rlabel polysilicon 107 -1333 107 -1333 0 3
rlabel polysilicon 114 -1327 114 -1327 0 1
rlabel polysilicon 114 -1333 114 -1333 0 3
rlabel polysilicon 121 -1327 121 -1327 0 1
rlabel polysilicon 121 -1333 121 -1333 0 3
rlabel polysilicon 131 -1327 131 -1327 0 2
rlabel polysilicon 131 -1333 131 -1333 0 4
rlabel polysilicon 135 -1327 135 -1327 0 1
rlabel polysilicon 138 -1327 138 -1327 0 2
rlabel polysilicon 138 -1333 138 -1333 0 4
rlabel polysilicon 142 -1327 142 -1327 0 1
rlabel polysilicon 142 -1333 142 -1333 0 3
rlabel polysilicon 152 -1333 152 -1333 0 4
rlabel polysilicon 156 -1327 156 -1327 0 1
rlabel polysilicon 156 -1333 156 -1333 0 3
rlabel polysilicon 163 -1327 163 -1327 0 1
rlabel polysilicon 163 -1333 163 -1333 0 3
rlabel polysilicon 170 -1333 170 -1333 0 3
rlabel polysilicon 173 -1333 173 -1333 0 4
rlabel polysilicon 177 -1327 177 -1327 0 1
rlabel polysilicon 180 -1327 180 -1327 0 2
rlabel polysilicon 177 -1333 177 -1333 0 3
rlabel polysilicon 184 -1327 184 -1327 0 1
rlabel polysilicon 184 -1333 184 -1333 0 3
rlabel polysilicon 191 -1327 191 -1327 0 1
rlabel polysilicon 191 -1333 191 -1333 0 3
rlabel polysilicon 198 -1327 198 -1327 0 1
rlabel polysilicon 198 -1333 198 -1333 0 3
rlabel polysilicon 205 -1327 205 -1327 0 1
rlabel polysilicon 208 -1327 208 -1327 0 2
rlabel polysilicon 212 -1327 212 -1327 0 1
rlabel polysilicon 212 -1333 212 -1333 0 3
rlabel polysilicon 219 -1327 219 -1327 0 1
rlabel polysilicon 219 -1333 219 -1333 0 3
rlabel polysilicon 226 -1327 226 -1327 0 1
rlabel polysilicon 226 -1333 226 -1333 0 3
rlabel polysilicon 233 -1327 233 -1327 0 1
rlabel polysilicon 236 -1327 236 -1327 0 2
rlabel polysilicon 233 -1333 233 -1333 0 3
rlabel polysilicon 240 -1327 240 -1327 0 1
rlabel polysilicon 240 -1333 240 -1333 0 3
rlabel polysilicon 247 -1327 247 -1327 0 1
rlabel polysilicon 247 -1333 247 -1333 0 3
rlabel polysilicon 254 -1327 254 -1327 0 1
rlabel polysilicon 254 -1333 254 -1333 0 3
rlabel polysilicon 261 -1327 261 -1327 0 1
rlabel polysilicon 261 -1333 261 -1333 0 3
rlabel polysilicon 268 -1327 268 -1327 0 1
rlabel polysilicon 268 -1333 268 -1333 0 3
rlabel polysilicon 275 -1327 275 -1327 0 1
rlabel polysilicon 275 -1333 275 -1333 0 3
rlabel polysilicon 282 -1327 282 -1327 0 1
rlabel polysilicon 285 -1327 285 -1327 0 2
rlabel polysilicon 282 -1333 282 -1333 0 3
rlabel polysilicon 285 -1333 285 -1333 0 4
rlabel polysilicon 289 -1327 289 -1327 0 1
rlabel polysilicon 289 -1333 289 -1333 0 3
rlabel polysilicon 296 -1327 296 -1327 0 1
rlabel polysilicon 296 -1333 296 -1333 0 3
rlabel polysilicon 299 -1333 299 -1333 0 4
rlabel polysilicon 303 -1327 303 -1327 0 1
rlabel polysilicon 306 -1327 306 -1327 0 2
rlabel polysilicon 310 -1327 310 -1327 0 1
rlabel polysilicon 310 -1333 310 -1333 0 3
rlabel polysilicon 317 -1327 317 -1327 0 1
rlabel polysilicon 317 -1333 317 -1333 0 3
rlabel polysilicon 324 -1327 324 -1327 0 1
rlabel polysilicon 324 -1333 324 -1333 0 3
rlabel polysilicon 327 -1333 327 -1333 0 4
rlabel polysilicon 331 -1327 331 -1327 0 1
rlabel polysilicon 331 -1333 331 -1333 0 3
rlabel polysilicon 338 -1333 338 -1333 0 3
rlabel polysilicon 341 -1333 341 -1333 0 4
rlabel polysilicon 345 -1327 345 -1327 0 1
rlabel polysilicon 345 -1333 345 -1333 0 3
rlabel polysilicon 352 -1327 352 -1327 0 1
rlabel polysilicon 355 -1327 355 -1327 0 2
rlabel polysilicon 352 -1333 352 -1333 0 3
rlabel polysilicon 362 -1327 362 -1327 0 2
rlabel polysilicon 362 -1333 362 -1333 0 4
rlabel polysilicon 366 -1327 366 -1327 0 1
rlabel polysilicon 369 -1327 369 -1327 0 2
rlabel polysilicon 366 -1333 366 -1333 0 3
rlabel polysilicon 369 -1333 369 -1333 0 4
rlabel polysilicon 373 -1327 373 -1327 0 1
rlabel polysilicon 380 -1327 380 -1327 0 1
rlabel polysilicon 380 -1333 380 -1333 0 3
rlabel polysilicon 383 -1333 383 -1333 0 4
rlabel polysilicon 390 -1327 390 -1327 0 2
rlabel polysilicon 387 -1333 387 -1333 0 3
rlabel polysilicon 390 -1333 390 -1333 0 4
rlabel polysilicon 394 -1327 394 -1327 0 1
rlabel polysilicon 397 -1327 397 -1327 0 2
rlabel polysilicon 397 -1333 397 -1333 0 4
rlabel polysilicon 401 -1327 401 -1327 0 1
rlabel polysilicon 401 -1333 401 -1333 0 3
rlabel polysilicon 408 -1327 408 -1327 0 1
rlabel polysilicon 408 -1333 408 -1333 0 3
rlabel polysilicon 415 -1327 415 -1327 0 1
rlabel polysilicon 415 -1333 415 -1333 0 3
rlabel polysilicon 422 -1327 422 -1327 0 1
rlabel polysilicon 422 -1333 422 -1333 0 3
rlabel polysilicon 425 -1333 425 -1333 0 4
rlabel polysilicon 429 -1327 429 -1327 0 1
rlabel polysilicon 429 -1333 429 -1333 0 3
rlabel polysilicon 436 -1327 436 -1327 0 1
rlabel polysilicon 436 -1333 436 -1333 0 3
rlabel polysilicon 443 -1327 443 -1327 0 1
rlabel polysilicon 443 -1333 443 -1333 0 3
rlabel polysilicon 450 -1327 450 -1327 0 1
rlabel polysilicon 457 -1327 457 -1327 0 1
rlabel polysilicon 457 -1333 457 -1333 0 3
rlabel polysilicon 464 -1327 464 -1327 0 1
rlabel polysilicon 474 -1327 474 -1327 0 2
rlabel polysilicon 471 -1333 471 -1333 0 3
rlabel polysilicon 474 -1333 474 -1333 0 4
rlabel polysilicon 478 -1327 478 -1327 0 1
rlabel polysilicon 481 -1333 481 -1333 0 4
rlabel polysilicon 485 -1327 485 -1327 0 1
rlabel polysilicon 485 -1333 485 -1333 0 3
rlabel polysilicon 492 -1327 492 -1327 0 1
rlabel polysilicon 492 -1333 492 -1333 0 3
rlabel polysilicon 499 -1327 499 -1327 0 1
rlabel polysilicon 502 -1327 502 -1327 0 2
rlabel polysilicon 499 -1333 499 -1333 0 3
rlabel polysilicon 506 -1327 506 -1327 0 1
rlabel polysilicon 506 -1333 506 -1333 0 3
rlabel polysilicon 513 -1327 513 -1327 0 1
rlabel polysilicon 513 -1333 513 -1333 0 3
rlabel polysilicon 520 -1327 520 -1327 0 1
rlabel polysilicon 520 -1333 520 -1333 0 3
rlabel polysilicon 527 -1327 527 -1327 0 1
rlabel polysilicon 527 -1333 527 -1333 0 3
rlabel polysilicon 534 -1327 534 -1327 0 1
rlabel polysilicon 534 -1333 534 -1333 0 3
rlabel polysilicon 541 -1327 541 -1327 0 1
rlabel polysilicon 541 -1333 541 -1333 0 3
rlabel polysilicon 548 -1327 548 -1327 0 1
rlabel polysilicon 548 -1333 548 -1333 0 3
rlabel polysilicon 555 -1327 555 -1327 0 1
rlabel polysilicon 555 -1333 555 -1333 0 3
rlabel polysilicon 562 -1327 562 -1327 0 1
rlabel polysilicon 562 -1333 562 -1333 0 3
rlabel polysilicon 569 -1327 569 -1327 0 1
rlabel polysilicon 569 -1333 569 -1333 0 3
rlabel polysilicon 576 -1327 576 -1327 0 1
rlabel polysilicon 576 -1333 576 -1333 0 3
rlabel polysilicon 583 -1327 583 -1327 0 1
rlabel polysilicon 583 -1333 583 -1333 0 3
rlabel polysilicon 590 -1327 590 -1327 0 1
rlabel polysilicon 590 -1333 590 -1333 0 3
rlabel polysilicon 597 -1327 597 -1327 0 1
rlabel polysilicon 597 -1333 597 -1333 0 3
rlabel polysilicon 604 -1327 604 -1327 0 1
rlabel polysilicon 604 -1333 604 -1333 0 3
rlabel polysilicon 611 -1327 611 -1327 0 1
rlabel polysilicon 611 -1333 611 -1333 0 3
rlabel polysilicon 618 -1327 618 -1327 0 1
rlabel polysilicon 618 -1333 618 -1333 0 3
rlabel polysilicon 625 -1327 625 -1327 0 1
rlabel polysilicon 625 -1333 625 -1333 0 3
rlabel polysilicon 632 -1327 632 -1327 0 1
rlabel polysilicon 632 -1333 632 -1333 0 3
rlabel polysilicon 639 -1327 639 -1327 0 1
rlabel polysilicon 639 -1333 639 -1333 0 3
rlabel polysilicon 646 -1333 646 -1333 0 3
rlabel polysilicon 653 -1327 653 -1327 0 1
rlabel polysilicon 653 -1333 653 -1333 0 3
rlabel polysilicon 660 -1327 660 -1327 0 1
rlabel polysilicon 667 -1327 667 -1327 0 1
rlabel polysilicon 670 -1327 670 -1327 0 2
rlabel polysilicon 670 -1333 670 -1333 0 4
rlabel polysilicon 674 -1327 674 -1327 0 1
rlabel polysilicon 674 -1333 674 -1333 0 3
rlabel polysilicon 681 -1327 681 -1327 0 1
rlabel polysilicon 681 -1333 681 -1333 0 3
rlabel polysilicon 702 -1327 702 -1327 0 1
rlabel polysilicon 702 -1333 702 -1333 0 3
rlabel polysilicon 33 -1392 33 -1392 0 4
rlabel polysilicon 37 -1386 37 -1386 0 1
rlabel polysilicon 37 -1392 37 -1392 0 3
rlabel polysilicon 44 -1386 44 -1386 0 1
rlabel polysilicon 44 -1392 44 -1392 0 3
rlabel polysilicon 51 -1386 51 -1386 0 1
rlabel polysilicon 51 -1392 51 -1392 0 3
rlabel polysilicon 58 -1386 58 -1386 0 1
rlabel polysilicon 58 -1392 58 -1392 0 3
rlabel polysilicon 65 -1386 65 -1386 0 1
rlabel polysilicon 65 -1392 65 -1392 0 3
rlabel polysilicon 72 -1386 72 -1386 0 1
rlabel polysilicon 72 -1392 72 -1392 0 3
rlabel polysilicon 79 -1386 79 -1386 0 1
rlabel polysilicon 79 -1392 79 -1392 0 3
rlabel polysilicon 86 -1386 86 -1386 0 1
rlabel polysilicon 86 -1392 86 -1392 0 3
rlabel polysilicon 93 -1386 93 -1386 0 1
rlabel polysilicon 93 -1392 93 -1392 0 3
rlabel polysilicon 100 -1386 100 -1386 0 1
rlabel polysilicon 103 -1392 103 -1392 0 4
rlabel polysilicon 107 -1386 107 -1386 0 1
rlabel polysilicon 107 -1392 107 -1392 0 3
rlabel polysilicon 114 -1386 114 -1386 0 1
rlabel polysilicon 114 -1392 114 -1392 0 3
rlabel polysilicon 121 -1386 121 -1386 0 1
rlabel polysilicon 124 -1386 124 -1386 0 2
rlabel polysilicon 128 -1386 128 -1386 0 1
rlabel polysilicon 128 -1392 128 -1392 0 3
rlabel polysilicon 135 -1386 135 -1386 0 1
rlabel polysilicon 138 -1386 138 -1386 0 2
rlabel polysilicon 138 -1392 138 -1392 0 4
rlabel polysilicon 145 -1386 145 -1386 0 2
rlabel polysilicon 145 -1392 145 -1392 0 4
rlabel polysilicon 149 -1386 149 -1386 0 1
rlabel polysilicon 149 -1392 149 -1392 0 3
rlabel polysilicon 159 -1386 159 -1386 0 2
rlabel polysilicon 156 -1392 156 -1392 0 3
rlabel polysilicon 163 -1386 163 -1386 0 1
rlabel polysilicon 163 -1392 163 -1392 0 3
rlabel polysilicon 170 -1386 170 -1386 0 1
rlabel polysilicon 170 -1392 170 -1392 0 3
rlabel polysilicon 177 -1386 177 -1386 0 1
rlabel polysilicon 177 -1392 177 -1392 0 3
rlabel polysilicon 184 -1386 184 -1386 0 1
rlabel polysilicon 184 -1392 184 -1392 0 3
rlabel polysilicon 187 -1392 187 -1392 0 4
rlabel polysilicon 191 -1386 191 -1386 0 1
rlabel polysilicon 191 -1392 191 -1392 0 3
rlabel polysilicon 198 -1386 198 -1386 0 1
rlabel polysilicon 201 -1386 201 -1386 0 2
rlabel polysilicon 201 -1392 201 -1392 0 4
rlabel polysilicon 205 -1386 205 -1386 0 1
rlabel polysilicon 208 -1386 208 -1386 0 2
rlabel polysilicon 205 -1392 205 -1392 0 3
rlabel polysilicon 212 -1386 212 -1386 0 1
rlabel polysilicon 212 -1392 212 -1392 0 3
rlabel polysilicon 219 -1386 219 -1386 0 1
rlabel polysilicon 222 -1386 222 -1386 0 2
rlabel polysilicon 219 -1392 219 -1392 0 3
rlabel polysilicon 226 -1386 226 -1386 0 1
rlabel polysilicon 226 -1392 226 -1392 0 3
rlabel polysilicon 233 -1392 233 -1392 0 3
rlabel polysilicon 236 -1392 236 -1392 0 4
rlabel polysilicon 240 -1386 240 -1386 0 1
rlabel polysilicon 243 -1386 243 -1386 0 2
rlabel polysilicon 243 -1392 243 -1392 0 4
rlabel polysilicon 247 -1386 247 -1386 0 1
rlabel polysilicon 250 -1386 250 -1386 0 2
rlabel polysilicon 247 -1392 247 -1392 0 3
rlabel polysilicon 254 -1386 254 -1386 0 1
rlabel polysilicon 254 -1392 254 -1392 0 3
rlabel polysilicon 261 -1386 261 -1386 0 1
rlabel polysilicon 261 -1392 261 -1392 0 3
rlabel polysilicon 268 -1386 268 -1386 0 1
rlabel polysilicon 268 -1392 268 -1392 0 3
rlabel polysilicon 275 -1386 275 -1386 0 1
rlabel polysilicon 275 -1392 275 -1392 0 3
rlabel polysilicon 282 -1386 282 -1386 0 1
rlabel polysilicon 285 -1386 285 -1386 0 2
rlabel polysilicon 282 -1392 282 -1392 0 3
rlabel polysilicon 285 -1392 285 -1392 0 4
rlabel polysilicon 289 -1386 289 -1386 0 1
rlabel polysilicon 289 -1392 289 -1392 0 3
rlabel polysilicon 296 -1386 296 -1386 0 1
rlabel polysilicon 296 -1392 296 -1392 0 3
rlabel polysilicon 303 -1386 303 -1386 0 1
rlabel polysilicon 303 -1392 303 -1392 0 3
rlabel polysilicon 310 -1386 310 -1386 0 1
rlabel polysilicon 310 -1392 310 -1392 0 3
rlabel polysilicon 317 -1386 317 -1386 0 1
rlabel polysilicon 317 -1392 317 -1392 0 3
rlabel polysilicon 324 -1386 324 -1386 0 1
rlabel polysilicon 324 -1392 324 -1392 0 3
rlabel polysilicon 331 -1386 331 -1386 0 1
rlabel polysilicon 331 -1392 331 -1392 0 3
rlabel polysilicon 338 -1386 338 -1386 0 1
rlabel polysilicon 338 -1392 338 -1392 0 3
rlabel polysilicon 345 -1386 345 -1386 0 1
rlabel polysilicon 348 -1386 348 -1386 0 2
rlabel polysilicon 352 -1386 352 -1386 0 1
rlabel polysilicon 352 -1392 352 -1392 0 3
rlabel polysilicon 359 -1386 359 -1386 0 1
rlabel polysilicon 362 -1386 362 -1386 0 2
rlabel polysilicon 366 -1386 366 -1386 0 1
rlabel polysilicon 369 -1386 369 -1386 0 2
rlabel polysilicon 366 -1392 366 -1392 0 3
rlabel polysilicon 369 -1392 369 -1392 0 4
rlabel polysilicon 373 -1386 373 -1386 0 1
rlabel polysilicon 373 -1392 373 -1392 0 3
rlabel polysilicon 383 -1386 383 -1386 0 2
rlabel polysilicon 380 -1392 380 -1392 0 3
rlabel polysilicon 383 -1392 383 -1392 0 4
rlabel polysilicon 390 -1386 390 -1386 0 2
rlabel polysilicon 387 -1392 387 -1392 0 3
rlabel polysilicon 394 -1386 394 -1386 0 1
rlabel polysilicon 394 -1392 394 -1392 0 3
rlabel polysilicon 404 -1386 404 -1386 0 2
rlabel polysilicon 401 -1392 401 -1392 0 3
rlabel polysilicon 404 -1392 404 -1392 0 4
rlabel polysilicon 408 -1386 408 -1386 0 1
rlabel polysilicon 408 -1392 408 -1392 0 3
rlabel polysilicon 418 -1386 418 -1386 0 2
rlabel polysilicon 418 -1392 418 -1392 0 4
rlabel polysilicon 425 -1386 425 -1386 0 2
rlabel polysilicon 425 -1392 425 -1392 0 4
rlabel polysilicon 429 -1392 429 -1392 0 3
rlabel polysilicon 432 -1392 432 -1392 0 4
rlabel polysilicon 436 -1386 436 -1386 0 1
rlabel polysilicon 436 -1392 436 -1392 0 3
rlabel polysilicon 443 -1386 443 -1386 0 1
rlabel polysilicon 443 -1392 443 -1392 0 3
rlabel polysilicon 450 -1386 450 -1386 0 1
rlabel polysilicon 450 -1392 450 -1392 0 3
rlabel polysilicon 460 -1386 460 -1386 0 2
rlabel polysilicon 460 -1392 460 -1392 0 4
rlabel polysilicon 464 -1386 464 -1386 0 1
rlabel polysilicon 464 -1392 464 -1392 0 3
rlabel polysilicon 471 -1386 471 -1386 0 1
rlabel polysilicon 471 -1392 471 -1392 0 3
rlabel polysilicon 478 -1386 478 -1386 0 1
rlabel polysilicon 481 -1386 481 -1386 0 2
rlabel polysilicon 485 -1386 485 -1386 0 1
rlabel polysilicon 485 -1392 485 -1392 0 3
rlabel polysilicon 492 -1386 492 -1386 0 1
rlabel polysilicon 492 -1392 492 -1392 0 3
rlabel polysilicon 499 -1386 499 -1386 0 1
rlabel polysilicon 499 -1392 499 -1392 0 3
rlabel polysilicon 506 -1386 506 -1386 0 1
rlabel polysilicon 506 -1392 506 -1392 0 3
rlabel polysilicon 513 -1386 513 -1386 0 1
rlabel polysilicon 513 -1392 513 -1392 0 3
rlabel polysilicon 520 -1386 520 -1386 0 1
rlabel polysilicon 520 -1392 520 -1392 0 3
rlabel polysilicon 527 -1386 527 -1386 0 1
rlabel polysilicon 527 -1392 527 -1392 0 3
rlabel polysilicon 534 -1386 534 -1386 0 1
rlabel polysilicon 534 -1392 534 -1392 0 3
rlabel polysilicon 541 -1386 541 -1386 0 1
rlabel polysilicon 541 -1392 541 -1392 0 3
rlabel polysilicon 548 -1386 548 -1386 0 1
rlabel polysilicon 548 -1392 548 -1392 0 3
rlabel polysilicon 555 -1386 555 -1386 0 1
rlabel polysilicon 555 -1392 555 -1392 0 3
rlabel polysilicon 562 -1386 562 -1386 0 1
rlabel polysilicon 562 -1392 562 -1392 0 3
rlabel polysilicon 569 -1386 569 -1386 0 1
rlabel polysilicon 569 -1392 569 -1392 0 3
rlabel polysilicon 576 -1386 576 -1386 0 1
rlabel polysilicon 576 -1392 576 -1392 0 3
rlabel polysilicon 583 -1386 583 -1386 0 1
rlabel polysilicon 583 -1392 583 -1392 0 3
rlabel polysilicon 590 -1386 590 -1386 0 1
rlabel polysilicon 590 -1392 590 -1392 0 3
rlabel polysilicon 600 -1386 600 -1386 0 2
rlabel polysilicon 600 -1392 600 -1392 0 4
rlabel polysilicon 604 -1386 604 -1386 0 1
rlabel polysilicon 604 -1392 604 -1392 0 3
rlabel polysilicon 611 -1386 611 -1386 0 1
rlabel polysilicon 611 -1392 611 -1392 0 3
rlabel polysilicon 621 -1386 621 -1386 0 2
rlabel polysilicon 621 -1392 621 -1392 0 4
rlabel polysilicon 625 -1386 625 -1386 0 1
rlabel polysilicon 625 -1392 625 -1392 0 3
rlabel polysilicon 635 -1392 635 -1392 0 4
rlabel polysilicon 639 -1386 639 -1386 0 1
rlabel polysilicon 639 -1392 639 -1392 0 3
rlabel polysilicon 646 -1386 646 -1386 0 1
rlabel polysilicon 646 -1392 646 -1392 0 3
rlabel polysilicon 653 -1386 653 -1386 0 1
rlabel polysilicon 656 -1386 656 -1386 0 2
rlabel polysilicon 660 -1386 660 -1386 0 1
rlabel polysilicon 660 -1392 660 -1392 0 3
rlabel polysilicon 667 -1386 667 -1386 0 1
rlabel polysilicon 667 -1392 667 -1392 0 3
rlabel polysilicon 702 -1386 702 -1386 0 1
rlabel polysilicon 705 -1392 705 -1392 0 4
rlabel polysilicon 37 -1445 37 -1445 0 1
rlabel polysilicon 37 -1451 37 -1451 0 3
rlabel polysilicon 44 -1445 44 -1445 0 1
rlabel polysilicon 44 -1451 44 -1451 0 3
rlabel polysilicon 51 -1445 51 -1445 0 1
rlabel polysilicon 51 -1451 51 -1451 0 3
rlabel polysilicon 58 -1445 58 -1445 0 1
rlabel polysilicon 58 -1451 58 -1451 0 3
rlabel polysilicon 65 -1445 65 -1445 0 1
rlabel polysilicon 65 -1451 65 -1451 0 3
rlabel polysilicon 72 -1445 72 -1445 0 1
rlabel polysilicon 72 -1451 72 -1451 0 3
rlabel polysilicon 79 -1445 79 -1445 0 1
rlabel polysilicon 79 -1451 79 -1451 0 3
rlabel polysilicon 86 -1445 86 -1445 0 1
rlabel polysilicon 86 -1451 86 -1451 0 3
rlabel polysilicon 93 -1445 93 -1445 0 1
rlabel polysilicon 93 -1451 93 -1451 0 3
rlabel polysilicon 103 -1445 103 -1445 0 2
rlabel polysilicon 107 -1445 107 -1445 0 1
rlabel polysilicon 107 -1451 107 -1451 0 3
rlabel polysilicon 117 -1445 117 -1445 0 2
rlabel polysilicon 117 -1451 117 -1451 0 4
rlabel polysilicon 121 -1445 121 -1445 0 1
rlabel polysilicon 124 -1445 124 -1445 0 2
rlabel polysilicon 128 -1445 128 -1445 0 1
rlabel polysilicon 128 -1451 128 -1451 0 3
rlabel polysilicon 135 -1445 135 -1445 0 1
rlabel polysilicon 138 -1445 138 -1445 0 2
rlabel polysilicon 135 -1451 135 -1451 0 3
rlabel polysilicon 145 -1445 145 -1445 0 2
rlabel polysilicon 142 -1451 142 -1451 0 3
rlabel polysilicon 149 -1445 149 -1445 0 1
rlabel polysilicon 149 -1451 149 -1451 0 3
rlabel polysilicon 156 -1451 156 -1451 0 3
rlabel polysilicon 159 -1451 159 -1451 0 4
rlabel polysilicon 163 -1445 163 -1445 0 1
rlabel polysilicon 163 -1451 163 -1451 0 3
rlabel polysilicon 170 -1445 170 -1445 0 1
rlabel polysilicon 170 -1451 170 -1451 0 3
rlabel polysilicon 177 -1445 177 -1445 0 1
rlabel polysilicon 177 -1451 177 -1451 0 3
rlabel polysilicon 184 -1451 184 -1451 0 3
rlabel polysilicon 191 -1445 191 -1445 0 1
rlabel polysilicon 191 -1451 191 -1451 0 3
rlabel polysilicon 198 -1451 198 -1451 0 3
rlabel polysilicon 205 -1445 205 -1445 0 1
rlabel polysilicon 205 -1451 205 -1451 0 3
rlabel polysilicon 212 -1445 212 -1445 0 1
rlabel polysilicon 215 -1445 215 -1445 0 2
rlabel polysilicon 215 -1451 215 -1451 0 4
rlabel polysilicon 219 -1445 219 -1445 0 1
rlabel polysilicon 219 -1451 219 -1451 0 3
rlabel polysilicon 226 -1445 226 -1445 0 1
rlabel polysilicon 229 -1451 229 -1451 0 4
rlabel polysilicon 233 -1445 233 -1445 0 1
rlabel polysilicon 233 -1451 233 -1451 0 3
rlabel polysilicon 240 -1445 240 -1445 0 1
rlabel polysilicon 240 -1451 240 -1451 0 3
rlabel polysilicon 243 -1451 243 -1451 0 4
rlabel polysilicon 247 -1445 247 -1445 0 1
rlabel polysilicon 247 -1451 247 -1451 0 3
rlabel polysilicon 254 -1445 254 -1445 0 1
rlabel polysilicon 254 -1451 254 -1451 0 3
rlabel polysilicon 261 -1445 261 -1445 0 1
rlabel polysilicon 261 -1451 261 -1451 0 3
rlabel polysilicon 268 -1445 268 -1445 0 1
rlabel polysilicon 271 -1445 271 -1445 0 2
rlabel polysilicon 271 -1451 271 -1451 0 4
rlabel polysilicon 275 -1445 275 -1445 0 1
rlabel polysilicon 275 -1451 275 -1451 0 3
rlabel polysilicon 282 -1445 282 -1445 0 1
rlabel polysilicon 282 -1451 282 -1451 0 3
rlabel polysilicon 289 -1445 289 -1445 0 1
rlabel polysilicon 289 -1451 289 -1451 0 3
rlabel polysilicon 296 -1445 296 -1445 0 1
rlabel polysilicon 296 -1451 296 -1451 0 3
rlabel polysilicon 303 -1445 303 -1445 0 1
rlabel polysilicon 303 -1451 303 -1451 0 3
rlabel polysilicon 310 -1445 310 -1445 0 1
rlabel polysilicon 310 -1451 310 -1451 0 3
rlabel polysilicon 317 -1445 317 -1445 0 1
rlabel polysilicon 317 -1451 317 -1451 0 3
rlabel polysilicon 327 -1445 327 -1445 0 2
rlabel polysilicon 324 -1451 324 -1451 0 3
rlabel polysilicon 327 -1451 327 -1451 0 4
rlabel polysilicon 331 -1445 331 -1445 0 1
rlabel polysilicon 331 -1451 331 -1451 0 3
rlabel polysilicon 338 -1445 338 -1445 0 1
rlabel polysilicon 338 -1451 338 -1451 0 3
rlabel polysilicon 345 -1445 345 -1445 0 1
rlabel polysilicon 345 -1451 345 -1451 0 3
rlabel polysilicon 355 -1445 355 -1445 0 2
rlabel polysilicon 359 -1445 359 -1445 0 1
rlabel polysilicon 359 -1451 359 -1451 0 3
rlabel polysilicon 366 -1445 366 -1445 0 1
rlabel polysilicon 369 -1445 369 -1445 0 2
rlabel polysilicon 373 -1445 373 -1445 0 1
rlabel polysilicon 376 -1445 376 -1445 0 2
rlabel polysilicon 380 -1445 380 -1445 0 1
rlabel polysilicon 380 -1451 380 -1451 0 3
rlabel polysilicon 387 -1445 387 -1445 0 1
rlabel polysilicon 390 -1445 390 -1445 0 2
rlabel polysilicon 387 -1451 387 -1451 0 3
rlabel polysilicon 390 -1451 390 -1451 0 4
rlabel polysilicon 394 -1445 394 -1445 0 1
rlabel polysilicon 397 -1445 397 -1445 0 2
rlabel polysilicon 401 -1445 401 -1445 0 1
rlabel polysilicon 401 -1451 401 -1451 0 3
rlabel polysilicon 408 -1445 408 -1445 0 1
rlabel polysilicon 408 -1451 408 -1451 0 3
rlabel polysilicon 415 -1445 415 -1445 0 1
rlabel polysilicon 415 -1451 415 -1451 0 3
rlabel polysilicon 422 -1445 422 -1445 0 1
rlabel polysilicon 422 -1451 422 -1451 0 3
rlabel polysilicon 429 -1445 429 -1445 0 1
rlabel polysilicon 429 -1451 429 -1451 0 3
rlabel polysilicon 436 -1445 436 -1445 0 1
rlabel polysilicon 439 -1445 439 -1445 0 2
rlabel polysilicon 439 -1451 439 -1451 0 4
rlabel polysilicon 443 -1445 443 -1445 0 1
rlabel polysilicon 446 -1445 446 -1445 0 2
rlabel polysilicon 443 -1451 443 -1451 0 3
rlabel polysilicon 446 -1451 446 -1451 0 4
rlabel polysilicon 450 -1445 450 -1445 0 1
rlabel polysilicon 453 -1445 453 -1445 0 2
rlabel polysilicon 457 -1445 457 -1445 0 1
rlabel polysilicon 457 -1451 457 -1451 0 3
rlabel polysilicon 464 -1445 464 -1445 0 1
rlabel polysilicon 464 -1451 464 -1451 0 3
rlabel polysilicon 471 -1445 471 -1445 0 1
rlabel polysilicon 471 -1451 471 -1451 0 3
rlabel polysilicon 478 -1451 478 -1451 0 3
rlabel polysilicon 485 -1445 485 -1445 0 1
rlabel polysilicon 485 -1451 485 -1451 0 3
rlabel polysilicon 492 -1445 492 -1445 0 1
rlabel polysilicon 492 -1451 492 -1451 0 3
rlabel polysilicon 499 -1445 499 -1445 0 1
rlabel polysilicon 499 -1451 499 -1451 0 3
rlabel polysilicon 506 -1445 506 -1445 0 1
rlabel polysilicon 506 -1451 506 -1451 0 3
rlabel polysilicon 513 -1445 513 -1445 0 1
rlabel polysilicon 513 -1451 513 -1451 0 3
rlabel polysilicon 520 -1445 520 -1445 0 1
rlabel polysilicon 520 -1451 520 -1451 0 3
rlabel polysilicon 527 -1445 527 -1445 0 1
rlabel polysilicon 527 -1451 527 -1451 0 3
rlabel polysilicon 534 -1445 534 -1445 0 1
rlabel polysilicon 534 -1451 534 -1451 0 3
rlabel polysilicon 541 -1445 541 -1445 0 1
rlabel polysilicon 541 -1451 541 -1451 0 3
rlabel polysilicon 548 -1445 548 -1445 0 1
rlabel polysilicon 551 -1445 551 -1445 0 2
rlabel polysilicon 555 -1445 555 -1445 0 1
rlabel polysilicon 555 -1451 555 -1451 0 3
rlabel polysilicon 565 -1445 565 -1445 0 2
rlabel polysilicon 562 -1451 562 -1451 0 3
rlabel polysilicon 565 -1451 565 -1451 0 4
rlabel polysilicon 569 -1451 569 -1451 0 3
rlabel polysilicon 572 -1451 572 -1451 0 4
rlabel polysilicon 576 -1445 576 -1445 0 1
rlabel polysilicon 576 -1451 576 -1451 0 3
rlabel polysilicon 583 -1445 583 -1445 0 1
rlabel polysilicon 583 -1451 583 -1451 0 3
rlabel polysilicon 590 -1445 590 -1445 0 1
rlabel polysilicon 590 -1451 590 -1451 0 3
rlabel polysilicon 597 -1445 597 -1445 0 1
rlabel polysilicon 597 -1451 597 -1451 0 3
rlabel polysilicon 604 -1445 604 -1445 0 1
rlabel polysilicon 604 -1451 604 -1451 0 3
rlabel polysilicon 646 -1445 646 -1445 0 1
rlabel polysilicon 705 -1445 705 -1445 0 2
rlabel polysilicon 702 -1451 702 -1451 0 3
rlabel polysilicon 712 -1451 712 -1451 0 4
rlabel polysilicon 16 -1498 16 -1498 0 1
rlabel polysilicon 16 -1504 16 -1504 0 3
rlabel polysilicon 23 -1504 23 -1504 0 3
rlabel polysilicon 30 -1498 30 -1498 0 1
rlabel polysilicon 30 -1504 30 -1504 0 3
rlabel polysilicon 37 -1498 37 -1498 0 1
rlabel polysilicon 37 -1504 37 -1504 0 3
rlabel polysilicon 44 -1498 44 -1498 0 1
rlabel polysilicon 51 -1498 51 -1498 0 1
rlabel polysilicon 51 -1504 51 -1504 0 3
rlabel polysilicon 54 -1504 54 -1504 0 4
rlabel polysilicon 58 -1498 58 -1498 0 1
rlabel polysilicon 58 -1504 58 -1504 0 3
rlabel polysilicon 65 -1498 65 -1498 0 1
rlabel polysilicon 65 -1504 65 -1504 0 3
rlabel polysilicon 72 -1498 72 -1498 0 1
rlabel polysilicon 72 -1504 72 -1504 0 3
rlabel polysilicon 79 -1498 79 -1498 0 1
rlabel polysilicon 79 -1504 79 -1504 0 3
rlabel polysilicon 86 -1498 86 -1498 0 1
rlabel polysilicon 89 -1504 89 -1504 0 4
rlabel polysilicon 93 -1498 93 -1498 0 1
rlabel polysilicon 93 -1504 93 -1504 0 3
rlabel polysilicon 100 -1498 100 -1498 0 1
rlabel polysilicon 100 -1504 100 -1504 0 3
rlabel polysilicon 107 -1498 107 -1498 0 1
rlabel polysilicon 110 -1498 110 -1498 0 2
rlabel polysilicon 114 -1498 114 -1498 0 1
rlabel polysilicon 114 -1504 114 -1504 0 3
rlabel polysilicon 124 -1498 124 -1498 0 2
rlabel polysilicon 121 -1504 121 -1504 0 3
rlabel polysilicon 128 -1498 128 -1498 0 1
rlabel polysilicon 128 -1504 128 -1504 0 3
rlabel polysilicon 135 -1498 135 -1498 0 1
rlabel polysilicon 135 -1504 135 -1504 0 3
rlabel polysilicon 142 -1498 142 -1498 0 1
rlabel polysilicon 142 -1504 142 -1504 0 3
rlabel polysilicon 149 -1504 149 -1504 0 3
rlabel polysilicon 152 -1504 152 -1504 0 4
rlabel polysilicon 156 -1498 156 -1498 0 1
rlabel polysilicon 156 -1504 156 -1504 0 3
rlabel polysilicon 163 -1498 163 -1498 0 1
rlabel polysilicon 166 -1498 166 -1498 0 2
rlabel polysilicon 170 -1504 170 -1504 0 3
rlabel polysilicon 173 -1504 173 -1504 0 4
rlabel polysilicon 177 -1498 177 -1498 0 1
rlabel polysilicon 180 -1498 180 -1498 0 2
rlabel polysilicon 180 -1504 180 -1504 0 4
rlabel polysilicon 184 -1504 184 -1504 0 3
rlabel polysilicon 187 -1504 187 -1504 0 4
rlabel polysilicon 191 -1498 191 -1498 0 1
rlabel polysilicon 191 -1504 191 -1504 0 3
rlabel polysilicon 198 -1498 198 -1498 0 1
rlabel polysilicon 198 -1504 198 -1504 0 3
rlabel polysilicon 205 -1504 205 -1504 0 3
rlabel polysilicon 208 -1504 208 -1504 0 4
rlabel polysilicon 212 -1498 212 -1498 0 1
rlabel polysilicon 212 -1504 212 -1504 0 3
rlabel polysilicon 219 -1498 219 -1498 0 1
rlabel polysilicon 219 -1504 219 -1504 0 3
rlabel polysilicon 226 -1498 226 -1498 0 1
rlabel polysilicon 229 -1504 229 -1504 0 4
rlabel polysilicon 233 -1498 233 -1498 0 1
rlabel polysilicon 236 -1504 236 -1504 0 4
rlabel polysilicon 240 -1498 240 -1498 0 1
rlabel polysilicon 240 -1504 240 -1504 0 3
rlabel polysilicon 250 -1498 250 -1498 0 2
rlabel polysilicon 247 -1504 247 -1504 0 3
rlabel polysilicon 254 -1498 254 -1498 0 1
rlabel polysilicon 254 -1504 254 -1504 0 3
rlabel polysilicon 261 -1498 261 -1498 0 1
rlabel polysilicon 261 -1504 261 -1504 0 3
rlabel polysilicon 268 -1498 268 -1498 0 1
rlabel polysilicon 271 -1498 271 -1498 0 2
rlabel polysilicon 275 -1498 275 -1498 0 1
rlabel polysilicon 275 -1504 275 -1504 0 3
rlabel polysilicon 282 -1498 282 -1498 0 1
rlabel polysilicon 282 -1504 282 -1504 0 3
rlabel polysilicon 289 -1498 289 -1498 0 1
rlabel polysilicon 292 -1498 292 -1498 0 2
rlabel polysilicon 289 -1504 289 -1504 0 3
rlabel polysilicon 292 -1504 292 -1504 0 4
rlabel polysilicon 296 -1498 296 -1498 0 1
rlabel polysilicon 296 -1504 296 -1504 0 3
rlabel polysilicon 306 -1498 306 -1498 0 2
rlabel polysilicon 303 -1504 303 -1504 0 3
rlabel polysilicon 310 -1498 310 -1498 0 1
rlabel polysilicon 310 -1504 310 -1504 0 3
rlabel polysilicon 313 -1504 313 -1504 0 4
rlabel polysilicon 317 -1504 317 -1504 0 3
rlabel polysilicon 320 -1504 320 -1504 0 4
rlabel polysilicon 324 -1498 324 -1498 0 1
rlabel polysilicon 331 -1498 331 -1498 0 1
rlabel polysilicon 331 -1504 331 -1504 0 3
rlabel polysilicon 338 -1498 338 -1498 0 1
rlabel polysilicon 338 -1504 338 -1504 0 3
rlabel polysilicon 345 -1498 345 -1498 0 1
rlabel polysilicon 345 -1504 345 -1504 0 3
rlabel polysilicon 352 -1498 352 -1498 0 1
rlabel polysilicon 352 -1504 352 -1504 0 3
rlabel polysilicon 359 -1498 359 -1498 0 1
rlabel polysilicon 359 -1504 359 -1504 0 3
rlabel polysilicon 366 -1498 366 -1498 0 1
rlabel polysilicon 369 -1498 369 -1498 0 2
rlabel polysilicon 373 -1498 373 -1498 0 1
rlabel polysilicon 373 -1504 373 -1504 0 3
rlabel polysilicon 380 -1498 380 -1498 0 1
rlabel polysilicon 380 -1504 380 -1504 0 3
rlabel polysilicon 387 -1498 387 -1498 0 1
rlabel polysilicon 387 -1504 387 -1504 0 3
rlabel polysilicon 394 -1498 394 -1498 0 1
rlabel polysilicon 394 -1504 394 -1504 0 3
rlabel polysilicon 401 -1498 401 -1498 0 1
rlabel polysilicon 401 -1504 401 -1504 0 3
rlabel polysilicon 408 -1498 408 -1498 0 1
rlabel polysilicon 408 -1504 408 -1504 0 3
rlabel polysilicon 415 -1498 415 -1498 0 1
rlabel polysilicon 415 -1504 415 -1504 0 3
rlabel polysilicon 425 -1498 425 -1498 0 2
rlabel polysilicon 422 -1504 422 -1504 0 3
rlabel polysilicon 429 -1498 429 -1498 0 1
rlabel polysilicon 432 -1498 432 -1498 0 2
rlabel polysilicon 429 -1504 429 -1504 0 3
rlabel polysilicon 436 -1498 436 -1498 0 1
rlabel polysilicon 436 -1504 436 -1504 0 3
rlabel polysilicon 443 -1498 443 -1498 0 1
rlabel polysilicon 443 -1504 443 -1504 0 3
rlabel polysilicon 450 -1498 450 -1498 0 1
rlabel polysilicon 450 -1504 450 -1504 0 3
rlabel polysilicon 457 -1498 457 -1498 0 1
rlabel polysilicon 457 -1504 457 -1504 0 3
rlabel polysilicon 464 -1498 464 -1498 0 1
rlabel polysilicon 464 -1504 464 -1504 0 3
rlabel polysilicon 471 -1498 471 -1498 0 1
rlabel polysilicon 471 -1504 471 -1504 0 3
rlabel polysilicon 478 -1498 478 -1498 0 1
rlabel polysilicon 485 -1498 485 -1498 0 1
rlabel polysilicon 485 -1504 485 -1504 0 3
rlabel polysilicon 492 -1498 492 -1498 0 1
rlabel polysilicon 492 -1504 492 -1504 0 3
rlabel polysilicon 499 -1498 499 -1498 0 1
rlabel polysilicon 499 -1504 499 -1504 0 3
rlabel polysilicon 506 -1498 506 -1498 0 1
rlabel polysilicon 506 -1504 506 -1504 0 3
rlabel polysilicon 513 -1498 513 -1498 0 1
rlabel polysilicon 513 -1504 513 -1504 0 3
rlabel polysilicon 520 -1498 520 -1498 0 1
rlabel polysilicon 520 -1504 520 -1504 0 3
rlabel polysilicon 527 -1498 527 -1498 0 1
rlabel polysilicon 527 -1504 527 -1504 0 3
rlabel polysilicon 534 -1498 534 -1498 0 1
rlabel polysilicon 534 -1504 534 -1504 0 3
rlabel polysilicon 541 -1498 541 -1498 0 1
rlabel polysilicon 541 -1504 541 -1504 0 3
rlabel polysilicon 548 -1498 548 -1498 0 1
rlabel polysilicon 548 -1504 548 -1504 0 3
rlabel polysilicon 555 -1498 555 -1498 0 1
rlabel polysilicon 555 -1504 555 -1504 0 3
rlabel polysilicon 562 -1498 562 -1498 0 1
rlabel polysilicon 565 -1498 565 -1498 0 2
rlabel polysilicon 562 -1504 562 -1504 0 3
rlabel polysilicon 565 -1504 565 -1504 0 4
rlabel polysilicon 569 -1498 569 -1498 0 1
rlabel polysilicon 569 -1504 569 -1504 0 3
rlabel polysilicon 576 -1498 576 -1498 0 1
rlabel polysilicon 576 -1504 576 -1504 0 3
rlabel polysilicon 579 -1504 579 -1504 0 4
rlabel polysilicon 583 -1498 583 -1498 0 1
rlabel polysilicon 583 -1504 583 -1504 0 3
rlabel polysilicon 590 -1498 590 -1498 0 1
rlabel polysilicon 590 -1504 590 -1504 0 3
rlabel polysilicon 51 -1547 51 -1547 0 1
rlabel polysilicon 51 -1553 51 -1553 0 3
rlabel polysilicon 58 -1547 58 -1547 0 1
rlabel polysilicon 65 -1547 65 -1547 0 1
rlabel polysilicon 65 -1553 65 -1553 0 3
rlabel polysilicon 72 -1553 72 -1553 0 3
rlabel polysilicon 75 -1553 75 -1553 0 4
rlabel polysilicon 79 -1547 79 -1547 0 1
rlabel polysilicon 79 -1553 79 -1553 0 3
rlabel polysilicon 86 -1547 86 -1547 0 1
rlabel polysilicon 86 -1553 86 -1553 0 3
rlabel polysilicon 96 -1547 96 -1547 0 2
rlabel polysilicon 96 -1553 96 -1553 0 4
rlabel polysilicon 103 -1553 103 -1553 0 4
rlabel polysilicon 110 -1547 110 -1547 0 2
rlabel polysilicon 107 -1553 107 -1553 0 3
rlabel polysilicon 114 -1547 114 -1547 0 1
rlabel polysilicon 114 -1553 114 -1553 0 3
rlabel polysilicon 121 -1547 121 -1547 0 1
rlabel polysilicon 121 -1553 121 -1553 0 3
rlabel polysilicon 128 -1547 128 -1547 0 1
rlabel polysilicon 128 -1553 128 -1553 0 3
rlabel polysilicon 135 -1547 135 -1547 0 1
rlabel polysilicon 135 -1553 135 -1553 0 3
rlabel polysilicon 142 -1547 142 -1547 0 1
rlabel polysilicon 142 -1553 142 -1553 0 3
rlabel polysilicon 152 -1547 152 -1547 0 2
rlabel polysilicon 149 -1553 149 -1553 0 3
rlabel polysilicon 152 -1553 152 -1553 0 4
rlabel polysilicon 156 -1547 156 -1547 0 1
rlabel polysilicon 156 -1553 156 -1553 0 3
rlabel polysilicon 159 -1553 159 -1553 0 4
rlabel polysilicon 163 -1547 163 -1547 0 1
rlabel polysilicon 163 -1553 163 -1553 0 3
rlabel polysilicon 170 -1547 170 -1547 0 1
rlabel polysilicon 173 -1553 173 -1553 0 4
rlabel polysilicon 177 -1547 177 -1547 0 1
rlabel polysilicon 177 -1553 177 -1553 0 3
rlabel polysilicon 184 -1547 184 -1547 0 1
rlabel polysilicon 184 -1553 184 -1553 0 3
rlabel polysilicon 191 -1553 191 -1553 0 3
rlabel polysilicon 194 -1553 194 -1553 0 4
rlabel polysilicon 198 -1547 198 -1547 0 1
rlabel polysilicon 201 -1547 201 -1547 0 2
rlabel polysilicon 205 -1547 205 -1547 0 1
rlabel polysilicon 205 -1553 205 -1553 0 3
rlabel polysilicon 212 -1547 212 -1547 0 1
rlabel polysilicon 212 -1553 212 -1553 0 3
rlabel polysilicon 222 -1553 222 -1553 0 4
rlabel polysilicon 229 -1547 229 -1547 0 2
rlabel polysilicon 236 -1547 236 -1547 0 2
rlabel polysilicon 236 -1553 236 -1553 0 4
rlabel polysilicon 240 -1547 240 -1547 0 1
rlabel polysilicon 240 -1553 240 -1553 0 3
rlabel polysilicon 243 -1553 243 -1553 0 4
rlabel polysilicon 247 -1547 247 -1547 0 1
rlabel polysilicon 247 -1553 247 -1553 0 3
rlabel polysilicon 254 -1547 254 -1547 0 1
rlabel polysilicon 254 -1553 254 -1553 0 3
rlabel polysilicon 261 -1547 261 -1547 0 1
rlabel polysilicon 261 -1553 261 -1553 0 3
rlabel polysilicon 268 -1547 268 -1547 0 1
rlabel polysilicon 268 -1553 268 -1553 0 3
rlabel polysilicon 275 -1547 275 -1547 0 1
rlabel polysilicon 275 -1553 275 -1553 0 3
rlabel polysilicon 282 -1547 282 -1547 0 1
rlabel polysilicon 285 -1553 285 -1553 0 4
rlabel polysilicon 292 -1553 292 -1553 0 4
rlabel polysilicon 296 -1547 296 -1547 0 1
rlabel polysilicon 296 -1553 296 -1553 0 3
rlabel polysilicon 303 -1547 303 -1547 0 1
rlabel polysilicon 303 -1553 303 -1553 0 3
rlabel polysilicon 310 -1547 310 -1547 0 1
rlabel polysilicon 310 -1553 310 -1553 0 3
rlabel polysilicon 317 -1547 317 -1547 0 1
rlabel polysilicon 317 -1553 317 -1553 0 3
rlabel polysilicon 327 -1547 327 -1547 0 2
rlabel polysilicon 327 -1553 327 -1553 0 4
rlabel polysilicon 331 -1547 331 -1547 0 1
rlabel polysilicon 331 -1553 331 -1553 0 3
rlabel polysilicon 338 -1547 338 -1547 0 1
rlabel polysilicon 338 -1553 338 -1553 0 3
rlabel polysilicon 345 -1547 345 -1547 0 1
rlabel polysilicon 345 -1553 345 -1553 0 3
rlabel polysilicon 352 -1547 352 -1547 0 1
rlabel polysilicon 352 -1553 352 -1553 0 3
rlabel polysilicon 359 -1547 359 -1547 0 1
rlabel polysilicon 359 -1553 359 -1553 0 3
rlabel polysilicon 369 -1547 369 -1547 0 2
rlabel polysilicon 366 -1553 366 -1553 0 3
rlabel polysilicon 369 -1553 369 -1553 0 4
rlabel polysilicon 373 -1547 373 -1547 0 1
rlabel polysilicon 373 -1553 373 -1553 0 3
rlabel polysilicon 380 -1547 380 -1547 0 1
rlabel polysilicon 383 -1547 383 -1547 0 2
rlabel polysilicon 380 -1553 380 -1553 0 3
rlabel polysilicon 387 -1547 387 -1547 0 1
rlabel polysilicon 387 -1553 387 -1553 0 3
rlabel polysilicon 394 -1547 394 -1547 0 1
rlabel polysilicon 394 -1553 394 -1553 0 3
rlabel polysilicon 401 -1547 401 -1547 0 1
rlabel polysilicon 401 -1553 401 -1553 0 3
rlabel polysilicon 408 -1547 408 -1547 0 1
rlabel polysilicon 408 -1553 408 -1553 0 3
rlabel polysilicon 415 -1553 415 -1553 0 3
rlabel polysilicon 425 -1547 425 -1547 0 2
rlabel polysilicon 422 -1553 422 -1553 0 3
rlabel polysilicon 429 -1547 429 -1547 0 1
rlabel polysilicon 429 -1553 429 -1553 0 3
rlabel polysilicon 436 -1547 436 -1547 0 1
rlabel polysilicon 436 -1553 436 -1553 0 3
rlabel polysilicon 443 -1547 443 -1547 0 1
rlabel polysilicon 443 -1553 443 -1553 0 3
rlabel polysilicon 450 -1547 450 -1547 0 1
rlabel polysilicon 450 -1553 450 -1553 0 3
rlabel polysilicon 457 -1547 457 -1547 0 1
rlabel polysilicon 457 -1553 457 -1553 0 3
rlabel polysilicon 464 -1547 464 -1547 0 1
rlabel polysilicon 464 -1553 464 -1553 0 3
rlabel polysilicon 474 -1547 474 -1547 0 2
rlabel polysilicon 478 -1547 478 -1547 0 1
rlabel polysilicon 478 -1553 478 -1553 0 3
rlabel polysilicon 488 -1547 488 -1547 0 2
rlabel polysilicon 492 -1547 492 -1547 0 1
rlabel polysilicon 492 -1553 492 -1553 0 3
rlabel polysilicon 499 -1547 499 -1547 0 1
rlabel polysilicon 499 -1553 499 -1553 0 3
rlabel polysilicon 502 -1553 502 -1553 0 4
rlabel polysilicon 506 -1547 506 -1547 0 1
rlabel polysilicon 506 -1553 506 -1553 0 3
rlabel polysilicon 513 -1547 513 -1547 0 1
rlabel polysilicon 513 -1553 513 -1553 0 3
rlabel polysilicon 520 -1547 520 -1547 0 1
rlabel polysilicon 520 -1553 520 -1553 0 3
rlabel polysilicon 527 -1547 527 -1547 0 1
rlabel polysilicon 527 -1553 527 -1553 0 3
rlabel polysilicon 586 -1553 586 -1553 0 4
rlabel polysilicon 590 -1547 590 -1547 0 1
rlabel polysilicon 590 -1553 590 -1553 0 3
rlabel polysilicon 75 -1590 75 -1590 0 4
rlabel polysilicon 79 -1584 79 -1584 0 1
rlabel polysilicon 79 -1590 79 -1590 0 3
rlabel polysilicon 128 -1584 128 -1584 0 1
rlabel polysilicon 128 -1590 128 -1590 0 3
rlabel polysilicon 135 -1584 135 -1584 0 1
rlabel polysilicon 135 -1590 135 -1590 0 3
rlabel polysilicon 142 -1584 142 -1584 0 1
rlabel polysilicon 145 -1590 145 -1590 0 4
rlabel polysilicon 152 -1584 152 -1584 0 2
rlabel polysilicon 152 -1590 152 -1590 0 4
rlabel polysilicon 159 -1584 159 -1584 0 2
rlabel polysilicon 156 -1590 156 -1590 0 3
rlabel polysilicon 163 -1584 163 -1584 0 1
rlabel polysilicon 163 -1590 163 -1590 0 3
rlabel polysilicon 170 -1584 170 -1584 0 1
rlabel polysilicon 170 -1590 170 -1590 0 3
rlabel polysilicon 177 -1584 177 -1584 0 1
rlabel polysilicon 177 -1590 177 -1590 0 3
rlabel polysilicon 184 -1584 184 -1584 0 1
rlabel polysilicon 184 -1590 184 -1590 0 3
rlabel polysilicon 191 -1584 191 -1584 0 1
rlabel polysilicon 194 -1584 194 -1584 0 2
rlabel polysilicon 191 -1590 191 -1590 0 3
rlabel polysilicon 194 -1590 194 -1590 0 4
rlabel polysilicon 198 -1584 198 -1584 0 1
rlabel polysilicon 201 -1584 201 -1584 0 2
rlabel polysilicon 205 -1590 205 -1590 0 3
rlabel polysilicon 208 -1590 208 -1590 0 4
rlabel polysilicon 212 -1584 212 -1584 0 1
rlabel polysilicon 212 -1590 212 -1590 0 3
rlabel polysilicon 219 -1584 219 -1584 0 1
rlabel polysilicon 222 -1584 222 -1584 0 2
rlabel polysilicon 226 -1584 226 -1584 0 1
rlabel polysilicon 229 -1584 229 -1584 0 2
rlabel polysilicon 226 -1590 226 -1590 0 3
rlabel polysilicon 233 -1584 233 -1584 0 1
rlabel polysilicon 233 -1590 233 -1590 0 3
rlabel polysilicon 240 -1590 240 -1590 0 3
rlabel polysilicon 243 -1590 243 -1590 0 4
rlabel polysilicon 247 -1584 247 -1584 0 1
rlabel polysilicon 247 -1590 247 -1590 0 3
rlabel polysilicon 254 -1584 254 -1584 0 1
rlabel polysilicon 254 -1590 254 -1590 0 3
rlabel polysilicon 261 -1584 261 -1584 0 1
rlabel polysilicon 261 -1590 261 -1590 0 3
rlabel polysilicon 271 -1584 271 -1584 0 2
rlabel polysilicon 268 -1590 268 -1590 0 3
rlabel polysilicon 275 -1584 275 -1584 0 1
rlabel polysilicon 275 -1590 275 -1590 0 3
rlabel polysilicon 282 -1584 282 -1584 0 1
rlabel polysilicon 282 -1590 282 -1590 0 3
rlabel polysilicon 289 -1584 289 -1584 0 1
rlabel polysilicon 289 -1590 289 -1590 0 3
rlabel polysilicon 296 -1584 296 -1584 0 1
rlabel polysilicon 296 -1590 296 -1590 0 3
rlabel polysilicon 303 -1584 303 -1584 0 1
rlabel polysilicon 303 -1590 303 -1590 0 3
rlabel polysilicon 313 -1584 313 -1584 0 2
rlabel polysilicon 310 -1590 310 -1590 0 3
rlabel polysilicon 317 -1584 317 -1584 0 1
rlabel polysilicon 317 -1590 317 -1590 0 3
rlabel polysilicon 320 -1590 320 -1590 0 4
rlabel polysilicon 324 -1584 324 -1584 0 1
rlabel polysilicon 324 -1590 324 -1590 0 3
rlabel polysilicon 331 -1584 331 -1584 0 1
rlabel polysilicon 331 -1590 331 -1590 0 3
rlabel polysilicon 338 -1590 338 -1590 0 3
rlabel polysilicon 345 -1590 345 -1590 0 3
rlabel polysilicon 352 -1584 352 -1584 0 1
rlabel polysilicon 352 -1590 352 -1590 0 3
rlabel polysilicon 359 -1584 359 -1584 0 1
rlabel polysilicon 359 -1590 359 -1590 0 3
rlabel polysilicon 366 -1584 366 -1584 0 1
rlabel polysilicon 369 -1584 369 -1584 0 2
rlabel polysilicon 369 -1590 369 -1590 0 4
rlabel polysilicon 373 -1584 373 -1584 0 1
rlabel polysilicon 373 -1590 373 -1590 0 3
rlabel polysilicon 380 -1584 380 -1584 0 1
rlabel polysilicon 390 -1584 390 -1584 0 2
rlabel polysilicon 387 -1590 387 -1590 0 3
rlabel polysilicon 394 -1584 394 -1584 0 1
rlabel polysilicon 394 -1590 394 -1590 0 3
rlabel polysilicon 401 -1584 401 -1584 0 1
rlabel polysilicon 401 -1590 401 -1590 0 3
rlabel polysilicon 422 -1590 422 -1590 0 3
rlabel polysilicon 429 -1584 429 -1584 0 1
rlabel polysilicon 429 -1590 429 -1590 0 3
rlabel polysilicon 436 -1584 436 -1584 0 1
rlabel polysilicon 436 -1590 436 -1590 0 3
rlabel polysilicon 464 -1584 464 -1584 0 1
rlabel polysilicon 464 -1590 464 -1590 0 3
rlabel polysilicon 471 -1584 471 -1584 0 1
rlabel polysilicon 471 -1590 471 -1590 0 3
rlabel polysilicon 485 -1584 485 -1584 0 1
rlabel polysilicon 485 -1590 485 -1590 0 3
rlabel polysilicon 492 -1584 492 -1584 0 1
rlabel polysilicon 492 -1590 492 -1590 0 3
rlabel polysilicon 506 -1590 506 -1590 0 3
rlabel polysilicon 513 -1584 513 -1584 0 1
rlabel polysilicon 513 -1590 513 -1590 0 3
rlabel polysilicon 33 -1623 33 -1623 0 4
rlabel polysilicon 72 -1617 72 -1617 0 1
rlabel polysilicon 72 -1623 72 -1623 0 3
rlabel polysilicon 82 -1617 82 -1617 0 2
rlabel polysilicon 89 -1617 89 -1617 0 2
rlabel polysilicon 86 -1623 86 -1623 0 3
rlabel polysilicon 89 -1623 89 -1623 0 4
rlabel polysilicon 93 -1617 93 -1617 0 1
rlabel polysilicon 93 -1623 93 -1623 0 3
rlabel polysilicon 100 -1623 100 -1623 0 3
rlabel polysilicon 114 -1617 114 -1617 0 1
rlabel polysilicon 114 -1623 114 -1623 0 3
rlabel polysilicon 121 -1623 121 -1623 0 3
rlabel polysilicon 124 -1623 124 -1623 0 4
rlabel polysilicon 131 -1617 131 -1617 0 2
rlabel polysilicon 135 -1617 135 -1617 0 1
rlabel polysilicon 135 -1623 135 -1623 0 3
rlabel polysilicon 142 -1617 142 -1617 0 1
rlabel polysilicon 142 -1623 142 -1623 0 3
rlabel polysilicon 152 -1617 152 -1617 0 2
rlabel polysilicon 149 -1623 149 -1623 0 3
rlabel polysilicon 156 -1617 156 -1617 0 1
rlabel polysilicon 156 -1623 156 -1623 0 3
rlabel polysilicon 163 -1617 163 -1617 0 1
rlabel polysilicon 163 -1623 163 -1623 0 3
rlabel polysilicon 170 -1617 170 -1617 0 1
rlabel polysilicon 170 -1623 170 -1623 0 3
rlabel polysilicon 177 -1623 177 -1623 0 3
rlabel polysilicon 180 -1623 180 -1623 0 4
rlabel polysilicon 191 -1617 191 -1617 0 1
rlabel polysilicon 201 -1617 201 -1617 0 2
rlabel polysilicon 198 -1623 198 -1623 0 3
rlabel polysilicon 205 -1617 205 -1617 0 1
rlabel polysilicon 205 -1623 205 -1623 0 3
rlabel polysilicon 215 -1617 215 -1617 0 2
rlabel polysilicon 212 -1623 212 -1623 0 3
rlabel polysilicon 215 -1623 215 -1623 0 4
rlabel polysilicon 219 -1617 219 -1617 0 1
rlabel polysilicon 219 -1623 219 -1623 0 3
rlabel polysilicon 226 -1617 226 -1617 0 1
rlabel polysilicon 226 -1623 226 -1623 0 3
rlabel polysilicon 236 -1617 236 -1617 0 2
rlabel polysilicon 236 -1623 236 -1623 0 4
rlabel polysilicon 240 -1617 240 -1617 0 1
rlabel polysilicon 243 -1617 243 -1617 0 2
rlabel polysilicon 240 -1623 240 -1623 0 3
rlabel polysilicon 250 -1617 250 -1617 0 2
rlabel polysilicon 254 -1617 254 -1617 0 1
rlabel polysilicon 254 -1623 254 -1623 0 3
rlabel polysilicon 261 -1617 261 -1617 0 1
rlabel polysilicon 264 -1623 264 -1623 0 4
rlabel polysilicon 268 -1617 268 -1617 0 1
rlabel polysilicon 275 -1617 275 -1617 0 1
rlabel polysilicon 278 -1617 278 -1617 0 2
rlabel polysilicon 275 -1623 275 -1623 0 3
rlabel polysilicon 278 -1623 278 -1623 0 4
rlabel polysilicon 282 -1617 282 -1617 0 1
rlabel polysilicon 289 -1617 289 -1617 0 1
rlabel polysilicon 289 -1623 289 -1623 0 3
rlabel polysilicon 296 -1617 296 -1617 0 1
rlabel polysilicon 299 -1617 299 -1617 0 2
rlabel polysilicon 296 -1623 296 -1623 0 3
rlabel polysilicon 303 -1617 303 -1617 0 1
rlabel polysilicon 303 -1623 303 -1623 0 3
rlabel polysilicon 310 -1617 310 -1617 0 1
rlabel polysilicon 310 -1623 310 -1623 0 3
rlabel polysilicon 317 -1617 317 -1617 0 1
rlabel polysilicon 317 -1623 317 -1623 0 3
rlabel polysilicon 324 -1617 324 -1617 0 1
rlabel polysilicon 324 -1623 324 -1623 0 3
rlabel polysilicon 334 -1617 334 -1617 0 2
rlabel polysilicon 334 -1623 334 -1623 0 4
rlabel polysilicon 338 -1617 338 -1617 0 1
rlabel polysilicon 341 -1617 341 -1617 0 2
rlabel polysilicon 345 -1617 345 -1617 0 1
rlabel polysilicon 345 -1623 345 -1623 0 3
rlabel polysilicon 352 -1617 352 -1617 0 1
rlabel polysilicon 352 -1623 352 -1623 0 3
rlabel polysilicon 359 -1617 359 -1617 0 1
rlabel polysilicon 359 -1623 359 -1623 0 3
rlabel polysilicon 366 -1617 366 -1617 0 1
rlabel polysilicon 366 -1623 366 -1623 0 3
rlabel polysilicon 380 -1617 380 -1617 0 1
rlabel polysilicon 383 -1617 383 -1617 0 2
rlabel polysilicon 387 -1617 387 -1617 0 1
rlabel polysilicon 387 -1623 387 -1623 0 3
rlabel polysilicon 394 -1617 394 -1617 0 1
rlabel polysilicon 394 -1623 394 -1623 0 3
rlabel polysilicon 443 -1617 443 -1617 0 1
rlabel polysilicon 443 -1623 443 -1623 0 3
rlabel polysilicon 467 -1623 467 -1623 0 4
rlabel polysilicon 471 -1617 471 -1617 0 1
rlabel polysilicon 471 -1623 471 -1623 0 3
rlabel polysilicon 485 -1617 485 -1617 0 1
rlabel polysilicon 488 -1623 488 -1623 0 4
rlabel polysilicon 492 -1617 492 -1617 0 1
rlabel polysilicon 492 -1623 492 -1623 0 3
rlabel polysilicon 30 -1646 30 -1646 0 1
rlabel polysilicon 37 -1646 37 -1646 0 1
rlabel polysilicon 37 -1652 37 -1652 0 3
rlabel polysilicon 44 -1646 44 -1646 0 1
rlabel polysilicon 44 -1652 44 -1652 0 3
rlabel polysilicon 51 -1646 51 -1646 0 1
rlabel polysilicon 51 -1652 51 -1652 0 3
rlabel polysilicon 58 -1646 58 -1646 0 1
rlabel polysilicon 65 -1646 65 -1646 0 1
rlabel polysilicon 65 -1652 65 -1652 0 3
rlabel polysilicon 72 -1646 72 -1646 0 1
rlabel polysilicon 72 -1652 72 -1652 0 3
rlabel polysilicon 79 -1646 79 -1646 0 1
rlabel polysilicon 79 -1652 79 -1652 0 3
rlabel polysilicon 86 -1646 86 -1646 0 1
rlabel polysilicon 86 -1652 86 -1652 0 3
rlabel polysilicon 93 -1652 93 -1652 0 3
rlabel polysilicon 96 -1652 96 -1652 0 4
rlabel polysilicon 100 -1646 100 -1646 0 1
rlabel polysilicon 100 -1652 100 -1652 0 3
rlabel polysilicon 107 -1646 107 -1646 0 1
rlabel polysilicon 110 -1646 110 -1646 0 2
rlabel polysilicon 114 -1646 114 -1646 0 1
rlabel polysilicon 114 -1652 114 -1652 0 3
rlabel polysilicon 117 -1652 117 -1652 0 4
rlabel polysilicon 124 -1646 124 -1646 0 2
rlabel polysilicon 121 -1652 121 -1652 0 3
rlabel polysilicon 124 -1652 124 -1652 0 4
rlabel polysilicon 131 -1646 131 -1646 0 2
rlabel polysilicon 128 -1652 128 -1652 0 3
rlabel polysilicon 135 -1646 135 -1646 0 1
rlabel polysilicon 138 -1646 138 -1646 0 2
rlabel polysilicon 138 -1652 138 -1652 0 4
rlabel polysilicon 145 -1646 145 -1646 0 2
rlabel polysilicon 145 -1652 145 -1652 0 4
rlabel polysilicon 149 -1646 149 -1646 0 1
rlabel polysilicon 149 -1652 149 -1652 0 3
rlabel polysilicon 156 -1646 156 -1646 0 1
rlabel polysilicon 156 -1652 156 -1652 0 3
rlabel polysilicon 163 -1646 163 -1646 0 1
rlabel polysilicon 163 -1652 163 -1652 0 3
rlabel polysilicon 170 -1646 170 -1646 0 1
rlabel polysilicon 170 -1652 170 -1652 0 3
rlabel polysilicon 177 -1646 177 -1646 0 1
rlabel polysilicon 177 -1652 177 -1652 0 3
rlabel polysilicon 184 -1652 184 -1652 0 3
rlabel polysilicon 191 -1646 191 -1646 0 1
rlabel polysilicon 191 -1652 191 -1652 0 3
rlabel polysilicon 198 -1646 198 -1646 0 1
rlabel polysilicon 201 -1646 201 -1646 0 2
rlabel polysilicon 205 -1646 205 -1646 0 1
rlabel polysilicon 205 -1652 205 -1652 0 3
rlabel polysilicon 208 -1652 208 -1652 0 4
rlabel polysilicon 212 -1652 212 -1652 0 3
rlabel polysilicon 215 -1652 215 -1652 0 4
rlabel polysilicon 219 -1646 219 -1646 0 1
rlabel polysilicon 222 -1646 222 -1646 0 2
rlabel polysilicon 219 -1652 219 -1652 0 3
rlabel polysilicon 222 -1652 222 -1652 0 4
rlabel polysilicon 226 -1646 226 -1646 0 1
rlabel polysilicon 229 -1646 229 -1646 0 2
rlabel polysilicon 226 -1652 226 -1652 0 3
rlabel polysilicon 233 -1646 233 -1646 0 1
rlabel polysilicon 236 -1652 236 -1652 0 4
rlabel polysilicon 240 -1646 240 -1646 0 1
rlabel polysilicon 240 -1652 240 -1652 0 3
rlabel polysilicon 243 -1652 243 -1652 0 4
rlabel polysilicon 247 -1646 247 -1646 0 1
rlabel polysilicon 247 -1652 247 -1652 0 3
rlabel polysilicon 254 -1646 254 -1646 0 1
rlabel polysilicon 254 -1652 254 -1652 0 3
rlabel polysilicon 261 -1646 261 -1646 0 1
rlabel polysilicon 261 -1652 261 -1652 0 3
rlabel polysilicon 271 -1646 271 -1646 0 2
rlabel polysilicon 268 -1652 268 -1652 0 3
rlabel polysilicon 271 -1652 271 -1652 0 4
rlabel polysilicon 275 -1646 275 -1646 0 1
rlabel polysilicon 275 -1652 275 -1652 0 3
rlabel polysilicon 282 -1646 282 -1646 0 1
rlabel polysilicon 282 -1652 282 -1652 0 3
rlabel polysilicon 289 -1646 289 -1646 0 1
rlabel polysilicon 289 -1652 289 -1652 0 3
rlabel polysilicon 296 -1646 296 -1646 0 1
rlabel polysilicon 296 -1652 296 -1652 0 3
rlabel polysilicon 303 -1646 303 -1646 0 1
rlabel polysilicon 310 -1646 310 -1646 0 1
rlabel polysilicon 310 -1652 310 -1652 0 3
rlabel polysilicon 317 -1646 317 -1646 0 1
rlabel polysilicon 317 -1652 317 -1652 0 3
rlabel polysilicon 327 -1646 327 -1646 0 2
rlabel polysilicon 324 -1652 324 -1652 0 3
rlabel polysilicon 331 -1646 331 -1646 0 1
rlabel polysilicon 331 -1652 331 -1652 0 3
rlabel polysilicon 338 -1646 338 -1646 0 1
rlabel polysilicon 338 -1652 338 -1652 0 3
rlabel polysilicon 345 -1646 345 -1646 0 1
rlabel polysilicon 345 -1652 345 -1652 0 3
rlabel polysilicon 352 -1646 352 -1646 0 1
rlabel polysilicon 352 -1652 352 -1652 0 3
rlabel polysilicon 359 -1646 359 -1646 0 1
rlabel polysilicon 359 -1652 359 -1652 0 3
rlabel polysilicon 366 -1646 366 -1646 0 1
rlabel polysilicon 366 -1652 366 -1652 0 3
rlabel polysilicon 373 -1646 373 -1646 0 1
rlabel polysilicon 373 -1652 373 -1652 0 3
rlabel polysilicon 380 -1646 380 -1646 0 1
rlabel polysilicon 380 -1652 380 -1652 0 3
rlabel polysilicon 387 -1646 387 -1646 0 1
rlabel polysilicon 387 -1652 387 -1652 0 3
rlabel polysilicon 394 -1646 394 -1646 0 1
rlabel polysilicon 394 -1652 394 -1652 0 3
rlabel polysilicon 401 -1646 401 -1646 0 1
rlabel polysilicon 404 -1646 404 -1646 0 2
rlabel polysilicon 2 -1687 2 -1687 0 3
rlabel polysilicon 19 -1681 19 -1681 0 2
rlabel polysilicon 23 -1681 23 -1681 0 1
rlabel polysilicon 23 -1687 23 -1687 0 3
rlabel polysilicon 33 -1687 33 -1687 0 4
rlabel polysilicon 79 -1687 79 -1687 0 3
rlabel polysilicon 103 -1681 103 -1681 0 2
rlabel polysilicon 107 -1681 107 -1681 0 1
rlabel polysilicon 107 -1687 107 -1687 0 3
rlabel polysilicon 114 -1687 114 -1687 0 3
rlabel polysilicon 121 -1681 121 -1681 0 1
rlabel polysilicon 121 -1687 121 -1687 0 3
rlabel polysilicon 131 -1687 131 -1687 0 4
rlabel polysilicon 135 -1681 135 -1681 0 1
rlabel polysilicon 135 -1687 135 -1687 0 3
rlabel polysilicon 145 -1681 145 -1681 0 2
rlabel polysilicon 149 -1681 149 -1681 0 1
rlabel polysilicon 149 -1687 149 -1687 0 3
rlabel polysilicon 156 -1681 156 -1681 0 1
rlabel polysilicon 156 -1687 156 -1687 0 3
rlabel polysilicon 163 -1681 163 -1681 0 1
rlabel polysilicon 163 -1687 163 -1687 0 3
rlabel polysilicon 170 -1687 170 -1687 0 3
rlabel polysilicon 173 -1687 173 -1687 0 4
rlabel polysilicon 177 -1687 177 -1687 0 3
rlabel polysilicon 184 -1687 184 -1687 0 3
rlabel polysilicon 191 -1681 191 -1681 0 1
rlabel polysilicon 191 -1687 191 -1687 0 3
rlabel polysilicon 198 -1681 198 -1681 0 1
rlabel polysilicon 198 -1687 198 -1687 0 3
rlabel polysilicon 205 -1681 205 -1681 0 1
rlabel polysilicon 205 -1687 205 -1687 0 3
rlabel polysilicon 212 -1681 212 -1681 0 1
rlabel polysilicon 212 -1687 212 -1687 0 3
rlabel polysilicon 222 -1681 222 -1681 0 2
rlabel polysilicon 219 -1687 219 -1687 0 3
rlabel polysilicon 226 -1681 226 -1681 0 1
rlabel polysilicon 229 -1681 229 -1681 0 2
rlabel polysilicon 226 -1687 226 -1687 0 3
rlabel polysilicon 229 -1687 229 -1687 0 4
rlabel polysilicon 233 -1681 233 -1681 0 1
rlabel polysilicon 233 -1687 233 -1687 0 3
rlabel polysilicon 240 -1681 240 -1681 0 1
rlabel polysilicon 243 -1687 243 -1687 0 4
rlabel polysilicon 247 -1681 247 -1681 0 1
rlabel polysilicon 247 -1687 247 -1687 0 3
rlabel polysilicon 254 -1687 254 -1687 0 3
rlabel polysilicon 261 -1681 261 -1681 0 1
rlabel polysilicon 264 -1687 264 -1687 0 4
rlabel polysilicon 268 -1681 268 -1681 0 1
rlabel polysilicon 268 -1687 268 -1687 0 3
rlabel polysilicon 275 -1687 275 -1687 0 3
rlabel polysilicon 285 -1681 285 -1681 0 2
rlabel polysilicon 285 -1687 285 -1687 0 4
rlabel polysilicon 289 -1687 289 -1687 0 3
rlabel polysilicon 296 -1681 296 -1681 0 1
rlabel polysilicon 296 -1687 296 -1687 0 3
rlabel polysilicon 303 -1681 303 -1681 0 1
rlabel polysilicon 303 -1687 303 -1687 0 3
rlabel polysilicon 310 -1681 310 -1681 0 1
rlabel polysilicon 310 -1687 310 -1687 0 3
rlabel polysilicon 320 -1681 320 -1681 0 2
rlabel polysilicon 317 -1687 317 -1687 0 3
rlabel polysilicon 324 -1681 324 -1681 0 1
rlabel polysilicon 324 -1687 324 -1687 0 3
rlabel polysilicon 331 -1681 331 -1681 0 1
rlabel polysilicon 331 -1687 331 -1687 0 3
rlabel polysilicon 338 -1681 338 -1681 0 1
rlabel polysilicon 338 -1687 338 -1687 0 3
rlabel polysilicon 348 -1681 348 -1681 0 2
rlabel polysilicon 352 -1681 352 -1681 0 1
rlabel polysilicon 352 -1687 352 -1687 0 3
rlabel polysilicon 359 -1687 359 -1687 0 3
rlabel polysilicon 366 -1681 366 -1681 0 1
rlabel polysilicon 373 -1681 373 -1681 0 1
rlabel polysilicon 373 -1687 373 -1687 0 3
rlabel polysilicon 380 -1681 380 -1681 0 1
rlabel polysilicon 380 -1687 380 -1687 0 3
rlabel polysilicon 390 -1681 390 -1681 0 2
rlabel polysilicon 394 -1681 394 -1681 0 1
rlabel polysilicon 394 -1687 394 -1687 0 3
rlabel polysilicon 401 -1681 401 -1681 0 1
rlabel polysilicon 401 -1687 401 -1687 0 3
rlabel polysilicon 5 -1710 5 -1710 0 4
rlabel polysilicon 9 -1704 9 -1704 0 1
rlabel polysilicon 9 -1710 9 -1710 0 3
rlabel polysilicon 16 -1704 16 -1704 0 1
rlabel polysilicon 30 -1704 30 -1704 0 1
rlabel polysilicon 79 -1704 79 -1704 0 1
rlabel polysilicon 89 -1704 89 -1704 0 2
rlabel polysilicon 96 -1704 96 -1704 0 2
rlabel polysilicon 100 -1704 100 -1704 0 1
rlabel polysilicon 117 -1704 117 -1704 0 2
rlabel polysilicon 121 -1704 121 -1704 0 1
rlabel polysilicon 128 -1704 128 -1704 0 1
rlabel polysilicon 131 -1704 131 -1704 0 2
rlabel polysilicon 128 -1710 128 -1710 0 3
rlabel polysilicon 135 -1704 135 -1704 0 1
rlabel polysilicon 135 -1710 135 -1710 0 3
rlabel polysilicon 142 -1710 142 -1710 0 3
rlabel polysilicon 152 -1710 152 -1710 0 4
rlabel polysilicon 156 -1704 156 -1704 0 1
rlabel polysilicon 156 -1710 156 -1710 0 3
rlabel polysilicon 163 -1704 163 -1704 0 1
rlabel polysilicon 163 -1710 163 -1710 0 3
rlabel polysilicon 170 -1704 170 -1704 0 1
rlabel polysilicon 170 -1710 170 -1710 0 3
rlabel polysilicon 177 -1704 177 -1704 0 1
rlabel polysilicon 177 -1710 177 -1710 0 3
rlabel polysilicon 187 -1710 187 -1710 0 4
rlabel polysilicon 194 -1704 194 -1704 0 2
rlabel polysilicon 201 -1704 201 -1704 0 2
rlabel polysilicon 201 -1710 201 -1710 0 4
rlabel polysilicon 205 -1704 205 -1704 0 1
rlabel polysilicon 205 -1710 205 -1710 0 3
rlabel polysilicon 212 -1704 212 -1704 0 1
rlabel polysilicon 212 -1710 212 -1710 0 3
rlabel polysilicon 222 -1704 222 -1704 0 2
rlabel polysilicon 219 -1710 219 -1710 0 3
rlabel polysilicon 226 -1704 226 -1704 0 1
rlabel polysilicon 226 -1710 226 -1710 0 3
rlabel polysilicon 233 -1704 233 -1704 0 1
rlabel polysilicon 233 -1710 233 -1710 0 3
rlabel polysilicon 243 -1710 243 -1710 0 4
rlabel polysilicon 257 -1704 257 -1704 0 2
rlabel polysilicon 278 -1704 278 -1704 0 2
rlabel polysilicon 285 -1704 285 -1704 0 2
rlabel polysilicon 292 -1704 292 -1704 0 2
rlabel polysilicon 296 -1704 296 -1704 0 1
rlabel polysilicon 303 -1710 303 -1710 0 3
rlabel polysilicon 310 -1704 310 -1704 0 1
rlabel polysilicon 310 -1710 310 -1710 0 3
rlabel polysilicon 317 -1710 317 -1710 0 3
rlabel polysilicon 324 -1704 324 -1704 0 1
rlabel polysilicon 324 -1710 324 -1710 0 3
rlabel polysilicon 352 -1704 352 -1704 0 1
rlabel metal2 177 1 177 1 0 net=1571
rlabel metal2 198 1 198 1 0 net=2635
rlabel metal2 208 1 208 1 0 net=16
rlabel metal2 240 1 240 1 0 net=2475
rlabel metal2 275 1 275 1 0 net=3633
rlabel metal2 289 1 289 1 0 net=2207
rlabel metal2 215 -1 215 -1 0 net=1619
rlabel metal2 243 -1 243 -1 0 net=3757
rlabel metal2 107 -12 107 -12 0 net=896
rlabel metal2 142 -12 142 -12 0 net=1959
rlabel metal2 177 -12 177 -12 0 net=1572
rlabel metal2 219 -12 219 -12 0 net=1620
rlabel metal2 254 -12 254 -12 0 net=3759
rlabel metal2 289 -12 289 -12 0 net=2208
rlabel metal2 149 -14 149 -14 0 net=2697
rlabel metal2 163 -14 163 -14 0 net=392
rlabel metal2 208 -14 208 -14 0 net=3113
rlabel metal2 226 -14 226 -14 0 net=2476
rlabel metal2 264 -14 264 -14 0 net=3119
rlabel metal2 282 -14 282 -14 0 net=3634
rlabel metal2 292 -14 292 -14 0 net=4307
rlabel metal2 184 -16 184 -16 0 net=3251
rlabel metal2 240 -16 240 -16 0 net=1075
rlabel metal2 296 -16 296 -16 0 net=3639
rlabel metal2 191 -18 191 -18 0 net=2636
rlabel metal2 198 -20 198 -20 0 net=3385
rlabel metal2 135 -31 135 -31 0 net=1891
rlabel metal2 149 -31 149 -31 0 net=2698
rlabel metal2 149 -31 149 -31 0 net=2698
rlabel metal2 152 -31 152 -31 0 net=1011
rlabel metal2 177 -31 177 -31 0 net=169
rlabel metal2 233 -31 233 -31 0 net=2759
rlabel metal2 247 -31 247 -31 0 net=2983
rlabel metal2 275 -31 275 -31 0 net=3121
rlabel metal2 275 -31 275 -31 0 net=3121
rlabel metal2 282 -31 282 -31 0 net=4017
rlabel metal2 296 -31 296 -31 0 net=3640
rlabel metal2 310 -31 310 -31 0 net=4309
rlabel metal2 478 -31 478 -31 0 net=3427
rlabel metal2 579 -31 579 -31 0 net=3861
rlabel metal2 142 -33 142 -33 0 net=1960
rlabel metal2 184 -33 184 -33 0 net=3253
rlabel metal2 184 -33 184 -33 0 net=3253
rlabel metal2 191 -33 191 -33 0 net=3386
rlabel metal2 212 -33 212 -33 0 net=3114
rlabel metal2 240 -33 240 -33 0 net=1077
rlabel metal2 257 -33 257 -33 0 net=3760
rlabel metal2 285 -33 285 -33 0 net=64
rlabel metal2 296 -33 296 -33 0 net=3825
rlabel metal2 317 -33 317 -33 0 net=3183
rlabel metal2 79 -44 79 -44 0 net=664
rlabel metal2 135 -44 135 -44 0 net=1892
rlabel metal2 156 -44 156 -44 0 net=1013
rlabel metal2 156 -44 156 -44 0 net=1013
rlabel metal2 170 -44 170 -44 0 net=1095
rlabel metal2 184 -44 184 -44 0 net=3254
rlabel metal2 212 -44 212 -44 0 net=435
rlabel metal2 219 -44 219 -44 0 net=2761
rlabel metal2 240 -44 240 -44 0 net=4018
rlabel metal2 289 -44 289 -44 0 net=1365
rlabel metal2 338 -44 338 -44 0 net=4099
rlabel metal2 352 -44 352 -44 0 net=3919
rlabel metal2 467 -44 467 -44 0 net=3923
rlabel metal2 478 -44 478 -44 0 net=3429
rlabel metal2 576 -44 576 -44 0 net=3863
rlabel metal2 149 -46 149 -46 0 net=3793
rlabel metal2 149 -46 149 -46 0 net=3793
rlabel metal2 177 -46 177 -46 0 net=795
rlabel metal2 212 -46 212 -46 0 net=426
rlabel metal2 247 -46 247 -46 0 net=853
rlabel metal2 292 -46 292 -46 0 net=3184
rlabel metal2 184 -48 184 -48 0 net=1475
rlabel metal2 222 -48 222 -48 0 net=2095
rlabel metal2 233 -48 233 -48 0 net=2984
rlabel metal2 296 -48 296 -48 0 net=3827
rlabel metal2 296 -48 296 -48 0 net=3827
rlabel metal2 310 -48 310 -48 0 net=4310
rlabel metal2 229 -50 229 -50 0 net=2555
rlabel metal2 317 -50 317 -50 0 net=459
rlabel metal2 247 -52 247 -52 0 net=1721
rlabel metal2 324 -52 324 -52 0 net=2153
rlabel metal2 250 -54 250 -54 0 net=3122
rlabel metal2 254 -56 254 -56 0 net=1079
rlabel metal2 254 -56 254 -56 0 net=1079
rlabel metal2 275 -56 275 -56 0 net=3479
rlabel metal2 142 -67 142 -67 0 net=3794
rlabel metal2 170 -67 170 -67 0 net=1097
rlabel metal2 170 -67 170 -67 0 net=1097
rlabel metal2 177 -67 177 -67 0 net=1091
rlabel metal2 177 -67 177 -67 0 net=1091
rlabel metal2 198 -67 198 -67 0 net=904
rlabel metal2 198 -67 198 -67 0 net=904
rlabel metal2 205 -67 205 -67 0 net=1477
rlabel metal2 219 -67 219 -67 0 net=2762
rlabel metal2 247 -67 247 -67 0 net=2556
rlabel metal2 268 -67 268 -67 0 net=1723
rlabel metal2 324 -67 324 -67 0 net=2154
rlabel metal2 324 -67 324 -67 0 net=2154
rlabel metal2 338 -67 338 -67 0 net=4101
rlabel metal2 471 -67 471 -67 0 net=3924
rlabel metal2 471 -67 471 -67 0 net=3924
rlabel metal2 474 -67 474 -67 0 net=3531
rlabel metal2 576 -67 576 -67 0 net=3865
rlabel metal2 576 -67 576 -67 0 net=3865
rlabel metal2 138 -69 138 -69 0 net=2863
rlabel metal2 226 -69 226 -69 0 net=2097
rlabel metal2 240 -69 240 -69 0 net=1366
rlabel metal2 345 -69 345 -69 0 net=3920
rlabel metal2 478 -69 478 -69 0 net=3431
rlabel metal2 478 -69 478 -69 0 net=3431
rlabel metal2 142 -71 142 -71 0 net=3403
rlabel metal2 166 -71 166 -71 0 net=483
rlabel metal2 226 -71 226 -71 0 net=3481
rlabel metal2 278 -71 278 -71 0 net=3828
rlabel metal2 320 -71 320 -71 0 net=3273
rlabel metal2 149 -73 149 -73 0 net=1015
rlabel metal2 236 -73 236 -73 0 net=741
rlabel metal2 296 -73 296 -73 0 net=2197
rlabel metal2 247 -75 247 -75 0 net=1081
rlabel metal2 261 -75 261 -75 0 net=2419
rlabel metal2 240 -77 240 -77 0 net=1597
rlabel metal2 268 -77 268 -77 0 net=747
rlabel metal2 275 -79 275 -79 0 net=3963
rlabel metal2 121 -90 121 -90 0 net=515
rlabel metal2 121 -90 121 -90 0 net=515
rlabel metal2 128 -90 128 -90 0 net=1329
rlabel metal2 142 -90 142 -90 0 net=3404
rlabel metal2 149 -90 149 -90 0 net=1016
rlabel metal2 163 -90 163 -90 0 net=3483
rlabel metal2 233 -90 233 -90 0 net=2099
rlabel metal2 271 -90 271 -90 0 net=3211
rlabel metal2 397 -90 397 -90 0 net=4053
rlabel metal2 481 -90 481 -90 0 net=3532
rlabel metal2 576 -90 576 -90 0 net=3867
rlabel metal2 107 -92 107 -92 0 net=1833
rlabel metal2 152 -92 152 -92 0 net=1565
rlabel metal2 166 -92 166 -92 0 net=1098
rlabel metal2 177 -92 177 -92 0 net=1093
rlabel metal2 187 -92 187 -92 0 net=1001
rlabel metal2 205 -92 205 -92 0 net=560
rlabel metal2 257 -92 257 -92 0 net=2420
rlabel metal2 289 -92 289 -92 0 net=1815
rlabel metal2 338 -92 338 -92 0 net=4102
rlabel metal2 352 -92 352 -92 0 net=3275
rlabel metal2 478 -92 478 -92 0 net=3433
rlabel metal2 576 -92 576 -92 0 net=2303
rlabel metal2 191 -94 191 -94 0 net=4339
rlabel metal2 219 -94 219 -94 0 net=2865
rlabel metal2 310 -94 310 -94 0 net=3149
rlabel metal2 478 -94 478 -94 0 net=1049
rlabel metal2 194 -96 194 -96 0 net=1347
rlabel metal2 240 -96 240 -96 0 net=3964
rlabel metal2 341 -96 341 -96 0 net=716
rlabel metal2 212 -98 212 -98 0 net=1478
rlabel metal2 222 -98 222 -98 0 net=3047
rlabel metal2 212 -100 212 -100 0 net=3501
rlabel metal2 243 -100 243 -100 0 net=1082
rlabel metal2 250 -100 250 -100 0 net=3013
rlabel metal2 338 -100 338 -100 0 net=2345
rlabel metal2 254 -102 254 -102 0 net=1599
rlabel metal2 275 -102 275 -102 0 net=2189
rlabel metal2 317 -102 317 -102 0 net=4107
rlabel metal2 254 -104 254 -104 0 net=228
rlabel metal2 296 -106 296 -106 0 net=2199
rlabel metal2 282 -108 282 -108 0 net=1725
rlabel metal2 180 -110 180 -110 0 net=2357
rlabel metal2 65 -121 65 -121 0 net=1835
rlabel metal2 131 -121 131 -121 0 net=1330
rlabel metal2 145 -121 145 -121 0 net=914
rlabel metal2 173 -121 173 -121 0 net=1094
rlabel metal2 191 -121 191 -121 0 net=4340
rlabel metal2 208 -121 208 -121 0 net=1615
rlabel metal2 264 -121 264 -121 0 net=266
rlabel metal2 289 -121 289 -121 0 net=1817
rlabel metal2 324 -121 324 -121 0 net=3015
rlabel metal2 345 -121 345 -121 0 net=2347
rlabel metal2 345 -121 345 -121 0 net=2347
rlabel metal2 359 -121 359 -121 0 net=3213
rlabel metal2 422 -121 422 -121 0 net=4055
rlabel metal2 478 -121 478 -121 0 net=3434
rlabel metal2 492 -121 492 -121 0 net=1051
rlabel metal2 576 -121 576 -121 0 net=3868
rlabel metal2 590 -121 590 -121 0 net=2305
rlabel metal2 590 -121 590 -121 0 net=2305
rlabel metal2 72 -123 72 -123 0 net=2137
rlabel metal2 107 -123 107 -123 0 net=1569
rlabel metal2 128 -123 128 -123 0 net=1003
rlabel metal2 149 -123 149 -123 0 net=1567
rlabel metal2 163 -123 163 -123 0 net=3484
rlabel metal2 243 -123 243 -123 0 net=2190
rlabel metal2 331 -123 331 -123 0 net=2201
rlabel metal2 86 -125 86 -125 0 net=1635
rlabel metal2 170 -125 170 -125 0 net=1393
rlabel metal2 219 -125 219 -125 0 net=3150
rlabel metal2 380 -125 380 -125 0 net=3277
rlabel metal2 93 -127 93 -127 0 net=3549
rlabel metal2 275 -127 275 -127 0 net=4108
rlabel metal2 387 -127 387 -127 0 net=3893
rlabel metal2 156 -129 156 -129 0 net=2039
rlabel metal2 222 -129 222 -129 0 net=3502
rlabel metal2 282 -129 282 -129 0 net=2359
rlabel metal2 334 -129 334 -129 0 net=3771
rlabel metal2 394 -129 394 -129 0 net=4193
rlabel metal2 177 -131 177 -131 0 net=1733
rlabel metal2 299 -131 299 -131 0 net=3469
rlabel metal2 184 -133 184 -133 0 net=1215
rlabel metal2 303 -133 303 -133 0 net=2867
rlabel metal2 191 -135 191 -135 0 net=1349
rlabel metal2 229 -135 229 -135 0 net=3591
rlabel metal2 352 -135 352 -135 0 net=3049
rlabel metal2 198 -137 198 -137 0 net=1002
rlabel metal2 222 -137 222 -137 0 net=2823
rlabel metal2 352 -137 352 -137 0 net=3855
rlabel metal2 198 -139 198 -139 0 net=1601
rlabel metal2 205 -141 205 -141 0 net=1301
rlabel metal2 261 -141 261 -141 0 net=1726
rlabel metal2 226 -143 226 -143 0 net=2100
rlabel metal2 240 -145 240 -145 0 net=2743
rlabel metal2 240 -147 240 -147 0 net=2185
rlabel metal2 257 -149 257 -149 0 net=3687
rlabel metal2 19 -160 19 -160 0 net=678
rlabel metal2 65 -160 65 -160 0 net=1836
rlabel metal2 131 -160 131 -160 0 net=558
rlabel metal2 163 -160 163 -160 0 net=1302
rlabel metal2 264 -160 264 -160 0 net=2360
rlabel metal2 317 -160 317 -160 0 net=1818
rlabel metal2 352 -160 352 -160 0 net=3278
rlabel metal2 499 -160 499 -160 0 net=1053
rlabel metal2 590 -160 590 -160 0 net=2307
rlabel metal2 590 -160 590 -160 0 net=2307
rlabel metal2 72 -162 72 -162 0 net=2138
rlabel metal2 135 -162 135 -162 0 net=1005
rlabel metal2 135 -162 135 -162 0 net=1005
rlabel metal2 149 -162 149 -162 0 net=1568
rlabel metal2 208 -162 208 -162 0 net=3214
rlabel metal2 79 -164 79 -164 0 net=434
rlabel metal2 149 -164 149 -164 0 net=2041
rlabel metal2 219 -164 219 -164 0 net=1507
rlabel metal2 320 -164 320 -164 0 net=3894
rlabel metal2 79 -166 79 -166 0 net=4215
rlabel metal2 128 -166 128 -166 0 net=1217
rlabel metal2 226 -166 226 -166 0 net=1383
rlabel metal2 268 -166 268 -166 0 net=3689
rlabel metal2 86 -168 86 -168 0 net=1636
rlabel metal2 226 -168 226 -168 0 net=1675
rlabel metal2 345 -168 345 -168 0 net=2349
rlabel metal2 93 -170 93 -170 0 net=3550
rlabel metal2 236 -170 236 -170 0 net=1119
rlabel metal2 278 -170 278 -170 0 net=73
rlabel metal2 100 -172 100 -172 0 net=1735
rlabel metal2 243 -172 243 -172 0 net=3016
rlabel metal2 352 -172 352 -172 0 net=3069
rlabel metal2 103 -174 103 -174 0 net=380
rlabel metal2 177 -174 177 -174 0 net=2191
rlabel metal2 212 -174 212 -174 0 net=2567
rlabel metal2 359 -174 359 -174 0 net=3471
rlabel metal2 86 -176 86 -176 0 net=3843
rlabel metal2 212 -176 212 -176 0 net=776
rlabel metal2 299 -176 299 -176 0 net=2202
rlabel metal2 107 -178 107 -178 0 net=1570
rlabel metal2 282 -178 282 -178 0 net=2993
rlabel metal2 324 -178 324 -178 0 net=2825
rlabel metal2 366 -178 366 -178 0 net=3773
rlabel metal2 366 -178 366 -178 0 net=3773
rlabel metal2 373 -178 373 -178 0 net=2869
rlabel metal2 107 -180 107 -180 0 net=1603
rlabel metal2 254 -180 254 -180 0 net=1617
rlabel metal2 373 -180 373 -180 0 net=3059
rlabel metal2 422 -180 422 -180 0 net=4056
rlabel metal2 114 -182 114 -182 0 net=1395
rlabel metal2 191 -182 191 -182 0 net=1351
rlabel metal2 299 -182 299 -182 0 net=3849
rlabel metal2 401 -182 401 -182 0 net=4195
rlabel metal2 93 -184 93 -184 0 net=882
rlabel metal2 243 -184 243 -184 0 net=3845
rlabel metal2 121 -186 121 -186 0 net=898
rlabel metal2 303 -186 303 -186 0 net=2745
rlabel metal2 394 -186 394 -186 0 net=3857
rlabel metal2 191 -188 191 -188 0 net=1409
rlabel metal2 380 -188 380 -188 0 net=3051
rlabel metal2 261 -190 261 -190 0 net=3245
rlabel metal2 240 -192 240 -192 0 net=1337
rlabel metal2 240 -194 240 -194 0 net=2186
rlabel metal2 275 -196 275 -196 0 net=3592
rlabel metal2 233 -198 233 -198 0 net=448
rlabel metal2 12 -209 12 -209 0 net=466
rlabel metal2 12 -209 12 -209 0 net=466
rlabel metal2 79 -209 79 -209 0 net=4216
rlabel metal2 243 -209 243 -209 0 net=1618
rlabel metal2 348 -209 348 -209 0 net=3472
rlabel metal2 443 -209 443 -209 0 net=3846
rlabel metal2 506 -209 506 -209 0 net=1054
rlabel metal2 562 -209 562 -209 0 net=894
rlabel metal2 590 -209 590 -209 0 net=2309
rlabel metal2 590 -209 590 -209 0 net=2309
rlabel metal2 86 -211 86 -211 0 net=3844
rlabel metal2 219 -211 219 -211 0 net=2568
rlabel metal2 380 -211 380 -211 0 net=3247
rlabel metal2 450 -211 450 -211 0 net=4285
rlabel metal2 100 -213 100 -213 0 net=1736
rlabel metal2 268 -213 268 -213 0 net=1121
rlabel metal2 268 -213 268 -213 0 net=1121
rlabel metal2 278 -213 278 -213 0 net=3690
rlabel metal2 107 -215 107 -215 0 net=1604
rlabel metal2 240 -215 240 -215 0 net=1352
rlabel metal2 296 -215 296 -215 0 net=3060
rlabel metal2 383 -215 383 -215 0 net=3052
rlabel metal2 401 -215 401 -215 0 net=3859
rlabel metal2 401 -215 401 -215 0 net=3859
rlabel metal2 408 -215 408 -215 0 net=4197
rlabel metal2 408 -215 408 -215 0 net=4197
rlabel metal2 114 -217 114 -217 0 net=1396
rlabel metal2 222 -217 222 -217 0 net=2870
rlabel metal2 114 -219 114 -219 0 net=2995
rlabel metal2 236 -219 236 -219 0 net=2994
rlabel metal2 317 -219 317 -219 0 net=3070
rlabel metal2 359 -219 359 -219 0 net=2747
rlabel metal2 128 -221 128 -221 0 net=1218
rlabel metal2 212 -221 212 -221 0 net=447
rlabel metal2 320 -221 320 -221 0 net=4271
rlabel metal2 135 -223 135 -223 0 net=1006
rlabel metal2 149 -223 149 -223 0 net=2043
rlabel metal2 149 -223 149 -223 0 net=2043
rlabel metal2 156 -223 156 -223 0 net=633
rlabel metal2 243 -223 243 -223 0 net=4033
rlabel metal2 128 -225 128 -225 0 net=1369
rlabel metal2 163 -225 163 -225 0 net=2473
rlabel metal2 282 -225 282 -225 0 net=1411
rlabel metal2 324 -225 324 -225 0 net=2827
rlabel metal2 135 -227 135 -227 0 net=1643
rlabel metal2 173 -227 173 -227 0 net=607
rlabel metal2 289 -227 289 -227 0 net=2437
rlabel metal2 331 -227 331 -227 0 net=1677
rlabel metal2 142 -229 142 -229 0 net=2565
rlabel metal2 191 -229 191 -229 0 net=1385
rlabel metal2 254 -229 254 -229 0 net=1339
rlabel metal2 292 -229 292 -229 0 net=1981
rlabel metal2 338 -229 338 -229 0 net=3775
rlabel metal2 177 -231 177 -231 0 net=4315
rlabel metal2 226 -231 226 -231 0 net=1033
rlabel metal2 261 -231 261 -231 0 net=3195
rlabel metal2 184 -233 184 -233 0 net=2193
rlabel metal2 212 -233 212 -233 0 net=250
rlabel metal2 296 -233 296 -233 0 net=3551
rlabel metal2 198 -235 198 -235 0 net=1509
rlabel metal2 345 -235 345 -235 0 net=2350
rlabel metal2 278 -237 278 -237 0 net=2243
rlabel metal2 352 -237 352 -237 0 net=2461
rlabel metal2 387 -237 387 -237 0 net=3851
rlabel metal2 275 -239 275 -239 0 net=4239
rlabel metal2 65 -250 65 -250 0 net=3699
rlabel metal2 107 -250 107 -250 0 net=2763
rlabel metal2 124 -250 124 -250 0 net=323
rlabel metal2 177 -250 177 -250 0 net=4316
rlabel metal2 198 -250 198 -250 0 net=1511
rlabel metal2 268 -250 268 -250 0 net=1123
rlabel metal2 268 -250 268 -250 0 net=1123
rlabel metal2 292 -250 292 -250 0 net=2019
rlabel metal2 366 -250 366 -250 0 net=3860
rlabel metal2 415 -250 415 -250 0 net=4273
rlabel metal2 502 -250 502 -250 0 net=3969
rlabel metal2 562 -250 562 -250 0 net=2369
rlabel metal2 562 -250 562 -250 0 net=2369
rlabel metal2 590 -250 590 -250 0 net=2310
rlabel metal2 600 -250 600 -250 0 net=3053
rlabel metal2 646 -250 646 -250 0 net=4127
rlabel metal2 646 -250 646 -250 0 net=4127
rlabel metal2 79 -252 79 -252 0 net=3841
rlabel metal2 320 -252 320 -252 0 net=3776
rlabel metal2 422 -252 422 -252 0 net=3249
rlabel metal2 471 -252 471 -252 0 net=3279
rlabel metal2 506 -252 506 -252 0 net=1521
rlabel metal2 86 -254 86 -254 0 net=1371
rlabel metal2 135 -254 135 -254 0 net=1644
rlabel metal2 303 -254 303 -254 0 net=2439
rlabel metal2 429 -254 429 -254 0 net=3853
rlabel metal2 114 -256 114 -256 0 net=2996
rlabel metal2 338 -256 338 -256 0 net=3879
rlabel metal2 443 -256 443 -256 0 net=1679
rlabel metal2 443 -256 443 -256 0 net=1679
rlabel metal2 450 -256 450 -256 0 net=4287
rlabel metal2 114 -258 114 -258 0 net=1441
rlabel metal2 135 -258 135 -258 0 net=1653
rlabel metal2 173 -258 173 -258 0 net=1823
rlabel metal2 184 -258 184 -258 0 net=2194
rlabel metal2 247 -258 247 -258 0 net=1035
rlabel metal2 247 -258 247 -258 0 net=1035
rlabel metal2 254 -258 254 -258 0 net=1340
rlabel metal2 320 -258 320 -258 0 net=4198
rlabel metal2 464 -258 464 -258 0 net=3267
rlabel metal2 142 -260 142 -260 0 net=2566
rlabel metal2 257 -260 257 -260 0 net=2828
rlabel metal2 348 -260 348 -260 0 net=2291
rlabel metal2 436 -260 436 -260 0 net=4035
rlabel metal2 142 -262 142 -262 0 net=1243
rlabel metal2 187 -262 187 -262 0 net=425
rlabel metal2 324 -262 324 -262 0 net=3552
rlabel metal2 373 -262 373 -262 0 net=2749
rlabel metal2 149 -264 149 -264 0 net=2044
rlabel metal2 163 -264 163 -264 0 net=2474
rlabel metal2 191 -264 191 -264 0 net=1386
rlabel metal2 303 -264 303 -264 0 net=2259
rlabel metal2 380 -264 380 -264 0 net=3903
rlabel metal2 149 -266 149 -266 0 net=2327
rlabel metal2 208 -266 208 -266 0 net=738
rlabel metal2 236 -266 236 -266 0 net=373
rlabel metal2 352 -266 352 -266 0 net=2463
rlabel metal2 387 -266 387 -266 0 net=4241
rlabel metal2 156 -268 156 -268 0 net=1953
rlabel metal2 222 -268 222 -268 0 net=2244
rlabel metal2 317 -268 317 -268 0 net=2441
rlabel metal2 394 -268 394 -268 0 net=3197
rlabel metal2 163 -270 163 -270 0 net=1151
rlabel metal2 331 -270 331 -270 0 net=1983
rlabel metal2 201 -272 201 -272 0 net=510
rlabel metal2 299 -272 299 -272 0 net=2559
rlabel metal2 208 -274 208 -274 0 net=2287
rlabel metal2 219 -276 219 -276 0 net=1343
rlabel metal2 226 -278 226 -278 0 net=1413
rlabel metal2 275 -280 275 -280 0 net=1445
rlabel metal2 75 -291 75 -291 0 net=263
rlabel metal2 257 -291 257 -291 0 net=2873
rlabel metal2 324 -291 324 -291 0 net=3854
rlabel metal2 516 -291 516 -291 0 net=3355
rlabel metal2 562 -291 562 -291 0 net=2371
rlabel metal2 562 -291 562 -291 0 net=2371
rlabel metal2 604 -291 604 -291 0 net=3055
rlabel metal2 646 -291 646 -291 0 net=4129
rlabel metal2 674 -291 674 -291 0 net=3885
rlabel metal2 79 -293 79 -293 0 net=3842
rlabel metal2 219 -293 219 -293 0 net=1345
rlabel metal2 303 -293 303 -293 0 net=2440
rlabel metal2 425 -293 425 -293 0 net=3250
rlabel metal2 464 -293 464 -293 0 net=4037
rlabel metal2 520 -293 520 -293 0 net=3970
rlabel metal2 649 -293 649 -293 0 net=2837
rlabel metal2 79 -295 79 -295 0 net=2765
rlabel metal2 114 -295 114 -295 0 net=1955
rlabel metal2 170 -295 170 -295 0 net=1825
rlabel metal2 187 -295 187 -295 0 net=281
rlabel metal2 205 -295 205 -295 0 net=1893
rlabel metal2 289 -295 289 -295 0 net=3280
rlabel metal2 527 -295 527 -295 0 net=1522
rlabel metal2 86 -297 86 -297 0 net=1372
rlabel metal2 212 -297 212 -297 0 net=1819
rlabel metal2 236 -297 236 -297 0 net=909
rlabel metal2 390 -297 390 -297 0 net=4274
rlabel metal2 506 -297 506 -297 0 net=3269
rlabel metal2 86 -299 86 -299 0 net=1245
rlabel metal2 219 -299 219 -299 0 net=3337
rlabel metal2 485 -299 485 -299 0 net=4289
rlabel metal2 93 -301 93 -301 0 net=3700
rlabel metal2 247 -301 247 -301 0 net=1036
rlabel metal2 324 -301 324 -301 0 net=2750
rlabel metal2 436 -301 436 -301 0 net=4243
rlabel metal2 93 -303 93 -303 0 net=2329
rlabel metal2 247 -303 247 -303 0 net=2021
rlabel metal2 348 -303 348 -303 0 net=1984
rlabel metal2 394 -303 394 -303 0 net=2661
rlabel metal2 100 -305 100 -305 0 net=1131
rlabel metal2 128 -305 128 -305 0 net=1443
rlabel metal2 254 -305 254 -305 0 net=1125
rlabel metal2 275 -305 275 -305 0 net=1447
rlabel metal2 275 -305 275 -305 0 net=1447
rlabel metal2 282 -305 282 -305 0 net=3875
rlabel metal2 103 -307 103 -307 0 net=1333
rlabel metal2 135 -307 135 -307 0 net=1654
rlabel metal2 261 -307 261 -307 0 net=1512
rlabel metal2 289 -307 289 -307 0 net=2477
rlabel metal2 341 -307 341 -307 0 net=1680
rlabel metal2 107 -309 107 -309 0 net=1153
rlabel metal2 198 -309 198 -309 0 net=1415
rlabel metal2 303 -309 303 -309 0 net=2293
rlabel metal2 443 -309 443 -309 0 net=3329
rlabel metal2 128 -311 128 -311 0 net=1787
rlabel metal2 163 -311 163 -311 0 net=4207
rlabel metal2 191 -311 191 -311 0 net=2079
rlabel metal2 313 -311 313 -311 0 net=3503
rlabel metal2 345 -313 345 -313 0 net=3198
rlabel metal2 352 -315 352 -315 0 net=2443
rlabel metal2 408 -315 408 -315 0 net=3905
rlabel metal2 331 -317 331 -317 0 net=2561
rlabel metal2 366 -317 366 -317 0 net=2289
rlabel metal2 408 -317 408 -317 0 net=2841
rlabel metal2 331 -319 331 -319 0 net=2351
rlabel metal2 415 -319 415 -319 0 net=3881
rlabel metal2 240 -321 240 -321 0 net=2715
rlabel metal2 422 -321 422 -321 0 net=4175
rlabel metal2 229 -323 229 -323 0 net=1313
rlabel metal2 366 -323 366 -323 0 net=2973
rlabel metal2 373 -325 373 -325 0 net=2465
rlabel metal2 359 -327 359 -327 0 net=2261
rlabel metal2 359 -329 359 -329 0 net=3359
rlabel metal2 44 -340 44 -340 0 net=4021
rlabel metal2 338 -340 338 -340 0 net=3270
rlabel metal2 541 -340 541 -340 0 net=4109
rlabel metal2 583 -340 583 -340 0 net=3057
rlabel metal2 642 -340 642 -340 0 net=2547
rlabel metal2 51 -342 51 -342 0 net=1957
rlabel metal2 128 -342 128 -342 0 net=1444
rlabel metal2 166 -342 166 -342 0 net=316
rlabel metal2 243 -342 243 -342 0 net=2131
rlabel metal2 264 -342 264 -342 0 net=4181
rlabel metal2 649 -342 649 -342 0 net=4130
rlabel metal2 660 -342 660 -342 0 net=2839
rlabel metal2 58 -344 58 -344 0 net=2479
rlabel metal2 296 -344 296 -344 0 net=1346
rlabel metal2 341 -344 341 -344 0 net=2662
rlabel metal2 471 -344 471 -344 0 net=3505
rlabel metal2 523 -344 523 -344 0 net=4123
rlabel metal2 667 -344 667 -344 0 net=3887
rlabel metal2 79 -346 79 -346 0 net=2766
rlabel metal2 233 -346 233 -346 0 net=2681
rlabel metal2 359 -346 359 -346 0 net=3997
rlabel metal2 79 -348 79 -348 0 net=1827
rlabel metal2 177 -348 177 -348 0 net=4208
rlabel metal2 233 -348 233 -348 0 net=2562
rlabel metal2 362 -348 362 -348 0 net=4244
rlabel metal2 544 -348 544 -348 0 net=411
rlabel metal2 86 -350 86 -350 0 net=1246
rlabel metal2 177 -350 177 -350 0 net=1029
rlabel metal2 222 -350 222 -350 0 net=782
rlabel metal2 366 -350 366 -350 0 net=4159
rlabel metal2 86 -352 86 -352 0 net=2023
rlabel metal2 254 -352 254 -352 0 net=1127
rlabel metal2 275 -352 275 -352 0 net=1449
rlabel metal2 341 -352 341 -352 0 net=3601
rlabel metal2 548 -352 548 -352 0 net=3357
rlabel metal2 93 -354 93 -354 0 net=2330
rlabel metal2 159 -354 159 -354 0 net=1061
rlabel metal2 292 -354 292 -354 0 net=2485
rlabel metal2 380 -354 380 -354 0 net=2290
rlabel metal2 411 -354 411 -354 0 net=2974
rlabel metal2 460 -354 460 -354 0 net=3589
rlabel metal2 558 -354 558 -354 0 net=2372
rlabel metal2 72 -356 72 -356 0 net=972
rlabel metal2 205 -356 205 -356 0 net=1894
rlabel metal2 327 -356 327 -356 0 net=2791
rlabel metal2 562 -356 562 -356 0 net=4347
rlabel metal2 72 -358 72 -358 0 net=1821
rlabel metal2 236 -358 236 -358 0 net=500
rlabel metal2 327 -358 327 -358 0 net=2955
rlabel metal2 415 -358 415 -358 0 net=2717
rlabel metal2 471 -358 471 -358 0 net=2853
rlabel metal2 93 -360 93 -360 0 net=1133
rlabel metal2 114 -360 114 -360 0 net=2445
rlabel metal2 415 -360 415 -360 0 net=2423
rlabel metal2 478 -360 478 -360 0 net=4039
rlabel metal2 100 -362 100 -362 0 net=1335
rlabel metal2 128 -362 128 -362 0 net=1789
rlabel metal2 142 -362 142 -362 0 net=1159
rlabel metal2 373 -362 373 -362 0 net=2263
rlabel metal2 485 -362 485 -362 0 net=3877
rlabel metal2 68 -364 68 -364 0 net=965
rlabel metal2 152 -364 152 -364 0 net=859
rlabel metal2 380 -364 380 -364 0 net=2237
rlabel metal2 394 -364 394 -364 0 net=2467
rlabel metal2 422 -364 422 -364 0 net=3609
rlabel metal2 107 -366 107 -366 0 net=1154
rlabel metal2 205 -366 205 -366 0 net=1315
rlabel metal2 317 -366 317 -366 0 net=2875
rlabel metal2 422 -366 422 -366 0 net=3360
rlabel metal2 107 -368 107 -368 0 net=2245
rlabel metal2 317 -368 317 -368 0 net=2843
rlabel metal2 492 -368 492 -368 0 net=3883
rlabel metal2 110 -370 110 -370 0 net=3623
rlabel metal2 443 -370 443 -370 0 net=3331
rlabel metal2 499 -370 499 -370 0 net=4177
rlabel metal2 121 -372 121 -372 0 net=2081
rlabel metal2 303 -372 303 -372 0 net=2295
rlabel metal2 450 -372 450 -372 0 net=3907
rlabel metal2 506 -372 506 -372 0 net=4291
rlabel metal2 170 -374 170 -374 0 net=1257
rlabel metal2 303 -374 303 -374 0 net=1807
rlabel metal2 348 -374 348 -374 0 net=4057
rlabel metal2 184 -376 184 -376 0 net=2275
rlabel metal2 310 -376 310 -376 0 net=1573
rlabel metal2 429 -376 429 -376 0 net=3221
rlabel metal2 464 -376 464 -376 0 net=3339
rlabel metal2 184 -378 184 -378 0 net=1417
rlabel metal2 331 -378 331 -378 0 net=2353
rlabel metal2 138 -380 138 -380 0 net=1765
rlabel metal2 282 -380 282 -380 0 net=1373
rlabel metal2 2 -391 2 -391 0 net=3123
rlabel metal2 205 -391 205 -391 0 net=1317
rlabel metal2 233 -391 233 -391 0 net=1574
rlabel metal2 317 -391 317 -391 0 net=2844
rlabel metal2 359 -391 359 -391 0 net=3998
rlabel metal2 628 -391 628 -391 0 net=1715
rlabel metal2 649 -391 649 -391 0 net=2840
rlabel metal2 16 -393 16 -393 0 net=3087
rlabel metal2 303 -393 303 -393 0 net=1809
rlabel metal2 355 -393 355 -393 0 net=2613
rlabel metal2 373 -393 373 -393 0 net=3625
rlabel metal2 597 -393 597 -393 0 net=4125
rlabel metal2 667 -393 667 -393 0 net=3888
rlabel metal2 30 -395 30 -395 0 net=2777
rlabel metal2 44 -395 44 -395 0 net=4022
rlabel metal2 240 -395 240 -395 0 net=2354
rlabel metal2 485 -395 485 -395 0 net=3333
rlabel metal2 485 -395 485 -395 0 net=3333
rlabel metal2 513 -395 513 -395 0 net=3507
rlabel metal2 513 -395 513 -395 0 net=3507
rlabel metal2 527 -395 527 -395 0 net=3603
rlabel metal2 527 -395 527 -395 0 net=3603
rlabel metal2 597 -395 597 -395 0 net=4183
rlabel metal2 667 -395 667 -395 0 net=2549
rlabel metal2 44 -397 44 -397 0 net=2945
rlabel metal2 401 -397 401 -397 0 net=2469
rlabel metal2 436 -397 436 -397 0 net=2719
rlabel metal2 450 -397 450 -397 0 net=3358
rlabel metal2 51 -399 51 -399 0 net=1958
rlabel metal2 149 -399 149 -399 0 net=2277
rlabel metal2 215 -399 215 -399 0 net=2876
rlabel metal2 401 -399 401 -399 0 net=4292
rlabel metal2 51 -401 51 -401 0 net=2195
rlabel metal2 163 -401 163 -401 0 net=1419
rlabel metal2 219 -401 219 -401 0 net=2395
rlabel metal2 436 -401 436 -401 0 net=3590
rlabel metal2 576 -401 576 -401 0 net=3610
rlabel metal2 58 -403 58 -403 0 net=2480
rlabel metal2 373 -403 373 -403 0 net=3345
rlabel metal2 460 -403 460 -403 0 net=2792
rlabel metal2 558 -403 558 -403 0 net=2913
rlabel metal2 583 -403 583 -403 0 net=3058
rlabel metal2 58 -405 58 -405 0 net=2257
rlabel metal2 268 -405 268 -405 0 net=1128
rlabel metal2 317 -405 317 -405 0 net=2487
rlabel metal2 376 -405 376 -405 0 net=2424
rlabel metal2 439 -405 439 -405 0 net=3884
rlabel metal2 65 -407 65 -407 0 net=1041
rlabel metal2 334 -407 334 -407 0 net=3878
rlabel metal2 604 -407 604 -407 0 net=4349
rlabel metal2 72 -409 72 -409 0 net=1822
rlabel metal2 341 -409 341 -409 0 net=2264
rlabel metal2 492 -409 492 -409 0 net=3909
rlabel metal2 569 -409 569 -409 0 net=4111
rlabel metal2 653 -409 653 -409 0 net=3891
rlabel metal2 72 -411 72 -411 0 net=2539
rlabel metal2 254 -411 254 -411 0 net=1063
rlabel metal2 285 -411 285 -411 0 net=1450
rlabel metal2 369 -411 369 -411 0 net=3317
rlabel metal2 541 -411 541 -411 0 net=4041
rlabel metal2 79 -413 79 -413 0 net=1828
rlabel metal2 247 -413 247 -413 0 net=2247
rlabel metal2 380 -413 380 -413 0 net=2239
rlabel metal2 380 -413 380 -413 0 net=2239
rlabel metal2 387 -413 387 -413 0 net=4160
rlabel metal2 79 -415 79 -415 0 net=3701
rlabel metal2 247 -415 247 -415 0 net=2133
rlabel metal2 289 -415 289 -415 0 net=1227
rlabel metal2 387 -415 387 -415 0 net=2297
rlabel metal2 467 -415 467 -415 0 net=4161
rlabel metal2 86 -417 86 -417 0 net=2024
rlabel metal2 345 -417 345 -417 0 net=2683
rlabel metal2 471 -417 471 -417 0 net=2855
rlabel metal2 499 -417 499 -417 0 net=4059
rlabel metal2 555 -417 555 -417 0 net=4179
rlabel metal2 93 -419 93 -419 0 net=1135
rlabel metal2 93 -419 93 -419 0 net=1135
rlabel metal2 100 -419 100 -419 0 net=1336
rlabel metal2 184 -419 184 -419 0 net=2025
rlabel metal2 236 -419 236 -419 0 net=1627
rlabel metal2 408 -419 408 -419 0 net=2957
rlabel metal2 100 -421 100 -421 0 net=1239
rlabel metal2 159 -421 159 -421 0 net=3815
rlabel metal2 107 -423 107 -423 0 net=1767
rlabel metal2 236 -423 236 -423 0 net=80
rlabel metal2 324 -423 324 -423 0 net=3340
rlabel metal2 114 -425 114 -425 0 net=2447
rlabel metal2 408 -425 408 -425 0 net=3685
rlabel metal2 114 -427 114 -427 0 net=1790
rlabel metal2 135 -427 135 -427 0 net=576
rlabel metal2 198 -427 198 -427 0 net=3915
rlabel metal2 121 -429 121 -429 0 net=2083
rlabel metal2 415 -429 415 -429 0 net=3223
rlabel metal2 86 -431 86 -431 0 net=1813
rlabel metal2 128 -431 128 -431 0 net=1259
rlabel metal2 261 -431 261 -431 0 net=1375
rlabel metal2 338 -431 338 -431 0 net=2883
rlabel metal2 142 -433 142 -433 0 net=1161
rlabel metal2 170 -435 170 -435 0 net=1031
rlabel metal2 205 -435 205 -435 0 net=1503
rlabel metal2 23 -437 23 -437 0 net=2949
rlabel metal2 9 -448 9 -448 0 net=21
rlabel metal2 131 -448 131 -448 0 net=3816
rlabel metal2 541 -448 541 -448 0 net=4061
rlabel metal2 558 -448 558 -448 0 net=4112
rlabel metal2 611 -448 611 -448 0 net=4126
rlabel metal2 635 -448 635 -448 0 net=3892
rlabel metal2 660 -448 660 -448 0 net=2551
rlabel metal2 9 -450 9 -450 0 net=4293
rlabel metal2 369 -450 369 -450 0 net=3910
rlabel metal2 583 -450 583 -450 0 net=4351
rlabel metal2 646 -450 646 -450 0 net=4199
rlabel metal2 646 -450 646 -450 0 net=4199
rlabel metal2 653 -450 653 -450 0 net=4283
rlabel metal2 16 -452 16 -452 0 net=3088
rlabel metal2 247 -452 247 -452 0 net=2134
rlabel metal2 292 -452 292 -452 0 net=3224
rlabel metal2 418 -452 418 -452 0 net=3747
rlabel metal2 16 -454 16 -454 0 net=4031
rlabel metal2 142 -454 142 -454 0 net=1032
rlabel metal2 208 -454 208 -454 0 net=1228
rlabel metal2 373 -454 373 -454 0 net=2958
rlabel metal2 520 -454 520 -454 0 net=3627
rlabel metal2 23 -456 23 -456 0 net=2950
rlabel metal2 215 -456 215 -456 0 net=1376
rlabel metal2 275 -456 275 -456 0 net=2449
rlabel metal2 376 -456 376 -456 0 net=3508
rlabel metal2 23 -458 23 -458 0 net=3557
rlabel metal2 107 -458 107 -458 0 net=1769
rlabel metal2 177 -458 177 -458 0 net=3171
rlabel metal2 397 -458 397 -458 0 net=2856
rlabel metal2 499 -458 499 -458 0 net=3917
rlabel metal2 513 -458 513 -458 0 net=3605
rlabel metal2 30 -460 30 -460 0 net=3167
rlabel metal2 142 -460 142 -460 0 net=2249
rlabel metal2 317 -460 317 -460 0 net=2489
rlabel metal2 317 -460 317 -460 0 net=2489
rlabel metal2 324 -460 324 -460 0 net=1551
rlabel metal2 436 -460 436 -460 0 net=3953
rlabel metal2 33 -462 33 -462 0 net=2778
rlabel metal2 44 -462 44 -462 0 net=2946
rlabel metal2 159 -462 159 -462 0 net=2614
rlabel metal2 408 -462 408 -462 0 net=2471
rlabel metal2 436 -462 436 -462 0 net=4180
rlabel metal2 37 -464 37 -464 0 net=2651
rlabel metal2 121 -464 121 -464 0 net=1814
rlabel metal2 163 -464 163 -464 0 net=1420
rlabel metal2 226 -464 226 -464 0 net=1319
rlabel metal2 226 -464 226 -464 0 net=1319
rlabel metal2 233 -464 233 -464 0 net=2139
rlabel metal2 359 -464 359 -464 0 net=2299
rlabel metal2 457 -464 457 -464 0 net=3686
rlabel metal2 576 -464 576 -464 0 net=2915
rlabel metal2 44 -466 44 -466 0 net=2279
rlabel metal2 163 -466 163 -466 0 net=1628
rlabel metal2 387 -466 387 -466 0 net=2720
rlabel metal2 478 -466 478 -466 0 net=3319
rlabel metal2 576 -466 576 -466 0 net=4185
rlabel metal2 51 -468 51 -468 0 net=2196
rlabel metal2 219 -468 219 -468 0 net=2397
rlabel metal2 243 -468 243 -468 0 net=3823
rlabel metal2 597 -468 597 -468 0 net=4143
rlabel metal2 2 -470 2 -470 0 net=3124
rlabel metal2 247 -470 247 -470 0 net=4091
rlabel metal2 485 -470 485 -470 0 net=3335
rlabel metal2 51 -472 51 -472 0 net=1241
rlabel metal2 121 -472 121 -472 0 net=2015
rlabel metal2 275 -472 275 -472 0 net=1811
rlabel metal2 397 -472 397 -472 0 net=4145
rlabel metal2 58 -474 58 -474 0 net=2258
rlabel metal2 166 -474 166 -474 0 net=2127
rlabel metal2 205 -474 205 -474 0 net=1505
rlabel metal2 254 -474 254 -474 0 net=1162
rlabel metal2 296 -474 296 -474 0 net=1667
rlabel metal2 58 -476 58 -476 0 net=3281
rlabel metal2 429 -476 429 -476 0 net=2885
rlabel metal2 632 -476 632 -476 0 net=1717
rlabel metal2 65 -478 65 -478 0 net=1042
rlabel metal2 429 -478 429 -478 0 net=2685
rlabel metal2 450 -478 450 -478 0 net=3347
rlabel metal2 590 -478 590 -478 0 net=4163
rlabel metal2 65 -480 65 -480 0 net=3916
rlabel metal2 72 -482 72 -482 0 net=2540
rlabel metal2 212 -482 212 -482 0 net=1543
rlabel metal2 268 -482 268 -482 0 net=1065
rlabel metal2 345 -482 345 -482 0 net=2045
rlabel metal2 548 -482 548 -482 0 net=4043
rlabel metal2 72 -484 72 -484 0 net=1261
rlabel metal2 177 -484 177 -484 0 net=2027
rlabel metal2 215 -484 215 -484 0 net=119
rlabel metal2 390 -484 390 -484 0 net=2593
rlabel metal2 79 -486 79 -486 0 net=3703
rlabel metal2 79 -488 79 -488 0 net=1137
rlabel metal2 100 -488 100 -488 0 net=2229
rlabel metal2 282 -488 282 -488 0 net=3653
rlabel metal2 86 -490 86 -490 0 net=2515
rlabel metal2 128 -490 128 -490 0 net=2389
rlabel metal2 282 -490 282 -490 0 net=2085
rlabel metal2 352 -490 352 -490 0 net=3485
rlabel metal2 310 -492 310 -492 0 net=2241
rlabel metal2 380 -494 380 -494 0 net=3847
rlabel metal2 5 -505 5 -505 0 net=329
rlabel metal2 198 -505 198 -505 0 net=32
rlabel metal2 366 -505 366 -505 0 net=2093
rlabel metal2 618 -505 618 -505 0 net=2916
rlabel metal2 632 -505 632 -505 0 net=1719
rlabel metal2 632 -505 632 -505 0 net=1719
rlabel metal2 653 -505 653 -505 0 net=4284
rlabel metal2 681 -505 681 -505 0 net=3209
rlabel metal2 9 -507 9 -507 0 net=4294
rlabel metal2 121 -507 121 -507 0 net=2017
rlabel metal2 152 -507 152 -507 0 net=1812
rlabel metal2 285 -507 285 -507 0 net=3848
rlabel metal2 583 -507 583 -507 0 net=4353
rlabel metal2 628 -507 628 -507 0 net=4200
rlabel metal2 660 -507 660 -507 0 net=2553
rlabel metal2 660 -507 660 -507 0 net=2553
rlabel metal2 667 -507 667 -507 0 net=4337
rlabel metal2 9 -509 9 -509 0 net=3925
rlabel metal2 65 -509 65 -509 0 net=2517
rlabel metal2 93 -509 93 -509 0 net=2230
rlabel metal2 121 -509 121 -509 0 net=4093
rlabel metal2 254 -509 254 -509 0 net=1545
rlabel metal2 254 -509 254 -509 0 net=1545
rlabel metal2 268 -509 268 -509 0 net=1669
rlabel metal2 310 -509 310 -509 0 net=2242
rlabel metal2 383 -509 383 -509 0 net=3824
rlabel metal2 499 -509 499 -509 0 net=3918
rlabel metal2 604 -509 604 -509 0 net=78
rlabel metal2 618 -509 618 -509 0 net=4023
rlabel metal2 23 -511 23 -511 0 net=3558
rlabel metal2 68 -511 68 -511 0 net=586
rlabel metal2 219 -511 219 -511 0 net=1506
rlabel metal2 289 -511 289 -511 0 net=1066
rlabel metal2 338 -511 338 -511 0 net=2450
rlabel metal2 369 -511 369 -511 0 net=4261
rlabel metal2 639 -511 639 -511 0 net=4165
rlabel metal2 23 -513 23 -513 0 net=3567
rlabel metal2 243 -513 243 -513 0 net=3320
rlabel metal2 576 -513 576 -513 0 net=4187
rlabel metal2 30 -515 30 -515 0 net=3168
rlabel metal2 212 -515 212 -515 0 net=1321
rlabel metal2 243 -515 243 -515 0 net=3977
rlabel metal2 390 -515 390 -515 0 net=3954
rlabel metal2 555 -515 555 -515 0 net=4063
rlabel metal2 30 -517 30 -517 0 net=2947
rlabel metal2 278 -517 278 -517 0 net=3829
rlabel metal2 37 -519 37 -519 0 net=2652
rlabel metal2 163 -519 163 -519 0 net=2155
rlabel metal2 450 -519 450 -519 0 net=3487
rlabel metal2 502 -519 502 -519 0 net=3606
rlabel metal2 37 -521 37 -521 0 net=2251
rlabel metal2 149 -521 149 -521 0 net=3577
rlabel metal2 292 -521 292 -521 0 net=1307
rlabel metal2 478 -521 478 -521 0 net=3943
rlabel metal2 16 -523 16 -523 0 net=4032
rlabel metal2 156 -523 156 -523 0 net=2399
rlabel metal2 296 -523 296 -523 0 net=2141
rlabel metal2 331 -523 331 -523 0 net=3533
rlabel metal2 16 -525 16 -525 0 net=1043
rlabel metal2 86 -525 86 -525 0 net=2887
rlabel metal2 114 -525 114 -525 0 net=3869
rlabel metal2 44 -527 44 -527 0 net=2280
rlabel metal2 303 -527 303 -527 0 net=1553
rlabel metal2 341 -527 341 -527 0 net=3419
rlabel metal2 457 -527 457 -527 0 net=2886
rlabel metal2 485 -527 485 -527 0 net=4147
rlabel metal2 44 -529 44 -529 0 net=3085
rlabel metal2 324 -529 324 -529 0 net=2047
rlabel metal2 373 -529 373 -529 0 net=3172
rlabel metal2 397 -529 397 -529 0 net=4144
rlabel metal2 72 -531 72 -531 0 net=1262
rlabel metal2 170 -531 170 -531 0 net=1771
rlabel metal2 345 -531 345 -531 0 net=2519
rlabel metal2 415 -531 415 -531 0 net=3336
rlabel metal2 548 -531 548 -531 0 net=4045
rlabel metal2 51 -533 51 -533 0 net=1242
rlabel metal2 93 -533 93 -533 0 net=2391
rlabel metal2 205 -533 205 -533 0 net=1547
rlabel metal2 359 -533 359 -533 0 net=2301
rlabel metal2 415 -533 415 -533 0 net=2687
rlabel metal2 471 -533 471 -533 0 net=3349
rlabel metal2 499 -533 499 -533 0 net=3635
rlabel metal2 534 -533 534 -533 0 net=3749
rlabel metal2 51 -535 51 -535 0 net=1139
rlabel metal2 107 -535 107 -535 0 net=1027
rlabel metal2 170 -535 170 -535 0 net=2087
rlabel metal2 401 -535 401 -535 0 net=3283
rlabel metal2 506 -535 506 -535 0 net=3629
rlabel metal2 107 -537 107 -537 0 net=2129
rlabel metal2 208 -537 208 -537 0 net=3025
rlabel metal2 464 -537 464 -537 0 net=3655
rlabel metal2 261 -539 261 -539 0 net=1101
rlabel metal2 422 -539 422 -539 0 net=3705
rlabel metal2 128 -541 128 -541 0 net=3239
rlabel metal2 355 -541 355 -541 0 net=3107
rlabel metal2 513 -541 513 -541 0 net=3291
rlabel metal2 131 -543 131 -543 0 net=213
rlabel metal2 313 -543 313 -543 0 net=3509
rlabel metal2 159 -545 159 -545 0 net=3443
rlabel metal2 355 -545 355 -545 0 net=2472
rlabel metal2 177 -547 177 -547 0 net=2029
rlabel metal2 408 -547 408 -547 0 net=2595
rlabel metal2 317 -549 317 -549 0 net=2491
rlabel metal2 271 -551 271 -551 0 net=615
rlabel metal2 2 -562 2 -562 0 net=1671
rlabel metal2 275 -562 275 -562 0 net=363
rlabel metal2 345 -562 345 -562 0 net=2699
rlabel metal2 436 -562 436 -562 0 net=1308
rlabel metal2 646 -562 646 -562 0 net=4024
rlabel metal2 670 -562 670 -562 0 net=512
rlabel metal2 688 -562 688 -562 0 net=3210
rlabel metal2 688 -562 688 -562 0 net=3210
rlabel metal2 19 -564 19 -564 0 net=935
rlabel metal2 310 -564 310 -564 0 net=2302
rlabel metal2 401 -564 401 -564 0 net=1720
rlabel metal2 653 -564 653 -564 0 net=4167
rlabel metal2 674 -564 674 -564 0 net=4338
rlabel metal2 23 -566 23 -566 0 net=3568
rlabel metal2 107 -566 107 -566 0 net=2130
rlabel metal2 296 -566 296 -566 0 net=2142
rlabel metal2 380 -566 380 -566 0 net=2521
rlabel metal2 404 -566 404 -566 0 net=4046
rlabel metal2 618 -566 618 -566 0 net=4087
rlabel metal2 653 -566 653 -566 0 net=2554
rlabel metal2 23 -568 23 -568 0 net=4095
rlabel metal2 128 -568 128 -568 0 net=3578
rlabel metal2 233 -568 233 -568 0 net=1549
rlabel metal2 278 -568 278 -568 0 net=3534
rlabel metal2 576 -568 576 -568 0 net=3871
rlabel metal2 576 -568 576 -568 0 net=3871
rlabel metal2 590 -568 590 -568 0 net=4189
rlabel metal2 9 -570 9 -570 0 net=3926
rlabel metal2 131 -570 131 -570 0 net=4262
rlabel metal2 9 -572 9 -572 0 net=4355
rlabel metal2 180 -572 180 -572 0 net=3284
rlabel metal2 478 -572 478 -572 0 net=4113
rlabel metal2 604 -572 604 -572 0 net=4151
rlabel metal2 30 -574 30 -574 0 net=2948
rlabel metal2 107 -574 107 -574 0 net=2089
rlabel metal2 243 -574 243 -574 0 net=3706
rlabel metal2 30 -576 30 -576 0 net=3889
rlabel metal2 247 -576 247 -576 0 net=2018
rlabel metal2 383 -576 383 -576 0 net=3157
rlabel metal2 499 -576 499 -576 0 net=3293
rlabel metal2 534 -576 534 -576 0 net=3657
rlabel metal2 562 -576 562 -576 0 net=4065
rlabel metal2 37 -578 37 -578 0 net=2252
rlabel metal2 345 -578 345 -578 0 net=2111
rlabel metal2 355 -578 355 -578 0 net=2492
rlabel metal2 457 -578 457 -578 0 net=3488
rlabel metal2 40 -580 40 -580 0 net=324
rlabel metal2 184 -580 184 -580 0 net=3445
rlabel metal2 254 -580 254 -580 0 net=1546
rlabel metal2 485 -580 485 -580 0 net=3351
rlabel metal2 44 -582 44 -582 0 net=3086
rlabel metal2 149 -582 149 -582 0 net=2877
rlabel metal2 149 -582 149 -582 0 net=2877
rlabel metal2 163 -582 163 -582 0 net=2157
rlabel metal2 285 -582 285 -582 0 net=2899
rlabel metal2 366 -582 366 -582 0 net=2094
rlabel metal2 387 -582 387 -582 0 net=3979
rlabel metal2 51 -584 51 -584 0 net=1140
rlabel metal2 65 -584 65 -584 0 net=2518
rlabel metal2 93 -584 93 -584 0 net=2393
rlabel metal2 317 -584 317 -584 0 net=3944
rlabel metal2 16 -586 16 -586 0 net=1044
rlabel metal2 100 -586 100 -586 0 net=14
rlabel metal2 121 -586 121 -586 0 net=2231
rlabel metal2 212 -586 212 -586 0 net=1323
rlabel metal2 289 -586 289 -586 0 net=3569
rlabel metal2 548 -586 548 -586 0 net=3751
rlabel metal2 51 -588 51 -588 0 net=2889
rlabel metal2 114 -588 114 -588 0 net=2400
rlabel metal2 163 -588 163 -588 0 net=1772
rlabel metal2 236 -588 236 -588 0 net=1857
rlabel metal2 366 -588 366 -588 0 net=4263
rlabel metal2 58 -590 58 -590 0 net=2975
rlabel metal2 131 -590 131 -590 0 net=530
rlabel metal2 289 -590 289 -590 0 net=2159
rlabel metal2 471 -590 471 -590 0 net=4354
rlabel metal2 656 -590 656 -590 0 net=1
rlabel metal2 65 -592 65 -592 0 net=3125
rlabel metal2 135 -592 135 -592 0 net=1028
rlabel metal2 198 -592 198 -592 0 net=2031
rlabel metal2 282 -592 282 -592 0 net=1555
rlabel metal2 373 -592 373 -592 0 net=2891
rlabel metal2 485 -592 485 -592 0 net=3511
rlabel metal2 583 -592 583 -592 0 net=4149
rlabel metal2 75 -594 75 -594 0 net=1761
rlabel metal2 359 -594 359 -594 0 net=3927
rlabel metal2 79 -596 79 -596 0 net=1523
rlabel metal2 198 -596 198 -596 0 net=1247
rlabel metal2 303 -596 303 -596 0 net=3830
rlabel metal2 135 -598 135 -598 0 net=1103
rlabel metal2 359 -598 359 -598 0 net=3097
rlabel metal2 429 -598 429 -598 0 net=3027
rlabel metal2 460 -598 460 -598 0 net=3141
rlabel metal2 527 -598 527 -598 0 net=3637
rlabel metal2 142 -600 142 -600 0 net=2271
rlabel metal2 205 -600 205 -600 0 net=2731
rlabel metal2 450 -600 450 -600 0 net=3421
rlabel metal2 170 -602 170 -602 0 net=1221
rlabel metal2 205 -602 205 -602 0 net=1421
rlabel metal2 373 -602 373 -602 0 net=2315
rlabel metal2 408 -602 408 -602 0 net=2597
rlabel metal2 408 -602 408 -602 0 net=2597
rlabel metal2 415 -602 415 -602 0 net=2689
rlabel metal2 415 -602 415 -602 0 net=2689
rlabel metal2 450 -602 450 -602 0 net=3108
rlabel metal2 506 -602 506 -602 0 net=3631
rlabel metal2 212 -604 212 -604 0 net=2217
rlabel metal2 331 -604 331 -604 0 net=3241
rlabel metal2 324 -606 324 -606 0 net=2049
rlabel metal2 387 -606 387 -606 0 net=2829
rlabel metal2 464 -606 464 -606 0 net=3831
rlabel metal2 72 -608 72 -608 0 net=3405
rlabel metal2 2 -619 2 -619 0 net=1672
rlabel metal2 411 -619 411 -619 0 net=4114
rlabel metal2 632 -619 632 -619 0 net=4265
rlabel metal2 716 -619 716 -619 0 net=4277
rlabel metal2 2 -621 2 -621 0 net=3311
rlabel metal2 51 -621 51 -621 0 net=2890
rlabel metal2 159 -621 159 -621 0 net=3446
rlabel metal2 285 -621 285 -621 0 net=3045
rlabel metal2 492 -621 492 -621 0 net=4066
rlabel metal2 653 -621 653 -621 0 net=4168
rlabel metal2 681 -621 681 -621 0 net=1129
rlabel metal2 695 -621 695 -621 0 net=3457
rlabel metal2 9 -623 9 -623 0 net=4356
rlabel metal2 194 -623 194 -623 0 net=2160
rlabel metal2 296 -623 296 -623 0 net=2394
rlabel metal2 355 -623 355 -623 0 net=3098
rlabel metal2 376 -623 376 -623 0 net=3142
rlabel metal2 527 -623 527 -623 0 net=3423
rlabel metal2 618 -623 618 -623 0 net=4089
rlabel metal2 9 -625 9 -625 0 net=3265
rlabel metal2 93 -625 93 -625 0 net=846
rlabel metal2 107 -625 107 -625 0 net=2091
rlabel metal2 380 -625 380 -625 0 net=4297
rlabel metal2 23 -627 23 -627 0 net=4096
rlabel metal2 107 -627 107 -627 0 net=2879
rlabel metal2 166 -627 166 -627 0 net=1201
rlabel metal2 177 -627 177 -627 0 net=303
rlabel metal2 390 -627 390 -627 0 net=3872
rlabel metal2 583 -627 583 -627 0 net=3929
rlabel metal2 23 -629 23 -629 0 net=3109
rlabel metal2 177 -629 177 -629 0 net=2219
rlabel metal2 226 -629 226 -629 0 net=2033
rlabel metal2 289 -629 289 -629 0 net=2317
rlabel metal2 383 -629 383 -629 0 net=3752
rlabel metal2 30 -631 30 -631 0 net=3890
rlabel metal2 394 -631 394 -631 0 net=2599
rlabel metal2 425 -631 425 -631 0 net=3632
rlabel metal2 562 -631 562 -631 0 net=3833
rlabel metal2 30 -633 30 -633 0 net=2361
rlabel metal2 184 -633 184 -633 0 net=539
rlabel metal2 317 -633 317 -633 0 net=1859
rlabel metal2 317 -633 317 -633 0 net=1859
rlabel metal2 331 -633 331 -633 0 net=2051
rlabel metal2 331 -633 331 -633 0 net=2051
rlabel metal2 345 -633 345 -633 0 net=2113
rlabel metal2 453 -633 453 -633 0 net=4119
rlabel metal2 16 -635 16 -635 0 net=921
rlabel metal2 345 -635 345 -635 0 net=2923
rlabel metal2 495 -635 495 -635 0 net=3255
rlabel metal2 37 -637 37 -637 0 net=1539
rlabel metal2 65 -637 65 -637 0 net=3127
rlabel metal2 65 -637 65 -637 0 net=3127
rlabel metal2 72 -637 72 -637 0 net=2233
rlabel metal2 128 -637 128 -637 0 net=675
rlabel metal2 212 -637 212 -637 0 net=2158
rlabel metal2 240 -637 240 -637 0 net=1324
rlabel metal2 366 -637 366 -637 0 net=4249
rlabel metal2 44 -639 44 -639 0 net=1363
rlabel metal2 93 -639 93 -639 0 net=3215
rlabel metal2 541 -639 541 -639 0 net=3659
rlabel metal2 54 -641 54 -641 0 net=2311
rlabel metal2 303 -641 303 -641 0 net=2665
rlabel metal2 369 -641 369 -641 0 net=3638
rlabel metal2 58 -643 58 -643 0 net=2976
rlabel metal2 114 -643 114 -643 0 net=2101
rlabel metal2 240 -643 240 -643 0 net=1550
rlabel metal2 324 -643 324 -643 0 net=3407
rlabel metal2 117 -645 117 -645 0 net=834
rlabel metal2 229 -645 229 -645 0 net=2331
rlabel metal2 324 -645 324 -645 0 net=2523
rlabel metal2 453 -645 453 -645 0 net=3563
rlabel metal2 121 -647 121 -647 0 net=1997
rlabel metal2 149 -647 149 -647 0 net=1423
rlabel metal2 243 -647 243 -647 0 net=1556
rlabel metal2 310 -647 310 -647 0 net=1763
rlabel metal2 464 -647 464 -647 0 net=4150
rlabel metal2 79 -649 79 -649 0 net=1525
rlabel metal2 387 -649 387 -649 0 net=1311
rlabel metal2 474 -649 474 -649 0 net=4007
rlabel metal2 79 -651 79 -651 0 net=2005
rlabel metal2 135 -651 135 -651 0 net=1105
rlabel metal2 282 -651 282 -651 0 net=3375
rlabel metal2 142 -653 142 -653 0 net=2273
rlabel metal2 506 -653 506 -653 0 net=3243
rlabel metal2 534 -653 534 -653 0 net=3571
rlabel metal2 142 -655 142 -655 0 net=3512
rlabel metal2 499 -655 499 -655 0 net=3295
rlabel metal2 156 -657 156 -657 0 net=1801
rlabel metal2 243 -657 243 -657 0 net=3089
rlabel metal2 513 -657 513 -657 0 net=3353
rlabel metal2 198 -659 198 -659 0 net=1249
rlabel metal2 338 -659 338 -659 0 net=2901
rlabel metal2 135 -661 135 -661 0 net=1287
rlabel metal2 457 -661 457 -661 0 net=3029
rlabel metal2 191 -663 191 -663 0 net=1223
rlabel metal2 457 -663 457 -663 0 net=4190
rlabel metal2 191 -665 191 -665 0 net=670
rlabel metal2 478 -667 478 -667 0 net=3159
rlabel metal2 625 -667 625 -667 0 net=4153
rlabel metal2 443 -669 443 -669 0 net=2893
rlabel metal2 597 -669 597 -669 0 net=3981
rlabel metal2 299 -671 299 -671 0 net=3945
rlabel metal2 429 -673 429 -673 0 net=2733
rlabel metal2 415 -675 415 -675 0 net=2691
rlabel metal2 415 -677 415 -677 0 net=2831
rlabel metal2 422 -679 422 -679 0 net=2701
rlabel metal2 422 -681 422 -681 0 net=3671
rlabel metal2 2 -692 2 -692 0 net=3312
rlabel metal2 82 -692 82 -692 0 net=2702
rlabel metal2 450 -692 450 -692 0 net=3354
rlabel metal2 632 -692 632 -692 0 net=3565
rlabel metal2 730 -692 730 -692 0 net=4278
rlabel metal2 800 -692 800 -692 0 net=3381
rlabel metal2 9 -694 9 -694 0 net=3266
rlabel metal2 215 -694 215 -694 0 net=1526
rlabel metal2 341 -694 341 -694 0 net=3046
rlabel metal2 478 -694 478 -694 0 net=2895
rlabel metal2 478 -694 478 -694 0 net=2895
rlabel metal2 534 -694 534 -694 0 net=3297
rlabel metal2 16 -696 16 -696 0 net=2525
rlabel metal2 345 -696 345 -696 0 net=3244
rlabel metal2 674 -696 674 -696 0 net=3458
rlabel metal2 702 -696 702 -696 0 net=4267
rlabel metal2 19 -698 19 -698 0 net=413
rlabel metal2 121 -698 121 -698 0 net=1999
rlabel metal2 219 -698 219 -698 0 net=1107
rlabel metal2 219 -698 219 -698 0 net=1107
rlabel metal2 226 -698 226 -698 0 net=2034
rlabel metal2 278 -698 278 -698 0 net=3376
rlabel metal2 653 -698 653 -698 0 net=4299
rlabel metal2 9 -700 9 -700 0 net=3387
rlabel metal2 236 -700 236 -700 0 net=637
rlabel metal2 464 -700 464 -700 0 net=3572
rlabel metal2 646 -700 646 -700 0 net=4155
rlabel metal2 23 -702 23 -702 0 net=3110
rlabel metal2 254 -702 254 -702 0 net=2312
rlabel metal2 422 -702 422 -702 0 net=1130
rlabel metal2 23 -704 23 -704 0 net=2669
rlabel metal2 201 -704 201 -704 0 net=3935
rlabel metal2 429 -704 429 -704 0 net=2693
rlabel metal2 499 -704 499 -704 0 net=3031
rlabel metal2 569 -704 569 -704 0 net=4251
rlabel metal2 30 -706 30 -706 0 net=2362
rlabel metal2 254 -706 254 -706 0 net=2319
rlabel metal2 296 -706 296 -706 0 net=1764
rlabel metal2 408 -706 408 -706 0 net=3983
rlabel metal2 30 -708 30 -708 0 net=2253
rlabel metal2 100 -708 100 -708 0 net=1312
rlabel metal2 401 -708 401 -708 0 net=2177
rlabel metal2 467 -708 467 -708 0 net=4343
rlabel metal2 576 -708 576 -708 0 net=3673
rlabel metal2 37 -710 37 -710 0 net=1540
rlabel metal2 93 -710 93 -710 0 net=1803
rlabel metal2 240 -710 240 -710 0 net=2541
rlabel metal2 432 -710 432 -710 0 net=3982
rlabel metal2 2 -712 2 -712 0 net=3543
rlabel metal2 100 -712 100 -712 0 net=683
rlabel metal2 40 -714 40 -714 0 net=2666
rlabel metal2 310 -714 310 -714 0 net=2053
rlabel metal2 352 -714 352 -714 0 net=2092
rlabel metal2 366 -714 366 -714 0 net=3930
rlabel metal2 44 -716 44 -716 0 net=1364
rlabel metal2 233 -716 233 -716 0 net=1877
rlabel metal2 359 -716 359 -716 0 net=4229
rlabel metal2 44 -718 44 -718 0 net=1781
rlabel metal2 128 -718 128 -718 0 net=2007
rlabel metal2 128 -718 128 -718 0 net=2007
rlabel metal2 135 -718 135 -718 0 net=1037
rlabel metal2 247 -718 247 -718 0 net=2274
rlabel metal2 373 -718 373 -718 0 net=4157
rlabel metal2 408 -718 408 -718 0 net=3424
rlabel metal2 58 -720 58 -720 0 net=3129
rlabel metal2 72 -720 72 -720 0 net=2235
rlabel metal2 72 -720 72 -720 0 net=2235
rlabel metal2 142 -720 142 -720 0 net=3377
rlabel metal2 317 -720 317 -720 0 net=1861
rlabel metal2 373 -720 373 -720 0 net=3019
rlabel metal2 548 -720 548 -720 0 net=3257
rlabel metal2 583 -720 583 -720 0 net=3731
rlabel metal2 65 -722 65 -722 0 net=2601
rlabel metal2 415 -722 415 -722 0 net=2833
rlabel metal2 562 -722 562 -722 0 net=3661
rlabel metal2 142 -724 142 -724 0 net=1285
rlabel metal2 296 -724 296 -724 0 net=2121
rlabel metal2 436 -724 436 -724 0 net=3217
rlabel metal2 565 -724 565 -724 0 net=4257
rlabel metal2 149 -726 149 -726 0 net=1425
rlabel metal2 247 -726 247 -726 0 net=4120
rlabel metal2 114 -728 114 -728 0 net=2103
rlabel metal2 156 -728 156 -728 0 net=1175
rlabel metal2 443 -728 443 -728 0 net=2735
rlabel metal2 492 -728 492 -728 0 net=2925
rlabel metal2 590 -728 590 -728 0 net=3835
rlabel metal2 114 -730 114 -730 0 net=1251
rlabel metal2 261 -730 261 -730 0 net=1609
rlabel metal2 184 -732 184 -732 0 net=1533
rlabel metal2 278 -732 278 -732 0 net=179
rlabel metal2 331 -732 331 -732 0 net=2115
rlabel metal2 450 -732 450 -732 0 net=2637
rlabel metal2 492 -732 492 -732 0 net=3263
rlabel metal2 597 -732 597 -732 0 net=3947
rlabel metal2 639 -732 639 -732 0 net=4009
rlabel metal2 170 -734 170 -734 0 net=1203
rlabel metal2 191 -734 191 -734 0 net=2333
rlabel metal2 299 -734 299 -734 0 net=1224
rlabel metal2 348 -734 348 -734 0 net=2407
rlabel metal2 453 -734 453 -734 0 net=4090
rlabel metal2 107 -736 107 -736 0 net=2881
rlabel metal2 317 -736 317 -736 0 net=1561
rlabel metal2 366 -736 366 -736 0 net=2653
rlabel metal2 107 -738 107 -738 0 net=2221
rlabel metal2 243 -738 243 -738 0 net=3745
rlabel metal2 170 -740 170 -740 0 net=1289
rlabel metal2 376 -740 376 -740 0 net=2871
rlabel metal2 506 -740 506 -740 0 net=3091
rlabel metal2 555 -740 555 -740 0 net=3409
rlabel metal2 51 -742 51 -742 0 net=3707
rlabel metal2 380 -742 380 -742 0 net=4253
rlabel metal2 177 -744 177 -744 0 net=1479
rlabel metal2 485 -746 485 -746 0 net=2903
rlabel metal2 513 -746 513 -746 0 net=3161
rlabel metal2 485 -748 485 -748 0 net=3451
rlabel metal2 30 -759 30 -759 0 net=2254
rlabel metal2 429 -759 429 -759 0 net=1589
rlabel metal2 807 -759 807 -759 0 net=3383
rlabel metal2 807 -759 807 -759 0 net=3383
rlabel metal2 30 -761 30 -761 0 net=332
rlabel metal2 89 -761 89 -761 0 net=2104
rlabel metal2 177 -761 177 -761 0 net=1480
rlabel metal2 243 -761 243 -761 0 net=2203
rlabel metal2 289 -761 289 -761 0 net=2054
rlabel metal2 327 -761 327 -761 0 net=3746
rlabel metal2 674 -761 674 -761 0 net=4231
rlabel metal2 733 -761 733 -761 0 net=4268
rlabel metal2 2 -763 2 -763 0 net=3544
rlabel metal2 107 -763 107 -763 0 net=2222
rlabel metal2 226 -763 226 -763 0 net=1862
rlabel metal2 387 -763 387 -763 0 net=3298
rlabel metal2 723 -763 723 -763 0 net=3566
rlabel metal2 23 -765 23 -765 0 net=2670
rlabel metal2 390 -765 390 -765 0 net=3264
rlabel metal2 604 -765 604 -765 0 net=4259
rlabel metal2 23 -767 23 -767 0 net=19
rlabel metal2 58 -767 58 -767 0 net=3130
rlabel metal2 100 -767 100 -767 0 net=467
rlabel metal2 121 -767 121 -767 0 net=173
rlabel metal2 142 -767 142 -767 0 net=1286
rlabel metal2 299 -767 299 -767 0 net=2209
rlabel metal2 422 -767 422 -767 0 net=3937
rlabel metal2 37 -769 37 -769 0 net=1805
rlabel metal2 100 -769 100 -769 0 net=2321
rlabel metal2 261 -769 261 -769 0 net=1611
rlabel metal2 334 -769 334 -769 0 net=3452
rlabel metal2 527 -769 527 -769 0 net=3662
rlabel metal2 632 -769 632 -769 0 net=3985
rlabel metal2 51 -771 51 -771 0 net=3709
rlabel metal2 702 -771 702 -771 0 net=4255
rlabel metal2 58 -773 58 -773 0 net=2335
rlabel metal2 247 -773 247 -773 0 net=2151
rlabel metal2 341 -773 341 -773 0 net=2872
rlabel metal2 495 -773 495 -773 0 net=3836
rlabel metal2 712 -773 712 -773 0 net=4359
rlabel metal2 65 -775 65 -775 0 net=2602
rlabel metal2 390 -775 390 -775 0 net=2409
rlabel metal2 436 -775 436 -775 0 net=3219
rlabel metal2 65 -777 65 -777 0 net=1513
rlabel metal2 93 -777 93 -777 0 net=1173
rlabel metal2 345 -777 345 -777 0 net=1879
rlabel metal2 373 -777 373 -777 0 net=3021
rlabel metal2 541 -777 541 -777 0 net=4156
rlabel metal2 72 -779 72 -779 0 net=2236
rlabel metal2 121 -779 121 -779 0 net=4135
rlabel metal2 72 -781 72 -781 0 net=1045
rlabel metal2 247 -781 247 -781 0 net=1563
rlabel metal2 352 -781 352 -781 0 net=1869
rlabel metal2 439 -781 439 -781 0 net=1007
rlabel metal2 79 -783 79 -783 0 net=790
rlabel metal2 303 -783 303 -783 0 net=3379
rlabel metal2 124 -785 124 -785 0 net=2000
rlabel metal2 170 -785 170 -785 0 net=1291
rlabel metal2 373 -785 373 -785 0 net=2589
rlabel metal2 383 -785 383 -785 0 net=4295
rlabel metal2 2 -787 2 -787 0 net=2481
rlabel metal2 170 -787 170 -787 0 net=1163
rlabel metal2 303 -787 303 -787 0 net=2117
rlabel metal2 380 -787 380 -787 0 net=3071
rlabel metal2 611 -787 611 -787 0 net=3675
rlabel metal2 632 -787 632 -787 0 net=4011
rlabel metal2 9 -789 9 -789 0 net=3388
rlabel metal2 149 -789 149 -789 0 net=2543
rlabel metal2 394 -789 394 -789 0 net=1941
rlabel metal2 464 -789 464 -789 0 net=2695
rlabel metal2 544 -789 544 -789 0 net=3789
rlabel metal2 9 -791 9 -791 0 net=2009
rlabel metal2 156 -791 156 -791 0 net=1177
rlabel metal2 240 -791 240 -791 0 net=4369
rlabel metal2 16 -793 16 -793 0 net=2526
rlabel metal2 362 -793 362 -793 0 net=3553
rlabel metal2 488 -793 488 -793 0 net=2991
rlabel metal2 16 -795 16 -795 0 net=1039
rlabel metal2 156 -795 156 -795 0 net=2067
rlabel metal2 397 -795 397 -795 0 net=697
rlabel metal2 453 -795 453 -795 0 net=3711
rlabel metal2 44 -797 44 -797 0 net=1782
rlabel metal2 177 -797 177 -797 0 net=2387
rlabel metal2 212 -797 212 -797 0 net=1427
rlabel metal2 366 -797 366 -797 0 net=2655
rlabel metal2 548 -797 548 -797 0 net=2926
rlabel metal2 586 -797 586 -797 0 net=4252
rlabel metal2 44 -799 44 -799 0 net=2647
rlabel metal2 404 -799 404 -799 0 net=4329
rlabel metal2 590 -799 590 -799 0 net=3411
rlabel metal2 618 -799 618 -799 0 net=3949
rlabel metal2 128 -801 128 -801 0 net=1109
rlabel metal2 222 -801 222 -801 0 net=3513
rlabel metal2 411 -801 411 -801 0 net=2959
rlabel metal2 534 -801 534 -801 0 net=3033
rlabel metal2 681 -801 681 -801 0 net=3733
rlabel metal2 103 -803 103 -803 0 net=2667
rlabel metal2 555 -803 555 -803 0 net=3163
rlabel metal2 184 -805 184 -805 0 net=1204
rlabel metal2 219 -805 219 -805 0 net=2882
rlabel metal2 415 -805 415 -805 0 net=2408
rlabel metal2 520 -805 520 -805 0 net=3093
rlabel metal2 562 -805 562 -805 0 net=4300
rlabel metal2 114 -807 114 -807 0 net=1253
rlabel metal2 198 -807 198 -807 0 net=4158
rlabel metal2 695 -807 695 -807 0 net=3785
rlabel metal2 110 -809 110 -809 0 net=1629
rlabel metal2 233 -809 233 -809 0 net=1919
rlabel metal2 436 -809 436 -809 0 net=3593
rlabel metal2 205 -811 205 -811 0 net=1535
rlabel metal2 268 -811 268 -811 0 net=2179
rlabel metal2 499 -811 499 -811 0 net=2835
rlabel metal2 569 -811 569 -811 0 net=4345
rlabel metal2 205 -813 205 -813 0 net=1145
rlabel metal2 359 -813 359 -813 0 net=3225
rlabel metal2 576 -813 576 -813 0 net=3259
rlabel metal2 296 -815 296 -815 0 net=2123
rlabel metal2 499 -815 499 -815 0 net=2905
rlabel metal2 520 -815 520 -815 0 net=153
rlabel metal2 296 -817 296 -817 0 net=2721
rlabel metal2 471 -819 471 -819 0 net=2639
rlabel metal2 523 -819 523 -819 0 net=3101
rlabel metal2 457 -821 457 -821 0 net=2737
rlabel metal2 530 -821 530 -821 0 net=3439
rlabel metal2 457 -823 457 -823 0 net=2896
rlabel metal2 478 -825 478 -825 0 net=2569
rlabel metal2 9 -836 9 -836 0 net=2010
rlabel metal2 278 -836 278 -836 0 net=4370
rlabel metal2 803 -836 803 -836 0 net=3384
rlabel metal2 9 -838 9 -838 0 net=2545
rlabel metal2 159 -838 159 -838 0 net=199
rlabel metal2 460 -838 460 -838 0 net=4260
rlabel metal2 16 -840 16 -840 0 net=1040
rlabel metal2 184 -840 184 -840 0 net=1254
rlabel metal2 366 -840 366 -840 0 net=1920
rlabel metal2 439 -840 439 -840 0 net=4346
rlabel metal2 16 -842 16 -842 0 net=3099
rlabel metal2 184 -842 184 -842 0 net=1871
rlabel metal2 359 -842 359 -842 0 net=2125
rlabel metal2 460 -842 460 -842 0 net=3938
rlabel metal2 751 -842 751 -842 0 net=1590
rlabel metal2 23 -844 23 -844 0 net=2971
rlabel metal2 149 -844 149 -844 0 net=768
rlabel metal2 404 -844 404 -844 0 net=2836
rlabel metal2 625 -844 625 -844 0 net=3677
rlabel metal2 625 -844 625 -844 0 net=3677
rlabel metal2 688 -844 688 -844 0 net=3735
rlabel metal2 688 -844 688 -844 0 net=3735
rlabel metal2 730 -844 730 -844 0 net=4233
rlabel metal2 751 -844 751 -844 0 net=4313
rlabel metal2 30 -846 30 -846 0 net=2969
rlabel metal2 240 -846 240 -846 0 net=1564
rlabel metal2 268 -846 268 -846 0 net=2181
rlabel metal2 366 -846 366 -846 0 net=1837
rlabel metal2 390 -846 390 -846 0 net=4360
rlabel metal2 37 -848 37 -848 0 net=1806
rlabel metal2 107 -848 107 -848 0 net=2069
rlabel metal2 166 -848 166 -848 0 net=632
rlabel metal2 215 -848 215 -848 0 net=3710
rlabel metal2 716 -848 716 -848 0 net=4137
rlabel metal2 786 -848 786 -848 0 net=3067
rlabel metal2 44 -850 44 -850 0 net=2648
rlabel metal2 142 -850 142 -850 0 net=1099
rlabel metal2 142 -850 142 -850 0 net=1099
rlabel metal2 156 -850 156 -850 0 net=2668
rlabel metal2 667 -850 667 -850 0 net=3713
rlabel metal2 54 -852 54 -852 0 net=4296
rlabel metal2 58 -854 58 -854 0 net=2336
rlabel metal2 338 -854 338 -854 0 net=3515
rlabel metal2 72 -856 72 -856 0 net=1047
rlabel metal2 268 -856 268 -856 0 net=1429
rlabel metal2 373 -856 373 -856 0 net=2591
rlabel metal2 646 -856 646 -856 0 net=2992
rlabel metal2 51 -858 51 -858 0 net=1889
rlabel metal2 82 -858 82 -858 0 net=1008
rlabel metal2 128 -860 128 -860 0 net=1111
rlabel metal2 219 -860 219 -860 0 net=943
rlabel metal2 275 -860 275 -860 0 net=2205
rlabel metal2 383 -860 383 -860 0 net=4341
rlabel metal2 2 -862 2 -862 0 net=2482
rlabel metal2 282 -862 282 -862 0 net=1255
rlabel metal2 397 -862 397 -862 0 net=3072
rlabel metal2 44 -864 44 -864 0 net=1219
rlabel metal2 135 -864 135 -864 0 net=2861
rlabel metal2 467 -864 467 -864 0 net=3164
rlabel metal2 170 -866 170 -866 0 net=1165
rlabel metal2 201 -866 201 -866 0 net=2427
rlabel metal2 401 -866 401 -866 0 net=1785
rlabel metal2 418 -866 418 -866 0 net=3034
rlabel metal2 93 -868 93 -868 0 net=1174
rlabel metal2 205 -868 205 -868 0 net=1147
rlabel metal2 205 -868 205 -868 0 net=1147
rlabel metal2 226 -868 226 -868 0 net=1179
rlabel metal2 292 -868 292 -868 0 net=4139
rlabel metal2 58 -870 58 -870 0 net=1009
rlabel metal2 229 -870 229 -870 0 net=3440
rlabel metal2 93 -872 93 -872 0 net=1631
rlabel metal2 170 -872 170 -872 0 net=2152
rlabel metal2 282 -872 282 -872 0 net=1753
rlabel metal2 411 -872 411 -872 0 net=3389
rlabel metal2 114 -874 114 -874 0 net=1193
rlabel metal2 177 -874 177 -874 0 net=2388
rlabel metal2 233 -874 233 -874 0 net=1537
rlabel metal2 296 -874 296 -874 0 net=1293
rlabel metal2 334 -874 334 -874 0 net=3285
rlabel metal2 488 -874 488 -874 0 net=3790
rlabel metal2 37 -876 37 -876 0 net=2405
rlabel metal2 303 -876 303 -876 0 net=2119
rlabel metal2 348 -876 348 -876 0 net=3817
rlabel metal2 65 -878 65 -878 0 net=1515
rlabel metal2 177 -878 177 -878 0 net=3380
rlabel metal2 65 -880 65 -880 0 net=2147
rlabel metal2 303 -880 303 -880 0 net=1943
rlabel metal2 422 -880 422 -880 0 net=2411
rlabel metal2 506 -880 506 -880 0 net=2641
rlabel metal2 523 -880 523 -880 0 net=3986
rlabel metal2 324 -882 324 -882 0 net=1613
rlabel metal2 488 -882 488 -882 0 net=3220
rlabel metal2 191 -884 191 -884 0 net=1273
rlabel metal2 394 -884 394 -884 0 net=2696
rlabel metal2 569 -884 569 -884 0 net=3227
rlabel metal2 653 -884 653 -884 0 net=3787
rlabel metal2 450 -886 450 -886 0 net=2657
rlabel metal2 576 -886 576 -886 0 net=3103
rlabel metal2 611 -886 611 -886 0 net=3261
rlabel metal2 695 -886 695 -886 0 net=3951
rlabel metal2 450 -888 450 -888 0 net=4256
rlabel metal2 464 -890 464 -890 0 net=3555
rlabel metal2 618 -890 618 -890 0 net=4013
rlabel metal2 152 -892 152 -892 0 net=3115
rlabel metal2 464 -894 464 -894 0 net=2493
rlabel metal2 583 -894 583 -894 0 net=4331
rlabel metal2 495 -896 495 -896 0 net=3795
rlabel metal2 499 -898 499 -898 0 net=2907
rlabel metal2 513 -898 513 -898 0 net=3023
rlabel metal2 583 -898 583 -898 0 net=3413
rlabel metal2 478 -900 478 -900 0 net=2571
rlabel metal2 527 -900 527 -900 0 net=4269
rlabel metal2 100 -902 100 -902 0 net=2323
rlabel metal2 499 -902 499 -902 0 net=3131
rlabel metal2 79 -904 79 -904 0 net=3313
rlabel metal2 443 -904 443 -904 0 net=2961
rlabel metal2 530 -904 530 -904 0 net=2722
rlabel metal2 590 -904 590 -904 0 net=3595
rlabel metal2 79 -906 79 -906 0 net=1881
rlabel metal2 485 -906 485 -906 0 net=2727
rlabel metal2 555 -906 555 -906 0 net=3095
rlabel metal2 331 -908 331 -908 0 net=2143
rlabel metal2 471 -908 471 -908 0 net=2739
rlabel metal2 331 -910 331 -910 0 net=1185
rlabel metal2 408 -910 408 -910 0 net=2211
rlabel metal2 408 -912 408 -912 0 net=4077
rlabel metal2 9 -923 9 -923 0 net=2546
rlabel metal2 229 -923 229 -923 0 net=2206
rlabel metal2 348 -923 348 -923 0 net=3556
rlabel metal2 688 -923 688 -923 0 net=3737
rlabel metal2 688 -923 688 -923 0 net=3737
rlabel metal2 723 -923 723 -923 0 net=4078
rlabel metal2 779 -923 779 -923 0 net=3068
rlabel metal2 9 -925 9 -925 0 net=2183
rlabel metal2 366 -925 366 -925 0 net=2144
rlabel metal2 446 -925 446 -925 0 net=4138
rlabel metal2 751 -925 751 -925 0 net=4314
rlabel metal2 16 -927 16 -927 0 net=3100
rlabel metal2 121 -927 121 -927 0 net=1517
rlabel metal2 142 -927 142 -927 0 net=1100
rlabel metal2 159 -927 159 -927 0 net=981
rlabel metal2 432 -927 432 -927 0 net=2572
rlabel metal2 548 -927 548 -927 0 net=2729
rlabel metal2 548 -927 548 -927 0 net=2729
rlabel metal2 576 -927 576 -927 0 net=4245
rlabel metal2 16 -929 16 -929 0 net=3315
rlabel metal2 107 -929 107 -929 0 net=2071
rlabel metal2 149 -929 149 -929 0 net=1754
rlabel metal2 408 -929 408 -929 0 net=2592
rlabel metal2 576 -929 576 -929 0 net=3229
rlabel metal2 723 -929 723 -929 0 net=4221
rlabel metal2 23 -931 23 -931 0 net=2972
rlabel metal2 236 -931 236 -931 0 net=3788
rlabel metal2 23 -933 23 -933 0 net=1875
rlabel metal2 107 -933 107 -933 0 net=1697
rlabel metal2 285 -933 285 -933 0 net=1614
rlabel metal2 460 -933 460 -933 0 net=4234
rlabel metal2 30 -935 30 -935 0 net=2970
rlabel metal2 415 -935 415 -935 0 net=3761
rlabel metal2 499 -935 499 -935 0 net=3952
rlabel metal2 30 -937 30 -937 0 net=1873
rlabel metal2 191 -937 191 -937 0 net=919
rlabel metal2 201 -937 201 -937 0 net=67
rlabel metal2 513 -937 513 -937 0 net=2741
rlabel metal2 579 -937 579 -937 0 net=3104
rlabel metal2 681 -937 681 -937 0 net=3262
rlabel metal2 37 -939 37 -939 0 net=2406
rlabel metal2 86 -939 86 -939 0 net=272
rlabel metal2 275 -939 275 -939 0 net=1945
rlabel metal2 310 -939 310 -939 0 net=2120
rlabel metal2 317 -939 317 -939 0 net=1256
rlabel metal2 418 -939 418 -939 0 net=3096
rlabel metal2 604 -939 604 -939 0 net=3679
rlabel metal2 674 -939 674 -939 0 net=3715
rlabel metal2 37 -941 37 -941 0 net=1731
rlabel metal2 86 -941 86 -941 0 net=1157
rlabel metal2 114 -941 114 -941 0 net=1195
rlabel metal2 135 -941 135 -941 0 net=2862
rlabel metal2 243 -941 243 -941 0 net=1538
rlabel metal2 296 -941 296 -941 0 net=1295
rlabel metal2 348 -941 348 -941 0 net=1786
rlabel metal2 418 -941 418 -941 0 net=2401
rlabel metal2 527 -941 527 -941 0 net=2963
rlabel metal2 44 -943 44 -943 0 net=1220
rlabel metal2 464 -943 464 -943 0 net=4342
rlabel metal2 51 -945 51 -945 0 net=1890
rlabel metal2 114 -945 114 -945 0 net=3643
rlabel metal2 51 -947 51 -947 0 net=1633
rlabel metal2 149 -947 149 -947 0 net=1973
rlabel metal2 359 -947 359 -947 0 net=2429
rlabel metal2 467 -947 467 -947 0 net=4270
rlabel metal2 65 -949 65 -949 0 net=1181
rlabel metal2 397 -949 397 -949 0 net=2126
rlabel metal2 471 -949 471 -949 0 net=2213
rlabel metal2 618 -949 618 -949 0 net=4015
rlabel metal2 79 -951 79 -951 0 net=1883
rlabel metal2 163 -951 163 -951 0 net=2149
rlabel metal2 488 -951 488 -951 0 net=3765
rlabel metal2 44 -953 44 -953 0 net=1541
rlabel metal2 89 -953 89 -953 0 net=3024
rlabel metal2 590 -953 590 -953 0 net=3597
rlabel metal2 163 -955 163 -955 0 net=1113
rlabel metal2 226 -955 226 -955 0 net=1527
rlabel metal2 429 -955 429 -955 0 net=3287
rlabel metal2 597 -955 597 -955 0 net=3391
rlabel metal2 58 -957 58 -957 0 net=1010
rlabel metal2 506 -957 506 -957 0 net=2909
rlabel metal2 618 -957 618 -957 0 net=3473
rlabel metal2 58 -959 58 -959 0 net=1773
rlabel metal2 478 -959 478 -959 0 net=2325
rlabel metal2 520 -959 520 -959 0 net=2643
rlabel metal2 534 -959 534 -959 0 net=4332
rlabel metal2 170 -961 170 -961 0 net=1483
rlabel metal2 457 -961 457 -961 0 net=3299
rlabel metal2 555 -961 555 -961 0 net=2495
rlabel metal2 632 -961 632 -961 0 net=3117
rlabel metal2 177 -963 177 -963 0 net=1229
rlabel metal2 390 -963 390 -963 0 net=2779
rlabel metal2 583 -963 583 -963 0 net=3415
rlabel metal2 180 -965 180 -965 0 net=3447
rlabel metal2 457 -965 457 -965 0 net=2413
rlabel metal2 583 -965 583 -965 0 net=3133
rlabel metal2 184 -967 184 -967 0 net=1431
rlabel metal2 278 -967 278 -967 0 net=1155
rlabel metal2 191 -969 191 -969 0 net=1149
rlabel metal2 212 -969 212 -969 0 net=1279
rlabel metal2 226 -969 226 -969 0 net=1083
rlabel metal2 471 -969 471 -969 0 net=2629
rlabel metal2 639 -969 639 -969 0 net=3517
rlabel metal2 205 -971 205 -971 0 net=2077
rlabel metal2 243 -971 243 -971 0 net=1186
rlabel metal2 492 -971 492 -971 0 net=2659
rlabel metal2 667 -971 667 -971 0 net=3797
rlabel metal2 198 -973 198 -973 0 net=1213
rlabel metal2 702 -973 702 -973 0 net=3819
rlabel metal2 219 -975 219 -975 0 net=2563
rlabel metal2 268 -975 268 -975 0 net=1275
rlabel metal2 709 -975 709 -975 0 net=4141
rlabel metal2 247 -977 247 -977 0 net=1048
rlabel metal2 394 -977 394 -977 0 net=3987
rlabel metal2 236 -979 236 -979 0 net=2011
rlabel metal2 254 -979 254 -979 0 net=1166
rlabel metal2 254 -981 254 -981 0 net=2785
rlabel metal2 289 -983 289 -983 0 net=2173
rlabel metal2 296 -985 296 -985 0 net=1965
rlabel metal2 310 -987 310 -987 0 net=2373
rlabel metal2 324 -989 324 -989 0 net=1839
rlabel metal2 9 -1000 9 -1000 0 net=2184
rlabel metal2 334 -1000 334 -1000 0 net=2150
rlabel metal2 411 -1000 411 -1000 0 net=2742
rlabel metal2 604 -1000 604 -1000 0 net=3681
rlabel metal2 604 -1000 604 -1000 0 net=3681
rlabel metal2 688 -1000 688 -1000 0 net=3738
rlabel metal2 688 -1000 688 -1000 0 net=3738
rlabel metal2 737 -1000 737 -1000 0 net=147
rlabel metal2 16 -1002 16 -1002 0 net=3316
rlabel metal2 198 -1002 198 -1002 0 net=848
rlabel metal2 373 -1002 373 -1002 0 net=3367
rlabel metal2 394 -1002 394 -1002 0 net=2577
rlabel metal2 408 -1002 408 -1002 0 net=2813
rlabel metal2 471 -1002 471 -1002 0 net=4016
rlabel metal2 740 -1002 740 -1002 0 net=1156
rlabel metal2 23 -1004 23 -1004 0 net=1876
rlabel metal2 243 -1004 243 -1004 0 net=2457
rlabel metal2 362 -1004 362 -1004 0 net=3230
rlabel metal2 23 -1006 23 -1006 0 net=1975
rlabel metal2 166 -1006 166 -1006 0 net=460
rlabel metal2 233 -1006 233 -1006 0 net=1214
rlabel metal2 338 -1006 338 -1006 0 net=1529
rlabel metal2 373 -1006 373 -1006 0 net=2497
rlabel metal2 576 -1006 576 -1006 0 net=2977
rlabel metal2 30 -1008 30 -1008 0 net=1874
rlabel metal2 250 -1008 250 -1008 0 net=2564
rlabel metal2 268 -1008 268 -1008 0 net=1277
rlabel metal2 338 -1008 338 -1008 0 net=2403
rlabel metal2 33 -1010 33 -1010 0 net=986
rlabel metal2 191 -1010 191 -1010 0 net=1150
rlabel metal2 247 -1010 247 -1010 0 net=2013
rlabel metal2 282 -1010 282 -1010 0 net=3518
rlabel metal2 37 -1012 37 -1012 0 net=1732
rlabel metal2 107 -1012 107 -1012 0 net=1698
rlabel metal2 345 -1012 345 -1012 0 net=4246
rlabel metal2 37 -1014 37 -1014 0 net=4219
rlabel metal2 114 -1014 114 -1014 0 net=715
rlabel metal2 44 -1016 44 -1016 0 net=1542
rlabel metal2 65 -1016 65 -1016 0 net=1183
rlabel metal2 114 -1016 114 -1016 0 net=1197
rlabel metal2 142 -1016 142 -1016 0 net=2072
rlabel metal2 170 -1016 170 -1016 0 net=1485
rlabel metal2 296 -1016 296 -1016 0 net=1967
rlabel metal2 348 -1016 348 -1016 0 net=236
rlabel metal2 443 -1016 443 -1016 0 net=2730
rlabel metal2 562 -1016 562 -1016 0 net=2911
rlabel metal2 51 -1018 51 -1018 0 net=1634
rlabel metal2 121 -1018 121 -1018 0 net=1433
rlabel metal2 205 -1018 205 -1018 0 net=2078
rlabel metal2 275 -1018 275 -1018 0 net=1947
rlabel metal2 303 -1018 303 -1018 0 net=1297
rlabel metal2 303 -1018 303 -1018 0 net=1297
rlabel metal2 352 -1018 352 -1018 0 net=3474
rlabel metal2 51 -1020 51 -1020 0 net=2607
rlabel metal2 135 -1020 135 -1020 0 net=1885
rlabel metal2 149 -1020 149 -1020 0 net=1647
rlabel metal2 352 -1020 352 -1020 0 net=1639
rlabel metal2 376 -1020 376 -1020 0 net=2326
rlabel metal2 590 -1020 590 -1020 0 net=3289
rlabel metal2 58 -1022 58 -1022 0 net=1775
rlabel metal2 191 -1022 191 -1022 0 net=1187
rlabel metal2 212 -1022 212 -1022 0 net=1281
rlabel metal2 380 -1022 380 -1022 0 net=3449
rlabel metal2 415 -1022 415 -1022 0 net=3118
rlabel metal2 65 -1024 65 -1024 0 net=2713
rlabel metal2 135 -1024 135 -1024 0 net=1331
rlabel metal2 163 -1024 163 -1024 0 net=1115
rlabel metal2 380 -1024 380 -1024 0 net=3135
rlabel metal2 590 -1024 590 -1024 0 net=3393
rlabel metal2 72 -1026 72 -1026 0 net=1158
rlabel metal2 170 -1026 170 -1026 0 net=1085
rlabel metal2 597 -1026 597 -1026 0 net=3645
rlabel metal2 44 -1028 44 -1028 0 net=3873
rlabel metal2 156 -1028 156 -1028 0 net=2167
rlabel metal2 310 -1028 310 -1028 0 net=3801
rlabel metal2 75 -1030 75 -1030 0 net=118
rlabel metal2 397 -1030 397 -1030 0 net=3739
rlabel metal2 79 -1032 79 -1032 0 net=1519
rlabel metal2 156 -1032 156 -1032 0 net=1231
rlabel metal2 418 -1032 418 -1032 0 net=2414
rlabel metal2 478 -1032 478 -1032 0 net=3301
rlabel metal2 128 -1034 128 -1034 0 net=2175
rlabel metal2 401 -1034 401 -1034 0 net=2431
rlabel metal2 478 -1034 478 -1034 0 net=4142
rlabel metal2 177 -1036 177 -1036 0 net=2711
rlabel metal2 289 -1036 289 -1036 0 net=1841
rlabel metal2 401 -1036 401 -1036 0 net=2964
rlabel metal2 646 -1036 646 -1036 0 net=3599
rlabel metal2 324 -1038 324 -1038 0 net=2631
rlabel metal2 625 -1038 625 -1038 0 net=3767
rlabel metal2 313 -1040 313 -1040 0 net=4067
rlabel metal2 212 -1042 212 -1042 0 net=2061
rlabel metal2 425 -1042 425 -1042 0 net=4169
rlabel metal2 432 -1044 432 -1044 0 net=3999
rlabel metal2 436 -1046 436 -1046 0 net=2375
rlabel metal2 446 -1046 446 -1046 0 net=2660
rlabel metal2 495 -1046 495 -1046 0 net=2847
rlabel metal2 520 -1046 520 -1046 0 net=995
rlabel metal2 646 -1046 646 -1046 0 net=3821
rlabel metal2 450 -1048 450 -1048 0 net=2214
rlabel metal2 702 -1048 702 -1048 0 net=4223
rlabel metal2 453 -1050 453 -1050 0 net=3798
rlabel metal2 467 -1052 467 -1052 0 net=1587
rlabel metal2 667 -1052 667 -1052 0 net=3989
rlabel metal2 485 -1054 485 -1054 0 net=3763
rlabel metal2 716 -1054 716 -1054 0 net=3615
rlabel metal2 278 -1056 278 -1056 0 net=3683
rlabel metal2 492 -1056 492 -1056 0 net=2780
rlabel metal2 499 -1058 499 -1058 0 net=2645
rlabel metal2 541 -1058 541 -1058 0 net=2787
rlabel metal2 425 -1060 425 -1060 0 net=2965
rlabel metal2 569 -1060 569 -1060 0 net=3417
rlabel metal2 429 -1062 429 -1062 0 net=2223
rlabel metal2 632 -1062 632 -1062 0 net=3717
rlabel metal2 681 -1064 681 -1064 0 net=4275
rlabel metal2 9 -1075 9 -1075 0 net=1435
rlabel metal2 128 -1075 128 -1075 0 net=2176
rlabel metal2 243 -1075 243 -1075 0 net=38
rlabel metal2 387 -1075 387 -1075 0 net=3450
rlabel metal2 418 -1075 418 -1075 0 net=4170
rlabel metal2 677 -1075 677 -1075 0 net=4235
rlabel metal2 702 -1075 702 -1075 0 net=4225
rlabel metal2 702 -1075 702 -1075 0 net=4225
rlabel metal2 16 -1077 16 -1077 0 net=2897
rlabel metal2 37 -1077 37 -1077 0 net=4220
rlabel metal2 187 -1077 187 -1077 0 net=2014
rlabel metal2 278 -1077 278 -1077 0 net=1298
rlabel metal2 313 -1077 313 -1077 0 net=1977
rlabel metal2 415 -1077 415 -1077 0 net=2433
rlabel metal2 478 -1077 478 -1077 0 net=569
rlabel metal2 44 -1079 44 -1079 0 net=3874
rlabel metal2 128 -1079 128 -1079 0 net=2063
rlabel metal2 254 -1079 254 -1079 0 net=1116
rlabel metal2 324 -1079 324 -1079 0 net=2632
rlabel metal2 394 -1079 394 -1079 0 net=2579
rlabel metal2 443 -1079 443 -1079 0 net=2377
rlabel metal2 443 -1079 443 -1079 0 net=2377
rlabel metal2 485 -1079 485 -1079 0 net=3684
rlabel metal2 51 -1081 51 -1081 0 net=2608
rlabel metal2 166 -1081 166 -1081 0 net=648
rlabel metal2 282 -1081 282 -1081 0 net=1283
rlabel metal2 310 -1081 310 -1081 0 net=4276
rlabel metal2 51 -1083 51 -1083 0 net=3933
rlabel metal2 86 -1083 86 -1083 0 net=2073
rlabel metal2 282 -1083 282 -1083 0 net=1531
rlabel metal2 401 -1083 401 -1083 0 net=3007
rlabel metal2 495 -1083 495 -1083 0 net=3718
rlabel metal2 65 -1085 65 -1085 0 net=2714
rlabel metal2 194 -1085 194 -1085 0 net=1278
rlabel metal2 324 -1085 324 -1085 0 net=1657
rlabel metal2 352 -1085 352 -1085 0 net=1641
rlabel metal2 352 -1085 352 -1085 0 net=1641
rlabel metal2 359 -1085 359 -1085 0 net=2459
rlabel metal2 464 -1085 464 -1085 0 net=2815
rlabel metal2 499 -1085 499 -1085 0 net=2646
rlabel metal2 527 -1085 527 -1085 0 net=2967
rlabel metal2 527 -1085 527 -1085 0 net=2967
rlabel metal2 534 -1085 534 -1085 0 net=3394
rlabel metal2 611 -1085 611 -1085 0 net=1588
rlabel metal2 58 -1087 58 -1087 0 net=1309
rlabel metal2 72 -1087 72 -1087 0 net=1233
rlabel metal2 177 -1087 177 -1087 0 net=1583
rlabel metal2 289 -1087 289 -1087 0 net=1843
rlabel metal2 334 -1087 334 -1087 0 net=3290
rlabel metal2 632 -1087 632 -1087 0 net=4001
rlabel metal2 79 -1089 79 -1089 0 net=1520
rlabel metal2 198 -1089 198 -1089 0 net=2404
rlabel metal2 345 -1089 345 -1089 0 net=1969
rlabel metal2 422 -1089 422 -1089 0 net=2912
rlabel metal2 23 -1091 23 -1091 0 net=1976
rlabel metal2 289 -1091 289 -1091 0 net=2225
rlabel metal2 439 -1091 439 -1091 0 net=3791
rlabel metal2 506 -1091 506 -1091 0 net=3418
rlabel metal2 583 -1091 583 -1091 0 net=3741
rlabel metal2 611 -1091 611 -1091 0 net=3991
rlabel metal2 93 -1093 93 -1093 0 net=1184
rlabel metal2 422 -1093 422 -1093 0 net=2793
rlabel metal2 513 -1093 513 -1093 0 net=2849
rlabel metal2 537 -1093 537 -1093 0 net=784
rlabel metal2 37 -1095 37 -1095 0 net=1341
rlabel metal2 100 -1095 100 -1095 0 net=1887
rlabel metal2 145 -1095 145 -1095 0 net=1299
rlabel metal2 268 -1095 268 -1095 0 net=2712
rlabel metal2 453 -1095 453 -1095 0 net=4371
rlabel metal2 107 -1097 107 -1097 0 net=1087
rlabel metal2 268 -1097 268 -1097 0 net=1117
rlabel metal2 513 -1097 513 -1097 0 net=2979
rlabel metal2 583 -1097 583 -1097 0 net=3647
rlabel metal2 618 -1097 618 -1097 0 net=4069
rlabel metal2 114 -1099 114 -1099 0 net=1199
rlabel metal2 114 -1099 114 -1099 0 net=1199
rlabel metal2 135 -1099 135 -1099 0 net=1332
rlabel metal2 296 -1099 296 -1099 0 net=1948
rlabel metal2 523 -1099 523 -1099 0 net=4305
rlabel metal2 576 -1099 576 -1099 0 net=2789
rlabel metal2 135 -1101 135 -1101 0 net=2169
rlabel metal2 296 -1101 296 -1101 0 net=1305
rlabel metal2 565 -1101 565 -1101 0 net=3682
rlabel metal2 684 -1101 684 -1101 0 net=2753
rlabel metal2 142 -1103 142 -1103 0 net=3136
rlabel metal2 523 -1103 523 -1103 0 net=4335
rlabel metal2 149 -1105 149 -1105 0 net=1649
rlabel metal2 275 -1105 275 -1105 0 net=3897
rlabel metal2 184 -1107 184 -1107 0 net=1777
rlabel metal2 338 -1107 338 -1107 0 net=1933
rlabel metal2 541 -1107 541 -1107 0 net=3822
rlabel metal2 23 -1109 23 -1109 0 net=3309
rlabel metal2 219 -1109 219 -1109 0 net=1487
rlabel metal2 247 -1109 247 -1109 0 net=3489
rlabel metal2 555 -1109 555 -1109 0 net=3369
rlabel metal2 597 -1109 597 -1109 0 net=3803
rlabel metal2 68 -1111 68 -1111 0 net=4333
rlabel metal2 205 -1113 205 -1113 0 net=1189
rlabel metal2 373 -1113 373 -1113 0 net=2499
rlabel metal2 548 -1113 548 -1113 0 net=3303
rlabel metal2 205 -1115 205 -1115 0 net=1829
rlabel metal2 380 -1115 380 -1115 0 net=3764
rlabel metal2 376 -1117 376 -1117 0 net=4327
rlabel metal2 425 -1119 425 -1119 0 net=3691
rlabel metal2 548 -1119 548 -1119 0 net=3769
rlabel metal2 425 -1121 425 -1121 0 net=3600
rlabel metal2 450 -1123 450 -1123 0 net=4115
rlabel metal2 709 -1123 709 -1123 0 net=3617
rlabel metal2 411 -1125 411 -1125 0 net=2703
rlabel metal2 474 -1125 474 -1125 0 net=3169
rlabel metal2 2 -1136 2 -1136 0 net=2065
rlabel metal2 145 -1136 145 -1136 0 net=13
rlabel metal2 159 -1136 159 -1136 0 net=1118
rlabel metal2 275 -1136 275 -1136 0 net=1306
rlabel metal2 303 -1136 303 -1136 0 net=1284
rlabel metal2 317 -1136 317 -1136 0 net=1845
rlabel metal2 369 -1136 369 -1136 0 net=4328
rlabel metal2 646 -1136 646 -1136 0 net=4334
rlabel metal2 677 -1136 677 -1136 0 net=3618
rlabel metal2 9 -1138 9 -1138 0 net=1436
rlabel metal2 170 -1138 170 -1138 0 net=3370
rlabel metal2 646 -1138 646 -1138 0 net=4117
rlabel metal2 677 -1138 677 -1138 0 net=3435
rlabel metal2 688 -1138 688 -1138 0 net=4237
rlabel metal2 688 -1138 688 -1138 0 net=4237
rlabel metal2 695 -1138 695 -1138 0 net=2755
rlabel metal2 9 -1140 9 -1140 0 net=3005
rlabel metal2 250 -1140 250 -1140 0 net=2460
rlabel metal2 464 -1140 464 -1140 0 net=2500
rlabel metal2 464 -1140 464 -1140 0 net=2500
rlabel metal2 506 -1140 506 -1140 0 net=3323
rlabel metal2 523 -1140 523 -1140 0 net=2968
rlabel metal2 530 -1140 530 -1140 0 net=2850
rlabel metal2 544 -1140 544 -1140 0 net=4079
rlabel metal2 702 -1140 702 -1140 0 net=4227
rlabel metal2 702 -1140 702 -1140 0 net=4227
rlabel metal2 16 -1142 16 -1142 0 net=2898
rlabel metal2 47 -1142 47 -1142 0 net=1310
rlabel metal2 72 -1142 72 -1142 0 net=1234
rlabel metal2 219 -1142 219 -1142 0 net=1191
rlabel metal2 261 -1142 261 -1142 0 net=1584
rlabel metal2 380 -1142 380 -1142 0 net=1971
rlabel metal2 429 -1142 429 -1142 0 net=3304
rlabel metal2 562 -1142 562 -1142 0 net=4071
rlabel metal2 37 -1144 37 -1144 0 net=1342
rlabel metal2 79 -1144 79 -1144 0 net=1621
rlabel metal2 334 -1144 334 -1144 0 net=2378
rlabel metal2 478 -1144 478 -1144 0 net=3009
rlabel metal2 590 -1144 590 -1144 0 net=3743
rlabel metal2 37 -1146 37 -1146 0 net=1405
rlabel metal2 331 -1146 331 -1146 0 net=3490
rlabel metal2 583 -1146 583 -1146 0 net=3649
rlabel metal2 44 -1148 44 -1148 0 net=2573
rlabel metal2 226 -1148 226 -1148 0 net=1779
rlabel metal2 278 -1148 278 -1148 0 net=3170
rlabel metal2 51 -1150 51 -1150 0 net=3934
rlabel metal2 93 -1150 93 -1150 0 net=482
rlabel metal2 184 -1150 184 -1150 0 net=1300
rlabel metal2 282 -1150 282 -1150 0 net=1532
rlabel metal2 429 -1150 429 -1150 0 net=2581
rlabel metal2 471 -1150 471 -1150 0 net=2795
rlabel metal2 492 -1150 492 -1150 0 net=2981
rlabel metal2 541 -1150 541 -1150 0 net=3693
rlabel metal2 604 -1150 604 -1150 0 net=3899
rlabel metal2 51 -1152 51 -1152 0 net=1651
rlabel metal2 156 -1152 156 -1152 0 net=3189
rlabel metal2 289 -1152 289 -1152 0 net=2227
rlabel metal2 289 -1152 289 -1152 0 net=2227
rlabel metal2 310 -1152 310 -1152 0 net=1659
rlabel metal2 345 -1152 345 -1152 0 net=3792
rlabel metal2 19 -1154 19 -1154 0 net=858
rlabel metal2 348 -1154 348 -1154 0 net=4306
rlabel metal2 58 -1156 58 -1156 0 net=1831
rlabel metal2 226 -1156 226 -1156 0 net=1353
rlabel metal2 317 -1156 317 -1156 0 net=4372
rlabel metal2 82 -1158 82 -1158 0 net=1755
rlabel metal2 100 -1158 100 -1158 0 net=1888
rlabel metal2 205 -1158 205 -1158 0 net=1685
rlabel metal2 233 -1158 233 -1158 0 net=1489
rlabel metal2 348 -1158 348 -1158 0 net=1642
rlabel metal2 373 -1158 373 -1158 0 net=1979
rlabel metal2 415 -1158 415 -1158 0 net=2435
rlabel metal2 432 -1158 432 -1158 0 net=3777
rlabel metal2 569 -1158 569 -1158 0 net=4003
rlabel metal2 660 -1158 660 -1158 0 net=4336
rlabel metal2 86 -1160 86 -1160 0 net=2075
rlabel metal2 387 -1160 387 -1160 0 net=2313
rlabel metal2 443 -1160 443 -1160 0 net=3729
rlabel metal2 632 -1160 632 -1160 0 net=3975
rlabel metal2 30 -1162 30 -1162 0 net=1921
rlabel metal2 107 -1162 107 -1162 0 net=1088
rlabel metal2 236 -1162 236 -1162 0 net=1637
rlabel metal2 394 -1162 394 -1162 0 net=2583
rlabel metal2 450 -1162 450 -1162 0 net=2705
rlabel metal2 485 -1162 485 -1162 0 net=2817
rlabel metal2 107 -1164 107 -1164 0 net=1200
rlabel metal2 121 -1164 121 -1164 0 net=709
rlabel metal2 362 -1164 362 -1164 0 net=3539
rlabel metal2 397 -1164 397 -1164 0 net=2790
rlabel metal2 23 -1166 23 -1166 0 net=3310
rlabel metal2 121 -1166 121 -1166 0 net=1935
rlabel metal2 387 -1166 387 -1166 0 net=3547
rlabel metal2 110 -1168 110 -1168 0 net=2363
rlabel metal2 135 -1168 135 -1168 0 net=2171
rlabel metal2 450 -1168 450 -1168 0 net=3770
rlabel metal2 135 -1170 135 -1170 0 net=3525
rlabel metal2 156 -1170 156 -1170 0 net=1699
rlabel metal2 184 -1170 184 -1170 0 net=1663
rlabel metal2 338 -1170 338 -1170 0 net=3361
rlabel metal2 548 -1170 548 -1170 0 net=3805
rlabel metal2 142 -1172 142 -1172 0 net=4311
rlabel metal2 142 -1174 142 -1174 0 net=2709
rlabel metal2 485 -1174 485 -1174 0 net=2751
rlabel metal2 145 -1176 145 -1176 0 net=150
rlabel metal2 597 -1176 597 -1176 0 net=3993
rlabel metal2 163 -1178 163 -1178 0 net=1899
rlabel metal2 173 -1178 173 -1178 0 net=1263
rlabel metal2 366 -1178 366 -1178 0 net=2603
rlabel metal2 446 -1178 446 -1178 0 net=3073
rlabel metal2 166 -1180 166 -1180 0 net=3545
rlabel metal2 191 -1182 191 -1182 0 net=1471
rlabel metal2 390 -1182 390 -1182 0 net=3911
rlabel metal2 2 -1193 2 -1193 0 net=2066
rlabel metal2 156 -1193 156 -1193 0 net=1901
rlabel metal2 166 -1193 166 -1193 0 net=305
rlabel metal2 201 -1193 201 -1193 0 net=241
rlabel metal2 275 -1193 275 -1193 0 net=1638
rlabel metal2 303 -1193 303 -1193 0 net=2582
rlabel metal2 436 -1193 436 -1193 0 net=3548
rlabel metal2 667 -1193 667 -1193 0 net=3437
rlabel metal2 702 -1193 702 -1193 0 net=4228
rlabel metal2 709 -1193 709 -1193 0 net=2757
rlabel metal2 2 -1195 2 -1195 0 net=2611
rlabel metal2 110 -1195 110 -1195 0 net=317
rlabel metal2 215 -1195 215 -1195 0 net=1192
rlabel metal2 296 -1195 296 -1195 0 net=3011
rlabel metal2 530 -1195 530 -1195 0 net=3976
rlabel metal2 674 -1195 674 -1195 0 net=4238
rlabel metal2 9 -1197 9 -1197 0 net=3006
rlabel metal2 30 -1197 30 -1197 0 net=1923
rlabel metal2 306 -1197 306 -1197 0 net=2172
rlabel metal2 359 -1197 359 -1197 0 net=1847
rlabel metal2 359 -1197 359 -1197 0 net=1847
rlabel metal2 383 -1197 383 -1197 0 net=3173
rlabel metal2 541 -1197 541 -1197 0 net=3650
rlabel metal2 597 -1197 597 -1197 0 net=3995
rlabel metal2 9 -1199 9 -1199 0 net=2575
rlabel metal2 54 -1199 54 -1199 0 net=701
rlabel metal2 229 -1199 229 -1199 0 net=2076
rlabel metal2 289 -1199 289 -1199 0 net=2228
rlabel metal2 310 -1199 310 -1199 0 net=1661
rlabel metal2 320 -1199 320 -1199 0 net=3651
rlabel metal2 16 -1201 16 -1201 0 net=2627
rlabel metal2 89 -1201 89 -1201 0 net=3324
rlabel metal2 562 -1201 562 -1201 0 net=4073
rlabel metal2 23 -1203 23 -1203 0 net=1407
rlabel metal2 198 -1203 198 -1203 0 net=1473
rlabel metal2 310 -1203 310 -1203 0 net=4357
rlabel metal2 30 -1205 30 -1205 0 net=2807
rlabel metal2 117 -1205 117 -1205 0 net=2314
rlabel metal2 436 -1205 436 -1205 0 net=2707
rlabel metal2 478 -1205 478 -1205 0 net=2797
rlabel metal2 562 -1205 562 -1205 0 net=3231
rlabel metal2 37 -1207 37 -1207 0 net=1406
rlabel metal2 142 -1207 142 -1207 0 net=2999
rlabel metal2 569 -1207 569 -1207 0 net=4005
rlabel metal2 37 -1209 37 -1209 0 net=1665
rlabel metal2 219 -1209 219 -1209 0 net=1687
rlabel metal2 324 -1209 324 -1209 0 net=1980
rlabel metal2 387 -1209 387 -1209 0 net=2436
rlabel metal2 443 -1209 443 -1209 0 net=3546
rlabel metal2 597 -1209 597 -1209 0 net=3075
rlabel metal2 58 -1211 58 -1211 0 net=1832
rlabel metal2 233 -1211 233 -1211 0 net=4312
rlabel metal2 58 -1213 58 -1213 0 net=1071
rlabel metal2 93 -1213 93 -1213 0 net=1757
rlabel metal2 93 -1213 93 -1213 0 net=1757
rlabel metal2 100 -1213 100 -1213 0 net=2710
rlabel metal2 460 -1213 460 -1213 0 net=3719
rlabel metal2 65 -1215 65 -1215 0 net=2135
rlabel metal2 100 -1215 100 -1215 0 net=2281
rlabel metal2 121 -1215 121 -1215 0 net=1937
rlabel metal2 240 -1215 240 -1215 0 net=1265
rlabel metal2 341 -1215 341 -1215 0 net=1972
rlabel metal2 387 -1215 387 -1215 0 net=1985
rlabel metal2 499 -1215 499 -1215 0 net=2819
rlabel metal2 548 -1215 548 -1215 0 net=3807
rlabel metal2 72 -1217 72 -1217 0 net=772
rlabel metal2 194 -1217 194 -1217 0 net=1387
rlabel metal2 247 -1217 247 -1217 0 net=3900
rlabel metal2 145 -1219 145 -1219 0 net=312
rlabel metal2 327 -1219 327 -1219 0 net=2752
rlabel metal2 513 -1219 513 -1219 0 net=3363
rlabel metal2 149 -1221 149 -1221 0 net=1701
rlabel metal2 254 -1221 254 -1221 0 net=3191
rlabel metal2 513 -1221 513 -1221 0 net=4209
rlabel metal2 51 -1223 51 -1223 0 net=1652
rlabel metal2 327 -1223 327 -1223 0 net=3730
rlabel metal2 334 -1225 334 -1225 0 net=2673
rlabel metal2 604 -1225 604 -1225 0 net=4081
rlabel metal2 348 -1227 348 -1227 0 net=3641
rlabel metal2 352 -1229 352 -1229 0 net=2633
rlabel metal2 583 -1229 583 -1229 0 net=3695
rlabel metal2 366 -1231 366 -1231 0 net=2605
rlabel metal2 429 -1231 429 -1231 0 net=3177
rlabel metal2 135 -1233 135 -1233 0 net=3527
rlabel metal2 373 -1233 373 -1233 0 net=2337
rlabel metal2 401 -1233 401 -1233 0 net=2585
rlabel metal2 432 -1233 432 -1233 0 net=2145
rlabel metal2 446 -1233 446 -1233 0 net=4047
rlabel metal2 79 -1235 79 -1235 0 net=1623
rlabel metal2 380 -1235 380 -1235 0 net=3744
rlabel metal2 79 -1237 79 -1237 0 net=2365
rlabel metal2 331 -1237 331 -1237 0 net=3401
rlabel metal2 128 -1239 128 -1239 0 net=1355
rlabel metal2 394 -1239 394 -1239 0 net=3541
rlabel metal2 226 -1241 226 -1241 0 net=1780
rlabel metal2 401 -1241 401 -1241 0 net=3035
rlabel metal2 534 -1241 534 -1241 0 net=3779
rlabel metal2 254 -1243 254 -1243 0 net=214
rlabel metal2 450 -1243 450 -1243 0 net=4118
rlabel metal2 261 -1245 261 -1245 0 net=1491
rlabel metal2 415 -1245 415 -1245 0 net=3913
rlabel metal2 170 -1247 170 -1247 0 net=1019
rlabel metal2 345 -1247 345 -1247 0 net=2285
rlabel metal2 450 -1247 450 -1247 0 net=1575
rlabel metal2 345 -1249 345 -1249 0 net=1709
rlabel metal2 453 -1249 453 -1249 0 net=2982
rlabel metal2 534 -1249 534 -1249 0 net=3151
rlabel metal2 457 -1251 457 -1251 0 net=2781
rlabel metal2 492 -1253 492 -1253 0 net=2985
rlabel metal2 16 -1264 16 -1264 0 net=2628
rlabel metal2 72 -1264 72 -1264 0 net=4358
rlabel metal2 712 -1264 712 -1264 0 net=2758
rlabel metal2 2 -1266 2 -1266 0 net=2612
rlabel metal2 93 -1266 93 -1266 0 net=1758
rlabel metal2 107 -1266 107 -1266 0 net=1463
rlabel metal2 317 -1266 317 -1266 0 net=1662
rlabel metal2 394 -1266 394 -1266 0 net=4006
rlabel metal2 2 -1268 2 -1268 0 net=1625
rlabel metal2 142 -1268 142 -1268 0 net=1903
rlabel metal2 177 -1268 177 -1268 0 net=826
rlabel metal2 254 -1268 254 -1268 0 net=1492
rlabel metal2 271 -1268 271 -1268 0 net=2986
rlabel metal2 667 -1268 667 -1268 0 net=3438
rlabel metal2 9 -1270 9 -1270 0 net=2576
rlabel metal2 145 -1270 145 -1270 0 net=1474
rlabel metal2 303 -1270 303 -1270 0 net=410
rlabel metal2 9 -1272 9 -1272 0 net=3105
rlabel metal2 194 -1272 194 -1272 0 net=3528
rlabel metal2 397 -1272 397 -1272 0 net=3542
rlabel metal2 667 -1272 667 -1272 0 net=1576
rlabel metal2 702 -1272 702 -1272 0 net=3467
rlabel metal2 23 -1274 23 -1274 0 net=1408
rlabel metal2 208 -1274 208 -1274 0 net=3
rlabel metal2 222 -1274 222 -1274 0 net=2771
rlabel metal2 257 -1274 257 -1274 0 net=1557
rlabel metal2 303 -1274 303 -1274 0 net=2146
rlabel metal2 460 -1274 460 -1274 0 net=3111
rlabel metal2 23 -1276 23 -1276 0 net=2367
rlabel metal2 86 -1276 86 -1276 0 net=1073
rlabel metal2 100 -1276 100 -1276 0 net=2283
rlabel metal2 128 -1276 128 -1276 0 net=1357
rlabel metal2 212 -1276 212 -1276 0 net=1089
rlabel metal2 212 -1276 212 -1276 0 net=1089
rlabel metal2 215 -1276 215 -1276 0 net=1266
rlabel metal2 345 -1276 345 -1276 0 net=1711
rlabel metal2 345 -1276 345 -1276 0 net=1711
rlabel metal2 352 -1276 352 -1276 0 net=3076
rlabel metal2 30 -1278 30 -1278 0 net=2809
rlabel metal2 114 -1278 114 -1278 0 net=1327
rlabel metal2 236 -1278 236 -1278 0 net=1171
rlabel metal2 324 -1278 324 -1278 0 net=2606
rlabel metal2 429 -1278 429 -1278 0 net=3153
rlabel metal2 576 -1278 576 -1278 0 net=3721
rlabel metal2 37 -1280 37 -1280 0 net=1666
rlabel metal2 362 -1280 362 -1280 0 net=2820
rlabel metal2 534 -1280 534 -1280 0 net=3809
rlabel metal2 569 -1280 569 -1280 0 net=3365
rlabel metal2 40 -1282 40 -1282 0 net=2136
rlabel metal2 131 -1282 131 -1282 0 net=137
rlabel metal2 240 -1282 240 -1282 0 net=1389
rlabel metal2 240 -1282 240 -1282 0 net=1389
rlabel metal2 285 -1282 285 -1282 0 net=3642
rlabel metal2 44 -1284 44 -1284 0 net=833
rlabel metal2 149 -1284 149 -1284 0 net=1703
rlabel metal2 177 -1284 177 -1284 0 net=3914
rlabel metal2 44 -1286 44 -1286 0 net=1939
rlabel metal2 219 -1286 219 -1286 0 net=1017
rlabel metal2 495 -1286 495 -1286 0 net=4191
rlabel metal2 47 -1288 47 -1288 0 net=2674
rlabel metal2 506 -1288 506 -1288 0 net=3001
rlabel metal2 51 -1290 51 -1290 0 net=2355
rlabel metal2 180 -1290 180 -1290 0 net=2105
rlabel metal2 226 -1290 226 -1290 0 net=1451
rlabel metal2 310 -1290 310 -1290 0 net=3753
rlabel metal2 366 -1290 366 -1290 0 net=3143
rlabel metal2 58 -1292 58 -1292 0 net=2987
rlabel metal2 163 -1292 163 -1292 0 net=1925
rlabel metal2 327 -1292 327 -1292 0 net=2927
rlabel metal2 380 -1292 380 -1292 0 net=3799
rlabel metal2 65 -1294 65 -1294 0 net=3307
rlabel metal2 233 -1294 233 -1294 0 net=25
rlabel metal2 478 -1294 478 -1294 0 net=3573
rlabel metal2 513 -1294 513 -1294 0 net=3696
rlabel metal2 121 -1296 121 -1296 0 net=1991
rlabel metal2 184 -1296 184 -1296 0 net=3012
rlabel metal2 380 -1296 380 -1296 0 net=2286
rlabel metal2 422 -1296 422 -1296 0 net=2587
rlabel metal2 639 -1296 639 -1296 0 net=4211
rlabel metal2 170 -1298 170 -1298 0 net=1021
rlabel metal2 247 -1298 247 -1298 0 net=3519
rlabel metal2 373 -1298 373 -1298 0 net=2339
rlabel metal2 432 -1298 432 -1298 0 net=2708
rlabel metal2 443 -1298 443 -1298 0 net=2615
rlabel metal2 520 -1298 520 -1298 0 net=3233
rlabel metal2 632 -1298 632 -1298 0 net=3652
rlabel metal2 268 -1300 268 -1300 0 net=750
rlabel metal2 436 -1300 436 -1300 0 net=3193
rlabel metal2 562 -1300 562 -1300 0 net=4083
rlabel metal2 268 -1302 268 -1302 0 net=1689
rlabel metal2 296 -1302 296 -1302 0 net=1986
rlabel metal2 397 -1302 397 -1302 0 net=2997
rlabel metal2 464 -1302 464 -1302 0 net=3175
rlabel metal2 261 -1304 261 -1304 0 net=1745
rlabel metal2 306 -1304 306 -1304 0 net=1848
rlabel metal2 373 -1304 373 -1304 0 net=3077
rlabel metal2 590 -1304 590 -1304 0 net=4049
rlabel metal2 275 -1306 275 -1306 0 net=1673
rlabel metal2 401 -1306 401 -1306 0 net=3037
rlabel metal2 324 -1308 324 -1308 0 net=3535
rlabel metal2 390 -1310 390 -1310 0 net=2267
rlabel metal2 408 -1310 408 -1310 0 net=2634
rlabel metal2 485 -1310 485 -1310 0 net=3179
rlabel metal2 464 -1312 464 -1312 0 net=3402
rlabel metal2 548 -1314 548 -1314 0 net=3781
rlabel metal2 618 -1314 618 -1314 0 net=4075
rlabel metal2 180 -1316 180 -1316 0 net=3955
rlabel metal2 499 -1318 499 -1318 0 net=2783
rlabel metal2 499 -1320 499 -1320 0 net=3996
rlabel metal2 541 -1322 541 -1322 0 net=2799
rlabel metal2 450 -1324 450 -1324 0 net=3325
rlabel metal2 2 -1335 2 -1335 0 net=1626
rlabel metal2 208 -1335 208 -1335 0 net=1690
rlabel metal2 303 -1335 303 -1335 0 net=2507
rlabel metal2 404 -1335 404 -1335 0 net=2998
rlabel metal2 460 -1335 460 -1335 0 net=3176
rlabel metal2 653 -1335 653 -1335 0 net=2784
rlabel metal2 702 -1335 702 -1335 0 net=3468
rlabel metal2 702 -1335 702 -1335 0 net=3468
rlabel metal2 9 -1337 9 -1337 0 net=3106
rlabel metal2 212 -1337 212 -1337 0 net=1090
rlabel metal2 338 -1337 338 -1337 0 net=3536
rlabel metal2 646 -1337 646 -1337 0 net=851
rlabel metal2 667 -1337 667 -1337 0 net=3003
rlabel metal2 19 -1339 19 -1339 0 net=1328
rlabel metal2 135 -1339 135 -1339 0 net=545
rlabel metal2 254 -1339 254 -1339 0 net=2772
rlabel metal2 366 -1339 366 -1339 0 net=3722
rlabel metal2 646 -1339 646 -1339 0 net=4217
rlabel metal2 33 -1341 33 -1341 0 net=591
rlabel metal2 138 -1341 138 -1341 0 net=865
rlabel metal2 338 -1341 338 -1341 0 net=2341
rlabel metal2 422 -1341 422 -1341 0 net=3366
rlabel metal2 590 -1341 590 -1341 0 net=4213
rlabel metal2 44 -1343 44 -1343 0 net=1940
rlabel metal2 373 -1343 373 -1343 0 net=3079
rlabel metal2 576 -1343 576 -1343 0 net=4051
rlabel metal2 51 -1345 51 -1345 0 net=2356
rlabel metal2 261 -1345 261 -1345 0 net=1747
rlabel metal2 275 -1345 275 -1345 0 net=1674
rlabel metal2 352 -1345 352 -1345 0 net=136
rlabel metal2 58 -1347 58 -1347 0 net=2988
rlabel metal2 86 -1347 86 -1347 0 net=2811
rlabel metal2 86 -1347 86 -1347 0 net=2811
rlabel metal2 100 -1347 100 -1347 0 net=2284
rlabel metal2 149 -1347 149 -1347 0 net=1705
rlabel metal2 159 -1347 159 -1347 0 net=98
rlabel metal2 366 -1347 366 -1347 0 net=2588
rlabel metal2 58 -1349 58 -1349 0 net=1927
rlabel metal2 177 -1349 177 -1349 0 net=1023
rlabel metal2 219 -1349 219 -1349 0 net=1018
rlabel metal2 380 -1349 380 -1349 0 net=2767
rlabel metal2 408 -1349 408 -1349 0 net=2845
rlabel metal2 37 -1351 37 -1351 0 net=4121
rlabel metal2 222 -1351 222 -1351 0 net=362
rlabel metal2 450 -1351 450 -1351 0 net=3327
rlabel metal2 51 -1353 51 -1353 0 net=3147
rlabel metal2 226 -1353 226 -1353 0 net=1453
rlabel metal2 261 -1353 261 -1353 0 net=1713
rlabel metal2 348 -1353 348 -1353 0 net=3453
rlabel metal2 425 -1353 425 -1353 0 net=3800
rlabel metal2 65 -1355 65 -1355 0 net=3308
rlabel metal2 383 -1355 383 -1355 0 net=3112
rlabel metal2 541 -1355 541 -1355 0 net=2801
rlabel metal2 65 -1357 65 -1357 0 net=1795
rlabel metal2 163 -1357 163 -1357 0 net=1359
rlabel metal2 226 -1357 226 -1357 0 net=1499
rlabel metal2 285 -1357 285 -1357 0 net=115
rlabel metal2 383 -1357 383 -1357 0 net=403
rlabel metal2 474 -1357 474 -1357 0 net=4076
rlabel metal2 72 -1359 72 -1359 0 net=1303
rlabel metal2 240 -1359 240 -1359 0 net=1391
rlabel metal2 289 -1359 289 -1359 0 net=1559
rlabel metal2 387 -1359 387 -1359 0 net=3194
rlabel metal2 478 -1359 478 -1359 0 net=3144
rlabel metal2 583 -1359 583 -1359 0 net=3957
rlabel metal2 44 -1361 44 -1361 0 net=3529
rlabel metal2 285 -1361 285 -1361 0 net=1469
rlabel metal2 436 -1361 436 -1361 0 net=2617
rlabel metal2 481 -1361 481 -1361 0 net=4192
rlabel metal2 75 -1363 75 -1363 0 net=1074
rlabel metal2 100 -1363 100 -1363 0 net=391
rlabel metal2 401 -1363 401 -1363 0 net=2269
rlabel metal2 481 -1363 481 -1363 0 net=4131
rlabel metal2 79 -1365 79 -1365 0 net=3521
rlabel metal2 485 -1365 485 -1365 0 net=3181
rlabel metal2 485 -1365 485 -1365 0 net=3181
rlabel metal2 492 -1365 492 -1365 0 net=3575
rlabel metal2 548 -1365 548 -1365 0 net=3783
rlabel metal2 600 -1365 600 -1365 0 net=4201
rlabel metal2 93 -1367 93 -1367 0 net=1993
rlabel metal2 124 -1367 124 -1367 0 net=1909
rlabel metal2 429 -1367 429 -1367 0 net=3155
rlabel metal2 562 -1367 562 -1367 0 net=4085
rlabel metal2 107 -1369 107 -1369 0 net=1464
rlabel metal2 212 -1369 212 -1369 0 net=1267
rlabel metal2 310 -1369 310 -1369 0 net=3755
rlabel metal2 107 -1371 107 -1371 0 net=2529
rlabel metal2 310 -1371 310 -1371 0 net=1579
rlabel metal2 492 -1371 492 -1371 0 net=3039
rlabel metal2 513 -1371 513 -1371 0 net=3811
rlabel metal2 114 -1373 114 -1373 0 net=1905
rlabel metal2 170 -1373 170 -1373 0 net=2107
rlabel metal2 362 -1373 362 -1373 0 net=3491
rlabel metal2 23 -1375 23 -1375 0 net=2368
rlabel metal2 471 -1375 471 -1375 0 net=3725
rlabel metal2 121 -1377 121 -1377 0 net=1172
rlabel metal2 331 -1377 331 -1377 0 net=2929
rlabel metal2 499 -1377 499 -1377 0 net=2425
rlabel metal2 128 -1379 128 -1379 0 net=1693
rlabel metal2 296 -1379 296 -1379 0 net=2451
rlabel metal2 369 -1379 369 -1379 0 net=4317
rlabel metal2 506 -1379 506 -1379 0 net=3235
rlabel metal2 296 -1381 296 -1381 0 net=2989
rlabel metal2 464 -1381 464 -1381 0 net=3305
rlabel metal2 317 -1383 317 -1383 0 net=1691
rlabel metal2 33 -1394 33 -1394 0 net=379
rlabel metal2 233 -1394 233 -1394 0 net=2990
rlabel metal2 317 -1394 317 -1394 0 net=1692
rlabel metal2 366 -1394 366 -1394 0 net=3328
rlabel metal2 453 -1394 453 -1394 0 net=3784
rlabel metal2 600 -1394 600 -1394 0 net=3004
rlabel metal2 705 -1394 705 -1394 0 net=740
rlabel metal2 705 -1394 705 -1394 0 net=740
rlabel metal2 37 -1396 37 -1396 0 net=4122
rlabel metal2 233 -1396 233 -1396 0 net=3306
rlabel metal2 551 -1396 551 -1396 0 net=4214
rlabel metal2 604 -1396 604 -1396 0 net=4133
rlabel metal2 604 -1396 604 -1396 0 net=4133
rlabel metal2 621 -1396 621 -1396 0 net=2426
rlabel metal2 646 -1396 646 -1396 0 net=4218
rlabel metal2 646 -1396 646 -1396 0 net=4218
rlabel metal2 37 -1398 37 -1398 0 net=1581
rlabel metal2 317 -1398 317 -1398 0 net=1585
rlabel metal2 373 -1398 373 -1398 0 net=3080
rlabel metal2 390 -1398 390 -1398 0 net=2270
rlabel metal2 460 -1398 460 -1398 0 net=2265
rlabel metal2 635 -1398 635 -1398 0 net=2846
rlabel metal2 44 -1400 44 -1400 0 net=3530
rlabel metal2 380 -1400 380 -1400 0 net=3182
rlabel metal2 499 -1400 499 -1400 0 net=4319
rlabel metal2 44 -1402 44 -1402 0 net=3901
rlabel metal2 184 -1402 184 -1402 0 net=1560
rlabel metal2 369 -1402 369 -1402 0 net=3756
rlabel metal2 51 -1404 51 -1404 0 net=3148
rlabel metal2 275 -1404 275 -1404 0 net=1392
rlabel metal2 296 -1404 296 -1404 0 net=1911
rlabel metal2 331 -1404 331 -1404 0 net=2453
rlabel metal2 387 -1404 387 -1404 0 net=509
rlabel metal2 432 -1404 432 -1404 0 net=3726
rlabel metal2 51 -1406 51 -1406 0 net=1907
rlabel metal2 124 -1406 124 -1406 0 net=420
rlabel metal2 201 -1406 201 -1406 0 net=627
rlabel metal2 404 -1406 404 -1406 0 net=3065
rlabel metal2 436 -1406 436 -1406 0 net=2619
rlabel metal2 464 -1406 464 -1406 0 net=3236
rlabel metal2 513 -1406 513 -1406 0 net=3813
rlabel metal2 58 -1408 58 -1408 0 net=1928
rlabel metal2 247 -1408 247 -1408 0 net=3156
rlabel metal2 58 -1410 58 -1410 0 net=1361
rlabel metal2 247 -1410 247 -1410 0 net=1791
rlabel metal2 464 -1410 464 -1410 0 net=4086
rlabel metal2 72 -1412 72 -1412 0 net=1304
rlabel metal2 261 -1412 261 -1412 0 net=1714
rlabel metal2 394 -1412 394 -1412 0 net=2769
rlabel metal2 418 -1412 418 -1412 0 net=3576
rlabel metal2 583 -1412 583 -1412 0 net=4203
rlabel metal2 72 -1414 72 -1414 0 net=1707
rlabel metal2 163 -1414 163 -1414 0 net=1025
rlabel metal2 187 -1414 187 -1414 0 net=128
rlabel metal2 401 -1414 401 -1414 0 net=2857
rlabel metal2 485 -1414 485 -1414 0 net=2803
rlabel metal2 86 -1416 86 -1416 0 net=2812
rlabel metal2 107 -1416 107 -1416 0 net=2531
rlabel metal2 397 -1416 397 -1416 0 net=4281
rlabel metal2 79 -1418 79 -1418 0 net=3523
rlabel metal2 93 -1418 93 -1418 0 net=1995
rlabel metal2 93 -1418 93 -1418 0 net=1995
rlabel metal2 103 -1418 103 -1418 0 net=1470
rlabel metal2 310 -1418 310 -1418 0 net=3727
rlabel metal2 422 -1418 422 -1418 0 net=2535
rlabel metal2 79 -1420 79 -1420 0 net=1501
rlabel metal2 243 -1420 243 -1420 0 net=3611
rlabel metal2 107 -1422 107 -1422 0 net=3203
rlabel metal2 138 -1422 138 -1422 0 net=1591
rlabel metal2 177 -1422 177 -1422 0 net=1949
rlabel metal2 425 -1422 425 -1422 0 net=3237
rlabel metal2 205 -1424 205 -1424 0 net=1397
rlabel metal2 254 -1424 254 -1424 0 net=1455
rlabel metal2 268 -1424 268 -1424 0 net=1748
rlabel metal2 436 -1424 436 -1424 0 net=4052
rlabel metal2 219 -1426 219 -1426 0 net=1851
rlabel metal2 275 -1426 275 -1426 0 net=2055
rlabel metal2 492 -1426 492 -1426 0 net=3041
rlabel metal2 513 -1426 513 -1426 0 net=3493
rlabel metal2 576 -1426 576 -1426 0 net=3959
rlabel metal2 191 -1428 191 -1428 0 net=3965
rlabel metal2 191 -1430 191 -1430 0 net=1269
rlabel metal2 240 -1430 240 -1430 0 net=1849
rlabel metal2 282 -1430 282 -1430 0 net=2939
rlabel metal2 65 -1432 65 -1432 0 net=1796
rlabel metal2 215 -1432 215 -1432 0 net=2671
rlabel metal2 289 -1432 289 -1432 0 net=2509
rlabel metal2 331 -1432 331 -1432 0 net=2343
rlabel metal2 471 -1432 471 -1432 0 net=2931
rlabel metal2 65 -1434 65 -1434 0 net=2109
rlabel metal2 338 -1434 338 -1434 0 net=1207
rlabel metal2 128 -1436 128 -1436 0 net=1695
rlabel metal2 439 -1436 439 -1436 0 net=2675
rlabel metal2 117 -1438 117 -1438 0 net=1235
rlabel metal2 145 -1438 145 -1438 0 net=1403
rlabel metal2 145 -1440 145 -1440 0 net=3454
rlabel metal2 408 -1442 408 -1442 0 net=2483
rlabel metal2 16 -1453 16 -1453 0 net=1951
rlabel metal2 215 -1453 215 -1453 0 net=37
rlabel metal2 429 -1453 429 -1453 0 net=3066
rlabel metal2 702 -1453 702 -1453 0 net=188
rlabel metal2 44 -1455 44 -1455 0 net=3902
rlabel metal2 163 -1455 163 -1455 0 net=1026
rlabel metal2 254 -1455 254 -1455 0 net=1850
rlabel metal2 310 -1455 310 -1455 0 net=3728
rlabel metal2 443 -1455 443 -1455 0 net=3814
rlabel metal2 548 -1455 548 -1455 0 net=4321
rlabel metal2 51 -1457 51 -1457 0 net=1908
rlabel metal2 254 -1457 254 -1457 0 net=1167
rlabel metal2 327 -1457 327 -1457 0 net=2344
rlabel metal2 359 -1457 359 -1457 0 net=2770
rlabel metal2 422 -1457 422 -1457 0 net=2537
rlabel metal2 450 -1457 450 -1457 0 net=2933
rlabel metal2 562 -1457 562 -1457 0 net=4134
rlabel metal2 65 -1459 65 -1459 0 net=2110
rlabel metal2 268 -1459 268 -1459 0 net=2917
rlabel metal2 432 -1459 432 -1459 0 net=2804
rlabel metal2 492 -1459 492 -1459 0 net=3613
rlabel metal2 565 -1459 565 -1459 0 net=2266
rlabel metal2 51 -1461 51 -1461 0 net=1493
rlabel metal2 72 -1461 72 -1461 0 net=1708
rlabel metal2 271 -1461 271 -1461 0 net=2484
rlabel metal2 436 -1461 436 -1461 0 net=3043
rlabel metal2 534 -1461 534 -1461 0 net=3921
rlabel metal2 569 -1461 569 -1461 0 net=4205
rlabel metal2 72 -1463 72 -1463 0 net=1271
rlabel metal2 212 -1463 212 -1463 0 net=1055
rlabel metal2 240 -1463 240 -1463 0 net=4361
rlabel metal2 478 -1463 478 -1463 0 net=3238
rlabel metal2 572 -1463 572 -1463 0 net=4027
rlabel metal2 58 -1465 58 -1465 0 net=1362
rlabel metal2 271 -1465 271 -1465 0 net=1696
rlabel metal2 331 -1465 331 -1465 0 net=2621
rlabel metal2 478 -1465 478 -1465 0 net=4282
rlabel metal2 58 -1467 58 -1467 0 net=1793
rlabel metal2 282 -1467 282 -1467 0 net=2672
rlabel metal2 401 -1467 401 -1467 0 net=2859
rlabel metal2 506 -1467 506 -1467 0 net=3663
rlabel metal2 79 -1469 79 -1469 0 net=1502
rlabel metal2 250 -1469 250 -1469 0 net=3017
rlabel metal2 457 -1469 457 -1469 0 net=2941
rlabel metal2 520 -1469 520 -1469 0 net=3961
rlabel metal2 79 -1471 79 -1471 0 net=1853
rlabel metal2 261 -1471 261 -1471 0 net=1457
rlabel metal2 289 -1471 289 -1471 0 net=2511
rlabel metal2 429 -1471 429 -1471 0 net=3581
rlabel metal2 541 -1471 541 -1471 0 net=3967
rlabel metal2 576 -1471 576 -1471 0 net=4171
rlabel metal2 37 -1473 37 -1473 0 net=1582
rlabel metal2 292 -1473 292 -1473 0 net=2501
rlabel metal2 37 -1475 37 -1475 0 net=2255
rlabel metal2 86 -1475 86 -1475 0 net=3524
rlabel metal2 163 -1475 163 -1475 0 net=771
rlabel metal2 261 -1475 261 -1475 0 net=1209
rlabel metal2 345 -1475 345 -1475 0 net=2533
rlabel metal2 30 -1477 30 -1477 0 net=2527
rlabel metal2 93 -1477 93 -1477 0 net=1996
rlabel metal2 142 -1477 142 -1477 0 net=3931
rlabel metal2 205 -1477 205 -1477 0 net=1399
rlabel metal2 296 -1477 296 -1477 0 net=1913
rlabel metal2 359 -1477 359 -1477 0 net=2455
rlabel metal2 93 -1479 93 -1479 0 net=3205
rlabel metal2 110 -1479 110 -1479 0 net=4301
rlabel metal2 149 -1479 149 -1479 0 net=1593
rlabel metal2 296 -1479 296 -1479 0 net=1377
rlabel metal2 100 -1481 100 -1481 0 net=1437
rlabel metal2 107 -1483 107 -1483 0 net=503
rlabel metal2 170 -1483 170 -1483 0 net=1404
rlabel metal2 338 -1483 338 -1483 0 net=2677
rlabel metal2 114 -1485 114 -1485 0 net=1237
rlabel metal2 135 -1485 135 -1485 0 net=2057
rlabel metal2 369 -1485 369 -1485 0 net=3971
rlabel metal2 128 -1487 128 -1487 0 net=1655
rlabel metal2 177 -1487 177 -1487 0 net=3459
rlabel metal2 380 -1487 380 -1487 0 net=2379
rlabel metal2 471 -1487 471 -1487 0 net=3495
rlabel metal2 124 -1489 124 -1489 0 net=3837
rlabel metal2 156 -1491 156 -1491 0 net=4103
rlabel metal2 275 -1493 275 -1493 0 net=3145
rlabel metal2 390 -1493 390 -1493 0 net=3425
rlabel metal2 317 -1495 317 -1495 0 net=1586
rlabel metal2 16 -1506 16 -1506 0 net=1952
rlabel metal2 173 -1506 173 -1506 0 net=3932
rlabel metal2 205 -1506 205 -1506 0 net=3146
rlabel metal2 292 -1506 292 -1506 0 net=2538
rlabel metal2 464 -1506 464 -1506 0 net=3426
rlabel metal2 478 -1506 478 -1506 0 net=3839
rlabel metal2 565 -1506 565 -1506 0 net=4206
rlabel metal2 579 -1506 579 -1506 0 net=4028
rlabel metal2 590 -1506 590 -1506 0 net=4173
rlabel metal2 590 -1506 590 -1506 0 net=4173
rlabel metal2 23 -1508 23 -1508 0 net=624
rlabel metal2 58 -1508 58 -1508 0 net=1794
rlabel metal2 142 -1508 142 -1508 0 net=4303
rlabel metal2 184 -1508 184 -1508 0 net=2456
rlabel metal2 369 -1508 369 -1508 0 net=3044
rlabel metal2 443 -1508 443 -1508 0 net=2935
rlabel metal2 488 -1508 488 -1508 0 net=3972
rlabel metal2 30 -1510 30 -1510 0 net=2528
rlabel metal2 72 -1510 72 -1510 0 net=1272
rlabel metal2 152 -1510 152 -1510 0 net=680
rlabel metal2 184 -1510 184 -1510 0 net=3061
rlabel metal2 313 -1510 313 -1510 0 net=2534
rlabel metal2 422 -1510 422 -1510 0 net=3962
rlabel metal2 37 -1512 37 -1512 0 net=2256
rlabel metal2 79 -1512 79 -1512 0 net=1855
rlabel metal2 152 -1512 152 -1512 0 net=166
rlabel metal2 240 -1512 240 -1512 0 net=3968
rlabel metal2 51 -1514 51 -1514 0 net=3207
rlabel metal2 100 -1514 100 -1514 0 net=1439
rlabel metal2 163 -1514 163 -1514 0 net=3137
rlabel metal2 247 -1514 247 -1514 0 net=142
rlabel metal2 320 -1514 320 -1514 0 net=3614
rlabel metal2 506 -1514 506 -1514 0 net=3665
rlabel metal2 506 -1514 506 -1514 0 net=3665
rlabel metal2 513 -1514 513 -1514 0 net=4323
rlabel metal2 65 -1516 65 -1516 0 net=1495
rlabel metal2 86 -1516 86 -1516 0 net=1169
rlabel metal2 268 -1516 268 -1516 0 net=1459
rlabel metal2 303 -1516 303 -1516 0 net=1915
rlabel metal2 401 -1516 401 -1516 0 net=3018
rlabel metal2 429 -1516 429 -1516 0 net=4365
rlabel metal2 492 -1516 492 -1516 0 net=4105
rlabel metal2 65 -1518 65 -1518 0 net=3895
rlabel metal2 275 -1518 275 -1518 0 net=2503
rlabel metal2 387 -1518 387 -1518 0 net=2513
rlabel metal2 89 -1520 89 -1520 0 net=77
rlabel metal2 187 -1520 187 -1520 0 net=4019
rlabel metal2 282 -1520 282 -1520 0 net=377
rlabel metal2 327 -1520 327 -1520 0 net=2860
rlabel metal2 520 -1520 520 -1520 0 net=4247
rlabel metal2 110 -1522 110 -1522 0 net=1656
rlabel metal2 135 -1522 135 -1522 0 net=2059
rlabel metal2 261 -1522 261 -1522 0 net=1211
rlabel metal2 331 -1522 331 -1522 0 net=2623
rlabel metal2 373 -1522 373 -1522 0 net=2381
rlabel metal2 383 -1522 383 -1522 0 net=592
rlabel metal2 436 -1522 436 -1522 0 net=2943
rlabel metal2 114 -1524 114 -1524 0 net=1238
rlabel metal2 191 -1524 191 -1524 0 net=1595
rlabel metal2 229 -1524 229 -1524 0 net=1963
rlabel metal2 380 -1524 380 -1524 0 net=3559
rlabel metal2 450 -1524 450 -1524 0 net=3497
rlabel metal2 96 -1526 96 -1526 0 net=1481
rlabel metal2 128 -1526 128 -1526 0 net=1401
rlabel metal2 236 -1526 236 -1526 0 net=1681
rlabel metal2 457 -1526 457 -1526 0 net=3583
rlabel metal2 135 -1528 135 -1528 0 net=1379
rlabel metal2 499 -1528 499 -1528 0 net=3922
rlabel metal2 156 -1530 156 -1530 0 net=3607
rlabel metal2 198 -1532 198 -1532 0 net=1056
rlabel metal2 236 -1532 236 -1532 0 net=2035
rlabel metal2 212 -1534 212 -1534 0 net=1367
rlabel metal2 296 -1534 296 -1534 0 net=1645
rlabel metal2 317 -1536 317 -1536 0 net=4363
rlabel metal2 352 -1538 352 -1538 0 net=3461
rlabel metal2 352 -1540 352 -1540 0 net=2919
rlabel metal2 338 -1542 338 -1542 0 net=2679
rlabel metal2 338 -1544 338 -1544 0 net=1497
rlabel metal2 51 -1555 51 -1555 0 net=3208
rlabel metal2 121 -1555 121 -1555 0 net=1856
rlabel metal2 261 -1555 261 -1555 0 net=1964
rlabel metal2 289 -1555 289 -1555 0 net=2037
rlabel metal2 352 -1555 352 -1555 0 net=2921
rlabel metal2 352 -1555 352 -1555 0 net=2921
rlabel metal2 359 -1555 359 -1555 0 net=2624
rlabel metal2 401 -1555 401 -1555 0 net=3561
rlabel metal2 401 -1555 401 -1555 0 net=3561
rlabel metal2 415 -1555 415 -1555 0 net=2944
rlabel metal2 450 -1555 450 -1555 0 net=3499
rlabel metal2 485 -1555 485 -1555 0 net=4248
rlabel metal2 586 -1555 586 -1555 0 net=4174
rlabel metal2 72 -1557 72 -1557 0 net=1496
rlabel metal2 86 -1557 86 -1557 0 net=1170
rlabel metal2 226 -1557 226 -1557 0 net=2161
rlabel metal2 236 -1557 236 -1557 0 net=2060
rlabel metal2 261 -1557 261 -1557 0 net=1461
rlabel metal2 271 -1557 271 -1557 0 net=3199
rlabel metal2 380 -1557 380 -1557 0 net=4106
rlabel metal2 513 -1557 513 -1557 0 net=4325
rlabel metal2 513 -1557 513 -1557 0 net=4325
rlabel metal2 75 -1559 75 -1559 0 net=3455
rlabel metal2 96 -1559 96 -1559 0 net=383
rlabel metal2 422 -1559 422 -1559 0 net=418
rlabel metal2 103 -1561 103 -1561 0 net=1482
rlabel metal2 128 -1561 128 -1561 0 net=1402
rlabel metal2 331 -1561 331 -1561 0 net=1683
rlabel metal2 331 -1561 331 -1561 0 net=1683
rlabel metal2 429 -1561 429 -1561 0 net=3608
rlabel metal2 149 -1563 149 -1563 0 net=4304
rlabel metal2 194 -1563 194 -1563 0 net=1646
rlabel metal2 303 -1563 303 -1563 0 net=1917
rlabel metal2 303 -1563 303 -1563 0 net=1917
rlabel metal2 310 -1563 310 -1563 0 net=1212
rlabel metal2 429 -1563 429 -1563 0 net=4367
rlabel metal2 492 -1563 492 -1563 0 net=3667
rlabel metal2 142 -1565 142 -1565 0 net=1440
rlabel metal2 198 -1565 198 -1565 0 net=245
rlabel metal2 240 -1565 240 -1565 0 net=1498
rlabel metal2 369 -1565 369 -1565 0 net=2680
rlabel metal2 436 -1565 436 -1565 0 net=2937
rlabel metal2 457 -1565 457 -1565 0 net=3585
rlabel metal2 142 -1567 142 -1567 0 net=176
rlabel metal2 205 -1567 205 -1567 0 net=1596
rlabel metal2 247 -1567 247 -1567 0 net=3081
rlabel metal2 317 -1567 317 -1567 0 net=4364
rlabel metal2 128 -1569 128 -1569 0 net=1325
rlabel metal2 219 -1569 219 -1569 0 net=4020
rlabel metal2 275 -1569 275 -1569 0 net=2505
rlabel metal2 317 -1569 317 -1569 0 net=3840
rlabel metal2 159 -1571 159 -1571 0 net=1368
rlabel metal2 254 -1571 254 -1571 0 net=2773
rlabel metal2 292 -1571 292 -1571 0 net=2514
rlabel metal2 65 -1573 65 -1573 0 net=3896
rlabel metal2 163 -1573 163 -1573 0 net=3139
rlabel metal2 173 -1573 173 -1573 0 net=101
rlabel metal2 275 -1573 275 -1573 0 net=1737
rlabel metal2 373 -1573 373 -1573 0 net=2383
rlabel metal2 135 -1575 135 -1575 0 net=1381
rlabel metal2 324 -1575 324 -1575 0 net=3697
rlabel metal2 135 -1577 135 -1577 0 net=3441
rlabel metal2 163 -1577 163 -1577 0 net=3063
rlabel metal2 373 -1577 373 -1577 0 net=3463
rlabel metal2 152 -1579 152 -1579 0 net=473
rlabel metal2 156 -1581 156 -1581 0 net=359
rlabel metal2 72 -1592 72 -1592 0 net=2663
rlabel metal2 89 -1592 89 -1592 0 net=1577
rlabel metal2 128 -1592 128 -1592 0 net=1326
rlabel metal2 163 -1592 163 -1592 0 net=3064
rlabel metal2 219 -1592 219 -1592 0 net=1057
rlabel metal2 243 -1592 243 -1592 0 net=1462
rlabel metal2 282 -1592 282 -1592 0 net=2038
rlabel metal2 296 -1592 296 -1592 0 net=2506
rlabel metal2 320 -1592 320 -1592 0 net=127
rlabel metal2 345 -1592 345 -1592 0 net=2922
rlabel metal2 366 -1592 366 -1592 0 net=3465
rlabel metal2 383 -1592 383 -1592 0 net=4368
rlabel metal2 471 -1592 471 -1592 0 net=3500
rlabel metal2 492 -1592 492 -1592 0 net=3669
rlabel metal2 492 -1592 492 -1592 0 net=3669
rlabel metal2 506 -1592 506 -1592 0 net=4326
rlabel metal2 75 -1594 75 -1594 0 net=3456
rlabel metal2 135 -1594 135 -1594 0 net=3442
rlabel metal2 163 -1594 163 -1594 0 net=3271
rlabel metal2 205 -1594 205 -1594 0 net=3083
rlabel metal2 254 -1594 254 -1594 0 net=2774
rlabel metal2 387 -1594 387 -1594 0 net=3341
rlabel metal2 387 -1594 387 -1594 0 net=3341
rlabel metal2 394 -1594 394 -1594 0 net=2385
rlabel metal2 394 -1594 394 -1594 0 net=2385
rlabel metal2 422 -1594 422 -1594 0 net=2938
rlabel metal2 443 -1594 443 -1594 0 net=4097
rlabel metal2 114 -1596 114 -1596 0 net=1895
rlabel metal2 170 -1596 170 -1596 0 net=3140
rlabel metal2 170 -1596 170 -1596 0 net=3140
rlabel metal2 177 -1596 177 -1596 0 net=978
rlabel metal2 275 -1596 275 -1596 0 net=1739
rlabel metal2 317 -1596 317 -1596 0 net=3185
rlabel metal2 352 -1596 352 -1596 0 net=1727
rlabel metal2 464 -1596 464 -1596 0 net=3587
rlabel metal2 131 -1598 131 -1598 0 net=2851
rlabel metal2 142 -1598 142 -1598 0 net=2649
rlabel metal2 156 -1598 156 -1598 0 net=3619
rlabel metal2 282 -1598 282 -1598 0 net=2821
rlabel metal2 317 -1598 317 -1598 0 net=3201
rlabel metal2 184 -1600 184 -1600 0 net=157
rlabel metal2 226 -1600 226 -1600 0 net=3698
rlabel metal2 331 -1600 331 -1600 0 net=1684
rlabel metal2 338 -1600 338 -1600 0 net=3562
rlabel metal2 191 -1602 191 -1602 0 net=440
rlabel metal2 212 -1602 212 -1602 0 net=1382
rlabel metal2 299 -1602 299 -1602 0 net=3475
rlabel metal2 191 -1604 191 -1604 0 net=66
rlabel metal2 226 -1604 226 -1604 0 net=1465
rlabel metal2 233 -1606 233 -1606 0 net=2163
rlabel metal2 261 -1606 261 -1606 0 net=1918
rlabel metal2 236 -1608 236 -1608 0 net=630
rlabel metal2 240 -1610 240 -1610 0 net=844
rlabel metal2 243 -1612 243 -1612 0 net=4029
rlabel metal2 250 -1614 250 -1614 0 net=2415
rlabel metal2 30 -1625 30 -1625 0 net=723
rlabel metal2 37 -1625 37 -1625 0 net=3723
rlabel metal2 198 -1625 198 -1625 0 net=294
rlabel metal2 233 -1625 233 -1625 0 net=57
rlabel metal2 240 -1625 240 -1625 0 net=72
rlabel metal2 275 -1625 275 -1625 0 net=3202
rlabel metal2 334 -1625 334 -1625 0 net=3466
rlabel metal2 387 -1625 387 -1625 0 net=3343
rlabel metal2 387 -1625 387 -1625 0 net=3343
rlabel metal2 394 -1625 394 -1625 0 net=2386
rlabel metal2 394 -1625 394 -1625 0 net=2386
rlabel metal2 401 -1625 401 -1625 0 net=4098
rlabel metal2 467 -1625 467 -1625 0 net=3588
rlabel metal2 488 -1625 488 -1625 0 net=3670
rlabel metal2 44 -1627 44 -1627 0 net=3621
rlabel metal2 177 -1627 177 -1627 0 net=1058
rlabel metal2 254 -1627 254 -1627 0 net=2165
rlabel metal2 261 -1627 261 -1627 0 net=1729
rlabel metal2 359 -1627 359 -1627 0 net=3477
rlabel metal2 51 -1629 51 -1629 0 net=3579
rlabel metal2 93 -1629 93 -1629 0 net=1578
rlabel metal2 121 -1629 121 -1629 0 net=2650
rlabel metal2 149 -1629 149 -1629 0 net=3272
rlabel metal2 177 -1629 177 -1629 0 net=2001
rlabel metal2 205 -1629 205 -1629 0 net=3084
rlabel metal2 205 -1629 205 -1629 0 net=3084
rlabel metal2 212 -1629 212 -1629 0 net=1749
rlabel metal2 254 -1629 254 -1629 0 net=1741
rlabel metal2 296 -1629 296 -1629 0 net=4030
rlabel metal2 327 -1629 327 -1629 0 net=2215
rlabel metal2 65 -1631 65 -1631 0 net=2775
rlabel metal2 124 -1631 124 -1631 0 net=2852
rlabel metal2 138 -1631 138 -1631 0 net=475
rlabel metal2 191 -1631 191 -1631 0 net=1067
rlabel metal2 303 -1631 303 -1631 0 net=2417
rlabel metal2 72 -1633 72 -1633 0 net=2664
rlabel metal2 100 -1633 100 -1633 0 net=1863
rlabel metal2 135 -1633 135 -1633 0 net=1141
rlabel metal2 163 -1633 163 -1633 0 net=1467
rlabel metal2 264 -1633 264 -1633 0 net=1797
rlabel metal2 345 -1633 345 -1633 0 net=3187
rlabel metal2 72 -1635 72 -1635 0 net=2609
rlabel metal2 170 -1635 170 -1635 0 net=1605
rlabel metal2 275 -1635 275 -1635 0 net=1961
rlabel metal2 345 -1635 345 -1635 0 net=2951
rlabel metal2 79 -1637 79 -1637 0 net=1897
rlabel metal2 198 -1637 198 -1637 0 net=822
rlabel metal2 226 -1637 226 -1637 0 net=1987
rlabel metal2 303 -1637 303 -1637 0 net=2822
rlabel metal2 58 -1639 58 -1639 0 net=767
rlabel metal2 219 -1639 219 -1639 0 net=3939
rlabel metal2 86 -1641 86 -1641 0 net=1759
rlabel metal2 278 -1641 278 -1641 0 net=3321
rlabel metal2 107 -1643 107 -1643 0 net=1205
rlabel metal2 282 -1643 282 -1643 0 net=1225
rlabel metal2 19 -1654 19 -1654 0 net=3373
rlabel metal2 37 -1654 37 -1654 0 net=3724
rlabel metal2 226 -1654 226 -1654 0 net=3188
rlabel metal2 387 -1654 387 -1654 0 net=3344
rlabel metal2 44 -1656 44 -1656 0 net=3622
rlabel metal2 149 -1656 149 -1656 0 net=1206
rlabel metal2 219 -1656 219 -1656 0 net=580
rlabel metal2 243 -1656 243 -1656 0 net=1730
rlabel metal2 268 -1656 268 -1656 0 net=1226
rlabel metal2 317 -1656 317 -1656 0 net=1799
rlabel metal2 51 -1658 51 -1658 0 net=3580
rlabel metal2 163 -1658 163 -1658 0 net=1468
rlabel metal2 191 -1658 191 -1658 0 net=1069
rlabel metal2 212 -1658 212 -1658 0 net=2166
rlabel metal2 296 -1658 296 -1658 0 net=1989
rlabel metal2 324 -1658 324 -1658 0 net=3322
rlabel metal2 65 -1660 65 -1660 0 net=2776
rlabel metal2 100 -1660 100 -1660 0 net=1865
rlabel metal2 156 -1660 156 -1660 0 net=1143
rlabel metal2 212 -1660 212 -1660 0 net=2421
rlabel metal2 331 -1660 331 -1660 0 net=3941
rlabel metal2 72 -1662 72 -1662 0 net=2610
rlabel metal2 103 -1662 103 -1662 0 net=3395
rlabel metal2 117 -1662 117 -1662 0 net=239
rlabel metal2 226 -1662 226 -1662 0 net=2557
rlabel metal2 331 -1662 331 -1662 0 net=2953
rlabel metal2 366 -1662 366 -1662 0 net=3478
rlabel metal2 79 -1664 79 -1664 0 net=1898
rlabel metal2 156 -1664 156 -1664 0 net=1607
rlabel metal2 222 -1664 222 -1664 0 net=3973
rlabel metal2 86 -1666 86 -1666 0 net=1760
rlabel metal2 121 -1666 121 -1666 0 net=764
rlabel metal2 229 -1666 229 -1666 0 net=563
rlabel metal2 338 -1666 338 -1666 0 net=1962
rlabel metal2 121 -1668 121 -1668 0 net=2003
rlabel metal2 205 -1668 205 -1668 0 net=2805
rlabel metal2 145 -1670 145 -1670 0 net=1929
rlabel metal2 205 -1670 205 -1670 0 net=998
rlabel metal2 282 -1670 282 -1670 0 net=2216
rlabel metal2 233 -1672 233 -1672 0 net=1751
rlabel metal2 254 -1672 254 -1672 0 net=1743
rlabel metal2 285 -1672 285 -1672 0 net=3397
rlabel metal2 348 -1672 348 -1672 0 net=3537
rlabel metal2 208 -1674 208 -1674 0 net=1783
rlabel metal2 261 -1674 261 -1674 0 net=2723
rlabel metal2 236 -1676 236 -1676 0 net=2418
rlabel metal2 240 -1678 240 -1678 0 net=946
rlabel metal2 2 -1689 2 -1689 0 net=3371
rlabel metal2 16 -1689 16 -1689 0 net=3374
rlabel metal2 30 -1689 30 -1689 0 net=22
rlabel metal2 79 -1689 79 -1689 0 net=465
rlabel metal2 79 -1689 79 -1689 0 net=465
rlabel metal2 89 -1689 89 -1689 0 net=167
rlabel metal2 100 -1689 100 -1689 0 net=3396
rlabel metal2 114 -1689 114 -1689 0 net=299
rlabel metal2 222 -1689 222 -1689 0 net=991
rlabel metal2 254 -1689 254 -1689 0 net=1800
rlabel metal2 121 -1691 121 -1691 0 net=2004
rlabel metal2 226 -1691 226 -1691 0 net=1752
rlabel metal2 257 -1691 257 -1691 0 net=2422
rlabel metal2 317 -1691 317 -1691 0 net=2954
rlabel metal2 352 -1691 352 -1691 0 net=3538
rlabel metal2 352 -1691 352 -1691 0 net=3538
rlabel metal2 359 -1691 359 -1691 0 net=3942
rlabel metal2 121 -1693 121 -1693 0 net=682
rlabel metal2 156 -1693 156 -1693 0 net=1608
rlabel metal2 191 -1693 191 -1693 0 net=1784
rlabel metal2 264 -1693 264 -1693 0 net=1990
rlabel metal2 135 -1695 135 -1695 0 net=1867
rlabel metal2 163 -1695 163 -1695 0 net=1144
rlabel metal2 194 -1695 194 -1695 0 net=4279
rlabel metal2 226 -1695 226 -1695 0 net=2558
rlabel metal2 131 -1697 131 -1697 0 net=4025
rlabel metal2 149 -1697 149 -1697 0 net=1931
rlabel metal2 170 -1697 170 -1697 0 net=2187
rlabel metal2 198 -1697 198 -1697 0 net=1070
rlabel metal2 229 -1697 229 -1697 0 net=1059
rlabel metal2 268 -1697 268 -1697 0 net=1744
rlabel metal2 292 -1697 292 -1697 0 net=3974
rlabel metal2 117 -1699 117 -1699 0 net=412
rlabel metal2 173 -1699 173 -1699 0 net=2625
rlabel metal2 201 -1699 201 -1699 0 net=3165
rlabel metal2 275 -1699 275 -1699 0 net=279
rlabel metal2 285 -1699 285 -1699 0 net=507
rlabel metal2 296 -1699 296 -1699 0 net=2806
rlabel metal2 303 -1701 303 -1701 0 net=2725
rlabel metal2 324 -1701 324 -1701 0 net=3399
rlabel metal2 5 -1712 5 -1712 0 net=3372
rlabel metal2 128 -1712 128 -1712 0 net=4026
rlabel metal2 142 -1712 142 -1712 0 net=1932
rlabel metal2 170 -1712 170 -1712 0 net=2188
rlabel metal2 212 -1712 212 -1712 0 net=3166
rlabel metal2 233 -1712 233 -1712 0 net=1060
rlabel metal2 303 -1712 303 -1712 0 net=2726
rlabel metal2 317 -1712 317 -1712 0 net=3400
rlabel metal2 152 -1714 152 -1714 0 net=1868
rlabel metal2 177 -1714 177 -1714 0 net=2626
rlabel metal2 187 -1716 187 -1716 0 net=4280
<< end >>
