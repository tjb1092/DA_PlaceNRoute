magic
tech scmos
timestamp 1555016892 
<< pdiffusion >>
rect 1 -6 7 0
rect 8 -6 14 0
rect 43 -6 49 0
rect 50 -6 56 0
rect 85 -6 91 0
rect 1 -17 7 -11
rect 22 -17 28 -11
rect 29 -17 32 -11
rect 36 -17 42 -11
rect 57 -17 60 -11
rect 64 -17 70 -11
rect 85 -17 91 -11
rect 92 -17 95 -11
rect 8 -32 14 -26
rect 15 -32 18 -26
rect 22 -32 28 -26
rect 29 -32 35 -26
rect 36 -32 39 -26
rect 43 -32 46 -26
rect 50 -32 56 -26
rect 57 -32 60 -26
rect 64 -32 67 -26
rect 71 -32 77 -26
rect 78 -32 84 -26
rect 85 -32 88 -26
rect 92 -32 95 -26
rect 15 -53 18 -47
rect 22 -53 25 -47
rect 29 -53 35 -47
rect 36 -53 42 -47
rect 43 -53 49 -47
rect 50 -53 53 -47
rect 57 -53 60 -47
rect 64 -53 70 -47
rect 71 -53 77 -47
rect 78 -53 81 -47
rect 85 -53 88 -47
rect 92 -53 95 -47
rect 99 -53 102 -47
rect 8 -74 14 -68
rect 15 -74 18 -68
rect 22 -74 25 -68
rect 29 -74 35 -68
rect 36 -74 42 -68
rect 43 -74 46 -68
rect 50 -74 56 -68
rect 57 -74 63 -68
rect 64 -74 70 -68
rect 71 -74 77 -68
rect 78 -74 81 -68
rect 85 -74 88 -68
rect 92 -74 95 -68
rect 99 -74 102 -68
rect 106 -74 109 -68
rect 113 -74 119 -68
rect 1 -101 4 -95
rect 8 -101 11 -95
rect 15 -101 21 -95
rect 22 -101 28 -95
rect 29 -101 35 -95
rect 36 -101 39 -95
rect 43 -101 49 -95
rect 50 -101 56 -95
rect 57 -101 63 -95
rect 64 -101 70 -95
rect 71 -101 74 -95
rect 78 -101 84 -95
rect 85 -101 88 -95
rect 92 -101 95 -95
rect 99 -101 102 -95
rect 106 -101 109 -95
rect 113 -101 116 -95
rect 120 -101 123 -95
rect 15 -126 18 -120
rect 22 -126 28 -120
rect 29 -126 32 -120
rect 36 -126 39 -120
rect 43 -126 49 -120
rect 50 -126 56 -120
rect 57 -126 63 -120
rect 64 -126 70 -120
rect 71 -126 74 -120
rect 78 -126 81 -120
rect 85 -126 91 -120
rect 92 -126 95 -120
rect 99 -126 105 -120
rect 1 -147 4 -141
rect 8 -147 11 -141
rect 15 -147 21 -141
rect 22 -147 28 -141
rect 29 -147 35 -141
rect 36 -147 39 -141
rect 43 -147 49 -141
rect 50 -147 56 -141
rect 57 -147 60 -141
rect 64 -147 67 -141
rect 71 -147 74 -141
rect 78 -147 84 -141
rect 85 -147 88 -141
<< polysilicon >>
rect 44 -7 45 -5
rect 47 -7 48 -5
rect 54 -7 55 -5
rect 86 -7 87 -5
rect 26 -18 27 -16
rect 30 -12 31 -10
rect 30 -18 31 -16
rect 37 -12 38 -10
rect 40 -12 41 -10
rect 40 -18 41 -16
rect 58 -12 59 -10
rect 58 -18 59 -16
rect 68 -12 69 -10
rect 86 -18 87 -16
rect 89 -18 90 -16
rect 93 -12 94 -10
rect 93 -18 94 -16
rect 9 -27 10 -25
rect 16 -27 17 -25
rect 16 -33 17 -31
rect 26 -27 27 -25
rect 23 -33 24 -31
rect 26 -33 27 -31
rect 30 -27 31 -25
rect 30 -33 31 -31
rect 33 -33 34 -31
rect 37 -27 38 -25
rect 37 -33 38 -31
rect 44 -27 45 -25
rect 44 -33 45 -31
rect 51 -33 52 -31
rect 54 -33 55 -31
rect 58 -27 59 -25
rect 58 -33 59 -31
rect 65 -27 66 -25
rect 65 -33 66 -31
rect 72 -33 73 -31
rect 75 -33 76 -31
rect 82 -27 83 -25
rect 79 -33 80 -31
rect 86 -27 87 -25
rect 86 -33 87 -31
rect 93 -27 94 -25
rect 93 -33 94 -31
rect 16 -48 17 -46
rect 16 -54 17 -52
rect 23 -48 24 -46
rect 23 -54 24 -52
rect 30 -48 31 -46
rect 33 -48 34 -46
rect 30 -54 31 -52
rect 37 -54 38 -52
rect 40 -54 41 -52
rect 44 -48 45 -46
rect 44 -54 45 -52
rect 51 -48 52 -46
rect 51 -54 52 -52
rect 58 -48 59 -46
rect 58 -54 59 -52
rect 68 -48 69 -46
rect 65 -54 66 -52
rect 68 -54 69 -52
rect 72 -48 73 -46
rect 75 -48 76 -46
rect 79 -48 80 -46
rect 79 -54 80 -52
rect 86 -48 87 -46
rect 86 -54 87 -52
rect 93 -48 94 -46
rect 93 -54 94 -52
rect 100 -48 101 -46
rect 100 -54 101 -52
rect 12 -69 13 -67
rect 16 -69 17 -67
rect 16 -75 17 -73
rect 23 -69 24 -67
rect 23 -75 24 -73
rect 30 -69 31 -67
rect 33 -69 34 -67
rect 30 -75 31 -73
rect 33 -75 34 -73
rect 37 -69 38 -67
rect 40 -69 41 -67
rect 44 -69 45 -67
rect 44 -75 45 -73
rect 51 -69 52 -67
rect 54 -69 55 -67
rect 51 -75 52 -73
rect 54 -75 55 -73
rect 61 -69 62 -67
rect 58 -75 59 -73
rect 65 -69 66 -67
rect 68 -75 69 -73
rect 75 -69 76 -67
rect 75 -75 76 -73
rect 79 -69 80 -67
rect 79 -75 80 -73
rect 86 -69 87 -67
rect 86 -75 87 -73
rect 93 -69 94 -67
rect 93 -75 94 -73
rect 100 -69 101 -67
rect 100 -75 101 -73
rect 107 -69 108 -67
rect 107 -75 108 -73
rect 114 -69 115 -67
rect 117 -69 118 -67
rect 114 -75 115 -73
rect 2 -96 3 -94
rect 2 -102 3 -100
rect 9 -96 10 -94
rect 9 -102 10 -100
rect 16 -96 17 -94
rect 19 -96 20 -94
rect 23 -96 24 -94
rect 23 -102 24 -100
rect 30 -102 31 -100
rect 33 -102 34 -100
rect 37 -96 38 -94
rect 37 -102 38 -100
rect 44 -102 45 -100
rect 47 -102 48 -100
rect 54 -96 55 -94
rect 51 -102 52 -100
rect 54 -102 55 -100
rect 58 -96 59 -94
rect 61 -96 62 -94
rect 58 -102 59 -100
rect 65 -96 66 -94
rect 68 -96 69 -94
rect 65 -102 66 -100
rect 68 -102 69 -100
rect 72 -96 73 -94
rect 72 -102 73 -100
rect 79 -102 80 -100
rect 86 -96 87 -94
rect 86 -102 87 -100
rect 93 -96 94 -94
rect 93 -102 94 -100
rect 100 -96 101 -94
rect 100 -102 101 -100
rect 107 -96 108 -94
rect 107 -102 108 -100
rect 114 -96 115 -94
rect 114 -102 115 -100
rect 121 -96 122 -94
rect 121 -102 122 -100
rect 16 -121 17 -119
rect 16 -127 17 -125
rect 26 -127 27 -125
rect 30 -121 31 -119
rect 30 -127 31 -125
rect 37 -121 38 -119
rect 37 -127 38 -125
rect 44 -121 45 -119
rect 47 -121 48 -119
rect 51 -121 52 -119
rect 54 -121 55 -119
rect 61 -121 62 -119
rect 58 -127 59 -125
rect 65 -121 66 -119
rect 68 -121 69 -119
rect 65 -127 66 -125
rect 68 -127 69 -125
rect 72 -121 73 -119
rect 72 -127 73 -125
rect 79 -121 80 -119
rect 79 -127 80 -125
rect 86 -121 87 -119
rect 93 -121 94 -119
rect 93 -127 94 -125
rect 103 -121 104 -119
rect 100 -127 101 -125
rect 2 -142 3 -140
rect 2 -148 3 -146
rect 9 -142 10 -140
rect 9 -148 10 -146
rect 19 -142 20 -140
rect 26 -142 27 -140
rect 23 -148 24 -146
rect 30 -142 31 -140
rect 33 -148 34 -146
rect 37 -142 38 -140
rect 37 -148 38 -146
rect 44 -142 45 -140
rect 44 -148 45 -146
rect 51 -148 52 -146
rect 54 -148 55 -146
rect 58 -142 59 -140
rect 58 -148 59 -146
rect 65 -142 66 -140
rect 65 -148 66 -146
rect 72 -142 73 -140
rect 72 -148 73 -146
rect 79 -148 80 -146
rect 82 -148 83 -146
rect 86 -142 87 -140
rect 86 -148 87 -146
<< metal1 >>
rect 30 -9 38 -8
rect 40 -9 45 -8
rect 47 -9 55 -8
rect 58 -9 69 -8
rect 86 -9 94 -8
rect 9 -20 38 -19
rect 40 -20 45 -19
rect 58 -20 66 -19
rect 89 -20 94 -19
rect 16 -22 31 -21
rect 58 -22 83 -21
rect 86 -22 94 -21
rect 30 -24 87 -23
rect 26 -35 31 -34
rect 51 -35 66 -34
rect 72 -35 101 -34
rect 16 -37 31 -36
rect 44 -37 52 -36
rect 54 -37 59 -36
rect 75 -37 87 -36
rect 16 -39 24 -38
rect 33 -39 45 -38
rect 75 -39 87 -38
rect 23 -41 34 -40
rect 37 -41 59 -40
rect 79 -41 94 -40
rect 68 -43 94 -42
rect 72 -45 80 -44
rect 12 -56 55 -55
rect 61 -56 87 -55
rect 16 -58 38 -57
rect 40 -58 52 -57
rect 65 -58 101 -57
rect 16 -60 24 -59
rect 30 -60 34 -59
rect 37 -60 69 -59
rect 75 -60 108 -59
rect 23 -62 31 -61
rect 51 -62 59 -61
rect 65 -62 94 -61
rect 100 -62 118 -61
rect 79 -64 94 -63
rect 40 -66 80 -65
rect 86 -66 115 -65
rect 2 -77 17 -76
rect 19 -77 24 -76
rect 30 -77 38 -76
rect 51 -77 101 -76
rect 107 -77 115 -76
rect 9 -79 34 -78
rect 54 -79 122 -78
rect 16 -81 87 -80
rect 23 -83 55 -82
rect 58 -83 69 -82
rect 75 -83 94 -82
rect 44 -85 94 -84
rect 58 -87 73 -86
rect 79 -87 108 -86
rect 61 -89 101 -88
rect 65 -91 87 -90
rect 68 -93 115 -92
rect 2 -104 24 -103
rect 37 -104 45 -103
rect 47 -104 73 -103
rect 79 -104 101 -103
rect 9 -106 34 -105
rect 37 -106 87 -105
rect 16 -108 59 -107
rect 65 -108 80 -107
rect 86 -108 115 -107
rect 44 -110 55 -109
rect 61 -110 66 -109
rect 68 -110 73 -109
rect 30 -112 55 -111
rect 68 -112 108 -111
rect 30 -114 48 -113
rect 51 -114 122 -113
rect 51 -116 94 -115
rect 93 -118 104 -117
rect 2 -129 20 -128
rect 65 -129 80 -128
rect 86 -129 101 -128
rect 16 -131 27 -130
rect 30 -131 66 -130
rect 68 -131 94 -130
rect 9 -133 31 -132
rect 26 -135 59 -134
rect 37 -137 59 -136
rect 37 -139 45 -138
rect 2 -150 24 -149
rect 33 -150 38 -149
rect 44 -150 66 -149
rect 72 -150 83 -149
rect 9 -152 52 -151
rect 54 -152 59 -151
rect 79 -152 87 -151
<< m2contact >>
rect 30 -9 31 -8
rect 37 -9 38 -8
rect 40 -9 41 -8
rect 44 -9 45 -8
rect 47 -9 48 -8
rect 54 -9 55 -8
rect 58 -9 59 -8
rect 68 -9 69 -8
rect 86 -9 87 -8
rect 93 -9 94 -8
rect 9 -20 10 -19
rect 37 -20 38 -19
rect 40 -20 41 -19
rect 44 -20 45 -19
rect 58 -20 59 -19
rect 65 -20 66 -19
rect 89 -20 90 -19
rect 93 -20 94 -19
rect 16 -22 17 -21
rect 30 -22 31 -21
rect 58 -22 59 -21
rect 82 -22 83 -21
rect 86 -22 87 -21
rect 93 -22 94 -21
rect 30 -24 31 -23
rect 86 -24 87 -23
rect 26 -35 27 -34
rect 30 -35 31 -34
rect 51 -35 52 -34
rect 65 -35 66 -34
rect 72 -35 73 -34
rect 100 -35 101 -34
rect 16 -37 17 -36
rect 30 -37 31 -36
rect 44 -37 45 -36
rect 51 -37 52 -36
rect 54 -37 55 -36
rect 58 -37 59 -36
rect 75 -37 76 -36
rect 86 -37 87 -36
rect 16 -39 17 -38
rect 23 -39 24 -38
rect 33 -39 34 -38
rect 44 -39 45 -38
rect 75 -39 76 -38
rect 86 -39 87 -38
rect 23 -41 24 -40
rect 33 -41 34 -40
rect 37 -41 38 -40
rect 58 -41 59 -40
rect 79 -41 80 -40
rect 93 -41 94 -40
rect 68 -43 69 -42
rect 93 -43 94 -42
rect 72 -45 73 -44
rect 79 -45 80 -44
rect 12 -56 13 -55
rect 54 -56 55 -55
rect 61 -56 62 -55
rect 86 -56 87 -55
rect 16 -58 17 -57
rect 37 -58 38 -57
rect 40 -58 41 -57
rect 51 -58 52 -57
rect 65 -58 66 -57
rect 100 -58 101 -57
rect 16 -60 17 -59
rect 23 -60 24 -59
rect 30 -60 31 -59
rect 33 -60 34 -59
rect 37 -60 38 -59
rect 68 -60 69 -59
rect 75 -60 76 -59
rect 107 -60 108 -59
rect 23 -62 24 -61
rect 30 -62 31 -61
rect 51 -62 52 -61
rect 58 -62 59 -61
rect 65 -62 66 -61
rect 93 -62 94 -61
rect 100 -62 101 -61
rect 117 -62 118 -61
rect 79 -64 80 -63
rect 93 -64 94 -63
rect 40 -66 41 -65
rect 79 -66 80 -65
rect 86 -66 87 -65
rect 114 -66 115 -65
rect 2 -77 3 -76
rect 16 -77 17 -76
rect 19 -77 20 -76
rect 23 -77 24 -76
rect 30 -77 31 -76
rect 37 -77 38 -76
rect 51 -77 52 -76
rect 100 -77 101 -76
rect 107 -77 108 -76
rect 114 -77 115 -76
rect 9 -79 10 -78
rect 33 -79 34 -78
rect 54 -79 55 -78
rect 121 -79 122 -78
rect 16 -81 17 -80
rect 86 -81 87 -80
rect 23 -83 24 -82
rect 54 -83 55 -82
rect 58 -83 59 -82
rect 68 -83 69 -82
rect 75 -83 76 -82
rect 93 -83 94 -82
rect 44 -85 45 -84
rect 93 -85 94 -84
rect 58 -87 59 -86
rect 72 -87 73 -86
rect 79 -87 80 -86
rect 107 -87 108 -86
rect 61 -89 62 -88
rect 100 -89 101 -88
rect 65 -91 66 -90
rect 86 -91 87 -90
rect 68 -93 69 -92
rect 114 -93 115 -92
rect 2 -104 3 -103
rect 23 -104 24 -103
rect 37 -104 38 -103
rect 44 -104 45 -103
rect 47 -104 48 -103
rect 72 -104 73 -103
rect 79 -104 80 -103
rect 100 -104 101 -103
rect 9 -106 10 -105
rect 33 -106 34 -105
rect 37 -106 38 -105
rect 86 -106 87 -105
rect 16 -108 17 -107
rect 58 -108 59 -107
rect 65 -108 66 -107
rect 79 -108 80 -107
rect 86 -108 87 -107
rect 114 -108 115 -107
rect 44 -110 45 -109
rect 54 -110 55 -109
rect 61 -110 62 -109
rect 65 -110 66 -109
rect 68 -110 69 -109
rect 72 -110 73 -109
rect 30 -112 31 -111
rect 54 -112 55 -111
rect 68 -112 69 -111
rect 107 -112 108 -111
rect 30 -114 31 -113
rect 47 -114 48 -113
rect 51 -114 52 -113
rect 121 -114 122 -113
rect 51 -116 52 -115
rect 93 -116 94 -115
rect 93 -118 94 -117
rect 103 -118 104 -117
rect 2 -129 3 -128
rect 19 -129 20 -128
rect 65 -129 66 -128
rect 79 -129 80 -128
rect 86 -129 87 -128
rect 100 -129 101 -128
rect 16 -131 17 -130
rect 26 -131 27 -130
rect 30 -131 31 -130
rect 65 -131 66 -130
rect 68 -131 69 -130
rect 93 -131 94 -130
rect 9 -133 10 -132
rect 30 -133 31 -132
rect 26 -135 27 -134
rect 58 -135 59 -134
rect 37 -137 38 -136
rect 58 -137 59 -136
rect 37 -139 38 -138
rect 44 -139 45 -138
rect 2 -150 3 -149
rect 23 -150 24 -149
rect 33 -150 34 -149
rect 37 -150 38 -149
rect 44 -150 45 -149
rect 65 -150 66 -149
rect 72 -150 73 -149
rect 82 -150 83 -149
rect 9 -152 10 -151
rect 51 -152 52 -151
rect 54 -152 55 -151
rect 58 -152 59 -151
rect 79 -152 80 -151
rect 86 -152 87 -151
<< metal2 >>
rect 30 -10 31 -8
rect 37 -10 38 -8
rect 40 -10 41 -8
rect 44 -9 45 -7
rect 47 -9 48 -7
rect 54 -9 55 -7
rect 58 -10 59 -8
rect 68 -10 69 -8
rect 86 -9 87 -7
rect 93 -10 94 -8
rect 9 -25 10 -19
rect 37 -25 38 -19
rect 40 -20 41 -18
rect 44 -25 45 -19
rect 58 -20 59 -18
rect 65 -25 66 -19
rect 89 -20 90 -18
rect 93 -20 94 -18
rect 16 -25 17 -21
rect 30 -22 31 -18
rect 58 -25 59 -21
rect 82 -25 83 -21
rect 86 -22 87 -18
rect 93 -25 94 -21
rect 26 -24 27 -18
rect 26 -25 27 -23
rect 26 -24 27 -18
rect 26 -25 27 -23
rect 30 -25 31 -23
rect 86 -25 87 -23
rect 26 -35 27 -33
rect 30 -35 31 -33
rect 51 -35 52 -33
rect 65 -35 66 -33
rect 72 -35 73 -33
rect 100 -46 101 -34
rect 16 -37 17 -33
rect 30 -46 31 -36
rect 44 -37 45 -33
rect 51 -46 52 -36
rect 54 -37 55 -33
rect 58 -37 59 -33
rect 75 -37 76 -33
rect 86 -37 87 -33
rect 16 -46 17 -38
rect 23 -39 24 -33
rect 33 -39 34 -33
rect 44 -46 45 -38
rect 75 -46 76 -38
rect 86 -46 87 -38
rect 23 -46 24 -40
rect 33 -46 34 -40
rect 37 -41 38 -33
rect 58 -46 59 -40
rect 79 -41 80 -33
rect 93 -41 94 -33
rect 68 -46 69 -42
rect 93 -46 94 -42
rect 72 -46 73 -44
rect 79 -46 80 -44
rect 12 -67 13 -55
rect 54 -67 55 -55
rect 61 -67 62 -55
rect 86 -56 87 -54
rect 16 -58 17 -54
rect 37 -58 38 -54
rect 40 -58 41 -54
rect 51 -58 52 -54
rect 65 -58 66 -54
rect 100 -58 101 -54
rect 16 -67 17 -59
rect 23 -60 24 -54
rect 30 -60 31 -54
rect 33 -67 34 -59
rect 37 -67 38 -59
rect 68 -60 69 -54
rect 75 -67 76 -59
rect 107 -67 108 -59
rect 23 -67 24 -61
rect 30 -67 31 -61
rect 44 -62 45 -54
rect 44 -67 45 -61
rect 44 -62 45 -54
rect 44 -67 45 -61
rect 51 -67 52 -61
rect 58 -62 59 -54
rect 65 -67 66 -61
rect 93 -62 94 -54
rect 100 -67 101 -61
rect 117 -67 118 -61
rect 79 -64 80 -54
rect 93 -67 94 -63
rect 40 -67 41 -65
rect 79 -67 80 -65
rect 86 -67 87 -65
rect 114 -67 115 -65
rect 2 -94 3 -76
rect 16 -77 17 -75
rect 19 -94 20 -76
rect 23 -77 24 -75
rect 30 -77 31 -75
rect 37 -94 38 -76
rect 51 -77 52 -75
rect 100 -77 101 -75
rect 107 -77 108 -75
rect 114 -77 115 -75
rect 9 -94 10 -78
rect 33 -79 34 -75
rect 54 -79 55 -75
rect 121 -94 122 -78
rect 16 -94 17 -80
rect 86 -81 87 -75
rect 23 -94 24 -82
rect 54 -94 55 -82
rect 58 -83 59 -75
rect 68 -83 69 -75
rect 75 -83 76 -75
rect 93 -83 94 -75
rect 44 -85 45 -75
rect 93 -94 94 -84
rect 58 -94 59 -86
rect 72 -94 73 -86
rect 79 -87 80 -75
rect 107 -94 108 -86
rect 61 -94 62 -88
rect 100 -94 101 -88
rect 65 -94 66 -90
rect 86 -94 87 -90
rect 68 -94 69 -92
rect 114 -94 115 -92
rect 2 -104 3 -102
rect 23 -104 24 -102
rect 37 -104 38 -102
rect 44 -104 45 -102
rect 47 -104 48 -102
rect 72 -104 73 -102
rect 79 -104 80 -102
rect 100 -104 101 -102
rect 9 -106 10 -102
rect 33 -106 34 -102
rect 37 -119 38 -105
rect 86 -106 87 -102
rect 16 -119 17 -107
rect 58 -108 59 -102
rect 65 -108 66 -102
rect 79 -119 80 -107
rect 86 -119 87 -107
rect 114 -108 115 -102
rect 44 -119 45 -109
rect 54 -110 55 -102
rect 61 -119 62 -109
rect 65 -119 66 -109
rect 68 -110 69 -102
rect 72 -119 73 -109
rect 30 -112 31 -102
rect 54 -119 55 -111
rect 68 -119 69 -111
rect 107 -112 108 -102
rect 30 -119 31 -113
rect 47 -119 48 -113
rect 51 -114 52 -102
rect 121 -114 122 -102
rect 51 -119 52 -115
rect 93 -116 94 -102
rect 93 -119 94 -117
rect 103 -119 104 -117
rect 2 -140 3 -128
rect 19 -140 20 -128
rect 65 -129 66 -127
rect 79 -129 80 -127
rect 86 -140 87 -128
rect 100 -129 101 -127
rect 16 -131 17 -127
rect 26 -131 27 -127
rect 30 -131 31 -127
rect 65 -140 66 -130
rect 68 -131 69 -127
rect 93 -131 94 -127
rect 9 -140 10 -132
rect 30 -140 31 -132
rect 72 -133 73 -127
rect 72 -140 73 -132
rect 72 -133 73 -127
rect 72 -140 73 -132
rect 26 -140 27 -134
rect 58 -135 59 -127
rect 37 -137 38 -127
rect 58 -140 59 -136
rect 37 -140 38 -138
rect 44 -140 45 -138
rect 2 -150 3 -148
rect 23 -150 24 -148
rect 33 -150 34 -148
rect 37 -150 38 -148
rect 44 -150 45 -148
rect 65 -150 66 -148
rect 72 -150 73 -148
rect 82 -150 83 -148
rect 9 -152 10 -148
rect 51 -152 52 -148
rect 54 -152 55 -148
rect 58 -152 59 -148
rect 79 -152 80 -148
rect 86 -152 87 -148
<< labels >>
rlabel pdiffusion 3 -4 3 -4 0 cellNo=19
rlabel pdiffusion 10 -4 10 -4 0 cellNo=35
rlabel pdiffusion 45 -4 45 -4 0 cellNo=6
rlabel pdiffusion 52 -4 52 -4 0 cellNo=27
rlabel pdiffusion 87 -4 87 -4 0 cellNo=7
rlabel pdiffusion 3 -15 3 -15 0 cellNo=25
rlabel pdiffusion 24 -15 24 -15 0 cellNo=22
rlabel pdiffusion 31 -15 31 -15 0 feedthrough
rlabel pdiffusion 38 -15 38 -15 0 cellNo=50
rlabel pdiffusion 59 -15 59 -15 0 feedthrough
rlabel pdiffusion 66 -15 66 -15 0 cellNo=8
rlabel pdiffusion 87 -15 87 -15 0 cellNo=46
rlabel pdiffusion 94 -15 94 -15 0 feedthrough
rlabel pdiffusion 10 -30 10 -30 0 cellNo=21
rlabel pdiffusion 17 -30 17 -30 0 feedthrough
rlabel pdiffusion 24 -30 24 -30 0 cellNo=28
rlabel pdiffusion 31 -30 31 -30 0 cellNo=20
rlabel pdiffusion 38 -30 38 -30 0 feedthrough
rlabel pdiffusion 45 -30 45 -30 0 feedthrough
rlabel pdiffusion 52 -30 52 -30 0 cellNo=2
rlabel pdiffusion 59 -30 59 -30 0 feedthrough
rlabel pdiffusion 66 -30 66 -30 0 feedthrough
rlabel pdiffusion 73 -30 73 -30 0 cellNo=1
rlabel pdiffusion 80 -30 80 -30 0 cellNo=9
rlabel pdiffusion 87 -30 87 -30 0 feedthrough
rlabel pdiffusion 94 -30 94 -30 0 feedthrough
rlabel pdiffusion 17 -51 17 -51 0 feedthrough
rlabel pdiffusion 24 -51 24 -51 0 feedthrough
rlabel pdiffusion 31 -51 31 -51 0 cellNo=5
rlabel pdiffusion 38 -51 38 -51 0 cellNo=17
rlabel pdiffusion 45 -51 45 -51 0 cellNo=29
rlabel pdiffusion 52 -51 52 -51 0 feedthrough
rlabel pdiffusion 59 -51 59 -51 0 feedthrough
rlabel pdiffusion 66 -51 66 -51 0 cellNo=13
rlabel pdiffusion 73 -51 73 -51 0 cellNo=47
rlabel pdiffusion 80 -51 80 -51 0 feedthrough
rlabel pdiffusion 87 -51 87 -51 0 feedthrough
rlabel pdiffusion 94 -51 94 -51 0 feedthrough
rlabel pdiffusion 101 -51 101 -51 0 feedthrough
rlabel pdiffusion 10 -72 10 -72 0 cellNo=12
rlabel pdiffusion 17 -72 17 -72 0 feedthrough
rlabel pdiffusion 24 -72 24 -72 0 feedthrough
rlabel pdiffusion 31 -72 31 -72 0 cellNo=44
rlabel pdiffusion 38 -72 38 -72 0 cellNo=26
rlabel pdiffusion 45 -72 45 -72 0 feedthrough
rlabel pdiffusion 52 -72 52 -72 0 cellNo=33
rlabel pdiffusion 59 -72 59 -72 0 cellNo=31
rlabel pdiffusion 66 -72 66 -72 0 cellNo=15
rlabel pdiffusion 73 -72 73 -72 0 cellNo=3
rlabel pdiffusion 80 -72 80 -72 0 feedthrough
rlabel pdiffusion 87 -72 87 -72 0 feedthrough
rlabel pdiffusion 94 -72 94 -72 0 feedthrough
rlabel pdiffusion 101 -72 101 -72 0 feedthrough
rlabel pdiffusion 108 -72 108 -72 0 feedthrough
rlabel pdiffusion 115 -72 115 -72 0 cellNo=14
rlabel pdiffusion 3 -99 3 -99 0 feedthrough
rlabel pdiffusion 10 -99 10 -99 0 feedthrough
rlabel pdiffusion 17 -99 17 -99 0 cellNo=34
rlabel pdiffusion 24 -99 24 -99 0 cellNo=30
rlabel pdiffusion 31 -99 31 -99 0 cellNo=43
rlabel pdiffusion 38 -99 38 -99 0 feedthrough
rlabel pdiffusion 45 -99 45 -99 0 cellNo=42
rlabel pdiffusion 52 -99 52 -99 0 cellNo=38
rlabel pdiffusion 59 -99 59 -99 0 cellNo=11
rlabel pdiffusion 66 -99 66 -99 0 cellNo=39
rlabel pdiffusion 73 -99 73 -99 0 feedthrough
rlabel pdiffusion 80 -99 80 -99 0 cellNo=48
rlabel pdiffusion 87 -99 87 -99 0 feedthrough
rlabel pdiffusion 94 -99 94 -99 0 feedthrough
rlabel pdiffusion 101 -99 101 -99 0 feedthrough
rlabel pdiffusion 108 -99 108 -99 0 feedthrough
rlabel pdiffusion 115 -99 115 -99 0 feedthrough
rlabel pdiffusion 122 -99 122 -99 0 feedthrough
rlabel pdiffusion 17 -124 17 -124 0 feedthrough
rlabel pdiffusion 24 -124 24 -124 0 cellNo=23
rlabel pdiffusion 31 -124 31 -124 0 feedthrough
rlabel pdiffusion 38 -124 38 -124 0 feedthrough
rlabel pdiffusion 45 -124 45 -124 0 cellNo=41
rlabel pdiffusion 52 -124 52 -124 0 cellNo=32
rlabel pdiffusion 59 -124 59 -124 0 cellNo=24
rlabel pdiffusion 66 -124 66 -124 0 cellNo=16
rlabel pdiffusion 73 -124 73 -124 0 feedthrough
rlabel pdiffusion 80 -124 80 -124 0 feedthrough
rlabel pdiffusion 87 -124 87 -124 0 cellNo=49
rlabel pdiffusion 94 -124 94 -124 0 feedthrough
rlabel pdiffusion 101 -124 101 -124 0 cellNo=37
rlabel pdiffusion 3 -145 3 -145 0 feedthrough
rlabel pdiffusion 10 -145 10 -145 0 feedthrough
rlabel pdiffusion 17 -145 17 -145 0 cellNo=10
rlabel pdiffusion 24 -145 24 -145 0 cellNo=36
rlabel pdiffusion 31 -145 31 -145 0 cellNo=18
rlabel pdiffusion 38 -145 38 -145 0 feedthrough
rlabel pdiffusion 45 -145 45 -145 0 cellNo=40
rlabel pdiffusion 52 -145 52 -145 0 cellNo=45
rlabel pdiffusion 59 -145 59 -145 0 feedthrough
rlabel pdiffusion 66 -145 66 -145 0 feedthrough
rlabel pdiffusion 73 -145 73 -145 0 feedthrough
rlabel pdiffusion 80 -145 80 -145 0 cellNo=4
rlabel pdiffusion 87 -145 87 -145 0 feedthrough
rlabel polysilicon 44 -6 44 -6 0 3
rlabel polysilicon 47 -6 47 -6 0 4
rlabel polysilicon 54 -6 54 -6 0 4
rlabel polysilicon 86 -6 86 -6 0 3
rlabel polysilicon 26 -17 26 -17 0 4
rlabel polysilicon 30 -11 30 -11 0 1
rlabel polysilicon 30 -17 30 -17 0 3
rlabel polysilicon 37 -11 37 -11 0 1
rlabel polysilicon 40 -11 40 -11 0 2
rlabel polysilicon 40 -17 40 -17 0 4
rlabel polysilicon 58 -11 58 -11 0 1
rlabel polysilicon 58 -17 58 -17 0 3
rlabel polysilicon 68 -11 68 -11 0 2
rlabel polysilicon 86 -17 86 -17 0 3
rlabel polysilicon 89 -17 89 -17 0 4
rlabel polysilicon 93 -11 93 -11 0 1
rlabel polysilicon 93 -17 93 -17 0 3
rlabel polysilicon 9 -26 9 -26 0 1
rlabel polysilicon 16 -26 16 -26 0 1
rlabel polysilicon 16 -32 16 -32 0 3
rlabel polysilicon 26 -26 26 -26 0 2
rlabel polysilicon 23 -32 23 -32 0 3
rlabel polysilicon 26 -32 26 -32 0 4
rlabel polysilicon 30 -26 30 -26 0 1
rlabel polysilicon 30 -32 30 -32 0 3
rlabel polysilicon 33 -32 33 -32 0 4
rlabel polysilicon 37 -26 37 -26 0 1
rlabel polysilicon 37 -32 37 -32 0 3
rlabel polysilicon 44 -26 44 -26 0 1
rlabel polysilicon 44 -32 44 -32 0 3
rlabel polysilicon 51 -32 51 -32 0 3
rlabel polysilicon 54 -32 54 -32 0 4
rlabel polysilicon 58 -26 58 -26 0 1
rlabel polysilicon 58 -32 58 -32 0 3
rlabel polysilicon 65 -26 65 -26 0 1
rlabel polysilicon 65 -32 65 -32 0 3
rlabel polysilicon 72 -32 72 -32 0 3
rlabel polysilicon 75 -32 75 -32 0 4
rlabel polysilicon 82 -26 82 -26 0 2
rlabel polysilicon 79 -32 79 -32 0 3
rlabel polysilicon 86 -26 86 -26 0 1
rlabel polysilicon 86 -32 86 -32 0 3
rlabel polysilicon 93 -26 93 -26 0 1
rlabel polysilicon 93 -32 93 -32 0 3
rlabel polysilicon 16 -47 16 -47 0 1
rlabel polysilicon 16 -53 16 -53 0 3
rlabel polysilicon 23 -47 23 -47 0 1
rlabel polysilicon 23 -53 23 -53 0 3
rlabel polysilicon 30 -47 30 -47 0 1
rlabel polysilicon 33 -47 33 -47 0 2
rlabel polysilicon 30 -53 30 -53 0 3
rlabel polysilicon 37 -53 37 -53 0 3
rlabel polysilicon 40 -53 40 -53 0 4
rlabel polysilicon 44 -47 44 -47 0 1
rlabel polysilicon 44 -53 44 -53 0 3
rlabel polysilicon 51 -47 51 -47 0 1
rlabel polysilicon 51 -53 51 -53 0 3
rlabel polysilicon 58 -47 58 -47 0 1
rlabel polysilicon 58 -53 58 -53 0 3
rlabel polysilicon 68 -47 68 -47 0 2
rlabel polysilicon 65 -53 65 -53 0 3
rlabel polysilicon 68 -53 68 -53 0 4
rlabel polysilicon 72 -47 72 -47 0 1
rlabel polysilicon 75 -47 75 -47 0 2
rlabel polysilicon 79 -47 79 -47 0 1
rlabel polysilicon 79 -53 79 -53 0 3
rlabel polysilicon 86 -47 86 -47 0 1
rlabel polysilicon 86 -53 86 -53 0 3
rlabel polysilicon 93 -47 93 -47 0 1
rlabel polysilicon 93 -53 93 -53 0 3
rlabel polysilicon 100 -47 100 -47 0 1
rlabel polysilicon 100 -53 100 -53 0 3
rlabel polysilicon 12 -68 12 -68 0 2
rlabel polysilicon 16 -68 16 -68 0 1
rlabel polysilicon 16 -74 16 -74 0 3
rlabel polysilicon 23 -68 23 -68 0 1
rlabel polysilicon 23 -74 23 -74 0 3
rlabel polysilicon 30 -68 30 -68 0 1
rlabel polysilicon 33 -68 33 -68 0 2
rlabel polysilicon 30 -74 30 -74 0 3
rlabel polysilicon 33 -74 33 -74 0 4
rlabel polysilicon 37 -68 37 -68 0 1
rlabel polysilicon 40 -68 40 -68 0 2
rlabel polysilicon 44 -68 44 -68 0 1
rlabel polysilicon 44 -74 44 -74 0 3
rlabel polysilicon 51 -68 51 -68 0 1
rlabel polysilicon 54 -68 54 -68 0 2
rlabel polysilicon 51 -74 51 -74 0 3
rlabel polysilicon 54 -74 54 -74 0 4
rlabel polysilicon 61 -68 61 -68 0 2
rlabel polysilicon 58 -74 58 -74 0 3
rlabel polysilicon 65 -68 65 -68 0 1
rlabel polysilicon 68 -74 68 -74 0 4
rlabel polysilicon 75 -68 75 -68 0 2
rlabel polysilicon 75 -74 75 -74 0 4
rlabel polysilicon 79 -68 79 -68 0 1
rlabel polysilicon 79 -74 79 -74 0 3
rlabel polysilicon 86 -68 86 -68 0 1
rlabel polysilicon 86 -74 86 -74 0 3
rlabel polysilicon 93 -68 93 -68 0 1
rlabel polysilicon 93 -74 93 -74 0 3
rlabel polysilicon 100 -68 100 -68 0 1
rlabel polysilicon 100 -74 100 -74 0 3
rlabel polysilicon 107 -68 107 -68 0 1
rlabel polysilicon 107 -74 107 -74 0 3
rlabel polysilicon 114 -68 114 -68 0 1
rlabel polysilicon 117 -68 117 -68 0 2
rlabel polysilicon 114 -74 114 -74 0 3
rlabel polysilicon 2 -95 2 -95 0 1
rlabel polysilicon 2 -101 2 -101 0 3
rlabel polysilicon 9 -95 9 -95 0 1
rlabel polysilicon 9 -101 9 -101 0 3
rlabel polysilicon 16 -95 16 -95 0 1
rlabel polysilicon 19 -95 19 -95 0 2
rlabel polysilicon 23 -95 23 -95 0 1
rlabel polysilicon 23 -101 23 -101 0 3
rlabel polysilicon 30 -101 30 -101 0 3
rlabel polysilicon 33 -101 33 -101 0 4
rlabel polysilicon 37 -95 37 -95 0 1
rlabel polysilicon 37 -101 37 -101 0 3
rlabel polysilicon 44 -101 44 -101 0 3
rlabel polysilicon 47 -101 47 -101 0 4
rlabel polysilicon 54 -95 54 -95 0 2
rlabel polysilicon 51 -101 51 -101 0 3
rlabel polysilicon 54 -101 54 -101 0 4
rlabel polysilicon 58 -95 58 -95 0 1
rlabel polysilicon 61 -95 61 -95 0 2
rlabel polysilicon 58 -101 58 -101 0 3
rlabel polysilicon 65 -95 65 -95 0 1
rlabel polysilicon 68 -95 68 -95 0 2
rlabel polysilicon 65 -101 65 -101 0 3
rlabel polysilicon 68 -101 68 -101 0 4
rlabel polysilicon 72 -95 72 -95 0 1
rlabel polysilicon 72 -101 72 -101 0 3
rlabel polysilicon 79 -101 79 -101 0 3
rlabel polysilicon 86 -95 86 -95 0 1
rlabel polysilicon 86 -101 86 -101 0 3
rlabel polysilicon 93 -95 93 -95 0 1
rlabel polysilicon 93 -101 93 -101 0 3
rlabel polysilicon 100 -95 100 -95 0 1
rlabel polysilicon 100 -101 100 -101 0 3
rlabel polysilicon 107 -95 107 -95 0 1
rlabel polysilicon 107 -101 107 -101 0 3
rlabel polysilicon 114 -95 114 -95 0 1
rlabel polysilicon 114 -101 114 -101 0 3
rlabel polysilicon 121 -95 121 -95 0 1
rlabel polysilicon 121 -101 121 -101 0 3
rlabel polysilicon 16 -120 16 -120 0 1
rlabel polysilicon 16 -126 16 -126 0 3
rlabel polysilicon 26 -126 26 -126 0 4
rlabel polysilicon 30 -120 30 -120 0 1
rlabel polysilicon 30 -126 30 -126 0 3
rlabel polysilicon 37 -120 37 -120 0 1
rlabel polysilicon 37 -126 37 -126 0 3
rlabel polysilicon 44 -120 44 -120 0 1
rlabel polysilicon 47 -120 47 -120 0 2
rlabel polysilicon 51 -120 51 -120 0 1
rlabel polysilicon 54 -120 54 -120 0 2
rlabel polysilicon 61 -120 61 -120 0 2
rlabel polysilicon 58 -126 58 -126 0 3
rlabel polysilicon 65 -120 65 -120 0 1
rlabel polysilicon 68 -120 68 -120 0 2
rlabel polysilicon 65 -126 65 -126 0 3
rlabel polysilicon 68 -126 68 -126 0 4
rlabel polysilicon 72 -120 72 -120 0 1
rlabel polysilicon 72 -126 72 -126 0 3
rlabel polysilicon 79 -120 79 -120 0 1
rlabel polysilicon 79 -126 79 -126 0 3
rlabel polysilicon 86 -120 86 -120 0 1
rlabel polysilicon 93 -120 93 -120 0 1
rlabel polysilicon 93 -126 93 -126 0 3
rlabel polysilicon 103 -120 103 -120 0 2
rlabel polysilicon 100 -126 100 -126 0 3
rlabel polysilicon 2 -141 2 -141 0 1
rlabel polysilicon 2 -147 2 -147 0 3
rlabel polysilicon 9 -141 9 -141 0 1
rlabel polysilicon 9 -147 9 -147 0 3
rlabel polysilicon 19 -141 19 -141 0 2
rlabel polysilicon 26 -141 26 -141 0 2
rlabel polysilicon 23 -147 23 -147 0 3
rlabel polysilicon 30 -141 30 -141 0 1
rlabel polysilicon 33 -147 33 -147 0 4
rlabel polysilicon 37 -141 37 -141 0 1
rlabel polysilicon 37 -147 37 -147 0 3
rlabel polysilicon 44 -141 44 -141 0 1
rlabel polysilicon 44 -147 44 -147 0 3
rlabel polysilicon 51 -147 51 -147 0 3
rlabel polysilicon 54 -147 54 -147 0 4
rlabel polysilicon 58 -141 58 -141 0 1
rlabel polysilicon 58 -147 58 -147 0 3
rlabel polysilicon 65 -141 65 -141 0 1
rlabel polysilicon 65 -147 65 -147 0 3
rlabel polysilicon 72 -141 72 -141 0 1
rlabel polysilicon 72 -147 72 -147 0 3
rlabel polysilicon 79 -147 79 -147 0 3
rlabel polysilicon 82 -147 82 -147 0 4
rlabel polysilicon 86 -141 86 -141 0 1
rlabel polysilicon 86 -147 86 -147 0 3
rlabel metal2 30 -8 30 -8 0 net=81
rlabel metal2 40 -8 40 -8 0 net=49
rlabel metal2 47 -8 47 -8 0 net=44
rlabel metal2 58 -8 58 -8 0 net=63
rlabel metal2 86 -8 86 -8 0 net=95
rlabel metal2 9 -19 9 -19 0 net=69
rlabel metal2 40 -19 40 -19 0 net=125
rlabel metal2 58 -19 58 -19 0 net=65
rlabel metal2 89 -19 89 -19 0 net=96
rlabel metal2 16 -21 16 -21 0 net=83
rlabel metal2 58 -21 58 -21 0 net=99
rlabel metal2 86 -21 86 -21 0 net=131
rlabel metal2 26 -23 26 -23 0 net=20
rlabel metal2 26 -23 26 -23 0 net=20
rlabel metal2 30 -23 30 -23 0 net=103
rlabel metal2 26 -34 26 -34 0 net=25
rlabel metal2 51 -34 51 -34 0 net=66
rlabel metal2 72 -34 72 -34 0 net=135
rlabel metal2 16 -36 16 -36 0 net=84
rlabel metal2 44 -36 44 -36 0 net=127
rlabel metal2 54 -36 54 -36 0 net=100
rlabel metal2 75 -36 75 -36 0 net=104
rlabel metal2 16 -38 16 -38 0 net=85
rlabel metal2 33 -38 33 -38 0 net=27
rlabel metal2 75 -38 75 -38 0 net=101
rlabel metal2 23 -40 23 -40 0 net=57
rlabel metal2 37 -40 37 -40 0 net=71
rlabel metal2 79 -40 79 -40 0 net=132
rlabel metal2 68 -42 68 -42 0 net=133
rlabel metal2 72 -44 72 -44 0 net=115
rlabel metal2 12 -55 12 -55 0 net=46
rlabel metal2 61 -55 61 -55 0 net=102
rlabel metal2 16 -57 16 -57 0 net=86
rlabel metal2 40 -57 40 -57 0 net=128
rlabel metal2 65 -57 65 -57 0 net=136
rlabel metal2 16 -59 16 -59 0 net=59
rlabel metal2 30 -59 30 -59 0 net=13
rlabel metal2 37 -59 37 -59 0 net=42
rlabel metal2 75 -59 75 -59 0 net=141
rlabel metal2 23 -61 23 -61 0 net=53
rlabel metal2 44 -61 44 -61 0 net=87
rlabel metal2 44 -61 44 -61 0 net=87
rlabel metal2 51 -61 51 -61 0 net=72
rlabel metal2 65 -61 65 -61 0 net=134
rlabel metal2 100 -61 100 -61 0 net=139
rlabel metal2 79 -63 79 -63 0 net=117
rlabel metal2 40 -65 40 -65 0 net=105
rlabel metal2 86 -65 86 -65 0 net=111
rlabel metal2 2 -76 2 -76 0 net=61
rlabel metal2 19 -76 19 -76 0 net=54
rlabel metal2 30 -76 30 -76 0 net=51
rlabel metal2 51 -76 51 -76 0 net=140
rlabel metal2 107 -76 107 -76 0 net=142
rlabel metal2 9 -78 9 -78 0 net=73
rlabel metal2 54 -78 54 -78 0 net=113
rlabel metal2 16 -80 16 -80 0 net=112
rlabel metal2 23 -82 23 -82 0 net=45
rlabel metal2 58 -82 58 -82 0 net=1
rlabel metal2 75 -82 75 -82 0 net=118
rlabel metal2 44 -84 44 -84 0 net=89
rlabel metal2 58 -86 58 -86 0 net=67
rlabel metal2 79 -86 79 -86 0 net=107
rlabel metal2 61 -88 61 -88 0 net=97
rlabel metal2 65 -90 65 -90 0 net=75
rlabel metal2 68 -92 68 -92 0 net=109
rlabel metal2 2 -103 2 -103 0 net=62
rlabel metal2 37 -103 37 -103 0 net=52
rlabel metal2 47 -103 47 -103 0 net=68
rlabel metal2 79 -103 79 -103 0 net=98
rlabel metal2 9 -105 9 -105 0 net=74
rlabel metal2 37 -105 37 -105 0 net=77
rlabel metal2 16 -107 16 -107 0 net=91
rlabel metal2 65 -107 65 -107 0 net=123
rlabel metal2 86 -107 86 -107 0 net=110
rlabel metal2 44 -109 44 -109 0 net=24
rlabel metal2 61 -109 61 -109 0 net=40
rlabel metal2 68 -109 68 -109 0 net=119
rlabel metal2 30 -111 30 -111 0 net=36
rlabel metal2 68 -111 68 -111 0 net=108
rlabel metal2 30 -113 30 -113 0 net=145
rlabel metal2 51 -113 51 -113 0 net=114
rlabel metal2 51 -115 51 -115 0 net=90
rlabel metal2 93 -117 93 -117 0 net=129
rlabel metal2 2 -128 2 -128 0 net=137
rlabel metal2 65 -128 65 -128 0 net=124
rlabel metal2 86 -128 86 -128 0 net=55
rlabel metal2 16 -130 16 -130 0 net=92
rlabel metal2 30 -130 30 -130 0 net=147
rlabel metal2 68 -130 68 -130 0 net=130
rlabel metal2 9 -132 9 -132 0 net=143
rlabel metal2 72 -132 72 -132 0 net=121
rlabel metal2 72 -132 72 -132 0 net=121
rlabel metal2 26 -134 26 -134 0 net=23
rlabel metal2 37 -136 37 -136 0 net=79
rlabel metal2 37 -138 37 -138 0 net=93
rlabel metal2 2 -149 2 -149 0 net=138
rlabel metal2 33 -149 33 -149 0 net=94
rlabel metal2 44 -149 44 -149 0 net=148
rlabel metal2 72 -149 72 -149 0 net=122
rlabel metal2 9 -151 9 -151 0 net=144
rlabel metal2 54 -151 54 -151 0 net=80
rlabel metal2 79 -151 79 -151 0 net=56
<< end >>
