magic
tech scmos
timestamp 1555071791 
<< pdiffusion >>
rect 1 -10 7 -4
rect 8 -10 14 -4
rect 15 -10 21 -4
rect 22 -10 28 -4
rect 29 -10 35 -4
rect 36 -10 42 -4
rect 176 -10 179 -4
rect 183 -10 189 -4
rect 190 -10 196 -4
rect 197 -10 203 -4
rect 204 -10 210 -4
rect 211 -10 214 -4
rect 253 -10 259 -4
rect 267 -10 273 -4
rect 274 -10 277 -4
rect 281 -10 284 -4
rect 309 -10 312 -4
rect 344 -10 350 -4
rect 358 -10 364 -4
rect 365 -10 368 -4
rect 1 -27 7 -21
rect 8 -27 14 -21
rect 15 -27 21 -21
rect 22 -27 28 -21
rect 29 -27 35 -21
rect 155 -27 161 -21
rect 197 -27 203 -21
rect 211 -27 217 -21
rect 218 -27 221 -21
rect 232 -27 235 -21
rect 239 -27 242 -21
rect 246 -27 252 -21
rect 253 -27 256 -21
rect 260 -27 263 -21
rect 267 -27 273 -21
rect 281 -27 284 -21
rect 295 -27 301 -21
rect 302 -27 305 -21
rect 330 -27 336 -21
rect 337 -27 343 -21
rect 365 -27 368 -21
rect 372 -27 375 -21
rect 379 -27 385 -21
rect 386 -27 389 -21
rect 393 -27 396 -21
rect 1 -48 7 -42
rect 8 -48 14 -42
rect 15 -48 21 -42
rect 22 -48 28 -42
rect 99 -48 105 -42
rect 106 -48 112 -42
rect 155 -48 158 -42
rect 162 -48 168 -42
rect 169 -48 175 -42
rect 176 -48 179 -42
rect 183 -48 189 -42
rect 190 -48 196 -42
rect 197 -48 200 -42
rect 204 -48 207 -42
rect 211 -48 217 -42
rect 218 -48 221 -42
rect 225 -48 228 -42
rect 232 -48 238 -42
rect 239 -48 242 -42
rect 246 -48 249 -42
rect 253 -48 259 -42
rect 260 -48 263 -42
rect 267 -48 270 -42
rect 274 -48 277 -42
rect 281 -48 284 -42
rect 288 -48 291 -42
rect 295 -48 301 -42
rect 302 -48 308 -42
rect 309 -48 312 -42
rect 316 -48 319 -42
rect 323 -48 326 -42
rect 330 -48 333 -42
rect 337 -48 343 -42
rect 344 -48 347 -42
rect 351 -48 354 -42
rect 358 -48 364 -42
rect 365 -48 368 -42
rect 372 -48 378 -42
rect 379 -48 385 -42
rect 386 -48 389 -42
rect 393 -48 396 -42
rect 400 -48 406 -42
rect 407 -48 413 -42
rect 414 -48 417 -42
rect 421 -48 424 -42
rect 428 -48 431 -42
rect 435 -48 441 -42
rect 442 -48 448 -42
rect 449 -48 452 -42
rect 1 -85 7 -79
rect 8 -85 14 -79
rect 15 -85 21 -79
rect 22 -85 28 -79
rect 85 -85 88 -79
rect 92 -85 95 -79
rect 99 -85 102 -79
rect 106 -85 112 -79
rect 113 -85 119 -79
rect 120 -85 126 -79
rect 127 -85 130 -79
rect 134 -85 137 -79
rect 141 -85 144 -79
rect 148 -85 151 -79
rect 155 -85 161 -79
rect 162 -85 165 -79
rect 169 -85 172 -79
rect 176 -85 179 -79
rect 183 -85 189 -79
rect 190 -85 193 -79
rect 197 -85 203 -79
rect 204 -85 207 -79
rect 211 -85 217 -79
rect 218 -85 224 -79
rect 225 -85 228 -79
rect 232 -85 238 -79
rect 239 -85 245 -79
rect 246 -85 249 -79
rect 253 -85 259 -79
rect 260 -85 263 -79
rect 267 -85 270 -79
rect 274 -85 277 -79
rect 281 -85 284 -79
rect 288 -85 291 -79
rect 295 -85 298 -79
rect 302 -85 305 -79
rect 309 -85 315 -79
rect 316 -85 319 -79
rect 323 -85 326 -79
rect 330 -85 333 -79
rect 337 -85 343 -79
rect 344 -85 350 -79
rect 351 -85 357 -79
rect 358 -85 364 -79
rect 365 -85 371 -79
rect 372 -85 375 -79
rect 379 -85 382 -79
rect 386 -85 389 -79
rect 393 -85 396 -79
rect 400 -85 403 -79
rect 407 -85 410 -79
rect 414 -85 417 -79
rect 421 -85 424 -79
rect 428 -85 431 -79
rect 435 -85 438 -79
rect 442 -85 445 -79
rect 449 -85 452 -79
rect 456 -85 459 -79
rect 463 -85 466 -79
rect 470 -85 473 -79
rect 477 -85 480 -79
rect 484 -85 487 -79
rect 491 -85 497 -79
rect 498 -85 501 -79
rect 505 -85 511 -79
rect 561 -85 567 -79
rect 575 -85 581 -79
rect 582 -85 585 -79
rect 1 -140 7 -134
rect 8 -140 14 -134
rect 15 -140 21 -134
rect 50 -140 56 -134
rect 57 -140 60 -134
rect 64 -140 67 -134
rect 71 -140 74 -134
rect 78 -140 81 -134
rect 85 -140 88 -134
rect 92 -140 95 -134
rect 99 -140 105 -134
rect 106 -140 109 -134
rect 113 -140 116 -134
rect 120 -140 123 -134
rect 127 -140 130 -134
rect 134 -140 137 -134
rect 141 -140 144 -134
rect 148 -140 151 -134
rect 155 -140 158 -134
rect 162 -140 165 -134
rect 169 -140 172 -134
rect 176 -140 182 -134
rect 183 -140 189 -134
rect 190 -140 196 -134
rect 197 -140 200 -134
rect 204 -140 207 -134
rect 211 -140 217 -134
rect 218 -140 224 -134
rect 225 -140 231 -134
rect 232 -140 235 -134
rect 239 -140 245 -134
rect 246 -140 249 -134
rect 253 -140 256 -134
rect 260 -140 263 -134
rect 267 -140 270 -134
rect 274 -140 277 -134
rect 281 -140 287 -134
rect 288 -140 291 -134
rect 295 -140 301 -134
rect 302 -140 308 -134
rect 309 -140 312 -134
rect 316 -140 319 -134
rect 323 -140 326 -134
rect 330 -140 336 -134
rect 337 -140 343 -134
rect 344 -140 347 -134
rect 351 -140 357 -134
rect 358 -140 364 -134
rect 365 -140 371 -134
rect 372 -140 378 -134
rect 379 -140 385 -134
rect 386 -140 392 -134
rect 393 -140 396 -134
rect 400 -140 403 -134
rect 407 -140 410 -134
rect 414 -140 417 -134
rect 421 -140 427 -134
rect 428 -140 431 -134
rect 435 -140 438 -134
rect 442 -140 445 -134
rect 449 -140 452 -134
rect 456 -140 459 -134
rect 463 -140 466 -134
rect 470 -140 473 -134
rect 477 -140 480 -134
rect 484 -140 487 -134
rect 491 -140 494 -134
rect 498 -140 501 -134
rect 505 -140 508 -134
rect 512 -140 515 -134
rect 519 -140 522 -134
rect 526 -140 529 -134
rect 533 -140 536 -134
rect 540 -140 543 -134
rect 547 -140 553 -134
rect 554 -140 557 -134
rect 561 -140 564 -134
rect 568 -140 571 -134
rect 575 -140 578 -134
rect 582 -140 585 -134
rect 589 -140 595 -134
rect 596 -140 599 -134
rect 617 -140 620 -134
rect 1 -199 7 -193
rect 8 -199 14 -193
rect 64 -199 67 -193
rect 71 -199 77 -193
rect 78 -199 81 -193
rect 85 -199 88 -193
rect 92 -199 95 -193
rect 99 -199 102 -193
rect 106 -199 109 -193
rect 113 -199 116 -193
rect 120 -199 123 -193
rect 127 -199 130 -193
rect 134 -199 140 -193
rect 141 -199 147 -193
rect 148 -199 151 -193
rect 155 -199 158 -193
rect 162 -199 165 -193
rect 169 -199 175 -193
rect 176 -199 179 -193
rect 183 -199 189 -193
rect 190 -199 196 -193
rect 197 -199 200 -193
rect 204 -199 210 -193
rect 211 -199 217 -193
rect 218 -199 221 -193
rect 225 -199 228 -193
rect 232 -199 238 -193
rect 239 -199 242 -193
rect 246 -199 249 -193
rect 253 -199 256 -193
rect 260 -199 263 -193
rect 267 -199 270 -193
rect 274 -199 277 -193
rect 281 -199 284 -193
rect 288 -199 291 -193
rect 295 -199 301 -193
rect 302 -199 308 -193
rect 309 -199 312 -193
rect 316 -199 322 -193
rect 323 -199 326 -193
rect 330 -199 333 -193
rect 337 -199 340 -193
rect 344 -199 347 -193
rect 351 -199 357 -193
rect 358 -199 364 -193
rect 365 -199 368 -193
rect 372 -199 378 -193
rect 379 -199 382 -193
rect 386 -199 389 -193
rect 393 -199 399 -193
rect 400 -199 406 -193
rect 407 -199 410 -193
rect 414 -199 417 -193
rect 421 -199 424 -193
rect 428 -199 431 -193
rect 435 -199 441 -193
rect 442 -199 445 -193
rect 449 -199 452 -193
rect 456 -199 462 -193
rect 463 -199 466 -193
rect 470 -199 473 -193
rect 477 -199 480 -193
rect 484 -199 487 -193
rect 491 -199 494 -193
rect 498 -199 501 -193
rect 505 -199 511 -193
rect 512 -199 515 -193
rect 519 -199 522 -193
rect 526 -199 529 -193
rect 533 -199 536 -193
rect 540 -199 546 -193
rect 547 -199 550 -193
rect 554 -199 557 -193
rect 561 -199 564 -193
rect 568 -199 574 -193
rect 575 -199 578 -193
rect 582 -199 585 -193
rect 589 -199 592 -193
rect 631 -199 634 -193
rect 638 -199 644 -193
rect 645 -199 648 -193
rect 1 -256 7 -250
rect 15 -256 18 -250
rect 22 -256 25 -250
rect 29 -256 32 -250
rect 36 -256 39 -250
rect 43 -256 46 -250
rect 50 -256 56 -250
rect 57 -256 60 -250
rect 64 -256 67 -250
rect 71 -256 74 -250
rect 78 -256 81 -250
rect 85 -256 88 -250
rect 92 -256 95 -250
rect 99 -256 105 -250
rect 106 -256 112 -250
rect 113 -256 116 -250
rect 120 -256 123 -250
rect 127 -256 133 -250
rect 134 -256 140 -250
rect 141 -256 147 -250
rect 148 -256 151 -250
rect 155 -256 161 -250
rect 162 -256 165 -250
rect 169 -256 172 -250
rect 176 -256 179 -250
rect 183 -256 186 -250
rect 190 -256 196 -250
rect 197 -256 200 -250
rect 204 -256 210 -250
rect 211 -256 217 -250
rect 218 -256 224 -250
rect 225 -256 231 -250
rect 232 -256 235 -250
rect 239 -256 242 -250
rect 246 -256 249 -250
rect 253 -256 256 -250
rect 260 -256 263 -250
rect 267 -256 273 -250
rect 274 -256 277 -250
rect 281 -256 284 -250
rect 288 -256 291 -250
rect 295 -256 298 -250
rect 302 -256 305 -250
rect 309 -256 312 -250
rect 316 -256 319 -250
rect 323 -256 326 -250
rect 330 -256 333 -250
rect 337 -256 343 -250
rect 344 -256 347 -250
rect 351 -256 354 -250
rect 358 -256 361 -250
rect 365 -256 368 -250
rect 372 -256 375 -250
rect 379 -256 382 -250
rect 386 -256 392 -250
rect 393 -256 399 -250
rect 400 -256 403 -250
rect 407 -256 413 -250
rect 414 -256 420 -250
rect 421 -256 424 -250
rect 428 -256 431 -250
rect 435 -256 438 -250
rect 442 -256 445 -250
rect 449 -256 452 -250
rect 456 -256 462 -250
rect 463 -256 469 -250
rect 470 -256 473 -250
rect 477 -256 483 -250
rect 484 -256 487 -250
rect 491 -256 494 -250
rect 498 -256 501 -250
rect 505 -256 511 -250
rect 512 -256 515 -250
rect 519 -256 522 -250
rect 526 -256 529 -250
rect 533 -256 536 -250
rect 540 -256 543 -250
rect 547 -256 550 -250
rect 554 -256 557 -250
rect 561 -256 564 -250
rect 568 -256 574 -250
rect 575 -256 578 -250
rect 582 -256 585 -250
rect 589 -256 592 -250
rect 596 -256 599 -250
rect 603 -256 606 -250
rect 610 -256 613 -250
rect 617 -256 620 -250
rect 624 -256 627 -250
rect 631 -256 634 -250
rect 638 -256 641 -250
rect 645 -256 648 -250
rect 652 -256 655 -250
rect 659 -256 662 -250
rect 666 -256 672 -250
rect 673 -256 676 -250
rect 680 -256 683 -250
rect 687 -256 690 -250
rect 694 -256 697 -250
rect 750 -256 753 -250
rect 855 -256 861 -250
rect 29 -309 32 -303
rect 36 -309 39 -303
rect 43 -309 49 -303
rect 50 -309 53 -303
rect 57 -309 60 -303
rect 64 -309 70 -303
rect 71 -309 74 -303
rect 78 -309 84 -303
rect 85 -309 88 -303
rect 92 -309 95 -303
rect 99 -309 105 -303
rect 106 -309 109 -303
rect 113 -309 119 -303
rect 120 -309 123 -303
rect 127 -309 130 -303
rect 134 -309 140 -303
rect 141 -309 144 -303
rect 148 -309 151 -303
rect 155 -309 158 -303
rect 162 -309 165 -303
rect 169 -309 172 -303
rect 176 -309 182 -303
rect 183 -309 186 -303
rect 190 -309 193 -303
rect 197 -309 200 -303
rect 204 -309 207 -303
rect 211 -309 217 -303
rect 218 -309 224 -303
rect 225 -309 228 -303
rect 232 -309 238 -303
rect 239 -309 245 -303
rect 246 -309 252 -303
rect 253 -309 259 -303
rect 260 -309 263 -303
rect 267 -309 270 -303
rect 274 -309 277 -303
rect 281 -309 284 -303
rect 288 -309 294 -303
rect 295 -309 301 -303
rect 302 -309 305 -303
rect 309 -309 312 -303
rect 316 -309 319 -303
rect 323 -309 326 -303
rect 330 -309 336 -303
rect 337 -309 343 -303
rect 344 -309 347 -303
rect 351 -309 354 -303
rect 358 -309 361 -303
rect 365 -309 368 -303
rect 372 -309 378 -303
rect 379 -309 382 -303
rect 386 -309 389 -303
rect 393 -309 399 -303
rect 400 -309 406 -303
rect 407 -309 410 -303
rect 414 -309 417 -303
rect 421 -309 427 -303
rect 428 -309 431 -303
rect 435 -309 441 -303
rect 442 -309 448 -303
rect 449 -309 452 -303
rect 456 -309 459 -303
rect 463 -309 466 -303
rect 470 -309 473 -303
rect 477 -309 480 -303
rect 484 -309 487 -303
rect 491 -309 494 -303
rect 498 -309 501 -303
rect 505 -309 508 -303
rect 512 -309 515 -303
rect 519 -309 522 -303
rect 526 -309 529 -303
rect 533 -309 536 -303
rect 540 -309 546 -303
rect 547 -309 550 -303
rect 554 -309 557 -303
rect 561 -309 567 -303
rect 568 -309 571 -303
rect 575 -309 578 -303
rect 582 -309 585 -303
rect 589 -309 592 -303
rect 596 -309 599 -303
rect 603 -309 606 -303
rect 610 -309 613 -303
rect 617 -309 620 -303
rect 624 -309 627 -303
rect 631 -309 634 -303
rect 638 -309 641 -303
rect 645 -309 648 -303
rect 652 -309 655 -303
rect 659 -309 662 -303
rect 666 -309 669 -303
rect 673 -309 679 -303
rect 680 -309 683 -303
rect 687 -309 690 -303
rect 694 -309 697 -303
rect 701 -309 704 -303
rect 708 -309 711 -303
rect 715 -309 718 -303
rect 722 -309 728 -303
rect 729 -309 732 -303
rect 736 -309 739 -303
rect 743 -309 746 -303
rect 750 -309 753 -303
rect 827 -309 830 -303
rect 855 -309 858 -303
rect 1 -380 4 -374
rect 8 -380 11 -374
rect 15 -380 18 -374
rect 22 -380 25 -374
rect 29 -380 32 -374
rect 36 -380 39 -374
rect 43 -380 46 -374
rect 50 -380 53 -374
rect 57 -380 60 -374
rect 64 -380 67 -374
rect 71 -380 77 -374
rect 78 -380 81 -374
rect 85 -380 88 -374
rect 92 -380 98 -374
rect 99 -380 102 -374
rect 106 -380 112 -374
rect 113 -380 116 -374
rect 120 -380 123 -374
rect 127 -380 133 -374
rect 134 -380 140 -374
rect 141 -380 147 -374
rect 148 -380 154 -374
rect 155 -380 158 -374
rect 162 -380 165 -374
rect 169 -380 172 -374
rect 176 -380 179 -374
rect 183 -380 186 -374
rect 190 -380 193 -374
rect 197 -380 203 -374
rect 204 -380 210 -374
rect 211 -380 217 -374
rect 218 -380 221 -374
rect 225 -380 228 -374
rect 232 -380 238 -374
rect 239 -380 242 -374
rect 246 -380 249 -374
rect 253 -380 256 -374
rect 260 -380 263 -374
rect 267 -380 270 -374
rect 274 -380 280 -374
rect 281 -380 284 -374
rect 288 -380 291 -374
rect 295 -380 298 -374
rect 302 -380 305 -374
rect 309 -380 312 -374
rect 316 -380 319 -374
rect 323 -380 329 -374
rect 330 -380 336 -374
rect 337 -380 340 -374
rect 344 -380 347 -374
rect 351 -380 354 -374
rect 358 -380 364 -374
rect 365 -380 371 -374
rect 372 -380 378 -374
rect 379 -380 382 -374
rect 386 -380 389 -374
rect 393 -380 396 -374
rect 400 -380 406 -374
rect 407 -380 410 -374
rect 414 -380 417 -374
rect 421 -380 427 -374
rect 428 -380 434 -374
rect 435 -380 438 -374
rect 442 -380 445 -374
rect 449 -380 452 -374
rect 456 -380 459 -374
rect 463 -380 466 -374
rect 470 -380 476 -374
rect 477 -380 480 -374
rect 484 -380 487 -374
rect 491 -380 497 -374
rect 498 -380 501 -374
rect 505 -380 511 -374
rect 512 -380 518 -374
rect 519 -380 522 -374
rect 526 -380 529 -374
rect 533 -380 536 -374
rect 540 -380 543 -374
rect 547 -380 550 -374
rect 554 -380 557 -374
rect 561 -380 564 -374
rect 568 -380 571 -374
rect 575 -380 578 -374
rect 582 -380 588 -374
rect 589 -380 592 -374
rect 596 -380 599 -374
rect 603 -380 609 -374
rect 610 -380 613 -374
rect 617 -380 620 -374
rect 624 -380 627 -374
rect 631 -380 634 -374
rect 638 -380 641 -374
rect 645 -380 648 -374
rect 652 -380 655 -374
rect 659 -380 662 -374
rect 666 -380 669 -374
rect 673 -380 676 -374
rect 680 -380 683 -374
rect 687 -380 690 -374
rect 694 -380 697 -374
rect 701 -380 704 -374
rect 708 -380 711 -374
rect 715 -380 718 -374
rect 722 -380 725 -374
rect 729 -380 732 -374
rect 736 -380 739 -374
rect 743 -380 746 -374
rect 750 -380 753 -374
rect 757 -380 760 -374
rect 764 -380 767 -374
rect 771 -380 774 -374
rect 778 -380 781 -374
rect 785 -380 788 -374
rect 792 -380 795 -374
rect 799 -380 802 -374
rect 806 -380 809 -374
rect 813 -380 816 -374
rect 820 -380 823 -374
rect 827 -380 830 -374
rect 834 -380 837 -374
rect 841 -380 844 -374
rect 848 -380 854 -374
rect 855 -380 858 -374
rect 862 -380 865 -374
rect 869 -380 872 -374
rect 876 -380 882 -374
rect 883 -380 889 -374
rect 890 -380 893 -374
rect 1 -469 4 -463
rect 8 -469 11 -463
rect 15 -469 18 -463
rect 22 -469 25 -463
rect 29 -469 32 -463
rect 36 -469 39 -463
rect 43 -469 49 -463
rect 50 -469 56 -463
rect 57 -469 60 -463
rect 64 -469 67 -463
rect 71 -469 74 -463
rect 78 -469 84 -463
rect 85 -469 88 -463
rect 92 -469 95 -463
rect 99 -469 105 -463
rect 106 -469 112 -463
rect 113 -469 119 -463
rect 120 -469 123 -463
rect 127 -469 130 -463
rect 134 -469 137 -463
rect 141 -469 144 -463
rect 148 -469 154 -463
rect 155 -469 161 -463
rect 162 -469 168 -463
rect 169 -469 172 -463
rect 176 -469 179 -463
rect 183 -469 186 -463
rect 190 -469 196 -463
rect 197 -469 203 -463
rect 204 -469 207 -463
rect 211 -469 217 -463
rect 218 -469 224 -463
rect 225 -469 228 -463
rect 232 -469 235 -463
rect 239 -469 245 -463
rect 246 -469 249 -463
rect 253 -469 256 -463
rect 260 -469 263 -463
rect 267 -469 270 -463
rect 274 -469 277 -463
rect 281 -469 284 -463
rect 288 -469 291 -463
rect 295 -469 301 -463
rect 302 -469 308 -463
rect 309 -469 312 -463
rect 316 -469 319 -463
rect 323 -469 326 -463
rect 330 -469 333 -463
rect 337 -469 340 -463
rect 344 -469 350 -463
rect 351 -469 354 -463
rect 358 -469 361 -463
rect 365 -469 371 -463
rect 372 -469 375 -463
rect 379 -469 385 -463
rect 386 -469 392 -463
rect 393 -469 396 -463
rect 400 -469 403 -463
rect 407 -469 410 -463
rect 414 -469 420 -463
rect 421 -469 424 -463
rect 428 -469 434 -463
rect 435 -469 441 -463
rect 442 -469 445 -463
rect 449 -469 452 -463
rect 456 -469 462 -463
rect 463 -469 466 -463
rect 470 -469 473 -463
rect 477 -469 480 -463
rect 484 -469 490 -463
rect 491 -469 494 -463
rect 498 -469 504 -463
rect 505 -469 511 -463
rect 512 -469 515 -463
rect 519 -469 525 -463
rect 526 -469 529 -463
rect 533 -469 536 -463
rect 540 -469 543 -463
rect 547 -469 550 -463
rect 554 -469 557 -463
rect 561 -469 564 -463
rect 568 -469 571 -463
rect 575 -469 578 -463
rect 582 -469 585 -463
rect 589 -469 592 -463
rect 596 -469 599 -463
rect 603 -469 606 -463
rect 610 -469 613 -463
rect 617 -469 623 -463
rect 624 -469 627 -463
rect 631 -469 634 -463
rect 638 -469 641 -463
rect 645 -469 648 -463
rect 652 -469 655 -463
rect 659 -469 662 -463
rect 666 -469 669 -463
rect 673 -469 676 -463
rect 680 -469 683 -463
rect 687 -469 690 -463
rect 694 -469 697 -463
rect 701 -469 704 -463
rect 708 -469 711 -463
rect 715 -469 718 -463
rect 722 -469 725 -463
rect 729 -469 732 -463
rect 736 -469 739 -463
rect 743 -469 746 -463
rect 750 -469 753 -463
rect 757 -469 760 -463
rect 764 -469 767 -463
rect 771 -469 774 -463
rect 778 -469 781 -463
rect 785 -469 788 -463
rect 792 -469 795 -463
rect 799 -469 802 -463
rect 806 -469 809 -463
rect 813 -469 816 -463
rect 820 -469 823 -463
rect 827 -469 830 -463
rect 834 -469 837 -463
rect 841 -469 844 -463
rect 848 -469 851 -463
rect 855 -469 858 -463
rect 862 -469 865 -463
rect 869 -469 872 -463
rect 876 -469 879 -463
rect 883 -469 886 -463
rect 890 -469 893 -463
rect 897 -469 900 -463
rect 904 -469 907 -463
rect 911 -469 914 -463
rect 918 -469 921 -463
rect 925 -469 928 -463
rect 932 -469 935 -463
rect 939 -469 942 -463
rect 946 -469 949 -463
rect 1 -556 4 -550
rect 8 -556 11 -550
rect 15 -556 18 -550
rect 22 -556 28 -550
rect 29 -556 32 -550
rect 36 -556 39 -550
rect 43 -556 49 -550
rect 50 -556 53 -550
rect 57 -556 60 -550
rect 64 -556 67 -550
rect 71 -556 74 -550
rect 78 -556 81 -550
rect 85 -556 88 -550
rect 92 -556 98 -550
rect 99 -556 102 -550
rect 106 -556 109 -550
rect 113 -556 116 -550
rect 120 -556 123 -550
rect 127 -556 130 -550
rect 134 -556 137 -550
rect 141 -556 147 -550
rect 148 -556 151 -550
rect 155 -556 161 -550
rect 162 -556 168 -550
rect 169 -556 172 -550
rect 176 -556 182 -550
rect 183 -556 186 -550
rect 190 -556 193 -550
rect 197 -556 200 -550
rect 204 -556 210 -550
rect 211 -556 217 -550
rect 218 -556 221 -550
rect 225 -556 228 -550
rect 232 -556 235 -550
rect 239 -556 245 -550
rect 246 -556 249 -550
rect 253 -556 256 -550
rect 260 -556 266 -550
rect 267 -556 270 -550
rect 274 -556 277 -550
rect 281 -556 284 -550
rect 288 -556 291 -550
rect 295 -556 298 -550
rect 302 -556 305 -550
rect 309 -556 315 -550
rect 316 -556 322 -550
rect 323 -556 326 -550
rect 330 -556 336 -550
rect 337 -556 343 -550
rect 344 -556 347 -550
rect 351 -556 354 -550
rect 358 -556 364 -550
rect 365 -556 368 -550
rect 372 -556 375 -550
rect 379 -556 382 -550
rect 386 -556 392 -550
rect 393 -556 396 -550
rect 400 -556 403 -550
rect 407 -556 410 -550
rect 414 -556 420 -550
rect 421 -556 427 -550
rect 428 -556 431 -550
rect 435 -556 438 -550
rect 442 -556 445 -550
rect 449 -556 455 -550
rect 456 -556 459 -550
rect 463 -556 466 -550
rect 470 -556 473 -550
rect 477 -556 483 -550
rect 484 -556 487 -550
rect 491 -556 497 -550
rect 498 -556 504 -550
rect 505 -556 511 -550
rect 512 -556 515 -550
rect 519 -556 525 -550
rect 526 -556 529 -550
rect 533 -556 536 -550
rect 540 -556 546 -550
rect 547 -556 550 -550
rect 554 -556 557 -550
rect 561 -556 564 -550
rect 568 -556 571 -550
rect 575 -556 578 -550
rect 582 -556 585 -550
rect 589 -556 592 -550
rect 596 -556 599 -550
rect 603 -556 609 -550
rect 610 -556 613 -550
rect 617 -556 620 -550
rect 624 -556 627 -550
rect 631 -556 634 -550
rect 638 -556 641 -550
rect 645 -556 651 -550
rect 652 -556 655 -550
rect 659 -556 662 -550
rect 666 -556 669 -550
rect 673 -556 676 -550
rect 680 -556 683 -550
rect 687 -556 690 -550
rect 694 -556 697 -550
rect 701 -556 704 -550
rect 708 -556 711 -550
rect 715 -556 718 -550
rect 722 -556 728 -550
rect 729 -556 732 -550
rect 736 -556 739 -550
rect 743 -556 746 -550
rect 750 -556 756 -550
rect 757 -556 760 -550
rect 764 -556 767 -550
rect 771 -556 774 -550
rect 778 -556 781 -550
rect 785 -556 788 -550
rect 792 -556 798 -550
rect 799 -556 802 -550
rect 806 -556 809 -550
rect 813 -556 816 -550
rect 820 -556 823 -550
rect 834 -556 837 -550
rect 855 -556 858 -550
rect 1 -639 4 -633
rect 8 -639 11 -633
rect 15 -639 18 -633
rect 22 -639 25 -633
rect 29 -639 32 -633
rect 36 -639 42 -633
rect 43 -639 46 -633
rect 50 -639 53 -633
rect 57 -639 63 -633
rect 64 -639 67 -633
rect 71 -639 74 -633
rect 78 -639 81 -633
rect 85 -639 91 -633
rect 92 -639 95 -633
rect 99 -639 105 -633
rect 106 -639 109 -633
rect 113 -639 116 -633
rect 120 -639 126 -633
rect 127 -639 133 -633
rect 134 -639 140 -633
rect 141 -639 147 -633
rect 148 -639 151 -633
rect 155 -639 158 -633
rect 162 -639 165 -633
rect 169 -639 175 -633
rect 176 -639 179 -633
rect 183 -639 186 -633
rect 190 -639 193 -633
rect 197 -639 200 -633
rect 204 -639 207 -633
rect 211 -639 217 -633
rect 218 -639 221 -633
rect 225 -639 231 -633
rect 232 -639 238 -633
rect 239 -639 245 -633
rect 246 -639 249 -633
rect 253 -639 256 -633
rect 260 -639 263 -633
rect 267 -639 270 -633
rect 274 -639 277 -633
rect 281 -639 284 -633
rect 288 -639 291 -633
rect 295 -639 298 -633
rect 302 -639 308 -633
rect 309 -639 315 -633
rect 316 -639 319 -633
rect 323 -639 326 -633
rect 330 -639 336 -633
rect 337 -639 343 -633
rect 344 -639 350 -633
rect 351 -639 354 -633
rect 358 -639 361 -633
rect 365 -639 368 -633
rect 372 -639 375 -633
rect 379 -639 382 -633
rect 386 -639 389 -633
rect 393 -639 396 -633
rect 400 -639 406 -633
rect 407 -639 410 -633
rect 414 -639 417 -633
rect 421 -639 424 -633
rect 428 -639 431 -633
rect 435 -639 438 -633
rect 442 -639 445 -633
rect 449 -639 455 -633
rect 456 -639 459 -633
rect 463 -639 469 -633
rect 470 -639 476 -633
rect 477 -639 480 -633
rect 484 -639 487 -633
rect 491 -639 494 -633
rect 498 -639 501 -633
rect 505 -639 508 -633
rect 512 -639 515 -633
rect 519 -639 525 -633
rect 526 -639 529 -633
rect 533 -639 539 -633
rect 540 -639 546 -633
rect 547 -639 550 -633
rect 554 -639 557 -633
rect 561 -639 564 -633
rect 568 -639 571 -633
rect 575 -639 578 -633
rect 582 -639 585 -633
rect 589 -639 595 -633
rect 596 -639 602 -633
rect 603 -639 606 -633
rect 610 -639 616 -633
rect 617 -639 623 -633
rect 624 -639 627 -633
rect 631 -639 634 -633
rect 638 -639 641 -633
rect 645 -639 648 -633
rect 652 -639 655 -633
rect 659 -639 662 -633
rect 666 -639 669 -633
rect 673 -639 676 -633
rect 680 -639 683 -633
rect 687 -639 690 -633
rect 694 -639 700 -633
rect 701 -639 704 -633
rect 708 -639 711 -633
rect 715 -639 718 -633
rect 722 -639 725 -633
rect 729 -639 732 -633
rect 736 -639 739 -633
rect 743 -639 746 -633
rect 750 -639 753 -633
rect 757 -639 760 -633
rect 764 -639 767 -633
rect 771 -639 774 -633
rect 778 -639 781 -633
rect 785 -639 788 -633
rect 792 -639 795 -633
rect 799 -639 802 -633
rect 806 -639 809 -633
rect 813 -639 816 -633
rect 820 -639 823 -633
rect 827 -639 830 -633
rect 834 -639 837 -633
rect 841 -639 844 -633
rect 848 -639 851 -633
rect 855 -639 858 -633
rect 862 -639 865 -633
rect 869 -639 872 -633
rect 876 -639 879 -633
rect 883 -639 886 -633
rect 890 -639 893 -633
rect 897 -639 900 -633
rect 904 -639 907 -633
rect 911 -639 914 -633
rect 918 -639 924 -633
rect 925 -639 928 -633
rect 946 -639 949 -633
rect 1 -718 4 -712
rect 8 -718 11 -712
rect 15 -718 18 -712
rect 22 -718 28 -712
rect 29 -718 35 -712
rect 36 -718 39 -712
rect 43 -718 46 -712
rect 50 -718 53 -712
rect 57 -718 60 -712
rect 64 -718 67 -712
rect 71 -718 74 -712
rect 78 -718 81 -712
rect 85 -718 91 -712
rect 92 -718 95 -712
rect 99 -718 105 -712
rect 106 -718 112 -712
rect 113 -718 116 -712
rect 120 -718 123 -712
rect 127 -718 133 -712
rect 134 -718 137 -712
rect 141 -718 147 -712
rect 148 -718 151 -712
rect 155 -718 158 -712
rect 162 -718 165 -712
rect 169 -718 172 -712
rect 176 -718 179 -712
rect 183 -718 186 -712
rect 190 -718 193 -712
rect 197 -718 200 -712
rect 204 -718 210 -712
rect 211 -718 217 -712
rect 218 -718 221 -712
rect 225 -718 231 -712
rect 232 -718 235 -712
rect 239 -718 245 -712
rect 246 -718 252 -712
rect 253 -718 256 -712
rect 260 -718 263 -712
rect 267 -718 270 -712
rect 274 -718 280 -712
rect 281 -718 284 -712
rect 288 -718 291 -712
rect 295 -718 298 -712
rect 302 -718 305 -712
rect 309 -718 312 -712
rect 316 -718 319 -712
rect 323 -718 326 -712
rect 330 -718 336 -712
rect 337 -718 340 -712
rect 344 -718 350 -712
rect 351 -718 354 -712
rect 358 -718 361 -712
rect 365 -718 368 -712
rect 372 -718 378 -712
rect 379 -718 382 -712
rect 386 -718 392 -712
rect 393 -718 399 -712
rect 400 -718 403 -712
rect 407 -718 413 -712
rect 414 -718 420 -712
rect 421 -718 424 -712
rect 428 -718 431 -712
rect 435 -718 438 -712
rect 442 -718 445 -712
rect 449 -718 452 -712
rect 456 -718 459 -712
rect 463 -718 466 -712
rect 470 -718 476 -712
rect 477 -718 483 -712
rect 484 -718 490 -712
rect 491 -718 494 -712
rect 498 -718 504 -712
rect 505 -718 508 -712
rect 512 -718 518 -712
rect 519 -718 522 -712
rect 526 -718 529 -712
rect 533 -718 536 -712
rect 540 -718 546 -712
rect 547 -718 553 -712
rect 554 -718 560 -712
rect 561 -718 567 -712
rect 568 -718 571 -712
rect 575 -718 578 -712
rect 582 -718 585 -712
rect 589 -718 595 -712
rect 596 -718 599 -712
rect 603 -718 606 -712
rect 610 -718 613 -712
rect 617 -718 620 -712
rect 624 -718 630 -712
rect 631 -718 634 -712
rect 638 -718 641 -712
rect 645 -718 648 -712
rect 652 -718 655 -712
rect 659 -718 662 -712
rect 666 -718 669 -712
rect 673 -718 676 -712
rect 680 -718 683 -712
rect 687 -718 690 -712
rect 694 -718 697 -712
rect 701 -718 704 -712
rect 708 -718 711 -712
rect 715 -718 718 -712
rect 722 -718 725 -712
rect 729 -718 732 -712
rect 736 -718 739 -712
rect 743 -718 746 -712
rect 750 -718 753 -712
rect 757 -718 760 -712
rect 764 -718 767 -712
rect 771 -718 774 -712
rect 778 -718 781 -712
rect 785 -718 788 -712
rect 792 -718 795 -712
rect 799 -718 802 -712
rect 806 -718 809 -712
rect 813 -718 816 -712
rect 820 -718 823 -712
rect 827 -718 830 -712
rect 834 -718 837 -712
rect 841 -718 844 -712
rect 848 -718 851 -712
rect 855 -718 858 -712
rect 862 -718 865 -712
rect 869 -718 872 -712
rect 876 -718 879 -712
rect 883 -718 889 -712
rect 890 -718 893 -712
rect 897 -718 900 -712
rect 904 -718 907 -712
rect 911 -718 914 -712
rect 918 -718 921 -712
rect 925 -718 928 -712
rect 953 -718 956 -712
rect 1030 -718 1033 -712
rect 22 -789 25 -783
rect 29 -789 32 -783
rect 36 -789 39 -783
rect 43 -789 46 -783
rect 50 -789 56 -783
rect 57 -789 60 -783
rect 64 -789 70 -783
rect 71 -789 77 -783
rect 78 -789 81 -783
rect 85 -789 88 -783
rect 92 -789 95 -783
rect 99 -789 102 -783
rect 106 -789 112 -783
rect 113 -789 119 -783
rect 120 -789 123 -783
rect 127 -789 130 -783
rect 134 -789 137 -783
rect 141 -789 144 -783
rect 148 -789 151 -783
rect 155 -789 158 -783
rect 162 -789 165 -783
rect 169 -789 172 -783
rect 176 -789 179 -783
rect 183 -789 189 -783
rect 190 -789 193 -783
rect 197 -789 200 -783
rect 204 -789 207 -783
rect 211 -789 217 -783
rect 218 -789 221 -783
rect 225 -789 231 -783
rect 232 -789 238 -783
rect 239 -789 245 -783
rect 246 -789 249 -783
rect 253 -789 256 -783
rect 260 -789 266 -783
rect 267 -789 270 -783
rect 274 -789 277 -783
rect 281 -789 284 -783
rect 288 -789 291 -783
rect 295 -789 298 -783
rect 302 -789 305 -783
rect 309 -789 315 -783
rect 316 -789 319 -783
rect 323 -789 326 -783
rect 330 -789 333 -783
rect 337 -789 343 -783
rect 344 -789 347 -783
rect 351 -789 357 -783
rect 358 -789 361 -783
rect 365 -789 368 -783
rect 372 -789 378 -783
rect 379 -789 382 -783
rect 386 -789 392 -783
rect 393 -789 396 -783
rect 400 -789 406 -783
rect 407 -789 410 -783
rect 414 -789 420 -783
rect 421 -789 427 -783
rect 428 -789 431 -783
rect 435 -789 438 -783
rect 442 -789 445 -783
rect 449 -789 452 -783
rect 456 -789 459 -783
rect 463 -789 466 -783
rect 470 -789 473 -783
rect 477 -789 480 -783
rect 484 -789 487 -783
rect 491 -789 497 -783
rect 498 -789 501 -783
rect 505 -789 508 -783
rect 512 -789 518 -783
rect 519 -789 522 -783
rect 526 -789 532 -783
rect 533 -789 536 -783
rect 540 -789 546 -783
rect 547 -789 550 -783
rect 554 -789 560 -783
rect 561 -789 567 -783
rect 568 -789 571 -783
rect 575 -789 581 -783
rect 582 -789 585 -783
rect 589 -789 592 -783
rect 596 -789 599 -783
rect 603 -789 606 -783
rect 610 -789 613 -783
rect 617 -789 623 -783
rect 624 -789 627 -783
rect 631 -789 634 -783
rect 638 -789 641 -783
rect 645 -789 648 -783
rect 652 -789 655 -783
rect 659 -789 662 -783
rect 666 -789 672 -783
rect 673 -789 676 -783
rect 680 -789 683 -783
rect 687 -789 690 -783
rect 694 -789 697 -783
rect 701 -789 704 -783
rect 708 -789 711 -783
rect 715 -789 718 -783
rect 722 -789 725 -783
rect 729 -789 732 -783
rect 736 -789 739 -783
rect 743 -789 746 -783
rect 750 -789 753 -783
rect 757 -789 760 -783
rect 764 -789 767 -783
rect 771 -789 774 -783
rect 778 -789 781 -783
rect 785 -789 788 -783
rect 792 -789 795 -783
rect 799 -789 802 -783
rect 806 -789 809 -783
rect 813 -789 816 -783
rect 820 -789 823 -783
rect 827 -789 830 -783
rect 834 -789 837 -783
rect 841 -789 844 -783
rect 848 -789 851 -783
rect 855 -789 858 -783
rect 862 -789 865 -783
rect 869 -789 872 -783
rect 876 -789 879 -783
rect 883 -789 886 -783
rect 890 -789 896 -783
rect 897 -789 900 -783
rect 904 -789 910 -783
rect 911 -789 917 -783
rect 918 -789 921 -783
rect 960 -789 963 -783
rect 974 -789 977 -783
rect 988 -789 994 -783
rect 1002 -789 1008 -783
rect 1009 -789 1012 -783
rect 1016 -789 1019 -783
rect 1065 -789 1068 -783
rect 1 -886 4 -880
rect 8 -886 14 -880
rect 15 -886 18 -880
rect 22 -886 25 -880
rect 29 -886 32 -880
rect 36 -886 39 -880
rect 43 -886 49 -880
rect 50 -886 53 -880
rect 57 -886 60 -880
rect 64 -886 70 -880
rect 71 -886 74 -880
rect 78 -886 81 -880
rect 85 -886 88 -880
rect 92 -886 95 -880
rect 99 -886 102 -880
rect 106 -886 112 -880
rect 113 -886 119 -880
rect 120 -886 123 -880
rect 127 -886 133 -880
rect 134 -886 140 -880
rect 141 -886 144 -880
rect 148 -886 151 -880
rect 155 -886 158 -880
rect 162 -886 165 -880
rect 169 -886 175 -880
rect 176 -886 182 -880
rect 183 -886 186 -880
rect 190 -886 193 -880
rect 197 -886 200 -880
rect 204 -886 210 -880
rect 211 -886 217 -880
rect 218 -886 224 -880
rect 225 -886 231 -880
rect 232 -886 235 -880
rect 239 -886 245 -880
rect 246 -886 249 -880
rect 253 -886 256 -880
rect 260 -886 263 -880
rect 267 -886 270 -880
rect 274 -886 277 -880
rect 281 -886 284 -880
rect 288 -886 291 -880
rect 295 -886 298 -880
rect 302 -886 305 -880
rect 309 -886 312 -880
rect 316 -886 319 -880
rect 323 -886 326 -880
rect 330 -886 333 -880
rect 337 -886 340 -880
rect 344 -886 347 -880
rect 351 -886 357 -880
rect 358 -886 364 -880
rect 365 -886 371 -880
rect 372 -886 375 -880
rect 379 -886 382 -880
rect 386 -886 389 -880
rect 393 -886 396 -880
rect 400 -886 403 -880
rect 407 -886 413 -880
rect 414 -886 420 -880
rect 421 -886 424 -880
rect 428 -886 431 -880
rect 435 -886 441 -880
rect 442 -886 445 -880
rect 449 -886 452 -880
rect 456 -886 459 -880
rect 463 -886 469 -880
rect 470 -886 473 -880
rect 477 -886 480 -880
rect 484 -886 487 -880
rect 491 -886 497 -880
rect 498 -886 504 -880
rect 505 -886 508 -880
rect 512 -886 515 -880
rect 519 -886 525 -880
rect 526 -886 529 -880
rect 533 -886 539 -880
rect 540 -886 546 -880
rect 547 -886 553 -880
rect 554 -886 557 -880
rect 561 -886 567 -880
rect 568 -886 574 -880
rect 575 -886 578 -880
rect 582 -886 585 -880
rect 589 -886 592 -880
rect 596 -886 599 -880
rect 603 -886 606 -880
rect 610 -886 613 -880
rect 617 -886 620 -880
rect 624 -886 627 -880
rect 631 -886 634 -880
rect 638 -886 641 -880
rect 645 -886 648 -880
rect 652 -886 655 -880
rect 659 -886 662 -880
rect 666 -886 672 -880
rect 673 -886 676 -880
rect 680 -886 683 -880
rect 687 -886 690 -880
rect 694 -886 697 -880
rect 701 -886 704 -880
rect 708 -886 711 -880
rect 715 -886 718 -880
rect 722 -886 725 -880
rect 729 -886 732 -880
rect 736 -886 739 -880
rect 743 -886 746 -880
rect 750 -886 753 -880
rect 757 -886 760 -880
rect 764 -886 767 -880
rect 771 -886 774 -880
rect 778 -886 781 -880
rect 785 -886 788 -880
rect 792 -886 795 -880
rect 799 -886 802 -880
rect 806 -886 809 -880
rect 813 -886 819 -880
rect 820 -886 823 -880
rect 827 -886 830 -880
rect 834 -886 837 -880
rect 841 -886 844 -880
rect 848 -886 851 -880
rect 855 -886 858 -880
rect 862 -886 865 -880
rect 869 -886 872 -880
rect 876 -886 879 -880
rect 883 -886 886 -880
rect 890 -886 893 -880
rect 897 -886 900 -880
rect 904 -886 907 -880
rect 911 -886 914 -880
rect 918 -886 921 -880
rect 925 -886 928 -880
rect 932 -886 935 -880
rect 939 -886 942 -880
rect 946 -886 949 -880
rect 953 -886 956 -880
rect 960 -886 963 -880
rect 967 -886 970 -880
rect 974 -886 977 -880
rect 981 -886 984 -880
rect 988 -886 994 -880
rect 995 -886 998 -880
rect 1002 -886 1005 -880
rect 1009 -886 1015 -880
rect 1016 -886 1019 -880
rect 1023 -886 1026 -880
rect 1037 -886 1040 -880
rect 1079 -886 1082 -880
rect 8 -967 14 -961
rect 15 -967 18 -961
rect 22 -967 25 -961
rect 29 -967 32 -961
rect 36 -967 39 -961
rect 43 -967 46 -961
rect 50 -967 53 -961
rect 57 -967 60 -961
rect 64 -967 67 -961
rect 71 -967 74 -961
rect 78 -967 81 -961
rect 85 -967 88 -961
rect 92 -967 95 -961
rect 99 -967 102 -961
rect 106 -967 109 -961
rect 113 -967 116 -961
rect 120 -967 123 -961
rect 127 -967 133 -961
rect 134 -967 137 -961
rect 141 -967 144 -961
rect 148 -967 151 -961
rect 155 -967 158 -961
rect 162 -967 165 -961
rect 169 -967 172 -961
rect 176 -967 182 -961
rect 183 -967 186 -961
rect 190 -967 193 -961
rect 197 -967 200 -961
rect 204 -967 207 -961
rect 211 -967 217 -961
rect 218 -967 224 -961
rect 225 -967 231 -961
rect 232 -967 238 -961
rect 239 -967 245 -961
rect 246 -967 249 -961
rect 253 -967 256 -961
rect 260 -967 263 -961
rect 267 -967 270 -961
rect 274 -967 280 -961
rect 281 -967 287 -961
rect 288 -967 291 -961
rect 295 -967 298 -961
rect 302 -967 305 -961
rect 309 -967 312 -961
rect 316 -967 319 -961
rect 323 -967 329 -961
rect 330 -967 333 -961
rect 337 -967 340 -961
rect 344 -967 347 -961
rect 351 -967 354 -961
rect 358 -967 364 -961
rect 365 -967 368 -961
rect 372 -967 375 -961
rect 379 -967 385 -961
rect 386 -967 389 -961
rect 393 -967 399 -961
rect 400 -967 403 -961
rect 407 -967 410 -961
rect 414 -967 420 -961
rect 421 -967 424 -961
rect 428 -967 431 -961
rect 435 -967 441 -961
rect 442 -967 445 -961
rect 449 -967 455 -961
rect 456 -967 459 -961
rect 463 -967 466 -961
rect 470 -967 476 -961
rect 477 -967 483 -961
rect 484 -967 487 -961
rect 491 -967 497 -961
rect 498 -967 501 -961
rect 505 -967 508 -961
rect 512 -967 518 -961
rect 519 -967 522 -961
rect 526 -967 532 -961
rect 533 -967 536 -961
rect 540 -967 543 -961
rect 547 -967 550 -961
rect 554 -967 557 -961
rect 561 -967 567 -961
rect 568 -967 571 -961
rect 575 -967 578 -961
rect 582 -967 585 -961
rect 589 -967 592 -961
rect 596 -967 602 -961
rect 603 -967 609 -961
rect 610 -967 613 -961
rect 617 -967 623 -961
rect 624 -967 630 -961
rect 631 -967 637 -961
rect 638 -967 641 -961
rect 645 -967 648 -961
rect 652 -967 658 -961
rect 659 -967 662 -961
rect 666 -967 669 -961
rect 673 -967 676 -961
rect 680 -967 683 -961
rect 687 -967 690 -961
rect 694 -967 700 -961
rect 701 -967 704 -961
rect 708 -967 711 -961
rect 715 -967 718 -961
rect 722 -967 725 -961
rect 729 -967 732 -961
rect 736 -967 739 -961
rect 743 -967 746 -961
rect 750 -967 753 -961
rect 757 -967 760 -961
rect 764 -967 767 -961
rect 771 -967 774 -961
rect 778 -967 781 -961
rect 785 -967 788 -961
rect 792 -967 795 -961
rect 799 -967 802 -961
rect 806 -967 809 -961
rect 813 -967 816 -961
rect 820 -967 823 -961
rect 827 -967 830 -961
rect 834 -967 837 -961
rect 841 -967 844 -961
rect 848 -967 851 -961
rect 855 -967 858 -961
rect 862 -967 865 -961
rect 869 -967 872 -961
rect 876 -967 879 -961
rect 883 -967 886 -961
rect 890 -967 893 -961
rect 897 -967 900 -961
rect 904 -967 907 -961
rect 911 -967 917 -961
rect 918 -967 924 -961
rect 925 -967 931 -961
rect 932 -967 938 -961
rect 939 -967 945 -961
rect 946 -967 949 -961
rect 953 -967 956 -961
rect 960 -967 963 -961
rect 967 -967 970 -961
rect 981 -967 984 -961
rect 1009 -967 1012 -961
rect 1037 -967 1040 -961
rect 1058 -967 1061 -961
rect 1086 -967 1089 -961
rect 8 -1060 11 -1054
rect 15 -1060 18 -1054
rect 22 -1060 25 -1054
rect 29 -1060 32 -1054
rect 36 -1060 42 -1054
rect 43 -1060 46 -1054
rect 50 -1060 53 -1054
rect 57 -1060 63 -1054
rect 64 -1060 67 -1054
rect 71 -1060 74 -1054
rect 78 -1060 81 -1054
rect 85 -1060 88 -1054
rect 92 -1060 95 -1054
rect 99 -1060 102 -1054
rect 106 -1060 109 -1054
rect 113 -1060 116 -1054
rect 120 -1060 123 -1054
rect 127 -1060 133 -1054
rect 134 -1060 137 -1054
rect 141 -1060 147 -1054
rect 148 -1060 151 -1054
rect 155 -1060 158 -1054
rect 162 -1060 168 -1054
rect 169 -1060 175 -1054
rect 176 -1060 182 -1054
rect 183 -1060 186 -1054
rect 190 -1060 193 -1054
rect 197 -1060 200 -1054
rect 204 -1060 210 -1054
rect 211 -1060 214 -1054
rect 218 -1060 224 -1054
rect 225 -1060 228 -1054
rect 232 -1060 235 -1054
rect 239 -1060 242 -1054
rect 246 -1060 249 -1054
rect 253 -1060 259 -1054
rect 260 -1060 263 -1054
rect 267 -1060 270 -1054
rect 274 -1060 277 -1054
rect 281 -1060 284 -1054
rect 288 -1060 291 -1054
rect 295 -1060 301 -1054
rect 302 -1060 305 -1054
rect 309 -1060 312 -1054
rect 316 -1060 319 -1054
rect 323 -1060 326 -1054
rect 330 -1060 333 -1054
rect 337 -1060 340 -1054
rect 344 -1060 347 -1054
rect 351 -1060 357 -1054
rect 358 -1060 361 -1054
rect 365 -1060 368 -1054
rect 372 -1060 375 -1054
rect 379 -1060 382 -1054
rect 386 -1060 389 -1054
rect 393 -1060 396 -1054
rect 400 -1060 403 -1054
rect 407 -1060 413 -1054
rect 414 -1060 417 -1054
rect 421 -1060 424 -1054
rect 428 -1060 434 -1054
rect 435 -1060 438 -1054
rect 442 -1060 448 -1054
rect 449 -1060 455 -1054
rect 456 -1060 459 -1054
rect 463 -1060 466 -1054
rect 470 -1060 476 -1054
rect 477 -1060 483 -1054
rect 484 -1060 490 -1054
rect 491 -1060 497 -1054
rect 498 -1060 501 -1054
rect 505 -1060 508 -1054
rect 512 -1060 518 -1054
rect 519 -1060 522 -1054
rect 526 -1060 529 -1054
rect 533 -1060 539 -1054
rect 540 -1060 543 -1054
rect 547 -1060 553 -1054
rect 554 -1060 557 -1054
rect 561 -1060 564 -1054
rect 568 -1060 574 -1054
rect 575 -1060 581 -1054
rect 582 -1060 588 -1054
rect 589 -1060 592 -1054
rect 596 -1060 599 -1054
rect 603 -1060 609 -1054
rect 610 -1060 613 -1054
rect 617 -1060 620 -1054
rect 624 -1060 630 -1054
rect 631 -1060 634 -1054
rect 638 -1060 641 -1054
rect 645 -1060 651 -1054
rect 652 -1060 655 -1054
rect 659 -1060 662 -1054
rect 666 -1060 669 -1054
rect 673 -1060 676 -1054
rect 680 -1060 683 -1054
rect 687 -1060 693 -1054
rect 694 -1060 697 -1054
rect 701 -1060 704 -1054
rect 708 -1060 711 -1054
rect 715 -1060 718 -1054
rect 722 -1060 725 -1054
rect 729 -1060 735 -1054
rect 736 -1060 739 -1054
rect 743 -1060 746 -1054
rect 750 -1060 753 -1054
rect 757 -1060 760 -1054
rect 764 -1060 767 -1054
rect 771 -1060 774 -1054
rect 778 -1060 781 -1054
rect 785 -1060 788 -1054
rect 792 -1060 795 -1054
rect 799 -1060 802 -1054
rect 806 -1060 809 -1054
rect 813 -1060 816 -1054
rect 820 -1060 823 -1054
rect 827 -1060 830 -1054
rect 834 -1060 837 -1054
rect 841 -1060 844 -1054
rect 848 -1060 851 -1054
rect 855 -1060 858 -1054
rect 862 -1060 865 -1054
rect 869 -1060 872 -1054
rect 876 -1060 879 -1054
rect 883 -1060 886 -1054
rect 890 -1060 893 -1054
rect 897 -1060 900 -1054
rect 904 -1060 907 -1054
rect 911 -1060 914 -1054
rect 918 -1060 921 -1054
rect 925 -1060 928 -1054
rect 932 -1060 935 -1054
rect 939 -1060 942 -1054
rect 946 -1060 949 -1054
rect 953 -1060 956 -1054
rect 960 -1060 963 -1054
rect 967 -1060 970 -1054
rect 974 -1060 977 -1054
rect 981 -1060 984 -1054
rect 988 -1060 991 -1054
rect 995 -1060 998 -1054
rect 1002 -1060 1005 -1054
rect 1009 -1060 1012 -1054
rect 1016 -1060 1019 -1054
rect 1023 -1060 1029 -1054
rect 1030 -1060 1033 -1054
rect 1037 -1060 1040 -1054
rect 1044 -1060 1047 -1054
rect 1051 -1060 1054 -1054
rect 1058 -1060 1061 -1054
rect 1065 -1060 1071 -1054
rect 1072 -1060 1078 -1054
rect 1079 -1060 1085 -1054
rect 1086 -1060 1089 -1054
rect 1093 -1060 1096 -1054
rect 1100 -1060 1103 -1054
rect 1 -1159 4 -1153
rect 8 -1159 14 -1153
rect 15 -1159 21 -1153
rect 22 -1159 25 -1153
rect 29 -1159 35 -1153
rect 36 -1159 39 -1153
rect 43 -1159 46 -1153
rect 50 -1159 53 -1153
rect 57 -1159 60 -1153
rect 64 -1159 67 -1153
rect 71 -1159 74 -1153
rect 78 -1159 84 -1153
rect 85 -1159 88 -1153
rect 92 -1159 95 -1153
rect 99 -1159 102 -1153
rect 106 -1159 109 -1153
rect 113 -1159 116 -1153
rect 120 -1159 123 -1153
rect 127 -1159 133 -1153
rect 134 -1159 137 -1153
rect 141 -1159 147 -1153
rect 148 -1159 151 -1153
rect 155 -1159 158 -1153
rect 162 -1159 165 -1153
rect 169 -1159 172 -1153
rect 176 -1159 179 -1153
rect 183 -1159 189 -1153
rect 190 -1159 193 -1153
rect 197 -1159 200 -1153
rect 204 -1159 207 -1153
rect 211 -1159 214 -1153
rect 218 -1159 221 -1153
rect 225 -1159 231 -1153
rect 232 -1159 238 -1153
rect 239 -1159 245 -1153
rect 246 -1159 249 -1153
rect 253 -1159 256 -1153
rect 260 -1159 266 -1153
rect 267 -1159 270 -1153
rect 274 -1159 277 -1153
rect 281 -1159 284 -1153
rect 288 -1159 291 -1153
rect 295 -1159 298 -1153
rect 302 -1159 308 -1153
rect 309 -1159 312 -1153
rect 316 -1159 319 -1153
rect 323 -1159 326 -1153
rect 330 -1159 336 -1153
rect 337 -1159 340 -1153
rect 344 -1159 347 -1153
rect 351 -1159 357 -1153
rect 358 -1159 361 -1153
rect 365 -1159 371 -1153
rect 372 -1159 375 -1153
rect 379 -1159 382 -1153
rect 386 -1159 389 -1153
rect 393 -1159 396 -1153
rect 400 -1159 403 -1153
rect 407 -1159 410 -1153
rect 414 -1159 417 -1153
rect 421 -1159 424 -1153
rect 428 -1159 431 -1153
rect 435 -1159 441 -1153
rect 442 -1159 448 -1153
rect 449 -1159 452 -1153
rect 456 -1159 459 -1153
rect 463 -1159 469 -1153
rect 470 -1159 476 -1153
rect 477 -1159 480 -1153
rect 484 -1159 487 -1153
rect 491 -1159 497 -1153
rect 498 -1159 501 -1153
rect 505 -1159 511 -1153
rect 512 -1159 515 -1153
rect 519 -1159 522 -1153
rect 526 -1159 532 -1153
rect 533 -1159 536 -1153
rect 540 -1159 543 -1153
rect 547 -1159 550 -1153
rect 554 -1159 557 -1153
rect 561 -1159 564 -1153
rect 568 -1159 571 -1153
rect 575 -1159 578 -1153
rect 582 -1159 588 -1153
rect 589 -1159 595 -1153
rect 596 -1159 602 -1153
rect 603 -1159 609 -1153
rect 610 -1159 613 -1153
rect 617 -1159 623 -1153
rect 624 -1159 630 -1153
rect 631 -1159 634 -1153
rect 638 -1159 644 -1153
rect 645 -1159 648 -1153
rect 652 -1159 655 -1153
rect 659 -1159 665 -1153
rect 666 -1159 669 -1153
rect 673 -1159 679 -1153
rect 680 -1159 683 -1153
rect 687 -1159 693 -1153
rect 694 -1159 697 -1153
rect 701 -1159 704 -1153
rect 708 -1159 711 -1153
rect 715 -1159 718 -1153
rect 722 -1159 728 -1153
rect 729 -1159 735 -1153
rect 736 -1159 739 -1153
rect 743 -1159 746 -1153
rect 750 -1159 753 -1153
rect 757 -1159 760 -1153
rect 764 -1159 767 -1153
rect 771 -1159 774 -1153
rect 778 -1159 781 -1153
rect 785 -1159 788 -1153
rect 792 -1159 795 -1153
rect 799 -1159 802 -1153
rect 806 -1159 809 -1153
rect 813 -1159 816 -1153
rect 820 -1159 823 -1153
rect 827 -1159 830 -1153
rect 834 -1159 837 -1153
rect 841 -1159 844 -1153
rect 848 -1159 851 -1153
rect 855 -1159 858 -1153
rect 862 -1159 865 -1153
rect 869 -1159 872 -1153
rect 876 -1159 879 -1153
rect 883 -1159 886 -1153
rect 890 -1159 893 -1153
rect 897 -1159 900 -1153
rect 904 -1159 907 -1153
rect 911 -1159 914 -1153
rect 918 -1159 921 -1153
rect 925 -1159 928 -1153
rect 932 -1159 935 -1153
rect 939 -1159 942 -1153
rect 946 -1159 949 -1153
rect 953 -1159 956 -1153
rect 960 -1159 963 -1153
rect 967 -1159 970 -1153
rect 974 -1159 977 -1153
rect 981 -1159 984 -1153
rect 988 -1159 991 -1153
rect 995 -1159 998 -1153
rect 1002 -1159 1005 -1153
rect 1009 -1159 1012 -1153
rect 1016 -1159 1019 -1153
rect 1023 -1159 1026 -1153
rect 1030 -1159 1033 -1153
rect 1037 -1159 1040 -1153
rect 1044 -1159 1047 -1153
rect 1051 -1159 1054 -1153
rect 1058 -1159 1061 -1153
rect 1065 -1159 1068 -1153
rect 1072 -1159 1075 -1153
rect 1079 -1159 1082 -1153
rect 1086 -1159 1092 -1153
rect 1093 -1159 1096 -1153
rect 1100 -1159 1103 -1153
rect 1 -1262 4 -1256
rect 8 -1262 11 -1256
rect 15 -1262 21 -1256
rect 22 -1262 28 -1256
rect 29 -1262 32 -1256
rect 36 -1262 39 -1256
rect 43 -1262 46 -1256
rect 50 -1262 56 -1256
rect 57 -1262 60 -1256
rect 64 -1262 67 -1256
rect 71 -1262 74 -1256
rect 78 -1262 84 -1256
rect 85 -1262 88 -1256
rect 92 -1262 95 -1256
rect 99 -1262 102 -1256
rect 106 -1262 109 -1256
rect 113 -1262 119 -1256
rect 120 -1262 123 -1256
rect 127 -1262 130 -1256
rect 134 -1262 137 -1256
rect 141 -1262 144 -1256
rect 148 -1262 151 -1256
rect 155 -1262 158 -1256
rect 162 -1262 168 -1256
rect 169 -1262 175 -1256
rect 176 -1262 179 -1256
rect 183 -1262 189 -1256
rect 190 -1262 196 -1256
rect 197 -1262 203 -1256
rect 204 -1262 207 -1256
rect 211 -1262 217 -1256
rect 218 -1262 224 -1256
rect 225 -1262 228 -1256
rect 232 -1262 235 -1256
rect 239 -1262 242 -1256
rect 246 -1262 249 -1256
rect 253 -1262 256 -1256
rect 260 -1262 263 -1256
rect 267 -1262 270 -1256
rect 274 -1262 277 -1256
rect 281 -1262 284 -1256
rect 288 -1262 294 -1256
rect 295 -1262 298 -1256
rect 302 -1262 305 -1256
rect 309 -1262 312 -1256
rect 316 -1262 319 -1256
rect 323 -1262 326 -1256
rect 330 -1262 333 -1256
rect 337 -1262 340 -1256
rect 344 -1262 347 -1256
rect 351 -1262 354 -1256
rect 358 -1262 361 -1256
rect 365 -1262 368 -1256
rect 372 -1262 375 -1256
rect 379 -1262 382 -1256
rect 386 -1262 389 -1256
rect 393 -1262 396 -1256
rect 400 -1262 403 -1256
rect 407 -1262 410 -1256
rect 414 -1262 417 -1256
rect 421 -1262 427 -1256
rect 428 -1262 434 -1256
rect 435 -1262 438 -1256
rect 442 -1262 445 -1256
rect 449 -1262 452 -1256
rect 456 -1262 462 -1256
rect 463 -1262 466 -1256
rect 470 -1262 476 -1256
rect 477 -1262 480 -1256
rect 484 -1262 487 -1256
rect 491 -1262 497 -1256
rect 498 -1262 504 -1256
rect 505 -1262 508 -1256
rect 512 -1262 518 -1256
rect 519 -1262 525 -1256
rect 526 -1262 529 -1256
rect 533 -1262 539 -1256
rect 540 -1262 546 -1256
rect 547 -1262 553 -1256
rect 554 -1262 557 -1256
rect 561 -1262 567 -1256
rect 568 -1262 571 -1256
rect 575 -1262 578 -1256
rect 582 -1262 588 -1256
rect 589 -1262 595 -1256
rect 596 -1262 599 -1256
rect 603 -1262 609 -1256
rect 610 -1262 613 -1256
rect 617 -1262 620 -1256
rect 624 -1262 627 -1256
rect 631 -1262 634 -1256
rect 638 -1262 641 -1256
rect 645 -1262 648 -1256
rect 652 -1262 658 -1256
rect 659 -1262 662 -1256
rect 666 -1262 669 -1256
rect 673 -1262 676 -1256
rect 680 -1262 686 -1256
rect 687 -1262 690 -1256
rect 694 -1262 697 -1256
rect 701 -1262 704 -1256
rect 708 -1262 711 -1256
rect 715 -1262 721 -1256
rect 722 -1262 725 -1256
rect 729 -1262 732 -1256
rect 736 -1262 739 -1256
rect 743 -1262 746 -1256
rect 750 -1262 753 -1256
rect 757 -1262 760 -1256
rect 764 -1262 767 -1256
rect 771 -1262 774 -1256
rect 778 -1262 784 -1256
rect 785 -1262 788 -1256
rect 792 -1262 795 -1256
rect 799 -1262 802 -1256
rect 806 -1262 809 -1256
rect 813 -1262 819 -1256
rect 820 -1262 823 -1256
rect 827 -1262 830 -1256
rect 834 -1262 837 -1256
rect 841 -1262 844 -1256
rect 848 -1262 851 -1256
rect 855 -1262 858 -1256
rect 862 -1262 865 -1256
rect 869 -1262 872 -1256
rect 876 -1262 879 -1256
rect 883 -1262 886 -1256
rect 890 -1262 893 -1256
rect 897 -1262 900 -1256
rect 904 -1262 907 -1256
rect 911 -1262 914 -1256
rect 918 -1262 921 -1256
rect 925 -1262 928 -1256
rect 932 -1262 935 -1256
rect 939 -1262 942 -1256
rect 946 -1262 949 -1256
rect 953 -1262 956 -1256
rect 960 -1262 963 -1256
rect 967 -1262 970 -1256
rect 974 -1262 977 -1256
rect 981 -1262 984 -1256
rect 988 -1262 991 -1256
rect 995 -1262 998 -1256
rect 1002 -1262 1005 -1256
rect 1009 -1262 1012 -1256
rect 1016 -1262 1019 -1256
rect 1023 -1262 1026 -1256
rect 1030 -1262 1036 -1256
rect 1037 -1262 1043 -1256
rect 1044 -1262 1047 -1256
rect 1051 -1262 1054 -1256
rect 1058 -1262 1061 -1256
rect 1065 -1262 1068 -1256
rect 1072 -1262 1075 -1256
rect 8 -1341 11 -1335
rect 15 -1341 18 -1335
rect 22 -1341 25 -1335
rect 29 -1341 32 -1335
rect 36 -1341 39 -1335
rect 43 -1341 46 -1335
rect 50 -1341 53 -1335
rect 57 -1341 60 -1335
rect 64 -1341 67 -1335
rect 71 -1341 74 -1335
rect 78 -1341 84 -1335
rect 85 -1341 91 -1335
rect 92 -1341 95 -1335
rect 99 -1341 102 -1335
rect 106 -1341 109 -1335
rect 113 -1341 119 -1335
rect 120 -1341 123 -1335
rect 127 -1341 133 -1335
rect 134 -1341 140 -1335
rect 141 -1341 144 -1335
rect 148 -1341 151 -1335
rect 155 -1341 161 -1335
rect 162 -1341 165 -1335
rect 169 -1341 175 -1335
rect 176 -1341 182 -1335
rect 183 -1341 186 -1335
rect 190 -1341 196 -1335
rect 197 -1341 200 -1335
rect 204 -1341 207 -1335
rect 211 -1341 214 -1335
rect 218 -1341 224 -1335
rect 225 -1341 228 -1335
rect 232 -1341 235 -1335
rect 239 -1341 242 -1335
rect 246 -1341 249 -1335
rect 253 -1341 256 -1335
rect 260 -1341 263 -1335
rect 267 -1341 270 -1335
rect 274 -1341 277 -1335
rect 281 -1341 284 -1335
rect 288 -1341 294 -1335
rect 295 -1341 298 -1335
rect 302 -1341 305 -1335
rect 309 -1341 312 -1335
rect 316 -1341 322 -1335
rect 323 -1341 329 -1335
rect 330 -1341 333 -1335
rect 337 -1341 340 -1335
rect 344 -1341 347 -1335
rect 351 -1341 357 -1335
rect 358 -1341 361 -1335
rect 365 -1341 371 -1335
rect 372 -1341 375 -1335
rect 379 -1341 382 -1335
rect 386 -1341 389 -1335
rect 393 -1341 396 -1335
rect 400 -1341 403 -1335
rect 407 -1341 410 -1335
rect 414 -1341 417 -1335
rect 421 -1341 424 -1335
rect 428 -1341 434 -1335
rect 435 -1341 438 -1335
rect 442 -1341 445 -1335
rect 449 -1341 452 -1335
rect 456 -1341 462 -1335
rect 463 -1341 466 -1335
rect 470 -1341 476 -1335
rect 477 -1341 480 -1335
rect 484 -1341 487 -1335
rect 491 -1341 497 -1335
rect 498 -1341 501 -1335
rect 505 -1341 511 -1335
rect 512 -1341 515 -1335
rect 519 -1341 522 -1335
rect 526 -1341 529 -1335
rect 533 -1341 539 -1335
rect 540 -1341 543 -1335
rect 547 -1341 550 -1335
rect 554 -1341 557 -1335
rect 561 -1341 564 -1335
rect 568 -1341 571 -1335
rect 575 -1341 581 -1335
rect 582 -1341 588 -1335
rect 589 -1341 592 -1335
rect 596 -1341 602 -1335
rect 603 -1341 606 -1335
rect 610 -1341 613 -1335
rect 617 -1341 623 -1335
rect 624 -1341 627 -1335
rect 631 -1341 634 -1335
rect 638 -1341 641 -1335
rect 645 -1341 651 -1335
rect 652 -1341 655 -1335
rect 659 -1341 662 -1335
rect 666 -1341 669 -1335
rect 673 -1341 679 -1335
rect 680 -1341 683 -1335
rect 687 -1341 690 -1335
rect 694 -1341 697 -1335
rect 701 -1341 707 -1335
rect 708 -1341 711 -1335
rect 715 -1341 718 -1335
rect 722 -1341 725 -1335
rect 729 -1341 732 -1335
rect 736 -1341 742 -1335
rect 743 -1341 746 -1335
rect 750 -1341 753 -1335
rect 757 -1341 763 -1335
rect 764 -1341 767 -1335
rect 771 -1341 774 -1335
rect 778 -1341 781 -1335
rect 785 -1341 788 -1335
rect 792 -1341 795 -1335
rect 799 -1341 802 -1335
rect 806 -1341 809 -1335
rect 813 -1341 816 -1335
rect 820 -1341 823 -1335
rect 827 -1341 830 -1335
rect 834 -1341 837 -1335
rect 841 -1341 844 -1335
rect 848 -1341 851 -1335
rect 855 -1341 858 -1335
rect 862 -1341 865 -1335
rect 869 -1341 872 -1335
rect 876 -1341 879 -1335
rect 883 -1341 886 -1335
rect 890 -1341 893 -1335
rect 897 -1341 900 -1335
rect 904 -1341 907 -1335
rect 911 -1341 914 -1335
rect 918 -1341 921 -1335
rect 925 -1341 928 -1335
rect 932 -1341 935 -1335
rect 939 -1341 942 -1335
rect 946 -1341 949 -1335
rect 953 -1341 956 -1335
rect 960 -1341 963 -1335
rect 967 -1341 970 -1335
rect 974 -1341 977 -1335
rect 981 -1341 984 -1335
rect 988 -1341 991 -1335
rect 995 -1341 998 -1335
rect 1002 -1341 1005 -1335
rect 1009 -1341 1012 -1335
rect 1016 -1341 1019 -1335
rect 1023 -1341 1029 -1335
rect 1030 -1341 1036 -1335
rect 1037 -1341 1043 -1335
rect 1044 -1341 1050 -1335
rect 1051 -1341 1054 -1335
rect 1058 -1341 1064 -1335
rect 1065 -1341 1068 -1335
rect 1072 -1341 1075 -1335
rect 1079 -1341 1082 -1335
rect 15 -1418 18 -1412
rect 22 -1418 25 -1412
rect 29 -1418 32 -1412
rect 36 -1418 39 -1412
rect 43 -1418 46 -1412
rect 50 -1418 56 -1412
rect 57 -1418 63 -1412
rect 64 -1418 67 -1412
rect 71 -1418 74 -1412
rect 78 -1418 81 -1412
rect 85 -1418 91 -1412
rect 92 -1418 95 -1412
rect 99 -1418 102 -1412
rect 106 -1418 109 -1412
rect 113 -1418 116 -1412
rect 120 -1418 123 -1412
rect 127 -1418 130 -1412
rect 134 -1418 140 -1412
rect 141 -1418 147 -1412
rect 148 -1418 151 -1412
rect 155 -1418 161 -1412
rect 162 -1418 168 -1412
rect 169 -1418 172 -1412
rect 176 -1418 179 -1412
rect 183 -1418 186 -1412
rect 190 -1418 193 -1412
rect 197 -1418 200 -1412
rect 204 -1418 210 -1412
rect 211 -1418 214 -1412
rect 218 -1418 224 -1412
rect 225 -1418 228 -1412
rect 232 -1418 235 -1412
rect 239 -1418 245 -1412
rect 246 -1418 249 -1412
rect 253 -1418 256 -1412
rect 260 -1418 263 -1412
rect 267 -1418 270 -1412
rect 274 -1418 277 -1412
rect 281 -1418 284 -1412
rect 288 -1418 291 -1412
rect 295 -1418 298 -1412
rect 302 -1418 308 -1412
rect 309 -1418 312 -1412
rect 316 -1418 319 -1412
rect 323 -1418 326 -1412
rect 330 -1418 333 -1412
rect 337 -1418 340 -1412
rect 344 -1418 347 -1412
rect 351 -1418 357 -1412
rect 358 -1418 364 -1412
rect 365 -1418 368 -1412
rect 372 -1418 375 -1412
rect 379 -1418 382 -1412
rect 386 -1418 392 -1412
rect 393 -1418 396 -1412
rect 400 -1418 406 -1412
rect 407 -1418 413 -1412
rect 414 -1418 417 -1412
rect 421 -1418 424 -1412
rect 428 -1418 431 -1412
rect 435 -1418 438 -1412
rect 442 -1418 445 -1412
rect 449 -1418 452 -1412
rect 456 -1418 459 -1412
rect 463 -1418 466 -1412
rect 470 -1418 473 -1412
rect 477 -1418 480 -1412
rect 484 -1418 487 -1412
rect 491 -1418 494 -1412
rect 498 -1418 501 -1412
rect 505 -1418 511 -1412
rect 512 -1418 518 -1412
rect 519 -1418 525 -1412
rect 526 -1418 529 -1412
rect 533 -1418 536 -1412
rect 540 -1418 543 -1412
rect 547 -1418 550 -1412
rect 554 -1418 557 -1412
rect 561 -1418 567 -1412
rect 568 -1418 574 -1412
rect 575 -1418 581 -1412
rect 582 -1418 588 -1412
rect 589 -1418 592 -1412
rect 596 -1418 599 -1412
rect 603 -1418 606 -1412
rect 610 -1418 613 -1412
rect 617 -1418 620 -1412
rect 624 -1418 627 -1412
rect 631 -1418 634 -1412
rect 638 -1418 641 -1412
rect 645 -1418 648 -1412
rect 652 -1418 655 -1412
rect 659 -1418 665 -1412
rect 666 -1418 669 -1412
rect 673 -1418 676 -1412
rect 680 -1418 686 -1412
rect 687 -1418 690 -1412
rect 694 -1418 697 -1412
rect 701 -1418 707 -1412
rect 708 -1418 714 -1412
rect 715 -1418 718 -1412
rect 722 -1418 725 -1412
rect 729 -1418 732 -1412
rect 736 -1418 742 -1412
rect 743 -1418 746 -1412
rect 750 -1418 753 -1412
rect 757 -1418 760 -1412
rect 764 -1418 770 -1412
rect 771 -1418 774 -1412
rect 778 -1418 781 -1412
rect 785 -1418 788 -1412
rect 792 -1418 795 -1412
rect 799 -1418 802 -1412
rect 806 -1418 809 -1412
rect 813 -1418 816 -1412
rect 820 -1418 823 -1412
rect 827 -1418 830 -1412
rect 834 -1418 837 -1412
rect 841 -1418 844 -1412
rect 848 -1418 851 -1412
rect 855 -1418 858 -1412
rect 862 -1418 865 -1412
rect 869 -1418 872 -1412
rect 876 -1418 879 -1412
rect 883 -1418 886 -1412
rect 890 -1418 893 -1412
rect 897 -1418 900 -1412
rect 904 -1418 907 -1412
rect 911 -1418 914 -1412
rect 918 -1418 921 -1412
rect 925 -1418 931 -1412
rect 932 -1418 935 -1412
rect 939 -1418 942 -1412
rect 946 -1418 952 -1412
rect 953 -1418 956 -1412
rect 960 -1418 963 -1412
rect 967 -1418 973 -1412
rect 974 -1418 977 -1412
rect 981 -1418 984 -1412
rect 988 -1418 991 -1412
rect 995 -1418 998 -1412
rect 1002 -1418 1008 -1412
rect 1009 -1418 1012 -1412
rect 1016 -1418 1019 -1412
rect 1023 -1418 1026 -1412
rect 1030 -1418 1033 -1412
rect 1037 -1418 1043 -1412
rect 1044 -1418 1047 -1412
rect 1051 -1418 1054 -1412
rect 1072 -1418 1075 -1412
rect 22 -1499 28 -1493
rect 29 -1499 32 -1493
rect 36 -1499 39 -1493
rect 43 -1499 46 -1493
rect 50 -1499 56 -1493
rect 57 -1499 60 -1493
rect 64 -1499 67 -1493
rect 71 -1499 77 -1493
rect 78 -1499 81 -1493
rect 85 -1499 91 -1493
rect 92 -1499 95 -1493
rect 99 -1499 102 -1493
rect 106 -1499 109 -1493
rect 113 -1499 116 -1493
rect 120 -1499 126 -1493
rect 127 -1499 133 -1493
rect 134 -1499 137 -1493
rect 141 -1499 144 -1493
rect 148 -1499 151 -1493
rect 155 -1499 158 -1493
rect 162 -1499 165 -1493
rect 169 -1499 172 -1493
rect 176 -1499 182 -1493
rect 183 -1499 189 -1493
rect 190 -1499 193 -1493
rect 197 -1499 200 -1493
rect 204 -1499 207 -1493
rect 211 -1499 214 -1493
rect 218 -1499 224 -1493
rect 225 -1499 231 -1493
rect 232 -1499 235 -1493
rect 239 -1499 245 -1493
rect 246 -1499 249 -1493
rect 253 -1499 256 -1493
rect 260 -1499 263 -1493
rect 267 -1499 270 -1493
rect 274 -1499 277 -1493
rect 281 -1499 284 -1493
rect 288 -1499 294 -1493
rect 295 -1499 298 -1493
rect 302 -1499 308 -1493
rect 309 -1499 315 -1493
rect 316 -1499 322 -1493
rect 323 -1499 326 -1493
rect 330 -1499 333 -1493
rect 337 -1499 340 -1493
rect 344 -1499 347 -1493
rect 351 -1499 354 -1493
rect 358 -1499 361 -1493
rect 365 -1499 368 -1493
rect 372 -1499 375 -1493
rect 379 -1499 382 -1493
rect 386 -1499 389 -1493
rect 393 -1499 399 -1493
rect 400 -1499 403 -1493
rect 407 -1499 410 -1493
rect 414 -1499 420 -1493
rect 421 -1499 424 -1493
rect 428 -1499 431 -1493
rect 435 -1499 441 -1493
rect 442 -1499 445 -1493
rect 449 -1499 452 -1493
rect 456 -1499 459 -1493
rect 463 -1499 466 -1493
rect 470 -1499 473 -1493
rect 477 -1499 480 -1493
rect 484 -1499 487 -1493
rect 491 -1499 494 -1493
rect 498 -1499 504 -1493
rect 505 -1499 508 -1493
rect 512 -1499 515 -1493
rect 519 -1499 522 -1493
rect 526 -1499 529 -1493
rect 533 -1499 539 -1493
rect 540 -1499 546 -1493
rect 547 -1499 550 -1493
rect 554 -1499 560 -1493
rect 561 -1499 567 -1493
rect 568 -1499 571 -1493
rect 575 -1499 581 -1493
rect 582 -1499 585 -1493
rect 589 -1499 592 -1493
rect 596 -1499 599 -1493
rect 603 -1499 606 -1493
rect 610 -1499 613 -1493
rect 617 -1499 623 -1493
rect 624 -1499 627 -1493
rect 631 -1499 637 -1493
rect 638 -1499 641 -1493
rect 645 -1499 648 -1493
rect 652 -1499 658 -1493
rect 659 -1499 662 -1493
rect 666 -1499 669 -1493
rect 673 -1499 676 -1493
rect 680 -1499 686 -1493
rect 687 -1499 690 -1493
rect 694 -1499 697 -1493
rect 701 -1499 704 -1493
rect 708 -1499 711 -1493
rect 715 -1499 718 -1493
rect 722 -1499 728 -1493
rect 729 -1499 732 -1493
rect 736 -1499 739 -1493
rect 743 -1499 746 -1493
rect 750 -1499 753 -1493
rect 757 -1499 760 -1493
rect 764 -1499 767 -1493
rect 771 -1499 774 -1493
rect 778 -1499 781 -1493
rect 785 -1499 788 -1493
rect 792 -1499 795 -1493
rect 799 -1499 805 -1493
rect 806 -1499 809 -1493
rect 813 -1499 816 -1493
rect 820 -1499 823 -1493
rect 827 -1499 830 -1493
rect 834 -1499 837 -1493
rect 841 -1499 844 -1493
rect 848 -1499 851 -1493
rect 855 -1499 858 -1493
rect 862 -1499 865 -1493
rect 869 -1499 872 -1493
rect 876 -1499 879 -1493
rect 883 -1499 886 -1493
rect 890 -1499 893 -1493
rect 897 -1499 900 -1493
rect 904 -1499 907 -1493
rect 911 -1499 914 -1493
rect 918 -1499 924 -1493
rect 925 -1499 928 -1493
rect 932 -1499 935 -1493
rect 939 -1499 945 -1493
rect 946 -1499 949 -1493
rect 953 -1499 956 -1493
rect 960 -1499 966 -1493
rect 967 -1499 973 -1493
rect 974 -1499 977 -1493
rect 981 -1499 984 -1493
rect 988 -1499 991 -1493
rect 995 -1499 998 -1493
rect 1002 -1499 1005 -1493
rect 1037 -1499 1040 -1493
rect 1065 -1499 1071 -1493
rect 1 -1596 4 -1590
rect 8 -1596 11 -1590
rect 15 -1596 18 -1590
rect 22 -1596 25 -1590
rect 29 -1596 32 -1590
rect 36 -1596 39 -1590
rect 43 -1596 49 -1590
rect 50 -1596 53 -1590
rect 57 -1596 60 -1590
rect 64 -1596 67 -1590
rect 71 -1596 77 -1590
rect 78 -1596 84 -1590
rect 85 -1596 88 -1590
rect 92 -1596 95 -1590
rect 99 -1596 102 -1590
rect 106 -1596 109 -1590
rect 113 -1596 116 -1590
rect 120 -1596 126 -1590
rect 127 -1596 130 -1590
rect 134 -1596 137 -1590
rect 141 -1596 144 -1590
rect 148 -1596 151 -1590
rect 155 -1596 158 -1590
rect 162 -1596 165 -1590
rect 169 -1596 172 -1590
rect 176 -1596 179 -1590
rect 183 -1596 186 -1590
rect 190 -1596 196 -1590
rect 197 -1596 200 -1590
rect 204 -1596 207 -1590
rect 211 -1596 214 -1590
rect 218 -1596 224 -1590
rect 225 -1596 231 -1590
rect 232 -1596 238 -1590
rect 239 -1596 245 -1590
rect 246 -1596 252 -1590
rect 253 -1596 256 -1590
rect 260 -1596 263 -1590
rect 267 -1596 270 -1590
rect 274 -1596 277 -1590
rect 281 -1596 284 -1590
rect 288 -1596 291 -1590
rect 295 -1596 298 -1590
rect 302 -1596 305 -1590
rect 309 -1596 312 -1590
rect 316 -1596 319 -1590
rect 323 -1596 329 -1590
rect 330 -1596 333 -1590
rect 337 -1596 343 -1590
rect 344 -1596 347 -1590
rect 351 -1596 357 -1590
rect 358 -1596 364 -1590
rect 365 -1596 368 -1590
rect 372 -1596 378 -1590
rect 379 -1596 382 -1590
rect 386 -1596 389 -1590
rect 393 -1596 399 -1590
rect 400 -1596 406 -1590
rect 407 -1596 410 -1590
rect 414 -1596 420 -1590
rect 421 -1596 424 -1590
rect 428 -1596 431 -1590
rect 435 -1596 441 -1590
rect 442 -1596 445 -1590
rect 449 -1596 455 -1590
rect 456 -1596 462 -1590
rect 463 -1596 466 -1590
rect 470 -1596 476 -1590
rect 477 -1596 480 -1590
rect 484 -1596 487 -1590
rect 491 -1596 497 -1590
rect 498 -1596 501 -1590
rect 505 -1596 511 -1590
rect 512 -1596 518 -1590
rect 519 -1596 522 -1590
rect 526 -1596 529 -1590
rect 533 -1596 539 -1590
rect 540 -1596 546 -1590
rect 547 -1596 550 -1590
rect 554 -1596 557 -1590
rect 561 -1596 564 -1590
rect 568 -1596 571 -1590
rect 575 -1596 578 -1590
rect 582 -1596 585 -1590
rect 589 -1596 592 -1590
rect 596 -1596 599 -1590
rect 603 -1596 606 -1590
rect 610 -1596 613 -1590
rect 617 -1596 620 -1590
rect 624 -1596 627 -1590
rect 631 -1596 634 -1590
rect 638 -1596 641 -1590
rect 645 -1596 648 -1590
rect 652 -1596 655 -1590
rect 659 -1596 665 -1590
rect 666 -1596 669 -1590
rect 673 -1596 676 -1590
rect 680 -1596 686 -1590
rect 687 -1596 690 -1590
rect 694 -1596 697 -1590
rect 701 -1596 704 -1590
rect 708 -1596 714 -1590
rect 715 -1596 718 -1590
rect 722 -1596 725 -1590
rect 729 -1596 735 -1590
rect 736 -1596 739 -1590
rect 743 -1596 746 -1590
rect 750 -1596 753 -1590
rect 757 -1596 763 -1590
rect 764 -1596 767 -1590
rect 771 -1596 774 -1590
rect 778 -1596 781 -1590
rect 785 -1596 788 -1590
rect 792 -1596 795 -1590
rect 799 -1596 805 -1590
rect 806 -1596 809 -1590
rect 813 -1596 816 -1590
rect 820 -1596 823 -1590
rect 827 -1596 830 -1590
rect 834 -1596 837 -1590
rect 841 -1596 844 -1590
rect 848 -1596 851 -1590
rect 855 -1596 858 -1590
rect 862 -1596 865 -1590
rect 869 -1596 872 -1590
rect 876 -1596 879 -1590
rect 883 -1596 886 -1590
rect 890 -1596 893 -1590
rect 897 -1596 900 -1590
rect 904 -1596 907 -1590
rect 911 -1596 914 -1590
rect 918 -1596 921 -1590
rect 925 -1596 928 -1590
rect 932 -1596 935 -1590
rect 939 -1596 942 -1590
rect 946 -1596 949 -1590
rect 953 -1596 956 -1590
rect 960 -1596 963 -1590
rect 967 -1596 970 -1590
rect 974 -1596 977 -1590
rect 981 -1596 984 -1590
rect 988 -1596 991 -1590
rect 995 -1596 998 -1590
rect 1002 -1596 1005 -1590
rect 1009 -1596 1012 -1590
rect 1016 -1596 1019 -1590
rect 1023 -1596 1026 -1590
rect 1030 -1596 1033 -1590
rect 1037 -1596 1040 -1590
rect 1044 -1596 1047 -1590
rect 1051 -1596 1054 -1590
rect 1058 -1596 1061 -1590
rect 1065 -1596 1068 -1590
rect 1072 -1596 1075 -1590
rect 1079 -1596 1082 -1590
rect 1086 -1596 1089 -1590
rect 1093 -1596 1096 -1590
rect 1100 -1596 1103 -1590
rect 1107 -1596 1113 -1590
rect 1 -1683 4 -1677
rect 8 -1683 11 -1677
rect 15 -1683 18 -1677
rect 22 -1683 25 -1677
rect 29 -1683 32 -1677
rect 36 -1683 39 -1677
rect 43 -1683 46 -1677
rect 50 -1683 53 -1677
rect 57 -1683 63 -1677
rect 64 -1683 67 -1677
rect 71 -1683 74 -1677
rect 78 -1683 84 -1677
rect 85 -1683 88 -1677
rect 92 -1683 98 -1677
rect 99 -1683 102 -1677
rect 106 -1683 109 -1677
rect 113 -1683 116 -1677
rect 120 -1683 123 -1677
rect 127 -1683 130 -1677
rect 134 -1683 140 -1677
rect 141 -1683 144 -1677
rect 148 -1683 154 -1677
rect 155 -1683 161 -1677
rect 162 -1683 165 -1677
rect 169 -1683 172 -1677
rect 176 -1683 179 -1677
rect 183 -1683 186 -1677
rect 190 -1683 196 -1677
rect 197 -1683 203 -1677
rect 204 -1683 207 -1677
rect 211 -1683 217 -1677
rect 218 -1683 224 -1677
rect 225 -1683 231 -1677
rect 232 -1683 238 -1677
rect 239 -1683 242 -1677
rect 246 -1683 249 -1677
rect 253 -1683 256 -1677
rect 260 -1683 263 -1677
rect 267 -1683 270 -1677
rect 274 -1683 277 -1677
rect 281 -1683 287 -1677
rect 288 -1683 294 -1677
rect 295 -1683 301 -1677
rect 302 -1683 305 -1677
rect 309 -1683 312 -1677
rect 316 -1683 319 -1677
rect 323 -1683 326 -1677
rect 330 -1683 333 -1677
rect 337 -1683 340 -1677
rect 344 -1683 350 -1677
rect 351 -1683 354 -1677
rect 358 -1683 361 -1677
rect 365 -1683 371 -1677
rect 372 -1683 375 -1677
rect 379 -1683 385 -1677
rect 386 -1683 392 -1677
rect 393 -1683 396 -1677
rect 400 -1683 403 -1677
rect 407 -1683 410 -1677
rect 414 -1683 417 -1677
rect 421 -1683 424 -1677
rect 428 -1683 431 -1677
rect 435 -1683 438 -1677
rect 442 -1683 445 -1677
rect 449 -1683 455 -1677
rect 456 -1683 459 -1677
rect 463 -1683 469 -1677
rect 470 -1683 476 -1677
rect 477 -1683 483 -1677
rect 484 -1683 490 -1677
rect 491 -1683 497 -1677
rect 498 -1683 501 -1677
rect 505 -1683 508 -1677
rect 512 -1683 515 -1677
rect 519 -1683 522 -1677
rect 526 -1683 529 -1677
rect 533 -1683 539 -1677
rect 540 -1683 543 -1677
rect 547 -1683 553 -1677
rect 554 -1683 560 -1677
rect 561 -1683 567 -1677
rect 568 -1683 571 -1677
rect 575 -1683 578 -1677
rect 582 -1683 585 -1677
rect 589 -1683 592 -1677
rect 596 -1683 599 -1677
rect 603 -1683 606 -1677
rect 610 -1683 613 -1677
rect 617 -1683 620 -1677
rect 624 -1683 627 -1677
rect 631 -1683 634 -1677
rect 638 -1683 641 -1677
rect 645 -1683 648 -1677
rect 652 -1683 655 -1677
rect 659 -1683 662 -1677
rect 666 -1683 669 -1677
rect 673 -1683 676 -1677
rect 680 -1683 683 -1677
rect 687 -1683 690 -1677
rect 694 -1683 697 -1677
rect 701 -1683 704 -1677
rect 708 -1683 711 -1677
rect 715 -1683 718 -1677
rect 722 -1683 725 -1677
rect 729 -1683 735 -1677
rect 736 -1683 739 -1677
rect 743 -1683 746 -1677
rect 750 -1683 753 -1677
rect 757 -1683 760 -1677
rect 764 -1683 767 -1677
rect 771 -1683 774 -1677
rect 778 -1683 781 -1677
rect 785 -1683 788 -1677
rect 792 -1683 795 -1677
rect 799 -1683 802 -1677
rect 806 -1683 809 -1677
rect 813 -1683 816 -1677
rect 820 -1683 826 -1677
rect 827 -1683 830 -1677
rect 834 -1683 837 -1677
rect 841 -1683 844 -1677
rect 848 -1683 851 -1677
rect 855 -1683 858 -1677
rect 862 -1683 865 -1677
rect 869 -1683 872 -1677
rect 876 -1683 879 -1677
rect 883 -1683 889 -1677
rect 890 -1683 896 -1677
rect 897 -1683 900 -1677
rect 904 -1683 907 -1677
rect 911 -1683 917 -1677
rect 918 -1683 921 -1677
rect 925 -1683 928 -1677
rect 932 -1683 935 -1677
rect 939 -1683 942 -1677
rect 946 -1683 949 -1677
rect 953 -1683 956 -1677
rect 960 -1683 963 -1677
rect 974 -1683 977 -1677
rect 981 -1683 984 -1677
rect 1002 -1683 1005 -1677
rect 1023 -1683 1029 -1677
rect 1051 -1683 1054 -1677
rect 1 -1778 4 -1772
rect 8 -1778 14 -1772
rect 15 -1778 21 -1772
rect 22 -1778 25 -1772
rect 29 -1778 32 -1772
rect 36 -1778 39 -1772
rect 43 -1778 46 -1772
rect 50 -1778 56 -1772
rect 57 -1778 63 -1772
rect 64 -1778 67 -1772
rect 71 -1778 74 -1772
rect 78 -1778 81 -1772
rect 85 -1778 88 -1772
rect 92 -1778 95 -1772
rect 99 -1778 105 -1772
rect 106 -1778 112 -1772
rect 113 -1778 116 -1772
rect 120 -1778 123 -1772
rect 127 -1778 130 -1772
rect 134 -1778 137 -1772
rect 141 -1778 144 -1772
rect 148 -1778 154 -1772
rect 155 -1778 158 -1772
rect 162 -1778 168 -1772
rect 169 -1778 172 -1772
rect 176 -1778 182 -1772
rect 183 -1778 189 -1772
rect 190 -1778 193 -1772
rect 197 -1778 200 -1772
rect 204 -1778 207 -1772
rect 211 -1778 217 -1772
rect 218 -1778 224 -1772
rect 225 -1778 228 -1772
rect 232 -1778 235 -1772
rect 239 -1778 245 -1772
rect 246 -1778 249 -1772
rect 253 -1778 256 -1772
rect 260 -1778 263 -1772
rect 267 -1778 270 -1772
rect 274 -1778 277 -1772
rect 281 -1778 284 -1772
rect 288 -1778 291 -1772
rect 295 -1778 298 -1772
rect 302 -1778 305 -1772
rect 309 -1778 315 -1772
rect 316 -1778 319 -1772
rect 323 -1778 329 -1772
rect 330 -1778 333 -1772
rect 337 -1778 340 -1772
rect 344 -1778 347 -1772
rect 351 -1778 354 -1772
rect 358 -1778 361 -1772
rect 365 -1778 371 -1772
rect 372 -1778 378 -1772
rect 379 -1778 385 -1772
rect 386 -1778 389 -1772
rect 393 -1778 396 -1772
rect 400 -1778 406 -1772
rect 407 -1778 413 -1772
rect 414 -1778 417 -1772
rect 421 -1778 427 -1772
rect 428 -1778 431 -1772
rect 435 -1778 438 -1772
rect 442 -1778 445 -1772
rect 449 -1778 452 -1772
rect 456 -1778 459 -1772
rect 463 -1778 469 -1772
rect 470 -1778 473 -1772
rect 477 -1778 483 -1772
rect 484 -1778 487 -1772
rect 491 -1778 494 -1772
rect 498 -1778 501 -1772
rect 505 -1778 508 -1772
rect 512 -1778 518 -1772
rect 519 -1778 522 -1772
rect 526 -1778 529 -1772
rect 533 -1778 536 -1772
rect 540 -1778 546 -1772
rect 547 -1778 550 -1772
rect 554 -1778 557 -1772
rect 561 -1778 564 -1772
rect 568 -1778 571 -1772
rect 575 -1778 578 -1772
rect 582 -1778 585 -1772
rect 589 -1778 595 -1772
rect 596 -1778 599 -1772
rect 603 -1778 606 -1772
rect 610 -1778 616 -1772
rect 617 -1778 623 -1772
rect 624 -1778 627 -1772
rect 631 -1778 637 -1772
rect 638 -1778 641 -1772
rect 645 -1778 651 -1772
rect 652 -1778 658 -1772
rect 659 -1778 662 -1772
rect 666 -1778 669 -1772
rect 673 -1778 679 -1772
rect 680 -1778 683 -1772
rect 687 -1778 690 -1772
rect 694 -1778 697 -1772
rect 701 -1778 704 -1772
rect 708 -1778 711 -1772
rect 715 -1778 718 -1772
rect 722 -1778 725 -1772
rect 729 -1778 732 -1772
rect 736 -1778 739 -1772
rect 743 -1778 746 -1772
rect 750 -1778 753 -1772
rect 757 -1778 760 -1772
rect 764 -1778 767 -1772
rect 771 -1778 774 -1772
rect 778 -1778 781 -1772
rect 785 -1778 788 -1772
rect 792 -1778 795 -1772
rect 799 -1778 805 -1772
rect 806 -1778 809 -1772
rect 813 -1778 816 -1772
rect 820 -1778 823 -1772
rect 827 -1778 830 -1772
rect 834 -1778 837 -1772
rect 841 -1778 844 -1772
rect 848 -1778 851 -1772
rect 855 -1778 858 -1772
rect 862 -1778 865 -1772
rect 869 -1778 872 -1772
rect 876 -1778 879 -1772
rect 883 -1778 886 -1772
rect 890 -1778 893 -1772
rect 897 -1778 900 -1772
rect 904 -1778 907 -1772
rect 911 -1778 914 -1772
rect 918 -1778 921 -1772
rect 925 -1778 928 -1772
rect 932 -1778 935 -1772
rect 939 -1778 942 -1772
rect 946 -1778 949 -1772
rect 953 -1778 956 -1772
rect 960 -1778 963 -1772
rect 967 -1778 970 -1772
rect 974 -1778 977 -1772
rect 981 -1778 984 -1772
rect 988 -1778 991 -1772
rect 995 -1778 1001 -1772
rect 1002 -1778 1008 -1772
rect 1009 -1778 1012 -1772
rect 1016 -1778 1019 -1772
rect 1023 -1778 1026 -1772
rect 50 -1869 53 -1863
rect 57 -1869 60 -1863
rect 64 -1869 67 -1863
rect 71 -1869 74 -1863
rect 78 -1869 81 -1863
rect 85 -1869 88 -1863
rect 92 -1869 95 -1863
rect 99 -1869 102 -1863
rect 106 -1869 109 -1863
rect 113 -1869 116 -1863
rect 120 -1869 123 -1863
rect 127 -1869 133 -1863
rect 134 -1869 137 -1863
rect 141 -1869 144 -1863
rect 148 -1869 151 -1863
rect 155 -1869 158 -1863
rect 162 -1869 168 -1863
rect 169 -1869 172 -1863
rect 176 -1869 179 -1863
rect 183 -1869 186 -1863
rect 190 -1869 196 -1863
rect 197 -1869 203 -1863
rect 204 -1869 210 -1863
rect 211 -1869 217 -1863
rect 218 -1869 224 -1863
rect 225 -1869 231 -1863
rect 232 -1869 235 -1863
rect 239 -1869 245 -1863
rect 246 -1869 249 -1863
rect 253 -1869 256 -1863
rect 260 -1869 263 -1863
rect 267 -1869 270 -1863
rect 274 -1869 277 -1863
rect 281 -1869 284 -1863
rect 288 -1869 291 -1863
rect 295 -1869 298 -1863
rect 302 -1869 305 -1863
rect 309 -1869 312 -1863
rect 316 -1869 319 -1863
rect 323 -1869 326 -1863
rect 330 -1869 333 -1863
rect 337 -1869 340 -1863
rect 344 -1869 350 -1863
rect 351 -1869 354 -1863
rect 358 -1869 364 -1863
rect 365 -1869 371 -1863
rect 372 -1869 375 -1863
rect 379 -1869 382 -1863
rect 386 -1869 389 -1863
rect 393 -1869 396 -1863
rect 400 -1869 403 -1863
rect 407 -1869 413 -1863
rect 414 -1869 420 -1863
rect 421 -1869 427 -1863
rect 428 -1869 431 -1863
rect 435 -1869 438 -1863
rect 442 -1869 445 -1863
rect 449 -1869 452 -1863
rect 456 -1869 462 -1863
rect 463 -1869 466 -1863
rect 470 -1869 473 -1863
rect 477 -1869 480 -1863
rect 484 -1869 487 -1863
rect 491 -1869 494 -1863
rect 498 -1869 501 -1863
rect 505 -1869 511 -1863
rect 512 -1869 515 -1863
rect 519 -1869 525 -1863
rect 526 -1869 532 -1863
rect 533 -1869 536 -1863
rect 540 -1869 543 -1863
rect 547 -1869 553 -1863
rect 554 -1869 557 -1863
rect 561 -1869 567 -1863
rect 568 -1869 574 -1863
rect 575 -1869 578 -1863
rect 582 -1869 585 -1863
rect 589 -1869 592 -1863
rect 596 -1869 599 -1863
rect 603 -1869 606 -1863
rect 610 -1869 613 -1863
rect 617 -1869 620 -1863
rect 624 -1869 630 -1863
rect 631 -1869 637 -1863
rect 638 -1869 644 -1863
rect 645 -1869 648 -1863
rect 652 -1869 655 -1863
rect 659 -1869 665 -1863
rect 666 -1869 669 -1863
rect 673 -1869 676 -1863
rect 680 -1869 683 -1863
rect 687 -1869 690 -1863
rect 694 -1869 697 -1863
rect 701 -1869 707 -1863
rect 708 -1869 711 -1863
rect 715 -1869 718 -1863
rect 722 -1869 728 -1863
rect 729 -1869 732 -1863
rect 736 -1869 739 -1863
rect 743 -1869 746 -1863
rect 750 -1869 753 -1863
rect 757 -1869 760 -1863
rect 764 -1869 767 -1863
rect 771 -1869 774 -1863
rect 778 -1869 781 -1863
rect 785 -1869 788 -1863
rect 792 -1869 795 -1863
rect 799 -1869 802 -1863
rect 806 -1869 809 -1863
rect 813 -1869 819 -1863
rect 820 -1869 823 -1863
rect 827 -1869 830 -1863
rect 834 -1869 840 -1863
rect 841 -1869 847 -1863
rect 848 -1869 854 -1863
rect 855 -1869 858 -1863
rect 862 -1869 865 -1863
rect 869 -1869 872 -1863
rect 876 -1869 879 -1863
rect 897 -1869 900 -1863
rect 911 -1869 917 -1863
rect 946 -1869 952 -1863
rect 15 -1940 18 -1934
rect 22 -1940 25 -1934
rect 29 -1940 35 -1934
rect 36 -1940 42 -1934
rect 43 -1940 49 -1934
rect 50 -1940 53 -1934
rect 57 -1940 60 -1934
rect 64 -1940 67 -1934
rect 71 -1940 74 -1934
rect 78 -1940 81 -1934
rect 85 -1940 88 -1934
rect 92 -1940 95 -1934
rect 99 -1940 102 -1934
rect 106 -1940 109 -1934
rect 113 -1940 116 -1934
rect 120 -1940 126 -1934
rect 127 -1940 130 -1934
rect 134 -1940 137 -1934
rect 141 -1940 147 -1934
rect 148 -1940 151 -1934
rect 155 -1940 161 -1934
rect 162 -1940 165 -1934
rect 169 -1940 172 -1934
rect 176 -1940 182 -1934
rect 183 -1940 189 -1934
rect 190 -1940 196 -1934
rect 197 -1940 200 -1934
rect 204 -1940 207 -1934
rect 211 -1940 214 -1934
rect 218 -1940 224 -1934
rect 225 -1940 231 -1934
rect 232 -1940 238 -1934
rect 239 -1940 245 -1934
rect 246 -1940 249 -1934
rect 253 -1940 256 -1934
rect 260 -1940 263 -1934
rect 267 -1940 270 -1934
rect 274 -1940 277 -1934
rect 281 -1940 287 -1934
rect 288 -1940 291 -1934
rect 295 -1940 298 -1934
rect 302 -1940 305 -1934
rect 309 -1940 312 -1934
rect 316 -1940 322 -1934
rect 323 -1940 326 -1934
rect 330 -1940 336 -1934
rect 337 -1940 340 -1934
rect 344 -1940 347 -1934
rect 351 -1940 354 -1934
rect 358 -1940 361 -1934
rect 365 -1940 368 -1934
rect 372 -1940 375 -1934
rect 379 -1940 382 -1934
rect 386 -1940 389 -1934
rect 393 -1940 399 -1934
rect 400 -1940 403 -1934
rect 407 -1940 413 -1934
rect 414 -1940 420 -1934
rect 421 -1940 424 -1934
rect 428 -1940 431 -1934
rect 435 -1940 441 -1934
rect 442 -1940 445 -1934
rect 449 -1940 455 -1934
rect 456 -1940 462 -1934
rect 463 -1940 466 -1934
rect 470 -1940 476 -1934
rect 477 -1940 480 -1934
rect 484 -1940 487 -1934
rect 491 -1940 494 -1934
rect 498 -1940 504 -1934
rect 505 -1940 508 -1934
rect 512 -1940 515 -1934
rect 519 -1940 522 -1934
rect 526 -1940 529 -1934
rect 533 -1940 536 -1934
rect 540 -1940 543 -1934
rect 547 -1940 550 -1934
rect 554 -1940 557 -1934
rect 561 -1940 564 -1934
rect 568 -1940 571 -1934
rect 575 -1940 581 -1934
rect 582 -1940 585 -1934
rect 589 -1940 595 -1934
rect 596 -1940 599 -1934
rect 603 -1940 609 -1934
rect 610 -1940 613 -1934
rect 617 -1940 620 -1934
rect 624 -1940 627 -1934
rect 631 -1940 634 -1934
rect 638 -1940 641 -1934
rect 645 -1940 648 -1934
rect 652 -1940 655 -1934
rect 659 -1940 662 -1934
rect 666 -1940 669 -1934
rect 673 -1940 676 -1934
rect 680 -1940 686 -1934
rect 687 -1940 690 -1934
rect 694 -1940 697 -1934
rect 701 -1940 704 -1934
rect 708 -1940 711 -1934
rect 715 -1940 718 -1934
rect 722 -1940 725 -1934
rect 729 -1940 732 -1934
rect 736 -1940 739 -1934
rect 743 -1940 746 -1934
rect 750 -1940 753 -1934
rect 757 -1940 763 -1934
rect 764 -1940 767 -1934
rect 771 -1940 774 -1934
rect 778 -1940 784 -1934
rect 785 -1940 788 -1934
rect 792 -1940 795 -1934
rect 813 -1940 816 -1934
rect 820 -1940 823 -1934
rect 36 -1999 39 -1993
rect 43 -1999 46 -1993
rect 50 -1999 53 -1993
rect 57 -1999 60 -1993
rect 64 -1999 67 -1993
rect 71 -1999 74 -1993
rect 78 -1999 81 -1993
rect 85 -1999 88 -1993
rect 92 -1999 95 -1993
rect 99 -1999 102 -1993
rect 106 -1999 109 -1993
rect 113 -1999 116 -1993
rect 120 -1999 123 -1993
rect 127 -1999 133 -1993
rect 134 -1999 140 -1993
rect 141 -1999 144 -1993
rect 148 -1999 154 -1993
rect 155 -1999 161 -1993
rect 162 -1999 165 -1993
rect 169 -1999 172 -1993
rect 176 -1999 179 -1993
rect 183 -1999 186 -1993
rect 190 -1999 193 -1993
rect 197 -1999 203 -1993
rect 204 -1999 207 -1993
rect 211 -1999 214 -1993
rect 218 -1999 221 -1993
rect 225 -1999 231 -1993
rect 232 -1999 235 -1993
rect 239 -1999 245 -1993
rect 246 -1999 249 -1993
rect 253 -1999 256 -1993
rect 260 -1999 266 -1993
rect 267 -1999 273 -1993
rect 274 -1999 277 -1993
rect 281 -1999 284 -1993
rect 288 -1999 294 -1993
rect 295 -1999 298 -1993
rect 302 -1999 305 -1993
rect 309 -1999 315 -1993
rect 316 -1999 319 -1993
rect 323 -1999 326 -1993
rect 330 -1999 333 -1993
rect 337 -1999 340 -1993
rect 344 -1999 347 -1993
rect 351 -1999 354 -1993
rect 358 -1999 361 -1993
rect 365 -1999 371 -1993
rect 372 -1999 375 -1993
rect 379 -1999 385 -1993
rect 386 -1999 389 -1993
rect 393 -1999 396 -1993
rect 400 -1999 403 -1993
rect 407 -1999 410 -1993
rect 414 -1999 417 -1993
rect 421 -1999 424 -1993
rect 428 -1999 434 -1993
rect 435 -1999 441 -1993
rect 442 -1999 448 -1993
rect 449 -1999 452 -1993
rect 456 -1999 459 -1993
rect 463 -1999 466 -1993
rect 470 -1999 473 -1993
rect 477 -1999 480 -1993
rect 484 -1999 487 -1993
rect 491 -1999 497 -1993
rect 498 -1999 501 -1993
rect 505 -1999 508 -1993
rect 512 -1999 518 -1993
rect 519 -1999 522 -1993
rect 526 -1999 529 -1993
rect 533 -1999 536 -1993
rect 540 -1999 543 -1993
rect 547 -1999 550 -1993
rect 554 -1999 557 -1993
rect 561 -1999 564 -1993
rect 568 -1999 571 -1993
rect 575 -1999 578 -1993
rect 582 -1999 588 -1993
rect 589 -1999 595 -1993
rect 596 -1999 602 -1993
rect 603 -1999 606 -1993
rect 610 -1999 613 -1993
rect 617 -1999 620 -1993
rect 624 -1999 627 -1993
rect 631 -1999 634 -1993
rect 638 -1999 641 -1993
rect 645 -1999 648 -1993
rect 652 -1999 655 -1993
rect 659 -1999 665 -1993
rect 666 -1999 669 -1993
rect 673 -1999 679 -1993
rect 680 -1999 683 -1993
rect 687 -1999 693 -1993
rect 694 -1999 697 -1993
rect 701 -1999 704 -1993
rect 708 -1999 711 -1993
rect 715 -1999 718 -1993
rect 722 -1999 728 -1993
rect 729 -1999 732 -1993
rect 736 -1999 739 -1993
rect 743 -1999 749 -1993
rect 750 -1999 753 -1993
rect 757 -1999 760 -1993
rect 764 -1999 767 -1993
rect 771 -1999 774 -1993
rect 778 -1999 784 -1993
rect 785 -1999 788 -1993
rect 792 -1999 798 -1993
rect 799 -1999 802 -1993
rect 806 -1999 809 -1993
rect 813 -1999 816 -1993
rect 15 -2062 18 -2056
rect 22 -2062 25 -2056
rect 29 -2062 32 -2056
rect 36 -2062 39 -2056
rect 43 -2062 46 -2056
rect 50 -2062 53 -2056
rect 57 -2062 60 -2056
rect 64 -2062 67 -2056
rect 71 -2062 74 -2056
rect 78 -2062 81 -2056
rect 85 -2062 88 -2056
rect 92 -2062 95 -2056
rect 99 -2062 102 -2056
rect 106 -2062 109 -2056
rect 113 -2062 116 -2056
rect 120 -2062 126 -2056
rect 127 -2062 133 -2056
rect 134 -2062 137 -2056
rect 141 -2062 147 -2056
rect 148 -2062 151 -2056
rect 155 -2062 158 -2056
rect 162 -2062 168 -2056
rect 169 -2062 172 -2056
rect 176 -2062 182 -2056
rect 183 -2062 189 -2056
rect 190 -2062 193 -2056
rect 197 -2062 200 -2056
rect 204 -2062 207 -2056
rect 211 -2062 214 -2056
rect 218 -2062 221 -2056
rect 225 -2062 231 -2056
rect 232 -2062 238 -2056
rect 239 -2062 245 -2056
rect 246 -2062 249 -2056
rect 253 -2062 259 -2056
rect 260 -2062 263 -2056
rect 267 -2062 270 -2056
rect 274 -2062 277 -2056
rect 281 -2062 284 -2056
rect 288 -2062 291 -2056
rect 295 -2062 298 -2056
rect 302 -2062 305 -2056
rect 309 -2062 312 -2056
rect 316 -2062 319 -2056
rect 323 -2062 326 -2056
rect 330 -2062 333 -2056
rect 337 -2062 340 -2056
rect 344 -2062 350 -2056
rect 351 -2062 357 -2056
rect 358 -2062 361 -2056
rect 365 -2062 368 -2056
rect 372 -2062 375 -2056
rect 379 -2062 382 -2056
rect 386 -2062 389 -2056
rect 393 -2062 399 -2056
rect 400 -2062 406 -2056
rect 407 -2062 410 -2056
rect 414 -2062 420 -2056
rect 421 -2062 424 -2056
rect 428 -2062 434 -2056
rect 435 -2062 438 -2056
rect 442 -2062 445 -2056
rect 449 -2062 452 -2056
rect 456 -2062 462 -2056
rect 463 -2062 466 -2056
rect 470 -2062 476 -2056
rect 477 -2062 483 -2056
rect 484 -2062 490 -2056
rect 491 -2062 494 -2056
rect 498 -2062 501 -2056
rect 505 -2062 511 -2056
rect 512 -2062 518 -2056
rect 519 -2062 522 -2056
rect 526 -2062 529 -2056
rect 533 -2062 536 -2056
rect 540 -2062 543 -2056
rect 547 -2062 550 -2056
rect 554 -2062 557 -2056
rect 561 -2062 567 -2056
rect 568 -2062 574 -2056
rect 575 -2062 578 -2056
rect 582 -2062 585 -2056
rect 589 -2062 592 -2056
rect 596 -2062 599 -2056
rect 603 -2062 606 -2056
rect 610 -2062 613 -2056
rect 617 -2062 620 -2056
rect 624 -2062 627 -2056
rect 631 -2062 634 -2056
rect 638 -2062 641 -2056
rect 645 -2062 648 -2056
rect 652 -2062 658 -2056
rect 659 -2062 662 -2056
rect 666 -2062 672 -2056
rect 673 -2062 676 -2056
rect 680 -2062 683 -2056
rect 687 -2062 690 -2056
rect 694 -2062 697 -2056
rect 701 -2062 704 -2056
rect 708 -2062 711 -2056
rect 715 -2062 718 -2056
rect 722 -2062 728 -2056
rect 729 -2062 732 -2056
rect 736 -2062 739 -2056
rect 743 -2062 746 -2056
rect 750 -2062 753 -2056
rect 757 -2062 760 -2056
rect 764 -2062 767 -2056
rect 771 -2062 774 -2056
rect 778 -2062 781 -2056
rect 785 -2062 788 -2056
rect 15 -2127 18 -2121
rect 22 -2127 25 -2121
rect 29 -2127 32 -2121
rect 36 -2127 42 -2121
rect 43 -2127 46 -2121
rect 50 -2127 53 -2121
rect 57 -2127 60 -2121
rect 64 -2127 67 -2121
rect 71 -2127 74 -2121
rect 78 -2127 81 -2121
rect 85 -2127 88 -2121
rect 92 -2127 98 -2121
rect 99 -2127 105 -2121
rect 106 -2127 109 -2121
rect 113 -2127 116 -2121
rect 120 -2127 123 -2121
rect 127 -2127 133 -2121
rect 134 -2127 140 -2121
rect 141 -2127 144 -2121
rect 148 -2127 151 -2121
rect 155 -2127 161 -2121
rect 162 -2127 165 -2121
rect 169 -2127 175 -2121
rect 176 -2127 182 -2121
rect 183 -2127 189 -2121
rect 190 -2127 193 -2121
rect 197 -2127 203 -2121
rect 204 -2127 210 -2121
rect 211 -2127 214 -2121
rect 218 -2127 224 -2121
rect 225 -2127 231 -2121
rect 232 -2127 235 -2121
rect 239 -2127 242 -2121
rect 246 -2127 252 -2121
rect 253 -2127 256 -2121
rect 260 -2127 263 -2121
rect 267 -2127 270 -2121
rect 274 -2127 277 -2121
rect 281 -2127 284 -2121
rect 288 -2127 294 -2121
rect 295 -2127 298 -2121
rect 302 -2127 305 -2121
rect 309 -2127 312 -2121
rect 316 -2127 322 -2121
rect 323 -2127 326 -2121
rect 330 -2127 333 -2121
rect 337 -2127 340 -2121
rect 344 -2127 350 -2121
rect 351 -2127 354 -2121
rect 358 -2127 364 -2121
rect 365 -2127 368 -2121
rect 372 -2127 375 -2121
rect 379 -2127 385 -2121
rect 386 -2127 389 -2121
rect 393 -2127 396 -2121
rect 400 -2127 403 -2121
rect 407 -2127 413 -2121
rect 414 -2127 417 -2121
rect 421 -2127 424 -2121
rect 428 -2127 431 -2121
rect 435 -2127 441 -2121
rect 442 -2127 445 -2121
rect 449 -2127 452 -2121
rect 456 -2127 462 -2121
rect 463 -2127 469 -2121
rect 470 -2127 476 -2121
rect 477 -2127 480 -2121
rect 484 -2127 487 -2121
rect 491 -2127 494 -2121
rect 498 -2127 501 -2121
rect 505 -2127 511 -2121
rect 512 -2127 515 -2121
rect 519 -2127 522 -2121
rect 526 -2127 529 -2121
rect 533 -2127 536 -2121
rect 540 -2127 543 -2121
rect 547 -2127 550 -2121
rect 554 -2127 557 -2121
rect 561 -2127 564 -2121
rect 568 -2127 571 -2121
rect 575 -2127 578 -2121
rect 582 -2127 585 -2121
rect 589 -2127 595 -2121
rect 596 -2127 599 -2121
rect 603 -2127 606 -2121
rect 610 -2127 613 -2121
rect 617 -2127 620 -2121
rect 624 -2127 627 -2121
rect 631 -2127 634 -2121
rect 638 -2127 641 -2121
rect 645 -2127 648 -2121
rect 652 -2127 655 -2121
rect 659 -2127 662 -2121
rect 666 -2127 669 -2121
rect 673 -2127 676 -2121
rect 680 -2127 683 -2121
rect 687 -2127 690 -2121
rect 694 -2127 697 -2121
rect 701 -2127 704 -2121
rect 708 -2127 711 -2121
rect 715 -2127 718 -2121
rect 722 -2127 725 -2121
rect 729 -2127 735 -2121
rect 736 -2127 739 -2121
rect 85 -2178 88 -2172
rect 99 -2178 102 -2172
rect 106 -2178 109 -2172
rect 113 -2178 116 -2172
rect 120 -2178 123 -2172
rect 127 -2178 133 -2172
rect 134 -2178 140 -2172
rect 141 -2178 144 -2172
rect 148 -2178 154 -2172
rect 155 -2178 161 -2172
rect 162 -2178 165 -2172
rect 169 -2178 172 -2172
rect 176 -2178 179 -2172
rect 183 -2178 186 -2172
rect 190 -2178 193 -2172
rect 197 -2178 200 -2172
rect 204 -2178 207 -2172
rect 211 -2178 217 -2172
rect 218 -2178 224 -2172
rect 225 -2178 231 -2172
rect 232 -2178 235 -2172
rect 239 -2178 245 -2172
rect 246 -2178 249 -2172
rect 253 -2178 256 -2172
rect 260 -2178 263 -2172
rect 267 -2178 270 -2172
rect 274 -2178 277 -2172
rect 281 -2178 287 -2172
rect 288 -2178 291 -2172
rect 295 -2178 301 -2172
rect 302 -2178 305 -2172
rect 309 -2178 315 -2172
rect 316 -2178 319 -2172
rect 323 -2178 326 -2172
rect 330 -2178 336 -2172
rect 337 -2178 340 -2172
rect 344 -2178 347 -2172
rect 351 -2178 354 -2172
rect 358 -2178 361 -2172
rect 365 -2178 368 -2172
rect 372 -2178 375 -2172
rect 379 -2178 382 -2172
rect 386 -2178 392 -2172
rect 393 -2178 396 -2172
rect 400 -2178 403 -2172
rect 407 -2178 413 -2172
rect 414 -2178 417 -2172
rect 421 -2178 424 -2172
rect 428 -2178 434 -2172
rect 435 -2178 438 -2172
rect 442 -2178 445 -2172
rect 449 -2178 455 -2172
rect 456 -2178 462 -2172
rect 463 -2178 466 -2172
rect 470 -2178 473 -2172
rect 477 -2178 480 -2172
rect 484 -2178 487 -2172
rect 491 -2178 497 -2172
rect 498 -2178 501 -2172
rect 505 -2178 511 -2172
rect 512 -2178 515 -2172
rect 519 -2178 522 -2172
rect 526 -2178 529 -2172
rect 533 -2178 536 -2172
rect 540 -2178 543 -2172
rect 547 -2178 550 -2172
rect 554 -2178 560 -2172
rect 561 -2178 564 -2172
rect 568 -2178 574 -2172
rect 575 -2178 581 -2172
rect 582 -2178 588 -2172
rect 589 -2178 592 -2172
rect 596 -2178 599 -2172
rect 603 -2178 606 -2172
rect 610 -2178 613 -2172
rect 617 -2178 620 -2172
rect 624 -2178 627 -2172
rect 631 -2178 634 -2172
rect 638 -2178 641 -2172
rect 645 -2178 648 -2172
rect 652 -2178 655 -2172
rect 659 -2178 662 -2172
rect 666 -2178 672 -2172
rect 673 -2178 676 -2172
rect 680 -2178 686 -2172
rect 687 -2178 690 -2172
rect 694 -2178 700 -2172
rect 701 -2178 704 -2172
rect 708 -2178 711 -2172
rect 715 -2178 718 -2172
rect 722 -2178 725 -2172
rect 85 -2231 91 -2225
rect 106 -2231 109 -2225
rect 113 -2231 116 -2225
rect 120 -2231 126 -2225
rect 127 -2231 133 -2225
rect 134 -2231 140 -2225
rect 141 -2231 144 -2225
rect 148 -2231 151 -2225
rect 155 -2231 158 -2225
rect 162 -2231 168 -2225
rect 169 -2231 175 -2225
rect 176 -2231 182 -2225
rect 183 -2231 186 -2225
rect 190 -2231 193 -2225
rect 197 -2231 203 -2225
rect 204 -2231 210 -2225
rect 211 -2231 214 -2225
rect 218 -2231 221 -2225
rect 225 -2231 231 -2225
rect 232 -2231 235 -2225
rect 239 -2231 242 -2225
rect 246 -2231 249 -2225
rect 253 -2231 256 -2225
rect 260 -2231 263 -2225
rect 267 -2231 270 -2225
rect 274 -2231 277 -2225
rect 281 -2231 287 -2225
rect 288 -2231 291 -2225
rect 295 -2231 298 -2225
rect 302 -2231 308 -2225
rect 309 -2231 312 -2225
rect 316 -2231 319 -2225
rect 323 -2231 326 -2225
rect 330 -2231 333 -2225
rect 337 -2231 340 -2225
rect 344 -2231 347 -2225
rect 351 -2231 354 -2225
rect 358 -2231 364 -2225
rect 365 -2231 368 -2225
rect 372 -2231 378 -2225
rect 379 -2231 382 -2225
rect 386 -2231 392 -2225
rect 393 -2231 396 -2225
rect 400 -2231 403 -2225
rect 407 -2231 410 -2225
rect 414 -2231 417 -2225
rect 421 -2231 427 -2225
rect 428 -2231 431 -2225
rect 435 -2231 438 -2225
rect 442 -2231 448 -2225
rect 449 -2231 452 -2225
rect 456 -2231 459 -2225
rect 463 -2231 469 -2225
rect 470 -2231 473 -2225
rect 477 -2231 480 -2225
rect 484 -2231 487 -2225
rect 491 -2231 494 -2225
rect 498 -2231 501 -2225
rect 505 -2231 508 -2225
rect 512 -2231 515 -2225
rect 519 -2231 522 -2225
rect 526 -2231 529 -2225
rect 533 -2231 536 -2225
rect 540 -2231 543 -2225
rect 547 -2231 550 -2225
rect 554 -2231 557 -2225
rect 561 -2231 567 -2225
rect 568 -2231 571 -2225
rect 575 -2231 581 -2225
rect 582 -2231 585 -2225
rect 589 -2231 592 -2225
rect 596 -2231 599 -2225
rect 603 -2231 609 -2225
rect 610 -2231 616 -2225
rect 617 -2231 623 -2225
rect 624 -2231 630 -2225
rect 631 -2231 634 -2225
rect 638 -2231 641 -2225
rect 659 -2231 662 -2225
rect 113 -2268 116 -2262
rect 120 -2268 126 -2262
rect 127 -2268 133 -2262
rect 134 -2268 137 -2262
rect 141 -2268 147 -2262
rect 148 -2268 154 -2262
rect 155 -2268 158 -2262
rect 162 -2268 165 -2262
rect 169 -2268 172 -2262
rect 176 -2268 179 -2262
rect 183 -2268 186 -2262
rect 190 -2268 196 -2262
rect 197 -2268 200 -2262
rect 204 -2268 207 -2262
rect 211 -2268 217 -2262
rect 218 -2268 221 -2262
rect 225 -2268 228 -2262
rect 232 -2268 238 -2262
rect 239 -2268 245 -2262
rect 246 -2268 249 -2262
rect 253 -2268 256 -2262
rect 260 -2268 263 -2262
rect 267 -2268 270 -2262
rect 274 -2268 277 -2262
rect 281 -2268 287 -2262
rect 288 -2268 291 -2262
rect 295 -2268 298 -2262
rect 302 -2268 308 -2262
rect 309 -2268 315 -2262
rect 316 -2268 319 -2262
rect 323 -2268 329 -2262
rect 330 -2268 333 -2262
rect 337 -2268 340 -2262
rect 344 -2268 347 -2262
rect 351 -2268 354 -2262
rect 358 -2268 364 -2262
rect 365 -2268 368 -2262
rect 372 -2268 378 -2262
rect 379 -2268 382 -2262
rect 386 -2268 392 -2262
rect 393 -2268 399 -2262
rect 400 -2268 403 -2262
rect 407 -2268 413 -2262
rect 414 -2268 417 -2262
rect 421 -2268 424 -2262
rect 428 -2268 434 -2262
rect 435 -2268 438 -2262
rect 442 -2268 445 -2262
rect 449 -2268 452 -2262
rect 456 -2268 459 -2262
rect 463 -2268 466 -2262
rect 470 -2268 476 -2262
rect 477 -2268 480 -2262
rect 484 -2268 487 -2262
rect 491 -2268 494 -2262
rect 498 -2268 501 -2262
rect 505 -2268 508 -2262
rect 512 -2268 515 -2262
rect 519 -2268 522 -2262
rect 526 -2268 529 -2262
rect 533 -2268 536 -2262
rect 540 -2268 543 -2262
rect 547 -2268 550 -2262
rect 554 -2268 557 -2262
rect 561 -2268 567 -2262
rect 568 -2268 574 -2262
rect 575 -2268 578 -2262
rect 582 -2268 585 -2262
rect 638 -2268 641 -2262
rect 120 -2295 126 -2289
rect 176 -2295 179 -2289
rect 211 -2295 214 -2289
rect 218 -2295 224 -2289
rect 225 -2295 228 -2289
rect 232 -2295 235 -2289
rect 239 -2295 245 -2289
rect 246 -2295 252 -2289
rect 253 -2295 256 -2289
rect 267 -2295 270 -2289
rect 274 -2295 277 -2289
rect 281 -2295 284 -2289
rect 288 -2295 294 -2289
rect 295 -2295 298 -2289
rect 302 -2295 308 -2289
rect 309 -2295 312 -2289
rect 316 -2295 319 -2289
rect 323 -2295 329 -2289
rect 330 -2295 333 -2289
rect 337 -2295 343 -2289
rect 344 -2295 347 -2289
rect 365 -2295 368 -2289
rect 379 -2295 382 -2289
rect 400 -2295 406 -2289
rect 414 -2295 417 -2289
rect 421 -2295 424 -2289
rect 428 -2295 434 -2289
rect 435 -2295 441 -2289
rect 442 -2295 448 -2289
rect 449 -2295 452 -2289
rect 456 -2295 459 -2289
rect 463 -2295 466 -2289
rect 470 -2295 476 -2289
rect 477 -2295 483 -2289
rect 498 -2295 504 -2289
rect 505 -2295 508 -2289
rect 512 -2295 515 -2289
rect 519 -2295 522 -2289
rect 526 -2295 532 -2289
rect 533 -2295 539 -2289
rect 540 -2295 543 -2289
rect 547 -2295 553 -2289
rect 568 -2295 574 -2289
rect 575 -2295 578 -2289
rect 638 -2295 641 -2289
rect 169 -2312 175 -2306
rect 176 -2312 179 -2306
rect 211 -2312 217 -2306
rect 225 -2312 228 -2306
rect 232 -2312 235 -2306
rect 239 -2312 245 -2306
rect 246 -2312 249 -2306
rect 253 -2312 256 -2306
rect 260 -2312 266 -2306
rect 267 -2312 273 -2306
rect 274 -2312 280 -2306
rect 281 -2312 287 -2306
rect 288 -2312 294 -2306
rect 295 -2312 298 -2306
rect 302 -2312 308 -2306
rect 309 -2312 315 -2306
rect 316 -2312 319 -2306
rect 365 -2312 371 -2306
rect 379 -2312 382 -2306
rect 386 -2312 392 -2306
rect 400 -2312 406 -2306
rect 407 -2312 410 -2306
rect 505 -2312 511 -2306
rect 526 -2312 529 -2306
rect 533 -2312 539 -2306
rect 596 -2312 599 -2306
rect 603 -2312 609 -2306
rect 610 -2312 616 -2306
rect 638 -2312 644 -2306
rect 645 -2312 648 -2306
<< polysilicon >>
rect 177 -5 178 -3
rect 177 -11 178 -9
rect 184 -11 185 -9
rect 187 -11 188 -9
rect 191 -5 192 -3
rect 194 -11 195 -9
rect 198 -11 199 -9
rect 201 -11 202 -9
rect 205 -5 206 -3
rect 208 -11 209 -9
rect 212 -5 213 -3
rect 212 -11 213 -9
rect 257 -5 258 -3
rect 254 -11 255 -9
rect 271 -5 272 -3
rect 275 -5 276 -3
rect 275 -11 276 -9
rect 282 -5 283 -3
rect 282 -11 283 -9
rect 310 -5 311 -3
rect 310 -11 311 -9
rect 348 -5 349 -3
rect 348 -11 349 -9
rect 359 -5 360 -3
rect 366 -5 367 -3
rect 366 -11 367 -9
rect 156 -28 157 -26
rect 198 -22 199 -20
rect 215 -22 216 -20
rect 212 -28 213 -26
rect 215 -28 216 -26
rect 219 -22 220 -20
rect 219 -28 220 -26
rect 233 -22 234 -20
rect 233 -28 234 -26
rect 240 -22 241 -20
rect 240 -28 241 -26
rect 250 -22 251 -20
rect 254 -22 255 -20
rect 254 -28 255 -26
rect 261 -22 262 -20
rect 261 -28 262 -26
rect 271 -28 272 -26
rect 282 -22 283 -20
rect 282 -28 283 -26
rect 296 -28 297 -26
rect 303 -22 304 -20
rect 303 -28 304 -26
rect 334 -28 335 -26
rect 341 -22 342 -20
rect 341 -28 342 -26
rect 366 -22 367 -20
rect 366 -28 367 -26
rect 373 -22 374 -20
rect 373 -28 374 -26
rect 383 -22 384 -20
rect 380 -28 381 -26
rect 387 -22 388 -20
rect 387 -28 388 -26
rect 394 -22 395 -20
rect 394 -28 395 -26
rect 100 -49 101 -47
rect 107 -49 108 -47
rect 156 -43 157 -41
rect 156 -49 157 -47
rect 166 -43 167 -41
rect 170 -49 171 -47
rect 177 -43 178 -41
rect 177 -49 178 -47
rect 187 -49 188 -47
rect 194 -43 195 -41
rect 198 -43 199 -41
rect 198 -49 199 -47
rect 205 -43 206 -41
rect 205 -49 206 -47
rect 212 -43 213 -41
rect 215 -49 216 -47
rect 219 -43 220 -41
rect 219 -49 220 -47
rect 226 -43 227 -41
rect 226 -49 227 -47
rect 233 -43 234 -41
rect 240 -43 241 -41
rect 240 -49 241 -47
rect 247 -43 248 -41
rect 247 -49 248 -47
rect 254 -43 255 -41
rect 261 -43 262 -41
rect 261 -49 262 -47
rect 268 -43 269 -41
rect 268 -49 269 -47
rect 275 -43 276 -41
rect 275 -49 276 -47
rect 282 -43 283 -41
rect 282 -49 283 -47
rect 289 -43 290 -41
rect 289 -49 290 -47
rect 296 -43 297 -41
rect 299 -43 300 -41
rect 303 -49 304 -47
rect 310 -43 311 -41
rect 310 -49 311 -47
rect 317 -43 318 -41
rect 317 -49 318 -47
rect 324 -43 325 -41
rect 324 -49 325 -47
rect 331 -43 332 -41
rect 331 -49 332 -47
rect 338 -43 339 -41
rect 338 -49 339 -47
rect 345 -43 346 -41
rect 345 -49 346 -47
rect 352 -43 353 -41
rect 352 -49 353 -47
rect 362 -49 363 -47
rect 366 -43 367 -41
rect 366 -49 367 -47
rect 373 -43 374 -41
rect 376 -49 377 -47
rect 380 -43 381 -41
rect 387 -43 388 -41
rect 387 -49 388 -47
rect 394 -43 395 -41
rect 394 -49 395 -47
rect 401 -49 402 -47
rect 411 -43 412 -41
rect 415 -43 416 -41
rect 415 -49 416 -47
rect 422 -43 423 -41
rect 422 -49 423 -47
rect 429 -43 430 -41
rect 429 -49 430 -47
rect 436 -49 437 -47
rect 443 -49 444 -47
rect 450 -43 451 -41
rect 450 -49 451 -47
rect 86 -80 87 -78
rect 86 -86 87 -84
rect 93 -80 94 -78
rect 93 -86 94 -84
rect 100 -80 101 -78
rect 100 -86 101 -84
rect 107 -80 108 -78
rect 114 -86 115 -84
rect 117 -86 118 -84
rect 121 -80 122 -78
rect 124 -86 125 -84
rect 128 -80 129 -78
rect 128 -86 129 -84
rect 135 -80 136 -78
rect 135 -86 136 -84
rect 142 -80 143 -78
rect 142 -86 143 -84
rect 149 -80 150 -78
rect 149 -86 150 -84
rect 156 -80 157 -78
rect 156 -86 157 -84
rect 163 -80 164 -78
rect 163 -86 164 -84
rect 170 -80 171 -78
rect 170 -86 171 -84
rect 177 -80 178 -78
rect 177 -86 178 -84
rect 184 -86 185 -84
rect 191 -80 192 -78
rect 191 -86 192 -84
rect 198 -80 199 -78
rect 205 -80 206 -78
rect 205 -86 206 -84
rect 215 -80 216 -78
rect 219 -80 220 -78
rect 222 -86 223 -84
rect 226 -80 227 -78
rect 226 -86 227 -84
rect 233 -80 234 -78
rect 233 -86 234 -84
rect 243 -80 244 -78
rect 243 -86 244 -84
rect 247 -80 248 -78
rect 247 -86 248 -84
rect 254 -86 255 -84
rect 261 -80 262 -78
rect 261 -86 262 -84
rect 268 -80 269 -78
rect 268 -86 269 -84
rect 275 -80 276 -78
rect 275 -86 276 -84
rect 282 -80 283 -78
rect 282 -86 283 -84
rect 289 -80 290 -78
rect 289 -86 290 -84
rect 296 -80 297 -78
rect 296 -86 297 -84
rect 303 -80 304 -78
rect 303 -86 304 -84
rect 310 -80 311 -78
rect 313 -86 314 -84
rect 317 -80 318 -78
rect 317 -86 318 -84
rect 324 -80 325 -78
rect 324 -86 325 -84
rect 331 -80 332 -78
rect 331 -86 332 -84
rect 338 -80 339 -78
rect 341 -80 342 -78
rect 348 -80 349 -78
rect 345 -86 346 -84
rect 348 -86 349 -84
rect 355 -80 356 -78
rect 355 -86 356 -84
rect 362 -80 363 -78
rect 362 -86 363 -84
rect 369 -80 370 -78
rect 366 -86 367 -84
rect 373 -80 374 -78
rect 373 -86 374 -84
rect 380 -80 381 -78
rect 380 -86 381 -84
rect 387 -80 388 -78
rect 387 -86 388 -84
rect 394 -80 395 -78
rect 394 -86 395 -84
rect 401 -80 402 -78
rect 401 -86 402 -84
rect 408 -80 409 -78
rect 408 -86 409 -84
rect 415 -80 416 -78
rect 415 -86 416 -84
rect 422 -80 423 -78
rect 422 -86 423 -84
rect 429 -80 430 -78
rect 429 -86 430 -84
rect 436 -80 437 -78
rect 436 -86 437 -84
rect 443 -80 444 -78
rect 443 -86 444 -84
rect 450 -80 451 -78
rect 450 -86 451 -84
rect 457 -80 458 -78
rect 457 -86 458 -84
rect 464 -80 465 -78
rect 464 -86 465 -84
rect 471 -80 472 -78
rect 471 -86 472 -84
rect 478 -80 479 -78
rect 478 -86 479 -84
rect 485 -80 486 -78
rect 485 -86 486 -84
rect 495 -80 496 -78
rect 499 -80 500 -78
rect 499 -86 500 -84
rect 506 -86 507 -84
rect 562 -86 563 -84
rect 565 -86 566 -84
rect 579 -80 580 -78
rect 583 -80 584 -78
rect 583 -86 584 -84
rect 51 -141 52 -139
rect 58 -135 59 -133
rect 58 -141 59 -139
rect 65 -135 66 -133
rect 65 -141 66 -139
rect 72 -135 73 -133
rect 72 -141 73 -139
rect 79 -135 80 -133
rect 79 -141 80 -139
rect 86 -135 87 -133
rect 86 -141 87 -139
rect 93 -135 94 -133
rect 93 -141 94 -139
rect 100 -135 101 -133
rect 107 -135 108 -133
rect 107 -141 108 -139
rect 114 -135 115 -133
rect 114 -141 115 -139
rect 121 -135 122 -133
rect 121 -141 122 -139
rect 128 -135 129 -133
rect 128 -141 129 -139
rect 135 -135 136 -133
rect 135 -141 136 -139
rect 142 -135 143 -133
rect 142 -141 143 -139
rect 149 -135 150 -133
rect 149 -141 150 -139
rect 156 -135 157 -133
rect 156 -141 157 -139
rect 163 -135 164 -133
rect 163 -141 164 -139
rect 170 -135 171 -133
rect 170 -141 171 -139
rect 177 -135 178 -133
rect 180 -135 181 -133
rect 177 -141 178 -139
rect 180 -141 181 -139
rect 184 -135 185 -133
rect 187 -135 188 -133
rect 187 -141 188 -139
rect 191 -141 192 -139
rect 194 -141 195 -139
rect 198 -135 199 -133
rect 198 -141 199 -139
rect 205 -135 206 -133
rect 205 -141 206 -139
rect 212 -141 213 -139
rect 215 -141 216 -139
rect 222 -135 223 -133
rect 222 -141 223 -139
rect 226 -135 227 -133
rect 226 -141 227 -139
rect 229 -141 230 -139
rect 233 -135 234 -133
rect 233 -141 234 -139
rect 240 -135 241 -133
rect 243 -135 244 -133
rect 243 -141 244 -139
rect 247 -135 248 -133
rect 247 -141 248 -139
rect 254 -135 255 -133
rect 254 -141 255 -139
rect 261 -135 262 -133
rect 261 -141 262 -139
rect 268 -135 269 -133
rect 268 -141 269 -139
rect 275 -135 276 -133
rect 275 -141 276 -139
rect 282 -135 283 -133
rect 285 -135 286 -133
rect 282 -141 283 -139
rect 285 -141 286 -139
rect 289 -135 290 -133
rect 289 -141 290 -139
rect 296 -135 297 -133
rect 299 -135 300 -133
rect 296 -141 297 -139
rect 299 -141 300 -139
rect 303 -135 304 -133
rect 306 -135 307 -133
rect 310 -135 311 -133
rect 310 -141 311 -139
rect 317 -135 318 -133
rect 317 -141 318 -139
rect 324 -135 325 -133
rect 324 -141 325 -139
rect 331 -135 332 -133
rect 334 -135 335 -133
rect 331 -141 332 -139
rect 338 -141 339 -139
rect 341 -141 342 -139
rect 345 -135 346 -133
rect 345 -141 346 -139
rect 352 -135 353 -133
rect 352 -141 353 -139
rect 355 -141 356 -139
rect 359 -135 360 -133
rect 362 -135 363 -133
rect 359 -141 360 -139
rect 362 -141 363 -139
rect 366 -135 367 -133
rect 369 -135 370 -133
rect 366 -141 367 -139
rect 373 -135 374 -133
rect 376 -135 377 -133
rect 376 -141 377 -139
rect 383 -135 384 -133
rect 380 -141 381 -139
rect 387 -135 388 -133
rect 387 -141 388 -139
rect 390 -141 391 -139
rect 394 -135 395 -133
rect 394 -141 395 -139
rect 401 -135 402 -133
rect 401 -141 402 -139
rect 408 -135 409 -133
rect 408 -141 409 -139
rect 415 -135 416 -133
rect 415 -141 416 -139
rect 422 -135 423 -133
rect 422 -141 423 -139
rect 429 -135 430 -133
rect 429 -141 430 -139
rect 436 -135 437 -133
rect 436 -141 437 -139
rect 443 -135 444 -133
rect 443 -141 444 -139
rect 450 -135 451 -133
rect 450 -141 451 -139
rect 457 -135 458 -133
rect 457 -141 458 -139
rect 464 -135 465 -133
rect 464 -141 465 -139
rect 471 -135 472 -133
rect 471 -141 472 -139
rect 478 -135 479 -133
rect 478 -141 479 -139
rect 485 -135 486 -133
rect 485 -141 486 -139
rect 492 -135 493 -133
rect 492 -141 493 -139
rect 499 -135 500 -133
rect 499 -141 500 -139
rect 506 -135 507 -133
rect 506 -141 507 -139
rect 513 -135 514 -133
rect 513 -141 514 -139
rect 520 -135 521 -133
rect 520 -141 521 -139
rect 527 -135 528 -133
rect 527 -141 528 -139
rect 534 -135 535 -133
rect 534 -141 535 -139
rect 541 -135 542 -133
rect 541 -141 542 -139
rect 551 -141 552 -139
rect 555 -135 556 -133
rect 555 -141 556 -139
rect 562 -135 563 -133
rect 562 -141 563 -139
rect 569 -135 570 -133
rect 569 -141 570 -139
rect 576 -135 577 -133
rect 576 -141 577 -139
rect 583 -135 584 -133
rect 583 -141 584 -139
rect 590 -135 591 -133
rect 590 -141 591 -139
rect 597 -135 598 -133
rect 597 -141 598 -139
rect 618 -135 619 -133
rect 618 -141 619 -139
rect 65 -194 66 -192
rect 65 -200 66 -198
rect 72 -200 73 -198
rect 79 -194 80 -192
rect 79 -200 80 -198
rect 86 -194 87 -192
rect 86 -200 87 -198
rect 93 -194 94 -192
rect 93 -200 94 -198
rect 100 -194 101 -192
rect 100 -200 101 -198
rect 107 -194 108 -192
rect 107 -200 108 -198
rect 114 -194 115 -192
rect 114 -200 115 -198
rect 121 -194 122 -192
rect 121 -200 122 -198
rect 128 -194 129 -192
rect 128 -200 129 -198
rect 135 -194 136 -192
rect 138 -194 139 -192
rect 138 -200 139 -198
rect 142 -194 143 -192
rect 142 -200 143 -198
rect 149 -194 150 -192
rect 149 -200 150 -198
rect 156 -194 157 -192
rect 156 -200 157 -198
rect 163 -194 164 -192
rect 163 -200 164 -198
rect 170 -194 171 -192
rect 173 -194 174 -192
rect 173 -200 174 -198
rect 177 -194 178 -192
rect 177 -200 178 -198
rect 187 -194 188 -192
rect 184 -200 185 -198
rect 187 -200 188 -198
rect 191 -200 192 -198
rect 198 -194 199 -192
rect 198 -200 199 -198
rect 205 -194 206 -192
rect 208 -194 209 -192
rect 205 -200 206 -198
rect 208 -200 209 -198
rect 212 -194 213 -192
rect 215 -194 216 -192
rect 219 -194 220 -192
rect 219 -200 220 -198
rect 226 -194 227 -192
rect 226 -200 227 -198
rect 233 -194 234 -192
rect 236 -194 237 -192
rect 233 -200 234 -198
rect 236 -200 237 -198
rect 240 -194 241 -192
rect 240 -200 241 -198
rect 247 -194 248 -192
rect 247 -200 248 -198
rect 254 -194 255 -192
rect 254 -200 255 -198
rect 261 -194 262 -192
rect 261 -200 262 -198
rect 268 -194 269 -192
rect 268 -200 269 -198
rect 275 -194 276 -192
rect 275 -200 276 -198
rect 282 -194 283 -192
rect 282 -200 283 -198
rect 289 -194 290 -192
rect 289 -200 290 -198
rect 296 -194 297 -192
rect 296 -200 297 -198
rect 299 -200 300 -198
rect 306 -194 307 -192
rect 303 -200 304 -198
rect 310 -194 311 -192
rect 310 -200 311 -198
rect 317 -194 318 -192
rect 320 -194 321 -192
rect 317 -200 318 -198
rect 320 -200 321 -198
rect 324 -194 325 -192
rect 324 -200 325 -198
rect 331 -194 332 -192
rect 331 -200 332 -198
rect 338 -194 339 -192
rect 338 -200 339 -198
rect 345 -194 346 -192
rect 345 -200 346 -198
rect 352 -194 353 -192
rect 355 -194 356 -192
rect 355 -200 356 -198
rect 359 -194 360 -192
rect 362 -194 363 -192
rect 366 -194 367 -192
rect 366 -200 367 -198
rect 373 -194 374 -192
rect 376 -194 377 -192
rect 373 -200 374 -198
rect 376 -200 377 -198
rect 380 -194 381 -192
rect 380 -200 381 -198
rect 387 -194 388 -192
rect 387 -200 388 -198
rect 394 -200 395 -198
rect 397 -200 398 -198
rect 404 -194 405 -192
rect 404 -200 405 -198
rect 408 -194 409 -192
rect 408 -200 409 -198
rect 415 -194 416 -192
rect 415 -200 416 -198
rect 422 -194 423 -192
rect 422 -200 423 -198
rect 429 -194 430 -192
rect 429 -200 430 -198
rect 439 -194 440 -192
rect 439 -200 440 -198
rect 443 -194 444 -192
rect 443 -200 444 -198
rect 450 -194 451 -192
rect 450 -200 451 -198
rect 457 -194 458 -192
rect 460 -200 461 -198
rect 464 -194 465 -192
rect 464 -200 465 -198
rect 471 -194 472 -192
rect 471 -200 472 -198
rect 478 -194 479 -192
rect 478 -200 479 -198
rect 485 -194 486 -192
rect 485 -200 486 -198
rect 492 -194 493 -192
rect 492 -200 493 -198
rect 499 -194 500 -192
rect 499 -200 500 -198
rect 506 -200 507 -198
rect 509 -200 510 -198
rect 513 -194 514 -192
rect 513 -200 514 -198
rect 520 -194 521 -192
rect 520 -200 521 -198
rect 527 -194 528 -192
rect 527 -200 528 -198
rect 534 -194 535 -192
rect 534 -200 535 -198
rect 544 -194 545 -192
rect 544 -200 545 -198
rect 548 -194 549 -192
rect 548 -200 549 -198
rect 555 -194 556 -192
rect 555 -200 556 -198
rect 562 -194 563 -192
rect 562 -200 563 -198
rect 572 -194 573 -192
rect 569 -200 570 -198
rect 576 -194 577 -192
rect 576 -200 577 -198
rect 583 -194 584 -192
rect 583 -200 584 -198
rect 590 -194 591 -192
rect 590 -200 591 -198
rect 632 -194 633 -192
rect 632 -200 633 -198
rect 642 -194 643 -192
rect 646 -194 647 -192
rect 646 -200 647 -198
rect 16 -251 17 -249
rect 16 -257 17 -255
rect 23 -251 24 -249
rect 23 -257 24 -255
rect 30 -251 31 -249
rect 30 -257 31 -255
rect 37 -251 38 -249
rect 37 -257 38 -255
rect 44 -251 45 -249
rect 44 -257 45 -255
rect 51 -251 52 -249
rect 58 -251 59 -249
rect 58 -257 59 -255
rect 65 -251 66 -249
rect 65 -257 66 -255
rect 72 -251 73 -249
rect 72 -257 73 -255
rect 79 -251 80 -249
rect 79 -257 80 -255
rect 86 -251 87 -249
rect 86 -257 87 -255
rect 93 -251 94 -249
rect 93 -257 94 -255
rect 100 -251 101 -249
rect 100 -257 101 -255
rect 103 -257 104 -255
rect 107 -251 108 -249
rect 107 -257 108 -255
rect 114 -251 115 -249
rect 114 -257 115 -255
rect 121 -251 122 -249
rect 121 -257 122 -255
rect 128 -251 129 -249
rect 131 -251 132 -249
rect 138 -251 139 -249
rect 138 -257 139 -255
rect 142 -251 143 -249
rect 145 -251 146 -249
rect 149 -251 150 -249
rect 149 -257 150 -255
rect 156 -257 157 -255
rect 159 -257 160 -255
rect 163 -251 164 -249
rect 163 -257 164 -255
rect 170 -251 171 -249
rect 170 -257 171 -255
rect 177 -251 178 -249
rect 177 -257 178 -255
rect 184 -251 185 -249
rect 184 -257 185 -255
rect 191 -251 192 -249
rect 194 -251 195 -249
rect 194 -257 195 -255
rect 198 -251 199 -249
rect 198 -257 199 -255
rect 208 -251 209 -249
rect 205 -257 206 -255
rect 212 -251 213 -249
rect 215 -257 216 -255
rect 219 -251 220 -249
rect 222 -251 223 -249
rect 226 -251 227 -249
rect 229 -251 230 -249
rect 226 -257 227 -255
rect 229 -257 230 -255
rect 233 -251 234 -249
rect 233 -257 234 -255
rect 240 -251 241 -249
rect 240 -257 241 -255
rect 247 -251 248 -249
rect 247 -257 248 -255
rect 254 -251 255 -249
rect 254 -257 255 -255
rect 261 -251 262 -249
rect 261 -257 262 -255
rect 268 -251 269 -249
rect 268 -257 269 -255
rect 271 -257 272 -255
rect 275 -251 276 -249
rect 275 -257 276 -255
rect 282 -251 283 -249
rect 282 -257 283 -255
rect 289 -251 290 -249
rect 289 -257 290 -255
rect 296 -251 297 -249
rect 296 -257 297 -255
rect 303 -251 304 -249
rect 303 -257 304 -255
rect 310 -251 311 -249
rect 310 -257 311 -255
rect 317 -251 318 -249
rect 317 -257 318 -255
rect 324 -251 325 -249
rect 324 -257 325 -255
rect 331 -251 332 -249
rect 331 -257 332 -255
rect 338 -251 339 -249
rect 338 -257 339 -255
rect 341 -257 342 -255
rect 345 -251 346 -249
rect 345 -257 346 -255
rect 352 -251 353 -249
rect 352 -257 353 -255
rect 359 -251 360 -249
rect 359 -257 360 -255
rect 366 -251 367 -249
rect 366 -257 367 -255
rect 373 -251 374 -249
rect 373 -257 374 -255
rect 380 -251 381 -249
rect 380 -257 381 -255
rect 390 -251 391 -249
rect 387 -257 388 -255
rect 390 -257 391 -255
rect 394 -251 395 -249
rect 397 -251 398 -249
rect 397 -257 398 -255
rect 401 -251 402 -249
rect 401 -257 402 -255
rect 408 -251 409 -249
rect 411 -251 412 -249
rect 411 -257 412 -255
rect 415 -251 416 -249
rect 418 -251 419 -249
rect 422 -251 423 -249
rect 422 -257 423 -255
rect 429 -251 430 -249
rect 429 -257 430 -255
rect 436 -251 437 -249
rect 436 -257 437 -255
rect 443 -251 444 -249
rect 443 -257 444 -255
rect 450 -251 451 -249
rect 450 -257 451 -255
rect 457 -251 458 -249
rect 460 -257 461 -255
rect 464 -251 465 -249
rect 467 -251 468 -249
rect 471 -251 472 -249
rect 471 -257 472 -255
rect 478 -251 479 -249
rect 481 -257 482 -255
rect 485 -251 486 -249
rect 485 -257 486 -255
rect 492 -251 493 -249
rect 492 -257 493 -255
rect 499 -251 500 -249
rect 499 -257 500 -255
rect 509 -251 510 -249
rect 506 -257 507 -255
rect 513 -251 514 -249
rect 520 -251 521 -249
rect 520 -257 521 -255
rect 527 -251 528 -249
rect 527 -257 528 -255
rect 534 -251 535 -249
rect 534 -257 535 -255
rect 541 -251 542 -249
rect 541 -257 542 -255
rect 548 -251 549 -249
rect 548 -257 549 -255
rect 555 -251 556 -249
rect 555 -257 556 -255
rect 562 -251 563 -249
rect 562 -257 563 -255
rect 569 -251 570 -249
rect 572 -257 573 -255
rect 576 -251 577 -249
rect 576 -257 577 -255
rect 583 -251 584 -249
rect 583 -257 584 -255
rect 590 -251 591 -249
rect 590 -257 591 -255
rect 597 -251 598 -249
rect 597 -257 598 -255
rect 600 -257 601 -255
rect 604 -251 605 -249
rect 604 -257 605 -255
rect 611 -251 612 -249
rect 611 -257 612 -255
rect 618 -251 619 -249
rect 618 -257 619 -255
rect 625 -251 626 -249
rect 625 -257 626 -255
rect 632 -251 633 -249
rect 632 -257 633 -255
rect 639 -251 640 -249
rect 639 -257 640 -255
rect 646 -251 647 -249
rect 646 -257 647 -255
rect 653 -251 654 -249
rect 653 -257 654 -255
rect 660 -251 661 -249
rect 660 -257 661 -255
rect 667 -251 668 -249
rect 670 -251 671 -249
rect 667 -257 668 -255
rect 670 -257 671 -255
rect 674 -251 675 -249
rect 674 -257 675 -255
rect 681 -251 682 -249
rect 681 -257 682 -255
rect 688 -251 689 -249
rect 688 -257 689 -255
rect 695 -251 696 -249
rect 695 -257 696 -255
rect 751 -251 752 -249
rect 751 -257 752 -255
rect 859 -257 860 -255
rect 30 -304 31 -302
rect 30 -310 31 -308
rect 37 -304 38 -302
rect 37 -310 38 -308
rect 44 -310 45 -308
rect 51 -304 52 -302
rect 51 -310 52 -308
rect 58 -304 59 -302
rect 58 -310 59 -308
rect 68 -304 69 -302
rect 65 -310 66 -308
rect 72 -304 73 -302
rect 72 -310 73 -308
rect 79 -304 80 -302
rect 79 -310 80 -308
rect 86 -304 87 -302
rect 86 -310 87 -308
rect 93 -304 94 -302
rect 93 -310 94 -308
rect 100 -304 101 -302
rect 100 -310 101 -308
rect 107 -304 108 -302
rect 107 -310 108 -308
rect 117 -304 118 -302
rect 114 -310 115 -308
rect 121 -304 122 -302
rect 121 -310 122 -308
rect 128 -304 129 -302
rect 128 -310 129 -308
rect 135 -304 136 -302
rect 138 -310 139 -308
rect 142 -304 143 -302
rect 142 -310 143 -308
rect 149 -304 150 -302
rect 149 -310 150 -308
rect 156 -304 157 -302
rect 156 -310 157 -308
rect 163 -304 164 -302
rect 163 -310 164 -308
rect 170 -304 171 -302
rect 170 -310 171 -308
rect 177 -304 178 -302
rect 180 -304 181 -302
rect 177 -310 178 -308
rect 184 -304 185 -302
rect 184 -310 185 -308
rect 191 -304 192 -302
rect 191 -310 192 -308
rect 198 -304 199 -302
rect 205 -304 206 -302
rect 205 -310 206 -308
rect 215 -304 216 -302
rect 212 -310 213 -308
rect 215 -310 216 -308
rect 222 -304 223 -302
rect 219 -310 220 -308
rect 222 -310 223 -308
rect 226 -304 227 -302
rect 226 -310 227 -308
rect 236 -304 237 -302
rect 233 -310 234 -308
rect 236 -310 237 -308
rect 240 -304 241 -302
rect 243 -304 244 -302
rect 240 -310 241 -308
rect 247 -310 248 -308
rect 254 -304 255 -302
rect 254 -310 255 -308
rect 257 -310 258 -308
rect 261 -304 262 -302
rect 261 -310 262 -308
rect 268 -304 269 -302
rect 268 -310 269 -308
rect 275 -304 276 -302
rect 275 -310 276 -308
rect 282 -304 283 -302
rect 282 -310 283 -308
rect 289 -310 290 -308
rect 296 -304 297 -302
rect 299 -304 300 -302
rect 299 -310 300 -308
rect 303 -304 304 -302
rect 303 -310 304 -308
rect 310 -304 311 -302
rect 310 -310 311 -308
rect 317 -304 318 -302
rect 317 -310 318 -308
rect 324 -304 325 -302
rect 324 -310 325 -308
rect 331 -304 332 -302
rect 334 -304 335 -302
rect 331 -310 332 -308
rect 334 -310 335 -308
rect 338 -304 339 -302
rect 338 -310 339 -308
rect 341 -310 342 -308
rect 345 -304 346 -302
rect 345 -310 346 -308
rect 352 -304 353 -302
rect 352 -310 353 -308
rect 359 -304 360 -302
rect 359 -310 360 -308
rect 366 -304 367 -302
rect 366 -310 367 -308
rect 373 -304 374 -302
rect 380 -304 381 -302
rect 380 -310 381 -308
rect 387 -304 388 -302
rect 387 -310 388 -308
rect 394 -304 395 -302
rect 397 -304 398 -302
rect 394 -310 395 -308
rect 401 -304 402 -302
rect 404 -304 405 -302
rect 401 -310 402 -308
rect 408 -304 409 -302
rect 408 -310 409 -308
rect 415 -304 416 -302
rect 415 -310 416 -308
rect 422 -304 423 -302
rect 425 -304 426 -302
rect 429 -304 430 -302
rect 429 -310 430 -308
rect 439 -304 440 -302
rect 436 -310 437 -308
rect 439 -310 440 -308
rect 446 -304 447 -302
rect 450 -304 451 -302
rect 450 -310 451 -308
rect 453 -310 454 -308
rect 457 -304 458 -302
rect 457 -310 458 -308
rect 464 -304 465 -302
rect 464 -310 465 -308
rect 471 -304 472 -302
rect 471 -310 472 -308
rect 478 -304 479 -302
rect 478 -310 479 -308
rect 485 -304 486 -302
rect 485 -310 486 -308
rect 492 -304 493 -302
rect 492 -310 493 -308
rect 499 -304 500 -302
rect 499 -310 500 -308
rect 506 -304 507 -302
rect 506 -310 507 -308
rect 513 -310 514 -308
rect 520 -304 521 -302
rect 520 -310 521 -308
rect 527 -304 528 -302
rect 527 -310 528 -308
rect 534 -304 535 -302
rect 534 -310 535 -308
rect 541 -304 542 -302
rect 544 -304 545 -302
rect 544 -310 545 -308
rect 548 -304 549 -302
rect 548 -310 549 -308
rect 555 -304 556 -302
rect 555 -310 556 -308
rect 562 -304 563 -302
rect 565 -304 566 -302
rect 562 -310 563 -308
rect 569 -304 570 -302
rect 569 -310 570 -308
rect 576 -304 577 -302
rect 576 -310 577 -308
rect 583 -304 584 -302
rect 583 -310 584 -308
rect 590 -304 591 -302
rect 590 -310 591 -308
rect 597 -304 598 -302
rect 600 -304 601 -302
rect 597 -310 598 -308
rect 604 -304 605 -302
rect 604 -310 605 -308
rect 611 -304 612 -302
rect 611 -310 612 -308
rect 618 -304 619 -302
rect 618 -310 619 -308
rect 625 -304 626 -302
rect 625 -310 626 -308
rect 632 -304 633 -302
rect 632 -310 633 -308
rect 639 -304 640 -302
rect 639 -310 640 -308
rect 646 -304 647 -302
rect 646 -310 647 -308
rect 653 -304 654 -302
rect 653 -310 654 -308
rect 660 -304 661 -302
rect 660 -310 661 -308
rect 667 -304 668 -302
rect 667 -310 668 -308
rect 677 -310 678 -308
rect 681 -304 682 -302
rect 681 -310 682 -308
rect 688 -304 689 -302
rect 688 -310 689 -308
rect 695 -304 696 -302
rect 695 -310 696 -308
rect 702 -304 703 -302
rect 702 -310 703 -308
rect 709 -304 710 -302
rect 709 -310 710 -308
rect 716 -304 717 -302
rect 716 -310 717 -308
rect 723 -304 724 -302
rect 726 -310 727 -308
rect 730 -304 731 -302
rect 730 -310 731 -308
rect 737 -304 738 -302
rect 737 -310 738 -308
rect 744 -304 745 -302
rect 744 -310 745 -308
rect 751 -304 752 -302
rect 751 -310 752 -308
rect 828 -304 829 -302
rect 828 -310 829 -308
rect 856 -304 857 -302
rect 856 -310 857 -308
rect 2 -375 3 -373
rect 2 -381 3 -379
rect 9 -375 10 -373
rect 9 -381 10 -379
rect 16 -375 17 -373
rect 16 -381 17 -379
rect 23 -375 24 -373
rect 23 -381 24 -379
rect 30 -375 31 -373
rect 30 -381 31 -379
rect 37 -375 38 -373
rect 37 -381 38 -379
rect 44 -375 45 -373
rect 44 -381 45 -379
rect 51 -375 52 -373
rect 51 -381 52 -379
rect 58 -375 59 -373
rect 58 -381 59 -379
rect 65 -375 66 -373
rect 65 -381 66 -379
rect 75 -375 76 -373
rect 72 -381 73 -379
rect 75 -381 76 -379
rect 79 -375 80 -373
rect 79 -381 80 -379
rect 86 -375 87 -373
rect 86 -381 87 -379
rect 93 -375 94 -373
rect 96 -375 97 -373
rect 96 -381 97 -379
rect 100 -375 101 -373
rect 100 -381 101 -379
rect 107 -375 108 -373
rect 107 -381 108 -379
rect 114 -375 115 -373
rect 114 -381 115 -379
rect 121 -375 122 -373
rect 121 -381 122 -379
rect 128 -375 129 -373
rect 131 -375 132 -373
rect 128 -381 129 -379
rect 131 -381 132 -379
rect 135 -375 136 -373
rect 135 -381 136 -379
rect 142 -375 143 -373
rect 145 -375 146 -373
rect 142 -381 143 -379
rect 145 -381 146 -379
rect 152 -375 153 -373
rect 149 -381 150 -379
rect 152 -381 153 -379
rect 156 -375 157 -373
rect 156 -381 157 -379
rect 163 -375 164 -373
rect 163 -381 164 -379
rect 170 -375 171 -373
rect 170 -381 171 -379
rect 177 -375 178 -373
rect 177 -381 178 -379
rect 184 -375 185 -373
rect 184 -381 185 -379
rect 191 -375 192 -373
rect 191 -381 192 -379
rect 198 -381 199 -379
rect 201 -381 202 -379
rect 205 -375 206 -373
rect 205 -381 206 -379
rect 215 -375 216 -373
rect 212 -381 213 -379
rect 219 -375 220 -373
rect 219 -381 220 -379
rect 226 -375 227 -373
rect 226 -381 227 -379
rect 233 -375 234 -373
rect 233 -381 234 -379
rect 240 -375 241 -373
rect 240 -381 241 -379
rect 247 -375 248 -373
rect 247 -381 248 -379
rect 254 -375 255 -373
rect 254 -381 255 -379
rect 261 -375 262 -373
rect 261 -381 262 -379
rect 268 -375 269 -373
rect 268 -381 269 -379
rect 275 -375 276 -373
rect 278 -381 279 -379
rect 282 -375 283 -373
rect 282 -381 283 -379
rect 289 -375 290 -373
rect 289 -381 290 -379
rect 296 -375 297 -373
rect 296 -381 297 -379
rect 303 -375 304 -373
rect 303 -381 304 -379
rect 310 -375 311 -373
rect 310 -381 311 -379
rect 317 -375 318 -373
rect 317 -381 318 -379
rect 324 -375 325 -373
rect 327 -375 328 -373
rect 331 -375 332 -373
rect 334 -375 335 -373
rect 331 -381 332 -379
rect 334 -381 335 -379
rect 338 -375 339 -373
rect 338 -381 339 -379
rect 345 -375 346 -373
rect 345 -381 346 -379
rect 352 -375 353 -373
rect 352 -381 353 -379
rect 359 -375 360 -373
rect 362 -375 363 -373
rect 359 -381 360 -379
rect 362 -381 363 -379
rect 366 -375 367 -373
rect 369 -375 370 -373
rect 366 -381 367 -379
rect 369 -381 370 -379
rect 373 -375 374 -373
rect 373 -381 374 -379
rect 376 -381 377 -379
rect 380 -375 381 -373
rect 380 -381 381 -379
rect 387 -375 388 -373
rect 387 -381 388 -379
rect 394 -375 395 -373
rect 394 -381 395 -379
rect 401 -375 402 -373
rect 404 -375 405 -373
rect 401 -381 402 -379
rect 404 -381 405 -379
rect 408 -375 409 -373
rect 408 -381 409 -379
rect 415 -375 416 -373
rect 415 -381 416 -379
rect 422 -375 423 -373
rect 425 -375 426 -373
rect 422 -381 423 -379
rect 425 -381 426 -379
rect 429 -375 430 -373
rect 432 -375 433 -373
rect 429 -381 430 -379
rect 432 -381 433 -379
rect 436 -375 437 -373
rect 436 -381 437 -379
rect 443 -375 444 -373
rect 443 -381 444 -379
rect 450 -375 451 -373
rect 453 -375 454 -373
rect 450 -381 451 -379
rect 457 -375 458 -373
rect 457 -381 458 -379
rect 464 -375 465 -373
rect 464 -381 465 -379
rect 471 -375 472 -373
rect 474 -375 475 -373
rect 471 -381 472 -379
rect 478 -375 479 -373
rect 478 -381 479 -379
rect 485 -375 486 -373
rect 485 -381 486 -379
rect 495 -375 496 -373
rect 495 -381 496 -379
rect 499 -375 500 -373
rect 499 -381 500 -379
rect 506 -381 507 -379
rect 509 -381 510 -379
rect 513 -375 514 -373
rect 516 -375 517 -373
rect 513 -381 514 -379
rect 516 -381 517 -379
rect 520 -375 521 -373
rect 520 -381 521 -379
rect 527 -375 528 -373
rect 527 -381 528 -379
rect 534 -375 535 -373
rect 534 -381 535 -379
rect 541 -375 542 -373
rect 541 -381 542 -379
rect 548 -375 549 -373
rect 548 -381 549 -379
rect 555 -375 556 -373
rect 555 -381 556 -379
rect 562 -375 563 -373
rect 562 -381 563 -379
rect 569 -375 570 -373
rect 569 -381 570 -379
rect 576 -375 577 -373
rect 576 -381 577 -379
rect 583 -375 584 -373
rect 586 -375 587 -373
rect 590 -375 591 -373
rect 590 -381 591 -379
rect 597 -375 598 -373
rect 597 -381 598 -379
rect 604 -375 605 -373
rect 604 -381 605 -379
rect 611 -375 612 -373
rect 611 -381 612 -379
rect 618 -375 619 -373
rect 618 -381 619 -379
rect 625 -375 626 -373
rect 625 -381 626 -379
rect 632 -375 633 -373
rect 632 -381 633 -379
rect 639 -375 640 -373
rect 639 -381 640 -379
rect 646 -375 647 -373
rect 646 -381 647 -379
rect 653 -375 654 -373
rect 653 -381 654 -379
rect 660 -375 661 -373
rect 660 -381 661 -379
rect 667 -375 668 -373
rect 667 -381 668 -379
rect 674 -375 675 -373
rect 674 -381 675 -379
rect 681 -375 682 -373
rect 681 -381 682 -379
rect 688 -375 689 -373
rect 688 -381 689 -379
rect 695 -375 696 -373
rect 695 -381 696 -379
rect 702 -375 703 -373
rect 702 -381 703 -379
rect 709 -375 710 -373
rect 709 -381 710 -379
rect 716 -375 717 -373
rect 716 -381 717 -379
rect 723 -375 724 -373
rect 723 -381 724 -379
rect 730 -375 731 -373
rect 730 -381 731 -379
rect 737 -375 738 -373
rect 737 -381 738 -379
rect 744 -375 745 -373
rect 744 -381 745 -379
rect 751 -375 752 -373
rect 751 -381 752 -379
rect 758 -375 759 -373
rect 758 -381 759 -379
rect 765 -375 766 -373
rect 765 -381 766 -379
rect 772 -375 773 -373
rect 772 -381 773 -379
rect 779 -375 780 -373
rect 779 -381 780 -379
rect 786 -375 787 -373
rect 786 -381 787 -379
rect 793 -375 794 -373
rect 793 -381 794 -379
rect 800 -375 801 -373
rect 800 -381 801 -379
rect 807 -375 808 -373
rect 807 -381 808 -379
rect 814 -375 815 -373
rect 814 -381 815 -379
rect 821 -375 822 -373
rect 821 -381 822 -379
rect 828 -375 829 -373
rect 828 -381 829 -379
rect 835 -375 836 -373
rect 835 -381 836 -379
rect 842 -375 843 -373
rect 842 -381 843 -379
rect 849 -375 850 -373
rect 852 -375 853 -373
rect 849 -381 850 -379
rect 852 -381 853 -379
rect 856 -375 857 -373
rect 856 -381 857 -379
rect 863 -375 864 -373
rect 863 -381 864 -379
rect 870 -375 871 -373
rect 870 -381 871 -379
rect 877 -375 878 -373
rect 884 -381 885 -379
rect 891 -375 892 -373
rect 891 -381 892 -379
rect 2 -464 3 -462
rect 2 -470 3 -468
rect 9 -464 10 -462
rect 9 -470 10 -468
rect 16 -464 17 -462
rect 16 -470 17 -468
rect 23 -464 24 -462
rect 23 -470 24 -468
rect 30 -464 31 -462
rect 30 -470 31 -468
rect 37 -464 38 -462
rect 37 -470 38 -468
rect 44 -464 45 -462
rect 54 -464 55 -462
rect 51 -470 52 -468
rect 54 -470 55 -468
rect 58 -464 59 -462
rect 58 -470 59 -468
rect 65 -464 66 -462
rect 65 -470 66 -468
rect 72 -464 73 -462
rect 72 -470 73 -468
rect 79 -464 80 -462
rect 79 -470 80 -468
rect 82 -470 83 -468
rect 86 -464 87 -462
rect 86 -470 87 -468
rect 93 -464 94 -462
rect 93 -470 94 -468
rect 103 -464 104 -462
rect 100 -470 101 -468
rect 107 -464 108 -462
rect 110 -464 111 -462
rect 107 -470 108 -468
rect 114 -464 115 -462
rect 117 -464 118 -462
rect 117 -470 118 -468
rect 121 -464 122 -462
rect 121 -470 122 -468
rect 128 -464 129 -462
rect 128 -470 129 -468
rect 135 -464 136 -462
rect 135 -470 136 -468
rect 142 -464 143 -462
rect 142 -470 143 -468
rect 149 -464 150 -462
rect 149 -470 150 -468
rect 156 -464 157 -462
rect 159 -464 160 -462
rect 163 -464 164 -462
rect 163 -470 164 -468
rect 166 -470 167 -468
rect 170 -464 171 -462
rect 170 -470 171 -468
rect 177 -464 178 -462
rect 177 -470 178 -468
rect 184 -464 185 -462
rect 184 -470 185 -468
rect 191 -464 192 -462
rect 191 -470 192 -468
rect 194 -470 195 -468
rect 198 -464 199 -462
rect 198 -470 199 -468
rect 201 -470 202 -468
rect 205 -464 206 -462
rect 205 -470 206 -468
rect 212 -464 213 -462
rect 215 -464 216 -462
rect 212 -470 213 -468
rect 222 -464 223 -462
rect 219 -470 220 -468
rect 226 -464 227 -462
rect 226 -470 227 -468
rect 233 -464 234 -462
rect 233 -470 234 -468
rect 240 -464 241 -462
rect 243 -464 244 -462
rect 240 -470 241 -468
rect 243 -470 244 -468
rect 247 -464 248 -462
rect 247 -470 248 -468
rect 254 -464 255 -462
rect 254 -470 255 -468
rect 261 -464 262 -462
rect 261 -470 262 -468
rect 268 -464 269 -462
rect 268 -470 269 -468
rect 275 -464 276 -462
rect 275 -470 276 -468
rect 282 -464 283 -462
rect 282 -470 283 -468
rect 289 -464 290 -462
rect 289 -470 290 -468
rect 296 -464 297 -462
rect 299 -464 300 -462
rect 296 -470 297 -468
rect 303 -464 304 -462
rect 306 -464 307 -462
rect 303 -470 304 -468
rect 306 -470 307 -468
rect 310 -464 311 -462
rect 310 -470 311 -468
rect 317 -464 318 -462
rect 317 -470 318 -468
rect 324 -464 325 -462
rect 324 -470 325 -468
rect 331 -464 332 -462
rect 331 -470 332 -468
rect 338 -464 339 -462
rect 338 -470 339 -468
rect 348 -464 349 -462
rect 345 -470 346 -468
rect 348 -470 349 -468
rect 352 -464 353 -462
rect 352 -470 353 -468
rect 359 -464 360 -462
rect 359 -470 360 -468
rect 366 -464 367 -462
rect 369 -464 370 -462
rect 366 -470 367 -468
rect 369 -470 370 -468
rect 373 -464 374 -462
rect 373 -470 374 -468
rect 383 -464 384 -462
rect 380 -470 381 -468
rect 383 -470 384 -468
rect 387 -464 388 -462
rect 390 -464 391 -462
rect 387 -470 388 -468
rect 394 -464 395 -462
rect 394 -470 395 -468
rect 401 -464 402 -462
rect 401 -470 402 -468
rect 408 -464 409 -462
rect 408 -470 409 -468
rect 415 -464 416 -462
rect 418 -464 419 -462
rect 415 -470 416 -468
rect 418 -470 419 -468
rect 422 -464 423 -462
rect 422 -470 423 -468
rect 429 -464 430 -462
rect 432 -464 433 -462
rect 429 -470 430 -468
rect 432 -470 433 -468
rect 436 -464 437 -462
rect 436 -470 437 -468
rect 439 -470 440 -468
rect 443 -464 444 -462
rect 443 -470 444 -468
rect 450 -464 451 -462
rect 450 -470 451 -468
rect 457 -464 458 -462
rect 457 -470 458 -468
rect 460 -470 461 -468
rect 464 -464 465 -462
rect 464 -470 465 -468
rect 471 -464 472 -462
rect 471 -470 472 -468
rect 478 -464 479 -462
rect 478 -470 479 -468
rect 485 -464 486 -462
rect 485 -470 486 -468
rect 488 -470 489 -468
rect 492 -464 493 -462
rect 492 -470 493 -468
rect 499 -464 500 -462
rect 502 -464 503 -462
rect 499 -470 500 -468
rect 509 -464 510 -462
rect 506 -470 507 -468
rect 513 -464 514 -462
rect 513 -470 514 -468
rect 520 -464 521 -462
rect 523 -464 524 -462
rect 520 -470 521 -468
rect 523 -470 524 -468
rect 527 -464 528 -462
rect 527 -470 528 -468
rect 534 -464 535 -462
rect 534 -470 535 -468
rect 541 -464 542 -462
rect 541 -470 542 -468
rect 548 -464 549 -462
rect 548 -470 549 -468
rect 555 -464 556 -462
rect 555 -470 556 -468
rect 562 -464 563 -462
rect 562 -470 563 -468
rect 569 -464 570 -462
rect 569 -470 570 -468
rect 576 -464 577 -462
rect 576 -470 577 -468
rect 583 -464 584 -462
rect 583 -470 584 -468
rect 590 -464 591 -462
rect 590 -470 591 -468
rect 597 -464 598 -462
rect 597 -470 598 -468
rect 604 -464 605 -462
rect 604 -470 605 -468
rect 611 -464 612 -462
rect 611 -470 612 -468
rect 618 -464 619 -462
rect 621 -464 622 -462
rect 625 -464 626 -462
rect 625 -470 626 -468
rect 632 -464 633 -462
rect 632 -470 633 -468
rect 639 -464 640 -462
rect 639 -470 640 -468
rect 646 -464 647 -462
rect 646 -470 647 -468
rect 653 -464 654 -462
rect 653 -470 654 -468
rect 660 -464 661 -462
rect 660 -470 661 -468
rect 667 -464 668 -462
rect 667 -470 668 -468
rect 674 -464 675 -462
rect 674 -470 675 -468
rect 681 -464 682 -462
rect 681 -470 682 -468
rect 688 -464 689 -462
rect 688 -470 689 -468
rect 695 -464 696 -462
rect 695 -470 696 -468
rect 702 -464 703 -462
rect 702 -470 703 -468
rect 709 -464 710 -462
rect 709 -470 710 -468
rect 716 -464 717 -462
rect 716 -470 717 -468
rect 723 -464 724 -462
rect 723 -470 724 -468
rect 730 -464 731 -462
rect 730 -470 731 -468
rect 737 -464 738 -462
rect 737 -470 738 -468
rect 744 -464 745 -462
rect 744 -470 745 -468
rect 751 -464 752 -462
rect 751 -470 752 -468
rect 758 -464 759 -462
rect 758 -470 759 -468
rect 765 -464 766 -462
rect 765 -470 766 -468
rect 772 -464 773 -462
rect 772 -470 773 -468
rect 779 -464 780 -462
rect 779 -470 780 -468
rect 786 -464 787 -462
rect 786 -470 787 -468
rect 793 -464 794 -462
rect 793 -470 794 -468
rect 800 -464 801 -462
rect 800 -470 801 -468
rect 807 -464 808 -462
rect 807 -470 808 -468
rect 814 -464 815 -462
rect 814 -470 815 -468
rect 821 -464 822 -462
rect 821 -470 822 -468
rect 828 -464 829 -462
rect 828 -470 829 -468
rect 835 -464 836 -462
rect 835 -470 836 -468
rect 842 -464 843 -462
rect 842 -470 843 -468
rect 849 -464 850 -462
rect 849 -470 850 -468
rect 856 -464 857 -462
rect 856 -470 857 -468
rect 863 -464 864 -462
rect 863 -470 864 -468
rect 870 -464 871 -462
rect 870 -470 871 -468
rect 877 -464 878 -462
rect 877 -470 878 -468
rect 884 -464 885 -462
rect 884 -470 885 -468
rect 891 -464 892 -462
rect 891 -470 892 -468
rect 898 -464 899 -462
rect 898 -470 899 -468
rect 905 -464 906 -462
rect 905 -470 906 -468
rect 912 -464 913 -462
rect 912 -470 913 -468
rect 919 -464 920 -462
rect 919 -470 920 -468
rect 926 -464 927 -462
rect 926 -470 927 -468
rect 933 -464 934 -462
rect 933 -470 934 -468
rect 940 -464 941 -462
rect 940 -470 941 -468
rect 947 -464 948 -462
rect 947 -470 948 -468
rect 2 -551 3 -549
rect 2 -557 3 -555
rect 9 -551 10 -549
rect 9 -557 10 -555
rect 16 -551 17 -549
rect 16 -557 17 -555
rect 23 -557 24 -555
rect 30 -551 31 -549
rect 30 -557 31 -555
rect 37 -551 38 -549
rect 37 -557 38 -555
rect 44 -551 45 -549
rect 51 -551 52 -549
rect 51 -557 52 -555
rect 58 -551 59 -549
rect 58 -557 59 -555
rect 65 -551 66 -549
rect 65 -557 66 -555
rect 72 -551 73 -549
rect 72 -557 73 -555
rect 79 -551 80 -549
rect 79 -557 80 -555
rect 86 -551 87 -549
rect 86 -557 87 -555
rect 93 -551 94 -549
rect 96 -551 97 -549
rect 93 -557 94 -555
rect 96 -557 97 -555
rect 100 -551 101 -549
rect 100 -557 101 -555
rect 107 -551 108 -549
rect 107 -557 108 -555
rect 114 -551 115 -549
rect 114 -557 115 -555
rect 121 -551 122 -549
rect 121 -557 122 -555
rect 128 -551 129 -549
rect 128 -557 129 -555
rect 135 -551 136 -549
rect 135 -557 136 -555
rect 145 -551 146 -549
rect 145 -557 146 -555
rect 149 -551 150 -549
rect 149 -557 150 -555
rect 156 -551 157 -549
rect 159 -557 160 -555
rect 163 -551 164 -549
rect 166 -551 167 -549
rect 166 -557 167 -555
rect 170 -551 171 -549
rect 170 -557 171 -555
rect 180 -551 181 -549
rect 177 -557 178 -555
rect 180 -557 181 -555
rect 184 -551 185 -549
rect 184 -557 185 -555
rect 191 -551 192 -549
rect 191 -557 192 -555
rect 198 -551 199 -549
rect 198 -557 199 -555
rect 205 -551 206 -549
rect 205 -557 206 -555
rect 212 -557 213 -555
rect 215 -557 216 -555
rect 219 -551 220 -549
rect 219 -557 220 -555
rect 226 -551 227 -549
rect 226 -557 227 -555
rect 233 -551 234 -549
rect 233 -557 234 -555
rect 240 -551 241 -549
rect 243 -551 244 -549
rect 243 -557 244 -555
rect 247 -551 248 -549
rect 247 -557 248 -555
rect 254 -551 255 -549
rect 254 -557 255 -555
rect 261 -551 262 -549
rect 264 -551 265 -549
rect 261 -557 262 -555
rect 264 -557 265 -555
rect 268 -551 269 -549
rect 268 -557 269 -555
rect 275 -551 276 -549
rect 275 -557 276 -555
rect 282 -551 283 -549
rect 282 -557 283 -555
rect 289 -551 290 -549
rect 289 -557 290 -555
rect 296 -551 297 -549
rect 296 -557 297 -555
rect 303 -551 304 -549
rect 303 -557 304 -555
rect 310 -551 311 -549
rect 313 -551 314 -549
rect 313 -557 314 -555
rect 320 -551 321 -549
rect 317 -557 318 -555
rect 324 -551 325 -549
rect 324 -557 325 -555
rect 334 -551 335 -549
rect 331 -557 332 -555
rect 341 -551 342 -549
rect 338 -557 339 -555
rect 341 -557 342 -555
rect 345 -551 346 -549
rect 345 -557 346 -555
rect 352 -551 353 -549
rect 352 -557 353 -555
rect 359 -557 360 -555
rect 362 -557 363 -555
rect 366 -551 367 -549
rect 366 -557 367 -555
rect 373 -551 374 -549
rect 373 -557 374 -555
rect 380 -551 381 -549
rect 380 -557 381 -555
rect 387 -551 388 -549
rect 390 -551 391 -549
rect 387 -557 388 -555
rect 390 -557 391 -555
rect 394 -551 395 -549
rect 394 -557 395 -555
rect 401 -551 402 -549
rect 401 -557 402 -555
rect 408 -551 409 -549
rect 408 -557 409 -555
rect 415 -551 416 -549
rect 422 -551 423 -549
rect 425 -551 426 -549
rect 422 -557 423 -555
rect 425 -557 426 -555
rect 429 -551 430 -549
rect 429 -557 430 -555
rect 436 -551 437 -549
rect 436 -557 437 -555
rect 443 -551 444 -549
rect 443 -557 444 -555
rect 450 -551 451 -549
rect 453 -551 454 -549
rect 450 -557 451 -555
rect 453 -557 454 -555
rect 457 -551 458 -549
rect 457 -557 458 -555
rect 464 -551 465 -549
rect 464 -557 465 -555
rect 471 -551 472 -549
rect 471 -557 472 -555
rect 478 -551 479 -549
rect 481 -551 482 -549
rect 481 -557 482 -555
rect 485 -551 486 -549
rect 485 -557 486 -555
rect 495 -551 496 -549
rect 492 -557 493 -555
rect 495 -557 496 -555
rect 499 -551 500 -549
rect 502 -551 503 -549
rect 499 -557 500 -555
rect 502 -557 503 -555
rect 509 -551 510 -549
rect 509 -557 510 -555
rect 513 -551 514 -549
rect 513 -557 514 -555
rect 520 -551 521 -549
rect 520 -557 521 -555
rect 527 -551 528 -549
rect 527 -557 528 -555
rect 534 -551 535 -549
rect 534 -557 535 -555
rect 541 -551 542 -549
rect 544 -551 545 -549
rect 544 -557 545 -555
rect 548 -551 549 -549
rect 548 -557 549 -555
rect 555 -551 556 -549
rect 555 -557 556 -555
rect 562 -551 563 -549
rect 562 -557 563 -555
rect 569 -551 570 -549
rect 569 -557 570 -555
rect 576 -551 577 -549
rect 576 -557 577 -555
rect 583 -551 584 -549
rect 583 -557 584 -555
rect 590 -551 591 -549
rect 590 -557 591 -555
rect 597 -551 598 -549
rect 597 -557 598 -555
rect 607 -551 608 -549
rect 607 -557 608 -555
rect 611 -551 612 -549
rect 611 -557 612 -555
rect 618 -551 619 -549
rect 618 -557 619 -555
rect 625 -551 626 -549
rect 625 -557 626 -555
rect 632 -551 633 -549
rect 632 -557 633 -555
rect 639 -551 640 -549
rect 639 -557 640 -555
rect 646 -551 647 -549
rect 646 -557 647 -555
rect 653 -551 654 -549
rect 653 -557 654 -555
rect 660 -551 661 -549
rect 660 -557 661 -555
rect 667 -551 668 -549
rect 667 -557 668 -555
rect 674 -551 675 -549
rect 674 -557 675 -555
rect 681 -551 682 -549
rect 681 -557 682 -555
rect 688 -551 689 -549
rect 688 -557 689 -555
rect 695 -551 696 -549
rect 695 -557 696 -555
rect 702 -551 703 -549
rect 702 -557 703 -555
rect 709 -551 710 -549
rect 709 -557 710 -555
rect 716 -551 717 -549
rect 716 -557 717 -555
rect 723 -551 724 -549
rect 726 -551 727 -549
rect 723 -557 724 -555
rect 726 -557 727 -555
rect 730 -551 731 -549
rect 730 -557 731 -555
rect 737 -551 738 -549
rect 737 -557 738 -555
rect 744 -551 745 -549
rect 744 -557 745 -555
rect 754 -551 755 -549
rect 751 -557 752 -555
rect 754 -557 755 -555
rect 758 -551 759 -549
rect 758 -557 759 -555
rect 765 -551 766 -549
rect 765 -557 766 -555
rect 772 -551 773 -549
rect 772 -557 773 -555
rect 779 -551 780 -549
rect 779 -557 780 -555
rect 786 -551 787 -549
rect 786 -557 787 -555
rect 796 -551 797 -549
rect 793 -557 794 -555
rect 800 -551 801 -549
rect 800 -557 801 -555
rect 807 -551 808 -549
rect 807 -557 808 -555
rect 814 -551 815 -549
rect 814 -557 815 -555
rect 821 -551 822 -549
rect 821 -557 822 -555
rect 835 -551 836 -549
rect 835 -557 836 -555
rect 856 -551 857 -549
rect 856 -557 857 -555
rect 2 -634 3 -632
rect 2 -640 3 -638
rect 9 -634 10 -632
rect 9 -640 10 -638
rect 16 -634 17 -632
rect 16 -640 17 -638
rect 23 -634 24 -632
rect 23 -640 24 -638
rect 30 -634 31 -632
rect 30 -640 31 -638
rect 40 -634 41 -632
rect 44 -634 45 -632
rect 44 -640 45 -638
rect 51 -634 52 -632
rect 51 -640 52 -638
rect 61 -634 62 -632
rect 58 -640 59 -638
rect 61 -640 62 -638
rect 65 -634 66 -632
rect 65 -640 66 -638
rect 72 -634 73 -632
rect 72 -640 73 -638
rect 79 -634 80 -632
rect 79 -640 80 -638
rect 86 -634 87 -632
rect 86 -640 87 -638
rect 93 -634 94 -632
rect 93 -640 94 -638
rect 103 -634 104 -632
rect 100 -640 101 -638
rect 103 -640 104 -638
rect 107 -634 108 -632
rect 107 -640 108 -638
rect 114 -634 115 -632
rect 114 -640 115 -638
rect 124 -634 125 -632
rect 121 -640 122 -638
rect 131 -634 132 -632
rect 128 -640 129 -638
rect 135 -634 136 -632
rect 135 -640 136 -638
rect 138 -640 139 -638
rect 142 -640 143 -638
rect 145 -640 146 -638
rect 149 -634 150 -632
rect 149 -640 150 -638
rect 156 -634 157 -632
rect 156 -640 157 -638
rect 163 -634 164 -632
rect 163 -640 164 -638
rect 173 -634 174 -632
rect 170 -640 171 -638
rect 173 -640 174 -638
rect 177 -634 178 -632
rect 177 -640 178 -638
rect 184 -634 185 -632
rect 184 -640 185 -638
rect 191 -634 192 -632
rect 191 -640 192 -638
rect 198 -634 199 -632
rect 198 -640 199 -638
rect 205 -634 206 -632
rect 205 -640 206 -638
rect 212 -634 213 -632
rect 212 -640 213 -638
rect 219 -634 220 -632
rect 219 -640 220 -638
rect 226 -634 227 -632
rect 226 -640 227 -638
rect 233 -634 234 -632
rect 236 -634 237 -632
rect 236 -640 237 -638
rect 240 -634 241 -632
rect 240 -640 241 -638
rect 243 -640 244 -638
rect 247 -634 248 -632
rect 247 -640 248 -638
rect 254 -634 255 -632
rect 254 -640 255 -638
rect 261 -634 262 -632
rect 261 -640 262 -638
rect 268 -634 269 -632
rect 268 -640 269 -638
rect 275 -634 276 -632
rect 275 -640 276 -638
rect 282 -634 283 -632
rect 282 -640 283 -638
rect 289 -634 290 -632
rect 289 -640 290 -638
rect 296 -634 297 -632
rect 296 -640 297 -638
rect 306 -634 307 -632
rect 303 -640 304 -638
rect 310 -634 311 -632
rect 313 -634 314 -632
rect 310 -640 311 -638
rect 317 -634 318 -632
rect 317 -640 318 -638
rect 324 -634 325 -632
rect 324 -640 325 -638
rect 331 -634 332 -632
rect 334 -634 335 -632
rect 331 -640 332 -638
rect 338 -634 339 -632
rect 341 -634 342 -632
rect 338 -640 339 -638
rect 341 -640 342 -638
rect 345 -634 346 -632
rect 348 -634 349 -632
rect 352 -634 353 -632
rect 352 -640 353 -638
rect 359 -634 360 -632
rect 359 -640 360 -638
rect 366 -634 367 -632
rect 366 -640 367 -638
rect 373 -634 374 -632
rect 373 -640 374 -638
rect 380 -634 381 -632
rect 380 -640 381 -638
rect 387 -634 388 -632
rect 387 -640 388 -638
rect 394 -634 395 -632
rect 394 -640 395 -638
rect 401 -634 402 -632
rect 404 -634 405 -632
rect 401 -640 402 -638
rect 404 -640 405 -638
rect 408 -634 409 -632
rect 408 -640 409 -638
rect 415 -634 416 -632
rect 415 -640 416 -638
rect 422 -634 423 -632
rect 422 -640 423 -638
rect 429 -634 430 -632
rect 429 -640 430 -638
rect 436 -634 437 -632
rect 436 -640 437 -638
rect 443 -634 444 -632
rect 443 -640 444 -638
rect 450 -634 451 -632
rect 453 -640 454 -638
rect 457 -634 458 -632
rect 457 -640 458 -638
rect 464 -634 465 -632
rect 467 -634 468 -632
rect 464 -640 465 -638
rect 467 -640 468 -638
rect 471 -634 472 -632
rect 474 -634 475 -632
rect 471 -640 472 -638
rect 474 -640 475 -638
rect 478 -634 479 -632
rect 478 -640 479 -638
rect 485 -634 486 -632
rect 485 -640 486 -638
rect 492 -634 493 -632
rect 492 -640 493 -638
rect 499 -634 500 -632
rect 499 -640 500 -638
rect 506 -634 507 -632
rect 506 -640 507 -638
rect 513 -634 514 -632
rect 513 -640 514 -638
rect 523 -634 524 -632
rect 520 -640 521 -638
rect 523 -640 524 -638
rect 527 -634 528 -632
rect 527 -640 528 -638
rect 537 -634 538 -632
rect 537 -640 538 -638
rect 541 -634 542 -632
rect 544 -634 545 -632
rect 541 -640 542 -638
rect 548 -634 549 -632
rect 548 -640 549 -638
rect 555 -634 556 -632
rect 555 -640 556 -638
rect 562 -634 563 -632
rect 562 -640 563 -638
rect 569 -634 570 -632
rect 569 -640 570 -638
rect 576 -634 577 -632
rect 576 -640 577 -638
rect 583 -634 584 -632
rect 583 -640 584 -638
rect 590 -634 591 -632
rect 593 -634 594 -632
rect 593 -640 594 -638
rect 597 -634 598 -632
rect 597 -640 598 -638
rect 604 -634 605 -632
rect 604 -640 605 -638
rect 611 -634 612 -632
rect 611 -640 612 -638
rect 614 -640 615 -638
rect 621 -640 622 -638
rect 625 -634 626 -632
rect 625 -640 626 -638
rect 632 -634 633 -632
rect 632 -640 633 -638
rect 639 -634 640 -632
rect 639 -640 640 -638
rect 646 -634 647 -632
rect 646 -640 647 -638
rect 653 -634 654 -632
rect 653 -640 654 -638
rect 660 -634 661 -632
rect 660 -640 661 -638
rect 667 -634 668 -632
rect 667 -640 668 -638
rect 674 -634 675 -632
rect 674 -640 675 -638
rect 681 -634 682 -632
rect 681 -640 682 -638
rect 688 -634 689 -632
rect 688 -640 689 -638
rect 698 -634 699 -632
rect 702 -634 703 -632
rect 702 -640 703 -638
rect 709 -634 710 -632
rect 709 -640 710 -638
rect 716 -634 717 -632
rect 716 -640 717 -638
rect 723 -634 724 -632
rect 723 -640 724 -638
rect 730 -634 731 -632
rect 730 -640 731 -638
rect 737 -634 738 -632
rect 737 -640 738 -638
rect 744 -634 745 -632
rect 744 -640 745 -638
rect 751 -634 752 -632
rect 751 -640 752 -638
rect 758 -634 759 -632
rect 758 -640 759 -638
rect 765 -634 766 -632
rect 765 -640 766 -638
rect 772 -634 773 -632
rect 772 -640 773 -638
rect 779 -634 780 -632
rect 779 -640 780 -638
rect 786 -634 787 -632
rect 786 -640 787 -638
rect 793 -634 794 -632
rect 793 -640 794 -638
rect 800 -634 801 -632
rect 800 -640 801 -638
rect 807 -634 808 -632
rect 807 -640 808 -638
rect 814 -634 815 -632
rect 814 -640 815 -638
rect 821 -634 822 -632
rect 821 -640 822 -638
rect 828 -634 829 -632
rect 828 -640 829 -638
rect 835 -634 836 -632
rect 835 -640 836 -638
rect 842 -634 843 -632
rect 842 -640 843 -638
rect 849 -634 850 -632
rect 849 -640 850 -638
rect 856 -634 857 -632
rect 856 -640 857 -638
rect 863 -634 864 -632
rect 863 -640 864 -638
rect 870 -634 871 -632
rect 870 -640 871 -638
rect 877 -634 878 -632
rect 877 -640 878 -638
rect 884 -634 885 -632
rect 884 -640 885 -638
rect 891 -634 892 -632
rect 891 -640 892 -638
rect 898 -634 899 -632
rect 898 -640 899 -638
rect 905 -634 906 -632
rect 905 -640 906 -638
rect 912 -634 913 -632
rect 912 -640 913 -638
rect 919 -640 920 -638
rect 926 -634 927 -632
rect 926 -640 927 -638
rect 947 -634 948 -632
rect 947 -640 948 -638
rect 2 -713 3 -711
rect 2 -719 3 -717
rect 9 -713 10 -711
rect 9 -719 10 -717
rect 16 -713 17 -711
rect 16 -719 17 -717
rect 26 -719 27 -717
rect 30 -719 31 -717
rect 33 -719 34 -717
rect 37 -713 38 -711
rect 37 -719 38 -717
rect 44 -713 45 -711
rect 44 -719 45 -717
rect 51 -713 52 -711
rect 51 -719 52 -717
rect 58 -713 59 -711
rect 58 -719 59 -717
rect 65 -713 66 -711
rect 65 -719 66 -717
rect 72 -713 73 -711
rect 72 -719 73 -717
rect 79 -713 80 -711
rect 79 -719 80 -717
rect 86 -713 87 -711
rect 89 -713 90 -711
rect 86 -719 87 -717
rect 89 -719 90 -717
rect 93 -713 94 -711
rect 93 -719 94 -717
rect 100 -713 101 -711
rect 103 -713 104 -711
rect 100 -719 101 -717
rect 103 -719 104 -717
rect 110 -713 111 -711
rect 107 -719 108 -717
rect 110 -719 111 -717
rect 114 -713 115 -711
rect 114 -719 115 -717
rect 121 -713 122 -711
rect 121 -719 122 -717
rect 128 -719 129 -717
rect 131 -719 132 -717
rect 135 -713 136 -711
rect 135 -719 136 -717
rect 145 -713 146 -711
rect 142 -719 143 -717
rect 145 -719 146 -717
rect 149 -713 150 -711
rect 149 -719 150 -717
rect 156 -713 157 -711
rect 156 -719 157 -717
rect 163 -713 164 -711
rect 163 -719 164 -717
rect 170 -713 171 -711
rect 170 -719 171 -717
rect 177 -713 178 -711
rect 177 -719 178 -717
rect 184 -713 185 -711
rect 184 -719 185 -717
rect 191 -713 192 -711
rect 191 -719 192 -717
rect 198 -713 199 -711
rect 198 -719 199 -717
rect 205 -713 206 -711
rect 205 -719 206 -717
rect 212 -713 213 -711
rect 212 -719 213 -717
rect 219 -713 220 -711
rect 219 -719 220 -717
rect 229 -713 230 -711
rect 229 -719 230 -717
rect 233 -713 234 -711
rect 233 -719 234 -717
rect 240 -713 241 -711
rect 243 -713 244 -711
rect 240 -719 241 -717
rect 243 -719 244 -717
rect 250 -713 251 -711
rect 250 -719 251 -717
rect 254 -713 255 -711
rect 254 -719 255 -717
rect 261 -713 262 -711
rect 261 -719 262 -717
rect 268 -713 269 -711
rect 268 -719 269 -717
rect 275 -713 276 -711
rect 275 -719 276 -717
rect 282 -713 283 -711
rect 282 -719 283 -717
rect 289 -713 290 -711
rect 289 -719 290 -717
rect 296 -713 297 -711
rect 296 -719 297 -717
rect 303 -713 304 -711
rect 303 -719 304 -717
rect 310 -713 311 -711
rect 310 -719 311 -717
rect 317 -713 318 -711
rect 317 -719 318 -717
rect 324 -713 325 -711
rect 324 -719 325 -717
rect 334 -713 335 -711
rect 338 -713 339 -711
rect 338 -719 339 -717
rect 345 -713 346 -711
rect 348 -713 349 -711
rect 345 -719 346 -717
rect 348 -719 349 -717
rect 352 -713 353 -711
rect 352 -719 353 -717
rect 359 -713 360 -711
rect 359 -719 360 -717
rect 366 -713 367 -711
rect 366 -719 367 -717
rect 373 -719 374 -717
rect 376 -719 377 -717
rect 380 -713 381 -711
rect 380 -719 381 -717
rect 390 -713 391 -711
rect 387 -719 388 -717
rect 394 -713 395 -711
rect 394 -719 395 -717
rect 401 -713 402 -711
rect 401 -719 402 -717
rect 408 -713 409 -711
rect 411 -713 412 -711
rect 408 -719 409 -717
rect 415 -713 416 -711
rect 418 -713 419 -711
rect 415 -719 416 -717
rect 418 -719 419 -717
rect 422 -713 423 -711
rect 422 -719 423 -717
rect 429 -713 430 -711
rect 429 -719 430 -717
rect 436 -713 437 -711
rect 436 -719 437 -717
rect 443 -713 444 -711
rect 443 -719 444 -717
rect 450 -713 451 -711
rect 450 -719 451 -717
rect 457 -713 458 -711
rect 457 -719 458 -717
rect 464 -713 465 -711
rect 464 -719 465 -717
rect 471 -713 472 -711
rect 474 -713 475 -711
rect 478 -713 479 -711
rect 481 -713 482 -711
rect 478 -719 479 -717
rect 481 -719 482 -717
rect 485 -713 486 -711
rect 488 -713 489 -711
rect 485 -719 486 -717
rect 488 -719 489 -717
rect 492 -713 493 -711
rect 492 -719 493 -717
rect 502 -713 503 -711
rect 499 -719 500 -717
rect 502 -719 503 -717
rect 506 -713 507 -711
rect 506 -719 507 -717
rect 513 -719 514 -717
rect 516 -719 517 -717
rect 520 -713 521 -711
rect 520 -719 521 -717
rect 527 -713 528 -711
rect 527 -719 528 -717
rect 534 -713 535 -711
rect 534 -719 535 -717
rect 541 -713 542 -711
rect 544 -713 545 -711
rect 541 -719 542 -717
rect 544 -719 545 -717
rect 548 -713 549 -711
rect 551 -713 552 -711
rect 551 -719 552 -717
rect 555 -713 556 -711
rect 558 -713 559 -711
rect 558 -719 559 -717
rect 562 -713 563 -711
rect 565 -713 566 -711
rect 562 -719 563 -717
rect 569 -713 570 -711
rect 569 -719 570 -717
rect 576 -713 577 -711
rect 576 -719 577 -717
rect 583 -713 584 -711
rect 583 -719 584 -717
rect 590 -713 591 -711
rect 593 -713 594 -711
rect 590 -719 591 -717
rect 597 -713 598 -711
rect 597 -719 598 -717
rect 604 -713 605 -711
rect 604 -719 605 -717
rect 611 -713 612 -711
rect 611 -719 612 -717
rect 618 -713 619 -711
rect 618 -719 619 -717
rect 625 -713 626 -711
rect 628 -713 629 -711
rect 625 -719 626 -717
rect 628 -719 629 -717
rect 632 -713 633 -711
rect 632 -719 633 -717
rect 639 -713 640 -711
rect 639 -719 640 -717
rect 646 -713 647 -711
rect 646 -719 647 -717
rect 653 -713 654 -711
rect 653 -719 654 -717
rect 660 -713 661 -711
rect 660 -719 661 -717
rect 667 -713 668 -711
rect 667 -719 668 -717
rect 674 -713 675 -711
rect 674 -719 675 -717
rect 681 -713 682 -711
rect 681 -719 682 -717
rect 688 -713 689 -711
rect 688 -719 689 -717
rect 695 -713 696 -711
rect 695 -719 696 -717
rect 702 -713 703 -711
rect 702 -719 703 -717
rect 709 -713 710 -711
rect 709 -719 710 -717
rect 716 -713 717 -711
rect 716 -719 717 -717
rect 723 -713 724 -711
rect 723 -719 724 -717
rect 730 -713 731 -711
rect 730 -719 731 -717
rect 737 -713 738 -711
rect 737 -719 738 -717
rect 744 -713 745 -711
rect 744 -719 745 -717
rect 751 -713 752 -711
rect 751 -719 752 -717
rect 758 -713 759 -711
rect 758 -719 759 -717
rect 765 -713 766 -711
rect 765 -719 766 -717
rect 772 -713 773 -711
rect 772 -719 773 -717
rect 779 -713 780 -711
rect 779 -719 780 -717
rect 786 -713 787 -711
rect 786 -719 787 -717
rect 793 -713 794 -711
rect 793 -719 794 -717
rect 800 -713 801 -711
rect 800 -719 801 -717
rect 807 -713 808 -711
rect 807 -719 808 -717
rect 814 -713 815 -711
rect 814 -719 815 -717
rect 821 -713 822 -711
rect 821 -719 822 -717
rect 828 -713 829 -711
rect 828 -719 829 -717
rect 835 -713 836 -711
rect 835 -719 836 -717
rect 842 -713 843 -711
rect 842 -719 843 -717
rect 849 -713 850 -711
rect 849 -719 850 -717
rect 856 -713 857 -711
rect 856 -719 857 -717
rect 863 -713 864 -711
rect 863 -719 864 -717
rect 870 -713 871 -711
rect 870 -719 871 -717
rect 877 -713 878 -711
rect 877 -719 878 -717
rect 887 -713 888 -711
rect 891 -713 892 -711
rect 891 -719 892 -717
rect 898 -713 899 -711
rect 898 -719 899 -717
rect 905 -713 906 -711
rect 905 -719 906 -717
rect 912 -713 913 -711
rect 912 -719 913 -717
rect 919 -713 920 -711
rect 919 -719 920 -717
rect 926 -713 927 -711
rect 926 -719 927 -717
rect 954 -713 955 -711
rect 954 -719 955 -717
rect 1031 -713 1032 -711
rect 1031 -719 1032 -717
rect 23 -784 24 -782
rect 23 -790 24 -788
rect 30 -784 31 -782
rect 30 -790 31 -788
rect 37 -784 38 -782
rect 37 -790 38 -788
rect 44 -784 45 -782
rect 44 -790 45 -788
rect 51 -784 52 -782
rect 58 -784 59 -782
rect 58 -790 59 -788
rect 65 -790 66 -788
rect 72 -790 73 -788
rect 79 -784 80 -782
rect 79 -790 80 -788
rect 86 -784 87 -782
rect 86 -790 87 -788
rect 93 -784 94 -782
rect 93 -790 94 -788
rect 100 -784 101 -782
rect 100 -790 101 -788
rect 107 -784 108 -782
rect 110 -784 111 -782
rect 110 -790 111 -788
rect 114 -784 115 -782
rect 117 -784 118 -782
rect 114 -790 115 -788
rect 121 -784 122 -782
rect 121 -790 122 -788
rect 128 -784 129 -782
rect 128 -790 129 -788
rect 135 -784 136 -782
rect 135 -790 136 -788
rect 142 -784 143 -782
rect 142 -790 143 -788
rect 149 -784 150 -782
rect 149 -790 150 -788
rect 156 -784 157 -782
rect 156 -790 157 -788
rect 163 -784 164 -782
rect 163 -790 164 -788
rect 170 -784 171 -782
rect 170 -790 171 -788
rect 177 -784 178 -782
rect 177 -790 178 -788
rect 184 -784 185 -782
rect 187 -784 188 -782
rect 184 -790 185 -788
rect 191 -784 192 -782
rect 191 -790 192 -788
rect 198 -784 199 -782
rect 198 -790 199 -788
rect 205 -784 206 -782
rect 205 -790 206 -788
rect 212 -784 213 -782
rect 212 -790 213 -788
rect 219 -784 220 -782
rect 219 -790 220 -788
rect 226 -790 227 -788
rect 229 -790 230 -788
rect 236 -784 237 -782
rect 233 -790 234 -788
rect 236 -790 237 -788
rect 243 -784 244 -782
rect 240 -790 241 -788
rect 247 -784 248 -782
rect 247 -790 248 -788
rect 254 -784 255 -782
rect 254 -790 255 -788
rect 261 -784 262 -782
rect 264 -784 265 -782
rect 261 -790 262 -788
rect 268 -784 269 -782
rect 268 -790 269 -788
rect 275 -784 276 -782
rect 275 -790 276 -788
rect 282 -784 283 -782
rect 282 -790 283 -788
rect 289 -784 290 -782
rect 289 -790 290 -788
rect 296 -784 297 -782
rect 296 -790 297 -788
rect 303 -784 304 -782
rect 303 -790 304 -788
rect 310 -784 311 -782
rect 313 -790 314 -788
rect 317 -784 318 -782
rect 317 -790 318 -788
rect 324 -784 325 -782
rect 324 -790 325 -788
rect 331 -784 332 -782
rect 331 -790 332 -788
rect 338 -784 339 -782
rect 345 -784 346 -782
rect 345 -790 346 -788
rect 352 -784 353 -782
rect 355 -784 356 -782
rect 352 -790 353 -788
rect 355 -790 356 -788
rect 359 -784 360 -782
rect 359 -790 360 -788
rect 366 -784 367 -782
rect 366 -790 367 -788
rect 373 -784 374 -782
rect 373 -790 374 -788
rect 380 -784 381 -782
rect 380 -790 381 -788
rect 387 -784 388 -782
rect 390 -784 391 -782
rect 387 -790 388 -788
rect 394 -784 395 -782
rect 394 -790 395 -788
rect 401 -784 402 -782
rect 404 -784 405 -782
rect 408 -784 409 -782
rect 408 -790 409 -788
rect 415 -784 416 -782
rect 415 -790 416 -788
rect 422 -790 423 -788
rect 425 -790 426 -788
rect 429 -784 430 -782
rect 429 -790 430 -788
rect 436 -784 437 -782
rect 436 -790 437 -788
rect 443 -784 444 -782
rect 443 -790 444 -788
rect 450 -784 451 -782
rect 450 -790 451 -788
rect 457 -784 458 -782
rect 457 -790 458 -788
rect 464 -784 465 -782
rect 464 -790 465 -788
rect 471 -784 472 -782
rect 471 -790 472 -788
rect 478 -784 479 -782
rect 478 -790 479 -788
rect 485 -784 486 -782
rect 485 -790 486 -788
rect 492 -784 493 -782
rect 495 -784 496 -782
rect 492 -790 493 -788
rect 499 -784 500 -782
rect 499 -790 500 -788
rect 506 -784 507 -782
rect 506 -790 507 -788
rect 513 -784 514 -782
rect 513 -790 514 -788
rect 516 -790 517 -788
rect 520 -784 521 -782
rect 520 -790 521 -788
rect 527 -784 528 -782
rect 530 -784 531 -782
rect 527 -790 528 -788
rect 530 -790 531 -788
rect 534 -784 535 -782
rect 534 -790 535 -788
rect 541 -784 542 -782
rect 548 -784 549 -782
rect 548 -790 549 -788
rect 555 -784 556 -782
rect 555 -790 556 -788
rect 565 -784 566 -782
rect 562 -790 563 -788
rect 565 -790 566 -788
rect 569 -784 570 -782
rect 569 -790 570 -788
rect 576 -784 577 -782
rect 579 -784 580 -782
rect 576 -790 577 -788
rect 579 -790 580 -788
rect 583 -784 584 -782
rect 583 -790 584 -788
rect 590 -784 591 -782
rect 590 -790 591 -788
rect 597 -784 598 -782
rect 597 -790 598 -788
rect 604 -784 605 -782
rect 604 -790 605 -788
rect 611 -784 612 -782
rect 611 -790 612 -788
rect 618 -784 619 -782
rect 621 -784 622 -782
rect 618 -790 619 -788
rect 621 -790 622 -788
rect 625 -784 626 -782
rect 625 -790 626 -788
rect 632 -784 633 -782
rect 632 -790 633 -788
rect 639 -784 640 -782
rect 639 -790 640 -788
rect 646 -784 647 -782
rect 646 -790 647 -788
rect 653 -784 654 -782
rect 653 -790 654 -788
rect 660 -784 661 -782
rect 660 -790 661 -788
rect 667 -784 668 -782
rect 670 -784 671 -782
rect 667 -790 668 -788
rect 674 -784 675 -782
rect 674 -790 675 -788
rect 681 -784 682 -782
rect 681 -790 682 -788
rect 688 -784 689 -782
rect 688 -790 689 -788
rect 695 -784 696 -782
rect 695 -790 696 -788
rect 702 -784 703 -782
rect 702 -790 703 -788
rect 709 -784 710 -782
rect 709 -790 710 -788
rect 716 -784 717 -782
rect 716 -790 717 -788
rect 723 -784 724 -782
rect 723 -790 724 -788
rect 730 -784 731 -782
rect 730 -790 731 -788
rect 737 -784 738 -782
rect 737 -790 738 -788
rect 744 -784 745 -782
rect 744 -790 745 -788
rect 751 -784 752 -782
rect 751 -790 752 -788
rect 758 -784 759 -782
rect 758 -790 759 -788
rect 765 -784 766 -782
rect 765 -790 766 -788
rect 772 -784 773 -782
rect 772 -790 773 -788
rect 779 -784 780 -782
rect 779 -790 780 -788
rect 786 -784 787 -782
rect 786 -790 787 -788
rect 793 -784 794 -782
rect 793 -790 794 -788
rect 800 -784 801 -782
rect 800 -790 801 -788
rect 807 -784 808 -782
rect 807 -790 808 -788
rect 814 -784 815 -782
rect 814 -790 815 -788
rect 821 -784 822 -782
rect 821 -790 822 -788
rect 828 -784 829 -782
rect 828 -790 829 -788
rect 835 -784 836 -782
rect 835 -790 836 -788
rect 842 -784 843 -782
rect 842 -790 843 -788
rect 849 -784 850 -782
rect 849 -790 850 -788
rect 856 -784 857 -782
rect 856 -790 857 -788
rect 863 -784 864 -782
rect 863 -790 864 -788
rect 870 -784 871 -782
rect 870 -790 871 -788
rect 877 -784 878 -782
rect 877 -790 878 -788
rect 884 -784 885 -782
rect 884 -790 885 -788
rect 891 -784 892 -782
rect 891 -790 892 -788
rect 894 -790 895 -788
rect 898 -784 899 -782
rect 898 -790 899 -788
rect 908 -784 909 -782
rect 905 -790 906 -788
rect 908 -790 909 -788
rect 912 -784 913 -782
rect 915 -784 916 -782
rect 915 -790 916 -788
rect 919 -784 920 -782
rect 919 -790 920 -788
rect 961 -784 962 -782
rect 961 -790 962 -788
rect 975 -784 976 -782
rect 975 -790 976 -788
rect 989 -790 990 -788
rect 1006 -784 1007 -782
rect 1010 -784 1011 -782
rect 1010 -790 1011 -788
rect 1017 -784 1018 -782
rect 1017 -790 1018 -788
rect 1066 -784 1067 -782
rect 1066 -790 1067 -788
rect 2 -881 3 -879
rect 2 -887 3 -885
rect 12 -881 13 -879
rect 16 -881 17 -879
rect 16 -887 17 -885
rect 23 -881 24 -879
rect 23 -887 24 -885
rect 30 -881 31 -879
rect 30 -887 31 -885
rect 37 -881 38 -879
rect 37 -887 38 -885
rect 47 -881 48 -879
rect 44 -887 45 -885
rect 51 -881 52 -879
rect 51 -887 52 -885
rect 58 -881 59 -879
rect 58 -887 59 -885
rect 68 -881 69 -879
rect 72 -881 73 -879
rect 72 -887 73 -885
rect 79 -881 80 -879
rect 79 -887 80 -885
rect 86 -881 87 -879
rect 86 -887 87 -885
rect 93 -881 94 -879
rect 93 -887 94 -885
rect 100 -881 101 -879
rect 100 -887 101 -885
rect 110 -881 111 -879
rect 107 -887 108 -885
rect 110 -887 111 -885
rect 114 -881 115 -879
rect 117 -881 118 -879
rect 114 -887 115 -885
rect 121 -881 122 -879
rect 121 -887 122 -885
rect 131 -881 132 -879
rect 131 -887 132 -885
rect 135 -881 136 -879
rect 138 -881 139 -879
rect 142 -881 143 -879
rect 142 -887 143 -885
rect 149 -881 150 -879
rect 149 -887 150 -885
rect 156 -881 157 -879
rect 156 -887 157 -885
rect 163 -881 164 -879
rect 163 -887 164 -885
rect 170 -881 171 -879
rect 173 -881 174 -879
rect 170 -887 171 -885
rect 173 -887 174 -885
rect 177 -881 178 -879
rect 180 -881 181 -879
rect 180 -887 181 -885
rect 184 -881 185 -879
rect 184 -887 185 -885
rect 191 -881 192 -879
rect 191 -887 192 -885
rect 198 -881 199 -879
rect 198 -887 199 -885
rect 205 -881 206 -879
rect 208 -881 209 -879
rect 208 -887 209 -885
rect 212 -881 213 -879
rect 215 -887 216 -885
rect 219 -881 220 -879
rect 222 -887 223 -885
rect 229 -881 230 -879
rect 229 -887 230 -885
rect 233 -881 234 -879
rect 233 -887 234 -885
rect 240 -881 241 -879
rect 243 -881 244 -879
rect 240 -887 241 -885
rect 243 -887 244 -885
rect 247 -881 248 -879
rect 247 -887 248 -885
rect 254 -881 255 -879
rect 254 -887 255 -885
rect 261 -881 262 -879
rect 261 -887 262 -885
rect 268 -881 269 -879
rect 268 -887 269 -885
rect 275 -881 276 -879
rect 275 -887 276 -885
rect 282 -881 283 -879
rect 282 -887 283 -885
rect 289 -881 290 -879
rect 289 -887 290 -885
rect 296 -881 297 -879
rect 296 -887 297 -885
rect 303 -881 304 -879
rect 303 -887 304 -885
rect 310 -881 311 -879
rect 310 -887 311 -885
rect 317 -881 318 -879
rect 317 -887 318 -885
rect 324 -881 325 -879
rect 324 -887 325 -885
rect 331 -881 332 -879
rect 331 -887 332 -885
rect 338 -881 339 -879
rect 338 -887 339 -885
rect 345 -881 346 -879
rect 345 -887 346 -885
rect 352 -881 353 -879
rect 355 -881 356 -879
rect 352 -887 353 -885
rect 355 -887 356 -885
rect 359 -881 360 -879
rect 362 -881 363 -879
rect 366 -881 367 -879
rect 369 -881 370 -879
rect 366 -887 367 -885
rect 369 -887 370 -885
rect 373 -881 374 -879
rect 373 -887 374 -885
rect 380 -881 381 -879
rect 380 -887 381 -885
rect 387 -881 388 -879
rect 387 -887 388 -885
rect 394 -881 395 -879
rect 394 -887 395 -885
rect 401 -881 402 -879
rect 401 -887 402 -885
rect 408 -881 409 -879
rect 411 -881 412 -879
rect 408 -887 409 -885
rect 411 -887 412 -885
rect 415 -881 416 -879
rect 415 -887 416 -885
rect 422 -881 423 -879
rect 422 -887 423 -885
rect 429 -881 430 -879
rect 429 -887 430 -885
rect 436 -881 437 -879
rect 439 -881 440 -879
rect 436 -887 437 -885
rect 439 -887 440 -885
rect 443 -881 444 -879
rect 443 -887 444 -885
rect 450 -881 451 -879
rect 450 -887 451 -885
rect 457 -881 458 -879
rect 457 -887 458 -885
rect 464 -881 465 -879
rect 467 -881 468 -879
rect 467 -887 468 -885
rect 471 -881 472 -879
rect 471 -887 472 -885
rect 478 -881 479 -879
rect 478 -887 479 -885
rect 485 -881 486 -879
rect 485 -887 486 -885
rect 492 -881 493 -879
rect 492 -887 493 -885
rect 499 -887 500 -885
rect 502 -887 503 -885
rect 506 -881 507 -879
rect 506 -887 507 -885
rect 513 -881 514 -879
rect 513 -887 514 -885
rect 520 -881 521 -879
rect 523 -881 524 -879
rect 520 -887 521 -885
rect 523 -887 524 -885
rect 527 -881 528 -879
rect 527 -887 528 -885
rect 534 -881 535 -879
rect 537 -881 538 -879
rect 534 -887 535 -885
rect 537 -887 538 -885
rect 541 -881 542 -879
rect 544 -881 545 -879
rect 548 -881 549 -879
rect 551 -881 552 -879
rect 548 -887 549 -885
rect 551 -887 552 -885
rect 555 -881 556 -879
rect 555 -887 556 -885
rect 562 -881 563 -879
rect 565 -881 566 -879
rect 562 -887 563 -885
rect 572 -881 573 -879
rect 569 -887 570 -885
rect 572 -887 573 -885
rect 576 -881 577 -879
rect 576 -887 577 -885
rect 583 -881 584 -879
rect 583 -887 584 -885
rect 590 -881 591 -879
rect 590 -887 591 -885
rect 597 -881 598 -879
rect 597 -887 598 -885
rect 604 -881 605 -879
rect 604 -887 605 -885
rect 611 -881 612 -879
rect 611 -887 612 -885
rect 618 -881 619 -879
rect 618 -887 619 -885
rect 625 -881 626 -879
rect 625 -887 626 -885
rect 632 -881 633 -879
rect 632 -887 633 -885
rect 639 -881 640 -879
rect 639 -887 640 -885
rect 646 -881 647 -879
rect 646 -887 647 -885
rect 653 -881 654 -879
rect 653 -887 654 -885
rect 660 -881 661 -879
rect 660 -887 661 -885
rect 667 -881 668 -879
rect 670 -881 671 -879
rect 674 -881 675 -879
rect 674 -887 675 -885
rect 681 -881 682 -879
rect 681 -887 682 -885
rect 688 -881 689 -879
rect 688 -887 689 -885
rect 695 -881 696 -879
rect 695 -887 696 -885
rect 702 -881 703 -879
rect 702 -887 703 -885
rect 709 -881 710 -879
rect 709 -887 710 -885
rect 716 -881 717 -879
rect 716 -887 717 -885
rect 723 -881 724 -879
rect 723 -887 724 -885
rect 730 -881 731 -879
rect 730 -887 731 -885
rect 737 -881 738 -879
rect 737 -887 738 -885
rect 744 -881 745 -879
rect 744 -887 745 -885
rect 751 -881 752 -879
rect 751 -887 752 -885
rect 758 -881 759 -879
rect 758 -887 759 -885
rect 765 -881 766 -879
rect 765 -887 766 -885
rect 772 -881 773 -879
rect 772 -887 773 -885
rect 779 -881 780 -879
rect 779 -887 780 -885
rect 786 -881 787 -879
rect 786 -887 787 -885
rect 793 -881 794 -879
rect 793 -887 794 -885
rect 800 -881 801 -879
rect 800 -887 801 -885
rect 807 -881 808 -879
rect 807 -887 808 -885
rect 814 -881 815 -879
rect 817 -881 818 -879
rect 817 -887 818 -885
rect 821 -881 822 -879
rect 821 -887 822 -885
rect 828 -881 829 -879
rect 828 -887 829 -885
rect 835 -881 836 -879
rect 835 -887 836 -885
rect 842 -881 843 -879
rect 842 -887 843 -885
rect 849 -881 850 -879
rect 849 -887 850 -885
rect 856 -881 857 -879
rect 856 -887 857 -885
rect 863 -881 864 -879
rect 863 -887 864 -885
rect 870 -881 871 -879
rect 870 -887 871 -885
rect 877 -881 878 -879
rect 877 -887 878 -885
rect 884 -881 885 -879
rect 884 -887 885 -885
rect 891 -881 892 -879
rect 891 -887 892 -885
rect 898 -881 899 -879
rect 898 -887 899 -885
rect 905 -881 906 -879
rect 905 -887 906 -885
rect 912 -881 913 -879
rect 912 -887 913 -885
rect 919 -881 920 -879
rect 919 -887 920 -885
rect 926 -881 927 -879
rect 926 -887 927 -885
rect 933 -881 934 -879
rect 933 -887 934 -885
rect 940 -881 941 -879
rect 940 -887 941 -885
rect 947 -881 948 -879
rect 947 -887 948 -885
rect 954 -881 955 -879
rect 954 -887 955 -885
rect 961 -881 962 -879
rect 961 -887 962 -885
rect 968 -881 969 -879
rect 968 -887 969 -885
rect 975 -881 976 -879
rect 975 -887 976 -885
rect 982 -881 983 -879
rect 982 -887 983 -885
rect 989 -881 990 -879
rect 992 -881 993 -879
rect 989 -887 990 -885
rect 992 -887 993 -885
rect 996 -881 997 -879
rect 996 -887 997 -885
rect 1003 -881 1004 -879
rect 1003 -887 1004 -885
rect 1013 -881 1014 -879
rect 1010 -887 1011 -885
rect 1013 -887 1014 -885
rect 1017 -881 1018 -879
rect 1017 -887 1018 -885
rect 1024 -881 1025 -879
rect 1024 -887 1025 -885
rect 1038 -881 1039 -879
rect 1038 -887 1039 -885
rect 1080 -881 1081 -879
rect 1080 -887 1081 -885
rect 12 -968 13 -966
rect 16 -962 17 -960
rect 16 -968 17 -966
rect 23 -962 24 -960
rect 23 -968 24 -966
rect 30 -962 31 -960
rect 30 -968 31 -966
rect 37 -962 38 -960
rect 37 -968 38 -966
rect 44 -962 45 -960
rect 44 -968 45 -966
rect 51 -962 52 -960
rect 51 -968 52 -966
rect 58 -962 59 -960
rect 58 -968 59 -966
rect 65 -962 66 -960
rect 65 -968 66 -966
rect 72 -962 73 -960
rect 72 -968 73 -966
rect 79 -962 80 -960
rect 79 -968 80 -966
rect 86 -962 87 -960
rect 86 -968 87 -966
rect 93 -962 94 -960
rect 93 -968 94 -966
rect 100 -962 101 -960
rect 100 -968 101 -966
rect 107 -962 108 -960
rect 107 -968 108 -966
rect 114 -962 115 -960
rect 114 -968 115 -966
rect 121 -962 122 -960
rect 121 -968 122 -966
rect 128 -968 129 -966
rect 131 -968 132 -966
rect 135 -962 136 -960
rect 135 -968 136 -966
rect 142 -962 143 -960
rect 142 -968 143 -966
rect 149 -962 150 -960
rect 149 -968 150 -966
rect 156 -962 157 -960
rect 156 -968 157 -966
rect 163 -962 164 -960
rect 163 -968 164 -966
rect 170 -962 171 -960
rect 170 -968 171 -966
rect 180 -962 181 -960
rect 177 -968 178 -966
rect 180 -968 181 -966
rect 184 -962 185 -960
rect 184 -968 185 -966
rect 191 -962 192 -960
rect 191 -968 192 -966
rect 198 -962 199 -960
rect 198 -968 199 -966
rect 205 -962 206 -960
rect 205 -968 206 -966
rect 212 -962 213 -960
rect 215 -962 216 -960
rect 219 -962 220 -960
rect 222 -962 223 -960
rect 222 -968 223 -966
rect 226 -962 227 -960
rect 226 -968 227 -966
rect 233 -962 234 -960
rect 236 -962 237 -960
rect 240 -962 241 -960
rect 240 -968 241 -966
rect 243 -968 244 -966
rect 247 -962 248 -960
rect 247 -968 248 -966
rect 254 -962 255 -960
rect 254 -968 255 -966
rect 261 -962 262 -960
rect 261 -968 262 -966
rect 268 -962 269 -960
rect 268 -968 269 -966
rect 275 -962 276 -960
rect 278 -962 279 -960
rect 282 -962 283 -960
rect 285 -962 286 -960
rect 285 -968 286 -966
rect 289 -962 290 -960
rect 289 -968 290 -966
rect 296 -962 297 -960
rect 296 -968 297 -966
rect 303 -962 304 -960
rect 303 -968 304 -966
rect 310 -962 311 -960
rect 310 -968 311 -966
rect 317 -962 318 -960
rect 317 -968 318 -966
rect 324 -962 325 -960
rect 324 -968 325 -966
rect 327 -968 328 -966
rect 331 -962 332 -960
rect 331 -968 332 -966
rect 338 -962 339 -960
rect 338 -968 339 -966
rect 345 -962 346 -960
rect 345 -968 346 -966
rect 352 -962 353 -960
rect 352 -968 353 -966
rect 359 -962 360 -960
rect 359 -968 360 -966
rect 362 -968 363 -966
rect 366 -962 367 -960
rect 366 -968 367 -966
rect 373 -962 374 -960
rect 373 -968 374 -966
rect 380 -968 381 -966
rect 383 -968 384 -966
rect 387 -962 388 -960
rect 387 -968 388 -966
rect 397 -968 398 -966
rect 401 -962 402 -960
rect 401 -968 402 -966
rect 408 -962 409 -960
rect 408 -968 409 -966
rect 415 -962 416 -960
rect 418 -962 419 -960
rect 418 -968 419 -966
rect 422 -962 423 -960
rect 422 -968 423 -966
rect 429 -962 430 -960
rect 429 -968 430 -966
rect 439 -962 440 -960
rect 436 -968 437 -966
rect 439 -968 440 -966
rect 443 -962 444 -960
rect 443 -968 444 -966
rect 450 -968 451 -966
rect 453 -968 454 -966
rect 457 -962 458 -960
rect 457 -968 458 -966
rect 464 -962 465 -960
rect 464 -968 465 -966
rect 471 -962 472 -960
rect 474 -962 475 -960
rect 471 -968 472 -966
rect 474 -968 475 -966
rect 478 -962 479 -960
rect 478 -968 479 -966
rect 481 -968 482 -966
rect 485 -962 486 -960
rect 485 -968 486 -966
rect 492 -962 493 -960
rect 492 -968 493 -966
rect 495 -968 496 -966
rect 499 -962 500 -960
rect 499 -968 500 -966
rect 506 -962 507 -960
rect 506 -968 507 -966
rect 513 -962 514 -960
rect 520 -962 521 -960
rect 520 -968 521 -966
rect 530 -962 531 -960
rect 530 -968 531 -966
rect 534 -962 535 -960
rect 534 -968 535 -966
rect 541 -962 542 -960
rect 541 -968 542 -966
rect 548 -962 549 -960
rect 548 -968 549 -966
rect 555 -962 556 -960
rect 555 -968 556 -966
rect 562 -962 563 -960
rect 562 -968 563 -966
rect 565 -968 566 -966
rect 569 -962 570 -960
rect 569 -968 570 -966
rect 576 -962 577 -960
rect 576 -968 577 -966
rect 583 -962 584 -960
rect 583 -968 584 -966
rect 590 -962 591 -960
rect 590 -968 591 -966
rect 597 -962 598 -960
rect 600 -962 601 -960
rect 597 -968 598 -966
rect 600 -968 601 -966
rect 604 -962 605 -960
rect 604 -968 605 -966
rect 607 -968 608 -966
rect 611 -962 612 -960
rect 611 -968 612 -966
rect 618 -962 619 -960
rect 618 -968 619 -966
rect 628 -962 629 -960
rect 625 -968 626 -966
rect 635 -962 636 -960
rect 632 -968 633 -966
rect 635 -968 636 -966
rect 639 -962 640 -960
rect 639 -968 640 -966
rect 646 -962 647 -960
rect 646 -968 647 -966
rect 656 -962 657 -960
rect 653 -968 654 -966
rect 660 -962 661 -960
rect 660 -968 661 -966
rect 667 -962 668 -960
rect 667 -968 668 -966
rect 674 -962 675 -960
rect 674 -968 675 -966
rect 681 -962 682 -960
rect 681 -968 682 -966
rect 688 -962 689 -960
rect 688 -968 689 -966
rect 695 -962 696 -960
rect 695 -968 696 -966
rect 698 -968 699 -966
rect 702 -962 703 -960
rect 702 -968 703 -966
rect 709 -962 710 -960
rect 709 -968 710 -966
rect 716 -962 717 -960
rect 716 -968 717 -966
rect 723 -962 724 -960
rect 723 -968 724 -966
rect 730 -962 731 -960
rect 730 -968 731 -966
rect 737 -962 738 -960
rect 737 -968 738 -966
rect 744 -962 745 -960
rect 744 -968 745 -966
rect 751 -962 752 -960
rect 751 -968 752 -966
rect 758 -962 759 -960
rect 758 -968 759 -966
rect 765 -962 766 -960
rect 765 -968 766 -966
rect 772 -962 773 -960
rect 772 -968 773 -966
rect 779 -962 780 -960
rect 779 -968 780 -966
rect 786 -962 787 -960
rect 786 -968 787 -966
rect 793 -962 794 -960
rect 793 -968 794 -966
rect 800 -962 801 -960
rect 800 -968 801 -966
rect 807 -962 808 -960
rect 807 -968 808 -966
rect 814 -962 815 -960
rect 814 -968 815 -966
rect 821 -962 822 -960
rect 821 -968 822 -966
rect 828 -962 829 -960
rect 828 -968 829 -966
rect 835 -962 836 -960
rect 835 -968 836 -966
rect 842 -962 843 -960
rect 842 -968 843 -966
rect 849 -962 850 -960
rect 849 -968 850 -966
rect 856 -962 857 -960
rect 856 -968 857 -966
rect 863 -962 864 -960
rect 863 -968 864 -966
rect 870 -962 871 -960
rect 870 -968 871 -966
rect 877 -962 878 -960
rect 877 -968 878 -966
rect 884 -962 885 -960
rect 884 -968 885 -966
rect 891 -962 892 -960
rect 891 -968 892 -966
rect 898 -962 899 -960
rect 898 -968 899 -966
rect 905 -962 906 -960
rect 905 -968 906 -966
rect 912 -962 913 -960
rect 915 -962 916 -960
rect 915 -968 916 -966
rect 922 -962 923 -960
rect 919 -968 920 -966
rect 922 -968 923 -966
rect 929 -962 930 -960
rect 926 -968 927 -966
rect 929 -968 930 -966
rect 933 -962 934 -960
rect 933 -968 934 -966
rect 943 -962 944 -960
rect 943 -968 944 -966
rect 947 -962 948 -960
rect 947 -968 948 -966
rect 954 -962 955 -960
rect 954 -968 955 -966
rect 961 -962 962 -960
rect 961 -968 962 -966
rect 968 -962 969 -960
rect 968 -968 969 -966
rect 982 -962 983 -960
rect 982 -968 983 -966
rect 1010 -962 1011 -960
rect 1010 -968 1011 -966
rect 1038 -962 1039 -960
rect 1038 -968 1039 -966
rect 1059 -962 1060 -960
rect 1059 -968 1060 -966
rect 1087 -962 1088 -960
rect 1087 -968 1088 -966
rect 9 -1055 10 -1053
rect 9 -1061 10 -1059
rect 16 -1055 17 -1053
rect 16 -1061 17 -1059
rect 23 -1055 24 -1053
rect 23 -1061 24 -1059
rect 30 -1055 31 -1053
rect 30 -1061 31 -1059
rect 40 -1055 41 -1053
rect 44 -1055 45 -1053
rect 44 -1061 45 -1059
rect 51 -1055 52 -1053
rect 51 -1061 52 -1059
rect 61 -1055 62 -1053
rect 58 -1061 59 -1059
rect 65 -1055 66 -1053
rect 65 -1061 66 -1059
rect 72 -1055 73 -1053
rect 72 -1061 73 -1059
rect 79 -1055 80 -1053
rect 79 -1061 80 -1059
rect 86 -1055 87 -1053
rect 86 -1061 87 -1059
rect 93 -1055 94 -1053
rect 93 -1061 94 -1059
rect 100 -1055 101 -1053
rect 100 -1061 101 -1059
rect 107 -1055 108 -1053
rect 107 -1061 108 -1059
rect 114 -1055 115 -1053
rect 114 -1061 115 -1059
rect 121 -1055 122 -1053
rect 121 -1061 122 -1059
rect 131 -1055 132 -1053
rect 135 -1055 136 -1053
rect 135 -1061 136 -1059
rect 142 -1055 143 -1053
rect 145 -1055 146 -1053
rect 142 -1061 143 -1059
rect 149 -1055 150 -1053
rect 149 -1061 150 -1059
rect 156 -1055 157 -1053
rect 156 -1061 157 -1059
rect 163 -1055 164 -1053
rect 166 -1061 167 -1059
rect 170 -1061 171 -1059
rect 173 -1061 174 -1059
rect 180 -1055 181 -1053
rect 180 -1061 181 -1059
rect 184 -1055 185 -1053
rect 184 -1061 185 -1059
rect 191 -1055 192 -1053
rect 191 -1061 192 -1059
rect 198 -1055 199 -1053
rect 198 -1061 199 -1059
rect 205 -1055 206 -1053
rect 208 -1055 209 -1053
rect 205 -1061 206 -1059
rect 212 -1055 213 -1053
rect 219 -1055 220 -1053
rect 222 -1061 223 -1059
rect 226 -1055 227 -1053
rect 226 -1061 227 -1059
rect 233 -1055 234 -1053
rect 233 -1061 234 -1059
rect 240 -1055 241 -1053
rect 240 -1061 241 -1059
rect 247 -1055 248 -1053
rect 247 -1061 248 -1059
rect 257 -1055 258 -1053
rect 261 -1055 262 -1053
rect 261 -1061 262 -1059
rect 268 -1055 269 -1053
rect 268 -1061 269 -1059
rect 275 -1055 276 -1053
rect 275 -1061 276 -1059
rect 282 -1055 283 -1053
rect 282 -1061 283 -1059
rect 289 -1055 290 -1053
rect 289 -1061 290 -1059
rect 296 -1055 297 -1053
rect 299 -1055 300 -1053
rect 299 -1061 300 -1059
rect 303 -1055 304 -1053
rect 303 -1061 304 -1059
rect 310 -1055 311 -1053
rect 310 -1061 311 -1059
rect 317 -1055 318 -1053
rect 317 -1061 318 -1059
rect 324 -1055 325 -1053
rect 324 -1061 325 -1059
rect 331 -1055 332 -1053
rect 331 -1061 332 -1059
rect 338 -1055 339 -1053
rect 338 -1061 339 -1059
rect 345 -1055 346 -1053
rect 345 -1061 346 -1059
rect 352 -1055 353 -1053
rect 355 -1055 356 -1053
rect 352 -1061 353 -1059
rect 355 -1061 356 -1059
rect 359 -1055 360 -1053
rect 359 -1061 360 -1059
rect 366 -1055 367 -1053
rect 366 -1061 367 -1059
rect 373 -1055 374 -1053
rect 373 -1061 374 -1059
rect 380 -1055 381 -1053
rect 380 -1061 381 -1059
rect 387 -1055 388 -1053
rect 387 -1061 388 -1059
rect 394 -1055 395 -1053
rect 394 -1061 395 -1059
rect 401 -1055 402 -1053
rect 401 -1061 402 -1059
rect 411 -1055 412 -1053
rect 408 -1061 409 -1059
rect 411 -1061 412 -1059
rect 415 -1055 416 -1053
rect 415 -1061 416 -1059
rect 422 -1055 423 -1053
rect 422 -1061 423 -1059
rect 429 -1055 430 -1053
rect 432 -1055 433 -1053
rect 429 -1061 430 -1059
rect 436 -1055 437 -1053
rect 436 -1061 437 -1059
rect 443 -1055 444 -1053
rect 446 -1055 447 -1053
rect 443 -1061 444 -1059
rect 446 -1061 447 -1059
rect 450 -1055 451 -1053
rect 453 -1055 454 -1053
rect 453 -1061 454 -1059
rect 457 -1055 458 -1053
rect 457 -1061 458 -1059
rect 464 -1055 465 -1053
rect 464 -1061 465 -1059
rect 471 -1055 472 -1053
rect 474 -1055 475 -1053
rect 478 -1055 479 -1053
rect 478 -1061 479 -1059
rect 488 -1055 489 -1053
rect 485 -1061 486 -1059
rect 492 -1055 493 -1053
rect 492 -1061 493 -1059
rect 495 -1061 496 -1059
rect 499 -1055 500 -1053
rect 499 -1061 500 -1059
rect 506 -1055 507 -1053
rect 506 -1061 507 -1059
rect 516 -1055 517 -1053
rect 513 -1061 514 -1059
rect 520 -1055 521 -1053
rect 520 -1061 521 -1059
rect 527 -1055 528 -1053
rect 527 -1061 528 -1059
rect 537 -1055 538 -1053
rect 534 -1061 535 -1059
rect 537 -1061 538 -1059
rect 541 -1055 542 -1053
rect 541 -1061 542 -1059
rect 548 -1055 549 -1053
rect 551 -1055 552 -1053
rect 551 -1061 552 -1059
rect 555 -1055 556 -1053
rect 555 -1061 556 -1059
rect 562 -1055 563 -1053
rect 562 -1061 563 -1059
rect 569 -1055 570 -1053
rect 569 -1061 570 -1059
rect 572 -1061 573 -1059
rect 576 -1055 577 -1053
rect 576 -1061 577 -1059
rect 579 -1061 580 -1059
rect 583 -1055 584 -1053
rect 586 -1055 587 -1053
rect 583 -1061 584 -1059
rect 590 -1055 591 -1053
rect 590 -1061 591 -1059
rect 597 -1055 598 -1053
rect 597 -1061 598 -1059
rect 604 -1055 605 -1053
rect 607 -1055 608 -1053
rect 611 -1055 612 -1053
rect 611 -1061 612 -1059
rect 618 -1055 619 -1053
rect 618 -1061 619 -1059
rect 628 -1055 629 -1053
rect 628 -1061 629 -1059
rect 632 -1055 633 -1053
rect 632 -1061 633 -1059
rect 639 -1055 640 -1053
rect 639 -1061 640 -1059
rect 646 -1055 647 -1053
rect 649 -1055 650 -1053
rect 646 -1061 647 -1059
rect 649 -1061 650 -1059
rect 653 -1055 654 -1053
rect 653 -1061 654 -1059
rect 660 -1055 661 -1053
rect 660 -1061 661 -1059
rect 667 -1055 668 -1053
rect 667 -1061 668 -1059
rect 674 -1055 675 -1053
rect 674 -1061 675 -1059
rect 681 -1055 682 -1053
rect 681 -1061 682 -1059
rect 691 -1055 692 -1053
rect 688 -1061 689 -1059
rect 695 -1055 696 -1053
rect 695 -1061 696 -1059
rect 702 -1055 703 -1053
rect 702 -1061 703 -1059
rect 709 -1055 710 -1053
rect 709 -1061 710 -1059
rect 716 -1055 717 -1053
rect 716 -1061 717 -1059
rect 723 -1055 724 -1053
rect 723 -1061 724 -1059
rect 730 -1055 731 -1053
rect 733 -1055 734 -1053
rect 730 -1061 731 -1059
rect 737 -1055 738 -1053
rect 737 -1061 738 -1059
rect 744 -1055 745 -1053
rect 744 -1061 745 -1059
rect 751 -1055 752 -1053
rect 751 -1061 752 -1059
rect 758 -1055 759 -1053
rect 758 -1061 759 -1059
rect 765 -1055 766 -1053
rect 765 -1061 766 -1059
rect 772 -1055 773 -1053
rect 772 -1061 773 -1059
rect 779 -1055 780 -1053
rect 779 -1061 780 -1059
rect 786 -1055 787 -1053
rect 786 -1061 787 -1059
rect 793 -1055 794 -1053
rect 793 -1061 794 -1059
rect 800 -1055 801 -1053
rect 800 -1061 801 -1059
rect 807 -1055 808 -1053
rect 807 -1061 808 -1059
rect 814 -1055 815 -1053
rect 814 -1061 815 -1059
rect 821 -1055 822 -1053
rect 821 -1061 822 -1059
rect 828 -1055 829 -1053
rect 828 -1061 829 -1059
rect 835 -1055 836 -1053
rect 835 -1061 836 -1059
rect 842 -1055 843 -1053
rect 842 -1061 843 -1059
rect 849 -1055 850 -1053
rect 849 -1061 850 -1059
rect 856 -1055 857 -1053
rect 856 -1061 857 -1059
rect 863 -1055 864 -1053
rect 863 -1061 864 -1059
rect 870 -1055 871 -1053
rect 870 -1061 871 -1059
rect 877 -1055 878 -1053
rect 877 -1061 878 -1059
rect 884 -1055 885 -1053
rect 884 -1061 885 -1059
rect 891 -1055 892 -1053
rect 891 -1061 892 -1059
rect 898 -1055 899 -1053
rect 898 -1061 899 -1059
rect 905 -1055 906 -1053
rect 905 -1061 906 -1059
rect 912 -1055 913 -1053
rect 912 -1061 913 -1059
rect 919 -1055 920 -1053
rect 919 -1061 920 -1059
rect 926 -1055 927 -1053
rect 926 -1061 927 -1059
rect 933 -1055 934 -1053
rect 933 -1061 934 -1059
rect 940 -1055 941 -1053
rect 940 -1061 941 -1059
rect 947 -1055 948 -1053
rect 947 -1061 948 -1059
rect 954 -1055 955 -1053
rect 954 -1061 955 -1059
rect 961 -1055 962 -1053
rect 961 -1061 962 -1059
rect 968 -1055 969 -1053
rect 968 -1061 969 -1059
rect 975 -1055 976 -1053
rect 975 -1061 976 -1059
rect 982 -1055 983 -1053
rect 982 -1061 983 -1059
rect 989 -1055 990 -1053
rect 989 -1061 990 -1059
rect 996 -1055 997 -1053
rect 996 -1061 997 -1059
rect 1003 -1055 1004 -1053
rect 1003 -1061 1004 -1059
rect 1010 -1055 1011 -1053
rect 1010 -1061 1011 -1059
rect 1017 -1055 1018 -1053
rect 1017 -1061 1018 -1059
rect 1027 -1061 1028 -1059
rect 1031 -1055 1032 -1053
rect 1031 -1061 1032 -1059
rect 1038 -1055 1039 -1053
rect 1038 -1061 1039 -1059
rect 1045 -1055 1046 -1053
rect 1045 -1061 1046 -1059
rect 1052 -1055 1053 -1053
rect 1052 -1061 1053 -1059
rect 1059 -1055 1060 -1053
rect 1059 -1061 1060 -1059
rect 1066 -1055 1067 -1053
rect 1069 -1055 1070 -1053
rect 1069 -1061 1070 -1059
rect 1073 -1055 1074 -1053
rect 1076 -1055 1077 -1053
rect 1076 -1061 1077 -1059
rect 1080 -1061 1081 -1059
rect 1083 -1061 1084 -1059
rect 1087 -1055 1088 -1053
rect 1087 -1061 1088 -1059
rect 1094 -1055 1095 -1053
rect 1094 -1061 1095 -1059
rect 1097 -1061 1098 -1059
rect 1101 -1055 1102 -1053
rect 1101 -1061 1102 -1059
rect 2 -1154 3 -1152
rect 2 -1160 3 -1158
rect 9 -1160 10 -1158
rect 19 -1154 20 -1152
rect 23 -1154 24 -1152
rect 23 -1160 24 -1158
rect 30 -1160 31 -1158
rect 33 -1160 34 -1158
rect 37 -1154 38 -1152
rect 37 -1160 38 -1158
rect 44 -1154 45 -1152
rect 44 -1160 45 -1158
rect 51 -1154 52 -1152
rect 51 -1160 52 -1158
rect 58 -1154 59 -1152
rect 58 -1160 59 -1158
rect 65 -1154 66 -1152
rect 65 -1160 66 -1158
rect 72 -1154 73 -1152
rect 72 -1160 73 -1158
rect 79 -1160 80 -1158
rect 82 -1160 83 -1158
rect 86 -1154 87 -1152
rect 86 -1160 87 -1158
rect 93 -1154 94 -1152
rect 93 -1160 94 -1158
rect 100 -1154 101 -1152
rect 100 -1160 101 -1158
rect 107 -1154 108 -1152
rect 107 -1160 108 -1158
rect 114 -1154 115 -1152
rect 114 -1160 115 -1158
rect 121 -1154 122 -1152
rect 121 -1160 122 -1158
rect 128 -1154 129 -1152
rect 131 -1154 132 -1152
rect 128 -1160 129 -1158
rect 135 -1154 136 -1152
rect 135 -1160 136 -1158
rect 145 -1154 146 -1152
rect 142 -1160 143 -1158
rect 149 -1154 150 -1152
rect 149 -1160 150 -1158
rect 156 -1154 157 -1152
rect 156 -1160 157 -1158
rect 163 -1154 164 -1152
rect 163 -1160 164 -1158
rect 170 -1154 171 -1152
rect 170 -1160 171 -1158
rect 177 -1154 178 -1152
rect 177 -1160 178 -1158
rect 187 -1154 188 -1152
rect 184 -1160 185 -1158
rect 187 -1160 188 -1158
rect 191 -1154 192 -1152
rect 191 -1160 192 -1158
rect 198 -1154 199 -1152
rect 198 -1160 199 -1158
rect 205 -1154 206 -1152
rect 205 -1160 206 -1158
rect 212 -1160 213 -1158
rect 219 -1154 220 -1152
rect 219 -1160 220 -1158
rect 226 -1154 227 -1152
rect 229 -1154 230 -1152
rect 226 -1160 227 -1158
rect 229 -1160 230 -1158
rect 236 -1154 237 -1152
rect 233 -1160 234 -1158
rect 236 -1160 237 -1158
rect 240 -1154 241 -1152
rect 243 -1154 244 -1152
rect 240 -1160 241 -1158
rect 243 -1160 244 -1158
rect 247 -1154 248 -1152
rect 247 -1160 248 -1158
rect 254 -1154 255 -1152
rect 254 -1160 255 -1158
rect 261 -1154 262 -1152
rect 264 -1154 265 -1152
rect 264 -1160 265 -1158
rect 268 -1154 269 -1152
rect 268 -1160 269 -1158
rect 275 -1154 276 -1152
rect 275 -1160 276 -1158
rect 282 -1154 283 -1152
rect 282 -1160 283 -1158
rect 289 -1154 290 -1152
rect 289 -1160 290 -1158
rect 296 -1154 297 -1152
rect 296 -1160 297 -1158
rect 306 -1160 307 -1158
rect 310 -1154 311 -1152
rect 310 -1160 311 -1158
rect 317 -1154 318 -1152
rect 317 -1160 318 -1158
rect 324 -1154 325 -1152
rect 324 -1160 325 -1158
rect 334 -1154 335 -1152
rect 331 -1160 332 -1158
rect 338 -1154 339 -1152
rect 338 -1160 339 -1158
rect 345 -1154 346 -1152
rect 345 -1160 346 -1158
rect 355 -1160 356 -1158
rect 359 -1154 360 -1152
rect 359 -1160 360 -1158
rect 366 -1154 367 -1152
rect 369 -1154 370 -1152
rect 366 -1160 367 -1158
rect 373 -1154 374 -1152
rect 373 -1160 374 -1158
rect 380 -1154 381 -1152
rect 380 -1160 381 -1158
rect 387 -1154 388 -1152
rect 387 -1160 388 -1158
rect 394 -1154 395 -1152
rect 394 -1160 395 -1158
rect 401 -1154 402 -1152
rect 401 -1160 402 -1158
rect 408 -1154 409 -1152
rect 408 -1160 409 -1158
rect 415 -1154 416 -1152
rect 415 -1160 416 -1158
rect 422 -1154 423 -1152
rect 422 -1160 423 -1158
rect 429 -1154 430 -1152
rect 429 -1160 430 -1158
rect 436 -1154 437 -1152
rect 439 -1154 440 -1152
rect 436 -1160 437 -1158
rect 439 -1160 440 -1158
rect 443 -1154 444 -1152
rect 446 -1154 447 -1152
rect 443 -1160 444 -1158
rect 446 -1160 447 -1158
rect 450 -1154 451 -1152
rect 450 -1160 451 -1158
rect 457 -1154 458 -1152
rect 457 -1160 458 -1158
rect 467 -1154 468 -1152
rect 464 -1160 465 -1158
rect 467 -1160 468 -1158
rect 474 -1154 475 -1152
rect 471 -1160 472 -1158
rect 474 -1160 475 -1158
rect 478 -1154 479 -1152
rect 478 -1160 479 -1158
rect 485 -1154 486 -1152
rect 485 -1160 486 -1158
rect 492 -1154 493 -1152
rect 495 -1154 496 -1152
rect 495 -1160 496 -1158
rect 499 -1154 500 -1152
rect 499 -1160 500 -1158
rect 506 -1154 507 -1152
rect 509 -1154 510 -1152
rect 509 -1160 510 -1158
rect 513 -1154 514 -1152
rect 513 -1160 514 -1158
rect 520 -1154 521 -1152
rect 520 -1160 521 -1158
rect 530 -1154 531 -1152
rect 530 -1160 531 -1158
rect 534 -1154 535 -1152
rect 534 -1160 535 -1158
rect 541 -1154 542 -1152
rect 541 -1160 542 -1158
rect 548 -1154 549 -1152
rect 548 -1160 549 -1158
rect 555 -1154 556 -1152
rect 555 -1160 556 -1158
rect 562 -1154 563 -1152
rect 562 -1160 563 -1158
rect 569 -1154 570 -1152
rect 569 -1160 570 -1158
rect 576 -1154 577 -1152
rect 576 -1160 577 -1158
rect 583 -1154 584 -1152
rect 586 -1154 587 -1152
rect 583 -1160 584 -1158
rect 586 -1160 587 -1158
rect 590 -1154 591 -1152
rect 593 -1154 594 -1152
rect 590 -1160 591 -1158
rect 593 -1160 594 -1158
rect 597 -1154 598 -1152
rect 600 -1154 601 -1152
rect 597 -1160 598 -1158
rect 600 -1160 601 -1158
rect 604 -1154 605 -1152
rect 607 -1154 608 -1152
rect 604 -1160 605 -1158
rect 611 -1154 612 -1152
rect 611 -1160 612 -1158
rect 621 -1154 622 -1152
rect 618 -1160 619 -1158
rect 621 -1160 622 -1158
rect 628 -1154 629 -1152
rect 625 -1160 626 -1158
rect 628 -1160 629 -1158
rect 632 -1154 633 -1152
rect 632 -1160 633 -1158
rect 642 -1154 643 -1152
rect 639 -1160 640 -1158
rect 642 -1160 643 -1158
rect 646 -1154 647 -1152
rect 646 -1160 647 -1158
rect 653 -1154 654 -1152
rect 653 -1160 654 -1158
rect 660 -1154 661 -1152
rect 660 -1160 661 -1158
rect 663 -1160 664 -1158
rect 667 -1154 668 -1152
rect 667 -1160 668 -1158
rect 674 -1154 675 -1152
rect 677 -1154 678 -1152
rect 677 -1160 678 -1158
rect 681 -1154 682 -1152
rect 681 -1160 682 -1158
rect 688 -1154 689 -1152
rect 691 -1160 692 -1158
rect 695 -1154 696 -1152
rect 695 -1160 696 -1158
rect 702 -1154 703 -1152
rect 702 -1160 703 -1158
rect 709 -1154 710 -1152
rect 709 -1160 710 -1158
rect 716 -1154 717 -1152
rect 716 -1160 717 -1158
rect 723 -1154 724 -1152
rect 726 -1154 727 -1152
rect 723 -1160 724 -1158
rect 730 -1154 731 -1152
rect 733 -1160 734 -1158
rect 737 -1154 738 -1152
rect 737 -1160 738 -1158
rect 744 -1154 745 -1152
rect 744 -1160 745 -1158
rect 751 -1154 752 -1152
rect 751 -1160 752 -1158
rect 758 -1154 759 -1152
rect 758 -1160 759 -1158
rect 765 -1154 766 -1152
rect 765 -1160 766 -1158
rect 772 -1154 773 -1152
rect 772 -1160 773 -1158
rect 779 -1154 780 -1152
rect 779 -1160 780 -1158
rect 786 -1154 787 -1152
rect 786 -1160 787 -1158
rect 793 -1154 794 -1152
rect 793 -1160 794 -1158
rect 800 -1154 801 -1152
rect 800 -1160 801 -1158
rect 807 -1154 808 -1152
rect 807 -1160 808 -1158
rect 814 -1154 815 -1152
rect 814 -1160 815 -1158
rect 821 -1154 822 -1152
rect 821 -1160 822 -1158
rect 828 -1154 829 -1152
rect 828 -1160 829 -1158
rect 835 -1154 836 -1152
rect 835 -1160 836 -1158
rect 842 -1154 843 -1152
rect 842 -1160 843 -1158
rect 849 -1154 850 -1152
rect 849 -1160 850 -1158
rect 856 -1154 857 -1152
rect 856 -1160 857 -1158
rect 863 -1154 864 -1152
rect 863 -1160 864 -1158
rect 870 -1154 871 -1152
rect 870 -1160 871 -1158
rect 877 -1154 878 -1152
rect 877 -1160 878 -1158
rect 884 -1154 885 -1152
rect 884 -1160 885 -1158
rect 891 -1154 892 -1152
rect 891 -1160 892 -1158
rect 898 -1154 899 -1152
rect 898 -1160 899 -1158
rect 905 -1154 906 -1152
rect 905 -1160 906 -1158
rect 912 -1154 913 -1152
rect 912 -1160 913 -1158
rect 919 -1154 920 -1152
rect 919 -1160 920 -1158
rect 926 -1154 927 -1152
rect 926 -1160 927 -1158
rect 933 -1154 934 -1152
rect 933 -1160 934 -1158
rect 940 -1154 941 -1152
rect 940 -1160 941 -1158
rect 947 -1154 948 -1152
rect 947 -1160 948 -1158
rect 954 -1154 955 -1152
rect 954 -1160 955 -1158
rect 961 -1154 962 -1152
rect 961 -1160 962 -1158
rect 968 -1154 969 -1152
rect 968 -1160 969 -1158
rect 975 -1154 976 -1152
rect 975 -1160 976 -1158
rect 982 -1154 983 -1152
rect 982 -1160 983 -1158
rect 989 -1154 990 -1152
rect 989 -1160 990 -1158
rect 996 -1154 997 -1152
rect 996 -1160 997 -1158
rect 1003 -1154 1004 -1152
rect 1003 -1160 1004 -1158
rect 1010 -1154 1011 -1152
rect 1010 -1160 1011 -1158
rect 1017 -1154 1018 -1152
rect 1017 -1160 1018 -1158
rect 1024 -1154 1025 -1152
rect 1024 -1160 1025 -1158
rect 1031 -1154 1032 -1152
rect 1031 -1160 1032 -1158
rect 1038 -1154 1039 -1152
rect 1038 -1160 1039 -1158
rect 1045 -1154 1046 -1152
rect 1045 -1160 1046 -1158
rect 1052 -1154 1053 -1152
rect 1052 -1160 1053 -1158
rect 1059 -1154 1060 -1152
rect 1059 -1160 1060 -1158
rect 1066 -1154 1067 -1152
rect 1066 -1160 1067 -1158
rect 1073 -1154 1074 -1152
rect 1073 -1160 1074 -1158
rect 1080 -1154 1081 -1152
rect 1080 -1160 1081 -1158
rect 1087 -1154 1088 -1152
rect 1087 -1160 1088 -1158
rect 1090 -1160 1091 -1158
rect 1094 -1154 1095 -1152
rect 1097 -1154 1098 -1152
rect 1094 -1160 1095 -1158
rect 1101 -1154 1102 -1152
rect 1101 -1160 1102 -1158
rect 2 -1257 3 -1255
rect 2 -1263 3 -1261
rect 9 -1257 10 -1255
rect 9 -1263 10 -1261
rect 16 -1257 17 -1255
rect 23 -1257 24 -1255
rect 26 -1257 27 -1255
rect 23 -1263 24 -1261
rect 30 -1257 31 -1255
rect 30 -1263 31 -1261
rect 37 -1257 38 -1255
rect 37 -1263 38 -1261
rect 44 -1257 45 -1255
rect 44 -1263 45 -1261
rect 51 -1257 52 -1255
rect 51 -1263 52 -1261
rect 54 -1263 55 -1261
rect 58 -1257 59 -1255
rect 58 -1263 59 -1261
rect 65 -1257 66 -1255
rect 65 -1263 66 -1261
rect 72 -1257 73 -1255
rect 72 -1263 73 -1261
rect 79 -1257 80 -1255
rect 82 -1257 83 -1255
rect 86 -1257 87 -1255
rect 86 -1263 87 -1261
rect 93 -1257 94 -1255
rect 93 -1263 94 -1261
rect 100 -1257 101 -1255
rect 100 -1263 101 -1261
rect 107 -1257 108 -1255
rect 107 -1263 108 -1261
rect 114 -1257 115 -1255
rect 117 -1257 118 -1255
rect 114 -1263 115 -1261
rect 117 -1263 118 -1261
rect 121 -1257 122 -1255
rect 121 -1263 122 -1261
rect 128 -1257 129 -1255
rect 128 -1263 129 -1261
rect 135 -1257 136 -1255
rect 135 -1263 136 -1261
rect 142 -1257 143 -1255
rect 142 -1263 143 -1261
rect 149 -1257 150 -1255
rect 149 -1263 150 -1261
rect 156 -1257 157 -1255
rect 156 -1263 157 -1261
rect 163 -1257 164 -1255
rect 166 -1257 167 -1255
rect 163 -1263 164 -1261
rect 166 -1263 167 -1261
rect 170 -1257 171 -1255
rect 170 -1263 171 -1261
rect 177 -1257 178 -1255
rect 177 -1263 178 -1261
rect 184 -1257 185 -1255
rect 187 -1257 188 -1255
rect 184 -1263 185 -1261
rect 187 -1263 188 -1261
rect 191 -1257 192 -1255
rect 194 -1257 195 -1255
rect 194 -1263 195 -1261
rect 198 -1257 199 -1255
rect 201 -1263 202 -1261
rect 205 -1257 206 -1255
rect 205 -1263 206 -1261
rect 215 -1257 216 -1255
rect 212 -1263 213 -1261
rect 215 -1263 216 -1261
rect 219 -1257 220 -1255
rect 219 -1263 220 -1261
rect 222 -1263 223 -1261
rect 226 -1257 227 -1255
rect 226 -1263 227 -1261
rect 233 -1257 234 -1255
rect 233 -1263 234 -1261
rect 240 -1257 241 -1255
rect 240 -1263 241 -1261
rect 247 -1257 248 -1255
rect 247 -1263 248 -1261
rect 254 -1257 255 -1255
rect 254 -1263 255 -1261
rect 261 -1257 262 -1255
rect 261 -1263 262 -1261
rect 268 -1257 269 -1255
rect 268 -1263 269 -1261
rect 275 -1257 276 -1255
rect 275 -1263 276 -1261
rect 282 -1257 283 -1255
rect 282 -1263 283 -1261
rect 289 -1257 290 -1255
rect 292 -1257 293 -1255
rect 289 -1263 290 -1261
rect 292 -1263 293 -1261
rect 296 -1257 297 -1255
rect 296 -1263 297 -1261
rect 303 -1257 304 -1255
rect 303 -1263 304 -1261
rect 310 -1257 311 -1255
rect 310 -1263 311 -1261
rect 317 -1257 318 -1255
rect 317 -1263 318 -1261
rect 324 -1257 325 -1255
rect 324 -1263 325 -1261
rect 331 -1257 332 -1255
rect 331 -1263 332 -1261
rect 338 -1257 339 -1255
rect 338 -1263 339 -1261
rect 345 -1257 346 -1255
rect 345 -1263 346 -1261
rect 352 -1257 353 -1255
rect 352 -1263 353 -1261
rect 359 -1257 360 -1255
rect 359 -1263 360 -1261
rect 366 -1257 367 -1255
rect 366 -1263 367 -1261
rect 373 -1257 374 -1255
rect 373 -1263 374 -1261
rect 380 -1257 381 -1255
rect 380 -1263 381 -1261
rect 387 -1257 388 -1255
rect 387 -1263 388 -1261
rect 394 -1257 395 -1255
rect 394 -1263 395 -1261
rect 401 -1257 402 -1255
rect 401 -1263 402 -1261
rect 408 -1257 409 -1255
rect 408 -1263 409 -1261
rect 415 -1257 416 -1255
rect 415 -1263 416 -1261
rect 422 -1257 423 -1255
rect 422 -1263 423 -1261
rect 425 -1263 426 -1261
rect 429 -1257 430 -1255
rect 432 -1263 433 -1261
rect 436 -1257 437 -1255
rect 436 -1263 437 -1261
rect 443 -1257 444 -1255
rect 443 -1263 444 -1261
rect 450 -1257 451 -1255
rect 450 -1263 451 -1261
rect 457 -1257 458 -1255
rect 460 -1257 461 -1255
rect 457 -1263 458 -1261
rect 464 -1257 465 -1255
rect 464 -1263 465 -1261
rect 471 -1257 472 -1255
rect 474 -1257 475 -1255
rect 471 -1263 472 -1261
rect 478 -1257 479 -1255
rect 478 -1263 479 -1261
rect 485 -1257 486 -1255
rect 485 -1263 486 -1261
rect 492 -1257 493 -1255
rect 495 -1257 496 -1255
rect 492 -1263 493 -1261
rect 495 -1263 496 -1261
rect 499 -1257 500 -1255
rect 502 -1257 503 -1255
rect 499 -1263 500 -1261
rect 502 -1263 503 -1261
rect 506 -1257 507 -1255
rect 506 -1263 507 -1261
rect 513 -1257 514 -1255
rect 516 -1257 517 -1255
rect 513 -1263 514 -1261
rect 516 -1263 517 -1261
rect 523 -1257 524 -1255
rect 520 -1263 521 -1261
rect 527 -1257 528 -1255
rect 527 -1263 528 -1261
rect 537 -1263 538 -1261
rect 541 -1257 542 -1255
rect 544 -1257 545 -1255
rect 541 -1263 542 -1261
rect 544 -1263 545 -1261
rect 548 -1257 549 -1255
rect 551 -1257 552 -1255
rect 548 -1263 549 -1261
rect 555 -1257 556 -1255
rect 555 -1263 556 -1261
rect 562 -1257 563 -1255
rect 565 -1257 566 -1255
rect 562 -1263 563 -1261
rect 565 -1263 566 -1261
rect 569 -1257 570 -1255
rect 569 -1263 570 -1261
rect 576 -1257 577 -1255
rect 576 -1263 577 -1261
rect 586 -1257 587 -1255
rect 583 -1263 584 -1261
rect 586 -1263 587 -1261
rect 590 -1257 591 -1255
rect 597 -1257 598 -1255
rect 597 -1263 598 -1261
rect 604 -1257 605 -1255
rect 607 -1257 608 -1255
rect 604 -1263 605 -1261
rect 607 -1263 608 -1261
rect 611 -1257 612 -1255
rect 611 -1263 612 -1261
rect 618 -1257 619 -1255
rect 618 -1263 619 -1261
rect 625 -1257 626 -1255
rect 625 -1263 626 -1261
rect 632 -1257 633 -1255
rect 632 -1263 633 -1261
rect 639 -1257 640 -1255
rect 639 -1263 640 -1261
rect 646 -1257 647 -1255
rect 646 -1263 647 -1261
rect 656 -1257 657 -1255
rect 653 -1263 654 -1261
rect 656 -1263 657 -1261
rect 660 -1257 661 -1255
rect 660 -1263 661 -1261
rect 667 -1257 668 -1255
rect 667 -1263 668 -1261
rect 674 -1257 675 -1255
rect 674 -1263 675 -1261
rect 681 -1257 682 -1255
rect 684 -1257 685 -1255
rect 688 -1257 689 -1255
rect 688 -1263 689 -1261
rect 695 -1257 696 -1255
rect 695 -1263 696 -1261
rect 702 -1257 703 -1255
rect 702 -1263 703 -1261
rect 709 -1257 710 -1255
rect 709 -1263 710 -1261
rect 716 -1257 717 -1255
rect 719 -1257 720 -1255
rect 716 -1263 717 -1261
rect 723 -1257 724 -1255
rect 723 -1263 724 -1261
rect 730 -1257 731 -1255
rect 730 -1263 731 -1261
rect 737 -1257 738 -1255
rect 737 -1263 738 -1261
rect 744 -1257 745 -1255
rect 744 -1263 745 -1261
rect 751 -1257 752 -1255
rect 751 -1263 752 -1261
rect 758 -1257 759 -1255
rect 758 -1263 759 -1261
rect 765 -1257 766 -1255
rect 765 -1263 766 -1261
rect 772 -1257 773 -1255
rect 772 -1263 773 -1261
rect 779 -1257 780 -1255
rect 782 -1257 783 -1255
rect 786 -1257 787 -1255
rect 786 -1263 787 -1261
rect 793 -1257 794 -1255
rect 793 -1263 794 -1261
rect 800 -1257 801 -1255
rect 800 -1263 801 -1261
rect 807 -1257 808 -1255
rect 807 -1263 808 -1261
rect 814 -1257 815 -1255
rect 817 -1263 818 -1261
rect 821 -1257 822 -1255
rect 821 -1263 822 -1261
rect 828 -1257 829 -1255
rect 828 -1263 829 -1261
rect 835 -1257 836 -1255
rect 835 -1263 836 -1261
rect 842 -1257 843 -1255
rect 842 -1263 843 -1261
rect 849 -1257 850 -1255
rect 849 -1263 850 -1261
rect 856 -1257 857 -1255
rect 856 -1263 857 -1261
rect 863 -1257 864 -1255
rect 863 -1263 864 -1261
rect 870 -1257 871 -1255
rect 870 -1263 871 -1261
rect 877 -1257 878 -1255
rect 877 -1263 878 -1261
rect 884 -1257 885 -1255
rect 884 -1263 885 -1261
rect 891 -1257 892 -1255
rect 891 -1263 892 -1261
rect 898 -1257 899 -1255
rect 898 -1263 899 -1261
rect 905 -1257 906 -1255
rect 905 -1263 906 -1261
rect 912 -1257 913 -1255
rect 912 -1263 913 -1261
rect 919 -1257 920 -1255
rect 919 -1263 920 -1261
rect 926 -1257 927 -1255
rect 933 -1257 934 -1255
rect 933 -1263 934 -1261
rect 940 -1257 941 -1255
rect 940 -1263 941 -1261
rect 947 -1257 948 -1255
rect 947 -1263 948 -1261
rect 954 -1257 955 -1255
rect 954 -1263 955 -1261
rect 961 -1257 962 -1255
rect 961 -1263 962 -1261
rect 968 -1257 969 -1255
rect 968 -1263 969 -1261
rect 975 -1257 976 -1255
rect 975 -1263 976 -1261
rect 982 -1257 983 -1255
rect 982 -1263 983 -1261
rect 989 -1257 990 -1255
rect 989 -1263 990 -1261
rect 996 -1257 997 -1255
rect 996 -1263 997 -1261
rect 1003 -1257 1004 -1255
rect 1003 -1263 1004 -1261
rect 1010 -1257 1011 -1255
rect 1010 -1263 1011 -1261
rect 1017 -1257 1018 -1255
rect 1017 -1263 1018 -1261
rect 1020 -1263 1021 -1261
rect 1024 -1257 1025 -1255
rect 1024 -1263 1025 -1261
rect 1031 -1257 1032 -1255
rect 1038 -1257 1039 -1255
rect 1041 -1257 1042 -1255
rect 1041 -1263 1042 -1261
rect 1045 -1257 1046 -1255
rect 1045 -1263 1046 -1261
rect 1052 -1257 1053 -1255
rect 1052 -1263 1053 -1261
rect 1059 -1257 1060 -1255
rect 1059 -1263 1060 -1261
rect 1066 -1257 1067 -1255
rect 1066 -1263 1067 -1261
rect 1073 -1257 1074 -1255
rect 1073 -1263 1074 -1261
rect 9 -1336 10 -1334
rect 9 -1342 10 -1340
rect 16 -1336 17 -1334
rect 16 -1342 17 -1340
rect 23 -1336 24 -1334
rect 23 -1342 24 -1340
rect 30 -1336 31 -1334
rect 30 -1342 31 -1340
rect 37 -1336 38 -1334
rect 37 -1342 38 -1340
rect 44 -1336 45 -1334
rect 44 -1342 45 -1340
rect 51 -1336 52 -1334
rect 51 -1342 52 -1340
rect 58 -1336 59 -1334
rect 58 -1342 59 -1340
rect 65 -1336 66 -1334
rect 65 -1342 66 -1340
rect 72 -1336 73 -1334
rect 72 -1342 73 -1340
rect 79 -1342 80 -1340
rect 86 -1336 87 -1334
rect 86 -1342 87 -1340
rect 93 -1336 94 -1334
rect 93 -1342 94 -1340
rect 100 -1336 101 -1334
rect 100 -1342 101 -1340
rect 107 -1336 108 -1334
rect 107 -1342 108 -1340
rect 117 -1336 118 -1334
rect 121 -1336 122 -1334
rect 121 -1342 122 -1340
rect 131 -1336 132 -1334
rect 128 -1342 129 -1340
rect 138 -1336 139 -1334
rect 138 -1342 139 -1340
rect 142 -1336 143 -1334
rect 142 -1342 143 -1340
rect 149 -1336 150 -1334
rect 149 -1342 150 -1340
rect 159 -1336 160 -1334
rect 159 -1342 160 -1340
rect 163 -1336 164 -1334
rect 163 -1342 164 -1340
rect 170 -1336 171 -1334
rect 173 -1336 174 -1334
rect 173 -1342 174 -1340
rect 177 -1342 178 -1340
rect 180 -1342 181 -1340
rect 184 -1336 185 -1334
rect 184 -1342 185 -1340
rect 191 -1336 192 -1334
rect 194 -1336 195 -1334
rect 194 -1342 195 -1340
rect 198 -1336 199 -1334
rect 198 -1342 199 -1340
rect 205 -1336 206 -1334
rect 205 -1342 206 -1340
rect 212 -1336 213 -1334
rect 212 -1342 213 -1340
rect 219 -1336 220 -1334
rect 222 -1336 223 -1334
rect 219 -1342 220 -1340
rect 222 -1342 223 -1340
rect 226 -1336 227 -1334
rect 226 -1342 227 -1340
rect 233 -1336 234 -1334
rect 233 -1342 234 -1340
rect 240 -1336 241 -1334
rect 240 -1342 241 -1340
rect 247 -1336 248 -1334
rect 247 -1342 248 -1340
rect 254 -1336 255 -1334
rect 254 -1342 255 -1340
rect 261 -1336 262 -1334
rect 261 -1342 262 -1340
rect 268 -1336 269 -1334
rect 268 -1342 269 -1340
rect 275 -1336 276 -1334
rect 275 -1342 276 -1340
rect 282 -1336 283 -1334
rect 282 -1342 283 -1340
rect 292 -1336 293 -1334
rect 292 -1342 293 -1340
rect 296 -1336 297 -1334
rect 296 -1342 297 -1340
rect 303 -1336 304 -1334
rect 303 -1342 304 -1340
rect 310 -1336 311 -1334
rect 310 -1342 311 -1340
rect 317 -1336 318 -1334
rect 320 -1336 321 -1334
rect 317 -1342 318 -1340
rect 327 -1336 328 -1334
rect 324 -1342 325 -1340
rect 327 -1342 328 -1340
rect 331 -1336 332 -1334
rect 331 -1342 332 -1340
rect 338 -1336 339 -1334
rect 338 -1342 339 -1340
rect 345 -1336 346 -1334
rect 345 -1342 346 -1340
rect 352 -1336 353 -1334
rect 355 -1336 356 -1334
rect 352 -1342 353 -1340
rect 355 -1342 356 -1340
rect 359 -1336 360 -1334
rect 359 -1342 360 -1340
rect 366 -1336 367 -1334
rect 369 -1336 370 -1334
rect 369 -1342 370 -1340
rect 373 -1336 374 -1334
rect 373 -1342 374 -1340
rect 380 -1336 381 -1334
rect 380 -1342 381 -1340
rect 387 -1336 388 -1334
rect 387 -1342 388 -1340
rect 394 -1336 395 -1334
rect 394 -1342 395 -1340
rect 401 -1336 402 -1334
rect 401 -1342 402 -1340
rect 408 -1336 409 -1334
rect 408 -1342 409 -1340
rect 415 -1336 416 -1334
rect 415 -1342 416 -1340
rect 422 -1336 423 -1334
rect 422 -1342 423 -1340
rect 432 -1336 433 -1334
rect 429 -1342 430 -1340
rect 432 -1342 433 -1340
rect 436 -1336 437 -1334
rect 436 -1342 437 -1340
rect 443 -1336 444 -1334
rect 443 -1342 444 -1340
rect 450 -1336 451 -1334
rect 450 -1342 451 -1340
rect 457 -1336 458 -1334
rect 460 -1336 461 -1334
rect 460 -1342 461 -1340
rect 464 -1336 465 -1334
rect 464 -1342 465 -1340
rect 474 -1336 475 -1334
rect 471 -1342 472 -1340
rect 478 -1336 479 -1334
rect 478 -1342 479 -1340
rect 485 -1336 486 -1334
rect 485 -1342 486 -1340
rect 492 -1336 493 -1334
rect 492 -1342 493 -1340
rect 495 -1342 496 -1340
rect 499 -1336 500 -1334
rect 499 -1342 500 -1340
rect 509 -1336 510 -1334
rect 506 -1342 507 -1340
rect 513 -1336 514 -1334
rect 513 -1342 514 -1340
rect 520 -1336 521 -1334
rect 520 -1342 521 -1340
rect 527 -1336 528 -1334
rect 527 -1342 528 -1340
rect 534 -1336 535 -1334
rect 537 -1336 538 -1334
rect 541 -1336 542 -1334
rect 541 -1342 542 -1340
rect 548 -1336 549 -1334
rect 548 -1342 549 -1340
rect 555 -1336 556 -1334
rect 555 -1342 556 -1340
rect 562 -1336 563 -1334
rect 562 -1342 563 -1340
rect 569 -1336 570 -1334
rect 569 -1342 570 -1340
rect 576 -1336 577 -1334
rect 579 -1336 580 -1334
rect 576 -1342 577 -1340
rect 579 -1342 580 -1340
rect 583 -1336 584 -1334
rect 583 -1342 584 -1340
rect 590 -1336 591 -1334
rect 590 -1342 591 -1340
rect 597 -1336 598 -1334
rect 597 -1342 598 -1340
rect 600 -1342 601 -1340
rect 604 -1336 605 -1334
rect 604 -1342 605 -1340
rect 611 -1336 612 -1334
rect 611 -1342 612 -1340
rect 621 -1336 622 -1334
rect 618 -1342 619 -1340
rect 625 -1336 626 -1334
rect 625 -1342 626 -1340
rect 632 -1336 633 -1334
rect 632 -1342 633 -1340
rect 639 -1336 640 -1334
rect 639 -1342 640 -1340
rect 646 -1336 647 -1334
rect 646 -1342 647 -1340
rect 649 -1342 650 -1340
rect 653 -1336 654 -1334
rect 653 -1342 654 -1340
rect 660 -1336 661 -1334
rect 660 -1342 661 -1340
rect 667 -1336 668 -1334
rect 667 -1342 668 -1340
rect 677 -1336 678 -1334
rect 674 -1342 675 -1340
rect 677 -1342 678 -1340
rect 681 -1336 682 -1334
rect 681 -1342 682 -1340
rect 688 -1336 689 -1334
rect 688 -1342 689 -1340
rect 695 -1336 696 -1334
rect 695 -1342 696 -1340
rect 702 -1342 703 -1340
rect 705 -1342 706 -1340
rect 709 -1336 710 -1334
rect 709 -1342 710 -1340
rect 716 -1336 717 -1334
rect 716 -1342 717 -1340
rect 723 -1336 724 -1334
rect 723 -1342 724 -1340
rect 730 -1336 731 -1334
rect 730 -1342 731 -1340
rect 737 -1342 738 -1340
rect 744 -1336 745 -1334
rect 744 -1342 745 -1340
rect 751 -1336 752 -1334
rect 751 -1342 752 -1340
rect 758 -1336 759 -1334
rect 761 -1336 762 -1334
rect 758 -1342 759 -1340
rect 765 -1336 766 -1334
rect 765 -1342 766 -1340
rect 772 -1336 773 -1334
rect 772 -1342 773 -1340
rect 779 -1336 780 -1334
rect 779 -1342 780 -1340
rect 786 -1336 787 -1334
rect 786 -1342 787 -1340
rect 793 -1336 794 -1334
rect 793 -1342 794 -1340
rect 800 -1336 801 -1334
rect 800 -1342 801 -1340
rect 807 -1336 808 -1334
rect 807 -1342 808 -1340
rect 814 -1336 815 -1334
rect 814 -1342 815 -1340
rect 821 -1336 822 -1334
rect 821 -1342 822 -1340
rect 828 -1336 829 -1334
rect 828 -1342 829 -1340
rect 835 -1336 836 -1334
rect 835 -1342 836 -1340
rect 842 -1336 843 -1334
rect 842 -1342 843 -1340
rect 849 -1336 850 -1334
rect 849 -1342 850 -1340
rect 856 -1336 857 -1334
rect 856 -1342 857 -1340
rect 863 -1336 864 -1334
rect 863 -1342 864 -1340
rect 870 -1336 871 -1334
rect 870 -1342 871 -1340
rect 877 -1336 878 -1334
rect 877 -1342 878 -1340
rect 884 -1336 885 -1334
rect 884 -1342 885 -1340
rect 891 -1336 892 -1334
rect 891 -1342 892 -1340
rect 898 -1336 899 -1334
rect 898 -1342 899 -1340
rect 905 -1336 906 -1334
rect 905 -1342 906 -1340
rect 912 -1336 913 -1334
rect 912 -1342 913 -1340
rect 919 -1336 920 -1334
rect 919 -1342 920 -1340
rect 926 -1342 927 -1340
rect 933 -1336 934 -1334
rect 933 -1342 934 -1340
rect 940 -1336 941 -1334
rect 940 -1342 941 -1340
rect 947 -1336 948 -1334
rect 947 -1342 948 -1340
rect 954 -1336 955 -1334
rect 954 -1342 955 -1340
rect 961 -1336 962 -1334
rect 961 -1342 962 -1340
rect 968 -1336 969 -1334
rect 968 -1342 969 -1340
rect 975 -1336 976 -1334
rect 975 -1342 976 -1340
rect 982 -1336 983 -1334
rect 982 -1342 983 -1340
rect 989 -1336 990 -1334
rect 989 -1342 990 -1340
rect 996 -1336 997 -1334
rect 996 -1342 997 -1340
rect 1003 -1336 1004 -1334
rect 1003 -1342 1004 -1340
rect 1010 -1336 1011 -1334
rect 1010 -1342 1011 -1340
rect 1017 -1336 1018 -1334
rect 1020 -1336 1021 -1334
rect 1017 -1342 1018 -1340
rect 1024 -1342 1025 -1340
rect 1031 -1336 1032 -1334
rect 1034 -1336 1035 -1334
rect 1031 -1342 1032 -1340
rect 1034 -1342 1035 -1340
rect 1038 -1336 1039 -1334
rect 1038 -1342 1039 -1340
rect 1045 -1336 1046 -1334
rect 1048 -1336 1049 -1334
rect 1048 -1342 1049 -1340
rect 1052 -1336 1053 -1334
rect 1052 -1342 1053 -1340
rect 1059 -1336 1060 -1334
rect 1062 -1336 1063 -1334
rect 1066 -1336 1067 -1334
rect 1066 -1342 1067 -1340
rect 1073 -1336 1074 -1334
rect 1073 -1342 1074 -1340
rect 1080 -1336 1081 -1334
rect 1080 -1342 1081 -1340
rect 16 -1413 17 -1411
rect 16 -1419 17 -1417
rect 23 -1413 24 -1411
rect 23 -1419 24 -1417
rect 30 -1413 31 -1411
rect 30 -1419 31 -1417
rect 37 -1413 38 -1411
rect 37 -1419 38 -1417
rect 44 -1413 45 -1411
rect 44 -1419 45 -1417
rect 54 -1413 55 -1411
rect 51 -1419 52 -1417
rect 61 -1413 62 -1411
rect 65 -1413 66 -1411
rect 65 -1419 66 -1417
rect 72 -1413 73 -1411
rect 72 -1419 73 -1417
rect 79 -1413 80 -1411
rect 79 -1419 80 -1417
rect 86 -1413 87 -1411
rect 89 -1413 90 -1411
rect 86 -1419 87 -1417
rect 89 -1419 90 -1417
rect 93 -1413 94 -1411
rect 93 -1419 94 -1417
rect 100 -1413 101 -1411
rect 100 -1419 101 -1417
rect 107 -1413 108 -1411
rect 107 -1419 108 -1417
rect 114 -1413 115 -1411
rect 114 -1419 115 -1417
rect 121 -1413 122 -1411
rect 121 -1419 122 -1417
rect 128 -1413 129 -1411
rect 128 -1419 129 -1417
rect 135 -1413 136 -1411
rect 138 -1419 139 -1417
rect 145 -1413 146 -1411
rect 142 -1419 143 -1417
rect 149 -1413 150 -1411
rect 149 -1419 150 -1417
rect 156 -1413 157 -1411
rect 159 -1419 160 -1417
rect 163 -1413 164 -1411
rect 163 -1419 164 -1417
rect 166 -1419 167 -1417
rect 170 -1413 171 -1411
rect 170 -1419 171 -1417
rect 177 -1413 178 -1411
rect 177 -1419 178 -1417
rect 184 -1413 185 -1411
rect 184 -1419 185 -1417
rect 191 -1413 192 -1411
rect 191 -1419 192 -1417
rect 198 -1413 199 -1411
rect 198 -1419 199 -1417
rect 205 -1413 206 -1411
rect 208 -1413 209 -1411
rect 205 -1419 206 -1417
rect 212 -1413 213 -1411
rect 212 -1419 213 -1417
rect 222 -1413 223 -1411
rect 219 -1419 220 -1417
rect 222 -1419 223 -1417
rect 226 -1413 227 -1411
rect 226 -1419 227 -1417
rect 233 -1413 234 -1411
rect 233 -1419 234 -1417
rect 240 -1419 241 -1417
rect 243 -1419 244 -1417
rect 247 -1413 248 -1411
rect 247 -1419 248 -1417
rect 254 -1413 255 -1411
rect 254 -1419 255 -1417
rect 261 -1413 262 -1411
rect 261 -1419 262 -1417
rect 268 -1413 269 -1411
rect 268 -1419 269 -1417
rect 275 -1413 276 -1411
rect 275 -1419 276 -1417
rect 282 -1413 283 -1411
rect 282 -1419 283 -1417
rect 289 -1413 290 -1411
rect 289 -1419 290 -1417
rect 296 -1413 297 -1411
rect 296 -1419 297 -1417
rect 303 -1413 304 -1411
rect 303 -1419 304 -1417
rect 306 -1419 307 -1417
rect 310 -1413 311 -1411
rect 310 -1419 311 -1417
rect 317 -1413 318 -1411
rect 317 -1419 318 -1417
rect 324 -1413 325 -1411
rect 324 -1419 325 -1417
rect 331 -1413 332 -1411
rect 331 -1419 332 -1417
rect 338 -1413 339 -1411
rect 338 -1419 339 -1417
rect 345 -1413 346 -1411
rect 345 -1419 346 -1417
rect 352 -1413 353 -1411
rect 355 -1413 356 -1411
rect 355 -1419 356 -1417
rect 359 -1413 360 -1411
rect 362 -1419 363 -1417
rect 366 -1413 367 -1411
rect 366 -1419 367 -1417
rect 373 -1413 374 -1411
rect 373 -1419 374 -1417
rect 380 -1413 381 -1411
rect 380 -1419 381 -1417
rect 387 -1413 388 -1411
rect 390 -1419 391 -1417
rect 394 -1413 395 -1411
rect 394 -1419 395 -1417
rect 401 -1413 402 -1411
rect 401 -1419 402 -1417
rect 408 -1413 409 -1411
rect 411 -1413 412 -1411
rect 408 -1419 409 -1417
rect 411 -1419 412 -1417
rect 415 -1413 416 -1411
rect 415 -1419 416 -1417
rect 422 -1413 423 -1411
rect 422 -1419 423 -1417
rect 429 -1413 430 -1411
rect 429 -1419 430 -1417
rect 436 -1413 437 -1411
rect 436 -1419 437 -1417
rect 443 -1413 444 -1411
rect 443 -1419 444 -1417
rect 450 -1413 451 -1411
rect 450 -1419 451 -1417
rect 457 -1413 458 -1411
rect 457 -1419 458 -1417
rect 464 -1413 465 -1411
rect 464 -1419 465 -1417
rect 471 -1413 472 -1411
rect 471 -1419 472 -1417
rect 478 -1413 479 -1411
rect 478 -1419 479 -1417
rect 485 -1413 486 -1411
rect 485 -1419 486 -1417
rect 492 -1413 493 -1411
rect 492 -1419 493 -1417
rect 499 -1413 500 -1411
rect 499 -1419 500 -1417
rect 506 -1413 507 -1411
rect 509 -1413 510 -1411
rect 506 -1419 507 -1417
rect 516 -1413 517 -1411
rect 513 -1419 514 -1417
rect 516 -1419 517 -1417
rect 520 -1413 521 -1411
rect 523 -1413 524 -1411
rect 523 -1419 524 -1417
rect 527 -1413 528 -1411
rect 527 -1419 528 -1417
rect 534 -1413 535 -1411
rect 534 -1419 535 -1417
rect 541 -1413 542 -1411
rect 541 -1419 542 -1417
rect 548 -1413 549 -1411
rect 548 -1419 549 -1417
rect 555 -1413 556 -1411
rect 555 -1419 556 -1417
rect 565 -1413 566 -1411
rect 562 -1419 563 -1417
rect 569 -1413 570 -1411
rect 572 -1413 573 -1411
rect 569 -1419 570 -1417
rect 576 -1413 577 -1411
rect 579 -1413 580 -1411
rect 576 -1419 577 -1417
rect 583 -1413 584 -1411
rect 586 -1413 587 -1411
rect 583 -1419 584 -1417
rect 586 -1419 587 -1417
rect 590 -1413 591 -1411
rect 590 -1419 591 -1417
rect 597 -1413 598 -1411
rect 597 -1419 598 -1417
rect 604 -1413 605 -1411
rect 604 -1419 605 -1417
rect 611 -1413 612 -1411
rect 611 -1419 612 -1417
rect 618 -1413 619 -1411
rect 618 -1419 619 -1417
rect 625 -1413 626 -1411
rect 625 -1419 626 -1417
rect 632 -1413 633 -1411
rect 632 -1419 633 -1417
rect 639 -1413 640 -1411
rect 639 -1419 640 -1417
rect 646 -1413 647 -1411
rect 646 -1419 647 -1417
rect 653 -1413 654 -1411
rect 653 -1419 654 -1417
rect 660 -1413 661 -1411
rect 663 -1413 664 -1411
rect 660 -1419 661 -1417
rect 663 -1419 664 -1417
rect 667 -1413 668 -1411
rect 667 -1419 668 -1417
rect 674 -1413 675 -1411
rect 674 -1419 675 -1417
rect 681 -1413 682 -1411
rect 684 -1413 685 -1411
rect 681 -1419 682 -1417
rect 688 -1413 689 -1411
rect 688 -1419 689 -1417
rect 695 -1413 696 -1411
rect 695 -1419 696 -1417
rect 705 -1413 706 -1411
rect 702 -1419 703 -1417
rect 709 -1413 710 -1411
rect 709 -1419 710 -1417
rect 712 -1419 713 -1417
rect 716 -1413 717 -1411
rect 716 -1419 717 -1417
rect 723 -1413 724 -1411
rect 723 -1419 724 -1417
rect 730 -1413 731 -1411
rect 730 -1419 731 -1417
rect 737 -1413 738 -1411
rect 744 -1413 745 -1411
rect 744 -1419 745 -1417
rect 751 -1413 752 -1411
rect 751 -1419 752 -1417
rect 758 -1413 759 -1411
rect 758 -1419 759 -1417
rect 765 -1419 766 -1417
rect 768 -1419 769 -1417
rect 772 -1413 773 -1411
rect 772 -1419 773 -1417
rect 779 -1413 780 -1411
rect 779 -1419 780 -1417
rect 786 -1413 787 -1411
rect 786 -1419 787 -1417
rect 793 -1413 794 -1411
rect 793 -1419 794 -1417
rect 800 -1413 801 -1411
rect 800 -1419 801 -1417
rect 807 -1413 808 -1411
rect 807 -1419 808 -1417
rect 814 -1413 815 -1411
rect 814 -1419 815 -1417
rect 821 -1413 822 -1411
rect 821 -1419 822 -1417
rect 828 -1413 829 -1411
rect 828 -1419 829 -1417
rect 835 -1413 836 -1411
rect 835 -1419 836 -1417
rect 842 -1413 843 -1411
rect 842 -1419 843 -1417
rect 849 -1413 850 -1411
rect 849 -1419 850 -1417
rect 856 -1413 857 -1411
rect 856 -1419 857 -1417
rect 863 -1413 864 -1411
rect 863 -1419 864 -1417
rect 870 -1413 871 -1411
rect 870 -1419 871 -1417
rect 877 -1413 878 -1411
rect 877 -1419 878 -1417
rect 884 -1413 885 -1411
rect 884 -1419 885 -1417
rect 891 -1413 892 -1411
rect 891 -1419 892 -1417
rect 898 -1413 899 -1411
rect 898 -1419 899 -1417
rect 905 -1413 906 -1411
rect 905 -1419 906 -1417
rect 912 -1413 913 -1411
rect 912 -1419 913 -1417
rect 919 -1413 920 -1411
rect 919 -1419 920 -1417
rect 926 -1419 927 -1417
rect 929 -1419 930 -1417
rect 933 -1413 934 -1411
rect 933 -1419 934 -1417
rect 940 -1413 941 -1411
rect 940 -1419 941 -1417
rect 950 -1413 951 -1411
rect 947 -1419 948 -1417
rect 950 -1419 951 -1417
rect 954 -1413 955 -1411
rect 954 -1419 955 -1417
rect 961 -1413 962 -1411
rect 961 -1419 962 -1417
rect 971 -1413 972 -1411
rect 968 -1419 969 -1417
rect 971 -1419 972 -1417
rect 975 -1413 976 -1411
rect 975 -1419 976 -1417
rect 982 -1413 983 -1411
rect 982 -1419 983 -1417
rect 989 -1413 990 -1411
rect 989 -1419 990 -1417
rect 996 -1413 997 -1411
rect 996 -1419 997 -1417
rect 1003 -1413 1004 -1411
rect 1006 -1419 1007 -1417
rect 1010 -1413 1011 -1411
rect 1010 -1419 1011 -1417
rect 1017 -1413 1018 -1411
rect 1017 -1419 1018 -1417
rect 1024 -1413 1025 -1411
rect 1024 -1419 1025 -1417
rect 1031 -1413 1032 -1411
rect 1031 -1419 1032 -1417
rect 1041 -1419 1042 -1417
rect 1045 -1413 1046 -1411
rect 1045 -1419 1046 -1417
rect 1052 -1413 1053 -1411
rect 1052 -1419 1053 -1417
rect 1073 -1413 1074 -1411
rect 1073 -1419 1074 -1417
rect 26 -1494 27 -1492
rect 30 -1494 31 -1492
rect 30 -1500 31 -1498
rect 37 -1494 38 -1492
rect 37 -1500 38 -1498
rect 44 -1494 45 -1492
rect 44 -1500 45 -1498
rect 51 -1494 52 -1492
rect 54 -1494 55 -1492
rect 58 -1494 59 -1492
rect 58 -1500 59 -1498
rect 65 -1494 66 -1492
rect 65 -1500 66 -1498
rect 72 -1494 73 -1492
rect 75 -1494 76 -1492
rect 75 -1500 76 -1498
rect 79 -1494 80 -1492
rect 79 -1500 80 -1498
rect 86 -1494 87 -1492
rect 86 -1500 87 -1498
rect 93 -1494 94 -1492
rect 93 -1500 94 -1498
rect 100 -1494 101 -1492
rect 100 -1500 101 -1498
rect 107 -1494 108 -1492
rect 107 -1500 108 -1498
rect 114 -1494 115 -1492
rect 114 -1500 115 -1498
rect 121 -1494 122 -1492
rect 124 -1494 125 -1492
rect 121 -1500 122 -1498
rect 128 -1494 129 -1492
rect 131 -1500 132 -1498
rect 135 -1494 136 -1492
rect 135 -1500 136 -1498
rect 142 -1494 143 -1492
rect 142 -1500 143 -1498
rect 149 -1494 150 -1492
rect 149 -1500 150 -1498
rect 156 -1494 157 -1492
rect 156 -1500 157 -1498
rect 163 -1494 164 -1492
rect 163 -1500 164 -1498
rect 170 -1494 171 -1492
rect 170 -1500 171 -1498
rect 177 -1494 178 -1492
rect 180 -1500 181 -1498
rect 184 -1494 185 -1492
rect 187 -1494 188 -1492
rect 187 -1500 188 -1498
rect 191 -1494 192 -1492
rect 191 -1500 192 -1498
rect 198 -1494 199 -1492
rect 198 -1500 199 -1498
rect 205 -1494 206 -1492
rect 205 -1500 206 -1498
rect 212 -1494 213 -1492
rect 212 -1500 213 -1498
rect 219 -1494 220 -1492
rect 219 -1500 220 -1498
rect 226 -1494 227 -1492
rect 226 -1500 227 -1498
rect 233 -1494 234 -1492
rect 233 -1500 234 -1498
rect 243 -1494 244 -1492
rect 240 -1500 241 -1498
rect 243 -1500 244 -1498
rect 247 -1494 248 -1492
rect 247 -1500 248 -1498
rect 254 -1494 255 -1492
rect 254 -1500 255 -1498
rect 261 -1494 262 -1492
rect 261 -1500 262 -1498
rect 268 -1494 269 -1492
rect 268 -1500 269 -1498
rect 275 -1494 276 -1492
rect 275 -1500 276 -1498
rect 282 -1494 283 -1492
rect 282 -1500 283 -1498
rect 289 -1494 290 -1492
rect 292 -1494 293 -1492
rect 292 -1500 293 -1498
rect 296 -1494 297 -1492
rect 296 -1500 297 -1498
rect 306 -1494 307 -1492
rect 303 -1500 304 -1498
rect 306 -1500 307 -1498
rect 310 -1494 311 -1492
rect 310 -1500 311 -1498
rect 313 -1500 314 -1498
rect 317 -1494 318 -1492
rect 320 -1494 321 -1492
rect 317 -1500 318 -1498
rect 324 -1494 325 -1492
rect 324 -1500 325 -1498
rect 331 -1494 332 -1492
rect 331 -1500 332 -1498
rect 338 -1494 339 -1492
rect 338 -1500 339 -1498
rect 345 -1494 346 -1492
rect 345 -1500 346 -1498
rect 352 -1494 353 -1492
rect 352 -1500 353 -1498
rect 359 -1494 360 -1492
rect 359 -1500 360 -1498
rect 366 -1494 367 -1492
rect 366 -1500 367 -1498
rect 373 -1494 374 -1492
rect 373 -1500 374 -1498
rect 380 -1494 381 -1492
rect 380 -1500 381 -1498
rect 387 -1494 388 -1492
rect 387 -1500 388 -1498
rect 394 -1494 395 -1492
rect 397 -1494 398 -1492
rect 394 -1500 395 -1498
rect 397 -1500 398 -1498
rect 401 -1494 402 -1492
rect 401 -1500 402 -1498
rect 408 -1494 409 -1492
rect 408 -1500 409 -1498
rect 415 -1494 416 -1492
rect 418 -1494 419 -1492
rect 415 -1500 416 -1498
rect 418 -1500 419 -1498
rect 422 -1494 423 -1492
rect 422 -1500 423 -1498
rect 429 -1494 430 -1492
rect 429 -1500 430 -1498
rect 436 -1494 437 -1492
rect 439 -1500 440 -1498
rect 443 -1494 444 -1492
rect 443 -1500 444 -1498
rect 450 -1494 451 -1492
rect 450 -1500 451 -1498
rect 457 -1494 458 -1492
rect 457 -1500 458 -1498
rect 464 -1494 465 -1492
rect 464 -1500 465 -1498
rect 471 -1494 472 -1492
rect 471 -1500 472 -1498
rect 478 -1494 479 -1492
rect 478 -1500 479 -1498
rect 485 -1494 486 -1492
rect 485 -1500 486 -1498
rect 492 -1494 493 -1492
rect 492 -1500 493 -1498
rect 499 -1494 500 -1492
rect 499 -1500 500 -1498
rect 506 -1494 507 -1492
rect 506 -1500 507 -1498
rect 513 -1494 514 -1492
rect 513 -1500 514 -1498
rect 520 -1494 521 -1492
rect 520 -1500 521 -1498
rect 527 -1494 528 -1492
rect 527 -1500 528 -1498
rect 537 -1494 538 -1492
rect 534 -1500 535 -1498
rect 537 -1500 538 -1498
rect 544 -1494 545 -1492
rect 544 -1500 545 -1498
rect 548 -1494 549 -1492
rect 548 -1500 549 -1498
rect 555 -1494 556 -1492
rect 558 -1494 559 -1492
rect 558 -1500 559 -1498
rect 562 -1494 563 -1492
rect 565 -1494 566 -1492
rect 562 -1500 563 -1498
rect 565 -1500 566 -1498
rect 569 -1494 570 -1492
rect 569 -1500 570 -1498
rect 579 -1494 580 -1492
rect 576 -1500 577 -1498
rect 579 -1500 580 -1498
rect 583 -1494 584 -1492
rect 583 -1500 584 -1498
rect 590 -1494 591 -1492
rect 590 -1500 591 -1498
rect 597 -1494 598 -1492
rect 597 -1500 598 -1498
rect 604 -1494 605 -1492
rect 604 -1500 605 -1498
rect 611 -1494 612 -1492
rect 611 -1500 612 -1498
rect 618 -1494 619 -1492
rect 618 -1500 619 -1498
rect 625 -1494 626 -1492
rect 625 -1500 626 -1498
rect 635 -1494 636 -1492
rect 639 -1494 640 -1492
rect 639 -1500 640 -1498
rect 646 -1494 647 -1492
rect 646 -1500 647 -1498
rect 656 -1494 657 -1492
rect 653 -1500 654 -1498
rect 656 -1500 657 -1498
rect 660 -1494 661 -1492
rect 660 -1500 661 -1498
rect 667 -1494 668 -1492
rect 667 -1500 668 -1498
rect 674 -1494 675 -1492
rect 674 -1500 675 -1498
rect 681 -1494 682 -1492
rect 684 -1494 685 -1492
rect 681 -1500 682 -1498
rect 684 -1500 685 -1498
rect 688 -1494 689 -1492
rect 688 -1500 689 -1498
rect 695 -1494 696 -1492
rect 695 -1500 696 -1498
rect 702 -1494 703 -1492
rect 702 -1500 703 -1498
rect 709 -1494 710 -1492
rect 709 -1500 710 -1498
rect 716 -1494 717 -1492
rect 716 -1500 717 -1498
rect 726 -1494 727 -1492
rect 723 -1500 724 -1498
rect 726 -1500 727 -1498
rect 730 -1494 731 -1492
rect 730 -1500 731 -1498
rect 737 -1494 738 -1492
rect 737 -1500 738 -1498
rect 744 -1494 745 -1492
rect 744 -1500 745 -1498
rect 751 -1494 752 -1492
rect 751 -1500 752 -1498
rect 758 -1494 759 -1492
rect 758 -1500 759 -1498
rect 765 -1494 766 -1492
rect 765 -1500 766 -1498
rect 772 -1494 773 -1492
rect 772 -1500 773 -1498
rect 779 -1494 780 -1492
rect 779 -1500 780 -1498
rect 786 -1494 787 -1492
rect 786 -1500 787 -1498
rect 793 -1494 794 -1492
rect 793 -1500 794 -1498
rect 800 -1500 801 -1498
rect 803 -1500 804 -1498
rect 807 -1494 808 -1492
rect 807 -1500 808 -1498
rect 814 -1494 815 -1492
rect 814 -1500 815 -1498
rect 821 -1494 822 -1492
rect 821 -1500 822 -1498
rect 828 -1494 829 -1492
rect 828 -1500 829 -1498
rect 835 -1494 836 -1492
rect 835 -1500 836 -1498
rect 842 -1494 843 -1492
rect 842 -1500 843 -1498
rect 849 -1494 850 -1492
rect 849 -1500 850 -1498
rect 856 -1494 857 -1492
rect 856 -1500 857 -1498
rect 863 -1494 864 -1492
rect 863 -1500 864 -1498
rect 870 -1494 871 -1492
rect 870 -1500 871 -1498
rect 877 -1494 878 -1492
rect 877 -1500 878 -1498
rect 884 -1494 885 -1492
rect 884 -1500 885 -1498
rect 891 -1494 892 -1492
rect 891 -1500 892 -1498
rect 898 -1494 899 -1492
rect 898 -1500 899 -1498
rect 905 -1494 906 -1492
rect 905 -1500 906 -1498
rect 912 -1494 913 -1492
rect 912 -1500 913 -1498
rect 919 -1494 920 -1492
rect 922 -1494 923 -1492
rect 922 -1500 923 -1498
rect 926 -1494 927 -1492
rect 926 -1500 927 -1498
rect 933 -1494 934 -1492
rect 933 -1500 934 -1498
rect 940 -1494 941 -1492
rect 943 -1494 944 -1492
rect 947 -1494 948 -1492
rect 947 -1500 948 -1498
rect 954 -1494 955 -1492
rect 954 -1500 955 -1498
rect 964 -1500 965 -1498
rect 971 -1494 972 -1492
rect 971 -1500 972 -1498
rect 975 -1494 976 -1492
rect 975 -1500 976 -1498
rect 982 -1494 983 -1492
rect 982 -1500 983 -1498
rect 989 -1494 990 -1492
rect 989 -1500 990 -1498
rect 996 -1494 997 -1492
rect 996 -1500 997 -1498
rect 1003 -1494 1004 -1492
rect 1003 -1500 1004 -1498
rect 1038 -1494 1039 -1492
rect 1038 -1500 1039 -1498
rect 1066 -1494 1067 -1492
rect 2 -1591 3 -1589
rect 2 -1597 3 -1595
rect 9 -1591 10 -1589
rect 9 -1597 10 -1595
rect 16 -1591 17 -1589
rect 16 -1597 17 -1595
rect 23 -1591 24 -1589
rect 23 -1597 24 -1595
rect 30 -1591 31 -1589
rect 30 -1597 31 -1595
rect 37 -1591 38 -1589
rect 37 -1597 38 -1595
rect 47 -1597 48 -1595
rect 51 -1591 52 -1589
rect 51 -1597 52 -1595
rect 58 -1591 59 -1589
rect 58 -1597 59 -1595
rect 65 -1591 66 -1589
rect 65 -1597 66 -1595
rect 72 -1591 73 -1589
rect 72 -1597 73 -1595
rect 75 -1597 76 -1595
rect 79 -1591 80 -1589
rect 82 -1591 83 -1589
rect 82 -1597 83 -1595
rect 86 -1591 87 -1589
rect 86 -1597 87 -1595
rect 93 -1591 94 -1589
rect 93 -1597 94 -1595
rect 100 -1591 101 -1589
rect 100 -1597 101 -1595
rect 107 -1591 108 -1589
rect 107 -1597 108 -1595
rect 114 -1591 115 -1589
rect 114 -1597 115 -1595
rect 124 -1591 125 -1589
rect 121 -1597 122 -1595
rect 124 -1597 125 -1595
rect 128 -1591 129 -1589
rect 128 -1597 129 -1595
rect 135 -1591 136 -1589
rect 135 -1597 136 -1595
rect 142 -1591 143 -1589
rect 142 -1597 143 -1595
rect 149 -1591 150 -1589
rect 149 -1597 150 -1595
rect 156 -1591 157 -1589
rect 156 -1597 157 -1595
rect 163 -1591 164 -1589
rect 163 -1597 164 -1595
rect 170 -1591 171 -1589
rect 170 -1597 171 -1595
rect 177 -1591 178 -1589
rect 177 -1597 178 -1595
rect 184 -1591 185 -1589
rect 184 -1597 185 -1595
rect 194 -1591 195 -1589
rect 194 -1597 195 -1595
rect 198 -1591 199 -1589
rect 198 -1597 199 -1595
rect 205 -1591 206 -1589
rect 205 -1597 206 -1595
rect 212 -1591 213 -1589
rect 212 -1597 213 -1595
rect 222 -1591 223 -1589
rect 222 -1597 223 -1595
rect 226 -1591 227 -1589
rect 229 -1591 230 -1589
rect 226 -1597 227 -1595
rect 233 -1591 234 -1589
rect 233 -1597 234 -1595
rect 240 -1591 241 -1589
rect 243 -1591 244 -1589
rect 243 -1597 244 -1595
rect 247 -1591 248 -1589
rect 247 -1597 248 -1595
rect 250 -1597 251 -1595
rect 254 -1591 255 -1589
rect 254 -1597 255 -1595
rect 261 -1591 262 -1589
rect 261 -1597 262 -1595
rect 268 -1591 269 -1589
rect 268 -1597 269 -1595
rect 275 -1591 276 -1589
rect 275 -1597 276 -1595
rect 282 -1591 283 -1589
rect 282 -1597 283 -1595
rect 289 -1591 290 -1589
rect 289 -1597 290 -1595
rect 296 -1591 297 -1589
rect 296 -1597 297 -1595
rect 303 -1591 304 -1589
rect 303 -1597 304 -1595
rect 310 -1591 311 -1589
rect 310 -1597 311 -1595
rect 317 -1591 318 -1589
rect 317 -1597 318 -1595
rect 324 -1591 325 -1589
rect 327 -1591 328 -1589
rect 331 -1591 332 -1589
rect 331 -1597 332 -1595
rect 338 -1591 339 -1589
rect 341 -1591 342 -1589
rect 338 -1597 339 -1595
rect 341 -1597 342 -1595
rect 345 -1591 346 -1589
rect 345 -1597 346 -1595
rect 352 -1591 353 -1589
rect 355 -1591 356 -1589
rect 355 -1597 356 -1595
rect 359 -1591 360 -1589
rect 362 -1591 363 -1589
rect 362 -1597 363 -1595
rect 366 -1591 367 -1589
rect 366 -1597 367 -1595
rect 373 -1591 374 -1589
rect 376 -1591 377 -1589
rect 373 -1597 374 -1595
rect 376 -1597 377 -1595
rect 380 -1591 381 -1589
rect 380 -1597 381 -1595
rect 387 -1591 388 -1589
rect 387 -1597 388 -1595
rect 394 -1591 395 -1589
rect 397 -1591 398 -1589
rect 394 -1597 395 -1595
rect 401 -1591 402 -1589
rect 401 -1597 402 -1595
rect 408 -1591 409 -1589
rect 408 -1597 409 -1595
rect 418 -1591 419 -1589
rect 422 -1591 423 -1589
rect 422 -1597 423 -1595
rect 429 -1591 430 -1589
rect 429 -1597 430 -1595
rect 436 -1591 437 -1589
rect 439 -1591 440 -1589
rect 436 -1597 437 -1595
rect 443 -1591 444 -1589
rect 443 -1597 444 -1595
rect 450 -1591 451 -1589
rect 450 -1597 451 -1595
rect 453 -1597 454 -1595
rect 457 -1591 458 -1589
rect 460 -1591 461 -1589
rect 457 -1597 458 -1595
rect 460 -1597 461 -1595
rect 464 -1591 465 -1589
rect 464 -1597 465 -1595
rect 471 -1591 472 -1589
rect 474 -1591 475 -1589
rect 471 -1597 472 -1595
rect 474 -1597 475 -1595
rect 478 -1591 479 -1589
rect 478 -1597 479 -1595
rect 485 -1591 486 -1589
rect 485 -1597 486 -1595
rect 495 -1591 496 -1589
rect 492 -1597 493 -1595
rect 499 -1591 500 -1589
rect 499 -1597 500 -1595
rect 506 -1591 507 -1589
rect 506 -1597 507 -1595
rect 513 -1591 514 -1589
rect 516 -1591 517 -1589
rect 513 -1597 514 -1595
rect 520 -1591 521 -1589
rect 520 -1597 521 -1595
rect 527 -1591 528 -1589
rect 527 -1597 528 -1595
rect 534 -1591 535 -1589
rect 537 -1597 538 -1595
rect 544 -1591 545 -1589
rect 544 -1597 545 -1595
rect 548 -1591 549 -1589
rect 548 -1597 549 -1595
rect 555 -1591 556 -1589
rect 555 -1597 556 -1595
rect 562 -1591 563 -1589
rect 562 -1597 563 -1595
rect 569 -1591 570 -1589
rect 569 -1597 570 -1595
rect 576 -1591 577 -1589
rect 576 -1597 577 -1595
rect 583 -1591 584 -1589
rect 583 -1597 584 -1595
rect 590 -1591 591 -1589
rect 590 -1597 591 -1595
rect 597 -1591 598 -1589
rect 597 -1597 598 -1595
rect 604 -1591 605 -1589
rect 604 -1597 605 -1595
rect 611 -1591 612 -1589
rect 611 -1597 612 -1595
rect 618 -1591 619 -1589
rect 618 -1597 619 -1595
rect 625 -1591 626 -1589
rect 625 -1597 626 -1595
rect 632 -1591 633 -1589
rect 632 -1597 633 -1595
rect 639 -1591 640 -1589
rect 639 -1597 640 -1595
rect 646 -1591 647 -1589
rect 646 -1597 647 -1595
rect 653 -1591 654 -1589
rect 653 -1597 654 -1595
rect 660 -1591 661 -1589
rect 663 -1591 664 -1589
rect 663 -1597 664 -1595
rect 667 -1591 668 -1589
rect 667 -1597 668 -1595
rect 674 -1591 675 -1589
rect 674 -1597 675 -1595
rect 681 -1591 682 -1589
rect 684 -1591 685 -1589
rect 684 -1597 685 -1595
rect 688 -1591 689 -1589
rect 688 -1597 689 -1595
rect 695 -1591 696 -1589
rect 695 -1597 696 -1595
rect 702 -1591 703 -1589
rect 702 -1597 703 -1595
rect 709 -1591 710 -1589
rect 712 -1591 713 -1589
rect 709 -1597 710 -1595
rect 716 -1591 717 -1589
rect 716 -1597 717 -1595
rect 723 -1591 724 -1589
rect 723 -1597 724 -1595
rect 733 -1591 734 -1589
rect 730 -1597 731 -1595
rect 733 -1597 734 -1595
rect 737 -1591 738 -1589
rect 737 -1597 738 -1595
rect 744 -1591 745 -1589
rect 744 -1597 745 -1595
rect 751 -1591 752 -1589
rect 751 -1597 752 -1595
rect 758 -1591 759 -1589
rect 758 -1597 759 -1595
rect 765 -1591 766 -1589
rect 765 -1597 766 -1595
rect 772 -1591 773 -1589
rect 772 -1597 773 -1595
rect 779 -1591 780 -1589
rect 779 -1597 780 -1595
rect 786 -1591 787 -1589
rect 786 -1597 787 -1595
rect 793 -1591 794 -1589
rect 793 -1597 794 -1595
rect 800 -1591 801 -1589
rect 803 -1591 804 -1589
rect 803 -1597 804 -1595
rect 807 -1591 808 -1589
rect 807 -1597 808 -1595
rect 814 -1591 815 -1589
rect 814 -1597 815 -1595
rect 821 -1591 822 -1589
rect 821 -1597 822 -1595
rect 828 -1591 829 -1589
rect 828 -1597 829 -1595
rect 835 -1591 836 -1589
rect 835 -1597 836 -1595
rect 842 -1591 843 -1589
rect 842 -1597 843 -1595
rect 849 -1591 850 -1589
rect 849 -1597 850 -1595
rect 856 -1591 857 -1589
rect 856 -1597 857 -1595
rect 863 -1591 864 -1589
rect 863 -1597 864 -1595
rect 870 -1591 871 -1589
rect 870 -1597 871 -1595
rect 877 -1591 878 -1589
rect 877 -1597 878 -1595
rect 884 -1591 885 -1589
rect 884 -1597 885 -1595
rect 891 -1591 892 -1589
rect 891 -1597 892 -1595
rect 898 -1591 899 -1589
rect 898 -1597 899 -1595
rect 905 -1591 906 -1589
rect 905 -1597 906 -1595
rect 912 -1591 913 -1589
rect 912 -1597 913 -1595
rect 919 -1591 920 -1589
rect 919 -1597 920 -1595
rect 926 -1591 927 -1589
rect 926 -1597 927 -1595
rect 933 -1591 934 -1589
rect 933 -1597 934 -1595
rect 940 -1591 941 -1589
rect 940 -1597 941 -1595
rect 947 -1591 948 -1589
rect 947 -1597 948 -1595
rect 954 -1591 955 -1589
rect 954 -1597 955 -1595
rect 961 -1591 962 -1589
rect 961 -1597 962 -1595
rect 968 -1591 969 -1589
rect 968 -1597 969 -1595
rect 975 -1591 976 -1589
rect 975 -1597 976 -1595
rect 982 -1591 983 -1589
rect 982 -1597 983 -1595
rect 989 -1591 990 -1589
rect 989 -1597 990 -1595
rect 996 -1591 997 -1589
rect 996 -1597 997 -1595
rect 1003 -1591 1004 -1589
rect 1003 -1597 1004 -1595
rect 1010 -1591 1011 -1589
rect 1010 -1597 1011 -1595
rect 1017 -1591 1018 -1589
rect 1017 -1597 1018 -1595
rect 1024 -1591 1025 -1589
rect 1024 -1597 1025 -1595
rect 1031 -1591 1032 -1589
rect 1031 -1597 1032 -1595
rect 1038 -1591 1039 -1589
rect 1038 -1597 1039 -1595
rect 1045 -1591 1046 -1589
rect 1045 -1597 1046 -1595
rect 1052 -1591 1053 -1589
rect 1052 -1597 1053 -1595
rect 1059 -1591 1060 -1589
rect 1059 -1597 1060 -1595
rect 1066 -1591 1067 -1589
rect 1066 -1597 1067 -1595
rect 1073 -1591 1074 -1589
rect 1073 -1597 1074 -1595
rect 1080 -1591 1081 -1589
rect 1080 -1597 1081 -1595
rect 1087 -1591 1088 -1589
rect 1087 -1597 1088 -1595
rect 1094 -1591 1095 -1589
rect 1094 -1597 1095 -1595
rect 1101 -1591 1102 -1589
rect 1101 -1597 1102 -1595
rect 1108 -1591 1109 -1589
rect 1111 -1591 1112 -1589
rect 1108 -1597 1109 -1595
rect 2 -1678 3 -1676
rect 2 -1684 3 -1682
rect 9 -1678 10 -1676
rect 9 -1684 10 -1682
rect 16 -1678 17 -1676
rect 16 -1684 17 -1682
rect 23 -1678 24 -1676
rect 23 -1684 24 -1682
rect 30 -1678 31 -1676
rect 30 -1684 31 -1682
rect 37 -1678 38 -1676
rect 37 -1684 38 -1682
rect 44 -1678 45 -1676
rect 44 -1684 45 -1682
rect 51 -1678 52 -1676
rect 51 -1684 52 -1682
rect 61 -1678 62 -1676
rect 65 -1678 66 -1676
rect 65 -1684 66 -1682
rect 72 -1678 73 -1676
rect 72 -1684 73 -1682
rect 79 -1678 80 -1676
rect 86 -1678 87 -1676
rect 86 -1684 87 -1682
rect 96 -1684 97 -1682
rect 100 -1678 101 -1676
rect 100 -1684 101 -1682
rect 107 -1678 108 -1676
rect 107 -1684 108 -1682
rect 114 -1678 115 -1676
rect 114 -1684 115 -1682
rect 121 -1678 122 -1676
rect 121 -1684 122 -1682
rect 128 -1678 129 -1676
rect 128 -1684 129 -1682
rect 135 -1678 136 -1676
rect 138 -1678 139 -1676
rect 138 -1684 139 -1682
rect 142 -1678 143 -1676
rect 142 -1684 143 -1682
rect 149 -1678 150 -1676
rect 149 -1684 150 -1682
rect 152 -1684 153 -1682
rect 159 -1678 160 -1676
rect 156 -1684 157 -1682
rect 163 -1678 164 -1676
rect 163 -1684 164 -1682
rect 170 -1678 171 -1676
rect 170 -1684 171 -1682
rect 177 -1678 178 -1676
rect 177 -1684 178 -1682
rect 184 -1678 185 -1676
rect 184 -1684 185 -1682
rect 194 -1678 195 -1676
rect 191 -1684 192 -1682
rect 194 -1684 195 -1682
rect 198 -1678 199 -1676
rect 198 -1684 199 -1682
rect 201 -1684 202 -1682
rect 205 -1678 206 -1676
rect 205 -1684 206 -1682
rect 212 -1678 213 -1676
rect 215 -1684 216 -1682
rect 222 -1678 223 -1676
rect 222 -1684 223 -1682
rect 226 -1678 227 -1676
rect 226 -1684 227 -1682
rect 229 -1684 230 -1682
rect 233 -1678 234 -1676
rect 236 -1678 237 -1676
rect 240 -1678 241 -1676
rect 240 -1684 241 -1682
rect 247 -1678 248 -1676
rect 247 -1684 248 -1682
rect 254 -1678 255 -1676
rect 254 -1684 255 -1682
rect 261 -1678 262 -1676
rect 261 -1684 262 -1682
rect 268 -1678 269 -1676
rect 268 -1684 269 -1682
rect 275 -1678 276 -1676
rect 275 -1684 276 -1682
rect 282 -1678 283 -1676
rect 285 -1684 286 -1682
rect 289 -1678 290 -1676
rect 289 -1684 290 -1682
rect 292 -1684 293 -1682
rect 296 -1678 297 -1676
rect 299 -1678 300 -1676
rect 299 -1684 300 -1682
rect 303 -1678 304 -1676
rect 303 -1684 304 -1682
rect 310 -1678 311 -1676
rect 310 -1684 311 -1682
rect 317 -1678 318 -1676
rect 317 -1684 318 -1682
rect 324 -1678 325 -1676
rect 324 -1684 325 -1682
rect 331 -1678 332 -1676
rect 331 -1684 332 -1682
rect 338 -1678 339 -1676
rect 338 -1684 339 -1682
rect 345 -1678 346 -1676
rect 345 -1684 346 -1682
rect 348 -1684 349 -1682
rect 352 -1678 353 -1676
rect 352 -1684 353 -1682
rect 359 -1678 360 -1676
rect 359 -1684 360 -1682
rect 366 -1678 367 -1676
rect 366 -1684 367 -1682
rect 369 -1684 370 -1682
rect 373 -1678 374 -1676
rect 373 -1684 374 -1682
rect 380 -1684 381 -1682
rect 383 -1684 384 -1682
rect 387 -1678 388 -1676
rect 390 -1678 391 -1676
rect 394 -1678 395 -1676
rect 394 -1684 395 -1682
rect 401 -1678 402 -1676
rect 401 -1684 402 -1682
rect 408 -1678 409 -1676
rect 408 -1684 409 -1682
rect 415 -1678 416 -1676
rect 415 -1684 416 -1682
rect 422 -1678 423 -1676
rect 422 -1684 423 -1682
rect 429 -1678 430 -1676
rect 429 -1684 430 -1682
rect 436 -1678 437 -1676
rect 436 -1684 437 -1682
rect 443 -1678 444 -1676
rect 443 -1684 444 -1682
rect 450 -1678 451 -1676
rect 453 -1678 454 -1676
rect 450 -1684 451 -1682
rect 453 -1684 454 -1682
rect 457 -1678 458 -1676
rect 457 -1684 458 -1682
rect 464 -1678 465 -1676
rect 467 -1678 468 -1676
rect 464 -1684 465 -1682
rect 467 -1684 468 -1682
rect 474 -1678 475 -1676
rect 471 -1684 472 -1682
rect 474 -1684 475 -1682
rect 478 -1678 479 -1676
rect 481 -1678 482 -1676
rect 478 -1684 479 -1682
rect 481 -1684 482 -1682
rect 488 -1678 489 -1676
rect 485 -1684 486 -1682
rect 488 -1684 489 -1682
rect 492 -1678 493 -1676
rect 492 -1684 493 -1682
rect 495 -1684 496 -1682
rect 499 -1678 500 -1676
rect 499 -1684 500 -1682
rect 506 -1678 507 -1676
rect 506 -1684 507 -1682
rect 513 -1678 514 -1676
rect 513 -1684 514 -1682
rect 520 -1678 521 -1676
rect 520 -1684 521 -1682
rect 527 -1678 528 -1676
rect 527 -1684 528 -1682
rect 534 -1678 535 -1676
rect 537 -1678 538 -1676
rect 541 -1678 542 -1676
rect 541 -1684 542 -1682
rect 548 -1678 549 -1676
rect 548 -1684 549 -1682
rect 551 -1684 552 -1682
rect 555 -1678 556 -1676
rect 558 -1678 559 -1676
rect 558 -1684 559 -1682
rect 565 -1678 566 -1676
rect 562 -1684 563 -1682
rect 565 -1684 566 -1682
rect 569 -1678 570 -1676
rect 569 -1684 570 -1682
rect 576 -1678 577 -1676
rect 576 -1684 577 -1682
rect 583 -1678 584 -1676
rect 583 -1684 584 -1682
rect 590 -1678 591 -1676
rect 590 -1684 591 -1682
rect 597 -1678 598 -1676
rect 597 -1684 598 -1682
rect 604 -1678 605 -1676
rect 604 -1684 605 -1682
rect 611 -1678 612 -1676
rect 611 -1684 612 -1682
rect 618 -1678 619 -1676
rect 618 -1684 619 -1682
rect 625 -1678 626 -1676
rect 625 -1684 626 -1682
rect 632 -1678 633 -1676
rect 632 -1684 633 -1682
rect 639 -1678 640 -1676
rect 639 -1684 640 -1682
rect 646 -1678 647 -1676
rect 646 -1684 647 -1682
rect 653 -1678 654 -1676
rect 653 -1684 654 -1682
rect 660 -1678 661 -1676
rect 660 -1684 661 -1682
rect 667 -1678 668 -1676
rect 667 -1684 668 -1682
rect 674 -1678 675 -1676
rect 674 -1684 675 -1682
rect 681 -1678 682 -1676
rect 681 -1684 682 -1682
rect 688 -1678 689 -1676
rect 688 -1684 689 -1682
rect 695 -1678 696 -1676
rect 695 -1684 696 -1682
rect 702 -1678 703 -1676
rect 702 -1684 703 -1682
rect 709 -1678 710 -1676
rect 709 -1684 710 -1682
rect 716 -1678 717 -1676
rect 716 -1684 717 -1682
rect 723 -1678 724 -1676
rect 723 -1684 724 -1682
rect 730 -1684 731 -1682
rect 733 -1684 734 -1682
rect 737 -1678 738 -1676
rect 737 -1684 738 -1682
rect 744 -1678 745 -1676
rect 744 -1684 745 -1682
rect 751 -1678 752 -1676
rect 751 -1684 752 -1682
rect 758 -1678 759 -1676
rect 758 -1684 759 -1682
rect 765 -1678 766 -1676
rect 765 -1684 766 -1682
rect 772 -1678 773 -1676
rect 772 -1684 773 -1682
rect 779 -1678 780 -1676
rect 779 -1684 780 -1682
rect 786 -1678 787 -1676
rect 786 -1684 787 -1682
rect 793 -1678 794 -1676
rect 793 -1684 794 -1682
rect 800 -1678 801 -1676
rect 800 -1684 801 -1682
rect 807 -1678 808 -1676
rect 807 -1684 808 -1682
rect 814 -1678 815 -1676
rect 814 -1684 815 -1682
rect 821 -1678 822 -1676
rect 824 -1678 825 -1676
rect 821 -1684 822 -1682
rect 828 -1678 829 -1676
rect 828 -1684 829 -1682
rect 835 -1678 836 -1676
rect 835 -1684 836 -1682
rect 842 -1678 843 -1676
rect 842 -1684 843 -1682
rect 849 -1678 850 -1676
rect 849 -1684 850 -1682
rect 856 -1678 857 -1676
rect 856 -1684 857 -1682
rect 863 -1678 864 -1676
rect 863 -1684 864 -1682
rect 870 -1678 871 -1676
rect 870 -1684 871 -1682
rect 877 -1678 878 -1676
rect 877 -1684 878 -1682
rect 887 -1678 888 -1676
rect 884 -1684 885 -1682
rect 887 -1684 888 -1682
rect 891 -1678 892 -1676
rect 894 -1678 895 -1676
rect 891 -1684 892 -1682
rect 894 -1684 895 -1682
rect 898 -1678 899 -1676
rect 898 -1684 899 -1682
rect 905 -1678 906 -1676
rect 905 -1684 906 -1682
rect 915 -1678 916 -1676
rect 912 -1684 913 -1682
rect 919 -1678 920 -1676
rect 919 -1684 920 -1682
rect 926 -1678 927 -1676
rect 926 -1684 927 -1682
rect 933 -1678 934 -1676
rect 933 -1684 934 -1682
rect 940 -1678 941 -1676
rect 940 -1684 941 -1682
rect 947 -1678 948 -1676
rect 947 -1684 948 -1682
rect 954 -1678 955 -1676
rect 954 -1684 955 -1682
rect 961 -1678 962 -1676
rect 961 -1684 962 -1682
rect 975 -1678 976 -1676
rect 975 -1684 976 -1682
rect 982 -1678 983 -1676
rect 982 -1684 983 -1682
rect 1003 -1678 1004 -1676
rect 1003 -1684 1004 -1682
rect 1024 -1684 1025 -1682
rect 1027 -1684 1028 -1682
rect 1052 -1678 1053 -1676
rect 1052 -1684 1053 -1682
rect 2 -1773 3 -1771
rect 2 -1779 3 -1777
rect 9 -1779 10 -1777
rect 16 -1773 17 -1771
rect 23 -1773 24 -1771
rect 23 -1779 24 -1777
rect 30 -1773 31 -1771
rect 30 -1779 31 -1777
rect 37 -1773 38 -1771
rect 37 -1779 38 -1777
rect 44 -1773 45 -1771
rect 44 -1779 45 -1777
rect 51 -1773 52 -1771
rect 54 -1773 55 -1771
rect 51 -1779 52 -1777
rect 54 -1779 55 -1777
rect 61 -1773 62 -1771
rect 65 -1773 66 -1771
rect 65 -1779 66 -1777
rect 72 -1773 73 -1771
rect 72 -1779 73 -1777
rect 79 -1773 80 -1771
rect 79 -1779 80 -1777
rect 86 -1773 87 -1771
rect 86 -1779 87 -1777
rect 93 -1773 94 -1771
rect 93 -1779 94 -1777
rect 100 -1773 101 -1771
rect 103 -1773 104 -1771
rect 100 -1779 101 -1777
rect 103 -1779 104 -1777
rect 107 -1773 108 -1771
rect 110 -1773 111 -1771
rect 110 -1779 111 -1777
rect 114 -1773 115 -1771
rect 114 -1779 115 -1777
rect 121 -1773 122 -1771
rect 121 -1779 122 -1777
rect 128 -1773 129 -1771
rect 128 -1779 129 -1777
rect 135 -1773 136 -1771
rect 135 -1779 136 -1777
rect 142 -1773 143 -1771
rect 142 -1779 143 -1777
rect 149 -1773 150 -1771
rect 149 -1779 150 -1777
rect 156 -1773 157 -1771
rect 156 -1779 157 -1777
rect 163 -1773 164 -1771
rect 166 -1773 167 -1771
rect 170 -1773 171 -1771
rect 170 -1779 171 -1777
rect 177 -1773 178 -1771
rect 180 -1773 181 -1771
rect 177 -1779 178 -1777
rect 187 -1773 188 -1771
rect 187 -1779 188 -1777
rect 191 -1773 192 -1771
rect 191 -1779 192 -1777
rect 198 -1773 199 -1771
rect 198 -1779 199 -1777
rect 205 -1773 206 -1771
rect 205 -1779 206 -1777
rect 215 -1779 216 -1777
rect 222 -1773 223 -1771
rect 219 -1779 220 -1777
rect 226 -1773 227 -1771
rect 226 -1779 227 -1777
rect 233 -1773 234 -1771
rect 233 -1779 234 -1777
rect 240 -1773 241 -1771
rect 243 -1773 244 -1771
rect 240 -1779 241 -1777
rect 243 -1779 244 -1777
rect 247 -1773 248 -1771
rect 247 -1779 248 -1777
rect 254 -1773 255 -1771
rect 254 -1779 255 -1777
rect 261 -1773 262 -1771
rect 261 -1779 262 -1777
rect 268 -1773 269 -1771
rect 268 -1779 269 -1777
rect 275 -1773 276 -1771
rect 275 -1779 276 -1777
rect 282 -1773 283 -1771
rect 282 -1779 283 -1777
rect 289 -1773 290 -1771
rect 289 -1779 290 -1777
rect 296 -1773 297 -1771
rect 296 -1779 297 -1777
rect 303 -1773 304 -1771
rect 303 -1779 304 -1777
rect 313 -1773 314 -1771
rect 310 -1779 311 -1777
rect 313 -1779 314 -1777
rect 317 -1773 318 -1771
rect 317 -1779 318 -1777
rect 324 -1773 325 -1771
rect 324 -1779 325 -1777
rect 327 -1779 328 -1777
rect 331 -1773 332 -1771
rect 331 -1779 332 -1777
rect 338 -1773 339 -1771
rect 338 -1779 339 -1777
rect 345 -1773 346 -1771
rect 345 -1779 346 -1777
rect 352 -1773 353 -1771
rect 352 -1779 353 -1777
rect 359 -1773 360 -1771
rect 359 -1779 360 -1777
rect 366 -1773 367 -1771
rect 369 -1773 370 -1771
rect 366 -1779 367 -1777
rect 369 -1779 370 -1777
rect 373 -1773 374 -1771
rect 376 -1773 377 -1771
rect 373 -1779 374 -1777
rect 376 -1779 377 -1777
rect 383 -1773 384 -1771
rect 380 -1779 381 -1777
rect 387 -1773 388 -1771
rect 387 -1779 388 -1777
rect 394 -1773 395 -1771
rect 394 -1779 395 -1777
rect 401 -1773 402 -1771
rect 404 -1773 405 -1771
rect 401 -1779 402 -1777
rect 408 -1773 409 -1771
rect 411 -1773 412 -1771
rect 408 -1779 409 -1777
rect 415 -1773 416 -1771
rect 415 -1779 416 -1777
rect 422 -1773 423 -1771
rect 425 -1773 426 -1771
rect 429 -1773 430 -1771
rect 429 -1779 430 -1777
rect 436 -1773 437 -1771
rect 436 -1779 437 -1777
rect 443 -1773 444 -1771
rect 443 -1779 444 -1777
rect 450 -1773 451 -1771
rect 450 -1779 451 -1777
rect 457 -1773 458 -1771
rect 457 -1779 458 -1777
rect 464 -1773 465 -1771
rect 467 -1773 468 -1771
rect 464 -1779 465 -1777
rect 467 -1779 468 -1777
rect 471 -1773 472 -1771
rect 471 -1779 472 -1777
rect 478 -1773 479 -1771
rect 481 -1773 482 -1771
rect 485 -1773 486 -1771
rect 485 -1779 486 -1777
rect 492 -1773 493 -1771
rect 492 -1779 493 -1777
rect 499 -1773 500 -1771
rect 499 -1779 500 -1777
rect 506 -1773 507 -1771
rect 506 -1779 507 -1777
rect 513 -1773 514 -1771
rect 516 -1773 517 -1771
rect 516 -1779 517 -1777
rect 520 -1773 521 -1771
rect 520 -1779 521 -1777
rect 527 -1773 528 -1771
rect 527 -1779 528 -1777
rect 534 -1773 535 -1771
rect 534 -1779 535 -1777
rect 541 -1773 542 -1771
rect 541 -1779 542 -1777
rect 548 -1773 549 -1771
rect 548 -1779 549 -1777
rect 555 -1773 556 -1771
rect 555 -1779 556 -1777
rect 562 -1773 563 -1771
rect 562 -1779 563 -1777
rect 569 -1773 570 -1771
rect 569 -1779 570 -1777
rect 576 -1773 577 -1771
rect 576 -1779 577 -1777
rect 583 -1773 584 -1771
rect 583 -1779 584 -1777
rect 593 -1773 594 -1771
rect 590 -1779 591 -1777
rect 593 -1779 594 -1777
rect 597 -1773 598 -1771
rect 597 -1779 598 -1777
rect 604 -1773 605 -1771
rect 604 -1779 605 -1777
rect 614 -1773 615 -1771
rect 611 -1779 612 -1777
rect 618 -1773 619 -1771
rect 621 -1773 622 -1771
rect 618 -1779 619 -1777
rect 621 -1779 622 -1777
rect 625 -1773 626 -1771
rect 625 -1779 626 -1777
rect 632 -1779 633 -1777
rect 635 -1779 636 -1777
rect 639 -1773 640 -1771
rect 639 -1779 640 -1777
rect 646 -1773 647 -1771
rect 649 -1773 650 -1771
rect 646 -1779 647 -1777
rect 653 -1773 654 -1771
rect 653 -1779 654 -1777
rect 656 -1779 657 -1777
rect 660 -1773 661 -1771
rect 660 -1779 661 -1777
rect 667 -1773 668 -1771
rect 667 -1779 668 -1777
rect 674 -1773 675 -1771
rect 677 -1773 678 -1771
rect 674 -1779 675 -1777
rect 677 -1779 678 -1777
rect 681 -1773 682 -1771
rect 681 -1779 682 -1777
rect 688 -1773 689 -1771
rect 688 -1779 689 -1777
rect 695 -1773 696 -1771
rect 695 -1779 696 -1777
rect 702 -1773 703 -1771
rect 702 -1779 703 -1777
rect 709 -1773 710 -1771
rect 709 -1779 710 -1777
rect 716 -1773 717 -1771
rect 716 -1779 717 -1777
rect 723 -1773 724 -1771
rect 723 -1779 724 -1777
rect 730 -1773 731 -1771
rect 730 -1779 731 -1777
rect 737 -1773 738 -1771
rect 737 -1779 738 -1777
rect 744 -1773 745 -1771
rect 744 -1779 745 -1777
rect 751 -1773 752 -1771
rect 751 -1779 752 -1777
rect 758 -1773 759 -1771
rect 758 -1779 759 -1777
rect 765 -1773 766 -1771
rect 765 -1779 766 -1777
rect 772 -1773 773 -1771
rect 772 -1779 773 -1777
rect 779 -1773 780 -1771
rect 779 -1779 780 -1777
rect 786 -1773 787 -1771
rect 786 -1779 787 -1777
rect 793 -1773 794 -1771
rect 793 -1779 794 -1777
rect 803 -1773 804 -1771
rect 807 -1773 808 -1771
rect 807 -1779 808 -1777
rect 814 -1773 815 -1771
rect 814 -1779 815 -1777
rect 821 -1773 822 -1771
rect 821 -1779 822 -1777
rect 828 -1773 829 -1771
rect 828 -1779 829 -1777
rect 835 -1773 836 -1771
rect 835 -1779 836 -1777
rect 842 -1773 843 -1771
rect 842 -1779 843 -1777
rect 849 -1773 850 -1771
rect 849 -1779 850 -1777
rect 856 -1773 857 -1771
rect 856 -1779 857 -1777
rect 863 -1773 864 -1771
rect 863 -1779 864 -1777
rect 870 -1773 871 -1771
rect 870 -1779 871 -1777
rect 877 -1773 878 -1771
rect 877 -1779 878 -1777
rect 884 -1773 885 -1771
rect 884 -1779 885 -1777
rect 891 -1773 892 -1771
rect 891 -1779 892 -1777
rect 898 -1773 899 -1771
rect 898 -1779 899 -1777
rect 905 -1773 906 -1771
rect 905 -1779 906 -1777
rect 912 -1773 913 -1771
rect 912 -1779 913 -1777
rect 919 -1773 920 -1771
rect 919 -1779 920 -1777
rect 926 -1773 927 -1771
rect 926 -1779 927 -1777
rect 933 -1773 934 -1771
rect 933 -1779 934 -1777
rect 940 -1773 941 -1771
rect 940 -1779 941 -1777
rect 947 -1773 948 -1771
rect 947 -1779 948 -1777
rect 954 -1773 955 -1771
rect 954 -1779 955 -1777
rect 961 -1773 962 -1771
rect 961 -1779 962 -1777
rect 968 -1773 969 -1771
rect 968 -1779 969 -1777
rect 975 -1773 976 -1771
rect 975 -1779 976 -1777
rect 982 -1773 983 -1771
rect 982 -1779 983 -1777
rect 989 -1773 990 -1771
rect 989 -1779 990 -1777
rect 996 -1779 997 -1777
rect 999 -1779 1000 -1777
rect 1006 -1773 1007 -1771
rect 1003 -1779 1004 -1777
rect 1010 -1773 1011 -1771
rect 1010 -1779 1011 -1777
rect 1017 -1773 1018 -1771
rect 1017 -1779 1018 -1777
rect 1024 -1773 1025 -1771
rect 1024 -1779 1025 -1777
rect 51 -1864 52 -1862
rect 51 -1870 52 -1868
rect 58 -1864 59 -1862
rect 58 -1870 59 -1868
rect 65 -1864 66 -1862
rect 65 -1870 66 -1868
rect 72 -1864 73 -1862
rect 72 -1870 73 -1868
rect 79 -1864 80 -1862
rect 79 -1870 80 -1868
rect 86 -1864 87 -1862
rect 86 -1870 87 -1868
rect 93 -1864 94 -1862
rect 93 -1870 94 -1868
rect 100 -1864 101 -1862
rect 100 -1870 101 -1868
rect 107 -1864 108 -1862
rect 107 -1870 108 -1868
rect 114 -1864 115 -1862
rect 114 -1870 115 -1868
rect 121 -1864 122 -1862
rect 121 -1870 122 -1868
rect 128 -1864 129 -1862
rect 131 -1870 132 -1868
rect 135 -1864 136 -1862
rect 135 -1870 136 -1868
rect 142 -1864 143 -1862
rect 142 -1870 143 -1868
rect 149 -1864 150 -1862
rect 149 -1870 150 -1868
rect 156 -1864 157 -1862
rect 156 -1870 157 -1868
rect 163 -1864 164 -1862
rect 163 -1870 164 -1868
rect 166 -1870 167 -1868
rect 170 -1864 171 -1862
rect 170 -1870 171 -1868
rect 177 -1864 178 -1862
rect 177 -1870 178 -1868
rect 184 -1864 185 -1862
rect 184 -1870 185 -1868
rect 194 -1864 195 -1862
rect 191 -1870 192 -1868
rect 201 -1864 202 -1862
rect 198 -1870 199 -1868
rect 205 -1870 206 -1868
rect 212 -1864 213 -1862
rect 215 -1864 216 -1862
rect 212 -1870 213 -1868
rect 215 -1870 216 -1868
rect 219 -1864 220 -1862
rect 219 -1870 220 -1868
rect 226 -1864 227 -1862
rect 229 -1864 230 -1862
rect 229 -1870 230 -1868
rect 233 -1864 234 -1862
rect 233 -1870 234 -1868
rect 240 -1870 241 -1868
rect 243 -1870 244 -1868
rect 247 -1864 248 -1862
rect 247 -1870 248 -1868
rect 254 -1864 255 -1862
rect 254 -1870 255 -1868
rect 261 -1864 262 -1862
rect 261 -1870 262 -1868
rect 268 -1864 269 -1862
rect 268 -1870 269 -1868
rect 275 -1864 276 -1862
rect 275 -1870 276 -1868
rect 282 -1864 283 -1862
rect 282 -1870 283 -1868
rect 289 -1864 290 -1862
rect 289 -1870 290 -1868
rect 296 -1864 297 -1862
rect 296 -1870 297 -1868
rect 303 -1864 304 -1862
rect 303 -1870 304 -1868
rect 310 -1864 311 -1862
rect 310 -1870 311 -1868
rect 317 -1864 318 -1862
rect 317 -1870 318 -1868
rect 324 -1864 325 -1862
rect 324 -1870 325 -1868
rect 331 -1864 332 -1862
rect 331 -1870 332 -1868
rect 338 -1864 339 -1862
rect 338 -1870 339 -1868
rect 345 -1864 346 -1862
rect 348 -1864 349 -1862
rect 345 -1870 346 -1868
rect 348 -1870 349 -1868
rect 352 -1864 353 -1862
rect 352 -1870 353 -1868
rect 362 -1870 363 -1868
rect 369 -1864 370 -1862
rect 373 -1864 374 -1862
rect 373 -1870 374 -1868
rect 380 -1864 381 -1862
rect 380 -1870 381 -1868
rect 387 -1864 388 -1862
rect 387 -1870 388 -1868
rect 394 -1864 395 -1862
rect 394 -1870 395 -1868
rect 401 -1864 402 -1862
rect 401 -1870 402 -1868
rect 408 -1864 409 -1862
rect 408 -1870 409 -1868
rect 411 -1870 412 -1868
rect 415 -1864 416 -1862
rect 418 -1864 419 -1862
rect 415 -1870 416 -1868
rect 418 -1870 419 -1868
rect 422 -1864 423 -1862
rect 425 -1864 426 -1862
rect 422 -1870 423 -1868
rect 429 -1864 430 -1862
rect 429 -1870 430 -1868
rect 436 -1864 437 -1862
rect 436 -1870 437 -1868
rect 443 -1864 444 -1862
rect 443 -1870 444 -1868
rect 450 -1864 451 -1862
rect 450 -1870 451 -1868
rect 457 -1864 458 -1862
rect 460 -1864 461 -1862
rect 457 -1870 458 -1868
rect 464 -1864 465 -1862
rect 464 -1870 465 -1868
rect 471 -1864 472 -1862
rect 471 -1870 472 -1868
rect 478 -1864 479 -1862
rect 478 -1870 479 -1868
rect 485 -1864 486 -1862
rect 485 -1870 486 -1868
rect 492 -1864 493 -1862
rect 492 -1870 493 -1868
rect 499 -1864 500 -1862
rect 499 -1870 500 -1868
rect 506 -1864 507 -1862
rect 506 -1870 507 -1868
rect 509 -1870 510 -1868
rect 513 -1864 514 -1862
rect 513 -1870 514 -1868
rect 520 -1864 521 -1862
rect 523 -1864 524 -1862
rect 523 -1870 524 -1868
rect 527 -1864 528 -1862
rect 530 -1870 531 -1868
rect 534 -1864 535 -1862
rect 534 -1870 535 -1868
rect 541 -1864 542 -1862
rect 541 -1870 542 -1868
rect 548 -1864 549 -1862
rect 551 -1864 552 -1862
rect 548 -1870 549 -1868
rect 551 -1870 552 -1868
rect 555 -1864 556 -1862
rect 555 -1870 556 -1868
rect 562 -1864 563 -1862
rect 565 -1864 566 -1862
rect 562 -1870 563 -1868
rect 569 -1864 570 -1862
rect 569 -1870 570 -1868
rect 576 -1864 577 -1862
rect 576 -1870 577 -1868
rect 583 -1864 584 -1862
rect 583 -1870 584 -1868
rect 590 -1864 591 -1862
rect 590 -1870 591 -1868
rect 597 -1864 598 -1862
rect 597 -1870 598 -1868
rect 604 -1864 605 -1862
rect 604 -1870 605 -1868
rect 611 -1864 612 -1862
rect 611 -1870 612 -1868
rect 618 -1864 619 -1862
rect 618 -1870 619 -1868
rect 628 -1864 629 -1862
rect 625 -1870 626 -1868
rect 628 -1870 629 -1868
rect 632 -1870 633 -1868
rect 642 -1864 643 -1862
rect 642 -1870 643 -1868
rect 646 -1864 647 -1862
rect 646 -1870 647 -1868
rect 653 -1864 654 -1862
rect 653 -1870 654 -1868
rect 660 -1864 661 -1862
rect 660 -1870 661 -1868
rect 663 -1870 664 -1868
rect 667 -1864 668 -1862
rect 667 -1870 668 -1868
rect 674 -1864 675 -1862
rect 674 -1870 675 -1868
rect 681 -1864 682 -1862
rect 681 -1870 682 -1868
rect 688 -1864 689 -1862
rect 688 -1870 689 -1868
rect 695 -1864 696 -1862
rect 695 -1870 696 -1868
rect 702 -1864 703 -1862
rect 702 -1870 703 -1868
rect 709 -1864 710 -1862
rect 709 -1870 710 -1868
rect 716 -1864 717 -1862
rect 716 -1870 717 -1868
rect 726 -1864 727 -1862
rect 723 -1870 724 -1868
rect 726 -1870 727 -1868
rect 730 -1864 731 -1862
rect 730 -1870 731 -1868
rect 737 -1864 738 -1862
rect 737 -1870 738 -1868
rect 744 -1864 745 -1862
rect 744 -1870 745 -1868
rect 751 -1864 752 -1862
rect 751 -1870 752 -1868
rect 758 -1864 759 -1862
rect 758 -1870 759 -1868
rect 765 -1864 766 -1862
rect 765 -1870 766 -1868
rect 772 -1864 773 -1862
rect 772 -1870 773 -1868
rect 779 -1864 780 -1862
rect 779 -1870 780 -1868
rect 786 -1864 787 -1862
rect 786 -1870 787 -1868
rect 793 -1864 794 -1862
rect 793 -1870 794 -1868
rect 800 -1864 801 -1862
rect 800 -1870 801 -1868
rect 807 -1864 808 -1862
rect 807 -1870 808 -1868
rect 814 -1864 815 -1862
rect 814 -1870 815 -1868
rect 817 -1870 818 -1868
rect 821 -1864 822 -1862
rect 821 -1870 822 -1868
rect 828 -1864 829 -1862
rect 828 -1870 829 -1868
rect 835 -1864 836 -1862
rect 838 -1864 839 -1862
rect 842 -1864 843 -1862
rect 845 -1864 846 -1862
rect 845 -1870 846 -1868
rect 849 -1864 850 -1862
rect 852 -1864 853 -1862
rect 856 -1864 857 -1862
rect 856 -1870 857 -1868
rect 863 -1864 864 -1862
rect 863 -1870 864 -1868
rect 870 -1864 871 -1862
rect 870 -1870 871 -1868
rect 877 -1864 878 -1862
rect 877 -1870 878 -1868
rect 898 -1864 899 -1862
rect 898 -1870 899 -1868
rect 915 -1864 916 -1862
rect 947 -1864 948 -1862
rect 950 -1864 951 -1862
rect 16 -1935 17 -1933
rect 16 -1941 17 -1939
rect 23 -1935 24 -1933
rect 23 -1941 24 -1939
rect 33 -1941 34 -1939
rect 37 -1941 38 -1939
rect 40 -1941 41 -1939
rect 44 -1935 45 -1933
rect 47 -1941 48 -1939
rect 51 -1935 52 -1933
rect 51 -1941 52 -1939
rect 58 -1935 59 -1933
rect 58 -1941 59 -1939
rect 65 -1935 66 -1933
rect 65 -1941 66 -1939
rect 72 -1935 73 -1933
rect 72 -1941 73 -1939
rect 79 -1935 80 -1933
rect 79 -1941 80 -1939
rect 86 -1935 87 -1933
rect 86 -1941 87 -1939
rect 93 -1935 94 -1933
rect 93 -1941 94 -1939
rect 100 -1935 101 -1933
rect 100 -1941 101 -1939
rect 107 -1935 108 -1933
rect 107 -1941 108 -1939
rect 114 -1935 115 -1933
rect 114 -1941 115 -1939
rect 121 -1935 122 -1933
rect 124 -1935 125 -1933
rect 128 -1935 129 -1933
rect 128 -1941 129 -1939
rect 135 -1935 136 -1933
rect 135 -1941 136 -1939
rect 142 -1935 143 -1933
rect 145 -1935 146 -1933
rect 142 -1941 143 -1939
rect 149 -1935 150 -1933
rect 149 -1941 150 -1939
rect 156 -1935 157 -1933
rect 159 -1935 160 -1933
rect 159 -1941 160 -1939
rect 163 -1935 164 -1933
rect 163 -1941 164 -1939
rect 170 -1935 171 -1933
rect 170 -1941 171 -1939
rect 177 -1935 178 -1933
rect 177 -1941 178 -1939
rect 180 -1941 181 -1939
rect 184 -1935 185 -1933
rect 184 -1941 185 -1939
rect 191 -1935 192 -1933
rect 194 -1935 195 -1933
rect 191 -1941 192 -1939
rect 194 -1941 195 -1939
rect 198 -1935 199 -1933
rect 198 -1941 199 -1939
rect 205 -1935 206 -1933
rect 205 -1941 206 -1939
rect 212 -1935 213 -1933
rect 212 -1941 213 -1939
rect 219 -1941 220 -1939
rect 222 -1941 223 -1939
rect 229 -1935 230 -1933
rect 226 -1941 227 -1939
rect 229 -1941 230 -1939
rect 233 -1941 234 -1939
rect 236 -1941 237 -1939
rect 240 -1935 241 -1933
rect 243 -1935 244 -1933
rect 240 -1941 241 -1939
rect 243 -1941 244 -1939
rect 247 -1935 248 -1933
rect 247 -1941 248 -1939
rect 254 -1935 255 -1933
rect 254 -1941 255 -1939
rect 261 -1935 262 -1933
rect 261 -1941 262 -1939
rect 268 -1935 269 -1933
rect 268 -1941 269 -1939
rect 275 -1935 276 -1933
rect 275 -1941 276 -1939
rect 282 -1935 283 -1933
rect 285 -1935 286 -1933
rect 282 -1941 283 -1939
rect 289 -1935 290 -1933
rect 289 -1941 290 -1939
rect 296 -1935 297 -1933
rect 296 -1941 297 -1939
rect 303 -1935 304 -1933
rect 303 -1941 304 -1939
rect 310 -1935 311 -1933
rect 310 -1941 311 -1939
rect 317 -1935 318 -1933
rect 317 -1941 318 -1939
rect 320 -1941 321 -1939
rect 324 -1935 325 -1933
rect 324 -1941 325 -1939
rect 331 -1935 332 -1933
rect 334 -1935 335 -1933
rect 331 -1941 332 -1939
rect 334 -1941 335 -1939
rect 338 -1935 339 -1933
rect 338 -1941 339 -1939
rect 345 -1935 346 -1933
rect 345 -1941 346 -1939
rect 352 -1935 353 -1933
rect 352 -1941 353 -1939
rect 359 -1935 360 -1933
rect 359 -1941 360 -1939
rect 366 -1935 367 -1933
rect 366 -1941 367 -1939
rect 373 -1935 374 -1933
rect 373 -1941 374 -1939
rect 380 -1935 381 -1933
rect 380 -1941 381 -1939
rect 387 -1935 388 -1933
rect 387 -1941 388 -1939
rect 394 -1935 395 -1933
rect 394 -1941 395 -1939
rect 401 -1935 402 -1933
rect 401 -1941 402 -1939
rect 408 -1935 409 -1933
rect 411 -1935 412 -1933
rect 408 -1941 409 -1939
rect 411 -1941 412 -1939
rect 418 -1935 419 -1933
rect 415 -1941 416 -1939
rect 418 -1941 419 -1939
rect 422 -1935 423 -1933
rect 422 -1941 423 -1939
rect 429 -1935 430 -1933
rect 429 -1941 430 -1939
rect 436 -1935 437 -1933
rect 439 -1935 440 -1933
rect 436 -1941 437 -1939
rect 439 -1941 440 -1939
rect 443 -1935 444 -1933
rect 443 -1941 444 -1939
rect 450 -1935 451 -1933
rect 453 -1935 454 -1933
rect 450 -1941 451 -1939
rect 453 -1941 454 -1939
rect 457 -1935 458 -1933
rect 460 -1935 461 -1933
rect 457 -1941 458 -1939
rect 460 -1941 461 -1939
rect 464 -1935 465 -1933
rect 464 -1941 465 -1939
rect 471 -1935 472 -1933
rect 474 -1941 475 -1939
rect 478 -1935 479 -1933
rect 478 -1941 479 -1939
rect 485 -1935 486 -1933
rect 485 -1941 486 -1939
rect 492 -1935 493 -1933
rect 492 -1941 493 -1939
rect 499 -1935 500 -1933
rect 499 -1941 500 -1939
rect 502 -1941 503 -1939
rect 506 -1935 507 -1933
rect 506 -1941 507 -1939
rect 513 -1935 514 -1933
rect 513 -1941 514 -1939
rect 520 -1935 521 -1933
rect 520 -1941 521 -1939
rect 527 -1935 528 -1933
rect 527 -1941 528 -1939
rect 534 -1935 535 -1933
rect 534 -1941 535 -1939
rect 541 -1935 542 -1933
rect 541 -1941 542 -1939
rect 548 -1935 549 -1933
rect 548 -1941 549 -1939
rect 555 -1935 556 -1933
rect 555 -1941 556 -1939
rect 562 -1935 563 -1933
rect 562 -1941 563 -1939
rect 569 -1935 570 -1933
rect 569 -1941 570 -1939
rect 576 -1935 577 -1933
rect 576 -1941 577 -1939
rect 579 -1941 580 -1939
rect 583 -1935 584 -1933
rect 583 -1941 584 -1939
rect 590 -1941 591 -1939
rect 593 -1941 594 -1939
rect 597 -1935 598 -1933
rect 597 -1941 598 -1939
rect 604 -1935 605 -1933
rect 604 -1941 605 -1939
rect 611 -1935 612 -1933
rect 611 -1941 612 -1939
rect 618 -1935 619 -1933
rect 618 -1941 619 -1939
rect 625 -1935 626 -1933
rect 625 -1941 626 -1939
rect 632 -1935 633 -1933
rect 632 -1941 633 -1939
rect 639 -1935 640 -1933
rect 639 -1941 640 -1939
rect 646 -1935 647 -1933
rect 646 -1941 647 -1939
rect 653 -1935 654 -1933
rect 653 -1941 654 -1939
rect 660 -1935 661 -1933
rect 660 -1941 661 -1939
rect 667 -1935 668 -1933
rect 667 -1941 668 -1939
rect 674 -1935 675 -1933
rect 674 -1941 675 -1939
rect 681 -1935 682 -1933
rect 681 -1941 682 -1939
rect 684 -1941 685 -1939
rect 688 -1935 689 -1933
rect 688 -1941 689 -1939
rect 695 -1935 696 -1933
rect 695 -1941 696 -1939
rect 702 -1935 703 -1933
rect 702 -1941 703 -1939
rect 709 -1935 710 -1933
rect 709 -1941 710 -1939
rect 716 -1935 717 -1933
rect 716 -1941 717 -1939
rect 723 -1935 724 -1933
rect 723 -1941 724 -1939
rect 730 -1935 731 -1933
rect 730 -1941 731 -1939
rect 737 -1935 738 -1933
rect 737 -1941 738 -1939
rect 744 -1935 745 -1933
rect 744 -1941 745 -1939
rect 751 -1935 752 -1933
rect 751 -1941 752 -1939
rect 758 -1935 759 -1933
rect 761 -1935 762 -1933
rect 758 -1941 759 -1939
rect 765 -1935 766 -1933
rect 765 -1941 766 -1939
rect 772 -1935 773 -1933
rect 772 -1941 773 -1939
rect 782 -1935 783 -1933
rect 779 -1941 780 -1939
rect 782 -1941 783 -1939
rect 786 -1935 787 -1933
rect 786 -1941 787 -1939
rect 793 -1935 794 -1933
rect 793 -1941 794 -1939
rect 814 -1935 815 -1933
rect 814 -1941 815 -1939
rect 821 -1935 822 -1933
rect 821 -1941 822 -1939
rect 37 -1994 38 -1992
rect 37 -2000 38 -1998
rect 44 -1994 45 -1992
rect 44 -2000 45 -1998
rect 51 -1994 52 -1992
rect 51 -2000 52 -1998
rect 58 -1994 59 -1992
rect 58 -2000 59 -1998
rect 65 -1994 66 -1992
rect 65 -2000 66 -1998
rect 72 -1994 73 -1992
rect 72 -2000 73 -1998
rect 79 -1994 80 -1992
rect 79 -2000 80 -1998
rect 86 -1994 87 -1992
rect 86 -2000 87 -1998
rect 93 -1994 94 -1992
rect 93 -2000 94 -1998
rect 100 -1994 101 -1992
rect 100 -2000 101 -1998
rect 107 -1994 108 -1992
rect 107 -2000 108 -1998
rect 114 -1994 115 -1992
rect 114 -2000 115 -1998
rect 121 -1994 122 -1992
rect 121 -2000 122 -1998
rect 128 -1994 129 -1992
rect 128 -2000 129 -1998
rect 135 -1994 136 -1992
rect 138 -1994 139 -1992
rect 135 -2000 136 -1998
rect 142 -1994 143 -1992
rect 142 -2000 143 -1998
rect 149 -1994 150 -1992
rect 149 -2000 150 -1998
rect 156 -1994 157 -1992
rect 159 -1994 160 -1992
rect 163 -1994 164 -1992
rect 163 -2000 164 -1998
rect 170 -1994 171 -1992
rect 170 -2000 171 -1998
rect 177 -1994 178 -1992
rect 177 -2000 178 -1998
rect 184 -1994 185 -1992
rect 184 -2000 185 -1998
rect 191 -1994 192 -1992
rect 191 -2000 192 -1998
rect 198 -1994 199 -1992
rect 198 -2000 199 -1998
rect 201 -2000 202 -1998
rect 205 -1994 206 -1992
rect 205 -2000 206 -1998
rect 212 -1994 213 -1992
rect 212 -2000 213 -1998
rect 219 -1994 220 -1992
rect 219 -2000 220 -1998
rect 229 -1994 230 -1992
rect 229 -2000 230 -1998
rect 233 -1994 234 -1992
rect 233 -2000 234 -1998
rect 240 -2000 241 -1998
rect 243 -2000 244 -1998
rect 247 -1994 248 -1992
rect 247 -2000 248 -1998
rect 254 -1994 255 -1992
rect 254 -2000 255 -1998
rect 261 -1994 262 -1992
rect 264 -1994 265 -1992
rect 261 -2000 262 -1998
rect 264 -2000 265 -1998
rect 268 -1994 269 -1992
rect 271 -1994 272 -1992
rect 271 -2000 272 -1998
rect 275 -1994 276 -1992
rect 275 -2000 276 -1998
rect 282 -1994 283 -1992
rect 282 -2000 283 -1998
rect 289 -2000 290 -1998
rect 292 -2000 293 -1998
rect 296 -1994 297 -1992
rect 296 -2000 297 -1998
rect 303 -1994 304 -1992
rect 303 -2000 304 -1998
rect 313 -2000 314 -1998
rect 317 -1994 318 -1992
rect 317 -2000 318 -1998
rect 324 -1994 325 -1992
rect 324 -2000 325 -1998
rect 331 -1994 332 -1992
rect 331 -2000 332 -1998
rect 338 -1994 339 -1992
rect 338 -2000 339 -1998
rect 345 -1994 346 -1992
rect 345 -2000 346 -1998
rect 352 -1994 353 -1992
rect 352 -2000 353 -1998
rect 359 -1994 360 -1992
rect 359 -2000 360 -1998
rect 369 -1994 370 -1992
rect 373 -1994 374 -1992
rect 373 -2000 374 -1998
rect 380 -1994 381 -1992
rect 380 -2000 381 -1998
rect 387 -1994 388 -1992
rect 387 -2000 388 -1998
rect 394 -1994 395 -1992
rect 394 -2000 395 -1998
rect 401 -1994 402 -1992
rect 401 -2000 402 -1998
rect 408 -1994 409 -1992
rect 408 -2000 409 -1998
rect 415 -1994 416 -1992
rect 415 -2000 416 -1998
rect 422 -1994 423 -1992
rect 422 -2000 423 -1998
rect 432 -1994 433 -1992
rect 429 -2000 430 -1998
rect 432 -2000 433 -1998
rect 436 -1994 437 -1992
rect 439 -1994 440 -1992
rect 446 -1994 447 -1992
rect 443 -2000 444 -1998
rect 446 -2000 447 -1998
rect 450 -1994 451 -1992
rect 450 -2000 451 -1998
rect 457 -1994 458 -1992
rect 457 -2000 458 -1998
rect 464 -1994 465 -1992
rect 464 -2000 465 -1998
rect 471 -1994 472 -1992
rect 471 -2000 472 -1998
rect 478 -1994 479 -1992
rect 478 -2000 479 -1998
rect 485 -1994 486 -1992
rect 485 -2000 486 -1998
rect 492 -1994 493 -1992
rect 495 -1994 496 -1992
rect 492 -2000 493 -1998
rect 499 -1994 500 -1992
rect 499 -2000 500 -1998
rect 506 -1994 507 -1992
rect 506 -2000 507 -1998
rect 516 -1994 517 -1992
rect 513 -2000 514 -1998
rect 520 -1994 521 -1992
rect 520 -2000 521 -1998
rect 527 -1994 528 -1992
rect 527 -2000 528 -1998
rect 534 -1994 535 -1992
rect 534 -2000 535 -1998
rect 541 -1994 542 -1992
rect 541 -2000 542 -1998
rect 548 -1994 549 -1992
rect 548 -2000 549 -1998
rect 555 -1994 556 -1992
rect 555 -2000 556 -1998
rect 562 -1994 563 -1992
rect 562 -2000 563 -1998
rect 569 -1994 570 -1992
rect 569 -2000 570 -1998
rect 576 -1994 577 -1992
rect 576 -2000 577 -1998
rect 583 -2000 584 -1998
rect 586 -2000 587 -1998
rect 593 -1994 594 -1992
rect 590 -2000 591 -1998
rect 593 -2000 594 -1998
rect 597 -1994 598 -1992
rect 597 -2000 598 -1998
rect 600 -2000 601 -1998
rect 604 -1994 605 -1992
rect 604 -2000 605 -1998
rect 611 -1994 612 -1992
rect 611 -2000 612 -1998
rect 618 -1994 619 -1992
rect 618 -2000 619 -1998
rect 625 -1994 626 -1992
rect 625 -2000 626 -1998
rect 632 -1994 633 -1992
rect 632 -2000 633 -1998
rect 639 -1994 640 -1992
rect 639 -2000 640 -1998
rect 646 -1994 647 -1992
rect 646 -2000 647 -1998
rect 653 -1994 654 -1992
rect 653 -2000 654 -1998
rect 660 -2000 661 -1998
rect 663 -2000 664 -1998
rect 667 -1994 668 -1992
rect 667 -2000 668 -1998
rect 674 -1994 675 -1992
rect 677 -1994 678 -1992
rect 674 -2000 675 -1998
rect 677 -2000 678 -1998
rect 681 -1994 682 -1992
rect 681 -2000 682 -1998
rect 688 -1994 689 -1992
rect 691 -2000 692 -1998
rect 695 -1994 696 -1992
rect 695 -2000 696 -1998
rect 702 -1994 703 -1992
rect 702 -2000 703 -1998
rect 709 -1994 710 -1992
rect 709 -2000 710 -1998
rect 716 -1994 717 -1992
rect 716 -2000 717 -1998
rect 723 -1994 724 -1992
rect 726 -1994 727 -1992
rect 730 -1994 731 -1992
rect 730 -2000 731 -1998
rect 737 -1994 738 -1992
rect 737 -2000 738 -1998
rect 744 -1994 745 -1992
rect 744 -2000 745 -1998
rect 751 -1994 752 -1992
rect 751 -2000 752 -1998
rect 758 -1994 759 -1992
rect 758 -2000 759 -1998
rect 765 -1994 766 -1992
rect 765 -2000 766 -1998
rect 772 -1994 773 -1992
rect 772 -2000 773 -1998
rect 779 -1994 780 -1992
rect 786 -1994 787 -1992
rect 786 -2000 787 -1998
rect 793 -2000 794 -1998
rect 796 -2000 797 -1998
rect 800 -1994 801 -1992
rect 800 -2000 801 -1998
rect 807 -1994 808 -1992
rect 807 -2000 808 -1998
rect 814 -1994 815 -1992
rect 814 -2000 815 -1998
rect 16 -2057 17 -2055
rect 16 -2063 17 -2061
rect 23 -2057 24 -2055
rect 23 -2063 24 -2061
rect 30 -2057 31 -2055
rect 30 -2063 31 -2061
rect 37 -2057 38 -2055
rect 37 -2063 38 -2061
rect 44 -2057 45 -2055
rect 44 -2063 45 -2061
rect 51 -2057 52 -2055
rect 51 -2063 52 -2061
rect 58 -2057 59 -2055
rect 58 -2063 59 -2061
rect 65 -2057 66 -2055
rect 65 -2063 66 -2061
rect 72 -2057 73 -2055
rect 72 -2063 73 -2061
rect 79 -2057 80 -2055
rect 79 -2063 80 -2061
rect 86 -2057 87 -2055
rect 86 -2063 87 -2061
rect 93 -2057 94 -2055
rect 93 -2063 94 -2061
rect 100 -2057 101 -2055
rect 100 -2063 101 -2061
rect 107 -2057 108 -2055
rect 107 -2063 108 -2061
rect 114 -2057 115 -2055
rect 114 -2063 115 -2061
rect 121 -2057 122 -2055
rect 124 -2063 125 -2061
rect 128 -2057 129 -2055
rect 128 -2063 129 -2061
rect 131 -2063 132 -2061
rect 135 -2057 136 -2055
rect 135 -2063 136 -2061
rect 142 -2057 143 -2055
rect 142 -2063 143 -2061
rect 145 -2063 146 -2061
rect 149 -2057 150 -2055
rect 149 -2063 150 -2061
rect 156 -2057 157 -2055
rect 156 -2063 157 -2061
rect 166 -2057 167 -2055
rect 163 -2063 164 -2061
rect 170 -2057 171 -2055
rect 170 -2063 171 -2061
rect 177 -2063 178 -2061
rect 180 -2063 181 -2061
rect 184 -2057 185 -2055
rect 187 -2057 188 -2055
rect 184 -2063 185 -2061
rect 187 -2063 188 -2061
rect 191 -2057 192 -2055
rect 191 -2063 192 -2061
rect 198 -2057 199 -2055
rect 198 -2063 199 -2061
rect 205 -2057 206 -2055
rect 205 -2063 206 -2061
rect 212 -2057 213 -2055
rect 212 -2063 213 -2061
rect 219 -2057 220 -2055
rect 219 -2063 220 -2061
rect 226 -2057 227 -2055
rect 229 -2057 230 -2055
rect 229 -2063 230 -2061
rect 233 -2057 234 -2055
rect 236 -2057 237 -2055
rect 233 -2063 234 -2061
rect 236 -2063 237 -2061
rect 243 -2057 244 -2055
rect 240 -2063 241 -2061
rect 243 -2063 244 -2061
rect 247 -2057 248 -2055
rect 247 -2063 248 -2061
rect 254 -2057 255 -2055
rect 257 -2057 258 -2055
rect 254 -2063 255 -2061
rect 257 -2063 258 -2061
rect 261 -2057 262 -2055
rect 261 -2063 262 -2061
rect 268 -2057 269 -2055
rect 268 -2063 269 -2061
rect 275 -2057 276 -2055
rect 275 -2063 276 -2061
rect 282 -2057 283 -2055
rect 282 -2063 283 -2061
rect 289 -2057 290 -2055
rect 289 -2063 290 -2061
rect 296 -2057 297 -2055
rect 296 -2063 297 -2061
rect 303 -2057 304 -2055
rect 303 -2063 304 -2061
rect 310 -2057 311 -2055
rect 310 -2063 311 -2061
rect 317 -2057 318 -2055
rect 317 -2063 318 -2061
rect 324 -2057 325 -2055
rect 324 -2063 325 -2061
rect 331 -2057 332 -2055
rect 331 -2063 332 -2061
rect 338 -2057 339 -2055
rect 338 -2063 339 -2061
rect 345 -2057 346 -2055
rect 348 -2057 349 -2055
rect 345 -2063 346 -2061
rect 352 -2057 353 -2055
rect 352 -2063 353 -2061
rect 359 -2057 360 -2055
rect 359 -2063 360 -2061
rect 366 -2057 367 -2055
rect 366 -2063 367 -2061
rect 373 -2057 374 -2055
rect 373 -2063 374 -2061
rect 380 -2057 381 -2055
rect 380 -2063 381 -2061
rect 387 -2057 388 -2055
rect 387 -2063 388 -2061
rect 394 -2057 395 -2055
rect 397 -2057 398 -2055
rect 394 -2063 395 -2061
rect 397 -2063 398 -2061
rect 401 -2057 402 -2055
rect 404 -2057 405 -2055
rect 408 -2057 409 -2055
rect 408 -2063 409 -2061
rect 415 -2057 416 -2055
rect 418 -2057 419 -2055
rect 415 -2063 416 -2061
rect 418 -2063 419 -2061
rect 422 -2057 423 -2055
rect 422 -2063 423 -2061
rect 432 -2057 433 -2055
rect 432 -2063 433 -2061
rect 436 -2057 437 -2055
rect 436 -2063 437 -2061
rect 443 -2057 444 -2055
rect 443 -2063 444 -2061
rect 450 -2057 451 -2055
rect 450 -2063 451 -2061
rect 457 -2057 458 -2055
rect 460 -2057 461 -2055
rect 457 -2063 458 -2061
rect 460 -2063 461 -2061
rect 464 -2057 465 -2055
rect 464 -2063 465 -2061
rect 474 -2057 475 -2055
rect 471 -2063 472 -2061
rect 474 -2063 475 -2061
rect 478 -2057 479 -2055
rect 478 -2063 479 -2061
rect 488 -2057 489 -2055
rect 485 -2063 486 -2061
rect 488 -2063 489 -2061
rect 492 -2057 493 -2055
rect 492 -2063 493 -2061
rect 499 -2057 500 -2055
rect 499 -2063 500 -2061
rect 506 -2063 507 -2061
rect 509 -2063 510 -2061
rect 513 -2057 514 -2055
rect 513 -2063 514 -2061
rect 516 -2063 517 -2061
rect 520 -2057 521 -2055
rect 520 -2063 521 -2061
rect 527 -2057 528 -2055
rect 527 -2063 528 -2061
rect 534 -2057 535 -2055
rect 534 -2063 535 -2061
rect 541 -2057 542 -2055
rect 541 -2063 542 -2061
rect 548 -2057 549 -2055
rect 548 -2063 549 -2061
rect 555 -2057 556 -2055
rect 555 -2063 556 -2061
rect 565 -2057 566 -2055
rect 562 -2063 563 -2061
rect 569 -2057 570 -2055
rect 569 -2063 570 -2061
rect 576 -2057 577 -2055
rect 576 -2063 577 -2061
rect 583 -2057 584 -2055
rect 583 -2063 584 -2061
rect 590 -2057 591 -2055
rect 590 -2063 591 -2061
rect 597 -2057 598 -2055
rect 597 -2063 598 -2061
rect 604 -2057 605 -2055
rect 604 -2063 605 -2061
rect 611 -2057 612 -2055
rect 611 -2063 612 -2061
rect 618 -2057 619 -2055
rect 618 -2063 619 -2061
rect 625 -2057 626 -2055
rect 625 -2063 626 -2061
rect 632 -2057 633 -2055
rect 632 -2063 633 -2061
rect 639 -2057 640 -2055
rect 639 -2063 640 -2061
rect 646 -2057 647 -2055
rect 646 -2063 647 -2061
rect 653 -2057 654 -2055
rect 660 -2057 661 -2055
rect 660 -2063 661 -2061
rect 667 -2057 668 -2055
rect 670 -2057 671 -2055
rect 670 -2063 671 -2061
rect 674 -2057 675 -2055
rect 674 -2063 675 -2061
rect 681 -2057 682 -2055
rect 681 -2063 682 -2061
rect 688 -2057 689 -2055
rect 688 -2063 689 -2061
rect 695 -2057 696 -2055
rect 695 -2063 696 -2061
rect 702 -2057 703 -2055
rect 702 -2063 703 -2061
rect 709 -2057 710 -2055
rect 709 -2063 710 -2061
rect 716 -2057 717 -2055
rect 716 -2063 717 -2061
rect 726 -2057 727 -2055
rect 723 -2063 724 -2061
rect 726 -2063 727 -2061
rect 730 -2057 731 -2055
rect 730 -2063 731 -2061
rect 737 -2057 738 -2055
rect 737 -2063 738 -2061
rect 744 -2057 745 -2055
rect 744 -2063 745 -2061
rect 751 -2057 752 -2055
rect 751 -2063 752 -2061
rect 758 -2057 759 -2055
rect 758 -2063 759 -2061
rect 765 -2057 766 -2055
rect 765 -2063 766 -2061
rect 772 -2057 773 -2055
rect 772 -2063 773 -2061
rect 779 -2057 780 -2055
rect 779 -2063 780 -2061
rect 786 -2057 787 -2055
rect 786 -2063 787 -2061
rect 16 -2122 17 -2120
rect 16 -2128 17 -2126
rect 23 -2122 24 -2120
rect 23 -2128 24 -2126
rect 30 -2122 31 -2120
rect 30 -2128 31 -2126
rect 40 -2128 41 -2126
rect 44 -2122 45 -2120
rect 44 -2128 45 -2126
rect 51 -2122 52 -2120
rect 51 -2128 52 -2126
rect 58 -2122 59 -2120
rect 58 -2128 59 -2126
rect 65 -2122 66 -2120
rect 65 -2128 66 -2126
rect 72 -2122 73 -2120
rect 72 -2128 73 -2126
rect 79 -2122 80 -2120
rect 79 -2128 80 -2126
rect 86 -2122 87 -2120
rect 86 -2128 87 -2126
rect 93 -2122 94 -2120
rect 96 -2122 97 -2120
rect 103 -2122 104 -2120
rect 100 -2128 101 -2126
rect 107 -2122 108 -2120
rect 107 -2128 108 -2126
rect 114 -2122 115 -2120
rect 114 -2128 115 -2126
rect 121 -2122 122 -2120
rect 121 -2128 122 -2126
rect 128 -2122 129 -2120
rect 128 -2128 129 -2126
rect 135 -2122 136 -2120
rect 138 -2122 139 -2120
rect 135 -2128 136 -2126
rect 142 -2122 143 -2120
rect 142 -2128 143 -2126
rect 149 -2122 150 -2120
rect 149 -2128 150 -2126
rect 156 -2122 157 -2120
rect 156 -2128 157 -2126
rect 159 -2128 160 -2126
rect 163 -2122 164 -2120
rect 163 -2128 164 -2126
rect 173 -2122 174 -2120
rect 170 -2128 171 -2126
rect 173 -2128 174 -2126
rect 177 -2122 178 -2120
rect 180 -2122 181 -2120
rect 177 -2128 178 -2126
rect 180 -2128 181 -2126
rect 184 -2122 185 -2120
rect 191 -2122 192 -2120
rect 191 -2128 192 -2126
rect 198 -2122 199 -2120
rect 198 -2128 199 -2126
rect 201 -2128 202 -2126
rect 205 -2122 206 -2120
rect 205 -2128 206 -2126
rect 208 -2128 209 -2126
rect 212 -2122 213 -2120
rect 212 -2128 213 -2126
rect 219 -2122 220 -2120
rect 219 -2128 220 -2126
rect 222 -2128 223 -2126
rect 229 -2122 230 -2120
rect 226 -2128 227 -2126
rect 233 -2122 234 -2120
rect 233 -2128 234 -2126
rect 240 -2122 241 -2120
rect 240 -2128 241 -2126
rect 247 -2122 248 -2120
rect 250 -2128 251 -2126
rect 254 -2122 255 -2120
rect 254 -2128 255 -2126
rect 261 -2122 262 -2120
rect 261 -2128 262 -2126
rect 268 -2122 269 -2120
rect 268 -2128 269 -2126
rect 275 -2122 276 -2120
rect 275 -2128 276 -2126
rect 282 -2122 283 -2120
rect 282 -2128 283 -2126
rect 289 -2122 290 -2120
rect 292 -2122 293 -2120
rect 296 -2122 297 -2120
rect 296 -2128 297 -2126
rect 303 -2122 304 -2120
rect 303 -2128 304 -2126
rect 310 -2122 311 -2120
rect 310 -2128 311 -2126
rect 317 -2122 318 -2120
rect 320 -2122 321 -2120
rect 320 -2128 321 -2126
rect 324 -2122 325 -2120
rect 324 -2128 325 -2126
rect 331 -2122 332 -2120
rect 331 -2128 332 -2126
rect 338 -2122 339 -2120
rect 338 -2128 339 -2126
rect 348 -2122 349 -2120
rect 345 -2128 346 -2126
rect 348 -2128 349 -2126
rect 352 -2122 353 -2120
rect 352 -2128 353 -2126
rect 362 -2122 363 -2120
rect 362 -2128 363 -2126
rect 366 -2122 367 -2120
rect 366 -2128 367 -2126
rect 373 -2122 374 -2120
rect 373 -2128 374 -2126
rect 383 -2122 384 -2120
rect 380 -2128 381 -2126
rect 387 -2122 388 -2120
rect 387 -2128 388 -2126
rect 394 -2122 395 -2120
rect 394 -2128 395 -2126
rect 401 -2122 402 -2120
rect 401 -2128 402 -2126
rect 411 -2122 412 -2120
rect 408 -2128 409 -2126
rect 411 -2128 412 -2126
rect 415 -2122 416 -2120
rect 415 -2128 416 -2126
rect 422 -2122 423 -2120
rect 422 -2128 423 -2126
rect 429 -2122 430 -2120
rect 429 -2128 430 -2126
rect 439 -2122 440 -2120
rect 439 -2128 440 -2126
rect 443 -2122 444 -2120
rect 443 -2128 444 -2126
rect 450 -2122 451 -2120
rect 450 -2128 451 -2126
rect 457 -2122 458 -2120
rect 460 -2122 461 -2120
rect 464 -2122 465 -2120
rect 464 -2128 465 -2126
rect 467 -2128 468 -2126
rect 474 -2122 475 -2120
rect 471 -2128 472 -2126
rect 474 -2128 475 -2126
rect 478 -2122 479 -2120
rect 478 -2128 479 -2126
rect 485 -2122 486 -2120
rect 485 -2128 486 -2126
rect 492 -2122 493 -2120
rect 492 -2128 493 -2126
rect 499 -2122 500 -2120
rect 499 -2128 500 -2126
rect 506 -2122 507 -2120
rect 506 -2128 507 -2126
rect 509 -2128 510 -2126
rect 513 -2122 514 -2120
rect 513 -2128 514 -2126
rect 520 -2122 521 -2120
rect 520 -2128 521 -2126
rect 527 -2122 528 -2120
rect 527 -2128 528 -2126
rect 534 -2122 535 -2120
rect 534 -2128 535 -2126
rect 541 -2122 542 -2120
rect 541 -2128 542 -2126
rect 548 -2122 549 -2120
rect 548 -2128 549 -2126
rect 555 -2122 556 -2120
rect 555 -2128 556 -2126
rect 562 -2122 563 -2120
rect 562 -2128 563 -2126
rect 569 -2122 570 -2120
rect 569 -2128 570 -2126
rect 576 -2122 577 -2120
rect 576 -2128 577 -2126
rect 583 -2122 584 -2120
rect 583 -2128 584 -2126
rect 593 -2122 594 -2120
rect 593 -2128 594 -2126
rect 597 -2122 598 -2120
rect 597 -2128 598 -2126
rect 604 -2122 605 -2120
rect 604 -2128 605 -2126
rect 611 -2122 612 -2120
rect 611 -2128 612 -2126
rect 618 -2122 619 -2120
rect 618 -2128 619 -2126
rect 625 -2122 626 -2120
rect 625 -2128 626 -2126
rect 632 -2122 633 -2120
rect 632 -2128 633 -2126
rect 639 -2122 640 -2120
rect 639 -2128 640 -2126
rect 646 -2122 647 -2120
rect 646 -2128 647 -2126
rect 653 -2122 654 -2120
rect 653 -2128 654 -2126
rect 660 -2122 661 -2120
rect 660 -2128 661 -2126
rect 667 -2122 668 -2120
rect 667 -2128 668 -2126
rect 674 -2122 675 -2120
rect 674 -2128 675 -2126
rect 681 -2122 682 -2120
rect 681 -2128 682 -2126
rect 688 -2122 689 -2120
rect 688 -2128 689 -2126
rect 695 -2122 696 -2120
rect 695 -2128 696 -2126
rect 702 -2122 703 -2120
rect 702 -2128 703 -2126
rect 709 -2122 710 -2120
rect 709 -2128 710 -2126
rect 716 -2122 717 -2120
rect 716 -2128 717 -2126
rect 723 -2122 724 -2120
rect 723 -2128 724 -2126
rect 730 -2128 731 -2126
rect 737 -2122 738 -2120
rect 737 -2128 738 -2126
rect 86 -2173 87 -2171
rect 86 -2179 87 -2177
rect 100 -2173 101 -2171
rect 100 -2179 101 -2177
rect 107 -2173 108 -2171
rect 107 -2179 108 -2177
rect 114 -2173 115 -2171
rect 114 -2179 115 -2177
rect 121 -2173 122 -2171
rect 121 -2179 122 -2177
rect 128 -2173 129 -2171
rect 128 -2179 129 -2177
rect 131 -2179 132 -2177
rect 135 -2173 136 -2171
rect 142 -2173 143 -2171
rect 142 -2179 143 -2177
rect 152 -2173 153 -2171
rect 152 -2179 153 -2177
rect 156 -2173 157 -2171
rect 159 -2173 160 -2171
rect 156 -2179 157 -2177
rect 163 -2173 164 -2171
rect 163 -2179 164 -2177
rect 170 -2173 171 -2171
rect 170 -2179 171 -2177
rect 177 -2173 178 -2171
rect 177 -2179 178 -2177
rect 184 -2173 185 -2171
rect 184 -2179 185 -2177
rect 191 -2173 192 -2171
rect 191 -2179 192 -2177
rect 198 -2173 199 -2171
rect 198 -2179 199 -2177
rect 205 -2173 206 -2171
rect 205 -2179 206 -2177
rect 212 -2173 213 -2171
rect 212 -2179 213 -2177
rect 219 -2173 220 -2171
rect 222 -2173 223 -2171
rect 219 -2179 220 -2177
rect 222 -2179 223 -2177
rect 226 -2173 227 -2171
rect 229 -2173 230 -2171
rect 233 -2173 234 -2171
rect 233 -2179 234 -2177
rect 240 -2179 241 -2177
rect 243 -2179 244 -2177
rect 247 -2173 248 -2171
rect 247 -2179 248 -2177
rect 254 -2173 255 -2171
rect 254 -2179 255 -2177
rect 261 -2173 262 -2171
rect 261 -2179 262 -2177
rect 268 -2173 269 -2171
rect 268 -2179 269 -2177
rect 275 -2173 276 -2171
rect 275 -2179 276 -2177
rect 282 -2173 283 -2171
rect 285 -2173 286 -2171
rect 282 -2179 283 -2177
rect 285 -2179 286 -2177
rect 289 -2173 290 -2171
rect 289 -2179 290 -2177
rect 296 -2173 297 -2171
rect 299 -2179 300 -2177
rect 303 -2173 304 -2171
rect 303 -2179 304 -2177
rect 310 -2173 311 -2171
rect 313 -2173 314 -2171
rect 310 -2179 311 -2177
rect 317 -2173 318 -2171
rect 317 -2179 318 -2177
rect 324 -2173 325 -2171
rect 324 -2179 325 -2177
rect 331 -2173 332 -2171
rect 334 -2173 335 -2171
rect 331 -2179 332 -2177
rect 338 -2173 339 -2171
rect 338 -2179 339 -2177
rect 345 -2173 346 -2171
rect 345 -2179 346 -2177
rect 352 -2173 353 -2171
rect 352 -2179 353 -2177
rect 359 -2173 360 -2171
rect 359 -2179 360 -2177
rect 366 -2173 367 -2171
rect 366 -2179 367 -2177
rect 373 -2173 374 -2171
rect 373 -2179 374 -2177
rect 380 -2173 381 -2171
rect 380 -2179 381 -2177
rect 387 -2173 388 -2171
rect 390 -2173 391 -2171
rect 390 -2179 391 -2177
rect 394 -2173 395 -2171
rect 394 -2179 395 -2177
rect 401 -2173 402 -2171
rect 401 -2179 402 -2177
rect 408 -2173 409 -2171
rect 411 -2179 412 -2177
rect 415 -2173 416 -2171
rect 415 -2179 416 -2177
rect 422 -2173 423 -2171
rect 422 -2179 423 -2177
rect 429 -2173 430 -2171
rect 429 -2179 430 -2177
rect 432 -2179 433 -2177
rect 436 -2173 437 -2171
rect 436 -2179 437 -2177
rect 443 -2173 444 -2171
rect 443 -2179 444 -2177
rect 453 -2173 454 -2171
rect 450 -2179 451 -2177
rect 457 -2173 458 -2171
rect 460 -2179 461 -2177
rect 464 -2173 465 -2171
rect 464 -2179 465 -2177
rect 471 -2173 472 -2171
rect 471 -2179 472 -2177
rect 478 -2173 479 -2171
rect 478 -2179 479 -2177
rect 485 -2173 486 -2171
rect 485 -2179 486 -2177
rect 492 -2179 493 -2177
rect 499 -2173 500 -2171
rect 499 -2179 500 -2177
rect 509 -2173 510 -2171
rect 509 -2179 510 -2177
rect 513 -2173 514 -2171
rect 513 -2179 514 -2177
rect 520 -2173 521 -2171
rect 520 -2179 521 -2177
rect 527 -2173 528 -2171
rect 527 -2179 528 -2177
rect 534 -2173 535 -2171
rect 534 -2179 535 -2177
rect 541 -2173 542 -2171
rect 541 -2179 542 -2177
rect 548 -2173 549 -2171
rect 548 -2179 549 -2177
rect 555 -2173 556 -2171
rect 558 -2173 559 -2171
rect 555 -2179 556 -2177
rect 558 -2179 559 -2177
rect 562 -2173 563 -2171
rect 562 -2179 563 -2177
rect 569 -2173 570 -2171
rect 569 -2179 570 -2177
rect 576 -2173 577 -2171
rect 579 -2173 580 -2171
rect 576 -2179 577 -2177
rect 583 -2179 584 -2177
rect 586 -2179 587 -2177
rect 590 -2173 591 -2171
rect 590 -2179 591 -2177
rect 597 -2173 598 -2171
rect 597 -2179 598 -2177
rect 604 -2173 605 -2171
rect 604 -2179 605 -2177
rect 611 -2173 612 -2171
rect 611 -2179 612 -2177
rect 618 -2173 619 -2171
rect 618 -2179 619 -2177
rect 625 -2173 626 -2171
rect 625 -2179 626 -2177
rect 632 -2173 633 -2171
rect 632 -2179 633 -2177
rect 639 -2173 640 -2171
rect 639 -2179 640 -2177
rect 646 -2173 647 -2171
rect 646 -2179 647 -2177
rect 653 -2173 654 -2171
rect 653 -2179 654 -2177
rect 660 -2173 661 -2171
rect 660 -2179 661 -2177
rect 667 -2173 668 -2171
rect 667 -2179 668 -2177
rect 670 -2179 671 -2177
rect 674 -2173 675 -2171
rect 674 -2179 675 -2177
rect 681 -2179 682 -2177
rect 688 -2173 689 -2171
rect 688 -2179 689 -2177
rect 695 -2173 696 -2171
rect 698 -2173 699 -2171
rect 702 -2173 703 -2171
rect 702 -2179 703 -2177
rect 709 -2173 710 -2171
rect 709 -2179 710 -2177
rect 716 -2173 717 -2171
rect 716 -2179 717 -2177
rect 723 -2173 724 -2171
rect 723 -2179 724 -2177
rect 89 -2226 90 -2224
rect 107 -2226 108 -2224
rect 107 -2232 108 -2230
rect 114 -2226 115 -2224
rect 114 -2232 115 -2230
rect 124 -2226 125 -2224
rect 124 -2232 125 -2230
rect 131 -2226 132 -2224
rect 128 -2232 129 -2230
rect 138 -2232 139 -2230
rect 142 -2226 143 -2224
rect 142 -2232 143 -2230
rect 149 -2226 150 -2224
rect 149 -2232 150 -2230
rect 156 -2226 157 -2224
rect 156 -2232 157 -2230
rect 163 -2232 164 -2230
rect 166 -2232 167 -2230
rect 170 -2226 171 -2224
rect 173 -2232 174 -2230
rect 177 -2226 178 -2224
rect 177 -2232 178 -2230
rect 180 -2232 181 -2230
rect 184 -2226 185 -2224
rect 184 -2232 185 -2230
rect 191 -2226 192 -2224
rect 191 -2232 192 -2230
rect 201 -2232 202 -2230
rect 205 -2226 206 -2224
rect 208 -2232 209 -2230
rect 212 -2226 213 -2224
rect 212 -2232 213 -2230
rect 219 -2226 220 -2224
rect 219 -2232 220 -2230
rect 226 -2232 227 -2230
rect 229 -2232 230 -2230
rect 233 -2226 234 -2224
rect 233 -2232 234 -2230
rect 240 -2226 241 -2224
rect 240 -2232 241 -2230
rect 247 -2226 248 -2224
rect 247 -2232 248 -2230
rect 254 -2226 255 -2224
rect 254 -2232 255 -2230
rect 261 -2226 262 -2224
rect 261 -2232 262 -2230
rect 268 -2226 269 -2224
rect 268 -2232 269 -2230
rect 275 -2226 276 -2224
rect 275 -2232 276 -2230
rect 285 -2226 286 -2224
rect 282 -2232 283 -2230
rect 289 -2226 290 -2224
rect 289 -2232 290 -2230
rect 296 -2226 297 -2224
rect 296 -2232 297 -2230
rect 306 -2226 307 -2224
rect 303 -2232 304 -2230
rect 306 -2232 307 -2230
rect 310 -2226 311 -2224
rect 310 -2232 311 -2230
rect 317 -2226 318 -2224
rect 317 -2232 318 -2230
rect 324 -2226 325 -2224
rect 324 -2232 325 -2230
rect 331 -2226 332 -2224
rect 331 -2232 332 -2230
rect 338 -2226 339 -2224
rect 338 -2232 339 -2230
rect 345 -2226 346 -2224
rect 345 -2232 346 -2230
rect 352 -2226 353 -2224
rect 352 -2232 353 -2230
rect 359 -2232 360 -2230
rect 366 -2226 367 -2224
rect 366 -2232 367 -2230
rect 373 -2232 374 -2230
rect 376 -2232 377 -2230
rect 380 -2226 381 -2224
rect 380 -2232 381 -2230
rect 387 -2226 388 -2224
rect 390 -2226 391 -2224
rect 390 -2232 391 -2230
rect 394 -2226 395 -2224
rect 394 -2232 395 -2230
rect 401 -2226 402 -2224
rect 401 -2232 402 -2230
rect 408 -2226 409 -2224
rect 408 -2232 409 -2230
rect 415 -2226 416 -2224
rect 415 -2232 416 -2230
rect 425 -2226 426 -2224
rect 425 -2232 426 -2230
rect 429 -2226 430 -2224
rect 429 -2232 430 -2230
rect 436 -2226 437 -2224
rect 436 -2232 437 -2230
rect 443 -2232 444 -2230
rect 446 -2232 447 -2230
rect 450 -2226 451 -2224
rect 450 -2232 451 -2230
rect 457 -2226 458 -2224
rect 457 -2232 458 -2230
rect 464 -2226 465 -2224
rect 464 -2232 465 -2230
rect 467 -2232 468 -2230
rect 471 -2226 472 -2224
rect 471 -2232 472 -2230
rect 478 -2226 479 -2224
rect 478 -2232 479 -2230
rect 485 -2226 486 -2224
rect 485 -2232 486 -2230
rect 492 -2226 493 -2224
rect 492 -2232 493 -2230
rect 499 -2226 500 -2224
rect 499 -2232 500 -2230
rect 506 -2226 507 -2224
rect 506 -2232 507 -2230
rect 513 -2226 514 -2224
rect 513 -2232 514 -2230
rect 520 -2226 521 -2224
rect 520 -2232 521 -2230
rect 527 -2226 528 -2224
rect 527 -2232 528 -2230
rect 534 -2226 535 -2224
rect 534 -2232 535 -2230
rect 541 -2226 542 -2224
rect 541 -2232 542 -2230
rect 548 -2226 549 -2224
rect 548 -2232 549 -2230
rect 555 -2226 556 -2224
rect 555 -2232 556 -2230
rect 562 -2226 563 -2224
rect 565 -2232 566 -2230
rect 569 -2226 570 -2224
rect 569 -2232 570 -2230
rect 579 -2226 580 -2224
rect 576 -2232 577 -2230
rect 579 -2232 580 -2230
rect 583 -2226 584 -2224
rect 583 -2232 584 -2230
rect 590 -2226 591 -2224
rect 590 -2232 591 -2230
rect 597 -2226 598 -2224
rect 597 -2232 598 -2230
rect 604 -2226 605 -2224
rect 607 -2232 608 -2230
rect 614 -2226 615 -2224
rect 611 -2232 612 -2230
rect 618 -2226 619 -2224
rect 621 -2226 622 -2224
rect 625 -2226 626 -2224
rect 632 -2226 633 -2224
rect 632 -2232 633 -2230
rect 639 -2226 640 -2224
rect 639 -2232 640 -2230
rect 660 -2226 661 -2224
rect 660 -2232 661 -2230
rect 114 -2263 115 -2261
rect 114 -2269 115 -2267
rect 121 -2263 122 -2261
rect 124 -2263 125 -2261
rect 124 -2269 125 -2267
rect 131 -2263 132 -2261
rect 131 -2269 132 -2267
rect 135 -2263 136 -2261
rect 135 -2269 136 -2267
rect 145 -2263 146 -2261
rect 142 -2269 143 -2267
rect 145 -2269 146 -2267
rect 149 -2263 150 -2261
rect 156 -2263 157 -2261
rect 156 -2269 157 -2267
rect 163 -2263 164 -2261
rect 163 -2269 164 -2267
rect 170 -2263 171 -2261
rect 170 -2269 171 -2267
rect 177 -2263 178 -2261
rect 177 -2269 178 -2267
rect 184 -2263 185 -2261
rect 184 -2269 185 -2267
rect 191 -2263 192 -2261
rect 194 -2263 195 -2261
rect 198 -2263 199 -2261
rect 198 -2269 199 -2267
rect 205 -2263 206 -2261
rect 205 -2269 206 -2267
rect 212 -2263 213 -2261
rect 212 -2269 213 -2267
rect 215 -2269 216 -2267
rect 219 -2263 220 -2261
rect 219 -2269 220 -2267
rect 226 -2263 227 -2261
rect 226 -2269 227 -2267
rect 236 -2263 237 -2261
rect 233 -2269 234 -2267
rect 240 -2263 241 -2261
rect 243 -2269 244 -2267
rect 247 -2263 248 -2261
rect 247 -2269 248 -2267
rect 254 -2263 255 -2261
rect 254 -2269 255 -2267
rect 261 -2263 262 -2261
rect 261 -2269 262 -2267
rect 268 -2263 269 -2261
rect 268 -2269 269 -2267
rect 275 -2263 276 -2261
rect 275 -2269 276 -2267
rect 282 -2263 283 -2261
rect 282 -2269 283 -2267
rect 289 -2263 290 -2261
rect 289 -2269 290 -2267
rect 296 -2263 297 -2261
rect 296 -2269 297 -2267
rect 303 -2263 304 -2261
rect 306 -2263 307 -2261
rect 303 -2269 304 -2267
rect 306 -2269 307 -2267
rect 313 -2263 314 -2261
rect 313 -2269 314 -2267
rect 317 -2263 318 -2261
rect 317 -2269 318 -2267
rect 324 -2263 325 -2261
rect 327 -2263 328 -2261
rect 331 -2263 332 -2261
rect 331 -2269 332 -2267
rect 338 -2263 339 -2261
rect 338 -2269 339 -2267
rect 345 -2263 346 -2261
rect 345 -2269 346 -2267
rect 352 -2263 353 -2261
rect 352 -2269 353 -2267
rect 359 -2263 360 -2261
rect 362 -2263 363 -2261
rect 359 -2269 360 -2267
rect 362 -2269 363 -2267
rect 366 -2263 367 -2261
rect 366 -2269 367 -2267
rect 373 -2263 374 -2261
rect 373 -2269 374 -2267
rect 380 -2263 381 -2261
rect 380 -2269 381 -2267
rect 390 -2263 391 -2261
rect 387 -2269 388 -2267
rect 394 -2263 395 -2261
rect 397 -2263 398 -2261
rect 401 -2263 402 -2261
rect 401 -2269 402 -2267
rect 408 -2263 409 -2261
rect 408 -2269 409 -2267
rect 415 -2263 416 -2261
rect 415 -2269 416 -2267
rect 422 -2263 423 -2261
rect 422 -2269 423 -2267
rect 432 -2263 433 -2261
rect 429 -2269 430 -2267
rect 432 -2269 433 -2267
rect 436 -2263 437 -2261
rect 436 -2269 437 -2267
rect 443 -2263 444 -2261
rect 443 -2269 444 -2267
rect 450 -2263 451 -2261
rect 450 -2269 451 -2267
rect 457 -2263 458 -2261
rect 457 -2269 458 -2267
rect 464 -2263 465 -2261
rect 464 -2269 465 -2267
rect 471 -2269 472 -2267
rect 474 -2269 475 -2267
rect 478 -2263 479 -2261
rect 478 -2269 479 -2267
rect 485 -2263 486 -2261
rect 485 -2269 486 -2267
rect 492 -2263 493 -2261
rect 492 -2269 493 -2267
rect 499 -2263 500 -2261
rect 499 -2269 500 -2267
rect 506 -2263 507 -2261
rect 506 -2269 507 -2267
rect 513 -2263 514 -2261
rect 513 -2269 514 -2267
rect 520 -2263 521 -2261
rect 520 -2269 521 -2267
rect 527 -2263 528 -2261
rect 527 -2269 528 -2267
rect 534 -2263 535 -2261
rect 534 -2269 535 -2267
rect 541 -2263 542 -2261
rect 541 -2269 542 -2267
rect 548 -2263 549 -2261
rect 548 -2269 549 -2267
rect 555 -2263 556 -2261
rect 555 -2269 556 -2267
rect 562 -2263 563 -2261
rect 565 -2263 566 -2261
rect 569 -2269 570 -2267
rect 576 -2263 577 -2261
rect 576 -2269 577 -2267
rect 583 -2263 584 -2261
rect 583 -2269 584 -2267
rect 639 -2263 640 -2261
rect 639 -2269 640 -2267
rect 121 -2290 122 -2288
rect 177 -2290 178 -2288
rect 177 -2296 178 -2294
rect 212 -2290 213 -2288
rect 212 -2296 213 -2294
rect 222 -2290 223 -2288
rect 226 -2290 227 -2288
rect 226 -2296 227 -2294
rect 233 -2290 234 -2288
rect 233 -2296 234 -2294
rect 240 -2290 241 -2288
rect 243 -2296 244 -2294
rect 250 -2290 251 -2288
rect 254 -2290 255 -2288
rect 254 -2296 255 -2294
rect 268 -2290 269 -2288
rect 268 -2296 269 -2294
rect 275 -2290 276 -2288
rect 275 -2296 276 -2294
rect 282 -2290 283 -2288
rect 282 -2296 283 -2294
rect 289 -2290 290 -2288
rect 289 -2296 290 -2294
rect 296 -2290 297 -2288
rect 296 -2296 297 -2294
rect 303 -2290 304 -2288
rect 306 -2296 307 -2294
rect 310 -2290 311 -2288
rect 310 -2296 311 -2294
rect 317 -2290 318 -2288
rect 317 -2296 318 -2294
rect 327 -2296 328 -2294
rect 331 -2290 332 -2288
rect 331 -2296 332 -2294
rect 338 -2296 339 -2294
rect 345 -2290 346 -2288
rect 345 -2296 346 -2294
rect 366 -2290 367 -2288
rect 366 -2296 367 -2294
rect 380 -2290 381 -2288
rect 380 -2296 381 -2294
rect 404 -2290 405 -2288
rect 415 -2290 416 -2288
rect 415 -2296 416 -2294
rect 422 -2290 423 -2288
rect 422 -2296 423 -2294
rect 432 -2296 433 -2294
rect 439 -2290 440 -2288
rect 439 -2296 440 -2294
rect 443 -2296 444 -2294
rect 446 -2296 447 -2294
rect 450 -2290 451 -2288
rect 450 -2296 451 -2294
rect 457 -2290 458 -2288
rect 457 -2296 458 -2294
rect 464 -2290 465 -2288
rect 464 -2296 465 -2294
rect 474 -2290 475 -2288
rect 478 -2290 479 -2288
rect 502 -2290 503 -2288
rect 502 -2296 503 -2294
rect 506 -2290 507 -2288
rect 506 -2296 507 -2294
rect 513 -2290 514 -2288
rect 513 -2296 514 -2294
rect 520 -2290 521 -2288
rect 520 -2296 521 -2294
rect 527 -2290 528 -2288
rect 530 -2290 531 -2288
rect 534 -2290 535 -2288
rect 534 -2296 535 -2294
rect 541 -2290 542 -2288
rect 541 -2296 542 -2294
rect 548 -2290 549 -2288
rect 572 -2290 573 -2288
rect 569 -2296 570 -2294
rect 576 -2290 577 -2288
rect 576 -2296 577 -2294
rect 639 -2290 640 -2288
rect 639 -2296 640 -2294
rect 170 -2313 171 -2311
rect 177 -2307 178 -2305
rect 177 -2313 178 -2311
rect 215 -2307 216 -2305
rect 226 -2307 227 -2305
rect 226 -2313 227 -2311
rect 233 -2307 234 -2305
rect 233 -2313 234 -2311
rect 240 -2313 241 -2311
rect 247 -2307 248 -2305
rect 247 -2313 248 -2311
rect 254 -2307 255 -2305
rect 254 -2313 255 -2311
rect 264 -2307 265 -2305
rect 268 -2313 269 -2311
rect 275 -2313 276 -2311
rect 278 -2313 279 -2311
rect 285 -2307 286 -2305
rect 282 -2313 283 -2311
rect 289 -2307 290 -2305
rect 296 -2307 297 -2305
rect 296 -2313 297 -2311
rect 306 -2313 307 -2311
rect 313 -2307 314 -2305
rect 317 -2307 318 -2305
rect 317 -2313 318 -2311
rect 369 -2307 370 -2305
rect 380 -2307 381 -2305
rect 380 -2313 381 -2311
rect 387 -2313 388 -2311
rect 404 -2313 405 -2311
rect 408 -2307 409 -2305
rect 408 -2313 409 -2311
rect 509 -2307 510 -2305
rect 527 -2307 528 -2305
rect 527 -2313 528 -2311
rect 534 -2313 535 -2311
rect 597 -2307 598 -2305
rect 597 -2313 598 -2311
rect 604 -2307 605 -2305
rect 614 -2307 615 -2305
rect 611 -2313 612 -2311
rect 639 -2307 640 -2305
rect 642 -2313 643 -2311
rect 646 -2307 647 -2305
rect 646 -2313 647 -2311
<< metal1 >>
rect 177 0 192 1
rect 205 0 213 1
rect 257 0 283 1
rect 310 0 349 1
rect 359 0 367 1
rect 271 -2 276 -1
rect 177 -13 188 -12
rect 194 -13 199 -12
rect 212 -13 220 -12
rect 233 -13 255 -12
rect 261 -13 276 -12
rect 303 -13 311 -12
rect 341 -13 395 -12
rect 184 -15 209 -14
rect 215 -15 255 -14
rect 348 -15 388 -14
rect 198 -17 202 -16
rect 240 -17 251 -16
rect 366 -17 374 -16
rect 366 -19 384 -18
rect 166 -30 199 -29
rect 205 -30 272 -29
rect 289 -30 297 -29
rect 299 -30 353 -29
rect 387 -30 430 -29
rect 177 -32 213 -31
rect 215 -32 220 -31
rect 226 -32 241 -31
rect 247 -32 262 -31
rect 268 -32 342 -31
rect 345 -32 367 -31
rect 380 -32 388 -31
rect 394 -32 423 -31
rect 194 -34 276 -33
rect 296 -34 332 -33
rect 373 -34 395 -33
rect 411 -34 451 -33
rect 212 -36 234 -35
rect 254 -36 311 -35
rect 317 -36 335 -35
rect 366 -36 374 -35
rect 380 -36 416 -35
rect 219 -38 255 -37
rect 261 -38 339 -37
rect 233 -40 241 -39
rect 303 -40 325 -39
rect 86 -51 108 -50
rect 121 -51 129 -50
rect 142 -51 171 -50
rect 177 -51 188 -50
rect 191 -51 220 -50
rect 233 -51 311 -50
rect 317 -51 465 -50
rect 579 -51 584 -50
rect 93 -53 101 -52
rect 107 -53 171 -52
rect 177 -53 227 -52
rect 247 -53 297 -52
rect 303 -53 353 -52
rect 355 -53 409 -52
rect 436 -53 486 -52
rect 135 -55 220 -54
rect 247 -55 262 -54
rect 275 -55 374 -54
rect 394 -55 437 -54
rect 443 -55 472 -54
rect 149 -57 244 -56
rect 275 -57 363 -56
rect 376 -57 395 -56
rect 429 -57 444 -56
rect 450 -57 458 -56
rect 163 -59 216 -58
rect 240 -59 262 -58
rect 303 -59 346 -58
rect 348 -59 479 -58
rect 205 -61 318 -60
rect 331 -61 370 -60
rect 422 -61 451 -60
rect 198 -63 206 -62
rect 215 -63 227 -62
rect 324 -63 332 -62
rect 338 -63 381 -62
rect 387 -63 423 -62
rect 100 -65 199 -64
rect 289 -65 388 -64
rect 282 -67 290 -66
rect 310 -67 325 -66
rect 338 -67 416 -66
rect 282 -69 402 -68
rect 341 -71 430 -70
rect 362 -73 500 -72
rect 366 -75 416 -74
rect 401 -77 496 -76
rect 58 -88 136 -87
rect 149 -88 234 -87
rect 282 -88 311 -87
rect 313 -88 416 -87
rect 436 -88 556 -87
rect 565 -88 619 -87
rect 65 -90 143 -89
rect 177 -90 234 -89
rect 247 -90 416 -89
rect 436 -90 507 -89
rect 583 -90 598 -89
rect 72 -92 255 -91
rect 282 -92 290 -91
rect 345 -92 402 -91
rect 450 -92 570 -91
rect 79 -94 115 -93
rect 121 -94 192 -93
rect 205 -94 255 -93
rect 268 -94 402 -93
rect 457 -94 542 -93
rect 86 -96 125 -95
rect 180 -96 528 -95
rect 86 -98 164 -97
rect 184 -98 199 -97
rect 205 -98 227 -97
rect 247 -98 297 -97
rect 317 -98 346 -97
rect 348 -98 465 -97
rect 478 -98 493 -97
rect 93 -100 118 -99
rect 149 -100 185 -99
rect 187 -100 241 -99
rect 268 -100 300 -99
rect 352 -100 430 -99
rect 485 -100 584 -99
rect 93 -102 157 -101
rect 163 -102 171 -101
rect 226 -102 297 -101
rect 331 -102 430 -101
rect 114 -104 244 -103
rect 275 -104 318 -103
rect 331 -104 577 -103
rect 170 -106 286 -105
rect 289 -106 304 -105
rect 355 -106 472 -105
rect 156 -108 304 -107
rect 306 -108 472 -107
rect 243 -110 591 -109
rect 261 -112 276 -111
rect 359 -112 500 -111
rect 222 -114 262 -113
rect 362 -114 384 -113
rect 387 -114 535 -113
rect 107 -116 363 -115
rect 366 -116 451 -115
rect 142 -118 223 -117
rect 369 -118 521 -117
rect 177 -120 367 -119
rect 373 -120 500 -119
rect 100 -122 374 -121
rect 376 -122 514 -121
rect 100 -124 136 -123
rect 387 -124 507 -123
rect 394 -126 458 -125
rect 334 -128 395 -127
rect 408 -128 465 -127
rect 380 -130 409 -129
rect 422 -130 486 -129
rect 422 -132 479 -131
rect 51 -143 188 -142
rect 208 -143 377 -142
rect 380 -143 472 -142
rect 544 -143 573 -142
rect 618 -143 633 -142
rect 642 -143 647 -142
rect 65 -145 195 -144
rect 222 -145 255 -144
rect 282 -145 430 -144
rect 439 -145 577 -144
rect 65 -147 108 -146
rect 121 -147 230 -146
rect 236 -147 276 -146
rect 282 -147 318 -146
rect 320 -147 402 -146
rect 457 -147 472 -146
rect 506 -147 577 -146
rect 72 -149 377 -148
rect 387 -149 570 -148
rect 79 -151 178 -150
rect 180 -151 363 -150
rect 366 -151 542 -150
rect 79 -153 136 -152
rect 138 -153 367 -152
rect 390 -153 563 -152
rect 86 -155 188 -154
rect 247 -155 255 -154
rect 285 -155 416 -154
rect 457 -155 563 -154
rect 86 -157 244 -156
rect 296 -157 535 -156
rect 100 -159 164 -158
rect 173 -159 241 -158
rect 296 -159 521 -158
rect 527 -159 535 -158
rect 107 -161 157 -160
rect 191 -161 248 -160
rect 317 -161 325 -160
rect 331 -161 500 -160
rect 527 -161 591 -160
rect 114 -163 332 -162
rect 341 -163 388 -162
rect 408 -163 416 -162
rect 464 -163 549 -162
rect 114 -165 129 -164
rect 135 -165 213 -164
rect 324 -165 405 -164
rect 408 -165 423 -164
rect 443 -165 465 -164
rect 478 -165 521 -164
rect 121 -167 171 -166
rect 177 -167 213 -166
rect 345 -167 381 -166
rect 394 -167 479 -166
rect 492 -167 500 -166
rect 513 -167 591 -166
rect 128 -169 311 -168
rect 338 -169 346 -168
rect 352 -169 430 -168
rect 436 -169 514 -168
rect 149 -171 307 -170
rect 359 -171 584 -170
rect 149 -173 300 -172
rect 362 -173 444 -172
rect 450 -173 493 -172
rect 583 -173 598 -172
rect 156 -175 206 -174
rect 261 -175 311 -174
rect 355 -175 451 -174
rect 163 -177 353 -176
rect 355 -177 556 -176
rect 170 -179 269 -178
rect 275 -179 360 -178
rect 551 -179 556 -178
rect 205 -181 423 -180
rect 226 -183 269 -182
rect 289 -183 339 -182
rect 198 -185 227 -184
rect 233 -185 262 -184
rect 289 -185 374 -184
rect 93 -187 234 -186
rect 93 -189 143 -188
rect 198 -189 216 -188
rect 58 -191 143 -190
rect 215 -191 220 -190
rect 16 -202 157 -201
rect 187 -202 276 -201
rect 303 -202 640 -201
rect 646 -202 689 -201
rect 37 -204 185 -203
rect 198 -204 297 -203
rect 320 -204 451 -203
rect 460 -204 661 -203
rect 670 -204 675 -203
rect 44 -206 132 -205
rect 205 -206 514 -205
rect 520 -206 654 -205
rect 65 -208 195 -207
rect 212 -208 220 -207
rect 233 -208 402 -207
rect 411 -208 440 -207
rect 467 -208 612 -207
rect 618 -208 633 -207
rect 65 -210 143 -209
rect 233 -210 241 -209
rect 261 -210 276 -209
rect 289 -210 304 -209
rect 331 -210 458 -209
rect 513 -210 549 -209
rect 562 -210 696 -209
rect 79 -212 220 -211
rect 236 -212 297 -211
rect 355 -212 563 -211
rect 569 -212 584 -211
rect 590 -212 633 -211
rect 51 -214 80 -213
rect 86 -214 139 -213
rect 173 -214 290 -213
rect 359 -214 381 -213
rect 390 -214 479 -213
rect 520 -214 556 -213
rect 569 -214 752 -213
rect 86 -216 150 -215
rect 222 -216 381 -215
rect 397 -216 465 -215
rect 471 -216 556 -215
rect 576 -216 682 -215
rect 93 -218 262 -217
rect 268 -218 332 -217
rect 373 -218 626 -217
rect 93 -220 146 -219
rect 198 -220 269 -219
rect 282 -220 374 -219
rect 376 -220 486 -219
rect 492 -220 577 -219
rect 597 -220 668 -219
rect 100 -222 185 -221
rect 240 -222 255 -221
rect 299 -222 472 -221
rect 527 -222 647 -221
rect 30 -224 101 -223
rect 107 -224 192 -223
rect 226 -224 255 -223
rect 397 -224 451 -223
rect 464 -224 535 -223
rect 544 -224 584 -223
rect 23 -226 108 -225
rect 121 -226 150 -225
rect 177 -226 283 -225
rect 324 -226 535 -225
rect 58 -228 227 -227
rect 310 -228 325 -227
rect 404 -228 479 -227
rect 509 -228 528 -227
rect 72 -230 192 -229
rect 247 -230 311 -229
rect 408 -230 549 -229
rect 72 -232 115 -231
rect 121 -232 143 -231
rect 163 -232 248 -231
rect 408 -232 500 -231
rect 114 -234 209 -233
rect 415 -234 437 -233
rect 443 -234 493 -233
rect 128 -236 353 -235
rect 366 -236 444 -235
rect 485 -236 510 -235
rect 128 -238 171 -237
rect 208 -238 542 -237
rect 138 -240 178 -239
rect 338 -240 367 -239
rect 422 -240 591 -239
rect 163 -242 230 -241
rect 338 -242 500 -241
rect 345 -244 416 -243
rect 418 -244 423 -243
rect 429 -244 507 -243
rect 345 -246 388 -245
rect 394 -246 430 -245
rect 394 -248 605 -247
rect 23 -259 136 -258
rect 142 -259 262 -258
rect 299 -259 426 -258
rect 439 -259 577 -258
rect 590 -259 594 -258
rect 597 -259 601 -258
rect 604 -259 671 -258
rect 674 -259 717 -258
rect 751 -259 829 -258
rect 856 -259 860 -258
rect 51 -261 59 -260
rect 65 -261 237 -260
rect 240 -261 272 -260
rect 334 -261 661 -260
rect 681 -261 738 -260
rect 16 -263 241 -262
rect 247 -263 398 -262
rect 401 -263 573 -262
rect 590 -263 640 -262
rect 646 -263 682 -262
rect 688 -263 745 -262
rect 58 -265 80 -264
rect 107 -265 122 -264
rect 128 -265 227 -264
rect 229 -265 255 -264
rect 261 -265 276 -264
rect 338 -265 353 -264
rect 359 -265 409 -264
rect 415 -265 423 -264
rect 443 -265 479 -264
rect 499 -265 503 -264
rect 534 -265 570 -264
rect 597 -265 612 -264
rect 618 -265 668 -264
rect 688 -265 724 -264
rect 44 -267 80 -266
rect 107 -267 157 -266
rect 191 -267 195 -266
rect 205 -267 227 -266
rect 268 -267 353 -266
rect 359 -267 402 -266
rect 446 -267 605 -266
rect 625 -267 710 -266
rect 68 -269 101 -268
rect 114 -269 160 -268
rect 184 -269 269 -268
rect 275 -269 311 -268
rect 341 -269 458 -268
rect 460 -269 731 -268
rect 72 -271 139 -270
rect 149 -271 157 -270
rect 177 -271 185 -270
rect 205 -271 297 -270
rect 310 -271 318 -270
rect 373 -271 398 -270
rect 481 -271 668 -270
rect 37 -273 178 -272
rect 215 -273 405 -272
rect 499 -273 514 -272
rect 520 -273 626 -272
rect 632 -273 647 -272
rect 30 -275 216 -274
rect 222 -275 283 -274
rect 296 -275 304 -274
rect 317 -275 325 -274
rect 373 -275 752 -274
rect 30 -277 87 -276
rect 100 -277 104 -276
rect 117 -277 633 -276
rect 639 -277 654 -276
rect 37 -279 94 -278
rect 121 -279 199 -278
rect 282 -279 332 -278
rect 380 -279 465 -278
rect 471 -279 521 -278
rect 541 -279 619 -278
rect 72 -281 164 -280
rect 180 -281 199 -280
rect 243 -281 381 -280
rect 390 -281 545 -280
rect 555 -281 661 -280
rect 86 -283 332 -282
rect 394 -283 535 -282
rect 562 -283 577 -282
rect 600 -283 612 -282
rect 93 -285 255 -284
rect 289 -285 304 -284
rect 324 -285 367 -284
rect 429 -285 472 -284
rect 527 -285 556 -284
rect 565 -285 703 -284
rect 149 -287 171 -286
rect 345 -287 367 -286
rect 411 -287 528 -286
rect 163 -289 542 -288
rect 170 -291 234 -290
rect 345 -291 549 -290
rect 387 -293 549 -292
rect 387 -295 696 -294
rect 429 -297 437 -296
rect 450 -297 563 -296
rect 422 -299 451 -298
rect 506 -299 696 -298
rect 338 -301 507 -300
rect 2 -312 101 -311
rect 107 -312 115 -311
rect 121 -312 125 -311
rect 128 -312 496 -311
rect 653 -312 836 -311
rect 849 -312 864 -311
rect 9 -314 66 -313
rect 72 -314 216 -313
rect 233 -314 346 -313
rect 352 -314 563 -313
rect 590 -314 654 -313
rect 674 -314 678 -313
rect 681 -314 724 -313
rect 726 -314 871 -313
rect 16 -316 80 -315
rect 114 -316 416 -315
rect 422 -316 493 -315
rect 534 -316 563 -315
rect 569 -316 591 -315
rect 695 -316 780 -315
rect 828 -316 892 -315
rect 23 -318 178 -317
rect 215 -318 248 -317
rect 257 -318 262 -317
rect 275 -318 342 -317
rect 352 -318 486 -317
rect 513 -318 535 -317
rect 548 -318 570 -317
rect 597 -318 696 -317
rect 702 -318 815 -317
rect 852 -318 857 -317
rect 30 -320 80 -319
rect 96 -320 178 -319
rect 219 -320 346 -319
rect 359 -320 433 -319
rect 450 -320 454 -319
rect 513 -320 521 -319
rect 544 -320 703 -319
rect 709 -320 759 -319
rect 44 -322 108 -321
rect 121 -322 395 -321
rect 401 -322 661 -321
rect 667 -322 710 -321
rect 730 -322 829 -321
rect 44 -324 237 -323
rect 240 -324 444 -323
rect 450 -324 472 -323
rect 520 -324 528 -323
rect 583 -324 598 -323
rect 618 -324 661 -323
rect 737 -324 808 -323
rect 51 -326 339 -325
rect 362 -326 801 -325
rect 51 -328 185 -327
rect 233 -328 794 -327
rect 37 -330 185 -329
rect 240 -330 283 -329
rect 289 -330 682 -329
rect 744 -330 787 -329
rect 58 -332 132 -331
rect 135 -332 223 -331
rect 247 -332 318 -331
rect 334 -332 409 -331
rect 471 -332 479 -331
rect 499 -332 528 -331
rect 583 -332 633 -331
rect 639 -332 731 -331
rect 751 -332 822 -331
rect 58 -334 150 -333
rect 212 -334 409 -333
rect 474 -334 619 -333
rect 639 -334 878 -333
rect 65 -336 192 -335
rect 261 -336 304 -335
rect 310 -336 339 -335
rect 373 -336 766 -335
rect 75 -338 153 -337
rect 170 -338 192 -337
rect 282 -338 325 -337
rect 380 -338 549 -337
rect 586 -338 857 -337
rect 86 -340 318 -339
rect 380 -340 388 -339
rect 394 -340 458 -339
rect 506 -340 633 -339
rect 646 -340 668 -339
rect 688 -340 752 -339
rect 86 -342 269 -341
rect 289 -342 325 -341
rect 401 -342 426 -341
rect 436 -342 689 -341
rect 93 -344 311 -343
rect 429 -344 437 -343
rect 457 -344 465 -343
rect 516 -344 745 -343
rect 93 -346 843 -345
rect 100 -348 360 -347
rect 429 -348 500 -347
rect 604 -348 738 -347
rect 128 -350 220 -349
rect 254 -350 388 -349
rect 604 -350 612 -349
rect 625 -350 647 -349
rect 138 -352 276 -351
rect 296 -352 405 -351
rect 576 -352 612 -351
rect 142 -354 370 -353
rect 555 -354 577 -353
rect 30 -356 143 -355
rect 145 -356 486 -355
rect 156 -358 171 -357
rect 198 -358 465 -357
rect 156 -360 164 -359
rect 254 -360 328 -359
rect 331 -360 556 -359
rect 37 -362 332 -361
rect 334 -362 626 -361
rect 163 -364 206 -363
rect 268 -364 440 -363
rect 453 -364 479 -363
rect 205 -366 416 -365
rect 299 -368 542 -367
rect 303 -370 367 -369
rect 366 -372 773 -371
rect 2 -383 199 -382
rect 205 -383 941 -382
rect 2 -385 199 -384
rect 261 -385 363 -384
rect 369 -385 535 -384
rect 621 -385 640 -384
rect 828 -385 878 -384
rect 16 -387 132 -386
rect 159 -387 906 -386
rect 16 -389 45 -388
rect 51 -389 216 -388
rect 261 -389 433 -388
rect 478 -389 514 -388
rect 516 -389 738 -388
rect 842 -389 899 -388
rect 23 -391 244 -390
rect 275 -391 433 -390
rect 436 -391 479 -390
rect 502 -391 808 -390
rect 852 -391 892 -390
rect 23 -393 178 -392
rect 282 -393 377 -392
rect 390 -393 780 -392
rect 807 -393 850 -392
rect 863 -393 885 -392
rect 37 -395 507 -394
rect 509 -395 934 -394
rect 37 -397 104 -396
rect 107 -397 223 -396
rect 310 -397 349 -396
rect 359 -397 654 -396
rect 716 -397 892 -396
rect 44 -399 178 -398
rect 184 -399 283 -398
rect 303 -399 311 -398
rect 317 -399 493 -398
rect 495 -399 885 -398
rect 54 -401 136 -400
rect 145 -401 864 -400
rect 870 -401 927 -400
rect 75 -403 269 -402
rect 303 -403 822 -402
rect 79 -405 97 -404
rect 100 -405 185 -404
rect 201 -405 269 -404
rect 324 -405 395 -404
rect 401 -405 458 -404
rect 520 -405 584 -404
rect 604 -405 640 -404
rect 674 -405 871 -404
rect 9 -407 80 -406
rect 86 -407 234 -406
rect 240 -407 360 -406
rect 373 -407 829 -406
rect 9 -409 220 -408
rect 240 -409 318 -408
rect 331 -409 353 -408
rect 408 -409 510 -408
rect 520 -409 752 -408
rect 772 -409 850 -408
rect 72 -411 353 -410
rect 369 -411 409 -410
rect 415 -411 535 -410
rect 555 -411 654 -410
rect 695 -411 773 -410
rect 814 -411 822 -410
rect 72 -413 164 -412
rect 170 -413 206 -412
rect 212 -413 780 -412
rect 86 -415 157 -414
rect 163 -415 570 -414
rect 576 -415 605 -414
rect 625 -415 696 -414
rect 716 -415 801 -414
rect 93 -417 248 -416
rect 254 -417 374 -416
rect 422 -417 843 -416
rect 65 -419 255 -418
rect 289 -419 395 -418
rect 422 -419 682 -418
rect 730 -419 815 -418
rect 58 -421 66 -420
rect 107 -421 367 -420
rect 425 -421 598 -420
rect 611 -421 626 -420
rect 646 -421 682 -420
rect 730 -421 766 -420
rect 58 -423 297 -422
rect 338 -423 948 -422
rect 110 -425 248 -424
rect 289 -425 381 -424
rect 436 -425 836 -424
rect 117 -427 384 -426
rect 450 -427 458 -426
rect 471 -427 801 -426
rect 835 -427 857 -426
rect 114 -429 472 -428
rect 485 -429 577 -428
rect 590 -429 675 -428
rect 688 -429 766 -428
rect 114 -431 570 -430
rect 632 -431 857 -430
rect 121 -433 402 -432
rect 418 -433 451 -432
rect 523 -433 920 -432
rect 121 -435 150 -434
rect 156 -435 335 -434
rect 345 -435 514 -434
rect 527 -435 591 -434
rect 646 -435 668 -434
rect 688 -435 710 -434
rect 751 -435 787 -434
rect 30 -437 150 -436
rect 212 -437 913 -436
rect 30 -439 129 -438
rect 135 -439 307 -438
rect 366 -439 598 -438
rect 618 -439 787 -438
rect 128 -441 192 -440
rect 233 -441 486 -440
rect 548 -441 633 -440
rect 667 -441 745 -440
rect 142 -443 171 -442
rect 191 -443 339 -442
rect 404 -443 528 -442
rect 555 -443 563 -442
rect 611 -443 619 -442
rect 702 -443 710 -442
rect 142 -445 430 -444
rect 443 -445 549 -444
rect 702 -445 794 -444
rect 152 -447 745 -446
rect 296 -449 738 -448
rect 331 -451 430 -450
rect 541 -451 563 -450
rect 723 -451 794 -450
rect 299 -453 724 -452
rect 387 -455 444 -454
rect 499 -455 542 -454
rect 278 -457 500 -456
rect 387 -459 465 -458
rect 415 -461 465 -460
rect 2 -472 265 -471
rect 268 -472 426 -471
rect 429 -472 815 -471
rect 2 -474 220 -473
rect 243 -474 514 -473
rect 544 -474 892 -473
rect 9 -476 521 -475
rect 607 -476 619 -475
rect 726 -476 822 -475
rect 9 -478 45 -477
rect 51 -478 146 -477
rect 180 -478 202 -477
rect 212 -478 941 -477
rect 30 -480 52 -479
rect 54 -480 696 -479
rect 814 -480 920 -479
rect 30 -482 38 -481
rect 58 -482 304 -481
rect 313 -482 948 -481
rect 37 -484 384 -483
rect 394 -484 419 -483
rect 439 -484 797 -483
rect 58 -486 136 -485
rect 184 -486 220 -485
rect 243 -486 283 -485
rect 303 -486 318 -485
rect 320 -486 549 -485
rect 695 -486 703 -485
rect 79 -488 97 -487
rect 100 -488 654 -487
rect 660 -488 703 -487
rect 23 -490 80 -489
rect 86 -490 199 -489
rect 324 -490 395 -489
rect 401 -490 822 -489
rect 86 -492 248 -491
rect 352 -492 433 -491
rect 460 -492 766 -491
rect 100 -494 108 -493
rect 114 -494 391 -493
rect 408 -494 430 -493
rect 464 -494 524 -493
rect 541 -494 549 -493
rect 639 -494 661 -493
rect 765 -494 836 -493
rect 82 -496 108 -495
rect 117 -496 675 -495
rect 835 -496 843 -495
rect 121 -498 409 -497
rect 415 -498 794 -497
rect 121 -500 346 -499
rect 359 -500 370 -499
rect 373 -500 402 -499
rect 415 -500 577 -499
rect 639 -500 668 -499
rect 674 -500 689 -499
rect 128 -502 297 -501
rect 324 -502 542 -501
rect 576 -502 605 -501
rect 646 -502 654 -501
rect 667 -502 755 -501
rect 16 -504 129 -503
rect 135 -504 311 -503
rect 366 -504 472 -503
rect 485 -504 780 -503
rect 16 -506 164 -505
rect 166 -506 486 -505
rect 488 -506 871 -505
rect 142 -508 353 -507
rect 373 -508 535 -507
rect 646 -508 850 -507
rect 149 -510 167 -509
rect 177 -510 283 -509
rect 296 -510 335 -509
rect 338 -510 367 -509
rect 380 -510 633 -509
rect 688 -510 738 -509
rect 779 -510 885 -509
rect 65 -512 150 -511
rect 156 -512 472 -511
rect 502 -512 899 -511
rect 65 -514 349 -513
rect 464 -514 482 -513
rect 506 -514 787 -513
rect 163 -516 423 -515
rect 509 -516 857 -515
rect 184 -518 227 -517
rect 247 -518 388 -517
rect 422 -518 584 -517
rect 632 -518 682 -517
rect 709 -518 738 -517
rect 786 -518 934 -517
rect 191 -520 773 -519
rect 856 -520 927 -519
rect 93 -522 192 -521
rect 194 -522 241 -521
rect 254 -522 346 -521
rect 387 -522 591 -521
rect 709 -522 801 -521
rect 93 -524 307 -523
rect 341 -524 535 -523
rect 569 -524 584 -523
rect 590 -524 598 -523
rect 751 -524 773 -523
rect 800 -524 913 -523
rect 198 -526 234 -525
rect 240 -526 906 -525
rect 226 -528 493 -527
rect 513 -528 528 -527
rect 597 -528 626 -527
rect 233 -530 500 -529
rect 520 -530 745 -529
rect 254 -532 276 -531
rect 289 -532 381 -531
rect 436 -532 570 -531
rect 611 -532 626 -531
rect 744 -532 759 -531
rect 205 -534 276 -533
rect 289 -534 332 -533
rect 453 -534 612 -533
rect 730 -534 759 -533
rect 72 -536 206 -535
rect 268 -536 311 -535
rect 457 -536 682 -535
rect 730 -536 829 -535
rect 72 -538 451 -537
rect 457 -538 479 -537
rect 499 -538 864 -537
rect 450 -540 496 -539
rect 527 -540 563 -539
rect 478 -542 724 -541
rect 555 -544 563 -543
rect 723 -544 878 -543
rect 261 -546 556 -545
rect 261 -548 437 -547
rect 2 -559 482 -558
rect 502 -559 577 -558
rect 583 -559 605 -558
rect 607 -559 626 -558
rect 681 -559 899 -558
rect 2 -561 31 -560
rect 37 -561 97 -560
rect 131 -561 164 -560
rect 177 -561 318 -560
rect 345 -561 363 -560
rect 373 -561 496 -560
rect 506 -561 538 -560
rect 541 -561 829 -560
rect 835 -561 843 -560
rect 9 -563 125 -562
rect 135 -563 332 -562
rect 373 -563 402 -562
rect 404 -563 885 -562
rect 9 -565 87 -564
rect 156 -565 244 -564
rect 317 -565 524 -564
rect 544 -565 906 -564
rect 23 -567 181 -566
rect 191 -567 342 -566
rect 401 -567 479 -566
rect 520 -567 626 -566
rect 646 -567 836 -566
rect 23 -569 52 -568
rect 58 -569 262 -568
rect 415 -569 451 -568
rect 453 -569 528 -568
rect 555 -569 727 -568
rect 744 -569 752 -568
rect 754 -569 927 -568
rect 30 -571 307 -570
rect 436 -571 510 -570
rect 562 -571 577 -570
rect 583 -571 598 -570
rect 660 -571 682 -570
rect 695 -571 752 -570
rect 765 -571 850 -570
rect 40 -573 342 -572
rect 429 -573 437 -572
rect 457 -573 556 -572
rect 597 -573 689 -572
rect 723 -573 948 -572
rect 44 -575 87 -574
rect 103 -575 262 -574
rect 348 -575 430 -574
rect 457 -575 514 -574
rect 548 -575 563 -574
rect 618 -575 724 -574
rect 744 -575 759 -574
rect 772 -575 892 -574
rect 51 -577 122 -576
rect 128 -577 549 -576
rect 653 -577 661 -576
rect 698 -577 773 -576
rect 786 -577 913 -576
rect 65 -579 69 -578
rect 79 -579 391 -578
rect 474 -579 633 -578
rect 702 -579 759 -578
rect 793 -579 857 -578
rect 65 -581 314 -580
rect 338 -581 787 -580
rect 800 -581 871 -580
rect 79 -583 185 -582
rect 191 -583 332 -582
rect 485 -583 766 -582
rect 779 -583 857 -582
rect 93 -585 794 -584
rect 800 -585 808 -584
rect 814 -585 864 -584
rect 93 -587 101 -586
rect 135 -587 689 -586
rect 730 -587 808 -586
rect 159 -589 241 -588
rect 264 -589 731 -588
rect 737 -589 815 -588
rect 166 -591 647 -590
rect 173 -593 178 -592
rect 184 -593 199 -592
rect 205 -593 878 -592
rect 198 -595 297 -594
rect 313 -595 444 -594
rect 471 -595 780 -594
rect 205 -597 220 -596
rect 226 -597 528 -596
rect 534 -597 654 -596
rect 212 -599 283 -598
rect 289 -599 444 -598
rect 471 -599 591 -598
rect 632 -599 668 -598
rect 16 -601 213 -600
rect 215 -601 346 -600
rect 359 -601 486 -600
rect 513 -601 545 -600
rect 569 -601 738 -600
rect 16 -603 62 -602
rect 219 -603 234 -602
rect 236 -603 423 -602
rect 425 -603 668 -602
rect 114 -605 423 -604
rect 590 -605 675 -604
rect 114 -607 171 -606
rect 226 -607 269 -606
rect 275 -607 297 -606
rect 359 -607 367 -606
rect 380 -607 570 -606
rect 639 -607 703 -606
rect 149 -609 234 -608
rect 247 -609 269 -608
rect 275 -609 500 -608
rect 611 -609 640 -608
rect 149 -611 325 -610
rect 338 -611 381 -610
rect 467 -611 500 -610
rect 611 -611 717 -610
rect 145 -613 325 -612
rect 366 -613 395 -612
rect 492 -613 675 -612
rect 709 -613 717 -612
rect 247 -615 388 -614
rect 450 -615 710 -614
rect 72 -617 388 -616
rect 72 -619 311 -618
rect 334 -619 493 -618
rect 282 -621 304 -620
rect 352 -621 395 -620
rect 289 -623 409 -622
rect 68 -625 409 -624
rect 352 -627 465 -626
rect 464 -629 822 -628
rect 593 -631 822 -630
rect 2 -642 59 -641
rect 61 -642 136 -641
rect 138 -642 454 -641
rect 464 -642 724 -641
rect 821 -642 955 -641
rect 2 -644 157 -643
rect 173 -644 283 -643
rect 289 -644 304 -643
rect 331 -644 570 -643
rect 590 -644 871 -643
rect 947 -644 1032 -643
rect 16 -646 87 -645
rect 93 -646 111 -645
rect 184 -646 412 -645
rect 436 -646 465 -645
rect 488 -646 584 -645
rect 593 -646 906 -645
rect 16 -648 150 -647
rect 184 -648 269 -647
rect 289 -648 395 -647
rect 404 -648 556 -647
rect 562 -648 570 -647
rect 583 -648 633 -647
rect 660 -648 696 -647
rect 793 -648 822 -647
rect 891 -648 906 -647
rect 37 -650 335 -649
rect 338 -650 367 -649
rect 387 -650 451 -649
rect 481 -650 594 -649
rect 604 -650 619 -649
rect 621 -650 759 -649
rect 786 -650 794 -649
rect 814 -650 871 -649
rect 51 -652 472 -651
rect 502 -652 808 -651
rect 828 -652 892 -651
rect 30 -654 472 -653
rect 513 -654 535 -653
rect 537 -654 766 -653
rect 779 -654 787 -653
rect 51 -656 479 -655
rect 520 -656 913 -655
rect 58 -658 178 -657
rect 198 -658 269 -657
rect 338 -658 475 -657
rect 506 -658 521 -657
rect 523 -658 598 -657
rect 611 -658 815 -657
rect 912 -658 927 -657
rect 65 -660 157 -659
rect 177 -660 276 -659
rect 341 -660 374 -659
rect 436 -660 545 -659
rect 551 -660 703 -659
rect 716 -660 780 -659
rect 65 -662 122 -661
rect 149 -662 192 -661
rect 198 -662 220 -661
rect 233 -662 318 -661
rect 345 -662 528 -661
rect 541 -662 710 -661
rect 730 -662 927 -661
rect 72 -664 318 -663
rect 359 -664 395 -663
rect 408 -664 528 -663
rect 541 -664 857 -663
rect 72 -666 444 -665
rect 474 -666 829 -665
rect 79 -668 244 -667
rect 247 -668 283 -667
rect 366 -668 402 -667
rect 443 -668 468 -667
rect 499 -668 507 -667
rect 555 -668 738 -667
rect 765 -668 836 -667
rect 9 -670 244 -669
rect 250 -670 255 -669
rect 275 -670 416 -669
rect 478 -670 738 -669
rect 9 -672 45 -671
rect 79 -672 381 -671
rect 390 -672 836 -671
rect 23 -674 45 -673
rect 86 -674 857 -673
rect 93 -676 146 -675
rect 170 -676 192 -675
rect 205 -676 304 -675
rect 324 -676 402 -675
rect 562 -676 850 -675
rect 100 -678 549 -677
rect 576 -678 605 -677
rect 614 -678 920 -677
rect 103 -680 612 -679
rect 625 -680 633 -679
rect 639 -680 661 -679
rect 667 -680 920 -679
rect 100 -682 668 -681
rect 674 -682 724 -681
rect 730 -682 801 -681
rect 842 -682 850 -681
rect 103 -684 143 -683
rect 170 -684 262 -683
rect 324 -684 430 -683
rect 576 -684 626 -683
rect 639 -684 888 -683
rect 107 -686 129 -685
rect 205 -686 255 -685
rect 261 -686 311 -685
rect 352 -686 416 -685
rect 422 -686 430 -685
rect 646 -686 675 -685
rect 688 -686 759 -685
rect 772 -686 801 -685
rect 842 -686 878 -685
rect 114 -688 311 -687
rect 352 -688 629 -687
rect 653 -688 703 -687
rect 751 -688 773 -687
rect 877 -688 899 -687
rect 89 -690 115 -689
rect 121 -690 164 -689
rect 212 -690 598 -689
rect 744 -690 752 -689
rect 863 -690 899 -689
rect 135 -692 213 -691
rect 219 -692 297 -691
rect 380 -692 458 -691
rect 485 -692 647 -691
rect 681 -692 745 -691
rect 863 -692 885 -691
rect 145 -694 689 -693
rect 163 -696 566 -695
rect 226 -698 409 -697
rect 422 -698 549 -697
rect 558 -698 682 -697
rect 229 -700 458 -699
rect 485 -700 717 -699
rect 236 -702 710 -701
rect 240 -704 360 -703
rect 492 -704 654 -703
rect 240 -706 808 -705
rect 296 -708 419 -707
rect 348 -710 493 -709
rect 16 -721 104 -720
rect 135 -721 391 -720
rect 415 -721 766 -720
rect 849 -721 885 -720
rect 908 -721 913 -720
rect 926 -721 976 -720
rect 1006 -721 1018 -720
rect 1031 -721 1067 -720
rect 23 -723 118 -722
rect 135 -723 150 -722
rect 170 -723 419 -722
rect 478 -723 545 -722
rect 551 -723 857 -722
rect 912 -723 962 -722
rect 26 -725 31 -724
rect 33 -725 671 -724
rect 716 -725 766 -724
rect 793 -725 850 -724
rect 954 -725 1011 -724
rect 30 -727 164 -726
rect 170 -727 188 -726
rect 229 -727 311 -726
rect 317 -727 388 -726
rect 464 -727 479 -726
rect 481 -727 584 -726
rect 590 -727 717 -726
rect 744 -727 794 -726
rect 807 -727 857 -726
rect 44 -729 111 -728
rect 128 -729 388 -728
rect 436 -729 465 -728
rect 488 -729 535 -728
rect 555 -729 836 -728
rect 2 -731 45 -730
rect 58 -731 206 -730
rect 240 -731 542 -730
rect 558 -731 892 -730
rect 58 -733 192 -732
rect 205 -733 234 -732
rect 247 -733 339 -732
rect 348 -733 493 -732
rect 516 -733 654 -732
rect 674 -733 745 -732
rect 779 -733 808 -732
rect 891 -733 916 -732
rect 86 -735 598 -734
rect 621 -735 906 -734
rect 86 -737 283 -736
rect 317 -737 500 -736
rect 506 -737 598 -736
rect 625 -737 899 -736
rect 51 -739 507 -738
rect 527 -739 549 -738
rect 565 -739 801 -738
rect 898 -739 920 -738
rect 65 -741 500 -740
rect 541 -741 675 -740
rect 723 -741 780 -740
rect 814 -741 920 -740
rect 89 -743 668 -742
rect 688 -743 724 -742
rect 737 -743 836 -742
rect 93 -745 244 -744
rect 254 -745 356 -744
rect 373 -745 822 -744
rect 51 -747 94 -746
rect 128 -747 496 -746
rect 569 -747 591 -746
rect 625 -747 640 -746
rect 667 -747 731 -746
rect 758 -747 801 -746
rect 821 -747 829 -746
rect 72 -749 374 -748
rect 394 -749 535 -748
rect 569 -749 577 -748
rect 579 -749 773 -748
rect 142 -751 220 -750
rect 261 -751 265 -750
rect 268 -751 283 -750
rect 331 -751 430 -750
rect 436 -751 458 -750
rect 485 -751 654 -750
rect 660 -751 731 -750
rect 9 -753 458 -752
rect 527 -753 829 -752
rect 107 -755 269 -754
rect 296 -755 430 -754
rect 576 -755 773 -754
rect 107 -757 115 -756
rect 142 -757 353 -756
rect 380 -757 486 -756
rect 583 -757 605 -756
rect 628 -757 871 -756
rect 100 -759 115 -758
rect 145 -759 150 -758
rect 156 -759 164 -758
rect 191 -759 251 -758
rect 254 -759 262 -758
rect 296 -759 346 -758
rect 359 -759 381 -758
rect 394 -759 402 -758
rect 415 -759 815 -758
rect 842 -759 871 -758
rect 100 -761 409 -760
rect 639 -761 647 -760
rect 688 -761 752 -760
rect 786 -761 843 -760
rect 156 -763 199 -762
rect 212 -763 220 -762
rect 236 -763 661 -762
rect 702 -763 738 -762
rect 751 -763 878 -762
rect 37 -765 213 -764
rect 243 -765 360 -764
rect 408 -765 444 -764
rect 450 -765 647 -764
rect 681 -765 703 -764
rect 709 -765 759 -764
rect 863 -765 878 -764
rect 37 -767 514 -766
rect 520 -767 682 -766
rect 695 -767 710 -766
rect 177 -769 199 -768
rect 275 -769 402 -768
rect 404 -769 444 -768
rect 450 -769 531 -768
rect 611 -769 696 -768
rect 79 -771 276 -770
rect 289 -771 521 -770
rect 562 -771 612 -770
rect 632 -771 787 -770
rect 79 -773 377 -772
rect 492 -773 864 -772
rect 177 -775 185 -774
rect 289 -775 304 -774
rect 324 -775 353 -774
rect 513 -775 605 -774
rect 618 -775 633 -774
rect 121 -777 185 -776
rect 310 -777 325 -776
rect 338 -777 367 -776
rect 471 -777 619 -776
rect 110 -779 122 -778
rect 131 -779 304 -778
rect 345 -779 503 -778
rect 366 -781 423 -780
rect 16 -792 66 -791
rect 68 -792 111 -791
rect 114 -792 244 -791
rect 310 -792 370 -791
rect 387 -792 948 -791
rect 961 -792 1014 -791
rect 1017 -792 1025 -791
rect 1066 -792 1081 -791
rect 23 -794 73 -793
rect 79 -794 181 -793
rect 233 -794 304 -793
rect 338 -794 451 -793
rect 492 -794 745 -793
rect 814 -794 955 -793
rect 975 -794 1018 -793
rect 23 -796 150 -795
rect 173 -796 363 -795
rect 411 -796 521 -795
rect 523 -796 850 -795
rect 863 -796 934 -795
rect 989 -796 993 -795
rect 1010 -796 1039 -795
rect 30 -798 314 -797
rect 380 -798 521 -797
rect 530 -798 640 -797
rect 653 -798 850 -797
rect 877 -798 997 -797
rect 37 -800 185 -799
rect 233 -800 297 -799
rect 380 -800 542 -799
rect 551 -800 654 -799
rect 695 -800 895 -799
rect 915 -800 1004 -799
rect 37 -802 227 -801
rect 240 -802 290 -801
rect 296 -802 577 -801
rect 618 -802 787 -801
rect 817 -802 962 -801
rect 44 -804 237 -803
rect 254 -804 577 -803
rect 621 -804 899 -803
rect 47 -806 262 -805
rect 268 -806 304 -805
rect 422 -806 969 -805
rect 51 -808 230 -807
rect 254 -808 318 -807
rect 422 -808 430 -807
rect 439 -808 913 -807
rect 30 -810 230 -809
rect 261 -810 528 -809
rect 537 -810 752 -809
rect 800 -810 899 -809
rect 58 -812 353 -811
rect 429 -812 738 -811
rect 751 -812 906 -811
rect 12 -814 59 -813
rect 72 -814 143 -813
rect 149 -814 220 -813
rect 282 -814 353 -813
rect 450 -814 479 -813
rect 485 -814 528 -813
rect 544 -814 619 -813
rect 639 -814 990 -813
rect 79 -816 468 -815
rect 471 -816 486 -815
rect 492 -816 745 -815
rect 821 -816 983 -815
rect 86 -818 426 -817
rect 443 -818 472 -817
rect 478 -818 668 -817
rect 681 -818 738 -817
rect 765 -818 822 -817
rect 828 -818 976 -817
rect 86 -820 94 -819
rect 114 -820 409 -819
rect 499 -820 682 -819
rect 695 -820 815 -819
rect 828 -820 885 -819
rect 93 -822 164 -821
rect 184 -822 346 -821
rect 513 -822 591 -821
rect 667 -822 689 -821
rect 716 -822 864 -821
rect 121 -824 402 -823
rect 513 -824 626 -823
rect 723 -824 766 -823
rect 835 -824 941 -823
rect 121 -826 136 -825
rect 138 -826 192 -825
rect 205 -826 283 -825
rect 289 -826 367 -825
rect 373 -826 724 -825
rect 730 -826 909 -825
rect 2 -828 206 -827
rect 219 -828 675 -827
rect 772 -828 836 -827
rect 128 -830 318 -829
rect 345 -830 416 -829
rect 516 -830 633 -829
rect 660 -830 675 -829
rect 772 -830 808 -829
rect 110 -832 661 -831
rect 670 -832 731 -831
rect 758 -832 808 -831
rect 117 -834 633 -833
rect 702 -834 759 -833
rect 131 -836 857 -835
rect 135 -838 878 -837
rect 142 -840 199 -839
rect 240 -840 444 -839
rect 534 -840 717 -839
rect 163 -842 171 -841
rect 191 -842 248 -841
rect 268 -842 409 -841
rect 415 -842 598 -841
rect 604 -842 689 -841
rect 156 -844 248 -843
rect 324 -844 605 -843
rect 611 -844 626 -843
rect 100 -846 325 -845
rect 355 -846 703 -845
rect 100 -848 332 -847
rect 355 -848 871 -847
rect 156 -850 209 -849
rect 331 -850 395 -849
rect 457 -850 598 -849
rect 793 -850 871 -849
rect 170 -852 178 -851
rect 198 -852 213 -851
rect 275 -852 395 -851
rect 457 -852 465 -851
rect 548 -852 794 -851
rect 177 -854 388 -853
rect 464 -854 927 -853
rect 212 -856 801 -855
rect 366 -858 573 -857
rect 579 -858 906 -857
rect 373 -860 535 -859
rect 548 -860 612 -859
rect 555 -862 857 -861
rect 359 -864 556 -863
rect 562 -864 885 -863
rect 275 -866 360 -865
rect 565 -866 787 -865
rect 565 -868 843 -867
rect 583 -870 591 -869
rect 779 -870 843 -869
rect 436 -872 584 -871
rect 436 -874 647 -873
rect 562 -876 780 -875
rect 569 -878 647 -877
rect 16 -889 115 -888
rect 135 -889 332 -888
rect 359 -889 584 -888
rect 600 -889 871 -888
rect 915 -889 920 -888
rect 954 -889 993 -888
rect 1013 -889 1025 -888
rect 1038 -889 1060 -888
rect 1080 -889 1088 -888
rect 16 -891 171 -890
rect 184 -891 356 -890
rect 366 -891 682 -890
rect 814 -891 822 -890
rect 870 -891 997 -890
rect 1010 -891 1039 -890
rect 23 -893 227 -892
rect 243 -893 276 -892
rect 289 -893 332 -892
rect 366 -893 423 -892
rect 429 -893 531 -892
rect 534 -893 780 -892
rect 817 -893 829 -892
rect 961 -893 1011 -892
rect 2 -895 24 -894
rect 51 -895 419 -894
rect 422 -895 524 -894
rect 534 -895 556 -894
rect 569 -895 899 -894
rect 961 -895 969 -894
rect 989 -895 1018 -894
rect 51 -897 150 -896
rect 156 -897 185 -896
rect 205 -897 276 -896
rect 289 -897 353 -896
rect 369 -897 514 -896
rect 520 -897 787 -896
rect 828 -897 850 -896
rect 891 -897 899 -896
rect 968 -897 976 -896
rect 58 -899 216 -898
rect 219 -899 738 -898
rect 765 -899 787 -898
rect 849 -899 885 -898
rect 891 -899 927 -898
rect 58 -901 388 -900
rect 408 -901 451 -900
rect 464 -901 472 -900
rect 474 -901 794 -900
rect 884 -901 934 -900
rect 65 -903 339 -902
rect 352 -903 374 -902
rect 387 -903 395 -902
rect 408 -903 577 -902
rect 628 -903 801 -902
rect 933 -903 941 -902
rect 72 -905 230 -904
rect 278 -905 521 -904
rect 527 -905 577 -904
rect 730 -905 822 -904
rect 72 -907 311 -906
rect 317 -907 493 -906
rect 499 -907 717 -906
rect 737 -907 745 -906
rect 751 -907 794 -906
rect 800 -907 843 -906
rect 93 -909 241 -908
rect 261 -909 318 -908
rect 324 -909 339 -908
rect 345 -909 493 -908
rect 499 -909 507 -908
rect 537 -909 542 -908
rect 548 -909 983 -908
rect 93 -911 598 -910
rect 635 -911 731 -910
rect 765 -911 836 -910
rect 842 -911 857 -910
rect 905 -911 983 -910
rect 107 -913 612 -912
rect 688 -913 717 -912
rect 723 -913 745 -912
rect 779 -913 944 -912
rect 107 -915 241 -914
rect 261 -915 304 -914
rect 310 -915 563 -914
rect 597 -915 668 -914
rect 702 -915 724 -914
rect 856 -915 864 -914
rect 905 -915 913 -914
rect 110 -917 255 -916
rect 285 -917 304 -916
rect 373 -917 573 -916
rect 604 -917 612 -916
rect 653 -917 703 -916
rect 709 -917 752 -916
rect 863 -917 878 -916
rect 912 -917 923 -916
rect 114 -919 192 -918
rect 198 -919 255 -918
rect 411 -919 710 -918
rect 149 -921 164 -920
rect 170 -921 237 -920
rect 429 -921 458 -920
rect 467 -921 647 -920
rect 660 -921 689 -920
rect 30 -923 164 -922
rect 180 -923 325 -922
rect 436 -923 549 -922
rect 551 -923 591 -922
rect 639 -923 647 -922
rect 660 -923 675 -922
rect 30 -925 216 -924
rect 439 -925 930 -924
rect 86 -927 181 -926
rect 191 -927 234 -926
rect 439 -927 507 -926
rect 513 -927 591 -926
rect 625 -927 675 -926
rect 86 -929 143 -928
rect 156 -929 269 -928
rect 443 -929 570 -928
rect 632 -929 640 -928
rect 37 -931 444 -930
rect 457 -931 486 -930
rect 502 -931 682 -930
rect 37 -933 132 -932
rect 142 -933 297 -932
rect 471 -933 584 -932
rect 173 -935 297 -934
rect 478 -935 486 -934
rect 555 -935 696 -934
rect 198 -937 605 -936
rect 695 -937 1004 -936
rect 208 -939 283 -938
rect 478 -939 878 -938
rect 44 -941 283 -940
rect 562 -941 836 -940
rect 44 -943 402 -942
rect 212 -945 223 -944
rect 233 -945 248 -944
rect 268 -945 381 -944
rect 401 -945 657 -944
rect 100 -947 248 -946
rect 79 -949 101 -948
rect 222 -949 346 -948
rect 79 -951 416 -950
rect 415 -953 759 -952
rect 758 -955 773 -954
rect 618 -957 773 -956
rect 618 -959 955 -958
rect 9 -970 374 -969
rect 380 -970 549 -969
rect 565 -970 822 -969
rect 835 -970 941 -969
rect 947 -970 997 -969
rect 1010 -970 1032 -969
rect 1038 -970 1074 -969
rect 1087 -970 1095 -969
rect 16 -972 472 -971
rect 474 -972 1077 -971
rect 16 -974 367 -973
rect 373 -974 402 -973
rect 408 -974 433 -973
rect 453 -974 465 -973
rect 481 -974 675 -973
rect 698 -974 871 -973
rect 891 -974 1046 -973
rect 1059 -974 1102 -973
rect 37 -976 209 -975
rect 226 -976 587 -975
rect 600 -976 731 -975
rect 751 -976 836 -975
rect 842 -976 948 -975
rect 954 -976 1088 -975
rect 58 -978 475 -977
rect 488 -978 577 -977
rect 607 -978 801 -977
rect 828 -978 843 -977
rect 863 -978 892 -977
rect 898 -978 990 -977
rect 30 -980 608 -979
rect 635 -980 1011 -979
rect 30 -982 199 -981
rect 240 -982 633 -981
rect 639 -982 675 -981
rect 681 -982 752 -981
rect 758 -982 913 -981
rect 919 -982 969 -981
rect 982 -982 1070 -981
rect 61 -984 633 -983
rect 653 -984 885 -983
rect 905 -984 1039 -983
rect 93 -986 244 -985
rect 247 -986 465 -985
rect 471 -986 955 -985
rect 100 -988 328 -987
rect 338 -988 412 -987
rect 418 -988 734 -987
rect 737 -988 829 -987
rect 856 -988 969 -987
rect 100 -990 220 -989
rect 247 -990 346 -989
rect 366 -990 458 -989
rect 492 -990 689 -989
rect 716 -990 759 -989
rect 765 -990 822 -989
rect 905 -990 916 -989
rect 929 -990 962 -989
rect 93 -992 493 -991
rect 495 -992 1018 -991
rect 114 -994 213 -993
rect 261 -994 346 -993
rect 380 -994 486 -993
rect 506 -994 682 -993
rect 730 -994 864 -993
rect 933 -994 983 -993
rect 114 -996 150 -995
rect 177 -996 356 -995
rect 383 -996 402 -995
rect 436 -996 766 -995
rect 793 -996 801 -995
rect 814 -996 885 -995
rect 943 -996 1060 -995
rect 121 -998 129 -997
rect 131 -998 976 -997
rect 72 -1000 122 -999
rect 131 -1000 227 -999
rect 261 -1000 423 -999
rect 457 -1000 542 -999
rect 548 -1000 871 -999
rect 65 -1002 423 -1001
rect 506 -1002 650 -1001
rect 660 -1002 738 -1001
rect 786 -1002 794 -1001
rect 814 -1002 1067 -1001
rect 65 -1004 157 -1003
rect 180 -1004 241 -1003
rect 282 -1004 563 -1003
rect 576 -1004 1053 -1003
rect 72 -1006 255 -1005
rect 285 -1006 780 -1005
rect 135 -1008 440 -1007
rect 450 -1008 780 -1007
rect 135 -1010 927 -1009
rect 142 -1012 531 -1011
rect 537 -1012 850 -1011
rect 44 -1014 143 -1013
rect 145 -1014 1004 -1013
rect 149 -1016 164 -1015
rect 180 -1016 276 -1015
rect 296 -1016 437 -1015
rect 450 -1016 927 -1015
rect 23 -1018 164 -1017
rect 191 -1018 234 -1017
rect 299 -1018 521 -1017
rect 527 -1018 668 -1017
rect 723 -1018 787 -1017
rect 849 -1018 878 -1017
rect 23 -1020 223 -1019
rect 303 -1020 563 -1019
rect 597 -1020 920 -1019
rect 40 -1022 192 -1021
rect 198 -1022 206 -1021
rect 257 -1022 598 -1021
rect 604 -1022 899 -1021
rect 51 -1024 297 -1023
rect 303 -1024 430 -1023
rect 443 -1024 668 -1023
rect 702 -1024 724 -1023
rect 807 -1024 878 -1023
rect 51 -1026 87 -1025
rect 156 -1026 206 -1025
rect 310 -1026 479 -1025
rect 499 -1026 521 -1025
rect 541 -1026 591 -1025
rect 604 -1026 934 -1025
rect 44 -1028 479 -1027
rect 499 -1028 923 -1027
rect 79 -1030 311 -1029
rect 317 -1030 339 -1029
rect 387 -1030 395 -1029
rect 397 -1030 416 -1029
rect 443 -1030 745 -1029
rect 79 -1032 360 -1031
rect 516 -1032 773 -1031
rect 268 -1034 318 -1033
rect 324 -1034 388 -1033
rect 429 -1034 773 -1033
rect 107 -1036 269 -1035
rect 331 -1036 360 -1035
rect 534 -1036 591 -1035
rect 611 -1036 654 -1035
rect 702 -1036 710 -1035
rect 107 -1038 171 -1037
rect 184 -1038 325 -1037
rect 331 -1038 353 -1037
rect 551 -1038 857 -1037
rect 12 -1040 353 -1039
rect 555 -1040 640 -1039
rect 646 -1040 661 -1039
rect 691 -1040 710 -1039
rect 184 -1042 290 -1041
rect 453 -1042 556 -1041
rect 569 -1042 612 -1041
rect 618 -1042 717 -1041
rect 289 -1044 363 -1043
rect 446 -1044 619 -1043
rect 625 -1044 962 -1043
rect 569 -1046 696 -1045
rect 583 -1048 745 -1047
rect 86 -1050 584 -1049
rect 628 -1050 808 -1049
rect 646 -1052 696 -1051
rect 16 -1063 451 -1062
rect 478 -1063 829 -1062
rect 961 -1063 1025 -1062
rect 1027 -1063 1053 -1062
rect 1059 -1063 1084 -1062
rect 1094 -1063 1098 -1062
rect 19 -1065 335 -1064
rect 338 -1065 444 -1064
rect 464 -1065 479 -1064
rect 495 -1065 878 -1064
rect 989 -1065 1060 -1064
rect 1094 -1065 1102 -1064
rect 30 -1067 38 -1066
rect 51 -1067 59 -1066
rect 65 -1067 146 -1066
rect 156 -1067 181 -1066
rect 191 -1067 195 -1066
rect 219 -1067 230 -1066
rect 275 -1067 549 -1066
rect 569 -1067 899 -1066
rect 996 -1067 1053 -1066
rect 51 -1069 132 -1068
rect 142 -1069 265 -1068
rect 282 -1069 475 -1068
rect 513 -1069 577 -1068
rect 579 -1069 871 -1068
rect 1017 -1069 1074 -1068
rect 58 -1071 356 -1070
rect 369 -1071 934 -1070
rect 65 -1073 262 -1072
rect 296 -1073 374 -1072
rect 387 -1073 514 -1072
rect 576 -1073 601 -1072
rect 604 -1073 829 -1072
rect 926 -1073 1018 -1072
rect 2 -1075 262 -1074
rect 303 -1075 468 -1074
rect 583 -1075 1046 -1074
rect 79 -1077 188 -1076
rect 191 -1077 213 -1076
rect 222 -1077 346 -1076
rect 352 -1077 941 -1076
rect 114 -1079 174 -1078
rect 177 -1079 199 -1078
rect 233 -1079 276 -1078
rect 310 -1079 496 -1078
rect 569 -1079 584 -1078
rect 586 -1079 913 -1078
rect 940 -1079 1088 -1078
rect 1097 -1079 1102 -1078
rect 93 -1081 115 -1080
rect 121 -1081 255 -1080
rect 317 -1081 444 -1080
rect 572 -1081 1046 -1080
rect 44 -1083 122 -1082
rect 156 -1083 290 -1082
rect 324 -1083 454 -1082
rect 593 -1083 955 -1082
rect 44 -1085 538 -1084
rect 597 -1085 608 -1084
rect 621 -1085 997 -1084
rect 93 -1087 244 -1086
rect 247 -1087 283 -1086
rect 289 -1087 332 -1086
rect 338 -1087 437 -1086
rect 439 -1087 542 -1086
rect 628 -1087 836 -1086
rect 863 -1087 927 -1086
rect 135 -1089 325 -1088
rect 345 -1089 591 -1088
rect 628 -1089 948 -1088
rect 107 -1091 136 -1090
rect 163 -1091 493 -1090
rect 509 -1091 948 -1090
rect 107 -1093 171 -1092
rect 184 -1093 318 -1092
rect 359 -1093 374 -1092
rect 387 -1093 402 -1092
rect 408 -1093 864 -1092
rect 912 -1093 983 -1092
rect 100 -1095 171 -1094
rect 198 -1095 381 -1094
rect 394 -1095 409 -1094
rect 411 -1095 447 -1094
rect 541 -1095 1070 -1094
rect 9 -1097 101 -1096
rect 166 -1097 962 -1096
rect 240 -1099 311 -1098
rect 359 -1099 447 -1098
rect 590 -1099 885 -1098
rect 919 -1099 955 -1098
rect 247 -1101 598 -1100
rect 646 -1101 678 -1100
rect 688 -1101 906 -1100
rect 919 -1101 1081 -1100
rect 380 -1103 507 -1102
rect 649 -1103 969 -1102
rect 1003 -1103 1081 -1102
rect 72 -1105 507 -1104
rect 688 -1105 983 -1104
rect 23 -1107 73 -1106
rect 394 -1107 563 -1106
rect 723 -1107 836 -1106
rect 849 -1107 969 -1106
rect 23 -1109 129 -1108
rect 401 -1109 535 -1108
rect 555 -1109 563 -1108
rect 639 -1109 724 -1108
rect 726 -1109 899 -1108
rect 422 -1111 552 -1110
rect 555 -1111 612 -1110
rect 730 -1111 990 -1110
rect 268 -1113 423 -1112
rect 429 -1113 668 -1112
rect 730 -1113 1039 -1112
rect 429 -1115 528 -1114
rect 611 -1115 633 -1114
rect 667 -1115 752 -1114
rect 765 -1115 850 -1114
rect 856 -1115 906 -1114
rect 1038 -1115 1077 -1114
rect 436 -1117 1067 -1116
rect 457 -1119 647 -1118
rect 779 -1119 871 -1118
rect 457 -1121 500 -1120
rect 520 -1121 535 -1120
rect 618 -1121 752 -1120
rect 786 -1121 1004 -1120
rect 226 -1123 500 -1122
rect 520 -1123 661 -1122
rect 716 -1123 780 -1122
rect 800 -1123 885 -1122
rect 226 -1125 269 -1124
rect 530 -1125 766 -1124
rect 800 -1125 815 -1124
rect 821 -1125 878 -1124
rect 632 -1127 738 -1126
rect 758 -1127 822 -1126
rect 653 -1129 787 -1128
rect 807 -1129 857 -1128
rect 653 -1131 745 -1130
rect 772 -1131 815 -1130
rect 240 -1133 745 -1132
rect 807 -1133 892 -1132
rect 660 -1135 1011 -1134
rect 681 -1137 717 -1136
rect 793 -1137 892 -1136
rect 1010 -1137 1032 -1136
rect 299 -1139 682 -1138
rect 695 -1139 738 -1138
rect 842 -1139 1032 -1138
rect 492 -1141 794 -1140
rect 842 -1141 976 -1140
rect 485 -1143 976 -1142
rect 366 -1145 486 -1144
rect 674 -1145 696 -1144
rect 702 -1145 773 -1144
rect 366 -1147 416 -1146
rect 642 -1147 703 -1146
rect 709 -1147 759 -1146
rect 149 -1149 416 -1148
rect 674 -1149 934 -1148
rect 149 -1151 237 -1150
rect 709 -1151 1088 -1150
rect 30 -1162 587 -1161
rect 590 -1162 622 -1161
rect 639 -1162 892 -1161
rect 1090 -1162 1102 -1161
rect 30 -1164 150 -1163
rect 156 -1164 237 -1163
rect 243 -1164 311 -1163
rect 331 -1164 920 -1163
rect 33 -1166 94 -1165
rect 121 -1166 150 -1165
rect 156 -1166 367 -1165
rect 429 -1166 461 -1165
rect 464 -1166 1081 -1165
rect 51 -1168 367 -1167
rect 436 -1168 1042 -1167
rect 58 -1170 83 -1169
rect 93 -1170 164 -1169
rect 194 -1170 241 -1169
rect 247 -1170 465 -1169
rect 471 -1170 1025 -1169
rect 58 -1172 87 -1171
rect 114 -1172 122 -1171
rect 128 -1172 388 -1171
rect 439 -1172 479 -1171
rect 495 -1172 850 -1171
rect 891 -1172 997 -1171
rect 51 -1174 87 -1173
rect 114 -1174 682 -1173
rect 684 -1174 1004 -1173
rect 82 -1176 101 -1175
rect 128 -1176 136 -1175
rect 163 -1176 955 -1175
rect 135 -1178 213 -1177
rect 226 -1178 626 -1177
rect 639 -1178 773 -1177
rect 842 -1178 1004 -1177
rect 117 -1180 626 -1179
rect 642 -1180 738 -1179
rect 772 -1180 829 -1179
rect 842 -1180 1088 -1179
rect 170 -1182 241 -1181
rect 247 -1182 395 -1181
rect 446 -1182 535 -1181
rect 544 -1182 801 -1181
rect 919 -1182 990 -1181
rect 184 -1184 990 -1183
rect 37 -1186 185 -1185
rect 198 -1186 479 -1185
rect 495 -1186 787 -1185
rect 954 -1186 1067 -1185
rect 37 -1188 167 -1187
rect 226 -1188 318 -1187
rect 331 -1188 346 -1187
rect 352 -1188 374 -1187
rect 380 -1188 437 -1187
rect 450 -1188 528 -1187
rect 548 -1188 552 -1187
rect 590 -1188 997 -1187
rect 79 -1190 346 -1189
rect 380 -1190 402 -1189
rect 450 -1190 486 -1189
rect 509 -1190 1018 -1189
rect 79 -1192 507 -1191
rect 513 -1192 584 -1191
rect 597 -1192 1032 -1191
rect 44 -1194 514 -1193
rect 516 -1194 850 -1193
rect 1010 -1194 1018 -1193
rect 44 -1196 171 -1195
rect 229 -1196 276 -1195
rect 282 -1196 566 -1195
rect 600 -1196 941 -1195
rect 72 -1198 598 -1197
rect 604 -1198 717 -1197
rect 723 -1198 1053 -1197
rect 26 -1200 605 -1199
rect 618 -1200 647 -1199
rect 660 -1200 829 -1199
rect 835 -1200 1053 -1199
rect 72 -1202 325 -1201
rect 387 -1202 570 -1201
rect 618 -1202 629 -1201
rect 660 -1202 696 -1201
rect 716 -1202 885 -1201
rect 912 -1202 1011 -1201
rect 107 -1204 325 -1203
rect 394 -1204 416 -1203
rect 485 -1204 710 -1203
rect 723 -1204 815 -1203
rect 884 -1204 983 -1203
rect 107 -1206 199 -1205
rect 233 -1206 307 -1205
rect 310 -1206 542 -1205
rect 555 -1206 647 -1205
rect 667 -1206 689 -1205
rect 691 -1206 1025 -1205
rect 219 -1208 234 -1207
rect 254 -1208 318 -1207
rect 401 -1208 409 -1207
rect 492 -1208 668 -1207
rect 677 -1208 1046 -1207
rect 16 -1210 255 -1209
rect 261 -1210 549 -1209
rect 555 -1210 577 -1209
rect 586 -1210 913 -1209
rect 1045 -1210 1074 -1209
rect 177 -1212 220 -1211
rect 264 -1212 675 -1211
rect 695 -1212 766 -1211
rect 814 -1212 1039 -1211
rect 1073 -1212 1095 -1211
rect 177 -1214 524 -1213
rect 541 -1214 1032 -1213
rect 1038 -1214 1067 -1213
rect 268 -1216 416 -1215
rect 502 -1216 836 -1215
rect 856 -1216 983 -1215
rect 268 -1218 472 -1217
rect 520 -1218 531 -1217
rect 562 -1218 577 -1217
rect 653 -1218 766 -1217
rect 807 -1218 857 -1217
rect 275 -1220 360 -1219
rect 408 -1220 475 -1219
rect 562 -1220 822 -1219
rect 282 -1222 657 -1221
rect 709 -1222 720 -1221
rect 730 -1222 878 -1221
rect 142 -1224 878 -1223
rect 2 -1226 143 -1225
rect 289 -1226 430 -1225
rect 457 -1226 475 -1225
rect 569 -1226 780 -1225
rect 807 -1226 906 -1225
rect 2 -1228 206 -1227
rect 292 -1228 734 -1227
rect 737 -1228 745 -1227
rect 758 -1228 801 -1227
rect 821 -1228 871 -1227
rect 9 -1230 290 -1229
rect 296 -1230 374 -1229
rect 663 -1230 906 -1229
rect 9 -1232 216 -1231
rect 296 -1232 500 -1231
rect 702 -1232 745 -1231
rect 751 -1232 759 -1231
rect 779 -1232 941 -1231
rect 23 -1234 458 -1233
rect 499 -1234 633 -1233
rect 681 -1234 703 -1233
rect 751 -1234 783 -1233
rect 870 -1234 948 -1233
rect 23 -1236 934 -1235
rect 947 -1236 976 -1235
rect 191 -1238 206 -1237
rect 303 -1238 468 -1237
rect 933 -1238 1060 -1237
rect 100 -1240 192 -1239
rect 338 -1240 360 -1239
rect 422 -1240 633 -1239
rect 793 -1240 1060 -1239
rect 338 -1242 594 -1241
rect 961 -1242 976 -1241
rect 355 -1244 423 -1243
rect 443 -1244 794 -1243
rect 961 -1244 969 -1243
rect 443 -1246 608 -1245
rect 898 -1246 969 -1245
rect 863 -1248 899 -1247
rect 863 -1250 927 -1249
rect 187 -1252 927 -1251
rect 187 -1254 787 -1253
rect 2 -1265 517 -1264
rect 520 -1265 801 -1264
rect 814 -1265 843 -1264
rect 870 -1265 874 -1264
rect 982 -1265 1063 -1264
rect 1066 -1265 1081 -1264
rect 9 -1267 17 -1266
rect 30 -1267 167 -1266
rect 170 -1267 241 -1266
rect 254 -1267 503 -1266
rect 513 -1267 822 -1266
rect 870 -1267 927 -1266
rect 947 -1267 983 -1266
rect 1017 -1267 1021 -1266
rect 9 -1269 59 -1268
rect 86 -1269 591 -1268
rect 604 -1269 780 -1268
rect 912 -1269 948 -1268
rect 1017 -1269 1053 -1268
rect 30 -1271 87 -1270
rect 93 -1271 216 -1270
rect 219 -1271 234 -1270
rect 240 -1271 262 -1270
rect 317 -1271 328 -1270
rect 331 -1271 461 -1270
rect 464 -1271 521 -1270
rect 541 -1271 1004 -1270
rect 1020 -1271 1053 -1270
rect 51 -1273 297 -1272
rect 320 -1273 479 -1272
rect 548 -1273 731 -1272
rect 751 -1273 1067 -1272
rect 51 -1275 150 -1274
rect 159 -1275 472 -1274
rect 478 -1275 696 -1274
rect 761 -1275 822 -1274
rect 884 -1275 913 -1274
rect 1003 -1275 1035 -1274
rect 54 -1277 311 -1276
rect 366 -1277 496 -1276
rect 576 -1277 584 -1276
rect 586 -1277 689 -1276
rect 884 -1277 892 -1276
rect 58 -1279 283 -1278
rect 292 -1279 731 -1278
rect 835 -1279 892 -1278
rect 65 -1281 150 -1280
rect 170 -1281 675 -1280
rect 677 -1281 1011 -1280
rect 65 -1283 339 -1282
rect 369 -1283 528 -1282
rect 555 -1283 577 -1282
rect 583 -1283 633 -1282
rect 639 -1283 696 -1282
rect 817 -1283 836 -1282
rect 954 -1283 1011 -1282
rect 93 -1285 101 -1284
rect 114 -1285 132 -1284
rect 135 -1285 318 -1284
rect 331 -1285 367 -1284
rect 422 -1285 549 -1284
rect 565 -1285 640 -1284
rect 653 -1285 962 -1284
rect 100 -1287 122 -1286
rect 142 -1287 290 -1286
rect 292 -1287 325 -1286
rect 338 -1287 353 -1286
rect 425 -1287 437 -1286
rect 443 -1287 542 -1286
rect 604 -1287 612 -1286
rect 625 -1287 633 -1286
rect 653 -1287 1060 -1286
rect 23 -1289 122 -1288
rect 142 -1289 227 -1288
rect 261 -1289 276 -1288
rect 282 -1289 360 -1288
rect 415 -1289 437 -1288
rect 443 -1289 475 -1288
rect 527 -1289 535 -1288
rect 537 -1289 556 -1288
rect 607 -1289 857 -1288
rect 940 -1289 962 -1288
rect 23 -1291 108 -1290
rect 117 -1291 738 -1290
rect 751 -1291 1060 -1290
rect 72 -1293 353 -1292
rect 359 -1293 766 -1292
rect 793 -1293 857 -1292
rect 919 -1293 941 -1292
rect 72 -1295 388 -1294
rect 464 -1295 507 -1294
rect 537 -1295 647 -1294
rect 656 -1295 990 -1294
rect 107 -1297 139 -1296
rect 163 -1297 626 -1296
rect 660 -1297 843 -1296
rect 849 -1297 920 -1296
rect 968 -1297 990 -1296
rect 117 -1299 311 -1298
rect 373 -1299 388 -1298
rect 611 -1299 619 -1298
rect 660 -1299 703 -1298
rect 716 -1299 766 -1298
rect 793 -1299 1039 -1298
rect 128 -1301 164 -1300
rect 173 -1301 1025 -1300
rect 187 -1303 997 -1302
rect 191 -1305 976 -1304
rect 996 -1305 1032 -1304
rect 194 -1307 248 -1306
rect 268 -1307 647 -1306
rect 667 -1307 801 -1306
rect 807 -1307 955 -1306
rect 194 -1309 255 -1308
rect 268 -1309 346 -1308
rect 373 -1309 486 -1308
rect 667 -1309 1042 -1308
rect 198 -1311 223 -1310
rect 247 -1311 451 -1310
rect 485 -1311 622 -1310
rect 681 -1311 773 -1310
rect 786 -1311 808 -1310
rect 905 -1311 969 -1310
rect 184 -1313 223 -1312
rect 275 -1313 545 -1312
rect 562 -1313 773 -1312
rect 933 -1313 976 -1312
rect 44 -1315 185 -1314
rect 201 -1315 395 -1314
rect 432 -1315 451 -1314
rect 509 -1315 563 -1314
rect 688 -1315 710 -1314
rect 716 -1315 759 -1314
rect 877 -1315 934 -1314
rect 44 -1317 178 -1316
rect 205 -1317 234 -1316
rect 296 -1317 500 -1316
rect 709 -1317 724 -1316
rect 758 -1317 906 -1316
rect 156 -1319 206 -1318
rect 212 -1319 227 -1318
rect 345 -1319 458 -1318
rect 499 -1319 1049 -1318
rect 212 -1321 304 -1320
rect 355 -1321 787 -1320
rect 828 -1321 878 -1320
rect 37 -1323 304 -1322
rect 380 -1323 395 -1322
rect 432 -1323 514 -1322
rect 597 -1323 724 -1322
rect 37 -1325 220 -1324
rect 380 -1325 402 -1324
rect 422 -1325 598 -1324
rect 401 -1327 409 -1326
rect 457 -1327 850 -1326
rect 408 -1329 570 -1328
rect 492 -1331 829 -1330
rect 415 -1333 493 -1332
rect 569 -1333 580 -1332
rect 16 -1344 80 -1343
rect 89 -1344 297 -1343
rect 303 -1344 328 -1343
rect 352 -1344 381 -1343
rect 387 -1344 433 -1343
rect 471 -1344 633 -1343
rect 646 -1344 906 -1343
rect 950 -1344 997 -1343
rect 1031 -1344 1053 -1343
rect 16 -1346 174 -1345
rect 222 -1346 283 -1345
rect 292 -1346 535 -1345
rect 576 -1346 843 -1345
rect 891 -1346 906 -1345
rect 1024 -1346 1032 -1345
rect 1038 -1346 1074 -1345
rect 23 -1348 87 -1347
rect 107 -1348 171 -1347
rect 222 -1348 311 -1347
rect 338 -1348 353 -1347
rect 366 -1348 451 -1347
rect 471 -1348 591 -1347
rect 597 -1348 913 -1347
rect 971 -1348 1025 -1347
rect 1045 -1348 1049 -1347
rect 1073 -1348 1081 -1347
rect 9 -1350 87 -1349
rect 107 -1350 332 -1349
rect 338 -1350 465 -1349
rect 495 -1350 724 -1349
rect 737 -1350 871 -1349
rect 30 -1352 62 -1351
rect 65 -1352 69 -1351
rect 79 -1352 356 -1351
rect 380 -1352 395 -1351
rect 411 -1352 563 -1351
rect 576 -1352 682 -1351
rect 705 -1352 745 -1351
rect 758 -1352 976 -1351
rect 30 -1354 101 -1353
rect 114 -1354 220 -1353
rect 254 -1354 311 -1353
rect 331 -1354 549 -1353
rect 579 -1354 941 -1353
rect 961 -1354 976 -1353
rect 37 -1356 136 -1355
rect 138 -1356 402 -1355
rect 415 -1356 458 -1355
rect 506 -1356 689 -1355
rect 705 -1356 1018 -1355
rect 37 -1358 45 -1357
rect 51 -1358 178 -1357
rect 254 -1358 507 -1357
rect 509 -1358 696 -1357
rect 723 -1358 787 -1357
rect 835 -1358 892 -1357
rect 44 -1360 346 -1359
rect 401 -1360 570 -1359
rect 590 -1360 605 -1359
rect 618 -1360 969 -1359
rect 54 -1362 601 -1361
rect 611 -1362 619 -1361
rect 632 -1362 752 -1361
rect 758 -1362 780 -1361
rect 835 -1362 857 -1361
rect 863 -1362 962 -1361
rect 65 -1364 94 -1363
rect 100 -1364 423 -1363
rect 429 -1364 997 -1363
rect 93 -1366 479 -1365
rect 523 -1366 605 -1365
rect 611 -1366 675 -1365
rect 684 -1366 941 -1365
rect 121 -1368 195 -1367
rect 247 -1368 346 -1367
rect 355 -1368 423 -1367
rect 429 -1368 517 -1367
rect 548 -1368 678 -1367
rect 688 -1368 703 -1367
rect 709 -1368 787 -1367
rect 842 -1368 899 -1367
rect 58 -1370 122 -1369
rect 128 -1370 514 -1369
rect 572 -1370 752 -1369
rect 765 -1370 1053 -1369
rect 128 -1372 209 -1371
rect 268 -1372 297 -1371
rect 303 -1372 710 -1371
rect 730 -1372 745 -1371
rect 779 -1372 801 -1371
rect 849 -1372 913 -1371
rect 145 -1374 157 -1373
rect 159 -1374 542 -1373
rect 579 -1374 864 -1373
rect 870 -1374 878 -1373
rect 884 -1374 899 -1373
rect 149 -1376 269 -1375
rect 275 -1376 395 -1375
rect 415 -1376 664 -1375
rect 674 -1376 717 -1375
rect 737 -1376 773 -1375
rect 800 -1376 808 -1375
rect 884 -1376 983 -1375
rect 149 -1378 181 -1377
rect 184 -1378 248 -1377
rect 261 -1378 276 -1377
rect 282 -1378 388 -1377
rect 450 -1378 500 -1377
rect 583 -1378 857 -1377
rect 982 -1378 990 -1377
rect 163 -1380 192 -1379
rect 205 -1380 262 -1379
rect 324 -1380 479 -1379
rect 492 -1380 808 -1379
rect 23 -1382 206 -1381
rect 324 -1382 374 -1381
rect 443 -1382 500 -1381
rect 583 -1382 955 -1381
rect 68 -1384 374 -1383
rect 443 -1384 486 -1383
rect 492 -1384 521 -1383
rect 586 -1384 990 -1383
rect 163 -1386 290 -1385
rect 359 -1386 731 -1385
rect 772 -1386 829 -1385
rect 947 -1386 955 -1385
rect 177 -1388 199 -1387
rect 359 -1388 437 -1387
rect 464 -1388 570 -1387
rect 597 -1388 1067 -1387
rect 184 -1390 318 -1389
rect 369 -1390 850 -1389
rect 198 -1392 234 -1391
rect 317 -1392 461 -1391
rect 485 -1392 556 -1391
rect 565 -1392 829 -1391
rect 72 -1394 556 -1393
rect 646 -1394 654 -1393
rect 660 -1394 717 -1393
rect 72 -1396 227 -1395
rect 408 -1396 521 -1395
rect 653 -1396 1035 -1395
rect 142 -1398 227 -1397
rect 408 -1398 542 -1397
rect 660 -1398 1011 -1397
rect 212 -1400 234 -1399
rect 436 -1400 528 -1399
rect 681 -1400 878 -1399
rect 1003 -1400 1011 -1399
rect 212 -1402 241 -1401
rect 527 -1402 626 -1401
rect 695 -1402 815 -1401
rect 1003 -1402 1018 -1401
rect 625 -1404 668 -1403
rect 814 -1404 934 -1403
rect 639 -1406 668 -1405
rect 926 -1406 934 -1405
rect 639 -1408 794 -1407
rect 649 -1410 794 -1409
rect 16 -1421 125 -1420
rect 135 -1421 297 -1420
rect 310 -1421 360 -1420
rect 390 -1421 451 -1420
rect 471 -1421 538 -1420
rect 569 -1421 675 -1420
rect 681 -1421 801 -1420
rect 828 -1421 832 -1420
rect 842 -1421 944 -1420
rect 971 -1421 1032 -1420
rect 1066 -1421 1074 -1420
rect 23 -1423 223 -1422
rect 268 -1423 307 -1422
rect 310 -1423 738 -1422
rect 793 -1423 951 -1422
rect 975 -1423 1004 -1422
rect 1010 -1423 1039 -1422
rect 30 -1425 160 -1424
rect 163 -1425 304 -1424
rect 338 -1425 563 -1424
rect 579 -1425 787 -1424
rect 793 -1425 822 -1424
rect 828 -1425 850 -1424
rect 877 -1425 969 -1424
rect 1024 -1425 1042 -1424
rect 30 -1427 52 -1426
rect 54 -1427 129 -1426
rect 138 -1427 143 -1426
rect 163 -1427 213 -1426
rect 219 -1427 654 -1426
rect 663 -1427 780 -1426
rect 821 -1427 906 -1426
rect 929 -1427 962 -1426
rect 44 -1429 129 -1428
rect 142 -1429 171 -1428
rect 205 -1429 892 -1428
rect 44 -1431 188 -1430
rect 205 -1431 241 -1430
rect 289 -1431 472 -1430
rect 499 -1431 514 -1430
rect 516 -1431 717 -1430
rect 744 -1431 976 -1430
rect 58 -1433 685 -1432
rect 688 -1433 717 -1432
rect 723 -1433 745 -1432
rect 772 -1433 787 -1432
rect 835 -1433 850 -1432
rect 877 -1433 927 -1432
rect 72 -1435 402 -1434
rect 408 -1435 521 -1434
rect 523 -1435 626 -1434
rect 635 -1435 808 -1434
rect 835 -1435 871 -1434
rect 884 -1435 923 -1434
rect 926 -1435 955 -1434
rect 37 -1437 73 -1436
rect 75 -1437 297 -1436
rect 338 -1437 587 -1436
rect 597 -1437 689 -1436
rect 712 -1437 815 -1436
rect 842 -1437 941 -1436
rect 954 -1437 1018 -1436
rect 37 -1439 150 -1438
rect 170 -1439 178 -1438
rect 212 -1439 318 -1438
rect 345 -1439 388 -1438
rect 394 -1439 409 -1438
rect 411 -1439 486 -1438
rect 513 -1439 710 -1438
rect 765 -1439 885 -1438
rect 86 -1441 780 -1440
rect 807 -1441 857 -1440
rect 870 -1441 990 -1440
rect 26 -1443 87 -1442
rect 89 -1443 773 -1442
rect 814 -1443 864 -1442
rect 947 -1443 990 -1442
rect 93 -1445 500 -1444
rect 555 -1445 570 -1444
rect 583 -1445 619 -1444
rect 639 -1445 675 -1444
rect 681 -1445 899 -1444
rect 912 -1445 948 -1444
rect 93 -1447 199 -1446
rect 219 -1447 262 -1446
rect 292 -1447 346 -1446
rect 352 -1447 542 -1446
rect 555 -1447 612 -1446
rect 632 -1447 640 -1446
rect 646 -1447 710 -1446
rect 726 -1447 899 -1446
rect 100 -1449 566 -1448
rect 604 -1449 769 -1448
rect 831 -1449 913 -1448
rect 79 -1451 101 -1450
rect 107 -1451 657 -1450
rect 660 -1451 892 -1450
rect 79 -1453 325 -1452
rect 362 -1453 598 -1452
rect 611 -1453 731 -1452
rect 751 -1453 766 -1452
rect 856 -1453 920 -1452
rect 107 -1455 577 -1454
rect 667 -1455 731 -1454
rect 863 -1455 934 -1454
rect 121 -1457 244 -1456
rect 247 -1457 325 -1456
rect 397 -1457 1053 -1456
rect 121 -1459 269 -1458
rect 317 -1459 416 -1458
rect 418 -1459 458 -1458
rect 478 -1459 605 -1458
rect 702 -1459 752 -1458
rect 919 -1459 1046 -1458
rect 149 -1461 430 -1460
rect 450 -1461 465 -1460
rect 478 -1461 591 -1460
rect 695 -1461 703 -1460
rect 933 -1461 997 -1460
rect 166 -1463 584 -1462
rect 590 -1463 1007 -1462
rect 177 -1465 192 -1464
rect 198 -1465 395 -1464
rect 401 -1465 559 -1464
rect 562 -1465 668 -1464
rect 695 -1465 941 -1464
rect 982 -1465 997 -1464
rect 184 -1467 262 -1466
rect 366 -1467 430 -1466
rect 457 -1467 535 -1466
rect 618 -1467 983 -1466
rect 184 -1469 332 -1468
rect 366 -1469 374 -1468
rect 415 -1469 626 -1468
rect 191 -1471 507 -1470
rect 527 -1471 647 -1470
rect 243 -1473 661 -1472
rect 247 -1475 307 -1474
rect 320 -1475 332 -1474
rect 355 -1475 374 -1474
rect 443 -1475 528 -1474
rect 51 -1477 444 -1476
rect 464 -1477 493 -1476
rect 506 -1477 549 -1476
rect 254 -1479 290 -1478
rect 422 -1479 493 -1478
rect 548 -1479 972 -1478
rect 233 -1481 255 -1480
rect 422 -1481 437 -1480
rect 485 -1481 545 -1480
rect 114 -1483 234 -1482
rect 436 -1483 906 -1482
rect 114 -1485 283 -1484
rect 275 -1487 283 -1486
rect 226 -1489 276 -1488
rect 156 -1491 227 -1490
rect 9 -1502 402 -1501
rect 418 -1502 493 -1501
rect 506 -1502 545 -1501
rect 558 -1502 766 -1501
rect 800 -1502 836 -1501
rect 856 -1502 969 -1501
rect 1038 -1502 1074 -1501
rect 16 -1504 150 -1503
rect 194 -1504 500 -1503
rect 506 -1504 713 -1503
rect 726 -1504 808 -1503
rect 835 -1504 1112 -1503
rect 23 -1506 164 -1505
rect 226 -1506 360 -1505
rect 394 -1506 1102 -1505
rect 30 -1508 244 -1507
rect 268 -1508 318 -1507
rect 327 -1508 626 -1507
rect 667 -1508 766 -1507
rect 870 -1508 1067 -1507
rect 30 -1510 143 -1509
rect 149 -1510 398 -1509
rect 418 -1510 521 -1509
rect 534 -1510 808 -1509
rect 870 -1510 983 -1509
rect 1003 -1510 1039 -1509
rect 37 -1512 241 -1511
rect 268 -1512 325 -1511
rect 341 -1512 829 -1511
rect 842 -1512 1004 -1511
rect 37 -1514 657 -1513
rect 681 -1514 885 -1513
rect 891 -1514 1109 -1513
rect 51 -1516 101 -1515
rect 121 -1516 941 -1515
rect 947 -1516 972 -1515
rect 58 -1518 125 -1517
rect 128 -1518 157 -1517
rect 163 -1518 213 -1517
rect 229 -1518 262 -1517
rect 275 -1518 304 -1517
rect 317 -1518 479 -1517
rect 513 -1518 556 -1517
rect 562 -1518 703 -1517
rect 733 -1518 1081 -1517
rect 58 -1520 377 -1519
rect 422 -1520 626 -1519
rect 646 -1520 983 -1519
rect 65 -1522 87 -1521
rect 93 -1522 314 -1521
rect 352 -1522 440 -1521
rect 450 -1522 514 -1521
rect 520 -1522 538 -1521
rect 562 -1522 598 -1521
rect 618 -1522 843 -1521
rect 877 -1522 1018 -1521
rect 44 -1524 66 -1523
rect 72 -1524 829 -1523
rect 877 -1524 934 -1523
rect 954 -1524 1095 -1523
rect 79 -1526 545 -1525
rect 565 -1526 815 -1525
rect 898 -1526 1025 -1525
rect 79 -1528 549 -1527
rect 618 -1528 696 -1527
rect 702 -1528 731 -1527
rect 744 -1528 857 -1527
rect 898 -1528 976 -1527
rect 82 -1530 479 -1529
rect 534 -1530 1088 -1529
rect 86 -1532 171 -1531
rect 177 -1532 227 -1531
rect 247 -1532 276 -1531
rect 282 -1532 353 -1531
rect 359 -1532 633 -1531
rect 646 -1532 801 -1531
rect 863 -1532 976 -1531
rect 93 -1534 416 -1533
rect 436 -1534 804 -1533
rect 905 -1534 1053 -1533
rect 100 -1536 241 -1535
rect 254 -1536 304 -1535
rect 306 -1536 906 -1535
rect 912 -1536 920 -1535
rect 922 -1536 962 -1535
rect 964 -1536 990 -1535
rect 135 -1538 395 -1537
rect 464 -1538 500 -1537
rect 548 -1538 612 -1537
rect 653 -1538 948 -1537
rect 135 -1540 458 -1539
rect 474 -1540 710 -1539
rect 716 -1540 815 -1539
rect 926 -1540 1032 -1539
rect 142 -1542 346 -1541
rect 362 -1542 955 -1541
rect 156 -1544 430 -1543
rect 569 -1544 612 -1543
rect 674 -1544 892 -1543
rect 180 -1546 213 -1545
rect 219 -1546 283 -1545
rect 289 -1546 577 -1545
rect 590 -1546 654 -1545
rect 660 -1546 675 -1545
rect 681 -1546 822 -1545
rect 184 -1548 325 -1547
rect 331 -1548 598 -1547
rect 604 -1548 717 -1547
rect 751 -1548 864 -1547
rect 107 -1550 332 -1549
rect 338 -1550 570 -1549
rect 590 -1550 689 -1549
rect 695 -1550 738 -1549
rect 758 -1550 1046 -1549
rect 107 -1552 115 -1551
rect 170 -1552 339 -1551
rect 345 -1552 444 -1551
rect 460 -1552 738 -1551
rect 758 -1552 913 -1551
rect 114 -1554 451 -1553
rect 485 -1554 752 -1553
rect 772 -1554 885 -1553
rect 187 -1556 440 -1555
rect 471 -1556 486 -1555
rect 663 -1556 689 -1555
rect 709 -1556 1011 -1555
rect 222 -1558 661 -1557
rect 684 -1558 990 -1557
rect 233 -1560 458 -1559
rect 723 -1560 773 -1559
rect 786 -1560 934 -1559
rect 233 -1562 668 -1561
rect 723 -1562 780 -1561
rect 793 -1562 927 -1561
rect 131 -1564 794 -1563
rect 803 -1564 1060 -1563
rect 243 -1566 577 -1565
rect 583 -1566 787 -1565
rect 821 -1566 850 -1565
rect 247 -1568 685 -1567
rect 254 -1570 293 -1569
rect 296 -1570 605 -1569
rect 639 -1570 780 -1569
rect 198 -1572 297 -1571
rect 310 -1572 745 -1571
rect 75 -1574 311 -1573
rect 373 -1574 465 -1573
rect 527 -1574 640 -1573
rect 2 -1576 374 -1575
rect 387 -1576 423 -1575
rect 495 -1576 528 -1575
rect 579 -1576 850 -1575
rect 198 -1578 206 -1577
rect 261 -1578 472 -1577
rect 191 -1580 206 -1579
rect 387 -1580 517 -1579
rect 397 -1582 444 -1581
rect 401 -1584 584 -1583
rect 408 -1586 430 -1585
rect 355 -1588 409 -1587
rect 2 -1599 300 -1598
rect 303 -1599 325 -1598
rect 355 -1599 787 -1598
rect 803 -1599 1032 -1598
rect 2 -1601 160 -1600
rect 163 -1601 342 -1600
rect 359 -1601 430 -1600
rect 453 -1601 983 -1600
rect 23 -1603 251 -1602
rect 261 -1603 353 -1602
rect 373 -1603 584 -1602
rect 660 -1603 689 -1602
rect 709 -1603 1095 -1602
rect 23 -1605 108 -1604
rect 121 -1605 794 -1604
rect 824 -1605 920 -1604
rect 982 -1605 1081 -1604
rect 30 -1607 234 -1606
rect 236 -1607 255 -1606
rect 282 -1607 416 -1606
rect 429 -1607 528 -1606
rect 555 -1607 710 -1606
rect 723 -1607 801 -1606
rect 849 -1607 916 -1606
rect 919 -1607 969 -1606
rect 30 -1609 486 -1608
rect 492 -1609 591 -1608
rect 663 -1609 892 -1608
rect 37 -1611 48 -1610
rect 61 -1611 451 -1610
rect 453 -1611 899 -1610
rect 37 -1613 129 -1612
rect 135 -1613 363 -1612
rect 376 -1613 381 -1612
rect 390 -1613 577 -1612
rect 583 -1613 612 -1612
rect 681 -1613 738 -1612
rect 758 -1613 1046 -1612
rect 72 -1615 829 -1614
rect 891 -1615 962 -1614
rect 72 -1617 444 -1616
rect 457 -1617 780 -1616
rect 786 -1617 836 -1616
rect 947 -1617 962 -1616
rect 75 -1619 241 -1618
rect 289 -1619 374 -1618
rect 460 -1619 542 -1618
rect 555 -1619 1004 -1618
rect 79 -1621 633 -1620
rect 688 -1621 703 -1620
rect 716 -1621 899 -1620
rect 996 -1621 1004 -1620
rect 58 -1623 633 -1622
rect 674 -1623 717 -1622
rect 723 -1623 766 -1622
rect 772 -1623 850 -1622
rect 877 -1623 948 -1622
rect 82 -1625 598 -1624
rect 611 -1625 640 -1624
rect 695 -1625 759 -1624
rect 765 -1625 857 -1624
rect 877 -1625 976 -1624
rect 86 -1627 244 -1626
rect 289 -1627 311 -1626
rect 317 -1627 538 -1626
rect 562 -1627 577 -1626
rect 590 -1627 619 -1626
rect 639 -1627 955 -1626
rect 975 -1627 1039 -1626
rect 107 -1629 339 -1628
rect 467 -1629 1053 -1628
rect 121 -1631 195 -1630
rect 205 -1631 262 -1630
rect 268 -1631 339 -1630
rect 471 -1631 696 -1630
rect 702 -1631 745 -1630
rect 751 -1631 955 -1630
rect 1052 -1631 1074 -1630
rect 9 -1633 206 -1632
rect 212 -1633 255 -1632
rect 303 -1633 409 -1632
rect 474 -1633 1109 -1632
rect 9 -1635 136 -1634
rect 138 -1635 269 -1634
rect 310 -1635 388 -1634
rect 408 -1635 647 -1634
rect 730 -1635 1018 -1634
rect 128 -1637 185 -1636
rect 212 -1637 843 -1636
rect 856 -1637 927 -1636
rect 142 -1639 402 -1638
rect 474 -1639 738 -1638
rect 744 -1639 815 -1638
rect 835 -1639 934 -1638
rect 65 -1641 402 -1640
rect 481 -1641 906 -1640
rect 926 -1641 1060 -1640
rect 65 -1643 125 -1642
rect 142 -1643 178 -1642
rect 222 -1643 297 -1642
rect 317 -1643 437 -1642
rect 492 -1643 829 -1642
rect 842 -1643 941 -1642
rect 149 -1645 185 -1644
rect 194 -1645 437 -1644
rect 499 -1645 528 -1644
rect 537 -1645 1088 -1644
rect 44 -1647 150 -1646
rect 156 -1647 444 -1646
rect 478 -1647 500 -1646
rect 513 -1647 1102 -1646
rect 170 -1649 535 -1648
rect 544 -1649 619 -1648
rect 684 -1649 941 -1648
rect 170 -1651 199 -1650
rect 222 -1651 276 -1650
rect 296 -1651 507 -1650
rect 513 -1651 888 -1650
rect 905 -1651 1011 -1650
rect 86 -1653 199 -1652
rect 226 -1653 871 -1652
rect 933 -1653 1025 -1652
rect 16 -1655 227 -1654
rect 233 -1655 283 -1654
rect 366 -1655 507 -1654
rect 520 -1655 675 -1654
rect 772 -1655 895 -1654
rect 16 -1657 52 -1656
rect 163 -1657 367 -1656
rect 387 -1657 451 -1656
rect 565 -1657 1067 -1656
rect 51 -1659 570 -1658
rect 597 -1659 626 -1658
rect 779 -1659 885 -1658
rect 177 -1661 423 -1660
rect 558 -1661 570 -1660
rect 604 -1661 752 -1660
rect 793 -1661 864 -1660
rect 100 -1663 423 -1662
rect 464 -1663 605 -1662
rect 625 -1663 654 -1662
rect 814 -1663 913 -1662
rect 100 -1665 248 -1664
rect 275 -1665 808 -1664
rect 821 -1665 871 -1664
rect 93 -1667 248 -1666
rect 345 -1667 521 -1666
rect 653 -1667 668 -1666
rect 733 -1667 808 -1666
rect 863 -1667 990 -1666
rect 345 -1669 458 -1668
rect 478 -1669 822 -1668
rect 394 -1671 647 -1670
rect 331 -1673 395 -1672
rect 488 -1673 668 -1672
rect 331 -1675 465 -1674
rect 2 -1686 377 -1685
rect 443 -1686 563 -1685
rect 593 -1686 1018 -1685
rect 1027 -1686 1053 -1685
rect 2 -1688 97 -1687
rect 110 -1688 129 -1687
rect 152 -1688 276 -1687
rect 282 -1688 395 -1687
rect 429 -1688 563 -1687
rect 621 -1688 717 -1687
rect 730 -1688 871 -1687
rect 887 -1688 962 -1687
rect 1003 -1688 1011 -1687
rect 9 -1690 192 -1689
rect 198 -1690 598 -1689
rect 649 -1690 857 -1689
rect 891 -1690 983 -1689
rect 16 -1692 216 -1691
rect 233 -1692 437 -1691
rect 443 -1692 678 -1691
rect 716 -1692 724 -1691
rect 730 -1692 759 -1691
rect 779 -1692 783 -1691
rect 803 -1692 808 -1691
rect 821 -1692 969 -1691
rect 23 -1694 195 -1693
rect 198 -1694 255 -1693
rect 275 -1694 734 -1693
rect 779 -1694 815 -1693
rect 835 -1694 871 -1693
rect 912 -1694 976 -1693
rect 23 -1696 223 -1695
rect 240 -1696 412 -1695
rect 415 -1696 437 -1695
rect 457 -1696 857 -1695
rect 898 -1696 976 -1695
rect 30 -1698 468 -1697
rect 471 -1698 752 -1697
rect 793 -1698 815 -1697
rect 835 -1698 941 -1697
rect 30 -1700 346 -1699
rect 348 -1700 388 -1699
rect 394 -1700 507 -1699
rect 548 -1700 808 -1699
rect 898 -1700 920 -1699
rect 926 -1700 962 -1699
rect 37 -1702 181 -1701
rect 184 -1702 192 -1701
rect 222 -1702 262 -1701
rect 285 -1702 409 -1701
rect 467 -1702 738 -1701
rect 793 -1702 829 -1701
rect 863 -1702 920 -1701
rect 940 -1702 1007 -1701
rect 37 -1704 293 -1703
rect 299 -1704 552 -1703
rect 555 -1704 619 -1703
rect 639 -1704 892 -1703
rect 44 -1706 62 -1705
rect 65 -1706 167 -1705
rect 170 -1706 297 -1705
rect 317 -1706 426 -1705
rect 464 -1706 640 -1705
rect 688 -1706 752 -1705
rect 782 -1706 829 -1705
rect 16 -1708 465 -1707
rect 471 -1708 566 -1707
rect 569 -1708 689 -1707
rect 723 -1708 745 -1707
rect 44 -1710 405 -1709
rect 408 -1710 710 -1709
rect 51 -1712 384 -1711
rect 478 -1712 535 -1711
rect 548 -1712 577 -1711
rect 597 -1712 633 -1711
rect 51 -1714 94 -1713
rect 128 -1714 482 -1713
rect 485 -1714 990 -1713
rect 54 -1716 255 -1715
rect 261 -1716 325 -1715
rect 338 -1716 346 -1715
rect 352 -1716 381 -1715
rect 481 -1716 612 -1715
rect 614 -1716 710 -1715
rect 65 -1718 230 -1717
rect 243 -1718 269 -1717
rect 289 -1718 514 -1717
rect 516 -1718 738 -1717
rect 72 -1720 451 -1719
rect 488 -1720 528 -1719
rect 576 -1720 591 -1719
rect 618 -1720 759 -1719
rect 72 -1722 164 -1721
rect 177 -1722 430 -1721
rect 450 -1722 661 -1721
rect 79 -1724 122 -1723
rect 135 -1724 479 -1723
rect 492 -1724 955 -1723
rect 86 -1726 745 -1725
rect 947 -1726 955 -1725
rect 86 -1728 104 -1727
rect 121 -1728 143 -1727
rect 149 -1728 384 -1727
rect 401 -1728 528 -1727
rect 541 -1728 661 -1727
rect 905 -1728 948 -1727
rect 138 -1730 927 -1729
rect 142 -1732 304 -1731
rect 317 -1732 475 -1731
rect 492 -1732 895 -1731
rect 149 -1734 241 -1733
rect 247 -1734 559 -1733
rect 156 -1736 202 -1735
rect 268 -1736 325 -1735
rect 331 -1736 339 -1735
rect 352 -1736 454 -1735
rect 495 -1736 675 -1735
rect 156 -1738 227 -1737
rect 289 -1738 360 -1737
rect 366 -1738 654 -1737
rect 674 -1738 878 -1737
rect 100 -1740 360 -1739
rect 366 -1740 983 -1739
rect 100 -1742 171 -1741
rect 177 -1742 248 -1741
rect 303 -1742 311 -1741
rect 369 -1742 521 -1741
rect 541 -1742 906 -1741
rect 114 -1744 521 -1743
rect 842 -1744 878 -1743
rect 107 -1746 115 -1745
rect 163 -1746 314 -1745
rect 331 -1746 370 -1745
rect 373 -1746 416 -1745
rect 485 -1746 654 -1745
rect 786 -1746 843 -1745
rect 107 -1748 822 -1747
rect 187 -1750 864 -1749
rect 226 -1752 626 -1751
rect 786 -1752 934 -1751
rect 401 -1754 458 -1753
rect 499 -1754 507 -1753
rect 513 -1754 584 -1753
rect 625 -1754 668 -1753
rect 884 -1754 934 -1753
rect 373 -1756 500 -1755
rect 583 -1756 703 -1755
rect 800 -1756 885 -1755
rect 604 -1758 703 -1757
rect 604 -1760 647 -1759
rect 667 -1760 682 -1759
rect 569 -1762 647 -1761
rect 681 -1762 696 -1761
rect 695 -1764 766 -1763
rect 765 -1766 773 -1765
rect 422 -1768 773 -1767
rect 422 -1770 913 -1769
rect 2 -1781 188 -1780
rect 205 -1781 524 -1780
rect 565 -1781 948 -1780
rect 975 -1781 1000 -1780
rect 9 -1783 31 -1782
rect 37 -1783 311 -1782
rect 313 -1783 500 -1782
rect 506 -1783 517 -1782
rect 590 -1783 962 -1782
rect 996 -1783 1011 -1782
rect 23 -1785 213 -1784
rect 215 -1785 297 -1784
rect 310 -1785 458 -1784
rect 460 -1785 920 -1784
rect 947 -1785 1025 -1784
rect 44 -1787 367 -1786
rect 369 -1787 395 -1786
rect 422 -1787 703 -1786
rect 726 -1787 955 -1786
rect 51 -1789 892 -1788
rect 915 -1789 934 -1788
rect 51 -1791 349 -1790
rect 369 -1791 388 -1790
rect 450 -1791 542 -1790
rect 590 -1791 605 -1790
rect 611 -1791 857 -1790
rect 54 -1793 73 -1792
rect 79 -1793 104 -1792
rect 107 -1793 192 -1792
rect 215 -1793 657 -1792
rect 674 -1793 815 -1792
rect 842 -1793 853 -1792
rect 58 -1795 122 -1794
rect 128 -1795 150 -1794
rect 177 -1795 230 -1794
rect 240 -1795 528 -1794
rect 541 -1795 629 -1794
rect 632 -1795 927 -1794
rect 65 -1797 328 -1796
rect 380 -1797 640 -1796
rect 642 -1797 990 -1796
rect 65 -1799 143 -1798
rect 149 -1799 157 -1798
rect 170 -1799 178 -1798
rect 226 -1799 402 -1798
rect 415 -1799 451 -1798
rect 464 -1799 549 -1798
rect 604 -1799 745 -1798
rect 814 -1799 899 -1798
rect 72 -1801 416 -1800
rect 464 -1801 563 -1800
rect 611 -1801 766 -1800
rect 898 -1801 951 -1800
rect 79 -1803 594 -1802
rect 618 -1803 752 -1802
rect 93 -1805 129 -1804
rect 135 -1805 185 -1804
rect 226 -1805 552 -1804
rect 618 -1805 724 -1804
rect 751 -1805 850 -1804
rect 93 -1807 115 -1806
rect 121 -1807 426 -1806
rect 467 -1807 514 -1806
rect 527 -1807 983 -1806
rect 100 -1809 402 -1808
rect 478 -1809 535 -1808
rect 548 -1809 766 -1808
rect 100 -1811 199 -1810
rect 243 -1811 388 -1810
rect 499 -1811 626 -1810
rect 635 -1811 829 -1810
rect 110 -1813 493 -1812
rect 506 -1813 773 -1812
rect 828 -1813 836 -1812
rect 86 -1815 493 -1814
rect 534 -1815 556 -1814
rect 576 -1815 836 -1814
rect 86 -1817 202 -1816
rect 254 -1817 563 -1816
rect 576 -1817 598 -1816
rect 621 -1817 745 -1816
rect 114 -1819 444 -1818
rect 555 -1819 668 -1818
rect 674 -1819 717 -1818
rect 135 -1821 164 -1820
rect 170 -1821 458 -1820
rect 646 -1821 857 -1820
rect 142 -1823 304 -1822
rect 380 -1823 521 -1822
rect 653 -1823 871 -1822
rect 156 -1825 220 -1824
rect 247 -1825 304 -1824
rect 418 -1825 647 -1824
rect 653 -1825 731 -1824
rect 194 -1827 220 -1826
rect 247 -1827 276 -1826
rect 282 -1827 395 -1826
rect 443 -1827 689 -1826
rect 702 -1827 1018 -1826
rect 254 -1829 325 -1828
rect 520 -1829 878 -1828
rect 268 -1831 374 -1830
rect 660 -1831 773 -1830
rect 786 -1831 878 -1830
rect 261 -1833 269 -1832
rect 275 -1833 678 -1832
rect 681 -1833 801 -1832
rect 233 -1835 262 -1834
rect 282 -1835 339 -1834
rect 373 -1835 409 -1834
rect 597 -1835 661 -1834
rect 667 -1835 941 -1834
rect 233 -1837 353 -1836
rect 408 -1837 850 -1836
rect 289 -1839 353 -1838
rect 681 -1839 696 -1838
rect 709 -1839 871 -1838
rect 289 -1841 332 -1840
rect 338 -1841 486 -1840
rect 688 -1841 780 -1840
rect 786 -1841 864 -1840
rect 296 -1843 377 -1842
rect 695 -1843 794 -1842
rect 838 -1843 864 -1842
rect 317 -1845 486 -1844
rect 709 -1845 759 -1844
rect 793 -1845 843 -1844
rect 317 -1847 346 -1846
rect 716 -1847 808 -1846
rect 324 -1849 437 -1848
rect 730 -1849 822 -1848
rect 331 -1851 570 -1850
rect 737 -1851 780 -1850
rect 807 -1851 969 -1850
rect 345 -1853 1004 -1852
rect 429 -1855 437 -1854
rect 569 -1855 885 -1854
rect 429 -1857 472 -1856
rect 737 -1857 913 -1856
rect 359 -1859 472 -1858
rect 758 -1859 846 -1858
rect 821 -1861 906 -1860
rect 16 -1872 52 -1871
rect 58 -1872 164 -1871
rect 184 -1872 199 -1871
rect 219 -1872 262 -1871
rect 285 -1872 871 -1871
rect 23 -1874 185 -1873
rect 194 -1874 199 -1873
rect 229 -1874 241 -1873
rect 243 -1874 318 -1873
rect 324 -1874 412 -1873
rect 415 -1874 451 -1873
rect 464 -1874 468 -1873
rect 509 -1874 738 -1873
rect 782 -1874 878 -1873
rect 51 -1876 192 -1875
rect 247 -1876 325 -1875
rect 334 -1876 710 -1875
rect 845 -1876 899 -1875
rect 58 -1878 297 -1877
rect 348 -1878 353 -1877
rect 359 -1878 440 -1877
rect 443 -1878 640 -1877
rect 702 -1878 822 -1877
rect 65 -1880 160 -1879
rect 177 -1880 244 -1879
rect 247 -1880 388 -1879
rect 411 -1880 461 -1879
rect 464 -1880 479 -1879
rect 520 -1880 584 -1879
rect 618 -1880 664 -1879
rect 702 -1880 759 -1879
rect 821 -1880 864 -1879
rect 65 -1882 125 -1881
rect 128 -1882 150 -1881
rect 177 -1882 458 -1881
rect 471 -1882 738 -1881
rect 758 -1882 794 -1881
rect 72 -1884 241 -1883
rect 296 -1884 402 -1883
rect 418 -1884 619 -1883
rect 628 -1884 675 -1883
rect 709 -1884 762 -1883
rect 793 -1884 857 -1883
rect 72 -1886 146 -1885
rect 191 -1886 276 -1885
rect 338 -1886 353 -1885
rect 362 -1886 486 -1885
rect 527 -1886 815 -1885
rect 79 -1888 230 -1887
rect 289 -1888 339 -1887
rect 366 -1888 524 -1887
rect 530 -1888 598 -1887
rect 632 -1888 787 -1887
rect 814 -1888 829 -1887
rect 79 -1890 283 -1889
rect 289 -1890 318 -1889
rect 373 -1890 633 -1889
rect 674 -1890 717 -1889
rect 751 -1890 787 -1889
rect 44 -1892 283 -1891
rect 310 -1892 374 -1891
rect 387 -1892 451 -1891
rect 471 -1892 773 -1891
rect 100 -1894 262 -1893
rect 394 -1894 402 -1893
rect 408 -1894 598 -1893
rect 646 -1894 717 -1893
rect 751 -1894 780 -1893
rect 100 -1896 115 -1895
rect 121 -1896 164 -1895
rect 215 -1896 419 -1895
rect 422 -1896 643 -1895
rect 646 -1896 689 -1895
rect 86 -1898 122 -1897
rect 142 -1898 276 -1897
rect 408 -1898 668 -1897
rect 681 -1898 689 -1897
rect 86 -1900 234 -1899
rect 380 -1900 668 -1899
rect 681 -1900 773 -1899
rect 93 -1902 143 -1901
rect 212 -1902 381 -1901
rect 422 -1902 724 -1901
rect 93 -1904 332 -1903
rect 429 -1904 444 -1903
rect 478 -1904 493 -1903
rect 548 -1904 727 -1903
rect 107 -1906 206 -1905
rect 212 -1906 269 -1905
rect 310 -1906 332 -1905
rect 429 -1906 514 -1905
rect 548 -1906 605 -1905
rect 625 -1906 724 -1905
rect 107 -1908 136 -1907
rect 166 -1908 206 -1907
rect 268 -1908 304 -1907
rect 457 -1908 514 -1907
rect 551 -1908 801 -1907
rect 114 -1910 157 -1909
rect 254 -1910 304 -1909
rect 485 -1910 507 -1909
rect 583 -1910 661 -1909
rect 135 -1912 171 -1911
rect 254 -1912 570 -1911
rect 604 -1912 808 -1911
rect 131 -1914 171 -1913
rect 492 -1914 500 -1913
rect 506 -1914 542 -1913
rect 562 -1914 661 -1913
rect 149 -1916 157 -1915
rect 394 -1916 563 -1915
rect 625 -1916 696 -1915
rect 499 -1918 577 -1917
rect 653 -1918 696 -1917
rect 467 -1920 577 -1919
rect 611 -1920 654 -1919
rect 453 -1922 612 -1921
rect 534 -1924 570 -1923
rect 534 -1926 591 -1925
rect 541 -1928 556 -1927
rect 555 -1930 731 -1929
rect 730 -1932 818 -1931
rect 33 -1943 38 -1942
rect 40 -1943 48 -1942
rect 51 -1943 395 -1942
rect 418 -1943 668 -1942
rect 677 -1943 689 -1942
rect 695 -1943 801 -1942
rect 37 -1945 115 -1944
rect 121 -1945 178 -1944
rect 191 -1945 549 -1944
rect 576 -1945 731 -1944
rect 782 -1945 822 -1944
rect 44 -1947 136 -1946
rect 138 -1947 265 -1946
rect 275 -1947 332 -1946
rect 373 -1947 412 -1946
rect 446 -1947 493 -1946
rect 495 -1947 542 -1946
rect 593 -1947 626 -1946
rect 653 -1947 759 -1946
rect 786 -1947 808 -1946
rect 58 -1949 237 -1948
rect 243 -1949 388 -1948
rect 394 -1949 780 -1948
rect 72 -1951 76 -1950
rect 93 -1951 433 -1950
rect 439 -1951 626 -1950
rect 653 -1951 675 -1950
rect 684 -1951 752 -1950
rect 772 -1951 780 -1950
rect 72 -1953 108 -1952
rect 114 -1953 143 -1952
rect 170 -1953 178 -1952
rect 219 -1953 290 -1952
rect 296 -1953 605 -1952
rect 611 -1953 752 -1952
rect 75 -1955 108 -1954
rect 128 -1955 185 -1954
rect 229 -1955 262 -1954
rect 275 -1955 335 -1954
rect 352 -1955 388 -1954
rect 439 -1955 465 -1954
rect 499 -1955 696 -1954
rect 709 -1955 787 -1954
rect 51 -1957 230 -1956
rect 233 -1957 269 -1956
rect 296 -1957 475 -1956
rect 478 -1957 500 -1956
rect 506 -1957 549 -1956
rect 583 -1957 612 -1956
rect 618 -1957 759 -1956
rect 58 -1959 129 -1958
rect 142 -1959 195 -1958
rect 205 -1959 262 -1958
rect 317 -1959 465 -1958
rect 506 -1959 514 -1958
rect 516 -1959 773 -1958
rect 86 -1961 220 -1960
rect 254 -1961 332 -1960
rect 352 -1961 409 -1960
rect 415 -1961 710 -1960
rect 86 -1963 283 -1962
rect 317 -1963 346 -1962
rect 359 -1963 374 -1962
rect 408 -1963 423 -1962
rect 450 -1963 556 -1962
rect 579 -1963 619 -1962
rect 660 -1963 668 -1962
rect 688 -1963 766 -1962
rect 93 -1965 181 -1964
rect 184 -1965 311 -1964
rect 320 -1965 402 -1964
rect 415 -1965 461 -1964
rect 527 -1965 542 -1964
rect 555 -1965 563 -1964
rect 593 -1965 731 -1964
rect 744 -1965 766 -1964
rect 100 -1967 157 -1966
rect 163 -1967 171 -1966
rect 205 -1967 227 -1966
rect 247 -1967 255 -1966
rect 271 -1967 451 -1966
rect 453 -1967 738 -1966
rect 100 -1969 136 -1968
rect 149 -1969 269 -1968
rect 282 -1969 493 -1968
rect 527 -1969 727 -1968
rect 149 -1971 223 -1970
rect 303 -1971 360 -1970
rect 366 -1971 479 -1970
rect 534 -1971 591 -1970
rect 597 -1971 605 -1970
rect 723 -1971 738 -1970
rect 159 -1973 304 -1972
rect 324 -1973 346 -1972
rect 369 -1973 535 -1972
rect 562 -1973 640 -1972
rect 723 -1973 794 -1972
rect 79 -1975 325 -1974
rect 401 -1975 486 -1974
rect 576 -1975 745 -1974
rect 65 -1977 80 -1976
rect 159 -1977 164 -1976
rect 198 -1977 248 -1976
rect 422 -1977 503 -1976
rect 597 -1977 647 -1976
rect 16 -1979 66 -1978
rect 191 -1979 199 -1978
rect 212 -1979 234 -1978
rect 443 -1979 486 -1978
rect 632 -1979 640 -1978
rect 646 -1979 675 -1978
rect 212 -1981 241 -1980
rect 457 -1981 521 -1980
rect 569 -1981 633 -1980
rect 338 -1983 458 -1982
rect 520 -1983 682 -1982
rect 338 -1985 381 -1984
rect 429 -1985 570 -1984
rect 681 -1985 703 -1984
rect 380 -1987 472 -1986
rect 702 -1987 717 -1986
rect 436 -1989 717 -1988
rect 23 -1991 437 -1990
rect 16 -2002 94 -2001
rect 156 -2002 188 -2001
rect 201 -2002 227 -2001
rect 229 -2002 339 -2001
rect 387 -2002 405 -2001
rect 432 -2002 570 -2001
rect 586 -2002 640 -2001
rect 646 -2002 664 -2001
rect 670 -2002 787 -2001
rect 796 -2002 815 -2001
rect 30 -2004 80 -2003
rect 177 -2004 311 -2003
rect 313 -2004 325 -2003
rect 331 -2004 398 -2003
rect 488 -2004 514 -2003
rect 548 -2004 780 -2003
rect 37 -2006 150 -2005
rect 229 -2006 269 -2005
rect 271 -2006 360 -2005
rect 387 -2006 493 -2005
rect 513 -2006 633 -2005
rect 639 -2006 696 -2005
rect 744 -2006 808 -2005
rect 37 -2008 185 -2007
rect 233 -2008 241 -2007
rect 247 -2008 381 -2007
rect 492 -2008 556 -2007
rect 569 -2008 794 -2007
rect 44 -2010 199 -2009
rect 236 -2010 549 -2009
rect 555 -2010 619 -2009
rect 660 -2010 703 -2009
rect 744 -2010 752 -2009
rect 758 -2010 787 -2009
rect 44 -2012 108 -2011
rect 149 -2012 171 -2011
rect 191 -2012 199 -2011
rect 247 -2012 255 -2011
rect 264 -2012 633 -2011
rect 653 -2012 661 -2011
rect 674 -2012 696 -2011
rect 751 -2012 773 -2011
rect 51 -2014 167 -2013
rect 170 -2014 258 -2013
rect 289 -2014 353 -2013
rect 359 -2014 374 -2013
rect 380 -2014 409 -2013
rect 464 -2014 675 -2013
rect 688 -2014 731 -2013
rect 758 -2014 766 -2013
rect 51 -2016 591 -2015
rect 593 -2016 801 -2015
rect 58 -2018 244 -2017
rect 289 -2018 349 -2017
rect 352 -2018 423 -2017
rect 464 -2018 479 -2017
rect 562 -2018 619 -2017
rect 691 -2018 738 -2017
rect 58 -2020 115 -2019
rect 191 -2020 213 -2019
rect 243 -2020 283 -2019
rect 292 -2020 433 -2019
rect 471 -2020 703 -2019
rect 716 -2020 731 -2019
rect 65 -2022 234 -2021
rect 296 -2022 367 -2021
rect 373 -2022 451 -2021
rect 565 -2022 738 -2021
rect 65 -2024 461 -2023
rect 583 -2024 654 -2023
rect 709 -2024 717 -2023
rect 72 -2026 136 -2025
rect 163 -2026 297 -2025
rect 303 -2026 437 -2025
rect 450 -2026 598 -2025
rect 681 -2026 710 -2025
rect 72 -2028 101 -2027
rect 107 -2028 255 -2027
rect 303 -2028 475 -2027
rect 541 -2028 598 -2027
rect 667 -2028 682 -2027
rect 79 -2030 318 -2029
rect 324 -2030 395 -2029
rect 401 -2030 766 -2029
rect 86 -2032 136 -2031
rect 219 -2032 283 -2031
rect 317 -2032 458 -2031
rect 527 -2032 542 -2031
rect 583 -2032 612 -2031
rect 646 -2032 668 -2031
rect 86 -2034 521 -2033
rect 590 -2034 727 -2033
rect 100 -2036 122 -2035
rect 128 -2036 213 -2035
rect 261 -2036 528 -2035
rect 611 -2036 678 -2035
rect 23 -2038 129 -2037
rect 205 -2038 220 -2037
rect 261 -2038 346 -2037
rect 394 -2038 773 -2037
rect 114 -2040 143 -2039
rect 205 -2040 447 -2039
rect 457 -2040 605 -2039
rect 93 -2042 143 -2041
rect 331 -2042 402 -2041
rect 408 -2042 416 -2041
rect 418 -2042 605 -2041
rect 121 -2044 185 -2043
rect 338 -2044 601 -2043
rect 345 -2046 444 -2045
rect 506 -2046 521 -2045
rect 415 -2048 535 -2047
rect 422 -2050 500 -2049
rect 429 -2052 444 -2051
rect 478 -2052 500 -2051
rect 485 -2054 535 -2053
rect 23 -2065 398 -2064
rect 411 -2065 514 -2064
rect 534 -2065 538 -2064
rect 541 -2065 594 -2064
rect 653 -2065 738 -2064
rect 23 -2067 241 -2066
rect 254 -2067 283 -2066
rect 292 -2067 367 -2066
rect 373 -2067 402 -2066
rect 418 -2067 500 -2066
rect 534 -2067 556 -2066
rect 569 -2067 633 -2066
rect 667 -2067 682 -2066
rect 723 -2067 759 -2066
rect 30 -2069 146 -2068
rect 184 -2069 237 -2068
rect 240 -2069 276 -2068
rect 345 -2069 423 -2068
rect 436 -2069 514 -2068
rect 537 -2069 556 -2068
rect 569 -2069 584 -2068
rect 632 -2069 647 -2068
rect 670 -2069 787 -2068
rect 30 -2071 472 -2070
rect 474 -2071 619 -2070
rect 646 -2071 731 -2070
rect 37 -2073 230 -2072
rect 257 -2073 430 -2072
rect 457 -2073 780 -2072
rect 44 -2075 178 -2074
rect 212 -2075 283 -2074
rect 296 -2075 423 -2074
rect 457 -2075 584 -2074
rect 618 -2075 661 -2074
rect 681 -2075 773 -2074
rect 44 -2077 171 -2076
rect 212 -2077 349 -2076
rect 352 -2077 563 -2076
rect 660 -2077 675 -2076
rect 709 -2077 724 -2076
rect 726 -2077 738 -2076
rect 51 -2079 125 -2078
rect 135 -2079 178 -2078
rect 219 -2079 255 -2078
rect 275 -2079 311 -2078
rect 324 -2079 353 -2078
rect 373 -2079 486 -2078
rect 488 -2079 493 -2078
rect 499 -2079 591 -2078
rect 709 -2079 752 -2078
rect 51 -2081 150 -2080
rect 268 -2081 311 -2080
rect 317 -2081 325 -2080
rect 359 -2081 486 -2080
rect 492 -2081 549 -2080
rect 562 -2081 598 -2080
rect 58 -2083 132 -2082
rect 135 -2083 339 -2082
rect 380 -2083 416 -2082
rect 464 -2083 510 -2082
rect 527 -2083 675 -2082
rect 58 -2085 129 -2084
rect 142 -2085 363 -2084
rect 366 -2085 465 -2084
rect 474 -2085 577 -2084
rect 65 -2087 139 -2086
rect 142 -2087 157 -2086
rect 233 -2087 269 -2086
rect 296 -2087 332 -2086
rect 338 -2087 461 -2086
rect 478 -2087 703 -2086
rect 65 -2089 244 -2088
rect 317 -2089 598 -2088
rect 688 -2089 703 -2088
rect 72 -2091 104 -2090
rect 107 -2091 185 -2090
rect 233 -2091 290 -2090
rect 331 -2091 388 -2090
rect 415 -2091 451 -2090
rect 460 -2091 766 -2090
rect 72 -2093 262 -2092
rect 320 -2093 451 -2092
rect 478 -2093 517 -2092
rect 520 -2093 528 -2092
rect 576 -2093 626 -2092
rect 688 -2093 717 -2092
rect 79 -2095 440 -2094
rect 506 -2095 549 -2094
rect 625 -2095 640 -2094
rect 716 -2095 745 -2094
rect 79 -2097 174 -2096
rect 247 -2097 290 -2096
rect 387 -2097 507 -2096
rect 520 -2097 605 -2096
rect 86 -2099 188 -2098
rect 261 -2099 433 -2098
rect 604 -2099 696 -2098
rect 86 -2101 97 -2100
rect 100 -2101 108 -2100
rect 121 -2101 304 -2100
rect 394 -2101 640 -2100
rect 93 -2103 230 -2102
rect 303 -2103 384 -2102
rect 394 -2103 409 -2102
rect 16 -2105 94 -2104
rect 128 -2105 542 -2104
rect 149 -2107 192 -2106
rect 163 -2109 248 -2108
rect 156 -2111 164 -2110
rect 180 -2111 696 -2110
rect 180 -2113 199 -2112
rect 191 -2115 206 -2114
rect 16 -2117 206 -2116
rect 198 -2119 220 -2118
rect 16 -2130 475 -2129
rect 506 -2130 626 -2129
rect 688 -2130 699 -2129
rect 40 -2132 153 -2131
rect 163 -2132 174 -2131
rect 184 -2132 255 -2131
rect 261 -2132 454 -2131
rect 457 -2132 689 -2131
rect 695 -2132 731 -2131
rect 44 -2134 230 -2133
rect 254 -2134 339 -2133
rect 345 -2134 598 -2133
rect 625 -2134 710 -2133
rect 51 -2136 220 -2135
rect 226 -2136 241 -2135
rect 261 -2136 353 -2135
rect 359 -2136 430 -2135
rect 436 -2136 468 -2135
rect 509 -2136 542 -2135
rect 558 -2136 717 -2135
rect 58 -2138 101 -2137
rect 121 -2138 248 -2137
rect 268 -2138 346 -2137
rect 348 -2138 412 -2137
rect 439 -2138 612 -2137
rect 660 -2138 717 -2137
rect 65 -2140 321 -2139
rect 324 -2140 353 -2139
rect 380 -2140 395 -2139
rect 408 -2140 514 -2139
rect 534 -2140 710 -2139
rect 72 -2142 335 -2141
rect 362 -2142 381 -2141
rect 390 -2142 493 -2141
rect 513 -2142 521 -2141
rect 541 -2142 549 -2141
rect 579 -2142 703 -2141
rect 100 -2144 115 -2143
rect 128 -2144 157 -2143
rect 170 -2144 416 -2143
rect 464 -2144 563 -2143
rect 583 -2144 591 -2143
rect 593 -2144 696 -2143
rect 30 -2146 129 -2145
rect 135 -2146 164 -2145
rect 198 -2146 451 -2145
rect 464 -2146 500 -2145
rect 520 -2146 528 -2145
rect 548 -2146 570 -2145
rect 597 -2146 605 -2145
rect 611 -2146 654 -2145
rect 107 -2148 136 -2147
rect 142 -2148 160 -2147
rect 198 -2148 223 -2147
rect 226 -2148 269 -2147
rect 282 -2148 290 -2147
rect 296 -2148 339 -2147
rect 373 -2148 395 -2147
rect 408 -2148 535 -2147
rect 555 -2148 703 -2147
rect 23 -2150 160 -2149
rect 170 -2150 556 -2149
rect 604 -2150 619 -2149
rect 639 -2150 661 -2149
rect 107 -2152 178 -2151
rect 201 -2152 276 -2151
rect 282 -2152 325 -2151
rect 331 -2152 430 -2151
rect 471 -2152 563 -2151
rect 639 -2152 682 -2151
rect 114 -2154 286 -2153
rect 296 -2154 388 -2153
rect 443 -2154 472 -2153
rect 485 -2154 619 -2153
rect 646 -2154 654 -2153
rect 121 -2156 388 -2155
rect 443 -2156 479 -2155
rect 499 -2156 510 -2155
rect 646 -2156 675 -2155
rect 142 -2158 234 -2157
rect 275 -2158 304 -2157
rect 313 -2158 738 -2157
rect 149 -2160 206 -2159
rect 212 -2160 234 -2159
rect 303 -2160 311 -2159
rect 331 -2160 528 -2159
rect 667 -2160 675 -2159
rect 79 -2162 213 -2161
rect 219 -2162 416 -2161
rect 478 -2162 570 -2161
rect 667 -2162 724 -2161
rect 156 -2164 311 -2163
rect 366 -2164 486 -2163
rect 576 -2164 724 -2163
rect 177 -2166 181 -2165
rect 191 -2166 206 -2165
rect 222 -2166 318 -2165
rect 366 -2166 423 -2165
rect 191 -2168 209 -2167
rect 373 -2168 402 -2167
rect 422 -2168 577 -2167
rect 250 -2170 402 -2169
rect 86 -2181 90 -2180
rect 114 -2181 307 -2180
rect 380 -2181 493 -2180
rect 506 -2181 528 -2180
rect 534 -2181 671 -2180
rect 674 -2181 682 -2180
rect 114 -2183 185 -2182
rect 205 -2183 220 -2182
rect 222 -2183 577 -2182
rect 579 -2183 724 -2182
rect 121 -2185 150 -2184
rect 163 -2185 185 -2184
rect 205 -2185 300 -2184
rect 324 -2185 381 -2184
rect 401 -2185 461 -2184
rect 492 -2185 559 -2184
rect 569 -2185 717 -2184
rect 124 -2187 255 -2186
rect 282 -2187 367 -2186
rect 401 -2187 423 -2186
rect 425 -2187 563 -2186
rect 583 -2187 689 -2186
rect 128 -2189 412 -2188
rect 429 -2189 619 -2188
rect 639 -2189 668 -2188
rect 142 -2191 220 -2190
rect 240 -2191 514 -2190
rect 555 -2191 612 -2190
rect 170 -2193 241 -2192
rect 243 -2193 255 -2192
rect 285 -2193 391 -2192
rect 394 -2193 563 -2192
rect 569 -2193 619 -2192
rect 142 -2195 171 -2194
rect 198 -2195 395 -2194
rect 408 -2195 444 -2194
rect 450 -2195 465 -2194
rect 499 -2195 528 -2194
rect 555 -2195 633 -2194
rect 212 -2197 346 -2196
rect 366 -2197 374 -2196
rect 387 -2197 465 -2196
rect 513 -2197 549 -2196
rect 583 -2197 654 -2196
rect 152 -2199 213 -2198
rect 285 -2199 451 -2198
rect 548 -2199 591 -2198
rect 597 -2199 640 -2198
rect 296 -2201 615 -2200
rect 632 -2201 703 -2200
rect 317 -2203 346 -2202
rect 415 -2203 500 -2202
rect 586 -2203 605 -2202
rect 317 -2205 472 -2204
rect 509 -2205 605 -2204
rect 324 -2207 353 -2206
rect 359 -2207 416 -2206
rect 429 -2207 479 -2206
rect 590 -2207 626 -2206
rect 268 -2209 353 -2208
rect 432 -2209 458 -2208
rect 478 -2209 622 -2208
rect 268 -2211 311 -2210
rect 331 -2211 472 -2210
rect 485 -2211 626 -2210
rect 261 -2213 332 -2212
rect 436 -2213 535 -2212
rect 597 -2213 647 -2212
rect 261 -2215 339 -2214
rect 390 -2215 437 -2214
rect 485 -2215 521 -2214
rect 156 -2217 339 -2216
rect 520 -2217 542 -2216
rect 156 -2219 178 -2218
rect 289 -2219 311 -2218
rect 541 -2219 661 -2218
rect 131 -2221 178 -2220
rect 247 -2221 290 -2220
rect 660 -2221 710 -2220
rect 100 -2223 132 -2222
rect 247 -2223 304 -2222
rect 107 -2234 230 -2233
rect 275 -2234 283 -2233
rect 306 -2234 479 -2233
rect 534 -2234 612 -2233
rect 114 -2236 195 -2235
rect 198 -2236 237 -2235
rect 254 -2236 276 -2235
rect 313 -2236 402 -2235
rect 415 -2236 426 -2235
rect 443 -2236 479 -2235
rect 527 -2236 535 -2235
rect 562 -2236 591 -2235
rect 607 -2236 661 -2235
rect 114 -2238 143 -2237
rect 149 -2238 171 -2237
rect 173 -2238 192 -2237
rect 201 -2238 213 -2237
rect 219 -2238 255 -2237
rect 324 -2238 360 -2237
rect 366 -2238 377 -2237
rect 390 -2238 416 -2237
rect 422 -2238 430 -2237
rect 446 -2238 542 -2237
rect 565 -2238 633 -2237
rect 121 -2240 125 -2239
rect 128 -2240 139 -2239
rect 149 -2240 209 -2239
rect 212 -2240 220 -2239
rect 261 -2240 325 -2239
rect 327 -2240 363 -2239
rect 366 -2240 381 -2239
rect 397 -2240 472 -2239
rect 513 -2240 542 -2239
rect 124 -2242 146 -2241
rect 156 -2242 192 -2241
rect 205 -2242 307 -2241
rect 331 -2242 391 -2241
rect 401 -2242 409 -2241
rect 464 -2242 521 -2241
rect 527 -2242 556 -2241
rect 131 -2244 136 -2243
rect 156 -2244 178 -2243
rect 261 -2244 409 -2243
rect 467 -2244 507 -2243
rect 513 -2244 577 -2243
rect 163 -2246 269 -2245
rect 296 -2246 332 -2245
rect 338 -2246 566 -2245
rect 576 -2246 598 -2245
rect 163 -2248 181 -2247
rect 247 -2248 297 -2247
rect 310 -2248 339 -2247
rect 345 -2248 465 -2247
rect 492 -2248 521 -2247
rect 555 -2248 570 -2247
rect 166 -2250 433 -2249
rect 485 -2250 493 -2249
rect 506 -2250 580 -2249
rect 177 -2252 185 -2251
rect 240 -2252 248 -2251
rect 268 -2252 283 -2251
rect 303 -2252 346 -2251
rect 359 -2252 444 -2251
rect 184 -2254 241 -2253
rect 373 -2254 437 -2253
rect 352 -2256 374 -2255
rect 394 -2256 486 -2255
rect 226 -2258 353 -2257
rect 380 -2258 395 -2257
rect 436 -2258 451 -2257
rect 226 -2260 234 -2259
rect 303 -2260 451 -2259
rect 114 -2271 132 -2270
rect 135 -2271 146 -2270
rect 163 -2271 307 -2270
rect 317 -2271 374 -2270
rect 401 -2271 440 -2270
rect 450 -2271 573 -2270
rect 121 -2273 125 -2272
rect 142 -2273 157 -2272
rect 170 -2273 213 -2272
rect 215 -2273 223 -2272
rect 240 -2273 251 -2272
rect 275 -2273 283 -2272
rect 289 -2273 311 -2272
rect 352 -2273 388 -2272
rect 404 -2273 416 -2272
rect 429 -2273 531 -2272
rect 541 -2273 570 -2272
rect 184 -2275 234 -2274
rect 243 -2275 479 -2274
rect 485 -2275 503 -2274
rect 534 -2275 542 -2274
rect 198 -2277 314 -2276
rect 359 -2277 465 -2276
rect 471 -2277 500 -2276
rect 534 -2277 556 -2276
rect 212 -2279 220 -2278
rect 226 -2279 234 -2278
rect 261 -2279 276 -2278
rect 289 -2279 318 -2278
rect 408 -2279 521 -2278
rect 205 -2281 227 -2280
rect 268 -2281 283 -2280
rect 303 -2281 332 -2280
rect 415 -2281 437 -2280
rect 457 -2281 465 -2280
rect 474 -2281 479 -2280
rect 513 -2281 521 -2280
rect 247 -2283 269 -2282
rect 303 -2283 367 -2282
rect 432 -2283 507 -2282
rect 513 -2283 528 -2282
rect 331 -2285 339 -2284
rect 362 -2285 367 -2284
rect 443 -2285 458 -2284
rect 492 -2285 507 -2284
rect 527 -2285 577 -2284
rect 450 -2287 475 -2286
rect 576 -2287 584 -2286
rect 212 -2298 216 -2297
rect 226 -2298 244 -2297
rect 247 -2298 255 -2297
rect 275 -2298 328 -2297
rect 338 -2298 346 -2297
rect 366 -2298 370 -2297
rect 408 -2298 416 -2297
rect 422 -2298 440 -2297
rect 443 -2298 465 -2297
rect 502 -2298 514 -2297
rect 520 -2298 528 -2297
rect 534 -2298 542 -2297
rect 569 -2298 577 -2297
rect 597 -2298 605 -2297
rect 639 -2298 647 -2297
rect 226 -2300 265 -2299
rect 282 -2300 290 -2299
rect 296 -2300 307 -2299
rect 313 -2300 318 -2299
rect 432 -2300 458 -2299
rect 506 -2300 510 -2299
rect 614 -2300 640 -2299
rect 254 -2302 286 -2301
rect 289 -2302 311 -2301
rect 317 -2302 332 -2301
rect 446 -2302 451 -2301
rect 268 -2304 297 -2303
rect 170 -2315 178 -2314
rect 226 -2315 283 -2314
rect 296 -2315 307 -2314
rect 380 -2315 388 -2314
rect 404 -2315 409 -2314
rect 527 -2315 535 -2314
rect 597 -2315 612 -2314
rect 642 -2315 647 -2314
rect 233 -2317 241 -2316
rect 247 -2317 269 -2316
rect 278 -2317 318 -2316
rect 254 -2319 276 -2318
<< m2contact >>
rect 177 0 178 1
rect 191 0 192 1
rect 205 0 206 1
rect 212 0 213 1
rect 257 0 258 1
rect 282 0 283 1
rect 310 0 311 1
rect 348 0 349 1
rect 359 0 360 1
rect 366 0 367 1
rect 271 -2 272 -1
rect 275 -2 276 -1
rect 177 -13 178 -12
rect 187 -13 188 -12
rect 194 -13 195 -12
rect 198 -13 199 -12
rect 212 -13 213 -12
rect 219 -13 220 -12
rect 233 -13 234 -12
rect 254 -13 255 -12
rect 261 -13 262 -12
rect 275 -13 276 -12
rect 303 -13 304 -12
rect 310 -13 311 -12
rect 341 -13 342 -12
rect 394 -13 395 -12
rect 184 -15 185 -14
rect 208 -15 209 -14
rect 215 -15 216 -14
rect 254 -15 255 -14
rect 348 -15 349 -14
rect 387 -15 388 -14
rect 198 -17 199 -16
rect 201 -17 202 -16
rect 240 -17 241 -16
rect 250 -17 251 -16
rect 366 -17 367 -16
rect 373 -17 374 -16
rect 366 -19 367 -18
rect 383 -19 384 -18
rect 166 -30 167 -29
rect 198 -30 199 -29
rect 205 -30 206 -29
rect 271 -30 272 -29
rect 289 -30 290 -29
rect 296 -30 297 -29
rect 299 -30 300 -29
rect 352 -30 353 -29
rect 387 -30 388 -29
rect 429 -30 430 -29
rect 177 -32 178 -31
rect 212 -32 213 -31
rect 215 -32 216 -31
rect 219 -32 220 -31
rect 226 -32 227 -31
rect 240 -32 241 -31
rect 247 -32 248 -31
rect 261 -32 262 -31
rect 268 -32 269 -31
rect 341 -32 342 -31
rect 345 -32 346 -31
rect 366 -32 367 -31
rect 380 -32 381 -31
rect 387 -32 388 -31
rect 394 -32 395 -31
rect 422 -32 423 -31
rect 194 -34 195 -33
rect 275 -34 276 -33
rect 296 -34 297 -33
rect 331 -34 332 -33
rect 373 -34 374 -33
rect 394 -34 395 -33
rect 411 -34 412 -33
rect 450 -34 451 -33
rect 212 -36 213 -35
rect 233 -36 234 -35
rect 254 -36 255 -35
rect 310 -36 311 -35
rect 317 -36 318 -35
rect 334 -36 335 -35
rect 366 -36 367 -35
rect 373 -36 374 -35
rect 380 -36 381 -35
rect 415 -36 416 -35
rect 219 -38 220 -37
rect 254 -38 255 -37
rect 261 -38 262 -37
rect 338 -38 339 -37
rect 233 -40 234 -39
rect 240 -40 241 -39
rect 303 -40 304 -39
rect 324 -40 325 -39
rect 86 -51 87 -50
rect 107 -51 108 -50
rect 121 -51 122 -50
rect 128 -51 129 -50
rect 142 -51 143 -50
rect 170 -51 171 -50
rect 177 -51 178 -50
rect 187 -51 188 -50
rect 191 -51 192 -50
rect 219 -51 220 -50
rect 233 -51 234 -50
rect 310 -51 311 -50
rect 317 -51 318 -50
rect 464 -51 465 -50
rect 579 -51 580 -50
rect 583 -51 584 -50
rect 93 -53 94 -52
rect 100 -53 101 -52
rect 107 -53 108 -52
rect 170 -53 171 -52
rect 177 -53 178 -52
rect 226 -53 227 -52
rect 247 -53 248 -52
rect 296 -53 297 -52
rect 303 -53 304 -52
rect 352 -53 353 -52
rect 355 -53 356 -52
rect 408 -53 409 -52
rect 436 -53 437 -52
rect 485 -53 486 -52
rect 135 -55 136 -54
rect 219 -55 220 -54
rect 247 -55 248 -54
rect 261 -55 262 -54
rect 275 -55 276 -54
rect 373 -55 374 -54
rect 394 -55 395 -54
rect 436 -55 437 -54
rect 443 -55 444 -54
rect 471 -55 472 -54
rect 149 -57 150 -56
rect 243 -57 244 -56
rect 275 -57 276 -56
rect 362 -57 363 -56
rect 376 -57 377 -56
rect 394 -57 395 -56
rect 429 -57 430 -56
rect 443 -57 444 -56
rect 450 -57 451 -56
rect 457 -57 458 -56
rect 163 -59 164 -58
rect 215 -59 216 -58
rect 240 -59 241 -58
rect 261 -59 262 -58
rect 303 -59 304 -58
rect 345 -59 346 -58
rect 348 -59 349 -58
rect 478 -59 479 -58
rect 205 -61 206 -60
rect 317 -61 318 -60
rect 331 -61 332 -60
rect 369 -61 370 -60
rect 422 -61 423 -60
rect 450 -61 451 -60
rect 198 -63 199 -62
rect 205 -63 206 -62
rect 215 -63 216 -62
rect 226 -63 227 -62
rect 324 -63 325 -62
rect 331 -63 332 -62
rect 338 -63 339 -62
rect 380 -63 381 -62
rect 387 -63 388 -62
rect 422 -63 423 -62
rect 100 -65 101 -64
rect 198 -65 199 -64
rect 289 -65 290 -64
rect 387 -65 388 -64
rect 282 -67 283 -66
rect 289 -67 290 -66
rect 310 -67 311 -66
rect 324 -67 325 -66
rect 338 -67 339 -66
rect 415 -67 416 -66
rect 282 -69 283 -68
rect 401 -69 402 -68
rect 341 -71 342 -70
rect 429 -71 430 -70
rect 362 -73 363 -72
rect 499 -73 500 -72
rect 366 -75 367 -74
rect 415 -75 416 -74
rect 401 -77 402 -76
rect 495 -77 496 -76
rect 58 -88 59 -87
rect 135 -88 136 -87
rect 149 -88 150 -87
rect 233 -88 234 -87
rect 282 -88 283 -87
rect 310 -88 311 -87
rect 313 -88 314 -87
rect 415 -88 416 -87
rect 436 -88 437 -87
rect 555 -88 556 -87
rect 565 -88 566 -87
rect 618 -88 619 -87
rect 65 -90 66 -89
rect 142 -90 143 -89
rect 177 -90 178 -89
rect 233 -90 234 -89
rect 247 -90 248 -89
rect 415 -90 416 -89
rect 436 -90 437 -89
rect 506 -90 507 -89
rect 583 -90 584 -89
rect 597 -90 598 -89
rect 72 -92 73 -91
rect 254 -92 255 -91
rect 282 -92 283 -91
rect 289 -92 290 -91
rect 345 -92 346 -91
rect 401 -92 402 -91
rect 450 -92 451 -91
rect 569 -92 570 -91
rect 79 -94 80 -93
rect 114 -94 115 -93
rect 121 -94 122 -93
rect 191 -94 192 -93
rect 205 -94 206 -93
rect 254 -94 255 -93
rect 268 -94 269 -93
rect 401 -94 402 -93
rect 457 -94 458 -93
rect 541 -94 542 -93
rect 86 -96 87 -95
rect 124 -96 125 -95
rect 180 -96 181 -95
rect 527 -96 528 -95
rect 86 -98 87 -97
rect 163 -98 164 -97
rect 184 -98 185 -97
rect 198 -98 199 -97
rect 205 -98 206 -97
rect 226 -98 227 -97
rect 247 -98 248 -97
rect 296 -98 297 -97
rect 317 -98 318 -97
rect 345 -98 346 -97
rect 348 -98 349 -97
rect 464 -98 465 -97
rect 478 -98 479 -97
rect 492 -98 493 -97
rect 93 -100 94 -99
rect 117 -100 118 -99
rect 149 -100 150 -99
rect 184 -100 185 -99
rect 187 -100 188 -99
rect 240 -100 241 -99
rect 268 -100 269 -99
rect 299 -100 300 -99
rect 352 -100 353 -99
rect 429 -100 430 -99
rect 485 -100 486 -99
rect 583 -100 584 -99
rect 93 -102 94 -101
rect 156 -102 157 -101
rect 163 -102 164 -101
rect 170 -102 171 -101
rect 226 -102 227 -101
rect 296 -102 297 -101
rect 331 -102 332 -101
rect 429 -102 430 -101
rect 114 -104 115 -103
rect 243 -104 244 -103
rect 275 -104 276 -103
rect 317 -104 318 -103
rect 331 -104 332 -103
rect 576 -104 577 -103
rect 170 -106 171 -105
rect 285 -106 286 -105
rect 289 -106 290 -105
rect 303 -106 304 -105
rect 355 -106 356 -105
rect 471 -106 472 -105
rect 156 -108 157 -107
rect 303 -108 304 -107
rect 306 -108 307 -107
rect 471 -108 472 -107
rect 243 -110 244 -109
rect 590 -110 591 -109
rect 261 -112 262 -111
rect 275 -112 276 -111
rect 359 -112 360 -111
rect 499 -112 500 -111
rect 222 -114 223 -113
rect 261 -114 262 -113
rect 362 -114 363 -113
rect 383 -114 384 -113
rect 387 -114 388 -113
rect 534 -114 535 -113
rect 107 -116 108 -115
rect 362 -116 363 -115
rect 366 -116 367 -115
rect 450 -116 451 -115
rect 142 -118 143 -117
rect 222 -118 223 -117
rect 369 -118 370 -117
rect 520 -118 521 -117
rect 177 -120 178 -119
rect 366 -120 367 -119
rect 373 -120 374 -119
rect 499 -120 500 -119
rect 100 -122 101 -121
rect 373 -122 374 -121
rect 376 -122 377 -121
rect 513 -122 514 -121
rect 100 -124 101 -123
rect 135 -124 136 -123
rect 387 -124 388 -123
rect 506 -124 507 -123
rect 394 -126 395 -125
rect 457 -126 458 -125
rect 334 -128 335 -127
rect 394 -128 395 -127
rect 408 -128 409 -127
rect 464 -128 465 -127
rect 380 -130 381 -129
rect 408 -130 409 -129
rect 422 -130 423 -129
rect 485 -130 486 -129
rect 422 -132 423 -131
rect 478 -132 479 -131
rect 51 -143 52 -142
rect 187 -143 188 -142
rect 208 -143 209 -142
rect 376 -143 377 -142
rect 380 -143 381 -142
rect 471 -143 472 -142
rect 544 -143 545 -142
rect 572 -143 573 -142
rect 618 -143 619 -142
rect 632 -143 633 -142
rect 642 -143 643 -142
rect 646 -143 647 -142
rect 65 -145 66 -144
rect 194 -145 195 -144
rect 222 -145 223 -144
rect 254 -145 255 -144
rect 282 -145 283 -144
rect 429 -145 430 -144
rect 439 -145 440 -144
rect 576 -145 577 -144
rect 65 -147 66 -146
rect 107 -147 108 -146
rect 121 -147 122 -146
rect 229 -147 230 -146
rect 236 -147 237 -146
rect 275 -147 276 -146
rect 282 -147 283 -146
rect 317 -147 318 -146
rect 320 -147 321 -146
rect 401 -147 402 -146
rect 457 -147 458 -146
rect 471 -147 472 -146
rect 506 -147 507 -146
rect 576 -147 577 -146
rect 72 -149 73 -148
rect 376 -149 377 -148
rect 387 -149 388 -148
rect 569 -149 570 -148
rect 79 -151 80 -150
rect 177 -151 178 -150
rect 180 -151 181 -150
rect 362 -151 363 -150
rect 366 -151 367 -150
rect 541 -151 542 -150
rect 79 -153 80 -152
rect 135 -153 136 -152
rect 138 -153 139 -152
rect 366 -153 367 -152
rect 390 -153 391 -152
rect 562 -153 563 -152
rect 86 -155 87 -154
rect 187 -155 188 -154
rect 247 -155 248 -154
rect 254 -155 255 -154
rect 285 -155 286 -154
rect 415 -155 416 -154
rect 457 -155 458 -154
rect 562 -155 563 -154
rect 86 -157 87 -156
rect 243 -157 244 -156
rect 296 -157 297 -156
rect 534 -157 535 -156
rect 100 -159 101 -158
rect 163 -159 164 -158
rect 173 -159 174 -158
rect 240 -159 241 -158
rect 296 -159 297 -158
rect 520 -159 521 -158
rect 527 -159 528 -158
rect 534 -159 535 -158
rect 107 -161 108 -160
rect 156 -161 157 -160
rect 191 -161 192 -160
rect 247 -161 248 -160
rect 317 -161 318 -160
rect 324 -161 325 -160
rect 331 -161 332 -160
rect 499 -161 500 -160
rect 527 -161 528 -160
rect 590 -161 591 -160
rect 114 -163 115 -162
rect 331 -163 332 -162
rect 341 -163 342 -162
rect 387 -163 388 -162
rect 408 -163 409 -162
rect 415 -163 416 -162
rect 464 -163 465 -162
rect 548 -163 549 -162
rect 114 -165 115 -164
rect 128 -165 129 -164
rect 135 -165 136 -164
rect 212 -165 213 -164
rect 324 -165 325 -164
rect 404 -165 405 -164
rect 408 -165 409 -164
rect 422 -165 423 -164
rect 443 -165 444 -164
rect 464 -165 465 -164
rect 478 -165 479 -164
rect 520 -165 521 -164
rect 121 -167 122 -166
rect 170 -167 171 -166
rect 177 -167 178 -166
rect 212 -167 213 -166
rect 345 -167 346 -166
rect 380 -167 381 -166
rect 394 -167 395 -166
rect 478 -167 479 -166
rect 492 -167 493 -166
rect 499 -167 500 -166
rect 513 -167 514 -166
rect 590 -167 591 -166
rect 128 -169 129 -168
rect 310 -169 311 -168
rect 338 -169 339 -168
rect 345 -169 346 -168
rect 352 -169 353 -168
rect 429 -169 430 -168
rect 436 -169 437 -168
rect 513 -169 514 -168
rect 149 -171 150 -170
rect 306 -171 307 -170
rect 359 -171 360 -170
rect 583 -171 584 -170
rect 149 -173 150 -172
rect 299 -173 300 -172
rect 362 -173 363 -172
rect 443 -173 444 -172
rect 450 -173 451 -172
rect 492 -173 493 -172
rect 583 -173 584 -172
rect 597 -173 598 -172
rect 156 -175 157 -174
rect 205 -175 206 -174
rect 261 -175 262 -174
rect 310 -175 311 -174
rect 355 -175 356 -174
rect 450 -175 451 -174
rect 163 -177 164 -176
rect 352 -177 353 -176
rect 355 -177 356 -176
rect 555 -177 556 -176
rect 170 -179 171 -178
rect 268 -179 269 -178
rect 275 -179 276 -178
rect 359 -179 360 -178
rect 551 -179 552 -178
rect 555 -179 556 -178
rect 205 -181 206 -180
rect 422 -181 423 -180
rect 226 -183 227 -182
rect 268 -183 269 -182
rect 289 -183 290 -182
rect 338 -183 339 -182
rect 198 -185 199 -184
rect 226 -185 227 -184
rect 233 -185 234 -184
rect 261 -185 262 -184
rect 289 -185 290 -184
rect 373 -185 374 -184
rect 93 -187 94 -186
rect 233 -187 234 -186
rect 93 -189 94 -188
rect 142 -189 143 -188
rect 198 -189 199 -188
rect 215 -189 216 -188
rect 58 -191 59 -190
rect 142 -191 143 -190
rect 215 -191 216 -190
rect 219 -191 220 -190
rect 16 -202 17 -201
rect 156 -202 157 -201
rect 187 -202 188 -201
rect 275 -202 276 -201
rect 303 -202 304 -201
rect 639 -202 640 -201
rect 646 -202 647 -201
rect 688 -202 689 -201
rect 37 -204 38 -203
rect 184 -204 185 -203
rect 198 -204 199 -203
rect 296 -204 297 -203
rect 320 -204 321 -203
rect 450 -204 451 -203
rect 460 -204 461 -203
rect 660 -204 661 -203
rect 670 -204 671 -203
rect 674 -204 675 -203
rect 44 -206 45 -205
rect 131 -206 132 -205
rect 205 -206 206 -205
rect 513 -206 514 -205
rect 520 -206 521 -205
rect 653 -206 654 -205
rect 65 -208 66 -207
rect 194 -208 195 -207
rect 212 -208 213 -207
rect 219 -208 220 -207
rect 233 -208 234 -207
rect 401 -208 402 -207
rect 411 -208 412 -207
rect 439 -208 440 -207
rect 467 -208 468 -207
rect 611 -208 612 -207
rect 618 -208 619 -207
rect 632 -208 633 -207
rect 65 -210 66 -209
rect 142 -210 143 -209
rect 233 -210 234 -209
rect 240 -210 241 -209
rect 261 -210 262 -209
rect 275 -210 276 -209
rect 289 -210 290 -209
rect 303 -210 304 -209
rect 331 -210 332 -209
rect 457 -210 458 -209
rect 513 -210 514 -209
rect 548 -210 549 -209
rect 562 -210 563 -209
rect 695 -210 696 -209
rect 79 -212 80 -211
rect 219 -212 220 -211
rect 236 -212 237 -211
rect 296 -212 297 -211
rect 355 -212 356 -211
rect 562 -212 563 -211
rect 569 -212 570 -211
rect 583 -212 584 -211
rect 590 -212 591 -211
rect 632 -212 633 -211
rect 51 -214 52 -213
rect 79 -214 80 -213
rect 86 -214 87 -213
rect 138 -214 139 -213
rect 173 -214 174 -213
rect 289 -214 290 -213
rect 359 -214 360 -213
rect 380 -214 381 -213
rect 390 -214 391 -213
rect 478 -214 479 -213
rect 520 -214 521 -213
rect 555 -214 556 -213
rect 569 -214 570 -213
rect 751 -214 752 -213
rect 86 -216 87 -215
rect 149 -216 150 -215
rect 222 -216 223 -215
rect 380 -216 381 -215
rect 397 -216 398 -215
rect 464 -216 465 -215
rect 471 -216 472 -215
rect 555 -216 556 -215
rect 576 -216 577 -215
rect 681 -216 682 -215
rect 93 -218 94 -217
rect 261 -218 262 -217
rect 268 -218 269 -217
rect 331 -218 332 -217
rect 373 -218 374 -217
rect 625 -218 626 -217
rect 93 -220 94 -219
rect 145 -220 146 -219
rect 198 -220 199 -219
rect 268 -220 269 -219
rect 282 -220 283 -219
rect 373 -220 374 -219
rect 376 -220 377 -219
rect 485 -220 486 -219
rect 492 -220 493 -219
rect 576 -220 577 -219
rect 597 -220 598 -219
rect 667 -220 668 -219
rect 100 -222 101 -221
rect 184 -222 185 -221
rect 240 -222 241 -221
rect 254 -222 255 -221
rect 299 -222 300 -221
rect 471 -222 472 -221
rect 527 -222 528 -221
rect 646 -222 647 -221
rect 30 -224 31 -223
rect 100 -224 101 -223
rect 107 -224 108 -223
rect 191 -224 192 -223
rect 226 -224 227 -223
rect 254 -224 255 -223
rect 397 -224 398 -223
rect 450 -224 451 -223
rect 464 -224 465 -223
rect 534 -224 535 -223
rect 544 -224 545 -223
rect 583 -224 584 -223
rect 23 -226 24 -225
rect 107 -226 108 -225
rect 121 -226 122 -225
rect 149 -226 150 -225
rect 177 -226 178 -225
rect 282 -226 283 -225
rect 324 -226 325 -225
rect 534 -226 535 -225
rect 58 -228 59 -227
rect 226 -228 227 -227
rect 310 -228 311 -227
rect 324 -228 325 -227
rect 404 -228 405 -227
rect 478 -228 479 -227
rect 509 -228 510 -227
rect 527 -228 528 -227
rect 72 -230 73 -229
rect 191 -230 192 -229
rect 247 -230 248 -229
rect 310 -230 311 -229
rect 408 -230 409 -229
rect 548 -230 549 -229
rect 72 -232 73 -231
rect 114 -232 115 -231
rect 121 -232 122 -231
rect 142 -232 143 -231
rect 163 -232 164 -231
rect 247 -232 248 -231
rect 408 -232 409 -231
rect 499 -232 500 -231
rect 114 -234 115 -233
rect 208 -234 209 -233
rect 415 -234 416 -233
rect 436 -234 437 -233
rect 443 -234 444 -233
rect 492 -234 493 -233
rect 128 -236 129 -235
rect 352 -236 353 -235
rect 366 -236 367 -235
rect 443 -236 444 -235
rect 485 -236 486 -235
rect 509 -236 510 -235
rect 128 -238 129 -237
rect 170 -238 171 -237
rect 208 -238 209 -237
rect 541 -238 542 -237
rect 138 -240 139 -239
rect 177 -240 178 -239
rect 338 -240 339 -239
rect 366 -240 367 -239
rect 422 -240 423 -239
rect 590 -240 591 -239
rect 163 -242 164 -241
rect 229 -242 230 -241
rect 338 -242 339 -241
rect 499 -242 500 -241
rect 345 -244 346 -243
rect 415 -244 416 -243
rect 418 -244 419 -243
rect 422 -244 423 -243
rect 429 -244 430 -243
rect 506 -244 507 -243
rect 345 -246 346 -245
rect 387 -246 388 -245
rect 394 -246 395 -245
rect 429 -246 430 -245
rect 394 -248 395 -247
rect 604 -248 605 -247
rect 23 -259 24 -258
rect 135 -259 136 -258
rect 142 -259 143 -258
rect 261 -259 262 -258
rect 299 -259 300 -258
rect 425 -259 426 -258
rect 439 -259 440 -258
rect 576 -259 577 -258
rect 590 -259 591 -258
rect 593 -259 594 -258
rect 597 -259 598 -258
rect 600 -259 601 -258
rect 604 -259 605 -258
rect 670 -259 671 -258
rect 674 -259 675 -258
rect 716 -259 717 -258
rect 751 -259 752 -258
rect 828 -259 829 -258
rect 856 -259 857 -258
rect 859 -259 860 -258
rect 51 -261 52 -260
rect 58 -261 59 -260
rect 65 -261 66 -260
rect 236 -261 237 -260
rect 240 -261 241 -260
rect 271 -261 272 -260
rect 334 -261 335 -260
rect 660 -261 661 -260
rect 681 -261 682 -260
rect 737 -261 738 -260
rect 16 -263 17 -262
rect 240 -263 241 -262
rect 247 -263 248 -262
rect 397 -263 398 -262
rect 401 -263 402 -262
rect 572 -263 573 -262
rect 590 -263 591 -262
rect 639 -263 640 -262
rect 646 -263 647 -262
rect 681 -263 682 -262
rect 688 -263 689 -262
rect 744 -263 745 -262
rect 58 -265 59 -264
rect 79 -265 80 -264
rect 107 -265 108 -264
rect 121 -265 122 -264
rect 128 -265 129 -264
rect 226 -265 227 -264
rect 229 -265 230 -264
rect 254 -265 255 -264
rect 261 -265 262 -264
rect 275 -265 276 -264
rect 338 -265 339 -264
rect 352 -265 353 -264
rect 359 -265 360 -264
rect 408 -265 409 -264
rect 415 -265 416 -264
rect 422 -265 423 -264
rect 443 -265 444 -264
rect 478 -265 479 -264
rect 499 -265 500 -264
rect 502 -265 503 -264
rect 534 -265 535 -264
rect 569 -265 570 -264
rect 597 -265 598 -264
rect 611 -265 612 -264
rect 618 -265 619 -264
rect 667 -265 668 -264
rect 688 -265 689 -264
rect 723 -265 724 -264
rect 44 -267 45 -266
rect 79 -267 80 -266
rect 107 -267 108 -266
rect 156 -267 157 -266
rect 191 -267 192 -266
rect 194 -267 195 -266
rect 205 -267 206 -266
rect 226 -267 227 -266
rect 268 -267 269 -266
rect 352 -267 353 -266
rect 359 -267 360 -266
rect 401 -267 402 -266
rect 446 -267 447 -266
rect 604 -267 605 -266
rect 625 -267 626 -266
rect 709 -267 710 -266
rect 68 -269 69 -268
rect 100 -269 101 -268
rect 114 -269 115 -268
rect 159 -269 160 -268
rect 184 -269 185 -268
rect 268 -269 269 -268
rect 275 -269 276 -268
rect 310 -269 311 -268
rect 341 -269 342 -268
rect 457 -269 458 -268
rect 460 -269 461 -268
rect 730 -269 731 -268
rect 72 -271 73 -270
rect 138 -271 139 -270
rect 149 -271 150 -270
rect 156 -271 157 -270
rect 177 -271 178 -270
rect 184 -271 185 -270
rect 205 -271 206 -270
rect 296 -271 297 -270
rect 310 -271 311 -270
rect 317 -271 318 -270
rect 373 -271 374 -270
rect 397 -271 398 -270
rect 481 -271 482 -270
rect 667 -271 668 -270
rect 37 -273 38 -272
rect 177 -273 178 -272
rect 215 -273 216 -272
rect 404 -273 405 -272
rect 499 -273 500 -272
rect 513 -273 514 -272
rect 520 -273 521 -272
rect 625 -273 626 -272
rect 632 -273 633 -272
rect 646 -273 647 -272
rect 30 -275 31 -274
rect 215 -275 216 -274
rect 222 -275 223 -274
rect 282 -275 283 -274
rect 296 -275 297 -274
rect 303 -275 304 -274
rect 317 -275 318 -274
rect 324 -275 325 -274
rect 373 -275 374 -274
rect 751 -275 752 -274
rect 30 -277 31 -276
rect 86 -277 87 -276
rect 100 -277 101 -276
rect 103 -277 104 -276
rect 117 -277 118 -276
rect 632 -277 633 -276
rect 639 -277 640 -276
rect 653 -277 654 -276
rect 37 -279 38 -278
rect 93 -279 94 -278
rect 121 -279 122 -278
rect 198 -279 199 -278
rect 282 -279 283 -278
rect 331 -279 332 -278
rect 380 -279 381 -278
rect 464 -279 465 -278
rect 471 -279 472 -278
rect 520 -279 521 -278
rect 541 -279 542 -278
rect 618 -279 619 -278
rect 72 -281 73 -280
rect 163 -281 164 -280
rect 180 -281 181 -280
rect 198 -281 199 -280
rect 243 -281 244 -280
rect 380 -281 381 -280
rect 390 -281 391 -280
rect 544 -281 545 -280
rect 555 -281 556 -280
rect 660 -281 661 -280
rect 86 -283 87 -282
rect 331 -283 332 -282
rect 394 -283 395 -282
rect 534 -283 535 -282
rect 562 -283 563 -282
rect 576 -283 577 -282
rect 600 -283 601 -282
rect 611 -283 612 -282
rect 93 -285 94 -284
rect 254 -285 255 -284
rect 289 -285 290 -284
rect 303 -285 304 -284
rect 324 -285 325 -284
rect 366 -285 367 -284
rect 429 -285 430 -284
rect 471 -285 472 -284
rect 527 -285 528 -284
rect 555 -285 556 -284
rect 565 -285 566 -284
rect 702 -285 703 -284
rect 149 -287 150 -286
rect 170 -287 171 -286
rect 345 -287 346 -286
rect 366 -287 367 -286
rect 411 -287 412 -286
rect 527 -287 528 -286
rect 163 -289 164 -288
rect 541 -289 542 -288
rect 170 -291 171 -290
rect 233 -291 234 -290
rect 345 -291 346 -290
rect 548 -291 549 -290
rect 387 -293 388 -292
rect 548 -293 549 -292
rect 387 -295 388 -294
rect 695 -295 696 -294
rect 429 -297 430 -296
rect 436 -297 437 -296
rect 450 -297 451 -296
rect 562 -297 563 -296
rect 422 -299 423 -298
rect 450 -299 451 -298
rect 506 -299 507 -298
rect 695 -299 696 -298
rect 338 -301 339 -300
rect 506 -301 507 -300
rect 2 -312 3 -311
rect 100 -312 101 -311
rect 107 -312 108 -311
rect 114 -312 115 -311
rect 121 -312 122 -311
rect 124 -312 125 -311
rect 128 -312 129 -311
rect 495 -312 496 -311
rect 653 -312 654 -311
rect 835 -312 836 -311
rect 849 -312 850 -311
rect 863 -312 864 -311
rect 9 -314 10 -313
rect 65 -314 66 -313
rect 72 -314 73 -313
rect 215 -314 216 -313
rect 233 -314 234 -313
rect 345 -314 346 -313
rect 352 -314 353 -313
rect 562 -314 563 -313
rect 590 -314 591 -313
rect 653 -314 654 -313
rect 674 -314 675 -313
rect 677 -314 678 -313
rect 681 -314 682 -313
rect 723 -314 724 -313
rect 726 -314 727 -313
rect 870 -314 871 -313
rect 16 -316 17 -315
rect 79 -316 80 -315
rect 114 -316 115 -315
rect 415 -316 416 -315
rect 422 -316 423 -315
rect 492 -316 493 -315
rect 534 -316 535 -315
rect 562 -316 563 -315
rect 569 -316 570 -315
rect 590 -316 591 -315
rect 695 -316 696 -315
rect 779 -316 780 -315
rect 828 -316 829 -315
rect 891 -316 892 -315
rect 23 -318 24 -317
rect 177 -318 178 -317
rect 215 -318 216 -317
rect 247 -318 248 -317
rect 257 -318 258 -317
rect 261 -318 262 -317
rect 275 -318 276 -317
rect 341 -318 342 -317
rect 352 -318 353 -317
rect 485 -318 486 -317
rect 513 -318 514 -317
rect 534 -318 535 -317
rect 548 -318 549 -317
rect 569 -318 570 -317
rect 597 -318 598 -317
rect 695 -318 696 -317
rect 702 -318 703 -317
rect 814 -318 815 -317
rect 852 -318 853 -317
rect 856 -318 857 -317
rect 30 -320 31 -319
rect 79 -320 80 -319
rect 96 -320 97 -319
rect 177 -320 178 -319
rect 219 -320 220 -319
rect 345 -320 346 -319
rect 359 -320 360 -319
rect 432 -320 433 -319
rect 450 -320 451 -319
rect 453 -320 454 -319
rect 513 -320 514 -319
rect 520 -320 521 -319
rect 544 -320 545 -319
rect 702 -320 703 -319
rect 709 -320 710 -319
rect 758 -320 759 -319
rect 44 -322 45 -321
rect 107 -322 108 -321
rect 121 -322 122 -321
rect 394 -322 395 -321
rect 401 -322 402 -321
rect 660 -322 661 -321
rect 667 -322 668 -321
rect 709 -322 710 -321
rect 730 -322 731 -321
rect 828 -322 829 -321
rect 44 -324 45 -323
rect 236 -324 237 -323
rect 240 -324 241 -323
rect 443 -324 444 -323
rect 450 -324 451 -323
rect 471 -324 472 -323
rect 520 -324 521 -323
rect 527 -324 528 -323
rect 583 -324 584 -323
rect 597 -324 598 -323
rect 618 -324 619 -323
rect 660 -324 661 -323
rect 737 -324 738 -323
rect 807 -324 808 -323
rect 51 -326 52 -325
rect 338 -326 339 -325
rect 362 -326 363 -325
rect 800 -326 801 -325
rect 51 -328 52 -327
rect 184 -328 185 -327
rect 233 -328 234 -327
rect 793 -328 794 -327
rect 37 -330 38 -329
rect 184 -330 185 -329
rect 240 -330 241 -329
rect 282 -330 283 -329
rect 289 -330 290 -329
rect 681 -330 682 -329
rect 744 -330 745 -329
rect 786 -330 787 -329
rect 58 -332 59 -331
rect 131 -332 132 -331
rect 135 -332 136 -331
rect 222 -332 223 -331
rect 247 -332 248 -331
rect 317 -332 318 -331
rect 334 -332 335 -331
rect 408 -332 409 -331
rect 471 -332 472 -331
rect 478 -332 479 -331
rect 499 -332 500 -331
rect 527 -332 528 -331
rect 583 -332 584 -331
rect 632 -332 633 -331
rect 639 -332 640 -331
rect 730 -332 731 -331
rect 751 -332 752 -331
rect 821 -332 822 -331
rect 58 -334 59 -333
rect 149 -334 150 -333
rect 212 -334 213 -333
rect 408 -334 409 -333
rect 474 -334 475 -333
rect 618 -334 619 -333
rect 639 -334 640 -333
rect 877 -334 878 -333
rect 65 -336 66 -335
rect 191 -336 192 -335
rect 261 -336 262 -335
rect 303 -336 304 -335
rect 310 -336 311 -335
rect 338 -336 339 -335
rect 373 -336 374 -335
rect 765 -336 766 -335
rect 75 -338 76 -337
rect 152 -338 153 -337
rect 170 -338 171 -337
rect 191 -338 192 -337
rect 282 -338 283 -337
rect 324 -338 325 -337
rect 380 -338 381 -337
rect 548 -338 549 -337
rect 586 -338 587 -337
rect 856 -338 857 -337
rect 86 -340 87 -339
rect 317 -340 318 -339
rect 380 -340 381 -339
rect 387 -340 388 -339
rect 394 -340 395 -339
rect 457 -340 458 -339
rect 506 -340 507 -339
rect 632 -340 633 -339
rect 646 -340 647 -339
rect 667 -340 668 -339
rect 688 -340 689 -339
rect 751 -340 752 -339
rect 86 -342 87 -341
rect 268 -342 269 -341
rect 289 -342 290 -341
rect 324 -342 325 -341
rect 401 -342 402 -341
rect 425 -342 426 -341
rect 436 -342 437 -341
rect 688 -342 689 -341
rect 93 -344 94 -343
rect 310 -344 311 -343
rect 429 -344 430 -343
rect 436 -344 437 -343
rect 457 -344 458 -343
rect 464 -344 465 -343
rect 516 -344 517 -343
rect 744 -344 745 -343
rect 93 -346 94 -345
rect 842 -346 843 -345
rect 100 -348 101 -347
rect 359 -348 360 -347
rect 429 -348 430 -347
rect 499 -348 500 -347
rect 604 -348 605 -347
rect 737 -348 738 -347
rect 128 -350 129 -349
rect 219 -350 220 -349
rect 254 -350 255 -349
rect 387 -350 388 -349
rect 604 -350 605 -349
rect 611 -350 612 -349
rect 625 -350 626 -349
rect 646 -350 647 -349
rect 138 -352 139 -351
rect 275 -352 276 -351
rect 296 -352 297 -351
rect 404 -352 405 -351
rect 576 -352 577 -351
rect 611 -352 612 -351
rect 142 -354 143 -353
rect 369 -354 370 -353
rect 555 -354 556 -353
rect 576 -354 577 -353
rect 30 -356 31 -355
rect 142 -356 143 -355
rect 145 -356 146 -355
rect 485 -356 486 -355
rect 156 -358 157 -357
rect 170 -358 171 -357
rect 198 -358 199 -357
rect 464 -358 465 -357
rect 156 -360 157 -359
rect 163 -360 164 -359
rect 254 -360 255 -359
rect 327 -360 328 -359
rect 331 -360 332 -359
rect 555 -360 556 -359
rect 37 -362 38 -361
rect 331 -362 332 -361
rect 334 -362 335 -361
rect 625 -362 626 -361
rect 163 -364 164 -363
rect 205 -364 206 -363
rect 268 -364 269 -363
rect 439 -364 440 -363
rect 453 -364 454 -363
rect 478 -364 479 -363
rect 205 -366 206 -365
rect 415 -366 416 -365
rect 299 -368 300 -367
rect 541 -368 542 -367
rect 303 -370 304 -369
rect 366 -370 367 -369
rect 366 -372 367 -371
rect 772 -372 773 -371
rect 2 -383 3 -382
rect 198 -383 199 -382
rect 205 -383 206 -382
rect 940 -383 941 -382
rect 2 -385 3 -384
rect 198 -385 199 -384
rect 261 -385 262 -384
rect 362 -385 363 -384
rect 369 -385 370 -384
rect 534 -385 535 -384
rect 621 -385 622 -384
rect 639 -385 640 -384
rect 828 -385 829 -384
rect 877 -385 878 -384
rect 16 -387 17 -386
rect 131 -387 132 -386
rect 159 -387 160 -386
rect 905 -387 906 -386
rect 16 -389 17 -388
rect 44 -389 45 -388
rect 51 -389 52 -388
rect 215 -389 216 -388
rect 261 -389 262 -388
rect 432 -389 433 -388
rect 478 -389 479 -388
rect 513 -389 514 -388
rect 516 -389 517 -388
rect 737 -389 738 -388
rect 842 -389 843 -388
rect 898 -389 899 -388
rect 23 -391 24 -390
rect 243 -391 244 -390
rect 275 -391 276 -390
rect 432 -391 433 -390
rect 436 -391 437 -390
rect 478 -391 479 -390
rect 502 -391 503 -390
rect 807 -391 808 -390
rect 852 -391 853 -390
rect 891 -391 892 -390
rect 23 -393 24 -392
rect 177 -393 178 -392
rect 282 -393 283 -392
rect 376 -393 377 -392
rect 390 -393 391 -392
rect 779 -393 780 -392
rect 807 -393 808 -392
rect 849 -393 850 -392
rect 863 -393 864 -392
rect 884 -393 885 -392
rect 37 -395 38 -394
rect 506 -395 507 -394
rect 509 -395 510 -394
rect 933 -395 934 -394
rect 37 -397 38 -396
rect 103 -397 104 -396
rect 107 -397 108 -396
rect 222 -397 223 -396
rect 310 -397 311 -396
rect 348 -397 349 -396
rect 359 -397 360 -396
rect 653 -397 654 -396
rect 716 -397 717 -396
rect 891 -397 892 -396
rect 44 -399 45 -398
rect 177 -399 178 -398
rect 184 -399 185 -398
rect 282 -399 283 -398
rect 303 -399 304 -398
rect 310 -399 311 -398
rect 317 -399 318 -398
rect 492 -399 493 -398
rect 495 -399 496 -398
rect 884 -399 885 -398
rect 54 -401 55 -400
rect 135 -401 136 -400
rect 145 -401 146 -400
rect 863 -401 864 -400
rect 870 -401 871 -400
rect 926 -401 927 -400
rect 75 -403 76 -402
rect 268 -403 269 -402
rect 303 -403 304 -402
rect 821 -403 822 -402
rect 79 -405 80 -404
rect 96 -405 97 -404
rect 100 -405 101 -404
rect 184 -405 185 -404
rect 201 -405 202 -404
rect 268 -405 269 -404
rect 324 -405 325 -404
rect 394 -405 395 -404
rect 401 -405 402 -404
rect 457 -405 458 -404
rect 520 -405 521 -404
rect 583 -405 584 -404
rect 604 -405 605 -404
rect 639 -405 640 -404
rect 674 -405 675 -404
rect 870 -405 871 -404
rect 9 -407 10 -406
rect 79 -407 80 -406
rect 86 -407 87 -406
rect 233 -407 234 -406
rect 240 -407 241 -406
rect 359 -407 360 -406
rect 373 -407 374 -406
rect 828 -407 829 -406
rect 9 -409 10 -408
rect 219 -409 220 -408
rect 240 -409 241 -408
rect 317 -409 318 -408
rect 331 -409 332 -408
rect 352 -409 353 -408
rect 408 -409 409 -408
rect 509 -409 510 -408
rect 520 -409 521 -408
rect 751 -409 752 -408
rect 772 -409 773 -408
rect 849 -409 850 -408
rect 72 -411 73 -410
rect 352 -411 353 -410
rect 369 -411 370 -410
rect 408 -411 409 -410
rect 415 -411 416 -410
rect 534 -411 535 -410
rect 555 -411 556 -410
rect 653 -411 654 -410
rect 695 -411 696 -410
rect 772 -411 773 -410
rect 814 -411 815 -410
rect 821 -411 822 -410
rect 72 -413 73 -412
rect 163 -413 164 -412
rect 170 -413 171 -412
rect 205 -413 206 -412
rect 212 -413 213 -412
rect 779 -413 780 -412
rect 86 -415 87 -414
rect 156 -415 157 -414
rect 163 -415 164 -414
rect 569 -415 570 -414
rect 576 -415 577 -414
rect 604 -415 605 -414
rect 625 -415 626 -414
rect 695 -415 696 -414
rect 716 -415 717 -414
rect 800 -415 801 -414
rect 93 -417 94 -416
rect 247 -417 248 -416
rect 254 -417 255 -416
rect 373 -417 374 -416
rect 422 -417 423 -416
rect 842 -417 843 -416
rect 65 -419 66 -418
rect 254 -419 255 -418
rect 289 -419 290 -418
rect 394 -419 395 -418
rect 422 -419 423 -418
rect 681 -419 682 -418
rect 730 -419 731 -418
rect 814 -419 815 -418
rect 58 -421 59 -420
rect 65 -421 66 -420
rect 107 -421 108 -420
rect 366 -421 367 -420
rect 425 -421 426 -420
rect 597 -421 598 -420
rect 611 -421 612 -420
rect 625 -421 626 -420
rect 646 -421 647 -420
rect 681 -421 682 -420
rect 730 -421 731 -420
rect 765 -421 766 -420
rect 58 -423 59 -422
rect 296 -423 297 -422
rect 338 -423 339 -422
rect 947 -423 948 -422
rect 110 -425 111 -424
rect 247 -425 248 -424
rect 289 -425 290 -424
rect 380 -425 381 -424
rect 436 -425 437 -424
rect 835 -425 836 -424
rect 117 -427 118 -426
rect 383 -427 384 -426
rect 450 -427 451 -426
rect 457 -427 458 -426
rect 471 -427 472 -426
rect 800 -427 801 -426
rect 835 -427 836 -426
rect 856 -427 857 -426
rect 114 -429 115 -428
rect 471 -429 472 -428
rect 485 -429 486 -428
rect 576 -429 577 -428
rect 590 -429 591 -428
rect 674 -429 675 -428
rect 688 -429 689 -428
rect 765 -429 766 -428
rect 114 -431 115 -430
rect 569 -431 570 -430
rect 632 -431 633 -430
rect 856 -431 857 -430
rect 121 -433 122 -432
rect 401 -433 402 -432
rect 418 -433 419 -432
rect 450 -433 451 -432
rect 523 -433 524 -432
rect 919 -433 920 -432
rect 121 -435 122 -434
rect 149 -435 150 -434
rect 156 -435 157 -434
rect 334 -435 335 -434
rect 345 -435 346 -434
rect 513 -435 514 -434
rect 527 -435 528 -434
rect 590 -435 591 -434
rect 646 -435 647 -434
rect 667 -435 668 -434
rect 688 -435 689 -434
rect 709 -435 710 -434
rect 751 -435 752 -434
rect 786 -435 787 -434
rect 30 -437 31 -436
rect 149 -437 150 -436
rect 212 -437 213 -436
rect 912 -437 913 -436
rect 30 -439 31 -438
rect 128 -439 129 -438
rect 135 -439 136 -438
rect 306 -439 307 -438
rect 366 -439 367 -438
rect 597 -439 598 -438
rect 618 -439 619 -438
rect 786 -439 787 -438
rect 128 -441 129 -440
rect 191 -441 192 -440
rect 233 -441 234 -440
rect 485 -441 486 -440
rect 548 -441 549 -440
rect 632 -441 633 -440
rect 667 -441 668 -440
rect 744 -441 745 -440
rect 142 -443 143 -442
rect 170 -443 171 -442
rect 191 -443 192 -442
rect 338 -443 339 -442
rect 404 -443 405 -442
rect 527 -443 528 -442
rect 555 -443 556 -442
rect 562 -443 563 -442
rect 611 -443 612 -442
rect 618 -443 619 -442
rect 702 -443 703 -442
rect 709 -443 710 -442
rect 142 -445 143 -444
rect 429 -445 430 -444
rect 443 -445 444 -444
rect 548 -445 549 -444
rect 702 -445 703 -444
rect 793 -445 794 -444
rect 152 -447 153 -446
rect 744 -447 745 -446
rect 296 -449 297 -448
rect 737 -449 738 -448
rect 331 -451 332 -450
rect 429 -451 430 -450
rect 541 -451 542 -450
rect 562 -451 563 -450
rect 723 -451 724 -450
rect 793 -451 794 -450
rect 299 -453 300 -452
rect 723 -453 724 -452
rect 387 -455 388 -454
rect 443 -455 444 -454
rect 499 -455 500 -454
rect 541 -455 542 -454
rect 278 -457 279 -456
rect 499 -457 500 -456
rect 387 -459 388 -458
rect 464 -459 465 -458
rect 415 -461 416 -460
rect 464 -461 465 -460
rect 2 -472 3 -471
rect 264 -472 265 -471
rect 268 -472 269 -471
rect 425 -472 426 -471
rect 429 -472 430 -471
rect 814 -472 815 -471
rect 2 -474 3 -473
rect 219 -474 220 -473
rect 243 -474 244 -473
rect 513 -474 514 -473
rect 544 -474 545 -473
rect 891 -474 892 -473
rect 9 -476 10 -475
rect 520 -476 521 -475
rect 607 -476 608 -475
rect 618 -476 619 -475
rect 726 -476 727 -475
rect 821 -476 822 -475
rect 9 -478 10 -477
rect 44 -478 45 -477
rect 51 -478 52 -477
rect 145 -478 146 -477
rect 180 -478 181 -477
rect 201 -478 202 -477
rect 212 -478 213 -477
rect 940 -478 941 -477
rect 30 -480 31 -479
rect 51 -480 52 -479
rect 54 -480 55 -479
rect 695 -480 696 -479
rect 814 -480 815 -479
rect 919 -480 920 -479
rect 30 -482 31 -481
rect 37 -482 38 -481
rect 58 -482 59 -481
rect 303 -482 304 -481
rect 313 -482 314 -481
rect 947 -482 948 -481
rect 37 -484 38 -483
rect 383 -484 384 -483
rect 394 -484 395 -483
rect 418 -484 419 -483
rect 439 -484 440 -483
rect 796 -484 797 -483
rect 58 -486 59 -485
rect 135 -486 136 -485
rect 184 -486 185 -485
rect 219 -486 220 -485
rect 243 -486 244 -485
rect 282 -486 283 -485
rect 303 -486 304 -485
rect 317 -486 318 -485
rect 320 -486 321 -485
rect 548 -486 549 -485
rect 695 -486 696 -485
rect 702 -486 703 -485
rect 79 -488 80 -487
rect 96 -488 97 -487
rect 100 -488 101 -487
rect 653 -488 654 -487
rect 660 -488 661 -487
rect 702 -488 703 -487
rect 23 -490 24 -489
rect 79 -490 80 -489
rect 86 -490 87 -489
rect 198 -490 199 -489
rect 324 -490 325 -489
rect 394 -490 395 -489
rect 401 -490 402 -489
rect 821 -490 822 -489
rect 86 -492 87 -491
rect 247 -492 248 -491
rect 352 -492 353 -491
rect 432 -492 433 -491
rect 460 -492 461 -491
rect 765 -492 766 -491
rect 100 -494 101 -493
rect 107 -494 108 -493
rect 114 -494 115 -493
rect 390 -494 391 -493
rect 408 -494 409 -493
rect 429 -494 430 -493
rect 464 -494 465 -493
rect 523 -494 524 -493
rect 541 -494 542 -493
rect 548 -494 549 -493
rect 639 -494 640 -493
rect 660 -494 661 -493
rect 765 -494 766 -493
rect 835 -494 836 -493
rect 82 -496 83 -495
rect 107 -496 108 -495
rect 117 -496 118 -495
rect 674 -496 675 -495
rect 835 -496 836 -495
rect 842 -496 843 -495
rect 121 -498 122 -497
rect 408 -498 409 -497
rect 415 -498 416 -497
rect 793 -498 794 -497
rect 121 -500 122 -499
rect 345 -500 346 -499
rect 359 -500 360 -499
rect 369 -500 370 -499
rect 373 -500 374 -499
rect 401 -500 402 -499
rect 415 -500 416 -499
rect 576 -500 577 -499
rect 639 -500 640 -499
rect 667 -500 668 -499
rect 674 -500 675 -499
rect 688 -500 689 -499
rect 128 -502 129 -501
rect 296 -502 297 -501
rect 324 -502 325 -501
rect 541 -502 542 -501
rect 576 -502 577 -501
rect 604 -502 605 -501
rect 646 -502 647 -501
rect 653 -502 654 -501
rect 667 -502 668 -501
rect 754 -502 755 -501
rect 16 -504 17 -503
rect 128 -504 129 -503
rect 135 -504 136 -503
rect 310 -504 311 -503
rect 366 -504 367 -503
rect 471 -504 472 -503
rect 485 -504 486 -503
rect 779 -504 780 -503
rect 16 -506 17 -505
rect 163 -506 164 -505
rect 166 -506 167 -505
rect 485 -506 486 -505
rect 488 -506 489 -505
rect 870 -506 871 -505
rect 142 -508 143 -507
rect 352 -508 353 -507
rect 373 -508 374 -507
rect 534 -508 535 -507
rect 646 -508 647 -507
rect 849 -508 850 -507
rect 149 -510 150 -509
rect 166 -510 167 -509
rect 177 -510 178 -509
rect 282 -510 283 -509
rect 296 -510 297 -509
rect 334 -510 335 -509
rect 338 -510 339 -509
rect 366 -510 367 -509
rect 380 -510 381 -509
rect 632 -510 633 -509
rect 688 -510 689 -509
rect 737 -510 738 -509
rect 779 -510 780 -509
rect 884 -510 885 -509
rect 65 -512 66 -511
rect 149 -512 150 -511
rect 156 -512 157 -511
rect 471 -512 472 -511
rect 502 -512 503 -511
rect 898 -512 899 -511
rect 65 -514 66 -513
rect 348 -514 349 -513
rect 464 -514 465 -513
rect 481 -514 482 -513
rect 506 -514 507 -513
rect 786 -514 787 -513
rect 163 -516 164 -515
rect 422 -516 423 -515
rect 509 -516 510 -515
rect 856 -516 857 -515
rect 184 -518 185 -517
rect 226 -518 227 -517
rect 247 -518 248 -517
rect 387 -518 388 -517
rect 422 -518 423 -517
rect 583 -518 584 -517
rect 632 -518 633 -517
rect 681 -518 682 -517
rect 709 -518 710 -517
rect 737 -518 738 -517
rect 786 -518 787 -517
rect 933 -518 934 -517
rect 191 -520 192 -519
rect 772 -520 773 -519
rect 856 -520 857 -519
rect 926 -520 927 -519
rect 93 -522 94 -521
rect 191 -522 192 -521
rect 194 -522 195 -521
rect 240 -522 241 -521
rect 254 -522 255 -521
rect 345 -522 346 -521
rect 387 -522 388 -521
rect 590 -522 591 -521
rect 709 -522 710 -521
rect 800 -522 801 -521
rect 93 -524 94 -523
rect 306 -524 307 -523
rect 341 -524 342 -523
rect 534 -524 535 -523
rect 569 -524 570 -523
rect 583 -524 584 -523
rect 590 -524 591 -523
rect 597 -524 598 -523
rect 751 -524 752 -523
rect 772 -524 773 -523
rect 800 -524 801 -523
rect 912 -524 913 -523
rect 198 -526 199 -525
rect 233 -526 234 -525
rect 240 -526 241 -525
rect 905 -526 906 -525
rect 226 -528 227 -527
rect 492 -528 493 -527
rect 513 -528 514 -527
rect 527 -528 528 -527
rect 597 -528 598 -527
rect 625 -528 626 -527
rect 233 -530 234 -529
rect 499 -530 500 -529
rect 520 -530 521 -529
rect 744 -530 745 -529
rect 254 -532 255 -531
rect 275 -532 276 -531
rect 289 -532 290 -531
rect 380 -532 381 -531
rect 436 -532 437 -531
rect 569 -532 570 -531
rect 611 -532 612 -531
rect 625 -532 626 -531
rect 744 -532 745 -531
rect 758 -532 759 -531
rect 205 -534 206 -533
rect 275 -534 276 -533
rect 289 -534 290 -533
rect 331 -534 332 -533
rect 453 -534 454 -533
rect 611 -534 612 -533
rect 730 -534 731 -533
rect 758 -534 759 -533
rect 72 -536 73 -535
rect 205 -536 206 -535
rect 268 -536 269 -535
rect 310 -536 311 -535
rect 457 -536 458 -535
rect 681 -536 682 -535
rect 730 -536 731 -535
rect 828 -536 829 -535
rect 72 -538 73 -537
rect 450 -538 451 -537
rect 457 -538 458 -537
rect 478 -538 479 -537
rect 499 -538 500 -537
rect 863 -538 864 -537
rect 450 -540 451 -539
rect 495 -540 496 -539
rect 527 -540 528 -539
rect 562 -540 563 -539
rect 478 -542 479 -541
rect 723 -542 724 -541
rect 555 -544 556 -543
rect 562 -544 563 -543
rect 723 -544 724 -543
rect 877 -544 878 -543
rect 261 -546 262 -545
rect 555 -546 556 -545
rect 261 -548 262 -547
rect 436 -548 437 -547
rect 2 -559 3 -558
rect 481 -559 482 -558
rect 502 -559 503 -558
rect 576 -559 577 -558
rect 583 -559 584 -558
rect 604 -559 605 -558
rect 607 -559 608 -558
rect 625 -559 626 -558
rect 681 -559 682 -558
rect 898 -559 899 -558
rect 2 -561 3 -560
rect 30 -561 31 -560
rect 37 -561 38 -560
rect 96 -561 97 -560
rect 131 -561 132 -560
rect 163 -561 164 -560
rect 177 -561 178 -560
rect 317 -561 318 -560
rect 345 -561 346 -560
rect 362 -561 363 -560
rect 373 -561 374 -560
rect 495 -561 496 -560
rect 506 -561 507 -560
rect 537 -561 538 -560
rect 541 -561 542 -560
rect 828 -561 829 -560
rect 835 -561 836 -560
rect 842 -561 843 -560
rect 9 -563 10 -562
rect 124 -563 125 -562
rect 135 -563 136 -562
rect 331 -563 332 -562
rect 373 -563 374 -562
rect 401 -563 402 -562
rect 404 -563 405 -562
rect 884 -563 885 -562
rect 9 -565 10 -564
rect 86 -565 87 -564
rect 156 -565 157 -564
rect 243 -565 244 -564
rect 317 -565 318 -564
rect 523 -565 524 -564
rect 544 -565 545 -564
rect 905 -565 906 -564
rect 23 -567 24 -566
rect 180 -567 181 -566
rect 191 -567 192 -566
rect 341 -567 342 -566
rect 401 -567 402 -566
rect 478 -567 479 -566
rect 520 -567 521 -566
rect 625 -567 626 -566
rect 646 -567 647 -566
rect 835 -567 836 -566
rect 23 -569 24 -568
rect 51 -569 52 -568
rect 58 -569 59 -568
rect 261 -569 262 -568
rect 415 -569 416 -568
rect 450 -569 451 -568
rect 453 -569 454 -568
rect 527 -569 528 -568
rect 555 -569 556 -568
rect 726 -569 727 -568
rect 744 -569 745 -568
rect 751 -569 752 -568
rect 754 -569 755 -568
rect 926 -569 927 -568
rect 30 -571 31 -570
rect 306 -571 307 -570
rect 436 -571 437 -570
rect 509 -571 510 -570
rect 562 -571 563 -570
rect 576 -571 577 -570
rect 583 -571 584 -570
rect 597 -571 598 -570
rect 660 -571 661 -570
rect 681 -571 682 -570
rect 695 -571 696 -570
rect 751 -571 752 -570
rect 765 -571 766 -570
rect 849 -571 850 -570
rect 40 -573 41 -572
rect 341 -573 342 -572
rect 429 -573 430 -572
rect 436 -573 437 -572
rect 457 -573 458 -572
rect 555 -573 556 -572
rect 597 -573 598 -572
rect 688 -573 689 -572
rect 723 -573 724 -572
rect 947 -573 948 -572
rect 44 -575 45 -574
rect 86 -575 87 -574
rect 103 -575 104 -574
rect 261 -575 262 -574
rect 348 -575 349 -574
rect 429 -575 430 -574
rect 457 -575 458 -574
rect 513 -575 514 -574
rect 548 -575 549 -574
rect 562 -575 563 -574
rect 618 -575 619 -574
rect 723 -575 724 -574
rect 744 -575 745 -574
rect 758 -575 759 -574
rect 772 -575 773 -574
rect 891 -575 892 -574
rect 51 -577 52 -576
rect 121 -577 122 -576
rect 128 -577 129 -576
rect 548 -577 549 -576
rect 653 -577 654 -576
rect 660 -577 661 -576
rect 698 -577 699 -576
rect 772 -577 773 -576
rect 786 -577 787 -576
rect 912 -577 913 -576
rect 65 -579 66 -578
rect 68 -579 69 -578
rect 79 -579 80 -578
rect 390 -579 391 -578
rect 474 -579 475 -578
rect 632 -579 633 -578
rect 702 -579 703 -578
rect 758 -579 759 -578
rect 793 -579 794 -578
rect 856 -579 857 -578
rect 65 -581 66 -580
rect 313 -581 314 -580
rect 338 -581 339 -580
rect 786 -581 787 -580
rect 800 -581 801 -580
rect 870 -581 871 -580
rect 79 -583 80 -582
rect 184 -583 185 -582
rect 191 -583 192 -582
rect 331 -583 332 -582
rect 485 -583 486 -582
rect 765 -583 766 -582
rect 779 -583 780 -582
rect 856 -583 857 -582
rect 93 -585 94 -584
rect 793 -585 794 -584
rect 800 -585 801 -584
rect 807 -585 808 -584
rect 814 -585 815 -584
rect 863 -585 864 -584
rect 93 -587 94 -586
rect 100 -587 101 -586
rect 135 -587 136 -586
rect 688 -587 689 -586
rect 730 -587 731 -586
rect 807 -587 808 -586
rect 159 -589 160 -588
rect 240 -589 241 -588
rect 264 -589 265 -588
rect 730 -589 731 -588
rect 737 -589 738 -588
rect 814 -589 815 -588
rect 166 -591 167 -590
rect 646 -591 647 -590
rect 173 -593 174 -592
rect 177 -593 178 -592
rect 184 -593 185 -592
rect 198 -593 199 -592
rect 205 -593 206 -592
rect 877 -593 878 -592
rect 198 -595 199 -594
rect 296 -595 297 -594
rect 313 -595 314 -594
rect 443 -595 444 -594
rect 471 -595 472 -594
rect 779 -595 780 -594
rect 205 -597 206 -596
rect 219 -597 220 -596
rect 226 -597 227 -596
rect 527 -597 528 -596
rect 534 -597 535 -596
rect 653 -597 654 -596
rect 212 -599 213 -598
rect 282 -599 283 -598
rect 289 -599 290 -598
rect 443 -599 444 -598
rect 471 -599 472 -598
rect 590 -599 591 -598
rect 632 -599 633 -598
rect 667 -599 668 -598
rect 16 -601 17 -600
rect 212 -601 213 -600
rect 215 -601 216 -600
rect 345 -601 346 -600
rect 359 -601 360 -600
rect 485 -601 486 -600
rect 513 -601 514 -600
rect 544 -601 545 -600
rect 569 -601 570 -600
rect 737 -601 738 -600
rect 16 -603 17 -602
rect 61 -603 62 -602
rect 219 -603 220 -602
rect 233 -603 234 -602
rect 236 -603 237 -602
rect 422 -603 423 -602
rect 425 -603 426 -602
rect 667 -603 668 -602
rect 114 -605 115 -604
rect 422 -605 423 -604
rect 590 -605 591 -604
rect 674 -605 675 -604
rect 114 -607 115 -606
rect 170 -607 171 -606
rect 226 -607 227 -606
rect 268 -607 269 -606
rect 275 -607 276 -606
rect 296 -607 297 -606
rect 359 -607 360 -606
rect 366 -607 367 -606
rect 380 -607 381 -606
rect 569 -607 570 -606
rect 639 -607 640 -606
rect 702 -607 703 -606
rect 149 -609 150 -608
rect 233 -609 234 -608
rect 247 -609 248 -608
rect 268 -609 269 -608
rect 275 -609 276 -608
rect 499 -609 500 -608
rect 611 -609 612 -608
rect 639 -609 640 -608
rect 149 -611 150 -610
rect 324 -611 325 -610
rect 338 -611 339 -610
rect 380 -611 381 -610
rect 467 -611 468 -610
rect 499 -611 500 -610
rect 611 -611 612 -610
rect 716 -611 717 -610
rect 145 -613 146 -612
rect 324 -613 325 -612
rect 366 -613 367 -612
rect 394 -613 395 -612
rect 492 -613 493 -612
rect 674 -613 675 -612
rect 709 -613 710 -612
rect 716 -613 717 -612
rect 247 -615 248 -614
rect 387 -615 388 -614
rect 450 -615 451 -614
rect 709 -615 710 -614
rect 72 -617 73 -616
rect 387 -617 388 -616
rect 72 -619 73 -618
rect 310 -619 311 -618
rect 334 -619 335 -618
rect 492 -619 493 -618
rect 282 -621 283 -620
rect 303 -621 304 -620
rect 352 -621 353 -620
rect 394 -621 395 -620
rect 289 -623 290 -622
rect 408 -623 409 -622
rect 68 -625 69 -624
rect 408 -625 409 -624
rect 352 -627 353 -626
rect 464 -627 465 -626
rect 464 -629 465 -628
rect 821 -629 822 -628
rect 593 -631 594 -630
rect 821 -631 822 -630
rect 2 -642 3 -641
rect 58 -642 59 -641
rect 61 -642 62 -641
rect 135 -642 136 -641
rect 138 -642 139 -641
rect 453 -642 454 -641
rect 464 -642 465 -641
rect 723 -642 724 -641
rect 821 -642 822 -641
rect 954 -642 955 -641
rect 2 -644 3 -643
rect 156 -644 157 -643
rect 173 -644 174 -643
rect 282 -644 283 -643
rect 289 -644 290 -643
rect 303 -644 304 -643
rect 331 -644 332 -643
rect 569 -644 570 -643
rect 590 -644 591 -643
rect 870 -644 871 -643
rect 947 -644 948 -643
rect 1031 -644 1032 -643
rect 16 -646 17 -645
rect 86 -646 87 -645
rect 93 -646 94 -645
rect 110 -646 111 -645
rect 184 -646 185 -645
rect 411 -646 412 -645
rect 436 -646 437 -645
rect 464 -646 465 -645
rect 488 -646 489 -645
rect 583 -646 584 -645
rect 593 -646 594 -645
rect 905 -646 906 -645
rect 16 -648 17 -647
rect 149 -648 150 -647
rect 184 -648 185 -647
rect 268 -648 269 -647
rect 289 -648 290 -647
rect 394 -648 395 -647
rect 404 -648 405 -647
rect 555 -648 556 -647
rect 562 -648 563 -647
rect 569 -648 570 -647
rect 583 -648 584 -647
rect 632 -648 633 -647
rect 660 -648 661 -647
rect 695 -648 696 -647
rect 793 -648 794 -647
rect 821 -648 822 -647
rect 891 -648 892 -647
rect 905 -648 906 -647
rect 37 -650 38 -649
rect 334 -650 335 -649
rect 338 -650 339 -649
rect 366 -650 367 -649
rect 387 -650 388 -649
rect 450 -650 451 -649
rect 481 -650 482 -649
rect 593 -650 594 -649
rect 604 -650 605 -649
rect 618 -650 619 -649
rect 621 -650 622 -649
rect 758 -650 759 -649
rect 786 -650 787 -649
rect 793 -650 794 -649
rect 814 -650 815 -649
rect 870 -650 871 -649
rect 51 -652 52 -651
rect 471 -652 472 -651
rect 502 -652 503 -651
rect 807 -652 808 -651
rect 828 -652 829 -651
rect 891 -652 892 -651
rect 30 -654 31 -653
rect 471 -654 472 -653
rect 513 -654 514 -653
rect 534 -654 535 -653
rect 537 -654 538 -653
rect 765 -654 766 -653
rect 779 -654 780 -653
rect 786 -654 787 -653
rect 51 -656 52 -655
rect 478 -656 479 -655
rect 520 -656 521 -655
rect 912 -656 913 -655
rect 58 -658 59 -657
rect 177 -658 178 -657
rect 198 -658 199 -657
rect 268 -658 269 -657
rect 338 -658 339 -657
rect 474 -658 475 -657
rect 506 -658 507 -657
rect 520 -658 521 -657
rect 523 -658 524 -657
rect 597 -658 598 -657
rect 611 -658 612 -657
rect 814 -658 815 -657
rect 912 -658 913 -657
rect 926 -658 927 -657
rect 65 -660 66 -659
rect 156 -660 157 -659
rect 177 -660 178 -659
rect 275 -660 276 -659
rect 341 -660 342 -659
rect 373 -660 374 -659
rect 436 -660 437 -659
rect 544 -660 545 -659
rect 551 -660 552 -659
rect 702 -660 703 -659
rect 716 -660 717 -659
rect 779 -660 780 -659
rect 65 -662 66 -661
rect 121 -662 122 -661
rect 149 -662 150 -661
rect 191 -662 192 -661
rect 198 -662 199 -661
rect 219 -662 220 -661
rect 233 -662 234 -661
rect 317 -662 318 -661
rect 345 -662 346 -661
rect 527 -662 528 -661
rect 541 -662 542 -661
rect 709 -662 710 -661
rect 730 -662 731 -661
rect 926 -662 927 -661
rect 72 -664 73 -663
rect 317 -664 318 -663
rect 359 -664 360 -663
rect 394 -664 395 -663
rect 408 -664 409 -663
rect 527 -664 528 -663
rect 541 -664 542 -663
rect 856 -664 857 -663
rect 72 -666 73 -665
rect 443 -666 444 -665
rect 474 -666 475 -665
rect 828 -666 829 -665
rect 79 -668 80 -667
rect 243 -668 244 -667
rect 247 -668 248 -667
rect 282 -668 283 -667
rect 366 -668 367 -667
rect 401 -668 402 -667
rect 443 -668 444 -667
rect 467 -668 468 -667
rect 499 -668 500 -667
rect 506 -668 507 -667
rect 555 -668 556 -667
rect 737 -668 738 -667
rect 765 -668 766 -667
rect 835 -668 836 -667
rect 9 -670 10 -669
rect 243 -670 244 -669
rect 250 -670 251 -669
rect 254 -670 255 -669
rect 275 -670 276 -669
rect 415 -670 416 -669
rect 478 -670 479 -669
rect 737 -670 738 -669
rect 9 -672 10 -671
rect 44 -672 45 -671
rect 79 -672 80 -671
rect 380 -672 381 -671
rect 390 -672 391 -671
rect 835 -672 836 -671
rect 23 -674 24 -673
rect 44 -674 45 -673
rect 86 -674 87 -673
rect 856 -674 857 -673
rect 93 -676 94 -675
rect 145 -676 146 -675
rect 170 -676 171 -675
rect 191 -676 192 -675
rect 205 -676 206 -675
rect 303 -676 304 -675
rect 324 -676 325 -675
rect 401 -676 402 -675
rect 562 -676 563 -675
rect 849 -676 850 -675
rect 100 -678 101 -677
rect 548 -678 549 -677
rect 576 -678 577 -677
rect 604 -678 605 -677
rect 614 -678 615 -677
rect 919 -678 920 -677
rect 103 -680 104 -679
rect 611 -680 612 -679
rect 625 -680 626 -679
rect 632 -680 633 -679
rect 639 -680 640 -679
rect 660 -680 661 -679
rect 667 -680 668 -679
rect 919 -680 920 -679
rect 100 -682 101 -681
rect 667 -682 668 -681
rect 674 -682 675 -681
rect 723 -682 724 -681
rect 730 -682 731 -681
rect 800 -682 801 -681
rect 842 -682 843 -681
rect 849 -682 850 -681
rect 103 -684 104 -683
rect 142 -684 143 -683
rect 170 -684 171 -683
rect 261 -684 262 -683
rect 324 -684 325 -683
rect 429 -684 430 -683
rect 576 -684 577 -683
rect 625 -684 626 -683
rect 639 -684 640 -683
rect 887 -684 888 -683
rect 107 -686 108 -685
rect 128 -686 129 -685
rect 205 -686 206 -685
rect 254 -686 255 -685
rect 261 -686 262 -685
rect 310 -686 311 -685
rect 352 -686 353 -685
rect 415 -686 416 -685
rect 422 -686 423 -685
rect 429 -686 430 -685
rect 646 -686 647 -685
rect 674 -686 675 -685
rect 688 -686 689 -685
rect 758 -686 759 -685
rect 772 -686 773 -685
rect 800 -686 801 -685
rect 842 -686 843 -685
rect 877 -686 878 -685
rect 114 -688 115 -687
rect 310 -688 311 -687
rect 352 -688 353 -687
rect 628 -688 629 -687
rect 653 -688 654 -687
rect 702 -688 703 -687
rect 751 -688 752 -687
rect 772 -688 773 -687
rect 877 -688 878 -687
rect 898 -688 899 -687
rect 89 -690 90 -689
rect 114 -690 115 -689
rect 121 -690 122 -689
rect 163 -690 164 -689
rect 212 -690 213 -689
rect 597 -690 598 -689
rect 744 -690 745 -689
rect 751 -690 752 -689
rect 863 -690 864 -689
rect 898 -690 899 -689
rect 135 -692 136 -691
rect 212 -692 213 -691
rect 219 -692 220 -691
rect 296 -692 297 -691
rect 380 -692 381 -691
rect 457 -692 458 -691
rect 485 -692 486 -691
rect 646 -692 647 -691
rect 681 -692 682 -691
rect 744 -692 745 -691
rect 863 -692 864 -691
rect 884 -692 885 -691
rect 145 -694 146 -693
rect 688 -694 689 -693
rect 163 -696 164 -695
rect 565 -696 566 -695
rect 226 -698 227 -697
rect 408 -698 409 -697
rect 422 -698 423 -697
rect 548 -698 549 -697
rect 558 -698 559 -697
rect 681 -698 682 -697
rect 229 -700 230 -699
rect 457 -700 458 -699
rect 485 -700 486 -699
rect 716 -700 717 -699
rect 236 -702 237 -701
rect 709 -702 710 -701
rect 240 -704 241 -703
rect 359 -704 360 -703
rect 492 -704 493 -703
rect 653 -704 654 -703
rect 240 -706 241 -705
rect 807 -706 808 -705
rect 296 -708 297 -707
rect 418 -708 419 -707
rect 348 -710 349 -709
rect 492 -710 493 -709
rect 16 -721 17 -720
rect 103 -721 104 -720
rect 135 -721 136 -720
rect 390 -721 391 -720
rect 415 -721 416 -720
rect 765 -721 766 -720
rect 849 -721 850 -720
rect 884 -721 885 -720
rect 908 -721 909 -720
rect 912 -721 913 -720
rect 926 -721 927 -720
rect 975 -721 976 -720
rect 1006 -721 1007 -720
rect 1017 -721 1018 -720
rect 1031 -721 1032 -720
rect 1066 -721 1067 -720
rect 23 -723 24 -722
rect 117 -723 118 -722
rect 135 -723 136 -722
rect 149 -723 150 -722
rect 170 -723 171 -722
rect 418 -723 419 -722
rect 478 -723 479 -722
rect 544 -723 545 -722
rect 551 -723 552 -722
rect 856 -723 857 -722
rect 912 -723 913 -722
rect 961 -723 962 -722
rect 26 -725 27 -724
rect 30 -725 31 -724
rect 33 -725 34 -724
rect 670 -725 671 -724
rect 716 -725 717 -724
rect 765 -725 766 -724
rect 793 -725 794 -724
rect 849 -725 850 -724
rect 954 -725 955 -724
rect 1010 -725 1011 -724
rect 30 -727 31 -726
rect 163 -727 164 -726
rect 170 -727 171 -726
rect 187 -727 188 -726
rect 229 -727 230 -726
rect 310 -727 311 -726
rect 317 -727 318 -726
rect 387 -727 388 -726
rect 464 -727 465 -726
rect 478 -727 479 -726
rect 481 -727 482 -726
rect 583 -727 584 -726
rect 590 -727 591 -726
rect 716 -727 717 -726
rect 744 -727 745 -726
rect 793 -727 794 -726
rect 807 -727 808 -726
rect 856 -727 857 -726
rect 44 -729 45 -728
rect 110 -729 111 -728
rect 128 -729 129 -728
rect 387 -729 388 -728
rect 436 -729 437 -728
rect 464 -729 465 -728
rect 488 -729 489 -728
rect 534 -729 535 -728
rect 555 -729 556 -728
rect 835 -729 836 -728
rect 2 -731 3 -730
rect 44 -731 45 -730
rect 58 -731 59 -730
rect 205 -731 206 -730
rect 240 -731 241 -730
rect 541 -731 542 -730
rect 558 -731 559 -730
rect 891 -731 892 -730
rect 58 -733 59 -732
rect 191 -733 192 -732
rect 205 -733 206 -732
rect 233 -733 234 -732
rect 247 -733 248 -732
rect 338 -733 339 -732
rect 348 -733 349 -732
rect 492 -733 493 -732
rect 516 -733 517 -732
rect 653 -733 654 -732
rect 674 -733 675 -732
rect 744 -733 745 -732
rect 779 -733 780 -732
rect 807 -733 808 -732
rect 891 -733 892 -732
rect 915 -733 916 -732
rect 86 -735 87 -734
rect 597 -735 598 -734
rect 621 -735 622 -734
rect 905 -735 906 -734
rect 86 -737 87 -736
rect 282 -737 283 -736
rect 317 -737 318 -736
rect 499 -737 500 -736
rect 506 -737 507 -736
rect 597 -737 598 -736
rect 625 -737 626 -736
rect 898 -737 899 -736
rect 51 -739 52 -738
rect 506 -739 507 -738
rect 527 -739 528 -738
rect 548 -739 549 -738
rect 565 -739 566 -738
rect 800 -739 801 -738
rect 898 -739 899 -738
rect 919 -739 920 -738
rect 65 -741 66 -740
rect 499 -741 500 -740
rect 541 -741 542 -740
rect 674 -741 675 -740
rect 723 -741 724 -740
rect 779 -741 780 -740
rect 814 -741 815 -740
rect 919 -741 920 -740
rect 89 -743 90 -742
rect 667 -743 668 -742
rect 688 -743 689 -742
rect 723 -743 724 -742
rect 737 -743 738 -742
rect 835 -743 836 -742
rect 93 -745 94 -744
rect 243 -745 244 -744
rect 254 -745 255 -744
rect 355 -745 356 -744
rect 373 -745 374 -744
rect 821 -745 822 -744
rect 51 -747 52 -746
rect 93 -747 94 -746
rect 128 -747 129 -746
rect 495 -747 496 -746
rect 569 -747 570 -746
rect 590 -747 591 -746
rect 625 -747 626 -746
rect 639 -747 640 -746
rect 667 -747 668 -746
rect 730 -747 731 -746
rect 758 -747 759 -746
rect 800 -747 801 -746
rect 821 -747 822 -746
rect 828 -747 829 -746
rect 72 -749 73 -748
rect 373 -749 374 -748
rect 394 -749 395 -748
rect 534 -749 535 -748
rect 569 -749 570 -748
rect 576 -749 577 -748
rect 579 -749 580 -748
rect 772 -749 773 -748
rect 142 -751 143 -750
rect 219 -751 220 -750
rect 261 -751 262 -750
rect 264 -751 265 -750
rect 268 -751 269 -750
rect 282 -751 283 -750
rect 331 -751 332 -750
rect 429 -751 430 -750
rect 436 -751 437 -750
rect 457 -751 458 -750
rect 485 -751 486 -750
rect 653 -751 654 -750
rect 660 -751 661 -750
rect 730 -751 731 -750
rect 9 -753 10 -752
rect 457 -753 458 -752
rect 527 -753 528 -752
rect 828 -753 829 -752
rect 107 -755 108 -754
rect 268 -755 269 -754
rect 296 -755 297 -754
rect 429 -755 430 -754
rect 576 -755 577 -754
rect 772 -755 773 -754
rect 107 -757 108 -756
rect 114 -757 115 -756
rect 142 -757 143 -756
rect 352 -757 353 -756
rect 380 -757 381 -756
rect 485 -757 486 -756
rect 583 -757 584 -756
rect 604 -757 605 -756
rect 628 -757 629 -756
rect 870 -757 871 -756
rect 100 -759 101 -758
rect 114 -759 115 -758
rect 145 -759 146 -758
rect 149 -759 150 -758
rect 156 -759 157 -758
rect 163 -759 164 -758
rect 191 -759 192 -758
rect 250 -759 251 -758
rect 254 -759 255 -758
rect 261 -759 262 -758
rect 296 -759 297 -758
rect 345 -759 346 -758
rect 359 -759 360 -758
rect 380 -759 381 -758
rect 394 -759 395 -758
rect 401 -759 402 -758
rect 415 -759 416 -758
rect 814 -759 815 -758
rect 842 -759 843 -758
rect 870 -759 871 -758
rect 100 -761 101 -760
rect 408 -761 409 -760
rect 639 -761 640 -760
rect 646 -761 647 -760
rect 688 -761 689 -760
rect 751 -761 752 -760
rect 786 -761 787 -760
rect 842 -761 843 -760
rect 156 -763 157 -762
rect 198 -763 199 -762
rect 212 -763 213 -762
rect 219 -763 220 -762
rect 236 -763 237 -762
rect 660 -763 661 -762
rect 702 -763 703 -762
rect 737 -763 738 -762
rect 751 -763 752 -762
rect 877 -763 878 -762
rect 37 -765 38 -764
rect 212 -765 213 -764
rect 243 -765 244 -764
rect 359 -765 360 -764
rect 408 -765 409 -764
rect 443 -765 444 -764
rect 450 -765 451 -764
rect 646 -765 647 -764
rect 681 -765 682 -764
rect 702 -765 703 -764
rect 709 -765 710 -764
rect 758 -765 759 -764
rect 863 -765 864 -764
rect 877 -765 878 -764
rect 37 -767 38 -766
rect 513 -767 514 -766
rect 520 -767 521 -766
rect 681 -767 682 -766
rect 695 -767 696 -766
rect 709 -767 710 -766
rect 177 -769 178 -768
rect 198 -769 199 -768
rect 275 -769 276 -768
rect 401 -769 402 -768
rect 404 -769 405 -768
rect 443 -769 444 -768
rect 450 -769 451 -768
rect 530 -769 531 -768
rect 611 -769 612 -768
rect 695 -769 696 -768
rect 79 -771 80 -770
rect 275 -771 276 -770
rect 289 -771 290 -770
rect 520 -771 521 -770
rect 562 -771 563 -770
rect 611 -771 612 -770
rect 632 -771 633 -770
rect 786 -771 787 -770
rect 79 -773 80 -772
rect 376 -773 377 -772
rect 492 -773 493 -772
rect 863 -773 864 -772
rect 177 -775 178 -774
rect 184 -775 185 -774
rect 289 -775 290 -774
rect 303 -775 304 -774
rect 324 -775 325 -774
rect 352 -775 353 -774
rect 513 -775 514 -774
rect 604 -775 605 -774
rect 618 -775 619 -774
rect 632 -775 633 -774
rect 121 -777 122 -776
rect 184 -777 185 -776
rect 310 -777 311 -776
rect 324 -777 325 -776
rect 338 -777 339 -776
rect 366 -777 367 -776
rect 471 -777 472 -776
rect 618 -777 619 -776
rect 110 -779 111 -778
rect 121 -779 122 -778
rect 131 -779 132 -778
rect 303 -779 304 -778
rect 345 -779 346 -778
rect 502 -779 503 -778
rect 366 -781 367 -780
rect 422 -781 423 -780
rect 16 -792 17 -791
rect 65 -792 66 -791
rect 68 -792 69 -791
rect 110 -792 111 -791
rect 114 -792 115 -791
rect 243 -792 244 -791
rect 310 -792 311 -791
rect 369 -792 370 -791
rect 387 -792 388 -791
rect 947 -792 948 -791
rect 961 -792 962 -791
rect 1013 -792 1014 -791
rect 1017 -792 1018 -791
rect 1024 -792 1025 -791
rect 1066 -792 1067 -791
rect 1080 -792 1081 -791
rect 23 -794 24 -793
rect 72 -794 73 -793
rect 79 -794 80 -793
rect 180 -794 181 -793
rect 233 -794 234 -793
rect 303 -794 304 -793
rect 338 -794 339 -793
rect 450 -794 451 -793
rect 492 -794 493 -793
rect 744 -794 745 -793
rect 814 -794 815 -793
rect 954 -794 955 -793
rect 975 -794 976 -793
rect 1017 -794 1018 -793
rect 23 -796 24 -795
rect 149 -796 150 -795
rect 173 -796 174 -795
rect 362 -796 363 -795
rect 411 -796 412 -795
rect 520 -796 521 -795
rect 523 -796 524 -795
rect 849 -796 850 -795
rect 863 -796 864 -795
rect 933 -796 934 -795
rect 989 -796 990 -795
rect 992 -796 993 -795
rect 1010 -796 1011 -795
rect 1038 -796 1039 -795
rect 30 -798 31 -797
rect 313 -798 314 -797
rect 380 -798 381 -797
rect 520 -798 521 -797
rect 530 -798 531 -797
rect 639 -798 640 -797
rect 653 -798 654 -797
rect 849 -798 850 -797
rect 877 -798 878 -797
rect 996 -798 997 -797
rect 37 -800 38 -799
rect 184 -800 185 -799
rect 233 -800 234 -799
rect 296 -800 297 -799
rect 380 -800 381 -799
rect 541 -800 542 -799
rect 551 -800 552 -799
rect 653 -800 654 -799
rect 695 -800 696 -799
rect 894 -800 895 -799
rect 915 -800 916 -799
rect 1003 -800 1004 -799
rect 37 -802 38 -801
rect 226 -802 227 -801
rect 240 -802 241 -801
rect 289 -802 290 -801
rect 296 -802 297 -801
rect 576 -802 577 -801
rect 618 -802 619 -801
rect 786 -802 787 -801
rect 817 -802 818 -801
rect 961 -802 962 -801
rect 44 -804 45 -803
rect 236 -804 237 -803
rect 254 -804 255 -803
rect 576 -804 577 -803
rect 621 -804 622 -803
rect 898 -804 899 -803
rect 47 -806 48 -805
rect 261 -806 262 -805
rect 268 -806 269 -805
rect 303 -806 304 -805
rect 422 -806 423 -805
rect 968 -806 969 -805
rect 51 -808 52 -807
rect 229 -808 230 -807
rect 254 -808 255 -807
rect 317 -808 318 -807
rect 422 -808 423 -807
rect 429 -808 430 -807
rect 439 -808 440 -807
rect 912 -808 913 -807
rect 30 -810 31 -809
rect 229 -810 230 -809
rect 261 -810 262 -809
rect 527 -810 528 -809
rect 537 -810 538 -809
rect 751 -810 752 -809
rect 800 -810 801 -809
rect 898 -810 899 -809
rect 58 -812 59 -811
rect 352 -812 353 -811
rect 429 -812 430 -811
rect 737 -812 738 -811
rect 751 -812 752 -811
rect 905 -812 906 -811
rect 12 -814 13 -813
rect 58 -814 59 -813
rect 72 -814 73 -813
rect 142 -814 143 -813
rect 149 -814 150 -813
rect 219 -814 220 -813
rect 282 -814 283 -813
rect 352 -814 353 -813
rect 450 -814 451 -813
rect 478 -814 479 -813
rect 485 -814 486 -813
rect 527 -814 528 -813
rect 544 -814 545 -813
rect 618 -814 619 -813
rect 639 -814 640 -813
rect 989 -814 990 -813
rect 79 -816 80 -815
rect 467 -816 468 -815
rect 471 -816 472 -815
rect 485 -816 486 -815
rect 492 -816 493 -815
rect 744 -816 745 -815
rect 821 -816 822 -815
rect 982 -816 983 -815
rect 86 -818 87 -817
rect 425 -818 426 -817
rect 443 -818 444 -817
rect 471 -818 472 -817
rect 478 -818 479 -817
rect 667 -818 668 -817
rect 681 -818 682 -817
rect 737 -818 738 -817
rect 765 -818 766 -817
rect 821 -818 822 -817
rect 828 -818 829 -817
rect 975 -818 976 -817
rect 86 -820 87 -819
rect 93 -820 94 -819
rect 114 -820 115 -819
rect 408 -820 409 -819
rect 499 -820 500 -819
rect 681 -820 682 -819
rect 695 -820 696 -819
rect 814 -820 815 -819
rect 828 -820 829 -819
rect 884 -820 885 -819
rect 93 -822 94 -821
rect 163 -822 164 -821
rect 184 -822 185 -821
rect 345 -822 346 -821
rect 513 -822 514 -821
rect 590 -822 591 -821
rect 667 -822 668 -821
rect 688 -822 689 -821
rect 716 -822 717 -821
rect 863 -822 864 -821
rect 121 -824 122 -823
rect 401 -824 402 -823
rect 513 -824 514 -823
rect 625 -824 626 -823
rect 723 -824 724 -823
rect 765 -824 766 -823
rect 835 -824 836 -823
rect 940 -824 941 -823
rect 121 -826 122 -825
rect 135 -826 136 -825
rect 138 -826 139 -825
rect 191 -826 192 -825
rect 205 -826 206 -825
rect 282 -826 283 -825
rect 289 -826 290 -825
rect 366 -826 367 -825
rect 373 -826 374 -825
rect 723 -826 724 -825
rect 730 -826 731 -825
rect 908 -826 909 -825
rect 2 -828 3 -827
rect 205 -828 206 -827
rect 219 -828 220 -827
rect 674 -828 675 -827
rect 772 -828 773 -827
rect 835 -828 836 -827
rect 128 -830 129 -829
rect 317 -830 318 -829
rect 345 -830 346 -829
rect 415 -830 416 -829
rect 516 -830 517 -829
rect 632 -830 633 -829
rect 660 -830 661 -829
rect 674 -830 675 -829
rect 772 -830 773 -829
rect 807 -830 808 -829
rect 110 -832 111 -831
rect 660 -832 661 -831
rect 670 -832 671 -831
rect 730 -832 731 -831
rect 758 -832 759 -831
rect 807 -832 808 -831
rect 117 -834 118 -833
rect 632 -834 633 -833
rect 702 -834 703 -833
rect 758 -834 759 -833
rect 131 -836 132 -835
rect 856 -836 857 -835
rect 135 -838 136 -837
rect 877 -838 878 -837
rect 142 -840 143 -839
rect 198 -840 199 -839
rect 240 -840 241 -839
rect 443 -840 444 -839
rect 534 -840 535 -839
rect 716 -840 717 -839
rect 163 -842 164 -841
rect 170 -842 171 -841
rect 191 -842 192 -841
rect 247 -842 248 -841
rect 268 -842 269 -841
rect 408 -842 409 -841
rect 415 -842 416 -841
rect 597 -842 598 -841
rect 604 -842 605 -841
rect 688 -842 689 -841
rect 156 -844 157 -843
rect 247 -844 248 -843
rect 324 -844 325 -843
rect 604 -844 605 -843
rect 611 -844 612 -843
rect 625 -844 626 -843
rect 100 -846 101 -845
rect 324 -846 325 -845
rect 355 -846 356 -845
rect 702 -846 703 -845
rect 100 -848 101 -847
rect 331 -848 332 -847
rect 355 -848 356 -847
rect 870 -848 871 -847
rect 156 -850 157 -849
rect 208 -850 209 -849
rect 331 -850 332 -849
rect 394 -850 395 -849
rect 457 -850 458 -849
rect 597 -850 598 -849
rect 793 -850 794 -849
rect 870 -850 871 -849
rect 170 -852 171 -851
rect 177 -852 178 -851
rect 198 -852 199 -851
rect 212 -852 213 -851
rect 275 -852 276 -851
rect 394 -852 395 -851
rect 457 -852 458 -851
rect 464 -852 465 -851
rect 548 -852 549 -851
rect 793 -852 794 -851
rect 177 -854 178 -853
rect 387 -854 388 -853
rect 464 -854 465 -853
rect 926 -854 927 -853
rect 212 -856 213 -855
rect 800 -856 801 -855
rect 366 -858 367 -857
rect 572 -858 573 -857
rect 579 -858 580 -857
rect 905 -858 906 -857
rect 373 -860 374 -859
rect 534 -860 535 -859
rect 548 -860 549 -859
rect 611 -860 612 -859
rect 555 -862 556 -861
rect 856 -862 857 -861
rect 359 -864 360 -863
rect 555 -864 556 -863
rect 562 -864 563 -863
rect 884 -864 885 -863
rect 275 -866 276 -865
rect 359 -866 360 -865
rect 565 -866 566 -865
rect 786 -866 787 -865
rect 565 -868 566 -867
rect 842 -868 843 -867
rect 583 -870 584 -869
rect 590 -870 591 -869
rect 779 -870 780 -869
rect 842 -870 843 -869
rect 436 -872 437 -871
rect 583 -872 584 -871
rect 436 -874 437 -873
rect 646 -874 647 -873
rect 562 -876 563 -875
rect 779 -876 780 -875
rect 569 -878 570 -877
rect 646 -878 647 -877
rect 16 -889 17 -888
rect 114 -889 115 -888
rect 135 -889 136 -888
rect 331 -889 332 -888
rect 359 -889 360 -888
rect 583 -889 584 -888
rect 600 -889 601 -888
rect 870 -889 871 -888
rect 915 -889 916 -888
rect 919 -889 920 -888
rect 954 -889 955 -888
rect 992 -889 993 -888
rect 1013 -889 1014 -888
rect 1024 -889 1025 -888
rect 1038 -889 1039 -888
rect 1059 -889 1060 -888
rect 1080 -889 1081 -888
rect 1087 -889 1088 -888
rect 16 -891 17 -890
rect 170 -891 171 -890
rect 184 -891 185 -890
rect 355 -891 356 -890
rect 366 -891 367 -890
rect 681 -891 682 -890
rect 814 -891 815 -890
rect 821 -891 822 -890
rect 870 -891 871 -890
rect 996 -891 997 -890
rect 1010 -891 1011 -890
rect 1038 -891 1039 -890
rect 23 -893 24 -892
rect 226 -893 227 -892
rect 243 -893 244 -892
rect 275 -893 276 -892
rect 289 -893 290 -892
rect 331 -893 332 -892
rect 366 -893 367 -892
rect 422 -893 423 -892
rect 429 -893 430 -892
rect 530 -893 531 -892
rect 534 -893 535 -892
rect 779 -893 780 -892
rect 817 -893 818 -892
rect 828 -893 829 -892
rect 961 -893 962 -892
rect 1010 -893 1011 -892
rect 2 -895 3 -894
rect 23 -895 24 -894
rect 51 -895 52 -894
rect 418 -895 419 -894
rect 422 -895 423 -894
rect 523 -895 524 -894
rect 534 -895 535 -894
rect 555 -895 556 -894
rect 569 -895 570 -894
rect 898 -895 899 -894
rect 961 -895 962 -894
rect 968 -895 969 -894
rect 989 -895 990 -894
rect 1017 -895 1018 -894
rect 51 -897 52 -896
rect 149 -897 150 -896
rect 156 -897 157 -896
rect 184 -897 185 -896
rect 205 -897 206 -896
rect 275 -897 276 -896
rect 289 -897 290 -896
rect 352 -897 353 -896
rect 369 -897 370 -896
rect 513 -897 514 -896
rect 520 -897 521 -896
rect 786 -897 787 -896
rect 828 -897 829 -896
rect 849 -897 850 -896
rect 891 -897 892 -896
rect 898 -897 899 -896
rect 968 -897 969 -896
rect 975 -897 976 -896
rect 58 -899 59 -898
rect 215 -899 216 -898
rect 219 -899 220 -898
rect 737 -899 738 -898
rect 765 -899 766 -898
rect 786 -899 787 -898
rect 849 -899 850 -898
rect 884 -899 885 -898
rect 891 -899 892 -898
rect 926 -899 927 -898
rect 58 -901 59 -900
rect 387 -901 388 -900
rect 408 -901 409 -900
rect 450 -901 451 -900
rect 464 -901 465 -900
rect 471 -901 472 -900
rect 474 -901 475 -900
rect 793 -901 794 -900
rect 884 -901 885 -900
rect 933 -901 934 -900
rect 65 -903 66 -902
rect 338 -903 339 -902
rect 352 -903 353 -902
rect 373 -903 374 -902
rect 387 -903 388 -902
rect 394 -903 395 -902
rect 408 -903 409 -902
rect 576 -903 577 -902
rect 628 -903 629 -902
rect 800 -903 801 -902
rect 933 -903 934 -902
rect 940 -903 941 -902
rect 72 -905 73 -904
rect 229 -905 230 -904
rect 278 -905 279 -904
rect 520 -905 521 -904
rect 527 -905 528 -904
rect 576 -905 577 -904
rect 730 -905 731 -904
rect 821 -905 822 -904
rect 72 -907 73 -906
rect 310 -907 311 -906
rect 317 -907 318 -906
rect 492 -907 493 -906
rect 499 -907 500 -906
rect 716 -907 717 -906
rect 737 -907 738 -906
rect 744 -907 745 -906
rect 751 -907 752 -906
rect 793 -907 794 -906
rect 800 -907 801 -906
rect 842 -907 843 -906
rect 93 -909 94 -908
rect 240 -909 241 -908
rect 261 -909 262 -908
rect 317 -909 318 -908
rect 324 -909 325 -908
rect 338 -909 339 -908
rect 345 -909 346 -908
rect 492 -909 493 -908
rect 499 -909 500 -908
rect 506 -909 507 -908
rect 537 -909 538 -908
rect 541 -909 542 -908
rect 548 -909 549 -908
rect 982 -909 983 -908
rect 93 -911 94 -910
rect 597 -911 598 -910
rect 635 -911 636 -910
rect 730 -911 731 -910
rect 765 -911 766 -910
rect 835 -911 836 -910
rect 842 -911 843 -910
rect 856 -911 857 -910
rect 905 -911 906 -910
rect 982 -911 983 -910
rect 107 -913 108 -912
rect 611 -913 612 -912
rect 688 -913 689 -912
rect 716 -913 717 -912
rect 723 -913 724 -912
rect 744 -913 745 -912
rect 779 -913 780 -912
rect 943 -913 944 -912
rect 107 -915 108 -914
rect 240 -915 241 -914
rect 261 -915 262 -914
rect 303 -915 304 -914
rect 310 -915 311 -914
rect 562 -915 563 -914
rect 597 -915 598 -914
rect 667 -915 668 -914
rect 702 -915 703 -914
rect 723 -915 724 -914
rect 856 -915 857 -914
rect 863 -915 864 -914
rect 905 -915 906 -914
rect 912 -915 913 -914
rect 110 -917 111 -916
rect 254 -917 255 -916
rect 285 -917 286 -916
rect 303 -917 304 -916
rect 373 -917 374 -916
rect 572 -917 573 -916
rect 604 -917 605 -916
rect 611 -917 612 -916
rect 653 -917 654 -916
rect 702 -917 703 -916
rect 709 -917 710 -916
rect 751 -917 752 -916
rect 863 -917 864 -916
rect 877 -917 878 -916
rect 912 -917 913 -916
rect 922 -917 923 -916
rect 114 -919 115 -918
rect 191 -919 192 -918
rect 198 -919 199 -918
rect 254 -919 255 -918
rect 411 -919 412 -918
rect 709 -919 710 -918
rect 149 -921 150 -920
rect 163 -921 164 -920
rect 170 -921 171 -920
rect 236 -921 237 -920
rect 429 -921 430 -920
rect 457 -921 458 -920
rect 467 -921 468 -920
rect 646 -921 647 -920
rect 660 -921 661 -920
rect 688 -921 689 -920
rect 30 -923 31 -922
rect 163 -923 164 -922
rect 180 -923 181 -922
rect 324 -923 325 -922
rect 436 -923 437 -922
rect 548 -923 549 -922
rect 551 -923 552 -922
rect 590 -923 591 -922
rect 639 -923 640 -922
rect 646 -923 647 -922
rect 660 -923 661 -922
rect 674 -923 675 -922
rect 30 -925 31 -924
rect 215 -925 216 -924
rect 439 -925 440 -924
rect 929 -925 930 -924
rect 86 -927 87 -926
rect 180 -927 181 -926
rect 191 -927 192 -926
rect 233 -927 234 -926
rect 439 -927 440 -926
rect 506 -927 507 -926
rect 513 -927 514 -926
rect 590 -927 591 -926
rect 625 -927 626 -926
rect 674 -927 675 -926
rect 86 -929 87 -928
rect 142 -929 143 -928
rect 156 -929 157 -928
rect 268 -929 269 -928
rect 443 -929 444 -928
rect 569 -929 570 -928
rect 632 -929 633 -928
rect 639 -929 640 -928
rect 37 -931 38 -930
rect 443 -931 444 -930
rect 457 -931 458 -930
rect 485 -931 486 -930
rect 502 -931 503 -930
rect 681 -931 682 -930
rect 37 -933 38 -932
rect 131 -933 132 -932
rect 142 -933 143 -932
rect 296 -933 297 -932
rect 471 -933 472 -932
rect 583 -933 584 -932
rect 173 -935 174 -934
rect 296 -935 297 -934
rect 478 -935 479 -934
rect 485 -935 486 -934
rect 555 -935 556 -934
rect 695 -935 696 -934
rect 198 -937 199 -936
rect 604 -937 605 -936
rect 695 -937 696 -936
rect 1003 -937 1004 -936
rect 208 -939 209 -938
rect 282 -939 283 -938
rect 478 -939 479 -938
rect 877 -939 878 -938
rect 44 -941 45 -940
rect 282 -941 283 -940
rect 562 -941 563 -940
rect 835 -941 836 -940
rect 44 -943 45 -942
rect 401 -943 402 -942
rect 212 -945 213 -944
rect 222 -945 223 -944
rect 233 -945 234 -944
rect 247 -945 248 -944
rect 268 -945 269 -944
rect 380 -945 381 -944
rect 401 -945 402 -944
rect 656 -945 657 -944
rect 100 -947 101 -946
rect 247 -947 248 -946
rect 79 -949 80 -948
rect 100 -949 101 -948
rect 222 -949 223 -948
rect 345 -949 346 -948
rect 79 -951 80 -950
rect 415 -951 416 -950
rect 415 -953 416 -952
rect 758 -953 759 -952
rect 758 -955 759 -954
rect 772 -955 773 -954
rect 618 -957 619 -956
rect 772 -957 773 -956
rect 618 -959 619 -958
rect 954 -959 955 -958
rect 9 -970 10 -969
rect 373 -970 374 -969
rect 380 -970 381 -969
rect 548 -970 549 -969
rect 565 -970 566 -969
rect 821 -970 822 -969
rect 835 -970 836 -969
rect 940 -970 941 -969
rect 947 -970 948 -969
rect 996 -970 997 -969
rect 1010 -970 1011 -969
rect 1031 -970 1032 -969
rect 1038 -970 1039 -969
rect 1073 -970 1074 -969
rect 1087 -970 1088 -969
rect 1094 -970 1095 -969
rect 16 -972 17 -971
rect 471 -972 472 -971
rect 474 -972 475 -971
rect 1076 -972 1077 -971
rect 16 -974 17 -973
rect 366 -974 367 -973
rect 373 -974 374 -973
rect 401 -974 402 -973
rect 408 -974 409 -973
rect 432 -974 433 -973
rect 453 -974 454 -973
rect 464 -974 465 -973
rect 481 -974 482 -973
rect 674 -974 675 -973
rect 698 -974 699 -973
rect 870 -974 871 -973
rect 891 -974 892 -973
rect 1045 -974 1046 -973
rect 1059 -974 1060 -973
rect 1101 -974 1102 -973
rect 37 -976 38 -975
rect 208 -976 209 -975
rect 226 -976 227 -975
rect 586 -976 587 -975
rect 600 -976 601 -975
rect 730 -976 731 -975
rect 751 -976 752 -975
rect 835 -976 836 -975
rect 842 -976 843 -975
rect 947 -976 948 -975
rect 954 -976 955 -975
rect 1087 -976 1088 -975
rect 58 -978 59 -977
rect 474 -978 475 -977
rect 488 -978 489 -977
rect 576 -978 577 -977
rect 607 -978 608 -977
rect 800 -978 801 -977
rect 828 -978 829 -977
rect 842 -978 843 -977
rect 863 -978 864 -977
rect 891 -978 892 -977
rect 898 -978 899 -977
rect 989 -978 990 -977
rect 30 -980 31 -979
rect 607 -980 608 -979
rect 635 -980 636 -979
rect 1010 -980 1011 -979
rect 30 -982 31 -981
rect 198 -982 199 -981
rect 240 -982 241 -981
rect 632 -982 633 -981
rect 639 -982 640 -981
rect 674 -982 675 -981
rect 681 -982 682 -981
rect 751 -982 752 -981
rect 758 -982 759 -981
rect 912 -982 913 -981
rect 919 -982 920 -981
rect 968 -982 969 -981
rect 982 -982 983 -981
rect 1069 -982 1070 -981
rect 61 -984 62 -983
rect 632 -984 633 -983
rect 653 -984 654 -983
rect 884 -984 885 -983
rect 905 -984 906 -983
rect 1038 -984 1039 -983
rect 93 -986 94 -985
rect 243 -986 244 -985
rect 247 -986 248 -985
rect 464 -986 465 -985
rect 471 -986 472 -985
rect 954 -986 955 -985
rect 100 -988 101 -987
rect 327 -988 328 -987
rect 338 -988 339 -987
rect 411 -988 412 -987
rect 418 -988 419 -987
rect 733 -988 734 -987
rect 737 -988 738 -987
rect 828 -988 829 -987
rect 856 -988 857 -987
rect 968 -988 969 -987
rect 100 -990 101 -989
rect 219 -990 220 -989
rect 247 -990 248 -989
rect 345 -990 346 -989
rect 366 -990 367 -989
rect 457 -990 458 -989
rect 492 -990 493 -989
rect 688 -990 689 -989
rect 716 -990 717 -989
rect 758 -990 759 -989
rect 765 -990 766 -989
rect 821 -990 822 -989
rect 905 -990 906 -989
rect 915 -990 916 -989
rect 929 -990 930 -989
rect 961 -990 962 -989
rect 93 -992 94 -991
rect 492 -992 493 -991
rect 495 -992 496 -991
rect 1017 -992 1018 -991
rect 114 -994 115 -993
rect 212 -994 213 -993
rect 261 -994 262 -993
rect 345 -994 346 -993
rect 380 -994 381 -993
rect 485 -994 486 -993
rect 506 -994 507 -993
rect 681 -994 682 -993
rect 730 -994 731 -993
rect 863 -994 864 -993
rect 933 -994 934 -993
rect 982 -994 983 -993
rect 114 -996 115 -995
rect 149 -996 150 -995
rect 177 -996 178 -995
rect 355 -996 356 -995
rect 383 -996 384 -995
rect 401 -996 402 -995
rect 436 -996 437 -995
rect 765 -996 766 -995
rect 793 -996 794 -995
rect 800 -996 801 -995
rect 814 -996 815 -995
rect 884 -996 885 -995
rect 943 -996 944 -995
rect 1059 -996 1060 -995
rect 121 -998 122 -997
rect 128 -998 129 -997
rect 131 -998 132 -997
rect 975 -998 976 -997
rect 72 -1000 73 -999
rect 121 -1000 122 -999
rect 131 -1000 132 -999
rect 226 -1000 227 -999
rect 261 -1000 262 -999
rect 422 -1000 423 -999
rect 457 -1000 458 -999
rect 541 -1000 542 -999
rect 548 -1000 549 -999
rect 870 -1000 871 -999
rect 65 -1002 66 -1001
rect 422 -1002 423 -1001
rect 506 -1002 507 -1001
rect 649 -1002 650 -1001
rect 660 -1002 661 -1001
rect 737 -1002 738 -1001
rect 786 -1002 787 -1001
rect 793 -1002 794 -1001
rect 814 -1002 815 -1001
rect 1066 -1002 1067 -1001
rect 65 -1004 66 -1003
rect 156 -1004 157 -1003
rect 180 -1004 181 -1003
rect 240 -1004 241 -1003
rect 282 -1004 283 -1003
rect 562 -1004 563 -1003
rect 576 -1004 577 -1003
rect 1052 -1004 1053 -1003
rect 72 -1006 73 -1005
rect 254 -1006 255 -1005
rect 285 -1006 286 -1005
rect 779 -1006 780 -1005
rect 135 -1008 136 -1007
rect 439 -1008 440 -1007
rect 450 -1008 451 -1007
rect 779 -1008 780 -1007
rect 135 -1010 136 -1009
rect 926 -1010 927 -1009
rect 142 -1012 143 -1011
rect 530 -1012 531 -1011
rect 537 -1012 538 -1011
rect 849 -1012 850 -1011
rect 44 -1014 45 -1013
rect 142 -1014 143 -1013
rect 145 -1014 146 -1013
rect 1003 -1014 1004 -1013
rect 149 -1016 150 -1015
rect 163 -1016 164 -1015
rect 180 -1016 181 -1015
rect 275 -1016 276 -1015
rect 296 -1016 297 -1015
rect 436 -1016 437 -1015
rect 450 -1016 451 -1015
rect 926 -1016 927 -1015
rect 23 -1018 24 -1017
rect 163 -1018 164 -1017
rect 191 -1018 192 -1017
rect 233 -1018 234 -1017
rect 299 -1018 300 -1017
rect 520 -1018 521 -1017
rect 527 -1018 528 -1017
rect 667 -1018 668 -1017
rect 723 -1018 724 -1017
rect 786 -1018 787 -1017
rect 849 -1018 850 -1017
rect 877 -1018 878 -1017
rect 23 -1020 24 -1019
rect 222 -1020 223 -1019
rect 303 -1020 304 -1019
rect 562 -1020 563 -1019
rect 597 -1020 598 -1019
rect 919 -1020 920 -1019
rect 40 -1022 41 -1021
rect 191 -1022 192 -1021
rect 198 -1022 199 -1021
rect 205 -1022 206 -1021
rect 257 -1022 258 -1021
rect 597 -1022 598 -1021
rect 604 -1022 605 -1021
rect 898 -1022 899 -1021
rect 51 -1024 52 -1023
rect 296 -1024 297 -1023
rect 303 -1024 304 -1023
rect 429 -1024 430 -1023
rect 443 -1024 444 -1023
rect 667 -1024 668 -1023
rect 702 -1024 703 -1023
rect 723 -1024 724 -1023
rect 807 -1024 808 -1023
rect 877 -1024 878 -1023
rect 51 -1026 52 -1025
rect 86 -1026 87 -1025
rect 156 -1026 157 -1025
rect 205 -1026 206 -1025
rect 310 -1026 311 -1025
rect 478 -1026 479 -1025
rect 499 -1026 500 -1025
rect 520 -1026 521 -1025
rect 541 -1026 542 -1025
rect 590 -1026 591 -1025
rect 604 -1026 605 -1025
rect 933 -1026 934 -1025
rect 44 -1028 45 -1027
rect 478 -1028 479 -1027
rect 499 -1028 500 -1027
rect 922 -1028 923 -1027
rect 79 -1030 80 -1029
rect 310 -1030 311 -1029
rect 317 -1030 318 -1029
rect 338 -1030 339 -1029
rect 387 -1030 388 -1029
rect 394 -1030 395 -1029
rect 397 -1030 398 -1029
rect 415 -1030 416 -1029
rect 443 -1030 444 -1029
rect 744 -1030 745 -1029
rect 79 -1032 80 -1031
rect 359 -1032 360 -1031
rect 516 -1032 517 -1031
rect 772 -1032 773 -1031
rect 268 -1034 269 -1033
rect 317 -1034 318 -1033
rect 324 -1034 325 -1033
rect 387 -1034 388 -1033
rect 429 -1034 430 -1033
rect 772 -1034 773 -1033
rect 107 -1036 108 -1035
rect 268 -1036 269 -1035
rect 331 -1036 332 -1035
rect 359 -1036 360 -1035
rect 534 -1036 535 -1035
rect 590 -1036 591 -1035
rect 611 -1036 612 -1035
rect 653 -1036 654 -1035
rect 702 -1036 703 -1035
rect 709 -1036 710 -1035
rect 107 -1038 108 -1037
rect 170 -1038 171 -1037
rect 184 -1038 185 -1037
rect 324 -1038 325 -1037
rect 331 -1038 332 -1037
rect 352 -1038 353 -1037
rect 551 -1038 552 -1037
rect 856 -1038 857 -1037
rect 12 -1040 13 -1039
rect 352 -1040 353 -1039
rect 555 -1040 556 -1039
rect 639 -1040 640 -1039
rect 646 -1040 647 -1039
rect 660 -1040 661 -1039
rect 691 -1040 692 -1039
rect 709 -1040 710 -1039
rect 184 -1042 185 -1041
rect 289 -1042 290 -1041
rect 453 -1042 454 -1041
rect 555 -1042 556 -1041
rect 569 -1042 570 -1041
rect 611 -1042 612 -1041
rect 618 -1042 619 -1041
rect 716 -1042 717 -1041
rect 289 -1044 290 -1043
rect 362 -1044 363 -1043
rect 446 -1044 447 -1043
rect 618 -1044 619 -1043
rect 625 -1044 626 -1043
rect 961 -1044 962 -1043
rect 569 -1046 570 -1045
rect 695 -1046 696 -1045
rect 583 -1048 584 -1047
rect 744 -1048 745 -1047
rect 86 -1050 87 -1049
rect 583 -1050 584 -1049
rect 628 -1050 629 -1049
rect 807 -1050 808 -1049
rect 646 -1052 647 -1051
rect 695 -1052 696 -1051
rect 16 -1063 17 -1062
rect 450 -1063 451 -1062
rect 478 -1063 479 -1062
rect 828 -1063 829 -1062
rect 961 -1063 962 -1062
rect 1024 -1063 1025 -1062
rect 1027 -1063 1028 -1062
rect 1052 -1063 1053 -1062
rect 1059 -1063 1060 -1062
rect 1083 -1063 1084 -1062
rect 1094 -1063 1095 -1062
rect 1097 -1063 1098 -1062
rect 19 -1065 20 -1064
rect 334 -1065 335 -1064
rect 338 -1065 339 -1064
rect 443 -1065 444 -1064
rect 464 -1065 465 -1064
rect 478 -1065 479 -1064
rect 495 -1065 496 -1064
rect 877 -1065 878 -1064
rect 989 -1065 990 -1064
rect 1059 -1065 1060 -1064
rect 1094 -1065 1095 -1064
rect 1101 -1065 1102 -1064
rect 30 -1067 31 -1066
rect 37 -1067 38 -1066
rect 51 -1067 52 -1066
rect 58 -1067 59 -1066
rect 65 -1067 66 -1066
rect 145 -1067 146 -1066
rect 156 -1067 157 -1066
rect 180 -1067 181 -1066
rect 191 -1067 192 -1066
rect 194 -1067 195 -1066
rect 219 -1067 220 -1066
rect 229 -1067 230 -1066
rect 275 -1067 276 -1066
rect 548 -1067 549 -1066
rect 569 -1067 570 -1066
rect 898 -1067 899 -1066
rect 996 -1067 997 -1066
rect 1052 -1067 1053 -1066
rect 51 -1069 52 -1068
rect 131 -1069 132 -1068
rect 142 -1069 143 -1068
rect 264 -1069 265 -1068
rect 282 -1069 283 -1068
rect 474 -1069 475 -1068
rect 513 -1069 514 -1068
rect 576 -1069 577 -1068
rect 579 -1069 580 -1068
rect 870 -1069 871 -1068
rect 1017 -1069 1018 -1068
rect 1073 -1069 1074 -1068
rect 58 -1071 59 -1070
rect 355 -1071 356 -1070
rect 369 -1071 370 -1070
rect 933 -1071 934 -1070
rect 65 -1073 66 -1072
rect 261 -1073 262 -1072
rect 296 -1073 297 -1072
rect 373 -1073 374 -1072
rect 387 -1073 388 -1072
rect 513 -1073 514 -1072
rect 576 -1073 577 -1072
rect 600 -1073 601 -1072
rect 604 -1073 605 -1072
rect 828 -1073 829 -1072
rect 926 -1073 927 -1072
rect 1017 -1073 1018 -1072
rect 2 -1075 3 -1074
rect 261 -1075 262 -1074
rect 303 -1075 304 -1074
rect 467 -1075 468 -1074
rect 583 -1075 584 -1074
rect 1045 -1075 1046 -1074
rect 79 -1077 80 -1076
rect 187 -1077 188 -1076
rect 191 -1077 192 -1076
rect 212 -1077 213 -1076
rect 222 -1077 223 -1076
rect 345 -1077 346 -1076
rect 352 -1077 353 -1076
rect 940 -1077 941 -1076
rect 114 -1079 115 -1078
rect 173 -1079 174 -1078
rect 177 -1079 178 -1078
rect 198 -1079 199 -1078
rect 233 -1079 234 -1078
rect 275 -1079 276 -1078
rect 310 -1079 311 -1078
rect 495 -1079 496 -1078
rect 569 -1079 570 -1078
rect 583 -1079 584 -1078
rect 586 -1079 587 -1078
rect 912 -1079 913 -1078
rect 940 -1079 941 -1078
rect 1087 -1079 1088 -1078
rect 1097 -1079 1098 -1078
rect 1101 -1079 1102 -1078
rect 93 -1081 94 -1080
rect 114 -1081 115 -1080
rect 121 -1081 122 -1080
rect 254 -1081 255 -1080
rect 317 -1081 318 -1080
rect 443 -1081 444 -1080
rect 572 -1081 573 -1080
rect 1045 -1081 1046 -1080
rect 44 -1083 45 -1082
rect 121 -1083 122 -1082
rect 156 -1083 157 -1082
rect 289 -1083 290 -1082
rect 324 -1083 325 -1082
rect 453 -1083 454 -1082
rect 593 -1083 594 -1082
rect 954 -1083 955 -1082
rect 44 -1085 45 -1084
rect 537 -1085 538 -1084
rect 597 -1085 598 -1084
rect 607 -1085 608 -1084
rect 621 -1085 622 -1084
rect 996 -1085 997 -1084
rect 93 -1087 94 -1086
rect 243 -1087 244 -1086
rect 247 -1087 248 -1086
rect 282 -1087 283 -1086
rect 289 -1087 290 -1086
rect 331 -1087 332 -1086
rect 338 -1087 339 -1086
rect 436 -1087 437 -1086
rect 439 -1087 440 -1086
rect 541 -1087 542 -1086
rect 628 -1087 629 -1086
rect 835 -1087 836 -1086
rect 863 -1087 864 -1086
rect 926 -1087 927 -1086
rect 135 -1089 136 -1088
rect 324 -1089 325 -1088
rect 345 -1089 346 -1088
rect 590 -1089 591 -1088
rect 628 -1089 629 -1088
rect 947 -1089 948 -1088
rect 107 -1091 108 -1090
rect 135 -1091 136 -1090
rect 163 -1091 164 -1090
rect 492 -1091 493 -1090
rect 509 -1091 510 -1090
rect 947 -1091 948 -1090
rect 107 -1093 108 -1092
rect 170 -1093 171 -1092
rect 184 -1093 185 -1092
rect 317 -1093 318 -1092
rect 359 -1093 360 -1092
rect 373 -1093 374 -1092
rect 387 -1093 388 -1092
rect 401 -1093 402 -1092
rect 408 -1093 409 -1092
rect 863 -1093 864 -1092
rect 912 -1093 913 -1092
rect 982 -1093 983 -1092
rect 100 -1095 101 -1094
rect 170 -1095 171 -1094
rect 198 -1095 199 -1094
rect 380 -1095 381 -1094
rect 394 -1095 395 -1094
rect 408 -1095 409 -1094
rect 411 -1095 412 -1094
rect 446 -1095 447 -1094
rect 541 -1095 542 -1094
rect 1069 -1095 1070 -1094
rect 9 -1097 10 -1096
rect 100 -1097 101 -1096
rect 166 -1097 167 -1096
rect 961 -1097 962 -1096
rect 240 -1099 241 -1098
rect 310 -1099 311 -1098
rect 359 -1099 360 -1098
rect 446 -1099 447 -1098
rect 590 -1099 591 -1098
rect 884 -1099 885 -1098
rect 919 -1099 920 -1098
rect 954 -1099 955 -1098
rect 247 -1101 248 -1100
rect 597 -1101 598 -1100
rect 646 -1101 647 -1100
rect 677 -1101 678 -1100
rect 688 -1101 689 -1100
rect 905 -1101 906 -1100
rect 919 -1101 920 -1100
rect 1080 -1101 1081 -1100
rect 380 -1103 381 -1102
rect 506 -1103 507 -1102
rect 649 -1103 650 -1102
rect 968 -1103 969 -1102
rect 1003 -1103 1004 -1102
rect 1080 -1103 1081 -1102
rect 72 -1105 73 -1104
rect 506 -1105 507 -1104
rect 688 -1105 689 -1104
rect 982 -1105 983 -1104
rect 23 -1107 24 -1106
rect 72 -1107 73 -1106
rect 394 -1107 395 -1106
rect 562 -1107 563 -1106
rect 723 -1107 724 -1106
rect 835 -1107 836 -1106
rect 849 -1107 850 -1106
rect 968 -1107 969 -1106
rect 23 -1109 24 -1108
rect 128 -1109 129 -1108
rect 401 -1109 402 -1108
rect 534 -1109 535 -1108
rect 555 -1109 556 -1108
rect 562 -1109 563 -1108
rect 639 -1109 640 -1108
rect 723 -1109 724 -1108
rect 726 -1109 727 -1108
rect 898 -1109 899 -1108
rect 422 -1111 423 -1110
rect 551 -1111 552 -1110
rect 555 -1111 556 -1110
rect 611 -1111 612 -1110
rect 730 -1111 731 -1110
rect 989 -1111 990 -1110
rect 268 -1113 269 -1112
rect 422 -1113 423 -1112
rect 429 -1113 430 -1112
rect 667 -1113 668 -1112
rect 730 -1113 731 -1112
rect 1038 -1113 1039 -1112
rect 429 -1115 430 -1114
rect 527 -1115 528 -1114
rect 611 -1115 612 -1114
rect 632 -1115 633 -1114
rect 667 -1115 668 -1114
rect 751 -1115 752 -1114
rect 765 -1115 766 -1114
rect 849 -1115 850 -1114
rect 856 -1115 857 -1114
rect 905 -1115 906 -1114
rect 1038 -1115 1039 -1114
rect 1076 -1115 1077 -1114
rect 436 -1117 437 -1116
rect 1066 -1117 1067 -1116
rect 457 -1119 458 -1118
rect 646 -1119 647 -1118
rect 779 -1119 780 -1118
rect 870 -1119 871 -1118
rect 457 -1121 458 -1120
rect 499 -1121 500 -1120
rect 520 -1121 521 -1120
rect 534 -1121 535 -1120
rect 618 -1121 619 -1120
rect 751 -1121 752 -1120
rect 786 -1121 787 -1120
rect 1003 -1121 1004 -1120
rect 226 -1123 227 -1122
rect 499 -1123 500 -1122
rect 520 -1123 521 -1122
rect 660 -1123 661 -1122
rect 716 -1123 717 -1122
rect 779 -1123 780 -1122
rect 800 -1123 801 -1122
rect 884 -1123 885 -1122
rect 226 -1125 227 -1124
rect 268 -1125 269 -1124
rect 530 -1125 531 -1124
rect 765 -1125 766 -1124
rect 800 -1125 801 -1124
rect 814 -1125 815 -1124
rect 821 -1125 822 -1124
rect 877 -1125 878 -1124
rect 632 -1127 633 -1126
rect 737 -1127 738 -1126
rect 758 -1127 759 -1126
rect 821 -1127 822 -1126
rect 653 -1129 654 -1128
rect 786 -1129 787 -1128
rect 807 -1129 808 -1128
rect 856 -1129 857 -1128
rect 653 -1131 654 -1130
rect 744 -1131 745 -1130
rect 772 -1131 773 -1130
rect 814 -1131 815 -1130
rect 240 -1133 241 -1132
rect 744 -1133 745 -1132
rect 807 -1133 808 -1132
rect 891 -1133 892 -1132
rect 660 -1135 661 -1134
rect 1010 -1135 1011 -1134
rect 681 -1137 682 -1136
rect 716 -1137 717 -1136
rect 793 -1137 794 -1136
rect 891 -1137 892 -1136
rect 1010 -1137 1011 -1136
rect 1031 -1137 1032 -1136
rect 299 -1139 300 -1138
rect 681 -1139 682 -1138
rect 695 -1139 696 -1138
rect 737 -1139 738 -1138
rect 842 -1139 843 -1138
rect 1031 -1139 1032 -1138
rect 492 -1141 493 -1140
rect 793 -1141 794 -1140
rect 842 -1141 843 -1140
rect 975 -1141 976 -1140
rect 485 -1143 486 -1142
rect 975 -1143 976 -1142
rect 366 -1145 367 -1144
rect 485 -1145 486 -1144
rect 674 -1145 675 -1144
rect 695 -1145 696 -1144
rect 702 -1145 703 -1144
rect 772 -1145 773 -1144
rect 366 -1147 367 -1146
rect 415 -1147 416 -1146
rect 642 -1147 643 -1146
rect 702 -1147 703 -1146
rect 709 -1147 710 -1146
rect 758 -1147 759 -1146
rect 149 -1149 150 -1148
rect 415 -1149 416 -1148
rect 674 -1149 675 -1148
rect 933 -1149 934 -1148
rect 149 -1151 150 -1150
rect 236 -1151 237 -1150
rect 709 -1151 710 -1150
rect 1087 -1151 1088 -1150
rect 30 -1162 31 -1161
rect 586 -1162 587 -1161
rect 590 -1162 591 -1161
rect 621 -1162 622 -1161
rect 639 -1162 640 -1161
rect 891 -1162 892 -1161
rect 1090 -1162 1091 -1161
rect 1101 -1162 1102 -1161
rect 30 -1164 31 -1163
rect 149 -1164 150 -1163
rect 156 -1164 157 -1163
rect 236 -1164 237 -1163
rect 243 -1164 244 -1163
rect 310 -1164 311 -1163
rect 331 -1164 332 -1163
rect 919 -1164 920 -1163
rect 33 -1166 34 -1165
rect 93 -1166 94 -1165
rect 121 -1166 122 -1165
rect 149 -1166 150 -1165
rect 156 -1166 157 -1165
rect 366 -1166 367 -1165
rect 429 -1166 430 -1165
rect 460 -1166 461 -1165
rect 464 -1166 465 -1165
rect 1080 -1166 1081 -1165
rect 51 -1168 52 -1167
rect 366 -1168 367 -1167
rect 436 -1168 437 -1167
rect 1041 -1168 1042 -1167
rect 58 -1170 59 -1169
rect 82 -1170 83 -1169
rect 93 -1170 94 -1169
rect 163 -1170 164 -1169
rect 194 -1170 195 -1169
rect 240 -1170 241 -1169
rect 247 -1170 248 -1169
rect 464 -1170 465 -1169
rect 471 -1170 472 -1169
rect 1024 -1170 1025 -1169
rect 58 -1172 59 -1171
rect 86 -1172 87 -1171
rect 114 -1172 115 -1171
rect 121 -1172 122 -1171
rect 128 -1172 129 -1171
rect 387 -1172 388 -1171
rect 439 -1172 440 -1171
rect 478 -1172 479 -1171
rect 495 -1172 496 -1171
rect 849 -1172 850 -1171
rect 891 -1172 892 -1171
rect 996 -1172 997 -1171
rect 51 -1174 52 -1173
rect 86 -1174 87 -1173
rect 114 -1174 115 -1173
rect 681 -1174 682 -1173
rect 684 -1174 685 -1173
rect 1003 -1174 1004 -1173
rect 82 -1176 83 -1175
rect 100 -1176 101 -1175
rect 128 -1176 129 -1175
rect 135 -1176 136 -1175
rect 163 -1176 164 -1175
rect 954 -1176 955 -1175
rect 135 -1178 136 -1177
rect 212 -1178 213 -1177
rect 226 -1178 227 -1177
rect 625 -1178 626 -1177
rect 639 -1178 640 -1177
rect 772 -1178 773 -1177
rect 842 -1178 843 -1177
rect 1003 -1178 1004 -1177
rect 117 -1180 118 -1179
rect 625 -1180 626 -1179
rect 642 -1180 643 -1179
rect 737 -1180 738 -1179
rect 772 -1180 773 -1179
rect 828 -1180 829 -1179
rect 842 -1180 843 -1179
rect 1087 -1180 1088 -1179
rect 170 -1182 171 -1181
rect 240 -1182 241 -1181
rect 247 -1182 248 -1181
rect 394 -1182 395 -1181
rect 446 -1182 447 -1181
rect 534 -1182 535 -1181
rect 544 -1182 545 -1181
rect 800 -1182 801 -1181
rect 919 -1182 920 -1181
rect 989 -1182 990 -1181
rect 184 -1184 185 -1183
rect 989 -1184 990 -1183
rect 37 -1186 38 -1185
rect 184 -1186 185 -1185
rect 198 -1186 199 -1185
rect 478 -1186 479 -1185
rect 495 -1186 496 -1185
rect 786 -1186 787 -1185
rect 954 -1186 955 -1185
rect 1066 -1186 1067 -1185
rect 37 -1188 38 -1187
rect 166 -1188 167 -1187
rect 226 -1188 227 -1187
rect 317 -1188 318 -1187
rect 331 -1188 332 -1187
rect 345 -1188 346 -1187
rect 352 -1188 353 -1187
rect 373 -1188 374 -1187
rect 380 -1188 381 -1187
rect 436 -1188 437 -1187
rect 450 -1188 451 -1187
rect 527 -1188 528 -1187
rect 548 -1188 549 -1187
rect 551 -1188 552 -1187
rect 590 -1188 591 -1187
rect 996 -1188 997 -1187
rect 79 -1190 80 -1189
rect 345 -1190 346 -1189
rect 380 -1190 381 -1189
rect 401 -1190 402 -1189
rect 450 -1190 451 -1189
rect 485 -1190 486 -1189
rect 509 -1190 510 -1189
rect 1017 -1190 1018 -1189
rect 79 -1192 80 -1191
rect 506 -1192 507 -1191
rect 513 -1192 514 -1191
rect 583 -1192 584 -1191
rect 597 -1192 598 -1191
rect 1031 -1192 1032 -1191
rect 44 -1194 45 -1193
rect 513 -1194 514 -1193
rect 516 -1194 517 -1193
rect 849 -1194 850 -1193
rect 1010 -1194 1011 -1193
rect 1017 -1194 1018 -1193
rect 44 -1196 45 -1195
rect 170 -1196 171 -1195
rect 229 -1196 230 -1195
rect 275 -1196 276 -1195
rect 282 -1196 283 -1195
rect 565 -1196 566 -1195
rect 600 -1196 601 -1195
rect 940 -1196 941 -1195
rect 72 -1198 73 -1197
rect 597 -1198 598 -1197
rect 604 -1198 605 -1197
rect 716 -1198 717 -1197
rect 723 -1198 724 -1197
rect 1052 -1198 1053 -1197
rect 26 -1200 27 -1199
rect 604 -1200 605 -1199
rect 618 -1200 619 -1199
rect 646 -1200 647 -1199
rect 660 -1200 661 -1199
rect 828 -1200 829 -1199
rect 835 -1200 836 -1199
rect 1052 -1200 1053 -1199
rect 72 -1202 73 -1201
rect 324 -1202 325 -1201
rect 387 -1202 388 -1201
rect 569 -1202 570 -1201
rect 618 -1202 619 -1201
rect 628 -1202 629 -1201
rect 660 -1202 661 -1201
rect 695 -1202 696 -1201
rect 716 -1202 717 -1201
rect 884 -1202 885 -1201
rect 912 -1202 913 -1201
rect 1010 -1202 1011 -1201
rect 107 -1204 108 -1203
rect 324 -1204 325 -1203
rect 394 -1204 395 -1203
rect 415 -1204 416 -1203
rect 485 -1204 486 -1203
rect 709 -1204 710 -1203
rect 723 -1204 724 -1203
rect 814 -1204 815 -1203
rect 884 -1204 885 -1203
rect 982 -1204 983 -1203
rect 107 -1206 108 -1205
rect 198 -1206 199 -1205
rect 233 -1206 234 -1205
rect 306 -1206 307 -1205
rect 310 -1206 311 -1205
rect 541 -1206 542 -1205
rect 555 -1206 556 -1205
rect 646 -1206 647 -1205
rect 667 -1206 668 -1205
rect 688 -1206 689 -1205
rect 691 -1206 692 -1205
rect 1024 -1206 1025 -1205
rect 219 -1208 220 -1207
rect 233 -1208 234 -1207
rect 254 -1208 255 -1207
rect 317 -1208 318 -1207
rect 401 -1208 402 -1207
rect 408 -1208 409 -1207
rect 492 -1208 493 -1207
rect 667 -1208 668 -1207
rect 677 -1208 678 -1207
rect 1045 -1208 1046 -1207
rect 16 -1210 17 -1209
rect 254 -1210 255 -1209
rect 261 -1210 262 -1209
rect 548 -1210 549 -1209
rect 555 -1210 556 -1209
rect 576 -1210 577 -1209
rect 586 -1210 587 -1209
rect 912 -1210 913 -1209
rect 1045 -1210 1046 -1209
rect 1073 -1210 1074 -1209
rect 177 -1212 178 -1211
rect 219 -1212 220 -1211
rect 264 -1212 265 -1211
rect 674 -1212 675 -1211
rect 695 -1212 696 -1211
rect 765 -1212 766 -1211
rect 814 -1212 815 -1211
rect 1038 -1212 1039 -1211
rect 1073 -1212 1074 -1211
rect 1094 -1212 1095 -1211
rect 177 -1214 178 -1213
rect 523 -1214 524 -1213
rect 541 -1214 542 -1213
rect 1031 -1214 1032 -1213
rect 1038 -1214 1039 -1213
rect 1066 -1214 1067 -1213
rect 268 -1216 269 -1215
rect 415 -1216 416 -1215
rect 502 -1216 503 -1215
rect 835 -1216 836 -1215
rect 856 -1216 857 -1215
rect 982 -1216 983 -1215
rect 268 -1218 269 -1217
rect 471 -1218 472 -1217
rect 520 -1218 521 -1217
rect 530 -1218 531 -1217
rect 562 -1218 563 -1217
rect 576 -1218 577 -1217
rect 653 -1218 654 -1217
rect 765 -1218 766 -1217
rect 807 -1218 808 -1217
rect 856 -1218 857 -1217
rect 275 -1220 276 -1219
rect 359 -1220 360 -1219
rect 408 -1220 409 -1219
rect 474 -1220 475 -1219
rect 562 -1220 563 -1219
rect 821 -1220 822 -1219
rect 282 -1222 283 -1221
rect 656 -1222 657 -1221
rect 709 -1222 710 -1221
rect 719 -1222 720 -1221
rect 730 -1222 731 -1221
rect 877 -1222 878 -1221
rect 142 -1224 143 -1223
rect 877 -1224 878 -1223
rect 2 -1226 3 -1225
rect 142 -1226 143 -1225
rect 289 -1226 290 -1225
rect 429 -1226 430 -1225
rect 457 -1226 458 -1225
rect 474 -1226 475 -1225
rect 569 -1226 570 -1225
rect 779 -1226 780 -1225
rect 807 -1226 808 -1225
rect 905 -1226 906 -1225
rect 2 -1228 3 -1227
rect 205 -1228 206 -1227
rect 292 -1228 293 -1227
rect 733 -1228 734 -1227
rect 737 -1228 738 -1227
rect 744 -1228 745 -1227
rect 758 -1228 759 -1227
rect 800 -1228 801 -1227
rect 821 -1228 822 -1227
rect 870 -1228 871 -1227
rect 9 -1230 10 -1229
rect 289 -1230 290 -1229
rect 296 -1230 297 -1229
rect 373 -1230 374 -1229
rect 663 -1230 664 -1229
rect 905 -1230 906 -1229
rect 9 -1232 10 -1231
rect 215 -1232 216 -1231
rect 296 -1232 297 -1231
rect 499 -1232 500 -1231
rect 702 -1232 703 -1231
rect 744 -1232 745 -1231
rect 751 -1232 752 -1231
rect 758 -1232 759 -1231
rect 779 -1232 780 -1231
rect 940 -1232 941 -1231
rect 23 -1234 24 -1233
rect 457 -1234 458 -1233
rect 499 -1234 500 -1233
rect 632 -1234 633 -1233
rect 681 -1234 682 -1233
rect 702 -1234 703 -1233
rect 751 -1234 752 -1233
rect 782 -1234 783 -1233
rect 870 -1234 871 -1233
rect 947 -1234 948 -1233
rect 23 -1236 24 -1235
rect 933 -1236 934 -1235
rect 947 -1236 948 -1235
rect 975 -1236 976 -1235
rect 191 -1238 192 -1237
rect 205 -1238 206 -1237
rect 303 -1238 304 -1237
rect 467 -1238 468 -1237
rect 933 -1238 934 -1237
rect 1059 -1238 1060 -1237
rect 100 -1240 101 -1239
rect 191 -1240 192 -1239
rect 338 -1240 339 -1239
rect 359 -1240 360 -1239
rect 422 -1240 423 -1239
rect 632 -1240 633 -1239
rect 793 -1240 794 -1239
rect 1059 -1240 1060 -1239
rect 338 -1242 339 -1241
rect 593 -1242 594 -1241
rect 961 -1242 962 -1241
rect 975 -1242 976 -1241
rect 355 -1244 356 -1243
rect 422 -1244 423 -1243
rect 443 -1244 444 -1243
rect 793 -1244 794 -1243
rect 961 -1244 962 -1243
rect 968 -1244 969 -1243
rect 443 -1246 444 -1245
rect 607 -1246 608 -1245
rect 898 -1246 899 -1245
rect 968 -1246 969 -1245
rect 863 -1248 864 -1247
rect 898 -1248 899 -1247
rect 863 -1250 864 -1249
rect 926 -1250 927 -1249
rect 187 -1252 188 -1251
rect 926 -1252 927 -1251
rect 187 -1254 188 -1253
rect 786 -1254 787 -1253
rect 2 -1265 3 -1264
rect 516 -1265 517 -1264
rect 520 -1265 521 -1264
rect 800 -1265 801 -1264
rect 814 -1265 815 -1264
rect 842 -1265 843 -1264
rect 870 -1265 871 -1264
rect 873 -1265 874 -1264
rect 982 -1265 983 -1264
rect 1062 -1265 1063 -1264
rect 1066 -1265 1067 -1264
rect 1080 -1265 1081 -1264
rect 9 -1267 10 -1266
rect 16 -1267 17 -1266
rect 30 -1267 31 -1266
rect 166 -1267 167 -1266
rect 170 -1267 171 -1266
rect 240 -1267 241 -1266
rect 254 -1267 255 -1266
rect 502 -1267 503 -1266
rect 513 -1267 514 -1266
rect 821 -1267 822 -1266
rect 870 -1267 871 -1266
rect 926 -1267 927 -1266
rect 947 -1267 948 -1266
rect 982 -1267 983 -1266
rect 1017 -1267 1018 -1266
rect 1020 -1267 1021 -1266
rect 9 -1269 10 -1268
rect 58 -1269 59 -1268
rect 86 -1269 87 -1268
rect 590 -1269 591 -1268
rect 604 -1269 605 -1268
rect 779 -1269 780 -1268
rect 912 -1269 913 -1268
rect 947 -1269 948 -1268
rect 1017 -1269 1018 -1268
rect 1052 -1269 1053 -1268
rect 30 -1271 31 -1270
rect 86 -1271 87 -1270
rect 93 -1271 94 -1270
rect 215 -1271 216 -1270
rect 219 -1271 220 -1270
rect 233 -1271 234 -1270
rect 240 -1271 241 -1270
rect 261 -1271 262 -1270
rect 317 -1271 318 -1270
rect 327 -1271 328 -1270
rect 331 -1271 332 -1270
rect 460 -1271 461 -1270
rect 464 -1271 465 -1270
rect 520 -1271 521 -1270
rect 541 -1271 542 -1270
rect 1003 -1271 1004 -1270
rect 1020 -1271 1021 -1270
rect 1052 -1271 1053 -1270
rect 51 -1273 52 -1272
rect 296 -1273 297 -1272
rect 320 -1273 321 -1272
rect 478 -1273 479 -1272
rect 548 -1273 549 -1272
rect 730 -1273 731 -1272
rect 751 -1273 752 -1272
rect 1066 -1273 1067 -1272
rect 51 -1275 52 -1274
rect 149 -1275 150 -1274
rect 159 -1275 160 -1274
rect 471 -1275 472 -1274
rect 478 -1275 479 -1274
rect 695 -1275 696 -1274
rect 761 -1275 762 -1274
rect 821 -1275 822 -1274
rect 884 -1275 885 -1274
rect 912 -1275 913 -1274
rect 1003 -1275 1004 -1274
rect 1034 -1275 1035 -1274
rect 54 -1277 55 -1276
rect 310 -1277 311 -1276
rect 366 -1277 367 -1276
rect 495 -1277 496 -1276
rect 576 -1277 577 -1276
rect 583 -1277 584 -1276
rect 586 -1277 587 -1276
rect 688 -1277 689 -1276
rect 884 -1277 885 -1276
rect 891 -1277 892 -1276
rect 58 -1279 59 -1278
rect 282 -1279 283 -1278
rect 292 -1279 293 -1278
rect 730 -1279 731 -1278
rect 835 -1279 836 -1278
rect 891 -1279 892 -1278
rect 65 -1281 66 -1280
rect 149 -1281 150 -1280
rect 170 -1281 171 -1280
rect 674 -1281 675 -1280
rect 677 -1281 678 -1280
rect 1010 -1281 1011 -1280
rect 65 -1283 66 -1282
rect 338 -1283 339 -1282
rect 369 -1283 370 -1282
rect 527 -1283 528 -1282
rect 555 -1283 556 -1282
rect 576 -1283 577 -1282
rect 583 -1283 584 -1282
rect 632 -1283 633 -1282
rect 639 -1283 640 -1282
rect 695 -1283 696 -1282
rect 817 -1283 818 -1282
rect 835 -1283 836 -1282
rect 954 -1283 955 -1282
rect 1010 -1283 1011 -1282
rect 93 -1285 94 -1284
rect 100 -1285 101 -1284
rect 114 -1285 115 -1284
rect 131 -1285 132 -1284
rect 135 -1285 136 -1284
rect 317 -1285 318 -1284
rect 331 -1285 332 -1284
rect 366 -1285 367 -1284
rect 422 -1285 423 -1284
rect 548 -1285 549 -1284
rect 565 -1285 566 -1284
rect 639 -1285 640 -1284
rect 653 -1285 654 -1284
rect 961 -1285 962 -1284
rect 100 -1287 101 -1286
rect 121 -1287 122 -1286
rect 142 -1287 143 -1286
rect 289 -1287 290 -1286
rect 292 -1287 293 -1286
rect 324 -1287 325 -1286
rect 338 -1287 339 -1286
rect 352 -1287 353 -1286
rect 425 -1287 426 -1286
rect 436 -1287 437 -1286
rect 443 -1287 444 -1286
rect 541 -1287 542 -1286
rect 604 -1287 605 -1286
rect 611 -1287 612 -1286
rect 625 -1287 626 -1286
rect 632 -1287 633 -1286
rect 653 -1287 654 -1286
rect 1059 -1287 1060 -1286
rect 23 -1289 24 -1288
rect 121 -1289 122 -1288
rect 142 -1289 143 -1288
rect 226 -1289 227 -1288
rect 261 -1289 262 -1288
rect 275 -1289 276 -1288
rect 282 -1289 283 -1288
rect 359 -1289 360 -1288
rect 415 -1289 416 -1288
rect 436 -1289 437 -1288
rect 443 -1289 444 -1288
rect 474 -1289 475 -1288
rect 527 -1289 528 -1288
rect 534 -1289 535 -1288
rect 537 -1289 538 -1288
rect 555 -1289 556 -1288
rect 607 -1289 608 -1288
rect 856 -1289 857 -1288
rect 940 -1289 941 -1288
rect 961 -1289 962 -1288
rect 23 -1291 24 -1290
rect 107 -1291 108 -1290
rect 117 -1291 118 -1290
rect 737 -1291 738 -1290
rect 751 -1291 752 -1290
rect 1059 -1291 1060 -1290
rect 72 -1293 73 -1292
rect 352 -1293 353 -1292
rect 359 -1293 360 -1292
rect 765 -1293 766 -1292
rect 793 -1293 794 -1292
rect 856 -1293 857 -1292
rect 919 -1293 920 -1292
rect 940 -1293 941 -1292
rect 72 -1295 73 -1294
rect 387 -1295 388 -1294
rect 464 -1295 465 -1294
rect 506 -1295 507 -1294
rect 537 -1295 538 -1294
rect 646 -1295 647 -1294
rect 656 -1295 657 -1294
rect 989 -1295 990 -1294
rect 107 -1297 108 -1296
rect 138 -1297 139 -1296
rect 163 -1297 164 -1296
rect 625 -1297 626 -1296
rect 660 -1297 661 -1296
rect 842 -1297 843 -1296
rect 849 -1297 850 -1296
rect 919 -1297 920 -1296
rect 968 -1297 969 -1296
rect 989 -1297 990 -1296
rect 117 -1299 118 -1298
rect 310 -1299 311 -1298
rect 373 -1299 374 -1298
rect 387 -1299 388 -1298
rect 611 -1299 612 -1298
rect 618 -1299 619 -1298
rect 660 -1299 661 -1298
rect 702 -1299 703 -1298
rect 716 -1299 717 -1298
rect 765 -1299 766 -1298
rect 793 -1299 794 -1298
rect 1038 -1299 1039 -1298
rect 128 -1301 129 -1300
rect 163 -1301 164 -1300
rect 173 -1301 174 -1300
rect 1024 -1301 1025 -1300
rect 187 -1303 188 -1302
rect 996 -1303 997 -1302
rect 191 -1305 192 -1304
rect 975 -1305 976 -1304
rect 996 -1305 997 -1304
rect 1031 -1305 1032 -1304
rect 194 -1307 195 -1306
rect 247 -1307 248 -1306
rect 268 -1307 269 -1306
rect 646 -1307 647 -1306
rect 667 -1307 668 -1306
rect 800 -1307 801 -1306
rect 807 -1307 808 -1306
rect 954 -1307 955 -1306
rect 194 -1309 195 -1308
rect 254 -1309 255 -1308
rect 268 -1309 269 -1308
rect 345 -1309 346 -1308
rect 373 -1309 374 -1308
rect 485 -1309 486 -1308
rect 667 -1309 668 -1308
rect 1041 -1309 1042 -1308
rect 198 -1311 199 -1310
rect 222 -1311 223 -1310
rect 247 -1311 248 -1310
rect 450 -1311 451 -1310
rect 485 -1311 486 -1310
rect 621 -1311 622 -1310
rect 681 -1311 682 -1310
rect 772 -1311 773 -1310
rect 786 -1311 787 -1310
rect 807 -1311 808 -1310
rect 905 -1311 906 -1310
rect 968 -1311 969 -1310
rect 184 -1313 185 -1312
rect 222 -1313 223 -1312
rect 275 -1313 276 -1312
rect 544 -1313 545 -1312
rect 562 -1313 563 -1312
rect 772 -1313 773 -1312
rect 933 -1313 934 -1312
rect 975 -1313 976 -1312
rect 44 -1315 45 -1314
rect 184 -1315 185 -1314
rect 201 -1315 202 -1314
rect 394 -1315 395 -1314
rect 432 -1315 433 -1314
rect 450 -1315 451 -1314
rect 509 -1315 510 -1314
rect 562 -1315 563 -1314
rect 688 -1315 689 -1314
rect 709 -1315 710 -1314
rect 716 -1315 717 -1314
rect 758 -1315 759 -1314
rect 877 -1315 878 -1314
rect 933 -1315 934 -1314
rect 44 -1317 45 -1316
rect 177 -1317 178 -1316
rect 205 -1317 206 -1316
rect 233 -1317 234 -1316
rect 296 -1317 297 -1316
rect 499 -1317 500 -1316
rect 709 -1317 710 -1316
rect 723 -1317 724 -1316
rect 758 -1317 759 -1316
rect 905 -1317 906 -1316
rect 156 -1319 157 -1318
rect 205 -1319 206 -1318
rect 212 -1319 213 -1318
rect 226 -1319 227 -1318
rect 345 -1319 346 -1318
rect 457 -1319 458 -1318
rect 499 -1319 500 -1318
rect 1048 -1319 1049 -1318
rect 212 -1321 213 -1320
rect 303 -1321 304 -1320
rect 355 -1321 356 -1320
rect 786 -1321 787 -1320
rect 828 -1321 829 -1320
rect 877 -1321 878 -1320
rect 37 -1323 38 -1322
rect 303 -1323 304 -1322
rect 380 -1323 381 -1322
rect 394 -1323 395 -1322
rect 432 -1323 433 -1322
rect 513 -1323 514 -1322
rect 597 -1323 598 -1322
rect 723 -1323 724 -1322
rect 37 -1325 38 -1324
rect 219 -1325 220 -1324
rect 380 -1325 381 -1324
rect 401 -1325 402 -1324
rect 422 -1325 423 -1324
rect 597 -1325 598 -1324
rect 401 -1327 402 -1326
rect 408 -1327 409 -1326
rect 457 -1327 458 -1326
rect 849 -1327 850 -1326
rect 408 -1329 409 -1328
rect 569 -1329 570 -1328
rect 492 -1331 493 -1330
rect 828 -1331 829 -1330
rect 415 -1333 416 -1332
rect 492 -1333 493 -1332
rect 569 -1333 570 -1332
rect 579 -1333 580 -1332
rect 16 -1344 17 -1343
rect 79 -1344 80 -1343
rect 89 -1344 90 -1343
rect 296 -1344 297 -1343
rect 303 -1344 304 -1343
rect 327 -1344 328 -1343
rect 352 -1344 353 -1343
rect 380 -1344 381 -1343
rect 387 -1344 388 -1343
rect 432 -1344 433 -1343
rect 471 -1344 472 -1343
rect 632 -1344 633 -1343
rect 646 -1344 647 -1343
rect 905 -1344 906 -1343
rect 950 -1344 951 -1343
rect 996 -1344 997 -1343
rect 1031 -1344 1032 -1343
rect 1052 -1344 1053 -1343
rect 16 -1346 17 -1345
rect 173 -1346 174 -1345
rect 222 -1346 223 -1345
rect 282 -1346 283 -1345
rect 292 -1346 293 -1345
rect 534 -1346 535 -1345
rect 576 -1346 577 -1345
rect 842 -1346 843 -1345
rect 891 -1346 892 -1345
rect 905 -1346 906 -1345
rect 1024 -1346 1025 -1345
rect 1031 -1346 1032 -1345
rect 1038 -1346 1039 -1345
rect 1073 -1346 1074 -1345
rect 23 -1348 24 -1347
rect 86 -1348 87 -1347
rect 107 -1348 108 -1347
rect 170 -1348 171 -1347
rect 222 -1348 223 -1347
rect 310 -1348 311 -1347
rect 338 -1348 339 -1347
rect 352 -1348 353 -1347
rect 366 -1348 367 -1347
rect 450 -1348 451 -1347
rect 471 -1348 472 -1347
rect 590 -1348 591 -1347
rect 597 -1348 598 -1347
rect 912 -1348 913 -1347
rect 971 -1348 972 -1347
rect 1024 -1348 1025 -1347
rect 1045 -1348 1046 -1347
rect 1048 -1348 1049 -1347
rect 1073 -1348 1074 -1347
rect 1080 -1348 1081 -1347
rect 9 -1350 10 -1349
rect 86 -1350 87 -1349
rect 107 -1350 108 -1349
rect 331 -1350 332 -1349
rect 338 -1350 339 -1349
rect 464 -1350 465 -1349
rect 495 -1350 496 -1349
rect 723 -1350 724 -1349
rect 737 -1350 738 -1349
rect 870 -1350 871 -1349
rect 30 -1352 31 -1351
rect 61 -1352 62 -1351
rect 65 -1352 66 -1351
rect 68 -1352 69 -1351
rect 79 -1352 80 -1351
rect 355 -1352 356 -1351
rect 380 -1352 381 -1351
rect 394 -1352 395 -1351
rect 411 -1352 412 -1351
rect 562 -1352 563 -1351
rect 576 -1352 577 -1351
rect 681 -1352 682 -1351
rect 705 -1352 706 -1351
rect 744 -1352 745 -1351
rect 758 -1352 759 -1351
rect 975 -1352 976 -1351
rect 30 -1354 31 -1353
rect 100 -1354 101 -1353
rect 114 -1354 115 -1353
rect 219 -1354 220 -1353
rect 254 -1354 255 -1353
rect 310 -1354 311 -1353
rect 331 -1354 332 -1353
rect 548 -1354 549 -1353
rect 579 -1354 580 -1353
rect 940 -1354 941 -1353
rect 961 -1354 962 -1353
rect 975 -1354 976 -1353
rect 37 -1356 38 -1355
rect 135 -1356 136 -1355
rect 138 -1356 139 -1355
rect 401 -1356 402 -1355
rect 415 -1356 416 -1355
rect 457 -1356 458 -1355
rect 506 -1356 507 -1355
rect 688 -1356 689 -1355
rect 705 -1356 706 -1355
rect 1017 -1356 1018 -1355
rect 37 -1358 38 -1357
rect 44 -1358 45 -1357
rect 51 -1358 52 -1357
rect 177 -1358 178 -1357
rect 254 -1358 255 -1357
rect 506 -1358 507 -1357
rect 509 -1358 510 -1357
rect 695 -1358 696 -1357
rect 723 -1358 724 -1357
rect 786 -1358 787 -1357
rect 835 -1358 836 -1357
rect 891 -1358 892 -1357
rect 44 -1360 45 -1359
rect 345 -1360 346 -1359
rect 401 -1360 402 -1359
rect 569 -1360 570 -1359
rect 590 -1360 591 -1359
rect 604 -1360 605 -1359
rect 618 -1360 619 -1359
rect 968 -1360 969 -1359
rect 54 -1362 55 -1361
rect 600 -1362 601 -1361
rect 611 -1362 612 -1361
rect 618 -1362 619 -1361
rect 632 -1362 633 -1361
rect 751 -1362 752 -1361
rect 758 -1362 759 -1361
rect 779 -1362 780 -1361
rect 835 -1362 836 -1361
rect 856 -1362 857 -1361
rect 863 -1362 864 -1361
rect 961 -1362 962 -1361
rect 65 -1364 66 -1363
rect 93 -1364 94 -1363
rect 100 -1364 101 -1363
rect 422 -1364 423 -1363
rect 429 -1364 430 -1363
rect 996 -1364 997 -1363
rect 93 -1366 94 -1365
rect 478 -1366 479 -1365
rect 523 -1366 524 -1365
rect 604 -1366 605 -1365
rect 611 -1366 612 -1365
rect 674 -1366 675 -1365
rect 684 -1366 685 -1365
rect 940 -1366 941 -1365
rect 121 -1368 122 -1367
rect 194 -1368 195 -1367
rect 247 -1368 248 -1367
rect 345 -1368 346 -1367
rect 355 -1368 356 -1367
rect 422 -1368 423 -1367
rect 429 -1368 430 -1367
rect 516 -1368 517 -1367
rect 548 -1368 549 -1367
rect 677 -1368 678 -1367
rect 688 -1368 689 -1367
rect 702 -1368 703 -1367
rect 709 -1368 710 -1367
rect 786 -1368 787 -1367
rect 842 -1368 843 -1367
rect 898 -1368 899 -1367
rect 58 -1370 59 -1369
rect 121 -1370 122 -1369
rect 128 -1370 129 -1369
rect 513 -1370 514 -1369
rect 572 -1370 573 -1369
rect 751 -1370 752 -1369
rect 765 -1370 766 -1369
rect 1052 -1370 1053 -1369
rect 128 -1372 129 -1371
rect 208 -1372 209 -1371
rect 268 -1372 269 -1371
rect 296 -1372 297 -1371
rect 303 -1372 304 -1371
rect 709 -1372 710 -1371
rect 730 -1372 731 -1371
rect 744 -1372 745 -1371
rect 779 -1372 780 -1371
rect 800 -1372 801 -1371
rect 849 -1372 850 -1371
rect 912 -1372 913 -1371
rect 145 -1374 146 -1373
rect 156 -1374 157 -1373
rect 159 -1374 160 -1373
rect 541 -1374 542 -1373
rect 579 -1374 580 -1373
rect 863 -1374 864 -1373
rect 870 -1374 871 -1373
rect 877 -1374 878 -1373
rect 884 -1374 885 -1373
rect 898 -1374 899 -1373
rect 149 -1376 150 -1375
rect 268 -1376 269 -1375
rect 275 -1376 276 -1375
rect 394 -1376 395 -1375
rect 415 -1376 416 -1375
rect 663 -1376 664 -1375
rect 674 -1376 675 -1375
rect 716 -1376 717 -1375
rect 737 -1376 738 -1375
rect 772 -1376 773 -1375
rect 800 -1376 801 -1375
rect 807 -1376 808 -1375
rect 884 -1376 885 -1375
rect 982 -1376 983 -1375
rect 149 -1378 150 -1377
rect 180 -1378 181 -1377
rect 184 -1378 185 -1377
rect 247 -1378 248 -1377
rect 261 -1378 262 -1377
rect 275 -1378 276 -1377
rect 282 -1378 283 -1377
rect 387 -1378 388 -1377
rect 450 -1378 451 -1377
rect 499 -1378 500 -1377
rect 583 -1378 584 -1377
rect 856 -1378 857 -1377
rect 982 -1378 983 -1377
rect 989 -1378 990 -1377
rect 163 -1380 164 -1379
rect 191 -1380 192 -1379
rect 205 -1380 206 -1379
rect 261 -1380 262 -1379
rect 324 -1380 325 -1379
rect 478 -1380 479 -1379
rect 492 -1380 493 -1379
rect 807 -1380 808 -1379
rect 23 -1382 24 -1381
rect 205 -1382 206 -1381
rect 324 -1382 325 -1381
rect 373 -1382 374 -1381
rect 443 -1382 444 -1381
rect 499 -1382 500 -1381
rect 583 -1382 584 -1381
rect 954 -1382 955 -1381
rect 68 -1384 69 -1383
rect 373 -1384 374 -1383
rect 443 -1384 444 -1383
rect 485 -1384 486 -1383
rect 492 -1384 493 -1383
rect 520 -1384 521 -1383
rect 586 -1384 587 -1383
rect 989 -1384 990 -1383
rect 163 -1386 164 -1385
rect 289 -1386 290 -1385
rect 359 -1386 360 -1385
rect 730 -1386 731 -1385
rect 772 -1386 773 -1385
rect 828 -1386 829 -1385
rect 947 -1386 948 -1385
rect 954 -1386 955 -1385
rect 177 -1388 178 -1387
rect 198 -1388 199 -1387
rect 359 -1388 360 -1387
rect 436 -1388 437 -1387
rect 464 -1388 465 -1387
rect 569 -1388 570 -1387
rect 597 -1388 598 -1387
rect 1066 -1388 1067 -1387
rect 184 -1390 185 -1389
rect 317 -1390 318 -1389
rect 369 -1390 370 -1389
rect 849 -1390 850 -1389
rect 198 -1392 199 -1391
rect 233 -1392 234 -1391
rect 317 -1392 318 -1391
rect 460 -1392 461 -1391
rect 485 -1392 486 -1391
rect 555 -1392 556 -1391
rect 565 -1392 566 -1391
rect 828 -1392 829 -1391
rect 72 -1394 73 -1393
rect 555 -1394 556 -1393
rect 646 -1394 647 -1393
rect 653 -1394 654 -1393
rect 660 -1394 661 -1393
rect 716 -1394 717 -1393
rect 72 -1396 73 -1395
rect 226 -1396 227 -1395
rect 408 -1396 409 -1395
rect 520 -1396 521 -1395
rect 653 -1396 654 -1395
rect 1034 -1396 1035 -1395
rect 142 -1398 143 -1397
rect 226 -1398 227 -1397
rect 408 -1398 409 -1397
rect 541 -1398 542 -1397
rect 660 -1398 661 -1397
rect 1010 -1398 1011 -1397
rect 212 -1400 213 -1399
rect 233 -1400 234 -1399
rect 436 -1400 437 -1399
rect 527 -1400 528 -1399
rect 681 -1400 682 -1399
rect 877 -1400 878 -1399
rect 1003 -1400 1004 -1399
rect 1010 -1400 1011 -1399
rect 212 -1402 213 -1401
rect 240 -1402 241 -1401
rect 527 -1402 528 -1401
rect 625 -1402 626 -1401
rect 695 -1402 696 -1401
rect 814 -1402 815 -1401
rect 1003 -1402 1004 -1401
rect 1017 -1402 1018 -1401
rect 625 -1404 626 -1403
rect 667 -1404 668 -1403
rect 814 -1404 815 -1403
rect 933 -1404 934 -1403
rect 639 -1406 640 -1405
rect 667 -1406 668 -1405
rect 926 -1406 927 -1405
rect 933 -1406 934 -1405
rect 639 -1408 640 -1407
rect 793 -1408 794 -1407
rect 649 -1410 650 -1409
rect 793 -1410 794 -1409
rect 16 -1421 17 -1420
rect 124 -1421 125 -1420
rect 135 -1421 136 -1420
rect 296 -1421 297 -1420
rect 310 -1421 311 -1420
rect 359 -1421 360 -1420
rect 390 -1421 391 -1420
rect 450 -1421 451 -1420
rect 471 -1421 472 -1420
rect 537 -1421 538 -1420
rect 569 -1421 570 -1420
rect 674 -1421 675 -1420
rect 681 -1421 682 -1420
rect 800 -1421 801 -1420
rect 828 -1421 829 -1420
rect 831 -1421 832 -1420
rect 842 -1421 843 -1420
rect 943 -1421 944 -1420
rect 971 -1421 972 -1420
rect 1031 -1421 1032 -1420
rect 1066 -1421 1067 -1420
rect 1073 -1421 1074 -1420
rect 23 -1423 24 -1422
rect 222 -1423 223 -1422
rect 268 -1423 269 -1422
rect 306 -1423 307 -1422
rect 310 -1423 311 -1422
rect 737 -1423 738 -1422
rect 793 -1423 794 -1422
rect 950 -1423 951 -1422
rect 975 -1423 976 -1422
rect 1003 -1423 1004 -1422
rect 1010 -1423 1011 -1422
rect 1038 -1423 1039 -1422
rect 30 -1425 31 -1424
rect 159 -1425 160 -1424
rect 163 -1425 164 -1424
rect 303 -1425 304 -1424
rect 338 -1425 339 -1424
rect 562 -1425 563 -1424
rect 579 -1425 580 -1424
rect 786 -1425 787 -1424
rect 793 -1425 794 -1424
rect 821 -1425 822 -1424
rect 828 -1425 829 -1424
rect 849 -1425 850 -1424
rect 877 -1425 878 -1424
rect 968 -1425 969 -1424
rect 1024 -1425 1025 -1424
rect 1041 -1425 1042 -1424
rect 30 -1427 31 -1426
rect 51 -1427 52 -1426
rect 54 -1427 55 -1426
rect 128 -1427 129 -1426
rect 138 -1427 139 -1426
rect 142 -1427 143 -1426
rect 163 -1427 164 -1426
rect 212 -1427 213 -1426
rect 219 -1427 220 -1426
rect 653 -1427 654 -1426
rect 663 -1427 664 -1426
rect 779 -1427 780 -1426
rect 821 -1427 822 -1426
rect 905 -1427 906 -1426
rect 929 -1427 930 -1426
rect 961 -1427 962 -1426
rect 44 -1429 45 -1428
rect 128 -1429 129 -1428
rect 142 -1429 143 -1428
rect 170 -1429 171 -1428
rect 205 -1429 206 -1428
rect 891 -1429 892 -1428
rect 44 -1431 45 -1430
rect 187 -1431 188 -1430
rect 205 -1431 206 -1430
rect 240 -1431 241 -1430
rect 289 -1431 290 -1430
rect 471 -1431 472 -1430
rect 499 -1431 500 -1430
rect 513 -1431 514 -1430
rect 516 -1431 517 -1430
rect 716 -1431 717 -1430
rect 744 -1431 745 -1430
rect 975 -1431 976 -1430
rect 58 -1433 59 -1432
rect 684 -1433 685 -1432
rect 688 -1433 689 -1432
rect 716 -1433 717 -1432
rect 723 -1433 724 -1432
rect 744 -1433 745 -1432
rect 772 -1433 773 -1432
rect 786 -1433 787 -1432
rect 835 -1433 836 -1432
rect 849 -1433 850 -1432
rect 877 -1433 878 -1432
rect 926 -1433 927 -1432
rect 72 -1435 73 -1434
rect 401 -1435 402 -1434
rect 408 -1435 409 -1434
rect 520 -1435 521 -1434
rect 523 -1435 524 -1434
rect 625 -1435 626 -1434
rect 635 -1435 636 -1434
rect 807 -1435 808 -1434
rect 835 -1435 836 -1434
rect 870 -1435 871 -1434
rect 884 -1435 885 -1434
rect 922 -1435 923 -1434
rect 926 -1435 927 -1434
rect 954 -1435 955 -1434
rect 37 -1437 38 -1436
rect 72 -1437 73 -1436
rect 75 -1437 76 -1436
rect 296 -1437 297 -1436
rect 338 -1437 339 -1436
rect 586 -1437 587 -1436
rect 597 -1437 598 -1436
rect 688 -1437 689 -1436
rect 712 -1437 713 -1436
rect 814 -1437 815 -1436
rect 842 -1437 843 -1436
rect 940 -1437 941 -1436
rect 954 -1437 955 -1436
rect 1017 -1437 1018 -1436
rect 37 -1439 38 -1438
rect 149 -1439 150 -1438
rect 170 -1439 171 -1438
rect 177 -1439 178 -1438
rect 212 -1439 213 -1438
rect 317 -1439 318 -1438
rect 345 -1439 346 -1438
rect 387 -1439 388 -1438
rect 394 -1439 395 -1438
rect 408 -1439 409 -1438
rect 411 -1439 412 -1438
rect 485 -1439 486 -1438
rect 513 -1439 514 -1438
rect 709 -1439 710 -1438
rect 765 -1439 766 -1438
rect 884 -1439 885 -1438
rect 86 -1441 87 -1440
rect 779 -1441 780 -1440
rect 807 -1441 808 -1440
rect 856 -1441 857 -1440
rect 870 -1441 871 -1440
rect 989 -1441 990 -1440
rect 26 -1443 27 -1442
rect 86 -1443 87 -1442
rect 89 -1443 90 -1442
rect 772 -1443 773 -1442
rect 814 -1443 815 -1442
rect 863 -1443 864 -1442
rect 947 -1443 948 -1442
rect 989 -1443 990 -1442
rect 93 -1445 94 -1444
rect 499 -1445 500 -1444
rect 555 -1445 556 -1444
rect 569 -1445 570 -1444
rect 583 -1445 584 -1444
rect 618 -1445 619 -1444
rect 639 -1445 640 -1444
rect 674 -1445 675 -1444
rect 681 -1445 682 -1444
rect 898 -1445 899 -1444
rect 912 -1445 913 -1444
rect 947 -1445 948 -1444
rect 93 -1447 94 -1446
rect 198 -1447 199 -1446
rect 219 -1447 220 -1446
rect 261 -1447 262 -1446
rect 292 -1447 293 -1446
rect 345 -1447 346 -1446
rect 352 -1447 353 -1446
rect 541 -1447 542 -1446
rect 555 -1447 556 -1446
rect 611 -1447 612 -1446
rect 632 -1447 633 -1446
rect 639 -1447 640 -1446
rect 646 -1447 647 -1446
rect 709 -1447 710 -1446
rect 726 -1447 727 -1446
rect 898 -1447 899 -1446
rect 100 -1449 101 -1448
rect 565 -1449 566 -1448
rect 604 -1449 605 -1448
rect 768 -1449 769 -1448
rect 831 -1449 832 -1448
rect 912 -1449 913 -1448
rect 79 -1451 80 -1450
rect 100 -1451 101 -1450
rect 107 -1451 108 -1450
rect 656 -1451 657 -1450
rect 660 -1451 661 -1450
rect 891 -1451 892 -1450
rect 79 -1453 80 -1452
rect 324 -1453 325 -1452
rect 362 -1453 363 -1452
rect 597 -1453 598 -1452
rect 611 -1453 612 -1452
rect 730 -1453 731 -1452
rect 751 -1453 752 -1452
rect 765 -1453 766 -1452
rect 856 -1453 857 -1452
rect 919 -1453 920 -1452
rect 107 -1455 108 -1454
rect 576 -1455 577 -1454
rect 667 -1455 668 -1454
rect 730 -1455 731 -1454
rect 863 -1455 864 -1454
rect 933 -1455 934 -1454
rect 121 -1457 122 -1456
rect 243 -1457 244 -1456
rect 247 -1457 248 -1456
rect 324 -1457 325 -1456
rect 397 -1457 398 -1456
rect 1052 -1457 1053 -1456
rect 121 -1459 122 -1458
rect 268 -1459 269 -1458
rect 317 -1459 318 -1458
rect 415 -1459 416 -1458
rect 418 -1459 419 -1458
rect 457 -1459 458 -1458
rect 478 -1459 479 -1458
rect 604 -1459 605 -1458
rect 702 -1459 703 -1458
rect 751 -1459 752 -1458
rect 919 -1459 920 -1458
rect 1045 -1459 1046 -1458
rect 149 -1461 150 -1460
rect 429 -1461 430 -1460
rect 450 -1461 451 -1460
rect 464 -1461 465 -1460
rect 478 -1461 479 -1460
rect 590 -1461 591 -1460
rect 695 -1461 696 -1460
rect 702 -1461 703 -1460
rect 933 -1461 934 -1460
rect 996 -1461 997 -1460
rect 166 -1463 167 -1462
rect 583 -1463 584 -1462
rect 590 -1463 591 -1462
rect 1006 -1463 1007 -1462
rect 177 -1465 178 -1464
rect 191 -1465 192 -1464
rect 198 -1465 199 -1464
rect 394 -1465 395 -1464
rect 401 -1465 402 -1464
rect 558 -1465 559 -1464
rect 562 -1465 563 -1464
rect 667 -1465 668 -1464
rect 695 -1465 696 -1464
rect 940 -1465 941 -1464
rect 982 -1465 983 -1464
rect 996 -1465 997 -1464
rect 184 -1467 185 -1466
rect 261 -1467 262 -1466
rect 366 -1467 367 -1466
rect 429 -1467 430 -1466
rect 457 -1467 458 -1466
rect 534 -1467 535 -1466
rect 618 -1467 619 -1466
rect 982 -1467 983 -1466
rect 184 -1469 185 -1468
rect 331 -1469 332 -1468
rect 366 -1469 367 -1468
rect 373 -1469 374 -1468
rect 415 -1469 416 -1468
rect 625 -1469 626 -1468
rect 191 -1471 192 -1470
rect 506 -1471 507 -1470
rect 527 -1471 528 -1470
rect 646 -1471 647 -1470
rect 243 -1473 244 -1472
rect 660 -1473 661 -1472
rect 247 -1475 248 -1474
rect 306 -1475 307 -1474
rect 320 -1475 321 -1474
rect 331 -1475 332 -1474
rect 355 -1475 356 -1474
rect 373 -1475 374 -1474
rect 443 -1475 444 -1474
rect 527 -1475 528 -1474
rect 51 -1477 52 -1476
rect 443 -1477 444 -1476
rect 464 -1477 465 -1476
rect 492 -1477 493 -1476
rect 506 -1477 507 -1476
rect 548 -1477 549 -1476
rect 254 -1479 255 -1478
rect 289 -1479 290 -1478
rect 422 -1479 423 -1478
rect 492 -1479 493 -1478
rect 548 -1479 549 -1478
rect 971 -1479 972 -1478
rect 233 -1481 234 -1480
rect 254 -1481 255 -1480
rect 422 -1481 423 -1480
rect 436 -1481 437 -1480
rect 485 -1481 486 -1480
rect 544 -1481 545 -1480
rect 114 -1483 115 -1482
rect 233 -1483 234 -1482
rect 436 -1483 437 -1482
rect 905 -1483 906 -1482
rect 114 -1485 115 -1484
rect 282 -1485 283 -1484
rect 275 -1487 276 -1486
rect 282 -1487 283 -1486
rect 226 -1489 227 -1488
rect 275 -1489 276 -1488
rect 156 -1491 157 -1490
rect 226 -1491 227 -1490
rect 9 -1502 10 -1501
rect 401 -1502 402 -1501
rect 418 -1502 419 -1501
rect 492 -1502 493 -1501
rect 506 -1502 507 -1501
rect 544 -1502 545 -1501
rect 558 -1502 559 -1501
rect 765 -1502 766 -1501
rect 800 -1502 801 -1501
rect 835 -1502 836 -1501
rect 856 -1502 857 -1501
rect 968 -1502 969 -1501
rect 1038 -1502 1039 -1501
rect 1073 -1502 1074 -1501
rect 16 -1504 17 -1503
rect 149 -1504 150 -1503
rect 194 -1504 195 -1503
rect 499 -1504 500 -1503
rect 506 -1504 507 -1503
rect 712 -1504 713 -1503
rect 726 -1504 727 -1503
rect 807 -1504 808 -1503
rect 835 -1504 836 -1503
rect 1111 -1504 1112 -1503
rect 23 -1506 24 -1505
rect 163 -1506 164 -1505
rect 226 -1506 227 -1505
rect 359 -1506 360 -1505
rect 394 -1506 395 -1505
rect 1101 -1506 1102 -1505
rect 30 -1508 31 -1507
rect 243 -1508 244 -1507
rect 268 -1508 269 -1507
rect 317 -1508 318 -1507
rect 327 -1508 328 -1507
rect 625 -1508 626 -1507
rect 667 -1508 668 -1507
rect 765 -1508 766 -1507
rect 870 -1508 871 -1507
rect 1066 -1508 1067 -1507
rect 30 -1510 31 -1509
rect 142 -1510 143 -1509
rect 149 -1510 150 -1509
rect 397 -1510 398 -1509
rect 418 -1510 419 -1509
rect 520 -1510 521 -1509
rect 534 -1510 535 -1509
rect 807 -1510 808 -1509
rect 870 -1510 871 -1509
rect 982 -1510 983 -1509
rect 1003 -1510 1004 -1509
rect 1038 -1510 1039 -1509
rect 37 -1512 38 -1511
rect 240 -1512 241 -1511
rect 268 -1512 269 -1511
rect 324 -1512 325 -1511
rect 341 -1512 342 -1511
rect 828 -1512 829 -1511
rect 842 -1512 843 -1511
rect 1003 -1512 1004 -1511
rect 37 -1514 38 -1513
rect 656 -1514 657 -1513
rect 681 -1514 682 -1513
rect 884 -1514 885 -1513
rect 891 -1514 892 -1513
rect 1108 -1514 1109 -1513
rect 51 -1516 52 -1515
rect 100 -1516 101 -1515
rect 121 -1516 122 -1515
rect 940 -1516 941 -1515
rect 947 -1516 948 -1515
rect 971 -1516 972 -1515
rect 58 -1518 59 -1517
rect 124 -1518 125 -1517
rect 128 -1518 129 -1517
rect 156 -1518 157 -1517
rect 163 -1518 164 -1517
rect 212 -1518 213 -1517
rect 229 -1518 230 -1517
rect 261 -1518 262 -1517
rect 275 -1518 276 -1517
rect 303 -1518 304 -1517
rect 317 -1518 318 -1517
rect 478 -1518 479 -1517
rect 513 -1518 514 -1517
rect 555 -1518 556 -1517
rect 562 -1518 563 -1517
rect 702 -1518 703 -1517
rect 733 -1518 734 -1517
rect 1080 -1518 1081 -1517
rect 58 -1520 59 -1519
rect 376 -1520 377 -1519
rect 422 -1520 423 -1519
rect 625 -1520 626 -1519
rect 646 -1520 647 -1519
rect 982 -1520 983 -1519
rect 65 -1522 66 -1521
rect 86 -1522 87 -1521
rect 93 -1522 94 -1521
rect 313 -1522 314 -1521
rect 352 -1522 353 -1521
rect 439 -1522 440 -1521
rect 450 -1522 451 -1521
rect 513 -1522 514 -1521
rect 520 -1522 521 -1521
rect 537 -1522 538 -1521
rect 562 -1522 563 -1521
rect 597 -1522 598 -1521
rect 618 -1522 619 -1521
rect 842 -1522 843 -1521
rect 877 -1522 878 -1521
rect 1017 -1522 1018 -1521
rect 44 -1524 45 -1523
rect 65 -1524 66 -1523
rect 72 -1524 73 -1523
rect 828 -1524 829 -1523
rect 877 -1524 878 -1523
rect 933 -1524 934 -1523
rect 954 -1524 955 -1523
rect 1094 -1524 1095 -1523
rect 79 -1526 80 -1525
rect 544 -1526 545 -1525
rect 565 -1526 566 -1525
rect 814 -1526 815 -1525
rect 898 -1526 899 -1525
rect 1024 -1526 1025 -1525
rect 79 -1528 80 -1527
rect 548 -1528 549 -1527
rect 618 -1528 619 -1527
rect 695 -1528 696 -1527
rect 702 -1528 703 -1527
rect 730 -1528 731 -1527
rect 744 -1528 745 -1527
rect 856 -1528 857 -1527
rect 898 -1528 899 -1527
rect 975 -1528 976 -1527
rect 82 -1530 83 -1529
rect 478 -1530 479 -1529
rect 534 -1530 535 -1529
rect 1087 -1530 1088 -1529
rect 86 -1532 87 -1531
rect 170 -1532 171 -1531
rect 177 -1532 178 -1531
rect 226 -1532 227 -1531
rect 247 -1532 248 -1531
rect 275 -1532 276 -1531
rect 282 -1532 283 -1531
rect 352 -1532 353 -1531
rect 359 -1532 360 -1531
rect 632 -1532 633 -1531
rect 646 -1532 647 -1531
rect 800 -1532 801 -1531
rect 863 -1532 864 -1531
rect 975 -1532 976 -1531
rect 93 -1534 94 -1533
rect 415 -1534 416 -1533
rect 436 -1534 437 -1533
rect 803 -1534 804 -1533
rect 905 -1534 906 -1533
rect 1052 -1534 1053 -1533
rect 100 -1536 101 -1535
rect 240 -1536 241 -1535
rect 254 -1536 255 -1535
rect 303 -1536 304 -1535
rect 306 -1536 307 -1535
rect 905 -1536 906 -1535
rect 912 -1536 913 -1535
rect 919 -1536 920 -1535
rect 922 -1536 923 -1535
rect 961 -1536 962 -1535
rect 964 -1536 965 -1535
rect 989 -1536 990 -1535
rect 135 -1538 136 -1537
rect 394 -1538 395 -1537
rect 464 -1538 465 -1537
rect 499 -1538 500 -1537
rect 548 -1538 549 -1537
rect 611 -1538 612 -1537
rect 653 -1538 654 -1537
rect 947 -1538 948 -1537
rect 135 -1540 136 -1539
rect 457 -1540 458 -1539
rect 474 -1540 475 -1539
rect 709 -1540 710 -1539
rect 716 -1540 717 -1539
rect 814 -1540 815 -1539
rect 926 -1540 927 -1539
rect 1031 -1540 1032 -1539
rect 142 -1542 143 -1541
rect 345 -1542 346 -1541
rect 362 -1542 363 -1541
rect 954 -1542 955 -1541
rect 156 -1544 157 -1543
rect 429 -1544 430 -1543
rect 569 -1544 570 -1543
rect 611 -1544 612 -1543
rect 674 -1544 675 -1543
rect 891 -1544 892 -1543
rect 180 -1546 181 -1545
rect 212 -1546 213 -1545
rect 219 -1546 220 -1545
rect 282 -1546 283 -1545
rect 289 -1546 290 -1545
rect 576 -1546 577 -1545
rect 590 -1546 591 -1545
rect 653 -1546 654 -1545
rect 660 -1546 661 -1545
rect 674 -1546 675 -1545
rect 681 -1546 682 -1545
rect 821 -1546 822 -1545
rect 184 -1548 185 -1547
rect 324 -1548 325 -1547
rect 331 -1548 332 -1547
rect 597 -1548 598 -1547
rect 604 -1548 605 -1547
rect 716 -1548 717 -1547
rect 751 -1548 752 -1547
rect 863 -1548 864 -1547
rect 107 -1550 108 -1549
rect 331 -1550 332 -1549
rect 338 -1550 339 -1549
rect 569 -1550 570 -1549
rect 590 -1550 591 -1549
rect 688 -1550 689 -1549
rect 695 -1550 696 -1549
rect 737 -1550 738 -1549
rect 758 -1550 759 -1549
rect 1045 -1550 1046 -1549
rect 107 -1552 108 -1551
rect 114 -1552 115 -1551
rect 170 -1552 171 -1551
rect 338 -1552 339 -1551
rect 345 -1552 346 -1551
rect 443 -1552 444 -1551
rect 460 -1552 461 -1551
rect 737 -1552 738 -1551
rect 758 -1552 759 -1551
rect 912 -1552 913 -1551
rect 114 -1554 115 -1553
rect 450 -1554 451 -1553
rect 485 -1554 486 -1553
rect 751 -1554 752 -1553
rect 772 -1554 773 -1553
rect 884 -1554 885 -1553
rect 187 -1556 188 -1555
rect 439 -1556 440 -1555
rect 471 -1556 472 -1555
rect 485 -1556 486 -1555
rect 663 -1556 664 -1555
rect 688 -1556 689 -1555
rect 709 -1556 710 -1555
rect 1010 -1556 1011 -1555
rect 222 -1558 223 -1557
rect 660 -1558 661 -1557
rect 684 -1558 685 -1557
rect 989 -1558 990 -1557
rect 233 -1560 234 -1559
rect 457 -1560 458 -1559
rect 723 -1560 724 -1559
rect 772 -1560 773 -1559
rect 786 -1560 787 -1559
rect 933 -1560 934 -1559
rect 233 -1562 234 -1561
rect 667 -1562 668 -1561
rect 723 -1562 724 -1561
rect 779 -1562 780 -1561
rect 793 -1562 794 -1561
rect 926 -1562 927 -1561
rect 131 -1564 132 -1563
rect 793 -1564 794 -1563
rect 803 -1564 804 -1563
rect 1059 -1564 1060 -1563
rect 243 -1566 244 -1565
rect 576 -1566 577 -1565
rect 583 -1566 584 -1565
rect 786 -1566 787 -1565
rect 821 -1566 822 -1565
rect 849 -1566 850 -1565
rect 247 -1568 248 -1567
rect 684 -1568 685 -1567
rect 254 -1570 255 -1569
rect 292 -1570 293 -1569
rect 296 -1570 297 -1569
rect 604 -1570 605 -1569
rect 639 -1570 640 -1569
rect 779 -1570 780 -1569
rect 198 -1572 199 -1571
rect 296 -1572 297 -1571
rect 310 -1572 311 -1571
rect 744 -1572 745 -1571
rect 75 -1574 76 -1573
rect 310 -1574 311 -1573
rect 373 -1574 374 -1573
rect 464 -1574 465 -1573
rect 527 -1574 528 -1573
rect 639 -1574 640 -1573
rect 2 -1576 3 -1575
rect 373 -1576 374 -1575
rect 387 -1576 388 -1575
rect 422 -1576 423 -1575
rect 495 -1576 496 -1575
rect 527 -1576 528 -1575
rect 579 -1576 580 -1575
rect 849 -1576 850 -1575
rect 198 -1578 199 -1577
rect 205 -1578 206 -1577
rect 261 -1578 262 -1577
rect 471 -1578 472 -1577
rect 191 -1580 192 -1579
rect 205 -1580 206 -1579
rect 387 -1580 388 -1579
rect 516 -1580 517 -1579
rect 397 -1582 398 -1581
rect 443 -1582 444 -1581
rect 401 -1584 402 -1583
rect 583 -1584 584 -1583
rect 408 -1586 409 -1585
rect 429 -1586 430 -1585
rect 355 -1588 356 -1587
rect 408 -1588 409 -1587
rect 2 -1599 3 -1598
rect 299 -1599 300 -1598
rect 303 -1599 304 -1598
rect 324 -1599 325 -1598
rect 355 -1599 356 -1598
rect 786 -1599 787 -1598
rect 803 -1599 804 -1598
rect 1031 -1599 1032 -1598
rect 2 -1601 3 -1600
rect 159 -1601 160 -1600
rect 163 -1601 164 -1600
rect 341 -1601 342 -1600
rect 359 -1601 360 -1600
rect 429 -1601 430 -1600
rect 453 -1601 454 -1600
rect 982 -1601 983 -1600
rect 23 -1603 24 -1602
rect 250 -1603 251 -1602
rect 261 -1603 262 -1602
rect 352 -1603 353 -1602
rect 373 -1603 374 -1602
rect 583 -1603 584 -1602
rect 660 -1603 661 -1602
rect 688 -1603 689 -1602
rect 709 -1603 710 -1602
rect 1094 -1603 1095 -1602
rect 23 -1605 24 -1604
rect 107 -1605 108 -1604
rect 121 -1605 122 -1604
rect 793 -1605 794 -1604
rect 824 -1605 825 -1604
rect 919 -1605 920 -1604
rect 982 -1605 983 -1604
rect 1080 -1605 1081 -1604
rect 30 -1607 31 -1606
rect 233 -1607 234 -1606
rect 236 -1607 237 -1606
rect 254 -1607 255 -1606
rect 282 -1607 283 -1606
rect 415 -1607 416 -1606
rect 429 -1607 430 -1606
rect 527 -1607 528 -1606
rect 555 -1607 556 -1606
rect 709 -1607 710 -1606
rect 723 -1607 724 -1606
rect 800 -1607 801 -1606
rect 849 -1607 850 -1606
rect 915 -1607 916 -1606
rect 919 -1607 920 -1606
rect 968 -1607 969 -1606
rect 30 -1609 31 -1608
rect 485 -1609 486 -1608
rect 492 -1609 493 -1608
rect 590 -1609 591 -1608
rect 663 -1609 664 -1608
rect 891 -1609 892 -1608
rect 37 -1611 38 -1610
rect 47 -1611 48 -1610
rect 61 -1611 62 -1610
rect 450 -1611 451 -1610
rect 453 -1611 454 -1610
rect 898 -1611 899 -1610
rect 37 -1613 38 -1612
rect 128 -1613 129 -1612
rect 135 -1613 136 -1612
rect 362 -1613 363 -1612
rect 376 -1613 377 -1612
rect 380 -1613 381 -1612
rect 390 -1613 391 -1612
rect 576 -1613 577 -1612
rect 583 -1613 584 -1612
rect 611 -1613 612 -1612
rect 681 -1613 682 -1612
rect 737 -1613 738 -1612
rect 758 -1613 759 -1612
rect 1045 -1613 1046 -1612
rect 72 -1615 73 -1614
rect 828 -1615 829 -1614
rect 891 -1615 892 -1614
rect 961 -1615 962 -1614
rect 72 -1617 73 -1616
rect 443 -1617 444 -1616
rect 457 -1617 458 -1616
rect 779 -1617 780 -1616
rect 786 -1617 787 -1616
rect 835 -1617 836 -1616
rect 947 -1617 948 -1616
rect 961 -1617 962 -1616
rect 75 -1619 76 -1618
rect 240 -1619 241 -1618
rect 289 -1619 290 -1618
rect 373 -1619 374 -1618
rect 460 -1619 461 -1618
rect 541 -1619 542 -1618
rect 555 -1619 556 -1618
rect 1003 -1619 1004 -1618
rect 79 -1621 80 -1620
rect 632 -1621 633 -1620
rect 688 -1621 689 -1620
rect 702 -1621 703 -1620
rect 716 -1621 717 -1620
rect 898 -1621 899 -1620
rect 996 -1621 997 -1620
rect 1003 -1621 1004 -1620
rect 58 -1623 59 -1622
rect 632 -1623 633 -1622
rect 674 -1623 675 -1622
rect 716 -1623 717 -1622
rect 723 -1623 724 -1622
rect 765 -1623 766 -1622
rect 772 -1623 773 -1622
rect 849 -1623 850 -1622
rect 877 -1623 878 -1622
rect 947 -1623 948 -1622
rect 82 -1625 83 -1624
rect 597 -1625 598 -1624
rect 611 -1625 612 -1624
rect 639 -1625 640 -1624
rect 695 -1625 696 -1624
rect 758 -1625 759 -1624
rect 765 -1625 766 -1624
rect 856 -1625 857 -1624
rect 877 -1625 878 -1624
rect 975 -1625 976 -1624
rect 86 -1627 87 -1626
rect 243 -1627 244 -1626
rect 289 -1627 290 -1626
rect 310 -1627 311 -1626
rect 317 -1627 318 -1626
rect 537 -1627 538 -1626
rect 562 -1627 563 -1626
rect 576 -1627 577 -1626
rect 590 -1627 591 -1626
rect 618 -1627 619 -1626
rect 639 -1627 640 -1626
rect 954 -1627 955 -1626
rect 975 -1627 976 -1626
rect 1038 -1627 1039 -1626
rect 107 -1629 108 -1628
rect 338 -1629 339 -1628
rect 467 -1629 468 -1628
rect 1052 -1629 1053 -1628
rect 121 -1631 122 -1630
rect 194 -1631 195 -1630
rect 205 -1631 206 -1630
rect 261 -1631 262 -1630
rect 268 -1631 269 -1630
rect 338 -1631 339 -1630
rect 471 -1631 472 -1630
rect 695 -1631 696 -1630
rect 702 -1631 703 -1630
rect 744 -1631 745 -1630
rect 751 -1631 752 -1630
rect 954 -1631 955 -1630
rect 1052 -1631 1053 -1630
rect 1073 -1631 1074 -1630
rect 9 -1633 10 -1632
rect 205 -1633 206 -1632
rect 212 -1633 213 -1632
rect 254 -1633 255 -1632
rect 303 -1633 304 -1632
rect 408 -1633 409 -1632
rect 474 -1633 475 -1632
rect 1108 -1633 1109 -1632
rect 9 -1635 10 -1634
rect 135 -1635 136 -1634
rect 138 -1635 139 -1634
rect 268 -1635 269 -1634
rect 310 -1635 311 -1634
rect 387 -1635 388 -1634
rect 408 -1635 409 -1634
rect 646 -1635 647 -1634
rect 730 -1635 731 -1634
rect 1017 -1635 1018 -1634
rect 128 -1637 129 -1636
rect 184 -1637 185 -1636
rect 212 -1637 213 -1636
rect 842 -1637 843 -1636
rect 856 -1637 857 -1636
rect 926 -1637 927 -1636
rect 142 -1639 143 -1638
rect 401 -1639 402 -1638
rect 474 -1639 475 -1638
rect 737 -1639 738 -1638
rect 744 -1639 745 -1638
rect 814 -1639 815 -1638
rect 835 -1639 836 -1638
rect 933 -1639 934 -1638
rect 65 -1641 66 -1640
rect 401 -1641 402 -1640
rect 481 -1641 482 -1640
rect 905 -1641 906 -1640
rect 926 -1641 927 -1640
rect 1059 -1641 1060 -1640
rect 65 -1643 66 -1642
rect 124 -1643 125 -1642
rect 142 -1643 143 -1642
rect 177 -1643 178 -1642
rect 222 -1643 223 -1642
rect 296 -1643 297 -1642
rect 317 -1643 318 -1642
rect 436 -1643 437 -1642
rect 492 -1643 493 -1642
rect 828 -1643 829 -1642
rect 842 -1643 843 -1642
rect 940 -1643 941 -1642
rect 149 -1645 150 -1644
rect 184 -1645 185 -1644
rect 194 -1645 195 -1644
rect 436 -1645 437 -1644
rect 499 -1645 500 -1644
rect 527 -1645 528 -1644
rect 537 -1645 538 -1644
rect 1087 -1645 1088 -1644
rect 44 -1647 45 -1646
rect 149 -1647 150 -1646
rect 156 -1647 157 -1646
rect 443 -1647 444 -1646
rect 478 -1647 479 -1646
rect 499 -1647 500 -1646
rect 513 -1647 514 -1646
rect 1101 -1647 1102 -1646
rect 170 -1649 171 -1648
rect 534 -1649 535 -1648
rect 544 -1649 545 -1648
rect 618 -1649 619 -1648
rect 684 -1649 685 -1648
rect 940 -1649 941 -1648
rect 170 -1651 171 -1650
rect 198 -1651 199 -1650
rect 222 -1651 223 -1650
rect 275 -1651 276 -1650
rect 296 -1651 297 -1650
rect 506 -1651 507 -1650
rect 513 -1651 514 -1650
rect 887 -1651 888 -1650
rect 905 -1651 906 -1650
rect 1010 -1651 1011 -1650
rect 86 -1653 87 -1652
rect 198 -1653 199 -1652
rect 226 -1653 227 -1652
rect 870 -1653 871 -1652
rect 933 -1653 934 -1652
rect 1024 -1653 1025 -1652
rect 16 -1655 17 -1654
rect 226 -1655 227 -1654
rect 233 -1655 234 -1654
rect 282 -1655 283 -1654
rect 366 -1655 367 -1654
rect 506 -1655 507 -1654
rect 520 -1655 521 -1654
rect 674 -1655 675 -1654
rect 772 -1655 773 -1654
rect 894 -1655 895 -1654
rect 16 -1657 17 -1656
rect 51 -1657 52 -1656
rect 163 -1657 164 -1656
rect 366 -1657 367 -1656
rect 387 -1657 388 -1656
rect 450 -1657 451 -1656
rect 565 -1657 566 -1656
rect 1066 -1657 1067 -1656
rect 51 -1659 52 -1658
rect 569 -1659 570 -1658
rect 597 -1659 598 -1658
rect 625 -1659 626 -1658
rect 779 -1659 780 -1658
rect 884 -1659 885 -1658
rect 177 -1661 178 -1660
rect 422 -1661 423 -1660
rect 558 -1661 559 -1660
rect 569 -1661 570 -1660
rect 604 -1661 605 -1660
rect 751 -1661 752 -1660
rect 793 -1661 794 -1660
rect 863 -1661 864 -1660
rect 100 -1663 101 -1662
rect 422 -1663 423 -1662
rect 464 -1663 465 -1662
rect 604 -1663 605 -1662
rect 625 -1663 626 -1662
rect 653 -1663 654 -1662
rect 814 -1663 815 -1662
rect 912 -1663 913 -1662
rect 100 -1665 101 -1664
rect 247 -1665 248 -1664
rect 275 -1665 276 -1664
rect 807 -1665 808 -1664
rect 821 -1665 822 -1664
rect 870 -1665 871 -1664
rect 93 -1667 94 -1666
rect 247 -1667 248 -1666
rect 345 -1667 346 -1666
rect 520 -1667 521 -1666
rect 653 -1667 654 -1666
rect 667 -1667 668 -1666
rect 733 -1667 734 -1666
rect 807 -1667 808 -1666
rect 863 -1667 864 -1666
rect 989 -1667 990 -1666
rect 345 -1669 346 -1668
rect 457 -1669 458 -1668
rect 478 -1669 479 -1668
rect 821 -1669 822 -1668
rect 394 -1671 395 -1670
rect 646 -1671 647 -1670
rect 331 -1673 332 -1672
rect 394 -1673 395 -1672
rect 488 -1673 489 -1672
rect 667 -1673 668 -1672
rect 331 -1675 332 -1674
rect 464 -1675 465 -1674
rect 2 -1686 3 -1685
rect 376 -1686 377 -1685
rect 443 -1686 444 -1685
rect 562 -1686 563 -1685
rect 593 -1686 594 -1685
rect 1017 -1686 1018 -1685
rect 1027 -1686 1028 -1685
rect 1052 -1686 1053 -1685
rect 2 -1688 3 -1687
rect 96 -1688 97 -1687
rect 110 -1688 111 -1687
rect 128 -1688 129 -1687
rect 152 -1688 153 -1687
rect 275 -1688 276 -1687
rect 282 -1688 283 -1687
rect 394 -1688 395 -1687
rect 429 -1688 430 -1687
rect 562 -1688 563 -1687
rect 621 -1688 622 -1687
rect 716 -1688 717 -1687
rect 730 -1688 731 -1687
rect 870 -1688 871 -1687
rect 887 -1688 888 -1687
rect 961 -1688 962 -1687
rect 1003 -1688 1004 -1687
rect 1010 -1688 1011 -1687
rect 9 -1690 10 -1689
rect 191 -1690 192 -1689
rect 198 -1690 199 -1689
rect 597 -1690 598 -1689
rect 649 -1690 650 -1689
rect 856 -1690 857 -1689
rect 891 -1690 892 -1689
rect 982 -1690 983 -1689
rect 16 -1692 17 -1691
rect 215 -1692 216 -1691
rect 233 -1692 234 -1691
rect 436 -1692 437 -1691
rect 443 -1692 444 -1691
rect 677 -1692 678 -1691
rect 716 -1692 717 -1691
rect 723 -1692 724 -1691
rect 730 -1692 731 -1691
rect 758 -1692 759 -1691
rect 779 -1692 780 -1691
rect 782 -1692 783 -1691
rect 803 -1692 804 -1691
rect 807 -1692 808 -1691
rect 821 -1692 822 -1691
rect 968 -1692 969 -1691
rect 23 -1694 24 -1693
rect 194 -1694 195 -1693
rect 198 -1694 199 -1693
rect 254 -1694 255 -1693
rect 275 -1694 276 -1693
rect 733 -1694 734 -1693
rect 779 -1694 780 -1693
rect 814 -1694 815 -1693
rect 835 -1694 836 -1693
rect 870 -1694 871 -1693
rect 912 -1694 913 -1693
rect 975 -1694 976 -1693
rect 23 -1696 24 -1695
rect 222 -1696 223 -1695
rect 240 -1696 241 -1695
rect 411 -1696 412 -1695
rect 415 -1696 416 -1695
rect 436 -1696 437 -1695
rect 457 -1696 458 -1695
rect 856 -1696 857 -1695
rect 898 -1696 899 -1695
rect 975 -1696 976 -1695
rect 30 -1698 31 -1697
rect 467 -1698 468 -1697
rect 471 -1698 472 -1697
rect 751 -1698 752 -1697
rect 793 -1698 794 -1697
rect 814 -1698 815 -1697
rect 835 -1698 836 -1697
rect 940 -1698 941 -1697
rect 30 -1700 31 -1699
rect 345 -1700 346 -1699
rect 348 -1700 349 -1699
rect 387 -1700 388 -1699
rect 394 -1700 395 -1699
rect 506 -1700 507 -1699
rect 548 -1700 549 -1699
rect 807 -1700 808 -1699
rect 898 -1700 899 -1699
rect 919 -1700 920 -1699
rect 926 -1700 927 -1699
rect 961 -1700 962 -1699
rect 37 -1702 38 -1701
rect 180 -1702 181 -1701
rect 184 -1702 185 -1701
rect 191 -1702 192 -1701
rect 222 -1702 223 -1701
rect 261 -1702 262 -1701
rect 285 -1702 286 -1701
rect 408 -1702 409 -1701
rect 467 -1702 468 -1701
rect 737 -1702 738 -1701
rect 793 -1702 794 -1701
rect 828 -1702 829 -1701
rect 863 -1702 864 -1701
rect 919 -1702 920 -1701
rect 940 -1702 941 -1701
rect 1006 -1702 1007 -1701
rect 37 -1704 38 -1703
rect 292 -1704 293 -1703
rect 299 -1704 300 -1703
rect 551 -1704 552 -1703
rect 555 -1704 556 -1703
rect 618 -1704 619 -1703
rect 639 -1704 640 -1703
rect 891 -1704 892 -1703
rect 44 -1706 45 -1705
rect 61 -1706 62 -1705
rect 65 -1706 66 -1705
rect 166 -1706 167 -1705
rect 170 -1706 171 -1705
rect 296 -1706 297 -1705
rect 317 -1706 318 -1705
rect 425 -1706 426 -1705
rect 464 -1706 465 -1705
rect 639 -1706 640 -1705
rect 688 -1706 689 -1705
rect 751 -1706 752 -1705
rect 782 -1706 783 -1705
rect 828 -1706 829 -1705
rect 16 -1708 17 -1707
rect 464 -1708 465 -1707
rect 471 -1708 472 -1707
rect 565 -1708 566 -1707
rect 569 -1708 570 -1707
rect 688 -1708 689 -1707
rect 723 -1708 724 -1707
rect 744 -1708 745 -1707
rect 44 -1710 45 -1709
rect 404 -1710 405 -1709
rect 408 -1710 409 -1709
rect 709 -1710 710 -1709
rect 51 -1712 52 -1711
rect 383 -1712 384 -1711
rect 478 -1712 479 -1711
rect 534 -1712 535 -1711
rect 548 -1712 549 -1711
rect 576 -1712 577 -1711
rect 597 -1712 598 -1711
rect 632 -1712 633 -1711
rect 51 -1714 52 -1713
rect 93 -1714 94 -1713
rect 128 -1714 129 -1713
rect 481 -1714 482 -1713
rect 485 -1714 486 -1713
rect 989 -1714 990 -1713
rect 54 -1716 55 -1715
rect 254 -1716 255 -1715
rect 261 -1716 262 -1715
rect 324 -1716 325 -1715
rect 338 -1716 339 -1715
rect 345 -1716 346 -1715
rect 352 -1716 353 -1715
rect 380 -1716 381 -1715
rect 481 -1716 482 -1715
rect 611 -1716 612 -1715
rect 614 -1716 615 -1715
rect 709 -1716 710 -1715
rect 65 -1718 66 -1717
rect 229 -1718 230 -1717
rect 243 -1718 244 -1717
rect 268 -1718 269 -1717
rect 289 -1718 290 -1717
rect 513 -1718 514 -1717
rect 516 -1718 517 -1717
rect 737 -1718 738 -1717
rect 72 -1720 73 -1719
rect 450 -1720 451 -1719
rect 488 -1720 489 -1719
rect 527 -1720 528 -1719
rect 576 -1720 577 -1719
rect 590 -1720 591 -1719
rect 618 -1720 619 -1719
rect 758 -1720 759 -1719
rect 72 -1722 73 -1721
rect 163 -1722 164 -1721
rect 177 -1722 178 -1721
rect 429 -1722 430 -1721
rect 450 -1722 451 -1721
rect 660 -1722 661 -1721
rect 79 -1724 80 -1723
rect 121 -1724 122 -1723
rect 135 -1724 136 -1723
rect 478 -1724 479 -1723
rect 492 -1724 493 -1723
rect 954 -1724 955 -1723
rect 86 -1726 87 -1725
rect 744 -1726 745 -1725
rect 947 -1726 948 -1725
rect 954 -1726 955 -1725
rect 86 -1728 87 -1727
rect 103 -1728 104 -1727
rect 121 -1728 122 -1727
rect 142 -1728 143 -1727
rect 149 -1728 150 -1727
rect 383 -1728 384 -1727
rect 401 -1728 402 -1727
rect 527 -1728 528 -1727
rect 541 -1728 542 -1727
rect 660 -1728 661 -1727
rect 905 -1728 906 -1727
rect 947 -1728 948 -1727
rect 138 -1730 139 -1729
rect 926 -1730 927 -1729
rect 142 -1732 143 -1731
rect 303 -1732 304 -1731
rect 317 -1732 318 -1731
rect 474 -1732 475 -1731
rect 492 -1732 493 -1731
rect 894 -1732 895 -1731
rect 149 -1734 150 -1733
rect 240 -1734 241 -1733
rect 247 -1734 248 -1733
rect 558 -1734 559 -1733
rect 156 -1736 157 -1735
rect 201 -1736 202 -1735
rect 268 -1736 269 -1735
rect 324 -1736 325 -1735
rect 331 -1736 332 -1735
rect 338 -1736 339 -1735
rect 352 -1736 353 -1735
rect 453 -1736 454 -1735
rect 495 -1736 496 -1735
rect 674 -1736 675 -1735
rect 156 -1738 157 -1737
rect 226 -1738 227 -1737
rect 289 -1738 290 -1737
rect 359 -1738 360 -1737
rect 366 -1738 367 -1737
rect 653 -1738 654 -1737
rect 674 -1738 675 -1737
rect 877 -1738 878 -1737
rect 100 -1740 101 -1739
rect 359 -1740 360 -1739
rect 366 -1740 367 -1739
rect 982 -1740 983 -1739
rect 100 -1742 101 -1741
rect 170 -1742 171 -1741
rect 177 -1742 178 -1741
rect 247 -1742 248 -1741
rect 303 -1742 304 -1741
rect 310 -1742 311 -1741
rect 369 -1742 370 -1741
rect 520 -1742 521 -1741
rect 541 -1742 542 -1741
rect 905 -1742 906 -1741
rect 114 -1744 115 -1743
rect 520 -1744 521 -1743
rect 842 -1744 843 -1743
rect 877 -1744 878 -1743
rect 107 -1746 108 -1745
rect 114 -1746 115 -1745
rect 163 -1746 164 -1745
rect 313 -1746 314 -1745
rect 331 -1746 332 -1745
rect 369 -1746 370 -1745
rect 373 -1746 374 -1745
rect 415 -1746 416 -1745
rect 485 -1746 486 -1745
rect 653 -1746 654 -1745
rect 786 -1746 787 -1745
rect 842 -1746 843 -1745
rect 107 -1748 108 -1747
rect 821 -1748 822 -1747
rect 187 -1750 188 -1749
rect 863 -1750 864 -1749
rect 226 -1752 227 -1751
rect 625 -1752 626 -1751
rect 786 -1752 787 -1751
rect 933 -1752 934 -1751
rect 401 -1754 402 -1753
rect 457 -1754 458 -1753
rect 499 -1754 500 -1753
rect 506 -1754 507 -1753
rect 513 -1754 514 -1753
rect 583 -1754 584 -1753
rect 625 -1754 626 -1753
rect 667 -1754 668 -1753
rect 884 -1754 885 -1753
rect 933 -1754 934 -1753
rect 373 -1756 374 -1755
rect 499 -1756 500 -1755
rect 583 -1756 584 -1755
rect 702 -1756 703 -1755
rect 800 -1756 801 -1755
rect 884 -1756 885 -1755
rect 604 -1758 605 -1757
rect 702 -1758 703 -1757
rect 604 -1760 605 -1759
rect 646 -1760 647 -1759
rect 667 -1760 668 -1759
rect 681 -1760 682 -1759
rect 569 -1762 570 -1761
rect 646 -1762 647 -1761
rect 681 -1762 682 -1761
rect 695 -1762 696 -1761
rect 695 -1764 696 -1763
rect 765 -1764 766 -1763
rect 765 -1766 766 -1765
rect 772 -1766 773 -1765
rect 422 -1768 423 -1767
rect 772 -1768 773 -1767
rect 422 -1770 423 -1769
rect 912 -1770 913 -1769
rect 2 -1781 3 -1780
rect 187 -1781 188 -1780
rect 205 -1781 206 -1780
rect 523 -1781 524 -1780
rect 565 -1781 566 -1780
rect 947 -1781 948 -1780
rect 975 -1781 976 -1780
rect 999 -1781 1000 -1780
rect 9 -1783 10 -1782
rect 30 -1783 31 -1782
rect 37 -1783 38 -1782
rect 310 -1783 311 -1782
rect 313 -1783 314 -1782
rect 499 -1783 500 -1782
rect 506 -1783 507 -1782
rect 516 -1783 517 -1782
rect 590 -1783 591 -1782
rect 961 -1783 962 -1782
rect 996 -1783 997 -1782
rect 1010 -1783 1011 -1782
rect 23 -1785 24 -1784
rect 212 -1785 213 -1784
rect 215 -1785 216 -1784
rect 296 -1785 297 -1784
rect 310 -1785 311 -1784
rect 457 -1785 458 -1784
rect 460 -1785 461 -1784
rect 919 -1785 920 -1784
rect 947 -1785 948 -1784
rect 1024 -1785 1025 -1784
rect 44 -1787 45 -1786
rect 366 -1787 367 -1786
rect 369 -1787 370 -1786
rect 394 -1787 395 -1786
rect 422 -1787 423 -1786
rect 702 -1787 703 -1786
rect 726 -1787 727 -1786
rect 954 -1787 955 -1786
rect 51 -1789 52 -1788
rect 891 -1789 892 -1788
rect 915 -1789 916 -1788
rect 933 -1789 934 -1788
rect 51 -1791 52 -1790
rect 348 -1791 349 -1790
rect 369 -1791 370 -1790
rect 387 -1791 388 -1790
rect 450 -1791 451 -1790
rect 541 -1791 542 -1790
rect 590 -1791 591 -1790
rect 604 -1791 605 -1790
rect 611 -1791 612 -1790
rect 856 -1791 857 -1790
rect 54 -1793 55 -1792
rect 72 -1793 73 -1792
rect 79 -1793 80 -1792
rect 103 -1793 104 -1792
rect 107 -1793 108 -1792
rect 191 -1793 192 -1792
rect 215 -1793 216 -1792
rect 656 -1793 657 -1792
rect 674 -1793 675 -1792
rect 814 -1793 815 -1792
rect 842 -1793 843 -1792
rect 852 -1793 853 -1792
rect 58 -1795 59 -1794
rect 121 -1795 122 -1794
rect 128 -1795 129 -1794
rect 149 -1795 150 -1794
rect 177 -1795 178 -1794
rect 229 -1795 230 -1794
rect 240 -1795 241 -1794
rect 527 -1795 528 -1794
rect 541 -1795 542 -1794
rect 628 -1795 629 -1794
rect 632 -1795 633 -1794
rect 926 -1795 927 -1794
rect 65 -1797 66 -1796
rect 327 -1797 328 -1796
rect 380 -1797 381 -1796
rect 639 -1797 640 -1796
rect 642 -1797 643 -1796
rect 989 -1797 990 -1796
rect 65 -1799 66 -1798
rect 142 -1799 143 -1798
rect 149 -1799 150 -1798
rect 156 -1799 157 -1798
rect 170 -1799 171 -1798
rect 177 -1799 178 -1798
rect 226 -1799 227 -1798
rect 401 -1799 402 -1798
rect 415 -1799 416 -1798
rect 450 -1799 451 -1798
rect 464 -1799 465 -1798
rect 548 -1799 549 -1798
rect 604 -1799 605 -1798
rect 744 -1799 745 -1798
rect 814 -1799 815 -1798
rect 898 -1799 899 -1798
rect 72 -1801 73 -1800
rect 415 -1801 416 -1800
rect 464 -1801 465 -1800
rect 562 -1801 563 -1800
rect 611 -1801 612 -1800
rect 765 -1801 766 -1800
rect 898 -1801 899 -1800
rect 950 -1801 951 -1800
rect 79 -1803 80 -1802
rect 593 -1803 594 -1802
rect 618 -1803 619 -1802
rect 751 -1803 752 -1802
rect 93 -1805 94 -1804
rect 128 -1805 129 -1804
rect 135 -1805 136 -1804
rect 184 -1805 185 -1804
rect 226 -1805 227 -1804
rect 551 -1805 552 -1804
rect 618 -1805 619 -1804
rect 723 -1805 724 -1804
rect 751 -1805 752 -1804
rect 849 -1805 850 -1804
rect 93 -1807 94 -1806
rect 114 -1807 115 -1806
rect 121 -1807 122 -1806
rect 425 -1807 426 -1806
rect 467 -1807 468 -1806
rect 513 -1807 514 -1806
rect 527 -1807 528 -1806
rect 982 -1807 983 -1806
rect 100 -1809 101 -1808
rect 401 -1809 402 -1808
rect 478 -1809 479 -1808
rect 534 -1809 535 -1808
rect 548 -1809 549 -1808
rect 765 -1809 766 -1808
rect 100 -1811 101 -1810
rect 198 -1811 199 -1810
rect 243 -1811 244 -1810
rect 387 -1811 388 -1810
rect 499 -1811 500 -1810
rect 625 -1811 626 -1810
rect 635 -1811 636 -1810
rect 828 -1811 829 -1810
rect 110 -1813 111 -1812
rect 492 -1813 493 -1812
rect 506 -1813 507 -1812
rect 772 -1813 773 -1812
rect 828 -1813 829 -1812
rect 835 -1813 836 -1812
rect 86 -1815 87 -1814
rect 492 -1815 493 -1814
rect 534 -1815 535 -1814
rect 555 -1815 556 -1814
rect 576 -1815 577 -1814
rect 835 -1815 836 -1814
rect 86 -1817 87 -1816
rect 201 -1817 202 -1816
rect 254 -1817 255 -1816
rect 562 -1817 563 -1816
rect 576 -1817 577 -1816
rect 597 -1817 598 -1816
rect 621 -1817 622 -1816
rect 744 -1817 745 -1816
rect 114 -1819 115 -1818
rect 443 -1819 444 -1818
rect 555 -1819 556 -1818
rect 667 -1819 668 -1818
rect 674 -1819 675 -1818
rect 716 -1819 717 -1818
rect 135 -1821 136 -1820
rect 163 -1821 164 -1820
rect 170 -1821 171 -1820
rect 457 -1821 458 -1820
rect 646 -1821 647 -1820
rect 856 -1821 857 -1820
rect 142 -1823 143 -1822
rect 303 -1823 304 -1822
rect 380 -1823 381 -1822
rect 520 -1823 521 -1822
rect 653 -1823 654 -1822
rect 870 -1823 871 -1822
rect 156 -1825 157 -1824
rect 219 -1825 220 -1824
rect 247 -1825 248 -1824
rect 303 -1825 304 -1824
rect 418 -1825 419 -1824
rect 646 -1825 647 -1824
rect 653 -1825 654 -1824
rect 730 -1825 731 -1824
rect 194 -1827 195 -1826
rect 219 -1827 220 -1826
rect 247 -1827 248 -1826
rect 275 -1827 276 -1826
rect 282 -1827 283 -1826
rect 394 -1827 395 -1826
rect 443 -1827 444 -1826
rect 688 -1827 689 -1826
rect 702 -1827 703 -1826
rect 1017 -1827 1018 -1826
rect 254 -1829 255 -1828
rect 324 -1829 325 -1828
rect 520 -1829 521 -1828
rect 877 -1829 878 -1828
rect 268 -1831 269 -1830
rect 373 -1831 374 -1830
rect 660 -1831 661 -1830
rect 772 -1831 773 -1830
rect 786 -1831 787 -1830
rect 877 -1831 878 -1830
rect 261 -1833 262 -1832
rect 268 -1833 269 -1832
rect 275 -1833 276 -1832
rect 677 -1833 678 -1832
rect 681 -1833 682 -1832
rect 800 -1833 801 -1832
rect 233 -1835 234 -1834
rect 261 -1835 262 -1834
rect 282 -1835 283 -1834
rect 338 -1835 339 -1834
rect 373 -1835 374 -1834
rect 408 -1835 409 -1834
rect 597 -1835 598 -1834
rect 660 -1835 661 -1834
rect 667 -1835 668 -1834
rect 940 -1835 941 -1834
rect 233 -1837 234 -1836
rect 352 -1837 353 -1836
rect 408 -1837 409 -1836
rect 849 -1837 850 -1836
rect 289 -1839 290 -1838
rect 352 -1839 353 -1838
rect 681 -1839 682 -1838
rect 695 -1839 696 -1838
rect 709 -1839 710 -1838
rect 870 -1839 871 -1838
rect 289 -1841 290 -1840
rect 331 -1841 332 -1840
rect 338 -1841 339 -1840
rect 485 -1841 486 -1840
rect 688 -1841 689 -1840
rect 779 -1841 780 -1840
rect 786 -1841 787 -1840
rect 863 -1841 864 -1840
rect 296 -1843 297 -1842
rect 376 -1843 377 -1842
rect 695 -1843 696 -1842
rect 793 -1843 794 -1842
rect 838 -1843 839 -1842
rect 863 -1843 864 -1842
rect 317 -1845 318 -1844
rect 485 -1845 486 -1844
rect 709 -1845 710 -1844
rect 758 -1845 759 -1844
rect 793 -1845 794 -1844
rect 842 -1845 843 -1844
rect 317 -1847 318 -1846
rect 345 -1847 346 -1846
rect 716 -1847 717 -1846
rect 807 -1847 808 -1846
rect 324 -1849 325 -1848
rect 436 -1849 437 -1848
rect 730 -1849 731 -1848
rect 821 -1849 822 -1848
rect 331 -1851 332 -1850
rect 569 -1851 570 -1850
rect 737 -1851 738 -1850
rect 779 -1851 780 -1850
rect 807 -1851 808 -1850
rect 968 -1851 969 -1850
rect 345 -1853 346 -1852
rect 1003 -1853 1004 -1852
rect 429 -1855 430 -1854
rect 436 -1855 437 -1854
rect 569 -1855 570 -1854
rect 884 -1855 885 -1854
rect 429 -1857 430 -1856
rect 471 -1857 472 -1856
rect 737 -1857 738 -1856
rect 912 -1857 913 -1856
rect 359 -1859 360 -1858
rect 471 -1859 472 -1858
rect 758 -1859 759 -1858
rect 845 -1859 846 -1858
rect 821 -1861 822 -1860
rect 905 -1861 906 -1860
rect 16 -1872 17 -1871
rect 51 -1872 52 -1871
rect 58 -1872 59 -1871
rect 163 -1872 164 -1871
rect 184 -1872 185 -1871
rect 198 -1872 199 -1871
rect 219 -1872 220 -1871
rect 261 -1872 262 -1871
rect 285 -1872 286 -1871
rect 870 -1872 871 -1871
rect 23 -1874 24 -1873
rect 184 -1874 185 -1873
rect 194 -1874 195 -1873
rect 198 -1874 199 -1873
rect 229 -1874 230 -1873
rect 240 -1874 241 -1873
rect 243 -1874 244 -1873
rect 317 -1874 318 -1873
rect 324 -1874 325 -1873
rect 411 -1874 412 -1873
rect 415 -1874 416 -1873
rect 450 -1874 451 -1873
rect 464 -1874 465 -1873
rect 467 -1874 468 -1873
rect 509 -1874 510 -1873
rect 737 -1874 738 -1873
rect 782 -1874 783 -1873
rect 877 -1874 878 -1873
rect 51 -1876 52 -1875
rect 191 -1876 192 -1875
rect 247 -1876 248 -1875
rect 324 -1876 325 -1875
rect 334 -1876 335 -1875
rect 709 -1876 710 -1875
rect 845 -1876 846 -1875
rect 898 -1876 899 -1875
rect 58 -1878 59 -1877
rect 296 -1878 297 -1877
rect 348 -1878 349 -1877
rect 352 -1878 353 -1877
rect 359 -1878 360 -1877
rect 439 -1878 440 -1877
rect 443 -1878 444 -1877
rect 639 -1878 640 -1877
rect 702 -1878 703 -1877
rect 821 -1878 822 -1877
rect 65 -1880 66 -1879
rect 159 -1880 160 -1879
rect 177 -1880 178 -1879
rect 243 -1880 244 -1879
rect 247 -1880 248 -1879
rect 387 -1880 388 -1879
rect 411 -1880 412 -1879
rect 460 -1880 461 -1879
rect 464 -1880 465 -1879
rect 478 -1880 479 -1879
rect 520 -1880 521 -1879
rect 583 -1880 584 -1879
rect 618 -1880 619 -1879
rect 663 -1880 664 -1879
rect 702 -1880 703 -1879
rect 758 -1880 759 -1879
rect 821 -1880 822 -1879
rect 863 -1880 864 -1879
rect 65 -1882 66 -1881
rect 124 -1882 125 -1881
rect 128 -1882 129 -1881
rect 149 -1882 150 -1881
rect 177 -1882 178 -1881
rect 457 -1882 458 -1881
rect 471 -1882 472 -1881
rect 737 -1882 738 -1881
rect 758 -1882 759 -1881
rect 793 -1882 794 -1881
rect 72 -1884 73 -1883
rect 240 -1884 241 -1883
rect 296 -1884 297 -1883
rect 401 -1884 402 -1883
rect 418 -1884 419 -1883
rect 618 -1884 619 -1883
rect 628 -1884 629 -1883
rect 674 -1884 675 -1883
rect 709 -1884 710 -1883
rect 761 -1884 762 -1883
rect 793 -1884 794 -1883
rect 856 -1884 857 -1883
rect 72 -1886 73 -1885
rect 145 -1886 146 -1885
rect 191 -1886 192 -1885
rect 275 -1886 276 -1885
rect 338 -1886 339 -1885
rect 352 -1886 353 -1885
rect 362 -1886 363 -1885
rect 485 -1886 486 -1885
rect 527 -1886 528 -1885
rect 814 -1886 815 -1885
rect 79 -1888 80 -1887
rect 229 -1888 230 -1887
rect 289 -1888 290 -1887
rect 338 -1888 339 -1887
rect 366 -1888 367 -1887
rect 523 -1888 524 -1887
rect 530 -1888 531 -1887
rect 597 -1888 598 -1887
rect 632 -1888 633 -1887
rect 786 -1888 787 -1887
rect 814 -1888 815 -1887
rect 828 -1888 829 -1887
rect 79 -1890 80 -1889
rect 282 -1890 283 -1889
rect 289 -1890 290 -1889
rect 317 -1890 318 -1889
rect 373 -1890 374 -1889
rect 632 -1890 633 -1889
rect 674 -1890 675 -1889
rect 716 -1890 717 -1889
rect 751 -1890 752 -1889
rect 786 -1890 787 -1889
rect 44 -1892 45 -1891
rect 282 -1892 283 -1891
rect 310 -1892 311 -1891
rect 373 -1892 374 -1891
rect 387 -1892 388 -1891
rect 450 -1892 451 -1891
rect 471 -1892 472 -1891
rect 772 -1892 773 -1891
rect 100 -1894 101 -1893
rect 261 -1894 262 -1893
rect 394 -1894 395 -1893
rect 401 -1894 402 -1893
rect 408 -1894 409 -1893
rect 597 -1894 598 -1893
rect 646 -1894 647 -1893
rect 716 -1894 717 -1893
rect 751 -1894 752 -1893
rect 779 -1894 780 -1893
rect 100 -1896 101 -1895
rect 114 -1896 115 -1895
rect 121 -1896 122 -1895
rect 163 -1896 164 -1895
rect 215 -1896 216 -1895
rect 418 -1896 419 -1895
rect 422 -1896 423 -1895
rect 642 -1896 643 -1895
rect 646 -1896 647 -1895
rect 688 -1896 689 -1895
rect 86 -1898 87 -1897
rect 121 -1898 122 -1897
rect 142 -1898 143 -1897
rect 275 -1898 276 -1897
rect 408 -1898 409 -1897
rect 667 -1898 668 -1897
rect 681 -1898 682 -1897
rect 688 -1898 689 -1897
rect 86 -1900 87 -1899
rect 233 -1900 234 -1899
rect 380 -1900 381 -1899
rect 667 -1900 668 -1899
rect 681 -1900 682 -1899
rect 772 -1900 773 -1899
rect 93 -1902 94 -1901
rect 142 -1902 143 -1901
rect 212 -1902 213 -1901
rect 380 -1902 381 -1901
rect 422 -1902 423 -1901
rect 723 -1902 724 -1901
rect 93 -1904 94 -1903
rect 331 -1904 332 -1903
rect 429 -1904 430 -1903
rect 443 -1904 444 -1903
rect 478 -1904 479 -1903
rect 492 -1904 493 -1903
rect 548 -1904 549 -1903
rect 726 -1904 727 -1903
rect 107 -1906 108 -1905
rect 205 -1906 206 -1905
rect 212 -1906 213 -1905
rect 268 -1906 269 -1905
rect 310 -1906 311 -1905
rect 331 -1906 332 -1905
rect 429 -1906 430 -1905
rect 513 -1906 514 -1905
rect 548 -1906 549 -1905
rect 604 -1906 605 -1905
rect 625 -1906 626 -1905
rect 723 -1906 724 -1905
rect 107 -1908 108 -1907
rect 135 -1908 136 -1907
rect 166 -1908 167 -1907
rect 205 -1908 206 -1907
rect 268 -1908 269 -1907
rect 303 -1908 304 -1907
rect 457 -1908 458 -1907
rect 513 -1908 514 -1907
rect 551 -1908 552 -1907
rect 800 -1908 801 -1907
rect 114 -1910 115 -1909
rect 156 -1910 157 -1909
rect 254 -1910 255 -1909
rect 303 -1910 304 -1909
rect 485 -1910 486 -1909
rect 506 -1910 507 -1909
rect 583 -1910 584 -1909
rect 660 -1910 661 -1909
rect 135 -1912 136 -1911
rect 170 -1912 171 -1911
rect 254 -1912 255 -1911
rect 569 -1912 570 -1911
rect 604 -1912 605 -1911
rect 807 -1912 808 -1911
rect 131 -1914 132 -1913
rect 170 -1914 171 -1913
rect 492 -1914 493 -1913
rect 499 -1914 500 -1913
rect 506 -1914 507 -1913
rect 541 -1914 542 -1913
rect 562 -1914 563 -1913
rect 660 -1914 661 -1913
rect 149 -1916 150 -1915
rect 156 -1916 157 -1915
rect 394 -1916 395 -1915
rect 562 -1916 563 -1915
rect 625 -1916 626 -1915
rect 695 -1916 696 -1915
rect 499 -1918 500 -1917
rect 576 -1918 577 -1917
rect 653 -1918 654 -1917
rect 695 -1918 696 -1917
rect 467 -1920 468 -1919
rect 576 -1920 577 -1919
rect 611 -1920 612 -1919
rect 653 -1920 654 -1919
rect 453 -1922 454 -1921
rect 611 -1922 612 -1921
rect 534 -1924 535 -1923
rect 569 -1924 570 -1923
rect 534 -1926 535 -1925
rect 590 -1926 591 -1925
rect 541 -1928 542 -1927
rect 555 -1928 556 -1927
rect 555 -1930 556 -1929
rect 730 -1930 731 -1929
rect 730 -1932 731 -1931
rect 817 -1932 818 -1931
rect 33 -1943 34 -1942
rect 37 -1943 38 -1942
rect 40 -1943 41 -1942
rect 47 -1943 48 -1942
rect 51 -1943 52 -1942
rect 394 -1943 395 -1942
rect 418 -1943 419 -1942
rect 667 -1943 668 -1942
rect 677 -1943 678 -1942
rect 688 -1943 689 -1942
rect 695 -1943 696 -1942
rect 800 -1943 801 -1942
rect 37 -1945 38 -1944
rect 114 -1945 115 -1944
rect 121 -1945 122 -1944
rect 177 -1945 178 -1944
rect 191 -1945 192 -1944
rect 548 -1945 549 -1944
rect 576 -1945 577 -1944
rect 730 -1945 731 -1944
rect 782 -1945 783 -1944
rect 821 -1945 822 -1944
rect 44 -1947 45 -1946
rect 135 -1947 136 -1946
rect 138 -1947 139 -1946
rect 264 -1947 265 -1946
rect 275 -1947 276 -1946
rect 331 -1947 332 -1946
rect 373 -1947 374 -1946
rect 411 -1947 412 -1946
rect 446 -1947 447 -1946
rect 492 -1947 493 -1946
rect 495 -1947 496 -1946
rect 541 -1947 542 -1946
rect 593 -1947 594 -1946
rect 625 -1947 626 -1946
rect 653 -1947 654 -1946
rect 758 -1947 759 -1946
rect 786 -1947 787 -1946
rect 807 -1947 808 -1946
rect 58 -1949 59 -1948
rect 236 -1949 237 -1948
rect 243 -1949 244 -1948
rect 387 -1949 388 -1948
rect 394 -1949 395 -1948
rect 779 -1949 780 -1948
rect 72 -1951 73 -1950
rect 75 -1951 76 -1950
rect 93 -1951 94 -1950
rect 432 -1951 433 -1950
rect 439 -1951 440 -1950
rect 625 -1951 626 -1950
rect 653 -1951 654 -1950
rect 674 -1951 675 -1950
rect 684 -1951 685 -1950
rect 751 -1951 752 -1950
rect 772 -1951 773 -1950
rect 779 -1951 780 -1950
rect 72 -1953 73 -1952
rect 107 -1953 108 -1952
rect 114 -1953 115 -1952
rect 142 -1953 143 -1952
rect 170 -1953 171 -1952
rect 177 -1953 178 -1952
rect 219 -1953 220 -1952
rect 289 -1953 290 -1952
rect 296 -1953 297 -1952
rect 604 -1953 605 -1952
rect 611 -1953 612 -1952
rect 751 -1953 752 -1952
rect 75 -1955 76 -1954
rect 107 -1955 108 -1954
rect 128 -1955 129 -1954
rect 184 -1955 185 -1954
rect 229 -1955 230 -1954
rect 261 -1955 262 -1954
rect 275 -1955 276 -1954
rect 334 -1955 335 -1954
rect 352 -1955 353 -1954
rect 387 -1955 388 -1954
rect 439 -1955 440 -1954
rect 464 -1955 465 -1954
rect 499 -1955 500 -1954
rect 695 -1955 696 -1954
rect 709 -1955 710 -1954
rect 786 -1955 787 -1954
rect 51 -1957 52 -1956
rect 229 -1957 230 -1956
rect 233 -1957 234 -1956
rect 268 -1957 269 -1956
rect 296 -1957 297 -1956
rect 474 -1957 475 -1956
rect 478 -1957 479 -1956
rect 499 -1957 500 -1956
rect 506 -1957 507 -1956
rect 548 -1957 549 -1956
rect 583 -1957 584 -1956
rect 611 -1957 612 -1956
rect 618 -1957 619 -1956
rect 758 -1957 759 -1956
rect 58 -1959 59 -1958
rect 128 -1959 129 -1958
rect 142 -1959 143 -1958
rect 194 -1959 195 -1958
rect 205 -1959 206 -1958
rect 261 -1959 262 -1958
rect 317 -1959 318 -1958
rect 464 -1959 465 -1958
rect 506 -1959 507 -1958
rect 513 -1959 514 -1958
rect 516 -1959 517 -1958
rect 772 -1959 773 -1958
rect 86 -1961 87 -1960
rect 219 -1961 220 -1960
rect 254 -1961 255 -1960
rect 331 -1961 332 -1960
rect 352 -1961 353 -1960
rect 408 -1961 409 -1960
rect 415 -1961 416 -1960
rect 709 -1961 710 -1960
rect 86 -1963 87 -1962
rect 282 -1963 283 -1962
rect 317 -1963 318 -1962
rect 345 -1963 346 -1962
rect 359 -1963 360 -1962
rect 373 -1963 374 -1962
rect 408 -1963 409 -1962
rect 422 -1963 423 -1962
rect 450 -1963 451 -1962
rect 555 -1963 556 -1962
rect 579 -1963 580 -1962
rect 618 -1963 619 -1962
rect 660 -1963 661 -1962
rect 667 -1963 668 -1962
rect 688 -1963 689 -1962
rect 765 -1963 766 -1962
rect 93 -1965 94 -1964
rect 180 -1965 181 -1964
rect 184 -1965 185 -1964
rect 310 -1965 311 -1964
rect 320 -1965 321 -1964
rect 401 -1965 402 -1964
rect 415 -1965 416 -1964
rect 460 -1965 461 -1964
rect 527 -1965 528 -1964
rect 541 -1965 542 -1964
rect 555 -1965 556 -1964
rect 562 -1965 563 -1964
rect 593 -1965 594 -1964
rect 730 -1965 731 -1964
rect 744 -1965 745 -1964
rect 765 -1965 766 -1964
rect 100 -1967 101 -1966
rect 156 -1967 157 -1966
rect 163 -1967 164 -1966
rect 170 -1967 171 -1966
rect 205 -1967 206 -1966
rect 226 -1967 227 -1966
rect 247 -1967 248 -1966
rect 254 -1967 255 -1966
rect 271 -1967 272 -1966
rect 450 -1967 451 -1966
rect 453 -1967 454 -1966
rect 737 -1967 738 -1966
rect 100 -1969 101 -1968
rect 135 -1969 136 -1968
rect 149 -1969 150 -1968
rect 268 -1969 269 -1968
rect 282 -1969 283 -1968
rect 492 -1969 493 -1968
rect 527 -1969 528 -1968
rect 726 -1969 727 -1968
rect 149 -1971 150 -1970
rect 222 -1971 223 -1970
rect 303 -1971 304 -1970
rect 359 -1971 360 -1970
rect 366 -1971 367 -1970
rect 478 -1971 479 -1970
rect 534 -1971 535 -1970
rect 590 -1971 591 -1970
rect 597 -1971 598 -1970
rect 604 -1971 605 -1970
rect 723 -1971 724 -1970
rect 737 -1971 738 -1970
rect 159 -1973 160 -1972
rect 303 -1973 304 -1972
rect 324 -1973 325 -1972
rect 345 -1973 346 -1972
rect 369 -1973 370 -1972
rect 534 -1973 535 -1972
rect 562 -1973 563 -1972
rect 639 -1973 640 -1972
rect 723 -1973 724 -1972
rect 793 -1973 794 -1972
rect 79 -1975 80 -1974
rect 324 -1975 325 -1974
rect 401 -1975 402 -1974
rect 485 -1975 486 -1974
rect 576 -1975 577 -1974
rect 744 -1975 745 -1974
rect 65 -1977 66 -1976
rect 79 -1977 80 -1976
rect 159 -1977 160 -1976
rect 163 -1977 164 -1976
rect 198 -1977 199 -1976
rect 247 -1977 248 -1976
rect 422 -1977 423 -1976
rect 502 -1977 503 -1976
rect 597 -1977 598 -1976
rect 646 -1977 647 -1976
rect 16 -1979 17 -1978
rect 65 -1979 66 -1978
rect 191 -1979 192 -1978
rect 198 -1979 199 -1978
rect 212 -1979 213 -1978
rect 233 -1979 234 -1978
rect 443 -1979 444 -1978
rect 485 -1979 486 -1978
rect 632 -1979 633 -1978
rect 639 -1979 640 -1978
rect 646 -1979 647 -1978
rect 674 -1979 675 -1978
rect 212 -1981 213 -1980
rect 240 -1981 241 -1980
rect 457 -1981 458 -1980
rect 520 -1981 521 -1980
rect 569 -1981 570 -1980
rect 632 -1981 633 -1980
rect 338 -1983 339 -1982
rect 457 -1983 458 -1982
rect 520 -1983 521 -1982
rect 681 -1983 682 -1982
rect 338 -1985 339 -1984
rect 380 -1985 381 -1984
rect 429 -1985 430 -1984
rect 569 -1985 570 -1984
rect 681 -1985 682 -1984
rect 702 -1985 703 -1984
rect 380 -1987 381 -1986
rect 471 -1987 472 -1986
rect 702 -1987 703 -1986
rect 716 -1987 717 -1986
rect 436 -1989 437 -1988
rect 716 -1989 717 -1988
rect 23 -1991 24 -1990
rect 436 -1991 437 -1990
rect 16 -2002 17 -2001
rect 93 -2002 94 -2001
rect 156 -2002 157 -2001
rect 187 -2002 188 -2001
rect 201 -2002 202 -2001
rect 226 -2002 227 -2001
rect 229 -2002 230 -2001
rect 338 -2002 339 -2001
rect 387 -2002 388 -2001
rect 404 -2002 405 -2001
rect 432 -2002 433 -2001
rect 569 -2002 570 -2001
rect 586 -2002 587 -2001
rect 639 -2002 640 -2001
rect 646 -2002 647 -2001
rect 663 -2002 664 -2001
rect 670 -2002 671 -2001
rect 786 -2002 787 -2001
rect 796 -2002 797 -2001
rect 814 -2002 815 -2001
rect 30 -2004 31 -2003
rect 79 -2004 80 -2003
rect 177 -2004 178 -2003
rect 310 -2004 311 -2003
rect 313 -2004 314 -2003
rect 324 -2004 325 -2003
rect 331 -2004 332 -2003
rect 397 -2004 398 -2003
rect 488 -2004 489 -2003
rect 513 -2004 514 -2003
rect 548 -2004 549 -2003
rect 779 -2004 780 -2003
rect 37 -2006 38 -2005
rect 149 -2006 150 -2005
rect 229 -2006 230 -2005
rect 268 -2006 269 -2005
rect 271 -2006 272 -2005
rect 359 -2006 360 -2005
rect 387 -2006 388 -2005
rect 492 -2006 493 -2005
rect 513 -2006 514 -2005
rect 632 -2006 633 -2005
rect 639 -2006 640 -2005
rect 695 -2006 696 -2005
rect 744 -2006 745 -2005
rect 807 -2006 808 -2005
rect 37 -2008 38 -2007
rect 184 -2008 185 -2007
rect 233 -2008 234 -2007
rect 240 -2008 241 -2007
rect 247 -2008 248 -2007
rect 380 -2008 381 -2007
rect 492 -2008 493 -2007
rect 555 -2008 556 -2007
rect 569 -2008 570 -2007
rect 793 -2008 794 -2007
rect 44 -2010 45 -2009
rect 198 -2010 199 -2009
rect 236 -2010 237 -2009
rect 548 -2010 549 -2009
rect 555 -2010 556 -2009
rect 618 -2010 619 -2009
rect 660 -2010 661 -2009
rect 702 -2010 703 -2009
rect 744 -2010 745 -2009
rect 751 -2010 752 -2009
rect 758 -2010 759 -2009
rect 786 -2010 787 -2009
rect 44 -2012 45 -2011
rect 107 -2012 108 -2011
rect 149 -2012 150 -2011
rect 170 -2012 171 -2011
rect 191 -2012 192 -2011
rect 198 -2012 199 -2011
rect 247 -2012 248 -2011
rect 254 -2012 255 -2011
rect 264 -2012 265 -2011
rect 632 -2012 633 -2011
rect 653 -2012 654 -2011
rect 660 -2012 661 -2011
rect 674 -2012 675 -2011
rect 695 -2012 696 -2011
rect 751 -2012 752 -2011
rect 772 -2012 773 -2011
rect 51 -2014 52 -2013
rect 166 -2014 167 -2013
rect 170 -2014 171 -2013
rect 257 -2014 258 -2013
rect 289 -2014 290 -2013
rect 352 -2014 353 -2013
rect 359 -2014 360 -2013
rect 373 -2014 374 -2013
rect 380 -2014 381 -2013
rect 408 -2014 409 -2013
rect 464 -2014 465 -2013
rect 674 -2014 675 -2013
rect 688 -2014 689 -2013
rect 730 -2014 731 -2013
rect 758 -2014 759 -2013
rect 765 -2014 766 -2013
rect 51 -2016 52 -2015
rect 590 -2016 591 -2015
rect 593 -2016 594 -2015
rect 800 -2016 801 -2015
rect 58 -2018 59 -2017
rect 243 -2018 244 -2017
rect 289 -2018 290 -2017
rect 348 -2018 349 -2017
rect 352 -2018 353 -2017
rect 422 -2018 423 -2017
rect 464 -2018 465 -2017
rect 478 -2018 479 -2017
rect 562 -2018 563 -2017
rect 618 -2018 619 -2017
rect 691 -2018 692 -2017
rect 737 -2018 738 -2017
rect 58 -2020 59 -2019
rect 114 -2020 115 -2019
rect 191 -2020 192 -2019
rect 212 -2020 213 -2019
rect 243 -2020 244 -2019
rect 282 -2020 283 -2019
rect 292 -2020 293 -2019
rect 432 -2020 433 -2019
rect 471 -2020 472 -2019
rect 702 -2020 703 -2019
rect 716 -2020 717 -2019
rect 730 -2020 731 -2019
rect 65 -2022 66 -2021
rect 233 -2022 234 -2021
rect 296 -2022 297 -2021
rect 366 -2022 367 -2021
rect 373 -2022 374 -2021
rect 450 -2022 451 -2021
rect 565 -2022 566 -2021
rect 737 -2022 738 -2021
rect 65 -2024 66 -2023
rect 460 -2024 461 -2023
rect 583 -2024 584 -2023
rect 653 -2024 654 -2023
rect 709 -2024 710 -2023
rect 716 -2024 717 -2023
rect 72 -2026 73 -2025
rect 135 -2026 136 -2025
rect 163 -2026 164 -2025
rect 296 -2026 297 -2025
rect 303 -2026 304 -2025
rect 436 -2026 437 -2025
rect 450 -2026 451 -2025
rect 597 -2026 598 -2025
rect 681 -2026 682 -2025
rect 709 -2026 710 -2025
rect 72 -2028 73 -2027
rect 100 -2028 101 -2027
rect 107 -2028 108 -2027
rect 254 -2028 255 -2027
rect 303 -2028 304 -2027
rect 474 -2028 475 -2027
rect 541 -2028 542 -2027
rect 597 -2028 598 -2027
rect 667 -2028 668 -2027
rect 681 -2028 682 -2027
rect 79 -2030 80 -2029
rect 317 -2030 318 -2029
rect 324 -2030 325 -2029
rect 394 -2030 395 -2029
rect 401 -2030 402 -2029
rect 765 -2030 766 -2029
rect 86 -2032 87 -2031
rect 135 -2032 136 -2031
rect 219 -2032 220 -2031
rect 282 -2032 283 -2031
rect 317 -2032 318 -2031
rect 457 -2032 458 -2031
rect 527 -2032 528 -2031
rect 541 -2032 542 -2031
rect 583 -2032 584 -2031
rect 611 -2032 612 -2031
rect 646 -2032 647 -2031
rect 667 -2032 668 -2031
rect 86 -2034 87 -2033
rect 520 -2034 521 -2033
rect 590 -2034 591 -2033
rect 726 -2034 727 -2033
rect 100 -2036 101 -2035
rect 121 -2036 122 -2035
rect 128 -2036 129 -2035
rect 212 -2036 213 -2035
rect 261 -2036 262 -2035
rect 527 -2036 528 -2035
rect 611 -2036 612 -2035
rect 677 -2036 678 -2035
rect 23 -2038 24 -2037
rect 128 -2038 129 -2037
rect 205 -2038 206 -2037
rect 219 -2038 220 -2037
rect 261 -2038 262 -2037
rect 345 -2038 346 -2037
rect 394 -2038 395 -2037
rect 772 -2038 773 -2037
rect 114 -2040 115 -2039
rect 142 -2040 143 -2039
rect 205 -2040 206 -2039
rect 446 -2040 447 -2039
rect 457 -2040 458 -2039
rect 604 -2040 605 -2039
rect 93 -2042 94 -2041
rect 142 -2042 143 -2041
rect 331 -2042 332 -2041
rect 401 -2042 402 -2041
rect 408 -2042 409 -2041
rect 415 -2042 416 -2041
rect 418 -2042 419 -2041
rect 604 -2042 605 -2041
rect 121 -2044 122 -2043
rect 184 -2044 185 -2043
rect 338 -2044 339 -2043
rect 600 -2044 601 -2043
rect 345 -2046 346 -2045
rect 443 -2046 444 -2045
rect 506 -2046 507 -2045
rect 520 -2046 521 -2045
rect 415 -2048 416 -2047
rect 534 -2048 535 -2047
rect 422 -2050 423 -2049
rect 499 -2050 500 -2049
rect 429 -2052 430 -2051
rect 443 -2052 444 -2051
rect 478 -2052 479 -2051
rect 499 -2052 500 -2051
rect 485 -2054 486 -2053
rect 534 -2054 535 -2053
rect 23 -2065 24 -2064
rect 397 -2065 398 -2064
rect 411 -2065 412 -2064
rect 513 -2065 514 -2064
rect 534 -2065 535 -2064
rect 537 -2065 538 -2064
rect 541 -2065 542 -2064
rect 593 -2065 594 -2064
rect 653 -2065 654 -2064
rect 737 -2065 738 -2064
rect 23 -2067 24 -2066
rect 240 -2067 241 -2066
rect 254 -2067 255 -2066
rect 282 -2067 283 -2066
rect 292 -2067 293 -2066
rect 366 -2067 367 -2066
rect 373 -2067 374 -2066
rect 401 -2067 402 -2066
rect 418 -2067 419 -2066
rect 499 -2067 500 -2066
rect 534 -2067 535 -2066
rect 555 -2067 556 -2066
rect 569 -2067 570 -2066
rect 632 -2067 633 -2066
rect 667 -2067 668 -2066
rect 681 -2067 682 -2066
rect 723 -2067 724 -2066
rect 758 -2067 759 -2066
rect 30 -2069 31 -2068
rect 145 -2069 146 -2068
rect 184 -2069 185 -2068
rect 236 -2069 237 -2068
rect 240 -2069 241 -2068
rect 275 -2069 276 -2068
rect 345 -2069 346 -2068
rect 422 -2069 423 -2068
rect 436 -2069 437 -2068
rect 513 -2069 514 -2068
rect 537 -2069 538 -2068
rect 555 -2069 556 -2068
rect 569 -2069 570 -2068
rect 583 -2069 584 -2068
rect 632 -2069 633 -2068
rect 646 -2069 647 -2068
rect 670 -2069 671 -2068
rect 786 -2069 787 -2068
rect 30 -2071 31 -2070
rect 471 -2071 472 -2070
rect 474 -2071 475 -2070
rect 618 -2071 619 -2070
rect 646 -2071 647 -2070
rect 730 -2071 731 -2070
rect 37 -2073 38 -2072
rect 229 -2073 230 -2072
rect 257 -2073 258 -2072
rect 429 -2073 430 -2072
rect 457 -2073 458 -2072
rect 779 -2073 780 -2072
rect 44 -2075 45 -2074
rect 177 -2075 178 -2074
rect 212 -2075 213 -2074
rect 282 -2075 283 -2074
rect 296 -2075 297 -2074
rect 422 -2075 423 -2074
rect 457 -2075 458 -2074
rect 583 -2075 584 -2074
rect 618 -2075 619 -2074
rect 660 -2075 661 -2074
rect 681 -2075 682 -2074
rect 772 -2075 773 -2074
rect 44 -2077 45 -2076
rect 170 -2077 171 -2076
rect 212 -2077 213 -2076
rect 348 -2077 349 -2076
rect 352 -2077 353 -2076
rect 562 -2077 563 -2076
rect 660 -2077 661 -2076
rect 674 -2077 675 -2076
rect 709 -2077 710 -2076
rect 723 -2077 724 -2076
rect 726 -2077 727 -2076
rect 737 -2077 738 -2076
rect 51 -2079 52 -2078
rect 124 -2079 125 -2078
rect 135 -2079 136 -2078
rect 177 -2079 178 -2078
rect 219 -2079 220 -2078
rect 254 -2079 255 -2078
rect 275 -2079 276 -2078
rect 310 -2079 311 -2078
rect 324 -2079 325 -2078
rect 352 -2079 353 -2078
rect 373 -2079 374 -2078
rect 485 -2079 486 -2078
rect 488 -2079 489 -2078
rect 492 -2079 493 -2078
rect 499 -2079 500 -2078
rect 590 -2079 591 -2078
rect 709 -2079 710 -2078
rect 751 -2079 752 -2078
rect 51 -2081 52 -2080
rect 149 -2081 150 -2080
rect 268 -2081 269 -2080
rect 310 -2081 311 -2080
rect 317 -2081 318 -2080
rect 324 -2081 325 -2080
rect 359 -2081 360 -2080
rect 485 -2081 486 -2080
rect 492 -2081 493 -2080
rect 548 -2081 549 -2080
rect 562 -2081 563 -2080
rect 597 -2081 598 -2080
rect 58 -2083 59 -2082
rect 131 -2083 132 -2082
rect 135 -2083 136 -2082
rect 338 -2083 339 -2082
rect 380 -2083 381 -2082
rect 415 -2083 416 -2082
rect 464 -2083 465 -2082
rect 509 -2083 510 -2082
rect 527 -2083 528 -2082
rect 674 -2083 675 -2082
rect 58 -2085 59 -2084
rect 128 -2085 129 -2084
rect 142 -2085 143 -2084
rect 362 -2085 363 -2084
rect 366 -2085 367 -2084
rect 464 -2085 465 -2084
rect 474 -2085 475 -2084
rect 576 -2085 577 -2084
rect 65 -2087 66 -2086
rect 138 -2087 139 -2086
rect 142 -2087 143 -2086
rect 156 -2087 157 -2086
rect 233 -2087 234 -2086
rect 268 -2087 269 -2086
rect 296 -2087 297 -2086
rect 331 -2087 332 -2086
rect 338 -2087 339 -2086
rect 460 -2087 461 -2086
rect 478 -2087 479 -2086
rect 702 -2087 703 -2086
rect 65 -2089 66 -2088
rect 243 -2089 244 -2088
rect 317 -2089 318 -2088
rect 597 -2089 598 -2088
rect 688 -2089 689 -2088
rect 702 -2089 703 -2088
rect 72 -2091 73 -2090
rect 103 -2091 104 -2090
rect 107 -2091 108 -2090
rect 184 -2091 185 -2090
rect 233 -2091 234 -2090
rect 289 -2091 290 -2090
rect 331 -2091 332 -2090
rect 387 -2091 388 -2090
rect 415 -2091 416 -2090
rect 450 -2091 451 -2090
rect 460 -2091 461 -2090
rect 765 -2091 766 -2090
rect 72 -2093 73 -2092
rect 261 -2093 262 -2092
rect 320 -2093 321 -2092
rect 450 -2093 451 -2092
rect 478 -2093 479 -2092
rect 516 -2093 517 -2092
rect 520 -2093 521 -2092
rect 527 -2093 528 -2092
rect 576 -2093 577 -2092
rect 625 -2093 626 -2092
rect 688 -2093 689 -2092
rect 716 -2093 717 -2092
rect 79 -2095 80 -2094
rect 439 -2095 440 -2094
rect 506 -2095 507 -2094
rect 548 -2095 549 -2094
rect 625 -2095 626 -2094
rect 639 -2095 640 -2094
rect 716 -2095 717 -2094
rect 744 -2095 745 -2094
rect 79 -2097 80 -2096
rect 173 -2097 174 -2096
rect 247 -2097 248 -2096
rect 289 -2097 290 -2096
rect 387 -2097 388 -2096
rect 506 -2097 507 -2096
rect 520 -2097 521 -2096
rect 604 -2097 605 -2096
rect 86 -2099 87 -2098
rect 187 -2099 188 -2098
rect 261 -2099 262 -2098
rect 432 -2099 433 -2098
rect 604 -2099 605 -2098
rect 695 -2099 696 -2098
rect 86 -2101 87 -2100
rect 96 -2101 97 -2100
rect 100 -2101 101 -2100
rect 107 -2101 108 -2100
rect 121 -2101 122 -2100
rect 303 -2101 304 -2100
rect 394 -2101 395 -2100
rect 639 -2101 640 -2100
rect 93 -2103 94 -2102
rect 229 -2103 230 -2102
rect 303 -2103 304 -2102
rect 383 -2103 384 -2102
rect 394 -2103 395 -2102
rect 408 -2103 409 -2102
rect 16 -2105 17 -2104
rect 93 -2105 94 -2104
rect 128 -2105 129 -2104
rect 541 -2105 542 -2104
rect 149 -2107 150 -2106
rect 191 -2107 192 -2106
rect 163 -2109 164 -2108
rect 247 -2109 248 -2108
rect 156 -2111 157 -2110
rect 163 -2111 164 -2110
rect 180 -2111 181 -2110
rect 695 -2111 696 -2110
rect 180 -2113 181 -2112
rect 198 -2113 199 -2112
rect 191 -2115 192 -2114
rect 205 -2115 206 -2114
rect 16 -2117 17 -2116
rect 205 -2117 206 -2116
rect 198 -2119 199 -2118
rect 219 -2119 220 -2118
rect 16 -2130 17 -2129
rect 474 -2130 475 -2129
rect 506 -2130 507 -2129
rect 625 -2130 626 -2129
rect 688 -2130 689 -2129
rect 698 -2130 699 -2129
rect 40 -2132 41 -2131
rect 152 -2132 153 -2131
rect 163 -2132 164 -2131
rect 173 -2132 174 -2131
rect 184 -2132 185 -2131
rect 254 -2132 255 -2131
rect 261 -2132 262 -2131
rect 453 -2132 454 -2131
rect 457 -2132 458 -2131
rect 688 -2132 689 -2131
rect 695 -2132 696 -2131
rect 730 -2132 731 -2131
rect 44 -2134 45 -2133
rect 229 -2134 230 -2133
rect 254 -2134 255 -2133
rect 338 -2134 339 -2133
rect 345 -2134 346 -2133
rect 597 -2134 598 -2133
rect 625 -2134 626 -2133
rect 709 -2134 710 -2133
rect 51 -2136 52 -2135
rect 219 -2136 220 -2135
rect 226 -2136 227 -2135
rect 240 -2136 241 -2135
rect 261 -2136 262 -2135
rect 352 -2136 353 -2135
rect 359 -2136 360 -2135
rect 429 -2136 430 -2135
rect 436 -2136 437 -2135
rect 467 -2136 468 -2135
rect 509 -2136 510 -2135
rect 541 -2136 542 -2135
rect 558 -2136 559 -2135
rect 716 -2136 717 -2135
rect 58 -2138 59 -2137
rect 100 -2138 101 -2137
rect 121 -2138 122 -2137
rect 247 -2138 248 -2137
rect 268 -2138 269 -2137
rect 345 -2138 346 -2137
rect 348 -2138 349 -2137
rect 411 -2138 412 -2137
rect 439 -2138 440 -2137
rect 611 -2138 612 -2137
rect 660 -2138 661 -2137
rect 716 -2138 717 -2137
rect 65 -2140 66 -2139
rect 320 -2140 321 -2139
rect 324 -2140 325 -2139
rect 352 -2140 353 -2139
rect 380 -2140 381 -2139
rect 394 -2140 395 -2139
rect 408 -2140 409 -2139
rect 513 -2140 514 -2139
rect 534 -2140 535 -2139
rect 709 -2140 710 -2139
rect 72 -2142 73 -2141
rect 334 -2142 335 -2141
rect 362 -2142 363 -2141
rect 380 -2142 381 -2141
rect 390 -2142 391 -2141
rect 492 -2142 493 -2141
rect 513 -2142 514 -2141
rect 520 -2142 521 -2141
rect 541 -2142 542 -2141
rect 548 -2142 549 -2141
rect 579 -2142 580 -2141
rect 702 -2142 703 -2141
rect 100 -2144 101 -2143
rect 114 -2144 115 -2143
rect 128 -2144 129 -2143
rect 156 -2144 157 -2143
rect 170 -2144 171 -2143
rect 415 -2144 416 -2143
rect 464 -2144 465 -2143
rect 562 -2144 563 -2143
rect 583 -2144 584 -2143
rect 590 -2144 591 -2143
rect 593 -2144 594 -2143
rect 695 -2144 696 -2143
rect 30 -2146 31 -2145
rect 128 -2146 129 -2145
rect 135 -2146 136 -2145
rect 163 -2146 164 -2145
rect 198 -2146 199 -2145
rect 450 -2146 451 -2145
rect 464 -2146 465 -2145
rect 499 -2146 500 -2145
rect 520 -2146 521 -2145
rect 527 -2146 528 -2145
rect 548 -2146 549 -2145
rect 569 -2146 570 -2145
rect 597 -2146 598 -2145
rect 604 -2146 605 -2145
rect 611 -2146 612 -2145
rect 653 -2146 654 -2145
rect 107 -2148 108 -2147
rect 135 -2148 136 -2147
rect 142 -2148 143 -2147
rect 159 -2148 160 -2147
rect 198 -2148 199 -2147
rect 222 -2148 223 -2147
rect 226 -2148 227 -2147
rect 268 -2148 269 -2147
rect 282 -2148 283 -2147
rect 289 -2148 290 -2147
rect 296 -2148 297 -2147
rect 338 -2148 339 -2147
rect 373 -2148 374 -2147
rect 394 -2148 395 -2147
rect 408 -2148 409 -2147
rect 534 -2148 535 -2147
rect 555 -2148 556 -2147
rect 702 -2148 703 -2147
rect 23 -2150 24 -2149
rect 159 -2150 160 -2149
rect 170 -2150 171 -2149
rect 555 -2150 556 -2149
rect 604 -2150 605 -2149
rect 618 -2150 619 -2149
rect 639 -2150 640 -2149
rect 660 -2150 661 -2149
rect 107 -2152 108 -2151
rect 177 -2152 178 -2151
rect 201 -2152 202 -2151
rect 275 -2152 276 -2151
rect 282 -2152 283 -2151
rect 324 -2152 325 -2151
rect 331 -2152 332 -2151
rect 429 -2152 430 -2151
rect 471 -2152 472 -2151
rect 562 -2152 563 -2151
rect 639 -2152 640 -2151
rect 681 -2152 682 -2151
rect 114 -2154 115 -2153
rect 285 -2154 286 -2153
rect 296 -2154 297 -2153
rect 387 -2154 388 -2153
rect 443 -2154 444 -2153
rect 471 -2154 472 -2153
rect 485 -2154 486 -2153
rect 618 -2154 619 -2153
rect 646 -2154 647 -2153
rect 653 -2154 654 -2153
rect 121 -2156 122 -2155
rect 387 -2156 388 -2155
rect 443 -2156 444 -2155
rect 478 -2156 479 -2155
rect 499 -2156 500 -2155
rect 509 -2156 510 -2155
rect 646 -2156 647 -2155
rect 674 -2156 675 -2155
rect 142 -2158 143 -2157
rect 233 -2158 234 -2157
rect 275 -2158 276 -2157
rect 303 -2158 304 -2157
rect 313 -2158 314 -2157
rect 737 -2158 738 -2157
rect 149 -2160 150 -2159
rect 205 -2160 206 -2159
rect 212 -2160 213 -2159
rect 233 -2160 234 -2159
rect 303 -2160 304 -2159
rect 310 -2160 311 -2159
rect 331 -2160 332 -2159
rect 527 -2160 528 -2159
rect 667 -2160 668 -2159
rect 674 -2160 675 -2159
rect 79 -2162 80 -2161
rect 212 -2162 213 -2161
rect 219 -2162 220 -2161
rect 415 -2162 416 -2161
rect 478 -2162 479 -2161
rect 569 -2162 570 -2161
rect 667 -2162 668 -2161
rect 723 -2162 724 -2161
rect 156 -2164 157 -2163
rect 310 -2164 311 -2163
rect 366 -2164 367 -2163
rect 485 -2164 486 -2163
rect 576 -2164 577 -2163
rect 723 -2164 724 -2163
rect 177 -2166 178 -2165
rect 180 -2166 181 -2165
rect 191 -2166 192 -2165
rect 205 -2166 206 -2165
rect 222 -2166 223 -2165
rect 317 -2166 318 -2165
rect 366 -2166 367 -2165
rect 422 -2166 423 -2165
rect 191 -2168 192 -2167
rect 208 -2168 209 -2167
rect 373 -2168 374 -2167
rect 401 -2168 402 -2167
rect 422 -2168 423 -2167
rect 576 -2168 577 -2167
rect 250 -2170 251 -2169
rect 401 -2170 402 -2169
rect 86 -2181 87 -2180
rect 89 -2181 90 -2180
rect 114 -2181 115 -2180
rect 306 -2181 307 -2180
rect 380 -2181 381 -2180
rect 492 -2181 493 -2180
rect 506 -2181 507 -2180
rect 527 -2181 528 -2180
rect 534 -2181 535 -2180
rect 670 -2181 671 -2180
rect 674 -2181 675 -2180
rect 681 -2181 682 -2180
rect 114 -2183 115 -2182
rect 184 -2183 185 -2182
rect 205 -2183 206 -2182
rect 219 -2183 220 -2182
rect 222 -2183 223 -2182
rect 576 -2183 577 -2182
rect 579 -2183 580 -2182
rect 723 -2183 724 -2182
rect 121 -2185 122 -2184
rect 149 -2185 150 -2184
rect 163 -2185 164 -2184
rect 184 -2185 185 -2184
rect 205 -2185 206 -2184
rect 299 -2185 300 -2184
rect 324 -2185 325 -2184
rect 380 -2185 381 -2184
rect 401 -2185 402 -2184
rect 460 -2185 461 -2184
rect 492 -2185 493 -2184
rect 558 -2185 559 -2184
rect 569 -2185 570 -2184
rect 716 -2185 717 -2184
rect 124 -2187 125 -2186
rect 254 -2187 255 -2186
rect 282 -2187 283 -2186
rect 366 -2187 367 -2186
rect 401 -2187 402 -2186
rect 422 -2187 423 -2186
rect 425 -2187 426 -2186
rect 562 -2187 563 -2186
rect 583 -2187 584 -2186
rect 688 -2187 689 -2186
rect 128 -2189 129 -2188
rect 411 -2189 412 -2188
rect 429 -2189 430 -2188
rect 618 -2189 619 -2188
rect 639 -2189 640 -2188
rect 667 -2189 668 -2188
rect 142 -2191 143 -2190
rect 219 -2191 220 -2190
rect 240 -2191 241 -2190
rect 513 -2191 514 -2190
rect 555 -2191 556 -2190
rect 611 -2191 612 -2190
rect 170 -2193 171 -2192
rect 240 -2193 241 -2192
rect 243 -2193 244 -2192
rect 254 -2193 255 -2192
rect 285 -2193 286 -2192
rect 390 -2193 391 -2192
rect 394 -2193 395 -2192
rect 562 -2193 563 -2192
rect 569 -2193 570 -2192
rect 618 -2193 619 -2192
rect 142 -2195 143 -2194
rect 170 -2195 171 -2194
rect 198 -2195 199 -2194
rect 394 -2195 395 -2194
rect 408 -2195 409 -2194
rect 443 -2195 444 -2194
rect 450 -2195 451 -2194
rect 464 -2195 465 -2194
rect 499 -2195 500 -2194
rect 527 -2195 528 -2194
rect 555 -2195 556 -2194
rect 632 -2195 633 -2194
rect 212 -2197 213 -2196
rect 345 -2197 346 -2196
rect 366 -2197 367 -2196
rect 373 -2197 374 -2196
rect 387 -2197 388 -2196
rect 464 -2197 465 -2196
rect 513 -2197 514 -2196
rect 548 -2197 549 -2196
rect 583 -2197 584 -2196
rect 653 -2197 654 -2196
rect 152 -2199 153 -2198
rect 212 -2199 213 -2198
rect 285 -2199 286 -2198
rect 450 -2199 451 -2198
rect 548 -2199 549 -2198
rect 590 -2199 591 -2198
rect 597 -2199 598 -2198
rect 639 -2199 640 -2198
rect 296 -2201 297 -2200
rect 614 -2201 615 -2200
rect 632 -2201 633 -2200
rect 702 -2201 703 -2200
rect 317 -2203 318 -2202
rect 345 -2203 346 -2202
rect 415 -2203 416 -2202
rect 499 -2203 500 -2202
rect 586 -2203 587 -2202
rect 604 -2203 605 -2202
rect 317 -2205 318 -2204
rect 471 -2205 472 -2204
rect 509 -2205 510 -2204
rect 604 -2205 605 -2204
rect 324 -2207 325 -2206
rect 352 -2207 353 -2206
rect 359 -2207 360 -2206
rect 415 -2207 416 -2206
rect 429 -2207 430 -2206
rect 478 -2207 479 -2206
rect 590 -2207 591 -2206
rect 625 -2207 626 -2206
rect 268 -2209 269 -2208
rect 352 -2209 353 -2208
rect 432 -2209 433 -2208
rect 457 -2209 458 -2208
rect 478 -2209 479 -2208
rect 621 -2209 622 -2208
rect 268 -2211 269 -2210
rect 310 -2211 311 -2210
rect 331 -2211 332 -2210
rect 471 -2211 472 -2210
rect 485 -2211 486 -2210
rect 625 -2211 626 -2210
rect 261 -2213 262 -2212
rect 331 -2213 332 -2212
rect 436 -2213 437 -2212
rect 534 -2213 535 -2212
rect 597 -2213 598 -2212
rect 646 -2213 647 -2212
rect 261 -2215 262 -2214
rect 338 -2215 339 -2214
rect 390 -2215 391 -2214
rect 436 -2215 437 -2214
rect 485 -2215 486 -2214
rect 520 -2215 521 -2214
rect 156 -2217 157 -2216
rect 338 -2217 339 -2216
rect 520 -2217 521 -2216
rect 541 -2217 542 -2216
rect 156 -2219 157 -2218
rect 177 -2219 178 -2218
rect 289 -2219 290 -2218
rect 310 -2219 311 -2218
rect 541 -2219 542 -2218
rect 660 -2219 661 -2218
rect 131 -2221 132 -2220
rect 177 -2221 178 -2220
rect 247 -2221 248 -2220
rect 289 -2221 290 -2220
rect 660 -2221 661 -2220
rect 709 -2221 710 -2220
rect 100 -2223 101 -2222
rect 131 -2223 132 -2222
rect 247 -2223 248 -2222
rect 303 -2223 304 -2222
rect 107 -2234 108 -2233
rect 229 -2234 230 -2233
rect 275 -2234 276 -2233
rect 282 -2234 283 -2233
rect 306 -2234 307 -2233
rect 478 -2234 479 -2233
rect 534 -2234 535 -2233
rect 611 -2234 612 -2233
rect 114 -2236 115 -2235
rect 194 -2236 195 -2235
rect 198 -2236 199 -2235
rect 236 -2236 237 -2235
rect 254 -2236 255 -2235
rect 275 -2236 276 -2235
rect 313 -2236 314 -2235
rect 401 -2236 402 -2235
rect 415 -2236 416 -2235
rect 425 -2236 426 -2235
rect 443 -2236 444 -2235
rect 478 -2236 479 -2235
rect 527 -2236 528 -2235
rect 534 -2236 535 -2235
rect 562 -2236 563 -2235
rect 590 -2236 591 -2235
rect 607 -2236 608 -2235
rect 660 -2236 661 -2235
rect 114 -2238 115 -2237
rect 142 -2238 143 -2237
rect 149 -2238 150 -2237
rect 170 -2238 171 -2237
rect 173 -2238 174 -2237
rect 191 -2238 192 -2237
rect 201 -2238 202 -2237
rect 212 -2238 213 -2237
rect 219 -2238 220 -2237
rect 254 -2238 255 -2237
rect 324 -2238 325 -2237
rect 359 -2238 360 -2237
rect 366 -2238 367 -2237
rect 376 -2238 377 -2237
rect 390 -2238 391 -2237
rect 415 -2238 416 -2237
rect 422 -2238 423 -2237
rect 429 -2238 430 -2237
rect 446 -2238 447 -2237
rect 541 -2238 542 -2237
rect 565 -2238 566 -2237
rect 632 -2238 633 -2237
rect 121 -2240 122 -2239
rect 124 -2240 125 -2239
rect 128 -2240 129 -2239
rect 138 -2240 139 -2239
rect 149 -2240 150 -2239
rect 208 -2240 209 -2239
rect 212 -2240 213 -2239
rect 219 -2240 220 -2239
rect 261 -2240 262 -2239
rect 324 -2240 325 -2239
rect 327 -2240 328 -2239
rect 362 -2240 363 -2239
rect 366 -2240 367 -2239
rect 380 -2240 381 -2239
rect 397 -2240 398 -2239
rect 471 -2240 472 -2239
rect 513 -2240 514 -2239
rect 541 -2240 542 -2239
rect 124 -2242 125 -2241
rect 145 -2242 146 -2241
rect 156 -2242 157 -2241
rect 191 -2242 192 -2241
rect 205 -2242 206 -2241
rect 306 -2242 307 -2241
rect 331 -2242 332 -2241
rect 390 -2242 391 -2241
rect 401 -2242 402 -2241
rect 408 -2242 409 -2241
rect 464 -2242 465 -2241
rect 520 -2242 521 -2241
rect 527 -2242 528 -2241
rect 555 -2242 556 -2241
rect 131 -2244 132 -2243
rect 135 -2244 136 -2243
rect 156 -2244 157 -2243
rect 177 -2244 178 -2243
rect 261 -2244 262 -2243
rect 408 -2244 409 -2243
rect 467 -2244 468 -2243
rect 506 -2244 507 -2243
rect 513 -2244 514 -2243
rect 576 -2244 577 -2243
rect 163 -2246 164 -2245
rect 268 -2246 269 -2245
rect 296 -2246 297 -2245
rect 331 -2246 332 -2245
rect 338 -2246 339 -2245
rect 565 -2246 566 -2245
rect 576 -2246 577 -2245
rect 597 -2246 598 -2245
rect 163 -2248 164 -2247
rect 180 -2248 181 -2247
rect 247 -2248 248 -2247
rect 296 -2248 297 -2247
rect 310 -2248 311 -2247
rect 338 -2248 339 -2247
rect 345 -2248 346 -2247
rect 464 -2248 465 -2247
rect 492 -2248 493 -2247
rect 520 -2248 521 -2247
rect 555 -2248 556 -2247
rect 569 -2248 570 -2247
rect 166 -2250 167 -2249
rect 432 -2250 433 -2249
rect 485 -2250 486 -2249
rect 492 -2250 493 -2249
rect 506 -2250 507 -2249
rect 579 -2250 580 -2249
rect 177 -2252 178 -2251
rect 184 -2252 185 -2251
rect 240 -2252 241 -2251
rect 247 -2252 248 -2251
rect 268 -2252 269 -2251
rect 282 -2252 283 -2251
rect 303 -2252 304 -2251
rect 345 -2252 346 -2251
rect 359 -2252 360 -2251
rect 443 -2252 444 -2251
rect 184 -2254 185 -2253
rect 240 -2254 241 -2253
rect 373 -2254 374 -2253
rect 436 -2254 437 -2253
rect 352 -2256 353 -2255
rect 373 -2256 374 -2255
rect 394 -2256 395 -2255
rect 485 -2256 486 -2255
rect 226 -2258 227 -2257
rect 352 -2258 353 -2257
rect 380 -2258 381 -2257
rect 394 -2258 395 -2257
rect 436 -2258 437 -2257
rect 450 -2258 451 -2257
rect 226 -2260 227 -2259
rect 233 -2260 234 -2259
rect 303 -2260 304 -2259
rect 450 -2260 451 -2259
rect 114 -2271 115 -2270
rect 131 -2271 132 -2270
rect 135 -2271 136 -2270
rect 145 -2271 146 -2270
rect 163 -2271 164 -2270
rect 306 -2271 307 -2270
rect 317 -2271 318 -2270
rect 373 -2271 374 -2270
rect 401 -2271 402 -2270
rect 439 -2271 440 -2270
rect 450 -2271 451 -2270
rect 572 -2271 573 -2270
rect 121 -2273 122 -2272
rect 124 -2273 125 -2272
rect 142 -2273 143 -2272
rect 156 -2273 157 -2272
rect 170 -2273 171 -2272
rect 212 -2273 213 -2272
rect 215 -2273 216 -2272
rect 222 -2273 223 -2272
rect 240 -2273 241 -2272
rect 250 -2273 251 -2272
rect 275 -2273 276 -2272
rect 282 -2273 283 -2272
rect 289 -2273 290 -2272
rect 310 -2273 311 -2272
rect 352 -2273 353 -2272
rect 387 -2273 388 -2272
rect 404 -2273 405 -2272
rect 415 -2273 416 -2272
rect 429 -2273 430 -2272
rect 530 -2273 531 -2272
rect 541 -2273 542 -2272
rect 569 -2273 570 -2272
rect 184 -2275 185 -2274
rect 233 -2275 234 -2274
rect 243 -2275 244 -2274
rect 478 -2275 479 -2274
rect 485 -2275 486 -2274
rect 502 -2275 503 -2274
rect 534 -2275 535 -2274
rect 541 -2275 542 -2274
rect 198 -2277 199 -2276
rect 313 -2277 314 -2276
rect 359 -2277 360 -2276
rect 464 -2277 465 -2276
rect 471 -2277 472 -2276
rect 499 -2277 500 -2276
rect 534 -2277 535 -2276
rect 555 -2277 556 -2276
rect 212 -2279 213 -2278
rect 219 -2279 220 -2278
rect 226 -2279 227 -2278
rect 233 -2279 234 -2278
rect 261 -2279 262 -2278
rect 275 -2279 276 -2278
rect 289 -2279 290 -2278
rect 317 -2279 318 -2278
rect 408 -2279 409 -2278
rect 520 -2279 521 -2278
rect 205 -2281 206 -2280
rect 226 -2281 227 -2280
rect 268 -2281 269 -2280
rect 282 -2281 283 -2280
rect 303 -2281 304 -2280
rect 331 -2281 332 -2280
rect 415 -2281 416 -2280
rect 436 -2281 437 -2280
rect 457 -2281 458 -2280
rect 464 -2281 465 -2280
rect 474 -2281 475 -2280
rect 478 -2281 479 -2280
rect 513 -2281 514 -2280
rect 520 -2281 521 -2280
rect 247 -2283 248 -2282
rect 268 -2283 269 -2282
rect 303 -2283 304 -2282
rect 366 -2283 367 -2282
rect 432 -2283 433 -2282
rect 506 -2283 507 -2282
rect 513 -2283 514 -2282
rect 527 -2283 528 -2282
rect 331 -2285 332 -2284
rect 338 -2285 339 -2284
rect 362 -2285 363 -2284
rect 366 -2285 367 -2284
rect 443 -2285 444 -2284
rect 457 -2285 458 -2284
rect 492 -2285 493 -2284
rect 506 -2285 507 -2284
rect 527 -2285 528 -2284
rect 576 -2285 577 -2284
rect 450 -2287 451 -2286
rect 474 -2287 475 -2286
rect 576 -2287 577 -2286
rect 583 -2287 584 -2286
rect 212 -2298 213 -2297
rect 215 -2298 216 -2297
rect 226 -2298 227 -2297
rect 243 -2298 244 -2297
rect 247 -2298 248 -2297
rect 254 -2298 255 -2297
rect 275 -2298 276 -2297
rect 327 -2298 328 -2297
rect 338 -2298 339 -2297
rect 345 -2298 346 -2297
rect 366 -2298 367 -2297
rect 369 -2298 370 -2297
rect 408 -2298 409 -2297
rect 415 -2298 416 -2297
rect 422 -2298 423 -2297
rect 439 -2298 440 -2297
rect 443 -2298 444 -2297
rect 464 -2298 465 -2297
rect 502 -2298 503 -2297
rect 513 -2298 514 -2297
rect 520 -2298 521 -2297
rect 527 -2298 528 -2297
rect 534 -2298 535 -2297
rect 541 -2298 542 -2297
rect 569 -2298 570 -2297
rect 576 -2298 577 -2297
rect 597 -2298 598 -2297
rect 604 -2298 605 -2297
rect 639 -2298 640 -2297
rect 646 -2298 647 -2297
rect 226 -2300 227 -2299
rect 264 -2300 265 -2299
rect 282 -2300 283 -2299
rect 289 -2300 290 -2299
rect 296 -2300 297 -2299
rect 306 -2300 307 -2299
rect 313 -2300 314 -2299
rect 317 -2300 318 -2299
rect 432 -2300 433 -2299
rect 457 -2300 458 -2299
rect 506 -2300 507 -2299
rect 509 -2300 510 -2299
rect 614 -2300 615 -2299
rect 639 -2300 640 -2299
rect 254 -2302 255 -2301
rect 285 -2302 286 -2301
rect 289 -2302 290 -2301
rect 310 -2302 311 -2301
rect 317 -2302 318 -2301
rect 331 -2302 332 -2301
rect 446 -2302 447 -2301
rect 450 -2302 451 -2301
rect 268 -2304 269 -2303
rect 296 -2304 297 -2303
rect 170 -2315 171 -2314
rect 177 -2315 178 -2314
rect 226 -2315 227 -2314
rect 282 -2315 283 -2314
rect 296 -2315 297 -2314
rect 306 -2315 307 -2314
rect 380 -2315 381 -2314
rect 387 -2315 388 -2314
rect 404 -2315 405 -2314
rect 408 -2315 409 -2314
rect 527 -2315 528 -2314
rect 534 -2315 535 -2314
rect 597 -2315 598 -2314
rect 611 -2315 612 -2314
rect 642 -2315 643 -2314
rect 646 -2315 647 -2314
rect 233 -2317 234 -2316
rect 240 -2317 241 -2316
rect 247 -2317 248 -2316
rect 268 -2317 269 -2316
rect 278 -2317 279 -2316
rect 317 -2317 318 -2316
rect 254 -2319 255 -2318
rect 275 -2319 276 -2318
<< metal2 >>
rect 177 -3 178 1
rect 191 -3 192 1
rect 205 -3 206 1
rect 212 -3 213 1
rect 257 -3 258 1
rect 282 -3 283 1
rect 310 -3 311 1
rect 348 -3 349 1
rect 359 -3 360 1
rect 366 -3 367 1
rect 271 -3 272 -1
rect 275 -3 276 -1
rect 177 -13 178 -11
rect 187 -13 188 -11
rect 194 -13 195 -11
rect 198 -13 199 -11
rect 212 -13 213 -11
rect 219 -20 220 -12
rect 233 -20 234 -12
rect 254 -13 255 -11
rect 261 -20 262 -12
rect 275 -13 276 -11
rect 282 -13 283 -11
rect 282 -20 283 -12
rect 282 -13 283 -11
rect 282 -20 283 -12
rect 303 -20 304 -12
rect 310 -13 311 -11
rect 341 -20 342 -12
rect 394 -20 395 -12
rect 184 -15 185 -11
rect 208 -15 209 -11
rect 215 -20 216 -14
rect 254 -20 255 -14
rect 348 -15 349 -11
rect 387 -20 388 -14
rect 198 -20 199 -16
rect 201 -17 202 -11
rect 240 -20 241 -16
rect 250 -20 251 -16
rect 366 -17 367 -11
rect 373 -20 374 -16
rect 366 -20 367 -18
rect 383 -20 384 -18
rect 156 -30 157 -28
rect 156 -41 157 -29
rect 156 -30 157 -28
rect 156 -41 157 -29
rect 166 -41 167 -29
rect 198 -41 199 -29
rect 205 -41 206 -29
rect 271 -30 272 -28
rect 282 -30 283 -28
rect 282 -41 283 -29
rect 282 -30 283 -28
rect 282 -41 283 -29
rect 289 -41 290 -29
rect 296 -30 297 -28
rect 299 -41 300 -29
rect 352 -41 353 -29
rect 387 -30 388 -28
rect 429 -41 430 -29
rect 177 -41 178 -31
rect 212 -32 213 -28
rect 215 -32 216 -28
rect 219 -32 220 -28
rect 226 -41 227 -31
rect 240 -32 241 -28
rect 247 -41 248 -31
rect 261 -32 262 -28
rect 268 -41 269 -31
rect 341 -32 342 -28
rect 345 -41 346 -31
rect 366 -32 367 -28
rect 380 -32 381 -28
rect 387 -41 388 -31
rect 394 -32 395 -28
rect 422 -41 423 -31
rect 194 -41 195 -33
rect 275 -41 276 -33
rect 296 -41 297 -33
rect 331 -41 332 -33
rect 373 -34 374 -28
rect 394 -41 395 -33
rect 411 -41 412 -33
rect 450 -41 451 -33
rect 212 -41 213 -35
rect 233 -36 234 -28
rect 254 -36 255 -28
rect 310 -41 311 -35
rect 317 -41 318 -35
rect 334 -36 335 -28
rect 366 -41 367 -35
rect 373 -41 374 -35
rect 380 -41 381 -35
rect 415 -41 416 -35
rect 219 -41 220 -37
rect 254 -41 255 -37
rect 261 -41 262 -37
rect 338 -41 339 -37
rect 233 -41 234 -39
rect 240 -41 241 -39
rect 303 -40 304 -28
rect 324 -41 325 -39
rect 86 -78 87 -50
rect 107 -51 108 -49
rect 121 -78 122 -50
rect 128 -78 129 -50
rect 142 -78 143 -50
rect 170 -51 171 -49
rect 177 -51 178 -49
rect 187 -51 188 -49
rect 191 -78 192 -50
rect 219 -51 220 -49
rect 233 -78 234 -50
rect 310 -51 311 -49
rect 317 -51 318 -49
rect 464 -78 465 -50
rect 579 -78 580 -50
rect 583 -78 584 -50
rect 93 -78 94 -52
rect 100 -53 101 -49
rect 107 -78 108 -52
rect 170 -78 171 -52
rect 177 -78 178 -52
rect 226 -53 227 -49
rect 247 -53 248 -49
rect 296 -78 297 -52
rect 303 -53 304 -49
rect 352 -53 353 -49
rect 355 -78 356 -52
rect 408 -78 409 -52
rect 436 -53 437 -49
rect 485 -78 486 -52
rect 135 -78 136 -54
rect 219 -78 220 -54
rect 247 -78 248 -54
rect 261 -55 262 -49
rect 268 -55 269 -49
rect 268 -78 269 -54
rect 268 -55 269 -49
rect 268 -78 269 -54
rect 275 -55 276 -49
rect 373 -78 374 -54
rect 394 -55 395 -49
rect 436 -78 437 -54
rect 443 -55 444 -49
rect 471 -78 472 -54
rect 149 -78 150 -56
rect 243 -78 244 -56
rect 275 -78 276 -56
rect 362 -57 363 -49
rect 376 -57 377 -49
rect 394 -78 395 -56
rect 429 -57 430 -49
rect 443 -78 444 -56
rect 450 -57 451 -49
rect 457 -78 458 -56
rect 156 -59 157 -49
rect 156 -78 157 -58
rect 156 -59 157 -49
rect 156 -78 157 -58
rect 163 -78 164 -58
rect 215 -59 216 -49
rect 240 -59 241 -49
rect 261 -78 262 -58
rect 303 -78 304 -58
rect 345 -59 346 -49
rect 348 -78 349 -58
rect 478 -78 479 -58
rect 205 -61 206 -49
rect 317 -78 318 -60
rect 331 -61 332 -49
rect 369 -78 370 -60
rect 422 -61 423 -49
rect 450 -78 451 -60
rect 198 -63 199 -49
rect 205 -78 206 -62
rect 215 -78 216 -62
rect 226 -78 227 -62
rect 324 -63 325 -49
rect 331 -78 332 -62
rect 338 -63 339 -49
rect 380 -78 381 -62
rect 387 -63 388 -49
rect 422 -78 423 -62
rect 100 -78 101 -64
rect 198 -78 199 -64
rect 289 -65 290 -49
rect 387 -78 388 -64
rect 282 -67 283 -49
rect 289 -78 290 -66
rect 310 -78 311 -66
rect 324 -78 325 -66
rect 338 -78 339 -66
rect 415 -67 416 -49
rect 282 -78 283 -68
rect 401 -69 402 -49
rect 341 -78 342 -70
rect 429 -78 430 -70
rect 362 -78 363 -72
rect 499 -78 500 -72
rect 366 -75 367 -49
rect 415 -78 416 -74
rect 401 -78 402 -76
rect 495 -78 496 -76
rect 58 -133 59 -87
rect 135 -88 136 -86
rect 149 -88 150 -86
rect 233 -88 234 -86
rect 282 -88 283 -86
rect 310 -133 311 -87
rect 313 -88 314 -86
rect 415 -88 416 -86
rect 436 -88 437 -86
rect 555 -133 556 -87
rect 562 -88 563 -86
rect 562 -133 563 -87
rect 562 -88 563 -86
rect 562 -133 563 -87
rect 565 -88 566 -86
rect 618 -133 619 -87
rect 65 -133 66 -89
rect 142 -90 143 -86
rect 177 -90 178 -86
rect 233 -133 234 -89
rect 247 -90 248 -86
rect 415 -133 416 -89
rect 436 -133 437 -89
rect 506 -90 507 -86
rect 583 -90 584 -86
rect 597 -133 598 -89
rect 72 -133 73 -91
rect 254 -92 255 -86
rect 282 -133 283 -91
rect 289 -92 290 -86
rect 324 -92 325 -86
rect 324 -133 325 -91
rect 324 -92 325 -86
rect 324 -133 325 -91
rect 345 -92 346 -86
rect 401 -92 402 -86
rect 443 -92 444 -86
rect 443 -133 444 -91
rect 443 -92 444 -86
rect 443 -133 444 -91
rect 450 -92 451 -86
rect 569 -133 570 -91
rect 79 -133 80 -93
rect 114 -94 115 -86
rect 121 -133 122 -93
rect 191 -94 192 -86
rect 205 -94 206 -86
rect 254 -133 255 -93
rect 268 -94 269 -86
rect 401 -133 402 -93
rect 457 -94 458 -86
rect 541 -133 542 -93
rect 86 -96 87 -86
rect 124 -96 125 -86
rect 128 -96 129 -86
rect 128 -133 129 -95
rect 128 -96 129 -86
rect 128 -133 129 -95
rect 180 -133 181 -95
rect 527 -133 528 -95
rect 86 -133 87 -97
rect 163 -98 164 -86
rect 184 -98 185 -86
rect 198 -133 199 -97
rect 205 -133 206 -97
rect 226 -98 227 -86
rect 247 -133 248 -97
rect 296 -98 297 -86
rect 317 -98 318 -86
rect 345 -133 346 -97
rect 348 -98 349 -86
rect 464 -98 465 -86
rect 478 -98 479 -86
rect 492 -133 493 -97
rect 93 -100 94 -86
rect 117 -100 118 -86
rect 149 -133 150 -99
rect 184 -133 185 -99
rect 187 -133 188 -99
rect 240 -133 241 -99
rect 268 -133 269 -99
rect 299 -133 300 -99
rect 352 -133 353 -99
rect 429 -100 430 -86
rect 485 -100 486 -86
rect 583 -133 584 -99
rect 93 -133 94 -101
rect 156 -102 157 -86
rect 163 -133 164 -101
rect 170 -102 171 -86
rect 226 -133 227 -101
rect 296 -133 297 -101
rect 331 -102 332 -86
rect 429 -133 430 -101
rect 114 -133 115 -103
rect 243 -104 244 -86
rect 275 -104 276 -86
rect 317 -133 318 -103
rect 331 -133 332 -103
rect 576 -133 577 -103
rect 170 -133 171 -105
rect 285 -133 286 -105
rect 289 -133 290 -105
rect 303 -106 304 -86
rect 355 -106 356 -86
rect 471 -106 472 -86
rect 156 -133 157 -107
rect 303 -133 304 -107
rect 306 -133 307 -107
rect 471 -133 472 -107
rect 243 -133 244 -109
rect 590 -133 591 -109
rect 261 -112 262 -86
rect 275 -133 276 -111
rect 359 -133 360 -111
rect 499 -112 500 -86
rect 222 -114 223 -86
rect 261 -133 262 -113
rect 362 -114 363 -86
rect 383 -133 384 -113
rect 387 -114 388 -86
rect 534 -133 535 -113
rect 107 -133 108 -115
rect 362 -133 363 -115
rect 366 -116 367 -86
rect 450 -133 451 -115
rect 142 -133 143 -117
rect 222 -133 223 -117
rect 369 -133 370 -117
rect 520 -133 521 -117
rect 177 -133 178 -119
rect 366 -133 367 -119
rect 373 -120 374 -86
rect 499 -133 500 -119
rect 100 -122 101 -86
rect 373 -133 374 -121
rect 376 -133 377 -121
rect 513 -133 514 -121
rect 100 -133 101 -123
rect 135 -133 136 -123
rect 387 -133 388 -123
rect 506 -133 507 -123
rect 394 -126 395 -86
rect 457 -133 458 -125
rect 334 -133 335 -127
rect 394 -133 395 -127
rect 408 -128 409 -86
rect 464 -133 465 -127
rect 380 -130 381 -86
rect 408 -133 409 -129
rect 422 -130 423 -86
rect 485 -133 486 -129
rect 422 -133 423 -131
rect 478 -133 479 -131
rect 51 -143 52 -141
rect 187 -143 188 -141
rect 208 -192 209 -142
rect 376 -143 377 -141
rect 380 -143 381 -141
rect 471 -143 472 -141
rect 485 -143 486 -141
rect 485 -192 486 -142
rect 485 -143 486 -141
rect 485 -192 486 -142
rect 544 -192 545 -142
rect 572 -192 573 -142
rect 618 -143 619 -141
rect 632 -192 633 -142
rect 642 -192 643 -142
rect 646 -192 647 -142
rect 65 -145 66 -141
rect 194 -145 195 -141
rect 222 -145 223 -141
rect 254 -145 255 -141
rect 282 -145 283 -141
rect 429 -145 430 -141
rect 439 -192 440 -144
rect 576 -145 577 -141
rect 65 -192 66 -146
rect 107 -147 108 -141
rect 121 -147 122 -141
rect 229 -147 230 -141
rect 236 -192 237 -146
rect 275 -147 276 -141
rect 282 -192 283 -146
rect 317 -147 318 -141
rect 320 -192 321 -146
rect 401 -147 402 -141
rect 457 -147 458 -141
rect 471 -192 472 -146
rect 506 -147 507 -141
rect 576 -192 577 -146
rect 72 -149 73 -141
rect 376 -192 377 -148
rect 387 -149 388 -141
rect 569 -149 570 -141
rect 79 -151 80 -141
rect 177 -151 178 -141
rect 180 -151 181 -141
rect 362 -151 363 -141
rect 366 -151 367 -141
rect 541 -151 542 -141
rect 79 -192 80 -152
rect 135 -153 136 -141
rect 138 -192 139 -152
rect 366 -192 367 -152
rect 390 -153 391 -141
rect 562 -153 563 -141
rect 86 -155 87 -141
rect 187 -192 188 -154
rect 247 -155 248 -141
rect 254 -192 255 -154
rect 285 -155 286 -141
rect 415 -155 416 -141
rect 457 -192 458 -154
rect 562 -192 563 -154
rect 86 -192 87 -156
rect 243 -157 244 -141
rect 296 -157 297 -141
rect 534 -157 535 -141
rect 100 -192 101 -158
rect 163 -159 164 -141
rect 173 -192 174 -158
rect 240 -192 241 -158
rect 296 -192 297 -158
rect 520 -159 521 -141
rect 527 -159 528 -141
rect 534 -192 535 -158
rect 107 -192 108 -160
rect 156 -161 157 -141
rect 191 -161 192 -141
rect 247 -192 248 -160
rect 317 -192 318 -160
rect 324 -161 325 -141
rect 331 -161 332 -141
rect 499 -161 500 -141
rect 527 -192 528 -160
rect 590 -161 591 -141
rect 114 -163 115 -141
rect 331 -192 332 -162
rect 341 -163 342 -141
rect 387 -192 388 -162
rect 408 -163 409 -141
rect 415 -192 416 -162
rect 464 -163 465 -141
rect 548 -192 549 -162
rect 114 -192 115 -164
rect 128 -165 129 -141
rect 135 -192 136 -164
rect 212 -165 213 -141
rect 324 -192 325 -164
rect 404 -192 405 -164
rect 408 -192 409 -164
rect 422 -165 423 -141
rect 443 -165 444 -141
rect 464 -192 465 -164
rect 478 -165 479 -141
rect 520 -192 521 -164
rect 121 -192 122 -166
rect 170 -167 171 -141
rect 177 -192 178 -166
rect 212 -192 213 -166
rect 345 -167 346 -141
rect 380 -192 381 -166
rect 394 -167 395 -141
rect 478 -192 479 -166
rect 492 -167 493 -141
rect 499 -192 500 -166
rect 513 -167 514 -141
rect 590 -192 591 -166
rect 128 -192 129 -168
rect 310 -169 311 -141
rect 338 -169 339 -141
rect 345 -192 346 -168
rect 352 -169 353 -141
rect 429 -192 430 -168
rect 436 -169 437 -141
rect 513 -192 514 -168
rect 149 -171 150 -141
rect 306 -192 307 -170
rect 359 -171 360 -141
rect 583 -171 584 -141
rect 149 -192 150 -172
rect 299 -173 300 -141
rect 362 -192 363 -172
rect 443 -192 444 -172
rect 450 -173 451 -141
rect 492 -192 493 -172
rect 583 -192 584 -172
rect 597 -173 598 -141
rect 156 -192 157 -174
rect 205 -175 206 -141
rect 261 -175 262 -141
rect 310 -192 311 -174
rect 355 -175 356 -141
rect 450 -192 451 -174
rect 163 -192 164 -176
rect 352 -192 353 -176
rect 355 -192 356 -176
rect 555 -177 556 -141
rect 170 -192 171 -178
rect 268 -179 269 -141
rect 275 -192 276 -178
rect 359 -192 360 -178
rect 551 -179 552 -141
rect 555 -192 556 -178
rect 205 -192 206 -180
rect 422 -192 423 -180
rect 226 -183 227 -141
rect 268 -192 269 -182
rect 289 -183 290 -141
rect 338 -192 339 -182
rect 198 -185 199 -141
rect 226 -192 227 -184
rect 233 -185 234 -141
rect 261 -192 262 -184
rect 289 -192 290 -184
rect 373 -192 374 -184
rect 93 -187 94 -141
rect 233 -192 234 -186
rect 93 -192 94 -188
rect 142 -189 143 -141
rect 198 -192 199 -188
rect 215 -189 216 -141
rect 58 -191 59 -141
rect 142 -192 143 -190
rect 215 -192 216 -190
rect 219 -192 220 -190
rect 16 -249 17 -201
rect 156 -202 157 -200
rect 187 -202 188 -200
rect 275 -202 276 -200
rect 303 -202 304 -200
rect 639 -249 640 -201
rect 646 -202 647 -200
rect 688 -249 689 -201
rect 37 -249 38 -203
rect 184 -204 185 -200
rect 198 -204 199 -200
rect 296 -204 297 -200
rect 317 -204 318 -200
rect 317 -249 318 -203
rect 317 -204 318 -200
rect 317 -249 318 -203
rect 320 -204 321 -200
rect 450 -204 451 -200
rect 460 -204 461 -200
rect 660 -249 661 -203
rect 670 -249 671 -203
rect 674 -249 675 -203
rect 44 -249 45 -205
rect 131 -249 132 -205
rect 205 -206 206 -200
rect 513 -206 514 -200
rect 520 -206 521 -200
rect 653 -249 654 -205
rect 65 -208 66 -200
rect 194 -249 195 -207
rect 212 -249 213 -207
rect 219 -208 220 -200
rect 233 -208 234 -200
rect 401 -249 402 -207
rect 411 -249 412 -207
rect 439 -208 440 -200
rect 467 -249 468 -207
rect 611 -249 612 -207
rect 618 -249 619 -207
rect 632 -208 633 -200
rect 65 -249 66 -209
rect 142 -210 143 -200
rect 233 -249 234 -209
rect 240 -210 241 -200
rect 261 -210 262 -200
rect 275 -249 276 -209
rect 289 -210 290 -200
rect 303 -249 304 -209
rect 331 -210 332 -200
rect 457 -249 458 -209
rect 513 -249 514 -209
rect 548 -210 549 -200
rect 562 -210 563 -200
rect 695 -249 696 -209
rect 79 -212 80 -200
rect 219 -249 220 -211
rect 236 -212 237 -200
rect 296 -249 297 -211
rect 355 -212 356 -200
rect 562 -249 563 -211
rect 569 -212 570 -200
rect 583 -212 584 -200
rect 590 -212 591 -200
rect 632 -249 633 -211
rect 51 -249 52 -213
rect 79 -249 80 -213
rect 86 -214 87 -200
rect 138 -214 139 -200
rect 173 -214 174 -200
rect 289 -249 290 -213
rect 359 -249 360 -213
rect 380 -214 381 -200
rect 390 -249 391 -213
rect 478 -214 479 -200
rect 520 -249 521 -213
rect 555 -214 556 -200
rect 569 -249 570 -213
rect 751 -249 752 -213
rect 86 -249 87 -215
rect 149 -216 150 -200
rect 222 -249 223 -215
rect 380 -249 381 -215
rect 397 -216 398 -200
rect 464 -216 465 -200
rect 471 -216 472 -200
rect 555 -249 556 -215
rect 576 -216 577 -200
rect 681 -249 682 -215
rect 93 -218 94 -200
rect 261 -249 262 -217
rect 268 -218 269 -200
rect 331 -249 332 -217
rect 373 -218 374 -200
rect 625 -249 626 -217
rect 93 -249 94 -219
rect 145 -249 146 -219
rect 198 -249 199 -219
rect 268 -249 269 -219
rect 282 -220 283 -200
rect 373 -249 374 -219
rect 376 -220 377 -200
rect 485 -220 486 -200
rect 492 -220 493 -200
rect 576 -249 577 -219
rect 597 -249 598 -219
rect 667 -249 668 -219
rect 100 -222 101 -200
rect 184 -249 185 -221
rect 240 -249 241 -221
rect 254 -222 255 -200
rect 299 -222 300 -200
rect 471 -249 472 -221
rect 527 -222 528 -200
rect 646 -249 647 -221
rect 30 -249 31 -223
rect 100 -249 101 -223
rect 107 -224 108 -200
rect 191 -224 192 -200
rect 226 -224 227 -200
rect 254 -249 255 -223
rect 397 -249 398 -223
rect 450 -249 451 -223
rect 464 -249 465 -223
rect 534 -224 535 -200
rect 544 -224 545 -200
rect 583 -249 584 -223
rect 23 -249 24 -225
rect 107 -249 108 -225
rect 121 -226 122 -200
rect 149 -249 150 -225
rect 177 -226 178 -200
rect 282 -249 283 -225
rect 324 -226 325 -200
rect 534 -249 535 -225
rect 58 -249 59 -227
rect 226 -249 227 -227
rect 310 -228 311 -200
rect 324 -249 325 -227
rect 404 -228 405 -200
rect 478 -249 479 -227
rect 509 -228 510 -200
rect 527 -249 528 -227
rect 72 -230 73 -200
rect 191 -249 192 -229
rect 247 -230 248 -200
rect 310 -249 311 -229
rect 408 -230 409 -200
rect 548 -249 549 -229
rect 72 -249 73 -231
rect 114 -232 115 -200
rect 121 -249 122 -231
rect 142 -249 143 -231
rect 163 -232 164 -200
rect 247 -249 248 -231
rect 408 -249 409 -231
rect 499 -232 500 -200
rect 114 -249 115 -233
rect 208 -234 209 -200
rect 415 -234 416 -200
rect 436 -249 437 -233
rect 443 -234 444 -200
rect 492 -249 493 -233
rect 128 -236 129 -200
rect 352 -249 353 -235
rect 366 -236 367 -200
rect 443 -249 444 -235
rect 485 -249 486 -235
rect 509 -249 510 -235
rect 128 -249 129 -237
rect 170 -249 171 -237
rect 208 -249 209 -237
rect 541 -249 542 -237
rect 138 -249 139 -239
rect 177 -249 178 -239
rect 338 -240 339 -200
rect 366 -249 367 -239
rect 422 -240 423 -200
rect 590 -249 591 -239
rect 163 -249 164 -241
rect 229 -249 230 -241
rect 338 -249 339 -241
rect 499 -249 500 -241
rect 345 -244 346 -200
rect 415 -249 416 -243
rect 418 -249 419 -243
rect 422 -249 423 -243
rect 429 -244 430 -200
rect 506 -244 507 -200
rect 345 -249 346 -245
rect 387 -246 388 -200
rect 394 -246 395 -200
rect 429 -249 430 -245
rect 394 -249 395 -247
rect 604 -249 605 -247
rect 23 -259 24 -257
rect 135 -302 136 -258
rect 142 -302 143 -258
rect 261 -259 262 -257
rect 299 -302 300 -258
rect 425 -302 426 -258
rect 439 -302 440 -258
rect 576 -259 577 -257
rect 583 -259 584 -257
rect 583 -302 584 -258
rect 583 -259 584 -257
rect 583 -302 584 -258
rect 590 -259 591 -257
rect 593 -283 594 -258
rect 597 -259 598 -257
rect 600 -259 601 -257
rect 604 -259 605 -257
rect 670 -259 671 -257
rect 674 -259 675 -257
rect 716 -302 717 -258
rect 751 -259 752 -257
rect 828 -302 829 -258
rect 856 -302 857 -258
rect 859 -259 860 -257
rect 51 -302 52 -260
rect 58 -261 59 -257
rect 65 -261 66 -257
rect 236 -302 237 -260
rect 240 -261 241 -257
rect 271 -261 272 -257
rect 334 -302 335 -260
rect 660 -261 661 -257
rect 681 -261 682 -257
rect 737 -302 738 -260
rect 16 -263 17 -257
rect 240 -302 241 -262
rect 247 -263 248 -257
rect 397 -263 398 -257
rect 401 -263 402 -257
rect 572 -263 573 -257
rect 590 -302 591 -262
rect 639 -263 640 -257
rect 646 -263 647 -257
rect 681 -302 682 -262
rect 688 -263 689 -257
rect 744 -302 745 -262
rect 58 -302 59 -264
rect 79 -265 80 -257
rect 107 -265 108 -257
rect 121 -265 122 -257
rect 128 -302 129 -264
rect 226 -265 227 -257
rect 229 -265 230 -257
rect 254 -265 255 -257
rect 261 -302 262 -264
rect 275 -265 276 -257
rect 338 -265 339 -257
rect 352 -265 353 -257
rect 359 -265 360 -257
rect 408 -302 409 -264
rect 415 -302 416 -264
rect 422 -265 423 -257
rect 443 -265 444 -257
rect 478 -302 479 -264
rect 485 -265 486 -257
rect 485 -302 486 -264
rect 485 -265 486 -257
rect 485 -302 486 -264
rect 492 -265 493 -257
rect 492 -302 493 -264
rect 492 -265 493 -257
rect 492 -302 493 -264
rect 499 -265 500 -257
rect 502 -283 503 -264
rect 534 -265 535 -257
rect 569 -302 570 -264
rect 597 -302 598 -264
rect 611 -265 612 -257
rect 618 -265 619 -257
rect 667 -265 668 -257
rect 688 -302 689 -264
rect 723 -302 724 -264
rect 44 -267 45 -257
rect 79 -302 80 -266
rect 107 -302 108 -266
rect 156 -267 157 -257
rect 191 -302 192 -266
rect 194 -267 195 -257
rect 205 -267 206 -257
rect 226 -302 227 -266
rect 268 -267 269 -257
rect 352 -302 353 -266
rect 359 -302 360 -266
rect 401 -302 402 -266
rect 446 -302 447 -266
rect 604 -302 605 -266
rect 625 -267 626 -257
rect 709 -302 710 -266
rect 68 -302 69 -268
rect 100 -269 101 -257
rect 114 -269 115 -257
rect 159 -269 160 -257
rect 184 -269 185 -257
rect 268 -302 269 -268
rect 275 -302 276 -268
rect 310 -269 311 -257
rect 341 -269 342 -257
rect 457 -302 458 -268
rect 460 -269 461 -257
rect 730 -302 731 -268
rect 72 -271 73 -257
rect 138 -271 139 -257
rect 149 -271 150 -257
rect 156 -302 157 -270
rect 177 -271 178 -257
rect 184 -302 185 -270
rect 205 -302 206 -270
rect 296 -271 297 -257
rect 310 -302 311 -270
rect 317 -271 318 -257
rect 373 -271 374 -257
rect 397 -302 398 -270
rect 481 -271 482 -257
rect 667 -302 668 -270
rect 37 -273 38 -257
rect 177 -302 178 -272
rect 215 -273 216 -257
rect 404 -302 405 -272
rect 499 -302 500 -272
rect 520 -273 521 -257
rect 625 -302 626 -272
rect 632 -273 633 -257
rect 646 -302 647 -272
rect 30 -275 31 -257
rect 215 -302 216 -274
rect 222 -302 223 -274
rect 282 -275 283 -257
rect 296 -302 297 -274
rect 303 -275 304 -257
rect 317 -302 318 -274
rect 324 -275 325 -257
rect 373 -302 374 -274
rect 751 -302 752 -274
rect 30 -302 31 -276
rect 86 -277 87 -257
rect 100 -302 101 -276
rect 103 -277 104 -257
rect 117 -302 118 -276
rect 632 -302 633 -276
rect 639 -302 640 -276
rect 653 -277 654 -257
rect 37 -302 38 -278
rect 93 -279 94 -257
rect 121 -302 122 -278
rect 198 -279 199 -257
rect 282 -302 283 -278
rect 331 -279 332 -257
rect 380 -279 381 -257
rect 464 -302 465 -278
rect 471 -279 472 -257
rect 520 -302 521 -278
rect 541 -279 542 -257
rect 618 -302 619 -278
rect 72 -302 73 -280
rect 163 -281 164 -257
rect 180 -302 181 -280
rect 198 -302 199 -280
rect 243 -302 244 -280
rect 380 -302 381 -280
rect 390 -281 391 -257
rect 544 -302 545 -280
rect 555 -281 556 -257
rect 660 -302 661 -280
rect 86 -302 87 -282
rect 331 -302 332 -282
rect 394 -302 395 -282
rect 534 -302 535 -282
rect 562 -283 563 -257
rect 576 -302 577 -282
rect 600 -302 601 -282
rect 611 -302 612 -282
rect 93 -302 94 -284
rect 254 -302 255 -284
rect 289 -285 290 -257
rect 303 -302 304 -284
rect 324 -302 325 -284
rect 366 -285 367 -257
rect 429 -285 430 -257
rect 471 -302 472 -284
rect 527 -285 528 -257
rect 555 -302 556 -284
rect 565 -302 566 -284
rect 702 -302 703 -284
rect 149 -302 150 -286
rect 170 -287 171 -257
rect 345 -287 346 -257
rect 366 -302 367 -286
rect 411 -287 412 -257
rect 527 -302 528 -286
rect 163 -302 164 -288
rect 541 -302 542 -288
rect 170 -302 171 -290
rect 233 -291 234 -257
rect 345 -302 346 -290
rect 548 -291 549 -257
rect 387 -293 388 -257
rect 548 -302 549 -292
rect 387 -302 388 -294
rect 695 -295 696 -257
rect 429 -302 430 -296
rect 436 -297 437 -257
rect 450 -297 451 -257
rect 562 -302 563 -296
rect 422 -302 423 -298
rect 450 -302 451 -298
rect 506 -299 507 -257
rect 695 -302 696 -298
rect 338 -302 339 -300
rect 506 -302 507 -300
rect 2 -373 3 -311
rect 100 -312 101 -310
rect 107 -312 108 -310
rect 114 -312 115 -310
rect 121 -312 122 -310
rect 124 -364 125 -311
rect 128 -312 129 -310
rect 495 -373 496 -311
rect 653 -312 654 -310
rect 835 -373 836 -311
rect 849 -373 850 -311
rect 863 -373 864 -311
rect 9 -373 10 -313
rect 65 -314 66 -310
rect 72 -314 73 -310
rect 215 -314 216 -310
rect 226 -314 227 -310
rect 226 -373 227 -313
rect 226 -314 227 -310
rect 226 -373 227 -313
rect 233 -314 234 -310
rect 345 -314 346 -310
rect 352 -314 353 -310
rect 562 -314 563 -310
rect 590 -314 591 -310
rect 653 -373 654 -313
rect 674 -373 675 -313
rect 677 -314 678 -310
rect 681 -314 682 -310
rect 723 -373 724 -313
rect 726 -314 727 -310
rect 870 -373 871 -313
rect 16 -373 17 -315
rect 79 -316 80 -310
rect 114 -373 115 -315
rect 415 -316 416 -310
rect 422 -373 423 -315
rect 492 -316 493 -310
rect 534 -316 535 -310
rect 562 -373 563 -315
rect 569 -316 570 -310
rect 590 -373 591 -315
rect 695 -316 696 -310
rect 779 -373 780 -315
rect 828 -316 829 -310
rect 891 -373 892 -315
rect 23 -373 24 -317
rect 177 -318 178 -310
rect 215 -373 216 -317
rect 247 -318 248 -310
rect 257 -318 258 -310
rect 261 -318 262 -310
rect 275 -318 276 -310
rect 341 -318 342 -310
rect 352 -373 353 -317
rect 485 -318 486 -310
rect 513 -318 514 -310
rect 534 -373 535 -317
rect 548 -318 549 -310
rect 569 -373 570 -317
rect 597 -318 598 -310
rect 695 -373 696 -317
rect 702 -318 703 -310
rect 814 -373 815 -317
rect 852 -373 853 -317
rect 856 -318 857 -310
rect 30 -320 31 -310
rect 79 -373 80 -319
rect 96 -373 97 -319
rect 177 -373 178 -319
rect 219 -320 220 -310
rect 345 -373 346 -319
rect 359 -320 360 -310
rect 432 -373 433 -319
rect 450 -320 451 -310
rect 453 -320 454 -310
rect 513 -373 514 -319
rect 520 -320 521 -310
rect 544 -320 545 -310
rect 702 -373 703 -319
rect 709 -320 710 -310
rect 758 -373 759 -319
rect 44 -322 45 -310
rect 107 -373 108 -321
rect 121 -373 122 -321
rect 394 -322 395 -310
rect 401 -322 402 -310
rect 660 -322 661 -310
rect 667 -322 668 -310
rect 709 -373 710 -321
rect 716 -322 717 -310
rect 716 -373 717 -321
rect 716 -322 717 -310
rect 716 -373 717 -321
rect 730 -322 731 -310
rect 828 -373 829 -321
rect 44 -373 45 -323
rect 236 -324 237 -310
rect 240 -324 241 -310
rect 443 -373 444 -323
rect 450 -373 451 -323
rect 471 -324 472 -310
rect 520 -373 521 -323
rect 527 -324 528 -310
rect 583 -324 584 -310
rect 597 -373 598 -323
rect 618 -324 619 -310
rect 660 -373 661 -323
rect 737 -324 738 -310
rect 807 -373 808 -323
rect 51 -326 52 -310
rect 338 -326 339 -310
rect 362 -373 363 -325
rect 800 -373 801 -325
rect 51 -373 52 -327
rect 184 -328 185 -310
rect 233 -373 234 -327
rect 793 -373 794 -327
rect 37 -330 38 -310
rect 184 -373 185 -329
rect 240 -373 241 -329
rect 282 -330 283 -310
rect 289 -330 290 -310
rect 681 -373 682 -329
rect 744 -330 745 -310
rect 786 -373 787 -329
rect 58 -332 59 -310
rect 131 -373 132 -331
rect 135 -373 136 -331
rect 222 -332 223 -310
rect 247 -373 248 -331
rect 317 -332 318 -310
rect 334 -332 335 -310
rect 408 -332 409 -310
rect 471 -373 472 -331
rect 478 -332 479 -310
rect 499 -332 500 -310
rect 527 -373 528 -331
rect 583 -373 584 -331
rect 632 -332 633 -310
rect 639 -332 640 -310
rect 730 -373 731 -331
rect 751 -332 752 -310
rect 821 -373 822 -331
rect 58 -373 59 -333
rect 149 -334 150 -310
rect 212 -334 213 -310
rect 408 -373 409 -333
rect 474 -373 475 -333
rect 618 -373 619 -333
rect 639 -373 640 -333
rect 877 -373 878 -333
rect 65 -373 66 -335
rect 191 -336 192 -310
rect 261 -373 262 -335
rect 303 -336 304 -310
rect 310 -336 311 -310
rect 338 -373 339 -335
rect 373 -373 374 -335
rect 765 -373 766 -335
rect 75 -373 76 -337
rect 152 -373 153 -337
rect 170 -338 171 -310
rect 191 -373 192 -337
rect 282 -373 283 -337
rect 324 -338 325 -310
rect 380 -338 381 -310
rect 548 -373 549 -337
rect 586 -373 587 -337
rect 856 -373 857 -337
rect 86 -340 87 -310
rect 317 -373 318 -339
rect 380 -373 381 -339
rect 387 -340 388 -310
rect 394 -373 395 -339
rect 457 -340 458 -310
rect 506 -340 507 -310
rect 632 -373 633 -339
rect 646 -340 647 -310
rect 667 -373 668 -339
rect 688 -340 689 -310
rect 751 -373 752 -339
rect 86 -373 87 -341
rect 268 -342 269 -310
rect 289 -373 290 -341
rect 324 -373 325 -341
rect 401 -373 402 -341
rect 425 -373 426 -341
rect 436 -342 437 -310
rect 688 -373 689 -341
rect 93 -344 94 -310
rect 310 -373 311 -343
rect 429 -344 430 -310
rect 436 -373 437 -343
rect 457 -373 458 -343
rect 464 -344 465 -310
rect 516 -373 517 -343
rect 744 -373 745 -343
rect 93 -373 94 -345
rect 842 -373 843 -345
rect 100 -373 101 -347
rect 359 -373 360 -347
rect 429 -373 430 -347
rect 499 -373 500 -347
rect 604 -348 605 -310
rect 737 -373 738 -347
rect 128 -373 129 -349
rect 219 -373 220 -349
rect 254 -350 255 -310
rect 387 -373 388 -349
rect 604 -373 605 -349
rect 611 -350 612 -310
rect 625 -350 626 -310
rect 646 -373 647 -349
rect 138 -352 139 -310
rect 275 -373 276 -351
rect 296 -373 297 -351
rect 404 -373 405 -351
rect 576 -352 577 -310
rect 611 -373 612 -351
rect 142 -354 143 -310
rect 369 -373 370 -353
rect 555 -354 556 -310
rect 576 -373 577 -353
rect 30 -373 31 -355
rect 142 -373 143 -355
rect 145 -373 146 -355
rect 485 -373 486 -355
rect 156 -358 157 -310
rect 170 -373 171 -357
rect 464 -373 465 -357
rect 156 -373 157 -359
rect 163 -360 164 -310
rect 254 -373 255 -359
rect 327 -373 328 -359
rect 331 -360 332 -310
rect 555 -373 556 -359
rect 37 -373 38 -361
rect 331 -373 332 -361
rect 334 -373 335 -361
rect 625 -373 626 -361
rect 163 -373 164 -363
rect 205 -364 206 -310
rect 268 -373 269 -363
rect 439 -364 440 -310
rect 453 -373 454 -363
rect 478 -373 479 -363
rect 205 -373 206 -365
rect 415 -373 416 -365
rect 299 -368 300 -310
rect 541 -373 542 -367
rect 303 -373 304 -369
rect 366 -370 367 -310
rect 366 -373 367 -371
rect 772 -373 773 -371
rect 2 -383 3 -381
rect 198 -383 199 -381
rect 205 -383 206 -381
rect 940 -462 941 -382
rect 2 -462 3 -384
rect 198 -462 199 -384
rect 226 -385 227 -381
rect 226 -462 227 -384
rect 226 -385 227 -381
rect 226 -462 227 -384
rect 261 -385 262 -381
rect 362 -385 363 -381
rect 369 -385 370 -381
rect 534 -385 535 -381
rect 621 -462 622 -384
rect 639 -385 640 -381
rect 660 -385 661 -381
rect 660 -462 661 -384
rect 660 -385 661 -381
rect 660 -462 661 -384
rect 758 -385 759 -381
rect 758 -462 759 -384
rect 758 -385 759 -381
rect 758 -462 759 -384
rect 828 -385 829 -381
rect 877 -462 878 -384
rect 16 -387 17 -381
rect 131 -387 132 -381
rect 159 -462 160 -386
rect 905 -462 906 -386
rect 16 -462 17 -388
rect 44 -389 45 -381
rect 51 -389 52 -381
rect 215 -462 216 -388
rect 261 -462 262 -388
rect 432 -389 433 -381
rect 478 -389 479 -381
rect 513 -389 514 -381
rect 516 -389 517 -381
rect 737 -389 738 -381
rect 842 -389 843 -381
rect 898 -462 899 -388
rect 23 -391 24 -381
rect 243 -462 244 -390
rect 275 -462 276 -390
rect 432 -462 433 -390
rect 436 -391 437 -381
rect 478 -462 479 -390
rect 502 -462 503 -390
rect 807 -391 808 -381
rect 852 -391 853 -381
rect 891 -391 892 -381
rect 23 -462 24 -392
rect 177 -393 178 -381
rect 282 -393 283 -381
rect 376 -393 377 -381
rect 390 -462 391 -392
rect 779 -393 780 -381
rect 807 -462 808 -392
rect 849 -393 850 -381
rect 863 -393 864 -381
rect 884 -393 885 -381
rect 37 -395 38 -381
rect 506 -395 507 -381
rect 509 -395 510 -381
rect 933 -462 934 -394
rect 37 -462 38 -396
rect 103 -462 104 -396
rect 107 -397 108 -381
rect 222 -462 223 -396
rect 310 -397 311 -381
rect 348 -462 349 -396
rect 359 -397 360 -381
rect 653 -397 654 -381
rect 716 -397 717 -381
rect 891 -462 892 -396
rect 44 -462 45 -398
rect 177 -462 178 -398
rect 184 -399 185 -381
rect 282 -462 283 -398
rect 303 -399 304 -381
rect 310 -462 311 -398
rect 317 -399 318 -381
rect 492 -462 493 -398
rect 495 -399 496 -381
rect 884 -462 885 -398
rect 54 -462 55 -400
rect 135 -401 136 -381
rect 145 -401 146 -381
rect 863 -462 864 -400
rect 870 -401 871 -381
rect 926 -462 927 -400
rect 75 -403 76 -381
rect 268 -403 269 -381
rect 303 -462 304 -402
rect 821 -403 822 -381
rect 79 -405 80 -381
rect 96 -405 97 -381
rect 100 -405 101 -381
rect 184 -462 185 -404
rect 201 -405 202 -381
rect 268 -462 269 -404
rect 324 -462 325 -404
rect 394 -405 395 -381
rect 401 -405 402 -381
rect 457 -405 458 -381
rect 520 -405 521 -381
rect 583 -462 584 -404
rect 604 -405 605 -381
rect 639 -462 640 -404
rect 674 -405 675 -381
rect 870 -462 871 -404
rect 9 -407 10 -381
rect 79 -462 80 -406
rect 86 -407 87 -381
rect 233 -407 234 -381
rect 240 -407 241 -381
rect 359 -462 360 -406
rect 373 -407 374 -381
rect 828 -462 829 -406
rect 9 -462 10 -408
rect 219 -409 220 -381
rect 240 -462 241 -408
rect 317 -462 318 -408
rect 331 -409 332 -381
rect 352 -409 353 -381
rect 408 -409 409 -381
rect 509 -462 510 -408
rect 520 -462 521 -408
rect 751 -409 752 -381
rect 772 -409 773 -381
rect 849 -462 850 -408
rect 72 -411 73 -381
rect 352 -462 353 -410
rect 369 -462 370 -410
rect 408 -462 409 -410
rect 415 -411 416 -381
rect 534 -462 535 -410
rect 555 -411 556 -381
rect 653 -462 654 -410
rect 695 -411 696 -381
rect 772 -462 773 -410
rect 814 -411 815 -381
rect 821 -462 822 -410
rect 72 -462 73 -412
rect 163 -413 164 -381
rect 170 -413 171 -381
rect 205 -462 206 -412
rect 212 -413 213 -381
rect 779 -462 780 -412
rect 86 -462 87 -414
rect 156 -415 157 -381
rect 163 -462 164 -414
rect 569 -415 570 -381
rect 576 -415 577 -381
rect 604 -462 605 -414
rect 625 -415 626 -381
rect 695 -462 696 -414
rect 716 -462 717 -414
rect 800 -415 801 -381
rect 93 -462 94 -416
rect 247 -417 248 -381
rect 254 -417 255 -381
rect 373 -462 374 -416
rect 422 -417 423 -381
rect 842 -462 843 -416
rect 65 -419 66 -381
rect 254 -462 255 -418
rect 289 -419 290 -381
rect 394 -462 395 -418
rect 422 -462 423 -418
rect 681 -419 682 -381
rect 730 -419 731 -381
rect 814 -462 815 -418
rect 58 -421 59 -381
rect 65 -462 66 -420
rect 107 -462 108 -420
rect 366 -421 367 -381
rect 425 -421 426 -381
rect 597 -421 598 -381
rect 611 -421 612 -381
rect 625 -462 626 -420
rect 646 -421 647 -381
rect 681 -462 682 -420
rect 730 -462 731 -420
rect 765 -421 766 -381
rect 58 -462 59 -422
rect 296 -423 297 -381
rect 338 -423 339 -381
rect 947 -462 948 -422
rect 110 -462 111 -424
rect 247 -462 248 -424
rect 289 -462 290 -424
rect 380 -425 381 -381
rect 436 -462 437 -424
rect 835 -425 836 -381
rect 117 -462 118 -426
rect 383 -462 384 -426
rect 450 -427 451 -381
rect 457 -462 458 -426
rect 471 -427 472 -381
rect 800 -462 801 -426
rect 835 -462 836 -426
rect 856 -427 857 -381
rect 114 -429 115 -381
rect 471 -462 472 -428
rect 485 -429 486 -381
rect 576 -462 577 -428
rect 590 -429 591 -381
rect 674 -462 675 -428
rect 688 -429 689 -381
rect 765 -462 766 -428
rect 114 -462 115 -430
rect 569 -462 570 -430
rect 632 -431 633 -381
rect 856 -462 857 -430
rect 121 -433 122 -381
rect 401 -462 402 -432
rect 418 -462 419 -432
rect 450 -462 451 -432
rect 523 -462 524 -432
rect 919 -462 920 -432
rect 121 -462 122 -434
rect 149 -435 150 -381
rect 156 -462 157 -434
rect 334 -435 335 -381
rect 345 -435 346 -381
rect 513 -462 514 -434
rect 527 -435 528 -381
rect 590 -462 591 -434
rect 646 -462 647 -434
rect 667 -435 668 -381
rect 688 -462 689 -434
rect 709 -435 710 -381
rect 751 -462 752 -434
rect 786 -435 787 -381
rect 30 -437 31 -381
rect 149 -462 150 -436
rect 212 -462 213 -436
rect 912 -462 913 -436
rect 30 -462 31 -438
rect 128 -439 129 -381
rect 135 -462 136 -438
rect 306 -462 307 -438
rect 366 -462 367 -438
rect 597 -462 598 -438
rect 618 -439 619 -381
rect 786 -462 787 -438
rect 128 -462 129 -440
rect 191 -441 192 -381
rect 233 -462 234 -440
rect 485 -462 486 -440
rect 548 -441 549 -381
rect 632 -462 633 -440
rect 667 -462 668 -440
rect 744 -441 745 -381
rect 142 -443 143 -381
rect 170 -462 171 -442
rect 191 -462 192 -442
rect 338 -462 339 -442
rect 404 -443 405 -381
rect 527 -462 528 -442
rect 555 -462 556 -442
rect 562 -443 563 -381
rect 611 -462 612 -442
rect 618 -462 619 -442
rect 702 -443 703 -381
rect 709 -462 710 -442
rect 142 -462 143 -444
rect 429 -445 430 -381
rect 443 -445 444 -381
rect 548 -462 549 -444
rect 702 -462 703 -444
rect 793 -445 794 -381
rect 152 -447 153 -381
rect 744 -462 745 -446
rect 296 -462 297 -448
rect 737 -462 738 -448
rect 331 -462 332 -450
rect 429 -462 430 -450
rect 541 -451 542 -381
rect 562 -462 563 -450
rect 723 -451 724 -381
rect 793 -462 794 -450
rect 299 -462 300 -452
rect 723 -462 724 -452
rect 387 -455 388 -381
rect 443 -462 444 -454
rect 499 -455 500 -381
rect 541 -462 542 -454
rect 278 -457 279 -381
rect 499 -462 500 -456
rect 387 -462 388 -458
rect 464 -459 465 -381
rect 415 -462 416 -460
rect 464 -462 465 -460
rect 2 -472 3 -470
rect 264 -549 265 -471
rect 268 -472 269 -470
rect 425 -549 426 -471
rect 429 -472 430 -470
rect 814 -472 815 -470
rect 2 -549 3 -473
rect 219 -474 220 -470
rect 243 -474 244 -470
rect 513 -474 514 -470
rect 544 -549 545 -473
rect 891 -474 892 -470
rect 9 -476 10 -470
rect 520 -476 521 -470
rect 607 -549 608 -475
rect 618 -549 619 -475
rect 716 -476 717 -470
rect 716 -549 717 -475
rect 716 -476 717 -470
rect 716 -549 717 -475
rect 726 -549 727 -475
rect 821 -476 822 -470
rect 9 -549 10 -477
rect 44 -549 45 -477
rect 51 -478 52 -470
rect 145 -549 146 -477
rect 170 -478 171 -470
rect 170 -549 171 -477
rect 170 -478 171 -470
rect 170 -549 171 -477
rect 180 -549 181 -477
rect 201 -478 202 -470
rect 212 -478 213 -470
rect 940 -478 941 -470
rect 30 -480 31 -470
rect 51 -549 52 -479
rect 54 -480 55 -470
rect 695 -480 696 -470
rect 807 -480 808 -470
rect 807 -549 808 -479
rect 807 -480 808 -470
rect 807 -549 808 -479
rect 814 -549 815 -479
rect 919 -480 920 -470
rect 30 -549 31 -481
rect 37 -482 38 -470
rect 58 -482 59 -470
rect 303 -482 304 -470
rect 313 -549 314 -481
rect 947 -482 948 -470
rect 37 -549 38 -483
rect 383 -484 384 -470
rect 394 -484 395 -470
rect 418 -484 419 -470
rect 439 -484 440 -470
rect 796 -549 797 -483
rect 58 -549 59 -485
rect 135 -486 136 -470
rect 184 -486 185 -470
rect 219 -549 220 -485
rect 243 -549 244 -485
rect 282 -486 283 -470
rect 303 -549 304 -485
rect 317 -486 318 -470
rect 320 -549 321 -485
rect 548 -486 549 -470
rect 695 -549 696 -485
rect 702 -486 703 -470
rect 79 -488 80 -470
rect 96 -549 97 -487
rect 100 -488 101 -470
rect 653 -488 654 -470
rect 660 -488 661 -470
rect 702 -549 703 -487
rect 23 -490 24 -470
rect 79 -549 80 -489
rect 86 -490 87 -470
rect 198 -490 199 -470
rect 324 -490 325 -470
rect 394 -549 395 -489
rect 401 -490 402 -470
rect 821 -549 822 -489
rect 86 -549 87 -491
rect 247 -492 248 -470
rect 352 -492 353 -470
rect 432 -492 433 -470
rect 443 -492 444 -470
rect 443 -549 444 -491
rect 443 -492 444 -470
rect 443 -549 444 -491
rect 460 -492 461 -470
rect 765 -492 766 -470
rect 100 -549 101 -493
rect 107 -494 108 -470
rect 114 -549 115 -493
rect 390 -549 391 -493
rect 408 -494 409 -470
rect 429 -549 430 -493
rect 464 -494 465 -470
rect 523 -494 524 -470
rect 541 -494 542 -470
rect 548 -549 549 -493
rect 639 -494 640 -470
rect 660 -549 661 -493
rect 765 -549 766 -493
rect 835 -494 836 -470
rect 82 -496 83 -470
rect 107 -549 108 -495
rect 117 -496 118 -470
rect 674 -496 675 -470
rect 835 -549 836 -495
rect 842 -496 843 -470
rect 121 -498 122 -470
rect 408 -549 409 -497
rect 415 -498 416 -470
rect 793 -498 794 -470
rect 121 -549 122 -499
rect 345 -500 346 -470
rect 359 -500 360 -470
rect 369 -500 370 -470
rect 373 -500 374 -470
rect 401 -549 402 -499
rect 415 -549 416 -499
rect 576 -500 577 -470
rect 639 -549 640 -499
rect 667 -500 668 -470
rect 674 -549 675 -499
rect 688 -500 689 -470
rect 128 -502 129 -470
rect 296 -502 297 -470
rect 324 -549 325 -501
rect 541 -549 542 -501
rect 576 -549 577 -501
rect 604 -502 605 -470
rect 646 -502 647 -470
rect 653 -549 654 -501
rect 667 -549 668 -501
rect 754 -549 755 -501
rect 16 -504 17 -470
rect 128 -549 129 -503
rect 135 -549 136 -503
rect 310 -504 311 -470
rect 366 -504 367 -470
rect 471 -504 472 -470
rect 485 -504 486 -470
rect 779 -504 780 -470
rect 16 -549 17 -505
rect 163 -506 164 -470
rect 166 -506 167 -470
rect 485 -549 486 -505
rect 488 -506 489 -470
rect 870 -506 871 -470
rect 142 -508 143 -470
rect 352 -549 353 -507
rect 373 -549 374 -507
rect 534 -508 535 -470
rect 646 -549 647 -507
rect 849 -508 850 -470
rect 149 -510 150 -470
rect 166 -549 167 -509
rect 177 -510 178 -470
rect 282 -549 283 -509
rect 296 -549 297 -509
rect 334 -549 335 -509
rect 338 -510 339 -470
rect 366 -549 367 -509
rect 380 -510 381 -470
rect 632 -510 633 -470
rect 688 -549 689 -509
rect 737 -510 738 -470
rect 779 -549 780 -509
rect 884 -510 885 -470
rect 65 -512 66 -470
rect 149 -549 150 -511
rect 156 -549 157 -511
rect 471 -549 472 -511
rect 502 -549 503 -511
rect 898 -512 899 -470
rect 65 -549 66 -513
rect 348 -514 349 -470
rect 464 -549 465 -513
rect 481 -549 482 -513
rect 506 -514 507 -470
rect 786 -514 787 -470
rect 163 -549 164 -515
rect 422 -516 423 -470
rect 509 -549 510 -515
rect 856 -516 857 -470
rect 184 -549 185 -517
rect 226 -518 227 -470
rect 247 -549 248 -517
rect 387 -518 388 -470
rect 422 -549 423 -517
rect 583 -518 584 -470
rect 632 -549 633 -517
rect 681 -518 682 -470
rect 709 -518 710 -470
rect 737 -549 738 -517
rect 786 -549 787 -517
rect 933 -518 934 -470
rect 191 -520 192 -470
rect 772 -520 773 -470
rect 856 -549 857 -519
rect 926 -520 927 -470
rect 93 -522 94 -470
rect 191 -549 192 -521
rect 194 -522 195 -470
rect 240 -522 241 -470
rect 254 -522 255 -470
rect 345 -549 346 -521
rect 387 -549 388 -521
rect 590 -522 591 -470
rect 709 -549 710 -521
rect 800 -522 801 -470
rect 93 -549 94 -523
rect 306 -524 307 -470
rect 341 -549 342 -523
rect 534 -549 535 -523
rect 569 -524 570 -470
rect 583 -549 584 -523
rect 590 -549 591 -523
rect 597 -524 598 -470
rect 751 -524 752 -470
rect 772 -549 773 -523
rect 800 -549 801 -523
rect 912 -524 913 -470
rect 198 -549 199 -525
rect 233 -526 234 -470
rect 240 -549 241 -525
rect 905 -526 906 -470
rect 226 -549 227 -527
rect 492 -528 493 -470
rect 513 -549 514 -527
rect 527 -528 528 -470
rect 597 -549 598 -527
rect 625 -528 626 -470
rect 233 -549 234 -529
rect 499 -530 500 -470
rect 520 -549 521 -529
rect 744 -530 745 -470
rect 254 -549 255 -531
rect 275 -532 276 -470
rect 289 -532 290 -470
rect 380 -549 381 -531
rect 436 -532 437 -470
rect 569 -549 570 -531
rect 611 -532 612 -470
rect 625 -549 626 -531
rect 744 -549 745 -531
rect 758 -532 759 -470
rect 205 -534 206 -470
rect 275 -549 276 -533
rect 289 -549 290 -533
rect 331 -534 332 -470
rect 453 -549 454 -533
rect 611 -549 612 -533
rect 730 -534 731 -470
rect 758 -549 759 -533
rect 72 -536 73 -470
rect 205 -549 206 -535
rect 268 -549 269 -535
rect 310 -549 311 -535
rect 457 -536 458 -470
rect 681 -549 682 -535
rect 730 -549 731 -535
rect 828 -536 829 -470
rect 72 -549 73 -537
rect 450 -538 451 -470
rect 457 -549 458 -537
rect 478 -538 479 -470
rect 499 -549 500 -537
rect 863 -538 864 -470
rect 450 -549 451 -539
rect 495 -549 496 -539
rect 527 -549 528 -539
rect 562 -540 563 -470
rect 478 -549 479 -541
rect 723 -542 724 -470
rect 555 -544 556 -470
rect 562 -549 563 -543
rect 723 -549 724 -543
rect 877 -544 878 -470
rect 261 -546 262 -470
rect 555 -549 556 -545
rect 261 -549 262 -547
rect 436 -549 437 -547
rect 2 -559 3 -557
rect 481 -559 482 -557
rect 502 -559 503 -557
rect 576 -559 577 -557
rect 583 -559 584 -557
rect 604 -632 605 -558
rect 607 -559 608 -557
rect 625 -559 626 -557
rect 681 -559 682 -557
rect 898 -632 899 -558
rect 2 -632 3 -560
rect 30 -561 31 -557
rect 37 -561 38 -557
rect 96 -561 97 -557
rect 107 -561 108 -557
rect 107 -632 108 -560
rect 107 -561 108 -557
rect 107 -632 108 -560
rect 131 -632 132 -560
rect 163 -632 164 -560
rect 177 -561 178 -557
rect 317 -561 318 -557
rect 345 -561 346 -557
rect 362 -561 363 -557
rect 373 -561 374 -557
rect 495 -561 496 -557
rect 506 -632 507 -560
rect 537 -632 538 -560
rect 541 -632 542 -560
rect 828 -632 829 -560
rect 835 -561 836 -557
rect 842 -632 843 -560
rect 9 -563 10 -557
rect 124 -632 125 -562
rect 135 -563 136 -557
rect 331 -563 332 -557
rect 373 -632 374 -562
rect 401 -563 402 -557
rect 404 -632 405 -562
rect 884 -632 885 -562
rect 9 -632 10 -564
rect 86 -565 87 -557
rect 156 -632 157 -564
rect 243 -565 244 -557
rect 254 -565 255 -557
rect 254 -632 255 -564
rect 254 -565 255 -557
rect 254 -632 255 -564
rect 317 -632 318 -564
rect 523 -632 524 -564
rect 544 -565 545 -557
rect 905 -632 906 -564
rect 23 -567 24 -557
rect 180 -567 181 -557
rect 191 -567 192 -557
rect 341 -567 342 -557
rect 401 -632 402 -566
rect 478 -632 479 -566
rect 520 -567 521 -557
rect 625 -632 626 -566
rect 646 -567 647 -557
rect 835 -632 836 -566
rect 23 -632 24 -568
rect 51 -569 52 -557
rect 58 -569 59 -557
rect 261 -569 262 -557
rect 415 -632 416 -568
rect 450 -569 451 -557
rect 453 -569 454 -557
rect 527 -569 528 -557
rect 555 -569 556 -557
rect 726 -569 727 -557
rect 744 -569 745 -557
rect 751 -569 752 -557
rect 754 -569 755 -557
rect 926 -632 927 -568
rect 30 -632 31 -570
rect 306 -632 307 -570
rect 436 -571 437 -557
rect 509 -571 510 -557
rect 562 -571 563 -557
rect 576 -632 577 -570
rect 583 -632 584 -570
rect 597 -571 598 -557
rect 660 -571 661 -557
rect 681 -632 682 -570
rect 695 -571 696 -557
rect 751 -632 752 -570
rect 765 -571 766 -557
rect 849 -632 850 -570
rect 40 -632 41 -572
rect 341 -632 342 -572
rect 429 -573 430 -557
rect 436 -632 437 -572
rect 457 -573 458 -557
rect 555 -632 556 -572
rect 597 -632 598 -572
rect 688 -573 689 -557
rect 723 -573 724 -557
rect 947 -632 948 -572
rect 44 -632 45 -574
rect 86 -632 87 -574
rect 103 -632 104 -574
rect 261 -632 262 -574
rect 348 -632 349 -574
rect 429 -632 430 -574
rect 457 -632 458 -574
rect 513 -575 514 -557
rect 548 -575 549 -557
rect 562 -632 563 -574
rect 618 -575 619 -557
rect 723 -632 724 -574
rect 744 -632 745 -574
rect 758 -575 759 -557
rect 772 -575 773 -557
rect 891 -632 892 -574
rect 51 -632 52 -576
rect 121 -577 122 -557
rect 128 -577 129 -557
rect 548 -632 549 -576
rect 653 -577 654 -557
rect 660 -632 661 -576
rect 698 -632 699 -576
rect 772 -632 773 -576
rect 786 -577 787 -557
rect 912 -632 913 -576
rect 65 -579 66 -557
rect 68 -625 69 -578
rect 79 -579 80 -557
rect 390 -579 391 -557
rect 474 -632 475 -578
rect 632 -579 633 -557
rect 702 -579 703 -557
rect 758 -632 759 -578
rect 793 -579 794 -557
rect 856 -579 857 -557
rect 65 -632 66 -580
rect 313 -581 314 -557
rect 338 -581 339 -557
rect 786 -632 787 -580
rect 800 -581 801 -557
rect 870 -632 871 -580
rect 79 -632 80 -582
rect 184 -583 185 -557
rect 191 -632 192 -582
rect 331 -632 332 -582
rect 485 -583 486 -557
rect 765 -632 766 -582
rect 779 -583 780 -557
rect 856 -632 857 -582
rect 93 -585 94 -557
rect 793 -632 794 -584
rect 800 -632 801 -584
rect 807 -585 808 -557
rect 814 -585 815 -557
rect 863 -632 864 -584
rect 93 -632 94 -586
rect 100 -587 101 -557
rect 135 -632 136 -586
rect 688 -632 689 -586
rect 730 -587 731 -557
rect 807 -632 808 -586
rect 159 -589 160 -557
rect 240 -632 241 -588
rect 264 -589 265 -557
rect 730 -632 731 -588
rect 737 -589 738 -557
rect 814 -632 815 -588
rect 166 -591 167 -557
rect 646 -632 647 -590
rect 173 -632 174 -592
rect 177 -632 178 -592
rect 184 -632 185 -592
rect 198 -593 199 -557
rect 205 -593 206 -557
rect 877 -632 878 -592
rect 198 -632 199 -594
rect 296 -595 297 -557
rect 313 -632 314 -594
rect 443 -595 444 -557
rect 471 -595 472 -557
rect 779 -632 780 -594
rect 205 -632 206 -596
rect 219 -597 220 -557
rect 226 -597 227 -557
rect 527 -632 528 -596
rect 534 -597 535 -557
rect 653 -632 654 -596
rect 212 -599 213 -557
rect 282 -599 283 -557
rect 289 -599 290 -557
rect 443 -632 444 -598
rect 471 -632 472 -598
rect 590 -599 591 -557
rect 632 -632 633 -598
rect 667 -599 668 -557
rect 16 -601 17 -557
rect 212 -632 213 -600
rect 215 -601 216 -557
rect 345 -632 346 -600
rect 359 -601 360 -557
rect 485 -632 486 -600
rect 513 -632 514 -600
rect 544 -632 545 -600
rect 569 -601 570 -557
rect 737 -632 738 -600
rect 16 -632 17 -602
rect 61 -632 62 -602
rect 219 -632 220 -602
rect 233 -603 234 -557
rect 236 -632 237 -602
rect 422 -603 423 -557
rect 425 -603 426 -557
rect 667 -632 668 -602
rect 114 -605 115 -557
rect 422 -632 423 -604
rect 590 -632 591 -604
rect 674 -605 675 -557
rect 114 -632 115 -606
rect 170 -607 171 -557
rect 226 -632 227 -606
rect 268 -607 269 -557
rect 275 -607 276 -557
rect 296 -632 297 -606
rect 359 -632 360 -606
rect 366 -607 367 -557
rect 380 -607 381 -557
rect 569 -632 570 -606
rect 639 -607 640 -557
rect 702 -632 703 -606
rect 149 -609 150 -557
rect 233 -632 234 -608
rect 247 -609 248 -557
rect 268 -632 269 -608
rect 275 -632 276 -608
rect 499 -609 500 -557
rect 611 -609 612 -557
rect 639 -632 640 -608
rect 149 -632 150 -610
rect 324 -611 325 -557
rect 338 -632 339 -610
rect 380 -632 381 -610
rect 467 -632 468 -610
rect 499 -632 500 -610
rect 611 -632 612 -610
rect 716 -611 717 -557
rect 145 -613 146 -557
rect 324 -632 325 -612
rect 366 -632 367 -612
rect 394 -613 395 -557
rect 492 -613 493 -557
rect 674 -632 675 -612
rect 709 -613 710 -557
rect 716 -632 717 -612
rect 247 -632 248 -614
rect 387 -615 388 -557
rect 450 -632 451 -614
rect 709 -632 710 -614
rect 72 -617 73 -557
rect 387 -632 388 -616
rect 72 -632 73 -618
rect 310 -632 311 -618
rect 334 -632 335 -618
rect 492 -632 493 -618
rect 282 -632 283 -620
rect 303 -621 304 -557
rect 352 -621 353 -557
rect 394 -632 395 -620
rect 289 -632 290 -622
rect 408 -623 409 -557
rect 408 -632 409 -624
rect 352 -632 353 -626
rect 464 -627 465 -557
rect 464 -632 465 -628
rect 821 -629 822 -557
rect 593 -632 594 -630
rect 821 -632 822 -630
rect 2 -642 3 -640
rect 58 -642 59 -640
rect 61 -642 62 -640
rect 135 -642 136 -640
rect 138 -642 139 -640
rect 453 -642 454 -640
rect 464 -642 465 -640
rect 723 -642 724 -640
rect 821 -642 822 -640
rect 954 -711 955 -641
rect 2 -711 3 -643
rect 156 -644 157 -640
rect 173 -644 174 -640
rect 282 -644 283 -640
rect 289 -644 290 -640
rect 303 -644 304 -640
rect 331 -644 332 -640
rect 569 -644 570 -640
rect 590 -711 591 -643
rect 870 -644 871 -640
rect 947 -644 948 -640
rect 1031 -711 1032 -643
rect 16 -646 17 -640
rect 86 -646 87 -640
rect 93 -646 94 -640
rect 110 -711 111 -645
rect 184 -646 185 -640
rect 411 -711 412 -645
rect 436 -646 437 -640
rect 464 -711 465 -645
rect 488 -711 489 -645
rect 583 -646 584 -640
rect 593 -646 594 -640
rect 905 -646 906 -640
rect 16 -711 17 -647
rect 149 -648 150 -640
rect 184 -711 185 -647
rect 268 -648 269 -640
rect 289 -711 290 -647
rect 394 -648 395 -640
rect 404 -648 405 -640
rect 555 -648 556 -640
rect 562 -648 563 -640
rect 569 -711 570 -647
rect 583 -711 584 -647
rect 632 -648 633 -640
rect 660 -648 661 -640
rect 695 -711 696 -647
rect 793 -648 794 -640
rect 821 -711 822 -647
rect 891 -648 892 -640
rect 905 -711 906 -647
rect 37 -711 38 -649
rect 334 -711 335 -649
rect 338 -650 339 -640
rect 366 -650 367 -640
rect 387 -650 388 -640
rect 450 -711 451 -649
rect 481 -711 482 -649
rect 593 -711 594 -649
rect 604 -650 605 -640
rect 618 -711 619 -649
rect 621 -650 622 -640
rect 758 -650 759 -640
rect 786 -650 787 -640
rect 793 -711 794 -649
rect 814 -650 815 -640
rect 870 -711 871 -649
rect 51 -652 52 -640
rect 471 -652 472 -640
rect 502 -711 503 -651
rect 807 -652 808 -640
rect 828 -652 829 -640
rect 891 -711 892 -651
rect 30 -654 31 -640
rect 471 -711 472 -653
rect 513 -654 514 -640
rect 534 -711 535 -653
rect 537 -654 538 -640
rect 765 -654 766 -640
rect 779 -654 780 -640
rect 786 -711 787 -653
rect 51 -711 52 -655
rect 478 -656 479 -640
rect 520 -656 521 -640
rect 912 -656 913 -640
rect 58 -711 59 -657
rect 177 -658 178 -640
rect 198 -658 199 -640
rect 268 -711 269 -657
rect 338 -711 339 -657
rect 474 -658 475 -640
rect 506 -658 507 -640
rect 520 -711 521 -657
rect 523 -658 524 -640
rect 597 -658 598 -640
rect 611 -658 612 -640
rect 814 -711 815 -657
rect 912 -711 913 -657
rect 926 -658 927 -640
rect 65 -660 66 -640
rect 156 -711 157 -659
rect 177 -711 178 -659
rect 275 -660 276 -640
rect 341 -660 342 -640
rect 373 -660 374 -640
rect 436 -711 437 -659
rect 544 -711 545 -659
rect 551 -711 552 -659
rect 702 -660 703 -640
rect 716 -660 717 -640
rect 779 -711 780 -659
rect 65 -711 66 -661
rect 121 -662 122 -640
rect 149 -711 150 -661
rect 191 -662 192 -640
rect 198 -711 199 -661
rect 219 -662 220 -640
rect 233 -711 234 -661
rect 317 -662 318 -640
rect 345 -711 346 -661
rect 527 -662 528 -640
rect 541 -662 542 -640
rect 709 -662 710 -640
rect 730 -662 731 -640
rect 926 -711 927 -661
rect 72 -664 73 -640
rect 317 -711 318 -663
rect 359 -664 360 -640
rect 394 -711 395 -663
rect 408 -664 409 -640
rect 527 -711 528 -663
rect 541 -711 542 -663
rect 856 -664 857 -640
rect 72 -711 73 -665
rect 443 -666 444 -640
rect 474 -711 475 -665
rect 828 -711 829 -665
rect 79 -668 80 -640
rect 243 -668 244 -640
rect 247 -668 248 -640
rect 282 -711 283 -667
rect 366 -711 367 -667
rect 401 -668 402 -640
rect 443 -711 444 -667
rect 467 -668 468 -640
rect 499 -668 500 -640
rect 506 -711 507 -667
rect 555 -711 556 -667
rect 737 -668 738 -640
rect 765 -711 766 -667
rect 835 -668 836 -640
rect 9 -670 10 -640
rect 243 -711 244 -669
rect 250 -711 251 -669
rect 254 -670 255 -640
rect 275 -711 276 -669
rect 415 -670 416 -640
rect 478 -711 479 -669
rect 737 -711 738 -669
rect 9 -711 10 -671
rect 44 -672 45 -640
rect 79 -711 80 -671
rect 380 -672 381 -640
rect 390 -711 391 -671
rect 835 -711 836 -671
rect 23 -674 24 -640
rect 44 -711 45 -673
rect 86 -711 87 -673
rect 856 -711 857 -673
rect 93 -711 94 -675
rect 145 -676 146 -640
rect 170 -676 171 -640
rect 191 -711 192 -675
rect 205 -676 206 -640
rect 303 -711 304 -675
rect 324 -676 325 -640
rect 401 -711 402 -675
rect 562 -711 563 -675
rect 849 -676 850 -640
rect 100 -678 101 -640
rect 548 -678 549 -640
rect 576 -678 577 -640
rect 604 -711 605 -677
rect 614 -678 615 -640
rect 919 -678 920 -640
rect 103 -680 104 -640
rect 611 -711 612 -679
rect 625 -680 626 -640
rect 632 -711 633 -679
rect 639 -680 640 -640
rect 660 -711 661 -679
rect 667 -680 668 -640
rect 919 -711 920 -679
rect 100 -711 101 -681
rect 667 -711 668 -681
rect 674 -682 675 -640
rect 723 -711 724 -681
rect 730 -711 731 -681
rect 800 -682 801 -640
rect 842 -682 843 -640
rect 849 -711 850 -681
rect 103 -711 104 -683
rect 142 -684 143 -640
rect 170 -711 171 -683
rect 261 -684 262 -640
rect 324 -711 325 -683
rect 429 -684 430 -640
rect 576 -711 577 -683
rect 625 -711 626 -683
rect 639 -711 640 -683
rect 887 -711 888 -683
rect 107 -686 108 -640
rect 128 -686 129 -640
rect 205 -711 206 -685
rect 254 -711 255 -685
rect 261 -711 262 -685
rect 310 -686 311 -640
rect 352 -686 353 -640
rect 415 -711 416 -685
rect 422 -686 423 -640
rect 429 -711 430 -685
rect 646 -686 647 -640
rect 674 -711 675 -685
rect 688 -686 689 -640
rect 758 -711 759 -685
rect 772 -686 773 -640
rect 800 -711 801 -685
rect 842 -711 843 -685
rect 877 -686 878 -640
rect 114 -688 115 -640
rect 310 -711 311 -687
rect 352 -711 353 -687
rect 628 -711 629 -687
rect 653 -688 654 -640
rect 702 -711 703 -687
rect 751 -688 752 -640
rect 772 -711 773 -687
rect 877 -711 878 -687
rect 898 -688 899 -640
rect 89 -711 90 -689
rect 114 -711 115 -689
rect 121 -711 122 -689
rect 163 -690 164 -640
rect 212 -690 213 -640
rect 597 -711 598 -689
rect 744 -690 745 -640
rect 751 -711 752 -689
rect 863 -690 864 -640
rect 898 -711 899 -689
rect 135 -711 136 -691
rect 212 -711 213 -691
rect 219 -711 220 -691
rect 296 -692 297 -640
rect 380 -711 381 -691
rect 457 -692 458 -640
rect 485 -692 486 -640
rect 646 -711 647 -691
rect 681 -692 682 -640
rect 744 -711 745 -691
rect 863 -711 864 -691
rect 884 -692 885 -640
rect 145 -711 146 -693
rect 688 -711 689 -693
rect 163 -711 164 -695
rect 565 -711 566 -695
rect 226 -698 227 -640
rect 408 -711 409 -697
rect 422 -711 423 -697
rect 548 -711 549 -697
rect 558 -711 559 -697
rect 681 -711 682 -697
rect 229 -711 230 -699
rect 457 -711 458 -699
rect 485 -711 486 -699
rect 716 -711 717 -699
rect 236 -702 237 -640
rect 709 -711 710 -701
rect 240 -704 241 -640
rect 359 -711 360 -703
rect 492 -704 493 -640
rect 653 -711 654 -703
rect 240 -711 241 -705
rect 807 -711 808 -705
rect 296 -711 297 -707
rect 418 -711 419 -707
rect 348 -711 349 -709
rect 492 -711 493 -709
rect 16 -721 17 -719
rect 103 -721 104 -719
rect 135 -721 136 -719
rect 390 -782 391 -720
rect 415 -721 416 -719
rect 765 -721 766 -719
rect 849 -721 850 -719
rect 884 -782 885 -720
rect 908 -782 909 -720
rect 912 -721 913 -719
rect 926 -721 927 -719
rect 975 -782 976 -720
rect 1006 -782 1007 -720
rect 1017 -782 1018 -720
rect 1031 -721 1032 -719
rect 1066 -782 1067 -720
rect 23 -782 24 -722
rect 117 -782 118 -722
rect 135 -782 136 -722
rect 149 -723 150 -719
rect 170 -723 171 -719
rect 418 -723 419 -719
rect 478 -723 479 -719
rect 544 -723 545 -719
rect 551 -723 552 -719
rect 856 -723 857 -719
rect 912 -782 913 -722
rect 961 -782 962 -722
rect 26 -725 27 -719
rect 30 -725 31 -719
rect 33 -725 34 -719
rect 670 -782 671 -724
rect 716 -725 717 -719
rect 765 -782 766 -724
rect 793 -725 794 -719
rect 849 -782 850 -724
rect 954 -725 955 -719
rect 1010 -782 1011 -724
rect 30 -782 31 -726
rect 163 -727 164 -719
rect 170 -782 171 -726
rect 187 -782 188 -726
rect 229 -727 230 -719
rect 310 -727 311 -719
rect 317 -727 318 -719
rect 387 -727 388 -719
rect 464 -727 465 -719
rect 478 -782 479 -726
rect 481 -727 482 -719
rect 583 -727 584 -719
rect 590 -727 591 -719
rect 716 -782 717 -726
rect 744 -727 745 -719
rect 793 -782 794 -726
rect 807 -727 808 -719
rect 856 -782 857 -726
rect 44 -729 45 -719
rect 110 -729 111 -719
rect 128 -729 129 -719
rect 387 -782 388 -728
rect 436 -729 437 -719
rect 464 -782 465 -728
rect 488 -729 489 -719
rect 534 -729 535 -719
rect 555 -782 556 -728
rect 835 -729 836 -719
rect 2 -731 3 -719
rect 44 -782 45 -730
rect 58 -731 59 -719
rect 205 -731 206 -719
rect 240 -731 241 -719
rect 541 -731 542 -719
rect 558 -731 559 -719
rect 891 -731 892 -719
rect 58 -782 59 -732
rect 191 -733 192 -719
rect 205 -782 206 -732
rect 233 -733 234 -719
rect 247 -782 248 -732
rect 338 -733 339 -719
rect 348 -733 349 -719
rect 492 -733 493 -719
rect 516 -733 517 -719
rect 653 -733 654 -719
rect 674 -733 675 -719
rect 744 -782 745 -732
rect 779 -733 780 -719
rect 807 -782 808 -732
rect 891 -782 892 -732
rect 915 -782 916 -732
rect 86 -735 87 -719
rect 597 -735 598 -719
rect 621 -782 622 -734
rect 905 -735 906 -719
rect 86 -782 87 -736
rect 282 -737 283 -719
rect 317 -782 318 -736
rect 499 -737 500 -719
rect 506 -737 507 -719
rect 597 -782 598 -736
rect 625 -737 626 -719
rect 898 -737 899 -719
rect 51 -739 52 -719
rect 506 -782 507 -738
rect 527 -739 528 -719
rect 548 -782 549 -738
rect 565 -782 566 -738
rect 800 -739 801 -719
rect 898 -782 899 -738
rect 919 -739 920 -719
rect 65 -741 66 -719
rect 499 -782 500 -740
rect 541 -782 542 -740
rect 674 -782 675 -740
rect 723 -741 724 -719
rect 779 -782 780 -740
rect 814 -741 815 -719
rect 919 -782 920 -740
rect 89 -743 90 -719
rect 667 -743 668 -719
rect 688 -743 689 -719
rect 723 -782 724 -742
rect 737 -743 738 -719
rect 835 -782 836 -742
rect 93 -745 94 -719
rect 243 -745 244 -719
rect 254 -745 255 -719
rect 355 -782 356 -744
rect 373 -745 374 -719
rect 821 -745 822 -719
rect 51 -782 52 -746
rect 93 -782 94 -746
rect 128 -782 129 -746
rect 495 -782 496 -746
rect 569 -747 570 -719
rect 590 -782 591 -746
rect 625 -782 626 -746
rect 639 -747 640 -719
rect 667 -782 668 -746
rect 730 -747 731 -719
rect 758 -747 759 -719
rect 800 -782 801 -746
rect 821 -782 822 -746
rect 828 -747 829 -719
rect 72 -749 73 -719
rect 373 -782 374 -748
rect 394 -749 395 -719
rect 534 -782 535 -748
rect 569 -782 570 -748
rect 576 -749 577 -719
rect 579 -782 580 -748
rect 772 -749 773 -719
rect 142 -751 143 -719
rect 219 -751 220 -719
rect 261 -751 262 -719
rect 264 -782 265 -750
rect 268 -751 269 -719
rect 282 -782 283 -750
rect 331 -782 332 -750
rect 429 -751 430 -719
rect 436 -782 437 -750
rect 457 -751 458 -719
rect 485 -751 486 -719
rect 653 -782 654 -750
rect 660 -751 661 -719
rect 730 -782 731 -750
rect 9 -753 10 -719
rect 457 -782 458 -752
rect 527 -782 528 -752
rect 828 -782 829 -752
rect 107 -755 108 -719
rect 268 -782 269 -754
rect 296 -755 297 -719
rect 429 -782 430 -754
rect 576 -782 577 -754
rect 772 -782 773 -754
rect 107 -782 108 -756
rect 114 -757 115 -719
rect 142 -782 143 -756
rect 352 -757 353 -719
rect 380 -757 381 -719
rect 485 -782 486 -756
rect 583 -782 584 -756
rect 604 -757 605 -719
rect 628 -757 629 -719
rect 870 -757 871 -719
rect 100 -759 101 -719
rect 114 -782 115 -758
rect 145 -759 146 -719
rect 149 -782 150 -758
rect 156 -759 157 -719
rect 163 -782 164 -758
rect 191 -782 192 -758
rect 250 -759 251 -719
rect 254 -782 255 -758
rect 261 -782 262 -758
rect 296 -782 297 -758
rect 345 -759 346 -719
rect 359 -759 360 -719
rect 380 -782 381 -758
rect 394 -782 395 -758
rect 401 -759 402 -719
rect 415 -782 416 -758
rect 814 -782 815 -758
rect 842 -759 843 -719
rect 870 -782 871 -758
rect 100 -782 101 -760
rect 408 -761 409 -719
rect 639 -782 640 -760
rect 646 -761 647 -719
rect 688 -782 689 -760
rect 751 -761 752 -719
rect 786 -761 787 -719
rect 842 -782 843 -760
rect 156 -782 157 -762
rect 198 -763 199 -719
rect 212 -763 213 -719
rect 219 -782 220 -762
rect 236 -782 237 -762
rect 660 -782 661 -762
rect 702 -763 703 -719
rect 737 -782 738 -762
rect 751 -782 752 -762
rect 877 -763 878 -719
rect 37 -765 38 -719
rect 212 -782 213 -764
rect 243 -782 244 -764
rect 359 -782 360 -764
rect 408 -782 409 -764
rect 443 -765 444 -719
rect 450 -765 451 -719
rect 646 -782 647 -764
rect 681 -765 682 -719
rect 702 -782 703 -764
rect 709 -765 710 -719
rect 758 -782 759 -764
rect 863 -765 864 -719
rect 877 -782 878 -764
rect 37 -782 38 -766
rect 513 -767 514 -719
rect 520 -767 521 -719
rect 681 -782 682 -766
rect 695 -767 696 -719
rect 709 -782 710 -766
rect 177 -769 178 -719
rect 198 -782 199 -768
rect 275 -769 276 -719
rect 401 -782 402 -768
rect 404 -782 405 -768
rect 443 -782 444 -768
rect 450 -782 451 -768
rect 530 -782 531 -768
rect 611 -769 612 -719
rect 695 -782 696 -768
rect 79 -771 80 -719
rect 275 -782 276 -770
rect 289 -771 290 -719
rect 520 -782 521 -770
rect 562 -771 563 -719
rect 611 -782 612 -770
rect 632 -771 633 -719
rect 786 -782 787 -770
rect 79 -782 80 -772
rect 376 -773 377 -719
rect 492 -782 493 -772
rect 863 -782 864 -772
rect 177 -782 178 -774
rect 184 -775 185 -719
rect 289 -782 290 -774
rect 303 -775 304 -719
rect 324 -775 325 -719
rect 352 -782 353 -774
rect 513 -782 514 -774
rect 604 -782 605 -774
rect 618 -775 619 -719
rect 632 -782 633 -774
rect 121 -777 122 -719
rect 184 -782 185 -776
rect 310 -782 311 -776
rect 324 -782 325 -776
rect 338 -782 339 -776
rect 366 -777 367 -719
rect 471 -782 472 -776
rect 618 -782 619 -776
rect 110 -782 111 -778
rect 121 -782 122 -778
rect 131 -779 132 -719
rect 303 -782 304 -778
rect 345 -782 346 -778
rect 502 -779 503 -719
rect 366 -782 367 -780
rect 422 -781 423 -719
rect 16 -879 17 -791
rect 65 -792 66 -790
rect 68 -879 69 -791
rect 110 -792 111 -790
rect 114 -792 115 -790
rect 243 -879 244 -791
rect 310 -879 311 -791
rect 369 -879 370 -791
rect 387 -792 388 -790
rect 947 -879 948 -791
rect 961 -792 962 -790
rect 1013 -879 1014 -791
rect 1017 -792 1018 -790
rect 1024 -879 1025 -791
rect 1066 -792 1067 -790
rect 1080 -879 1081 -791
rect 23 -794 24 -790
rect 72 -794 73 -790
rect 79 -794 80 -790
rect 180 -879 181 -793
rect 233 -794 234 -790
rect 303 -794 304 -790
rect 338 -879 339 -793
rect 450 -794 451 -790
rect 492 -794 493 -790
rect 744 -794 745 -790
rect 814 -794 815 -790
rect 954 -879 955 -793
rect 975 -794 976 -790
rect 1017 -879 1018 -793
rect 23 -879 24 -795
rect 149 -796 150 -790
rect 173 -879 174 -795
rect 362 -879 363 -795
rect 411 -879 412 -795
rect 520 -796 521 -790
rect 523 -879 524 -795
rect 849 -796 850 -790
rect 863 -796 864 -790
rect 933 -879 934 -795
rect 989 -796 990 -790
rect 992 -879 993 -795
rect 1010 -796 1011 -790
rect 1038 -879 1039 -795
rect 30 -798 31 -790
rect 313 -798 314 -790
rect 380 -798 381 -790
rect 520 -879 521 -797
rect 530 -798 531 -790
rect 639 -798 640 -790
rect 653 -798 654 -790
rect 849 -879 850 -797
rect 877 -798 878 -790
rect 996 -879 997 -797
rect 37 -800 38 -790
rect 184 -800 185 -790
rect 233 -879 234 -799
rect 296 -800 297 -790
rect 380 -879 381 -799
rect 541 -879 542 -799
rect 551 -879 552 -799
rect 653 -879 654 -799
rect 695 -800 696 -790
rect 894 -800 895 -790
rect 915 -800 916 -790
rect 1003 -879 1004 -799
rect 37 -879 38 -801
rect 226 -802 227 -790
rect 240 -802 241 -790
rect 289 -802 290 -790
rect 296 -879 297 -801
rect 576 -802 577 -790
rect 618 -802 619 -790
rect 786 -802 787 -790
rect 817 -879 818 -801
rect 961 -879 962 -801
rect 44 -804 45 -790
rect 236 -804 237 -790
rect 254 -804 255 -790
rect 576 -879 577 -803
rect 621 -804 622 -790
rect 898 -804 899 -790
rect 919 -804 920 -790
rect 919 -879 920 -803
rect 919 -804 920 -790
rect 919 -879 920 -803
rect 47 -879 48 -805
rect 261 -806 262 -790
rect 268 -806 269 -790
rect 303 -879 304 -805
rect 422 -806 423 -790
rect 968 -879 969 -805
rect 51 -879 52 -807
rect 229 -808 230 -790
rect 254 -879 255 -807
rect 317 -808 318 -790
rect 422 -879 423 -807
rect 429 -808 430 -790
rect 439 -879 440 -807
rect 912 -879 913 -807
rect 30 -879 31 -809
rect 229 -879 230 -809
rect 261 -879 262 -809
rect 527 -810 528 -790
rect 537 -879 538 -809
rect 751 -810 752 -790
rect 800 -810 801 -790
rect 898 -879 899 -809
rect 58 -812 59 -790
rect 352 -812 353 -790
rect 429 -879 430 -811
rect 737 -812 738 -790
rect 751 -879 752 -811
rect 905 -812 906 -790
rect 12 -879 13 -813
rect 58 -879 59 -813
rect 72 -879 73 -813
rect 142 -814 143 -790
rect 149 -879 150 -813
rect 219 -814 220 -790
rect 282 -814 283 -790
rect 352 -879 353 -813
rect 450 -879 451 -813
rect 478 -814 479 -790
rect 485 -814 486 -790
rect 527 -879 528 -813
rect 544 -879 545 -813
rect 618 -879 619 -813
rect 639 -879 640 -813
rect 989 -879 990 -813
rect 79 -879 80 -815
rect 467 -879 468 -815
rect 471 -816 472 -790
rect 485 -879 486 -815
rect 492 -879 493 -815
rect 744 -879 745 -815
rect 821 -816 822 -790
rect 982 -879 983 -815
rect 86 -818 87 -790
rect 425 -818 426 -790
rect 443 -818 444 -790
rect 471 -879 472 -817
rect 478 -879 479 -817
rect 667 -818 668 -790
rect 681 -818 682 -790
rect 737 -879 738 -817
rect 765 -818 766 -790
rect 821 -879 822 -817
rect 828 -818 829 -790
rect 975 -879 976 -817
rect 86 -879 87 -819
rect 93 -820 94 -790
rect 114 -879 115 -819
rect 408 -820 409 -790
rect 499 -820 500 -790
rect 681 -879 682 -819
rect 695 -879 696 -819
rect 814 -879 815 -819
rect 828 -879 829 -819
rect 884 -820 885 -790
rect 891 -820 892 -790
rect 891 -879 892 -819
rect 891 -820 892 -790
rect 891 -879 892 -819
rect 93 -879 94 -821
rect 163 -822 164 -790
rect 184 -879 185 -821
rect 345 -822 346 -790
rect 506 -822 507 -790
rect 506 -879 507 -821
rect 506 -822 507 -790
rect 506 -879 507 -821
rect 513 -822 514 -790
rect 590 -822 591 -790
rect 667 -879 668 -821
rect 688 -822 689 -790
rect 709 -822 710 -790
rect 709 -879 710 -821
rect 709 -822 710 -790
rect 709 -879 710 -821
rect 716 -822 717 -790
rect 863 -879 864 -821
rect 121 -824 122 -790
rect 401 -879 402 -823
rect 513 -879 514 -823
rect 625 -824 626 -790
rect 723 -824 724 -790
rect 765 -879 766 -823
rect 835 -824 836 -790
rect 940 -879 941 -823
rect 121 -879 122 -825
rect 135 -826 136 -790
rect 138 -879 139 -825
rect 191 -826 192 -790
rect 205 -826 206 -790
rect 282 -879 283 -825
rect 289 -879 290 -825
rect 366 -826 367 -790
rect 373 -826 374 -790
rect 723 -879 724 -825
rect 730 -826 731 -790
rect 908 -826 909 -790
rect 2 -879 3 -827
rect 205 -879 206 -827
rect 219 -879 220 -827
rect 674 -828 675 -790
rect 772 -828 773 -790
rect 835 -879 836 -827
rect 128 -830 129 -790
rect 317 -879 318 -829
rect 345 -879 346 -829
rect 415 -830 416 -790
rect 516 -830 517 -790
rect 632 -830 633 -790
rect 660 -830 661 -790
rect 674 -879 675 -829
rect 772 -879 773 -829
rect 807 -830 808 -790
rect 110 -879 111 -831
rect 660 -879 661 -831
rect 670 -879 671 -831
rect 730 -879 731 -831
rect 758 -832 759 -790
rect 807 -879 808 -831
rect 117 -879 118 -833
rect 632 -879 633 -833
rect 702 -834 703 -790
rect 758 -879 759 -833
rect 131 -879 132 -835
rect 856 -836 857 -790
rect 135 -879 136 -837
rect 877 -879 878 -837
rect 142 -879 143 -839
rect 198 -840 199 -790
rect 240 -879 241 -839
rect 443 -879 444 -839
rect 534 -840 535 -790
rect 716 -879 717 -839
rect 163 -879 164 -841
rect 170 -842 171 -790
rect 191 -879 192 -841
rect 247 -842 248 -790
rect 268 -879 269 -841
rect 408 -879 409 -841
rect 415 -879 416 -841
rect 597 -842 598 -790
rect 604 -842 605 -790
rect 688 -879 689 -841
rect 156 -844 157 -790
rect 247 -879 248 -843
rect 324 -844 325 -790
rect 604 -879 605 -843
rect 611 -844 612 -790
rect 625 -879 626 -843
rect 100 -846 101 -790
rect 324 -879 325 -845
rect 355 -846 356 -790
rect 702 -879 703 -845
rect 100 -879 101 -847
rect 331 -848 332 -790
rect 355 -879 356 -847
rect 870 -848 871 -790
rect 156 -879 157 -849
rect 208 -879 209 -849
rect 331 -879 332 -849
rect 394 -850 395 -790
rect 457 -850 458 -790
rect 597 -879 598 -849
rect 793 -850 794 -790
rect 870 -879 871 -849
rect 170 -879 171 -851
rect 177 -852 178 -790
rect 198 -879 199 -851
rect 212 -852 213 -790
rect 275 -852 276 -790
rect 394 -879 395 -851
rect 457 -879 458 -851
rect 464 -852 465 -790
rect 548 -852 549 -790
rect 793 -879 794 -851
rect 177 -879 178 -853
rect 387 -879 388 -853
rect 464 -879 465 -853
rect 926 -879 927 -853
rect 212 -879 213 -855
rect 800 -879 801 -855
rect 366 -879 367 -857
rect 572 -879 573 -857
rect 579 -858 580 -790
rect 905 -879 906 -857
rect 373 -879 374 -859
rect 534 -879 535 -859
rect 548 -879 549 -859
rect 611 -879 612 -859
rect 555 -862 556 -790
rect 856 -879 857 -861
rect 359 -864 360 -790
rect 555 -879 556 -863
rect 562 -864 563 -790
rect 884 -879 885 -863
rect 275 -879 276 -865
rect 359 -879 360 -865
rect 565 -866 566 -790
rect 786 -879 787 -865
rect 565 -879 566 -867
rect 842 -868 843 -790
rect 583 -870 584 -790
rect 590 -879 591 -869
rect 779 -870 780 -790
rect 842 -879 843 -869
rect 436 -872 437 -790
rect 583 -879 584 -871
rect 436 -879 437 -873
rect 646 -874 647 -790
rect 562 -879 563 -875
rect 779 -879 780 -875
rect 569 -878 570 -790
rect 646 -879 647 -877
rect 16 -889 17 -887
rect 114 -889 115 -887
rect 121 -889 122 -887
rect 121 -960 122 -888
rect 121 -889 122 -887
rect 121 -960 122 -888
rect 135 -960 136 -888
rect 331 -889 332 -887
rect 359 -960 360 -888
rect 583 -889 584 -887
rect 600 -960 601 -888
rect 870 -889 871 -887
rect 915 -960 916 -888
rect 919 -889 920 -887
rect 947 -889 948 -887
rect 947 -960 948 -888
rect 947 -889 948 -887
rect 947 -960 948 -888
rect 954 -889 955 -887
rect 992 -889 993 -887
rect 1013 -889 1014 -887
rect 1024 -889 1025 -887
rect 1038 -889 1039 -887
rect 1059 -960 1060 -888
rect 1080 -889 1081 -887
rect 1087 -960 1088 -888
rect 16 -960 17 -890
rect 170 -891 171 -887
rect 184 -891 185 -887
rect 355 -891 356 -887
rect 366 -891 367 -887
rect 681 -891 682 -887
rect 807 -891 808 -887
rect 807 -960 808 -890
rect 807 -891 808 -887
rect 807 -960 808 -890
rect 814 -960 815 -890
rect 821 -891 822 -887
rect 870 -960 871 -890
rect 996 -891 997 -887
rect 1010 -891 1011 -887
rect 1038 -960 1039 -890
rect 23 -893 24 -887
rect 226 -960 227 -892
rect 243 -893 244 -887
rect 275 -893 276 -887
rect 289 -893 290 -887
rect 331 -960 332 -892
rect 366 -960 367 -892
rect 422 -893 423 -887
rect 429 -893 430 -887
rect 530 -960 531 -892
rect 534 -893 535 -887
rect 779 -893 780 -887
rect 817 -893 818 -887
rect 828 -893 829 -887
rect 961 -893 962 -887
rect 1010 -960 1011 -892
rect 2 -895 3 -887
rect 23 -960 24 -894
rect 51 -895 52 -887
rect 418 -960 419 -894
rect 422 -960 423 -894
rect 523 -895 524 -887
rect 534 -960 535 -894
rect 555 -895 556 -887
rect 569 -895 570 -887
rect 898 -895 899 -887
rect 961 -960 962 -894
rect 968 -895 969 -887
rect 989 -895 990 -887
rect 1017 -895 1018 -887
rect 51 -960 52 -896
rect 149 -897 150 -887
rect 156 -897 157 -887
rect 184 -960 185 -896
rect 205 -960 206 -896
rect 275 -960 276 -896
rect 289 -960 290 -896
rect 352 -897 353 -887
rect 369 -897 370 -887
rect 513 -897 514 -887
rect 520 -897 521 -887
rect 786 -897 787 -887
rect 828 -960 829 -896
rect 849 -897 850 -887
rect 891 -897 892 -887
rect 898 -960 899 -896
rect 968 -960 969 -896
rect 975 -897 976 -887
rect 58 -899 59 -887
rect 215 -899 216 -887
rect 219 -960 220 -898
rect 737 -899 738 -887
rect 765 -899 766 -887
rect 786 -960 787 -898
rect 849 -960 850 -898
rect 884 -899 885 -887
rect 891 -960 892 -898
rect 926 -899 927 -887
rect 58 -960 59 -900
rect 387 -901 388 -887
rect 408 -901 409 -887
rect 450 -901 451 -887
rect 464 -960 465 -900
rect 471 -901 472 -887
rect 474 -960 475 -900
rect 793 -901 794 -887
rect 884 -960 885 -900
rect 933 -901 934 -887
rect 65 -960 66 -902
rect 338 -903 339 -887
rect 352 -960 353 -902
rect 373 -903 374 -887
rect 387 -960 388 -902
rect 394 -903 395 -887
rect 408 -960 409 -902
rect 576 -903 577 -887
rect 628 -960 629 -902
rect 800 -903 801 -887
rect 933 -960 934 -902
rect 940 -903 941 -887
rect 72 -905 73 -887
rect 229 -905 230 -887
rect 278 -960 279 -904
rect 520 -960 521 -904
rect 527 -905 528 -887
rect 576 -960 577 -904
rect 730 -905 731 -887
rect 821 -960 822 -904
rect 72 -960 73 -906
rect 310 -907 311 -887
rect 317 -907 318 -887
rect 492 -907 493 -887
rect 499 -907 500 -887
rect 716 -907 717 -887
rect 737 -960 738 -906
rect 744 -907 745 -887
rect 751 -907 752 -887
rect 793 -960 794 -906
rect 800 -960 801 -906
rect 842 -907 843 -887
rect 93 -909 94 -887
rect 240 -909 241 -887
rect 261 -909 262 -887
rect 317 -960 318 -908
rect 324 -909 325 -887
rect 338 -960 339 -908
rect 345 -909 346 -887
rect 492 -960 493 -908
rect 499 -960 500 -908
rect 506 -909 507 -887
rect 537 -909 538 -887
rect 541 -960 542 -908
rect 548 -909 549 -887
rect 982 -909 983 -887
rect 93 -960 94 -910
rect 597 -911 598 -887
rect 635 -960 636 -910
rect 730 -960 731 -910
rect 765 -960 766 -910
rect 835 -911 836 -887
rect 842 -960 843 -910
rect 856 -911 857 -887
rect 905 -911 906 -887
rect 982 -960 983 -910
rect 107 -913 108 -887
rect 611 -913 612 -887
rect 688 -913 689 -887
rect 716 -960 717 -912
rect 723 -913 724 -887
rect 744 -960 745 -912
rect 779 -960 780 -912
rect 943 -960 944 -912
rect 107 -960 108 -914
rect 240 -960 241 -914
rect 261 -960 262 -914
rect 303 -915 304 -887
rect 310 -960 311 -914
rect 562 -915 563 -887
rect 597 -960 598 -914
rect 667 -960 668 -914
rect 702 -915 703 -887
rect 723 -960 724 -914
rect 856 -960 857 -914
rect 863 -915 864 -887
rect 905 -960 906 -914
rect 912 -915 913 -887
rect 110 -917 111 -887
rect 254 -917 255 -887
rect 285 -960 286 -916
rect 303 -960 304 -916
rect 373 -960 374 -916
rect 572 -917 573 -887
rect 604 -917 605 -887
rect 611 -960 612 -916
rect 653 -917 654 -887
rect 702 -960 703 -916
rect 709 -917 710 -887
rect 751 -960 752 -916
rect 863 -960 864 -916
rect 877 -917 878 -887
rect 912 -960 913 -916
rect 922 -960 923 -916
rect 114 -960 115 -918
rect 191 -919 192 -887
rect 198 -919 199 -887
rect 254 -960 255 -918
rect 411 -919 412 -887
rect 709 -960 710 -918
rect 149 -960 150 -920
rect 163 -921 164 -887
rect 170 -960 171 -920
rect 236 -960 237 -920
rect 429 -960 430 -920
rect 457 -921 458 -887
rect 467 -921 468 -887
rect 646 -921 647 -887
rect 660 -921 661 -887
rect 688 -960 689 -920
rect 30 -923 31 -887
rect 163 -960 164 -922
rect 180 -923 181 -887
rect 324 -960 325 -922
rect 436 -923 437 -887
rect 548 -960 549 -922
rect 551 -923 552 -887
rect 590 -923 591 -887
rect 639 -923 640 -887
rect 646 -960 647 -922
rect 660 -960 661 -922
rect 674 -923 675 -887
rect 30 -960 31 -924
rect 215 -960 216 -924
rect 439 -925 440 -887
rect 929 -960 930 -924
rect 86 -927 87 -887
rect 180 -960 181 -926
rect 191 -960 192 -926
rect 233 -927 234 -887
rect 439 -960 440 -926
rect 506 -960 507 -926
rect 513 -960 514 -926
rect 590 -960 591 -926
rect 625 -927 626 -887
rect 674 -960 675 -926
rect 86 -960 87 -928
rect 142 -929 143 -887
rect 156 -960 157 -928
rect 268 -929 269 -887
rect 443 -929 444 -887
rect 569 -960 570 -928
rect 632 -929 633 -887
rect 639 -960 640 -928
rect 37 -931 38 -887
rect 443 -960 444 -930
rect 457 -960 458 -930
rect 485 -931 486 -887
rect 502 -931 503 -887
rect 681 -960 682 -930
rect 37 -960 38 -932
rect 131 -933 132 -887
rect 142 -960 143 -932
rect 296 -933 297 -887
rect 471 -960 472 -932
rect 583 -960 584 -932
rect 173 -935 174 -887
rect 296 -960 297 -934
rect 478 -935 479 -887
rect 485 -960 486 -934
rect 555 -960 556 -934
rect 695 -935 696 -887
rect 198 -960 199 -936
rect 604 -960 605 -936
rect 695 -960 696 -936
rect 1003 -937 1004 -887
rect 208 -939 209 -887
rect 282 -939 283 -887
rect 478 -960 479 -938
rect 877 -960 878 -938
rect 44 -941 45 -887
rect 282 -960 283 -940
rect 562 -960 563 -940
rect 835 -960 836 -940
rect 44 -960 45 -942
rect 401 -943 402 -887
rect 212 -960 213 -944
rect 222 -945 223 -887
rect 233 -960 234 -944
rect 247 -945 248 -887
rect 268 -960 269 -944
rect 380 -945 381 -887
rect 401 -960 402 -944
rect 656 -960 657 -944
rect 100 -947 101 -887
rect 247 -960 248 -946
rect 79 -949 80 -887
rect 100 -960 101 -948
rect 222 -960 223 -948
rect 345 -960 346 -948
rect 79 -960 80 -950
rect 415 -951 416 -887
rect 415 -960 416 -952
rect 758 -953 759 -887
rect 758 -960 759 -954
rect 772 -955 773 -887
rect 618 -957 619 -887
rect 772 -960 773 -956
rect 618 -960 619 -958
rect 954 -960 955 -958
rect 9 -1053 10 -969
rect 373 -970 374 -968
rect 380 -970 381 -968
rect 548 -970 549 -968
rect 565 -970 566 -968
rect 821 -970 822 -968
rect 835 -970 836 -968
rect 940 -1053 941 -969
rect 947 -970 948 -968
rect 996 -1053 997 -969
rect 1010 -970 1011 -968
rect 1031 -1053 1032 -969
rect 1038 -970 1039 -968
rect 1073 -1053 1074 -969
rect 1087 -970 1088 -968
rect 1094 -1053 1095 -969
rect 16 -972 17 -968
rect 471 -972 472 -968
rect 474 -972 475 -968
rect 1076 -1053 1077 -971
rect 16 -1053 17 -973
rect 366 -974 367 -968
rect 373 -1053 374 -973
rect 401 -974 402 -968
rect 408 -974 409 -968
rect 432 -1053 433 -973
rect 453 -974 454 -968
rect 464 -974 465 -968
rect 481 -974 482 -968
rect 674 -974 675 -968
rect 698 -974 699 -968
rect 870 -974 871 -968
rect 891 -974 892 -968
rect 1045 -1053 1046 -973
rect 1059 -974 1060 -968
rect 1101 -1053 1102 -973
rect 37 -976 38 -968
rect 208 -1053 209 -975
rect 226 -976 227 -968
rect 586 -1053 587 -975
rect 600 -976 601 -968
rect 730 -976 731 -968
rect 751 -976 752 -968
rect 835 -1053 836 -975
rect 842 -976 843 -968
rect 947 -1053 948 -975
rect 954 -976 955 -968
rect 1087 -1053 1088 -975
rect 58 -978 59 -968
rect 474 -1053 475 -977
rect 488 -1053 489 -977
rect 576 -978 577 -968
rect 607 -978 608 -968
rect 800 -978 801 -968
rect 828 -978 829 -968
rect 842 -1053 843 -977
rect 863 -978 864 -968
rect 891 -1053 892 -977
rect 898 -978 899 -968
rect 989 -1053 990 -977
rect 30 -980 31 -968
rect 607 -1053 608 -979
rect 635 -980 636 -968
rect 1010 -1053 1011 -979
rect 30 -1053 31 -981
rect 198 -982 199 -968
rect 240 -982 241 -968
rect 632 -982 633 -968
rect 639 -982 640 -968
rect 674 -1053 675 -981
rect 681 -982 682 -968
rect 751 -1053 752 -981
rect 758 -982 759 -968
rect 912 -1053 913 -981
rect 919 -982 920 -968
rect 968 -982 969 -968
rect 982 -982 983 -968
rect 1069 -1053 1070 -981
rect 61 -1053 62 -983
rect 632 -1053 633 -983
rect 653 -984 654 -968
rect 884 -984 885 -968
rect 905 -984 906 -968
rect 1038 -1053 1039 -983
rect 93 -986 94 -968
rect 243 -986 244 -968
rect 247 -986 248 -968
rect 464 -1053 465 -985
rect 471 -1053 472 -985
rect 954 -1053 955 -985
rect 100 -988 101 -968
rect 327 -988 328 -968
rect 338 -988 339 -968
rect 411 -1053 412 -987
rect 418 -988 419 -968
rect 733 -1053 734 -987
rect 737 -988 738 -968
rect 828 -1053 829 -987
rect 856 -988 857 -968
rect 968 -1053 969 -987
rect 100 -1053 101 -989
rect 219 -1053 220 -989
rect 247 -1053 248 -989
rect 345 -990 346 -968
rect 366 -1053 367 -989
rect 457 -990 458 -968
rect 492 -990 493 -968
rect 688 -990 689 -968
rect 716 -990 717 -968
rect 758 -1053 759 -989
rect 765 -990 766 -968
rect 821 -1053 822 -989
rect 905 -1053 906 -989
rect 915 -990 916 -968
rect 929 -990 930 -968
rect 961 -990 962 -968
rect 93 -1053 94 -991
rect 492 -1053 493 -991
rect 495 -992 496 -968
rect 1017 -1053 1018 -991
rect 114 -994 115 -968
rect 212 -1053 213 -993
rect 261 -994 262 -968
rect 345 -1053 346 -993
rect 380 -1053 381 -993
rect 485 -994 486 -968
rect 506 -994 507 -968
rect 681 -1053 682 -993
rect 730 -1053 731 -993
rect 863 -1053 864 -993
rect 933 -994 934 -968
rect 982 -1053 983 -993
rect 114 -1053 115 -995
rect 149 -996 150 -968
rect 177 -996 178 -968
rect 355 -1053 356 -995
rect 383 -996 384 -968
rect 401 -1053 402 -995
rect 436 -996 437 -968
rect 765 -1053 766 -995
rect 793 -996 794 -968
rect 800 -1053 801 -995
rect 814 -996 815 -968
rect 884 -1053 885 -995
rect 943 -996 944 -968
rect 1059 -1053 1060 -995
rect 121 -998 122 -968
rect 128 -998 129 -968
rect 131 -998 132 -968
rect 975 -1053 976 -997
rect 72 -1000 73 -968
rect 121 -1053 122 -999
rect 131 -1053 132 -999
rect 226 -1053 227 -999
rect 261 -1053 262 -999
rect 422 -1000 423 -968
rect 457 -1053 458 -999
rect 541 -1000 542 -968
rect 548 -1053 549 -999
rect 870 -1053 871 -999
rect 65 -1002 66 -968
rect 422 -1053 423 -1001
rect 506 -1053 507 -1001
rect 649 -1053 650 -1001
rect 660 -1002 661 -968
rect 737 -1053 738 -1001
rect 786 -1002 787 -968
rect 793 -1053 794 -1001
rect 814 -1053 815 -1001
rect 1066 -1053 1067 -1001
rect 65 -1053 66 -1003
rect 156 -1004 157 -968
rect 180 -1004 181 -968
rect 240 -1053 241 -1003
rect 282 -1053 283 -1003
rect 562 -1004 563 -968
rect 576 -1053 577 -1003
rect 1052 -1053 1053 -1003
rect 72 -1053 73 -1005
rect 254 -1006 255 -968
rect 285 -1006 286 -968
rect 779 -1006 780 -968
rect 135 -1008 136 -968
rect 439 -1008 440 -968
rect 450 -1008 451 -968
rect 779 -1053 780 -1007
rect 135 -1053 136 -1009
rect 926 -1010 927 -968
rect 142 -1012 143 -968
rect 530 -1012 531 -968
rect 537 -1053 538 -1011
rect 849 -1012 850 -968
rect 44 -1014 45 -968
rect 142 -1053 143 -1013
rect 145 -1053 146 -1013
rect 1003 -1053 1004 -1013
rect 149 -1053 150 -1015
rect 163 -1016 164 -968
rect 180 -1053 181 -1015
rect 275 -1053 276 -1015
rect 296 -1016 297 -968
rect 436 -1053 437 -1015
rect 450 -1053 451 -1015
rect 926 -1053 927 -1015
rect 23 -1018 24 -968
rect 163 -1053 164 -1017
rect 191 -1018 192 -968
rect 233 -1053 234 -1017
rect 299 -1053 300 -1017
rect 520 -1018 521 -968
rect 527 -1053 528 -1017
rect 667 -1018 668 -968
rect 723 -1018 724 -968
rect 786 -1053 787 -1017
rect 849 -1053 850 -1017
rect 877 -1018 878 -968
rect 23 -1053 24 -1019
rect 222 -1020 223 -968
rect 303 -1020 304 -968
rect 562 -1053 563 -1019
rect 597 -1020 598 -968
rect 919 -1053 920 -1019
rect 40 -1053 41 -1021
rect 191 -1053 192 -1021
rect 198 -1053 199 -1021
rect 205 -1022 206 -968
rect 257 -1053 258 -1021
rect 597 -1053 598 -1021
rect 604 -1022 605 -968
rect 898 -1053 899 -1021
rect 51 -1024 52 -968
rect 296 -1053 297 -1023
rect 303 -1053 304 -1023
rect 429 -1024 430 -968
rect 443 -1024 444 -968
rect 667 -1053 668 -1023
rect 702 -1024 703 -968
rect 723 -1053 724 -1023
rect 807 -1024 808 -968
rect 877 -1053 878 -1023
rect 51 -1053 52 -1025
rect 86 -1026 87 -968
rect 156 -1053 157 -1025
rect 205 -1053 206 -1025
rect 310 -1026 311 -968
rect 478 -1026 479 -968
rect 499 -1026 500 -968
rect 520 -1053 521 -1025
rect 541 -1053 542 -1025
rect 590 -1026 591 -968
rect 604 -1053 605 -1025
rect 933 -1053 934 -1025
rect 44 -1053 45 -1027
rect 478 -1053 479 -1027
rect 499 -1053 500 -1027
rect 922 -1028 923 -968
rect 79 -1030 80 -968
rect 310 -1053 311 -1029
rect 317 -1030 318 -968
rect 338 -1053 339 -1029
rect 387 -1030 388 -968
rect 394 -1053 395 -1029
rect 397 -1030 398 -968
rect 415 -1053 416 -1029
rect 443 -1053 444 -1029
rect 744 -1030 745 -968
rect 79 -1053 80 -1031
rect 359 -1032 360 -968
rect 516 -1053 517 -1031
rect 772 -1032 773 -968
rect 268 -1034 269 -968
rect 317 -1053 318 -1033
rect 324 -1034 325 -968
rect 387 -1053 388 -1033
rect 429 -1053 430 -1033
rect 772 -1053 773 -1033
rect 107 -1036 108 -968
rect 268 -1053 269 -1035
rect 331 -1036 332 -968
rect 359 -1053 360 -1035
rect 534 -1036 535 -968
rect 590 -1053 591 -1035
rect 611 -1036 612 -968
rect 653 -1053 654 -1035
rect 702 -1053 703 -1035
rect 709 -1036 710 -968
rect 107 -1053 108 -1037
rect 170 -1038 171 -968
rect 184 -1038 185 -968
rect 324 -1053 325 -1037
rect 331 -1053 332 -1037
rect 352 -1038 353 -968
rect 551 -1053 552 -1037
rect 856 -1053 857 -1037
rect 12 -1040 13 -968
rect 352 -1053 353 -1039
rect 555 -1040 556 -968
rect 639 -1053 640 -1039
rect 646 -1040 647 -968
rect 660 -1053 661 -1039
rect 691 -1053 692 -1039
rect 709 -1053 710 -1039
rect 184 -1053 185 -1041
rect 289 -1042 290 -968
rect 453 -1053 454 -1041
rect 555 -1053 556 -1041
rect 569 -1042 570 -968
rect 611 -1053 612 -1041
rect 618 -1042 619 -968
rect 716 -1053 717 -1041
rect 289 -1053 290 -1043
rect 362 -1044 363 -968
rect 446 -1053 447 -1043
rect 618 -1053 619 -1043
rect 625 -1044 626 -968
rect 961 -1053 962 -1043
rect 569 -1053 570 -1045
rect 695 -1046 696 -968
rect 583 -1048 584 -968
rect 744 -1053 745 -1047
rect 86 -1053 87 -1049
rect 583 -1053 584 -1049
rect 628 -1053 629 -1049
rect 807 -1053 808 -1049
rect 646 -1053 647 -1051
rect 695 -1053 696 -1051
rect 16 -1063 17 -1061
rect 450 -1152 451 -1062
rect 478 -1063 479 -1061
rect 828 -1063 829 -1061
rect 961 -1063 962 -1061
rect 1024 -1152 1025 -1062
rect 1027 -1063 1028 -1061
rect 1052 -1063 1053 -1061
rect 1059 -1063 1060 -1061
rect 1083 -1063 1084 -1061
rect 1094 -1063 1095 -1061
rect 1097 -1063 1098 -1061
rect 19 -1152 20 -1064
rect 334 -1152 335 -1064
rect 338 -1065 339 -1061
rect 443 -1065 444 -1061
rect 464 -1065 465 -1061
rect 478 -1152 479 -1064
rect 495 -1065 496 -1061
rect 877 -1065 878 -1061
rect 989 -1065 990 -1061
rect 1059 -1152 1060 -1064
rect 1094 -1152 1095 -1064
rect 1101 -1065 1102 -1061
rect 30 -1067 31 -1061
rect 37 -1152 38 -1066
rect 51 -1067 52 -1061
rect 58 -1067 59 -1061
rect 65 -1067 66 -1061
rect 145 -1152 146 -1066
rect 156 -1067 157 -1061
rect 180 -1067 181 -1061
rect 191 -1067 192 -1061
rect 194 -1079 195 -1066
rect 205 -1067 206 -1061
rect 205 -1152 206 -1066
rect 205 -1067 206 -1061
rect 205 -1152 206 -1066
rect 219 -1152 220 -1066
rect 229 -1152 230 -1066
rect 275 -1067 276 -1061
rect 548 -1152 549 -1066
rect 569 -1067 570 -1061
rect 898 -1067 899 -1061
rect 996 -1067 997 -1061
rect 1052 -1152 1053 -1066
rect 51 -1152 52 -1068
rect 131 -1152 132 -1068
rect 142 -1069 143 -1061
rect 264 -1152 265 -1068
rect 282 -1069 283 -1061
rect 474 -1152 475 -1068
rect 513 -1069 514 -1061
rect 576 -1069 577 -1061
rect 579 -1069 580 -1061
rect 870 -1069 871 -1061
rect 1017 -1069 1018 -1061
rect 1073 -1152 1074 -1068
rect 58 -1152 59 -1070
rect 355 -1071 356 -1061
rect 369 -1152 370 -1070
rect 933 -1071 934 -1061
rect 65 -1152 66 -1072
rect 261 -1073 262 -1061
rect 296 -1152 297 -1072
rect 373 -1073 374 -1061
rect 387 -1073 388 -1061
rect 513 -1152 514 -1072
rect 576 -1152 577 -1072
rect 600 -1152 601 -1072
rect 604 -1152 605 -1072
rect 828 -1152 829 -1072
rect 926 -1073 927 -1061
rect 1017 -1152 1018 -1072
rect 2 -1152 3 -1074
rect 261 -1152 262 -1074
rect 303 -1075 304 -1061
rect 467 -1152 468 -1074
rect 583 -1075 584 -1061
rect 1045 -1075 1046 -1061
rect 79 -1077 80 -1061
rect 187 -1152 188 -1076
rect 191 -1152 192 -1076
rect 222 -1077 223 -1061
rect 345 -1077 346 -1061
rect 352 -1077 353 -1061
rect 940 -1077 941 -1061
rect 86 -1079 87 -1061
rect 86 -1152 87 -1078
rect 86 -1079 87 -1061
rect 86 -1152 87 -1078
rect 114 -1079 115 -1061
rect 173 -1079 174 -1061
rect 177 -1152 178 -1078
rect 198 -1079 199 -1061
rect 233 -1079 234 -1061
rect 275 -1152 276 -1078
rect 310 -1079 311 -1061
rect 495 -1152 496 -1078
rect 569 -1152 570 -1078
rect 583 -1152 584 -1078
rect 586 -1152 587 -1078
rect 912 -1079 913 -1061
rect 940 -1152 941 -1078
rect 1087 -1079 1088 -1061
rect 1097 -1152 1098 -1078
rect 1101 -1152 1102 -1078
rect 93 -1081 94 -1061
rect 114 -1152 115 -1080
rect 121 -1081 122 -1061
rect 254 -1152 255 -1080
rect 317 -1081 318 -1061
rect 443 -1152 444 -1080
rect 572 -1081 573 -1061
rect 1045 -1152 1046 -1080
rect 44 -1083 45 -1061
rect 121 -1152 122 -1082
rect 156 -1152 157 -1082
rect 289 -1083 290 -1061
rect 324 -1083 325 -1061
rect 453 -1083 454 -1061
rect 593 -1152 594 -1082
rect 954 -1083 955 -1061
rect 44 -1152 45 -1084
rect 537 -1085 538 -1061
rect 597 -1085 598 -1061
rect 607 -1152 608 -1084
rect 621 -1152 622 -1084
rect 996 -1152 997 -1084
rect 93 -1152 94 -1086
rect 243 -1152 244 -1086
rect 247 -1087 248 -1061
rect 282 -1152 283 -1086
rect 289 -1152 290 -1086
rect 331 -1087 332 -1061
rect 338 -1152 339 -1086
rect 436 -1087 437 -1061
rect 439 -1152 440 -1086
rect 541 -1087 542 -1061
rect 628 -1087 629 -1061
rect 835 -1087 836 -1061
rect 863 -1087 864 -1061
rect 926 -1152 927 -1086
rect 135 -1089 136 -1061
rect 324 -1152 325 -1088
rect 345 -1152 346 -1088
rect 590 -1089 591 -1061
rect 628 -1152 629 -1088
rect 947 -1089 948 -1061
rect 107 -1091 108 -1061
rect 135 -1152 136 -1090
rect 163 -1152 164 -1090
rect 492 -1091 493 -1061
rect 509 -1152 510 -1090
rect 947 -1152 948 -1090
rect 107 -1152 108 -1092
rect 170 -1093 171 -1061
rect 184 -1093 185 -1061
rect 317 -1152 318 -1092
rect 359 -1093 360 -1061
rect 373 -1152 374 -1092
rect 387 -1152 388 -1092
rect 401 -1093 402 -1061
rect 408 -1093 409 -1061
rect 863 -1152 864 -1092
rect 912 -1152 913 -1092
rect 982 -1093 983 -1061
rect 100 -1095 101 -1061
rect 170 -1152 171 -1094
rect 198 -1152 199 -1094
rect 380 -1095 381 -1061
rect 394 -1095 395 -1061
rect 408 -1152 409 -1094
rect 411 -1095 412 -1061
rect 446 -1095 447 -1061
rect 541 -1152 542 -1094
rect 1069 -1095 1070 -1061
rect 9 -1097 10 -1061
rect 100 -1152 101 -1096
rect 166 -1097 167 -1061
rect 961 -1152 962 -1096
rect 240 -1099 241 -1061
rect 310 -1152 311 -1098
rect 359 -1152 360 -1098
rect 446 -1152 447 -1098
rect 590 -1152 591 -1098
rect 884 -1099 885 -1061
rect 919 -1099 920 -1061
rect 954 -1152 955 -1098
rect 247 -1152 248 -1100
rect 597 -1152 598 -1100
rect 646 -1101 647 -1061
rect 677 -1152 678 -1100
rect 688 -1101 689 -1061
rect 905 -1101 906 -1061
rect 919 -1152 920 -1100
rect 1080 -1101 1081 -1061
rect 380 -1152 381 -1102
rect 506 -1103 507 -1061
rect 649 -1103 650 -1061
rect 968 -1103 969 -1061
rect 1003 -1103 1004 -1061
rect 1080 -1152 1081 -1102
rect 72 -1105 73 -1061
rect 506 -1152 507 -1104
rect 688 -1152 689 -1104
rect 982 -1152 983 -1104
rect 23 -1107 24 -1061
rect 72 -1152 73 -1106
rect 394 -1152 395 -1106
rect 562 -1107 563 -1061
rect 723 -1107 724 -1061
rect 835 -1152 836 -1106
rect 849 -1107 850 -1061
rect 968 -1152 969 -1106
rect 23 -1152 24 -1108
rect 128 -1152 129 -1108
rect 401 -1152 402 -1108
rect 534 -1109 535 -1061
rect 555 -1109 556 -1061
rect 562 -1152 563 -1108
rect 639 -1109 640 -1061
rect 723 -1152 724 -1108
rect 726 -1152 727 -1108
rect 898 -1152 899 -1108
rect 422 -1111 423 -1061
rect 551 -1111 552 -1061
rect 555 -1152 556 -1110
rect 611 -1111 612 -1061
rect 730 -1111 731 -1061
rect 989 -1152 990 -1110
rect 268 -1113 269 -1061
rect 422 -1152 423 -1112
rect 429 -1113 430 -1061
rect 667 -1113 668 -1061
rect 730 -1152 731 -1112
rect 1038 -1113 1039 -1061
rect 429 -1152 430 -1114
rect 527 -1115 528 -1061
rect 611 -1152 612 -1114
rect 632 -1115 633 -1061
rect 667 -1152 668 -1114
rect 751 -1115 752 -1061
rect 765 -1115 766 -1061
rect 849 -1152 850 -1114
rect 856 -1115 857 -1061
rect 905 -1152 906 -1114
rect 1038 -1152 1039 -1114
rect 1076 -1115 1077 -1061
rect 436 -1152 437 -1116
rect 1066 -1152 1067 -1116
rect 457 -1119 458 -1061
rect 646 -1152 647 -1118
rect 779 -1119 780 -1061
rect 870 -1152 871 -1118
rect 457 -1152 458 -1120
rect 499 -1121 500 -1061
rect 520 -1121 521 -1061
rect 534 -1152 535 -1120
rect 618 -1121 619 -1061
rect 751 -1152 752 -1120
rect 786 -1121 787 -1061
rect 1003 -1152 1004 -1120
rect 226 -1123 227 -1061
rect 499 -1152 500 -1122
rect 520 -1152 521 -1122
rect 660 -1123 661 -1061
rect 716 -1123 717 -1061
rect 779 -1152 780 -1122
rect 800 -1123 801 -1061
rect 884 -1152 885 -1122
rect 226 -1152 227 -1124
rect 268 -1152 269 -1124
rect 530 -1152 531 -1124
rect 765 -1152 766 -1124
rect 800 -1152 801 -1124
rect 814 -1125 815 -1061
rect 821 -1125 822 -1061
rect 877 -1152 878 -1124
rect 632 -1152 633 -1126
rect 737 -1127 738 -1061
rect 758 -1127 759 -1061
rect 821 -1152 822 -1126
rect 653 -1129 654 -1061
rect 786 -1152 787 -1128
rect 807 -1129 808 -1061
rect 856 -1152 857 -1128
rect 653 -1152 654 -1130
rect 744 -1131 745 -1061
rect 772 -1131 773 -1061
rect 814 -1152 815 -1130
rect 240 -1152 241 -1132
rect 744 -1152 745 -1132
rect 807 -1152 808 -1132
rect 891 -1133 892 -1061
rect 660 -1152 661 -1134
rect 1010 -1135 1011 -1061
rect 681 -1137 682 -1061
rect 716 -1152 717 -1136
rect 793 -1137 794 -1061
rect 891 -1152 892 -1136
rect 1010 -1152 1011 -1136
rect 1031 -1137 1032 -1061
rect 299 -1139 300 -1061
rect 681 -1152 682 -1138
rect 695 -1139 696 -1061
rect 737 -1152 738 -1138
rect 842 -1139 843 -1061
rect 1031 -1152 1032 -1138
rect 492 -1152 493 -1140
rect 793 -1152 794 -1140
rect 842 -1152 843 -1140
rect 975 -1141 976 -1061
rect 485 -1143 486 -1061
rect 975 -1152 976 -1142
rect 366 -1145 367 -1061
rect 485 -1152 486 -1144
rect 674 -1145 675 -1061
rect 695 -1152 696 -1144
rect 702 -1145 703 -1061
rect 772 -1152 773 -1144
rect 366 -1152 367 -1146
rect 415 -1147 416 -1061
rect 642 -1152 643 -1146
rect 702 -1152 703 -1146
rect 709 -1147 710 -1061
rect 758 -1152 759 -1146
rect 149 -1149 150 -1061
rect 415 -1152 416 -1148
rect 674 -1152 675 -1148
rect 933 -1152 934 -1148
rect 149 -1152 150 -1150
rect 236 -1152 237 -1150
rect 709 -1152 710 -1150
rect 1087 -1152 1088 -1150
rect 30 -1162 31 -1160
rect 586 -1162 587 -1160
rect 590 -1162 591 -1160
rect 621 -1162 622 -1160
rect 639 -1162 640 -1160
rect 891 -1162 892 -1160
rect 1090 -1162 1091 -1160
rect 1101 -1162 1102 -1160
rect 30 -1255 31 -1163
rect 149 -1164 150 -1160
rect 156 -1164 157 -1160
rect 236 -1164 237 -1160
rect 243 -1164 244 -1160
rect 310 -1164 311 -1160
rect 331 -1164 332 -1160
rect 919 -1164 920 -1160
rect 33 -1166 34 -1160
rect 93 -1166 94 -1160
rect 121 -1166 122 -1160
rect 149 -1255 150 -1165
rect 156 -1255 157 -1165
rect 366 -1166 367 -1160
rect 429 -1166 430 -1160
rect 460 -1255 461 -1165
rect 464 -1166 465 -1160
rect 1080 -1166 1081 -1160
rect 51 -1168 52 -1160
rect 366 -1255 367 -1167
rect 436 -1168 437 -1160
rect 1041 -1255 1042 -1167
rect 58 -1170 59 -1160
rect 82 -1170 83 -1160
rect 93 -1255 94 -1169
rect 163 -1170 164 -1160
rect 194 -1255 195 -1169
rect 240 -1170 241 -1160
rect 247 -1170 248 -1160
rect 464 -1255 465 -1169
rect 471 -1170 472 -1160
rect 1024 -1170 1025 -1160
rect 58 -1255 59 -1171
rect 86 -1172 87 -1160
rect 114 -1172 115 -1160
rect 121 -1255 122 -1171
rect 128 -1172 129 -1160
rect 387 -1172 388 -1160
rect 439 -1172 440 -1160
rect 478 -1172 479 -1160
rect 495 -1172 496 -1160
rect 849 -1172 850 -1160
rect 891 -1255 892 -1171
rect 996 -1172 997 -1160
rect 51 -1255 52 -1173
rect 86 -1255 87 -1173
rect 114 -1255 115 -1173
rect 681 -1174 682 -1160
rect 684 -1255 685 -1173
rect 1003 -1174 1004 -1160
rect 65 -1176 66 -1160
rect 65 -1255 66 -1175
rect 65 -1176 66 -1160
rect 65 -1255 66 -1175
rect 82 -1255 83 -1175
rect 100 -1176 101 -1160
rect 128 -1255 129 -1175
rect 135 -1176 136 -1160
rect 163 -1255 164 -1175
rect 954 -1176 955 -1160
rect 135 -1255 136 -1177
rect 212 -1178 213 -1160
rect 226 -1178 227 -1160
rect 625 -1178 626 -1160
rect 639 -1255 640 -1177
rect 772 -1178 773 -1160
rect 842 -1178 843 -1160
rect 1003 -1255 1004 -1177
rect 117 -1255 118 -1179
rect 625 -1255 626 -1179
rect 642 -1180 643 -1160
rect 737 -1180 738 -1160
rect 772 -1255 773 -1179
rect 828 -1180 829 -1160
rect 842 -1255 843 -1179
rect 1087 -1180 1088 -1160
rect 170 -1182 171 -1160
rect 240 -1255 241 -1181
rect 247 -1255 248 -1181
rect 394 -1182 395 -1160
rect 446 -1182 447 -1160
rect 534 -1182 535 -1160
rect 544 -1255 545 -1181
rect 800 -1182 801 -1160
rect 919 -1255 920 -1181
rect 989 -1182 990 -1160
rect 184 -1184 185 -1160
rect 989 -1255 990 -1183
rect 37 -1186 38 -1160
rect 184 -1255 185 -1185
rect 198 -1186 199 -1160
rect 478 -1255 479 -1185
rect 495 -1255 496 -1185
rect 786 -1186 787 -1160
rect 954 -1255 955 -1185
rect 1066 -1186 1067 -1160
rect 37 -1255 38 -1187
rect 166 -1255 167 -1187
rect 226 -1255 227 -1187
rect 317 -1188 318 -1160
rect 331 -1255 332 -1187
rect 345 -1188 346 -1160
rect 352 -1255 353 -1187
rect 373 -1188 374 -1160
rect 380 -1188 381 -1160
rect 436 -1255 437 -1187
rect 450 -1188 451 -1160
rect 527 -1255 528 -1187
rect 548 -1188 549 -1160
rect 551 -1255 552 -1187
rect 590 -1255 591 -1187
rect 996 -1255 997 -1187
rect 79 -1190 80 -1160
rect 345 -1255 346 -1189
rect 380 -1255 381 -1189
rect 401 -1190 402 -1160
rect 450 -1255 451 -1189
rect 485 -1190 486 -1160
rect 509 -1190 510 -1160
rect 1017 -1190 1018 -1160
rect 79 -1255 80 -1191
rect 506 -1255 507 -1191
rect 513 -1192 514 -1160
rect 583 -1192 584 -1160
rect 597 -1192 598 -1160
rect 1031 -1192 1032 -1160
rect 44 -1194 45 -1160
rect 513 -1255 514 -1193
rect 516 -1255 517 -1193
rect 849 -1255 850 -1193
rect 1010 -1194 1011 -1160
rect 1017 -1255 1018 -1193
rect 44 -1255 45 -1195
rect 170 -1255 171 -1195
rect 229 -1196 230 -1160
rect 275 -1196 276 -1160
rect 282 -1196 283 -1160
rect 565 -1255 566 -1195
rect 600 -1196 601 -1160
rect 940 -1196 941 -1160
rect 72 -1198 73 -1160
rect 597 -1255 598 -1197
rect 604 -1198 605 -1160
rect 716 -1198 717 -1160
rect 723 -1198 724 -1160
rect 1052 -1198 1053 -1160
rect 26 -1255 27 -1199
rect 604 -1255 605 -1199
rect 611 -1200 612 -1160
rect 611 -1255 612 -1199
rect 611 -1200 612 -1160
rect 611 -1255 612 -1199
rect 618 -1200 619 -1160
rect 646 -1200 647 -1160
rect 660 -1200 661 -1160
rect 828 -1255 829 -1199
rect 835 -1200 836 -1160
rect 1052 -1255 1053 -1199
rect 72 -1255 73 -1201
rect 324 -1202 325 -1160
rect 387 -1255 388 -1201
rect 569 -1202 570 -1160
rect 618 -1255 619 -1201
rect 628 -1202 629 -1160
rect 660 -1255 661 -1201
rect 695 -1202 696 -1160
rect 716 -1255 717 -1201
rect 884 -1202 885 -1160
rect 912 -1202 913 -1160
rect 1010 -1255 1011 -1201
rect 107 -1204 108 -1160
rect 324 -1255 325 -1203
rect 394 -1255 395 -1203
rect 415 -1204 416 -1160
rect 485 -1255 486 -1203
rect 709 -1204 710 -1160
rect 723 -1255 724 -1203
rect 814 -1204 815 -1160
rect 884 -1255 885 -1203
rect 982 -1204 983 -1160
rect 107 -1255 108 -1205
rect 198 -1255 199 -1205
rect 233 -1206 234 -1160
rect 306 -1206 307 -1160
rect 310 -1255 311 -1205
rect 541 -1206 542 -1160
rect 555 -1206 556 -1160
rect 646 -1255 647 -1205
rect 667 -1206 668 -1160
rect 688 -1255 689 -1205
rect 691 -1206 692 -1160
rect 1024 -1255 1025 -1205
rect 219 -1208 220 -1160
rect 233 -1255 234 -1207
rect 254 -1208 255 -1160
rect 317 -1255 318 -1207
rect 401 -1255 402 -1207
rect 408 -1208 409 -1160
rect 492 -1255 493 -1207
rect 667 -1255 668 -1207
rect 677 -1208 678 -1160
rect 1045 -1208 1046 -1160
rect 16 -1255 17 -1209
rect 254 -1255 255 -1209
rect 261 -1255 262 -1209
rect 548 -1255 549 -1209
rect 555 -1255 556 -1209
rect 576 -1210 577 -1160
rect 586 -1255 587 -1209
rect 912 -1255 913 -1209
rect 1045 -1255 1046 -1209
rect 1073 -1210 1074 -1160
rect 177 -1212 178 -1160
rect 219 -1255 220 -1211
rect 264 -1212 265 -1160
rect 674 -1255 675 -1211
rect 695 -1255 696 -1211
rect 765 -1212 766 -1160
rect 814 -1255 815 -1211
rect 1038 -1212 1039 -1160
rect 1073 -1255 1074 -1211
rect 1094 -1212 1095 -1160
rect 177 -1255 178 -1213
rect 523 -1255 524 -1213
rect 541 -1255 542 -1213
rect 1031 -1255 1032 -1213
rect 1038 -1255 1039 -1213
rect 1066 -1255 1067 -1213
rect 268 -1216 269 -1160
rect 415 -1255 416 -1215
rect 502 -1255 503 -1215
rect 835 -1255 836 -1215
rect 856 -1216 857 -1160
rect 982 -1255 983 -1215
rect 268 -1255 269 -1217
rect 471 -1255 472 -1217
rect 520 -1218 521 -1160
rect 530 -1218 531 -1160
rect 562 -1218 563 -1160
rect 576 -1255 577 -1217
rect 653 -1218 654 -1160
rect 765 -1255 766 -1217
rect 807 -1218 808 -1160
rect 856 -1255 857 -1217
rect 275 -1255 276 -1219
rect 359 -1220 360 -1160
rect 408 -1255 409 -1219
rect 474 -1220 475 -1160
rect 562 -1255 563 -1219
rect 821 -1220 822 -1160
rect 282 -1255 283 -1221
rect 656 -1255 657 -1221
rect 709 -1255 710 -1221
rect 719 -1255 720 -1221
rect 730 -1255 731 -1221
rect 877 -1222 878 -1160
rect 142 -1224 143 -1160
rect 877 -1255 878 -1223
rect 2 -1226 3 -1160
rect 142 -1255 143 -1225
rect 289 -1226 290 -1160
rect 429 -1255 430 -1225
rect 457 -1226 458 -1160
rect 474 -1255 475 -1225
rect 569 -1255 570 -1225
rect 779 -1226 780 -1160
rect 807 -1255 808 -1225
rect 905 -1226 906 -1160
rect 2 -1255 3 -1227
rect 205 -1228 206 -1160
rect 292 -1255 293 -1227
rect 733 -1228 734 -1160
rect 737 -1255 738 -1227
rect 744 -1228 745 -1160
rect 758 -1228 759 -1160
rect 800 -1255 801 -1227
rect 821 -1255 822 -1227
rect 870 -1228 871 -1160
rect 9 -1230 10 -1160
rect 289 -1255 290 -1229
rect 296 -1230 297 -1160
rect 373 -1255 374 -1229
rect 663 -1230 664 -1160
rect 905 -1255 906 -1229
rect 9 -1255 10 -1231
rect 215 -1255 216 -1231
rect 296 -1255 297 -1231
rect 499 -1232 500 -1160
rect 702 -1232 703 -1160
rect 744 -1255 745 -1231
rect 751 -1232 752 -1160
rect 758 -1255 759 -1231
rect 779 -1255 780 -1231
rect 940 -1255 941 -1231
rect 23 -1234 24 -1160
rect 457 -1255 458 -1233
rect 499 -1255 500 -1233
rect 632 -1234 633 -1160
rect 681 -1255 682 -1233
rect 702 -1255 703 -1233
rect 751 -1255 752 -1233
rect 782 -1255 783 -1233
rect 870 -1255 871 -1233
rect 947 -1234 948 -1160
rect 23 -1255 24 -1235
rect 933 -1236 934 -1160
rect 947 -1255 948 -1235
rect 975 -1236 976 -1160
rect 191 -1238 192 -1160
rect 205 -1255 206 -1237
rect 303 -1255 304 -1237
rect 467 -1238 468 -1160
rect 933 -1255 934 -1237
rect 1059 -1238 1060 -1160
rect 100 -1255 101 -1239
rect 191 -1255 192 -1239
rect 338 -1240 339 -1160
rect 359 -1255 360 -1239
rect 422 -1240 423 -1160
rect 632 -1255 633 -1239
rect 793 -1240 794 -1160
rect 1059 -1255 1060 -1239
rect 338 -1255 339 -1241
rect 593 -1242 594 -1160
rect 961 -1242 962 -1160
rect 975 -1255 976 -1241
rect 355 -1244 356 -1160
rect 422 -1255 423 -1243
rect 443 -1244 444 -1160
rect 793 -1255 794 -1243
rect 961 -1255 962 -1243
rect 968 -1244 969 -1160
rect 443 -1255 444 -1245
rect 607 -1255 608 -1245
rect 898 -1246 899 -1160
rect 968 -1255 969 -1245
rect 863 -1248 864 -1160
rect 898 -1255 899 -1247
rect 863 -1255 864 -1249
rect 926 -1250 927 -1160
rect 187 -1252 188 -1160
rect 926 -1255 927 -1251
rect 187 -1255 188 -1253
rect 786 -1255 787 -1253
rect 2 -1265 3 -1263
rect 516 -1265 517 -1263
rect 520 -1265 521 -1263
rect 800 -1265 801 -1263
rect 814 -1334 815 -1264
rect 842 -1265 843 -1263
rect 863 -1265 864 -1263
rect 863 -1334 864 -1264
rect 863 -1265 864 -1263
rect 863 -1334 864 -1264
rect 870 -1265 871 -1263
rect 873 -1271 874 -1264
rect 898 -1265 899 -1263
rect 898 -1334 899 -1264
rect 898 -1265 899 -1263
rect 898 -1334 899 -1264
rect 982 -1265 983 -1263
rect 1062 -1334 1063 -1264
rect 1066 -1265 1067 -1263
rect 1080 -1334 1081 -1264
rect 9 -1267 10 -1263
rect 16 -1334 17 -1266
rect 30 -1267 31 -1263
rect 166 -1267 167 -1263
rect 170 -1267 171 -1263
rect 240 -1267 241 -1263
rect 254 -1267 255 -1263
rect 502 -1267 503 -1263
rect 513 -1267 514 -1263
rect 821 -1267 822 -1263
rect 870 -1334 871 -1266
rect 947 -1267 948 -1263
rect 982 -1334 983 -1266
rect 1017 -1267 1018 -1263
rect 1020 -1267 1021 -1263
rect 1045 -1267 1046 -1263
rect 1045 -1334 1046 -1266
rect 1045 -1267 1046 -1263
rect 1045 -1334 1046 -1266
rect 1073 -1267 1074 -1263
rect 1073 -1334 1074 -1266
rect 1073 -1267 1074 -1263
rect 1073 -1334 1074 -1266
rect 9 -1334 10 -1268
rect 58 -1269 59 -1263
rect 86 -1269 87 -1263
rect 590 -1334 591 -1268
rect 604 -1269 605 -1263
rect 779 -1334 780 -1268
rect 912 -1269 913 -1263
rect 947 -1334 948 -1268
rect 1017 -1334 1018 -1268
rect 1052 -1269 1053 -1263
rect 30 -1334 31 -1270
rect 86 -1334 87 -1270
rect 93 -1271 94 -1263
rect 215 -1271 216 -1263
rect 219 -1271 220 -1263
rect 233 -1271 234 -1263
rect 240 -1334 241 -1270
rect 261 -1271 262 -1263
rect 317 -1271 318 -1263
rect 327 -1334 328 -1270
rect 331 -1271 332 -1263
rect 460 -1334 461 -1270
rect 464 -1271 465 -1263
rect 520 -1334 521 -1270
rect 541 -1271 542 -1263
rect 1003 -1271 1004 -1263
rect 1020 -1334 1021 -1270
rect 1052 -1334 1053 -1270
rect 51 -1273 52 -1263
rect 296 -1273 297 -1263
rect 320 -1334 321 -1272
rect 478 -1273 479 -1263
rect 548 -1273 549 -1263
rect 730 -1273 731 -1263
rect 744 -1273 745 -1263
rect 744 -1334 745 -1272
rect 744 -1273 745 -1263
rect 744 -1334 745 -1272
rect 751 -1273 752 -1263
rect 1066 -1334 1067 -1272
rect 51 -1334 52 -1274
rect 149 -1275 150 -1263
rect 159 -1334 160 -1274
rect 471 -1275 472 -1263
rect 478 -1334 479 -1274
rect 695 -1275 696 -1263
rect 761 -1334 762 -1274
rect 821 -1334 822 -1274
rect 884 -1275 885 -1263
rect 912 -1334 913 -1274
rect 1003 -1334 1004 -1274
rect 1034 -1334 1035 -1274
rect 54 -1277 55 -1263
rect 310 -1277 311 -1263
rect 366 -1277 367 -1263
rect 495 -1277 496 -1263
rect 576 -1277 577 -1263
rect 583 -1277 584 -1263
rect 586 -1277 587 -1263
rect 688 -1277 689 -1263
rect 884 -1334 885 -1276
rect 891 -1277 892 -1263
rect 58 -1334 59 -1278
rect 282 -1279 283 -1263
rect 292 -1279 293 -1263
rect 730 -1334 731 -1278
rect 835 -1279 836 -1263
rect 891 -1334 892 -1278
rect 65 -1281 66 -1263
rect 149 -1334 150 -1280
rect 170 -1334 171 -1280
rect 674 -1281 675 -1263
rect 677 -1334 678 -1280
rect 1010 -1281 1011 -1263
rect 65 -1334 66 -1282
rect 338 -1283 339 -1263
rect 369 -1334 370 -1282
rect 527 -1283 528 -1263
rect 555 -1283 556 -1263
rect 576 -1334 577 -1282
rect 583 -1334 584 -1282
rect 632 -1283 633 -1263
rect 639 -1283 640 -1263
rect 695 -1334 696 -1282
rect 817 -1283 818 -1263
rect 835 -1334 836 -1282
rect 954 -1283 955 -1263
rect 1010 -1334 1011 -1282
rect 93 -1334 94 -1284
rect 100 -1285 101 -1263
rect 114 -1285 115 -1263
rect 131 -1334 132 -1284
rect 135 -1285 136 -1263
rect 317 -1334 318 -1284
rect 331 -1334 332 -1284
rect 366 -1334 367 -1284
rect 422 -1285 423 -1263
rect 548 -1334 549 -1284
rect 565 -1285 566 -1263
rect 639 -1334 640 -1284
rect 653 -1285 654 -1263
rect 961 -1285 962 -1263
rect 100 -1334 101 -1286
rect 121 -1287 122 -1263
rect 142 -1287 143 -1263
rect 289 -1287 290 -1263
rect 292 -1334 293 -1286
rect 324 -1287 325 -1263
rect 338 -1334 339 -1286
rect 352 -1287 353 -1263
rect 425 -1287 426 -1263
rect 436 -1287 437 -1263
rect 443 -1287 444 -1263
rect 541 -1334 542 -1286
rect 604 -1334 605 -1286
rect 611 -1287 612 -1263
rect 625 -1287 626 -1263
rect 632 -1334 633 -1286
rect 653 -1334 654 -1286
rect 1059 -1287 1060 -1263
rect 23 -1289 24 -1263
rect 121 -1334 122 -1288
rect 142 -1334 143 -1288
rect 226 -1289 227 -1263
rect 261 -1334 262 -1288
rect 275 -1289 276 -1263
rect 282 -1334 283 -1288
rect 359 -1289 360 -1263
rect 415 -1289 416 -1263
rect 436 -1334 437 -1288
rect 443 -1334 444 -1288
rect 474 -1334 475 -1288
rect 527 -1334 528 -1288
rect 534 -1334 535 -1288
rect 537 -1289 538 -1263
rect 555 -1334 556 -1288
rect 607 -1289 608 -1263
rect 856 -1289 857 -1263
rect 940 -1289 941 -1263
rect 961 -1334 962 -1288
rect 23 -1334 24 -1290
rect 107 -1291 108 -1263
rect 117 -1291 118 -1263
rect 737 -1291 738 -1263
rect 751 -1334 752 -1290
rect 1059 -1334 1060 -1290
rect 72 -1293 73 -1263
rect 352 -1334 353 -1292
rect 359 -1334 360 -1292
rect 765 -1293 766 -1263
rect 793 -1293 794 -1263
rect 856 -1334 857 -1292
rect 919 -1293 920 -1263
rect 940 -1334 941 -1292
rect 72 -1334 73 -1294
rect 387 -1295 388 -1263
rect 464 -1334 465 -1294
rect 506 -1295 507 -1263
rect 537 -1334 538 -1294
rect 646 -1295 647 -1263
rect 656 -1295 657 -1263
rect 989 -1295 990 -1263
rect 107 -1334 108 -1296
rect 138 -1334 139 -1296
rect 163 -1297 164 -1263
rect 625 -1334 626 -1296
rect 660 -1297 661 -1263
rect 842 -1334 843 -1296
rect 849 -1297 850 -1263
rect 919 -1334 920 -1296
rect 968 -1297 969 -1263
rect 989 -1334 990 -1296
rect 117 -1334 118 -1298
rect 310 -1334 311 -1298
rect 373 -1299 374 -1263
rect 387 -1334 388 -1298
rect 611 -1334 612 -1298
rect 618 -1299 619 -1263
rect 660 -1334 661 -1298
rect 702 -1299 703 -1263
rect 716 -1299 717 -1263
rect 765 -1334 766 -1298
rect 793 -1334 794 -1298
rect 1038 -1334 1039 -1298
rect 128 -1301 129 -1263
rect 163 -1334 164 -1300
rect 173 -1334 174 -1300
rect 1024 -1301 1025 -1263
rect 187 -1303 188 -1263
rect 996 -1303 997 -1263
rect 191 -1334 192 -1304
rect 975 -1305 976 -1263
rect 996 -1334 997 -1304
rect 1031 -1334 1032 -1304
rect 194 -1307 195 -1263
rect 247 -1307 248 -1263
rect 268 -1307 269 -1263
rect 646 -1334 647 -1306
rect 667 -1307 668 -1263
rect 800 -1334 801 -1306
rect 807 -1307 808 -1263
rect 954 -1334 955 -1306
rect 194 -1334 195 -1308
rect 254 -1334 255 -1308
rect 268 -1334 269 -1308
rect 345 -1309 346 -1263
rect 373 -1334 374 -1308
rect 485 -1309 486 -1263
rect 667 -1334 668 -1308
rect 1041 -1309 1042 -1263
rect 198 -1334 199 -1310
rect 222 -1311 223 -1263
rect 247 -1334 248 -1310
rect 450 -1311 451 -1263
rect 485 -1334 486 -1310
rect 621 -1334 622 -1310
rect 681 -1334 682 -1310
rect 772 -1311 773 -1263
rect 786 -1311 787 -1263
rect 807 -1334 808 -1310
rect 905 -1311 906 -1263
rect 968 -1334 969 -1310
rect 184 -1313 185 -1263
rect 222 -1334 223 -1312
rect 275 -1334 276 -1312
rect 544 -1313 545 -1263
rect 562 -1313 563 -1263
rect 772 -1334 773 -1312
rect 933 -1313 934 -1263
rect 975 -1334 976 -1312
rect 44 -1315 45 -1263
rect 184 -1334 185 -1314
rect 201 -1315 202 -1263
rect 394 -1315 395 -1263
rect 432 -1315 433 -1263
rect 450 -1334 451 -1314
rect 509 -1334 510 -1314
rect 562 -1334 563 -1314
rect 688 -1334 689 -1314
rect 709 -1315 710 -1263
rect 716 -1334 717 -1314
rect 758 -1315 759 -1263
rect 877 -1315 878 -1263
rect 933 -1334 934 -1314
rect 44 -1334 45 -1316
rect 177 -1317 178 -1263
rect 205 -1317 206 -1263
rect 233 -1334 234 -1316
rect 296 -1334 297 -1316
rect 499 -1317 500 -1263
rect 709 -1334 710 -1316
rect 723 -1317 724 -1263
rect 758 -1334 759 -1316
rect 905 -1334 906 -1316
rect 156 -1319 157 -1263
rect 205 -1334 206 -1318
rect 212 -1319 213 -1263
rect 226 -1334 227 -1318
rect 345 -1334 346 -1318
rect 457 -1319 458 -1263
rect 499 -1334 500 -1318
rect 1048 -1334 1049 -1318
rect 212 -1334 213 -1320
rect 303 -1321 304 -1263
rect 355 -1334 356 -1320
rect 786 -1334 787 -1320
rect 828 -1321 829 -1263
rect 877 -1334 878 -1320
rect 37 -1323 38 -1263
rect 303 -1334 304 -1322
rect 380 -1323 381 -1263
rect 394 -1334 395 -1322
rect 432 -1334 433 -1322
rect 513 -1334 514 -1322
rect 597 -1323 598 -1263
rect 723 -1334 724 -1322
rect 37 -1334 38 -1324
rect 219 -1334 220 -1324
rect 380 -1334 381 -1324
rect 401 -1325 402 -1263
rect 422 -1334 423 -1324
rect 597 -1334 598 -1324
rect 401 -1334 402 -1326
rect 408 -1327 409 -1263
rect 457 -1334 458 -1326
rect 849 -1334 850 -1326
rect 408 -1334 409 -1328
rect 569 -1329 570 -1263
rect 492 -1331 493 -1263
rect 828 -1334 829 -1330
rect 415 -1334 416 -1332
rect 492 -1334 493 -1332
rect 569 -1334 570 -1332
rect 579 -1334 580 -1332
rect 16 -1344 17 -1342
rect 79 -1344 80 -1342
rect 89 -1411 90 -1343
rect 296 -1344 297 -1342
rect 303 -1344 304 -1342
rect 327 -1344 328 -1342
rect 352 -1344 353 -1342
rect 380 -1344 381 -1342
rect 387 -1344 388 -1342
rect 432 -1344 433 -1342
rect 471 -1344 472 -1342
rect 632 -1344 633 -1342
rect 646 -1344 647 -1342
rect 905 -1344 906 -1342
rect 919 -1344 920 -1342
rect 919 -1411 920 -1343
rect 919 -1344 920 -1342
rect 919 -1411 920 -1343
rect 950 -1411 951 -1343
rect 996 -1344 997 -1342
rect 1031 -1344 1032 -1342
rect 1052 -1344 1053 -1342
rect 16 -1411 17 -1345
rect 173 -1346 174 -1342
rect 222 -1346 223 -1342
rect 282 -1346 283 -1342
rect 292 -1346 293 -1342
rect 534 -1411 535 -1345
rect 576 -1346 577 -1342
rect 842 -1346 843 -1342
rect 891 -1346 892 -1342
rect 905 -1411 906 -1345
rect 1024 -1346 1025 -1342
rect 1031 -1411 1032 -1345
rect 1038 -1346 1039 -1342
rect 1073 -1346 1074 -1342
rect 23 -1348 24 -1342
rect 86 -1348 87 -1342
rect 107 -1348 108 -1342
rect 170 -1411 171 -1347
rect 222 -1411 223 -1347
rect 310 -1348 311 -1342
rect 338 -1348 339 -1342
rect 352 -1411 353 -1347
rect 366 -1411 367 -1347
rect 450 -1348 451 -1342
rect 471 -1411 472 -1347
rect 590 -1348 591 -1342
rect 597 -1348 598 -1342
rect 912 -1348 913 -1342
rect 971 -1411 972 -1347
rect 1024 -1411 1025 -1347
rect 1045 -1411 1046 -1347
rect 1048 -1348 1049 -1342
rect 1073 -1411 1074 -1347
rect 1080 -1348 1081 -1342
rect 9 -1350 10 -1342
rect 86 -1411 87 -1349
rect 107 -1411 108 -1349
rect 331 -1350 332 -1342
rect 338 -1411 339 -1349
rect 464 -1350 465 -1342
rect 495 -1350 496 -1342
rect 723 -1350 724 -1342
rect 737 -1350 738 -1342
rect 870 -1350 871 -1342
rect 30 -1352 31 -1342
rect 61 -1411 62 -1351
rect 65 -1352 66 -1342
rect 68 -1384 69 -1351
rect 79 -1411 80 -1351
rect 355 -1352 356 -1342
rect 380 -1411 381 -1351
rect 394 -1352 395 -1342
rect 411 -1411 412 -1351
rect 562 -1352 563 -1342
rect 576 -1411 577 -1351
rect 681 -1352 682 -1342
rect 705 -1352 706 -1342
rect 744 -1352 745 -1342
rect 758 -1352 759 -1342
rect 975 -1352 976 -1342
rect 30 -1411 31 -1353
rect 100 -1354 101 -1342
rect 114 -1411 115 -1353
rect 219 -1354 220 -1342
rect 254 -1354 255 -1342
rect 310 -1411 311 -1353
rect 331 -1411 332 -1353
rect 548 -1354 549 -1342
rect 579 -1354 580 -1342
rect 940 -1354 941 -1342
rect 961 -1354 962 -1342
rect 975 -1411 976 -1353
rect 37 -1356 38 -1342
rect 135 -1411 136 -1355
rect 138 -1356 139 -1342
rect 401 -1356 402 -1342
rect 415 -1356 416 -1342
rect 457 -1411 458 -1355
rect 506 -1356 507 -1342
rect 688 -1356 689 -1342
rect 705 -1411 706 -1355
rect 1017 -1356 1018 -1342
rect 37 -1411 38 -1357
rect 44 -1358 45 -1342
rect 51 -1358 52 -1342
rect 177 -1358 178 -1342
rect 254 -1411 255 -1357
rect 506 -1411 507 -1357
rect 509 -1411 510 -1357
rect 695 -1358 696 -1342
rect 723 -1411 724 -1357
rect 786 -1358 787 -1342
rect 821 -1358 822 -1342
rect 821 -1411 822 -1357
rect 821 -1358 822 -1342
rect 821 -1411 822 -1357
rect 835 -1358 836 -1342
rect 891 -1411 892 -1357
rect 44 -1411 45 -1359
rect 345 -1360 346 -1342
rect 401 -1411 402 -1359
rect 569 -1360 570 -1342
rect 590 -1411 591 -1359
rect 604 -1360 605 -1342
rect 618 -1360 619 -1342
rect 968 -1360 969 -1342
rect 54 -1411 55 -1361
rect 600 -1362 601 -1342
rect 611 -1362 612 -1342
rect 618 -1411 619 -1361
rect 632 -1411 633 -1361
rect 751 -1362 752 -1342
rect 758 -1411 759 -1361
rect 779 -1362 780 -1342
rect 835 -1411 836 -1361
rect 856 -1362 857 -1342
rect 863 -1362 864 -1342
rect 961 -1411 962 -1361
rect 65 -1411 66 -1363
rect 93 -1364 94 -1342
rect 100 -1411 101 -1363
rect 422 -1364 423 -1342
rect 429 -1364 430 -1342
rect 996 -1411 997 -1363
rect 93 -1411 94 -1365
rect 478 -1366 479 -1342
rect 523 -1411 524 -1365
rect 604 -1411 605 -1365
rect 611 -1411 612 -1365
rect 674 -1366 675 -1342
rect 684 -1411 685 -1365
rect 940 -1411 941 -1365
rect 121 -1368 122 -1342
rect 194 -1368 195 -1342
rect 247 -1368 248 -1342
rect 345 -1411 346 -1367
rect 355 -1411 356 -1367
rect 422 -1411 423 -1367
rect 429 -1411 430 -1367
rect 516 -1411 517 -1367
rect 548 -1411 549 -1367
rect 677 -1368 678 -1342
rect 688 -1411 689 -1367
rect 702 -1368 703 -1342
rect 709 -1368 710 -1342
rect 786 -1411 787 -1367
rect 842 -1411 843 -1367
rect 898 -1368 899 -1342
rect 58 -1370 59 -1342
rect 121 -1411 122 -1369
rect 128 -1370 129 -1342
rect 513 -1370 514 -1342
rect 572 -1411 573 -1369
rect 751 -1411 752 -1369
rect 765 -1370 766 -1342
rect 1052 -1411 1053 -1369
rect 128 -1411 129 -1371
rect 208 -1411 209 -1371
rect 268 -1372 269 -1342
rect 296 -1411 297 -1371
rect 303 -1411 304 -1371
rect 709 -1411 710 -1371
rect 730 -1372 731 -1342
rect 744 -1411 745 -1371
rect 779 -1411 780 -1371
rect 800 -1372 801 -1342
rect 849 -1372 850 -1342
rect 912 -1411 913 -1371
rect 145 -1411 146 -1373
rect 156 -1411 157 -1373
rect 159 -1374 160 -1342
rect 541 -1374 542 -1342
rect 579 -1411 580 -1373
rect 863 -1411 864 -1373
rect 870 -1411 871 -1373
rect 877 -1374 878 -1342
rect 884 -1374 885 -1342
rect 898 -1411 899 -1373
rect 149 -1376 150 -1342
rect 268 -1411 269 -1375
rect 275 -1376 276 -1342
rect 394 -1411 395 -1375
rect 415 -1411 416 -1375
rect 663 -1411 664 -1375
rect 674 -1411 675 -1375
rect 716 -1376 717 -1342
rect 737 -1411 738 -1375
rect 772 -1376 773 -1342
rect 800 -1411 801 -1375
rect 807 -1376 808 -1342
rect 884 -1411 885 -1375
rect 982 -1376 983 -1342
rect 149 -1411 150 -1377
rect 180 -1378 181 -1342
rect 184 -1378 185 -1342
rect 247 -1411 248 -1377
rect 261 -1378 262 -1342
rect 275 -1411 276 -1377
rect 282 -1411 283 -1377
rect 387 -1411 388 -1377
rect 450 -1411 451 -1377
rect 499 -1378 500 -1342
rect 583 -1378 584 -1342
rect 856 -1411 857 -1377
rect 982 -1411 983 -1377
rect 989 -1378 990 -1342
rect 163 -1380 164 -1342
rect 191 -1411 192 -1379
rect 205 -1380 206 -1342
rect 261 -1411 262 -1379
rect 324 -1380 325 -1342
rect 478 -1411 479 -1379
rect 492 -1380 493 -1342
rect 807 -1411 808 -1379
rect 23 -1411 24 -1381
rect 205 -1411 206 -1381
rect 324 -1411 325 -1381
rect 373 -1382 374 -1342
rect 443 -1382 444 -1342
rect 499 -1411 500 -1381
rect 583 -1411 584 -1381
rect 954 -1382 955 -1342
rect 373 -1411 374 -1383
rect 443 -1411 444 -1383
rect 485 -1384 486 -1342
rect 492 -1411 493 -1383
rect 520 -1384 521 -1342
rect 586 -1411 587 -1383
rect 989 -1411 990 -1383
rect 163 -1411 164 -1385
rect 289 -1411 290 -1385
rect 359 -1386 360 -1342
rect 730 -1411 731 -1385
rect 772 -1411 773 -1385
rect 828 -1386 829 -1342
rect 947 -1386 948 -1342
rect 954 -1411 955 -1385
rect 177 -1411 178 -1387
rect 198 -1388 199 -1342
rect 359 -1411 360 -1387
rect 436 -1388 437 -1342
rect 464 -1411 465 -1387
rect 569 -1411 570 -1387
rect 597 -1411 598 -1387
rect 1066 -1388 1067 -1342
rect 184 -1411 185 -1389
rect 317 -1390 318 -1342
rect 369 -1390 370 -1342
rect 849 -1411 850 -1389
rect 198 -1411 199 -1391
rect 233 -1392 234 -1342
rect 317 -1411 318 -1391
rect 460 -1392 461 -1342
rect 485 -1411 486 -1391
rect 555 -1392 556 -1342
rect 565 -1411 566 -1391
rect 828 -1411 829 -1391
rect 72 -1394 73 -1342
rect 555 -1411 556 -1393
rect 646 -1411 647 -1393
rect 653 -1394 654 -1342
rect 660 -1394 661 -1342
rect 716 -1411 717 -1393
rect 72 -1411 73 -1395
rect 226 -1396 227 -1342
rect 408 -1396 409 -1342
rect 520 -1411 521 -1395
rect 653 -1411 654 -1395
rect 1034 -1396 1035 -1342
rect 142 -1398 143 -1342
rect 226 -1411 227 -1397
rect 408 -1411 409 -1397
rect 541 -1411 542 -1397
rect 660 -1411 661 -1397
rect 1010 -1398 1011 -1342
rect 212 -1400 213 -1342
rect 233 -1411 234 -1399
rect 436 -1411 437 -1399
rect 527 -1400 528 -1342
rect 681 -1411 682 -1399
rect 877 -1411 878 -1399
rect 1003 -1400 1004 -1342
rect 1010 -1411 1011 -1399
rect 212 -1411 213 -1401
rect 240 -1402 241 -1342
rect 527 -1411 528 -1401
rect 625 -1402 626 -1342
rect 695 -1411 696 -1401
rect 814 -1402 815 -1342
rect 1003 -1411 1004 -1401
rect 1017 -1411 1018 -1401
rect 625 -1411 626 -1403
rect 667 -1404 668 -1342
rect 814 -1411 815 -1403
rect 933 -1404 934 -1342
rect 639 -1406 640 -1342
rect 667 -1411 668 -1405
rect 926 -1406 927 -1342
rect 933 -1411 934 -1405
rect 639 -1411 640 -1407
rect 793 -1408 794 -1342
rect 649 -1410 650 -1342
rect 793 -1411 794 -1409
rect 16 -1421 17 -1419
rect 124 -1492 125 -1420
rect 135 -1492 136 -1420
rect 296 -1421 297 -1419
rect 310 -1421 311 -1419
rect 359 -1492 360 -1420
rect 380 -1421 381 -1419
rect 380 -1492 381 -1420
rect 380 -1421 381 -1419
rect 380 -1492 381 -1420
rect 390 -1421 391 -1419
rect 450 -1421 451 -1419
rect 471 -1421 472 -1419
rect 537 -1492 538 -1420
rect 569 -1421 570 -1419
rect 674 -1421 675 -1419
rect 681 -1421 682 -1419
rect 800 -1421 801 -1419
rect 828 -1421 829 -1419
rect 831 -1449 832 -1420
rect 842 -1421 843 -1419
rect 943 -1492 944 -1420
rect 971 -1421 972 -1419
rect 1031 -1421 1032 -1419
rect 1066 -1492 1067 -1420
rect 1073 -1421 1074 -1419
rect 23 -1423 24 -1419
rect 222 -1423 223 -1419
rect 268 -1423 269 -1419
rect 306 -1423 307 -1419
rect 310 -1492 311 -1422
rect 737 -1492 738 -1422
rect 758 -1423 759 -1419
rect 758 -1492 759 -1422
rect 758 -1423 759 -1419
rect 758 -1492 759 -1422
rect 793 -1423 794 -1419
rect 950 -1423 951 -1419
rect 975 -1423 976 -1419
rect 1003 -1492 1004 -1422
rect 1010 -1423 1011 -1419
rect 1038 -1492 1039 -1422
rect 30 -1425 31 -1419
rect 159 -1425 160 -1419
rect 163 -1425 164 -1419
rect 303 -1425 304 -1419
rect 338 -1425 339 -1419
rect 562 -1425 563 -1419
rect 579 -1492 580 -1424
rect 786 -1425 787 -1419
rect 793 -1492 794 -1424
rect 821 -1425 822 -1419
rect 828 -1492 829 -1424
rect 849 -1425 850 -1419
rect 877 -1425 878 -1419
rect 968 -1425 969 -1419
rect 1024 -1425 1025 -1419
rect 1041 -1425 1042 -1419
rect 30 -1492 31 -1426
rect 51 -1427 52 -1419
rect 54 -1492 55 -1426
rect 128 -1427 129 -1419
rect 138 -1427 139 -1419
rect 142 -1427 143 -1419
rect 163 -1492 164 -1426
rect 212 -1427 213 -1419
rect 219 -1427 220 -1419
rect 653 -1427 654 -1419
rect 663 -1427 664 -1419
rect 779 -1427 780 -1419
rect 821 -1492 822 -1426
rect 905 -1427 906 -1419
rect 929 -1427 930 -1419
rect 961 -1427 962 -1419
rect 44 -1429 45 -1419
rect 128 -1492 129 -1428
rect 142 -1492 143 -1428
rect 170 -1429 171 -1419
rect 205 -1429 206 -1419
rect 891 -1429 892 -1419
rect 44 -1492 45 -1430
rect 187 -1492 188 -1430
rect 205 -1492 206 -1430
rect 240 -1431 241 -1419
rect 289 -1431 290 -1419
rect 471 -1492 472 -1430
rect 499 -1431 500 -1419
rect 513 -1431 514 -1419
rect 516 -1431 517 -1419
rect 716 -1431 717 -1419
rect 744 -1431 745 -1419
rect 975 -1492 976 -1430
rect 58 -1492 59 -1432
rect 684 -1492 685 -1432
rect 688 -1433 689 -1419
rect 716 -1492 717 -1432
rect 723 -1433 724 -1419
rect 744 -1492 745 -1432
rect 772 -1433 773 -1419
rect 786 -1492 787 -1432
rect 835 -1433 836 -1419
rect 849 -1492 850 -1432
rect 877 -1492 878 -1432
rect 926 -1433 927 -1419
rect 65 -1435 66 -1419
rect 65 -1492 66 -1434
rect 65 -1435 66 -1419
rect 65 -1492 66 -1434
rect 72 -1435 73 -1419
rect 401 -1435 402 -1419
rect 408 -1435 409 -1419
rect 520 -1492 521 -1434
rect 523 -1435 524 -1419
rect 625 -1435 626 -1419
rect 635 -1492 636 -1434
rect 807 -1435 808 -1419
rect 835 -1492 836 -1434
rect 870 -1435 871 -1419
rect 884 -1435 885 -1419
rect 922 -1492 923 -1434
rect 926 -1492 927 -1434
rect 954 -1435 955 -1419
rect 37 -1437 38 -1419
rect 72 -1492 73 -1436
rect 75 -1492 76 -1436
rect 296 -1492 297 -1436
rect 338 -1492 339 -1436
rect 586 -1437 587 -1419
rect 597 -1437 598 -1419
rect 688 -1492 689 -1436
rect 712 -1437 713 -1419
rect 814 -1437 815 -1419
rect 842 -1492 843 -1436
rect 940 -1437 941 -1419
rect 954 -1492 955 -1436
rect 1017 -1437 1018 -1419
rect 37 -1492 38 -1438
rect 149 -1439 150 -1419
rect 170 -1492 171 -1438
rect 177 -1439 178 -1419
rect 212 -1492 213 -1438
rect 317 -1439 318 -1419
rect 345 -1439 346 -1419
rect 387 -1492 388 -1438
rect 394 -1439 395 -1419
rect 408 -1492 409 -1438
rect 411 -1439 412 -1419
rect 485 -1439 486 -1419
rect 513 -1492 514 -1438
rect 709 -1439 710 -1419
rect 765 -1439 766 -1419
rect 884 -1492 885 -1438
rect 86 -1441 87 -1419
rect 779 -1492 780 -1440
rect 807 -1492 808 -1440
rect 856 -1441 857 -1419
rect 870 -1492 871 -1440
rect 989 -1441 990 -1419
rect 26 -1492 27 -1442
rect 86 -1492 87 -1442
rect 89 -1443 90 -1419
rect 772 -1492 773 -1442
rect 814 -1492 815 -1442
rect 863 -1443 864 -1419
rect 947 -1443 948 -1419
rect 989 -1492 990 -1442
rect 93 -1445 94 -1419
rect 499 -1492 500 -1444
rect 555 -1445 556 -1419
rect 569 -1492 570 -1444
rect 583 -1445 584 -1419
rect 618 -1445 619 -1419
rect 639 -1445 640 -1419
rect 674 -1492 675 -1444
rect 681 -1492 682 -1444
rect 898 -1445 899 -1419
rect 912 -1445 913 -1419
rect 947 -1492 948 -1444
rect 93 -1492 94 -1446
rect 198 -1447 199 -1419
rect 219 -1492 220 -1446
rect 261 -1447 262 -1419
rect 292 -1492 293 -1446
rect 345 -1492 346 -1446
rect 352 -1492 353 -1446
rect 541 -1447 542 -1419
rect 555 -1492 556 -1446
rect 611 -1447 612 -1419
rect 632 -1447 633 -1419
rect 639 -1492 640 -1446
rect 646 -1447 647 -1419
rect 709 -1492 710 -1446
rect 726 -1492 727 -1446
rect 898 -1492 899 -1446
rect 100 -1449 101 -1419
rect 565 -1492 566 -1448
rect 604 -1449 605 -1419
rect 768 -1449 769 -1419
rect 912 -1492 913 -1448
rect 79 -1451 80 -1419
rect 100 -1492 101 -1450
rect 107 -1451 108 -1419
rect 656 -1492 657 -1450
rect 660 -1451 661 -1419
rect 891 -1492 892 -1450
rect 79 -1492 80 -1452
rect 324 -1453 325 -1419
rect 362 -1453 363 -1419
rect 597 -1492 598 -1452
rect 611 -1492 612 -1452
rect 730 -1453 731 -1419
rect 751 -1453 752 -1419
rect 765 -1492 766 -1452
rect 856 -1492 857 -1452
rect 919 -1453 920 -1419
rect 107 -1492 108 -1454
rect 576 -1455 577 -1419
rect 667 -1455 668 -1419
rect 730 -1492 731 -1454
rect 863 -1492 864 -1454
rect 933 -1455 934 -1419
rect 121 -1457 122 -1419
rect 243 -1457 244 -1419
rect 247 -1457 248 -1419
rect 324 -1492 325 -1456
rect 397 -1492 398 -1456
rect 1052 -1457 1053 -1419
rect 121 -1492 122 -1458
rect 268 -1492 269 -1458
rect 317 -1492 318 -1458
rect 415 -1459 416 -1419
rect 418 -1492 419 -1458
rect 457 -1459 458 -1419
rect 478 -1459 479 -1419
rect 604 -1492 605 -1458
rect 702 -1459 703 -1419
rect 751 -1492 752 -1458
rect 919 -1492 920 -1458
rect 1045 -1459 1046 -1419
rect 149 -1492 150 -1460
rect 429 -1461 430 -1419
rect 450 -1492 451 -1460
rect 464 -1461 465 -1419
rect 478 -1492 479 -1460
rect 590 -1461 591 -1419
rect 695 -1461 696 -1419
rect 702 -1492 703 -1460
rect 933 -1492 934 -1460
rect 996 -1461 997 -1419
rect 166 -1463 167 -1419
rect 583 -1492 584 -1462
rect 590 -1492 591 -1462
rect 1006 -1463 1007 -1419
rect 177 -1492 178 -1464
rect 191 -1465 192 -1419
rect 198 -1492 199 -1464
rect 394 -1492 395 -1464
rect 401 -1492 402 -1464
rect 558 -1492 559 -1464
rect 562 -1492 563 -1464
rect 667 -1492 668 -1464
rect 695 -1492 696 -1464
rect 940 -1492 941 -1464
rect 982 -1465 983 -1419
rect 996 -1492 997 -1464
rect 184 -1467 185 -1419
rect 261 -1492 262 -1466
rect 366 -1467 367 -1419
rect 429 -1492 430 -1466
rect 457 -1492 458 -1466
rect 534 -1467 535 -1419
rect 618 -1492 619 -1466
rect 982 -1492 983 -1466
rect 184 -1492 185 -1468
rect 331 -1469 332 -1419
rect 366 -1492 367 -1468
rect 373 -1469 374 -1419
rect 415 -1492 416 -1468
rect 625 -1492 626 -1468
rect 191 -1492 192 -1470
rect 506 -1471 507 -1419
rect 527 -1471 528 -1419
rect 646 -1492 647 -1470
rect 243 -1492 244 -1472
rect 660 -1492 661 -1472
rect 247 -1492 248 -1474
rect 306 -1492 307 -1474
rect 320 -1492 321 -1474
rect 331 -1492 332 -1474
rect 355 -1475 356 -1419
rect 373 -1492 374 -1474
rect 443 -1475 444 -1419
rect 527 -1492 528 -1474
rect 51 -1492 52 -1476
rect 443 -1492 444 -1476
rect 464 -1492 465 -1476
rect 492 -1477 493 -1419
rect 506 -1492 507 -1476
rect 548 -1477 549 -1419
rect 254 -1479 255 -1419
rect 289 -1492 290 -1478
rect 422 -1479 423 -1419
rect 492 -1492 493 -1478
rect 548 -1492 549 -1478
rect 971 -1492 972 -1478
rect 233 -1481 234 -1419
rect 254 -1492 255 -1480
rect 422 -1492 423 -1480
rect 436 -1481 437 -1419
rect 485 -1492 486 -1480
rect 544 -1492 545 -1480
rect 114 -1483 115 -1419
rect 233 -1492 234 -1482
rect 436 -1492 437 -1482
rect 905 -1492 906 -1482
rect 114 -1492 115 -1484
rect 282 -1485 283 -1419
rect 275 -1487 276 -1419
rect 282 -1492 283 -1486
rect 226 -1489 227 -1419
rect 275 -1492 276 -1488
rect 156 -1492 157 -1490
rect 226 -1492 227 -1490
rect 9 -1589 10 -1501
rect 401 -1502 402 -1500
rect 418 -1502 419 -1500
rect 492 -1502 493 -1500
rect 506 -1502 507 -1500
rect 544 -1502 545 -1500
rect 558 -1502 559 -1500
rect 765 -1502 766 -1500
rect 800 -1502 801 -1500
rect 835 -1502 836 -1500
rect 856 -1502 857 -1500
rect 968 -1589 969 -1501
rect 996 -1502 997 -1500
rect 996 -1589 997 -1501
rect 996 -1502 997 -1500
rect 996 -1589 997 -1501
rect 1038 -1502 1039 -1500
rect 1073 -1589 1074 -1501
rect 16 -1589 17 -1503
rect 149 -1504 150 -1500
rect 194 -1589 195 -1503
rect 499 -1504 500 -1500
rect 506 -1589 507 -1503
rect 712 -1589 713 -1503
rect 726 -1504 727 -1500
rect 807 -1504 808 -1500
rect 835 -1589 836 -1503
rect 1111 -1589 1112 -1503
rect 23 -1589 24 -1505
rect 163 -1506 164 -1500
rect 226 -1506 227 -1500
rect 359 -1506 360 -1500
rect 366 -1506 367 -1500
rect 366 -1589 367 -1505
rect 366 -1506 367 -1500
rect 366 -1589 367 -1505
rect 380 -1506 381 -1500
rect 380 -1589 381 -1505
rect 380 -1506 381 -1500
rect 380 -1589 381 -1505
rect 394 -1506 395 -1500
rect 1101 -1589 1102 -1505
rect 30 -1508 31 -1500
rect 243 -1508 244 -1500
rect 268 -1508 269 -1500
rect 317 -1508 318 -1500
rect 327 -1589 328 -1507
rect 625 -1508 626 -1500
rect 667 -1508 668 -1500
rect 765 -1589 766 -1507
rect 870 -1508 871 -1500
rect 1066 -1589 1067 -1507
rect 30 -1589 31 -1509
rect 142 -1510 143 -1500
rect 149 -1589 150 -1509
rect 397 -1510 398 -1500
rect 418 -1589 419 -1509
rect 520 -1510 521 -1500
rect 534 -1510 535 -1500
rect 807 -1589 808 -1509
rect 870 -1589 871 -1509
rect 982 -1510 983 -1500
rect 1003 -1510 1004 -1500
rect 1038 -1589 1039 -1509
rect 37 -1512 38 -1500
rect 240 -1512 241 -1500
rect 268 -1589 269 -1511
rect 324 -1512 325 -1500
rect 341 -1589 342 -1511
rect 828 -1512 829 -1500
rect 842 -1512 843 -1500
rect 1003 -1589 1004 -1511
rect 37 -1589 38 -1513
rect 656 -1514 657 -1500
rect 681 -1514 682 -1500
rect 884 -1514 885 -1500
rect 891 -1514 892 -1500
rect 1108 -1589 1109 -1513
rect 51 -1589 52 -1515
rect 100 -1516 101 -1500
rect 121 -1516 122 -1500
rect 940 -1589 941 -1515
rect 947 -1516 948 -1500
rect 971 -1516 972 -1500
rect 58 -1518 59 -1500
rect 124 -1589 125 -1517
rect 128 -1589 129 -1517
rect 156 -1518 157 -1500
rect 163 -1589 164 -1517
rect 212 -1518 213 -1500
rect 229 -1589 230 -1517
rect 261 -1518 262 -1500
rect 275 -1518 276 -1500
rect 303 -1518 304 -1500
rect 317 -1589 318 -1517
rect 478 -1518 479 -1500
rect 513 -1518 514 -1500
rect 555 -1589 556 -1517
rect 562 -1518 563 -1500
rect 702 -1518 703 -1500
rect 733 -1589 734 -1517
rect 1080 -1589 1081 -1517
rect 58 -1589 59 -1519
rect 376 -1589 377 -1519
rect 422 -1520 423 -1500
rect 625 -1589 626 -1519
rect 646 -1520 647 -1500
rect 982 -1589 983 -1519
rect 65 -1522 66 -1500
rect 86 -1522 87 -1500
rect 93 -1522 94 -1500
rect 313 -1522 314 -1500
rect 352 -1522 353 -1500
rect 439 -1522 440 -1500
rect 450 -1522 451 -1500
rect 513 -1589 514 -1521
rect 520 -1589 521 -1521
rect 537 -1522 538 -1500
rect 562 -1589 563 -1521
rect 597 -1522 598 -1500
rect 618 -1522 619 -1500
rect 842 -1589 843 -1521
rect 877 -1522 878 -1500
rect 1017 -1589 1018 -1521
rect 44 -1524 45 -1500
rect 65 -1589 66 -1523
rect 72 -1589 73 -1523
rect 828 -1589 829 -1523
rect 877 -1589 878 -1523
rect 933 -1524 934 -1500
rect 954 -1524 955 -1500
rect 1094 -1589 1095 -1523
rect 79 -1526 80 -1500
rect 544 -1589 545 -1525
rect 565 -1526 566 -1500
rect 814 -1526 815 -1500
rect 898 -1526 899 -1500
rect 1024 -1589 1025 -1525
rect 79 -1589 80 -1527
rect 548 -1528 549 -1500
rect 618 -1589 619 -1527
rect 695 -1528 696 -1500
rect 702 -1589 703 -1527
rect 730 -1528 731 -1500
rect 744 -1528 745 -1500
rect 856 -1589 857 -1527
rect 898 -1589 899 -1527
rect 975 -1528 976 -1500
rect 82 -1589 83 -1529
rect 478 -1589 479 -1529
rect 534 -1589 535 -1529
rect 1087 -1589 1088 -1529
rect 86 -1589 87 -1531
rect 170 -1532 171 -1500
rect 177 -1589 178 -1531
rect 226 -1589 227 -1531
rect 247 -1532 248 -1500
rect 275 -1589 276 -1531
rect 282 -1532 283 -1500
rect 352 -1589 353 -1531
rect 359 -1589 360 -1531
rect 632 -1589 633 -1531
rect 646 -1589 647 -1531
rect 800 -1589 801 -1531
rect 863 -1532 864 -1500
rect 975 -1589 976 -1531
rect 93 -1589 94 -1533
rect 415 -1534 416 -1500
rect 436 -1589 437 -1533
rect 803 -1534 804 -1500
rect 905 -1534 906 -1500
rect 1052 -1589 1053 -1533
rect 100 -1589 101 -1535
rect 240 -1589 241 -1535
rect 254 -1536 255 -1500
rect 303 -1589 304 -1535
rect 306 -1536 307 -1500
rect 905 -1589 906 -1535
rect 912 -1536 913 -1500
rect 919 -1589 920 -1535
rect 922 -1536 923 -1500
rect 961 -1589 962 -1535
rect 964 -1536 965 -1500
rect 989 -1536 990 -1500
rect 135 -1538 136 -1500
rect 394 -1589 395 -1537
rect 464 -1538 465 -1500
rect 499 -1589 500 -1537
rect 548 -1589 549 -1537
rect 611 -1538 612 -1500
rect 653 -1538 654 -1500
rect 947 -1589 948 -1537
rect 135 -1589 136 -1539
rect 457 -1540 458 -1500
rect 474 -1589 475 -1539
rect 709 -1540 710 -1500
rect 716 -1540 717 -1500
rect 814 -1589 815 -1539
rect 926 -1540 927 -1500
rect 1031 -1589 1032 -1539
rect 142 -1589 143 -1541
rect 345 -1542 346 -1500
rect 362 -1589 363 -1541
rect 954 -1589 955 -1541
rect 156 -1589 157 -1543
rect 429 -1544 430 -1500
rect 569 -1544 570 -1500
rect 611 -1589 612 -1543
rect 674 -1544 675 -1500
rect 891 -1589 892 -1543
rect 180 -1546 181 -1500
rect 212 -1589 213 -1545
rect 219 -1546 220 -1500
rect 282 -1589 283 -1545
rect 289 -1589 290 -1545
rect 576 -1546 577 -1500
rect 590 -1546 591 -1500
rect 653 -1589 654 -1545
rect 660 -1546 661 -1500
rect 674 -1589 675 -1545
rect 681 -1589 682 -1545
rect 821 -1546 822 -1500
rect 184 -1589 185 -1547
rect 324 -1589 325 -1547
rect 331 -1548 332 -1500
rect 597 -1589 598 -1547
rect 604 -1548 605 -1500
rect 716 -1589 717 -1547
rect 751 -1548 752 -1500
rect 863 -1589 864 -1547
rect 107 -1550 108 -1500
rect 331 -1589 332 -1549
rect 338 -1550 339 -1500
rect 569 -1589 570 -1549
rect 590 -1589 591 -1549
rect 688 -1550 689 -1500
rect 695 -1589 696 -1549
rect 737 -1550 738 -1500
rect 758 -1550 759 -1500
rect 1045 -1589 1046 -1549
rect 107 -1589 108 -1551
rect 114 -1552 115 -1500
rect 170 -1589 171 -1551
rect 338 -1589 339 -1551
rect 345 -1589 346 -1551
rect 443 -1552 444 -1500
rect 460 -1589 461 -1551
rect 737 -1589 738 -1551
rect 758 -1589 759 -1551
rect 912 -1589 913 -1551
rect 114 -1589 115 -1553
rect 450 -1589 451 -1553
rect 485 -1554 486 -1500
rect 751 -1589 752 -1553
rect 772 -1554 773 -1500
rect 884 -1589 885 -1553
rect 187 -1556 188 -1500
rect 439 -1589 440 -1555
rect 471 -1556 472 -1500
rect 485 -1589 486 -1555
rect 663 -1589 664 -1555
rect 688 -1589 689 -1555
rect 709 -1589 710 -1555
rect 1010 -1589 1011 -1555
rect 222 -1589 223 -1557
rect 660 -1589 661 -1557
rect 684 -1558 685 -1500
rect 989 -1589 990 -1557
rect 233 -1560 234 -1500
rect 457 -1589 458 -1559
rect 723 -1560 724 -1500
rect 772 -1589 773 -1559
rect 786 -1560 787 -1500
rect 933 -1589 934 -1559
rect 233 -1589 234 -1561
rect 667 -1589 668 -1561
rect 723 -1589 724 -1561
rect 779 -1562 780 -1500
rect 793 -1562 794 -1500
rect 926 -1589 927 -1561
rect 131 -1564 132 -1500
rect 793 -1589 794 -1563
rect 803 -1589 804 -1563
rect 1059 -1589 1060 -1563
rect 243 -1589 244 -1565
rect 576 -1589 577 -1565
rect 583 -1566 584 -1500
rect 786 -1589 787 -1565
rect 821 -1589 822 -1565
rect 849 -1566 850 -1500
rect 247 -1589 248 -1567
rect 684 -1589 685 -1567
rect 254 -1589 255 -1569
rect 292 -1570 293 -1500
rect 296 -1570 297 -1500
rect 604 -1589 605 -1569
rect 639 -1570 640 -1500
rect 779 -1589 780 -1569
rect 198 -1572 199 -1500
rect 296 -1589 297 -1571
rect 310 -1572 311 -1500
rect 744 -1589 745 -1571
rect 75 -1574 76 -1500
rect 310 -1589 311 -1573
rect 373 -1574 374 -1500
rect 464 -1589 465 -1573
rect 527 -1574 528 -1500
rect 639 -1589 640 -1573
rect 2 -1589 3 -1575
rect 373 -1589 374 -1575
rect 387 -1576 388 -1500
rect 422 -1589 423 -1575
rect 495 -1589 496 -1575
rect 527 -1589 528 -1575
rect 579 -1576 580 -1500
rect 849 -1589 850 -1575
rect 198 -1589 199 -1577
rect 205 -1578 206 -1500
rect 261 -1589 262 -1577
rect 471 -1589 472 -1577
rect 191 -1580 192 -1500
rect 205 -1589 206 -1579
rect 387 -1589 388 -1579
rect 516 -1589 517 -1579
rect 397 -1589 398 -1581
rect 443 -1589 444 -1581
rect 401 -1589 402 -1583
rect 583 -1589 584 -1583
rect 408 -1586 409 -1500
rect 429 -1589 430 -1585
rect 355 -1589 356 -1587
rect 408 -1589 409 -1587
rect 2 -1599 3 -1597
rect 299 -1676 300 -1598
rect 303 -1599 304 -1597
rect 324 -1676 325 -1598
rect 355 -1599 356 -1597
rect 786 -1599 787 -1597
rect 803 -1599 804 -1597
rect 1031 -1599 1032 -1597
rect 2 -1676 3 -1600
rect 159 -1676 160 -1600
rect 163 -1601 164 -1597
rect 341 -1601 342 -1597
rect 359 -1676 360 -1600
rect 429 -1601 430 -1597
rect 453 -1601 454 -1597
rect 982 -1601 983 -1597
rect 23 -1603 24 -1597
rect 250 -1603 251 -1597
rect 261 -1603 262 -1597
rect 352 -1676 353 -1602
rect 373 -1603 374 -1597
rect 583 -1603 584 -1597
rect 660 -1676 661 -1602
rect 688 -1603 689 -1597
rect 709 -1603 710 -1597
rect 1094 -1603 1095 -1597
rect 23 -1676 24 -1604
rect 107 -1605 108 -1597
rect 114 -1605 115 -1597
rect 114 -1676 115 -1604
rect 114 -1605 115 -1597
rect 114 -1676 115 -1604
rect 121 -1605 122 -1597
rect 793 -1605 794 -1597
rect 824 -1676 825 -1604
rect 919 -1605 920 -1597
rect 982 -1676 983 -1604
rect 1080 -1605 1081 -1597
rect 30 -1607 31 -1597
rect 233 -1607 234 -1597
rect 236 -1676 237 -1606
rect 254 -1607 255 -1597
rect 282 -1607 283 -1597
rect 415 -1676 416 -1606
rect 429 -1676 430 -1606
rect 527 -1607 528 -1597
rect 548 -1607 549 -1597
rect 548 -1676 549 -1606
rect 548 -1607 549 -1597
rect 548 -1676 549 -1606
rect 555 -1607 556 -1597
rect 709 -1676 710 -1606
rect 723 -1607 724 -1597
rect 800 -1676 801 -1606
rect 849 -1607 850 -1597
rect 915 -1676 916 -1606
rect 919 -1676 920 -1606
rect 968 -1607 969 -1597
rect 30 -1676 31 -1608
rect 485 -1609 486 -1597
rect 492 -1609 493 -1597
rect 590 -1609 591 -1597
rect 663 -1609 664 -1597
rect 891 -1609 892 -1597
rect 37 -1611 38 -1597
rect 47 -1611 48 -1597
rect 61 -1676 62 -1610
rect 450 -1611 451 -1597
rect 453 -1676 454 -1610
rect 898 -1611 899 -1597
rect 37 -1676 38 -1612
rect 128 -1613 129 -1597
rect 135 -1613 136 -1597
rect 362 -1613 363 -1597
rect 376 -1613 377 -1597
rect 380 -1613 381 -1597
rect 390 -1676 391 -1612
rect 576 -1613 577 -1597
rect 583 -1676 584 -1612
rect 611 -1613 612 -1597
rect 681 -1676 682 -1612
rect 737 -1613 738 -1597
rect 758 -1613 759 -1597
rect 1045 -1613 1046 -1597
rect 72 -1615 73 -1597
rect 828 -1615 829 -1597
rect 891 -1676 892 -1614
rect 961 -1615 962 -1597
rect 72 -1676 73 -1616
rect 443 -1617 444 -1597
rect 457 -1617 458 -1597
rect 779 -1617 780 -1597
rect 786 -1676 787 -1616
rect 835 -1617 836 -1597
rect 947 -1617 948 -1597
rect 961 -1676 962 -1616
rect 75 -1619 76 -1597
rect 240 -1676 241 -1618
rect 289 -1619 290 -1597
rect 373 -1676 374 -1618
rect 460 -1619 461 -1597
rect 541 -1676 542 -1618
rect 555 -1676 556 -1618
rect 1003 -1619 1004 -1597
rect 79 -1676 80 -1620
rect 632 -1621 633 -1597
rect 688 -1676 689 -1620
rect 702 -1621 703 -1597
rect 716 -1621 717 -1597
rect 898 -1676 899 -1620
rect 996 -1621 997 -1597
rect 1003 -1676 1004 -1620
rect 58 -1623 59 -1597
rect 632 -1676 633 -1622
rect 674 -1623 675 -1597
rect 716 -1676 717 -1622
rect 723 -1676 724 -1622
rect 765 -1623 766 -1597
rect 772 -1623 773 -1597
rect 849 -1676 850 -1622
rect 877 -1623 878 -1597
rect 947 -1676 948 -1622
rect 82 -1625 83 -1597
rect 597 -1625 598 -1597
rect 611 -1676 612 -1624
rect 639 -1625 640 -1597
rect 695 -1625 696 -1597
rect 758 -1676 759 -1624
rect 765 -1676 766 -1624
rect 856 -1625 857 -1597
rect 877 -1676 878 -1624
rect 975 -1625 976 -1597
rect 86 -1627 87 -1597
rect 243 -1627 244 -1597
rect 289 -1676 290 -1626
rect 310 -1627 311 -1597
rect 317 -1627 318 -1597
rect 537 -1627 538 -1597
rect 562 -1627 563 -1597
rect 576 -1676 577 -1626
rect 590 -1676 591 -1626
rect 618 -1627 619 -1597
rect 639 -1676 640 -1626
rect 954 -1627 955 -1597
rect 975 -1676 976 -1626
rect 1038 -1627 1039 -1597
rect 107 -1676 108 -1628
rect 338 -1629 339 -1597
rect 467 -1676 468 -1628
rect 1052 -1629 1053 -1597
rect 121 -1676 122 -1630
rect 194 -1631 195 -1597
rect 205 -1631 206 -1597
rect 261 -1676 262 -1630
rect 268 -1631 269 -1597
rect 338 -1676 339 -1630
rect 471 -1631 472 -1597
rect 695 -1676 696 -1630
rect 702 -1676 703 -1630
rect 744 -1631 745 -1597
rect 751 -1631 752 -1597
rect 954 -1676 955 -1630
rect 1052 -1676 1053 -1630
rect 1073 -1631 1074 -1597
rect 9 -1633 10 -1597
rect 205 -1676 206 -1632
rect 212 -1633 213 -1597
rect 254 -1676 255 -1632
rect 303 -1676 304 -1632
rect 408 -1633 409 -1597
rect 474 -1633 475 -1597
rect 1108 -1633 1109 -1597
rect 9 -1676 10 -1634
rect 135 -1676 136 -1634
rect 138 -1676 139 -1634
rect 268 -1676 269 -1634
rect 310 -1676 311 -1634
rect 387 -1635 388 -1597
rect 408 -1676 409 -1634
rect 646 -1635 647 -1597
rect 730 -1635 731 -1597
rect 1017 -1635 1018 -1597
rect 128 -1676 129 -1636
rect 184 -1637 185 -1597
rect 212 -1676 213 -1636
rect 842 -1637 843 -1597
rect 856 -1676 857 -1636
rect 926 -1637 927 -1597
rect 142 -1639 143 -1597
rect 401 -1639 402 -1597
rect 474 -1676 475 -1638
rect 737 -1676 738 -1638
rect 744 -1676 745 -1638
rect 814 -1639 815 -1597
rect 835 -1676 836 -1638
rect 933 -1639 934 -1597
rect 65 -1641 66 -1597
rect 401 -1676 402 -1640
rect 481 -1676 482 -1640
rect 905 -1641 906 -1597
rect 926 -1676 927 -1640
rect 1059 -1641 1060 -1597
rect 65 -1676 66 -1642
rect 124 -1643 125 -1597
rect 142 -1676 143 -1642
rect 177 -1643 178 -1597
rect 222 -1643 223 -1597
rect 296 -1643 297 -1597
rect 317 -1676 318 -1642
rect 436 -1643 437 -1597
rect 492 -1676 493 -1642
rect 828 -1676 829 -1642
rect 842 -1676 843 -1642
rect 940 -1643 941 -1597
rect 149 -1645 150 -1597
rect 184 -1676 185 -1644
rect 194 -1676 195 -1644
rect 436 -1676 437 -1644
rect 499 -1645 500 -1597
rect 527 -1676 528 -1644
rect 537 -1676 538 -1644
rect 1087 -1645 1088 -1597
rect 44 -1676 45 -1646
rect 149 -1676 150 -1646
rect 156 -1647 157 -1597
rect 443 -1676 444 -1646
rect 478 -1647 479 -1597
rect 499 -1676 500 -1646
rect 513 -1647 514 -1597
rect 1101 -1647 1102 -1597
rect 170 -1649 171 -1597
rect 534 -1676 535 -1648
rect 544 -1649 545 -1597
rect 618 -1676 619 -1648
rect 684 -1649 685 -1597
rect 940 -1676 941 -1648
rect 170 -1676 171 -1650
rect 198 -1651 199 -1597
rect 222 -1676 223 -1650
rect 275 -1651 276 -1597
rect 296 -1676 297 -1650
rect 506 -1651 507 -1597
rect 513 -1676 514 -1650
rect 887 -1676 888 -1650
rect 905 -1676 906 -1650
rect 1010 -1651 1011 -1597
rect 86 -1676 87 -1652
rect 198 -1676 199 -1652
rect 226 -1653 227 -1597
rect 870 -1653 871 -1597
rect 933 -1676 934 -1652
rect 1024 -1653 1025 -1597
rect 16 -1655 17 -1597
rect 226 -1676 227 -1654
rect 233 -1676 234 -1654
rect 282 -1676 283 -1654
rect 366 -1655 367 -1597
rect 506 -1676 507 -1654
rect 520 -1655 521 -1597
rect 674 -1676 675 -1654
rect 772 -1676 773 -1654
rect 894 -1676 895 -1654
rect 16 -1676 17 -1656
rect 51 -1657 52 -1597
rect 163 -1676 164 -1656
rect 366 -1676 367 -1656
rect 387 -1676 388 -1656
rect 450 -1676 451 -1656
rect 565 -1676 566 -1656
rect 1066 -1657 1067 -1597
rect 51 -1676 52 -1658
rect 569 -1659 570 -1597
rect 597 -1676 598 -1658
rect 625 -1659 626 -1597
rect 779 -1676 780 -1658
rect 884 -1659 885 -1597
rect 177 -1676 178 -1660
rect 422 -1661 423 -1597
rect 558 -1676 559 -1660
rect 569 -1676 570 -1660
rect 604 -1661 605 -1597
rect 751 -1676 752 -1660
rect 793 -1676 794 -1660
rect 863 -1661 864 -1597
rect 100 -1663 101 -1597
rect 422 -1676 423 -1662
rect 464 -1663 465 -1597
rect 604 -1676 605 -1662
rect 625 -1676 626 -1662
rect 653 -1663 654 -1597
rect 814 -1676 815 -1662
rect 912 -1663 913 -1597
rect 100 -1676 101 -1664
rect 247 -1665 248 -1597
rect 275 -1676 276 -1664
rect 807 -1665 808 -1597
rect 821 -1665 822 -1597
rect 870 -1676 871 -1664
rect 93 -1667 94 -1597
rect 247 -1676 248 -1666
rect 345 -1667 346 -1597
rect 520 -1676 521 -1666
rect 653 -1676 654 -1666
rect 667 -1667 668 -1597
rect 733 -1667 734 -1597
rect 807 -1676 808 -1666
rect 863 -1676 864 -1666
rect 989 -1667 990 -1597
rect 345 -1676 346 -1668
rect 457 -1676 458 -1668
rect 478 -1676 479 -1668
rect 821 -1676 822 -1668
rect 394 -1671 395 -1597
rect 646 -1676 647 -1670
rect 331 -1673 332 -1597
rect 394 -1676 395 -1672
rect 488 -1676 489 -1672
rect 667 -1676 668 -1672
rect 331 -1676 332 -1674
rect 464 -1676 465 -1674
rect 2 -1686 3 -1684
rect 376 -1771 377 -1685
rect 443 -1686 444 -1684
rect 562 -1686 563 -1684
rect 593 -1771 594 -1685
rect 1017 -1771 1018 -1685
rect 1024 -1686 1025 -1684
rect 1024 -1771 1025 -1685
rect 1024 -1686 1025 -1684
rect 1024 -1771 1025 -1685
rect 1027 -1686 1028 -1684
rect 1052 -1686 1053 -1684
rect 2 -1771 3 -1687
rect 96 -1688 97 -1684
rect 110 -1771 111 -1687
rect 128 -1688 129 -1684
rect 152 -1688 153 -1684
rect 275 -1688 276 -1684
rect 282 -1771 283 -1687
rect 394 -1688 395 -1684
rect 429 -1688 430 -1684
rect 562 -1771 563 -1687
rect 621 -1771 622 -1687
rect 716 -1688 717 -1684
rect 730 -1688 731 -1684
rect 870 -1688 871 -1684
rect 887 -1688 888 -1684
rect 961 -1688 962 -1684
rect 1003 -1688 1004 -1684
rect 1010 -1771 1011 -1687
rect 9 -1690 10 -1684
rect 191 -1690 192 -1684
rect 198 -1690 199 -1684
rect 597 -1690 598 -1684
rect 649 -1771 650 -1689
rect 856 -1690 857 -1684
rect 891 -1690 892 -1684
rect 982 -1690 983 -1684
rect 16 -1692 17 -1684
rect 215 -1692 216 -1684
rect 233 -1771 234 -1691
rect 436 -1692 437 -1684
rect 443 -1771 444 -1691
rect 677 -1771 678 -1691
rect 716 -1771 717 -1691
rect 723 -1692 724 -1684
rect 730 -1771 731 -1691
rect 758 -1692 759 -1684
rect 779 -1692 780 -1684
rect 782 -1706 783 -1691
rect 803 -1771 804 -1691
rect 807 -1692 808 -1684
rect 821 -1692 822 -1684
rect 968 -1771 969 -1691
rect 23 -1694 24 -1684
rect 194 -1694 195 -1684
rect 198 -1771 199 -1693
rect 254 -1694 255 -1684
rect 275 -1771 276 -1693
rect 733 -1694 734 -1684
rect 779 -1771 780 -1693
rect 814 -1694 815 -1684
rect 835 -1694 836 -1684
rect 870 -1771 871 -1693
rect 912 -1694 913 -1684
rect 975 -1694 976 -1684
rect 23 -1771 24 -1695
rect 222 -1696 223 -1684
rect 240 -1696 241 -1684
rect 411 -1771 412 -1695
rect 415 -1696 416 -1684
rect 436 -1771 437 -1695
rect 457 -1696 458 -1684
rect 856 -1771 857 -1695
rect 898 -1696 899 -1684
rect 975 -1771 976 -1695
rect 30 -1698 31 -1684
rect 467 -1698 468 -1684
rect 471 -1698 472 -1684
rect 751 -1698 752 -1684
rect 793 -1698 794 -1684
rect 814 -1771 815 -1697
rect 835 -1771 836 -1697
rect 940 -1698 941 -1684
rect 30 -1771 31 -1699
rect 345 -1700 346 -1684
rect 348 -1700 349 -1684
rect 387 -1771 388 -1699
rect 394 -1771 395 -1699
rect 506 -1700 507 -1684
rect 548 -1700 549 -1684
rect 807 -1771 808 -1699
rect 849 -1700 850 -1684
rect 849 -1771 850 -1699
rect 849 -1700 850 -1684
rect 849 -1771 850 -1699
rect 898 -1771 899 -1699
rect 919 -1700 920 -1684
rect 926 -1700 927 -1684
rect 961 -1771 962 -1699
rect 37 -1702 38 -1684
rect 180 -1771 181 -1701
rect 184 -1702 185 -1684
rect 191 -1771 192 -1701
rect 205 -1702 206 -1684
rect 205 -1771 206 -1701
rect 205 -1702 206 -1684
rect 205 -1771 206 -1701
rect 222 -1771 223 -1701
rect 261 -1702 262 -1684
rect 285 -1702 286 -1684
rect 408 -1702 409 -1684
rect 467 -1771 468 -1701
rect 737 -1702 738 -1684
rect 793 -1771 794 -1701
rect 828 -1702 829 -1684
rect 863 -1702 864 -1684
rect 919 -1771 920 -1701
rect 940 -1771 941 -1701
rect 1006 -1771 1007 -1701
rect 37 -1771 38 -1703
rect 292 -1704 293 -1684
rect 299 -1704 300 -1684
rect 551 -1704 552 -1684
rect 555 -1771 556 -1703
rect 618 -1704 619 -1684
rect 639 -1704 640 -1684
rect 891 -1771 892 -1703
rect 44 -1706 45 -1684
rect 61 -1771 62 -1705
rect 65 -1706 66 -1684
rect 166 -1771 167 -1705
rect 170 -1706 171 -1684
rect 296 -1771 297 -1705
rect 317 -1706 318 -1684
rect 425 -1771 426 -1705
rect 464 -1706 465 -1684
rect 639 -1771 640 -1705
rect 688 -1706 689 -1684
rect 751 -1771 752 -1705
rect 828 -1771 829 -1705
rect 16 -1771 17 -1707
rect 464 -1771 465 -1707
rect 471 -1771 472 -1707
rect 565 -1708 566 -1684
rect 569 -1708 570 -1684
rect 688 -1771 689 -1707
rect 723 -1771 724 -1707
rect 744 -1708 745 -1684
rect 44 -1771 45 -1709
rect 404 -1771 405 -1709
rect 408 -1771 409 -1709
rect 709 -1710 710 -1684
rect 51 -1712 52 -1684
rect 383 -1712 384 -1684
rect 478 -1712 479 -1684
rect 534 -1771 535 -1711
rect 548 -1771 549 -1711
rect 576 -1712 577 -1684
rect 597 -1771 598 -1711
rect 632 -1712 633 -1684
rect 51 -1771 52 -1713
rect 93 -1771 94 -1713
rect 128 -1771 129 -1713
rect 481 -1714 482 -1684
rect 485 -1714 486 -1684
rect 989 -1771 990 -1713
rect 54 -1771 55 -1715
rect 254 -1771 255 -1715
rect 261 -1771 262 -1715
rect 324 -1716 325 -1684
rect 338 -1716 339 -1684
rect 345 -1771 346 -1715
rect 352 -1716 353 -1684
rect 380 -1716 381 -1684
rect 481 -1771 482 -1715
rect 611 -1716 612 -1684
rect 614 -1771 615 -1715
rect 709 -1771 710 -1715
rect 65 -1771 66 -1717
rect 229 -1718 230 -1684
rect 243 -1771 244 -1717
rect 268 -1718 269 -1684
rect 289 -1718 290 -1684
rect 513 -1718 514 -1684
rect 516 -1771 517 -1717
rect 737 -1771 738 -1717
rect 72 -1720 73 -1684
rect 450 -1720 451 -1684
rect 488 -1720 489 -1684
rect 527 -1720 528 -1684
rect 576 -1771 577 -1719
rect 590 -1720 591 -1684
rect 618 -1771 619 -1719
rect 758 -1771 759 -1719
rect 72 -1771 73 -1721
rect 163 -1722 164 -1684
rect 177 -1722 178 -1684
rect 429 -1771 430 -1721
rect 450 -1771 451 -1721
rect 660 -1722 661 -1684
rect 79 -1771 80 -1723
rect 121 -1724 122 -1684
rect 135 -1771 136 -1723
rect 478 -1771 479 -1723
rect 492 -1724 493 -1684
rect 954 -1724 955 -1684
rect 86 -1726 87 -1684
rect 744 -1771 745 -1725
rect 947 -1726 948 -1684
rect 954 -1771 955 -1725
rect 86 -1771 87 -1727
rect 103 -1771 104 -1727
rect 121 -1771 122 -1727
rect 142 -1728 143 -1684
rect 149 -1728 150 -1684
rect 383 -1771 384 -1727
rect 401 -1728 402 -1684
rect 527 -1771 528 -1727
rect 541 -1728 542 -1684
rect 660 -1771 661 -1727
rect 905 -1728 906 -1684
rect 947 -1771 948 -1727
rect 138 -1730 139 -1684
rect 926 -1771 927 -1729
rect 142 -1771 143 -1731
rect 303 -1732 304 -1684
rect 317 -1771 318 -1731
rect 474 -1732 475 -1684
rect 492 -1771 493 -1731
rect 894 -1732 895 -1684
rect 149 -1771 150 -1733
rect 240 -1771 241 -1733
rect 247 -1734 248 -1684
rect 558 -1734 559 -1684
rect 156 -1736 157 -1684
rect 201 -1736 202 -1684
rect 268 -1771 269 -1735
rect 324 -1771 325 -1735
rect 331 -1736 332 -1684
rect 338 -1771 339 -1735
rect 352 -1771 353 -1735
rect 453 -1736 454 -1684
rect 495 -1736 496 -1684
rect 674 -1736 675 -1684
rect 156 -1771 157 -1737
rect 226 -1738 227 -1684
rect 289 -1771 290 -1737
rect 359 -1738 360 -1684
rect 366 -1738 367 -1684
rect 653 -1738 654 -1684
rect 674 -1771 675 -1737
rect 877 -1738 878 -1684
rect 100 -1740 101 -1684
rect 359 -1771 360 -1739
rect 366 -1771 367 -1739
rect 982 -1771 983 -1739
rect 100 -1771 101 -1741
rect 170 -1771 171 -1741
rect 177 -1771 178 -1741
rect 247 -1771 248 -1741
rect 303 -1771 304 -1741
rect 310 -1742 311 -1684
rect 369 -1742 370 -1684
rect 520 -1742 521 -1684
rect 541 -1771 542 -1741
rect 905 -1771 906 -1741
rect 114 -1744 115 -1684
rect 520 -1771 521 -1743
rect 842 -1744 843 -1684
rect 877 -1771 878 -1743
rect 107 -1746 108 -1684
rect 114 -1771 115 -1745
rect 163 -1771 164 -1745
rect 313 -1771 314 -1745
rect 331 -1771 332 -1745
rect 369 -1771 370 -1745
rect 373 -1746 374 -1684
rect 415 -1771 416 -1745
rect 485 -1771 486 -1745
rect 653 -1771 654 -1745
rect 786 -1746 787 -1684
rect 842 -1771 843 -1745
rect 107 -1771 108 -1747
rect 821 -1771 822 -1747
rect 187 -1771 188 -1749
rect 863 -1771 864 -1749
rect 226 -1771 227 -1751
rect 625 -1752 626 -1684
rect 786 -1771 787 -1751
rect 933 -1752 934 -1684
rect 401 -1771 402 -1753
rect 457 -1771 458 -1753
rect 499 -1754 500 -1684
rect 506 -1771 507 -1753
rect 513 -1771 514 -1753
rect 583 -1754 584 -1684
rect 625 -1771 626 -1753
rect 667 -1754 668 -1684
rect 884 -1754 885 -1684
rect 933 -1771 934 -1753
rect 373 -1771 374 -1755
rect 499 -1771 500 -1755
rect 583 -1771 584 -1755
rect 702 -1756 703 -1684
rect 800 -1756 801 -1684
rect 884 -1771 885 -1755
rect 604 -1758 605 -1684
rect 702 -1771 703 -1757
rect 604 -1771 605 -1759
rect 646 -1760 647 -1684
rect 667 -1771 668 -1759
rect 681 -1760 682 -1684
rect 569 -1771 570 -1761
rect 646 -1771 647 -1761
rect 681 -1771 682 -1761
rect 695 -1762 696 -1684
rect 695 -1771 696 -1763
rect 765 -1764 766 -1684
rect 765 -1771 766 -1765
rect 772 -1766 773 -1684
rect 422 -1768 423 -1684
rect 772 -1771 773 -1767
rect 422 -1771 423 -1769
rect 912 -1771 913 -1769
rect 2 -1781 3 -1779
rect 187 -1781 188 -1779
rect 205 -1781 206 -1779
rect 523 -1862 524 -1780
rect 565 -1862 566 -1780
rect 947 -1781 948 -1779
rect 975 -1781 976 -1779
rect 999 -1781 1000 -1779
rect 9 -1783 10 -1779
rect 30 -1783 31 -1779
rect 37 -1783 38 -1779
rect 310 -1783 311 -1779
rect 313 -1783 314 -1779
rect 499 -1783 500 -1779
rect 506 -1783 507 -1779
rect 516 -1783 517 -1779
rect 583 -1783 584 -1779
rect 583 -1862 584 -1782
rect 583 -1783 584 -1779
rect 583 -1862 584 -1782
rect 590 -1783 591 -1779
rect 961 -1783 962 -1779
rect 996 -1783 997 -1779
rect 1010 -1783 1011 -1779
rect 23 -1785 24 -1779
rect 212 -1862 213 -1784
rect 215 -1785 216 -1779
rect 296 -1785 297 -1779
rect 310 -1862 311 -1784
rect 457 -1785 458 -1779
rect 460 -1862 461 -1784
rect 919 -1785 920 -1779
rect 947 -1862 948 -1784
rect 1024 -1785 1025 -1779
rect 44 -1787 45 -1779
rect 366 -1787 367 -1779
rect 369 -1787 370 -1779
rect 394 -1787 395 -1779
rect 422 -1862 423 -1786
rect 702 -1787 703 -1779
rect 726 -1862 727 -1786
rect 954 -1787 955 -1779
rect 51 -1789 52 -1779
rect 891 -1789 892 -1779
rect 915 -1862 916 -1788
rect 933 -1789 934 -1779
rect 51 -1862 52 -1790
rect 348 -1862 349 -1790
rect 369 -1862 370 -1790
rect 387 -1791 388 -1779
rect 450 -1791 451 -1779
rect 541 -1791 542 -1779
rect 590 -1862 591 -1790
rect 604 -1791 605 -1779
rect 611 -1791 612 -1779
rect 856 -1791 857 -1779
rect 54 -1793 55 -1779
rect 72 -1793 73 -1779
rect 79 -1793 80 -1779
rect 103 -1793 104 -1779
rect 107 -1862 108 -1792
rect 191 -1793 192 -1779
rect 215 -1862 216 -1792
rect 656 -1793 657 -1779
rect 674 -1793 675 -1779
rect 814 -1793 815 -1779
rect 842 -1793 843 -1779
rect 852 -1862 853 -1792
rect 58 -1862 59 -1794
rect 121 -1795 122 -1779
rect 128 -1795 129 -1779
rect 149 -1795 150 -1779
rect 177 -1795 178 -1779
rect 229 -1862 230 -1794
rect 240 -1795 241 -1779
rect 527 -1795 528 -1779
rect 541 -1862 542 -1794
rect 628 -1862 629 -1794
rect 632 -1795 633 -1779
rect 926 -1795 927 -1779
rect 65 -1797 66 -1779
rect 327 -1797 328 -1779
rect 380 -1797 381 -1779
rect 639 -1797 640 -1779
rect 642 -1862 643 -1796
rect 989 -1797 990 -1779
rect 65 -1862 66 -1798
rect 142 -1799 143 -1779
rect 149 -1862 150 -1798
rect 156 -1799 157 -1779
rect 170 -1799 171 -1779
rect 177 -1862 178 -1798
rect 226 -1799 227 -1779
rect 401 -1799 402 -1779
rect 415 -1799 416 -1779
rect 450 -1862 451 -1798
rect 464 -1799 465 -1779
rect 548 -1799 549 -1779
rect 604 -1862 605 -1798
rect 744 -1799 745 -1779
rect 814 -1862 815 -1798
rect 898 -1799 899 -1779
rect 72 -1862 73 -1800
rect 415 -1862 416 -1800
rect 464 -1862 465 -1800
rect 562 -1801 563 -1779
rect 611 -1862 612 -1800
rect 765 -1801 766 -1779
rect 898 -1862 899 -1800
rect 950 -1862 951 -1800
rect 79 -1862 80 -1802
rect 593 -1803 594 -1779
rect 618 -1803 619 -1779
rect 751 -1803 752 -1779
rect 93 -1805 94 -1779
rect 128 -1862 129 -1804
rect 135 -1805 136 -1779
rect 184 -1862 185 -1804
rect 226 -1862 227 -1804
rect 551 -1862 552 -1804
rect 618 -1862 619 -1804
rect 723 -1805 724 -1779
rect 751 -1862 752 -1804
rect 849 -1805 850 -1779
rect 93 -1862 94 -1806
rect 114 -1807 115 -1779
rect 121 -1862 122 -1806
rect 425 -1862 426 -1806
rect 467 -1807 468 -1779
rect 513 -1862 514 -1806
rect 527 -1862 528 -1806
rect 982 -1807 983 -1779
rect 100 -1809 101 -1779
rect 401 -1862 402 -1808
rect 478 -1862 479 -1808
rect 534 -1809 535 -1779
rect 548 -1862 549 -1808
rect 765 -1862 766 -1808
rect 100 -1862 101 -1810
rect 198 -1811 199 -1779
rect 243 -1811 244 -1779
rect 387 -1862 388 -1810
rect 499 -1862 500 -1810
rect 625 -1811 626 -1779
rect 635 -1811 636 -1779
rect 828 -1811 829 -1779
rect 110 -1813 111 -1779
rect 492 -1813 493 -1779
rect 506 -1862 507 -1812
rect 772 -1813 773 -1779
rect 828 -1862 829 -1812
rect 835 -1813 836 -1779
rect 86 -1815 87 -1779
rect 492 -1862 493 -1814
rect 534 -1862 535 -1814
rect 555 -1815 556 -1779
rect 576 -1815 577 -1779
rect 835 -1862 836 -1814
rect 86 -1862 87 -1816
rect 201 -1862 202 -1816
rect 254 -1817 255 -1779
rect 562 -1862 563 -1816
rect 576 -1862 577 -1816
rect 597 -1817 598 -1779
rect 621 -1817 622 -1779
rect 744 -1862 745 -1816
rect 114 -1862 115 -1818
rect 443 -1819 444 -1779
rect 555 -1862 556 -1818
rect 667 -1819 668 -1779
rect 674 -1862 675 -1818
rect 716 -1819 717 -1779
rect 135 -1862 136 -1820
rect 163 -1862 164 -1820
rect 170 -1862 171 -1820
rect 457 -1862 458 -1820
rect 646 -1821 647 -1779
rect 856 -1862 857 -1820
rect 142 -1862 143 -1822
rect 303 -1823 304 -1779
rect 380 -1862 381 -1822
rect 520 -1823 521 -1779
rect 653 -1823 654 -1779
rect 870 -1823 871 -1779
rect 156 -1862 157 -1824
rect 219 -1825 220 -1779
rect 247 -1825 248 -1779
rect 303 -1862 304 -1824
rect 418 -1862 419 -1824
rect 646 -1862 647 -1824
rect 653 -1862 654 -1824
rect 730 -1825 731 -1779
rect 194 -1862 195 -1826
rect 219 -1862 220 -1826
rect 247 -1862 248 -1826
rect 275 -1827 276 -1779
rect 282 -1827 283 -1779
rect 394 -1862 395 -1826
rect 443 -1862 444 -1826
rect 688 -1827 689 -1779
rect 702 -1862 703 -1826
rect 1017 -1827 1018 -1779
rect 254 -1862 255 -1828
rect 324 -1829 325 -1779
rect 520 -1862 521 -1828
rect 877 -1829 878 -1779
rect 268 -1831 269 -1779
rect 373 -1831 374 -1779
rect 660 -1831 661 -1779
rect 772 -1862 773 -1830
rect 786 -1831 787 -1779
rect 877 -1862 878 -1830
rect 261 -1833 262 -1779
rect 268 -1862 269 -1832
rect 275 -1862 276 -1832
rect 677 -1833 678 -1779
rect 681 -1833 682 -1779
rect 800 -1862 801 -1832
rect 233 -1835 234 -1779
rect 261 -1862 262 -1834
rect 282 -1862 283 -1834
rect 338 -1835 339 -1779
rect 373 -1862 374 -1834
rect 408 -1835 409 -1779
rect 597 -1862 598 -1834
rect 660 -1862 661 -1834
rect 667 -1862 668 -1834
rect 940 -1835 941 -1779
rect 233 -1862 234 -1836
rect 352 -1837 353 -1779
rect 408 -1862 409 -1836
rect 849 -1862 850 -1836
rect 289 -1839 290 -1779
rect 352 -1862 353 -1838
rect 681 -1862 682 -1838
rect 695 -1839 696 -1779
rect 709 -1839 710 -1779
rect 870 -1862 871 -1838
rect 289 -1862 290 -1840
rect 331 -1841 332 -1779
rect 338 -1862 339 -1840
rect 485 -1841 486 -1779
rect 688 -1862 689 -1840
rect 779 -1841 780 -1779
rect 786 -1862 787 -1840
rect 863 -1841 864 -1779
rect 296 -1862 297 -1842
rect 376 -1843 377 -1779
rect 695 -1862 696 -1842
rect 793 -1843 794 -1779
rect 838 -1862 839 -1842
rect 863 -1862 864 -1842
rect 317 -1845 318 -1779
rect 485 -1862 486 -1844
rect 709 -1862 710 -1844
rect 758 -1845 759 -1779
rect 793 -1862 794 -1844
rect 842 -1862 843 -1844
rect 317 -1862 318 -1846
rect 345 -1847 346 -1779
rect 716 -1862 717 -1846
rect 807 -1847 808 -1779
rect 324 -1862 325 -1848
rect 436 -1849 437 -1779
rect 730 -1862 731 -1848
rect 821 -1849 822 -1779
rect 331 -1862 332 -1850
rect 569 -1851 570 -1779
rect 737 -1851 738 -1779
rect 779 -1862 780 -1850
rect 807 -1862 808 -1850
rect 968 -1851 969 -1779
rect 345 -1862 346 -1852
rect 1003 -1853 1004 -1779
rect 429 -1855 430 -1779
rect 436 -1862 437 -1854
rect 569 -1862 570 -1854
rect 884 -1855 885 -1779
rect 429 -1862 430 -1856
rect 471 -1857 472 -1779
rect 737 -1862 738 -1856
rect 912 -1857 913 -1779
rect 359 -1859 360 -1779
rect 471 -1862 472 -1858
rect 758 -1862 759 -1858
rect 845 -1862 846 -1858
rect 821 -1862 822 -1860
rect 905 -1861 906 -1779
rect 16 -1933 17 -1871
rect 51 -1872 52 -1870
rect 58 -1872 59 -1870
rect 163 -1872 164 -1870
rect 184 -1872 185 -1870
rect 198 -1872 199 -1870
rect 219 -1872 220 -1870
rect 261 -1872 262 -1870
rect 285 -1933 286 -1871
rect 870 -1872 871 -1870
rect 23 -1933 24 -1873
rect 184 -1933 185 -1873
rect 194 -1933 195 -1873
rect 198 -1933 199 -1873
rect 229 -1874 230 -1870
rect 240 -1874 241 -1870
rect 243 -1874 244 -1870
rect 317 -1874 318 -1870
rect 324 -1874 325 -1870
rect 411 -1874 412 -1870
rect 415 -1874 416 -1870
rect 450 -1874 451 -1870
rect 464 -1874 465 -1870
rect 467 -1920 468 -1873
rect 509 -1874 510 -1870
rect 737 -1874 738 -1870
rect 744 -1874 745 -1870
rect 744 -1933 745 -1873
rect 744 -1874 745 -1870
rect 744 -1933 745 -1873
rect 765 -1874 766 -1870
rect 765 -1933 766 -1873
rect 765 -1874 766 -1870
rect 765 -1933 766 -1873
rect 782 -1933 783 -1873
rect 877 -1874 878 -1870
rect 51 -1933 52 -1875
rect 191 -1876 192 -1870
rect 247 -1876 248 -1870
rect 324 -1933 325 -1875
rect 334 -1933 335 -1875
rect 709 -1876 710 -1870
rect 845 -1876 846 -1870
rect 898 -1876 899 -1870
rect 58 -1933 59 -1877
rect 296 -1878 297 -1870
rect 345 -1878 346 -1870
rect 345 -1933 346 -1877
rect 345 -1878 346 -1870
rect 345 -1933 346 -1877
rect 348 -1878 349 -1870
rect 352 -1878 353 -1870
rect 359 -1933 360 -1877
rect 439 -1933 440 -1877
rect 443 -1878 444 -1870
rect 639 -1933 640 -1877
rect 702 -1878 703 -1870
rect 821 -1878 822 -1870
rect 65 -1880 66 -1870
rect 159 -1933 160 -1879
rect 177 -1880 178 -1870
rect 243 -1933 244 -1879
rect 247 -1933 248 -1879
rect 387 -1880 388 -1870
rect 411 -1933 412 -1879
rect 460 -1933 461 -1879
rect 464 -1933 465 -1879
rect 478 -1880 479 -1870
rect 520 -1933 521 -1879
rect 583 -1880 584 -1870
rect 618 -1880 619 -1870
rect 663 -1880 664 -1870
rect 702 -1933 703 -1879
rect 758 -1880 759 -1870
rect 821 -1933 822 -1879
rect 863 -1880 864 -1870
rect 65 -1933 66 -1881
rect 124 -1933 125 -1881
rect 128 -1933 129 -1881
rect 149 -1882 150 -1870
rect 177 -1933 178 -1881
rect 457 -1882 458 -1870
rect 471 -1882 472 -1870
rect 737 -1933 738 -1881
rect 758 -1933 759 -1881
rect 793 -1882 794 -1870
rect 72 -1884 73 -1870
rect 240 -1933 241 -1883
rect 296 -1933 297 -1883
rect 401 -1884 402 -1870
rect 418 -1884 419 -1870
rect 618 -1933 619 -1883
rect 628 -1884 629 -1870
rect 674 -1884 675 -1870
rect 709 -1933 710 -1883
rect 761 -1933 762 -1883
rect 793 -1933 794 -1883
rect 856 -1884 857 -1870
rect 72 -1933 73 -1885
rect 145 -1933 146 -1885
rect 191 -1933 192 -1885
rect 275 -1886 276 -1870
rect 338 -1886 339 -1870
rect 352 -1933 353 -1885
rect 362 -1886 363 -1870
rect 485 -1886 486 -1870
rect 527 -1933 528 -1885
rect 814 -1886 815 -1870
rect 79 -1888 80 -1870
rect 229 -1933 230 -1887
rect 289 -1888 290 -1870
rect 338 -1933 339 -1887
rect 366 -1933 367 -1887
rect 523 -1888 524 -1870
rect 530 -1888 531 -1870
rect 597 -1888 598 -1870
rect 632 -1888 633 -1870
rect 786 -1888 787 -1870
rect 814 -1933 815 -1887
rect 828 -1888 829 -1870
rect 79 -1933 80 -1889
rect 282 -1890 283 -1870
rect 289 -1933 290 -1889
rect 317 -1933 318 -1889
rect 373 -1890 374 -1870
rect 632 -1933 633 -1889
rect 674 -1933 675 -1889
rect 716 -1890 717 -1870
rect 751 -1890 752 -1870
rect 786 -1933 787 -1889
rect 44 -1933 45 -1891
rect 282 -1933 283 -1891
rect 310 -1892 311 -1870
rect 373 -1933 374 -1891
rect 387 -1933 388 -1891
rect 450 -1933 451 -1891
rect 471 -1933 472 -1891
rect 772 -1892 773 -1870
rect 100 -1894 101 -1870
rect 261 -1933 262 -1893
rect 394 -1894 395 -1870
rect 401 -1933 402 -1893
rect 408 -1894 409 -1870
rect 597 -1933 598 -1893
rect 646 -1894 647 -1870
rect 716 -1933 717 -1893
rect 751 -1933 752 -1893
rect 779 -1894 780 -1870
rect 100 -1933 101 -1895
rect 114 -1896 115 -1870
rect 121 -1896 122 -1870
rect 163 -1933 164 -1895
rect 215 -1896 216 -1870
rect 418 -1933 419 -1895
rect 422 -1896 423 -1870
rect 642 -1896 643 -1870
rect 646 -1933 647 -1895
rect 688 -1896 689 -1870
rect 86 -1898 87 -1870
rect 121 -1933 122 -1897
rect 142 -1898 143 -1870
rect 275 -1933 276 -1897
rect 408 -1933 409 -1897
rect 667 -1898 668 -1870
rect 681 -1898 682 -1870
rect 688 -1933 689 -1897
rect 86 -1933 87 -1899
rect 233 -1900 234 -1870
rect 380 -1900 381 -1870
rect 667 -1933 668 -1899
rect 681 -1933 682 -1899
rect 772 -1933 773 -1899
rect 93 -1902 94 -1870
rect 142 -1933 143 -1901
rect 212 -1902 213 -1870
rect 380 -1933 381 -1901
rect 422 -1933 423 -1901
rect 723 -1902 724 -1870
rect 93 -1933 94 -1903
rect 331 -1904 332 -1870
rect 429 -1904 430 -1870
rect 443 -1933 444 -1903
rect 478 -1933 479 -1903
rect 492 -1904 493 -1870
rect 548 -1904 549 -1870
rect 726 -1904 727 -1870
rect 107 -1906 108 -1870
rect 205 -1906 206 -1870
rect 212 -1933 213 -1905
rect 268 -1906 269 -1870
rect 310 -1933 311 -1905
rect 331 -1933 332 -1905
rect 429 -1933 430 -1905
rect 513 -1906 514 -1870
rect 548 -1933 549 -1905
rect 604 -1906 605 -1870
rect 625 -1906 626 -1870
rect 723 -1933 724 -1905
rect 107 -1933 108 -1907
rect 135 -1908 136 -1870
rect 166 -1908 167 -1870
rect 205 -1933 206 -1907
rect 268 -1933 269 -1907
rect 303 -1908 304 -1870
rect 436 -1908 437 -1870
rect 436 -1933 437 -1907
rect 436 -1908 437 -1870
rect 436 -1933 437 -1907
rect 457 -1933 458 -1907
rect 513 -1933 514 -1907
rect 551 -1908 552 -1870
rect 800 -1908 801 -1870
rect 114 -1933 115 -1909
rect 156 -1910 157 -1870
rect 254 -1910 255 -1870
rect 303 -1933 304 -1909
rect 485 -1933 486 -1909
rect 506 -1910 507 -1870
rect 583 -1933 584 -1909
rect 660 -1910 661 -1870
rect 135 -1933 136 -1911
rect 170 -1912 171 -1870
rect 254 -1933 255 -1911
rect 569 -1912 570 -1870
rect 604 -1933 605 -1911
rect 807 -1912 808 -1870
rect 131 -1914 132 -1870
rect 170 -1933 171 -1913
rect 492 -1933 493 -1913
rect 499 -1914 500 -1870
rect 506 -1933 507 -1913
rect 541 -1914 542 -1870
rect 562 -1914 563 -1870
rect 660 -1933 661 -1913
rect 149 -1933 150 -1915
rect 156 -1933 157 -1915
rect 394 -1933 395 -1915
rect 562 -1933 563 -1915
rect 625 -1933 626 -1915
rect 695 -1916 696 -1870
rect 499 -1933 500 -1917
rect 576 -1918 577 -1870
rect 653 -1918 654 -1870
rect 695 -1933 696 -1917
rect 576 -1933 577 -1919
rect 611 -1920 612 -1870
rect 653 -1933 654 -1919
rect 453 -1933 454 -1921
rect 611 -1933 612 -1921
rect 534 -1924 535 -1870
rect 569 -1933 570 -1923
rect 534 -1933 535 -1925
rect 590 -1926 591 -1870
rect 541 -1933 542 -1927
rect 555 -1928 556 -1870
rect 555 -1933 556 -1929
rect 730 -1930 731 -1870
rect 730 -1933 731 -1931
rect 817 -1932 818 -1870
rect 33 -1943 34 -1941
rect 37 -1943 38 -1941
rect 40 -1943 41 -1941
rect 47 -1943 48 -1941
rect 51 -1943 52 -1941
rect 394 -1943 395 -1941
rect 418 -1943 419 -1941
rect 667 -1943 668 -1941
rect 677 -1992 678 -1942
rect 688 -1943 689 -1941
rect 695 -1943 696 -1941
rect 800 -1992 801 -1942
rect 814 -1943 815 -1941
rect 814 -1992 815 -1942
rect 814 -1943 815 -1941
rect 814 -1992 815 -1942
rect 37 -1992 38 -1944
rect 114 -1945 115 -1941
rect 121 -1992 122 -1944
rect 177 -1945 178 -1941
rect 191 -1945 192 -1941
rect 548 -1945 549 -1941
rect 576 -1945 577 -1941
rect 730 -1945 731 -1941
rect 782 -1945 783 -1941
rect 821 -1945 822 -1941
rect 44 -1992 45 -1946
rect 135 -1947 136 -1941
rect 138 -1992 139 -1946
rect 264 -1992 265 -1946
rect 275 -1947 276 -1941
rect 331 -1947 332 -1941
rect 373 -1947 374 -1941
rect 411 -1947 412 -1941
rect 446 -1992 447 -1946
rect 492 -1947 493 -1941
rect 495 -1992 496 -1946
rect 541 -1947 542 -1941
rect 593 -1947 594 -1941
rect 625 -1947 626 -1941
rect 653 -1947 654 -1941
rect 758 -1947 759 -1941
rect 786 -1947 787 -1941
rect 807 -1992 808 -1946
rect 58 -1949 59 -1941
rect 236 -1949 237 -1941
rect 243 -1949 244 -1941
rect 387 -1949 388 -1941
rect 394 -1992 395 -1948
rect 779 -1949 780 -1941
rect 72 -1951 73 -1941
rect 75 -1955 76 -1950
rect 93 -1951 94 -1941
rect 432 -1992 433 -1950
rect 439 -1951 440 -1941
rect 625 -1992 626 -1950
rect 653 -1992 654 -1950
rect 674 -1951 675 -1941
rect 684 -1951 685 -1941
rect 751 -1951 752 -1941
rect 772 -1951 773 -1941
rect 779 -1992 780 -1950
rect 72 -1992 73 -1952
rect 107 -1953 108 -1941
rect 114 -1992 115 -1952
rect 142 -1953 143 -1941
rect 170 -1953 171 -1941
rect 177 -1992 178 -1952
rect 219 -1953 220 -1941
rect 289 -1953 290 -1941
rect 296 -1953 297 -1941
rect 604 -1953 605 -1941
rect 611 -1953 612 -1941
rect 751 -1992 752 -1952
rect 107 -1992 108 -1954
rect 128 -1955 129 -1941
rect 184 -1955 185 -1941
rect 229 -1955 230 -1941
rect 261 -1955 262 -1941
rect 275 -1992 276 -1954
rect 334 -1955 335 -1941
rect 352 -1955 353 -1941
rect 387 -1992 388 -1954
rect 439 -1992 440 -1954
rect 464 -1955 465 -1941
rect 499 -1955 500 -1941
rect 695 -1992 696 -1954
rect 709 -1955 710 -1941
rect 786 -1992 787 -1954
rect 51 -1992 52 -1956
rect 229 -1992 230 -1956
rect 233 -1957 234 -1941
rect 268 -1957 269 -1941
rect 296 -1992 297 -1956
rect 474 -1957 475 -1941
rect 478 -1957 479 -1941
rect 499 -1992 500 -1956
rect 506 -1957 507 -1941
rect 548 -1992 549 -1956
rect 583 -1957 584 -1941
rect 611 -1992 612 -1956
rect 618 -1957 619 -1941
rect 758 -1992 759 -1956
rect 58 -1992 59 -1958
rect 128 -1992 129 -1958
rect 142 -1992 143 -1958
rect 194 -1959 195 -1941
rect 205 -1959 206 -1941
rect 261 -1992 262 -1958
rect 317 -1959 318 -1941
rect 464 -1992 465 -1958
rect 506 -1992 507 -1958
rect 513 -1959 514 -1941
rect 516 -1992 517 -1958
rect 772 -1992 773 -1958
rect 86 -1961 87 -1941
rect 219 -1992 220 -1960
rect 254 -1961 255 -1941
rect 331 -1992 332 -1960
rect 352 -1992 353 -1960
rect 408 -1961 409 -1941
rect 415 -1961 416 -1941
rect 709 -1992 710 -1960
rect 86 -1992 87 -1962
rect 282 -1963 283 -1941
rect 317 -1992 318 -1962
rect 345 -1963 346 -1941
rect 359 -1963 360 -1941
rect 373 -1992 374 -1962
rect 408 -1992 409 -1962
rect 422 -1963 423 -1941
rect 450 -1963 451 -1941
rect 555 -1963 556 -1941
rect 579 -1963 580 -1941
rect 618 -1992 619 -1962
rect 660 -1963 661 -1941
rect 667 -1992 668 -1962
rect 688 -1992 689 -1962
rect 765 -1963 766 -1941
rect 93 -1992 94 -1964
rect 180 -1965 181 -1941
rect 184 -1992 185 -1964
rect 310 -1965 311 -1941
rect 320 -1965 321 -1941
rect 401 -1965 402 -1941
rect 415 -1992 416 -1964
rect 460 -1965 461 -1941
rect 527 -1965 528 -1941
rect 541 -1992 542 -1964
rect 555 -1992 556 -1964
rect 562 -1965 563 -1941
rect 593 -1992 594 -1964
rect 730 -1992 731 -1964
rect 744 -1965 745 -1941
rect 765 -1992 766 -1964
rect 100 -1967 101 -1941
rect 156 -1992 157 -1966
rect 163 -1967 164 -1941
rect 170 -1992 171 -1966
rect 205 -1992 206 -1966
rect 226 -1967 227 -1941
rect 247 -1967 248 -1941
rect 254 -1992 255 -1966
rect 271 -1992 272 -1966
rect 450 -1992 451 -1966
rect 453 -1967 454 -1941
rect 737 -1967 738 -1941
rect 100 -1992 101 -1968
rect 135 -1992 136 -1968
rect 149 -1969 150 -1941
rect 268 -1992 269 -1968
rect 282 -1992 283 -1968
rect 492 -1992 493 -1968
rect 527 -1992 528 -1968
rect 726 -1992 727 -1968
rect 149 -1992 150 -1970
rect 222 -1971 223 -1941
rect 303 -1971 304 -1941
rect 359 -1992 360 -1970
rect 366 -1971 367 -1941
rect 478 -1992 479 -1970
rect 534 -1971 535 -1941
rect 590 -1971 591 -1941
rect 597 -1971 598 -1941
rect 604 -1992 605 -1970
rect 723 -1971 724 -1941
rect 737 -1992 738 -1970
rect 159 -1973 160 -1941
rect 303 -1992 304 -1972
rect 324 -1973 325 -1941
rect 345 -1992 346 -1972
rect 369 -1992 370 -1972
rect 534 -1992 535 -1972
rect 562 -1992 563 -1972
rect 639 -1973 640 -1941
rect 723 -1992 724 -1972
rect 793 -1973 794 -1941
rect 79 -1975 80 -1941
rect 324 -1992 325 -1974
rect 401 -1992 402 -1974
rect 485 -1975 486 -1941
rect 576 -1992 577 -1974
rect 744 -1992 745 -1974
rect 65 -1977 66 -1941
rect 79 -1992 80 -1976
rect 159 -1992 160 -1976
rect 163 -1992 164 -1976
rect 198 -1977 199 -1941
rect 247 -1992 248 -1976
rect 422 -1992 423 -1976
rect 502 -1977 503 -1941
rect 597 -1992 598 -1976
rect 646 -1977 647 -1941
rect 16 -1979 17 -1941
rect 65 -1992 66 -1978
rect 191 -1992 192 -1978
rect 198 -1992 199 -1978
rect 212 -1979 213 -1941
rect 233 -1992 234 -1978
rect 443 -1979 444 -1941
rect 485 -1992 486 -1978
rect 632 -1979 633 -1941
rect 639 -1992 640 -1978
rect 646 -1992 647 -1978
rect 674 -1992 675 -1978
rect 212 -1992 213 -1980
rect 240 -1981 241 -1941
rect 457 -1981 458 -1941
rect 520 -1981 521 -1941
rect 569 -1981 570 -1941
rect 632 -1992 633 -1980
rect 338 -1983 339 -1941
rect 457 -1992 458 -1982
rect 520 -1992 521 -1982
rect 681 -1983 682 -1941
rect 338 -1992 339 -1984
rect 380 -1985 381 -1941
rect 429 -1985 430 -1941
rect 569 -1992 570 -1984
rect 681 -1992 682 -1984
rect 702 -1985 703 -1941
rect 380 -1992 381 -1986
rect 471 -1992 472 -1986
rect 702 -1992 703 -1986
rect 716 -1987 717 -1941
rect 436 -1989 437 -1941
rect 716 -1992 717 -1988
rect 23 -1991 24 -1941
rect 436 -1992 437 -1990
rect 16 -2055 17 -2001
rect 93 -2002 94 -2000
rect 156 -2055 157 -2001
rect 187 -2055 188 -2001
rect 201 -2002 202 -2000
rect 226 -2055 227 -2001
rect 229 -2002 230 -2000
rect 338 -2002 339 -2000
rect 387 -2002 388 -2000
rect 404 -2055 405 -2001
rect 432 -2002 433 -2000
rect 569 -2002 570 -2000
rect 576 -2002 577 -2000
rect 576 -2055 577 -2001
rect 576 -2002 577 -2000
rect 576 -2055 577 -2001
rect 586 -2002 587 -2000
rect 639 -2002 640 -2000
rect 646 -2002 647 -2000
rect 663 -2002 664 -2000
rect 670 -2055 671 -2001
rect 786 -2002 787 -2000
rect 796 -2002 797 -2000
rect 814 -2002 815 -2000
rect 30 -2055 31 -2003
rect 79 -2004 80 -2000
rect 177 -2004 178 -2000
rect 310 -2055 311 -2003
rect 313 -2004 314 -2000
rect 324 -2004 325 -2000
rect 331 -2004 332 -2000
rect 397 -2055 398 -2003
rect 488 -2055 489 -2003
rect 513 -2004 514 -2000
rect 548 -2004 549 -2000
rect 779 -2055 780 -2003
rect 37 -2006 38 -2000
rect 149 -2006 150 -2000
rect 229 -2055 230 -2005
rect 268 -2055 269 -2005
rect 271 -2006 272 -2000
rect 359 -2006 360 -2000
rect 387 -2055 388 -2005
rect 492 -2006 493 -2000
rect 513 -2055 514 -2005
rect 632 -2006 633 -2000
rect 639 -2055 640 -2005
rect 695 -2006 696 -2000
rect 744 -2006 745 -2000
rect 807 -2006 808 -2000
rect 37 -2055 38 -2007
rect 184 -2008 185 -2000
rect 233 -2008 234 -2000
rect 240 -2008 241 -2000
rect 247 -2008 248 -2000
rect 380 -2008 381 -2000
rect 492 -2055 493 -2007
rect 555 -2008 556 -2000
rect 569 -2055 570 -2007
rect 793 -2008 794 -2000
rect 44 -2010 45 -2000
rect 198 -2010 199 -2000
rect 236 -2055 237 -2009
rect 548 -2055 549 -2009
rect 555 -2055 556 -2009
rect 618 -2010 619 -2000
rect 625 -2010 626 -2000
rect 625 -2055 626 -2009
rect 625 -2010 626 -2000
rect 625 -2055 626 -2009
rect 660 -2010 661 -2000
rect 702 -2010 703 -2000
rect 744 -2055 745 -2009
rect 751 -2010 752 -2000
rect 758 -2010 759 -2000
rect 786 -2055 787 -2009
rect 44 -2055 45 -2011
rect 107 -2012 108 -2000
rect 149 -2055 150 -2011
rect 170 -2012 171 -2000
rect 191 -2012 192 -2000
rect 198 -2055 199 -2011
rect 247 -2055 248 -2011
rect 254 -2012 255 -2000
rect 264 -2012 265 -2000
rect 632 -2055 633 -2011
rect 653 -2012 654 -2000
rect 660 -2055 661 -2011
rect 674 -2012 675 -2000
rect 695 -2055 696 -2011
rect 751 -2055 752 -2011
rect 772 -2012 773 -2000
rect 51 -2014 52 -2000
rect 166 -2055 167 -2013
rect 170 -2055 171 -2013
rect 257 -2055 258 -2013
rect 275 -2014 276 -2000
rect 275 -2055 276 -2013
rect 275 -2014 276 -2000
rect 275 -2055 276 -2013
rect 289 -2014 290 -2000
rect 352 -2014 353 -2000
rect 359 -2055 360 -2013
rect 373 -2014 374 -2000
rect 380 -2055 381 -2013
rect 408 -2014 409 -2000
rect 464 -2014 465 -2000
rect 674 -2055 675 -2013
rect 688 -2055 689 -2013
rect 730 -2014 731 -2000
rect 758 -2055 759 -2013
rect 765 -2014 766 -2000
rect 51 -2055 52 -2015
rect 590 -2016 591 -2000
rect 593 -2016 594 -2000
rect 800 -2016 801 -2000
rect 58 -2018 59 -2000
rect 243 -2018 244 -2000
rect 289 -2055 290 -2017
rect 348 -2055 349 -2017
rect 352 -2055 353 -2017
rect 422 -2018 423 -2000
rect 464 -2055 465 -2017
rect 478 -2018 479 -2000
rect 562 -2018 563 -2000
rect 618 -2055 619 -2017
rect 691 -2018 692 -2000
rect 737 -2018 738 -2000
rect 58 -2055 59 -2019
rect 114 -2020 115 -2000
rect 191 -2055 192 -2019
rect 212 -2020 213 -2000
rect 243 -2055 244 -2019
rect 282 -2020 283 -2000
rect 292 -2020 293 -2000
rect 432 -2055 433 -2019
rect 471 -2020 472 -2000
rect 702 -2055 703 -2019
rect 716 -2020 717 -2000
rect 730 -2055 731 -2019
rect 65 -2022 66 -2000
rect 233 -2055 234 -2021
rect 296 -2022 297 -2000
rect 366 -2055 367 -2021
rect 373 -2055 374 -2021
rect 450 -2022 451 -2000
rect 565 -2055 566 -2021
rect 737 -2055 738 -2021
rect 65 -2055 66 -2023
rect 460 -2055 461 -2023
rect 583 -2024 584 -2000
rect 653 -2055 654 -2023
rect 709 -2024 710 -2000
rect 716 -2055 717 -2023
rect 72 -2026 73 -2000
rect 135 -2026 136 -2000
rect 163 -2026 164 -2000
rect 296 -2055 297 -2025
rect 303 -2026 304 -2000
rect 436 -2055 437 -2025
rect 450 -2055 451 -2025
rect 597 -2026 598 -2000
rect 681 -2026 682 -2000
rect 709 -2055 710 -2025
rect 72 -2055 73 -2027
rect 100 -2028 101 -2000
rect 107 -2055 108 -2027
rect 254 -2055 255 -2027
rect 303 -2055 304 -2027
rect 474 -2055 475 -2027
rect 541 -2028 542 -2000
rect 597 -2055 598 -2027
rect 667 -2028 668 -2000
rect 681 -2055 682 -2027
rect 79 -2055 80 -2029
rect 317 -2030 318 -2000
rect 324 -2055 325 -2029
rect 394 -2030 395 -2000
rect 401 -2030 402 -2000
rect 765 -2055 766 -2029
rect 86 -2032 87 -2000
rect 135 -2055 136 -2031
rect 219 -2032 220 -2000
rect 282 -2055 283 -2031
rect 317 -2055 318 -2031
rect 457 -2032 458 -2000
rect 527 -2032 528 -2000
rect 541 -2055 542 -2031
rect 583 -2055 584 -2031
rect 611 -2032 612 -2000
rect 646 -2055 647 -2031
rect 667 -2055 668 -2031
rect 86 -2055 87 -2033
rect 520 -2034 521 -2000
rect 590 -2055 591 -2033
rect 726 -2055 727 -2033
rect 100 -2055 101 -2035
rect 121 -2036 122 -2000
rect 128 -2036 129 -2000
rect 212 -2055 213 -2035
rect 261 -2036 262 -2000
rect 527 -2055 528 -2035
rect 611 -2055 612 -2035
rect 677 -2036 678 -2000
rect 23 -2055 24 -2037
rect 128 -2055 129 -2037
rect 205 -2038 206 -2000
rect 219 -2055 220 -2037
rect 261 -2055 262 -2037
rect 345 -2038 346 -2000
rect 394 -2055 395 -2037
rect 772 -2055 773 -2037
rect 114 -2055 115 -2039
rect 142 -2040 143 -2000
rect 205 -2055 206 -2039
rect 446 -2040 447 -2000
rect 457 -2055 458 -2039
rect 604 -2040 605 -2000
rect 93 -2055 94 -2041
rect 142 -2055 143 -2041
rect 331 -2055 332 -2041
rect 401 -2055 402 -2041
rect 408 -2055 409 -2041
rect 415 -2042 416 -2000
rect 418 -2055 419 -2041
rect 604 -2055 605 -2041
rect 121 -2055 122 -2043
rect 184 -2055 185 -2043
rect 338 -2055 339 -2043
rect 600 -2044 601 -2000
rect 345 -2055 346 -2045
rect 443 -2046 444 -2000
rect 506 -2046 507 -2000
rect 520 -2055 521 -2045
rect 415 -2055 416 -2047
rect 534 -2048 535 -2000
rect 422 -2055 423 -2049
rect 499 -2050 500 -2000
rect 429 -2052 430 -2000
rect 443 -2055 444 -2051
rect 478 -2055 479 -2051
rect 499 -2055 500 -2051
rect 485 -2054 486 -2000
rect 534 -2055 535 -2053
rect 23 -2065 24 -2063
rect 397 -2065 398 -2063
rect 411 -2120 412 -2064
rect 513 -2065 514 -2063
rect 534 -2065 535 -2063
rect 537 -2069 538 -2064
rect 541 -2065 542 -2063
rect 593 -2120 594 -2064
rect 611 -2065 612 -2063
rect 611 -2120 612 -2064
rect 611 -2065 612 -2063
rect 611 -2120 612 -2064
rect 653 -2120 654 -2064
rect 737 -2065 738 -2063
rect 23 -2120 24 -2066
rect 240 -2067 241 -2063
rect 254 -2067 255 -2063
rect 282 -2067 283 -2063
rect 292 -2120 293 -2066
rect 366 -2067 367 -2063
rect 373 -2067 374 -2063
rect 401 -2120 402 -2066
rect 418 -2067 419 -2063
rect 499 -2067 500 -2063
rect 534 -2120 535 -2066
rect 555 -2067 556 -2063
rect 569 -2067 570 -2063
rect 632 -2067 633 -2063
rect 667 -2120 668 -2066
rect 681 -2067 682 -2063
rect 723 -2067 724 -2063
rect 758 -2067 759 -2063
rect 30 -2069 31 -2063
rect 145 -2069 146 -2063
rect 184 -2069 185 -2063
rect 236 -2069 237 -2063
rect 240 -2120 241 -2068
rect 275 -2069 276 -2063
rect 345 -2069 346 -2063
rect 422 -2069 423 -2063
rect 436 -2069 437 -2063
rect 513 -2120 514 -2068
rect 555 -2120 556 -2068
rect 569 -2120 570 -2068
rect 583 -2069 584 -2063
rect 632 -2120 633 -2068
rect 646 -2069 647 -2063
rect 670 -2069 671 -2063
rect 786 -2069 787 -2063
rect 30 -2120 31 -2070
rect 471 -2071 472 -2063
rect 474 -2071 475 -2063
rect 618 -2071 619 -2063
rect 646 -2120 647 -2070
rect 730 -2071 731 -2063
rect 37 -2073 38 -2063
rect 229 -2073 230 -2063
rect 257 -2073 258 -2063
rect 429 -2120 430 -2072
rect 443 -2073 444 -2063
rect 443 -2120 444 -2072
rect 443 -2073 444 -2063
rect 443 -2120 444 -2072
rect 457 -2073 458 -2063
rect 779 -2073 780 -2063
rect 44 -2075 45 -2063
rect 177 -2075 178 -2063
rect 212 -2075 213 -2063
rect 282 -2120 283 -2074
rect 296 -2075 297 -2063
rect 422 -2120 423 -2074
rect 457 -2120 458 -2074
rect 583 -2120 584 -2074
rect 618 -2120 619 -2074
rect 660 -2075 661 -2063
rect 681 -2120 682 -2074
rect 772 -2075 773 -2063
rect 44 -2120 45 -2076
rect 170 -2077 171 -2063
rect 212 -2120 213 -2076
rect 348 -2120 349 -2076
rect 352 -2077 353 -2063
rect 562 -2077 563 -2063
rect 660 -2120 661 -2076
rect 674 -2077 675 -2063
rect 709 -2077 710 -2063
rect 723 -2120 724 -2076
rect 726 -2077 727 -2063
rect 737 -2120 738 -2076
rect 51 -2079 52 -2063
rect 124 -2079 125 -2063
rect 135 -2079 136 -2063
rect 177 -2120 178 -2078
rect 219 -2079 220 -2063
rect 254 -2120 255 -2078
rect 275 -2120 276 -2078
rect 310 -2079 311 -2063
rect 324 -2079 325 -2063
rect 352 -2120 353 -2078
rect 373 -2120 374 -2078
rect 485 -2079 486 -2063
rect 488 -2079 489 -2063
rect 492 -2079 493 -2063
rect 499 -2120 500 -2078
rect 590 -2079 591 -2063
rect 709 -2120 710 -2078
rect 751 -2079 752 -2063
rect 51 -2120 52 -2080
rect 149 -2081 150 -2063
rect 268 -2081 269 -2063
rect 310 -2120 311 -2080
rect 317 -2081 318 -2063
rect 324 -2120 325 -2080
rect 359 -2081 360 -2063
rect 485 -2120 486 -2080
rect 492 -2120 493 -2080
rect 548 -2081 549 -2063
rect 562 -2120 563 -2080
rect 597 -2081 598 -2063
rect 58 -2083 59 -2063
rect 131 -2083 132 -2063
rect 135 -2120 136 -2082
rect 338 -2083 339 -2063
rect 380 -2083 381 -2063
rect 415 -2083 416 -2063
rect 464 -2083 465 -2063
rect 509 -2083 510 -2063
rect 527 -2083 528 -2063
rect 674 -2120 675 -2082
rect 58 -2120 59 -2084
rect 128 -2085 129 -2063
rect 142 -2085 143 -2063
rect 362 -2120 363 -2084
rect 366 -2120 367 -2084
rect 464 -2120 465 -2084
rect 474 -2120 475 -2084
rect 576 -2085 577 -2063
rect 65 -2087 66 -2063
rect 138 -2120 139 -2086
rect 142 -2120 143 -2086
rect 156 -2087 157 -2063
rect 233 -2087 234 -2063
rect 268 -2120 269 -2086
rect 296 -2120 297 -2086
rect 331 -2087 332 -2063
rect 338 -2120 339 -2086
rect 460 -2087 461 -2063
rect 478 -2087 479 -2063
rect 702 -2087 703 -2063
rect 65 -2120 66 -2088
rect 243 -2089 244 -2063
rect 317 -2120 318 -2088
rect 597 -2120 598 -2088
rect 688 -2089 689 -2063
rect 702 -2120 703 -2088
rect 72 -2091 73 -2063
rect 103 -2120 104 -2090
rect 107 -2091 108 -2063
rect 184 -2120 185 -2090
rect 233 -2120 234 -2090
rect 289 -2091 290 -2063
rect 331 -2120 332 -2090
rect 387 -2091 388 -2063
rect 415 -2120 416 -2090
rect 450 -2091 451 -2063
rect 460 -2120 461 -2090
rect 765 -2091 766 -2063
rect 72 -2120 73 -2092
rect 261 -2093 262 -2063
rect 320 -2120 321 -2092
rect 450 -2120 451 -2092
rect 478 -2120 479 -2092
rect 516 -2093 517 -2063
rect 520 -2093 521 -2063
rect 527 -2120 528 -2092
rect 576 -2120 577 -2092
rect 625 -2093 626 -2063
rect 688 -2120 689 -2092
rect 716 -2093 717 -2063
rect 79 -2095 80 -2063
rect 439 -2120 440 -2094
rect 506 -2095 507 -2063
rect 548 -2120 549 -2094
rect 625 -2120 626 -2094
rect 639 -2095 640 -2063
rect 716 -2120 717 -2094
rect 744 -2095 745 -2063
rect 79 -2120 80 -2096
rect 173 -2120 174 -2096
rect 247 -2097 248 -2063
rect 289 -2120 290 -2096
rect 387 -2120 388 -2096
rect 506 -2120 507 -2096
rect 520 -2120 521 -2096
rect 604 -2097 605 -2063
rect 86 -2099 87 -2063
rect 187 -2099 188 -2063
rect 261 -2120 262 -2098
rect 432 -2099 433 -2063
rect 604 -2120 605 -2098
rect 695 -2099 696 -2063
rect 86 -2120 87 -2100
rect 96 -2120 97 -2100
rect 100 -2101 101 -2063
rect 107 -2120 108 -2100
rect 114 -2101 115 -2063
rect 114 -2120 115 -2100
rect 114 -2101 115 -2063
rect 114 -2120 115 -2100
rect 121 -2120 122 -2100
rect 303 -2101 304 -2063
rect 394 -2101 395 -2063
rect 639 -2120 640 -2100
rect 93 -2103 94 -2063
rect 229 -2120 230 -2102
rect 303 -2120 304 -2102
rect 383 -2120 384 -2102
rect 394 -2120 395 -2102
rect 408 -2103 409 -2063
rect 16 -2105 17 -2063
rect 93 -2120 94 -2104
rect 128 -2120 129 -2104
rect 541 -2120 542 -2104
rect 149 -2120 150 -2106
rect 191 -2107 192 -2063
rect 163 -2109 164 -2063
rect 247 -2120 248 -2108
rect 156 -2120 157 -2110
rect 163 -2120 164 -2110
rect 180 -2111 181 -2063
rect 695 -2120 696 -2110
rect 180 -2120 181 -2112
rect 198 -2113 199 -2063
rect 191 -2120 192 -2114
rect 205 -2115 206 -2063
rect 16 -2120 17 -2116
rect 205 -2120 206 -2116
rect 198 -2120 199 -2118
rect 219 -2120 220 -2118
rect 16 -2130 17 -2128
rect 474 -2130 475 -2128
rect 506 -2130 507 -2128
rect 625 -2130 626 -2128
rect 632 -2130 633 -2128
rect 632 -2171 633 -2129
rect 632 -2130 633 -2128
rect 632 -2171 633 -2129
rect 688 -2130 689 -2128
rect 698 -2171 699 -2129
rect 40 -2132 41 -2128
rect 152 -2171 153 -2131
rect 163 -2132 164 -2128
rect 173 -2132 174 -2128
rect 184 -2171 185 -2131
rect 254 -2132 255 -2128
rect 261 -2132 262 -2128
rect 453 -2171 454 -2131
rect 457 -2171 458 -2131
rect 688 -2171 689 -2131
rect 695 -2132 696 -2128
rect 730 -2132 731 -2128
rect 44 -2134 45 -2128
rect 229 -2171 230 -2133
rect 254 -2171 255 -2133
rect 338 -2134 339 -2128
rect 345 -2134 346 -2128
rect 597 -2134 598 -2128
rect 625 -2171 626 -2133
rect 709 -2134 710 -2128
rect 51 -2136 52 -2128
rect 219 -2136 220 -2128
rect 226 -2136 227 -2128
rect 240 -2136 241 -2128
rect 261 -2171 262 -2135
rect 352 -2136 353 -2128
rect 359 -2171 360 -2135
rect 429 -2136 430 -2128
rect 436 -2171 437 -2135
rect 467 -2136 468 -2128
rect 509 -2136 510 -2128
rect 541 -2136 542 -2128
rect 558 -2171 559 -2135
rect 716 -2136 717 -2128
rect 58 -2138 59 -2128
rect 100 -2138 101 -2128
rect 121 -2138 122 -2128
rect 247 -2171 248 -2137
rect 268 -2138 269 -2128
rect 345 -2171 346 -2137
rect 348 -2138 349 -2128
rect 411 -2138 412 -2128
rect 439 -2138 440 -2128
rect 611 -2138 612 -2128
rect 660 -2138 661 -2128
rect 716 -2171 717 -2137
rect 65 -2140 66 -2128
rect 320 -2140 321 -2128
rect 324 -2140 325 -2128
rect 352 -2171 353 -2139
rect 380 -2140 381 -2128
rect 394 -2140 395 -2128
rect 408 -2140 409 -2128
rect 513 -2140 514 -2128
rect 534 -2140 535 -2128
rect 709 -2171 710 -2139
rect 72 -2142 73 -2128
rect 334 -2171 335 -2141
rect 362 -2142 363 -2128
rect 380 -2171 381 -2141
rect 390 -2171 391 -2141
rect 492 -2142 493 -2128
rect 513 -2171 514 -2141
rect 520 -2142 521 -2128
rect 541 -2171 542 -2141
rect 548 -2142 549 -2128
rect 579 -2171 580 -2141
rect 702 -2142 703 -2128
rect 86 -2144 87 -2128
rect 86 -2171 87 -2143
rect 86 -2144 87 -2128
rect 86 -2171 87 -2143
rect 100 -2171 101 -2143
rect 114 -2144 115 -2128
rect 128 -2144 129 -2128
rect 156 -2144 157 -2128
rect 170 -2144 171 -2128
rect 415 -2144 416 -2128
rect 464 -2144 465 -2128
rect 562 -2144 563 -2128
rect 583 -2144 584 -2128
rect 590 -2171 591 -2143
rect 593 -2144 594 -2128
rect 695 -2171 696 -2143
rect 30 -2146 31 -2128
rect 128 -2171 129 -2145
rect 135 -2146 136 -2128
rect 163 -2171 164 -2145
rect 198 -2146 199 -2128
rect 450 -2146 451 -2128
rect 464 -2171 465 -2145
rect 499 -2146 500 -2128
rect 520 -2171 521 -2145
rect 527 -2146 528 -2128
rect 548 -2171 549 -2145
rect 569 -2146 570 -2128
rect 597 -2171 598 -2145
rect 604 -2146 605 -2128
rect 611 -2171 612 -2145
rect 653 -2146 654 -2128
rect 107 -2148 108 -2128
rect 135 -2171 136 -2147
rect 142 -2148 143 -2128
rect 159 -2148 160 -2128
rect 198 -2171 199 -2147
rect 222 -2148 223 -2128
rect 226 -2171 227 -2147
rect 268 -2171 269 -2147
rect 282 -2148 283 -2128
rect 289 -2171 290 -2147
rect 296 -2148 297 -2128
rect 338 -2171 339 -2147
rect 373 -2148 374 -2128
rect 394 -2171 395 -2147
rect 408 -2171 409 -2147
rect 534 -2171 535 -2147
rect 555 -2148 556 -2128
rect 702 -2171 703 -2147
rect 23 -2150 24 -2128
rect 159 -2171 160 -2149
rect 170 -2171 171 -2149
rect 555 -2171 556 -2149
rect 604 -2171 605 -2149
rect 618 -2150 619 -2128
rect 639 -2150 640 -2128
rect 660 -2171 661 -2149
rect 107 -2171 108 -2151
rect 177 -2152 178 -2128
rect 201 -2152 202 -2128
rect 275 -2152 276 -2128
rect 282 -2171 283 -2151
rect 324 -2171 325 -2151
rect 331 -2152 332 -2128
rect 429 -2171 430 -2151
rect 471 -2152 472 -2128
rect 562 -2171 563 -2151
rect 639 -2171 640 -2151
rect 681 -2152 682 -2128
rect 114 -2171 115 -2153
rect 285 -2171 286 -2153
rect 296 -2171 297 -2153
rect 387 -2154 388 -2128
rect 443 -2154 444 -2128
rect 471 -2171 472 -2153
rect 485 -2154 486 -2128
rect 618 -2171 619 -2153
rect 646 -2154 647 -2128
rect 653 -2171 654 -2153
rect 121 -2171 122 -2155
rect 387 -2171 388 -2155
rect 443 -2171 444 -2155
rect 478 -2156 479 -2128
rect 499 -2171 500 -2155
rect 509 -2171 510 -2155
rect 646 -2171 647 -2155
rect 674 -2156 675 -2128
rect 142 -2171 143 -2157
rect 233 -2158 234 -2128
rect 275 -2171 276 -2157
rect 303 -2158 304 -2128
rect 313 -2171 314 -2157
rect 737 -2158 738 -2128
rect 149 -2160 150 -2128
rect 205 -2160 206 -2128
rect 212 -2160 213 -2128
rect 233 -2171 234 -2159
rect 303 -2171 304 -2159
rect 310 -2160 311 -2128
rect 331 -2171 332 -2159
rect 527 -2171 528 -2159
rect 667 -2160 668 -2128
rect 674 -2171 675 -2159
rect 79 -2162 80 -2128
rect 212 -2171 213 -2161
rect 219 -2171 220 -2161
rect 415 -2171 416 -2161
rect 478 -2171 479 -2161
rect 569 -2171 570 -2161
rect 667 -2171 668 -2161
rect 723 -2162 724 -2128
rect 156 -2171 157 -2163
rect 310 -2171 311 -2163
rect 366 -2164 367 -2128
rect 485 -2171 486 -2163
rect 576 -2164 577 -2128
rect 723 -2171 724 -2163
rect 177 -2171 178 -2165
rect 180 -2166 181 -2128
rect 191 -2166 192 -2128
rect 205 -2171 206 -2165
rect 222 -2171 223 -2165
rect 317 -2171 318 -2165
rect 366 -2171 367 -2165
rect 422 -2166 423 -2128
rect 191 -2171 192 -2167
rect 208 -2168 209 -2128
rect 373 -2171 374 -2167
rect 401 -2168 402 -2128
rect 422 -2171 423 -2167
rect 576 -2171 577 -2167
rect 250 -2170 251 -2128
rect 401 -2171 402 -2169
rect 86 -2181 87 -2179
rect 89 -2224 90 -2180
rect 107 -2181 108 -2179
rect 107 -2224 108 -2180
rect 107 -2181 108 -2179
rect 107 -2224 108 -2180
rect 114 -2181 115 -2179
rect 306 -2224 307 -2180
rect 380 -2181 381 -2179
rect 492 -2181 493 -2179
rect 506 -2224 507 -2180
rect 527 -2181 528 -2179
rect 534 -2181 535 -2179
rect 670 -2181 671 -2179
rect 674 -2181 675 -2179
rect 681 -2181 682 -2179
rect 114 -2224 115 -2182
rect 184 -2183 185 -2179
rect 191 -2183 192 -2179
rect 191 -2224 192 -2182
rect 191 -2183 192 -2179
rect 191 -2224 192 -2182
rect 205 -2183 206 -2179
rect 219 -2183 220 -2179
rect 222 -2183 223 -2179
rect 576 -2183 577 -2179
rect 579 -2224 580 -2182
rect 723 -2183 724 -2179
rect 121 -2185 122 -2179
rect 149 -2224 150 -2184
rect 163 -2185 164 -2179
rect 184 -2224 185 -2184
rect 205 -2224 206 -2184
rect 299 -2185 300 -2179
rect 324 -2185 325 -2179
rect 380 -2224 381 -2184
rect 401 -2185 402 -2179
rect 460 -2185 461 -2179
rect 492 -2224 493 -2184
rect 558 -2185 559 -2179
rect 569 -2185 570 -2179
rect 716 -2185 717 -2179
rect 124 -2224 125 -2186
rect 254 -2187 255 -2179
rect 275 -2187 276 -2179
rect 275 -2224 276 -2186
rect 275 -2187 276 -2179
rect 275 -2224 276 -2186
rect 282 -2187 283 -2179
rect 366 -2187 367 -2179
rect 401 -2224 402 -2186
rect 422 -2187 423 -2179
rect 425 -2224 426 -2186
rect 562 -2187 563 -2179
rect 583 -2187 584 -2179
rect 688 -2187 689 -2179
rect 128 -2189 129 -2179
rect 411 -2189 412 -2179
rect 429 -2189 430 -2179
rect 618 -2189 619 -2179
rect 639 -2189 640 -2179
rect 667 -2189 668 -2179
rect 142 -2191 143 -2179
rect 219 -2224 220 -2190
rect 233 -2191 234 -2179
rect 233 -2224 234 -2190
rect 233 -2191 234 -2179
rect 233 -2224 234 -2190
rect 240 -2191 241 -2179
rect 513 -2191 514 -2179
rect 555 -2191 556 -2179
rect 611 -2191 612 -2179
rect 170 -2193 171 -2179
rect 240 -2224 241 -2192
rect 243 -2193 244 -2179
rect 254 -2224 255 -2192
rect 285 -2193 286 -2179
rect 390 -2193 391 -2179
rect 394 -2193 395 -2179
rect 562 -2224 563 -2192
rect 569 -2224 570 -2192
rect 618 -2224 619 -2192
rect 142 -2224 143 -2194
rect 170 -2224 171 -2194
rect 198 -2195 199 -2179
rect 394 -2224 395 -2194
rect 408 -2224 409 -2194
rect 443 -2195 444 -2179
rect 450 -2195 451 -2179
rect 464 -2195 465 -2179
rect 499 -2195 500 -2179
rect 527 -2224 528 -2194
rect 555 -2224 556 -2194
rect 632 -2195 633 -2179
rect 212 -2197 213 -2179
rect 345 -2197 346 -2179
rect 366 -2224 367 -2196
rect 373 -2197 374 -2179
rect 387 -2224 388 -2196
rect 464 -2224 465 -2196
rect 513 -2224 514 -2196
rect 548 -2197 549 -2179
rect 583 -2224 584 -2196
rect 653 -2197 654 -2179
rect 152 -2199 153 -2179
rect 212 -2224 213 -2198
rect 285 -2224 286 -2198
rect 450 -2224 451 -2198
rect 548 -2224 549 -2198
rect 590 -2199 591 -2179
rect 597 -2199 598 -2179
rect 639 -2224 640 -2198
rect 296 -2224 297 -2200
rect 614 -2224 615 -2200
rect 632 -2224 633 -2200
rect 702 -2201 703 -2179
rect 317 -2203 318 -2179
rect 345 -2224 346 -2202
rect 415 -2203 416 -2179
rect 499 -2224 500 -2202
rect 586 -2203 587 -2179
rect 604 -2203 605 -2179
rect 317 -2224 318 -2204
rect 471 -2205 472 -2179
rect 509 -2205 510 -2179
rect 604 -2224 605 -2204
rect 324 -2224 325 -2206
rect 352 -2207 353 -2179
rect 359 -2207 360 -2179
rect 415 -2224 416 -2206
rect 429 -2224 430 -2206
rect 478 -2207 479 -2179
rect 590 -2224 591 -2206
rect 625 -2207 626 -2179
rect 268 -2209 269 -2179
rect 352 -2224 353 -2208
rect 432 -2209 433 -2179
rect 457 -2224 458 -2208
rect 478 -2224 479 -2208
rect 621 -2224 622 -2208
rect 268 -2224 269 -2210
rect 310 -2211 311 -2179
rect 331 -2211 332 -2179
rect 471 -2224 472 -2210
rect 485 -2211 486 -2179
rect 625 -2224 626 -2210
rect 261 -2213 262 -2179
rect 331 -2224 332 -2212
rect 436 -2213 437 -2179
rect 534 -2224 535 -2212
rect 597 -2224 598 -2212
rect 646 -2213 647 -2179
rect 261 -2224 262 -2214
rect 338 -2215 339 -2179
rect 390 -2224 391 -2214
rect 436 -2224 437 -2214
rect 485 -2224 486 -2214
rect 520 -2215 521 -2179
rect 156 -2217 157 -2179
rect 338 -2224 339 -2216
rect 520 -2224 521 -2216
rect 541 -2217 542 -2179
rect 156 -2224 157 -2218
rect 177 -2219 178 -2179
rect 289 -2219 290 -2179
rect 310 -2224 311 -2218
rect 541 -2224 542 -2218
rect 660 -2219 661 -2179
rect 131 -2221 132 -2179
rect 177 -2224 178 -2220
rect 247 -2221 248 -2179
rect 289 -2224 290 -2220
rect 660 -2224 661 -2220
rect 709 -2221 710 -2179
rect 100 -2223 101 -2179
rect 131 -2224 132 -2222
rect 247 -2224 248 -2222
rect 303 -2223 304 -2179
rect 107 -2234 108 -2232
rect 229 -2234 230 -2232
rect 275 -2234 276 -2232
rect 282 -2234 283 -2232
rect 289 -2234 290 -2232
rect 289 -2261 290 -2233
rect 289 -2234 290 -2232
rect 289 -2261 290 -2233
rect 306 -2234 307 -2232
rect 478 -2234 479 -2232
rect 499 -2234 500 -2232
rect 499 -2261 500 -2233
rect 499 -2234 500 -2232
rect 499 -2261 500 -2233
rect 534 -2234 535 -2232
rect 611 -2234 612 -2232
rect 639 -2234 640 -2232
rect 639 -2261 640 -2233
rect 639 -2234 640 -2232
rect 639 -2261 640 -2233
rect 114 -2236 115 -2232
rect 194 -2261 195 -2235
rect 198 -2261 199 -2235
rect 236 -2261 237 -2235
rect 254 -2236 255 -2232
rect 275 -2261 276 -2235
rect 313 -2261 314 -2235
rect 401 -2236 402 -2232
rect 415 -2236 416 -2232
rect 425 -2236 426 -2232
rect 443 -2236 444 -2232
rect 478 -2261 479 -2235
rect 527 -2236 528 -2232
rect 534 -2261 535 -2235
rect 548 -2236 549 -2232
rect 548 -2261 549 -2235
rect 548 -2236 549 -2232
rect 548 -2261 549 -2235
rect 562 -2261 563 -2235
rect 590 -2236 591 -2232
rect 607 -2236 608 -2232
rect 660 -2236 661 -2232
rect 114 -2261 115 -2237
rect 142 -2238 143 -2232
rect 149 -2238 150 -2232
rect 170 -2261 171 -2237
rect 173 -2238 174 -2232
rect 191 -2238 192 -2232
rect 201 -2238 202 -2232
rect 212 -2238 213 -2232
rect 219 -2238 220 -2232
rect 254 -2261 255 -2237
rect 317 -2238 318 -2232
rect 317 -2261 318 -2237
rect 317 -2238 318 -2232
rect 317 -2261 318 -2237
rect 324 -2238 325 -2232
rect 359 -2238 360 -2232
rect 366 -2238 367 -2232
rect 376 -2238 377 -2232
rect 390 -2238 391 -2232
rect 415 -2261 416 -2237
rect 422 -2261 423 -2237
rect 429 -2238 430 -2232
rect 446 -2238 447 -2232
rect 541 -2238 542 -2232
rect 565 -2238 566 -2232
rect 632 -2238 633 -2232
rect 121 -2261 122 -2239
rect 124 -2240 125 -2232
rect 128 -2240 129 -2232
rect 138 -2240 139 -2232
rect 149 -2261 150 -2239
rect 208 -2240 209 -2232
rect 212 -2261 213 -2239
rect 219 -2261 220 -2239
rect 261 -2240 262 -2232
rect 324 -2261 325 -2239
rect 327 -2261 328 -2239
rect 362 -2261 363 -2239
rect 366 -2261 367 -2239
rect 380 -2240 381 -2232
rect 397 -2261 398 -2239
rect 471 -2240 472 -2232
rect 513 -2240 514 -2232
rect 541 -2261 542 -2239
rect 583 -2240 584 -2232
rect 583 -2261 584 -2239
rect 583 -2240 584 -2232
rect 583 -2261 584 -2239
rect 124 -2261 125 -2241
rect 145 -2261 146 -2241
rect 156 -2242 157 -2232
rect 191 -2261 192 -2241
rect 205 -2261 206 -2241
rect 306 -2261 307 -2241
rect 331 -2242 332 -2232
rect 390 -2261 391 -2241
rect 401 -2261 402 -2241
rect 408 -2242 409 -2232
rect 457 -2242 458 -2232
rect 457 -2261 458 -2241
rect 457 -2242 458 -2232
rect 457 -2261 458 -2241
rect 464 -2242 465 -2232
rect 520 -2242 521 -2232
rect 527 -2261 528 -2241
rect 555 -2242 556 -2232
rect 131 -2261 132 -2243
rect 135 -2261 136 -2243
rect 156 -2261 157 -2243
rect 177 -2244 178 -2232
rect 261 -2261 262 -2243
rect 408 -2261 409 -2243
rect 467 -2244 468 -2232
rect 506 -2244 507 -2232
rect 513 -2261 514 -2243
rect 576 -2244 577 -2232
rect 163 -2246 164 -2232
rect 268 -2246 269 -2232
rect 296 -2246 297 -2232
rect 331 -2261 332 -2245
rect 338 -2246 339 -2232
rect 565 -2261 566 -2245
rect 576 -2261 577 -2245
rect 597 -2246 598 -2232
rect 163 -2261 164 -2247
rect 180 -2248 181 -2232
rect 247 -2248 248 -2232
rect 296 -2261 297 -2247
rect 310 -2248 311 -2232
rect 338 -2261 339 -2247
rect 345 -2248 346 -2232
rect 464 -2261 465 -2247
rect 492 -2248 493 -2232
rect 520 -2261 521 -2247
rect 555 -2261 556 -2247
rect 569 -2248 570 -2232
rect 166 -2250 167 -2232
rect 432 -2261 433 -2249
rect 485 -2250 486 -2232
rect 492 -2261 493 -2249
rect 506 -2261 507 -2249
rect 579 -2250 580 -2232
rect 177 -2261 178 -2251
rect 184 -2252 185 -2232
rect 240 -2252 241 -2232
rect 247 -2261 248 -2251
rect 268 -2261 269 -2251
rect 282 -2261 283 -2251
rect 303 -2252 304 -2232
rect 345 -2261 346 -2251
rect 359 -2261 360 -2251
rect 443 -2261 444 -2251
rect 184 -2261 185 -2253
rect 240 -2261 241 -2253
rect 373 -2254 374 -2232
rect 436 -2254 437 -2232
rect 352 -2256 353 -2232
rect 373 -2261 374 -2255
rect 394 -2256 395 -2232
rect 485 -2261 486 -2255
rect 226 -2258 227 -2232
rect 352 -2261 353 -2257
rect 380 -2261 381 -2257
rect 394 -2261 395 -2257
rect 436 -2261 437 -2257
rect 450 -2258 451 -2232
rect 226 -2261 227 -2259
rect 233 -2260 234 -2232
rect 303 -2261 304 -2259
rect 450 -2261 451 -2259
rect 114 -2271 115 -2269
rect 131 -2271 132 -2269
rect 135 -2271 136 -2269
rect 145 -2271 146 -2269
rect 163 -2271 164 -2269
rect 306 -2271 307 -2269
rect 317 -2271 318 -2269
rect 373 -2271 374 -2269
rect 380 -2271 381 -2269
rect 380 -2288 381 -2270
rect 380 -2271 381 -2269
rect 380 -2288 381 -2270
rect 401 -2271 402 -2269
rect 439 -2288 440 -2270
rect 450 -2271 451 -2269
rect 572 -2288 573 -2270
rect 639 -2271 640 -2269
rect 639 -2288 640 -2270
rect 639 -2271 640 -2269
rect 639 -2288 640 -2270
rect 121 -2288 122 -2272
rect 124 -2273 125 -2269
rect 142 -2273 143 -2269
rect 156 -2273 157 -2269
rect 170 -2273 171 -2269
rect 212 -2273 213 -2269
rect 215 -2273 216 -2269
rect 222 -2288 223 -2272
rect 240 -2288 241 -2272
rect 250 -2288 251 -2272
rect 254 -2273 255 -2269
rect 254 -2288 255 -2272
rect 254 -2273 255 -2269
rect 254 -2288 255 -2272
rect 275 -2273 276 -2269
rect 282 -2273 283 -2269
rect 289 -2273 290 -2269
rect 310 -2288 311 -2272
rect 345 -2273 346 -2269
rect 345 -2288 346 -2272
rect 345 -2273 346 -2269
rect 345 -2288 346 -2272
rect 352 -2273 353 -2269
rect 387 -2273 388 -2269
rect 404 -2288 405 -2272
rect 415 -2273 416 -2269
rect 422 -2273 423 -2269
rect 422 -2288 423 -2272
rect 422 -2273 423 -2269
rect 422 -2288 423 -2272
rect 429 -2273 430 -2269
rect 530 -2288 531 -2272
rect 541 -2273 542 -2269
rect 569 -2273 570 -2269
rect 177 -2275 178 -2269
rect 177 -2288 178 -2274
rect 177 -2275 178 -2269
rect 177 -2288 178 -2274
rect 184 -2275 185 -2269
rect 233 -2275 234 -2269
rect 243 -2275 244 -2269
rect 478 -2275 479 -2269
rect 485 -2275 486 -2269
rect 502 -2288 503 -2274
rect 534 -2275 535 -2269
rect 541 -2288 542 -2274
rect 548 -2275 549 -2269
rect 548 -2288 549 -2274
rect 548 -2275 549 -2269
rect 548 -2288 549 -2274
rect 198 -2277 199 -2269
rect 313 -2277 314 -2269
rect 359 -2277 360 -2269
rect 464 -2277 465 -2269
rect 471 -2277 472 -2269
rect 499 -2277 500 -2269
rect 534 -2288 535 -2276
rect 555 -2277 556 -2269
rect 212 -2288 213 -2278
rect 219 -2279 220 -2269
rect 226 -2279 227 -2269
rect 233 -2288 234 -2278
rect 261 -2279 262 -2269
rect 275 -2288 276 -2278
rect 289 -2288 290 -2278
rect 317 -2288 318 -2278
rect 408 -2279 409 -2269
rect 520 -2279 521 -2269
rect 205 -2281 206 -2269
rect 226 -2288 227 -2280
rect 268 -2281 269 -2269
rect 282 -2288 283 -2280
rect 296 -2281 297 -2269
rect 296 -2288 297 -2280
rect 296 -2281 297 -2269
rect 296 -2288 297 -2280
rect 303 -2281 304 -2269
rect 331 -2281 332 -2269
rect 415 -2288 416 -2280
rect 436 -2281 437 -2269
rect 457 -2281 458 -2269
rect 464 -2288 465 -2280
rect 474 -2281 475 -2269
rect 478 -2288 479 -2280
rect 513 -2281 514 -2269
rect 520 -2288 521 -2280
rect 247 -2283 248 -2269
rect 268 -2288 269 -2282
rect 303 -2288 304 -2282
rect 366 -2283 367 -2269
rect 432 -2283 433 -2269
rect 506 -2283 507 -2269
rect 513 -2288 514 -2282
rect 527 -2283 528 -2269
rect 331 -2288 332 -2284
rect 338 -2285 339 -2269
rect 362 -2285 363 -2269
rect 366 -2288 367 -2284
rect 443 -2285 444 -2269
rect 457 -2288 458 -2284
rect 492 -2285 493 -2269
rect 506 -2288 507 -2284
rect 527 -2288 528 -2284
rect 576 -2285 577 -2269
rect 450 -2288 451 -2286
rect 474 -2288 475 -2286
rect 576 -2288 577 -2286
rect 583 -2287 584 -2269
rect 177 -2298 178 -2296
rect 177 -2305 178 -2297
rect 177 -2298 178 -2296
rect 177 -2305 178 -2297
rect 212 -2298 213 -2296
rect 215 -2305 216 -2297
rect 226 -2298 227 -2296
rect 243 -2298 244 -2296
rect 247 -2305 248 -2297
rect 254 -2298 255 -2296
rect 275 -2298 276 -2296
rect 327 -2298 328 -2296
rect 338 -2298 339 -2296
rect 345 -2298 346 -2296
rect 366 -2298 367 -2296
rect 369 -2305 370 -2297
rect 380 -2298 381 -2296
rect 380 -2305 381 -2297
rect 380 -2298 381 -2296
rect 380 -2305 381 -2297
rect 408 -2305 409 -2297
rect 415 -2298 416 -2296
rect 422 -2298 423 -2296
rect 439 -2298 440 -2296
rect 443 -2298 444 -2296
rect 464 -2298 465 -2296
rect 502 -2298 503 -2296
rect 513 -2298 514 -2296
rect 520 -2298 521 -2296
rect 527 -2305 528 -2297
rect 534 -2298 535 -2296
rect 541 -2298 542 -2296
rect 569 -2298 570 -2296
rect 576 -2298 577 -2296
rect 597 -2305 598 -2297
rect 604 -2305 605 -2297
rect 639 -2298 640 -2296
rect 646 -2305 647 -2297
rect 226 -2305 227 -2299
rect 264 -2305 265 -2299
rect 282 -2300 283 -2296
rect 289 -2300 290 -2296
rect 296 -2300 297 -2296
rect 306 -2300 307 -2296
rect 313 -2305 314 -2299
rect 317 -2300 318 -2296
rect 432 -2300 433 -2296
rect 457 -2300 458 -2296
rect 506 -2300 507 -2296
rect 509 -2305 510 -2299
rect 614 -2305 615 -2299
rect 639 -2305 640 -2299
rect 233 -2302 234 -2296
rect 233 -2305 234 -2301
rect 233 -2302 234 -2296
rect 233 -2305 234 -2301
rect 254 -2305 255 -2301
rect 285 -2305 286 -2301
rect 289 -2305 290 -2301
rect 310 -2302 311 -2296
rect 317 -2305 318 -2301
rect 331 -2302 332 -2296
rect 446 -2302 447 -2296
rect 450 -2302 451 -2296
rect 268 -2304 269 -2296
rect 296 -2305 297 -2303
rect 170 -2315 171 -2313
rect 177 -2315 178 -2313
rect 226 -2315 227 -2313
rect 282 -2315 283 -2313
rect 296 -2315 297 -2313
rect 306 -2315 307 -2313
rect 380 -2315 381 -2313
rect 387 -2315 388 -2313
rect 404 -2315 405 -2313
rect 408 -2315 409 -2313
rect 527 -2315 528 -2313
rect 534 -2315 535 -2313
rect 597 -2315 598 -2313
rect 611 -2315 612 -2313
rect 642 -2315 643 -2313
rect 646 -2315 647 -2313
rect 233 -2317 234 -2313
rect 240 -2317 241 -2313
rect 247 -2317 248 -2313
rect 268 -2317 269 -2313
rect 278 -2317 279 -2313
rect 317 -2317 318 -2313
rect 254 -2319 255 -2313
rect 275 -2319 276 -2313
<< labels >>
rlabel pdiffusion 3 -8 3 -8 0 cellNo=39
rlabel pdiffusion 10 -8 10 -8 0 cellNo=225
rlabel pdiffusion 17 -8 17 -8 0 cellNo=92
rlabel pdiffusion 24 -8 24 -8 0 cellNo=295
rlabel pdiffusion 31 -8 31 -8 0 cellNo=175
rlabel pdiffusion 38 -8 38 -8 0 cellNo=556
rlabel pdiffusion 178 -8 178 -8 0 feedthrough
rlabel pdiffusion 185 -8 185 -8 0 cellNo=852
rlabel pdiffusion 192 -8 192 -8 0 cellNo=622
rlabel pdiffusion 199 -8 199 -8 0 cellNo=895
rlabel pdiffusion 206 -8 206 -8 0 cellNo=62
rlabel pdiffusion 213 -8 213 -8 0 feedthrough
rlabel pdiffusion 255 -8 255 -8 0 cellNo=218
rlabel pdiffusion 269 -8 269 -8 0 cellNo=141
rlabel pdiffusion 276 -8 276 -8 0 feedthrough
rlabel pdiffusion 283 -8 283 -8 0 feedthrough
rlabel pdiffusion 311 -8 311 -8 0 feedthrough
rlabel pdiffusion 346 -8 346 -8 0 cellNo=667
rlabel pdiffusion 360 -8 360 -8 0 cellNo=968
rlabel pdiffusion 367 -8 367 -8 0 feedthrough
rlabel pdiffusion 3 -25 3 -25 0 cellNo=73
rlabel pdiffusion 10 -25 10 -25 0 cellNo=970
rlabel pdiffusion 17 -25 17 -25 0 cellNo=129
rlabel pdiffusion 24 -25 24 -25 0 cellNo=171
rlabel pdiffusion 31 -25 31 -25 0 cellNo=316
rlabel pdiffusion 157 -25 157 -25 0 cellNo=435
rlabel pdiffusion 199 -25 199 -25 0 cellNo=405
rlabel pdiffusion 213 -25 213 -25 0 cellNo=52
rlabel pdiffusion 220 -25 220 -25 0 feedthrough
rlabel pdiffusion 234 -25 234 -25 0 feedthrough
rlabel pdiffusion 241 -25 241 -25 0 feedthrough
rlabel pdiffusion 248 -25 248 -25 0 cellNo=876
rlabel pdiffusion 255 -25 255 -25 0 feedthrough
rlabel pdiffusion 262 -25 262 -25 0 feedthrough
rlabel pdiffusion 269 -25 269 -25 0 cellNo=50
rlabel pdiffusion 283 -25 283 -25 0 feedthrough
rlabel pdiffusion 297 -25 297 -25 0 cellNo=779
rlabel pdiffusion 304 -25 304 -25 0 feedthrough
rlabel pdiffusion 332 -25 332 -25 0 cellNo=278
rlabel pdiffusion 339 -25 339 -25 0 cellNo=602
rlabel pdiffusion 367 -25 367 -25 0 feedthrough
rlabel pdiffusion 374 -25 374 -25 0 feedthrough
rlabel pdiffusion 381 -25 381 -25 0 cellNo=934
rlabel pdiffusion 388 -25 388 -25 0 feedthrough
rlabel pdiffusion 395 -25 395 -25 0 feedthrough
rlabel pdiffusion 3 -46 3 -46 0 cellNo=148
rlabel pdiffusion 10 -46 10 -46 0 cellNo=159
rlabel pdiffusion 17 -46 17 -46 0 cellNo=448
rlabel pdiffusion 24 -46 24 -46 0 cellNo=302
rlabel pdiffusion 101 -46 101 -46 0 cellNo=46
rlabel pdiffusion 108 -46 108 -46 0 cellNo=742
rlabel pdiffusion 157 -46 157 -46 0 feedthrough
rlabel pdiffusion 164 -46 164 -46 0 cellNo=842
rlabel pdiffusion 171 -46 171 -46 0 cellNo=160
rlabel pdiffusion 178 -46 178 -46 0 feedthrough
rlabel pdiffusion 185 -46 185 -46 0 cellNo=760
rlabel pdiffusion 192 -46 192 -46 0 cellNo=745
rlabel pdiffusion 199 -46 199 -46 0 feedthrough
rlabel pdiffusion 206 -46 206 -46 0 feedthrough
rlabel pdiffusion 213 -46 213 -46 0 cellNo=154
rlabel pdiffusion 220 -46 220 -46 0 feedthrough
rlabel pdiffusion 227 -46 227 -46 0 feedthrough
rlabel pdiffusion 234 -46 234 -46 0 cellNo=31
rlabel pdiffusion 241 -46 241 -46 0 feedthrough
rlabel pdiffusion 248 -46 248 -46 0 feedthrough
rlabel pdiffusion 255 -46 255 -46 0 cellNo=377
rlabel pdiffusion 262 -46 262 -46 0 feedthrough
rlabel pdiffusion 269 -46 269 -46 0 feedthrough
rlabel pdiffusion 276 -46 276 -46 0 feedthrough
rlabel pdiffusion 283 -46 283 -46 0 feedthrough
rlabel pdiffusion 290 -46 290 -46 0 feedthrough
rlabel pdiffusion 297 -46 297 -46 0 cellNo=964
rlabel pdiffusion 304 -46 304 -46 0 cellNo=582
rlabel pdiffusion 311 -46 311 -46 0 feedthrough
rlabel pdiffusion 318 -46 318 -46 0 feedthrough
rlabel pdiffusion 325 -46 325 -46 0 feedthrough
rlabel pdiffusion 332 -46 332 -46 0 feedthrough
rlabel pdiffusion 339 -46 339 -46 0 cellNo=863
rlabel pdiffusion 346 -46 346 -46 0 feedthrough
rlabel pdiffusion 353 -46 353 -46 0 feedthrough
rlabel pdiffusion 360 -46 360 -46 0 cellNo=298
rlabel pdiffusion 367 -46 367 -46 0 feedthrough
rlabel pdiffusion 374 -46 374 -46 0 cellNo=618
rlabel pdiffusion 381 -46 381 -46 0 cellNo=321
rlabel pdiffusion 388 -46 388 -46 0 feedthrough
rlabel pdiffusion 395 -46 395 -46 0 feedthrough
rlabel pdiffusion 402 -46 402 -46 0 cellNo=713
rlabel pdiffusion 409 -46 409 -46 0 cellNo=336
rlabel pdiffusion 416 -46 416 -46 0 feedthrough
rlabel pdiffusion 423 -46 423 -46 0 feedthrough
rlabel pdiffusion 430 -46 430 -46 0 feedthrough
rlabel pdiffusion 437 -46 437 -46 0 cellNo=624
rlabel pdiffusion 444 -46 444 -46 0 cellNo=733
rlabel pdiffusion 451 -46 451 -46 0 feedthrough
rlabel pdiffusion 3 -83 3 -83 0 cellNo=121
rlabel pdiffusion 10 -83 10 -83 0 cellNo=710
rlabel pdiffusion 17 -83 17 -83 0 cellNo=190
rlabel pdiffusion 24 -83 24 -83 0 cellNo=899
rlabel pdiffusion 87 -83 87 -83 0 feedthrough
rlabel pdiffusion 94 -83 94 -83 0 feedthrough
rlabel pdiffusion 101 -83 101 -83 0 feedthrough
rlabel pdiffusion 108 -83 108 -83 0 cellNo=764
rlabel pdiffusion 115 -83 115 -83 0 cellNo=26
rlabel pdiffusion 122 -83 122 -83 0 cellNo=564
rlabel pdiffusion 129 -83 129 -83 0 feedthrough
rlabel pdiffusion 136 -83 136 -83 0 feedthrough
rlabel pdiffusion 143 -83 143 -83 0 feedthrough
rlabel pdiffusion 150 -83 150 -83 0 feedthrough
rlabel pdiffusion 157 -83 157 -83 0 cellNo=573
rlabel pdiffusion 164 -83 164 -83 0 feedthrough
rlabel pdiffusion 171 -83 171 -83 0 feedthrough
rlabel pdiffusion 178 -83 178 -83 0 feedthrough
rlabel pdiffusion 185 -83 185 -83 0 cellNo=490
rlabel pdiffusion 192 -83 192 -83 0 feedthrough
rlabel pdiffusion 199 -83 199 -83 0 cellNo=189
rlabel pdiffusion 206 -83 206 -83 0 feedthrough
rlabel pdiffusion 213 -83 213 -83 0 cellNo=471
rlabel pdiffusion 220 -83 220 -83 0 cellNo=694
rlabel pdiffusion 227 -83 227 -83 0 feedthrough
rlabel pdiffusion 234 -83 234 -83 0 cellNo=487
rlabel pdiffusion 241 -83 241 -83 0 cellNo=980
rlabel pdiffusion 248 -83 248 -83 0 feedthrough
rlabel pdiffusion 255 -83 255 -83 0 cellNo=855
rlabel pdiffusion 262 -83 262 -83 0 feedthrough
rlabel pdiffusion 269 -83 269 -83 0 feedthrough
rlabel pdiffusion 276 -83 276 -83 0 feedthrough
rlabel pdiffusion 283 -83 283 -83 0 feedthrough
rlabel pdiffusion 290 -83 290 -83 0 feedthrough
rlabel pdiffusion 297 -83 297 -83 0 feedthrough
rlabel pdiffusion 304 -83 304 -83 0 feedthrough
rlabel pdiffusion 311 -83 311 -83 0 cellNo=83
rlabel pdiffusion 318 -83 318 -83 0 feedthrough
rlabel pdiffusion 325 -83 325 -83 0 feedthrough
rlabel pdiffusion 332 -83 332 -83 0 feedthrough
rlabel pdiffusion 339 -83 339 -83 0 cellNo=608
rlabel pdiffusion 346 -83 346 -83 0 cellNo=507
rlabel pdiffusion 353 -83 353 -83 0 cellNo=771
rlabel pdiffusion 360 -83 360 -83 0 cellNo=238
rlabel pdiffusion 367 -83 367 -83 0 cellNo=844
rlabel pdiffusion 374 -83 374 -83 0 feedthrough
rlabel pdiffusion 381 -83 381 -83 0 feedthrough
rlabel pdiffusion 388 -83 388 -83 0 feedthrough
rlabel pdiffusion 395 -83 395 -83 0 feedthrough
rlabel pdiffusion 402 -83 402 -83 0 feedthrough
rlabel pdiffusion 409 -83 409 -83 0 feedthrough
rlabel pdiffusion 416 -83 416 -83 0 feedthrough
rlabel pdiffusion 423 -83 423 -83 0 feedthrough
rlabel pdiffusion 430 -83 430 -83 0 feedthrough
rlabel pdiffusion 437 -83 437 -83 0 feedthrough
rlabel pdiffusion 444 -83 444 -83 0 feedthrough
rlabel pdiffusion 451 -83 451 -83 0 feedthrough
rlabel pdiffusion 458 -83 458 -83 0 feedthrough
rlabel pdiffusion 465 -83 465 -83 0 feedthrough
rlabel pdiffusion 472 -83 472 -83 0 feedthrough
rlabel pdiffusion 479 -83 479 -83 0 feedthrough
rlabel pdiffusion 486 -83 486 -83 0 feedthrough
rlabel pdiffusion 493 -83 493 -83 0 cellNo=262
rlabel pdiffusion 500 -83 500 -83 0 feedthrough
rlabel pdiffusion 507 -83 507 -83 0 cellNo=609
rlabel pdiffusion 563 -83 563 -83 0 cellNo=887
rlabel pdiffusion 577 -83 577 -83 0 cellNo=535
rlabel pdiffusion 584 -83 584 -83 0 feedthrough
rlabel pdiffusion 3 -138 3 -138 0 cellNo=133
rlabel pdiffusion 10 -138 10 -138 0 cellNo=680
rlabel pdiffusion 17 -138 17 -138 0 cellNo=768
rlabel pdiffusion 52 -138 52 -138 0 cellNo=574
rlabel pdiffusion 59 -138 59 -138 0 feedthrough
rlabel pdiffusion 66 -138 66 -138 0 feedthrough
rlabel pdiffusion 73 -138 73 -138 0 feedthrough
rlabel pdiffusion 80 -138 80 -138 0 feedthrough
rlabel pdiffusion 87 -138 87 -138 0 feedthrough
rlabel pdiffusion 94 -138 94 -138 0 feedthrough
rlabel pdiffusion 101 -138 101 -138 0 cellNo=720
rlabel pdiffusion 108 -138 108 -138 0 feedthrough
rlabel pdiffusion 115 -138 115 -138 0 feedthrough
rlabel pdiffusion 122 -138 122 -138 0 feedthrough
rlabel pdiffusion 129 -138 129 -138 0 feedthrough
rlabel pdiffusion 136 -138 136 -138 0 feedthrough
rlabel pdiffusion 143 -138 143 -138 0 feedthrough
rlabel pdiffusion 150 -138 150 -138 0 feedthrough
rlabel pdiffusion 157 -138 157 -138 0 feedthrough
rlabel pdiffusion 164 -138 164 -138 0 feedthrough
rlabel pdiffusion 171 -138 171 -138 0 feedthrough
rlabel pdiffusion 178 -138 178 -138 0 cellNo=207
rlabel pdiffusion 185 -138 185 -138 0 cellNo=40
rlabel pdiffusion 192 -138 192 -138 0 cellNo=366
rlabel pdiffusion 199 -138 199 -138 0 feedthrough
rlabel pdiffusion 206 -138 206 -138 0 feedthrough
rlabel pdiffusion 213 -138 213 -138 0 cellNo=15
rlabel pdiffusion 220 -138 220 -138 0 cellNo=519
rlabel pdiffusion 227 -138 227 -138 0 cellNo=300
rlabel pdiffusion 234 -138 234 -138 0 feedthrough
rlabel pdiffusion 241 -138 241 -138 0 cellNo=607
rlabel pdiffusion 248 -138 248 -138 0 feedthrough
rlabel pdiffusion 255 -138 255 -138 0 feedthrough
rlabel pdiffusion 262 -138 262 -138 0 feedthrough
rlabel pdiffusion 269 -138 269 -138 0 feedthrough
rlabel pdiffusion 276 -138 276 -138 0 feedthrough
rlabel pdiffusion 283 -138 283 -138 0 cellNo=990
rlabel pdiffusion 290 -138 290 -138 0 feedthrough
rlabel pdiffusion 297 -138 297 -138 0 cellNo=597
rlabel pdiffusion 304 -138 304 -138 0 cellNo=224
rlabel pdiffusion 311 -138 311 -138 0 feedthrough
rlabel pdiffusion 318 -138 318 -138 0 feedthrough
rlabel pdiffusion 325 -138 325 -138 0 feedthrough
rlabel pdiffusion 332 -138 332 -138 0 cellNo=263
rlabel pdiffusion 339 -138 339 -138 0 cellNo=917
rlabel pdiffusion 346 -138 346 -138 0 feedthrough
rlabel pdiffusion 353 -138 353 -138 0 cellNo=635
rlabel pdiffusion 360 -138 360 -138 0 cellNo=798
rlabel pdiffusion 367 -138 367 -138 0 cellNo=580
rlabel pdiffusion 374 -138 374 -138 0 cellNo=339
rlabel pdiffusion 381 -138 381 -138 0 cellNo=699
rlabel pdiffusion 388 -138 388 -138 0 cellNo=891
rlabel pdiffusion 395 -138 395 -138 0 feedthrough
rlabel pdiffusion 402 -138 402 -138 0 feedthrough
rlabel pdiffusion 409 -138 409 -138 0 feedthrough
rlabel pdiffusion 416 -138 416 -138 0 feedthrough
rlabel pdiffusion 423 -138 423 -138 0 cellNo=384
rlabel pdiffusion 430 -138 430 -138 0 feedthrough
rlabel pdiffusion 437 -138 437 -138 0 feedthrough
rlabel pdiffusion 444 -138 444 -138 0 feedthrough
rlabel pdiffusion 451 -138 451 -138 0 feedthrough
rlabel pdiffusion 458 -138 458 -138 0 feedthrough
rlabel pdiffusion 465 -138 465 -138 0 feedthrough
rlabel pdiffusion 472 -138 472 -138 0 feedthrough
rlabel pdiffusion 479 -138 479 -138 0 feedthrough
rlabel pdiffusion 486 -138 486 -138 0 feedthrough
rlabel pdiffusion 493 -138 493 -138 0 feedthrough
rlabel pdiffusion 500 -138 500 -138 0 feedthrough
rlabel pdiffusion 507 -138 507 -138 0 feedthrough
rlabel pdiffusion 514 -138 514 -138 0 feedthrough
rlabel pdiffusion 521 -138 521 -138 0 feedthrough
rlabel pdiffusion 528 -138 528 -138 0 feedthrough
rlabel pdiffusion 535 -138 535 -138 0 feedthrough
rlabel pdiffusion 542 -138 542 -138 0 feedthrough
rlabel pdiffusion 549 -138 549 -138 0 cellNo=518
rlabel pdiffusion 556 -138 556 -138 0 feedthrough
rlabel pdiffusion 563 -138 563 -138 0 feedthrough
rlabel pdiffusion 570 -138 570 -138 0 feedthrough
rlabel pdiffusion 577 -138 577 -138 0 feedthrough
rlabel pdiffusion 584 -138 584 -138 0 feedthrough
rlabel pdiffusion 591 -138 591 -138 0 cellNo=719
rlabel pdiffusion 598 -138 598 -138 0 feedthrough
rlabel pdiffusion 619 -138 619 -138 0 feedthrough
rlabel pdiffusion 3 -197 3 -197 0 cellNo=178
rlabel pdiffusion 10 -197 10 -197 0 cellNo=696
rlabel pdiffusion 66 -197 66 -197 0 feedthrough
rlabel pdiffusion 73 -197 73 -197 0 cellNo=111
rlabel pdiffusion 80 -197 80 -197 0 feedthrough
rlabel pdiffusion 87 -197 87 -197 0 feedthrough
rlabel pdiffusion 94 -197 94 -197 0 feedthrough
rlabel pdiffusion 101 -197 101 -197 0 feedthrough
rlabel pdiffusion 108 -197 108 -197 0 feedthrough
rlabel pdiffusion 115 -197 115 -197 0 feedthrough
rlabel pdiffusion 122 -197 122 -197 0 feedthrough
rlabel pdiffusion 129 -197 129 -197 0 feedthrough
rlabel pdiffusion 136 -197 136 -197 0 cellNo=285
rlabel pdiffusion 143 -197 143 -197 0 cellNo=372
rlabel pdiffusion 150 -197 150 -197 0 feedthrough
rlabel pdiffusion 157 -197 157 -197 0 feedthrough
rlabel pdiffusion 164 -197 164 -197 0 feedthrough
rlabel pdiffusion 171 -197 171 -197 0 cellNo=605
rlabel pdiffusion 178 -197 178 -197 0 feedthrough
rlabel pdiffusion 185 -197 185 -197 0 cellNo=265
rlabel pdiffusion 192 -197 192 -197 0 cellNo=307
rlabel pdiffusion 199 -197 199 -197 0 feedthrough
rlabel pdiffusion 206 -197 206 -197 0 cellNo=746
rlabel pdiffusion 213 -197 213 -197 0 cellNo=850
rlabel pdiffusion 220 -197 220 -197 0 feedthrough
rlabel pdiffusion 227 -197 227 -197 0 feedthrough
rlabel pdiffusion 234 -197 234 -197 0 cellNo=213
rlabel pdiffusion 241 -197 241 -197 0 feedthrough
rlabel pdiffusion 248 -197 248 -197 0 feedthrough
rlabel pdiffusion 255 -197 255 -197 0 feedthrough
rlabel pdiffusion 262 -197 262 -197 0 feedthrough
rlabel pdiffusion 269 -197 269 -197 0 feedthrough
rlabel pdiffusion 276 -197 276 -197 0 feedthrough
rlabel pdiffusion 283 -197 283 -197 0 feedthrough
rlabel pdiffusion 290 -197 290 -197 0 feedthrough
rlabel pdiffusion 297 -197 297 -197 0 cellNo=115
rlabel pdiffusion 304 -197 304 -197 0 cellNo=791
rlabel pdiffusion 311 -197 311 -197 0 feedthrough
rlabel pdiffusion 318 -197 318 -197 0 cellNo=526
rlabel pdiffusion 325 -197 325 -197 0 feedthrough
rlabel pdiffusion 332 -197 332 -197 0 feedthrough
rlabel pdiffusion 339 -197 339 -197 0 feedthrough
rlabel pdiffusion 346 -197 346 -197 0 feedthrough
rlabel pdiffusion 353 -197 353 -197 0 cellNo=439
rlabel pdiffusion 360 -197 360 -197 0 cellNo=792
rlabel pdiffusion 367 -197 367 -197 0 feedthrough
rlabel pdiffusion 374 -197 374 -197 0 cellNo=22
rlabel pdiffusion 381 -197 381 -197 0 feedthrough
rlabel pdiffusion 388 -197 388 -197 0 feedthrough
rlabel pdiffusion 395 -197 395 -197 0 cellNo=347
rlabel pdiffusion 402 -197 402 -197 0 cellNo=98
rlabel pdiffusion 409 -197 409 -197 0 feedthrough
rlabel pdiffusion 416 -197 416 -197 0 feedthrough
rlabel pdiffusion 423 -197 423 -197 0 feedthrough
rlabel pdiffusion 430 -197 430 -197 0 feedthrough
rlabel pdiffusion 437 -197 437 -197 0 cellNo=795
rlabel pdiffusion 444 -197 444 -197 0 feedthrough
rlabel pdiffusion 451 -197 451 -197 0 feedthrough
rlabel pdiffusion 458 -197 458 -197 0 cellNo=456
rlabel pdiffusion 465 -197 465 -197 0 feedthrough
rlabel pdiffusion 472 -197 472 -197 0 feedthrough
rlabel pdiffusion 479 -197 479 -197 0 feedthrough
rlabel pdiffusion 486 -197 486 -197 0 feedthrough
rlabel pdiffusion 493 -197 493 -197 0 feedthrough
rlabel pdiffusion 500 -197 500 -197 0 feedthrough
rlabel pdiffusion 507 -197 507 -197 0 cellNo=464
rlabel pdiffusion 514 -197 514 -197 0 feedthrough
rlabel pdiffusion 521 -197 521 -197 0 feedthrough
rlabel pdiffusion 528 -197 528 -197 0 feedthrough
rlabel pdiffusion 535 -197 535 -197 0 feedthrough
rlabel pdiffusion 542 -197 542 -197 0 cellNo=783
rlabel pdiffusion 549 -197 549 -197 0 feedthrough
rlabel pdiffusion 556 -197 556 -197 0 feedthrough
rlabel pdiffusion 563 -197 563 -197 0 feedthrough
rlabel pdiffusion 570 -197 570 -197 0 cellNo=531
rlabel pdiffusion 577 -197 577 -197 0 feedthrough
rlabel pdiffusion 584 -197 584 -197 0 feedthrough
rlabel pdiffusion 591 -197 591 -197 0 feedthrough
rlabel pdiffusion 633 -197 633 -197 0 feedthrough
rlabel pdiffusion 640 -197 640 -197 0 cellNo=578
rlabel pdiffusion 647 -197 647 -197 0 feedthrough
rlabel pdiffusion 3 -254 3 -254 0 cellNo=557
rlabel pdiffusion 17 -254 17 -254 0 feedthrough
rlabel pdiffusion 24 -254 24 -254 0 feedthrough
rlabel pdiffusion 31 -254 31 -254 0 feedthrough
rlabel pdiffusion 38 -254 38 -254 0 feedthrough
rlabel pdiffusion 45 -254 45 -254 0 feedthrough
rlabel pdiffusion 52 -254 52 -254 0 cellNo=533
rlabel pdiffusion 59 -254 59 -254 0 feedthrough
rlabel pdiffusion 66 -254 66 -254 0 feedthrough
rlabel pdiffusion 73 -254 73 -254 0 feedthrough
rlabel pdiffusion 80 -254 80 -254 0 feedthrough
rlabel pdiffusion 87 -254 87 -254 0 feedthrough
rlabel pdiffusion 94 -254 94 -254 0 feedthrough
rlabel pdiffusion 101 -254 101 -254 0 cellNo=569
rlabel pdiffusion 108 -254 108 -254 0 cellNo=120
rlabel pdiffusion 115 -254 115 -254 0 feedthrough
rlabel pdiffusion 122 -254 122 -254 0 feedthrough
rlabel pdiffusion 129 -254 129 -254 0 cellNo=603
rlabel pdiffusion 136 -254 136 -254 0 cellNo=554
rlabel pdiffusion 143 -254 143 -254 0 cellNo=228
rlabel pdiffusion 150 -254 150 -254 0 feedthrough
rlabel pdiffusion 157 -254 157 -254 0 cellNo=652
rlabel pdiffusion 164 -254 164 -254 0 feedthrough
rlabel pdiffusion 171 -254 171 -254 0 feedthrough
rlabel pdiffusion 178 -254 178 -254 0 feedthrough
rlabel pdiffusion 185 -254 185 -254 0 feedthrough
rlabel pdiffusion 192 -254 192 -254 0 cellNo=323
rlabel pdiffusion 199 -254 199 -254 0 feedthrough
rlabel pdiffusion 206 -254 206 -254 0 cellNo=157
rlabel pdiffusion 213 -254 213 -254 0 cellNo=524
rlabel pdiffusion 220 -254 220 -254 0 cellNo=103
rlabel pdiffusion 227 -254 227 -254 0 cellNo=499
rlabel pdiffusion 234 -254 234 -254 0 feedthrough
rlabel pdiffusion 241 -254 241 -254 0 feedthrough
rlabel pdiffusion 248 -254 248 -254 0 feedthrough
rlabel pdiffusion 255 -254 255 -254 0 feedthrough
rlabel pdiffusion 262 -254 262 -254 0 feedthrough
rlabel pdiffusion 269 -254 269 -254 0 cellNo=201
rlabel pdiffusion 276 -254 276 -254 0 feedthrough
rlabel pdiffusion 283 -254 283 -254 0 feedthrough
rlabel pdiffusion 290 -254 290 -254 0 feedthrough
rlabel pdiffusion 297 -254 297 -254 0 feedthrough
rlabel pdiffusion 304 -254 304 -254 0 feedthrough
rlabel pdiffusion 311 -254 311 -254 0 feedthrough
rlabel pdiffusion 318 -254 318 -254 0 feedthrough
rlabel pdiffusion 325 -254 325 -254 0 feedthrough
rlabel pdiffusion 332 -254 332 -254 0 feedthrough
rlabel pdiffusion 339 -254 339 -254 0 cellNo=957
rlabel pdiffusion 346 -254 346 -254 0 feedthrough
rlabel pdiffusion 353 -254 353 -254 0 feedthrough
rlabel pdiffusion 360 -254 360 -254 0 feedthrough
rlabel pdiffusion 367 -254 367 -254 0 feedthrough
rlabel pdiffusion 374 -254 374 -254 0 feedthrough
rlabel pdiffusion 381 -254 381 -254 0 feedthrough
rlabel pdiffusion 388 -254 388 -254 0 cellNo=216
rlabel pdiffusion 395 -254 395 -254 0 cellNo=345
rlabel pdiffusion 402 -254 402 -254 0 feedthrough
rlabel pdiffusion 409 -254 409 -254 0 cellNo=41
rlabel pdiffusion 416 -254 416 -254 0 cellNo=286
rlabel pdiffusion 423 -254 423 -254 0 feedthrough
rlabel pdiffusion 430 -254 430 -254 0 feedthrough
rlabel pdiffusion 437 -254 437 -254 0 feedthrough
rlabel pdiffusion 444 -254 444 -254 0 feedthrough
rlabel pdiffusion 451 -254 451 -254 0 feedthrough
rlabel pdiffusion 458 -254 458 -254 0 cellNo=232
rlabel pdiffusion 465 -254 465 -254 0 cellNo=777
rlabel pdiffusion 472 -254 472 -254 0 feedthrough
rlabel pdiffusion 479 -254 479 -254 0 cellNo=633
rlabel pdiffusion 486 -254 486 -254 0 feedthrough
rlabel pdiffusion 493 -254 493 -254 0 feedthrough
rlabel pdiffusion 500 -254 500 -254 0 feedthrough
rlabel pdiffusion 507 -254 507 -254 0 cellNo=170
rlabel pdiffusion 514 -254 514 -254 0 feedthrough
rlabel pdiffusion 521 -254 521 -254 0 feedthrough
rlabel pdiffusion 528 -254 528 -254 0 feedthrough
rlabel pdiffusion 535 -254 535 -254 0 feedthrough
rlabel pdiffusion 542 -254 542 -254 0 feedthrough
rlabel pdiffusion 549 -254 549 -254 0 feedthrough
rlabel pdiffusion 556 -254 556 -254 0 feedthrough
rlabel pdiffusion 563 -254 563 -254 0 feedthrough
rlabel pdiffusion 570 -254 570 -254 0 cellNo=392
rlabel pdiffusion 577 -254 577 -254 0 feedthrough
rlabel pdiffusion 584 -254 584 -254 0 feedthrough
rlabel pdiffusion 591 -254 591 -254 0 feedthrough
rlabel pdiffusion 598 -254 598 -254 0 feedthrough
rlabel pdiffusion 605 -254 605 -254 0 feedthrough
rlabel pdiffusion 612 -254 612 -254 0 feedthrough
rlabel pdiffusion 619 -254 619 -254 0 feedthrough
rlabel pdiffusion 626 -254 626 -254 0 feedthrough
rlabel pdiffusion 633 -254 633 -254 0 feedthrough
rlabel pdiffusion 640 -254 640 -254 0 feedthrough
rlabel pdiffusion 647 -254 647 -254 0 feedthrough
rlabel pdiffusion 654 -254 654 -254 0 feedthrough
rlabel pdiffusion 661 -254 661 -254 0 feedthrough
rlabel pdiffusion 668 -254 668 -254 0 cellNo=806
rlabel pdiffusion 675 -254 675 -254 0 feedthrough
rlabel pdiffusion 682 -254 682 -254 0 feedthrough
rlabel pdiffusion 689 -254 689 -254 0 feedthrough
rlabel pdiffusion 696 -254 696 -254 0 feedthrough
rlabel pdiffusion 752 -254 752 -254 0 feedthrough
rlabel pdiffusion 857 -254 857 -254 0 cellNo=375
rlabel pdiffusion 31 -307 31 -307 0 feedthrough
rlabel pdiffusion 38 -307 38 -307 0 feedthrough
rlabel pdiffusion 45 -307 45 -307 0 cellNo=725
rlabel pdiffusion 52 -307 52 -307 0 feedthrough
rlabel pdiffusion 59 -307 59 -307 0 feedthrough
rlabel pdiffusion 66 -307 66 -307 0 cellNo=442
rlabel pdiffusion 73 -307 73 -307 0 feedthrough
rlabel pdiffusion 80 -307 80 -307 0 cellNo=997
rlabel pdiffusion 87 -307 87 -307 0 feedthrough
rlabel pdiffusion 94 -307 94 -307 0 feedthrough
rlabel pdiffusion 101 -307 101 -307 0 cellNo=346
rlabel pdiffusion 108 -307 108 -307 0 feedthrough
rlabel pdiffusion 115 -307 115 -307 0 cellNo=60
rlabel pdiffusion 122 -307 122 -307 0 feedthrough
rlabel pdiffusion 129 -307 129 -307 0 feedthrough
rlabel pdiffusion 136 -307 136 -307 0 cellNo=199
rlabel pdiffusion 143 -307 143 -307 0 feedthrough
rlabel pdiffusion 150 -307 150 -307 0 feedthrough
rlabel pdiffusion 157 -307 157 -307 0 feedthrough
rlabel pdiffusion 164 -307 164 -307 0 feedthrough
rlabel pdiffusion 171 -307 171 -307 0 feedthrough
rlabel pdiffusion 178 -307 178 -307 0 cellNo=803
rlabel pdiffusion 185 -307 185 -307 0 feedthrough
rlabel pdiffusion 192 -307 192 -307 0 feedthrough
rlabel pdiffusion 199 -307 199 -307 0 feedthrough
rlabel pdiffusion 206 -307 206 -307 0 feedthrough
rlabel pdiffusion 213 -307 213 -307 0 cellNo=469
rlabel pdiffusion 220 -307 220 -307 0 cellNo=679
rlabel pdiffusion 227 -307 227 -307 0 feedthrough
rlabel pdiffusion 234 -307 234 -307 0 cellNo=525
rlabel pdiffusion 241 -307 241 -307 0 cellNo=697
rlabel pdiffusion 248 -307 248 -307 0 cellNo=913
rlabel pdiffusion 255 -307 255 -307 0 cellNo=393
rlabel pdiffusion 262 -307 262 -307 0 feedthrough
rlabel pdiffusion 269 -307 269 -307 0 feedthrough
rlabel pdiffusion 276 -307 276 -307 0 feedthrough
rlabel pdiffusion 283 -307 283 -307 0 feedthrough
rlabel pdiffusion 290 -307 290 -307 0 cellNo=328
rlabel pdiffusion 297 -307 297 -307 0 cellNo=288
rlabel pdiffusion 304 -307 304 -307 0 feedthrough
rlabel pdiffusion 311 -307 311 -307 0 feedthrough
rlabel pdiffusion 318 -307 318 -307 0 feedthrough
rlabel pdiffusion 325 -307 325 -307 0 feedthrough
rlabel pdiffusion 332 -307 332 -307 0 cellNo=727
rlabel pdiffusion 339 -307 339 -307 0 cellNo=398
rlabel pdiffusion 346 -307 346 -307 0 feedthrough
rlabel pdiffusion 353 -307 353 -307 0 feedthrough
rlabel pdiffusion 360 -307 360 -307 0 feedthrough
rlabel pdiffusion 367 -307 367 -307 0 feedthrough
rlabel pdiffusion 374 -307 374 -307 0 cellNo=953
rlabel pdiffusion 381 -307 381 -307 0 feedthrough
rlabel pdiffusion 388 -307 388 -307 0 feedthrough
rlabel pdiffusion 395 -307 395 -307 0 cellNo=627
rlabel pdiffusion 402 -307 402 -307 0 cellNo=506
rlabel pdiffusion 409 -307 409 -307 0 feedthrough
rlabel pdiffusion 416 -307 416 -307 0 feedthrough
rlabel pdiffusion 423 -307 423 -307 0 cellNo=728
rlabel pdiffusion 430 -307 430 -307 0 feedthrough
rlabel pdiffusion 437 -307 437 -307 0 cellNo=317
rlabel pdiffusion 444 -307 444 -307 0 cellNo=192
rlabel pdiffusion 451 -307 451 -307 0 feedthrough
rlabel pdiffusion 458 -307 458 -307 0 feedthrough
rlabel pdiffusion 465 -307 465 -307 0 feedthrough
rlabel pdiffusion 472 -307 472 -307 0 feedthrough
rlabel pdiffusion 479 -307 479 -307 0 feedthrough
rlabel pdiffusion 486 -307 486 -307 0 feedthrough
rlabel pdiffusion 493 -307 493 -307 0 feedthrough
rlabel pdiffusion 500 -307 500 -307 0 feedthrough
rlabel pdiffusion 507 -307 507 -307 0 feedthrough
rlabel pdiffusion 514 -307 514 -307 0 feedthrough
rlabel pdiffusion 521 -307 521 -307 0 feedthrough
rlabel pdiffusion 528 -307 528 -307 0 feedthrough
rlabel pdiffusion 535 -307 535 -307 0 feedthrough
rlabel pdiffusion 542 -307 542 -307 0 cellNo=137
rlabel pdiffusion 549 -307 549 -307 0 feedthrough
rlabel pdiffusion 556 -307 556 -307 0 feedthrough
rlabel pdiffusion 563 -307 563 -307 0 cellNo=460
rlabel pdiffusion 570 -307 570 -307 0 feedthrough
rlabel pdiffusion 577 -307 577 -307 0 feedthrough
rlabel pdiffusion 584 -307 584 -307 0 feedthrough
rlabel pdiffusion 591 -307 591 -307 0 feedthrough
rlabel pdiffusion 598 -307 598 -307 0 feedthrough
rlabel pdiffusion 605 -307 605 -307 0 feedthrough
rlabel pdiffusion 612 -307 612 -307 0 feedthrough
rlabel pdiffusion 619 -307 619 -307 0 feedthrough
rlabel pdiffusion 626 -307 626 -307 0 feedthrough
rlabel pdiffusion 633 -307 633 -307 0 feedthrough
rlabel pdiffusion 640 -307 640 -307 0 feedthrough
rlabel pdiffusion 647 -307 647 -307 0 feedthrough
rlabel pdiffusion 654 -307 654 -307 0 feedthrough
rlabel pdiffusion 661 -307 661 -307 0 feedthrough
rlabel pdiffusion 668 -307 668 -307 0 feedthrough
rlabel pdiffusion 675 -307 675 -307 0 cellNo=780
rlabel pdiffusion 682 -307 682 -307 0 feedthrough
rlabel pdiffusion 689 -307 689 -307 0 feedthrough
rlabel pdiffusion 696 -307 696 -307 0 feedthrough
rlabel pdiffusion 703 -307 703 -307 0 feedthrough
rlabel pdiffusion 710 -307 710 -307 0 feedthrough
rlabel pdiffusion 717 -307 717 -307 0 feedthrough
rlabel pdiffusion 724 -307 724 -307 0 cellNo=104
rlabel pdiffusion 731 -307 731 -307 0 feedthrough
rlabel pdiffusion 738 -307 738 -307 0 feedthrough
rlabel pdiffusion 745 -307 745 -307 0 feedthrough
rlabel pdiffusion 752 -307 752 -307 0 feedthrough
rlabel pdiffusion 829 -307 829 -307 0 feedthrough
rlabel pdiffusion 857 -307 857 -307 0 feedthrough
rlabel pdiffusion 3 -378 3 -378 0 feedthrough
rlabel pdiffusion 10 -378 10 -378 0 feedthrough
rlabel pdiffusion 17 -378 17 -378 0 feedthrough
rlabel pdiffusion 24 -378 24 -378 0 feedthrough
rlabel pdiffusion 31 -378 31 -378 0 feedthrough
rlabel pdiffusion 38 -378 38 -378 0 feedthrough
rlabel pdiffusion 45 -378 45 -378 0 feedthrough
rlabel pdiffusion 52 -378 52 -378 0 feedthrough
rlabel pdiffusion 59 -378 59 -378 0 feedthrough
rlabel pdiffusion 66 -378 66 -378 0 feedthrough
rlabel pdiffusion 73 -378 73 -378 0 cellNo=311
rlabel pdiffusion 80 -378 80 -378 0 feedthrough
rlabel pdiffusion 87 -378 87 -378 0 feedthrough
rlabel pdiffusion 94 -378 94 -378 0 cellNo=403
rlabel pdiffusion 101 -378 101 -378 0 feedthrough
rlabel pdiffusion 108 -378 108 -378 0 cellNo=390
rlabel pdiffusion 115 -378 115 -378 0 feedthrough
rlabel pdiffusion 122 -378 122 -378 0 feedthrough
rlabel pdiffusion 129 -378 129 -378 0 cellNo=534
rlabel pdiffusion 136 -378 136 -378 0 cellNo=332
rlabel pdiffusion 143 -378 143 -378 0 cellNo=871
rlabel pdiffusion 150 -378 150 -378 0 cellNo=653
rlabel pdiffusion 157 -378 157 -378 0 feedthrough
rlabel pdiffusion 164 -378 164 -378 0 feedthrough
rlabel pdiffusion 171 -378 171 -378 0 feedthrough
rlabel pdiffusion 178 -378 178 -378 0 feedthrough
rlabel pdiffusion 185 -378 185 -378 0 feedthrough
rlabel pdiffusion 192 -378 192 -378 0 feedthrough
rlabel pdiffusion 199 -378 199 -378 0 cellNo=859
rlabel pdiffusion 206 -378 206 -378 0 cellNo=124
rlabel pdiffusion 213 -378 213 -378 0 cellNo=70
rlabel pdiffusion 220 -378 220 -378 0 feedthrough
rlabel pdiffusion 227 -378 227 -378 0 feedthrough
rlabel pdiffusion 234 -378 234 -378 0 cellNo=45
rlabel pdiffusion 241 -378 241 -378 0 feedthrough
rlabel pdiffusion 248 -378 248 -378 0 feedthrough
rlabel pdiffusion 255 -378 255 -378 0 feedthrough
rlabel pdiffusion 262 -378 262 -378 0 feedthrough
rlabel pdiffusion 269 -378 269 -378 0 feedthrough
rlabel pdiffusion 276 -378 276 -378 0 cellNo=543
rlabel pdiffusion 283 -378 283 -378 0 feedthrough
rlabel pdiffusion 290 -378 290 -378 0 feedthrough
rlabel pdiffusion 297 -378 297 -378 0 feedthrough
rlabel pdiffusion 304 -378 304 -378 0 feedthrough
rlabel pdiffusion 311 -378 311 -378 0 feedthrough
rlabel pdiffusion 318 -378 318 -378 0 feedthrough
rlabel pdiffusion 325 -378 325 -378 0 cellNo=29
rlabel pdiffusion 332 -378 332 -378 0 cellNo=867
rlabel pdiffusion 339 -378 339 -378 0 feedthrough
rlabel pdiffusion 346 -378 346 -378 0 feedthrough
rlabel pdiffusion 353 -378 353 -378 0 feedthrough
rlabel pdiffusion 360 -378 360 -378 0 cellNo=18
rlabel pdiffusion 367 -378 367 -378 0 cellNo=523
rlabel pdiffusion 374 -378 374 -378 0 cellNo=493
rlabel pdiffusion 381 -378 381 -378 0 feedthrough
rlabel pdiffusion 388 -378 388 -378 0 feedthrough
rlabel pdiffusion 395 -378 395 -378 0 feedthrough
rlabel pdiffusion 402 -378 402 -378 0 cellNo=306
rlabel pdiffusion 409 -378 409 -378 0 feedthrough
rlabel pdiffusion 416 -378 416 -378 0 feedthrough
rlabel pdiffusion 423 -378 423 -378 0 cellNo=358
rlabel pdiffusion 430 -378 430 -378 0 cellNo=362
rlabel pdiffusion 437 -378 437 -378 0 feedthrough
rlabel pdiffusion 444 -378 444 -378 0 feedthrough
rlabel pdiffusion 451 -378 451 -378 0 feedthrough
rlabel pdiffusion 458 -378 458 -378 0 feedthrough
rlabel pdiffusion 465 -378 465 -378 0 feedthrough
rlabel pdiffusion 472 -378 472 -378 0 cellNo=972
rlabel pdiffusion 479 -378 479 -378 0 feedthrough
rlabel pdiffusion 486 -378 486 -378 0 feedthrough
rlabel pdiffusion 493 -378 493 -378 0 cellNo=105
rlabel pdiffusion 500 -378 500 -378 0 feedthrough
rlabel pdiffusion 507 -378 507 -378 0 cellNo=44
rlabel pdiffusion 514 -378 514 -378 0 cellNo=271
rlabel pdiffusion 521 -378 521 -378 0 feedthrough
rlabel pdiffusion 528 -378 528 -378 0 feedthrough
rlabel pdiffusion 535 -378 535 -378 0 feedthrough
rlabel pdiffusion 542 -378 542 -378 0 feedthrough
rlabel pdiffusion 549 -378 549 -378 0 feedthrough
rlabel pdiffusion 556 -378 556 -378 0 feedthrough
rlabel pdiffusion 563 -378 563 -378 0 feedthrough
rlabel pdiffusion 570 -378 570 -378 0 feedthrough
rlabel pdiffusion 577 -378 577 -378 0 feedthrough
rlabel pdiffusion 584 -378 584 -378 0 cellNo=663
rlabel pdiffusion 591 -378 591 -378 0 feedthrough
rlabel pdiffusion 598 -378 598 -378 0 feedthrough
rlabel pdiffusion 605 -378 605 -378 0 cellNo=595
rlabel pdiffusion 612 -378 612 -378 0 feedthrough
rlabel pdiffusion 619 -378 619 -378 0 feedthrough
rlabel pdiffusion 626 -378 626 -378 0 feedthrough
rlabel pdiffusion 633 -378 633 -378 0 feedthrough
rlabel pdiffusion 640 -378 640 -378 0 feedthrough
rlabel pdiffusion 647 -378 647 -378 0 feedthrough
rlabel pdiffusion 654 -378 654 -378 0 feedthrough
rlabel pdiffusion 661 -378 661 -378 0 feedthrough
rlabel pdiffusion 668 -378 668 -378 0 feedthrough
rlabel pdiffusion 675 -378 675 -378 0 feedthrough
rlabel pdiffusion 682 -378 682 -378 0 feedthrough
rlabel pdiffusion 689 -378 689 -378 0 feedthrough
rlabel pdiffusion 696 -378 696 -378 0 feedthrough
rlabel pdiffusion 703 -378 703 -378 0 feedthrough
rlabel pdiffusion 710 -378 710 -378 0 feedthrough
rlabel pdiffusion 717 -378 717 -378 0 feedthrough
rlabel pdiffusion 724 -378 724 -378 0 feedthrough
rlabel pdiffusion 731 -378 731 -378 0 feedthrough
rlabel pdiffusion 738 -378 738 -378 0 feedthrough
rlabel pdiffusion 745 -378 745 -378 0 feedthrough
rlabel pdiffusion 752 -378 752 -378 0 feedthrough
rlabel pdiffusion 759 -378 759 -378 0 feedthrough
rlabel pdiffusion 766 -378 766 -378 0 feedthrough
rlabel pdiffusion 773 -378 773 -378 0 feedthrough
rlabel pdiffusion 780 -378 780 -378 0 feedthrough
rlabel pdiffusion 787 -378 787 -378 0 feedthrough
rlabel pdiffusion 794 -378 794 -378 0 feedthrough
rlabel pdiffusion 801 -378 801 -378 0 feedthrough
rlabel pdiffusion 808 -378 808 -378 0 feedthrough
rlabel pdiffusion 815 -378 815 -378 0 feedthrough
rlabel pdiffusion 822 -378 822 -378 0 feedthrough
rlabel pdiffusion 829 -378 829 -378 0 feedthrough
rlabel pdiffusion 836 -378 836 -378 0 feedthrough
rlabel pdiffusion 843 -378 843 -378 0 feedthrough
rlabel pdiffusion 850 -378 850 -378 0 cellNo=94
rlabel pdiffusion 857 -378 857 -378 0 feedthrough
rlabel pdiffusion 864 -378 864 -378 0 feedthrough
rlabel pdiffusion 871 -378 871 -378 0 feedthrough
rlabel pdiffusion 878 -378 878 -378 0 cellNo=807
rlabel pdiffusion 885 -378 885 -378 0 cellNo=695
rlabel pdiffusion 892 -378 892 -378 0 feedthrough
rlabel pdiffusion 3 -467 3 -467 0 feedthrough
rlabel pdiffusion 10 -467 10 -467 0 feedthrough
rlabel pdiffusion 17 -467 17 -467 0 feedthrough
rlabel pdiffusion 24 -467 24 -467 0 feedthrough
rlabel pdiffusion 31 -467 31 -467 0 feedthrough
rlabel pdiffusion 38 -467 38 -467 0 feedthrough
rlabel pdiffusion 45 -467 45 -467 0 cellNo=195
rlabel pdiffusion 52 -467 52 -467 0 cellNo=935
rlabel pdiffusion 59 -467 59 -467 0 feedthrough
rlabel pdiffusion 66 -467 66 -467 0 feedthrough
rlabel pdiffusion 73 -467 73 -467 0 feedthrough
rlabel pdiffusion 80 -467 80 -467 0 cellNo=150
rlabel pdiffusion 87 -467 87 -467 0 feedthrough
rlabel pdiffusion 94 -467 94 -467 0 feedthrough
rlabel pdiffusion 101 -467 101 -467 0 cellNo=542
rlabel pdiffusion 108 -467 108 -467 0 cellNo=820
rlabel pdiffusion 115 -467 115 -467 0 cellNo=833
rlabel pdiffusion 122 -467 122 -467 0 feedthrough
rlabel pdiffusion 129 -467 129 -467 0 feedthrough
rlabel pdiffusion 136 -467 136 -467 0 feedthrough
rlabel pdiffusion 143 -467 143 -467 0 feedthrough
rlabel pdiffusion 150 -467 150 -467 0 cellNo=512
rlabel pdiffusion 157 -467 157 -467 0 cellNo=21
rlabel pdiffusion 164 -467 164 -467 0 cellNo=945
rlabel pdiffusion 171 -467 171 -467 0 feedthrough
rlabel pdiffusion 178 -467 178 -467 0 feedthrough
rlabel pdiffusion 185 -467 185 -467 0 feedthrough
rlabel pdiffusion 192 -467 192 -467 0 cellNo=164
rlabel pdiffusion 199 -467 199 -467 0 cellNo=823
rlabel pdiffusion 206 -467 206 -467 0 feedthrough
rlabel pdiffusion 213 -467 213 -467 0 cellNo=724
rlabel pdiffusion 220 -467 220 -467 0 cellNo=907
rlabel pdiffusion 227 -467 227 -467 0 feedthrough
rlabel pdiffusion 234 -467 234 -467 0 feedthrough
rlabel pdiffusion 241 -467 241 -467 0 cellNo=550
rlabel pdiffusion 248 -467 248 -467 0 feedthrough
rlabel pdiffusion 255 -467 255 -467 0 feedthrough
rlabel pdiffusion 262 -467 262 -467 0 feedthrough
rlabel pdiffusion 269 -467 269 -467 0 feedthrough
rlabel pdiffusion 276 -467 276 -467 0 feedthrough
rlabel pdiffusion 283 -467 283 -467 0 feedthrough
rlabel pdiffusion 290 -467 290 -467 0 feedthrough
rlabel pdiffusion 297 -467 297 -467 0 cellNo=230
rlabel pdiffusion 304 -467 304 -467 0 cellNo=101
rlabel pdiffusion 311 -467 311 -467 0 feedthrough
rlabel pdiffusion 318 -467 318 -467 0 feedthrough
rlabel pdiffusion 325 -467 325 -467 0 feedthrough
rlabel pdiffusion 332 -467 332 -467 0 feedthrough
rlabel pdiffusion 339 -467 339 -467 0 feedthrough
rlabel pdiffusion 346 -467 346 -467 0 cellNo=223
rlabel pdiffusion 353 -467 353 -467 0 feedthrough
rlabel pdiffusion 360 -467 360 -467 0 feedthrough
rlabel pdiffusion 367 -467 367 -467 0 cellNo=8
rlabel pdiffusion 374 -467 374 -467 0 feedthrough
rlabel pdiffusion 381 -467 381 -467 0 cellNo=912
rlabel pdiffusion 388 -467 388 -467 0 cellNo=186
rlabel pdiffusion 395 -467 395 -467 0 feedthrough
rlabel pdiffusion 402 -467 402 -467 0 feedthrough
rlabel pdiffusion 409 -467 409 -467 0 feedthrough
rlabel pdiffusion 416 -467 416 -467 0 cellNo=177
rlabel pdiffusion 423 -467 423 -467 0 feedthrough
rlabel pdiffusion 430 -467 430 -467 0 cellNo=373
rlabel pdiffusion 437 -467 437 -467 0 cellNo=57
rlabel pdiffusion 444 -467 444 -467 0 feedthrough
rlabel pdiffusion 451 -467 451 -467 0 feedthrough
rlabel pdiffusion 458 -467 458 -467 0 cellNo=305
rlabel pdiffusion 465 -467 465 -467 0 feedthrough
rlabel pdiffusion 472 -467 472 -467 0 feedthrough
rlabel pdiffusion 479 -467 479 -467 0 feedthrough
rlabel pdiffusion 486 -467 486 -467 0 cellNo=601
rlabel pdiffusion 493 -467 493 -467 0 feedthrough
rlabel pdiffusion 500 -467 500 -467 0 cellNo=870
rlabel pdiffusion 507 -467 507 -467 0 cellNo=593
rlabel pdiffusion 514 -467 514 -467 0 feedthrough
rlabel pdiffusion 521 -467 521 -467 0 cellNo=16
rlabel pdiffusion 528 -467 528 -467 0 feedthrough
rlabel pdiffusion 535 -467 535 -467 0 feedthrough
rlabel pdiffusion 542 -467 542 -467 0 feedthrough
rlabel pdiffusion 549 -467 549 -467 0 feedthrough
rlabel pdiffusion 556 -467 556 -467 0 feedthrough
rlabel pdiffusion 563 -467 563 -467 0 feedthrough
rlabel pdiffusion 570 -467 570 -467 0 feedthrough
rlabel pdiffusion 577 -467 577 -467 0 feedthrough
rlabel pdiffusion 584 -467 584 -467 0 feedthrough
rlabel pdiffusion 591 -467 591 -467 0 feedthrough
rlabel pdiffusion 598 -467 598 -467 0 feedthrough
rlabel pdiffusion 605 -467 605 -467 0 feedthrough
rlabel pdiffusion 612 -467 612 -467 0 feedthrough
rlabel pdiffusion 619 -467 619 -467 0 cellNo=420
rlabel pdiffusion 626 -467 626 -467 0 feedthrough
rlabel pdiffusion 633 -467 633 -467 0 feedthrough
rlabel pdiffusion 640 -467 640 -467 0 feedthrough
rlabel pdiffusion 647 -467 647 -467 0 feedthrough
rlabel pdiffusion 654 -467 654 -467 0 feedthrough
rlabel pdiffusion 661 -467 661 -467 0 feedthrough
rlabel pdiffusion 668 -467 668 -467 0 feedthrough
rlabel pdiffusion 675 -467 675 -467 0 feedthrough
rlabel pdiffusion 682 -467 682 -467 0 feedthrough
rlabel pdiffusion 689 -467 689 -467 0 feedthrough
rlabel pdiffusion 696 -467 696 -467 0 feedthrough
rlabel pdiffusion 703 -467 703 -467 0 feedthrough
rlabel pdiffusion 710 -467 710 -467 0 feedthrough
rlabel pdiffusion 717 -467 717 -467 0 feedthrough
rlabel pdiffusion 724 -467 724 -467 0 feedthrough
rlabel pdiffusion 731 -467 731 -467 0 feedthrough
rlabel pdiffusion 738 -467 738 -467 0 feedthrough
rlabel pdiffusion 745 -467 745 -467 0 feedthrough
rlabel pdiffusion 752 -467 752 -467 0 feedthrough
rlabel pdiffusion 759 -467 759 -467 0 feedthrough
rlabel pdiffusion 766 -467 766 -467 0 feedthrough
rlabel pdiffusion 773 -467 773 -467 0 feedthrough
rlabel pdiffusion 780 -467 780 -467 0 feedthrough
rlabel pdiffusion 787 -467 787 -467 0 feedthrough
rlabel pdiffusion 794 -467 794 -467 0 feedthrough
rlabel pdiffusion 801 -467 801 -467 0 feedthrough
rlabel pdiffusion 808 -467 808 -467 0 feedthrough
rlabel pdiffusion 815 -467 815 -467 0 feedthrough
rlabel pdiffusion 822 -467 822 -467 0 feedthrough
rlabel pdiffusion 829 -467 829 -467 0 feedthrough
rlabel pdiffusion 836 -467 836 -467 0 feedthrough
rlabel pdiffusion 843 -467 843 -467 0 feedthrough
rlabel pdiffusion 850 -467 850 -467 0 feedthrough
rlabel pdiffusion 857 -467 857 -467 0 feedthrough
rlabel pdiffusion 864 -467 864 -467 0 feedthrough
rlabel pdiffusion 871 -467 871 -467 0 feedthrough
rlabel pdiffusion 878 -467 878 -467 0 feedthrough
rlabel pdiffusion 885 -467 885 -467 0 feedthrough
rlabel pdiffusion 892 -467 892 -467 0 feedthrough
rlabel pdiffusion 899 -467 899 -467 0 feedthrough
rlabel pdiffusion 906 -467 906 -467 0 feedthrough
rlabel pdiffusion 913 -467 913 -467 0 feedthrough
rlabel pdiffusion 920 -467 920 -467 0 feedthrough
rlabel pdiffusion 927 -467 927 -467 0 feedthrough
rlabel pdiffusion 934 -467 934 -467 0 feedthrough
rlabel pdiffusion 941 -467 941 -467 0 feedthrough
rlabel pdiffusion 948 -467 948 -467 0 feedthrough
rlabel pdiffusion 3 -554 3 -554 0 feedthrough
rlabel pdiffusion 10 -554 10 -554 0 feedthrough
rlabel pdiffusion 17 -554 17 -554 0 feedthrough
rlabel pdiffusion 24 -554 24 -554 0 cellNo=985
rlabel pdiffusion 31 -554 31 -554 0 feedthrough
rlabel pdiffusion 38 -554 38 -554 0 feedthrough
rlabel pdiffusion 45 -554 45 -554 0 cellNo=397
rlabel pdiffusion 52 -554 52 -554 0 feedthrough
rlabel pdiffusion 59 -554 59 -554 0 feedthrough
rlabel pdiffusion 66 -554 66 -554 0 feedthrough
rlabel pdiffusion 73 -554 73 -554 0 feedthrough
rlabel pdiffusion 80 -554 80 -554 0 feedthrough
rlabel pdiffusion 87 -554 87 -554 0 feedthrough
rlabel pdiffusion 94 -554 94 -554 0 cellNo=672
rlabel pdiffusion 101 -554 101 -554 0 feedthrough
rlabel pdiffusion 108 -554 108 -554 0 feedthrough
rlabel pdiffusion 115 -554 115 -554 0 feedthrough
rlabel pdiffusion 122 -554 122 -554 0 feedthrough
rlabel pdiffusion 129 -554 129 -554 0 feedthrough
rlabel pdiffusion 136 -554 136 -554 0 feedthrough
rlabel pdiffusion 143 -554 143 -554 0 cellNo=845
rlabel pdiffusion 150 -554 150 -554 0 feedthrough
rlabel pdiffusion 157 -554 157 -554 0 cellNo=77
rlabel pdiffusion 164 -554 164 -554 0 cellNo=158
rlabel pdiffusion 171 -554 171 -554 0 feedthrough
rlabel pdiffusion 178 -554 178 -554 0 cellNo=610
rlabel pdiffusion 185 -554 185 -554 0 feedthrough
rlabel pdiffusion 192 -554 192 -554 0 feedthrough
rlabel pdiffusion 199 -554 199 -554 0 feedthrough
rlabel pdiffusion 206 -554 206 -554 0 cellNo=76
rlabel pdiffusion 213 -554 213 -554 0 cellNo=414
rlabel pdiffusion 220 -554 220 -554 0 feedthrough
rlabel pdiffusion 227 -554 227 -554 0 feedthrough
rlabel pdiffusion 234 -554 234 -554 0 feedthrough
rlabel pdiffusion 241 -554 241 -554 0 cellNo=589
rlabel pdiffusion 248 -554 248 -554 0 feedthrough
rlabel pdiffusion 255 -554 255 -554 0 feedthrough
rlabel pdiffusion 262 -554 262 -554 0 cellNo=4
rlabel pdiffusion 269 -554 269 -554 0 feedthrough
rlabel pdiffusion 276 -554 276 -554 0 feedthrough
rlabel pdiffusion 283 -554 283 -554 0 feedthrough
rlabel pdiffusion 290 -554 290 -554 0 feedthrough
rlabel pdiffusion 297 -554 297 -554 0 feedthrough
rlabel pdiffusion 304 -554 304 -554 0 feedthrough
rlabel pdiffusion 311 -554 311 -554 0 cellNo=239
rlabel pdiffusion 318 -554 318 -554 0 cellNo=562
rlabel pdiffusion 325 -554 325 -554 0 feedthrough
rlabel pdiffusion 332 -554 332 -554 0 cellNo=284
rlabel pdiffusion 339 -554 339 -554 0 cellNo=690
rlabel pdiffusion 346 -554 346 -554 0 feedthrough
rlabel pdiffusion 353 -554 353 -554 0 feedthrough
rlabel pdiffusion 360 -554 360 -554 0 cellNo=586
rlabel pdiffusion 367 -554 367 -554 0 feedthrough
rlabel pdiffusion 374 -554 374 -554 0 feedthrough
rlabel pdiffusion 381 -554 381 -554 0 feedthrough
rlabel pdiffusion 388 -554 388 -554 0 cellNo=187
rlabel pdiffusion 395 -554 395 -554 0 feedthrough
rlabel pdiffusion 402 -554 402 -554 0 feedthrough
rlabel pdiffusion 409 -554 409 -554 0 feedthrough
rlabel pdiffusion 416 -554 416 -554 0 cellNo=212
rlabel pdiffusion 423 -554 423 -554 0 cellNo=79
rlabel pdiffusion 430 -554 430 -554 0 feedthrough
rlabel pdiffusion 437 -554 437 -554 0 feedthrough
rlabel pdiffusion 444 -554 444 -554 0 feedthrough
rlabel pdiffusion 451 -554 451 -554 0 cellNo=658
rlabel pdiffusion 458 -554 458 -554 0 feedthrough
rlabel pdiffusion 465 -554 465 -554 0 feedthrough
rlabel pdiffusion 472 -554 472 -554 0 feedthrough
rlabel pdiffusion 479 -554 479 -554 0 cellNo=596
rlabel pdiffusion 486 -554 486 -554 0 feedthrough
rlabel pdiffusion 493 -554 493 -554 0 cellNo=591
rlabel pdiffusion 500 -554 500 -554 0 cellNo=349
rlabel pdiffusion 507 -554 507 -554 0 cellNo=385
rlabel pdiffusion 514 -554 514 -554 0 feedthrough
rlabel pdiffusion 521 -554 521 -554 0 cellNo=47
rlabel pdiffusion 528 -554 528 -554 0 feedthrough
rlabel pdiffusion 535 -554 535 -554 0 feedthrough
rlabel pdiffusion 542 -554 542 -554 0 cellNo=548
rlabel pdiffusion 549 -554 549 -554 0 feedthrough
rlabel pdiffusion 556 -554 556 -554 0 feedthrough
rlabel pdiffusion 563 -554 563 -554 0 feedthrough
rlabel pdiffusion 570 -554 570 -554 0 feedthrough
rlabel pdiffusion 577 -554 577 -554 0 feedthrough
rlabel pdiffusion 584 -554 584 -554 0 feedthrough
rlabel pdiffusion 591 -554 591 -554 0 feedthrough
rlabel pdiffusion 598 -554 598 -554 0 feedthrough
rlabel pdiffusion 605 -554 605 -554 0 cellNo=726
rlabel pdiffusion 612 -554 612 -554 0 feedthrough
rlabel pdiffusion 619 -554 619 -554 0 feedthrough
rlabel pdiffusion 626 -554 626 -554 0 feedthrough
rlabel pdiffusion 633 -554 633 -554 0 feedthrough
rlabel pdiffusion 640 -554 640 -554 0 feedthrough
rlabel pdiffusion 647 -554 647 -554 0 cellNo=492
rlabel pdiffusion 654 -554 654 -554 0 feedthrough
rlabel pdiffusion 661 -554 661 -554 0 feedthrough
rlabel pdiffusion 668 -554 668 -554 0 feedthrough
rlabel pdiffusion 675 -554 675 -554 0 feedthrough
rlabel pdiffusion 682 -554 682 -554 0 feedthrough
rlabel pdiffusion 689 -554 689 -554 0 feedthrough
rlabel pdiffusion 696 -554 696 -554 0 feedthrough
rlabel pdiffusion 703 -554 703 -554 0 feedthrough
rlabel pdiffusion 710 -554 710 -554 0 feedthrough
rlabel pdiffusion 717 -554 717 -554 0 feedthrough
rlabel pdiffusion 724 -554 724 -554 0 cellNo=568
rlabel pdiffusion 731 -554 731 -554 0 feedthrough
rlabel pdiffusion 738 -554 738 -554 0 feedthrough
rlabel pdiffusion 745 -554 745 -554 0 feedthrough
rlabel pdiffusion 752 -554 752 -554 0 cellNo=810
rlabel pdiffusion 759 -554 759 -554 0 feedthrough
rlabel pdiffusion 766 -554 766 -554 0 feedthrough
rlabel pdiffusion 773 -554 773 -554 0 feedthrough
rlabel pdiffusion 780 -554 780 -554 0 feedthrough
rlabel pdiffusion 787 -554 787 -554 0 feedthrough
rlabel pdiffusion 794 -554 794 -554 0 cellNo=168
rlabel pdiffusion 801 -554 801 -554 0 feedthrough
rlabel pdiffusion 808 -554 808 -554 0 feedthrough
rlabel pdiffusion 815 -554 815 -554 0 feedthrough
rlabel pdiffusion 822 -554 822 -554 0 feedthrough
rlabel pdiffusion 836 -554 836 -554 0 feedthrough
rlabel pdiffusion 857 -554 857 -554 0 feedthrough
rlabel pdiffusion 3 -637 3 -637 0 feedthrough
rlabel pdiffusion 10 -637 10 -637 0 feedthrough
rlabel pdiffusion 17 -637 17 -637 0 feedthrough
rlabel pdiffusion 24 -637 24 -637 0 feedthrough
rlabel pdiffusion 31 -637 31 -637 0 feedthrough
rlabel pdiffusion 38 -637 38 -637 0 cellNo=61
rlabel pdiffusion 45 -637 45 -637 0 feedthrough
rlabel pdiffusion 52 -637 52 -637 0 feedthrough
rlabel pdiffusion 59 -637 59 -637 0 cellNo=510
rlabel pdiffusion 66 -637 66 -637 0 feedthrough
rlabel pdiffusion 73 -637 73 -637 0 feedthrough
rlabel pdiffusion 80 -637 80 -637 0 feedthrough
rlabel pdiffusion 87 -637 87 -637 0 cellNo=357
rlabel pdiffusion 94 -637 94 -637 0 feedthrough
rlabel pdiffusion 101 -637 101 -637 0 cellNo=409
rlabel pdiffusion 108 -637 108 -637 0 feedthrough
rlabel pdiffusion 115 -637 115 -637 0 feedthrough
rlabel pdiffusion 122 -637 122 -637 0 cellNo=162
rlabel pdiffusion 129 -637 129 -637 0 cellNo=715
rlabel pdiffusion 136 -637 136 -637 0 cellNo=222
rlabel pdiffusion 143 -637 143 -637 0 cellNo=176
rlabel pdiffusion 150 -637 150 -637 0 feedthrough
rlabel pdiffusion 157 -637 157 -637 0 feedthrough
rlabel pdiffusion 164 -637 164 -637 0 feedthrough
rlabel pdiffusion 171 -637 171 -637 0 cellNo=237
rlabel pdiffusion 178 -637 178 -637 0 feedthrough
rlabel pdiffusion 185 -637 185 -637 0 feedthrough
rlabel pdiffusion 192 -637 192 -637 0 feedthrough
rlabel pdiffusion 199 -637 199 -637 0 feedthrough
rlabel pdiffusion 206 -637 206 -637 0 feedthrough
rlabel pdiffusion 213 -637 213 -637 0 cellNo=769
rlabel pdiffusion 220 -637 220 -637 0 feedthrough
rlabel pdiffusion 227 -637 227 -637 0 cellNo=180
rlabel pdiffusion 234 -637 234 -637 0 cellNo=854
rlabel pdiffusion 241 -637 241 -637 0 cellNo=446
rlabel pdiffusion 248 -637 248 -637 0 feedthrough
rlabel pdiffusion 255 -637 255 -637 0 feedthrough
rlabel pdiffusion 262 -637 262 -637 0 feedthrough
rlabel pdiffusion 269 -637 269 -637 0 feedthrough
rlabel pdiffusion 276 -637 276 -637 0 feedthrough
rlabel pdiffusion 283 -637 283 -637 0 feedthrough
rlabel pdiffusion 290 -637 290 -637 0 feedthrough
rlabel pdiffusion 297 -637 297 -637 0 feedthrough
rlabel pdiffusion 304 -637 304 -637 0 cellNo=532
rlabel pdiffusion 311 -637 311 -637 0 cellNo=752
rlabel pdiffusion 318 -637 318 -637 0 feedthrough
rlabel pdiffusion 325 -637 325 -637 0 feedthrough
rlabel pdiffusion 332 -637 332 -637 0 cellNo=370
rlabel pdiffusion 339 -637 339 -637 0 cellNo=296
rlabel pdiffusion 346 -637 346 -637 0 cellNo=910
rlabel pdiffusion 353 -637 353 -637 0 feedthrough
rlabel pdiffusion 360 -637 360 -637 0 feedthrough
rlabel pdiffusion 367 -637 367 -637 0 feedthrough
rlabel pdiffusion 374 -637 374 -637 0 feedthrough
rlabel pdiffusion 381 -637 381 -637 0 feedthrough
rlabel pdiffusion 388 -637 388 -637 0 feedthrough
rlabel pdiffusion 395 -637 395 -637 0 feedthrough
rlabel pdiffusion 402 -637 402 -637 0 cellNo=630
rlabel pdiffusion 409 -637 409 -637 0 feedthrough
rlabel pdiffusion 416 -637 416 -637 0 feedthrough
rlabel pdiffusion 423 -637 423 -637 0 feedthrough
rlabel pdiffusion 430 -637 430 -637 0 feedthrough
rlabel pdiffusion 437 -637 437 -637 0 feedthrough
rlabel pdiffusion 444 -637 444 -637 0 feedthrough
rlabel pdiffusion 451 -637 451 -637 0 cellNo=33
rlabel pdiffusion 458 -637 458 -637 0 feedthrough
rlabel pdiffusion 465 -637 465 -637 0 cellNo=584
rlabel pdiffusion 472 -637 472 -637 0 cellNo=537
rlabel pdiffusion 479 -637 479 -637 0 feedthrough
rlabel pdiffusion 486 -637 486 -637 0 feedthrough
rlabel pdiffusion 493 -637 493 -637 0 feedthrough
rlabel pdiffusion 500 -637 500 -637 0 feedthrough
rlabel pdiffusion 507 -637 507 -637 0 feedthrough
rlabel pdiffusion 514 -637 514 -637 0 feedthrough
rlabel pdiffusion 521 -637 521 -637 0 cellNo=686
rlabel pdiffusion 528 -637 528 -637 0 feedthrough
rlabel pdiffusion 535 -637 535 -637 0 cellNo=805
rlabel pdiffusion 542 -637 542 -637 0 cellNo=758
rlabel pdiffusion 549 -637 549 -637 0 feedthrough
rlabel pdiffusion 556 -637 556 -637 0 feedthrough
rlabel pdiffusion 563 -637 563 -637 0 feedthrough
rlabel pdiffusion 570 -637 570 -637 0 feedthrough
rlabel pdiffusion 577 -637 577 -637 0 feedthrough
rlabel pdiffusion 584 -637 584 -637 0 feedthrough
rlabel pdiffusion 591 -637 591 -637 0 cellNo=269
rlabel pdiffusion 598 -637 598 -637 0 cellNo=318
rlabel pdiffusion 605 -637 605 -637 0 feedthrough
rlabel pdiffusion 612 -637 612 -637 0 cellNo=962
rlabel pdiffusion 619 -637 619 -637 0 cellNo=551
rlabel pdiffusion 626 -637 626 -637 0 feedthrough
rlabel pdiffusion 633 -637 633 -637 0 feedthrough
rlabel pdiffusion 640 -637 640 -637 0 feedthrough
rlabel pdiffusion 647 -637 647 -637 0 feedthrough
rlabel pdiffusion 654 -637 654 -637 0 feedthrough
rlabel pdiffusion 661 -637 661 -637 0 feedthrough
rlabel pdiffusion 668 -637 668 -637 0 feedthrough
rlabel pdiffusion 675 -637 675 -637 0 feedthrough
rlabel pdiffusion 682 -637 682 -637 0 feedthrough
rlabel pdiffusion 689 -637 689 -637 0 feedthrough
rlabel pdiffusion 696 -637 696 -637 0 cellNo=235
rlabel pdiffusion 703 -637 703 -637 0 feedthrough
rlabel pdiffusion 710 -637 710 -637 0 feedthrough
rlabel pdiffusion 717 -637 717 -637 0 feedthrough
rlabel pdiffusion 724 -637 724 -637 0 feedthrough
rlabel pdiffusion 731 -637 731 -637 0 feedthrough
rlabel pdiffusion 738 -637 738 -637 0 feedthrough
rlabel pdiffusion 745 -637 745 -637 0 feedthrough
rlabel pdiffusion 752 -637 752 -637 0 feedthrough
rlabel pdiffusion 759 -637 759 -637 0 feedthrough
rlabel pdiffusion 766 -637 766 -637 0 feedthrough
rlabel pdiffusion 773 -637 773 -637 0 feedthrough
rlabel pdiffusion 780 -637 780 -637 0 feedthrough
rlabel pdiffusion 787 -637 787 -637 0 feedthrough
rlabel pdiffusion 794 -637 794 -637 0 feedthrough
rlabel pdiffusion 801 -637 801 -637 0 feedthrough
rlabel pdiffusion 808 -637 808 -637 0 feedthrough
rlabel pdiffusion 815 -637 815 -637 0 feedthrough
rlabel pdiffusion 822 -637 822 -637 0 feedthrough
rlabel pdiffusion 829 -637 829 -637 0 feedthrough
rlabel pdiffusion 836 -637 836 -637 0 feedthrough
rlabel pdiffusion 843 -637 843 -637 0 feedthrough
rlabel pdiffusion 850 -637 850 -637 0 feedthrough
rlabel pdiffusion 857 -637 857 -637 0 feedthrough
rlabel pdiffusion 864 -637 864 -637 0 feedthrough
rlabel pdiffusion 871 -637 871 -637 0 feedthrough
rlabel pdiffusion 878 -637 878 -637 0 feedthrough
rlabel pdiffusion 885 -637 885 -637 0 feedthrough
rlabel pdiffusion 892 -637 892 -637 0 feedthrough
rlabel pdiffusion 899 -637 899 -637 0 feedthrough
rlabel pdiffusion 906 -637 906 -637 0 feedthrough
rlabel pdiffusion 913 -637 913 -637 0 feedthrough
rlabel pdiffusion 920 -637 920 -637 0 cellNo=136
rlabel pdiffusion 927 -637 927 -637 0 feedthrough
rlabel pdiffusion 948 -637 948 -637 0 feedthrough
rlabel pdiffusion 3 -716 3 -716 0 feedthrough
rlabel pdiffusion 10 -716 10 -716 0 feedthrough
rlabel pdiffusion 17 -716 17 -716 0 feedthrough
rlabel pdiffusion 24 -716 24 -716 0 cellNo=683
rlabel pdiffusion 31 -716 31 -716 0 cellNo=563
rlabel pdiffusion 38 -716 38 -716 0 feedthrough
rlabel pdiffusion 45 -716 45 -716 0 feedthrough
rlabel pdiffusion 52 -716 52 -716 0 feedthrough
rlabel pdiffusion 59 -716 59 -716 0 feedthrough
rlabel pdiffusion 66 -716 66 -716 0 feedthrough
rlabel pdiffusion 73 -716 73 -716 0 feedthrough
rlabel pdiffusion 80 -716 80 -716 0 feedthrough
rlabel pdiffusion 87 -716 87 -716 0 cellNo=979
rlabel pdiffusion 94 -716 94 -716 0 feedthrough
rlabel pdiffusion 101 -716 101 -716 0 cellNo=30
rlabel pdiffusion 108 -716 108 -716 0 cellNo=677
rlabel pdiffusion 115 -716 115 -716 0 feedthrough
rlabel pdiffusion 122 -716 122 -716 0 feedthrough
rlabel pdiffusion 129 -716 129 -716 0 cellNo=989
rlabel pdiffusion 136 -716 136 -716 0 feedthrough
rlabel pdiffusion 143 -716 143 -716 0 cellNo=459
rlabel pdiffusion 150 -716 150 -716 0 feedthrough
rlabel pdiffusion 157 -716 157 -716 0 feedthrough
rlabel pdiffusion 164 -716 164 -716 0 feedthrough
rlabel pdiffusion 171 -716 171 -716 0 feedthrough
rlabel pdiffusion 178 -716 178 -716 0 feedthrough
rlabel pdiffusion 185 -716 185 -716 0 feedthrough
rlabel pdiffusion 192 -716 192 -716 0 feedthrough
rlabel pdiffusion 199 -716 199 -716 0 feedthrough
rlabel pdiffusion 206 -716 206 -716 0 cellNo=326
rlabel pdiffusion 213 -716 213 -716 0 cellNo=333
rlabel pdiffusion 220 -716 220 -716 0 feedthrough
rlabel pdiffusion 227 -716 227 -716 0 cellNo=315
rlabel pdiffusion 234 -716 234 -716 0 feedthrough
rlabel pdiffusion 241 -716 241 -716 0 cellNo=410
rlabel pdiffusion 248 -716 248 -716 0 cellNo=11
rlabel pdiffusion 255 -716 255 -716 0 feedthrough
rlabel pdiffusion 262 -716 262 -716 0 feedthrough
rlabel pdiffusion 269 -716 269 -716 0 feedthrough
rlabel pdiffusion 276 -716 276 -716 0 cellNo=835
rlabel pdiffusion 283 -716 283 -716 0 feedthrough
rlabel pdiffusion 290 -716 290 -716 0 feedthrough
rlabel pdiffusion 297 -716 297 -716 0 feedthrough
rlabel pdiffusion 304 -716 304 -716 0 feedthrough
rlabel pdiffusion 311 -716 311 -716 0 feedthrough
rlabel pdiffusion 318 -716 318 -716 0 feedthrough
rlabel pdiffusion 325 -716 325 -716 0 feedthrough
rlabel pdiffusion 332 -716 332 -716 0 cellNo=540
rlabel pdiffusion 339 -716 339 -716 0 feedthrough
rlabel pdiffusion 346 -716 346 -716 0 cellNo=72
rlabel pdiffusion 353 -716 353 -716 0 feedthrough
rlabel pdiffusion 360 -716 360 -716 0 feedthrough
rlabel pdiffusion 367 -716 367 -716 0 feedthrough
rlabel pdiffusion 374 -716 374 -716 0 cellNo=485
rlabel pdiffusion 381 -716 381 -716 0 feedthrough
rlabel pdiffusion 388 -716 388 -716 0 cellNo=308
rlabel pdiffusion 395 -716 395 -716 0 cellNo=147
rlabel pdiffusion 402 -716 402 -716 0 feedthrough
rlabel pdiffusion 409 -716 409 -716 0 cellNo=862
rlabel pdiffusion 416 -716 416 -716 0 cellNo=502
rlabel pdiffusion 423 -716 423 -716 0 feedthrough
rlabel pdiffusion 430 -716 430 -716 0 feedthrough
rlabel pdiffusion 437 -716 437 -716 0 feedthrough
rlabel pdiffusion 444 -716 444 -716 0 feedthrough
rlabel pdiffusion 451 -716 451 -716 0 feedthrough
rlabel pdiffusion 458 -716 458 -716 0 feedthrough
rlabel pdiffusion 465 -716 465 -716 0 feedthrough
rlabel pdiffusion 472 -716 472 -716 0 cellNo=521
rlabel pdiffusion 479 -716 479 -716 0 cellNo=378
rlabel pdiffusion 486 -716 486 -716 0 cellNo=208
rlabel pdiffusion 493 -716 493 -716 0 feedthrough
rlabel pdiffusion 500 -716 500 -716 0 cellNo=243
rlabel pdiffusion 507 -716 507 -716 0 feedthrough
rlabel pdiffusion 514 -716 514 -716 0 cellNo=738
rlabel pdiffusion 521 -716 521 -716 0 feedthrough
rlabel pdiffusion 528 -716 528 -716 0 feedthrough
rlabel pdiffusion 535 -716 535 -716 0 feedthrough
rlabel pdiffusion 542 -716 542 -716 0 cellNo=325
rlabel pdiffusion 549 -716 549 -716 0 cellNo=939
rlabel pdiffusion 556 -716 556 -716 0 cellNo=276
rlabel pdiffusion 563 -716 563 -716 0 cellNo=227
rlabel pdiffusion 570 -716 570 -716 0 feedthrough
rlabel pdiffusion 577 -716 577 -716 0 feedthrough
rlabel pdiffusion 584 -716 584 -716 0 feedthrough
rlabel pdiffusion 591 -716 591 -716 0 cellNo=135
rlabel pdiffusion 598 -716 598 -716 0 feedthrough
rlabel pdiffusion 605 -716 605 -716 0 feedthrough
rlabel pdiffusion 612 -716 612 -716 0 feedthrough
rlabel pdiffusion 619 -716 619 -716 0 feedthrough
rlabel pdiffusion 626 -716 626 -716 0 cellNo=790
rlabel pdiffusion 633 -716 633 -716 0 feedthrough
rlabel pdiffusion 640 -716 640 -716 0 feedthrough
rlabel pdiffusion 647 -716 647 -716 0 feedthrough
rlabel pdiffusion 654 -716 654 -716 0 feedthrough
rlabel pdiffusion 661 -716 661 -716 0 feedthrough
rlabel pdiffusion 668 -716 668 -716 0 feedthrough
rlabel pdiffusion 675 -716 675 -716 0 feedthrough
rlabel pdiffusion 682 -716 682 -716 0 feedthrough
rlabel pdiffusion 689 -716 689 -716 0 feedthrough
rlabel pdiffusion 696 -716 696 -716 0 feedthrough
rlabel pdiffusion 703 -716 703 -716 0 feedthrough
rlabel pdiffusion 710 -716 710 -716 0 feedthrough
rlabel pdiffusion 717 -716 717 -716 0 feedthrough
rlabel pdiffusion 724 -716 724 -716 0 feedthrough
rlabel pdiffusion 731 -716 731 -716 0 feedthrough
rlabel pdiffusion 738 -716 738 -716 0 feedthrough
rlabel pdiffusion 745 -716 745 -716 0 feedthrough
rlabel pdiffusion 752 -716 752 -716 0 feedthrough
rlabel pdiffusion 759 -716 759 -716 0 feedthrough
rlabel pdiffusion 766 -716 766 -716 0 feedthrough
rlabel pdiffusion 773 -716 773 -716 0 feedthrough
rlabel pdiffusion 780 -716 780 -716 0 feedthrough
rlabel pdiffusion 787 -716 787 -716 0 feedthrough
rlabel pdiffusion 794 -716 794 -716 0 feedthrough
rlabel pdiffusion 801 -716 801 -716 0 feedthrough
rlabel pdiffusion 808 -716 808 -716 0 feedthrough
rlabel pdiffusion 815 -716 815 -716 0 feedthrough
rlabel pdiffusion 822 -716 822 -716 0 feedthrough
rlabel pdiffusion 829 -716 829 -716 0 feedthrough
rlabel pdiffusion 836 -716 836 -716 0 feedthrough
rlabel pdiffusion 843 -716 843 -716 0 feedthrough
rlabel pdiffusion 850 -716 850 -716 0 feedthrough
rlabel pdiffusion 857 -716 857 -716 0 feedthrough
rlabel pdiffusion 864 -716 864 -716 0 feedthrough
rlabel pdiffusion 871 -716 871 -716 0 feedthrough
rlabel pdiffusion 878 -716 878 -716 0 feedthrough
rlabel pdiffusion 885 -716 885 -716 0 cellNo=949
rlabel pdiffusion 892 -716 892 -716 0 feedthrough
rlabel pdiffusion 899 -716 899 -716 0 feedthrough
rlabel pdiffusion 906 -716 906 -716 0 feedthrough
rlabel pdiffusion 913 -716 913 -716 0 feedthrough
rlabel pdiffusion 920 -716 920 -716 0 feedthrough
rlabel pdiffusion 927 -716 927 -716 0 feedthrough
rlabel pdiffusion 955 -716 955 -716 0 feedthrough
rlabel pdiffusion 1032 -716 1032 -716 0 feedthrough
rlabel pdiffusion 24 -787 24 -787 0 feedthrough
rlabel pdiffusion 31 -787 31 -787 0 feedthrough
rlabel pdiffusion 38 -787 38 -787 0 feedthrough
rlabel pdiffusion 45 -787 45 -787 0 feedthrough
rlabel pdiffusion 52 -787 52 -787 0 cellNo=753
rlabel pdiffusion 59 -787 59 -787 0 feedthrough
rlabel pdiffusion 66 -787 66 -787 0 cellNo=351
rlabel pdiffusion 73 -787 73 -787 0 cellNo=662
rlabel pdiffusion 80 -787 80 -787 0 feedthrough
rlabel pdiffusion 87 -787 87 -787 0 feedthrough
rlabel pdiffusion 94 -787 94 -787 0 feedthrough
rlabel pdiffusion 101 -787 101 -787 0 feedthrough
rlabel pdiffusion 108 -787 108 -787 0 cellNo=671
rlabel pdiffusion 115 -787 115 -787 0 cellNo=146
rlabel pdiffusion 122 -787 122 -787 0 feedthrough
rlabel pdiffusion 129 -787 129 -787 0 feedthrough
rlabel pdiffusion 136 -787 136 -787 0 feedthrough
rlabel pdiffusion 143 -787 143 -787 0 feedthrough
rlabel pdiffusion 150 -787 150 -787 0 feedthrough
rlabel pdiffusion 157 -787 157 -787 0 feedthrough
rlabel pdiffusion 164 -787 164 -787 0 feedthrough
rlabel pdiffusion 171 -787 171 -787 0 feedthrough
rlabel pdiffusion 178 -787 178 -787 0 feedthrough
rlabel pdiffusion 185 -787 185 -787 0 cellNo=368
rlabel pdiffusion 192 -787 192 -787 0 feedthrough
rlabel pdiffusion 199 -787 199 -787 0 feedthrough
rlabel pdiffusion 206 -787 206 -787 0 feedthrough
rlabel pdiffusion 213 -787 213 -787 0 cellNo=97
rlabel pdiffusion 220 -787 220 -787 0 feedthrough
rlabel pdiffusion 227 -787 227 -787 0 cellNo=496
rlabel pdiffusion 234 -787 234 -787 0 cellNo=702
rlabel pdiffusion 241 -787 241 -787 0 cellNo=395
rlabel pdiffusion 248 -787 248 -787 0 feedthrough
rlabel pdiffusion 255 -787 255 -787 0 feedthrough
rlabel pdiffusion 262 -787 262 -787 0 cellNo=258
rlabel pdiffusion 269 -787 269 -787 0 feedthrough
rlabel pdiffusion 276 -787 276 -787 0 feedthrough
rlabel pdiffusion 283 -787 283 -787 0 feedthrough
rlabel pdiffusion 290 -787 290 -787 0 feedthrough
rlabel pdiffusion 297 -787 297 -787 0 feedthrough
rlabel pdiffusion 304 -787 304 -787 0 feedthrough
rlabel pdiffusion 311 -787 311 -787 0 cellNo=560
rlabel pdiffusion 318 -787 318 -787 0 feedthrough
rlabel pdiffusion 325 -787 325 -787 0 feedthrough
rlabel pdiffusion 332 -787 332 -787 0 feedthrough
rlabel pdiffusion 339 -787 339 -787 0 cellNo=261
rlabel pdiffusion 346 -787 346 -787 0 feedthrough
rlabel pdiffusion 353 -787 353 -787 0 cellNo=304
rlabel pdiffusion 360 -787 360 -787 0 feedthrough
rlabel pdiffusion 367 -787 367 -787 0 feedthrough
rlabel pdiffusion 374 -787 374 -787 0 cellNo=200
rlabel pdiffusion 381 -787 381 -787 0 feedthrough
rlabel pdiffusion 388 -787 388 -787 0 cellNo=140
rlabel pdiffusion 395 -787 395 -787 0 feedthrough
rlabel pdiffusion 402 -787 402 -787 0 cellNo=364
rlabel pdiffusion 409 -787 409 -787 0 feedthrough
rlabel pdiffusion 416 -787 416 -787 0 cellNo=566
rlabel pdiffusion 423 -787 423 -787 0 cellNo=973
rlabel pdiffusion 430 -787 430 -787 0 feedthrough
rlabel pdiffusion 437 -787 437 -787 0 feedthrough
rlabel pdiffusion 444 -787 444 -787 0 feedthrough
rlabel pdiffusion 451 -787 451 -787 0 feedthrough
rlabel pdiffusion 458 -787 458 -787 0 feedthrough
rlabel pdiffusion 465 -787 465 -787 0 feedthrough
rlabel pdiffusion 472 -787 472 -787 0 feedthrough
rlabel pdiffusion 479 -787 479 -787 0 feedthrough
rlabel pdiffusion 486 -787 486 -787 0 feedthrough
rlabel pdiffusion 493 -787 493 -787 0 cellNo=400
rlabel pdiffusion 500 -787 500 -787 0 feedthrough
rlabel pdiffusion 507 -787 507 -787 0 feedthrough
rlabel pdiffusion 514 -787 514 -787 0 cellNo=615
rlabel pdiffusion 521 -787 521 -787 0 feedthrough
rlabel pdiffusion 528 -787 528 -787 0 cellNo=866
rlabel pdiffusion 535 -787 535 -787 0 feedthrough
rlabel pdiffusion 542 -787 542 -787 0 cellNo=344
rlabel pdiffusion 549 -787 549 -787 0 feedthrough
rlabel pdiffusion 556 -787 556 -787 0 cellNo=234
rlabel pdiffusion 563 -787 563 -787 0 cellNo=172
rlabel pdiffusion 570 -787 570 -787 0 feedthrough
rlabel pdiffusion 577 -787 577 -787 0 cellNo=303
rlabel pdiffusion 584 -787 584 -787 0 feedthrough
rlabel pdiffusion 591 -787 591 -787 0 feedthrough
rlabel pdiffusion 598 -787 598 -787 0 feedthrough
rlabel pdiffusion 605 -787 605 -787 0 feedthrough
rlabel pdiffusion 612 -787 612 -787 0 feedthrough
rlabel pdiffusion 619 -787 619 -787 0 cellNo=389
rlabel pdiffusion 626 -787 626 -787 0 feedthrough
rlabel pdiffusion 633 -787 633 -787 0 feedthrough
rlabel pdiffusion 640 -787 640 -787 0 feedthrough
rlabel pdiffusion 647 -787 647 -787 0 feedthrough
rlabel pdiffusion 654 -787 654 -787 0 feedthrough
rlabel pdiffusion 661 -787 661 -787 0 feedthrough
rlabel pdiffusion 668 -787 668 -787 0 cellNo=815
rlabel pdiffusion 675 -787 675 -787 0 feedthrough
rlabel pdiffusion 682 -787 682 -787 0 feedthrough
rlabel pdiffusion 689 -787 689 -787 0 feedthrough
rlabel pdiffusion 696 -787 696 -787 0 feedthrough
rlabel pdiffusion 703 -787 703 -787 0 feedthrough
rlabel pdiffusion 710 -787 710 -787 0 feedthrough
rlabel pdiffusion 717 -787 717 -787 0 feedthrough
rlabel pdiffusion 724 -787 724 -787 0 feedthrough
rlabel pdiffusion 731 -787 731 -787 0 feedthrough
rlabel pdiffusion 738 -787 738 -787 0 feedthrough
rlabel pdiffusion 745 -787 745 -787 0 feedthrough
rlabel pdiffusion 752 -787 752 -787 0 feedthrough
rlabel pdiffusion 759 -787 759 -787 0 feedthrough
rlabel pdiffusion 766 -787 766 -787 0 feedthrough
rlabel pdiffusion 773 -787 773 -787 0 feedthrough
rlabel pdiffusion 780 -787 780 -787 0 feedthrough
rlabel pdiffusion 787 -787 787 -787 0 feedthrough
rlabel pdiffusion 794 -787 794 -787 0 feedthrough
rlabel pdiffusion 801 -787 801 -787 0 feedthrough
rlabel pdiffusion 808 -787 808 -787 0 feedthrough
rlabel pdiffusion 815 -787 815 -787 0 feedthrough
rlabel pdiffusion 822 -787 822 -787 0 feedthrough
rlabel pdiffusion 829 -787 829 -787 0 feedthrough
rlabel pdiffusion 836 -787 836 -787 0 feedthrough
rlabel pdiffusion 843 -787 843 -787 0 feedthrough
rlabel pdiffusion 850 -787 850 -787 0 feedthrough
rlabel pdiffusion 857 -787 857 -787 0 feedthrough
rlabel pdiffusion 864 -787 864 -787 0 feedthrough
rlabel pdiffusion 871 -787 871 -787 0 feedthrough
rlabel pdiffusion 878 -787 878 -787 0 feedthrough
rlabel pdiffusion 885 -787 885 -787 0 feedthrough
rlabel pdiffusion 892 -787 892 -787 0 cellNo=787
rlabel pdiffusion 899 -787 899 -787 0 feedthrough
rlabel pdiffusion 906 -787 906 -787 0 cellNo=402
rlabel pdiffusion 913 -787 913 -787 0 cellNo=360
rlabel pdiffusion 920 -787 920 -787 0 feedthrough
rlabel pdiffusion 962 -787 962 -787 0 feedthrough
rlabel pdiffusion 976 -787 976 -787 0 feedthrough
rlabel pdiffusion 990 -787 990 -787 0 cellNo=330
rlabel pdiffusion 1004 -787 1004 -787 0 cellNo=42
rlabel pdiffusion 1011 -787 1011 -787 0 feedthrough
rlabel pdiffusion 1018 -787 1018 -787 0 feedthrough
rlabel pdiffusion 1067 -787 1067 -787 0 feedthrough
rlabel pdiffusion 3 -884 3 -884 0 feedthrough
rlabel pdiffusion 10 -884 10 -884 0 cellNo=483
rlabel pdiffusion 17 -884 17 -884 0 feedthrough
rlabel pdiffusion 24 -884 24 -884 0 feedthrough
rlabel pdiffusion 31 -884 31 -884 0 feedthrough
rlabel pdiffusion 38 -884 38 -884 0 feedthrough
rlabel pdiffusion 45 -884 45 -884 0 cellNo=292
rlabel pdiffusion 52 -884 52 -884 0 feedthrough
rlabel pdiffusion 59 -884 59 -884 0 feedthrough
rlabel pdiffusion 66 -884 66 -884 0 cellNo=701
rlabel pdiffusion 73 -884 73 -884 0 feedthrough
rlabel pdiffusion 80 -884 80 -884 0 feedthrough
rlabel pdiffusion 87 -884 87 -884 0 feedthrough
rlabel pdiffusion 94 -884 94 -884 0 feedthrough
rlabel pdiffusion 101 -884 101 -884 0 feedthrough
rlabel pdiffusion 108 -884 108 -884 0 cellNo=655
rlabel pdiffusion 115 -884 115 -884 0 cellNo=71
rlabel pdiffusion 122 -884 122 -884 0 feedthrough
rlabel pdiffusion 129 -884 129 -884 0 cellNo=660
rlabel pdiffusion 136 -884 136 -884 0 cellNo=880
rlabel pdiffusion 143 -884 143 -884 0 feedthrough
rlabel pdiffusion 150 -884 150 -884 0 feedthrough
rlabel pdiffusion 157 -884 157 -884 0 feedthrough
rlabel pdiffusion 164 -884 164 -884 0 feedthrough
rlabel pdiffusion 171 -884 171 -884 0 cellNo=740
rlabel pdiffusion 178 -884 178 -884 0 cellNo=118
rlabel pdiffusion 185 -884 185 -884 0 feedthrough
rlabel pdiffusion 192 -884 192 -884 0 feedthrough
rlabel pdiffusion 199 -884 199 -884 0 feedthrough
rlabel pdiffusion 206 -884 206 -884 0 cellNo=909
rlabel pdiffusion 213 -884 213 -884 0 cellNo=38
rlabel pdiffusion 220 -884 220 -884 0 cellNo=53
rlabel pdiffusion 227 -884 227 -884 0 cellNo=881
rlabel pdiffusion 234 -884 234 -884 0 feedthrough
rlabel pdiffusion 241 -884 241 -884 0 cellNo=489
rlabel pdiffusion 248 -884 248 -884 0 feedthrough
rlabel pdiffusion 255 -884 255 -884 0 feedthrough
rlabel pdiffusion 262 -884 262 -884 0 feedthrough
rlabel pdiffusion 269 -884 269 -884 0 feedthrough
rlabel pdiffusion 276 -884 276 -884 0 feedthrough
rlabel pdiffusion 283 -884 283 -884 0 feedthrough
rlabel pdiffusion 290 -884 290 -884 0 feedthrough
rlabel pdiffusion 297 -884 297 -884 0 feedthrough
rlabel pdiffusion 304 -884 304 -884 0 feedthrough
rlabel pdiffusion 311 -884 311 -884 0 feedthrough
rlabel pdiffusion 318 -884 318 -884 0 feedthrough
rlabel pdiffusion 325 -884 325 -884 0 feedthrough
rlabel pdiffusion 332 -884 332 -884 0 feedthrough
rlabel pdiffusion 339 -884 339 -884 0 feedthrough
rlabel pdiffusion 346 -884 346 -884 0 feedthrough
rlabel pdiffusion 353 -884 353 -884 0 cellNo=594
rlabel pdiffusion 360 -884 360 -884 0 cellNo=832
rlabel pdiffusion 367 -884 367 -884 0 cellNo=514
rlabel pdiffusion 374 -884 374 -884 0 feedthrough
rlabel pdiffusion 381 -884 381 -884 0 feedthrough
rlabel pdiffusion 388 -884 388 -884 0 feedthrough
rlabel pdiffusion 395 -884 395 -884 0 feedthrough
rlabel pdiffusion 402 -884 402 -884 0 feedthrough
rlabel pdiffusion 409 -884 409 -884 0 cellNo=628
rlabel pdiffusion 416 -884 416 -884 0 cellNo=163
rlabel pdiffusion 423 -884 423 -884 0 feedthrough
rlabel pdiffusion 430 -884 430 -884 0 feedthrough
rlabel pdiffusion 437 -884 437 -884 0 cellNo=424
rlabel pdiffusion 444 -884 444 -884 0 feedthrough
rlabel pdiffusion 451 -884 451 -884 0 feedthrough
rlabel pdiffusion 458 -884 458 -884 0 feedthrough
rlabel pdiffusion 465 -884 465 -884 0 cellNo=536
rlabel pdiffusion 472 -884 472 -884 0 feedthrough
rlabel pdiffusion 479 -884 479 -884 0 feedthrough
rlabel pdiffusion 486 -884 486 -884 0 feedthrough
rlabel pdiffusion 493 -884 493 -884 0 cellNo=56
rlabel pdiffusion 500 -884 500 -884 0 cellNo=723
rlabel pdiffusion 507 -884 507 -884 0 feedthrough
rlabel pdiffusion 514 -884 514 -884 0 feedthrough
rlabel pdiffusion 521 -884 521 -884 0 cellNo=294
rlabel pdiffusion 528 -884 528 -884 0 feedthrough
rlabel pdiffusion 535 -884 535 -884 0 cellNo=337
rlabel pdiffusion 542 -884 542 -884 0 cellNo=974
rlabel pdiffusion 549 -884 549 -884 0 cellNo=848
rlabel pdiffusion 556 -884 556 -884 0 feedthrough
rlabel pdiffusion 563 -884 563 -884 0 cellNo=864
rlabel pdiffusion 570 -884 570 -884 0 cellNo=708
rlabel pdiffusion 577 -884 577 -884 0 feedthrough
rlabel pdiffusion 584 -884 584 -884 0 feedthrough
rlabel pdiffusion 591 -884 591 -884 0 feedthrough
rlabel pdiffusion 598 -884 598 -884 0 feedthrough
rlabel pdiffusion 605 -884 605 -884 0 feedthrough
rlabel pdiffusion 612 -884 612 -884 0 feedthrough
rlabel pdiffusion 619 -884 619 -884 0 feedthrough
rlabel pdiffusion 626 -884 626 -884 0 feedthrough
rlabel pdiffusion 633 -884 633 -884 0 feedthrough
rlabel pdiffusion 640 -884 640 -884 0 feedthrough
rlabel pdiffusion 647 -884 647 -884 0 feedthrough
rlabel pdiffusion 654 -884 654 -884 0 feedthrough
rlabel pdiffusion 661 -884 661 -884 0 feedthrough
rlabel pdiffusion 668 -884 668 -884 0 cellNo=558
rlabel pdiffusion 675 -884 675 -884 0 feedthrough
rlabel pdiffusion 682 -884 682 -884 0 feedthrough
rlabel pdiffusion 689 -884 689 -884 0 feedthrough
rlabel pdiffusion 696 -884 696 -884 0 feedthrough
rlabel pdiffusion 703 -884 703 -884 0 feedthrough
rlabel pdiffusion 710 -884 710 -884 0 feedthrough
rlabel pdiffusion 717 -884 717 -884 0 feedthrough
rlabel pdiffusion 724 -884 724 -884 0 feedthrough
rlabel pdiffusion 731 -884 731 -884 0 feedthrough
rlabel pdiffusion 738 -884 738 -884 0 feedthrough
rlabel pdiffusion 745 -884 745 -884 0 feedthrough
rlabel pdiffusion 752 -884 752 -884 0 feedthrough
rlabel pdiffusion 759 -884 759 -884 0 feedthrough
rlabel pdiffusion 766 -884 766 -884 0 feedthrough
rlabel pdiffusion 773 -884 773 -884 0 feedthrough
rlabel pdiffusion 780 -884 780 -884 0 feedthrough
rlabel pdiffusion 787 -884 787 -884 0 feedthrough
rlabel pdiffusion 794 -884 794 -884 0 feedthrough
rlabel pdiffusion 801 -884 801 -884 0 feedthrough
rlabel pdiffusion 808 -884 808 -884 0 feedthrough
rlabel pdiffusion 815 -884 815 -884 0 cellNo=804
rlabel pdiffusion 822 -884 822 -884 0 feedthrough
rlabel pdiffusion 829 -884 829 -884 0 feedthrough
rlabel pdiffusion 836 -884 836 -884 0 feedthrough
rlabel pdiffusion 843 -884 843 -884 0 feedthrough
rlabel pdiffusion 850 -884 850 -884 0 feedthrough
rlabel pdiffusion 857 -884 857 -884 0 feedthrough
rlabel pdiffusion 864 -884 864 -884 0 feedthrough
rlabel pdiffusion 871 -884 871 -884 0 feedthrough
rlabel pdiffusion 878 -884 878 -884 0 feedthrough
rlabel pdiffusion 885 -884 885 -884 0 feedthrough
rlabel pdiffusion 892 -884 892 -884 0 feedthrough
rlabel pdiffusion 899 -884 899 -884 0 feedthrough
rlabel pdiffusion 906 -884 906 -884 0 feedthrough
rlabel pdiffusion 913 -884 913 -884 0 feedthrough
rlabel pdiffusion 920 -884 920 -884 0 feedthrough
rlabel pdiffusion 927 -884 927 -884 0 feedthrough
rlabel pdiffusion 934 -884 934 -884 0 feedthrough
rlabel pdiffusion 941 -884 941 -884 0 feedthrough
rlabel pdiffusion 948 -884 948 -884 0 feedthrough
rlabel pdiffusion 955 -884 955 -884 0 feedthrough
rlabel pdiffusion 962 -884 962 -884 0 feedthrough
rlabel pdiffusion 969 -884 969 -884 0 feedthrough
rlabel pdiffusion 976 -884 976 -884 0 feedthrough
rlabel pdiffusion 983 -884 983 -884 0 feedthrough
rlabel pdiffusion 990 -884 990 -884 0 cellNo=122
rlabel pdiffusion 997 -884 997 -884 0 feedthrough
rlabel pdiffusion 1004 -884 1004 -884 0 feedthrough
rlabel pdiffusion 1011 -884 1011 -884 0 cellNo=943
rlabel pdiffusion 1018 -884 1018 -884 0 feedthrough
rlabel pdiffusion 1025 -884 1025 -884 0 feedthrough
rlabel pdiffusion 1039 -884 1039 -884 0 feedthrough
rlabel pdiffusion 1081 -884 1081 -884 0 feedthrough
rlabel pdiffusion 10 -965 10 -965 0 cellNo=457
rlabel pdiffusion 17 -965 17 -965 0 feedthrough
rlabel pdiffusion 24 -965 24 -965 0 feedthrough
rlabel pdiffusion 31 -965 31 -965 0 feedthrough
rlabel pdiffusion 38 -965 38 -965 0 feedthrough
rlabel pdiffusion 45 -965 45 -965 0 feedthrough
rlabel pdiffusion 52 -965 52 -965 0 feedthrough
rlabel pdiffusion 59 -965 59 -965 0 feedthrough
rlabel pdiffusion 66 -965 66 -965 0 feedthrough
rlabel pdiffusion 73 -965 73 -965 0 feedthrough
rlabel pdiffusion 80 -965 80 -965 0 feedthrough
rlabel pdiffusion 87 -965 87 -965 0 feedthrough
rlabel pdiffusion 94 -965 94 -965 0 feedthrough
rlabel pdiffusion 101 -965 101 -965 0 feedthrough
rlabel pdiffusion 108 -965 108 -965 0 feedthrough
rlabel pdiffusion 115 -965 115 -965 0 feedthrough
rlabel pdiffusion 122 -965 122 -965 0 feedthrough
rlabel pdiffusion 129 -965 129 -965 0 cellNo=929
rlabel pdiffusion 136 -965 136 -965 0 feedthrough
rlabel pdiffusion 143 -965 143 -965 0 feedthrough
rlabel pdiffusion 150 -965 150 -965 0 feedthrough
rlabel pdiffusion 157 -965 157 -965 0 feedthrough
rlabel pdiffusion 164 -965 164 -965 0 feedthrough
rlabel pdiffusion 171 -965 171 -965 0 feedthrough
rlabel pdiffusion 178 -965 178 -965 0 cellNo=153
rlabel pdiffusion 185 -965 185 -965 0 feedthrough
rlabel pdiffusion 192 -965 192 -965 0 feedthrough
rlabel pdiffusion 199 -965 199 -965 0 feedthrough
rlabel pdiffusion 206 -965 206 -965 0 feedthrough
rlabel pdiffusion 213 -965 213 -965 0 cellNo=313
rlabel pdiffusion 220 -965 220 -965 0 cellNo=836
rlabel pdiffusion 227 -965 227 -965 0 cellNo=905
rlabel pdiffusion 234 -965 234 -965 0 cellNo=693
rlabel pdiffusion 241 -965 241 -965 0 cellNo=911
rlabel pdiffusion 248 -965 248 -965 0 feedthrough
rlabel pdiffusion 255 -965 255 -965 0 feedthrough
rlabel pdiffusion 262 -965 262 -965 0 feedthrough
rlabel pdiffusion 269 -965 269 -965 0 feedthrough
rlabel pdiffusion 276 -965 276 -965 0 cellNo=684
rlabel pdiffusion 283 -965 283 -965 0 cellNo=598
rlabel pdiffusion 290 -965 290 -965 0 feedthrough
rlabel pdiffusion 297 -965 297 -965 0 feedthrough
rlabel pdiffusion 304 -965 304 -965 0 feedthrough
rlabel pdiffusion 311 -965 311 -965 0 feedthrough
rlabel pdiffusion 318 -965 318 -965 0 feedthrough
rlabel pdiffusion 325 -965 325 -965 0 cellNo=914
rlabel pdiffusion 332 -965 332 -965 0 feedthrough
rlabel pdiffusion 339 -965 339 -965 0 feedthrough
rlabel pdiffusion 346 -965 346 -965 0 feedthrough
rlabel pdiffusion 353 -965 353 -965 0 feedthrough
rlabel pdiffusion 360 -965 360 -965 0 cellNo=906
rlabel pdiffusion 367 -965 367 -965 0 feedthrough
rlabel pdiffusion 374 -965 374 -965 0 feedthrough
rlabel pdiffusion 381 -965 381 -965 0 cellNo=211
rlabel pdiffusion 388 -965 388 -965 0 feedthrough
rlabel pdiffusion 395 -965 395 -965 0 cellNo=273
rlabel pdiffusion 402 -965 402 -965 0 feedthrough
rlabel pdiffusion 409 -965 409 -965 0 feedthrough
rlabel pdiffusion 416 -965 416 -965 0 cellNo=193
rlabel pdiffusion 423 -965 423 -965 0 feedthrough
rlabel pdiffusion 430 -965 430 -965 0 feedthrough
rlabel pdiffusion 437 -965 437 -965 0 cellNo=513
rlabel pdiffusion 444 -965 444 -965 0 feedthrough
rlabel pdiffusion 451 -965 451 -965 0 cellNo=340
rlabel pdiffusion 458 -965 458 -965 0 feedthrough
rlabel pdiffusion 465 -965 465 -965 0 feedthrough
rlabel pdiffusion 472 -965 472 -965 0 cellNo=245
rlabel pdiffusion 479 -965 479 -965 0 cellNo=636
rlabel pdiffusion 486 -965 486 -965 0 feedthrough
rlabel pdiffusion 493 -965 493 -965 0 cellNo=544
rlabel pdiffusion 500 -965 500 -965 0 feedthrough
rlabel pdiffusion 507 -965 507 -965 0 feedthrough
rlabel pdiffusion 514 -965 514 -965 0 cellNo=119
rlabel pdiffusion 521 -965 521 -965 0 feedthrough
rlabel pdiffusion 528 -965 528 -965 0 cellNo=583
rlabel pdiffusion 535 -965 535 -965 0 feedthrough
rlabel pdiffusion 542 -965 542 -965 0 feedthrough
rlabel pdiffusion 549 -965 549 -965 0 feedthrough
rlabel pdiffusion 556 -965 556 -965 0 feedthrough
rlabel pdiffusion 563 -965 563 -965 0 cellNo=279
rlabel pdiffusion 570 -965 570 -965 0 feedthrough
rlabel pdiffusion 577 -965 577 -965 0 feedthrough
rlabel pdiffusion 584 -965 584 -965 0 feedthrough
rlabel pdiffusion 591 -965 591 -965 0 feedthrough
rlabel pdiffusion 598 -965 598 -965 0 cellNo=640
rlabel pdiffusion 605 -965 605 -965 0 cellNo=130
rlabel pdiffusion 612 -965 612 -965 0 feedthrough
rlabel pdiffusion 619 -965 619 -965 0 cellNo=567
rlabel pdiffusion 626 -965 626 -965 0 cellNo=879
rlabel pdiffusion 633 -965 633 -965 0 cellNo=481
rlabel pdiffusion 640 -965 640 -965 0 feedthrough
rlabel pdiffusion 647 -965 647 -965 0 feedthrough
rlabel pdiffusion 654 -965 654 -965 0 cellNo=824
rlabel pdiffusion 661 -965 661 -965 0 feedthrough
rlabel pdiffusion 668 -965 668 -965 0 feedthrough
rlabel pdiffusion 675 -965 675 -965 0 feedthrough
rlabel pdiffusion 682 -965 682 -965 0 feedthrough
rlabel pdiffusion 689 -965 689 -965 0 feedthrough
rlabel pdiffusion 696 -965 696 -965 0 cellNo=432
rlabel pdiffusion 703 -965 703 -965 0 feedthrough
rlabel pdiffusion 710 -965 710 -965 0 feedthrough
rlabel pdiffusion 717 -965 717 -965 0 feedthrough
rlabel pdiffusion 724 -965 724 -965 0 feedthrough
rlabel pdiffusion 731 -965 731 -965 0 feedthrough
rlabel pdiffusion 738 -965 738 -965 0 feedthrough
rlabel pdiffusion 745 -965 745 -965 0 feedthrough
rlabel pdiffusion 752 -965 752 -965 0 feedthrough
rlabel pdiffusion 759 -965 759 -965 0 feedthrough
rlabel pdiffusion 766 -965 766 -965 0 feedthrough
rlabel pdiffusion 773 -965 773 -965 0 feedthrough
rlabel pdiffusion 780 -965 780 -965 0 feedthrough
rlabel pdiffusion 787 -965 787 -965 0 feedthrough
rlabel pdiffusion 794 -965 794 -965 0 feedthrough
rlabel pdiffusion 801 -965 801 -965 0 feedthrough
rlabel pdiffusion 808 -965 808 -965 0 feedthrough
rlabel pdiffusion 815 -965 815 -965 0 feedthrough
rlabel pdiffusion 822 -965 822 -965 0 feedthrough
rlabel pdiffusion 829 -965 829 -965 0 feedthrough
rlabel pdiffusion 836 -965 836 -965 0 feedthrough
rlabel pdiffusion 843 -965 843 -965 0 feedthrough
rlabel pdiffusion 850 -965 850 -965 0 feedthrough
rlabel pdiffusion 857 -965 857 -965 0 feedthrough
rlabel pdiffusion 864 -965 864 -965 0 feedthrough
rlabel pdiffusion 871 -965 871 -965 0 feedthrough
rlabel pdiffusion 878 -965 878 -965 0 feedthrough
rlabel pdiffusion 885 -965 885 -965 0 feedthrough
rlabel pdiffusion 892 -965 892 -965 0 feedthrough
rlabel pdiffusion 899 -965 899 -965 0 feedthrough
rlabel pdiffusion 906 -965 906 -965 0 feedthrough
rlabel pdiffusion 913 -965 913 -965 0 cellNo=252
rlabel pdiffusion 920 -965 920 -965 0 cellNo=613
rlabel pdiffusion 927 -965 927 -965 0 cellNo=837
rlabel pdiffusion 934 -965 934 -965 0 cellNo=983
rlabel pdiffusion 941 -965 941 -965 0 cellNo=467
rlabel pdiffusion 948 -965 948 -965 0 feedthrough
rlabel pdiffusion 955 -965 955 -965 0 feedthrough
rlabel pdiffusion 962 -965 962 -965 0 feedthrough
rlabel pdiffusion 969 -965 969 -965 0 feedthrough
rlabel pdiffusion 983 -965 983 -965 0 feedthrough
rlabel pdiffusion 1011 -965 1011 -965 0 feedthrough
rlabel pdiffusion 1039 -965 1039 -965 0 feedthrough
rlabel pdiffusion 1060 -965 1060 -965 0 feedthrough
rlabel pdiffusion 1088 -965 1088 -965 0 feedthrough
rlabel pdiffusion 10 -1058 10 -1058 0 feedthrough
rlabel pdiffusion 17 -1058 17 -1058 0 feedthrough
rlabel pdiffusion 24 -1058 24 -1058 0 feedthrough
rlabel pdiffusion 31 -1058 31 -1058 0 feedthrough
rlabel pdiffusion 38 -1058 38 -1058 0 cellNo=181
rlabel pdiffusion 45 -1058 45 -1058 0 feedthrough
rlabel pdiffusion 52 -1058 52 -1058 0 feedthrough
rlabel pdiffusion 59 -1058 59 -1058 0 cellNo=32
rlabel pdiffusion 66 -1058 66 -1058 0 feedthrough
rlabel pdiffusion 73 -1058 73 -1058 0 feedthrough
rlabel pdiffusion 80 -1058 80 -1058 0 feedthrough
rlabel pdiffusion 87 -1058 87 -1058 0 feedthrough
rlabel pdiffusion 94 -1058 94 -1058 0 feedthrough
rlabel pdiffusion 101 -1058 101 -1058 0 feedthrough
rlabel pdiffusion 108 -1058 108 -1058 0 feedthrough
rlabel pdiffusion 115 -1058 115 -1058 0 feedthrough
rlabel pdiffusion 122 -1058 122 -1058 0 feedthrough
rlabel pdiffusion 129 -1058 129 -1058 0 cellNo=538
rlabel pdiffusion 136 -1058 136 -1058 0 feedthrough
rlabel pdiffusion 143 -1058 143 -1058 0 cellNo=416
rlabel pdiffusion 150 -1058 150 -1058 0 feedthrough
rlabel pdiffusion 157 -1058 157 -1058 0 feedthrough
rlabel pdiffusion 164 -1058 164 -1058 0 cellNo=125
rlabel pdiffusion 171 -1058 171 -1058 0 cellNo=106
rlabel pdiffusion 178 -1058 178 -1058 0 cellNo=901
rlabel pdiffusion 185 -1058 185 -1058 0 feedthrough
rlabel pdiffusion 192 -1058 192 -1058 0 feedthrough
rlabel pdiffusion 199 -1058 199 -1058 0 feedthrough
rlabel pdiffusion 206 -1058 206 -1058 0 cellNo=470
rlabel pdiffusion 213 -1058 213 -1058 0 feedthrough
rlabel pdiffusion 220 -1058 220 -1058 0 cellNo=167
rlabel pdiffusion 227 -1058 227 -1058 0 feedthrough
rlabel pdiffusion 234 -1058 234 -1058 0 feedthrough
rlabel pdiffusion 241 -1058 241 -1058 0 feedthrough
rlabel pdiffusion 248 -1058 248 -1058 0 feedthrough
rlabel pdiffusion 255 -1058 255 -1058 0 cellNo=277
rlabel pdiffusion 262 -1058 262 -1058 0 feedthrough
rlabel pdiffusion 269 -1058 269 -1058 0 feedthrough
rlabel pdiffusion 276 -1058 276 -1058 0 feedthrough
rlabel pdiffusion 283 -1058 283 -1058 0 feedthrough
rlabel pdiffusion 290 -1058 290 -1058 0 feedthrough
rlabel pdiffusion 297 -1058 297 -1058 0 cellNo=85
rlabel pdiffusion 304 -1058 304 -1058 0 feedthrough
rlabel pdiffusion 311 -1058 311 -1058 0 feedthrough
rlabel pdiffusion 318 -1058 318 -1058 0 feedthrough
rlabel pdiffusion 325 -1058 325 -1058 0 feedthrough
rlabel pdiffusion 332 -1058 332 -1058 0 feedthrough
rlabel pdiffusion 339 -1058 339 -1058 0 feedthrough
rlabel pdiffusion 346 -1058 346 -1058 0 feedthrough
rlabel pdiffusion 353 -1058 353 -1058 0 cellNo=352
rlabel pdiffusion 360 -1058 360 -1058 0 feedthrough
rlabel pdiffusion 367 -1058 367 -1058 0 feedthrough
rlabel pdiffusion 374 -1058 374 -1058 0 feedthrough
rlabel pdiffusion 381 -1058 381 -1058 0 feedthrough
rlabel pdiffusion 388 -1058 388 -1058 0 feedthrough
rlabel pdiffusion 395 -1058 395 -1058 0 feedthrough
rlabel pdiffusion 402 -1058 402 -1058 0 feedthrough
rlabel pdiffusion 409 -1058 409 -1058 0 cellNo=827
rlabel pdiffusion 416 -1058 416 -1058 0 feedthrough
rlabel pdiffusion 423 -1058 423 -1058 0 feedthrough
rlabel pdiffusion 430 -1058 430 -1058 0 cellNo=884
rlabel pdiffusion 437 -1058 437 -1058 0 feedthrough
rlabel pdiffusion 444 -1058 444 -1058 0 cellNo=639
rlabel pdiffusion 451 -1058 451 -1058 0 cellNo=451
rlabel pdiffusion 458 -1058 458 -1058 0 feedthrough
rlabel pdiffusion 465 -1058 465 -1058 0 feedthrough
rlabel pdiffusion 472 -1058 472 -1058 0 cellNo=184
rlabel pdiffusion 479 -1058 479 -1058 0 cellNo=754
rlabel pdiffusion 486 -1058 486 -1058 0 cellNo=89
rlabel pdiffusion 493 -1058 493 -1058 0 cellNo=650
rlabel pdiffusion 500 -1058 500 -1058 0 feedthrough
rlabel pdiffusion 507 -1058 507 -1058 0 feedthrough
rlabel pdiffusion 514 -1058 514 -1058 0 cellNo=718
rlabel pdiffusion 521 -1058 521 -1058 0 feedthrough
rlabel pdiffusion 528 -1058 528 -1058 0 feedthrough
rlabel pdiffusion 535 -1058 535 -1058 0 cellNo=971
rlabel pdiffusion 542 -1058 542 -1058 0 feedthrough
rlabel pdiffusion 549 -1058 549 -1058 0 cellNo=417
rlabel pdiffusion 556 -1058 556 -1058 0 feedthrough
rlabel pdiffusion 563 -1058 563 -1058 0 feedthrough
rlabel pdiffusion 570 -1058 570 -1058 0 cellNo=681
rlabel pdiffusion 577 -1058 577 -1058 0 cellNo=539
rlabel pdiffusion 584 -1058 584 -1058 0 cellNo=498
rlabel pdiffusion 591 -1058 591 -1058 0 feedthrough
rlabel pdiffusion 598 -1058 598 -1058 0 feedthrough
rlabel pdiffusion 605 -1058 605 -1058 0 cellNo=590
rlabel pdiffusion 612 -1058 612 -1058 0 feedthrough
rlabel pdiffusion 619 -1058 619 -1058 0 feedthrough
rlabel pdiffusion 626 -1058 626 -1058 0 cellNo=182
rlabel pdiffusion 633 -1058 633 -1058 0 feedthrough
rlabel pdiffusion 640 -1058 640 -1058 0 feedthrough
rlabel pdiffusion 647 -1058 647 -1058 0 cellNo=88
rlabel pdiffusion 654 -1058 654 -1058 0 feedthrough
rlabel pdiffusion 661 -1058 661 -1058 0 feedthrough
rlabel pdiffusion 668 -1058 668 -1058 0 feedthrough
rlabel pdiffusion 675 -1058 675 -1058 0 feedthrough
rlabel pdiffusion 682 -1058 682 -1058 0 feedthrough
rlabel pdiffusion 689 -1058 689 -1058 0 cellNo=604
rlabel pdiffusion 696 -1058 696 -1058 0 feedthrough
rlabel pdiffusion 703 -1058 703 -1058 0 feedthrough
rlabel pdiffusion 710 -1058 710 -1058 0 feedthrough
rlabel pdiffusion 717 -1058 717 -1058 0 feedthrough
rlabel pdiffusion 724 -1058 724 -1058 0 feedthrough
rlabel pdiffusion 731 -1058 731 -1058 0 cellNo=666
rlabel pdiffusion 738 -1058 738 -1058 0 feedthrough
rlabel pdiffusion 745 -1058 745 -1058 0 feedthrough
rlabel pdiffusion 752 -1058 752 -1058 0 feedthrough
rlabel pdiffusion 759 -1058 759 -1058 0 feedthrough
rlabel pdiffusion 766 -1058 766 -1058 0 feedthrough
rlabel pdiffusion 773 -1058 773 -1058 0 feedthrough
rlabel pdiffusion 780 -1058 780 -1058 0 feedthrough
rlabel pdiffusion 787 -1058 787 -1058 0 feedthrough
rlabel pdiffusion 794 -1058 794 -1058 0 feedthrough
rlabel pdiffusion 801 -1058 801 -1058 0 feedthrough
rlabel pdiffusion 808 -1058 808 -1058 0 feedthrough
rlabel pdiffusion 815 -1058 815 -1058 0 feedthrough
rlabel pdiffusion 822 -1058 822 -1058 0 feedthrough
rlabel pdiffusion 829 -1058 829 -1058 0 feedthrough
rlabel pdiffusion 836 -1058 836 -1058 0 feedthrough
rlabel pdiffusion 843 -1058 843 -1058 0 feedthrough
rlabel pdiffusion 850 -1058 850 -1058 0 feedthrough
rlabel pdiffusion 857 -1058 857 -1058 0 feedthrough
rlabel pdiffusion 864 -1058 864 -1058 0 feedthrough
rlabel pdiffusion 871 -1058 871 -1058 0 feedthrough
rlabel pdiffusion 878 -1058 878 -1058 0 feedthrough
rlabel pdiffusion 885 -1058 885 -1058 0 feedthrough
rlabel pdiffusion 892 -1058 892 -1058 0 feedthrough
rlabel pdiffusion 899 -1058 899 -1058 0 feedthrough
rlabel pdiffusion 906 -1058 906 -1058 0 feedthrough
rlabel pdiffusion 913 -1058 913 -1058 0 feedthrough
rlabel pdiffusion 920 -1058 920 -1058 0 feedthrough
rlabel pdiffusion 927 -1058 927 -1058 0 feedthrough
rlabel pdiffusion 934 -1058 934 -1058 0 feedthrough
rlabel pdiffusion 941 -1058 941 -1058 0 feedthrough
rlabel pdiffusion 948 -1058 948 -1058 0 feedthrough
rlabel pdiffusion 955 -1058 955 -1058 0 feedthrough
rlabel pdiffusion 962 -1058 962 -1058 0 feedthrough
rlabel pdiffusion 969 -1058 969 -1058 0 feedthrough
rlabel pdiffusion 976 -1058 976 -1058 0 feedthrough
rlabel pdiffusion 983 -1058 983 -1058 0 feedthrough
rlabel pdiffusion 990 -1058 990 -1058 0 feedthrough
rlabel pdiffusion 997 -1058 997 -1058 0 feedthrough
rlabel pdiffusion 1004 -1058 1004 -1058 0 feedthrough
rlabel pdiffusion 1011 -1058 1011 -1058 0 feedthrough
rlabel pdiffusion 1018 -1058 1018 -1058 0 feedthrough
rlabel pdiffusion 1025 -1058 1025 -1058 0 cellNo=445
rlabel pdiffusion 1032 -1058 1032 -1058 0 feedthrough
rlabel pdiffusion 1039 -1058 1039 -1058 0 feedthrough
rlabel pdiffusion 1046 -1058 1046 -1058 0 feedthrough
rlabel pdiffusion 1053 -1058 1053 -1058 0 feedthrough
rlabel pdiffusion 1060 -1058 1060 -1058 0 feedthrough
rlabel pdiffusion 1067 -1058 1067 -1058 0 cellNo=197
rlabel pdiffusion 1074 -1058 1074 -1058 0 cellNo=812
rlabel pdiffusion 1081 -1058 1081 -1058 0 cellNo=447
rlabel pdiffusion 1088 -1058 1088 -1058 0 feedthrough
rlabel pdiffusion 1095 -1058 1095 -1058 0 feedthrough
rlabel pdiffusion 1102 -1058 1102 -1058 0 feedthrough
rlabel pdiffusion 3 -1157 3 -1157 0 feedthrough
rlabel pdiffusion 10 -1157 10 -1157 0 cellNo=453
rlabel pdiffusion 17 -1157 17 -1157 0 cellNo=747
rlabel pdiffusion 24 -1157 24 -1157 0 feedthrough
rlabel pdiffusion 31 -1157 31 -1157 0 cellNo=282
rlabel pdiffusion 38 -1157 38 -1157 0 feedthrough
rlabel pdiffusion 45 -1157 45 -1157 0 feedthrough
rlabel pdiffusion 52 -1157 52 -1157 0 feedthrough
rlabel pdiffusion 59 -1157 59 -1157 0 feedthrough
rlabel pdiffusion 66 -1157 66 -1157 0 feedthrough
rlabel pdiffusion 73 -1157 73 -1157 0 feedthrough
rlabel pdiffusion 80 -1157 80 -1157 0 cellNo=84
rlabel pdiffusion 87 -1157 87 -1157 0 feedthrough
rlabel pdiffusion 94 -1157 94 -1157 0 feedthrough
rlabel pdiffusion 101 -1157 101 -1157 0 feedthrough
rlabel pdiffusion 108 -1157 108 -1157 0 feedthrough
rlabel pdiffusion 115 -1157 115 -1157 0 feedthrough
rlabel pdiffusion 122 -1157 122 -1157 0 feedthrough
rlabel pdiffusion 129 -1157 129 -1157 0 cellNo=984
rlabel pdiffusion 136 -1157 136 -1157 0 feedthrough
rlabel pdiffusion 143 -1157 143 -1157 0 cellNo=81
rlabel pdiffusion 150 -1157 150 -1157 0 feedthrough
rlabel pdiffusion 157 -1157 157 -1157 0 feedthrough
rlabel pdiffusion 164 -1157 164 -1157 0 feedthrough
rlabel pdiffusion 171 -1157 171 -1157 0 feedthrough
rlabel pdiffusion 178 -1157 178 -1157 0 feedthrough
rlabel pdiffusion 185 -1157 185 -1157 0 cellNo=112
rlabel pdiffusion 192 -1157 192 -1157 0 feedthrough
rlabel pdiffusion 199 -1157 199 -1157 0 feedthrough
rlabel pdiffusion 206 -1157 206 -1157 0 feedthrough
rlabel pdiffusion 213 -1157 213 -1157 0 feedthrough
rlabel pdiffusion 220 -1157 220 -1157 0 feedthrough
rlabel pdiffusion 227 -1157 227 -1157 0 cellNo=253
rlabel pdiffusion 234 -1157 234 -1157 0 cellNo=440
rlabel pdiffusion 241 -1157 241 -1157 0 cellNo=661
rlabel pdiffusion 248 -1157 248 -1157 0 feedthrough
rlabel pdiffusion 255 -1157 255 -1157 0 feedthrough
rlabel pdiffusion 262 -1157 262 -1157 0 cellNo=505
rlabel pdiffusion 269 -1157 269 -1157 0 feedthrough
rlabel pdiffusion 276 -1157 276 -1157 0 feedthrough
rlabel pdiffusion 283 -1157 283 -1157 0 feedthrough
rlabel pdiffusion 290 -1157 290 -1157 0 feedthrough
rlabel pdiffusion 297 -1157 297 -1157 0 feedthrough
rlabel pdiffusion 304 -1157 304 -1157 0 cellNo=751
rlabel pdiffusion 311 -1157 311 -1157 0 feedthrough
rlabel pdiffusion 318 -1157 318 -1157 0 feedthrough
rlabel pdiffusion 325 -1157 325 -1157 0 feedthrough
rlabel pdiffusion 332 -1157 332 -1157 0 cellNo=231
rlabel pdiffusion 339 -1157 339 -1157 0 feedthrough
rlabel pdiffusion 346 -1157 346 -1157 0 feedthrough
rlabel pdiffusion 353 -1157 353 -1157 0 cellNo=509
rlabel pdiffusion 360 -1157 360 -1157 0 feedthrough
rlabel pdiffusion 367 -1157 367 -1157 0 cellNo=637
rlabel pdiffusion 374 -1157 374 -1157 0 feedthrough
rlabel pdiffusion 381 -1157 381 -1157 0 feedthrough
rlabel pdiffusion 388 -1157 388 -1157 0 feedthrough
rlabel pdiffusion 395 -1157 395 -1157 0 feedthrough
rlabel pdiffusion 402 -1157 402 -1157 0 feedthrough
rlabel pdiffusion 409 -1157 409 -1157 0 feedthrough
rlabel pdiffusion 416 -1157 416 -1157 0 feedthrough
rlabel pdiffusion 423 -1157 423 -1157 0 feedthrough
rlabel pdiffusion 430 -1157 430 -1157 0 feedthrough
rlabel pdiffusion 437 -1157 437 -1157 0 cellNo=721
rlabel pdiffusion 444 -1157 444 -1157 0 cellNo=813
rlabel pdiffusion 451 -1157 451 -1157 0 feedthrough
rlabel pdiffusion 458 -1157 458 -1157 0 feedthrough
rlabel pdiffusion 465 -1157 465 -1157 0 cellNo=834
rlabel pdiffusion 472 -1157 472 -1157 0 cellNo=923
rlabel pdiffusion 479 -1157 479 -1157 0 feedthrough
rlabel pdiffusion 486 -1157 486 -1157 0 feedthrough
rlabel pdiffusion 493 -1157 493 -1157 0 cellNo=925
rlabel pdiffusion 500 -1157 500 -1157 0 feedthrough
rlabel pdiffusion 507 -1157 507 -1157 0 cellNo=861
rlabel pdiffusion 514 -1157 514 -1157 0 feedthrough
rlabel pdiffusion 521 -1157 521 -1157 0 feedthrough
rlabel pdiffusion 528 -1157 528 -1157 0 cellNo=986
rlabel pdiffusion 535 -1157 535 -1157 0 feedthrough
rlabel pdiffusion 542 -1157 542 -1157 0 feedthrough
rlabel pdiffusion 549 -1157 549 -1157 0 feedthrough
rlabel pdiffusion 556 -1157 556 -1157 0 feedthrough
rlabel pdiffusion 563 -1157 563 -1157 0 feedthrough
rlabel pdiffusion 570 -1157 570 -1157 0 feedthrough
rlabel pdiffusion 577 -1157 577 -1157 0 feedthrough
rlabel pdiffusion 584 -1157 584 -1157 0 cellNo=668
rlabel pdiffusion 591 -1157 591 -1157 0 cellNo=858
rlabel pdiffusion 598 -1157 598 -1157 0 cellNo=274
rlabel pdiffusion 605 -1157 605 -1157 0 cellNo=257
rlabel pdiffusion 612 -1157 612 -1157 0 feedthrough
rlabel pdiffusion 619 -1157 619 -1157 0 cellNo=877
rlabel pdiffusion 626 -1157 626 -1157 0 cellNo=581
rlabel pdiffusion 633 -1157 633 -1157 0 feedthrough
rlabel pdiffusion 640 -1157 640 -1157 0 cellNo=241
rlabel pdiffusion 647 -1157 647 -1157 0 feedthrough
rlabel pdiffusion 654 -1157 654 -1157 0 feedthrough
rlabel pdiffusion 661 -1157 661 -1157 0 cellNo=144
rlabel pdiffusion 668 -1157 668 -1157 0 feedthrough
rlabel pdiffusion 675 -1157 675 -1157 0 cellNo=215
rlabel pdiffusion 682 -1157 682 -1157 0 feedthrough
rlabel pdiffusion 689 -1157 689 -1157 0 cellNo=818
rlabel pdiffusion 696 -1157 696 -1157 0 feedthrough
rlabel pdiffusion 703 -1157 703 -1157 0 feedthrough
rlabel pdiffusion 710 -1157 710 -1157 0 feedthrough
rlabel pdiffusion 717 -1157 717 -1157 0 feedthrough
rlabel pdiffusion 724 -1157 724 -1157 0 cellNo=730
rlabel pdiffusion 731 -1157 731 -1157 0 cellNo=93
rlabel pdiffusion 738 -1157 738 -1157 0 feedthrough
rlabel pdiffusion 745 -1157 745 -1157 0 feedthrough
rlabel pdiffusion 752 -1157 752 -1157 0 feedthrough
rlabel pdiffusion 759 -1157 759 -1157 0 feedthrough
rlabel pdiffusion 766 -1157 766 -1157 0 feedthrough
rlabel pdiffusion 773 -1157 773 -1157 0 feedthrough
rlabel pdiffusion 780 -1157 780 -1157 0 feedthrough
rlabel pdiffusion 787 -1157 787 -1157 0 feedthrough
rlabel pdiffusion 794 -1157 794 -1157 0 feedthrough
rlabel pdiffusion 801 -1157 801 -1157 0 feedthrough
rlabel pdiffusion 808 -1157 808 -1157 0 feedthrough
rlabel pdiffusion 815 -1157 815 -1157 0 feedthrough
rlabel pdiffusion 822 -1157 822 -1157 0 feedthrough
rlabel pdiffusion 829 -1157 829 -1157 0 feedthrough
rlabel pdiffusion 836 -1157 836 -1157 0 feedthrough
rlabel pdiffusion 843 -1157 843 -1157 0 feedthrough
rlabel pdiffusion 850 -1157 850 -1157 0 feedthrough
rlabel pdiffusion 857 -1157 857 -1157 0 feedthrough
rlabel pdiffusion 864 -1157 864 -1157 0 feedthrough
rlabel pdiffusion 871 -1157 871 -1157 0 feedthrough
rlabel pdiffusion 878 -1157 878 -1157 0 feedthrough
rlabel pdiffusion 885 -1157 885 -1157 0 feedthrough
rlabel pdiffusion 892 -1157 892 -1157 0 feedthrough
rlabel pdiffusion 899 -1157 899 -1157 0 feedthrough
rlabel pdiffusion 906 -1157 906 -1157 0 feedthrough
rlabel pdiffusion 913 -1157 913 -1157 0 feedthrough
rlabel pdiffusion 920 -1157 920 -1157 0 feedthrough
rlabel pdiffusion 927 -1157 927 -1157 0 feedthrough
rlabel pdiffusion 934 -1157 934 -1157 0 feedthrough
rlabel pdiffusion 941 -1157 941 -1157 0 feedthrough
rlabel pdiffusion 948 -1157 948 -1157 0 feedthrough
rlabel pdiffusion 955 -1157 955 -1157 0 feedthrough
rlabel pdiffusion 962 -1157 962 -1157 0 feedthrough
rlabel pdiffusion 969 -1157 969 -1157 0 feedthrough
rlabel pdiffusion 976 -1157 976 -1157 0 feedthrough
rlabel pdiffusion 983 -1157 983 -1157 0 feedthrough
rlabel pdiffusion 990 -1157 990 -1157 0 feedthrough
rlabel pdiffusion 997 -1157 997 -1157 0 feedthrough
rlabel pdiffusion 1004 -1157 1004 -1157 0 feedthrough
rlabel pdiffusion 1011 -1157 1011 -1157 0 feedthrough
rlabel pdiffusion 1018 -1157 1018 -1157 0 feedthrough
rlabel pdiffusion 1025 -1157 1025 -1157 0 feedthrough
rlabel pdiffusion 1032 -1157 1032 -1157 0 feedthrough
rlabel pdiffusion 1039 -1157 1039 -1157 0 feedthrough
rlabel pdiffusion 1046 -1157 1046 -1157 0 feedthrough
rlabel pdiffusion 1053 -1157 1053 -1157 0 feedthrough
rlabel pdiffusion 1060 -1157 1060 -1157 0 feedthrough
rlabel pdiffusion 1067 -1157 1067 -1157 0 feedthrough
rlabel pdiffusion 1074 -1157 1074 -1157 0 feedthrough
rlabel pdiffusion 1081 -1157 1081 -1157 0 feedthrough
rlabel pdiffusion 1088 -1157 1088 -1157 0 cellNo=860
rlabel pdiffusion 1095 -1157 1095 -1157 0 feedthrough
rlabel pdiffusion 1102 -1157 1102 -1157 0 feedthrough
rlabel pdiffusion 3 -1260 3 -1260 0 feedthrough
rlabel pdiffusion 10 -1260 10 -1260 0 feedthrough
rlabel pdiffusion 17 -1260 17 -1260 0 cellNo=354
rlabel pdiffusion 24 -1260 24 -1260 0 cellNo=450
rlabel pdiffusion 31 -1260 31 -1260 0 feedthrough
rlabel pdiffusion 38 -1260 38 -1260 0 feedthrough
rlabel pdiffusion 45 -1260 45 -1260 0 feedthrough
rlabel pdiffusion 52 -1260 52 -1260 0 cellNo=220
rlabel pdiffusion 59 -1260 59 -1260 0 feedthrough
rlabel pdiffusion 66 -1260 66 -1260 0 feedthrough
rlabel pdiffusion 73 -1260 73 -1260 0 feedthrough
rlabel pdiffusion 80 -1260 80 -1260 0 cellNo=272
rlabel pdiffusion 87 -1260 87 -1260 0 feedthrough
rlabel pdiffusion 94 -1260 94 -1260 0 feedthrough
rlabel pdiffusion 101 -1260 101 -1260 0 feedthrough
rlabel pdiffusion 108 -1260 108 -1260 0 feedthrough
rlabel pdiffusion 115 -1260 115 -1260 0 cellNo=734
rlabel pdiffusion 122 -1260 122 -1260 0 feedthrough
rlabel pdiffusion 129 -1260 129 -1260 0 feedthrough
rlabel pdiffusion 136 -1260 136 -1260 0 feedthrough
rlabel pdiffusion 143 -1260 143 -1260 0 feedthrough
rlabel pdiffusion 150 -1260 150 -1260 0 feedthrough
rlabel pdiffusion 157 -1260 157 -1260 0 feedthrough
rlabel pdiffusion 164 -1260 164 -1260 0 cellNo=343
rlabel pdiffusion 171 -1260 171 -1260 0 cellNo=546
rlabel pdiffusion 178 -1260 178 -1260 0 feedthrough
rlabel pdiffusion 185 -1260 185 -1260 0 cellNo=2
rlabel pdiffusion 192 -1260 192 -1260 0 cellNo=717
rlabel pdiffusion 199 -1260 199 -1260 0 cellNo=255
rlabel pdiffusion 206 -1260 206 -1260 0 feedthrough
rlabel pdiffusion 213 -1260 213 -1260 0 cellNo=579
rlabel pdiffusion 220 -1260 220 -1260 0 cellNo=714
rlabel pdiffusion 227 -1260 227 -1260 0 feedthrough
rlabel pdiffusion 234 -1260 234 -1260 0 feedthrough
rlabel pdiffusion 241 -1260 241 -1260 0 feedthrough
rlabel pdiffusion 248 -1260 248 -1260 0 feedthrough
rlabel pdiffusion 255 -1260 255 -1260 0 feedthrough
rlabel pdiffusion 262 -1260 262 -1260 0 feedthrough
rlabel pdiffusion 269 -1260 269 -1260 0 feedthrough
rlabel pdiffusion 276 -1260 276 -1260 0 feedthrough
rlabel pdiffusion 283 -1260 283 -1260 0 feedthrough
rlabel pdiffusion 290 -1260 290 -1260 0 cellNo=123
rlabel pdiffusion 297 -1260 297 -1260 0 feedthrough
rlabel pdiffusion 304 -1260 304 -1260 0 feedthrough
rlabel pdiffusion 311 -1260 311 -1260 0 feedthrough
rlabel pdiffusion 318 -1260 318 -1260 0 feedthrough
rlabel pdiffusion 325 -1260 325 -1260 0 feedthrough
rlabel pdiffusion 332 -1260 332 -1260 0 feedthrough
rlabel pdiffusion 339 -1260 339 -1260 0 feedthrough
rlabel pdiffusion 346 -1260 346 -1260 0 feedthrough
rlabel pdiffusion 353 -1260 353 -1260 0 feedthrough
rlabel pdiffusion 360 -1260 360 -1260 0 feedthrough
rlabel pdiffusion 367 -1260 367 -1260 0 feedthrough
rlabel pdiffusion 374 -1260 374 -1260 0 feedthrough
rlabel pdiffusion 381 -1260 381 -1260 0 feedthrough
rlabel pdiffusion 388 -1260 388 -1260 0 feedthrough
rlabel pdiffusion 395 -1260 395 -1260 0 feedthrough
rlabel pdiffusion 402 -1260 402 -1260 0 feedthrough
rlabel pdiffusion 409 -1260 409 -1260 0 feedthrough
rlabel pdiffusion 416 -1260 416 -1260 0 feedthrough
rlabel pdiffusion 423 -1260 423 -1260 0 cellNo=12
rlabel pdiffusion 430 -1260 430 -1260 0 cellNo=280
rlabel pdiffusion 437 -1260 437 -1260 0 feedthrough
rlabel pdiffusion 444 -1260 444 -1260 0 feedthrough
rlabel pdiffusion 451 -1260 451 -1260 0 feedthrough
rlabel pdiffusion 458 -1260 458 -1260 0 cellNo=188
rlabel pdiffusion 465 -1260 465 -1260 0 feedthrough
rlabel pdiffusion 472 -1260 472 -1260 0 cellNo=462
rlabel pdiffusion 479 -1260 479 -1260 0 feedthrough
rlabel pdiffusion 486 -1260 486 -1260 0 feedthrough
rlabel pdiffusion 493 -1260 493 -1260 0 cellNo=641
rlabel pdiffusion 500 -1260 500 -1260 0 cellNo=401
rlabel pdiffusion 507 -1260 507 -1260 0 feedthrough
rlabel pdiffusion 514 -1260 514 -1260 0 cellNo=778
rlabel pdiffusion 521 -1260 521 -1260 0 cellNo=376
rlabel pdiffusion 528 -1260 528 -1260 0 feedthrough
rlabel pdiffusion 535 -1260 535 -1260 0 cellNo=247
rlabel pdiffusion 542 -1260 542 -1260 0 cellNo=645
rlabel pdiffusion 549 -1260 549 -1260 0 cellNo=789
rlabel pdiffusion 556 -1260 556 -1260 0 feedthrough
rlabel pdiffusion 563 -1260 563 -1260 0 cellNo=132
rlabel pdiffusion 570 -1260 570 -1260 0 feedthrough
rlabel pdiffusion 577 -1260 577 -1260 0 feedthrough
rlabel pdiffusion 584 -1260 584 -1260 0 cellNo=374
rlabel pdiffusion 591 -1260 591 -1260 0 cellNo=430
rlabel pdiffusion 598 -1260 598 -1260 0 feedthrough
rlabel pdiffusion 605 -1260 605 -1260 0 cellNo=194
rlabel pdiffusion 612 -1260 612 -1260 0 feedthrough
rlabel pdiffusion 619 -1260 619 -1260 0 feedthrough
rlabel pdiffusion 626 -1260 626 -1260 0 feedthrough
rlabel pdiffusion 633 -1260 633 -1260 0 feedthrough
rlabel pdiffusion 640 -1260 640 -1260 0 feedthrough
rlabel pdiffusion 647 -1260 647 -1260 0 feedthrough
rlabel pdiffusion 654 -1260 654 -1260 0 cellNo=501
rlabel pdiffusion 661 -1260 661 -1260 0 feedthrough
rlabel pdiffusion 668 -1260 668 -1260 0 feedthrough
rlabel pdiffusion 675 -1260 675 -1260 0 feedthrough
rlabel pdiffusion 682 -1260 682 -1260 0 cellNo=951
rlabel pdiffusion 689 -1260 689 -1260 0 feedthrough
rlabel pdiffusion 696 -1260 696 -1260 0 feedthrough
rlabel pdiffusion 703 -1260 703 -1260 0 feedthrough
rlabel pdiffusion 710 -1260 710 -1260 0 feedthrough
rlabel pdiffusion 717 -1260 717 -1260 0 cellNo=931
rlabel pdiffusion 724 -1260 724 -1260 0 feedthrough
rlabel pdiffusion 731 -1260 731 -1260 0 feedthrough
rlabel pdiffusion 738 -1260 738 -1260 0 feedthrough
rlabel pdiffusion 745 -1260 745 -1260 0 feedthrough
rlabel pdiffusion 752 -1260 752 -1260 0 feedthrough
rlabel pdiffusion 759 -1260 759 -1260 0 feedthrough
rlabel pdiffusion 766 -1260 766 -1260 0 feedthrough
rlabel pdiffusion 773 -1260 773 -1260 0 feedthrough
rlabel pdiffusion 780 -1260 780 -1260 0 cellNo=762
rlabel pdiffusion 787 -1260 787 -1260 0 feedthrough
rlabel pdiffusion 794 -1260 794 -1260 0 feedthrough
rlabel pdiffusion 801 -1260 801 -1260 0 feedthrough
rlabel pdiffusion 808 -1260 808 -1260 0 feedthrough
rlabel pdiffusion 815 -1260 815 -1260 0 cellNo=793
rlabel pdiffusion 822 -1260 822 -1260 0 feedthrough
rlabel pdiffusion 829 -1260 829 -1260 0 feedthrough
rlabel pdiffusion 836 -1260 836 -1260 0 feedthrough
rlabel pdiffusion 843 -1260 843 -1260 0 feedthrough
rlabel pdiffusion 850 -1260 850 -1260 0 feedthrough
rlabel pdiffusion 857 -1260 857 -1260 0 feedthrough
rlabel pdiffusion 864 -1260 864 -1260 0 feedthrough
rlabel pdiffusion 871 -1260 871 -1260 0 feedthrough
rlabel pdiffusion 878 -1260 878 -1260 0 feedthrough
rlabel pdiffusion 885 -1260 885 -1260 0 feedthrough
rlabel pdiffusion 892 -1260 892 -1260 0 feedthrough
rlabel pdiffusion 899 -1260 899 -1260 0 feedthrough
rlabel pdiffusion 906 -1260 906 -1260 0 feedthrough
rlabel pdiffusion 913 -1260 913 -1260 0 feedthrough
rlabel pdiffusion 920 -1260 920 -1260 0 feedthrough
rlabel pdiffusion 927 -1260 927 -1260 0 feedthrough
rlabel pdiffusion 934 -1260 934 -1260 0 feedthrough
rlabel pdiffusion 941 -1260 941 -1260 0 feedthrough
rlabel pdiffusion 948 -1260 948 -1260 0 feedthrough
rlabel pdiffusion 955 -1260 955 -1260 0 feedthrough
rlabel pdiffusion 962 -1260 962 -1260 0 feedthrough
rlabel pdiffusion 969 -1260 969 -1260 0 feedthrough
rlabel pdiffusion 976 -1260 976 -1260 0 feedthrough
rlabel pdiffusion 983 -1260 983 -1260 0 feedthrough
rlabel pdiffusion 990 -1260 990 -1260 0 feedthrough
rlabel pdiffusion 997 -1260 997 -1260 0 feedthrough
rlabel pdiffusion 1004 -1260 1004 -1260 0 feedthrough
rlabel pdiffusion 1011 -1260 1011 -1260 0 feedthrough
rlabel pdiffusion 1018 -1260 1018 -1260 0 feedthrough
rlabel pdiffusion 1025 -1260 1025 -1260 0 feedthrough
rlabel pdiffusion 1032 -1260 1032 -1260 0 cellNo=788
rlabel pdiffusion 1039 -1260 1039 -1260 0 cellNo=572
rlabel pdiffusion 1046 -1260 1046 -1260 0 feedthrough
rlabel pdiffusion 1053 -1260 1053 -1260 0 feedthrough
rlabel pdiffusion 1060 -1260 1060 -1260 0 feedthrough
rlabel pdiffusion 1067 -1260 1067 -1260 0 feedthrough
rlabel pdiffusion 1074 -1260 1074 -1260 0 feedthrough
rlabel pdiffusion 10 -1339 10 -1339 0 feedthrough
rlabel pdiffusion 17 -1339 17 -1339 0 feedthrough
rlabel pdiffusion 24 -1339 24 -1339 0 feedthrough
rlabel pdiffusion 31 -1339 31 -1339 0 feedthrough
rlabel pdiffusion 38 -1339 38 -1339 0 feedthrough
rlabel pdiffusion 45 -1339 45 -1339 0 feedthrough
rlabel pdiffusion 52 -1339 52 -1339 0 feedthrough
rlabel pdiffusion 59 -1339 59 -1339 0 feedthrough
rlabel pdiffusion 66 -1339 66 -1339 0 feedthrough
rlabel pdiffusion 73 -1339 73 -1339 0 feedthrough
rlabel pdiffusion 80 -1339 80 -1339 0 cellNo=287
rlabel pdiffusion 87 -1339 87 -1339 0 cellNo=7
rlabel pdiffusion 94 -1339 94 -1339 0 feedthrough
rlabel pdiffusion 101 -1339 101 -1339 0 feedthrough
rlabel pdiffusion 108 -1339 108 -1339 0 feedthrough
rlabel pdiffusion 115 -1339 115 -1339 0 cellNo=612
rlabel pdiffusion 122 -1339 122 -1339 0 feedthrough
rlabel pdiffusion 129 -1339 129 -1339 0 cellNo=27
rlabel pdiffusion 136 -1339 136 -1339 0 cellNo=599
rlabel pdiffusion 143 -1339 143 -1339 0 feedthrough
rlabel pdiffusion 150 -1339 150 -1339 0 feedthrough
rlabel pdiffusion 157 -1339 157 -1339 0 cellNo=616
rlabel pdiffusion 164 -1339 164 -1339 0 feedthrough
rlabel pdiffusion 171 -1339 171 -1339 0 cellNo=341
rlabel pdiffusion 178 -1339 178 -1339 0 cellNo=545
rlabel pdiffusion 185 -1339 185 -1339 0 feedthrough
rlabel pdiffusion 192 -1339 192 -1339 0 cellNo=565
rlabel pdiffusion 199 -1339 199 -1339 0 feedthrough
rlabel pdiffusion 206 -1339 206 -1339 0 feedthrough
rlabel pdiffusion 213 -1339 213 -1339 0 feedthrough
rlabel pdiffusion 220 -1339 220 -1339 0 cellNo=882
rlabel pdiffusion 227 -1339 227 -1339 0 feedthrough
rlabel pdiffusion 234 -1339 234 -1339 0 feedthrough
rlabel pdiffusion 241 -1339 241 -1339 0 feedthrough
rlabel pdiffusion 248 -1339 248 -1339 0 feedthrough
rlabel pdiffusion 255 -1339 255 -1339 0 feedthrough
rlabel pdiffusion 262 -1339 262 -1339 0 feedthrough
rlabel pdiffusion 269 -1339 269 -1339 0 feedthrough
rlabel pdiffusion 276 -1339 276 -1339 0 feedthrough
rlabel pdiffusion 283 -1339 283 -1339 0 feedthrough
rlabel pdiffusion 290 -1339 290 -1339 0 cellNo=999
rlabel pdiffusion 297 -1339 297 -1339 0 feedthrough
rlabel pdiffusion 304 -1339 304 -1339 0 feedthrough
rlabel pdiffusion 311 -1339 311 -1339 0 feedthrough
rlabel pdiffusion 318 -1339 318 -1339 0 cellNo=722
rlabel pdiffusion 325 -1339 325 -1339 0 cellNo=987
rlabel pdiffusion 332 -1339 332 -1339 0 feedthrough
rlabel pdiffusion 339 -1339 339 -1339 0 feedthrough
rlabel pdiffusion 346 -1339 346 -1339 0 feedthrough
rlabel pdiffusion 353 -1339 353 -1339 0 cellNo=707
rlabel pdiffusion 360 -1339 360 -1339 0 feedthrough
rlabel pdiffusion 367 -1339 367 -1339 0 cellNo=250
rlabel pdiffusion 374 -1339 374 -1339 0 feedthrough
rlabel pdiffusion 381 -1339 381 -1339 0 feedthrough
rlabel pdiffusion 388 -1339 388 -1339 0 feedthrough
rlabel pdiffusion 395 -1339 395 -1339 0 feedthrough
rlabel pdiffusion 402 -1339 402 -1339 0 feedthrough
rlabel pdiffusion 409 -1339 409 -1339 0 feedthrough
rlabel pdiffusion 416 -1339 416 -1339 0 feedthrough
rlabel pdiffusion 423 -1339 423 -1339 0 feedthrough
rlabel pdiffusion 430 -1339 430 -1339 0 cellNo=486
rlabel pdiffusion 437 -1339 437 -1339 0 feedthrough
rlabel pdiffusion 444 -1339 444 -1339 0 feedthrough
rlabel pdiffusion 451 -1339 451 -1339 0 feedthrough
rlabel pdiffusion 458 -1339 458 -1339 0 cellNo=14
rlabel pdiffusion 465 -1339 465 -1339 0 feedthrough
rlabel pdiffusion 472 -1339 472 -1339 0 cellNo=654
rlabel pdiffusion 479 -1339 479 -1339 0 feedthrough
rlabel pdiffusion 486 -1339 486 -1339 0 feedthrough
rlabel pdiffusion 493 -1339 493 -1339 0 cellNo=729
rlabel pdiffusion 500 -1339 500 -1339 0 feedthrough
rlabel pdiffusion 507 -1339 507 -1339 0 cellNo=13
rlabel pdiffusion 514 -1339 514 -1339 0 feedthrough
rlabel pdiffusion 521 -1339 521 -1339 0 feedthrough
rlabel pdiffusion 528 -1339 528 -1339 0 feedthrough
rlabel pdiffusion 535 -1339 535 -1339 0 cellNo=327
rlabel pdiffusion 542 -1339 542 -1339 0 feedthrough
rlabel pdiffusion 549 -1339 549 -1339 0 feedthrough
rlabel pdiffusion 556 -1339 556 -1339 0 feedthrough
rlabel pdiffusion 563 -1339 563 -1339 0 feedthrough
rlabel pdiffusion 570 -1339 570 -1339 0 feedthrough
rlabel pdiffusion 577 -1339 577 -1339 0 cellNo=826
rlabel pdiffusion 584 -1339 584 -1339 0 cellNo=108
rlabel pdiffusion 591 -1339 591 -1339 0 feedthrough
rlabel pdiffusion 598 -1339 598 -1339 0 cellNo=275
rlabel pdiffusion 605 -1339 605 -1339 0 feedthrough
rlabel pdiffusion 612 -1339 612 -1339 0 feedthrough
rlabel pdiffusion 619 -1339 619 -1339 0 cellNo=735
rlabel pdiffusion 626 -1339 626 -1339 0 feedthrough
rlabel pdiffusion 633 -1339 633 -1339 0 feedthrough
rlabel pdiffusion 640 -1339 640 -1339 0 feedthrough
rlabel pdiffusion 647 -1339 647 -1339 0 cellNo=427
rlabel pdiffusion 654 -1339 654 -1339 0 feedthrough
rlabel pdiffusion 661 -1339 661 -1339 0 feedthrough
rlabel pdiffusion 668 -1339 668 -1339 0 feedthrough
rlabel pdiffusion 675 -1339 675 -1339 0 cellNo=23
rlabel pdiffusion 682 -1339 682 -1339 0 feedthrough
rlabel pdiffusion 689 -1339 689 -1339 0 feedthrough
rlabel pdiffusion 696 -1339 696 -1339 0 feedthrough
rlabel pdiffusion 703 -1339 703 -1339 0 cellNo=310
rlabel pdiffusion 710 -1339 710 -1339 0 feedthrough
rlabel pdiffusion 717 -1339 717 -1339 0 feedthrough
rlabel pdiffusion 724 -1339 724 -1339 0 feedthrough
rlabel pdiffusion 731 -1339 731 -1339 0 feedthrough
rlabel pdiffusion 738 -1339 738 -1339 0 cellNo=631
rlabel pdiffusion 745 -1339 745 -1339 0 feedthrough
rlabel pdiffusion 752 -1339 752 -1339 0 feedthrough
rlabel pdiffusion 759 -1339 759 -1339 0 cellNo=43
rlabel pdiffusion 766 -1339 766 -1339 0 feedthrough
rlabel pdiffusion 773 -1339 773 -1339 0 feedthrough
rlabel pdiffusion 780 -1339 780 -1339 0 feedthrough
rlabel pdiffusion 787 -1339 787 -1339 0 feedthrough
rlabel pdiffusion 794 -1339 794 -1339 0 feedthrough
rlabel pdiffusion 801 -1339 801 -1339 0 feedthrough
rlabel pdiffusion 808 -1339 808 -1339 0 feedthrough
rlabel pdiffusion 815 -1339 815 -1339 0 feedthrough
rlabel pdiffusion 822 -1339 822 -1339 0 feedthrough
rlabel pdiffusion 829 -1339 829 -1339 0 feedthrough
rlabel pdiffusion 836 -1339 836 -1339 0 feedthrough
rlabel pdiffusion 843 -1339 843 -1339 0 feedthrough
rlabel pdiffusion 850 -1339 850 -1339 0 feedthrough
rlabel pdiffusion 857 -1339 857 -1339 0 feedthrough
rlabel pdiffusion 864 -1339 864 -1339 0 feedthrough
rlabel pdiffusion 871 -1339 871 -1339 0 feedthrough
rlabel pdiffusion 878 -1339 878 -1339 0 feedthrough
rlabel pdiffusion 885 -1339 885 -1339 0 feedthrough
rlabel pdiffusion 892 -1339 892 -1339 0 feedthrough
rlabel pdiffusion 899 -1339 899 -1339 0 feedthrough
rlabel pdiffusion 906 -1339 906 -1339 0 feedthrough
rlabel pdiffusion 913 -1339 913 -1339 0 feedthrough
rlabel pdiffusion 920 -1339 920 -1339 0 feedthrough
rlabel pdiffusion 927 -1339 927 -1339 0 feedthrough
rlabel pdiffusion 934 -1339 934 -1339 0 feedthrough
rlabel pdiffusion 941 -1339 941 -1339 0 feedthrough
rlabel pdiffusion 948 -1339 948 -1339 0 feedthrough
rlabel pdiffusion 955 -1339 955 -1339 0 feedthrough
rlabel pdiffusion 962 -1339 962 -1339 0 feedthrough
rlabel pdiffusion 969 -1339 969 -1339 0 feedthrough
rlabel pdiffusion 976 -1339 976 -1339 0 feedthrough
rlabel pdiffusion 983 -1339 983 -1339 0 feedthrough
rlabel pdiffusion 990 -1339 990 -1339 0 feedthrough
rlabel pdiffusion 997 -1339 997 -1339 0 feedthrough
rlabel pdiffusion 1004 -1339 1004 -1339 0 feedthrough
rlabel pdiffusion 1011 -1339 1011 -1339 0 feedthrough
rlabel pdiffusion 1018 -1339 1018 -1339 0 feedthrough
rlabel pdiffusion 1025 -1339 1025 -1339 0 cellNo=86
rlabel pdiffusion 1032 -1339 1032 -1339 0 cellNo=673
rlabel pdiffusion 1039 -1339 1039 -1339 0 cellNo=363
rlabel pdiffusion 1046 -1339 1046 -1339 0 cellNo=474
rlabel pdiffusion 1053 -1339 1053 -1339 0 feedthrough
rlabel pdiffusion 1060 -1339 1060 -1339 0 cellNo=576
rlabel pdiffusion 1067 -1339 1067 -1339 0 feedthrough
rlabel pdiffusion 1074 -1339 1074 -1339 0 feedthrough
rlabel pdiffusion 1081 -1339 1081 -1339 0 feedthrough
rlabel pdiffusion 17 -1416 17 -1416 0 feedthrough
rlabel pdiffusion 24 -1416 24 -1416 0 feedthrough
rlabel pdiffusion 31 -1416 31 -1416 0 feedthrough
rlabel pdiffusion 38 -1416 38 -1416 0 feedthrough
rlabel pdiffusion 45 -1416 45 -1416 0 feedthrough
rlabel pdiffusion 52 -1416 52 -1416 0 cellNo=80
rlabel pdiffusion 59 -1416 59 -1416 0 cellNo=856
rlabel pdiffusion 66 -1416 66 -1416 0 feedthrough
rlabel pdiffusion 73 -1416 73 -1416 0 feedthrough
rlabel pdiffusion 80 -1416 80 -1416 0 feedthrough
rlabel pdiffusion 87 -1416 87 -1416 0 cellNo=399
rlabel pdiffusion 94 -1416 94 -1416 0 feedthrough
rlabel pdiffusion 101 -1416 101 -1416 0 feedthrough
rlabel pdiffusion 108 -1416 108 -1416 0 feedthrough
rlabel pdiffusion 115 -1416 115 -1416 0 feedthrough
rlabel pdiffusion 122 -1416 122 -1416 0 feedthrough
rlabel pdiffusion 129 -1416 129 -1416 0 feedthrough
rlabel pdiffusion 136 -1416 136 -1416 0 cellNo=411
rlabel pdiffusion 143 -1416 143 -1416 0 cellNo=924
rlabel pdiffusion 150 -1416 150 -1416 0 feedthrough
rlabel pdiffusion 157 -1416 157 -1416 0 cellNo=382
rlabel pdiffusion 164 -1416 164 -1416 0 cellNo=948
rlabel pdiffusion 171 -1416 171 -1416 0 feedthrough
rlabel pdiffusion 178 -1416 178 -1416 0 feedthrough
rlabel pdiffusion 185 -1416 185 -1416 0 feedthrough
rlabel pdiffusion 192 -1416 192 -1416 0 feedthrough
rlabel pdiffusion 199 -1416 199 -1416 0 feedthrough
rlabel pdiffusion 206 -1416 206 -1416 0 cellNo=289
rlabel pdiffusion 213 -1416 213 -1416 0 feedthrough
rlabel pdiffusion 220 -1416 220 -1416 0 cellNo=643
rlabel pdiffusion 227 -1416 227 -1416 0 feedthrough
rlabel pdiffusion 234 -1416 234 -1416 0 feedthrough
rlabel pdiffusion 241 -1416 241 -1416 0 cellNo=894
rlabel pdiffusion 248 -1416 248 -1416 0 feedthrough
rlabel pdiffusion 255 -1416 255 -1416 0 feedthrough
rlabel pdiffusion 262 -1416 262 -1416 0 feedthrough
rlabel pdiffusion 269 -1416 269 -1416 0 feedthrough
rlabel pdiffusion 276 -1416 276 -1416 0 feedthrough
rlabel pdiffusion 283 -1416 283 -1416 0 feedthrough
rlabel pdiffusion 290 -1416 290 -1416 0 feedthrough
rlabel pdiffusion 297 -1416 297 -1416 0 feedthrough
rlabel pdiffusion 304 -1416 304 -1416 0 cellNo=396
rlabel pdiffusion 311 -1416 311 -1416 0 feedthrough
rlabel pdiffusion 318 -1416 318 -1416 0 feedthrough
rlabel pdiffusion 325 -1416 325 -1416 0 feedthrough
rlabel pdiffusion 332 -1416 332 -1416 0 feedthrough
rlabel pdiffusion 339 -1416 339 -1416 0 feedthrough
rlabel pdiffusion 346 -1416 346 -1416 0 feedthrough
rlabel pdiffusion 353 -1416 353 -1416 0 cellNo=246
rlabel pdiffusion 360 -1416 360 -1416 0 cellNo=66
rlabel pdiffusion 367 -1416 367 -1416 0 feedthrough
rlabel pdiffusion 374 -1416 374 -1416 0 feedthrough
rlabel pdiffusion 381 -1416 381 -1416 0 feedthrough
rlabel pdiffusion 388 -1416 388 -1416 0 cellNo=165
rlabel pdiffusion 395 -1416 395 -1416 0 feedthrough
rlabel pdiffusion 402 -1416 402 -1416 0 cellNo=226
rlabel pdiffusion 409 -1416 409 -1416 0 cellNo=491
rlabel pdiffusion 416 -1416 416 -1416 0 feedthrough
rlabel pdiffusion 423 -1416 423 -1416 0 feedthrough
rlabel pdiffusion 430 -1416 430 -1416 0 feedthrough
rlabel pdiffusion 437 -1416 437 -1416 0 feedthrough
rlabel pdiffusion 444 -1416 444 -1416 0 feedthrough
rlabel pdiffusion 451 -1416 451 -1416 0 feedthrough
rlabel pdiffusion 458 -1416 458 -1416 0 feedthrough
rlabel pdiffusion 465 -1416 465 -1416 0 feedthrough
rlabel pdiffusion 472 -1416 472 -1416 0 feedthrough
rlabel pdiffusion 479 -1416 479 -1416 0 feedthrough
rlabel pdiffusion 486 -1416 486 -1416 0 feedthrough
rlabel pdiffusion 493 -1416 493 -1416 0 feedthrough
rlabel pdiffusion 500 -1416 500 -1416 0 feedthrough
rlabel pdiffusion 507 -1416 507 -1416 0 cellNo=155
rlabel pdiffusion 514 -1416 514 -1416 0 cellNo=204
rlabel pdiffusion 521 -1416 521 -1416 0 cellNo=161
rlabel pdiffusion 528 -1416 528 -1416 0 feedthrough
rlabel pdiffusion 535 -1416 535 -1416 0 feedthrough
rlabel pdiffusion 542 -1416 542 -1416 0 feedthrough
rlabel pdiffusion 549 -1416 549 -1416 0 feedthrough
rlabel pdiffusion 556 -1416 556 -1416 0 feedthrough
rlabel pdiffusion 563 -1416 563 -1416 0 cellNo=503
rlabel pdiffusion 570 -1416 570 -1416 0 cellNo=415
rlabel pdiffusion 577 -1416 577 -1416 0 cellNo=214
rlabel pdiffusion 584 -1416 584 -1416 0 cellNo=621
rlabel pdiffusion 591 -1416 591 -1416 0 feedthrough
rlabel pdiffusion 598 -1416 598 -1416 0 feedthrough
rlabel pdiffusion 605 -1416 605 -1416 0 feedthrough
rlabel pdiffusion 612 -1416 612 -1416 0 feedthrough
rlabel pdiffusion 619 -1416 619 -1416 0 feedthrough
rlabel pdiffusion 626 -1416 626 -1416 0 feedthrough
rlabel pdiffusion 633 -1416 633 -1416 0 feedthrough
rlabel pdiffusion 640 -1416 640 -1416 0 feedthrough
rlabel pdiffusion 647 -1416 647 -1416 0 feedthrough
rlabel pdiffusion 654 -1416 654 -1416 0 feedthrough
rlabel pdiffusion 661 -1416 661 -1416 0 cellNo=991
rlabel pdiffusion 668 -1416 668 -1416 0 feedthrough
rlabel pdiffusion 675 -1416 675 -1416 0 feedthrough
rlabel pdiffusion 682 -1416 682 -1416 0 cellNo=28
rlabel pdiffusion 689 -1416 689 -1416 0 feedthrough
rlabel pdiffusion 696 -1416 696 -1416 0 feedthrough
rlabel pdiffusion 703 -1416 703 -1416 0 cellNo=320
rlabel pdiffusion 710 -1416 710 -1416 0 cellNo=386
rlabel pdiffusion 717 -1416 717 -1416 0 feedthrough
rlabel pdiffusion 724 -1416 724 -1416 0 feedthrough
rlabel pdiffusion 731 -1416 731 -1416 0 feedthrough
rlabel pdiffusion 738 -1416 738 -1416 0 cellNo=956
rlabel pdiffusion 745 -1416 745 -1416 0 feedthrough
rlabel pdiffusion 752 -1416 752 -1416 0 feedthrough
rlabel pdiffusion 759 -1416 759 -1416 0 feedthrough
rlabel pdiffusion 766 -1416 766 -1416 0 cellNo=620
rlabel pdiffusion 773 -1416 773 -1416 0 feedthrough
rlabel pdiffusion 780 -1416 780 -1416 0 feedthrough
rlabel pdiffusion 787 -1416 787 -1416 0 feedthrough
rlabel pdiffusion 794 -1416 794 -1416 0 feedthrough
rlabel pdiffusion 801 -1416 801 -1416 0 feedthrough
rlabel pdiffusion 808 -1416 808 -1416 0 feedthrough
rlabel pdiffusion 815 -1416 815 -1416 0 feedthrough
rlabel pdiffusion 822 -1416 822 -1416 0 feedthrough
rlabel pdiffusion 829 -1416 829 -1416 0 feedthrough
rlabel pdiffusion 836 -1416 836 -1416 0 feedthrough
rlabel pdiffusion 843 -1416 843 -1416 0 feedthrough
rlabel pdiffusion 850 -1416 850 -1416 0 feedthrough
rlabel pdiffusion 857 -1416 857 -1416 0 feedthrough
rlabel pdiffusion 864 -1416 864 -1416 0 feedthrough
rlabel pdiffusion 871 -1416 871 -1416 0 feedthrough
rlabel pdiffusion 878 -1416 878 -1416 0 feedthrough
rlabel pdiffusion 885 -1416 885 -1416 0 feedthrough
rlabel pdiffusion 892 -1416 892 -1416 0 feedthrough
rlabel pdiffusion 899 -1416 899 -1416 0 feedthrough
rlabel pdiffusion 906 -1416 906 -1416 0 feedthrough
rlabel pdiffusion 913 -1416 913 -1416 0 feedthrough
rlabel pdiffusion 920 -1416 920 -1416 0 feedthrough
rlabel pdiffusion 927 -1416 927 -1416 0 cellNo=91
rlabel pdiffusion 934 -1416 934 -1416 0 feedthrough
rlabel pdiffusion 941 -1416 941 -1416 0 feedthrough
rlabel pdiffusion 948 -1416 948 -1416 0 cellNo=371
rlabel pdiffusion 955 -1416 955 -1416 0 feedthrough
rlabel pdiffusion 962 -1416 962 -1416 0 feedthrough
rlabel pdiffusion 969 -1416 969 -1416 0 cellNo=592
rlabel pdiffusion 976 -1416 976 -1416 0 feedthrough
rlabel pdiffusion 983 -1416 983 -1416 0 feedthrough
rlabel pdiffusion 990 -1416 990 -1416 0 feedthrough
rlabel pdiffusion 997 -1416 997 -1416 0 feedthrough
rlabel pdiffusion 1004 -1416 1004 -1416 0 cellNo=878
rlabel pdiffusion 1011 -1416 1011 -1416 0 feedthrough
rlabel pdiffusion 1018 -1416 1018 -1416 0 feedthrough
rlabel pdiffusion 1025 -1416 1025 -1416 0 feedthrough
rlabel pdiffusion 1032 -1416 1032 -1416 0 feedthrough
rlabel pdiffusion 1039 -1416 1039 -1416 0 cellNo=449
rlabel pdiffusion 1046 -1416 1046 -1416 0 feedthrough
rlabel pdiffusion 1053 -1416 1053 -1416 0 feedthrough
rlabel pdiffusion 1074 -1416 1074 -1416 0 feedthrough
rlabel pdiffusion 24 -1497 24 -1497 0 cellNo=606
rlabel pdiffusion 31 -1497 31 -1497 0 feedthrough
rlabel pdiffusion 38 -1497 38 -1497 0 feedthrough
rlabel pdiffusion 45 -1497 45 -1497 0 feedthrough
rlabel pdiffusion 52 -1497 52 -1497 0 cellNo=431
rlabel pdiffusion 59 -1497 59 -1497 0 feedthrough
rlabel pdiffusion 66 -1497 66 -1497 0 feedthrough
rlabel pdiffusion 73 -1497 73 -1497 0 cellNo=765
rlabel pdiffusion 80 -1497 80 -1497 0 feedthrough
rlabel pdiffusion 87 -1497 87 -1497 0 cellNo=356
rlabel pdiffusion 94 -1497 94 -1497 0 feedthrough
rlabel pdiffusion 101 -1497 101 -1497 0 feedthrough
rlabel pdiffusion 108 -1497 108 -1497 0 feedthrough
rlabel pdiffusion 115 -1497 115 -1497 0 feedthrough
rlabel pdiffusion 122 -1497 122 -1497 0 cellNo=355
rlabel pdiffusion 129 -1497 129 -1497 0 cellNo=508
rlabel pdiffusion 136 -1497 136 -1497 0 feedthrough
rlabel pdiffusion 143 -1497 143 -1497 0 feedthrough
rlabel pdiffusion 150 -1497 150 -1497 0 feedthrough
rlabel pdiffusion 157 -1497 157 -1497 0 feedthrough
rlabel pdiffusion 164 -1497 164 -1497 0 feedthrough
rlabel pdiffusion 171 -1497 171 -1497 0 feedthrough
rlabel pdiffusion 178 -1497 178 -1497 0 cellNo=126
rlabel pdiffusion 185 -1497 185 -1497 0 cellNo=547
rlabel pdiffusion 192 -1497 192 -1497 0 feedthrough
rlabel pdiffusion 199 -1497 199 -1497 0 feedthrough
rlabel pdiffusion 206 -1497 206 -1497 0 feedthrough
rlabel pdiffusion 213 -1497 213 -1497 0 feedthrough
rlabel pdiffusion 220 -1497 220 -1497 0 cellNo=179
rlabel pdiffusion 227 -1497 227 -1497 0 cellNo=240
rlabel pdiffusion 234 -1497 234 -1497 0 feedthrough
rlabel pdiffusion 241 -1497 241 -1497 0 cellNo=966
rlabel pdiffusion 248 -1497 248 -1497 0 feedthrough
rlabel pdiffusion 255 -1497 255 -1497 0 feedthrough
rlabel pdiffusion 262 -1497 262 -1497 0 feedthrough
rlabel pdiffusion 269 -1497 269 -1497 0 feedthrough
rlabel pdiffusion 276 -1497 276 -1497 0 feedthrough
rlabel pdiffusion 283 -1497 283 -1497 0 feedthrough
rlabel pdiffusion 290 -1497 290 -1497 0 cellNo=700
rlabel pdiffusion 297 -1497 297 -1497 0 feedthrough
rlabel pdiffusion 304 -1497 304 -1497 0 cellNo=529
rlabel pdiffusion 311 -1497 311 -1497 0 cellNo=117
rlabel pdiffusion 318 -1497 318 -1497 0 cellNo=904
rlabel pdiffusion 325 -1497 325 -1497 0 feedthrough
rlabel pdiffusion 332 -1497 332 -1497 0 feedthrough
rlabel pdiffusion 339 -1497 339 -1497 0 feedthrough
rlabel pdiffusion 346 -1497 346 -1497 0 feedthrough
rlabel pdiffusion 353 -1497 353 -1497 0 feedthrough
rlabel pdiffusion 360 -1497 360 -1497 0 feedthrough
rlabel pdiffusion 367 -1497 367 -1497 0 feedthrough
rlabel pdiffusion 374 -1497 374 -1497 0 feedthrough
rlabel pdiffusion 381 -1497 381 -1497 0 feedthrough
rlabel pdiffusion 388 -1497 388 -1497 0 feedthrough
rlabel pdiffusion 395 -1497 395 -1497 0 cellNo=705
rlabel pdiffusion 402 -1497 402 -1497 0 feedthrough
rlabel pdiffusion 409 -1497 409 -1497 0 feedthrough
rlabel pdiffusion 416 -1497 416 -1497 0 cellNo=781
rlabel pdiffusion 423 -1497 423 -1497 0 feedthrough
rlabel pdiffusion 430 -1497 430 -1497 0 feedthrough
rlabel pdiffusion 437 -1497 437 -1497 0 cellNo=838
rlabel pdiffusion 444 -1497 444 -1497 0 feedthrough
rlabel pdiffusion 451 -1497 451 -1497 0 feedthrough
rlabel pdiffusion 458 -1497 458 -1497 0 feedthrough
rlabel pdiffusion 465 -1497 465 -1497 0 feedthrough
rlabel pdiffusion 472 -1497 472 -1497 0 feedthrough
rlabel pdiffusion 479 -1497 479 -1497 0 feedthrough
rlabel pdiffusion 486 -1497 486 -1497 0 feedthrough
rlabel pdiffusion 493 -1497 493 -1497 0 feedthrough
rlabel pdiffusion 500 -1497 500 -1497 0 cellNo=293
rlabel pdiffusion 507 -1497 507 -1497 0 feedthrough
rlabel pdiffusion 514 -1497 514 -1497 0 feedthrough
rlabel pdiffusion 521 -1497 521 -1497 0 feedthrough
rlabel pdiffusion 528 -1497 528 -1497 0 feedthrough
rlabel pdiffusion 535 -1497 535 -1497 0 cellNo=6
rlabel pdiffusion 542 -1497 542 -1497 0 cellNo=422
rlabel pdiffusion 549 -1497 549 -1497 0 feedthrough
rlabel pdiffusion 556 -1497 556 -1497 0 cellNo=632
rlabel pdiffusion 563 -1497 563 -1497 0 cellNo=342
rlabel pdiffusion 570 -1497 570 -1497 0 feedthrough
rlabel pdiffusion 577 -1497 577 -1497 0 cellNo=937
rlabel pdiffusion 584 -1497 584 -1497 0 feedthrough
rlabel pdiffusion 591 -1497 591 -1497 0 feedthrough
rlabel pdiffusion 598 -1497 598 -1497 0 feedthrough
rlabel pdiffusion 605 -1497 605 -1497 0 feedthrough
rlabel pdiffusion 612 -1497 612 -1497 0 feedthrough
rlabel pdiffusion 619 -1497 619 -1497 0 cellNo=676
rlabel pdiffusion 626 -1497 626 -1497 0 feedthrough
rlabel pdiffusion 633 -1497 633 -1497 0 cellNo=497
rlabel pdiffusion 640 -1497 640 -1497 0 feedthrough
rlabel pdiffusion 647 -1497 647 -1497 0 feedthrough
rlabel pdiffusion 654 -1497 654 -1497 0 cellNo=229
rlabel pdiffusion 661 -1497 661 -1497 0 feedthrough
rlabel pdiffusion 668 -1497 668 -1497 0 feedthrough
rlabel pdiffusion 675 -1497 675 -1497 0 feedthrough
rlabel pdiffusion 682 -1497 682 -1497 0 cellNo=847
rlabel pdiffusion 689 -1497 689 -1497 0 feedthrough
rlabel pdiffusion 696 -1497 696 -1497 0 feedthrough
rlabel pdiffusion 703 -1497 703 -1497 0 feedthrough
rlabel pdiffusion 710 -1497 710 -1497 0 feedthrough
rlabel pdiffusion 717 -1497 717 -1497 0 feedthrough
rlabel pdiffusion 724 -1497 724 -1497 0 cellNo=737
rlabel pdiffusion 731 -1497 731 -1497 0 feedthrough
rlabel pdiffusion 738 -1497 738 -1497 0 feedthrough
rlabel pdiffusion 745 -1497 745 -1497 0 feedthrough
rlabel pdiffusion 752 -1497 752 -1497 0 feedthrough
rlabel pdiffusion 759 -1497 759 -1497 0 feedthrough
rlabel pdiffusion 766 -1497 766 -1497 0 feedthrough
rlabel pdiffusion 773 -1497 773 -1497 0 feedthrough
rlabel pdiffusion 780 -1497 780 -1497 0 feedthrough
rlabel pdiffusion 787 -1497 787 -1497 0 feedthrough
rlabel pdiffusion 794 -1497 794 -1497 0 feedthrough
rlabel pdiffusion 801 -1497 801 -1497 0 cellNo=868
rlabel pdiffusion 808 -1497 808 -1497 0 feedthrough
rlabel pdiffusion 815 -1497 815 -1497 0 feedthrough
rlabel pdiffusion 822 -1497 822 -1497 0 feedthrough
rlabel pdiffusion 829 -1497 829 -1497 0 feedthrough
rlabel pdiffusion 836 -1497 836 -1497 0 feedthrough
rlabel pdiffusion 843 -1497 843 -1497 0 feedthrough
rlabel pdiffusion 850 -1497 850 -1497 0 feedthrough
rlabel pdiffusion 857 -1497 857 -1497 0 feedthrough
rlabel pdiffusion 864 -1497 864 -1497 0 feedthrough
rlabel pdiffusion 871 -1497 871 -1497 0 feedthrough
rlabel pdiffusion 878 -1497 878 -1497 0 feedthrough
rlabel pdiffusion 885 -1497 885 -1497 0 feedthrough
rlabel pdiffusion 892 -1497 892 -1497 0 feedthrough
rlabel pdiffusion 899 -1497 899 -1497 0 feedthrough
rlabel pdiffusion 906 -1497 906 -1497 0 feedthrough
rlabel pdiffusion 913 -1497 913 -1497 0 feedthrough
rlabel pdiffusion 920 -1497 920 -1497 0 cellNo=527
rlabel pdiffusion 927 -1497 927 -1497 0 feedthrough
rlabel pdiffusion 934 -1497 934 -1497 0 feedthrough
rlabel pdiffusion 941 -1497 941 -1497 0 cellNo=892
rlabel pdiffusion 948 -1497 948 -1497 0 feedthrough
rlabel pdiffusion 955 -1497 955 -1497 0 feedthrough
rlabel pdiffusion 962 -1497 962 -1497 0 cellNo=68
rlabel pdiffusion 969 -1497 969 -1497 0 cellNo=785
rlabel pdiffusion 976 -1497 976 -1497 0 feedthrough
rlabel pdiffusion 983 -1497 983 -1497 0 feedthrough
rlabel pdiffusion 990 -1497 990 -1497 0 feedthrough
rlabel pdiffusion 997 -1497 997 -1497 0 feedthrough
rlabel pdiffusion 1004 -1497 1004 -1497 0 feedthrough
rlabel pdiffusion 1039 -1497 1039 -1497 0 feedthrough
rlabel pdiffusion 1067 -1497 1067 -1497 0 cellNo=116
rlabel pdiffusion 3 -1594 3 -1594 0 feedthrough
rlabel pdiffusion 10 -1594 10 -1594 0 feedthrough
rlabel pdiffusion 17 -1594 17 -1594 0 feedthrough
rlabel pdiffusion 24 -1594 24 -1594 0 feedthrough
rlabel pdiffusion 31 -1594 31 -1594 0 feedthrough
rlabel pdiffusion 38 -1594 38 -1594 0 feedthrough
rlabel pdiffusion 45 -1594 45 -1594 0 cellNo=982
rlabel pdiffusion 52 -1594 52 -1594 0 feedthrough
rlabel pdiffusion 59 -1594 59 -1594 0 feedthrough
rlabel pdiffusion 66 -1594 66 -1594 0 feedthrough
rlabel pdiffusion 73 -1594 73 -1594 0 cellNo=206
rlabel pdiffusion 80 -1594 80 -1594 0 cellNo=516
rlabel pdiffusion 87 -1594 87 -1594 0 feedthrough
rlabel pdiffusion 94 -1594 94 -1594 0 feedthrough
rlabel pdiffusion 101 -1594 101 -1594 0 feedthrough
rlabel pdiffusion 108 -1594 108 -1594 0 feedthrough
rlabel pdiffusion 115 -1594 115 -1594 0 feedthrough
rlabel pdiffusion 122 -1594 122 -1594 0 cellNo=831
rlabel pdiffusion 129 -1594 129 -1594 0 feedthrough
rlabel pdiffusion 136 -1594 136 -1594 0 feedthrough
rlabel pdiffusion 143 -1594 143 -1594 0 feedthrough
rlabel pdiffusion 150 -1594 150 -1594 0 feedthrough
rlabel pdiffusion 157 -1594 157 -1594 0 feedthrough
rlabel pdiffusion 164 -1594 164 -1594 0 feedthrough
rlabel pdiffusion 171 -1594 171 -1594 0 feedthrough
rlabel pdiffusion 178 -1594 178 -1594 0 feedthrough
rlabel pdiffusion 185 -1594 185 -1594 0 feedthrough
rlabel pdiffusion 192 -1594 192 -1594 0 cellNo=704
rlabel pdiffusion 199 -1594 199 -1594 0 feedthrough
rlabel pdiffusion 206 -1594 206 -1594 0 feedthrough
rlabel pdiffusion 213 -1594 213 -1594 0 feedthrough
rlabel pdiffusion 220 -1594 220 -1594 0 cellNo=689
rlabel pdiffusion 227 -1594 227 -1594 0 cellNo=709
rlabel pdiffusion 234 -1594 234 -1594 0 cellNo=479
rlabel pdiffusion 241 -1594 241 -1594 0 cellNo=961
rlabel pdiffusion 248 -1594 248 -1594 0 cellNo=638
rlabel pdiffusion 255 -1594 255 -1594 0 feedthrough
rlabel pdiffusion 262 -1594 262 -1594 0 feedthrough
rlabel pdiffusion 269 -1594 269 -1594 0 feedthrough
rlabel pdiffusion 276 -1594 276 -1594 0 feedthrough
rlabel pdiffusion 283 -1594 283 -1594 0 feedthrough
rlabel pdiffusion 290 -1594 290 -1594 0 feedthrough
rlabel pdiffusion 297 -1594 297 -1594 0 feedthrough
rlabel pdiffusion 304 -1594 304 -1594 0 feedthrough
rlabel pdiffusion 311 -1594 311 -1594 0 feedthrough
rlabel pdiffusion 318 -1594 318 -1594 0 feedthrough
rlabel pdiffusion 325 -1594 325 -1594 0 cellNo=334
rlabel pdiffusion 332 -1594 332 -1594 0 feedthrough
rlabel pdiffusion 339 -1594 339 -1594 0 cellNo=87
rlabel pdiffusion 346 -1594 346 -1594 0 feedthrough
rlabel pdiffusion 353 -1594 353 -1594 0 cellNo=65
rlabel pdiffusion 360 -1594 360 -1594 0 cellNo=418
rlabel pdiffusion 367 -1594 367 -1594 0 feedthrough
rlabel pdiffusion 374 -1594 374 -1594 0 cellNo=873
rlabel pdiffusion 381 -1594 381 -1594 0 feedthrough
rlabel pdiffusion 388 -1594 388 -1594 0 feedthrough
rlabel pdiffusion 395 -1594 395 -1594 0 cellNo=388
rlabel pdiffusion 402 -1594 402 -1594 0 cellNo=290
rlabel pdiffusion 409 -1594 409 -1594 0 feedthrough
rlabel pdiffusion 416 -1594 416 -1594 0 cellNo=941
rlabel pdiffusion 423 -1594 423 -1594 0 feedthrough
rlabel pdiffusion 430 -1594 430 -1594 0 feedthrough
rlabel pdiffusion 437 -1594 437 -1594 0 cellNo=840
rlabel pdiffusion 444 -1594 444 -1594 0 feedthrough
rlabel pdiffusion 451 -1594 451 -1594 0 cellNo=930
rlabel pdiffusion 458 -1594 458 -1594 0 cellNo=711
rlabel pdiffusion 465 -1594 465 -1594 0 feedthrough
rlabel pdiffusion 472 -1594 472 -1594 0 cellNo=466
rlabel pdiffusion 479 -1594 479 -1594 0 feedthrough
rlabel pdiffusion 486 -1594 486 -1594 0 feedthrough
rlabel pdiffusion 493 -1594 493 -1594 0 cellNo=312
rlabel pdiffusion 500 -1594 500 -1594 0 feedthrough
rlabel pdiffusion 507 -1594 507 -1594 0 cellNo=419
rlabel pdiffusion 514 -1594 514 -1594 0 cellNo=114
rlabel pdiffusion 521 -1594 521 -1594 0 feedthrough
rlabel pdiffusion 528 -1594 528 -1594 0 feedthrough
rlabel pdiffusion 535 -1594 535 -1594 0 cellNo=799
rlabel pdiffusion 542 -1594 542 -1594 0 cellNo=748
rlabel pdiffusion 549 -1594 549 -1594 0 feedthrough
rlabel pdiffusion 556 -1594 556 -1594 0 feedthrough
rlabel pdiffusion 563 -1594 563 -1594 0 feedthrough
rlabel pdiffusion 570 -1594 570 -1594 0 feedthrough
rlabel pdiffusion 577 -1594 577 -1594 0 feedthrough
rlabel pdiffusion 584 -1594 584 -1594 0 feedthrough
rlabel pdiffusion 591 -1594 591 -1594 0 feedthrough
rlabel pdiffusion 598 -1594 598 -1594 0 feedthrough
rlabel pdiffusion 605 -1594 605 -1594 0 feedthrough
rlabel pdiffusion 612 -1594 612 -1594 0 feedthrough
rlabel pdiffusion 619 -1594 619 -1594 0 feedthrough
rlabel pdiffusion 626 -1594 626 -1594 0 feedthrough
rlabel pdiffusion 633 -1594 633 -1594 0 feedthrough
rlabel pdiffusion 640 -1594 640 -1594 0 feedthrough
rlabel pdiffusion 647 -1594 647 -1594 0 feedthrough
rlabel pdiffusion 654 -1594 654 -1594 0 feedthrough
rlabel pdiffusion 661 -1594 661 -1594 0 cellNo=99
rlabel pdiffusion 668 -1594 668 -1594 0 feedthrough
rlabel pdiffusion 675 -1594 675 -1594 0 feedthrough
rlabel pdiffusion 682 -1594 682 -1594 0 cellNo=149
rlabel pdiffusion 689 -1594 689 -1594 0 feedthrough
rlabel pdiffusion 696 -1594 696 -1594 0 feedthrough
rlabel pdiffusion 703 -1594 703 -1594 0 feedthrough
rlabel pdiffusion 710 -1594 710 -1594 0 cellNo=205
rlabel pdiffusion 717 -1594 717 -1594 0 feedthrough
rlabel pdiffusion 724 -1594 724 -1594 0 feedthrough
rlabel pdiffusion 731 -1594 731 -1594 0 cellNo=248
rlabel pdiffusion 738 -1594 738 -1594 0 feedthrough
rlabel pdiffusion 745 -1594 745 -1594 0 feedthrough
rlabel pdiffusion 752 -1594 752 -1594 0 feedthrough
rlabel pdiffusion 759 -1594 759 -1594 0 cellNo=131
rlabel pdiffusion 766 -1594 766 -1594 0 feedthrough
rlabel pdiffusion 773 -1594 773 -1594 0 feedthrough
rlabel pdiffusion 780 -1594 780 -1594 0 feedthrough
rlabel pdiffusion 787 -1594 787 -1594 0 feedthrough
rlabel pdiffusion 794 -1594 794 -1594 0 feedthrough
rlabel pdiffusion 801 -1594 801 -1594 0 cellNo=433
rlabel pdiffusion 808 -1594 808 -1594 0 feedthrough
rlabel pdiffusion 815 -1594 815 -1594 0 feedthrough
rlabel pdiffusion 822 -1594 822 -1594 0 feedthrough
rlabel pdiffusion 829 -1594 829 -1594 0 feedthrough
rlabel pdiffusion 836 -1594 836 -1594 0 feedthrough
rlabel pdiffusion 843 -1594 843 -1594 0 feedthrough
rlabel pdiffusion 850 -1594 850 -1594 0 feedthrough
rlabel pdiffusion 857 -1594 857 -1594 0 feedthrough
rlabel pdiffusion 864 -1594 864 -1594 0 feedthrough
rlabel pdiffusion 871 -1594 871 -1594 0 feedthrough
rlabel pdiffusion 878 -1594 878 -1594 0 feedthrough
rlabel pdiffusion 885 -1594 885 -1594 0 feedthrough
rlabel pdiffusion 892 -1594 892 -1594 0 feedthrough
rlabel pdiffusion 899 -1594 899 -1594 0 feedthrough
rlabel pdiffusion 906 -1594 906 -1594 0 feedthrough
rlabel pdiffusion 913 -1594 913 -1594 0 feedthrough
rlabel pdiffusion 920 -1594 920 -1594 0 feedthrough
rlabel pdiffusion 927 -1594 927 -1594 0 feedthrough
rlabel pdiffusion 934 -1594 934 -1594 0 feedthrough
rlabel pdiffusion 941 -1594 941 -1594 0 feedthrough
rlabel pdiffusion 948 -1594 948 -1594 0 feedthrough
rlabel pdiffusion 955 -1594 955 -1594 0 feedthrough
rlabel pdiffusion 962 -1594 962 -1594 0 feedthrough
rlabel pdiffusion 969 -1594 969 -1594 0 feedthrough
rlabel pdiffusion 976 -1594 976 -1594 0 feedthrough
rlabel pdiffusion 983 -1594 983 -1594 0 feedthrough
rlabel pdiffusion 990 -1594 990 -1594 0 feedthrough
rlabel pdiffusion 997 -1594 997 -1594 0 feedthrough
rlabel pdiffusion 1004 -1594 1004 -1594 0 feedthrough
rlabel pdiffusion 1011 -1594 1011 -1594 0 feedthrough
rlabel pdiffusion 1018 -1594 1018 -1594 0 feedthrough
rlabel pdiffusion 1025 -1594 1025 -1594 0 feedthrough
rlabel pdiffusion 1032 -1594 1032 -1594 0 feedthrough
rlabel pdiffusion 1039 -1594 1039 -1594 0 feedthrough
rlabel pdiffusion 1046 -1594 1046 -1594 0 feedthrough
rlabel pdiffusion 1053 -1594 1053 -1594 0 feedthrough
rlabel pdiffusion 1060 -1594 1060 -1594 0 feedthrough
rlabel pdiffusion 1067 -1594 1067 -1594 0 feedthrough
rlabel pdiffusion 1074 -1594 1074 -1594 0 feedthrough
rlabel pdiffusion 1081 -1594 1081 -1594 0 feedthrough
rlabel pdiffusion 1088 -1594 1088 -1594 0 feedthrough
rlabel pdiffusion 1095 -1594 1095 -1594 0 feedthrough
rlabel pdiffusion 1102 -1594 1102 -1594 0 feedthrough
rlabel pdiffusion 1109 -1594 1109 -1594 0 cellNo=299
rlabel pdiffusion 3 -1681 3 -1681 0 feedthrough
rlabel pdiffusion 10 -1681 10 -1681 0 feedthrough
rlabel pdiffusion 17 -1681 17 -1681 0 feedthrough
rlabel pdiffusion 24 -1681 24 -1681 0 feedthrough
rlabel pdiffusion 31 -1681 31 -1681 0 feedthrough
rlabel pdiffusion 38 -1681 38 -1681 0 feedthrough
rlabel pdiffusion 45 -1681 45 -1681 0 feedthrough
rlabel pdiffusion 52 -1681 52 -1681 0 feedthrough
rlabel pdiffusion 59 -1681 59 -1681 0 cellNo=829
rlabel pdiffusion 66 -1681 66 -1681 0 feedthrough
rlabel pdiffusion 73 -1681 73 -1681 0 feedthrough
rlabel pdiffusion 80 -1681 80 -1681 0 cellNo=152
rlabel pdiffusion 87 -1681 87 -1681 0 feedthrough
rlabel pdiffusion 94 -1681 94 -1681 0 cellNo=659
rlabel pdiffusion 101 -1681 101 -1681 0 feedthrough
rlabel pdiffusion 108 -1681 108 -1681 0 feedthrough
rlabel pdiffusion 115 -1681 115 -1681 0 feedthrough
rlabel pdiffusion 122 -1681 122 -1681 0 feedthrough
rlabel pdiffusion 129 -1681 129 -1681 0 feedthrough
rlabel pdiffusion 136 -1681 136 -1681 0 cellNo=872
rlabel pdiffusion 143 -1681 143 -1681 0 feedthrough
rlabel pdiffusion 150 -1681 150 -1681 0 cellNo=828
rlabel pdiffusion 157 -1681 157 -1681 0 cellNo=407
rlabel pdiffusion 164 -1681 164 -1681 0 feedthrough
rlabel pdiffusion 171 -1681 171 -1681 0 feedthrough
rlabel pdiffusion 178 -1681 178 -1681 0 feedthrough
rlabel pdiffusion 185 -1681 185 -1681 0 feedthrough
rlabel pdiffusion 192 -1681 192 -1681 0 cellNo=10
rlabel pdiffusion 199 -1681 199 -1681 0 cellNo=59
rlabel pdiffusion 206 -1681 206 -1681 0 feedthrough
rlabel pdiffusion 213 -1681 213 -1681 0 cellNo=928
rlabel pdiffusion 220 -1681 220 -1681 0 cellNo=90
rlabel pdiffusion 227 -1681 227 -1681 0 cellNo=954
rlabel pdiffusion 234 -1681 234 -1681 0 cellNo=678
rlabel pdiffusion 241 -1681 241 -1681 0 feedthrough
rlabel pdiffusion 248 -1681 248 -1681 0 feedthrough
rlabel pdiffusion 255 -1681 255 -1681 0 feedthrough
rlabel pdiffusion 262 -1681 262 -1681 0 feedthrough
rlabel pdiffusion 269 -1681 269 -1681 0 feedthrough
rlabel pdiffusion 276 -1681 276 -1681 0 feedthrough
rlabel pdiffusion 283 -1681 283 -1681 0 cellNo=811
rlabel pdiffusion 290 -1681 290 -1681 0 cellNo=169
rlabel pdiffusion 297 -1681 297 -1681 0 cellNo=54
rlabel pdiffusion 304 -1681 304 -1681 0 feedthrough
rlabel pdiffusion 311 -1681 311 -1681 0 feedthrough
rlabel pdiffusion 318 -1681 318 -1681 0 feedthrough
rlabel pdiffusion 325 -1681 325 -1681 0 feedthrough
rlabel pdiffusion 332 -1681 332 -1681 0 feedthrough
rlabel pdiffusion 339 -1681 339 -1681 0 feedthrough
rlabel pdiffusion 346 -1681 346 -1681 0 cellNo=9
rlabel pdiffusion 353 -1681 353 -1681 0 feedthrough
rlabel pdiffusion 360 -1681 360 -1681 0 feedthrough
rlabel pdiffusion 367 -1681 367 -1681 0 cellNo=750
rlabel pdiffusion 374 -1681 374 -1681 0 feedthrough
rlabel pdiffusion 381 -1681 381 -1681 0 cellNo=976
rlabel pdiffusion 388 -1681 388 -1681 0 cellNo=301
rlabel pdiffusion 395 -1681 395 -1681 0 feedthrough
rlabel pdiffusion 402 -1681 402 -1681 0 feedthrough
rlabel pdiffusion 409 -1681 409 -1681 0 feedthrough
rlabel pdiffusion 416 -1681 416 -1681 0 feedthrough
rlabel pdiffusion 423 -1681 423 -1681 0 feedthrough
rlabel pdiffusion 430 -1681 430 -1681 0 feedthrough
rlabel pdiffusion 437 -1681 437 -1681 0 feedthrough
rlabel pdiffusion 444 -1681 444 -1681 0 feedthrough
rlabel pdiffusion 451 -1681 451 -1681 0 cellNo=885
rlabel pdiffusion 458 -1681 458 -1681 0 feedthrough
rlabel pdiffusion 465 -1681 465 -1681 0 cellNo=244
rlabel pdiffusion 472 -1681 472 -1681 0 cellNo=977
rlabel pdiffusion 479 -1681 479 -1681 0 cellNo=145
rlabel pdiffusion 486 -1681 486 -1681 0 cellNo=965
rlabel pdiffusion 493 -1681 493 -1681 0 cellNo=875
rlabel pdiffusion 500 -1681 500 -1681 0 feedthrough
rlabel pdiffusion 507 -1681 507 -1681 0 feedthrough
rlabel pdiffusion 514 -1681 514 -1681 0 feedthrough
rlabel pdiffusion 521 -1681 521 -1681 0 feedthrough
rlabel pdiffusion 528 -1681 528 -1681 0 feedthrough
rlabel pdiffusion 535 -1681 535 -1681 0 cellNo=825
rlabel pdiffusion 542 -1681 542 -1681 0 feedthrough
rlabel pdiffusion 549 -1681 549 -1681 0 cellNo=185
rlabel pdiffusion 556 -1681 556 -1681 0 cellNo=665
rlabel pdiffusion 563 -1681 563 -1681 0 cellNo=802
rlabel pdiffusion 570 -1681 570 -1681 0 feedthrough
rlabel pdiffusion 577 -1681 577 -1681 0 feedthrough
rlabel pdiffusion 584 -1681 584 -1681 0 feedthrough
rlabel pdiffusion 591 -1681 591 -1681 0 feedthrough
rlabel pdiffusion 598 -1681 598 -1681 0 feedthrough
rlabel pdiffusion 605 -1681 605 -1681 0 feedthrough
rlabel pdiffusion 612 -1681 612 -1681 0 feedthrough
rlabel pdiffusion 619 -1681 619 -1681 0 feedthrough
rlabel pdiffusion 626 -1681 626 -1681 0 feedthrough
rlabel pdiffusion 633 -1681 633 -1681 0 feedthrough
rlabel pdiffusion 640 -1681 640 -1681 0 feedthrough
rlabel pdiffusion 647 -1681 647 -1681 0 feedthrough
rlabel pdiffusion 654 -1681 654 -1681 0 feedthrough
rlabel pdiffusion 661 -1681 661 -1681 0 feedthrough
rlabel pdiffusion 668 -1681 668 -1681 0 feedthrough
rlabel pdiffusion 675 -1681 675 -1681 0 feedthrough
rlabel pdiffusion 682 -1681 682 -1681 0 feedthrough
rlabel pdiffusion 689 -1681 689 -1681 0 feedthrough
rlabel pdiffusion 696 -1681 696 -1681 0 feedthrough
rlabel pdiffusion 703 -1681 703 -1681 0 feedthrough
rlabel pdiffusion 710 -1681 710 -1681 0 feedthrough
rlabel pdiffusion 717 -1681 717 -1681 0 feedthrough
rlabel pdiffusion 724 -1681 724 -1681 0 feedthrough
rlabel pdiffusion 731 -1681 731 -1681 0 cellNo=102
rlabel pdiffusion 738 -1681 738 -1681 0 feedthrough
rlabel pdiffusion 745 -1681 745 -1681 0 feedthrough
rlabel pdiffusion 752 -1681 752 -1681 0 feedthrough
rlabel pdiffusion 759 -1681 759 -1681 0 feedthrough
rlabel pdiffusion 766 -1681 766 -1681 0 feedthrough
rlabel pdiffusion 773 -1681 773 -1681 0 feedthrough
rlabel pdiffusion 780 -1681 780 -1681 0 feedthrough
rlabel pdiffusion 787 -1681 787 -1681 0 feedthrough
rlabel pdiffusion 794 -1681 794 -1681 0 feedthrough
rlabel pdiffusion 801 -1681 801 -1681 0 feedthrough
rlabel pdiffusion 808 -1681 808 -1681 0 feedthrough
rlabel pdiffusion 815 -1681 815 -1681 0 feedthrough
rlabel pdiffusion 822 -1681 822 -1681 0 cellNo=127
rlabel pdiffusion 829 -1681 829 -1681 0 feedthrough
rlabel pdiffusion 836 -1681 836 -1681 0 feedthrough
rlabel pdiffusion 843 -1681 843 -1681 0 feedthrough
rlabel pdiffusion 850 -1681 850 -1681 0 feedthrough
rlabel pdiffusion 857 -1681 857 -1681 0 feedthrough
rlabel pdiffusion 864 -1681 864 -1681 0 feedthrough
rlabel pdiffusion 871 -1681 871 -1681 0 feedthrough
rlabel pdiffusion 878 -1681 878 -1681 0 feedthrough
rlabel pdiffusion 885 -1681 885 -1681 0 cellNo=461
rlabel pdiffusion 892 -1681 892 -1681 0 cellNo=69
rlabel pdiffusion 899 -1681 899 -1681 0 feedthrough
rlabel pdiffusion 906 -1681 906 -1681 0 feedthrough
rlabel pdiffusion 913 -1681 913 -1681 0 cellNo=647
rlabel pdiffusion 920 -1681 920 -1681 0 feedthrough
rlabel pdiffusion 927 -1681 927 -1681 0 feedthrough
rlabel pdiffusion 934 -1681 934 -1681 0 feedthrough
rlabel pdiffusion 941 -1681 941 -1681 0 feedthrough
rlabel pdiffusion 948 -1681 948 -1681 0 feedthrough
rlabel pdiffusion 955 -1681 955 -1681 0 feedthrough
rlabel pdiffusion 962 -1681 962 -1681 0 feedthrough
rlabel pdiffusion 976 -1681 976 -1681 0 feedthrough
rlabel pdiffusion 983 -1681 983 -1681 0 feedthrough
rlabel pdiffusion 1004 -1681 1004 -1681 0 feedthrough
rlabel pdiffusion 1025 -1681 1025 -1681 0 cellNo=5
rlabel pdiffusion 1053 -1681 1053 -1681 0 feedthrough
rlabel pdiffusion 3 -1776 3 -1776 0 feedthrough
rlabel pdiffusion 10 -1776 10 -1776 0 cellNo=739
rlabel pdiffusion 17 -1776 17 -1776 0 cellNo=994
rlabel pdiffusion 24 -1776 24 -1776 0 feedthrough
rlabel pdiffusion 31 -1776 31 -1776 0 feedthrough
rlabel pdiffusion 38 -1776 38 -1776 0 feedthrough
rlabel pdiffusion 45 -1776 45 -1776 0 feedthrough
rlabel pdiffusion 52 -1776 52 -1776 0 cellNo=233
rlabel pdiffusion 59 -1776 59 -1776 0 cellNo=958
rlabel pdiffusion 66 -1776 66 -1776 0 feedthrough
rlabel pdiffusion 73 -1776 73 -1776 0 feedthrough
rlabel pdiffusion 80 -1776 80 -1776 0 feedthrough
rlabel pdiffusion 87 -1776 87 -1776 0 feedthrough
rlabel pdiffusion 94 -1776 94 -1776 0 feedthrough
rlabel pdiffusion 101 -1776 101 -1776 0 cellNo=839
rlabel pdiffusion 108 -1776 108 -1776 0 cellNo=685
rlabel pdiffusion 115 -1776 115 -1776 0 feedthrough
rlabel pdiffusion 122 -1776 122 -1776 0 feedthrough
rlabel pdiffusion 129 -1776 129 -1776 0 feedthrough
rlabel pdiffusion 136 -1776 136 -1776 0 feedthrough
rlabel pdiffusion 143 -1776 143 -1776 0 feedthrough
rlabel pdiffusion 150 -1776 150 -1776 0 cellNo=623
rlabel pdiffusion 157 -1776 157 -1776 0 feedthrough
rlabel pdiffusion 164 -1776 164 -1776 0 cellNo=646
rlabel pdiffusion 171 -1776 171 -1776 0 feedthrough
rlabel pdiffusion 178 -1776 178 -1776 0 cellNo=436
rlabel pdiffusion 185 -1776 185 -1776 0 cellNo=809
rlabel pdiffusion 192 -1776 192 -1776 0 feedthrough
rlabel pdiffusion 199 -1776 199 -1776 0 feedthrough
rlabel pdiffusion 206 -1776 206 -1776 0 feedthrough
rlabel pdiffusion 213 -1776 213 -1776 0 cellNo=143
rlabel pdiffusion 220 -1776 220 -1776 0 cellNo=644
rlabel pdiffusion 227 -1776 227 -1776 0 feedthrough
rlabel pdiffusion 234 -1776 234 -1776 0 feedthrough
rlabel pdiffusion 241 -1776 241 -1776 0 cellNo=142
rlabel pdiffusion 248 -1776 248 -1776 0 feedthrough
rlabel pdiffusion 255 -1776 255 -1776 0 feedthrough
rlabel pdiffusion 262 -1776 262 -1776 0 feedthrough
rlabel pdiffusion 269 -1776 269 -1776 0 feedthrough
rlabel pdiffusion 276 -1776 276 -1776 0 feedthrough
rlabel pdiffusion 283 -1776 283 -1776 0 feedthrough
rlabel pdiffusion 290 -1776 290 -1776 0 feedthrough
rlabel pdiffusion 297 -1776 297 -1776 0 feedthrough
rlabel pdiffusion 304 -1776 304 -1776 0 feedthrough
rlabel pdiffusion 311 -1776 311 -1776 0 cellNo=993
rlabel pdiffusion 318 -1776 318 -1776 0 feedthrough
rlabel pdiffusion 325 -1776 325 -1776 0 cellNo=78
rlabel pdiffusion 332 -1776 332 -1776 0 feedthrough
rlabel pdiffusion 339 -1776 339 -1776 0 feedthrough
rlabel pdiffusion 346 -1776 346 -1776 0 feedthrough
rlabel pdiffusion 353 -1776 353 -1776 0 feedthrough
rlabel pdiffusion 360 -1776 360 -1776 0 feedthrough
rlabel pdiffusion 367 -1776 367 -1776 0 cellNo=559
rlabel pdiffusion 374 -1776 374 -1776 0 cellNo=107
rlabel pdiffusion 381 -1776 381 -1776 0 cellNo=706
rlabel pdiffusion 388 -1776 388 -1776 0 feedthrough
rlabel pdiffusion 395 -1776 395 -1776 0 feedthrough
rlabel pdiffusion 402 -1776 402 -1776 0 cellNo=314
rlabel pdiffusion 409 -1776 409 -1776 0 cellNo=338
rlabel pdiffusion 416 -1776 416 -1776 0 feedthrough
rlabel pdiffusion 423 -1776 423 -1776 0 cellNo=441
rlabel pdiffusion 430 -1776 430 -1776 0 feedthrough
rlabel pdiffusion 437 -1776 437 -1776 0 feedthrough
rlabel pdiffusion 444 -1776 444 -1776 0 feedthrough
rlabel pdiffusion 451 -1776 451 -1776 0 feedthrough
rlabel pdiffusion 458 -1776 458 -1776 0 feedthrough
rlabel pdiffusion 465 -1776 465 -1776 0 cellNo=264
rlabel pdiffusion 472 -1776 472 -1776 0 feedthrough
rlabel pdiffusion 479 -1776 479 -1776 0 cellNo=617
rlabel pdiffusion 486 -1776 486 -1776 0 feedthrough
rlabel pdiffusion 493 -1776 493 -1776 0 feedthrough
rlabel pdiffusion 500 -1776 500 -1776 0 feedthrough
rlabel pdiffusion 507 -1776 507 -1776 0 feedthrough
rlabel pdiffusion 514 -1776 514 -1776 0 cellNo=998
rlabel pdiffusion 521 -1776 521 -1776 0 feedthrough
rlabel pdiffusion 528 -1776 528 -1776 0 feedthrough
rlabel pdiffusion 535 -1776 535 -1776 0 feedthrough
rlabel pdiffusion 542 -1776 542 -1776 0 cellNo=688
rlabel pdiffusion 549 -1776 549 -1776 0 feedthrough
rlabel pdiffusion 556 -1776 556 -1776 0 feedthrough
rlabel pdiffusion 563 -1776 563 -1776 0 feedthrough
rlabel pdiffusion 570 -1776 570 -1776 0 feedthrough
rlabel pdiffusion 577 -1776 577 -1776 0 feedthrough
rlabel pdiffusion 584 -1776 584 -1776 0 feedthrough
rlabel pdiffusion 591 -1776 591 -1776 0 cellNo=675
rlabel pdiffusion 598 -1776 598 -1776 0 feedthrough
rlabel pdiffusion 605 -1776 605 -1776 0 feedthrough
rlabel pdiffusion 612 -1776 612 -1776 0 cellNo=794
rlabel pdiffusion 619 -1776 619 -1776 0 cellNo=291
rlabel pdiffusion 626 -1776 626 -1776 0 feedthrough
rlabel pdiffusion 633 -1776 633 -1776 0 cellNo=350
rlabel pdiffusion 640 -1776 640 -1776 0 feedthrough
rlabel pdiffusion 647 -1776 647 -1776 0 cellNo=113
rlabel pdiffusion 654 -1776 654 -1776 0 cellNo=553
rlabel pdiffusion 661 -1776 661 -1776 0 feedthrough
rlabel pdiffusion 668 -1776 668 -1776 0 feedthrough
rlabel pdiffusion 675 -1776 675 -1776 0 cellNo=830
rlabel pdiffusion 682 -1776 682 -1776 0 feedthrough
rlabel pdiffusion 689 -1776 689 -1776 0 feedthrough
rlabel pdiffusion 696 -1776 696 -1776 0 feedthrough
rlabel pdiffusion 703 -1776 703 -1776 0 feedthrough
rlabel pdiffusion 710 -1776 710 -1776 0 feedthrough
rlabel pdiffusion 717 -1776 717 -1776 0 feedthrough
rlabel pdiffusion 724 -1776 724 -1776 0 feedthrough
rlabel pdiffusion 731 -1776 731 -1776 0 feedthrough
rlabel pdiffusion 738 -1776 738 -1776 0 feedthrough
rlabel pdiffusion 745 -1776 745 -1776 0 feedthrough
rlabel pdiffusion 752 -1776 752 -1776 0 feedthrough
rlabel pdiffusion 759 -1776 759 -1776 0 feedthrough
rlabel pdiffusion 766 -1776 766 -1776 0 feedthrough
rlabel pdiffusion 773 -1776 773 -1776 0 feedthrough
rlabel pdiffusion 780 -1776 780 -1776 0 feedthrough
rlabel pdiffusion 787 -1776 787 -1776 0 feedthrough
rlabel pdiffusion 794 -1776 794 -1776 0 feedthrough
rlabel pdiffusion 801 -1776 801 -1776 0 cellNo=656
rlabel pdiffusion 808 -1776 808 -1776 0 feedthrough
rlabel pdiffusion 815 -1776 815 -1776 0 feedthrough
rlabel pdiffusion 822 -1776 822 -1776 0 feedthrough
rlabel pdiffusion 829 -1776 829 -1776 0 feedthrough
rlabel pdiffusion 836 -1776 836 -1776 0 feedthrough
rlabel pdiffusion 843 -1776 843 -1776 0 feedthrough
rlabel pdiffusion 850 -1776 850 -1776 0 feedthrough
rlabel pdiffusion 857 -1776 857 -1776 0 feedthrough
rlabel pdiffusion 864 -1776 864 -1776 0 feedthrough
rlabel pdiffusion 871 -1776 871 -1776 0 feedthrough
rlabel pdiffusion 878 -1776 878 -1776 0 feedthrough
rlabel pdiffusion 885 -1776 885 -1776 0 feedthrough
rlabel pdiffusion 892 -1776 892 -1776 0 feedthrough
rlabel pdiffusion 899 -1776 899 -1776 0 feedthrough
rlabel pdiffusion 906 -1776 906 -1776 0 feedthrough
rlabel pdiffusion 913 -1776 913 -1776 0 feedthrough
rlabel pdiffusion 920 -1776 920 -1776 0 feedthrough
rlabel pdiffusion 927 -1776 927 -1776 0 feedthrough
rlabel pdiffusion 934 -1776 934 -1776 0 feedthrough
rlabel pdiffusion 941 -1776 941 -1776 0 feedthrough
rlabel pdiffusion 948 -1776 948 -1776 0 feedthrough
rlabel pdiffusion 955 -1776 955 -1776 0 feedthrough
rlabel pdiffusion 962 -1776 962 -1776 0 feedthrough
rlabel pdiffusion 969 -1776 969 -1776 0 feedthrough
rlabel pdiffusion 976 -1776 976 -1776 0 feedthrough
rlabel pdiffusion 983 -1776 983 -1776 0 feedthrough
rlabel pdiffusion 990 -1776 990 -1776 0 feedthrough
rlabel pdiffusion 997 -1776 997 -1776 0 cellNo=478
rlabel pdiffusion 1004 -1776 1004 -1776 0 cellNo=900
rlabel pdiffusion 1011 -1776 1011 -1776 0 feedthrough
rlabel pdiffusion 1018 -1776 1018 -1776 0 feedthrough
rlabel pdiffusion 1025 -1776 1025 -1776 0 feedthrough
rlabel pdiffusion 52 -1867 52 -1867 0 feedthrough
rlabel pdiffusion 59 -1867 59 -1867 0 feedthrough
rlabel pdiffusion 66 -1867 66 -1867 0 feedthrough
rlabel pdiffusion 73 -1867 73 -1867 0 feedthrough
rlabel pdiffusion 80 -1867 80 -1867 0 feedthrough
rlabel pdiffusion 87 -1867 87 -1867 0 feedthrough
rlabel pdiffusion 94 -1867 94 -1867 0 feedthrough
rlabel pdiffusion 101 -1867 101 -1867 0 feedthrough
rlabel pdiffusion 108 -1867 108 -1867 0 feedthrough
rlabel pdiffusion 115 -1867 115 -1867 0 feedthrough
rlabel pdiffusion 122 -1867 122 -1867 0 feedthrough
rlabel pdiffusion 129 -1867 129 -1867 0 cellNo=571
rlabel pdiffusion 136 -1867 136 -1867 0 feedthrough
rlabel pdiffusion 143 -1867 143 -1867 0 feedthrough
rlabel pdiffusion 150 -1867 150 -1867 0 feedthrough
rlabel pdiffusion 157 -1867 157 -1867 0 feedthrough
rlabel pdiffusion 164 -1867 164 -1867 0 cellNo=570
rlabel pdiffusion 171 -1867 171 -1867 0 feedthrough
rlabel pdiffusion 178 -1867 178 -1867 0 feedthrough
rlabel pdiffusion 185 -1867 185 -1867 0 feedthrough
rlabel pdiffusion 192 -1867 192 -1867 0 cellNo=260
rlabel pdiffusion 199 -1867 199 -1867 0 cellNo=249
rlabel pdiffusion 206 -1867 206 -1867 0 cellNo=270
rlabel pdiffusion 213 -1867 213 -1867 0 cellNo=139
rlabel pdiffusion 220 -1867 220 -1867 0 cellNo=886
rlabel pdiffusion 227 -1867 227 -1867 0 cellNo=766
rlabel pdiffusion 234 -1867 234 -1867 0 feedthrough
rlabel pdiffusion 241 -1867 241 -1867 0 cellNo=387
rlabel pdiffusion 248 -1867 248 -1867 0 feedthrough
rlabel pdiffusion 255 -1867 255 -1867 0 feedthrough
rlabel pdiffusion 262 -1867 262 -1867 0 feedthrough
rlabel pdiffusion 269 -1867 269 -1867 0 feedthrough
rlabel pdiffusion 276 -1867 276 -1867 0 feedthrough
rlabel pdiffusion 283 -1867 283 -1867 0 feedthrough
rlabel pdiffusion 290 -1867 290 -1867 0 feedthrough
rlabel pdiffusion 297 -1867 297 -1867 0 feedthrough
rlabel pdiffusion 304 -1867 304 -1867 0 feedthrough
rlabel pdiffusion 311 -1867 311 -1867 0 feedthrough
rlabel pdiffusion 318 -1867 318 -1867 0 feedthrough
rlabel pdiffusion 325 -1867 325 -1867 0 feedthrough
rlabel pdiffusion 332 -1867 332 -1867 0 feedthrough
rlabel pdiffusion 339 -1867 339 -1867 0 feedthrough
rlabel pdiffusion 346 -1867 346 -1867 0 cellNo=17
rlabel pdiffusion 353 -1867 353 -1867 0 feedthrough
rlabel pdiffusion 360 -1867 360 -1867 0 cellNo=406
rlabel pdiffusion 367 -1867 367 -1867 0 cellNo=674
rlabel pdiffusion 374 -1867 374 -1867 0 feedthrough
rlabel pdiffusion 381 -1867 381 -1867 0 feedthrough
rlabel pdiffusion 388 -1867 388 -1867 0 feedthrough
rlabel pdiffusion 395 -1867 395 -1867 0 feedthrough
rlabel pdiffusion 402 -1867 402 -1867 0 feedthrough
rlabel pdiffusion 409 -1867 409 -1867 0 cellNo=443
rlabel pdiffusion 416 -1867 416 -1867 0 cellNo=898
rlabel pdiffusion 423 -1867 423 -1867 0 cellNo=51
rlabel pdiffusion 430 -1867 430 -1867 0 feedthrough
rlabel pdiffusion 437 -1867 437 -1867 0 feedthrough
rlabel pdiffusion 444 -1867 444 -1867 0 feedthrough
rlabel pdiffusion 451 -1867 451 -1867 0 feedthrough
rlabel pdiffusion 458 -1867 458 -1867 0 cellNo=757
rlabel pdiffusion 465 -1867 465 -1867 0 feedthrough
rlabel pdiffusion 472 -1867 472 -1867 0 feedthrough
rlabel pdiffusion 479 -1867 479 -1867 0 feedthrough
rlabel pdiffusion 486 -1867 486 -1867 0 feedthrough
rlabel pdiffusion 493 -1867 493 -1867 0 feedthrough
rlabel pdiffusion 500 -1867 500 -1867 0 feedthrough
rlabel pdiffusion 507 -1867 507 -1867 0 cellNo=687
rlabel pdiffusion 514 -1867 514 -1867 0 feedthrough
rlabel pdiffusion 521 -1867 521 -1867 0 cellNo=55
rlabel pdiffusion 528 -1867 528 -1867 0 cellNo=703
rlabel pdiffusion 535 -1867 535 -1867 0 feedthrough
rlabel pdiffusion 542 -1867 542 -1867 0 feedthrough
rlabel pdiffusion 549 -1867 549 -1867 0 cellNo=156
rlabel pdiffusion 556 -1867 556 -1867 0 feedthrough
rlabel pdiffusion 563 -1867 563 -1867 0 cellNo=511
rlabel pdiffusion 570 -1867 570 -1867 0 cellNo=151
rlabel pdiffusion 577 -1867 577 -1867 0 feedthrough
rlabel pdiffusion 584 -1867 584 -1867 0 feedthrough
rlabel pdiffusion 591 -1867 591 -1867 0 feedthrough
rlabel pdiffusion 598 -1867 598 -1867 0 feedthrough
rlabel pdiffusion 605 -1867 605 -1867 0 feedthrough
rlabel pdiffusion 612 -1867 612 -1867 0 feedthrough
rlabel pdiffusion 619 -1867 619 -1867 0 feedthrough
rlabel pdiffusion 626 -1867 626 -1867 0 cellNo=770
rlabel pdiffusion 633 -1867 633 -1867 0 cellNo=669
rlabel pdiffusion 640 -1867 640 -1867 0 cellNo=915
rlabel pdiffusion 647 -1867 647 -1867 0 feedthrough
rlabel pdiffusion 654 -1867 654 -1867 0 feedthrough
rlabel pdiffusion 661 -1867 661 -1867 0 cellNo=963
rlabel pdiffusion 668 -1867 668 -1867 0 feedthrough
rlabel pdiffusion 675 -1867 675 -1867 0 feedthrough
rlabel pdiffusion 682 -1867 682 -1867 0 feedthrough
rlabel pdiffusion 689 -1867 689 -1867 0 feedthrough
rlabel pdiffusion 696 -1867 696 -1867 0 feedthrough
rlabel pdiffusion 703 -1867 703 -1867 0 cellNo=975
rlabel pdiffusion 710 -1867 710 -1867 0 feedthrough
rlabel pdiffusion 717 -1867 717 -1867 0 feedthrough
rlabel pdiffusion 724 -1867 724 -1867 0 cellNo=774
rlabel pdiffusion 731 -1867 731 -1867 0 feedthrough
rlabel pdiffusion 738 -1867 738 -1867 0 feedthrough
rlabel pdiffusion 745 -1867 745 -1867 0 feedthrough
rlabel pdiffusion 752 -1867 752 -1867 0 feedthrough
rlabel pdiffusion 759 -1867 759 -1867 0 feedthrough
rlabel pdiffusion 766 -1867 766 -1867 0 feedthrough
rlabel pdiffusion 773 -1867 773 -1867 0 feedthrough
rlabel pdiffusion 780 -1867 780 -1867 0 feedthrough
rlabel pdiffusion 787 -1867 787 -1867 0 feedthrough
rlabel pdiffusion 794 -1867 794 -1867 0 feedthrough
rlabel pdiffusion 801 -1867 801 -1867 0 feedthrough
rlabel pdiffusion 808 -1867 808 -1867 0 feedthrough
rlabel pdiffusion 815 -1867 815 -1867 0 cellNo=763
rlabel pdiffusion 822 -1867 822 -1867 0 feedthrough
rlabel pdiffusion 829 -1867 829 -1867 0 feedthrough
rlabel pdiffusion 836 -1867 836 -1867 0 cellNo=391
rlabel pdiffusion 843 -1867 843 -1867 0 cellNo=477
rlabel pdiffusion 850 -1867 850 -1867 0 cellNo=515
rlabel pdiffusion 857 -1867 857 -1867 0 feedthrough
rlabel pdiffusion 864 -1867 864 -1867 0 feedthrough
rlabel pdiffusion 871 -1867 871 -1867 0 feedthrough
rlabel pdiffusion 878 -1867 878 -1867 0 feedthrough
rlabel pdiffusion 899 -1867 899 -1867 0 feedthrough
rlabel pdiffusion 913 -1867 913 -1867 0 cellNo=219
rlabel pdiffusion 948 -1867 948 -1867 0 cellNo=995
rlabel pdiffusion 17 -1938 17 -1938 0 feedthrough
rlabel pdiffusion 24 -1938 24 -1938 0 feedthrough
rlabel pdiffusion 31 -1938 31 -1938 0 cellNo=784
rlabel pdiffusion 38 -1938 38 -1938 0 cellNo=600
rlabel pdiffusion 45 -1938 45 -1938 0 cellNo=67
rlabel pdiffusion 52 -1938 52 -1938 0 feedthrough
rlabel pdiffusion 59 -1938 59 -1938 0 feedthrough
rlabel pdiffusion 66 -1938 66 -1938 0 feedthrough
rlabel pdiffusion 73 -1938 73 -1938 0 feedthrough
rlabel pdiffusion 80 -1938 80 -1938 0 feedthrough
rlabel pdiffusion 87 -1938 87 -1938 0 feedthrough
rlabel pdiffusion 94 -1938 94 -1938 0 feedthrough
rlabel pdiffusion 101 -1938 101 -1938 0 feedthrough
rlabel pdiffusion 108 -1938 108 -1938 0 feedthrough
rlabel pdiffusion 115 -1938 115 -1938 0 feedthrough
rlabel pdiffusion 122 -1938 122 -1938 0 cellNo=191
rlabel pdiffusion 129 -1938 129 -1938 0 feedthrough
rlabel pdiffusion 136 -1938 136 -1938 0 feedthrough
rlabel pdiffusion 143 -1938 143 -1938 0 cellNo=841
rlabel pdiffusion 150 -1938 150 -1938 0 feedthrough
rlabel pdiffusion 157 -1938 157 -1938 0 cellNo=648
rlabel pdiffusion 164 -1938 164 -1938 0 feedthrough
rlabel pdiffusion 171 -1938 171 -1938 0 feedthrough
rlabel pdiffusion 178 -1938 178 -1938 0 cellNo=504
rlabel pdiffusion 185 -1938 185 -1938 0 cellNo=896
rlabel pdiffusion 192 -1938 192 -1938 0 cellNo=634
rlabel pdiffusion 199 -1938 199 -1938 0 feedthrough
rlabel pdiffusion 206 -1938 206 -1938 0 feedthrough
rlabel pdiffusion 213 -1938 213 -1938 0 feedthrough
rlabel pdiffusion 220 -1938 220 -1938 0 cellNo=575
rlabel pdiffusion 227 -1938 227 -1938 0 cellNo=74
rlabel pdiffusion 234 -1938 234 -1938 0 cellNo=988
rlabel pdiffusion 241 -1938 241 -1938 0 cellNo=128
rlabel pdiffusion 248 -1938 248 -1938 0 feedthrough
rlabel pdiffusion 255 -1938 255 -1938 0 feedthrough
rlabel pdiffusion 262 -1938 262 -1938 0 feedthrough
rlabel pdiffusion 269 -1938 269 -1938 0 feedthrough
rlabel pdiffusion 276 -1938 276 -1938 0 feedthrough
rlabel pdiffusion 283 -1938 283 -1938 0 cellNo=254
rlabel pdiffusion 290 -1938 290 -1938 0 feedthrough
rlabel pdiffusion 297 -1938 297 -1938 0 feedthrough
rlabel pdiffusion 304 -1938 304 -1938 0 feedthrough
rlabel pdiffusion 311 -1938 311 -1938 0 feedthrough
rlabel pdiffusion 318 -1938 318 -1938 0 cellNo=465
rlabel pdiffusion 325 -1938 325 -1938 0 feedthrough
rlabel pdiffusion 332 -1938 332 -1938 0 cellNo=883
rlabel pdiffusion 339 -1938 339 -1938 0 feedthrough
rlabel pdiffusion 346 -1938 346 -1938 0 feedthrough
rlabel pdiffusion 353 -1938 353 -1938 0 feedthrough
rlabel pdiffusion 360 -1938 360 -1938 0 feedthrough
rlabel pdiffusion 367 -1938 367 -1938 0 feedthrough
rlabel pdiffusion 374 -1938 374 -1938 0 feedthrough
rlabel pdiffusion 381 -1938 381 -1938 0 feedthrough
rlabel pdiffusion 388 -1938 388 -1938 0 feedthrough
rlabel pdiffusion 395 -1938 395 -1938 0 cellNo=259
rlabel pdiffusion 402 -1938 402 -1938 0 feedthrough
rlabel pdiffusion 409 -1938 409 -1938 0 cellNo=619
rlabel pdiffusion 416 -1938 416 -1938 0 cellNo=379
rlabel pdiffusion 423 -1938 423 -1938 0 feedthrough
rlabel pdiffusion 430 -1938 430 -1938 0 feedthrough
rlabel pdiffusion 437 -1938 437 -1938 0 cellNo=183
rlabel pdiffusion 444 -1938 444 -1938 0 feedthrough
rlabel pdiffusion 451 -1938 451 -1938 0 cellNo=221
rlabel pdiffusion 458 -1938 458 -1938 0 cellNo=756
rlabel pdiffusion 465 -1938 465 -1938 0 feedthrough
rlabel pdiffusion 472 -1938 472 -1938 0 cellNo=520
rlabel pdiffusion 479 -1938 479 -1938 0 feedthrough
rlabel pdiffusion 486 -1938 486 -1938 0 feedthrough
rlabel pdiffusion 493 -1938 493 -1938 0 feedthrough
rlabel pdiffusion 500 -1938 500 -1938 0 cellNo=851
rlabel pdiffusion 507 -1938 507 -1938 0 feedthrough
rlabel pdiffusion 514 -1938 514 -1938 0 feedthrough
rlabel pdiffusion 521 -1938 521 -1938 0 feedthrough
rlabel pdiffusion 528 -1938 528 -1938 0 feedthrough
rlabel pdiffusion 535 -1938 535 -1938 0 feedthrough
rlabel pdiffusion 542 -1938 542 -1938 0 feedthrough
rlabel pdiffusion 549 -1938 549 -1938 0 feedthrough
rlabel pdiffusion 556 -1938 556 -1938 0 feedthrough
rlabel pdiffusion 563 -1938 563 -1938 0 feedthrough
rlabel pdiffusion 570 -1938 570 -1938 0 feedthrough
rlabel pdiffusion 577 -1938 577 -1938 0 cellNo=458
rlabel pdiffusion 584 -1938 584 -1938 0 feedthrough
rlabel pdiffusion 591 -1938 591 -1938 0 cellNo=926
rlabel pdiffusion 598 -1938 598 -1938 0 feedthrough
rlabel pdiffusion 605 -1938 605 -1938 0 cellNo=95
rlabel pdiffusion 612 -1938 612 -1938 0 feedthrough
rlabel pdiffusion 619 -1938 619 -1938 0 feedthrough
rlabel pdiffusion 626 -1938 626 -1938 0 feedthrough
rlabel pdiffusion 633 -1938 633 -1938 0 feedthrough
rlabel pdiffusion 640 -1938 640 -1938 0 feedthrough
rlabel pdiffusion 647 -1938 647 -1938 0 feedthrough
rlabel pdiffusion 654 -1938 654 -1938 0 feedthrough
rlabel pdiffusion 661 -1938 661 -1938 0 feedthrough
rlabel pdiffusion 668 -1938 668 -1938 0 feedthrough
rlabel pdiffusion 675 -1938 675 -1938 0 feedthrough
rlabel pdiffusion 682 -1938 682 -1938 0 cellNo=381
rlabel pdiffusion 689 -1938 689 -1938 0 feedthrough
rlabel pdiffusion 696 -1938 696 -1938 0 feedthrough
rlabel pdiffusion 703 -1938 703 -1938 0 feedthrough
rlabel pdiffusion 710 -1938 710 -1938 0 feedthrough
rlabel pdiffusion 717 -1938 717 -1938 0 feedthrough
rlabel pdiffusion 724 -1938 724 -1938 0 feedthrough
rlabel pdiffusion 731 -1938 731 -1938 0 feedthrough
rlabel pdiffusion 738 -1938 738 -1938 0 feedthrough
rlabel pdiffusion 745 -1938 745 -1938 0 feedthrough
rlabel pdiffusion 752 -1938 752 -1938 0 feedthrough
rlabel pdiffusion 759 -1938 759 -1938 0 cellNo=664
rlabel pdiffusion 766 -1938 766 -1938 0 feedthrough
rlabel pdiffusion 773 -1938 773 -1938 0 feedthrough
rlabel pdiffusion 780 -1938 780 -1938 0 cellNo=49
rlabel pdiffusion 787 -1938 787 -1938 0 feedthrough
rlabel pdiffusion 794 -1938 794 -1938 0 feedthrough
rlabel pdiffusion 815 -1938 815 -1938 0 feedthrough
rlabel pdiffusion 822 -1938 822 -1938 0 feedthrough
rlabel pdiffusion 38 -1997 38 -1997 0 feedthrough
rlabel pdiffusion 45 -1997 45 -1997 0 feedthrough
rlabel pdiffusion 52 -1997 52 -1997 0 feedthrough
rlabel pdiffusion 59 -1997 59 -1997 0 feedthrough
rlabel pdiffusion 66 -1997 66 -1997 0 feedthrough
rlabel pdiffusion 73 -1997 73 -1997 0 feedthrough
rlabel pdiffusion 80 -1997 80 -1997 0 feedthrough
rlabel pdiffusion 87 -1997 87 -1997 0 feedthrough
rlabel pdiffusion 94 -1997 94 -1997 0 feedthrough
rlabel pdiffusion 101 -1997 101 -1997 0 feedthrough
rlabel pdiffusion 108 -1997 108 -1997 0 feedthrough
rlabel pdiffusion 115 -1997 115 -1997 0 feedthrough
rlabel pdiffusion 122 -1997 122 -1997 0 feedthrough
rlabel pdiffusion 129 -1997 129 -1997 0 cellNo=331
rlabel pdiffusion 136 -1997 136 -1997 0 cellNo=916
rlabel pdiffusion 143 -1997 143 -1997 0 feedthrough
rlabel pdiffusion 150 -1997 150 -1997 0 cellNo=942
rlabel pdiffusion 157 -1997 157 -1997 0 cellNo=36
rlabel pdiffusion 164 -1997 164 -1997 0 feedthrough
rlabel pdiffusion 171 -1997 171 -1997 0 feedthrough
rlabel pdiffusion 178 -1997 178 -1997 0 feedthrough
rlabel pdiffusion 185 -1997 185 -1997 0 feedthrough
rlabel pdiffusion 192 -1997 192 -1997 0 feedthrough
rlabel pdiffusion 199 -1997 199 -1997 0 cellNo=1
rlabel pdiffusion 206 -1997 206 -1997 0 feedthrough
rlabel pdiffusion 213 -1997 213 -1997 0 feedthrough
rlabel pdiffusion 220 -1997 220 -1997 0 feedthrough
rlabel pdiffusion 227 -1997 227 -1997 0 cellNo=952
rlabel pdiffusion 234 -1997 234 -1997 0 feedthrough
rlabel pdiffusion 241 -1997 241 -1997 0 cellNo=767
rlabel pdiffusion 248 -1997 248 -1997 0 feedthrough
rlabel pdiffusion 255 -1997 255 -1997 0 feedthrough
rlabel pdiffusion 262 -1997 262 -1997 0 cellNo=429
rlabel pdiffusion 269 -1997 269 -1997 0 cellNo=421
rlabel pdiffusion 276 -1997 276 -1997 0 feedthrough
rlabel pdiffusion 283 -1997 283 -1997 0 feedthrough
rlabel pdiffusion 290 -1997 290 -1997 0 cellNo=19
rlabel pdiffusion 297 -1997 297 -1997 0 feedthrough
rlabel pdiffusion 304 -1997 304 -1997 0 feedthrough
rlabel pdiffusion 311 -1997 311 -1997 0 cellNo=203
rlabel pdiffusion 318 -1997 318 -1997 0 feedthrough
rlabel pdiffusion 325 -1997 325 -1997 0 feedthrough
rlabel pdiffusion 332 -1997 332 -1997 0 feedthrough
rlabel pdiffusion 339 -1997 339 -1997 0 feedthrough
rlabel pdiffusion 346 -1997 346 -1997 0 feedthrough
rlabel pdiffusion 353 -1997 353 -1997 0 feedthrough
rlabel pdiffusion 360 -1997 360 -1997 0 feedthrough
rlabel pdiffusion 367 -1997 367 -1997 0 cellNo=369
rlabel pdiffusion 374 -1997 374 -1997 0 feedthrough
rlabel pdiffusion 381 -1997 381 -1997 0 cellNo=651
rlabel pdiffusion 388 -1997 388 -1997 0 feedthrough
rlabel pdiffusion 395 -1997 395 -1997 0 feedthrough
rlabel pdiffusion 402 -1997 402 -1997 0 feedthrough
rlabel pdiffusion 409 -1997 409 -1997 0 feedthrough
rlabel pdiffusion 416 -1997 416 -1997 0 feedthrough
rlabel pdiffusion 423 -1997 423 -1997 0 feedthrough
rlabel pdiffusion 430 -1997 430 -1997 0 cellNo=202
rlabel pdiffusion 437 -1997 437 -1997 0 cellNo=64
rlabel pdiffusion 444 -1997 444 -1997 0 cellNo=776
rlabel pdiffusion 451 -1997 451 -1997 0 feedthrough
rlabel pdiffusion 458 -1997 458 -1997 0 feedthrough
rlabel pdiffusion 465 -1997 465 -1997 0 feedthrough
rlabel pdiffusion 472 -1997 472 -1997 0 feedthrough
rlabel pdiffusion 479 -1997 479 -1997 0 feedthrough
rlabel pdiffusion 486 -1997 486 -1997 0 feedthrough
rlabel pdiffusion 493 -1997 493 -1997 0 cellNo=266
rlabel pdiffusion 500 -1997 500 -1997 0 feedthrough
rlabel pdiffusion 507 -1997 507 -1997 0 feedthrough
rlabel pdiffusion 514 -1997 514 -1997 0 cellNo=217
rlabel pdiffusion 521 -1997 521 -1997 0 feedthrough
rlabel pdiffusion 528 -1997 528 -1997 0 feedthrough
rlabel pdiffusion 535 -1997 535 -1997 0 feedthrough
rlabel pdiffusion 542 -1997 542 -1997 0 feedthrough
rlabel pdiffusion 549 -1997 549 -1997 0 feedthrough
rlabel pdiffusion 556 -1997 556 -1997 0 feedthrough
rlabel pdiffusion 563 -1997 563 -1997 0 feedthrough
rlabel pdiffusion 570 -1997 570 -1997 0 feedthrough
rlabel pdiffusion 577 -1997 577 -1997 0 feedthrough
rlabel pdiffusion 584 -1997 584 -1997 0 cellNo=773
rlabel pdiffusion 591 -1997 591 -1997 0 cellNo=625
rlabel pdiffusion 598 -1997 598 -1997 0 cellNo=268
rlabel pdiffusion 605 -1997 605 -1997 0 feedthrough
rlabel pdiffusion 612 -1997 612 -1997 0 feedthrough
rlabel pdiffusion 619 -1997 619 -1997 0 feedthrough
rlabel pdiffusion 626 -1997 626 -1997 0 feedthrough
rlabel pdiffusion 633 -1997 633 -1997 0 feedthrough
rlabel pdiffusion 640 -1997 640 -1997 0 feedthrough
rlabel pdiffusion 647 -1997 647 -1997 0 feedthrough
rlabel pdiffusion 654 -1997 654 -1997 0 feedthrough
rlabel pdiffusion 661 -1997 661 -1997 0 cellNo=134
rlabel pdiffusion 668 -1997 668 -1997 0 feedthrough
rlabel pdiffusion 675 -1997 675 -1997 0 cellNo=348
rlabel pdiffusion 682 -1997 682 -1997 0 feedthrough
rlabel pdiffusion 689 -1997 689 -1997 0 cellNo=324
rlabel pdiffusion 696 -1997 696 -1997 0 feedthrough
rlabel pdiffusion 703 -1997 703 -1997 0 feedthrough
rlabel pdiffusion 710 -1997 710 -1997 0 feedthrough
rlabel pdiffusion 717 -1997 717 -1997 0 feedthrough
rlabel pdiffusion 724 -1997 724 -1997 0 cellNo=138
rlabel pdiffusion 731 -1997 731 -1997 0 feedthrough
rlabel pdiffusion 738 -1997 738 -1997 0 feedthrough
rlabel pdiffusion 745 -1997 745 -1997 0 cellNo=3
rlabel pdiffusion 752 -1997 752 -1997 0 feedthrough
rlabel pdiffusion 759 -1997 759 -1997 0 feedthrough
rlabel pdiffusion 766 -1997 766 -1997 0 feedthrough
rlabel pdiffusion 773 -1997 773 -1997 0 feedthrough
rlabel pdiffusion 780 -1997 780 -1997 0 cellNo=209
rlabel pdiffusion 787 -1997 787 -1997 0 feedthrough
rlabel pdiffusion 794 -1997 794 -1997 0 cellNo=412
rlabel pdiffusion 801 -1997 801 -1997 0 feedthrough
rlabel pdiffusion 808 -1997 808 -1997 0 feedthrough
rlabel pdiffusion 815 -1997 815 -1997 0 feedthrough
rlabel pdiffusion 17 -2060 17 -2060 0 feedthrough
rlabel pdiffusion 24 -2060 24 -2060 0 feedthrough
rlabel pdiffusion 31 -2060 31 -2060 0 feedthrough
rlabel pdiffusion 38 -2060 38 -2060 0 feedthrough
rlabel pdiffusion 45 -2060 45 -2060 0 feedthrough
rlabel pdiffusion 52 -2060 52 -2060 0 feedthrough
rlabel pdiffusion 59 -2060 59 -2060 0 feedthrough
rlabel pdiffusion 66 -2060 66 -2060 0 feedthrough
rlabel pdiffusion 73 -2060 73 -2060 0 feedthrough
rlabel pdiffusion 80 -2060 80 -2060 0 feedthrough
rlabel pdiffusion 87 -2060 87 -2060 0 feedthrough
rlabel pdiffusion 94 -2060 94 -2060 0 feedthrough
rlabel pdiffusion 101 -2060 101 -2060 0 feedthrough
rlabel pdiffusion 108 -2060 108 -2060 0 feedthrough
rlabel pdiffusion 115 -2060 115 -2060 0 feedthrough
rlabel pdiffusion 122 -2060 122 -2060 0 cellNo=698
rlabel pdiffusion 129 -2060 129 -2060 0 cellNo=394
rlabel pdiffusion 136 -2060 136 -2060 0 feedthrough
rlabel pdiffusion 143 -2060 143 -2060 0 cellNo=380
rlabel pdiffusion 150 -2060 150 -2060 0 feedthrough
rlabel pdiffusion 157 -2060 157 -2060 0 feedthrough
rlabel pdiffusion 164 -2060 164 -2060 0 cellNo=495
rlabel pdiffusion 171 -2060 171 -2060 0 feedthrough
rlabel pdiffusion 178 -2060 178 -2060 0 cellNo=283
rlabel pdiffusion 185 -2060 185 -2060 0 cellNo=404
rlabel pdiffusion 192 -2060 192 -2060 0 feedthrough
rlabel pdiffusion 199 -2060 199 -2060 0 feedthrough
rlabel pdiffusion 206 -2060 206 -2060 0 feedthrough
rlabel pdiffusion 213 -2060 213 -2060 0 feedthrough
rlabel pdiffusion 220 -2060 220 -2060 0 feedthrough
rlabel pdiffusion 227 -2060 227 -2060 0 cellNo=452
rlabel pdiffusion 234 -2060 234 -2060 0 cellNo=981
rlabel pdiffusion 241 -2060 241 -2060 0 cellNo=874
rlabel pdiffusion 248 -2060 248 -2060 0 feedthrough
rlabel pdiffusion 255 -2060 255 -2060 0 cellNo=426
rlabel pdiffusion 262 -2060 262 -2060 0 feedthrough
rlabel pdiffusion 269 -2060 269 -2060 0 feedthrough
rlabel pdiffusion 276 -2060 276 -2060 0 feedthrough
rlabel pdiffusion 283 -2060 283 -2060 0 feedthrough
rlabel pdiffusion 290 -2060 290 -2060 0 feedthrough
rlabel pdiffusion 297 -2060 297 -2060 0 feedthrough
rlabel pdiffusion 304 -2060 304 -2060 0 feedthrough
rlabel pdiffusion 311 -2060 311 -2060 0 feedthrough
rlabel pdiffusion 318 -2060 318 -2060 0 feedthrough
rlabel pdiffusion 325 -2060 325 -2060 0 feedthrough
rlabel pdiffusion 332 -2060 332 -2060 0 feedthrough
rlabel pdiffusion 339 -2060 339 -2060 0 feedthrough
rlabel pdiffusion 346 -2060 346 -2060 0 cellNo=468
rlabel pdiffusion 353 -2060 353 -2060 0 cellNo=196
rlabel pdiffusion 360 -2060 360 -2060 0 feedthrough
rlabel pdiffusion 367 -2060 367 -2060 0 feedthrough
rlabel pdiffusion 374 -2060 374 -2060 0 feedthrough
rlabel pdiffusion 381 -2060 381 -2060 0 feedthrough
rlabel pdiffusion 388 -2060 388 -2060 0 feedthrough
rlabel pdiffusion 395 -2060 395 -2060 0 cellNo=434
rlabel pdiffusion 402 -2060 402 -2060 0 cellNo=522
rlabel pdiffusion 409 -2060 409 -2060 0 feedthrough
rlabel pdiffusion 416 -2060 416 -2060 0 cellNo=549
rlabel pdiffusion 423 -2060 423 -2060 0 feedthrough
rlabel pdiffusion 430 -2060 430 -2060 0 cellNo=25
rlabel pdiffusion 437 -2060 437 -2060 0 feedthrough
rlabel pdiffusion 444 -2060 444 -2060 0 feedthrough
rlabel pdiffusion 451 -2060 451 -2060 0 feedthrough
rlabel pdiffusion 458 -2060 458 -2060 0 cellNo=786
rlabel pdiffusion 465 -2060 465 -2060 0 feedthrough
rlabel pdiffusion 472 -2060 472 -2060 0 cellNo=814
rlabel pdiffusion 479 -2060 479 -2060 0 cellNo=335
rlabel pdiffusion 486 -2060 486 -2060 0 cellNo=927
rlabel pdiffusion 493 -2060 493 -2060 0 feedthrough
rlabel pdiffusion 500 -2060 500 -2060 0 feedthrough
rlabel pdiffusion 507 -2060 507 -2060 0 cellNo=808
rlabel pdiffusion 514 -2060 514 -2060 0 cellNo=577
rlabel pdiffusion 521 -2060 521 -2060 0 feedthrough
rlabel pdiffusion 528 -2060 528 -2060 0 feedthrough
rlabel pdiffusion 535 -2060 535 -2060 0 feedthrough
rlabel pdiffusion 542 -2060 542 -2060 0 feedthrough
rlabel pdiffusion 549 -2060 549 -2060 0 feedthrough
rlabel pdiffusion 556 -2060 556 -2060 0 feedthrough
rlabel pdiffusion 563 -2060 563 -2060 0 cellNo=359
rlabel pdiffusion 570 -2060 570 -2060 0 cellNo=797
rlabel pdiffusion 577 -2060 577 -2060 0 feedthrough
rlabel pdiffusion 584 -2060 584 -2060 0 feedthrough
rlabel pdiffusion 591 -2060 591 -2060 0 feedthrough
rlabel pdiffusion 598 -2060 598 -2060 0 feedthrough
rlabel pdiffusion 605 -2060 605 -2060 0 feedthrough
rlabel pdiffusion 612 -2060 612 -2060 0 feedthrough
rlabel pdiffusion 619 -2060 619 -2060 0 feedthrough
rlabel pdiffusion 626 -2060 626 -2060 0 feedthrough
rlabel pdiffusion 633 -2060 633 -2060 0 feedthrough
rlabel pdiffusion 640 -2060 640 -2060 0 feedthrough
rlabel pdiffusion 647 -2060 647 -2060 0 feedthrough
rlabel pdiffusion 654 -2060 654 -2060 0 cellNo=437
rlabel pdiffusion 661 -2060 661 -2060 0 feedthrough
rlabel pdiffusion 668 -2060 668 -2060 0 cellNo=587
rlabel pdiffusion 675 -2060 675 -2060 0 feedthrough
rlabel pdiffusion 682 -2060 682 -2060 0 feedthrough
rlabel pdiffusion 689 -2060 689 -2060 0 feedthrough
rlabel pdiffusion 696 -2060 696 -2060 0 feedthrough
rlabel pdiffusion 703 -2060 703 -2060 0 feedthrough
rlabel pdiffusion 710 -2060 710 -2060 0 feedthrough
rlabel pdiffusion 717 -2060 717 -2060 0 feedthrough
rlabel pdiffusion 724 -2060 724 -2060 0 cellNo=817
rlabel pdiffusion 731 -2060 731 -2060 0 feedthrough
rlabel pdiffusion 738 -2060 738 -2060 0 feedthrough
rlabel pdiffusion 745 -2060 745 -2060 0 feedthrough
rlabel pdiffusion 752 -2060 752 -2060 0 feedthrough
rlabel pdiffusion 759 -2060 759 -2060 0 feedthrough
rlabel pdiffusion 766 -2060 766 -2060 0 feedthrough
rlabel pdiffusion 773 -2060 773 -2060 0 feedthrough
rlabel pdiffusion 780 -2060 780 -2060 0 feedthrough
rlabel pdiffusion 787 -2060 787 -2060 0 feedthrough
rlabel pdiffusion 17 -2125 17 -2125 0 feedthrough
rlabel pdiffusion 24 -2125 24 -2125 0 feedthrough
rlabel pdiffusion 31 -2125 31 -2125 0 feedthrough
rlabel pdiffusion 38 -2125 38 -2125 0 cellNo=996
rlabel pdiffusion 45 -2125 45 -2125 0 feedthrough
rlabel pdiffusion 52 -2125 52 -2125 0 feedthrough
rlabel pdiffusion 59 -2125 59 -2125 0 feedthrough
rlabel pdiffusion 66 -2125 66 -2125 0 feedthrough
rlabel pdiffusion 73 -2125 73 -2125 0 feedthrough
rlabel pdiffusion 80 -2125 80 -2125 0 feedthrough
rlabel pdiffusion 87 -2125 87 -2125 0 feedthrough
rlabel pdiffusion 94 -2125 94 -2125 0 cellNo=736
rlabel pdiffusion 101 -2125 101 -2125 0 cellNo=857
rlabel pdiffusion 108 -2125 108 -2125 0 feedthrough
rlabel pdiffusion 115 -2125 115 -2125 0 feedthrough
rlabel pdiffusion 122 -2125 122 -2125 0 feedthrough
rlabel pdiffusion 129 -2125 129 -2125 0 cellNo=626
rlabel pdiffusion 136 -2125 136 -2125 0 cellNo=463
rlabel pdiffusion 143 -2125 143 -2125 0 feedthrough
rlabel pdiffusion 150 -2125 150 -2125 0 feedthrough
rlabel pdiffusion 157 -2125 157 -2125 0 cellNo=210
rlabel pdiffusion 164 -2125 164 -2125 0 feedthrough
rlabel pdiffusion 171 -2125 171 -2125 0 cellNo=682
rlabel pdiffusion 178 -2125 178 -2125 0 cellNo=63
rlabel pdiffusion 185 -2125 185 -2125 0 cellNo=992
rlabel pdiffusion 192 -2125 192 -2125 0 feedthrough
rlabel pdiffusion 199 -2125 199 -2125 0 cellNo=947
rlabel pdiffusion 206 -2125 206 -2125 0 cellNo=267
rlabel pdiffusion 213 -2125 213 -2125 0 feedthrough
rlabel pdiffusion 220 -2125 220 -2125 0 cellNo=741
rlabel pdiffusion 227 -2125 227 -2125 0 cellNo=438
rlabel pdiffusion 234 -2125 234 -2125 0 feedthrough
rlabel pdiffusion 241 -2125 241 -2125 0 feedthrough
rlabel pdiffusion 248 -2125 248 -2125 0 cellNo=35
rlabel pdiffusion 255 -2125 255 -2125 0 feedthrough
rlabel pdiffusion 262 -2125 262 -2125 0 feedthrough
rlabel pdiffusion 269 -2125 269 -2125 0 feedthrough
rlabel pdiffusion 276 -2125 276 -2125 0 feedthrough
rlabel pdiffusion 283 -2125 283 -2125 0 feedthrough
rlabel pdiffusion 290 -2125 290 -2125 0 cellNo=761
rlabel pdiffusion 297 -2125 297 -2125 0 feedthrough
rlabel pdiffusion 304 -2125 304 -2125 0 feedthrough
rlabel pdiffusion 311 -2125 311 -2125 0 feedthrough
rlabel pdiffusion 318 -2125 318 -2125 0 cellNo=743
rlabel pdiffusion 325 -2125 325 -2125 0 feedthrough
rlabel pdiffusion 332 -2125 332 -2125 0 feedthrough
rlabel pdiffusion 339 -2125 339 -2125 0 feedthrough
rlabel pdiffusion 346 -2125 346 -2125 0 cellNo=561
rlabel pdiffusion 353 -2125 353 -2125 0 feedthrough
rlabel pdiffusion 360 -2125 360 -2125 0 cellNo=585
rlabel pdiffusion 367 -2125 367 -2125 0 feedthrough
rlabel pdiffusion 374 -2125 374 -2125 0 feedthrough
rlabel pdiffusion 381 -2125 381 -2125 0 cellNo=82
rlabel pdiffusion 388 -2125 388 -2125 0 feedthrough
rlabel pdiffusion 395 -2125 395 -2125 0 feedthrough
rlabel pdiffusion 402 -2125 402 -2125 0 feedthrough
rlabel pdiffusion 409 -2125 409 -2125 0 cellNo=657
rlabel pdiffusion 416 -2125 416 -2125 0 feedthrough
rlabel pdiffusion 423 -2125 423 -2125 0 feedthrough
rlabel pdiffusion 430 -2125 430 -2125 0 feedthrough
rlabel pdiffusion 437 -2125 437 -2125 0 cellNo=166
rlabel pdiffusion 444 -2125 444 -2125 0 feedthrough
rlabel pdiffusion 451 -2125 451 -2125 0 feedthrough
rlabel pdiffusion 458 -2125 458 -2125 0 cellNo=174
rlabel pdiffusion 465 -2125 465 -2125 0 cellNo=476
rlabel pdiffusion 472 -2125 472 -2125 0 cellNo=319
rlabel pdiffusion 479 -2125 479 -2125 0 feedthrough
rlabel pdiffusion 486 -2125 486 -2125 0 feedthrough
rlabel pdiffusion 493 -2125 493 -2125 0 feedthrough
rlabel pdiffusion 500 -2125 500 -2125 0 feedthrough
rlabel pdiffusion 507 -2125 507 -2125 0 cellNo=890
rlabel pdiffusion 514 -2125 514 -2125 0 feedthrough
rlabel pdiffusion 521 -2125 521 -2125 0 feedthrough
rlabel pdiffusion 528 -2125 528 -2125 0 feedthrough
rlabel pdiffusion 535 -2125 535 -2125 0 feedthrough
rlabel pdiffusion 542 -2125 542 -2125 0 feedthrough
rlabel pdiffusion 549 -2125 549 -2125 0 feedthrough
rlabel pdiffusion 556 -2125 556 -2125 0 feedthrough
rlabel pdiffusion 563 -2125 563 -2125 0 feedthrough
rlabel pdiffusion 570 -2125 570 -2125 0 feedthrough
rlabel pdiffusion 577 -2125 577 -2125 0 feedthrough
rlabel pdiffusion 584 -2125 584 -2125 0 feedthrough
rlabel pdiffusion 591 -2125 591 -2125 0 cellNo=959
rlabel pdiffusion 598 -2125 598 -2125 0 feedthrough
rlabel pdiffusion 605 -2125 605 -2125 0 feedthrough
rlabel pdiffusion 612 -2125 612 -2125 0 feedthrough
rlabel pdiffusion 619 -2125 619 -2125 0 feedthrough
rlabel pdiffusion 626 -2125 626 -2125 0 feedthrough
rlabel pdiffusion 633 -2125 633 -2125 0 feedthrough
rlabel pdiffusion 640 -2125 640 -2125 0 feedthrough
rlabel pdiffusion 647 -2125 647 -2125 0 feedthrough
rlabel pdiffusion 654 -2125 654 -2125 0 feedthrough
rlabel pdiffusion 661 -2125 661 -2125 0 feedthrough
rlabel pdiffusion 668 -2125 668 -2125 0 feedthrough
rlabel pdiffusion 675 -2125 675 -2125 0 feedthrough
rlabel pdiffusion 682 -2125 682 -2125 0 feedthrough
rlabel pdiffusion 689 -2125 689 -2125 0 feedthrough
rlabel pdiffusion 696 -2125 696 -2125 0 feedthrough
rlabel pdiffusion 703 -2125 703 -2125 0 feedthrough
rlabel pdiffusion 710 -2125 710 -2125 0 feedthrough
rlabel pdiffusion 717 -2125 717 -2125 0 feedthrough
rlabel pdiffusion 724 -2125 724 -2125 0 feedthrough
rlabel pdiffusion 731 -2125 731 -2125 0 cellNo=423
rlabel pdiffusion 738 -2125 738 -2125 0 feedthrough
rlabel pdiffusion 87 -2176 87 -2176 0 feedthrough
rlabel pdiffusion 101 -2176 101 -2176 0 feedthrough
rlabel pdiffusion 108 -2176 108 -2176 0 feedthrough
rlabel pdiffusion 115 -2176 115 -2176 0 feedthrough
rlabel pdiffusion 122 -2176 122 -2176 0 feedthrough
rlabel pdiffusion 129 -2176 129 -2176 0 cellNo=58
rlabel pdiffusion 136 -2176 136 -2176 0 cellNo=256
rlabel pdiffusion 143 -2176 143 -2176 0 feedthrough
rlabel pdiffusion 150 -2176 150 -2176 0 cellNo=955
rlabel pdiffusion 157 -2176 157 -2176 0 cellNo=236
rlabel pdiffusion 164 -2176 164 -2176 0 feedthrough
rlabel pdiffusion 171 -2176 171 -2176 0 feedthrough
rlabel pdiffusion 178 -2176 178 -2176 0 feedthrough
rlabel pdiffusion 185 -2176 185 -2176 0 feedthrough
rlabel pdiffusion 192 -2176 192 -2176 0 feedthrough
rlabel pdiffusion 199 -2176 199 -2176 0 feedthrough
rlabel pdiffusion 206 -2176 206 -2176 0 feedthrough
rlabel pdiffusion 213 -2176 213 -2176 0 cellNo=173
rlabel pdiffusion 220 -2176 220 -2176 0 cellNo=482
rlabel pdiffusion 227 -2176 227 -2176 0 cellNo=716
rlabel pdiffusion 234 -2176 234 -2176 0 feedthrough
rlabel pdiffusion 241 -2176 241 -2176 0 cellNo=1000
rlabel pdiffusion 248 -2176 248 -2176 0 feedthrough
rlabel pdiffusion 255 -2176 255 -2176 0 feedthrough
rlabel pdiffusion 262 -2176 262 -2176 0 feedthrough
rlabel pdiffusion 269 -2176 269 -2176 0 feedthrough
rlabel pdiffusion 276 -2176 276 -2176 0 feedthrough
rlabel pdiffusion 283 -2176 283 -2176 0 cellNo=555
rlabel pdiffusion 290 -2176 290 -2176 0 feedthrough
rlabel pdiffusion 297 -2176 297 -2176 0 cellNo=712
rlabel pdiffusion 304 -2176 304 -2176 0 feedthrough
rlabel pdiffusion 311 -2176 311 -2176 0 cellNo=849
rlabel pdiffusion 318 -2176 318 -2176 0 feedthrough
rlabel pdiffusion 325 -2176 325 -2176 0 feedthrough
rlabel pdiffusion 332 -2176 332 -2176 0 cellNo=903
rlabel pdiffusion 339 -2176 339 -2176 0 feedthrough
rlabel pdiffusion 346 -2176 346 -2176 0 feedthrough
rlabel pdiffusion 353 -2176 353 -2176 0 feedthrough
rlabel pdiffusion 360 -2176 360 -2176 0 feedthrough
rlabel pdiffusion 367 -2176 367 -2176 0 feedthrough
rlabel pdiffusion 374 -2176 374 -2176 0 feedthrough
rlabel pdiffusion 381 -2176 381 -2176 0 feedthrough
rlabel pdiffusion 388 -2176 388 -2176 0 cellNo=20
rlabel pdiffusion 395 -2176 395 -2176 0 feedthrough
rlabel pdiffusion 402 -2176 402 -2176 0 feedthrough
rlabel pdiffusion 409 -2176 409 -2176 0 cellNo=475
rlabel pdiffusion 416 -2176 416 -2176 0 feedthrough
rlabel pdiffusion 423 -2176 423 -2176 0 feedthrough
rlabel pdiffusion 430 -2176 430 -2176 0 cellNo=425
rlabel pdiffusion 437 -2176 437 -2176 0 feedthrough
rlabel pdiffusion 444 -2176 444 -2176 0 feedthrough
rlabel pdiffusion 451 -2176 451 -2176 0 cellNo=800
rlabel pdiffusion 458 -2176 458 -2176 0 cellNo=629
rlabel pdiffusion 465 -2176 465 -2176 0 feedthrough
rlabel pdiffusion 472 -2176 472 -2176 0 feedthrough
rlabel pdiffusion 479 -2176 479 -2176 0 feedthrough
rlabel pdiffusion 486 -2176 486 -2176 0 feedthrough
rlabel pdiffusion 493 -2176 493 -2176 0 cellNo=897
rlabel pdiffusion 500 -2176 500 -2176 0 feedthrough
rlabel pdiffusion 507 -2176 507 -2176 0 cellNo=281
rlabel pdiffusion 514 -2176 514 -2176 0 feedthrough
rlabel pdiffusion 521 -2176 521 -2176 0 feedthrough
rlabel pdiffusion 528 -2176 528 -2176 0 feedthrough
rlabel pdiffusion 535 -2176 535 -2176 0 feedthrough
rlabel pdiffusion 542 -2176 542 -2176 0 feedthrough
rlabel pdiffusion 549 -2176 549 -2176 0 feedthrough
rlabel pdiffusion 556 -2176 556 -2176 0 cellNo=796
rlabel pdiffusion 563 -2176 563 -2176 0 feedthrough
rlabel pdiffusion 570 -2176 570 -2176 0 cellNo=365
rlabel pdiffusion 577 -2176 577 -2176 0 cellNo=918
rlabel pdiffusion 584 -2176 584 -2176 0 cellNo=775
rlabel pdiffusion 591 -2176 591 -2176 0 feedthrough
rlabel pdiffusion 598 -2176 598 -2176 0 feedthrough
rlabel pdiffusion 605 -2176 605 -2176 0 feedthrough
rlabel pdiffusion 612 -2176 612 -2176 0 feedthrough
rlabel pdiffusion 619 -2176 619 -2176 0 feedthrough
rlabel pdiffusion 626 -2176 626 -2176 0 feedthrough
rlabel pdiffusion 633 -2176 633 -2176 0 feedthrough
rlabel pdiffusion 640 -2176 640 -2176 0 feedthrough
rlabel pdiffusion 647 -2176 647 -2176 0 feedthrough
rlabel pdiffusion 654 -2176 654 -2176 0 feedthrough
rlabel pdiffusion 661 -2176 661 -2176 0 feedthrough
rlabel pdiffusion 668 -2176 668 -2176 0 cellNo=938
rlabel pdiffusion 675 -2176 675 -2176 0 feedthrough
rlabel pdiffusion 682 -2176 682 -2176 0 cellNo=528
rlabel pdiffusion 689 -2176 689 -2176 0 feedthrough
rlabel pdiffusion 696 -2176 696 -2176 0 cellNo=865
rlabel pdiffusion 703 -2176 703 -2176 0 feedthrough
rlabel pdiffusion 710 -2176 710 -2176 0 feedthrough
rlabel pdiffusion 717 -2176 717 -2176 0 feedthrough
rlabel pdiffusion 724 -2176 724 -2176 0 feedthrough
rlabel pdiffusion 87 -2229 87 -2229 0 cellNo=361
rlabel pdiffusion 108 -2229 108 -2229 0 feedthrough
rlabel pdiffusion 115 -2229 115 -2229 0 feedthrough
rlabel pdiffusion 122 -2229 122 -2229 0 cellNo=969
rlabel pdiffusion 129 -2229 129 -2229 0 cellNo=732
rlabel pdiffusion 136 -2229 136 -2229 0 cellNo=110
rlabel pdiffusion 143 -2229 143 -2229 0 feedthrough
rlabel pdiffusion 150 -2229 150 -2229 0 feedthrough
rlabel pdiffusion 157 -2229 157 -2229 0 feedthrough
rlabel pdiffusion 164 -2229 164 -2229 0 cellNo=444
rlabel pdiffusion 171 -2229 171 -2229 0 cellNo=454
rlabel pdiffusion 178 -2229 178 -2229 0 cellNo=919
rlabel pdiffusion 185 -2229 185 -2229 0 feedthrough
rlabel pdiffusion 192 -2229 192 -2229 0 feedthrough
rlabel pdiffusion 199 -2229 199 -2229 0 cellNo=846
rlabel pdiffusion 206 -2229 206 -2229 0 cellNo=297
rlabel pdiffusion 213 -2229 213 -2229 0 feedthrough
rlabel pdiffusion 220 -2229 220 -2229 0 feedthrough
rlabel pdiffusion 227 -2229 227 -2229 0 cellNo=588
rlabel pdiffusion 234 -2229 234 -2229 0 feedthrough
rlabel pdiffusion 241 -2229 241 -2229 0 feedthrough
rlabel pdiffusion 248 -2229 248 -2229 0 feedthrough
rlabel pdiffusion 255 -2229 255 -2229 0 feedthrough
rlabel pdiffusion 262 -2229 262 -2229 0 feedthrough
rlabel pdiffusion 269 -2229 269 -2229 0 feedthrough
rlabel pdiffusion 276 -2229 276 -2229 0 feedthrough
rlabel pdiffusion 283 -2229 283 -2229 0 cellNo=893
rlabel pdiffusion 290 -2229 290 -2229 0 feedthrough
rlabel pdiffusion 297 -2229 297 -2229 0 feedthrough
rlabel pdiffusion 304 -2229 304 -2229 0 cellNo=889
rlabel pdiffusion 311 -2229 311 -2229 0 feedthrough
rlabel pdiffusion 318 -2229 318 -2229 0 feedthrough
rlabel pdiffusion 325 -2229 325 -2229 0 feedthrough
rlabel pdiffusion 332 -2229 332 -2229 0 feedthrough
rlabel pdiffusion 339 -2229 339 -2229 0 feedthrough
rlabel pdiffusion 346 -2229 346 -2229 0 feedthrough
rlabel pdiffusion 353 -2229 353 -2229 0 feedthrough
rlabel pdiffusion 360 -2229 360 -2229 0 cellNo=691
rlabel pdiffusion 367 -2229 367 -2229 0 feedthrough
rlabel pdiffusion 374 -2229 374 -2229 0 cellNo=902
rlabel pdiffusion 381 -2229 381 -2229 0 feedthrough
rlabel pdiffusion 388 -2229 388 -2229 0 cellNo=960
rlabel pdiffusion 395 -2229 395 -2229 0 feedthrough
rlabel pdiffusion 402 -2229 402 -2229 0 feedthrough
rlabel pdiffusion 409 -2229 409 -2229 0 feedthrough
rlabel pdiffusion 416 -2229 416 -2229 0 feedthrough
rlabel pdiffusion 423 -2229 423 -2229 0 cellNo=670
rlabel pdiffusion 430 -2229 430 -2229 0 feedthrough
rlabel pdiffusion 437 -2229 437 -2229 0 feedthrough
rlabel pdiffusion 444 -2229 444 -2229 0 cellNo=772
rlabel pdiffusion 451 -2229 451 -2229 0 feedthrough
rlabel pdiffusion 458 -2229 458 -2229 0 feedthrough
rlabel pdiffusion 465 -2229 465 -2229 0 cellNo=96
rlabel pdiffusion 472 -2229 472 -2229 0 feedthrough
rlabel pdiffusion 479 -2229 479 -2229 0 feedthrough
rlabel pdiffusion 486 -2229 486 -2229 0 feedthrough
rlabel pdiffusion 493 -2229 493 -2229 0 feedthrough
rlabel pdiffusion 500 -2229 500 -2229 0 feedthrough
rlabel pdiffusion 507 -2229 507 -2229 0 feedthrough
rlabel pdiffusion 514 -2229 514 -2229 0 feedthrough
rlabel pdiffusion 521 -2229 521 -2229 0 feedthrough
rlabel pdiffusion 528 -2229 528 -2229 0 feedthrough
rlabel pdiffusion 535 -2229 535 -2229 0 feedthrough
rlabel pdiffusion 542 -2229 542 -2229 0 feedthrough
rlabel pdiffusion 549 -2229 549 -2229 0 feedthrough
rlabel pdiffusion 556 -2229 556 -2229 0 feedthrough
rlabel pdiffusion 563 -2229 563 -2229 0 cellNo=649
rlabel pdiffusion 570 -2229 570 -2229 0 feedthrough
rlabel pdiffusion 577 -2229 577 -2229 0 cellNo=34
rlabel pdiffusion 584 -2229 584 -2229 0 feedthrough
rlabel pdiffusion 591 -2229 591 -2229 0 feedthrough
rlabel pdiffusion 598 -2229 598 -2229 0 feedthrough
rlabel pdiffusion 605 -2229 605 -2229 0 cellNo=908
rlabel pdiffusion 612 -2229 612 -2229 0 cellNo=749
rlabel pdiffusion 619 -2229 619 -2229 0 cellNo=500
rlabel pdiffusion 626 -2229 626 -2229 0 cellNo=242
rlabel pdiffusion 633 -2229 633 -2229 0 feedthrough
rlabel pdiffusion 640 -2229 640 -2229 0 feedthrough
rlabel pdiffusion 661 -2229 661 -2229 0 feedthrough
rlabel pdiffusion 115 -2266 115 -2266 0 feedthrough
rlabel pdiffusion 122 -2266 122 -2266 0 cellNo=921
rlabel pdiffusion 129 -2266 129 -2266 0 cellNo=936
rlabel pdiffusion 136 -2266 136 -2266 0 feedthrough
rlabel pdiffusion 143 -2266 143 -2266 0 cellNo=920
rlabel pdiffusion 150 -2266 150 -2266 0 cellNo=309
rlabel pdiffusion 157 -2266 157 -2266 0 feedthrough
rlabel pdiffusion 164 -2266 164 -2266 0 feedthrough
rlabel pdiffusion 171 -2266 171 -2266 0 feedthrough
rlabel pdiffusion 178 -2266 178 -2266 0 feedthrough
rlabel pdiffusion 185 -2266 185 -2266 0 feedthrough
rlabel pdiffusion 192 -2266 192 -2266 0 cellNo=950
rlabel pdiffusion 199 -2266 199 -2266 0 feedthrough
rlabel pdiffusion 206 -2266 206 -2266 0 feedthrough
rlabel pdiffusion 213 -2266 213 -2266 0 cellNo=48
rlabel pdiffusion 220 -2266 220 -2266 0 feedthrough
rlabel pdiffusion 227 -2266 227 -2266 0 feedthrough
rlabel pdiffusion 234 -2266 234 -2266 0 cellNo=383
rlabel pdiffusion 241 -2266 241 -2266 0 cellNo=455
rlabel pdiffusion 248 -2266 248 -2266 0 feedthrough
rlabel pdiffusion 255 -2266 255 -2266 0 feedthrough
rlabel pdiffusion 262 -2266 262 -2266 0 feedthrough
rlabel pdiffusion 269 -2266 269 -2266 0 feedthrough
rlabel pdiffusion 276 -2266 276 -2266 0 feedthrough
rlabel pdiffusion 283 -2266 283 -2266 0 cellNo=731
rlabel pdiffusion 290 -2266 290 -2266 0 feedthrough
rlabel pdiffusion 297 -2266 297 -2266 0 feedthrough
rlabel pdiffusion 304 -2266 304 -2266 0 cellNo=413
rlabel pdiffusion 311 -2266 311 -2266 0 cellNo=109
rlabel pdiffusion 318 -2266 318 -2266 0 feedthrough
rlabel pdiffusion 325 -2266 325 -2266 0 cellNo=932
rlabel pdiffusion 332 -2266 332 -2266 0 feedthrough
rlabel pdiffusion 339 -2266 339 -2266 0 feedthrough
rlabel pdiffusion 346 -2266 346 -2266 0 feedthrough
rlabel pdiffusion 353 -2266 353 -2266 0 feedthrough
rlabel pdiffusion 360 -2266 360 -2266 0 cellNo=822
rlabel pdiffusion 367 -2266 367 -2266 0 feedthrough
rlabel pdiffusion 374 -2266 374 -2266 0 cellNo=744
rlabel pdiffusion 381 -2266 381 -2266 0 feedthrough
rlabel pdiffusion 388 -2266 388 -2266 0 cellNo=801
rlabel pdiffusion 395 -2266 395 -2266 0 cellNo=611
rlabel pdiffusion 402 -2266 402 -2266 0 feedthrough
rlabel pdiffusion 409 -2266 409 -2266 0 cellNo=888
rlabel pdiffusion 416 -2266 416 -2266 0 feedthrough
rlabel pdiffusion 423 -2266 423 -2266 0 feedthrough
rlabel pdiffusion 430 -2266 430 -2266 0 cellNo=552
rlabel pdiffusion 437 -2266 437 -2266 0 feedthrough
rlabel pdiffusion 444 -2266 444 -2266 0 feedthrough
rlabel pdiffusion 451 -2266 451 -2266 0 feedthrough
rlabel pdiffusion 458 -2266 458 -2266 0 feedthrough
rlabel pdiffusion 465 -2266 465 -2266 0 feedthrough
rlabel pdiffusion 472 -2266 472 -2266 0 cellNo=692
rlabel pdiffusion 479 -2266 479 -2266 0 feedthrough
rlabel pdiffusion 486 -2266 486 -2266 0 feedthrough
rlabel pdiffusion 493 -2266 493 -2266 0 feedthrough
rlabel pdiffusion 500 -2266 500 -2266 0 feedthrough
rlabel pdiffusion 507 -2266 507 -2266 0 feedthrough
rlabel pdiffusion 514 -2266 514 -2266 0 feedthrough
rlabel pdiffusion 521 -2266 521 -2266 0 feedthrough
rlabel pdiffusion 528 -2266 528 -2266 0 feedthrough
rlabel pdiffusion 535 -2266 535 -2266 0 feedthrough
rlabel pdiffusion 542 -2266 542 -2266 0 feedthrough
rlabel pdiffusion 549 -2266 549 -2266 0 feedthrough
rlabel pdiffusion 556 -2266 556 -2266 0 feedthrough
rlabel pdiffusion 563 -2266 563 -2266 0 cellNo=967
rlabel pdiffusion 570 -2266 570 -2266 0 cellNo=408
rlabel pdiffusion 577 -2266 577 -2266 0 feedthrough
rlabel pdiffusion 584 -2266 584 -2266 0 feedthrough
rlabel pdiffusion 640 -2266 640 -2266 0 feedthrough
rlabel pdiffusion 122 -2293 122 -2293 0 cellNo=322
rlabel pdiffusion 178 -2293 178 -2293 0 feedthrough
rlabel pdiffusion 213 -2293 213 -2293 0 feedthrough
rlabel pdiffusion 220 -2293 220 -2293 0 cellNo=329
rlabel pdiffusion 227 -2293 227 -2293 0 feedthrough
rlabel pdiffusion 234 -2293 234 -2293 0 feedthrough
rlabel pdiffusion 241 -2293 241 -2293 0 cellNo=530
rlabel pdiffusion 248 -2293 248 -2293 0 cellNo=922
rlabel pdiffusion 255 -2293 255 -2293 0 feedthrough
rlabel pdiffusion 269 -2293 269 -2293 0 feedthrough
rlabel pdiffusion 276 -2293 276 -2293 0 feedthrough
rlabel pdiffusion 283 -2293 283 -2293 0 feedthrough
rlabel pdiffusion 290 -2293 290 -2293 0 cellNo=816
rlabel pdiffusion 297 -2293 297 -2293 0 feedthrough
rlabel pdiffusion 304 -2293 304 -2293 0 cellNo=944
rlabel pdiffusion 311 -2293 311 -2293 0 feedthrough
rlabel pdiffusion 318 -2293 318 -2293 0 feedthrough
rlabel pdiffusion 325 -2293 325 -2293 0 cellNo=488
rlabel pdiffusion 332 -2293 332 -2293 0 feedthrough
rlabel pdiffusion 339 -2293 339 -2293 0 cellNo=367
rlabel pdiffusion 346 -2293 346 -2293 0 feedthrough
rlabel pdiffusion 367 -2293 367 -2293 0 feedthrough
rlabel pdiffusion 381 -2293 381 -2293 0 feedthrough
rlabel pdiffusion 402 -2293 402 -2293 0 cellNo=480
rlabel pdiffusion 416 -2293 416 -2293 0 feedthrough
rlabel pdiffusion 423 -2293 423 -2293 0 feedthrough
rlabel pdiffusion 430 -2293 430 -2293 0 cellNo=75
rlabel pdiffusion 437 -2293 437 -2293 0 cellNo=933
rlabel pdiffusion 444 -2293 444 -2293 0 cellNo=978
rlabel pdiffusion 451 -2293 451 -2293 0 feedthrough
rlabel pdiffusion 458 -2293 458 -2293 0 feedthrough
rlabel pdiffusion 465 -2293 465 -2293 0 feedthrough
rlabel pdiffusion 472 -2293 472 -2293 0 cellNo=473
rlabel pdiffusion 479 -2293 479 -2293 0 cellNo=541
rlabel pdiffusion 500 -2293 500 -2293 0 cellNo=819
rlabel pdiffusion 507 -2293 507 -2293 0 feedthrough
rlabel pdiffusion 514 -2293 514 -2293 0 feedthrough
rlabel pdiffusion 521 -2293 521 -2293 0 feedthrough
rlabel pdiffusion 528 -2293 528 -2293 0 cellNo=517
rlabel pdiffusion 535 -2293 535 -2293 0 cellNo=821
rlabel pdiffusion 542 -2293 542 -2293 0 feedthrough
rlabel pdiffusion 549 -2293 549 -2293 0 cellNo=472
rlabel pdiffusion 570 -2293 570 -2293 0 cellNo=484
rlabel pdiffusion 577 -2293 577 -2293 0 feedthrough
rlabel pdiffusion 640 -2293 640 -2293 0 feedthrough
rlabel pdiffusion 171 -2310 171 -2310 0 cellNo=251
rlabel pdiffusion 178 -2310 178 -2310 0 feedthrough
rlabel pdiffusion 213 -2310 213 -2310 0 cellNo=782
rlabel pdiffusion 227 -2310 227 -2310 0 feedthrough
rlabel pdiffusion 234 -2310 234 -2310 0 feedthrough
rlabel pdiffusion 241 -2310 241 -2310 0 cellNo=198
rlabel pdiffusion 248 -2310 248 -2310 0 feedthrough
rlabel pdiffusion 255 -2310 255 -2310 0 feedthrough
rlabel pdiffusion 262 -2310 262 -2310 0 cellNo=37
rlabel pdiffusion 269 -2310 269 -2310 0 cellNo=755
rlabel pdiffusion 276 -2310 276 -2310 0 cellNo=843
rlabel pdiffusion 283 -2310 283 -2310 0 cellNo=353
rlabel pdiffusion 290 -2310 290 -2310 0 cellNo=614
rlabel pdiffusion 297 -2310 297 -2310 0 feedthrough
rlabel pdiffusion 304 -2310 304 -2310 0 cellNo=869
rlabel pdiffusion 311 -2310 311 -2310 0 cellNo=100
rlabel pdiffusion 318 -2310 318 -2310 0 feedthrough
rlabel pdiffusion 367 -2310 367 -2310 0 cellNo=428
rlabel pdiffusion 381 -2310 381 -2310 0 feedthrough
rlabel pdiffusion 388 -2310 388 -2310 0 cellNo=24
rlabel pdiffusion 402 -2310 402 -2310 0 cellNo=946
rlabel pdiffusion 409 -2310 409 -2310 0 feedthrough
rlabel pdiffusion 507 -2310 507 -2310 0 cellNo=853
rlabel pdiffusion 528 -2310 528 -2310 0 feedthrough
rlabel pdiffusion 535 -2310 535 -2310 0 cellNo=494
rlabel pdiffusion 598 -2310 598 -2310 0 feedthrough
rlabel pdiffusion 605 -2310 605 -2310 0 cellNo=642
rlabel pdiffusion 612 -2310 612 -2310 0 cellNo=759
rlabel pdiffusion 640 -2310 640 -2310 0 cellNo=940
rlabel pdiffusion 647 -2310 647 -2310 0 feedthrough
rlabel polysilicon 177 -4 177 -4 0 1
rlabel polysilicon 177 -10 177 -10 0 3
rlabel polysilicon 184 -10 184 -10 0 3
rlabel polysilicon 187 -10 187 -10 0 4
rlabel polysilicon 191 -4 191 -4 0 1
rlabel polysilicon 194 -10 194 -10 0 4
rlabel polysilicon 198 -10 198 -10 0 3
rlabel polysilicon 201 -10 201 -10 0 4
rlabel polysilicon 205 -4 205 -4 0 1
rlabel polysilicon 208 -10 208 -10 0 4
rlabel polysilicon 212 -4 212 -4 0 1
rlabel polysilicon 212 -10 212 -10 0 3
rlabel polysilicon 257 -4 257 -4 0 2
rlabel polysilicon 254 -10 254 -10 0 3
rlabel polysilicon 271 -4 271 -4 0 2
rlabel polysilicon 275 -4 275 -4 0 1
rlabel polysilicon 275 -10 275 -10 0 3
rlabel polysilicon 282 -4 282 -4 0 1
rlabel polysilicon 282 -10 282 -10 0 3
rlabel polysilicon 310 -4 310 -4 0 1
rlabel polysilicon 310 -10 310 -10 0 3
rlabel polysilicon 348 -4 348 -4 0 2
rlabel polysilicon 348 -10 348 -10 0 4
rlabel polysilicon 359 -4 359 -4 0 1
rlabel polysilicon 366 -4 366 -4 0 1
rlabel polysilicon 366 -10 366 -10 0 3
rlabel polysilicon 156 -27 156 -27 0 3
rlabel polysilicon 198 -21 198 -21 0 1
rlabel polysilicon 215 -21 215 -21 0 2
rlabel polysilicon 212 -27 212 -27 0 3
rlabel polysilicon 215 -27 215 -27 0 4
rlabel polysilicon 219 -21 219 -21 0 1
rlabel polysilicon 219 -27 219 -27 0 3
rlabel polysilicon 233 -21 233 -21 0 1
rlabel polysilicon 233 -27 233 -27 0 3
rlabel polysilicon 240 -21 240 -21 0 1
rlabel polysilicon 240 -27 240 -27 0 3
rlabel polysilicon 250 -21 250 -21 0 2
rlabel polysilicon 254 -21 254 -21 0 1
rlabel polysilicon 254 -27 254 -27 0 3
rlabel polysilicon 261 -21 261 -21 0 1
rlabel polysilicon 261 -27 261 -27 0 3
rlabel polysilicon 271 -27 271 -27 0 4
rlabel polysilicon 282 -21 282 -21 0 1
rlabel polysilicon 282 -27 282 -27 0 3
rlabel polysilicon 296 -27 296 -27 0 3
rlabel polysilicon 303 -21 303 -21 0 1
rlabel polysilicon 303 -27 303 -27 0 3
rlabel polysilicon 334 -27 334 -27 0 4
rlabel polysilicon 341 -21 341 -21 0 2
rlabel polysilicon 341 -27 341 -27 0 4
rlabel polysilicon 366 -21 366 -21 0 1
rlabel polysilicon 366 -27 366 -27 0 3
rlabel polysilicon 373 -21 373 -21 0 1
rlabel polysilicon 373 -27 373 -27 0 3
rlabel polysilicon 383 -21 383 -21 0 2
rlabel polysilicon 380 -27 380 -27 0 3
rlabel polysilicon 387 -21 387 -21 0 1
rlabel polysilicon 387 -27 387 -27 0 3
rlabel polysilicon 394 -21 394 -21 0 1
rlabel polysilicon 394 -27 394 -27 0 3
rlabel polysilicon 100 -48 100 -48 0 3
rlabel polysilicon 107 -48 107 -48 0 3
rlabel polysilicon 156 -42 156 -42 0 1
rlabel polysilicon 156 -48 156 -48 0 3
rlabel polysilicon 166 -42 166 -42 0 2
rlabel polysilicon 170 -48 170 -48 0 3
rlabel polysilicon 177 -42 177 -42 0 1
rlabel polysilicon 177 -48 177 -48 0 3
rlabel polysilicon 187 -48 187 -48 0 4
rlabel polysilicon 194 -42 194 -42 0 2
rlabel polysilicon 198 -42 198 -42 0 1
rlabel polysilicon 198 -48 198 -48 0 3
rlabel polysilicon 205 -42 205 -42 0 1
rlabel polysilicon 205 -48 205 -48 0 3
rlabel polysilicon 212 -42 212 -42 0 1
rlabel polysilicon 215 -48 215 -48 0 4
rlabel polysilicon 219 -42 219 -42 0 1
rlabel polysilicon 219 -48 219 -48 0 3
rlabel polysilicon 226 -42 226 -42 0 1
rlabel polysilicon 226 -48 226 -48 0 3
rlabel polysilicon 233 -42 233 -42 0 1
rlabel polysilicon 240 -42 240 -42 0 1
rlabel polysilicon 240 -48 240 -48 0 3
rlabel polysilicon 247 -42 247 -42 0 1
rlabel polysilicon 247 -48 247 -48 0 3
rlabel polysilicon 254 -42 254 -42 0 1
rlabel polysilicon 261 -42 261 -42 0 1
rlabel polysilicon 261 -48 261 -48 0 3
rlabel polysilicon 268 -42 268 -42 0 1
rlabel polysilicon 268 -48 268 -48 0 3
rlabel polysilicon 275 -42 275 -42 0 1
rlabel polysilicon 275 -48 275 -48 0 3
rlabel polysilicon 282 -42 282 -42 0 1
rlabel polysilicon 282 -48 282 -48 0 3
rlabel polysilicon 289 -42 289 -42 0 1
rlabel polysilicon 289 -48 289 -48 0 3
rlabel polysilicon 296 -42 296 -42 0 1
rlabel polysilicon 299 -42 299 -42 0 2
rlabel polysilicon 303 -48 303 -48 0 3
rlabel polysilicon 310 -42 310 -42 0 1
rlabel polysilicon 310 -48 310 -48 0 3
rlabel polysilicon 317 -42 317 -42 0 1
rlabel polysilicon 317 -48 317 -48 0 3
rlabel polysilicon 324 -42 324 -42 0 1
rlabel polysilicon 324 -48 324 -48 0 3
rlabel polysilicon 331 -42 331 -42 0 1
rlabel polysilicon 331 -48 331 -48 0 3
rlabel polysilicon 338 -42 338 -42 0 1
rlabel polysilicon 338 -48 338 -48 0 3
rlabel polysilicon 345 -42 345 -42 0 1
rlabel polysilicon 345 -48 345 -48 0 3
rlabel polysilicon 352 -42 352 -42 0 1
rlabel polysilicon 352 -48 352 -48 0 3
rlabel polysilicon 362 -48 362 -48 0 4
rlabel polysilicon 366 -42 366 -42 0 1
rlabel polysilicon 366 -48 366 -48 0 3
rlabel polysilicon 373 -42 373 -42 0 1
rlabel polysilicon 376 -48 376 -48 0 4
rlabel polysilicon 380 -42 380 -42 0 1
rlabel polysilicon 387 -42 387 -42 0 1
rlabel polysilicon 387 -48 387 -48 0 3
rlabel polysilicon 394 -42 394 -42 0 1
rlabel polysilicon 394 -48 394 -48 0 3
rlabel polysilicon 401 -48 401 -48 0 3
rlabel polysilicon 411 -42 411 -42 0 2
rlabel polysilicon 415 -42 415 -42 0 1
rlabel polysilicon 415 -48 415 -48 0 3
rlabel polysilicon 422 -42 422 -42 0 1
rlabel polysilicon 422 -48 422 -48 0 3
rlabel polysilicon 429 -42 429 -42 0 1
rlabel polysilicon 429 -48 429 -48 0 3
rlabel polysilicon 436 -48 436 -48 0 3
rlabel polysilicon 443 -48 443 -48 0 3
rlabel polysilicon 450 -42 450 -42 0 1
rlabel polysilicon 450 -48 450 -48 0 3
rlabel polysilicon 86 -79 86 -79 0 1
rlabel polysilicon 86 -85 86 -85 0 3
rlabel polysilicon 93 -79 93 -79 0 1
rlabel polysilicon 93 -85 93 -85 0 3
rlabel polysilicon 100 -79 100 -79 0 1
rlabel polysilicon 100 -85 100 -85 0 3
rlabel polysilicon 107 -79 107 -79 0 1
rlabel polysilicon 114 -85 114 -85 0 3
rlabel polysilicon 117 -85 117 -85 0 4
rlabel polysilicon 121 -79 121 -79 0 1
rlabel polysilicon 124 -85 124 -85 0 4
rlabel polysilicon 128 -79 128 -79 0 1
rlabel polysilicon 128 -85 128 -85 0 3
rlabel polysilicon 135 -79 135 -79 0 1
rlabel polysilicon 135 -85 135 -85 0 3
rlabel polysilicon 142 -79 142 -79 0 1
rlabel polysilicon 142 -85 142 -85 0 3
rlabel polysilicon 149 -79 149 -79 0 1
rlabel polysilicon 149 -85 149 -85 0 3
rlabel polysilicon 156 -79 156 -79 0 1
rlabel polysilicon 156 -85 156 -85 0 3
rlabel polysilicon 163 -79 163 -79 0 1
rlabel polysilicon 163 -85 163 -85 0 3
rlabel polysilicon 170 -79 170 -79 0 1
rlabel polysilicon 170 -85 170 -85 0 3
rlabel polysilicon 177 -79 177 -79 0 1
rlabel polysilicon 177 -85 177 -85 0 3
rlabel polysilicon 184 -85 184 -85 0 3
rlabel polysilicon 191 -79 191 -79 0 1
rlabel polysilicon 191 -85 191 -85 0 3
rlabel polysilicon 198 -79 198 -79 0 1
rlabel polysilicon 205 -79 205 -79 0 1
rlabel polysilicon 205 -85 205 -85 0 3
rlabel polysilicon 215 -79 215 -79 0 2
rlabel polysilicon 219 -79 219 -79 0 1
rlabel polysilicon 222 -85 222 -85 0 4
rlabel polysilicon 226 -79 226 -79 0 1
rlabel polysilicon 226 -85 226 -85 0 3
rlabel polysilicon 233 -79 233 -79 0 1
rlabel polysilicon 233 -85 233 -85 0 3
rlabel polysilicon 243 -79 243 -79 0 2
rlabel polysilicon 243 -85 243 -85 0 4
rlabel polysilicon 247 -79 247 -79 0 1
rlabel polysilicon 247 -85 247 -85 0 3
rlabel polysilicon 254 -85 254 -85 0 3
rlabel polysilicon 261 -79 261 -79 0 1
rlabel polysilicon 261 -85 261 -85 0 3
rlabel polysilicon 268 -79 268 -79 0 1
rlabel polysilicon 268 -85 268 -85 0 3
rlabel polysilicon 275 -79 275 -79 0 1
rlabel polysilicon 275 -85 275 -85 0 3
rlabel polysilicon 282 -79 282 -79 0 1
rlabel polysilicon 282 -85 282 -85 0 3
rlabel polysilicon 289 -79 289 -79 0 1
rlabel polysilicon 289 -85 289 -85 0 3
rlabel polysilicon 296 -79 296 -79 0 1
rlabel polysilicon 296 -85 296 -85 0 3
rlabel polysilicon 303 -79 303 -79 0 1
rlabel polysilicon 303 -85 303 -85 0 3
rlabel polysilicon 310 -79 310 -79 0 1
rlabel polysilicon 313 -85 313 -85 0 4
rlabel polysilicon 317 -79 317 -79 0 1
rlabel polysilicon 317 -85 317 -85 0 3
rlabel polysilicon 324 -79 324 -79 0 1
rlabel polysilicon 324 -85 324 -85 0 3
rlabel polysilicon 331 -79 331 -79 0 1
rlabel polysilicon 331 -85 331 -85 0 3
rlabel polysilicon 338 -79 338 -79 0 1
rlabel polysilicon 341 -79 341 -79 0 2
rlabel polysilicon 348 -79 348 -79 0 2
rlabel polysilicon 345 -85 345 -85 0 3
rlabel polysilicon 348 -85 348 -85 0 4
rlabel polysilicon 355 -79 355 -79 0 2
rlabel polysilicon 355 -85 355 -85 0 4
rlabel polysilicon 362 -79 362 -79 0 2
rlabel polysilicon 362 -85 362 -85 0 4
rlabel polysilicon 369 -79 369 -79 0 2
rlabel polysilicon 366 -85 366 -85 0 3
rlabel polysilicon 373 -79 373 -79 0 1
rlabel polysilicon 373 -85 373 -85 0 3
rlabel polysilicon 380 -79 380 -79 0 1
rlabel polysilicon 380 -85 380 -85 0 3
rlabel polysilicon 387 -79 387 -79 0 1
rlabel polysilicon 387 -85 387 -85 0 3
rlabel polysilicon 394 -79 394 -79 0 1
rlabel polysilicon 394 -85 394 -85 0 3
rlabel polysilicon 401 -79 401 -79 0 1
rlabel polysilicon 401 -85 401 -85 0 3
rlabel polysilicon 408 -79 408 -79 0 1
rlabel polysilicon 408 -85 408 -85 0 3
rlabel polysilicon 415 -79 415 -79 0 1
rlabel polysilicon 415 -85 415 -85 0 3
rlabel polysilicon 422 -79 422 -79 0 1
rlabel polysilicon 422 -85 422 -85 0 3
rlabel polysilicon 429 -79 429 -79 0 1
rlabel polysilicon 429 -85 429 -85 0 3
rlabel polysilicon 436 -79 436 -79 0 1
rlabel polysilicon 436 -85 436 -85 0 3
rlabel polysilicon 443 -79 443 -79 0 1
rlabel polysilicon 443 -85 443 -85 0 3
rlabel polysilicon 450 -79 450 -79 0 1
rlabel polysilicon 450 -85 450 -85 0 3
rlabel polysilicon 457 -79 457 -79 0 1
rlabel polysilicon 457 -85 457 -85 0 3
rlabel polysilicon 464 -79 464 -79 0 1
rlabel polysilicon 464 -85 464 -85 0 3
rlabel polysilicon 471 -79 471 -79 0 1
rlabel polysilicon 471 -85 471 -85 0 3
rlabel polysilicon 478 -79 478 -79 0 1
rlabel polysilicon 478 -85 478 -85 0 3
rlabel polysilicon 485 -79 485 -79 0 1
rlabel polysilicon 485 -85 485 -85 0 3
rlabel polysilicon 495 -79 495 -79 0 2
rlabel polysilicon 499 -79 499 -79 0 1
rlabel polysilicon 499 -85 499 -85 0 3
rlabel polysilicon 506 -85 506 -85 0 3
rlabel polysilicon 562 -85 562 -85 0 3
rlabel polysilicon 565 -85 565 -85 0 4
rlabel polysilicon 579 -79 579 -79 0 2
rlabel polysilicon 583 -79 583 -79 0 1
rlabel polysilicon 583 -85 583 -85 0 3
rlabel polysilicon 51 -140 51 -140 0 3
rlabel polysilicon 58 -134 58 -134 0 1
rlabel polysilicon 58 -140 58 -140 0 3
rlabel polysilicon 65 -134 65 -134 0 1
rlabel polysilicon 65 -140 65 -140 0 3
rlabel polysilicon 72 -134 72 -134 0 1
rlabel polysilicon 72 -140 72 -140 0 3
rlabel polysilicon 79 -134 79 -134 0 1
rlabel polysilicon 79 -140 79 -140 0 3
rlabel polysilicon 86 -134 86 -134 0 1
rlabel polysilicon 86 -140 86 -140 0 3
rlabel polysilicon 93 -134 93 -134 0 1
rlabel polysilicon 93 -140 93 -140 0 3
rlabel polysilicon 100 -134 100 -134 0 1
rlabel polysilicon 107 -134 107 -134 0 1
rlabel polysilicon 107 -140 107 -140 0 3
rlabel polysilicon 114 -134 114 -134 0 1
rlabel polysilicon 114 -140 114 -140 0 3
rlabel polysilicon 121 -134 121 -134 0 1
rlabel polysilicon 121 -140 121 -140 0 3
rlabel polysilicon 128 -134 128 -134 0 1
rlabel polysilicon 128 -140 128 -140 0 3
rlabel polysilicon 135 -134 135 -134 0 1
rlabel polysilicon 135 -140 135 -140 0 3
rlabel polysilicon 142 -134 142 -134 0 1
rlabel polysilicon 142 -140 142 -140 0 3
rlabel polysilicon 149 -134 149 -134 0 1
rlabel polysilicon 149 -140 149 -140 0 3
rlabel polysilicon 156 -134 156 -134 0 1
rlabel polysilicon 156 -140 156 -140 0 3
rlabel polysilicon 163 -134 163 -134 0 1
rlabel polysilicon 163 -140 163 -140 0 3
rlabel polysilicon 170 -134 170 -134 0 1
rlabel polysilicon 170 -140 170 -140 0 3
rlabel polysilicon 177 -134 177 -134 0 1
rlabel polysilicon 180 -134 180 -134 0 2
rlabel polysilicon 177 -140 177 -140 0 3
rlabel polysilicon 180 -140 180 -140 0 4
rlabel polysilicon 184 -134 184 -134 0 1
rlabel polysilicon 187 -134 187 -134 0 2
rlabel polysilicon 187 -140 187 -140 0 4
rlabel polysilicon 191 -140 191 -140 0 3
rlabel polysilicon 194 -140 194 -140 0 4
rlabel polysilicon 198 -134 198 -134 0 1
rlabel polysilicon 198 -140 198 -140 0 3
rlabel polysilicon 205 -134 205 -134 0 1
rlabel polysilicon 205 -140 205 -140 0 3
rlabel polysilicon 212 -140 212 -140 0 3
rlabel polysilicon 215 -140 215 -140 0 4
rlabel polysilicon 222 -134 222 -134 0 2
rlabel polysilicon 222 -140 222 -140 0 4
rlabel polysilicon 226 -134 226 -134 0 1
rlabel polysilicon 226 -140 226 -140 0 3
rlabel polysilicon 229 -140 229 -140 0 4
rlabel polysilicon 233 -134 233 -134 0 1
rlabel polysilicon 233 -140 233 -140 0 3
rlabel polysilicon 240 -134 240 -134 0 1
rlabel polysilicon 243 -134 243 -134 0 2
rlabel polysilicon 243 -140 243 -140 0 4
rlabel polysilicon 247 -134 247 -134 0 1
rlabel polysilicon 247 -140 247 -140 0 3
rlabel polysilicon 254 -134 254 -134 0 1
rlabel polysilicon 254 -140 254 -140 0 3
rlabel polysilicon 261 -134 261 -134 0 1
rlabel polysilicon 261 -140 261 -140 0 3
rlabel polysilicon 268 -134 268 -134 0 1
rlabel polysilicon 268 -140 268 -140 0 3
rlabel polysilicon 275 -134 275 -134 0 1
rlabel polysilicon 275 -140 275 -140 0 3
rlabel polysilicon 282 -134 282 -134 0 1
rlabel polysilicon 285 -134 285 -134 0 2
rlabel polysilicon 282 -140 282 -140 0 3
rlabel polysilicon 285 -140 285 -140 0 4
rlabel polysilicon 289 -134 289 -134 0 1
rlabel polysilicon 289 -140 289 -140 0 3
rlabel polysilicon 296 -134 296 -134 0 1
rlabel polysilicon 299 -134 299 -134 0 2
rlabel polysilicon 296 -140 296 -140 0 3
rlabel polysilicon 299 -140 299 -140 0 4
rlabel polysilicon 303 -134 303 -134 0 1
rlabel polysilicon 306 -134 306 -134 0 2
rlabel polysilicon 310 -134 310 -134 0 1
rlabel polysilicon 310 -140 310 -140 0 3
rlabel polysilicon 317 -134 317 -134 0 1
rlabel polysilicon 317 -140 317 -140 0 3
rlabel polysilicon 324 -134 324 -134 0 1
rlabel polysilicon 324 -140 324 -140 0 3
rlabel polysilicon 331 -134 331 -134 0 1
rlabel polysilicon 334 -134 334 -134 0 2
rlabel polysilicon 331 -140 331 -140 0 3
rlabel polysilicon 338 -140 338 -140 0 3
rlabel polysilicon 341 -140 341 -140 0 4
rlabel polysilicon 345 -134 345 -134 0 1
rlabel polysilicon 345 -140 345 -140 0 3
rlabel polysilicon 352 -134 352 -134 0 1
rlabel polysilicon 352 -140 352 -140 0 3
rlabel polysilicon 355 -140 355 -140 0 4
rlabel polysilicon 359 -134 359 -134 0 1
rlabel polysilicon 362 -134 362 -134 0 2
rlabel polysilicon 359 -140 359 -140 0 3
rlabel polysilicon 362 -140 362 -140 0 4
rlabel polysilicon 366 -134 366 -134 0 1
rlabel polysilicon 369 -134 369 -134 0 2
rlabel polysilicon 366 -140 366 -140 0 3
rlabel polysilicon 373 -134 373 -134 0 1
rlabel polysilicon 376 -134 376 -134 0 2
rlabel polysilicon 376 -140 376 -140 0 4
rlabel polysilicon 383 -134 383 -134 0 2
rlabel polysilicon 380 -140 380 -140 0 3
rlabel polysilicon 387 -134 387 -134 0 1
rlabel polysilicon 387 -140 387 -140 0 3
rlabel polysilicon 390 -140 390 -140 0 4
rlabel polysilicon 394 -134 394 -134 0 1
rlabel polysilicon 394 -140 394 -140 0 3
rlabel polysilicon 401 -134 401 -134 0 1
rlabel polysilicon 401 -140 401 -140 0 3
rlabel polysilicon 408 -134 408 -134 0 1
rlabel polysilicon 408 -140 408 -140 0 3
rlabel polysilicon 415 -134 415 -134 0 1
rlabel polysilicon 415 -140 415 -140 0 3
rlabel polysilicon 422 -134 422 -134 0 1
rlabel polysilicon 422 -140 422 -140 0 3
rlabel polysilicon 429 -134 429 -134 0 1
rlabel polysilicon 429 -140 429 -140 0 3
rlabel polysilicon 436 -134 436 -134 0 1
rlabel polysilicon 436 -140 436 -140 0 3
rlabel polysilicon 443 -134 443 -134 0 1
rlabel polysilicon 443 -140 443 -140 0 3
rlabel polysilicon 450 -134 450 -134 0 1
rlabel polysilicon 450 -140 450 -140 0 3
rlabel polysilicon 457 -134 457 -134 0 1
rlabel polysilicon 457 -140 457 -140 0 3
rlabel polysilicon 464 -134 464 -134 0 1
rlabel polysilicon 464 -140 464 -140 0 3
rlabel polysilicon 471 -134 471 -134 0 1
rlabel polysilicon 471 -140 471 -140 0 3
rlabel polysilicon 478 -134 478 -134 0 1
rlabel polysilicon 478 -140 478 -140 0 3
rlabel polysilicon 485 -134 485 -134 0 1
rlabel polysilicon 485 -140 485 -140 0 3
rlabel polysilicon 492 -134 492 -134 0 1
rlabel polysilicon 492 -140 492 -140 0 3
rlabel polysilicon 499 -134 499 -134 0 1
rlabel polysilicon 499 -140 499 -140 0 3
rlabel polysilicon 506 -134 506 -134 0 1
rlabel polysilicon 506 -140 506 -140 0 3
rlabel polysilicon 513 -134 513 -134 0 1
rlabel polysilicon 513 -140 513 -140 0 3
rlabel polysilicon 520 -134 520 -134 0 1
rlabel polysilicon 520 -140 520 -140 0 3
rlabel polysilicon 527 -134 527 -134 0 1
rlabel polysilicon 527 -140 527 -140 0 3
rlabel polysilicon 534 -134 534 -134 0 1
rlabel polysilicon 534 -140 534 -140 0 3
rlabel polysilicon 541 -134 541 -134 0 1
rlabel polysilicon 541 -140 541 -140 0 3
rlabel polysilicon 551 -140 551 -140 0 4
rlabel polysilicon 555 -134 555 -134 0 1
rlabel polysilicon 555 -140 555 -140 0 3
rlabel polysilicon 562 -134 562 -134 0 1
rlabel polysilicon 562 -140 562 -140 0 3
rlabel polysilicon 569 -134 569 -134 0 1
rlabel polysilicon 569 -140 569 -140 0 3
rlabel polysilicon 576 -134 576 -134 0 1
rlabel polysilicon 576 -140 576 -140 0 3
rlabel polysilicon 583 -134 583 -134 0 1
rlabel polysilicon 583 -140 583 -140 0 3
rlabel polysilicon 590 -134 590 -134 0 1
rlabel polysilicon 590 -140 590 -140 0 3
rlabel polysilicon 597 -134 597 -134 0 1
rlabel polysilicon 597 -140 597 -140 0 3
rlabel polysilicon 618 -134 618 -134 0 1
rlabel polysilicon 618 -140 618 -140 0 3
rlabel polysilicon 65 -193 65 -193 0 1
rlabel polysilicon 65 -199 65 -199 0 3
rlabel polysilicon 72 -199 72 -199 0 3
rlabel polysilicon 79 -193 79 -193 0 1
rlabel polysilicon 79 -199 79 -199 0 3
rlabel polysilicon 86 -193 86 -193 0 1
rlabel polysilicon 86 -199 86 -199 0 3
rlabel polysilicon 93 -193 93 -193 0 1
rlabel polysilicon 93 -199 93 -199 0 3
rlabel polysilicon 100 -193 100 -193 0 1
rlabel polysilicon 100 -199 100 -199 0 3
rlabel polysilicon 107 -193 107 -193 0 1
rlabel polysilicon 107 -199 107 -199 0 3
rlabel polysilicon 114 -193 114 -193 0 1
rlabel polysilicon 114 -199 114 -199 0 3
rlabel polysilicon 121 -193 121 -193 0 1
rlabel polysilicon 121 -199 121 -199 0 3
rlabel polysilicon 128 -193 128 -193 0 1
rlabel polysilicon 128 -199 128 -199 0 3
rlabel polysilicon 135 -193 135 -193 0 1
rlabel polysilicon 138 -193 138 -193 0 2
rlabel polysilicon 138 -199 138 -199 0 4
rlabel polysilicon 142 -193 142 -193 0 1
rlabel polysilicon 142 -199 142 -199 0 3
rlabel polysilicon 149 -193 149 -193 0 1
rlabel polysilicon 149 -199 149 -199 0 3
rlabel polysilicon 156 -193 156 -193 0 1
rlabel polysilicon 156 -199 156 -199 0 3
rlabel polysilicon 163 -193 163 -193 0 1
rlabel polysilicon 163 -199 163 -199 0 3
rlabel polysilicon 170 -193 170 -193 0 1
rlabel polysilicon 173 -193 173 -193 0 2
rlabel polysilicon 173 -199 173 -199 0 4
rlabel polysilicon 177 -193 177 -193 0 1
rlabel polysilicon 177 -199 177 -199 0 3
rlabel polysilicon 187 -193 187 -193 0 2
rlabel polysilicon 184 -199 184 -199 0 3
rlabel polysilicon 187 -199 187 -199 0 4
rlabel polysilicon 191 -199 191 -199 0 3
rlabel polysilicon 198 -193 198 -193 0 1
rlabel polysilicon 198 -199 198 -199 0 3
rlabel polysilicon 205 -193 205 -193 0 1
rlabel polysilicon 208 -193 208 -193 0 2
rlabel polysilicon 205 -199 205 -199 0 3
rlabel polysilicon 208 -199 208 -199 0 4
rlabel polysilicon 212 -193 212 -193 0 1
rlabel polysilicon 215 -193 215 -193 0 2
rlabel polysilicon 219 -193 219 -193 0 1
rlabel polysilicon 219 -199 219 -199 0 3
rlabel polysilicon 226 -193 226 -193 0 1
rlabel polysilicon 226 -199 226 -199 0 3
rlabel polysilicon 233 -193 233 -193 0 1
rlabel polysilicon 236 -193 236 -193 0 2
rlabel polysilicon 233 -199 233 -199 0 3
rlabel polysilicon 236 -199 236 -199 0 4
rlabel polysilicon 240 -193 240 -193 0 1
rlabel polysilicon 240 -199 240 -199 0 3
rlabel polysilicon 247 -193 247 -193 0 1
rlabel polysilicon 247 -199 247 -199 0 3
rlabel polysilicon 254 -193 254 -193 0 1
rlabel polysilicon 254 -199 254 -199 0 3
rlabel polysilicon 261 -193 261 -193 0 1
rlabel polysilicon 261 -199 261 -199 0 3
rlabel polysilicon 268 -193 268 -193 0 1
rlabel polysilicon 268 -199 268 -199 0 3
rlabel polysilicon 275 -193 275 -193 0 1
rlabel polysilicon 275 -199 275 -199 0 3
rlabel polysilicon 282 -193 282 -193 0 1
rlabel polysilicon 282 -199 282 -199 0 3
rlabel polysilicon 289 -193 289 -193 0 1
rlabel polysilicon 289 -199 289 -199 0 3
rlabel polysilicon 296 -193 296 -193 0 1
rlabel polysilicon 296 -199 296 -199 0 3
rlabel polysilicon 299 -199 299 -199 0 4
rlabel polysilicon 306 -193 306 -193 0 2
rlabel polysilicon 303 -199 303 -199 0 3
rlabel polysilicon 310 -193 310 -193 0 1
rlabel polysilicon 310 -199 310 -199 0 3
rlabel polysilicon 317 -193 317 -193 0 1
rlabel polysilicon 320 -193 320 -193 0 2
rlabel polysilicon 317 -199 317 -199 0 3
rlabel polysilicon 320 -199 320 -199 0 4
rlabel polysilicon 324 -193 324 -193 0 1
rlabel polysilicon 324 -199 324 -199 0 3
rlabel polysilicon 331 -193 331 -193 0 1
rlabel polysilicon 331 -199 331 -199 0 3
rlabel polysilicon 338 -193 338 -193 0 1
rlabel polysilicon 338 -199 338 -199 0 3
rlabel polysilicon 345 -193 345 -193 0 1
rlabel polysilicon 345 -199 345 -199 0 3
rlabel polysilicon 352 -193 352 -193 0 1
rlabel polysilicon 355 -193 355 -193 0 2
rlabel polysilicon 355 -199 355 -199 0 4
rlabel polysilicon 359 -193 359 -193 0 1
rlabel polysilicon 362 -193 362 -193 0 2
rlabel polysilicon 366 -193 366 -193 0 1
rlabel polysilicon 366 -199 366 -199 0 3
rlabel polysilicon 373 -193 373 -193 0 1
rlabel polysilicon 376 -193 376 -193 0 2
rlabel polysilicon 373 -199 373 -199 0 3
rlabel polysilicon 376 -199 376 -199 0 4
rlabel polysilicon 380 -193 380 -193 0 1
rlabel polysilicon 380 -199 380 -199 0 3
rlabel polysilicon 387 -193 387 -193 0 1
rlabel polysilicon 387 -199 387 -199 0 3
rlabel polysilicon 394 -199 394 -199 0 3
rlabel polysilicon 397 -199 397 -199 0 4
rlabel polysilicon 404 -193 404 -193 0 2
rlabel polysilicon 404 -199 404 -199 0 4
rlabel polysilicon 408 -193 408 -193 0 1
rlabel polysilicon 408 -199 408 -199 0 3
rlabel polysilicon 415 -193 415 -193 0 1
rlabel polysilicon 415 -199 415 -199 0 3
rlabel polysilicon 422 -193 422 -193 0 1
rlabel polysilicon 422 -199 422 -199 0 3
rlabel polysilicon 429 -193 429 -193 0 1
rlabel polysilicon 429 -199 429 -199 0 3
rlabel polysilicon 439 -193 439 -193 0 2
rlabel polysilicon 439 -199 439 -199 0 4
rlabel polysilicon 443 -193 443 -193 0 1
rlabel polysilicon 443 -199 443 -199 0 3
rlabel polysilicon 450 -193 450 -193 0 1
rlabel polysilicon 450 -199 450 -199 0 3
rlabel polysilicon 457 -193 457 -193 0 1
rlabel polysilicon 460 -199 460 -199 0 4
rlabel polysilicon 464 -193 464 -193 0 1
rlabel polysilicon 464 -199 464 -199 0 3
rlabel polysilicon 471 -193 471 -193 0 1
rlabel polysilicon 471 -199 471 -199 0 3
rlabel polysilicon 478 -193 478 -193 0 1
rlabel polysilicon 478 -199 478 -199 0 3
rlabel polysilicon 485 -193 485 -193 0 1
rlabel polysilicon 485 -199 485 -199 0 3
rlabel polysilicon 492 -193 492 -193 0 1
rlabel polysilicon 492 -199 492 -199 0 3
rlabel polysilicon 499 -193 499 -193 0 1
rlabel polysilicon 499 -199 499 -199 0 3
rlabel polysilicon 506 -199 506 -199 0 3
rlabel polysilicon 509 -199 509 -199 0 4
rlabel polysilicon 513 -193 513 -193 0 1
rlabel polysilicon 513 -199 513 -199 0 3
rlabel polysilicon 520 -193 520 -193 0 1
rlabel polysilicon 520 -199 520 -199 0 3
rlabel polysilicon 527 -193 527 -193 0 1
rlabel polysilicon 527 -199 527 -199 0 3
rlabel polysilicon 534 -193 534 -193 0 1
rlabel polysilicon 534 -199 534 -199 0 3
rlabel polysilicon 544 -193 544 -193 0 2
rlabel polysilicon 544 -199 544 -199 0 4
rlabel polysilicon 548 -193 548 -193 0 1
rlabel polysilicon 548 -199 548 -199 0 3
rlabel polysilicon 555 -193 555 -193 0 1
rlabel polysilicon 555 -199 555 -199 0 3
rlabel polysilicon 562 -193 562 -193 0 1
rlabel polysilicon 562 -199 562 -199 0 3
rlabel polysilicon 572 -193 572 -193 0 2
rlabel polysilicon 569 -199 569 -199 0 3
rlabel polysilicon 576 -193 576 -193 0 1
rlabel polysilicon 576 -199 576 -199 0 3
rlabel polysilicon 583 -193 583 -193 0 1
rlabel polysilicon 583 -199 583 -199 0 3
rlabel polysilicon 590 -193 590 -193 0 1
rlabel polysilicon 590 -199 590 -199 0 3
rlabel polysilicon 632 -193 632 -193 0 1
rlabel polysilicon 632 -199 632 -199 0 3
rlabel polysilicon 642 -193 642 -193 0 2
rlabel polysilicon 646 -193 646 -193 0 1
rlabel polysilicon 646 -199 646 -199 0 3
rlabel polysilicon 16 -250 16 -250 0 1
rlabel polysilicon 16 -256 16 -256 0 3
rlabel polysilicon 23 -250 23 -250 0 1
rlabel polysilicon 23 -256 23 -256 0 3
rlabel polysilicon 30 -250 30 -250 0 1
rlabel polysilicon 30 -256 30 -256 0 3
rlabel polysilicon 37 -250 37 -250 0 1
rlabel polysilicon 37 -256 37 -256 0 3
rlabel polysilicon 44 -250 44 -250 0 1
rlabel polysilicon 44 -256 44 -256 0 3
rlabel polysilicon 51 -250 51 -250 0 1
rlabel polysilicon 58 -250 58 -250 0 1
rlabel polysilicon 58 -256 58 -256 0 3
rlabel polysilicon 65 -250 65 -250 0 1
rlabel polysilicon 65 -256 65 -256 0 3
rlabel polysilicon 72 -250 72 -250 0 1
rlabel polysilicon 72 -256 72 -256 0 3
rlabel polysilicon 79 -250 79 -250 0 1
rlabel polysilicon 79 -256 79 -256 0 3
rlabel polysilicon 86 -250 86 -250 0 1
rlabel polysilicon 86 -256 86 -256 0 3
rlabel polysilicon 93 -250 93 -250 0 1
rlabel polysilicon 93 -256 93 -256 0 3
rlabel polysilicon 100 -250 100 -250 0 1
rlabel polysilicon 100 -256 100 -256 0 3
rlabel polysilicon 103 -256 103 -256 0 4
rlabel polysilicon 107 -250 107 -250 0 1
rlabel polysilicon 107 -256 107 -256 0 3
rlabel polysilicon 114 -250 114 -250 0 1
rlabel polysilicon 114 -256 114 -256 0 3
rlabel polysilicon 121 -250 121 -250 0 1
rlabel polysilicon 121 -256 121 -256 0 3
rlabel polysilicon 128 -250 128 -250 0 1
rlabel polysilicon 131 -250 131 -250 0 2
rlabel polysilicon 138 -250 138 -250 0 2
rlabel polysilicon 138 -256 138 -256 0 4
rlabel polysilicon 142 -250 142 -250 0 1
rlabel polysilicon 145 -250 145 -250 0 2
rlabel polysilicon 149 -250 149 -250 0 1
rlabel polysilicon 149 -256 149 -256 0 3
rlabel polysilicon 156 -256 156 -256 0 3
rlabel polysilicon 159 -256 159 -256 0 4
rlabel polysilicon 163 -250 163 -250 0 1
rlabel polysilicon 163 -256 163 -256 0 3
rlabel polysilicon 170 -250 170 -250 0 1
rlabel polysilicon 170 -256 170 -256 0 3
rlabel polysilicon 177 -250 177 -250 0 1
rlabel polysilicon 177 -256 177 -256 0 3
rlabel polysilicon 184 -250 184 -250 0 1
rlabel polysilicon 184 -256 184 -256 0 3
rlabel polysilicon 191 -250 191 -250 0 1
rlabel polysilicon 194 -250 194 -250 0 2
rlabel polysilicon 194 -256 194 -256 0 4
rlabel polysilicon 198 -250 198 -250 0 1
rlabel polysilicon 198 -256 198 -256 0 3
rlabel polysilicon 208 -250 208 -250 0 2
rlabel polysilicon 205 -256 205 -256 0 3
rlabel polysilicon 212 -250 212 -250 0 1
rlabel polysilicon 215 -256 215 -256 0 4
rlabel polysilicon 219 -250 219 -250 0 1
rlabel polysilicon 222 -250 222 -250 0 2
rlabel polysilicon 226 -250 226 -250 0 1
rlabel polysilicon 229 -250 229 -250 0 2
rlabel polysilicon 226 -256 226 -256 0 3
rlabel polysilicon 229 -256 229 -256 0 4
rlabel polysilicon 233 -250 233 -250 0 1
rlabel polysilicon 233 -256 233 -256 0 3
rlabel polysilicon 240 -250 240 -250 0 1
rlabel polysilicon 240 -256 240 -256 0 3
rlabel polysilicon 247 -250 247 -250 0 1
rlabel polysilicon 247 -256 247 -256 0 3
rlabel polysilicon 254 -250 254 -250 0 1
rlabel polysilicon 254 -256 254 -256 0 3
rlabel polysilicon 261 -250 261 -250 0 1
rlabel polysilicon 261 -256 261 -256 0 3
rlabel polysilicon 268 -250 268 -250 0 1
rlabel polysilicon 268 -256 268 -256 0 3
rlabel polysilicon 271 -256 271 -256 0 4
rlabel polysilicon 275 -250 275 -250 0 1
rlabel polysilicon 275 -256 275 -256 0 3
rlabel polysilicon 282 -250 282 -250 0 1
rlabel polysilicon 282 -256 282 -256 0 3
rlabel polysilicon 289 -250 289 -250 0 1
rlabel polysilicon 289 -256 289 -256 0 3
rlabel polysilicon 296 -250 296 -250 0 1
rlabel polysilicon 296 -256 296 -256 0 3
rlabel polysilicon 303 -250 303 -250 0 1
rlabel polysilicon 303 -256 303 -256 0 3
rlabel polysilicon 310 -250 310 -250 0 1
rlabel polysilicon 310 -256 310 -256 0 3
rlabel polysilicon 317 -250 317 -250 0 1
rlabel polysilicon 317 -256 317 -256 0 3
rlabel polysilicon 324 -250 324 -250 0 1
rlabel polysilicon 324 -256 324 -256 0 3
rlabel polysilicon 331 -250 331 -250 0 1
rlabel polysilicon 331 -256 331 -256 0 3
rlabel polysilicon 338 -250 338 -250 0 1
rlabel polysilicon 338 -256 338 -256 0 3
rlabel polysilicon 341 -256 341 -256 0 4
rlabel polysilicon 345 -250 345 -250 0 1
rlabel polysilicon 345 -256 345 -256 0 3
rlabel polysilicon 352 -250 352 -250 0 1
rlabel polysilicon 352 -256 352 -256 0 3
rlabel polysilicon 359 -250 359 -250 0 1
rlabel polysilicon 359 -256 359 -256 0 3
rlabel polysilicon 366 -250 366 -250 0 1
rlabel polysilicon 366 -256 366 -256 0 3
rlabel polysilicon 373 -250 373 -250 0 1
rlabel polysilicon 373 -256 373 -256 0 3
rlabel polysilicon 380 -250 380 -250 0 1
rlabel polysilicon 380 -256 380 -256 0 3
rlabel polysilicon 390 -250 390 -250 0 2
rlabel polysilicon 387 -256 387 -256 0 3
rlabel polysilicon 390 -256 390 -256 0 4
rlabel polysilicon 394 -250 394 -250 0 1
rlabel polysilicon 397 -250 397 -250 0 2
rlabel polysilicon 397 -256 397 -256 0 4
rlabel polysilicon 401 -250 401 -250 0 1
rlabel polysilicon 401 -256 401 -256 0 3
rlabel polysilicon 408 -250 408 -250 0 1
rlabel polysilicon 411 -250 411 -250 0 2
rlabel polysilicon 411 -256 411 -256 0 4
rlabel polysilicon 415 -250 415 -250 0 1
rlabel polysilicon 418 -250 418 -250 0 2
rlabel polysilicon 422 -250 422 -250 0 1
rlabel polysilicon 422 -256 422 -256 0 3
rlabel polysilicon 429 -250 429 -250 0 1
rlabel polysilicon 429 -256 429 -256 0 3
rlabel polysilicon 436 -250 436 -250 0 1
rlabel polysilicon 436 -256 436 -256 0 3
rlabel polysilicon 443 -250 443 -250 0 1
rlabel polysilicon 443 -256 443 -256 0 3
rlabel polysilicon 450 -250 450 -250 0 1
rlabel polysilicon 450 -256 450 -256 0 3
rlabel polysilicon 457 -250 457 -250 0 1
rlabel polysilicon 460 -256 460 -256 0 4
rlabel polysilicon 464 -250 464 -250 0 1
rlabel polysilicon 467 -250 467 -250 0 2
rlabel polysilicon 471 -250 471 -250 0 1
rlabel polysilicon 471 -256 471 -256 0 3
rlabel polysilicon 478 -250 478 -250 0 1
rlabel polysilicon 481 -256 481 -256 0 4
rlabel polysilicon 485 -250 485 -250 0 1
rlabel polysilicon 485 -256 485 -256 0 3
rlabel polysilicon 492 -250 492 -250 0 1
rlabel polysilicon 492 -256 492 -256 0 3
rlabel polysilicon 499 -250 499 -250 0 1
rlabel polysilicon 499 -256 499 -256 0 3
rlabel polysilicon 509 -250 509 -250 0 2
rlabel polysilicon 506 -256 506 -256 0 3
rlabel polysilicon 513 -250 513 -250 0 1
rlabel polysilicon 520 -250 520 -250 0 1
rlabel polysilicon 520 -256 520 -256 0 3
rlabel polysilicon 527 -250 527 -250 0 1
rlabel polysilicon 527 -256 527 -256 0 3
rlabel polysilicon 534 -250 534 -250 0 1
rlabel polysilicon 534 -256 534 -256 0 3
rlabel polysilicon 541 -250 541 -250 0 1
rlabel polysilicon 541 -256 541 -256 0 3
rlabel polysilicon 548 -250 548 -250 0 1
rlabel polysilicon 548 -256 548 -256 0 3
rlabel polysilicon 555 -250 555 -250 0 1
rlabel polysilicon 555 -256 555 -256 0 3
rlabel polysilicon 562 -250 562 -250 0 1
rlabel polysilicon 562 -256 562 -256 0 3
rlabel polysilicon 569 -250 569 -250 0 1
rlabel polysilicon 572 -256 572 -256 0 4
rlabel polysilicon 576 -250 576 -250 0 1
rlabel polysilicon 576 -256 576 -256 0 3
rlabel polysilicon 583 -250 583 -250 0 1
rlabel polysilicon 583 -256 583 -256 0 3
rlabel polysilicon 590 -250 590 -250 0 1
rlabel polysilicon 590 -256 590 -256 0 3
rlabel polysilicon 597 -250 597 -250 0 1
rlabel polysilicon 597 -256 597 -256 0 3
rlabel polysilicon 600 -256 600 -256 0 4
rlabel polysilicon 604 -250 604 -250 0 1
rlabel polysilicon 604 -256 604 -256 0 3
rlabel polysilicon 611 -250 611 -250 0 1
rlabel polysilicon 611 -256 611 -256 0 3
rlabel polysilicon 618 -250 618 -250 0 1
rlabel polysilicon 618 -256 618 -256 0 3
rlabel polysilicon 625 -250 625 -250 0 1
rlabel polysilicon 625 -256 625 -256 0 3
rlabel polysilicon 632 -250 632 -250 0 1
rlabel polysilicon 632 -256 632 -256 0 3
rlabel polysilicon 639 -250 639 -250 0 1
rlabel polysilicon 639 -256 639 -256 0 3
rlabel polysilicon 646 -250 646 -250 0 1
rlabel polysilicon 646 -256 646 -256 0 3
rlabel polysilicon 653 -250 653 -250 0 1
rlabel polysilicon 653 -256 653 -256 0 3
rlabel polysilicon 660 -250 660 -250 0 1
rlabel polysilicon 660 -256 660 -256 0 3
rlabel polysilicon 667 -250 667 -250 0 1
rlabel polysilicon 670 -250 670 -250 0 2
rlabel polysilicon 667 -256 667 -256 0 3
rlabel polysilicon 670 -256 670 -256 0 4
rlabel polysilicon 674 -250 674 -250 0 1
rlabel polysilicon 674 -256 674 -256 0 3
rlabel polysilicon 681 -250 681 -250 0 1
rlabel polysilicon 681 -256 681 -256 0 3
rlabel polysilicon 688 -250 688 -250 0 1
rlabel polysilicon 688 -256 688 -256 0 3
rlabel polysilicon 695 -250 695 -250 0 1
rlabel polysilicon 695 -256 695 -256 0 3
rlabel polysilicon 751 -250 751 -250 0 1
rlabel polysilicon 751 -256 751 -256 0 3
rlabel polysilicon 859 -256 859 -256 0 4
rlabel polysilicon 30 -303 30 -303 0 1
rlabel polysilicon 30 -309 30 -309 0 3
rlabel polysilicon 37 -303 37 -303 0 1
rlabel polysilicon 37 -309 37 -309 0 3
rlabel polysilicon 44 -309 44 -309 0 3
rlabel polysilicon 51 -303 51 -303 0 1
rlabel polysilicon 51 -309 51 -309 0 3
rlabel polysilicon 58 -303 58 -303 0 1
rlabel polysilicon 58 -309 58 -309 0 3
rlabel polysilicon 68 -303 68 -303 0 2
rlabel polysilicon 65 -309 65 -309 0 3
rlabel polysilicon 72 -303 72 -303 0 1
rlabel polysilicon 72 -309 72 -309 0 3
rlabel polysilicon 79 -303 79 -303 0 1
rlabel polysilicon 79 -309 79 -309 0 3
rlabel polysilicon 86 -303 86 -303 0 1
rlabel polysilicon 86 -309 86 -309 0 3
rlabel polysilicon 93 -303 93 -303 0 1
rlabel polysilicon 93 -309 93 -309 0 3
rlabel polysilicon 100 -303 100 -303 0 1
rlabel polysilicon 100 -309 100 -309 0 3
rlabel polysilicon 107 -303 107 -303 0 1
rlabel polysilicon 107 -309 107 -309 0 3
rlabel polysilicon 117 -303 117 -303 0 2
rlabel polysilicon 114 -309 114 -309 0 3
rlabel polysilicon 121 -303 121 -303 0 1
rlabel polysilicon 121 -309 121 -309 0 3
rlabel polysilicon 128 -303 128 -303 0 1
rlabel polysilicon 128 -309 128 -309 0 3
rlabel polysilicon 135 -303 135 -303 0 1
rlabel polysilicon 138 -309 138 -309 0 4
rlabel polysilicon 142 -303 142 -303 0 1
rlabel polysilicon 142 -309 142 -309 0 3
rlabel polysilicon 149 -303 149 -303 0 1
rlabel polysilicon 149 -309 149 -309 0 3
rlabel polysilicon 156 -303 156 -303 0 1
rlabel polysilicon 156 -309 156 -309 0 3
rlabel polysilicon 163 -303 163 -303 0 1
rlabel polysilicon 163 -309 163 -309 0 3
rlabel polysilicon 170 -303 170 -303 0 1
rlabel polysilicon 170 -309 170 -309 0 3
rlabel polysilicon 177 -303 177 -303 0 1
rlabel polysilicon 180 -303 180 -303 0 2
rlabel polysilicon 177 -309 177 -309 0 3
rlabel polysilicon 184 -303 184 -303 0 1
rlabel polysilicon 184 -309 184 -309 0 3
rlabel polysilicon 191 -303 191 -303 0 1
rlabel polysilicon 191 -309 191 -309 0 3
rlabel polysilicon 198 -303 198 -303 0 1
rlabel polysilicon 205 -303 205 -303 0 1
rlabel polysilicon 205 -309 205 -309 0 3
rlabel polysilicon 215 -303 215 -303 0 2
rlabel polysilicon 212 -309 212 -309 0 3
rlabel polysilicon 215 -309 215 -309 0 4
rlabel polysilicon 222 -303 222 -303 0 2
rlabel polysilicon 219 -309 219 -309 0 3
rlabel polysilicon 222 -309 222 -309 0 4
rlabel polysilicon 226 -303 226 -303 0 1
rlabel polysilicon 226 -309 226 -309 0 3
rlabel polysilicon 236 -303 236 -303 0 2
rlabel polysilicon 233 -309 233 -309 0 3
rlabel polysilicon 236 -309 236 -309 0 4
rlabel polysilicon 240 -303 240 -303 0 1
rlabel polysilicon 243 -303 243 -303 0 2
rlabel polysilicon 240 -309 240 -309 0 3
rlabel polysilicon 247 -309 247 -309 0 3
rlabel polysilicon 254 -303 254 -303 0 1
rlabel polysilicon 254 -309 254 -309 0 3
rlabel polysilicon 257 -309 257 -309 0 4
rlabel polysilicon 261 -303 261 -303 0 1
rlabel polysilicon 261 -309 261 -309 0 3
rlabel polysilicon 268 -303 268 -303 0 1
rlabel polysilicon 268 -309 268 -309 0 3
rlabel polysilicon 275 -303 275 -303 0 1
rlabel polysilicon 275 -309 275 -309 0 3
rlabel polysilicon 282 -303 282 -303 0 1
rlabel polysilicon 282 -309 282 -309 0 3
rlabel polysilicon 289 -309 289 -309 0 3
rlabel polysilicon 296 -303 296 -303 0 1
rlabel polysilicon 299 -303 299 -303 0 2
rlabel polysilicon 299 -309 299 -309 0 4
rlabel polysilicon 303 -303 303 -303 0 1
rlabel polysilicon 303 -309 303 -309 0 3
rlabel polysilicon 310 -303 310 -303 0 1
rlabel polysilicon 310 -309 310 -309 0 3
rlabel polysilicon 317 -303 317 -303 0 1
rlabel polysilicon 317 -309 317 -309 0 3
rlabel polysilicon 324 -303 324 -303 0 1
rlabel polysilicon 324 -309 324 -309 0 3
rlabel polysilicon 331 -303 331 -303 0 1
rlabel polysilicon 334 -303 334 -303 0 2
rlabel polysilicon 331 -309 331 -309 0 3
rlabel polysilicon 334 -309 334 -309 0 4
rlabel polysilicon 338 -303 338 -303 0 1
rlabel polysilicon 338 -309 338 -309 0 3
rlabel polysilicon 341 -309 341 -309 0 4
rlabel polysilicon 345 -303 345 -303 0 1
rlabel polysilicon 345 -309 345 -309 0 3
rlabel polysilicon 352 -303 352 -303 0 1
rlabel polysilicon 352 -309 352 -309 0 3
rlabel polysilicon 359 -303 359 -303 0 1
rlabel polysilicon 359 -309 359 -309 0 3
rlabel polysilicon 366 -303 366 -303 0 1
rlabel polysilicon 366 -309 366 -309 0 3
rlabel polysilicon 373 -303 373 -303 0 1
rlabel polysilicon 380 -303 380 -303 0 1
rlabel polysilicon 380 -309 380 -309 0 3
rlabel polysilicon 387 -303 387 -303 0 1
rlabel polysilicon 387 -309 387 -309 0 3
rlabel polysilicon 394 -303 394 -303 0 1
rlabel polysilicon 397 -303 397 -303 0 2
rlabel polysilicon 394 -309 394 -309 0 3
rlabel polysilicon 401 -303 401 -303 0 1
rlabel polysilicon 404 -303 404 -303 0 2
rlabel polysilicon 401 -309 401 -309 0 3
rlabel polysilicon 408 -303 408 -303 0 1
rlabel polysilicon 408 -309 408 -309 0 3
rlabel polysilicon 415 -303 415 -303 0 1
rlabel polysilicon 415 -309 415 -309 0 3
rlabel polysilicon 422 -303 422 -303 0 1
rlabel polysilicon 425 -303 425 -303 0 2
rlabel polysilicon 429 -303 429 -303 0 1
rlabel polysilicon 429 -309 429 -309 0 3
rlabel polysilicon 439 -303 439 -303 0 2
rlabel polysilicon 436 -309 436 -309 0 3
rlabel polysilicon 439 -309 439 -309 0 4
rlabel polysilicon 446 -303 446 -303 0 2
rlabel polysilicon 450 -303 450 -303 0 1
rlabel polysilicon 450 -309 450 -309 0 3
rlabel polysilicon 453 -309 453 -309 0 4
rlabel polysilicon 457 -303 457 -303 0 1
rlabel polysilicon 457 -309 457 -309 0 3
rlabel polysilicon 464 -303 464 -303 0 1
rlabel polysilicon 464 -309 464 -309 0 3
rlabel polysilicon 471 -303 471 -303 0 1
rlabel polysilicon 471 -309 471 -309 0 3
rlabel polysilicon 478 -303 478 -303 0 1
rlabel polysilicon 478 -309 478 -309 0 3
rlabel polysilicon 485 -303 485 -303 0 1
rlabel polysilicon 485 -309 485 -309 0 3
rlabel polysilicon 492 -303 492 -303 0 1
rlabel polysilicon 492 -309 492 -309 0 3
rlabel polysilicon 499 -303 499 -303 0 1
rlabel polysilicon 499 -309 499 -309 0 3
rlabel polysilicon 506 -303 506 -303 0 1
rlabel polysilicon 506 -309 506 -309 0 3
rlabel polysilicon 513 -309 513 -309 0 3
rlabel polysilicon 520 -303 520 -303 0 1
rlabel polysilicon 520 -309 520 -309 0 3
rlabel polysilicon 527 -303 527 -303 0 1
rlabel polysilicon 527 -309 527 -309 0 3
rlabel polysilicon 534 -303 534 -303 0 1
rlabel polysilicon 534 -309 534 -309 0 3
rlabel polysilicon 541 -303 541 -303 0 1
rlabel polysilicon 544 -303 544 -303 0 2
rlabel polysilicon 544 -309 544 -309 0 4
rlabel polysilicon 548 -303 548 -303 0 1
rlabel polysilicon 548 -309 548 -309 0 3
rlabel polysilicon 555 -303 555 -303 0 1
rlabel polysilicon 555 -309 555 -309 0 3
rlabel polysilicon 562 -303 562 -303 0 1
rlabel polysilicon 565 -303 565 -303 0 2
rlabel polysilicon 562 -309 562 -309 0 3
rlabel polysilicon 569 -303 569 -303 0 1
rlabel polysilicon 569 -309 569 -309 0 3
rlabel polysilicon 576 -303 576 -303 0 1
rlabel polysilicon 576 -309 576 -309 0 3
rlabel polysilicon 583 -303 583 -303 0 1
rlabel polysilicon 583 -309 583 -309 0 3
rlabel polysilicon 590 -303 590 -303 0 1
rlabel polysilicon 590 -309 590 -309 0 3
rlabel polysilicon 597 -303 597 -303 0 1
rlabel polysilicon 600 -303 600 -303 0 2
rlabel polysilicon 597 -309 597 -309 0 3
rlabel polysilicon 604 -303 604 -303 0 1
rlabel polysilicon 604 -309 604 -309 0 3
rlabel polysilicon 611 -303 611 -303 0 1
rlabel polysilicon 611 -309 611 -309 0 3
rlabel polysilicon 618 -303 618 -303 0 1
rlabel polysilicon 618 -309 618 -309 0 3
rlabel polysilicon 625 -303 625 -303 0 1
rlabel polysilicon 625 -309 625 -309 0 3
rlabel polysilicon 632 -303 632 -303 0 1
rlabel polysilicon 632 -309 632 -309 0 3
rlabel polysilicon 639 -303 639 -303 0 1
rlabel polysilicon 639 -309 639 -309 0 3
rlabel polysilicon 646 -303 646 -303 0 1
rlabel polysilicon 646 -309 646 -309 0 3
rlabel polysilicon 653 -303 653 -303 0 1
rlabel polysilicon 653 -309 653 -309 0 3
rlabel polysilicon 660 -303 660 -303 0 1
rlabel polysilicon 660 -309 660 -309 0 3
rlabel polysilicon 667 -303 667 -303 0 1
rlabel polysilicon 667 -309 667 -309 0 3
rlabel polysilicon 677 -309 677 -309 0 4
rlabel polysilicon 681 -303 681 -303 0 1
rlabel polysilicon 681 -309 681 -309 0 3
rlabel polysilicon 688 -303 688 -303 0 1
rlabel polysilicon 688 -309 688 -309 0 3
rlabel polysilicon 695 -303 695 -303 0 1
rlabel polysilicon 695 -309 695 -309 0 3
rlabel polysilicon 702 -303 702 -303 0 1
rlabel polysilicon 702 -309 702 -309 0 3
rlabel polysilicon 709 -303 709 -303 0 1
rlabel polysilicon 709 -309 709 -309 0 3
rlabel polysilicon 716 -303 716 -303 0 1
rlabel polysilicon 716 -309 716 -309 0 3
rlabel polysilicon 723 -303 723 -303 0 1
rlabel polysilicon 726 -309 726 -309 0 4
rlabel polysilicon 730 -303 730 -303 0 1
rlabel polysilicon 730 -309 730 -309 0 3
rlabel polysilicon 737 -303 737 -303 0 1
rlabel polysilicon 737 -309 737 -309 0 3
rlabel polysilicon 744 -303 744 -303 0 1
rlabel polysilicon 744 -309 744 -309 0 3
rlabel polysilicon 751 -303 751 -303 0 1
rlabel polysilicon 751 -309 751 -309 0 3
rlabel polysilicon 828 -303 828 -303 0 1
rlabel polysilicon 828 -309 828 -309 0 3
rlabel polysilicon 856 -303 856 -303 0 1
rlabel polysilicon 856 -309 856 -309 0 3
rlabel polysilicon 2 -374 2 -374 0 1
rlabel polysilicon 2 -380 2 -380 0 3
rlabel polysilicon 9 -374 9 -374 0 1
rlabel polysilicon 9 -380 9 -380 0 3
rlabel polysilicon 16 -374 16 -374 0 1
rlabel polysilicon 16 -380 16 -380 0 3
rlabel polysilicon 23 -374 23 -374 0 1
rlabel polysilicon 23 -380 23 -380 0 3
rlabel polysilicon 30 -374 30 -374 0 1
rlabel polysilicon 30 -380 30 -380 0 3
rlabel polysilicon 37 -374 37 -374 0 1
rlabel polysilicon 37 -380 37 -380 0 3
rlabel polysilicon 44 -374 44 -374 0 1
rlabel polysilicon 44 -380 44 -380 0 3
rlabel polysilicon 51 -374 51 -374 0 1
rlabel polysilicon 51 -380 51 -380 0 3
rlabel polysilicon 58 -374 58 -374 0 1
rlabel polysilicon 58 -380 58 -380 0 3
rlabel polysilicon 65 -374 65 -374 0 1
rlabel polysilicon 65 -380 65 -380 0 3
rlabel polysilicon 75 -374 75 -374 0 2
rlabel polysilicon 72 -380 72 -380 0 3
rlabel polysilicon 75 -380 75 -380 0 4
rlabel polysilicon 79 -374 79 -374 0 1
rlabel polysilicon 79 -380 79 -380 0 3
rlabel polysilicon 86 -374 86 -374 0 1
rlabel polysilicon 86 -380 86 -380 0 3
rlabel polysilicon 93 -374 93 -374 0 1
rlabel polysilicon 96 -374 96 -374 0 2
rlabel polysilicon 96 -380 96 -380 0 4
rlabel polysilicon 100 -374 100 -374 0 1
rlabel polysilicon 100 -380 100 -380 0 3
rlabel polysilicon 107 -374 107 -374 0 1
rlabel polysilicon 107 -380 107 -380 0 3
rlabel polysilicon 114 -374 114 -374 0 1
rlabel polysilicon 114 -380 114 -380 0 3
rlabel polysilicon 121 -374 121 -374 0 1
rlabel polysilicon 121 -380 121 -380 0 3
rlabel polysilicon 128 -374 128 -374 0 1
rlabel polysilicon 131 -374 131 -374 0 2
rlabel polysilicon 128 -380 128 -380 0 3
rlabel polysilicon 131 -380 131 -380 0 4
rlabel polysilicon 135 -374 135 -374 0 1
rlabel polysilicon 135 -380 135 -380 0 3
rlabel polysilicon 142 -374 142 -374 0 1
rlabel polysilicon 145 -374 145 -374 0 2
rlabel polysilicon 142 -380 142 -380 0 3
rlabel polysilicon 145 -380 145 -380 0 4
rlabel polysilicon 152 -374 152 -374 0 2
rlabel polysilicon 149 -380 149 -380 0 3
rlabel polysilicon 152 -380 152 -380 0 4
rlabel polysilicon 156 -374 156 -374 0 1
rlabel polysilicon 156 -380 156 -380 0 3
rlabel polysilicon 163 -374 163 -374 0 1
rlabel polysilicon 163 -380 163 -380 0 3
rlabel polysilicon 170 -374 170 -374 0 1
rlabel polysilicon 170 -380 170 -380 0 3
rlabel polysilicon 177 -374 177 -374 0 1
rlabel polysilicon 177 -380 177 -380 0 3
rlabel polysilicon 184 -374 184 -374 0 1
rlabel polysilicon 184 -380 184 -380 0 3
rlabel polysilicon 191 -374 191 -374 0 1
rlabel polysilicon 191 -380 191 -380 0 3
rlabel polysilicon 198 -380 198 -380 0 3
rlabel polysilicon 201 -380 201 -380 0 4
rlabel polysilicon 205 -374 205 -374 0 1
rlabel polysilicon 205 -380 205 -380 0 3
rlabel polysilicon 215 -374 215 -374 0 2
rlabel polysilicon 212 -380 212 -380 0 3
rlabel polysilicon 219 -374 219 -374 0 1
rlabel polysilicon 219 -380 219 -380 0 3
rlabel polysilicon 226 -374 226 -374 0 1
rlabel polysilicon 226 -380 226 -380 0 3
rlabel polysilicon 233 -374 233 -374 0 1
rlabel polysilicon 233 -380 233 -380 0 3
rlabel polysilicon 240 -374 240 -374 0 1
rlabel polysilicon 240 -380 240 -380 0 3
rlabel polysilicon 247 -374 247 -374 0 1
rlabel polysilicon 247 -380 247 -380 0 3
rlabel polysilicon 254 -374 254 -374 0 1
rlabel polysilicon 254 -380 254 -380 0 3
rlabel polysilicon 261 -374 261 -374 0 1
rlabel polysilicon 261 -380 261 -380 0 3
rlabel polysilicon 268 -374 268 -374 0 1
rlabel polysilicon 268 -380 268 -380 0 3
rlabel polysilicon 275 -374 275 -374 0 1
rlabel polysilicon 278 -380 278 -380 0 4
rlabel polysilicon 282 -374 282 -374 0 1
rlabel polysilicon 282 -380 282 -380 0 3
rlabel polysilicon 289 -374 289 -374 0 1
rlabel polysilicon 289 -380 289 -380 0 3
rlabel polysilicon 296 -374 296 -374 0 1
rlabel polysilicon 296 -380 296 -380 0 3
rlabel polysilicon 303 -374 303 -374 0 1
rlabel polysilicon 303 -380 303 -380 0 3
rlabel polysilicon 310 -374 310 -374 0 1
rlabel polysilicon 310 -380 310 -380 0 3
rlabel polysilicon 317 -374 317 -374 0 1
rlabel polysilicon 317 -380 317 -380 0 3
rlabel polysilicon 324 -374 324 -374 0 1
rlabel polysilicon 327 -374 327 -374 0 2
rlabel polysilicon 331 -374 331 -374 0 1
rlabel polysilicon 334 -374 334 -374 0 2
rlabel polysilicon 331 -380 331 -380 0 3
rlabel polysilicon 334 -380 334 -380 0 4
rlabel polysilicon 338 -374 338 -374 0 1
rlabel polysilicon 338 -380 338 -380 0 3
rlabel polysilicon 345 -374 345 -374 0 1
rlabel polysilicon 345 -380 345 -380 0 3
rlabel polysilicon 352 -374 352 -374 0 1
rlabel polysilicon 352 -380 352 -380 0 3
rlabel polysilicon 359 -374 359 -374 0 1
rlabel polysilicon 362 -374 362 -374 0 2
rlabel polysilicon 359 -380 359 -380 0 3
rlabel polysilicon 362 -380 362 -380 0 4
rlabel polysilicon 366 -374 366 -374 0 1
rlabel polysilicon 369 -374 369 -374 0 2
rlabel polysilicon 366 -380 366 -380 0 3
rlabel polysilicon 369 -380 369 -380 0 4
rlabel polysilicon 373 -374 373 -374 0 1
rlabel polysilicon 373 -380 373 -380 0 3
rlabel polysilicon 376 -380 376 -380 0 4
rlabel polysilicon 380 -374 380 -374 0 1
rlabel polysilicon 380 -380 380 -380 0 3
rlabel polysilicon 387 -374 387 -374 0 1
rlabel polysilicon 387 -380 387 -380 0 3
rlabel polysilicon 394 -374 394 -374 0 1
rlabel polysilicon 394 -380 394 -380 0 3
rlabel polysilicon 401 -374 401 -374 0 1
rlabel polysilicon 404 -374 404 -374 0 2
rlabel polysilicon 401 -380 401 -380 0 3
rlabel polysilicon 404 -380 404 -380 0 4
rlabel polysilicon 408 -374 408 -374 0 1
rlabel polysilicon 408 -380 408 -380 0 3
rlabel polysilicon 415 -374 415 -374 0 1
rlabel polysilicon 415 -380 415 -380 0 3
rlabel polysilicon 422 -374 422 -374 0 1
rlabel polysilicon 425 -374 425 -374 0 2
rlabel polysilicon 422 -380 422 -380 0 3
rlabel polysilicon 425 -380 425 -380 0 4
rlabel polysilicon 429 -374 429 -374 0 1
rlabel polysilicon 432 -374 432 -374 0 2
rlabel polysilicon 429 -380 429 -380 0 3
rlabel polysilicon 432 -380 432 -380 0 4
rlabel polysilicon 436 -374 436 -374 0 1
rlabel polysilicon 436 -380 436 -380 0 3
rlabel polysilicon 443 -374 443 -374 0 1
rlabel polysilicon 443 -380 443 -380 0 3
rlabel polysilicon 450 -374 450 -374 0 1
rlabel polysilicon 453 -374 453 -374 0 2
rlabel polysilicon 450 -380 450 -380 0 3
rlabel polysilicon 457 -374 457 -374 0 1
rlabel polysilicon 457 -380 457 -380 0 3
rlabel polysilicon 464 -374 464 -374 0 1
rlabel polysilicon 464 -380 464 -380 0 3
rlabel polysilicon 471 -374 471 -374 0 1
rlabel polysilicon 474 -374 474 -374 0 2
rlabel polysilicon 471 -380 471 -380 0 3
rlabel polysilicon 478 -374 478 -374 0 1
rlabel polysilicon 478 -380 478 -380 0 3
rlabel polysilicon 485 -374 485 -374 0 1
rlabel polysilicon 485 -380 485 -380 0 3
rlabel polysilicon 495 -374 495 -374 0 2
rlabel polysilicon 495 -380 495 -380 0 4
rlabel polysilicon 499 -374 499 -374 0 1
rlabel polysilicon 499 -380 499 -380 0 3
rlabel polysilicon 506 -380 506 -380 0 3
rlabel polysilicon 509 -380 509 -380 0 4
rlabel polysilicon 513 -374 513 -374 0 1
rlabel polysilicon 516 -374 516 -374 0 2
rlabel polysilicon 513 -380 513 -380 0 3
rlabel polysilicon 516 -380 516 -380 0 4
rlabel polysilicon 520 -374 520 -374 0 1
rlabel polysilicon 520 -380 520 -380 0 3
rlabel polysilicon 527 -374 527 -374 0 1
rlabel polysilicon 527 -380 527 -380 0 3
rlabel polysilicon 534 -374 534 -374 0 1
rlabel polysilicon 534 -380 534 -380 0 3
rlabel polysilicon 541 -374 541 -374 0 1
rlabel polysilicon 541 -380 541 -380 0 3
rlabel polysilicon 548 -374 548 -374 0 1
rlabel polysilicon 548 -380 548 -380 0 3
rlabel polysilicon 555 -374 555 -374 0 1
rlabel polysilicon 555 -380 555 -380 0 3
rlabel polysilicon 562 -374 562 -374 0 1
rlabel polysilicon 562 -380 562 -380 0 3
rlabel polysilicon 569 -374 569 -374 0 1
rlabel polysilicon 569 -380 569 -380 0 3
rlabel polysilicon 576 -374 576 -374 0 1
rlabel polysilicon 576 -380 576 -380 0 3
rlabel polysilicon 583 -374 583 -374 0 1
rlabel polysilicon 586 -374 586 -374 0 2
rlabel polysilicon 590 -374 590 -374 0 1
rlabel polysilicon 590 -380 590 -380 0 3
rlabel polysilicon 597 -374 597 -374 0 1
rlabel polysilicon 597 -380 597 -380 0 3
rlabel polysilicon 604 -374 604 -374 0 1
rlabel polysilicon 604 -380 604 -380 0 3
rlabel polysilicon 611 -374 611 -374 0 1
rlabel polysilicon 611 -380 611 -380 0 3
rlabel polysilicon 618 -374 618 -374 0 1
rlabel polysilicon 618 -380 618 -380 0 3
rlabel polysilicon 625 -374 625 -374 0 1
rlabel polysilicon 625 -380 625 -380 0 3
rlabel polysilicon 632 -374 632 -374 0 1
rlabel polysilicon 632 -380 632 -380 0 3
rlabel polysilicon 639 -374 639 -374 0 1
rlabel polysilicon 639 -380 639 -380 0 3
rlabel polysilicon 646 -374 646 -374 0 1
rlabel polysilicon 646 -380 646 -380 0 3
rlabel polysilicon 653 -374 653 -374 0 1
rlabel polysilicon 653 -380 653 -380 0 3
rlabel polysilicon 660 -374 660 -374 0 1
rlabel polysilicon 660 -380 660 -380 0 3
rlabel polysilicon 667 -374 667 -374 0 1
rlabel polysilicon 667 -380 667 -380 0 3
rlabel polysilicon 674 -374 674 -374 0 1
rlabel polysilicon 674 -380 674 -380 0 3
rlabel polysilicon 681 -374 681 -374 0 1
rlabel polysilicon 681 -380 681 -380 0 3
rlabel polysilicon 688 -374 688 -374 0 1
rlabel polysilicon 688 -380 688 -380 0 3
rlabel polysilicon 695 -374 695 -374 0 1
rlabel polysilicon 695 -380 695 -380 0 3
rlabel polysilicon 702 -374 702 -374 0 1
rlabel polysilicon 702 -380 702 -380 0 3
rlabel polysilicon 709 -374 709 -374 0 1
rlabel polysilicon 709 -380 709 -380 0 3
rlabel polysilicon 716 -374 716 -374 0 1
rlabel polysilicon 716 -380 716 -380 0 3
rlabel polysilicon 723 -374 723 -374 0 1
rlabel polysilicon 723 -380 723 -380 0 3
rlabel polysilicon 730 -374 730 -374 0 1
rlabel polysilicon 730 -380 730 -380 0 3
rlabel polysilicon 737 -374 737 -374 0 1
rlabel polysilicon 737 -380 737 -380 0 3
rlabel polysilicon 744 -374 744 -374 0 1
rlabel polysilicon 744 -380 744 -380 0 3
rlabel polysilicon 751 -374 751 -374 0 1
rlabel polysilicon 751 -380 751 -380 0 3
rlabel polysilicon 758 -374 758 -374 0 1
rlabel polysilicon 758 -380 758 -380 0 3
rlabel polysilicon 765 -374 765 -374 0 1
rlabel polysilicon 765 -380 765 -380 0 3
rlabel polysilicon 772 -374 772 -374 0 1
rlabel polysilicon 772 -380 772 -380 0 3
rlabel polysilicon 779 -374 779 -374 0 1
rlabel polysilicon 779 -380 779 -380 0 3
rlabel polysilicon 786 -374 786 -374 0 1
rlabel polysilicon 786 -380 786 -380 0 3
rlabel polysilicon 793 -374 793 -374 0 1
rlabel polysilicon 793 -380 793 -380 0 3
rlabel polysilicon 800 -374 800 -374 0 1
rlabel polysilicon 800 -380 800 -380 0 3
rlabel polysilicon 807 -374 807 -374 0 1
rlabel polysilicon 807 -380 807 -380 0 3
rlabel polysilicon 814 -374 814 -374 0 1
rlabel polysilicon 814 -380 814 -380 0 3
rlabel polysilicon 821 -374 821 -374 0 1
rlabel polysilicon 821 -380 821 -380 0 3
rlabel polysilicon 828 -374 828 -374 0 1
rlabel polysilicon 828 -380 828 -380 0 3
rlabel polysilicon 835 -374 835 -374 0 1
rlabel polysilicon 835 -380 835 -380 0 3
rlabel polysilicon 842 -374 842 -374 0 1
rlabel polysilicon 842 -380 842 -380 0 3
rlabel polysilicon 849 -374 849 -374 0 1
rlabel polysilicon 852 -374 852 -374 0 2
rlabel polysilicon 849 -380 849 -380 0 3
rlabel polysilicon 852 -380 852 -380 0 4
rlabel polysilicon 856 -374 856 -374 0 1
rlabel polysilicon 856 -380 856 -380 0 3
rlabel polysilicon 863 -374 863 -374 0 1
rlabel polysilicon 863 -380 863 -380 0 3
rlabel polysilicon 870 -374 870 -374 0 1
rlabel polysilicon 870 -380 870 -380 0 3
rlabel polysilicon 877 -374 877 -374 0 1
rlabel polysilicon 884 -380 884 -380 0 3
rlabel polysilicon 891 -374 891 -374 0 1
rlabel polysilicon 891 -380 891 -380 0 3
rlabel polysilicon 2 -463 2 -463 0 1
rlabel polysilicon 2 -469 2 -469 0 3
rlabel polysilicon 9 -463 9 -463 0 1
rlabel polysilicon 9 -469 9 -469 0 3
rlabel polysilicon 16 -463 16 -463 0 1
rlabel polysilicon 16 -469 16 -469 0 3
rlabel polysilicon 23 -463 23 -463 0 1
rlabel polysilicon 23 -469 23 -469 0 3
rlabel polysilicon 30 -463 30 -463 0 1
rlabel polysilicon 30 -469 30 -469 0 3
rlabel polysilicon 37 -463 37 -463 0 1
rlabel polysilicon 37 -469 37 -469 0 3
rlabel polysilicon 44 -463 44 -463 0 1
rlabel polysilicon 54 -463 54 -463 0 2
rlabel polysilicon 51 -469 51 -469 0 3
rlabel polysilicon 54 -469 54 -469 0 4
rlabel polysilicon 58 -463 58 -463 0 1
rlabel polysilicon 58 -469 58 -469 0 3
rlabel polysilicon 65 -463 65 -463 0 1
rlabel polysilicon 65 -469 65 -469 0 3
rlabel polysilicon 72 -463 72 -463 0 1
rlabel polysilicon 72 -469 72 -469 0 3
rlabel polysilicon 79 -463 79 -463 0 1
rlabel polysilicon 79 -469 79 -469 0 3
rlabel polysilicon 82 -469 82 -469 0 4
rlabel polysilicon 86 -463 86 -463 0 1
rlabel polysilicon 86 -469 86 -469 0 3
rlabel polysilicon 93 -463 93 -463 0 1
rlabel polysilicon 93 -469 93 -469 0 3
rlabel polysilicon 103 -463 103 -463 0 2
rlabel polysilicon 100 -469 100 -469 0 3
rlabel polysilicon 107 -463 107 -463 0 1
rlabel polysilicon 110 -463 110 -463 0 2
rlabel polysilicon 107 -469 107 -469 0 3
rlabel polysilicon 114 -463 114 -463 0 1
rlabel polysilicon 117 -463 117 -463 0 2
rlabel polysilicon 117 -469 117 -469 0 4
rlabel polysilicon 121 -463 121 -463 0 1
rlabel polysilicon 121 -469 121 -469 0 3
rlabel polysilicon 128 -463 128 -463 0 1
rlabel polysilicon 128 -469 128 -469 0 3
rlabel polysilicon 135 -463 135 -463 0 1
rlabel polysilicon 135 -469 135 -469 0 3
rlabel polysilicon 142 -463 142 -463 0 1
rlabel polysilicon 142 -469 142 -469 0 3
rlabel polysilicon 149 -463 149 -463 0 1
rlabel polysilicon 149 -469 149 -469 0 3
rlabel polysilicon 156 -463 156 -463 0 1
rlabel polysilicon 159 -463 159 -463 0 2
rlabel polysilicon 163 -463 163 -463 0 1
rlabel polysilicon 163 -469 163 -469 0 3
rlabel polysilicon 166 -469 166 -469 0 4
rlabel polysilicon 170 -463 170 -463 0 1
rlabel polysilicon 170 -469 170 -469 0 3
rlabel polysilicon 177 -463 177 -463 0 1
rlabel polysilicon 177 -469 177 -469 0 3
rlabel polysilicon 184 -463 184 -463 0 1
rlabel polysilicon 184 -469 184 -469 0 3
rlabel polysilicon 191 -463 191 -463 0 1
rlabel polysilicon 191 -469 191 -469 0 3
rlabel polysilicon 194 -469 194 -469 0 4
rlabel polysilicon 198 -463 198 -463 0 1
rlabel polysilicon 198 -469 198 -469 0 3
rlabel polysilicon 201 -469 201 -469 0 4
rlabel polysilicon 205 -463 205 -463 0 1
rlabel polysilicon 205 -469 205 -469 0 3
rlabel polysilicon 212 -463 212 -463 0 1
rlabel polysilicon 215 -463 215 -463 0 2
rlabel polysilicon 212 -469 212 -469 0 3
rlabel polysilicon 222 -463 222 -463 0 2
rlabel polysilicon 219 -469 219 -469 0 3
rlabel polysilicon 226 -463 226 -463 0 1
rlabel polysilicon 226 -469 226 -469 0 3
rlabel polysilicon 233 -463 233 -463 0 1
rlabel polysilicon 233 -469 233 -469 0 3
rlabel polysilicon 240 -463 240 -463 0 1
rlabel polysilicon 243 -463 243 -463 0 2
rlabel polysilicon 240 -469 240 -469 0 3
rlabel polysilicon 243 -469 243 -469 0 4
rlabel polysilicon 247 -463 247 -463 0 1
rlabel polysilicon 247 -469 247 -469 0 3
rlabel polysilicon 254 -463 254 -463 0 1
rlabel polysilicon 254 -469 254 -469 0 3
rlabel polysilicon 261 -463 261 -463 0 1
rlabel polysilicon 261 -469 261 -469 0 3
rlabel polysilicon 268 -463 268 -463 0 1
rlabel polysilicon 268 -469 268 -469 0 3
rlabel polysilicon 275 -463 275 -463 0 1
rlabel polysilicon 275 -469 275 -469 0 3
rlabel polysilicon 282 -463 282 -463 0 1
rlabel polysilicon 282 -469 282 -469 0 3
rlabel polysilicon 289 -463 289 -463 0 1
rlabel polysilicon 289 -469 289 -469 0 3
rlabel polysilicon 296 -463 296 -463 0 1
rlabel polysilicon 299 -463 299 -463 0 2
rlabel polysilicon 296 -469 296 -469 0 3
rlabel polysilicon 303 -463 303 -463 0 1
rlabel polysilicon 306 -463 306 -463 0 2
rlabel polysilicon 303 -469 303 -469 0 3
rlabel polysilicon 306 -469 306 -469 0 4
rlabel polysilicon 310 -463 310 -463 0 1
rlabel polysilicon 310 -469 310 -469 0 3
rlabel polysilicon 317 -463 317 -463 0 1
rlabel polysilicon 317 -469 317 -469 0 3
rlabel polysilicon 324 -463 324 -463 0 1
rlabel polysilicon 324 -469 324 -469 0 3
rlabel polysilicon 331 -463 331 -463 0 1
rlabel polysilicon 331 -469 331 -469 0 3
rlabel polysilicon 338 -463 338 -463 0 1
rlabel polysilicon 338 -469 338 -469 0 3
rlabel polysilicon 348 -463 348 -463 0 2
rlabel polysilicon 345 -469 345 -469 0 3
rlabel polysilicon 348 -469 348 -469 0 4
rlabel polysilicon 352 -463 352 -463 0 1
rlabel polysilicon 352 -469 352 -469 0 3
rlabel polysilicon 359 -463 359 -463 0 1
rlabel polysilicon 359 -469 359 -469 0 3
rlabel polysilicon 366 -463 366 -463 0 1
rlabel polysilicon 369 -463 369 -463 0 2
rlabel polysilicon 366 -469 366 -469 0 3
rlabel polysilicon 369 -469 369 -469 0 4
rlabel polysilicon 373 -463 373 -463 0 1
rlabel polysilicon 373 -469 373 -469 0 3
rlabel polysilicon 383 -463 383 -463 0 2
rlabel polysilicon 380 -469 380 -469 0 3
rlabel polysilicon 383 -469 383 -469 0 4
rlabel polysilicon 387 -463 387 -463 0 1
rlabel polysilicon 390 -463 390 -463 0 2
rlabel polysilicon 387 -469 387 -469 0 3
rlabel polysilicon 394 -463 394 -463 0 1
rlabel polysilicon 394 -469 394 -469 0 3
rlabel polysilicon 401 -463 401 -463 0 1
rlabel polysilicon 401 -469 401 -469 0 3
rlabel polysilicon 408 -463 408 -463 0 1
rlabel polysilicon 408 -469 408 -469 0 3
rlabel polysilicon 415 -463 415 -463 0 1
rlabel polysilicon 418 -463 418 -463 0 2
rlabel polysilicon 415 -469 415 -469 0 3
rlabel polysilicon 418 -469 418 -469 0 4
rlabel polysilicon 422 -463 422 -463 0 1
rlabel polysilicon 422 -469 422 -469 0 3
rlabel polysilicon 429 -463 429 -463 0 1
rlabel polysilicon 432 -463 432 -463 0 2
rlabel polysilicon 429 -469 429 -469 0 3
rlabel polysilicon 432 -469 432 -469 0 4
rlabel polysilicon 436 -463 436 -463 0 1
rlabel polysilicon 436 -469 436 -469 0 3
rlabel polysilicon 439 -469 439 -469 0 4
rlabel polysilicon 443 -463 443 -463 0 1
rlabel polysilicon 443 -469 443 -469 0 3
rlabel polysilicon 450 -463 450 -463 0 1
rlabel polysilicon 450 -469 450 -469 0 3
rlabel polysilicon 457 -463 457 -463 0 1
rlabel polysilicon 457 -469 457 -469 0 3
rlabel polysilicon 460 -469 460 -469 0 4
rlabel polysilicon 464 -463 464 -463 0 1
rlabel polysilicon 464 -469 464 -469 0 3
rlabel polysilicon 471 -463 471 -463 0 1
rlabel polysilicon 471 -469 471 -469 0 3
rlabel polysilicon 478 -463 478 -463 0 1
rlabel polysilicon 478 -469 478 -469 0 3
rlabel polysilicon 485 -463 485 -463 0 1
rlabel polysilicon 485 -469 485 -469 0 3
rlabel polysilicon 488 -469 488 -469 0 4
rlabel polysilicon 492 -463 492 -463 0 1
rlabel polysilicon 492 -469 492 -469 0 3
rlabel polysilicon 499 -463 499 -463 0 1
rlabel polysilicon 502 -463 502 -463 0 2
rlabel polysilicon 499 -469 499 -469 0 3
rlabel polysilicon 509 -463 509 -463 0 2
rlabel polysilicon 506 -469 506 -469 0 3
rlabel polysilicon 513 -463 513 -463 0 1
rlabel polysilicon 513 -469 513 -469 0 3
rlabel polysilicon 520 -463 520 -463 0 1
rlabel polysilicon 523 -463 523 -463 0 2
rlabel polysilicon 520 -469 520 -469 0 3
rlabel polysilicon 523 -469 523 -469 0 4
rlabel polysilicon 527 -463 527 -463 0 1
rlabel polysilicon 527 -469 527 -469 0 3
rlabel polysilicon 534 -463 534 -463 0 1
rlabel polysilicon 534 -469 534 -469 0 3
rlabel polysilicon 541 -463 541 -463 0 1
rlabel polysilicon 541 -469 541 -469 0 3
rlabel polysilicon 548 -463 548 -463 0 1
rlabel polysilicon 548 -469 548 -469 0 3
rlabel polysilicon 555 -463 555 -463 0 1
rlabel polysilicon 555 -469 555 -469 0 3
rlabel polysilicon 562 -463 562 -463 0 1
rlabel polysilicon 562 -469 562 -469 0 3
rlabel polysilicon 569 -463 569 -463 0 1
rlabel polysilicon 569 -469 569 -469 0 3
rlabel polysilicon 576 -463 576 -463 0 1
rlabel polysilicon 576 -469 576 -469 0 3
rlabel polysilicon 583 -463 583 -463 0 1
rlabel polysilicon 583 -469 583 -469 0 3
rlabel polysilicon 590 -463 590 -463 0 1
rlabel polysilicon 590 -469 590 -469 0 3
rlabel polysilicon 597 -463 597 -463 0 1
rlabel polysilicon 597 -469 597 -469 0 3
rlabel polysilicon 604 -463 604 -463 0 1
rlabel polysilicon 604 -469 604 -469 0 3
rlabel polysilicon 611 -463 611 -463 0 1
rlabel polysilicon 611 -469 611 -469 0 3
rlabel polysilicon 618 -463 618 -463 0 1
rlabel polysilicon 621 -463 621 -463 0 2
rlabel polysilicon 625 -463 625 -463 0 1
rlabel polysilicon 625 -469 625 -469 0 3
rlabel polysilicon 632 -463 632 -463 0 1
rlabel polysilicon 632 -469 632 -469 0 3
rlabel polysilicon 639 -463 639 -463 0 1
rlabel polysilicon 639 -469 639 -469 0 3
rlabel polysilicon 646 -463 646 -463 0 1
rlabel polysilicon 646 -469 646 -469 0 3
rlabel polysilicon 653 -463 653 -463 0 1
rlabel polysilicon 653 -469 653 -469 0 3
rlabel polysilicon 660 -463 660 -463 0 1
rlabel polysilicon 660 -469 660 -469 0 3
rlabel polysilicon 667 -463 667 -463 0 1
rlabel polysilicon 667 -469 667 -469 0 3
rlabel polysilicon 674 -463 674 -463 0 1
rlabel polysilicon 674 -469 674 -469 0 3
rlabel polysilicon 681 -463 681 -463 0 1
rlabel polysilicon 681 -469 681 -469 0 3
rlabel polysilicon 688 -463 688 -463 0 1
rlabel polysilicon 688 -469 688 -469 0 3
rlabel polysilicon 695 -463 695 -463 0 1
rlabel polysilicon 695 -469 695 -469 0 3
rlabel polysilicon 702 -463 702 -463 0 1
rlabel polysilicon 702 -469 702 -469 0 3
rlabel polysilicon 709 -463 709 -463 0 1
rlabel polysilicon 709 -469 709 -469 0 3
rlabel polysilicon 716 -463 716 -463 0 1
rlabel polysilicon 716 -469 716 -469 0 3
rlabel polysilicon 723 -463 723 -463 0 1
rlabel polysilicon 723 -469 723 -469 0 3
rlabel polysilicon 730 -463 730 -463 0 1
rlabel polysilicon 730 -469 730 -469 0 3
rlabel polysilicon 737 -463 737 -463 0 1
rlabel polysilicon 737 -469 737 -469 0 3
rlabel polysilicon 744 -463 744 -463 0 1
rlabel polysilicon 744 -469 744 -469 0 3
rlabel polysilicon 751 -463 751 -463 0 1
rlabel polysilicon 751 -469 751 -469 0 3
rlabel polysilicon 758 -463 758 -463 0 1
rlabel polysilicon 758 -469 758 -469 0 3
rlabel polysilicon 765 -463 765 -463 0 1
rlabel polysilicon 765 -469 765 -469 0 3
rlabel polysilicon 772 -463 772 -463 0 1
rlabel polysilicon 772 -469 772 -469 0 3
rlabel polysilicon 779 -463 779 -463 0 1
rlabel polysilicon 779 -469 779 -469 0 3
rlabel polysilicon 786 -463 786 -463 0 1
rlabel polysilicon 786 -469 786 -469 0 3
rlabel polysilicon 793 -463 793 -463 0 1
rlabel polysilicon 793 -469 793 -469 0 3
rlabel polysilicon 800 -463 800 -463 0 1
rlabel polysilicon 800 -469 800 -469 0 3
rlabel polysilicon 807 -463 807 -463 0 1
rlabel polysilicon 807 -469 807 -469 0 3
rlabel polysilicon 814 -463 814 -463 0 1
rlabel polysilicon 814 -469 814 -469 0 3
rlabel polysilicon 821 -463 821 -463 0 1
rlabel polysilicon 821 -469 821 -469 0 3
rlabel polysilicon 828 -463 828 -463 0 1
rlabel polysilicon 828 -469 828 -469 0 3
rlabel polysilicon 835 -463 835 -463 0 1
rlabel polysilicon 835 -469 835 -469 0 3
rlabel polysilicon 842 -463 842 -463 0 1
rlabel polysilicon 842 -469 842 -469 0 3
rlabel polysilicon 849 -463 849 -463 0 1
rlabel polysilicon 849 -469 849 -469 0 3
rlabel polysilicon 856 -463 856 -463 0 1
rlabel polysilicon 856 -469 856 -469 0 3
rlabel polysilicon 863 -463 863 -463 0 1
rlabel polysilicon 863 -469 863 -469 0 3
rlabel polysilicon 870 -463 870 -463 0 1
rlabel polysilicon 870 -469 870 -469 0 3
rlabel polysilicon 877 -463 877 -463 0 1
rlabel polysilicon 877 -469 877 -469 0 3
rlabel polysilicon 884 -463 884 -463 0 1
rlabel polysilicon 884 -469 884 -469 0 3
rlabel polysilicon 891 -463 891 -463 0 1
rlabel polysilicon 891 -469 891 -469 0 3
rlabel polysilicon 898 -463 898 -463 0 1
rlabel polysilicon 898 -469 898 -469 0 3
rlabel polysilicon 905 -463 905 -463 0 1
rlabel polysilicon 905 -469 905 -469 0 3
rlabel polysilicon 912 -463 912 -463 0 1
rlabel polysilicon 912 -469 912 -469 0 3
rlabel polysilicon 919 -463 919 -463 0 1
rlabel polysilicon 919 -469 919 -469 0 3
rlabel polysilicon 926 -463 926 -463 0 1
rlabel polysilicon 926 -469 926 -469 0 3
rlabel polysilicon 933 -463 933 -463 0 1
rlabel polysilicon 933 -469 933 -469 0 3
rlabel polysilicon 940 -463 940 -463 0 1
rlabel polysilicon 940 -469 940 -469 0 3
rlabel polysilicon 947 -463 947 -463 0 1
rlabel polysilicon 947 -469 947 -469 0 3
rlabel polysilicon 2 -550 2 -550 0 1
rlabel polysilicon 2 -556 2 -556 0 3
rlabel polysilicon 9 -550 9 -550 0 1
rlabel polysilicon 9 -556 9 -556 0 3
rlabel polysilicon 16 -550 16 -550 0 1
rlabel polysilicon 16 -556 16 -556 0 3
rlabel polysilicon 23 -556 23 -556 0 3
rlabel polysilicon 30 -550 30 -550 0 1
rlabel polysilicon 30 -556 30 -556 0 3
rlabel polysilicon 37 -550 37 -550 0 1
rlabel polysilicon 37 -556 37 -556 0 3
rlabel polysilicon 44 -550 44 -550 0 1
rlabel polysilicon 51 -550 51 -550 0 1
rlabel polysilicon 51 -556 51 -556 0 3
rlabel polysilicon 58 -550 58 -550 0 1
rlabel polysilicon 58 -556 58 -556 0 3
rlabel polysilicon 65 -550 65 -550 0 1
rlabel polysilicon 65 -556 65 -556 0 3
rlabel polysilicon 72 -550 72 -550 0 1
rlabel polysilicon 72 -556 72 -556 0 3
rlabel polysilicon 79 -550 79 -550 0 1
rlabel polysilicon 79 -556 79 -556 0 3
rlabel polysilicon 86 -550 86 -550 0 1
rlabel polysilicon 86 -556 86 -556 0 3
rlabel polysilicon 93 -550 93 -550 0 1
rlabel polysilicon 96 -550 96 -550 0 2
rlabel polysilicon 93 -556 93 -556 0 3
rlabel polysilicon 96 -556 96 -556 0 4
rlabel polysilicon 100 -550 100 -550 0 1
rlabel polysilicon 100 -556 100 -556 0 3
rlabel polysilicon 107 -550 107 -550 0 1
rlabel polysilicon 107 -556 107 -556 0 3
rlabel polysilicon 114 -550 114 -550 0 1
rlabel polysilicon 114 -556 114 -556 0 3
rlabel polysilicon 121 -550 121 -550 0 1
rlabel polysilicon 121 -556 121 -556 0 3
rlabel polysilicon 128 -550 128 -550 0 1
rlabel polysilicon 128 -556 128 -556 0 3
rlabel polysilicon 135 -550 135 -550 0 1
rlabel polysilicon 135 -556 135 -556 0 3
rlabel polysilicon 145 -550 145 -550 0 2
rlabel polysilicon 145 -556 145 -556 0 4
rlabel polysilicon 149 -550 149 -550 0 1
rlabel polysilicon 149 -556 149 -556 0 3
rlabel polysilicon 156 -550 156 -550 0 1
rlabel polysilicon 159 -556 159 -556 0 4
rlabel polysilicon 163 -550 163 -550 0 1
rlabel polysilicon 166 -550 166 -550 0 2
rlabel polysilicon 166 -556 166 -556 0 4
rlabel polysilicon 170 -550 170 -550 0 1
rlabel polysilicon 170 -556 170 -556 0 3
rlabel polysilicon 180 -550 180 -550 0 2
rlabel polysilicon 177 -556 177 -556 0 3
rlabel polysilicon 180 -556 180 -556 0 4
rlabel polysilicon 184 -550 184 -550 0 1
rlabel polysilicon 184 -556 184 -556 0 3
rlabel polysilicon 191 -550 191 -550 0 1
rlabel polysilicon 191 -556 191 -556 0 3
rlabel polysilicon 198 -550 198 -550 0 1
rlabel polysilicon 198 -556 198 -556 0 3
rlabel polysilicon 205 -550 205 -550 0 1
rlabel polysilicon 205 -556 205 -556 0 3
rlabel polysilicon 212 -556 212 -556 0 3
rlabel polysilicon 215 -556 215 -556 0 4
rlabel polysilicon 219 -550 219 -550 0 1
rlabel polysilicon 219 -556 219 -556 0 3
rlabel polysilicon 226 -550 226 -550 0 1
rlabel polysilicon 226 -556 226 -556 0 3
rlabel polysilicon 233 -550 233 -550 0 1
rlabel polysilicon 233 -556 233 -556 0 3
rlabel polysilicon 240 -550 240 -550 0 1
rlabel polysilicon 243 -550 243 -550 0 2
rlabel polysilicon 243 -556 243 -556 0 4
rlabel polysilicon 247 -550 247 -550 0 1
rlabel polysilicon 247 -556 247 -556 0 3
rlabel polysilicon 254 -550 254 -550 0 1
rlabel polysilicon 254 -556 254 -556 0 3
rlabel polysilicon 261 -550 261 -550 0 1
rlabel polysilicon 264 -550 264 -550 0 2
rlabel polysilicon 261 -556 261 -556 0 3
rlabel polysilicon 264 -556 264 -556 0 4
rlabel polysilicon 268 -550 268 -550 0 1
rlabel polysilicon 268 -556 268 -556 0 3
rlabel polysilicon 275 -550 275 -550 0 1
rlabel polysilicon 275 -556 275 -556 0 3
rlabel polysilicon 282 -550 282 -550 0 1
rlabel polysilicon 282 -556 282 -556 0 3
rlabel polysilicon 289 -550 289 -550 0 1
rlabel polysilicon 289 -556 289 -556 0 3
rlabel polysilicon 296 -550 296 -550 0 1
rlabel polysilicon 296 -556 296 -556 0 3
rlabel polysilicon 303 -550 303 -550 0 1
rlabel polysilicon 303 -556 303 -556 0 3
rlabel polysilicon 310 -550 310 -550 0 1
rlabel polysilicon 313 -550 313 -550 0 2
rlabel polysilicon 313 -556 313 -556 0 4
rlabel polysilicon 320 -550 320 -550 0 2
rlabel polysilicon 317 -556 317 -556 0 3
rlabel polysilicon 324 -550 324 -550 0 1
rlabel polysilicon 324 -556 324 -556 0 3
rlabel polysilicon 334 -550 334 -550 0 2
rlabel polysilicon 331 -556 331 -556 0 3
rlabel polysilicon 341 -550 341 -550 0 2
rlabel polysilicon 338 -556 338 -556 0 3
rlabel polysilicon 341 -556 341 -556 0 4
rlabel polysilicon 345 -550 345 -550 0 1
rlabel polysilicon 345 -556 345 -556 0 3
rlabel polysilicon 352 -550 352 -550 0 1
rlabel polysilicon 352 -556 352 -556 0 3
rlabel polysilicon 359 -556 359 -556 0 3
rlabel polysilicon 362 -556 362 -556 0 4
rlabel polysilicon 366 -550 366 -550 0 1
rlabel polysilicon 366 -556 366 -556 0 3
rlabel polysilicon 373 -550 373 -550 0 1
rlabel polysilicon 373 -556 373 -556 0 3
rlabel polysilicon 380 -550 380 -550 0 1
rlabel polysilicon 380 -556 380 -556 0 3
rlabel polysilicon 387 -550 387 -550 0 1
rlabel polysilicon 390 -550 390 -550 0 2
rlabel polysilicon 387 -556 387 -556 0 3
rlabel polysilicon 390 -556 390 -556 0 4
rlabel polysilicon 394 -550 394 -550 0 1
rlabel polysilicon 394 -556 394 -556 0 3
rlabel polysilicon 401 -550 401 -550 0 1
rlabel polysilicon 401 -556 401 -556 0 3
rlabel polysilicon 408 -550 408 -550 0 1
rlabel polysilicon 408 -556 408 -556 0 3
rlabel polysilicon 415 -550 415 -550 0 1
rlabel polysilicon 422 -550 422 -550 0 1
rlabel polysilicon 425 -550 425 -550 0 2
rlabel polysilicon 422 -556 422 -556 0 3
rlabel polysilicon 425 -556 425 -556 0 4
rlabel polysilicon 429 -550 429 -550 0 1
rlabel polysilicon 429 -556 429 -556 0 3
rlabel polysilicon 436 -550 436 -550 0 1
rlabel polysilicon 436 -556 436 -556 0 3
rlabel polysilicon 443 -550 443 -550 0 1
rlabel polysilicon 443 -556 443 -556 0 3
rlabel polysilicon 450 -550 450 -550 0 1
rlabel polysilicon 453 -550 453 -550 0 2
rlabel polysilicon 450 -556 450 -556 0 3
rlabel polysilicon 453 -556 453 -556 0 4
rlabel polysilicon 457 -550 457 -550 0 1
rlabel polysilicon 457 -556 457 -556 0 3
rlabel polysilicon 464 -550 464 -550 0 1
rlabel polysilicon 464 -556 464 -556 0 3
rlabel polysilicon 471 -550 471 -550 0 1
rlabel polysilicon 471 -556 471 -556 0 3
rlabel polysilicon 478 -550 478 -550 0 1
rlabel polysilicon 481 -550 481 -550 0 2
rlabel polysilicon 481 -556 481 -556 0 4
rlabel polysilicon 485 -550 485 -550 0 1
rlabel polysilicon 485 -556 485 -556 0 3
rlabel polysilicon 495 -550 495 -550 0 2
rlabel polysilicon 492 -556 492 -556 0 3
rlabel polysilicon 495 -556 495 -556 0 4
rlabel polysilicon 499 -550 499 -550 0 1
rlabel polysilicon 502 -550 502 -550 0 2
rlabel polysilicon 499 -556 499 -556 0 3
rlabel polysilicon 502 -556 502 -556 0 4
rlabel polysilicon 509 -550 509 -550 0 2
rlabel polysilicon 509 -556 509 -556 0 4
rlabel polysilicon 513 -550 513 -550 0 1
rlabel polysilicon 513 -556 513 -556 0 3
rlabel polysilicon 520 -550 520 -550 0 1
rlabel polysilicon 520 -556 520 -556 0 3
rlabel polysilicon 527 -550 527 -550 0 1
rlabel polysilicon 527 -556 527 -556 0 3
rlabel polysilicon 534 -550 534 -550 0 1
rlabel polysilicon 534 -556 534 -556 0 3
rlabel polysilicon 541 -550 541 -550 0 1
rlabel polysilicon 544 -550 544 -550 0 2
rlabel polysilicon 544 -556 544 -556 0 4
rlabel polysilicon 548 -550 548 -550 0 1
rlabel polysilicon 548 -556 548 -556 0 3
rlabel polysilicon 555 -550 555 -550 0 1
rlabel polysilicon 555 -556 555 -556 0 3
rlabel polysilicon 562 -550 562 -550 0 1
rlabel polysilicon 562 -556 562 -556 0 3
rlabel polysilicon 569 -550 569 -550 0 1
rlabel polysilicon 569 -556 569 -556 0 3
rlabel polysilicon 576 -550 576 -550 0 1
rlabel polysilicon 576 -556 576 -556 0 3
rlabel polysilicon 583 -550 583 -550 0 1
rlabel polysilicon 583 -556 583 -556 0 3
rlabel polysilicon 590 -550 590 -550 0 1
rlabel polysilicon 590 -556 590 -556 0 3
rlabel polysilicon 597 -550 597 -550 0 1
rlabel polysilicon 597 -556 597 -556 0 3
rlabel polysilicon 607 -550 607 -550 0 2
rlabel polysilicon 607 -556 607 -556 0 4
rlabel polysilicon 611 -550 611 -550 0 1
rlabel polysilicon 611 -556 611 -556 0 3
rlabel polysilicon 618 -550 618 -550 0 1
rlabel polysilicon 618 -556 618 -556 0 3
rlabel polysilicon 625 -550 625 -550 0 1
rlabel polysilicon 625 -556 625 -556 0 3
rlabel polysilicon 632 -550 632 -550 0 1
rlabel polysilicon 632 -556 632 -556 0 3
rlabel polysilicon 639 -550 639 -550 0 1
rlabel polysilicon 639 -556 639 -556 0 3
rlabel polysilicon 646 -550 646 -550 0 1
rlabel polysilicon 646 -556 646 -556 0 3
rlabel polysilicon 653 -550 653 -550 0 1
rlabel polysilicon 653 -556 653 -556 0 3
rlabel polysilicon 660 -550 660 -550 0 1
rlabel polysilicon 660 -556 660 -556 0 3
rlabel polysilicon 667 -550 667 -550 0 1
rlabel polysilicon 667 -556 667 -556 0 3
rlabel polysilicon 674 -550 674 -550 0 1
rlabel polysilicon 674 -556 674 -556 0 3
rlabel polysilicon 681 -550 681 -550 0 1
rlabel polysilicon 681 -556 681 -556 0 3
rlabel polysilicon 688 -550 688 -550 0 1
rlabel polysilicon 688 -556 688 -556 0 3
rlabel polysilicon 695 -550 695 -550 0 1
rlabel polysilicon 695 -556 695 -556 0 3
rlabel polysilicon 702 -550 702 -550 0 1
rlabel polysilicon 702 -556 702 -556 0 3
rlabel polysilicon 709 -550 709 -550 0 1
rlabel polysilicon 709 -556 709 -556 0 3
rlabel polysilicon 716 -550 716 -550 0 1
rlabel polysilicon 716 -556 716 -556 0 3
rlabel polysilicon 723 -550 723 -550 0 1
rlabel polysilicon 726 -550 726 -550 0 2
rlabel polysilicon 723 -556 723 -556 0 3
rlabel polysilicon 726 -556 726 -556 0 4
rlabel polysilicon 730 -550 730 -550 0 1
rlabel polysilicon 730 -556 730 -556 0 3
rlabel polysilicon 737 -550 737 -550 0 1
rlabel polysilicon 737 -556 737 -556 0 3
rlabel polysilicon 744 -550 744 -550 0 1
rlabel polysilicon 744 -556 744 -556 0 3
rlabel polysilicon 754 -550 754 -550 0 2
rlabel polysilicon 751 -556 751 -556 0 3
rlabel polysilicon 754 -556 754 -556 0 4
rlabel polysilicon 758 -550 758 -550 0 1
rlabel polysilicon 758 -556 758 -556 0 3
rlabel polysilicon 765 -550 765 -550 0 1
rlabel polysilicon 765 -556 765 -556 0 3
rlabel polysilicon 772 -550 772 -550 0 1
rlabel polysilicon 772 -556 772 -556 0 3
rlabel polysilicon 779 -550 779 -550 0 1
rlabel polysilicon 779 -556 779 -556 0 3
rlabel polysilicon 786 -550 786 -550 0 1
rlabel polysilicon 786 -556 786 -556 0 3
rlabel polysilicon 796 -550 796 -550 0 2
rlabel polysilicon 793 -556 793 -556 0 3
rlabel polysilicon 800 -550 800 -550 0 1
rlabel polysilicon 800 -556 800 -556 0 3
rlabel polysilicon 807 -550 807 -550 0 1
rlabel polysilicon 807 -556 807 -556 0 3
rlabel polysilicon 814 -550 814 -550 0 1
rlabel polysilicon 814 -556 814 -556 0 3
rlabel polysilicon 821 -550 821 -550 0 1
rlabel polysilicon 821 -556 821 -556 0 3
rlabel polysilicon 835 -550 835 -550 0 1
rlabel polysilicon 835 -556 835 -556 0 3
rlabel polysilicon 856 -550 856 -550 0 1
rlabel polysilicon 856 -556 856 -556 0 3
rlabel polysilicon 2 -633 2 -633 0 1
rlabel polysilicon 2 -639 2 -639 0 3
rlabel polysilicon 9 -633 9 -633 0 1
rlabel polysilicon 9 -639 9 -639 0 3
rlabel polysilicon 16 -633 16 -633 0 1
rlabel polysilicon 16 -639 16 -639 0 3
rlabel polysilicon 23 -633 23 -633 0 1
rlabel polysilicon 23 -639 23 -639 0 3
rlabel polysilicon 30 -633 30 -633 0 1
rlabel polysilicon 30 -639 30 -639 0 3
rlabel polysilicon 40 -633 40 -633 0 2
rlabel polysilicon 44 -633 44 -633 0 1
rlabel polysilicon 44 -639 44 -639 0 3
rlabel polysilicon 51 -633 51 -633 0 1
rlabel polysilicon 51 -639 51 -639 0 3
rlabel polysilicon 61 -633 61 -633 0 2
rlabel polysilicon 58 -639 58 -639 0 3
rlabel polysilicon 61 -639 61 -639 0 4
rlabel polysilicon 65 -633 65 -633 0 1
rlabel polysilicon 65 -639 65 -639 0 3
rlabel polysilicon 72 -633 72 -633 0 1
rlabel polysilicon 72 -639 72 -639 0 3
rlabel polysilicon 79 -633 79 -633 0 1
rlabel polysilicon 79 -639 79 -639 0 3
rlabel polysilicon 86 -633 86 -633 0 1
rlabel polysilicon 86 -639 86 -639 0 3
rlabel polysilicon 93 -633 93 -633 0 1
rlabel polysilicon 93 -639 93 -639 0 3
rlabel polysilicon 103 -633 103 -633 0 2
rlabel polysilicon 100 -639 100 -639 0 3
rlabel polysilicon 103 -639 103 -639 0 4
rlabel polysilicon 107 -633 107 -633 0 1
rlabel polysilicon 107 -639 107 -639 0 3
rlabel polysilicon 114 -633 114 -633 0 1
rlabel polysilicon 114 -639 114 -639 0 3
rlabel polysilicon 124 -633 124 -633 0 2
rlabel polysilicon 121 -639 121 -639 0 3
rlabel polysilicon 131 -633 131 -633 0 2
rlabel polysilicon 128 -639 128 -639 0 3
rlabel polysilicon 135 -633 135 -633 0 1
rlabel polysilicon 135 -639 135 -639 0 3
rlabel polysilicon 138 -639 138 -639 0 4
rlabel polysilicon 142 -639 142 -639 0 3
rlabel polysilicon 145 -639 145 -639 0 4
rlabel polysilicon 149 -633 149 -633 0 1
rlabel polysilicon 149 -639 149 -639 0 3
rlabel polysilicon 156 -633 156 -633 0 1
rlabel polysilicon 156 -639 156 -639 0 3
rlabel polysilicon 163 -633 163 -633 0 1
rlabel polysilicon 163 -639 163 -639 0 3
rlabel polysilicon 173 -633 173 -633 0 2
rlabel polysilicon 170 -639 170 -639 0 3
rlabel polysilicon 173 -639 173 -639 0 4
rlabel polysilicon 177 -633 177 -633 0 1
rlabel polysilicon 177 -639 177 -639 0 3
rlabel polysilicon 184 -633 184 -633 0 1
rlabel polysilicon 184 -639 184 -639 0 3
rlabel polysilicon 191 -633 191 -633 0 1
rlabel polysilicon 191 -639 191 -639 0 3
rlabel polysilicon 198 -633 198 -633 0 1
rlabel polysilicon 198 -639 198 -639 0 3
rlabel polysilicon 205 -633 205 -633 0 1
rlabel polysilicon 205 -639 205 -639 0 3
rlabel polysilicon 212 -633 212 -633 0 1
rlabel polysilicon 212 -639 212 -639 0 3
rlabel polysilicon 219 -633 219 -633 0 1
rlabel polysilicon 219 -639 219 -639 0 3
rlabel polysilicon 226 -633 226 -633 0 1
rlabel polysilicon 226 -639 226 -639 0 3
rlabel polysilicon 233 -633 233 -633 0 1
rlabel polysilicon 236 -633 236 -633 0 2
rlabel polysilicon 236 -639 236 -639 0 4
rlabel polysilicon 240 -633 240 -633 0 1
rlabel polysilicon 240 -639 240 -639 0 3
rlabel polysilicon 243 -639 243 -639 0 4
rlabel polysilicon 247 -633 247 -633 0 1
rlabel polysilicon 247 -639 247 -639 0 3
rlabel polysilicon 254 -633 254 -633 0 1
rlabel polysilicon 254 -639 254 -639 0 3
rlabel polysilicon 261 -633 261 -633 0 1
rlabel polysilicon 261 -639 261 -639 0 3
rlabel polysilicon 268 -633 268 -633 0 1
rlabel polysilicon 268 -639 268 -639 0 3
rlabel polysilicon 275 -633 275 -633 0 1
rlabel polysilicon 275 -639 275 -639 0 3
rlabel polysilicon 282 -633 282 -633 0 1
rlabel polysilicon 282 -639 282 -639 0 3
rlabel polysilicon 289 -633 289 -633 0 1
rlabel polysilicon 289 -639 289 -639 0 3
rlabel polysilicon 296 -633 296 -633 0 1
rlabel polysilicon 296 -639 296 -639 0 3
rlabel polysilicon 306 -633 306 -633 0 2
rlabel polysilicon 303 -639 303 -639 0 3
rlabel polysilicon 310 -633 310 -633 0 1
rlabel polysilicon 313 -633 313 -633 0 2
rlabel polysilicon 310 -639 310 -639 0 3
rlabel polysilicon 317 -633 317 -633 0 1
rlabel polysilicon 317 -639 317 -639 0 3
rlabel polysilicon 324 -633 324 -633 0 1
rlabel polysilicon 324 -639 324 -639 0 3
rlabel polysilicon 331 -633 331 -633 0 1
rlabel polysilicon 334 -633 334 -633 0 2
rlabel polysilicon 331 -639 331 -639 0 3
rlabel polysilicon 338 -633 338 -633 0 1
rlabel polysilicon 341 -633 341 -633 0 2
rlabel polysilicon 338 -639 338 -639 0 3
rlabel polysilicon 341 -639 341 -639 0 4
rlabel polysilicon 345 -633 345 -633 0 1
rlabel polysilicon 348 -633 348 -633 0 2
rlabel polysilicon 352 -633 352 -633 0 1
rlabel polysilicon 352 -639 352 -639 0 3
rlabel polysilicon 359 -633 359 -633 0 1
rlabel polysilicon 359 -639 359 -639 0 3
rlabel polysilicon 366 -633 366 -633 0 1
rlabel polysilicon 366 -639 366 -639 0 3
rlabel polysilicon 373 -633 373 -633 0 1
rlabel polysilicon 373 -639 373 -639 0 3
rlabel polysilicon 380 -633 380 -633 0 1
rlabel polysilicon 380 -639 380 -639 0 3
rlabel polysilicon 387 -633 387 -633 0 1
rlabel polysilicon 387 -639 387 -639 0 3
rlabel polysilicon 394 -633 394 -633 0 1
rlabel polysilicon 394 -639 394 -639 0 3
rlabel polysilicon 401 -633 401 -633 0 1
rlabel polysilicon 404 -633 404 -633 0 2
rlabel polysilicon 401 -639 401 -639 0 3
rlabel polysilicon 404 -639 404 -639 0 4
rlabel polysilicon 408 -633 408 -633 0 1
rlabel polysilicon 408 -639 408 -639 0 3
rlabel polysilicon 415 -633 415 -633 0 1
rlabel polysilicon 415 -639 415 -639 0 3
rlabel polysilicon 422 -633 422 -633 0 1
rlabel polysilicon 422 -639 422 -639 0 3
rlabel polysilicon 429 -633 429 -633 0 1
rlabel polysilicon 429 -639 429 -639 0 3
rlabel polysilicon 436 -633 436 -633 0 1
rlabel polysilicon 436 -639 436 -639 0 3
rlabel polysilicon 443 -633 443 -633 0 1
rlabel polysilicon 443 -639 443 -639 0 3
rlabel polysilicon 450 -633 450 -633 0 1
rlabel polysilicon 453 -639 453 -639 0 4
rlabel polysilicon 457 -633 457 -633 0 1
rlabel polysilicon 457 -639 457 -639 0 3
rlabel polysilicon 464 -633 464 -633 0 1
rlabel polysilicon 467 -633 467 -633 0 2
rlabel polysilicon 464 -639 464 -639 0 3
rlabel polysilicon 467 -639 467 -639 0 4
rlabel polysilicon 471 -633 471 -633 0 1
rlabel polysilicon 474 -633 474 -633 0 2
rlabel polysilicon 471 -639 471 -639 0 3
rlabel polysilicon 474 -639 474 -639 0 4
rlabel polysilicon 478 -633 478 -633 0 1
rlabel polysilicon 478 -639 478 -639 0 3
rlabel polysilicon 485 -633 485 -633 0 1
rlabel polysilicon 485 -639 485 -639 0 3
rlabel polysilicon 492 -633 492 -633 0 1
rlabel polysilicon 492 -639 492 -639 0 3
rlabel polysilicon 499 -633 499 -633 0 1
rlabel polysilicon 499 -639 499 -639 0 3
rlabel polysilicon 506 -633 506 -633 0 1
rlabel polysilicon 506 -639 506 -639 0 3
rlabel polysilicon 513 -633 513 -633 0 1
rlabel polysilicon 513 -639 513 -639 0 3
rlabel polysilicon 523 -633 523 -633 0 2
rlabel polysilicon 520 -639 520 -639 0 3
rlabel polysilicon 523 -639 523 -639 0 4
rlabel polysilicon 527 -633 527 -633 0 1
rlabel polysilicon 527 -639 527 -639 0 3
rlabel polysilicon 537 -633 537 -633 0 2
rlabel polysilicon 537 -639 537 -639 0 4
rlabel polysilicon 541 -633 541 -633 0 1
rlabel polysilicon 544 -633 544 -633 0 2
rlabel polysilicon 541 -639 541 -639 0 3
rlabel polysilicon 548 -633 548 -633 0 1
rlabel polysilicon 548 -639 548 -639 0 3
rlabel polysilicon 555 -633 555 -633 0 1
rlabel polysilicon 555 -639 555 -639 0 3
rlabel polysilicon 562 -633 562 -633 0 1
rlabel polysilicon 562 -639 562 -639 0 3
rlabel polysilicon 569 -633 569 -633 0 1
rlabel polysilicon 569 -639 569 -639 0 3
rlabel polysilicon 576 -633 576 -633 0 1
rlabel polysilicon 576 -639 576 -639 0 3
rlabel polysilicon 583 -633 583 -633 0 1
rlabel polysilicon 583 -639 583 -639 0 3
rlabel polysilicon 590 -633 590 -633 0 1
rlabel polysilicon 593 -633 593 -633 0 2
rlabel polysilicon 593 -639 593 -639 0 4
rlabel polysilicon 597 -633 597 -633 0 1
rlabel polysilicon 597 -639 597 -639 0 3
rlabel polysilicon 604 -633 604 -633 0 1
rlabel polysilicon 604 -639 604 -639 0 3
rlabel polysilicon 611 -633 611 -633 0 1
rlabel polysilicon 611 -639 611 -639 0 3
rlabel polysilicon 614 -639 614 -639 0 4
rlabel polysilicon 621 -639 621 -639 0 4
rlabel polysilicon 625 -633 625 -633 0 1
rlabel polysilicon 625 -639 625 -639 0 3
rlabel polysilicon 632 -633 632 -633 0 1
rlabel polysilicon 632 -639 632 -639 0 3
rlabel polysilicon 639 -633 639 -633 0 1
rlabel polysilicon 639 -639 639 -639 0 3
rlabel polysilicon 646 -633 646 -633 0 1
rlabel polysilicon 646 -639 646 -639 0 3
rlabel polysilicon 653 -633 653 -633 0 1
rlabel polysilicon 653 -639 653 -639 0 3
rlabel polysilicon 660 -633 660 -633 0 1
rlabel polysilicon 660 -639 660 -639 0 3
rlabel polysilicon 667 -633 667 -633 0 1
rlabel polysilicon 667 -639 667 -639 0 3
rlabel polysilicon 674 -633 674 -633 0 1
rlabel polysilicon 674 -639 674 -639 0 3
rlabel polysilicon 681 -633 681 -633 0 1
rlabel polysilicon 681 -639 681 -639 0 3
rlabel polysilicon 688 -633 688 -633 0 1
rlabel polysilicon 688 -639 688 -639 0 3
rlabel polysilicon 698 -633 698 -633 0 2
rlabel polysilicon 702 -633 702 -633 0 1
rlabel polysilicon 702 -639 702 -639 0 3
rlabel polysilicon 709 -633 709 -633 0 1
rlabel polysilicon 709 -639 709 -639 0 3
rlabel polysilicon 716 -633 716 -633 0 1
rlabel polysilicon 716 -639 716 -639 0 3
rlabel polysilicon 723 -633 723 -633 0 1
rlabel polysilicon 723 -639 723 -639 0 3
rlabel polysilicon 730 -633 730 -633 0 1
rlabel polysilicon 730 -639 730 -639 0 3
rlabel polysilicon 737 -633 737 -633 0 1
rlabel polysilicon 737 -639 737 -639 0 3
rlabel polysilicon 744 -633 744 -633 0 1
rlabel polysilicon 744 -639 744 -639 0 3
rlabel polysilicon 751 -633 751 -633 0 1
rlabel polysilicon 751 -639 751 -639 0 3
rlabel polysilicon 758 -633 758 -633 0 1
rlabel polysilicon 758 -639 758 -639 0 3
rlabel polysilicon 765 -633 765 -633 0 1
rlabel polysilicon 765 -639 765 -639 0 3
rlabel polysilicon 772 -633 772 -633 0 1
rlabel polysilicon 772 -639 772 -639 0 3
rlabel polysilicon 779 -633 779 -633 0 1
rlabel polysilicon 779 -639 779 -639 0 3
rlabel polysilicon 786 -633 786 -633 0 1
rlabel polysilicon 786 -639 786 -639 0 3
rlabel polysilicon 793 -633 793 -633 0 1
rlabel polysilicon 793 -639 793 -639 0 3
rlabel polysilicon 800 -633 800 -633 0 1
rlabel polysilicon 800 -639 800 -639 0 3
rlabel polysilicon 807 -633 807 -633 0 1
rlabel polysilicon 807 -639 807 -639 0 3
rlabel polysilicon 814 -633 814 -633 0 1
rlabel polysilicon 814 -639 814 -639 0 3
rlabel polysilicon 821 -633 821 -633 0 1
rlabel polysilicon 821 -639 821 -639 0 3
rlabel polysilicon 828 -633 828 -633 0 1
rlabel polysilicon 828 -639 828 -639 0 3
rlabel polysilicon 835 -633 835 -633 0 1
rlabel polysilicon 835 -639 835 -639 0 3
rlabel polysilicon 842 -633 842 -633 0 1
rlabel polysilicon 842 -639 842 -639 0 3
rlabel polysilicon 849 -633 849 -633 0 1
rlabel polysilicon 849 -639 849 -639 0 3
rlabel polysilicon 856 -633 856 -633 0 1
rlabel polysilicon 856 -639 856 -639 0 3
rlabel polysilicon 863 -633 863 -633 0 1
rlabel polysilicon 863 -639 863 -639 0 3
rlabel polysilicon 870 -633 870 -633 0 1
rlabel polysilicon 870 -639 870 -639 0 3
rlabel polysilicon 877 -633 877 -633 0 1
rlabel polysilicon 877 -639 877 -639 0 3
rlabel polysilicon 884 -633 884 -633 0 1
rlabel polysilicon 884 -639 884 -639 0 3
rlabel polysilicon 891 -633 891 -633 0 1
rlabel polysilicon 891 -639 891 -639 0 3
rlabel polysilicon 898 -633 898 -633 0 1
rlabel polysilicon 898 -639 898 -639 0 3
rlabel polysilicon 905 -633 905 -633 0 1
rlabel polysilicon 905 -639 905 -639 0 3
rlabel polysilicon 912 -633 912 -633 0 1
rlabel polysilicon 912 -639 912 -639 0 3
rlabel polysilicon 919 -639 919 -639 0 3
rlabel polysilicon 926 -633 926 -633 0 1
rlabel polysilicon 926 -639 926 -639 0 3
rlabel polysilicon 947 -633 947 -633 0 1
rlabel polysilicon 947 -639 947 -639 0 3
rlabel polysilicon 2 -712 2 -712 0 1
rlabel polysilicon 2 -718 2 -718 0 3
rlabel polysilicon 9 -712 9 -712 0 1
rlabel polysilicon 9 -718 9 -718 0 3
rlabel polysilicon 16 -712 16 -712 0 1
rlabel polysilicon 16 -718 16 -718 0 3
rlabel polysilicon 26 -718 26 -718 0 4
rlabel polysilicon 30 -718 30 -718 0 3
rlabel polysilicon 33 -718 33 -718 0 4
rlabel polysilicon 37 -712 37 -712 0 1
rlabel polysilicon 37 -718 37 -718 0 3
rlabel polysilicon 44 -712 44 -712 0 1
rlabel polysilicon 44 -718 44 -718 0 3
rlabel polysilicon 51 -712 51 -712 0 1
rlabel polysilicon 51 -718 51 -718 0 3
rlabel polysilicon 58 -712 58 -712 0 1
rlabel polysilicon 58 -718 58 -718 0 3
rlabel polysilicon 65 -712 65 -712 0 1
rlabel polysilicon 65 -718 65 -718 0 3
rlabel polysilicon 72 -712 72 -712 0 1
rlabel polysilicon 72 -718 72 -718 0 3
rlabel polysilicon 79 -712 79 -712 0 1
rlabel polysilicon 79 -718 79 -718 0 3
rlabel polysilicon 86 -712 86 -712 0 1
rlabel polysilicon 89 -712 89 -712 0 2
rlabel polysilicon 86 -718 86 -718 0 3
rlabel polysilicon 89 -718 89 -718 0 4
rlabel polysilicon 93 -712 93 -712 0 1
rlabel polysilicon 93 -718 93 -718 0 3
rlabel polysilicon 100 -712 100 -712 0 1
rlabel polysilicon 103 -712 103 -712 0 2
rlabel polysilicon 100 -718 100 -718 0 3
rlabel polysilicon 103 -718 103 -718 0 4
rlabel polysilicon 110 -712 110 -712 0 2
rlabel polysilicon 107 -718 107 -718 0 3
rlabel polysilicon 110 -718 110 -718 0 4
rlabel polysilicon 114 -712 114 -712 0 1
rlabel polysilicon 114 -718 114 -718 0 3
rlabel polysilicon 121 -712 121 -712 0 1
rlabel polysilicon 121 -718 121 -718 0 3
rlabel polysilicon 128 -718 128 -718 0 3
rlabel polysilicon 131 -718 131 -718 0 4
rlabel polysilicon 135 -712 135 -712 0 1
rlabel polysilicon 135 -718 135 -718 0 3
rlabel polysilicon 145 -712 145 -712 0 2
rlabel polysilicon 142 -718 142 -718 0 3
rlabel polysilicon 145 -718 145 -718 0 4
rlabel polysilicon 149 -712 149 -712 0 1
rlabel polysilicon 149 -718 149 -718 0 3
rlabel polysilicon 156 -712 156 -712 0 1
rlabel polysilicon 156 -718 156 -718 0 3
rlabel polysilicon 163 -712 163 -712 0 1
rlabel polysilicon 163 -718 163 -718 0 3
rlabel polysilicon 170 -712 170 -712 0 1
rlabel polysilicon 170 -718 170 -718 0 3
rlabel polysilicon 177 -712 177 -712 0 1
rlabel polysilicon 177 -718 177 -718 0 3
rlabel polysilicon 184 -712 184 -712 0 1
rlabel polysilicon 184 -718 184 -718 0 3
rlabel polysilicon 191 -712 191 -712 0 1
rlabel polysilicon 191 -718 191 -718 0 3
rlabel polysilicon 198 -712 198 -712 0 1
rlabel polysilicon 198 -718 198 -718 0 3
rlabel polysilicon 205 -712 205 -712 0 1
rlabel polysilicon 205 -718 205 -718 0 3
rlabel polysilicon 212 -712 212 -712 0 1
rlabel polysilicon 212 -718 212 -718 0 3
rlabel polysilicon 219 -712 219 -712 0 1
rlabel polysilicon 219 -718 219 -718 0 3
rlabel polysilicon 229 -712 229 -712 0 2
rlabel polysilicon 229 -718 229 -718 0 4
rlabel polysilicon 233 -712 233 -712 0 1
rlabel polysilicon 233 -718 233 -718 0 3
rlabel polysilicon 240 -712 240 -712 0 1
rlabel polysilicon 243 -712 243 -712 0 2
rlabel polysilicon 240 -718 240 -718 0 3
rlabel polysilicon 243 -718 243 -718 0 4
rlabel polysilicon 250 -712 250 -712 0 2
rlabel polysilicon 250 -718 250 -718 0 4
rlabel polysilicon 254 -712 254 -712 0 1
rlabel polysilicon 254 -718 254 -718 0 3
rlabel polysilicon 261 -712 261 -712 0 1
rlabel polysilicon 261 -718 261 -718 0 3
rlabel polysilicon 268 -712 268 -712 0 1
rlabel polysilicon 268 -718 268 -718 0 3
rlabel polysilicon 275 -712 275 -712 0 1
rlabel polysilicon 275 -718 275 -718 0 3
rlabel polysilicon 282 -712 282 -712 0 1
rlabel polysilicon 282 -718 282 -718 0 3
rlabel polysilicon 289 -712 289 -712 0 1
rlabel polysilicon 289 -718 289 -718 0 3
rlabel polysilicon 296 -712 296 -712 0 1
rlabel polysilicon 296 -718 296 -718 0 3
rlabel polysilicon 303 -712 303 -712 0 1
rlabel polysilicon 303 -718 303 -718 0 3
rlabel polysilicon 310 -712 310 -712 0 1
rlabel polysilicon 310 -718 310 -718 0 3
rlabel polysilicon 317 -712 317 -712 0 1
rlabel polysilicon 317 -718 317 -718 0 3
rlabel polysilicon 324 -712 324 -712 0 1
rlabel polysilicon 324 -718 324 -718 0 3
rlabel polysilicon 334 -712 334 -712 0 2
rlabel polysilicon 338 -712 338 -712 0 1
rlabel polysilicon 338 -718 338 -718 0 3
rlabel polysilicon 345 -712 345 -712 0 1
rlabel polysilicon 348 -712 348 -712 0 2
rlabel polysilicon 345 -718 345 -718 0 3
rlabel polysilicon 348 -718 348 -718 0 4
rlabel polysilicon 352 -712 352 -712 0 1
rlabel polysilicon 352 -718 352 -718 0 3
rlabel polysilicon 359 -712 359 -712 0 1
rlabel polysilicon 359 -718 359 -718 0 3
rlabel polysilicon 366 -712 366 -712 0 1
rlabel polysilicon 366 -718 366 -718 0 3
rlabel polysilicon 373 -718 373 -718 0 3
rlabel polysilicon 376 -718 376 -718 0 4
rlabel polysilicon 380 -712 380 -712 0 1
rlabel polysilicon 380 -718 380 -718 0 3
rlabel polysilicon 390 -712 390 -712 0 2
rlabel polysilicon 387 -718 387 -718 0 3
rlabel polysilicon 394 -712 394 -712 0 1
rlabel polysilicon 394 -718 394 -718 0 3
rlabel polysilicon 401 -712 401 -712 0 1
rlabel polysilicon 401 -718 401 -718 0 3
rlabel polysilicon 408 -712 408 -712 0 1
rlabel polysilicon 411 -712 411 -712 0 2
rlabel polysilicon 408 -718 408 -718 0 3
rlabel polysilicon 415 -712 415 -712 0 1
rlabel polysilicon 418 -712 418 -712 0 2
rlabel polysilicon 415 -718 415 -718 0 3
rlabel polysilicon 418 -718 418 -718 0 4
rlabel polysilicon 422 -712 422 -712 0 1
rlabel polysilicon 422 -718 422 -718 0 3
rlabel polysilicon 429 -712 429 -712 0 1
rlabel polysilicon 429 -718 429 -718 0 3
rlabel polysilicon 436 -712 436 -712 0 1
rlabel polysilicon 436 -718 436 -718 0 3
rlabel polysilicon 443 -712 443 -712 0 1
rlabel polysilicon 443 -718 443 -718 0 3
rlabel polysilicon 450 -712 450 -712 0 1
rlabel polysilicon 450 -718 450 -718 0 3
rlabel polysilicon 457 -712 457 -712 0 1
rlabel polysilicon 457 -718 457 -718 0 3
rlabel polysilicon 464 -712 464 -712 0 1
rlabel polysilicon 464 -718 464 -718 0 3
rlabel polysilicon 471 -712 471 -712 0 1
rlabel polysilicon 474 -712 474 -712 0 2
rlabel polysilicon 478 -712 478 -712 0 1
rlabel polysilicon 481 -712 481 -712 0 2
rlabel polysilicon 478 -718 478 -718 0 3
rlabel polysilicon 481 -718 481 -718 0 4
rlabel polysilicon 485 -712 485 -712 0 1
rlabel polysilicon 488 -712 488 -712 0 2
rlabel polysilicon 485 -718 485 -718 0 3
rlabel polysilicon 488 -718 488 -718 0 4
rlabel polysilicon 492 -712 492 -712 0 1
rlabel polysilicon 492 -718 492 -718 0 3
rlabel polysilicon 502 -712 502 -712 0 2
rlabel polysilicon 499 -718 499 -718 0 3
rlabel polysilicon 502 -718 502 -718 0 4
rlabel polysilicon 506 -712 506 -712 0 1
rlabel polysilicon 506 -718 506 -718 0 3
rlabel polysilicon 513 -718 513 -718 0 3
rlabel polysilicon 516 -718 516 -718 0 4
rlabel polysilicon 520 -712 520 -712 0 1
rlabel polysilicon 520 -718 520 -718 0 3
rlabel polysilicon 527 -712 527 -712 0 1
rlabel polysilicon 527 -718 527 -718 0 3
rlabel polysilicon 534 -712 534 -712 0 1
rlabel polysilicon 534 -718 534 -718 0 3
rlabel polysilicon 541 -712 541 -712 0 1
rlabel polysilicon 544 -712 544 -712 0 2
rlabel polysilicon 541 -718 541 -718 0 3
rlabel polysilicon 544 -718 544 -718 0 4
rlabel polysilicon 548 -712 548 -712 0 1
rlabel polysilicon 551 -712 551 -712 0 2
rlabel polysilicon 551 -718 551 -718 0 4
rlabel polysilicon 555 -712 555 -712 0 1
rlabel polysilicon 558 -712 558 -712 0 2
rlabel polysilicon 558 -718 558 -718 0 4
rlabel polysilicon 562 -712 562 -712 0 1
rlabel polysilicon 565 -712 565 -712 0 2
rlabel polysilicon 562 -718 562 -718 0 3
rlabel polysilicon 569 -712 569 -712 0 1
rlabel polysilicon 569 -718 569 -718 0 3
rlabel polysilicon 576 -712 576 -712 0 1
rlabel polysilicon 576 -718 576 -718 0 3
rlabel polysilicon 583 -712 583 -712 0 1
rlabel polysilicon 583 -718 583 -718 0 3
rlabel polysilicon 590 -712 590 -712 0 1
rlabel polysilicon 593 -712 593 -712 0 2
rlabel polysilicon 590 -718 590 -718 0 3
rlabel polysilicon 597 -712 597 -712 0 1
rlabel polysilicon 597 -718 597 -718 0 3
rlabel polysilicon 604 -712 604 -712 0 1
rlabel polysilicon 604 -718 604 -718 0 3
rlabel polysilicon 611 -712 611 -712 0 1
rlabel polysilicon 611 -718 611 -718 0 3
rlabel polysilicon 618 -712 618 -712 0 1
rlabel polysilicon 618 -718 618 -718 0 3
rlabel polysilicon 625 -712 625 -712 0 1
rlabel polysilicon 628 -712 628 -712 0 2
rlabel polysilicon 625 -718 625 -718 0 3
rlabel polysilicon 628 -718 628 -718 0 4
rlabel polysilicon 632 -712 632 -712 0 1
rlabel polysilicon 632 -718 632 -718 0 3
rlabel polysilicon 639 -712 639 -712 0 1
rlabel polysilicon 639 -718 639 -718 0 3
rlabel polysilicon 646 -712 646 -712 0 1
rlabel polysilicon 646 -718 646 -718 0 3
rlabel polysilicon 653 -712 653 -712 0 1
rlabel polysilicon 653 -718 653 -718 0 3
rlabel polysilicon 660 -712 660 -712 0 1
rlabel polysilicon 660 -718 660 -718 0 3
rlabel polysilicon 667 -712 667 -712 0 1
rlabel polysilicon 667 -718 667 -718 0 3
rlabel polysilicon 674 -712 674 -712 0 1
rlabel polysilicon 674 -718 674 -718 0 3
rlabel polysilicon 681 -712 681 -712 0 1
rlabel polysilicon 681 -718 681 -718 0 3
rlabel polysilicon 688 -712 688 -712 0 1
rlabel polysilicon 688 -718 688 -718 0 3
rlabel polysilicon 695 -712 695 -712 0 1
rlabel polysilicon 695 -718 695 -718 0 3
rlabel polysilicon 702 -712 702 -712 0 1
rlabel polysilicon 702 -718 702 -718 0 3
rlabel polysilicon 709 -712 709 -712 0 1
rlabel polysilicon 709 -718 709 -718 0 3
rlabel polysilicon 716 -712 716 -712 0 1
rlabel polysilicon 716 -718 716 -718 0 3
rlabel polysilicon 723 -712 723 -712 0 1
rlabel polysilicon 723 -718 723 -718 0 3
rlabel polysilicon 730 -712 730 -712 0 1
rlabel polysilicon 730 -718 730 -718 0 3
rlabel polysilicon 737 -712 737 -712 0 1
rlabel polysilicon 737 -718 737 -718 0 3
rlabel polysilicon 744 -712 744 -712 0 1
rlabel polysilicon 744 -718 744 -718 0 3
rlabel polysilicon 751 -712 751 -712 0 1
rlabel polysilicon 751 -718 751 -718 0 3
rlabel polysilicon 758 -712 758 -712 0 1
rlabel polysilicon 758 -718 758 -718 0 3
rlabel polysilicon 765 -712 765 -712 0 1
rlabel polysilicon 765 -718 765 -718 0 3
rlabel polysilicon 772 -712 772 -712 0 1
rlabel polysilicon 772 -718 772 -718 0 3
rlabel polysilicon 779 -712 779 -712 0 1
rlabel polysilicon 779 -718 779 -718 0 3
rlabel polysilicon 786 -712 786 -712 0 1
rlabel polysilicon 786 -718 786 -718 0 3
rlabel polysilicon 793 -712 793 -712 0 1
rlabel polysilicon 793 -718 793 -718 0 3
rlabel polysilicon 800 -712 800 -712 0 1
rlabel polysilicon 800 -718 800 -718 0 3
rlabel polysilicon 807 -712 807 -712 0 1
rlabel polysilicon 807 -718 807 -718 0 3
rlabel polysilicon 814 -712 814 -712 0 1
rlabel polysilicon 814 -718 814 -718 0 3
rlabel polysilicon 821 -712 821 -712 0 1
rlabel polysilicon 821 -718 821 -718 0 3
rlabel polysilicon 828 -712 828 -712 0 1
rlabel polysilicon 828 -718 828 -718 0 3
rlabel polysilicon 835 -712 835 -712 0 1
rlabel polysilicon 835 -718 835 -718 0 3
rlabel polysilicon 842 -712 842 -712 0 1
rlabel polysilicon 842 -718 842 -718 0 3
rlabel polysilicon 849 -712 849 -712 0 1
rlabel polysilicon 849 -718 849 -718 0 3
rlabel polysilicon 856 -712 856 -712 0 1
rlabel polysilicon 856 -718 856 -718 0 3
rlabel polysilicon 863 -712 863 -712 0 1
rlabel polysilicon 863 -718 863 -718 0 3
rlabel polysilicon 870 -712 870 -712 0 1
rlabel polysilicon 870 -718 870 -718 0 3
rlabel polysilicon 877 -712 877 -712 0 1
rlabel polysilicon 877 -718 877 -718 0 3
rlabel polysilicon 887 -712 887 -712 0 2
rlabel polysilicon 891 -712 891 -712 0 1
rlabel polysilicon 891 -718 891 -718 0 3
rlabel polysilicon 898 -712 898 -712 0 1
rlabel polysilicon 898 -718 898 -718 0 3
rlabel polysilicon 905 -712 905 -712 0 1
rlabel polysilicon 905 -718 905 -718 0 3
rlabel polysilicon 912 -712 912 -712 0 1
rlabel polysilicon 912 -718 912 -718 0 3
rlabel polysilicon 919 -712 919 -712 0 1
rlabel polysilicon 919 -718 919 -718 0 3
rlabel polysilicon 926 -712 926 -712 0 1
rlabel polysilicon 926 -718 926 -718 0 3
rlabel polysilicon 954 -712 954 -712 0 1
rlabel polysilicon 954 -718 954 -718 0 3
rlabel polysilicon 1031 -712 1031 -712 0 1
rlabel polysilicon 1031 -718 1031 -718 0 3
rlabel polysilicon 23 -783 23 -783 0 1
rlabel polysilicon 23 -789 23 -789 0 3
rlabel polysilicon 30 -783 30 -783 0 1
rlabel polysilicon 30 -789 30 -789 0 3
rlabel polysilicon 37 -783 37 -783 0 1
rlabel polysilicon 37 -789 37 -789 0 3
rlabel polysilicon 44 -783 44 -783 0 1
rlabel polysilicon 44 -789 44 -789 0 3
rlabel polysilicon 51 -783 51 -783 0 1
rlabel polysilicon 58 -783 58 -783 0 1
rlabel polysilicon 58 -789 58 -789 0 3
rlabel polysilicon 65 -789 65 -789 0 3
rlabel polysilicon 72 -789 72 -789 0 3
rlabel polysilicon 79 -783 79 -783 0 1
rlabel polysilicon 79 -789 79 -789 0 3
rlabel polysilicon 86 -783 86 -783 0 1
rlabel polysilicon 86 -789 86 -789 0 3
rlabel polysilicon 93 -783 93 -783 0 1
rlabel polysilicon 93 -789 93 -789 0 3
rlabel polysilicon 100 -783 100 -783 0 1
rlabel polysilicon 100 -789 100 -789 0 3
rlabel polysilicon 107 -783 107 -783 0 1
rlabel polysilicon 110 -783 110 -783 0 2
rlabel polysilicon 110 -789 110 -789 0 4
rlabel polysilicon 114 -783 114 -783 0 1
rlabel polysilicon 117 -783 117 -783 0 2
rlabel polysilicon 114 -789 114 -789 0 3
rlabel polysilicon 121 -783 121 -783 0 1
rlabel polysilicon 121 -789 121 -789 0 3
rlabel polysilicon 128 -783 128 -783 0 1
rlabel polysilicon 128 -789 128 -789 0 3
rlabel polysilicon 135 -783 135 -783 0 1
rlabel polysilicon 135 -789 135 -789 0 3
rlabel polysilicon 142 -783 142 -783 0 1
rlabel polysilicon 142 -789 142 -789 0 3
rlabel polysilicon 149 -783 149 -783 0 1
rlabel polysilicon 149 -789 149 -789 0 3
rlabel polysilicon 156 -783 156 -783 0 1
rlabel polysilicon 156 -789 156 -789 0 3
rlabel polysilicon 163 -783 163 -783 0 1
rlabel polysilicon 163 -789 163 -789 0 3
rlabel polysilicon 170 -783 170 -783 0 1
rlabel polysilicon 170 -789 170 -789 0 3
rlabel polysilicon 177 -783 177 -783 0 1
rlabel polysilicon 177 -789 177 -789 0 3
rlabel polysilicon 184 -783 184 -783 0 1
rlabel polysilicon 187 -783 187 -783 0 2
rlabel polysilicon 184 -789 184 -789 0 3
rlabel polysilicon 191 -783 191 -783 0 1
rlabel polysilicon 191 -789 191 -789 0 3
rlabel polysilicon 198 -783 198 -783 0 1
rlabel polysilicon 198 -789 198 -789 0 3
rlabel polysilicon 205 -783 205 -783 0 1
rlabel polysilicon 205 -789 205 -789 0 3
rlabel polysilicon 212 -783 212 -783 0 1
rlabel polysilicon 212 -789 212 -789 0 3
rlabel polysilicon 219 -783 219 -783 0 1
rlabel polysilicon 219 -789 219 -789 0 3
rlabel polysilicon 226 -789 226 -789 0 3
rlabel polysilicon 229 -789 229 -789 0 4
rlabel polysilicon 236 -783 236 -783 0 2
rlabel polysilicon 233 -789 233 -789 0 3
rlabel polysilicon 236 -789 236 -789 0 4
rlabel polysilicon 243 -783 243 -783 0 2
rlabel polysilicon 240 -789 240 -789 0 3
rlabel polysilicon 247 -783 247 -783 0 1
rlabel polysilicon 247 -789 247 -789 0 3
rlabel polysilicon 254 -783 254 -783 0 1
rlabel polysilicon 254 -789 254 -789 0 3
rlabel polysilicon 261 -783 261 -783 0 1
rlabel polysilicon 264 -783 264 -783 0 2
rlabel polysilicon 261 -789 261 -789 0 3
rlabel polysilicon 268 -783 268 -783 0 1
rlabel polysilicon 268 -789 268 -789 0 3
rlabel polysilicon 275 -783 275 -783 0 1
rlabel polysilicon 275 -789 275 -789 0 3
rlabel polysilicon 282 -783 282 -783 0 1
rlabel polysilicon 282 -789 282 -789 0 3
rlabel polysilicon 289 -783 289 -783 0 1
rlabel polysilicon 289 -789 289 -789 0 3
rlabel polysilicon 296 -783 296 -783 0 1
rlabel polysilicon 296 -789 296 -789 0 3
rlabel polysilicon 303 -783 303 -783 0 1
rlabel polysilicon 303 -789 303 -789 0 3
rlabel polysilicon 310 -783 310 -783 0 1
rlabel polysilicon 313 -789 313 -789 0 4
rlabel polysilicon 317 -783 317 -783 0 1
rlabel polysilicon 317 -789 317 -789 0 3
rlabel polysilicon 324 -783 324 -783 0 1
rlabel polysilicon 324 -789 324 -789 0 3
rlabel polysilicon 331 -783 331 -783 0 1
rlabel polysilicon 331 -789 331 -789 0 3
rlabel polysilicon 338 -783 338 -783 0 1
rlabel polysilicon 345 -783 345 -783 0 1
rlabel polysilicon 345 -789 345 -789 0 3
rlabel polysilicon 352 -783 352 -783 0 1
rlabel polysilicon 355 -783 355 -783 0 2
rlabel polysilicon 352 -789 352 -789 0 3
rlabel polysilicon 355 -789 355 -789 0 4
rlabel polysilicon 359 -783 359 -783 0 1
rlabel polysilicon 359 -789 359 -789 0 3
rlabel polysilicon 366 -783 366 -783 0 1
rlabel polysilicon 366 -789 366 -789 0 3
rlabel polysilicon 373 -783 373 -783 0 1
rlabel polysilicon 373 -789 373 -789 0 3
rlabel polysilicon 380 -783 380 -783 0 1
rlabel polysilicon 380 -789 380 -789 0 3
rlabel polysilicon 387 -783 387 -783 0 1
rlabel polysilicon 390 -783 390 -783 0 2
rlabel polysilicon 387 -789 387 -789 0 3
rlabel polysilicon 394 -783 394 -783 0 1
rlabel polysilicon 394 -789 394 -789 0 3
rlabel polysilicon 401 -783 401 -783 0 1
rlabel polysilicon 404 -783 404 -783 0 2
rlabel polysilicon 408 -783 408 -783 0 1
rlabel polysilicon 408 -789 408 -789 0 3
rlabel polysilicon 415 -783 415 -783 0 1
rlabel polysilicon 415 -789 415 -789 0 3
rlabel polysilicon 422 -789 422 -789 0 3
rlabel polysilicon 425 -789 425 -789 0 4
rlabel polysilicon 429 -783 429 -783 0 1
rlabel polysilicon 429 -789 429 -789 0 3
rlabel polysilicon 436 -783 436 -783 0 1
rlabel polysilicon 436 -789 436 -789 0 3
rlabel polysilicon 443 -783 443 -783 0 1
rlabel polysilicon 443 -789 443 -789 0 3
rlabel polysilicon 450 -783 450 -783 0 1
rlabel polysilicon 450 -789 450 -789 0 3
rlabel polysilicon 457 -783 457 -783 0 1
rlabel polysilicon 457 -789 457 -789 0 3
rlabel polysilicon 464 -783 464 -783 0 1
rlabel polysilicon 464 -789 464 -789 0 3
rlabel polysilicon 471 -783 471 -783 0 1
rlabel polysilicon 471 -789 471 -789 0 3
rlabel polysilicon 478 -783 478 -783 0 1
rlabel polysilicon 478 -789 478 -789 0 3
rlabel polysilicon 485 -783 485 -783 0 1
rlabel polysilicon 485 -789 485 -789 0 3
rlabel polysilicon 492 -783 492 -783 0 1
rlabel polysilicon 495 -783 495 -783 0 2
rlabel polysilicon 492 -789 492 -789 0 3
rlabel polysilicon 499 -783 499 -783 0 1
rlabel polysilicon 499 -789 499 -789 0 3
rlabel polysilicon 506 -783 506 -783 0 1
rlabel polysilicon 506 -789 506 -789 0 3
rlabel polysilicon 513 -783 513 -783 0 1
rlabel polysilicon 513 -789 513 -789 0 3
rlabel polysilicon 516 -789 516 -789 0 4
rlabel polysilicon 520 -783 520 -783 0 1
rlabel polysilicon 520 -789 520 -789 0 3
rlabel polysilicon 527 -783 527 -783 0 1
rlabel polysilicon 530 -783 530 -783 0 2
rlabel polysilicon 527 -789 527 -789 0 3
rlabel polysilicon 530 -789 530 -789 0 4
rlabel polysilicon 534 -783 534 -783 0 1
rlabel polysilicon 534 -789 534 -789 0 3
rlabel polysilicon 541 -783 541 -783 0 1
rlabel polysilicon 548 -783 548 -783 0 1
rlabel polysilicon 548 -789 548 -789 0 3
rlabel polysilicon 555 -783 555 -783 0 1
rlabel polysilicon 555 -789 555 -789 0 3
rlabel polysilicon 565 -783 565 -783 0 2
rlabel polysilicon 562 -789 562 -789 0 3
rlabel polysilicon 565 -789 565 -789 0 4
rlabel polysilicon 569 -783 569 -783 0 1
rlabel polysilicon 569 -789 569 -789 0 3
rlabel polysilicon 576 -783 576 -783 0 1
rlabel polysilicon 579 -783 579 -783 0 2
rlabel polysilicon 576 -789 576 -789 0 3
rlabel polysilicon 579 -789 579 -789 0 4
rlabel polysilicon 583 -783 583 -783 0 1
rlabel polysilicon 583 -789 583 -789 0 3
rlabel polysilicon 590 -783 590 -783 0 1
rlabel polysilicon 590 -789 590 -789 0 3
rlabel polysilicon 597 -783 597 -783 0 1
rlabel polysilicon 597 -789 597 -789 0 3
rlabel polysilicon 604 -783 604 -783 0 1
rlabel polysilicon 604 -789 604 -789 0 3
rlabel polysilicon 611 -783 611 -783 0 1
rlabel polysilicon 611 -789 611 -789 0 3
rlabel polysilicon 618 -783 618 -783 0 1
rlabel polysilicon 621 -783 621 -783 0 2
rlabel polysilicon 618 -789 618 -789 0 3
rlabel polysilicon 621 -789 621 -789 0 4
rlabel polysilicon 625 -783 625 -783 0 1
rlabel polysilicon 625 -789 625 -789 0 3
rlabel polysilicon 632 -783 632 -783 0 1
rlabel polysilicon 632 -789 632 -789 0 3
rlabel polysilicon 639 -783 639 -783 0 1
rlabel polysilicon 639 -789 639 -789 0 3
rlabel polysilicon 646 -783 646 -783 0 1
rlabel polysilicon 646 -789 646 -789 0 3
rlabel polysilicon 653 -783 653 -783 0 1
rlabel polysilicon 653 -789 653 -789 0 3
rlabel polysilicon 660 -783 660 -783 0 1
rlabel polysilicon 660 -789 660 -789 0 3
rlabel polysilicon 667 -783 667 -783 0 1
rlabel polysilicon 670 -783 670 -783 0 2
rlabel polysilicon 667 -789 667 -789 0 3
rlabel polysilicon 674 -783 674 -783 0 1
rlabel polysilicon 674 -789 674 -789 0 3
rlabel polysilicon 681 -783 681 -783 0 1
rlabel polysilicon 681 -789 681 -789 0 3
rlabel polysilicon 688 -783 688 -783 0 1
rlabel polysilicon 688 -789 688 -789 0 3
rlabel polysilicon 695 -783 695 -783 0 1
rlabel polysilicon 695 -789 695 -789 0 3
rlabel polysilicon 702 -783 702 -783 0 1
rlabel polysilicon 702 -789 702 -789 0 3
rlabel polysilicon 709 -783 709 -783 0 1
rlabel polysilicon 709 -789 709 -789 0 3
rlabel polysilicon 716 -783 716 -783 0 1
rlabel polysilicon 716 -789 716 -789 0 3
rlabel polysilicon 723 -783 723 -783 0 1
rlabel polysilicon 723 -789 723 -789 0 3
rlabel polysilicon 730 -783 730 -783 0 1
rlabel polysilicon 730 -789 730 -789 0 3
rlabel polysilicon 737 -783 737 -783 0 1
rlabel polysilicon 737 -789 737 -789 0 3
rlabel polysilicon 744 -783 744 -783 0 1
rlabel polysilicon 744 -789 744 -789 0 3
rlabel polysilicon 751 -783 751 -783 0 1
rlabel polysilicon 751 -789 751 -789 0 3
rlabel polysilicon 758 -783 758 -783 0 1
rlabel polysilicon 758 -789 758 -789 0 3
rlabel polysilicon 765 -783 765 -783 0 1
rlabel polysilicon 765 -789 765 -789 0 3
rlabel polysilicon 772 -783 772 -783 0 1
rlabel polysilicon 772 -789 772 -789 0 3
rlabel polysilicon 779 -783 779 -783 0 1
rlabel polysilicon 779 -789 779 -789 0 3
rlabel polysilicon 786 -783 786 -783 0 1
rlabel polysilicon 786 -789 786 -789 0 3
rlabel polysilicon 793 -783 793 -783 0 1
rlabel polysilicon 793 -789 793 -789 0 3
rlabel polysilicon 800 -783 800 -783 0 1
rlabel polysilicon 800 -789 800 -789 0 3
rlabel polysilicon 807 -783 807 -783 0 1
rlabel polysilicon 807 -789 807 -789 0 3
rlabel polysilicon 814 -783 814 -783 0 1
rlabel polysilicon 814 -789 814 -789 0 3
rlabel polysilicon 821 -783 821 -783 0 1
rlabel polysilicon 821 -789 821 -789 0 3
rlabel polysilicon 828 -783 828 -783 0 1
rlabel polysilicon 828 -789 828 -789 0 3
rlabel polysilicon 835 -783 835 -783 0 1
rlabel polysilicon 835 -789 835 -789 0 3
rlabel polysilicon 842 -783 842 -783 0 1
rlabel polysilicon 842 -789 842 -789 0 3
rlabel polysilicon 849 -783 849 -783 0 1
rlabel polysilicon 849 -789 849 -789 0 3
rlabel polysilicon 856 -783 856 -783 0 1
rlabel polysilicon 856 -789 856 -789 0 3
rlabel polysilicon 863 -783 863 -783 0 1
rlabel polysilicon 863 -789 863 -789 0 3
rlabel polysilicon 870 -783 870 -783 0 1
rlabel polysilicon 870 -789 870 -789 0 3
rlabel polysilicon 877 -783 877 -783 0 1
rlabel polysilicon 877 -789 877 -789 0 3
rlabel polysilicon 884 -783 884 -783 0 1
rlabel polysilicon 884 -789 884 -789 0 3
rlabel polysilicon 891 -783 891 -783 0 1
rlabel polysilicon 891 -789 891 -789 0 3
rlabel polysilicon 894 -789 894 -789 0 4
rlabel polysilicon 898 -783 898 -783 0 1
rlabel polysilicon 898 -789 898 -789 0 3
rlabel polysilicon 908 -783 908 -783 0 2
rlabel polysilicon 905 -789 905 -789 0 3
rlabel polysilicon 908 -789 908 -789 0 4
rlabel polysilicon 912 -783 912 -783 0 1
rlabel polysilicon 915 -783 915 -783 0 2
rlabel polysilicon 915 -789 915 -789 0 4
rlabel polysilicon 919 -783 919 -783 0 1
rlabel polysilicon 919 -789 919 -789 0 3
rlabel polysilicon 961 -783 961 -783 0 1
rlabel polysilicon 961 -789 961 -789 0 3
rlabel polysilicon 975 -783 975 -783 0 1
rlabel polysilicon 975 -789 975 -789 0 3
rlabel polysilicon 989 -789 989 -789 0 3
rlabel polysilicon 1006 -783 1006 -783 0 2
rlabel polysilicon 1010 -783 1010 -783 0 1
rlabel polysilicon 1010 -789 1010 -789 0 3
rlabel polysilicon 1017 -783 1017 -783 0 1
rlabel polysilicon 1017 -789 1017 -789 0 3
rlabel polysilicon 1066 -783 1066 -783 0 1
rlabel polysilicon 1066 -789 1066 -789 0 3
rlabel polysilicon 2 -880 2 -880 0 1
rlabel polysilicon 2 -886 2 -886 0 3
rlabel polysilicon 12 -880 12 -880 0 2
rlabel polysilicon 16 -880 16 -880 0 1
rlabel polysilicon 16 -886 16 -886 0 3
rlabel polysilicon 23 -880 23 -880 0 1
rlabel polysilicon 23 -886 23 -886 0 3
rlabel polysilicon 30 -880 30 -880 0 1
rlabel polysilicon 30 -886 30 -886 0 3
rlabel polysilicon 37 -880 37 -880 0 1
rlabel polysilicon 37 -886 37 -886 0 3
rlabel polysilicon 47 -880 47 -880 0 2
rlabel polysilicon 44 -886 44 -886 0 3
rlabel polysilicon 51 -880 51 -880 0 1
rlabel polysilicon 51 -886 51 -886 0 3
rlabel polysilicon 58 -880 58 -880 0 1
rlabel polysilicon 58 -886 58 -886 0 3
rlabel polysilicon 68 -880 68 -880 0 2
rlabel polysilicon 72 -880 72 -880 0 1
rlabel polysilicon 72 -886 72 -886 0 3
rlabel polysilicon 79 -880 79 -880 0 1
rlabel polysilicon 79 -886 79 -886 0 3
rlabel polysilicon 86 -880 86 -880 0 1
rlabel polysilicon 86 -886 86 -886 0 3
rlabel polysilicon 93 -880 93 -880 0 1
rlabel polysilicon 93 -886 93 -886 0 3
rlabel polysilicon 100 -880 100 -880 0 1
rlabel polysilicon 100 -886 100 -886 0 3
rlabel polysilicon 110 -880 110 -880 0 2
rlabel polysilicon 107 -886 107 -886 0 3
rlabel polysilicon 110 -886 110 -886 0 4
rlabel polysilicon 114 -880 114 -880 0 1
rlabel polysilicon 117 -880 117 -880 0 2
rlabel polysilicon 114 -886 114 -886 0 3
rlabel polysilicon 121 -880 121 -880 0 1
rlabel polysilicon 121 -886 121 -886 0 3
rlabel polysilicon 131 -880 131 -880 0 2
rlabel polysilicon 131 -886 131 -886 0 4
rlabel polysilicon 135 -880 135 -880 0 1
rlabel polysilicon 138 -880 138 -880 0 2
rlabel polysilicon 142 -880 142 -880 0 1
rlabel polysilicon 142 -886 142 -886 0 3
rlabel polysilicon 149 -880 149 -880 0 1
rlabel polysilicon 149 -886 149 -886 0 3
rlabel polysilicon 156 -880 156 -880 0 1
rlabel polysilicon 156 -886 156 -886 0 3
rlabel polysilicon 163 -880 163 -880 0 1
rlabel polysilicon 163 -886 163 -886 0 3
rlabel polysilicon 170 -880 170 -880 0 1
rlabel polysilicon 173 -880 173 -880 0 2
rlabel polysilicon 170 -886 170 -886 0 3
rlabel polysilicon 173 -886 173 -886 0 4
rlabel polysilicon 177 -880 177 -880 0 1
rlabel polysilicon 180 -880 180 -880 0 2
rlabel polysilicon 180 -886 180 -886 0 4
rlabel polysilicon 184 -880 184 -880 0 1
rlabel polysilicon 184 -886 184 -886 0 3
rlabel polysilicon 191 -880 191 -880 0 1
rlabel polysilicon 191 -886 191 -886 0 3
rlabel polysilicon 198 -880 198 -880 0 1
rlabel polysilicon 198 -886 198 -886 0 3
rlabel polysilicon 205 -880 205 -880 0 1
rlabel polysilicon 208 -880 208 -880 0 2
rlabel polysilicon 208 -886 208 -886 0 4
rlabel polysilicon 212 -880 212 -880 0 1
rlabel polysilicon 215 -886 215 -886 0 4
rlabel polysilicon 219 -880 219 -880 0 1
rlabel polysilicon 222 -886 222 -886 0 4
rlabel polysilicon 229 -880 229 -880 0 2
rlabel polysilicon 229 -886 229 -886 0 4
rlabel polysilicon 233 -880 233 -880 0 1
rlabel polysilicon 233 -886 233 -886 0 3
rlabel polysilicon 240 -880 240 -880 0 1
rlabel polysilicon 243 -880 243 -880 0 2
rlabel polysilicon 240 -886 240 -886 0 3
rlabel polysilicon 243 -886 243 -886 0 4
rlabel polysilicon 247 -880 247 -880 0 1
rlabel polysilicon 247 -886 247 -886 0 3
rlabel polysilicon 254 -880 254 -880 0 1
rlabel polysilicon 254 -886 254 -886 0 3
rlabel polysilicon 261 -880 261 -880 0 1
rlabel polysilicon 261 -886 261 -886 0 3
rlabel polysilicon 268 -880 268 -880 0 1
rlabel polysilicon 268 -886 268 -886 0 3
rlabel polysilicon 275 -880 275 -880 0 1
rlabel polysilicon 275 -886 275 -886 0 3
rlabel polysilicon 282 -880 282 -880 0 1
rlabel polysilicon 282 -886 282 -886 0 3
rlabel polysilicon 289 -880 289 -880 0 1
rlabel polysilicon 289 -886 289 -886 0 3
rlabel polysilicon 296 -880 296 -880 0 1
rlabel polysilicon 296 -886 296 -886 0 3
rlabel polysilicon 303 -880 303 -880 0 1
rlabel polysilicon 303 -886 303 -886 0 3
rlabel polysilicon 310 -880 310 -880 0 1
rlabel polysilicon 310 -886 310 -886 0 3
rlabel polysilicon 317 -880 317 -880 0 1
rlabel polysilicon 317 -886 317 -886 0 3
rlabel polysilicon 324 -880 324 -880 0 1
rlabel polysilicon 324 -886 324 -886 0 3
rlabel polysilicon 331 -880 331 -880 0 1
rlabel polysilicon 331 -886 331 -886 0 3
rlabel polysilicon 338 -880 338 -880 0 1
rlabel polysilicon 338 -886 338 -886 0 3
rlabel polysilicon 345 -880 345 -880 0 1
rlabel polysilicon 345 -886 345 -886 0 3
rlabel polysilicon 352 -880 352 -880 0 1
rlabel polysilicon 355 -880 355 -880 0 2
rlabel polysilicon 352 -886 352 -886 0 3
rlabel polysilicon 355 -886 355 -886 0 4
rlabel polysilicon 359 -880 359 -880 0 1
rlabel polysilicon 362 -880 362 -880 0 2
rlabel polysilicon 366 -880 366 -880 0 1
rlabel polysilicon 369 -880 369 -880 0 2
rlabel polysilicon 366 -886 366 -886 0 3
rlabel polysilicon 369 -886 369 -886 0 4
rlabel polysilicon 373 -880 373 -880 0 1
rlabel polysilicon 373 -886 373 -886 0 3
rlabel polysilicon 380 -880 380 -880 0 1
rlabel polysilicon 380 -886 380 -886 0 3
rlabel polysilicon 387 -880 387 -880 0 1
rlabel polysilicon 387 -886 387 -886 0 3
rlabel polysilicon 394 -880 394 -880 0 1
rlabel polysilicon 394 -886 394 -886 0 3
rlabel polysilicon 401 -880 401 -880 0 1
rlabel polysilicon 401 -886 401 -886 0 3
rlabel polysilicon 408 -880 408 -880 0 1
rlabel polysilicon 411 -880 411 -880 0 2
rlabel polysilicon 408 -886 408 -886 0 3
rlabel polysilicon 411 -886 411 -886 0 4
rlabel polysilicon 415 -880 415 -880 0 1
rlabel polysilicon 415 -886 415 -886 0 3
rlabel polysilicon 422 -880 422 -880 0 1
rlabel polysilicon 422 -886 422 -886 0 3
rlabel polysilicon 429 -880 429 -880 0 1
rlabel polysilicon 429 -886 429 -886 0 3
rlabel polysilicon 436 -880 436 -880 0 1
rlabel polysilicon 439 -880 439 -880 0 2
rlabel polysilicon 436 -886 436 -886 0 3
rlabel polysilicon 439 -886 439 -886 0 4
rlabel polysilicon 443 -880 443 -880 0 1
rlabel polysilicon 443 -886 443 -886 0 3
rlabel polysilicon 450 -880 450 -880 0 1
rlabel polysilicon 450 -886 450 -886 0 3
rlabel polysilicon 457 -880 457 -880 0 1
rlabel polysilicon 457 -886 457 -886 0 3
rlabel polysilicon 464 -880 464 -880 0 1
rlabel polysilicon 467 -880 467 -880 0 2
rlabel polysilicon 467 -886 467 -886 0 4
rlabel polysilicon 471 -880 471 -880 0 1
rlabel polysilicon 471 -886 471 -886 0 3
rlabel polysilicon 478 -880 478 -880 0 1
rlabel polysilicon 478 -886 478 -886 0 3
rlabel polysilicon 485 -880 485 -880 0 1
rlabel polysilicon 485 -886 485 -886 0 3
rlabel polysilicon 492 -880 492 -880 0 1
rlabel polysilicon 492 -886 492 -886 0 3
rlabel polysilicon 499 -886 499 -886 0 3
rlabel polysilicon 502 -886 502 -886 0 4
rlabel polysilicon 506 -880 506 -880 0 1
rlabel polysilicon 506 -886 506 -886 0 3
rlabel polysilicon 513 -880 513 -880 0 1
rlabel polysilicon 513 -886 513 -886 0 3
rlabel polysilicon 520 -880 520 -880 0 1
rlabel polysilicon 523 -880 523 -880 0 2
rlabel polysilicon 520 -886 520 -886 0 3
rlabel polysilicon 523 -886 523 -886 0 4
rlabel polysilicon 527 -880 527 -880 0 1
rlabel polysilicon 527 -886 527 -886 0 3
rlabel polysilicon 534 -880 534 -880 0 1
rlabel polysilicon 537 -880 537 -880 0 2
rlabel polysilicon 534 -886 534 -886 0 3
rlabel polysilicon 537 -886 537 -886 0 4
rlabel polysilicon 541 -880 541 -880 0 1
rlabel polysilicon 544 -880 544 -880 0 2
rlabel polysilicon 548 -880 548 -880 0 1
rlabel polysilicon 551 -880 551 -880 0 2
rlabel polysilicon 548 -886 548 -886 0 3
rlabel polysilicon 551 -886 551 -886 0 4
rlabel polysilicon 555 -880 555 -880 0 1
rlabel polysilicon 555 -886 555 -886 0 3
rlabel polysilicon 562 -880 562 -880 0 1
rlabel polysilicon 565 -880 565 -880 0 2
rlabel polysilicon 562 -886 562 -886 0 3
rlabel polysilicon 572 -880 572 -880 0 2
rlabel polysilicon 569 -886 569 -886 0 3
rlabel polysilicon 572 -886 572 -886 0 4
rlabel polysilicon 576 -880 576 -880 0 1
rlabel polysilicon 576 -886 576 -886 0 3
rlabel polysilicon 583 -880 583 -880 0 1
rlabel polysilicon 583 -886 583 -886 0 3
rlabel polysilicon 590 -880 590 -880 0 1
rlabel polysilicon 590 -886 590 -886 0 3
rlabel polysilicon 597 -880 597 -880 0 1
rlabel polysilicon 597 -886 597 -886 0 3
rlabel polysilicon 604 -880 604 -880 0 1
rlabel polysilicon 604 -886 604 -886 0 3
rlabel polysilicon 611 -880 611 -880 0 1
rlabel polysilicon 611 -886 611 -886 0 3
rlabel polysilicon 618 -880 618 -880 0 1
rlabel polysilicon 618 -886 618 -886 0 3
rlabel polysilicon 625 -880 625 -880 0 1
rlabel polysilicon 625 -886 625 -886 0 3
rlabel polysilicon 632 -880 632 -880 0 1
rlabel polysilicon 632 -886 632 -886 0 3
rlabel polysilicon 639 -880 639 -880 0 1
rlabel polysilicon 639 -886 639 -886 0 3
rlabel polysilicon 646 -880 646 -880 0 1
rlabel polysilicon 646 -886 646 -886 0 3
rlabel polysilicon 653 -880 653 -880 0 1
rlabel polysilicon 653 -886 653 -886 0 3
rlabel polysilicon 660 -880 660 -880 0 1
rlabel polysilicon 660 -886 660 -886 0 3
rlabel polysilicon 667 -880 667 -880 0 1
rlabel polysilicon 670 -880 670 -880 0 2
rlabel polysilicon 674 -880 674 -880 0 1
rlabel polysilicon 674 -886 674 -886 0 3
rlabel polysilicon 681 -880 681 -880 0 1
rlabel polysilicon 681 -886 681 -886 0 3
rlabel polysilicon 688 -880 688 -880 0 1
rlabel polysilicon 688 -886 688 -886 0 3
rlabel polysilicon 695 -880 695 -880 0 1
rlabel polysilicon 695 -886 695 -886 0 3
rlabel polysilicon 702 -880 702 -880 0 1
rlabel polysilicon 702 -886 702 -886 0 3
rlabel polysilicon 709 -880 709 -880 0 1
rlabel polysilicon 709 -886 709 -886 0 3
rlabel polysilicon 716 -880 716 -880 0 1
rlabel polysilicon 716 -886 716 -886 0 3
rlabel polysilicon 723 -880 723 -880 0 1
rlabel polysilicon 723 -886 723 -886 0 3
rlabel polysilicon 730 -880 730 -880 0 1
rlabel polysilicon 730 -886 730 -886 0 3
rlabel polysilicon 737 -880 737 -880 0 1
rlabel polysilicon 737 -886 737 -886 0 3
rlabel polysilicon 744 -880 744 -880 0 1
rlabel polysilicon 744 -886 744 -886 0 3
rlabel polysilicon 751 -880 751 -880 0 1
rlabel polysilicon 751 -886 751 -886 0 3
rlabel polysilicon 758 -880 758 -880 0 1
rlabel polysilicon 758 -886 758 -886 0 3
rlabel polysilicon 765 -880 765 -880 0 1
rlabel polysilicon 765 -886 765 -886 0 3
rlabel polysilicon 772 -880 772 -880 0 1
rlabel polysilicon 772 -886 772 -886 0 3
rlabel polysilicon 779 -880 779 -880 0 1
rlabel polysilicon 779 -886 779 -886 0 3
rlabel polysilicon 786 -880 786 -880 0 1
rlabel polysilicon 786 -886 786 -886 0 3
rlabel polysilicon 793 -880 793 -880 0 1
rlabel polysilicon 793 -886 793 -886 0 3
rlabel polysilicon 800 -880 800 -880 0 1
rlabel polysilicon 800 -886 800 -886 0 3
rlabel polysilicon 807 -880 807 -880 0 1
rlabel polysilicon 807 -886 807 -886 0 3
rlabel polysilicon 814 -880 814 -880 0 1
rlabel polysilicon 817 -880 817 -880 0 2
rlabel polysilicon 817 -886 817 -886 0 4
rlabel polysilicon 821 -880 821 -880 0 1
rlabel polysilicon 821 -886 821 -886 0 3
rlabel polysilicon 828 -880 828 -880 0 1
rlabel polysilicon 828 -886 828 -886 0 3
rlabel polysilicon 835 -880 835 -880 0 1
rlabel polysilicon 835 -886 835 -886 0 3
rlabel polysilicon 842 -880 842 -880 0 1
rlabel polysilicon 842 -886 842 -886 0 3
rlabel polysilicon 849 -880 849 -880 0 1
rlabel polysilicon 849 -886 849 -886 0 3
rlabel polysilicon 856 -880 856 -880 0 1
rlabel polysilicon 856 -886 856 -886 0 3
rlabel polysilicon 863 -880 863 -880 0 1
rlabel polysilicon 863 -886 863 -886 0 3
rlabel polysilicon 870 -880 870 -880 0 1
rlabel polysilicon 870 -886 870 -886 0 3
rlabel polysilicon 877 -880 877 -880 0 1
rlabel polysilicon 877 -886 877 -886 0 3
rlabel polysilicon 884 -880 884 -880 0 1
rlabel polysilicon 884 -886 884 -886 0 3
rlabel polysilicon 891 -880 891 -880 0 1
rlabel polysilicon 891 -886 891 -886 0 3
rlabel polysilicon 898 -880 898 -880 0 1
rlabel polysilicon 898 -886 898 -886 0 3
rlabel polysilicon 905 -880 905 -880 0 1
rlabel polysilicon 905 -886 905 -886 0 3
rlabel polysilicon 912 -880 912 -880 0 1
rlabel polysilicon 912 -886 912 -886 0 3
rlabel polysilicon 919 -880 919 -880 0 1
rlabel polysilicon 919 -886 919 -886 0 3
rlabel polysilicon 926 -880 926 -880 0 1
rlabel polysilicon 926 -886 926 -886 0 3
rlabel polysilicon 933 -880 933 -880 0 1
rlabel polysilicon 933 -886 933 -886 0 3
rlabel polysilicon 940 -880 940 -880 0 1
rlabel polysilicon 940 -886 940 -886 0 3
rlabel polysilicon 947 -880 947 -880 0 1
rlabel polysilicon 947 -886 947 -886 0 3
rlabel polysilicon 954 -880 954 -880 0 1
rlabel polysilicon 954 -886 954 -886 0 3
rlabel polysilicon 961 -880 961 -880 0 1
rlabel polysilicon 961 -886 961 -886 0 3
rlabel polysilicon 968 -880 968 -880 0 1
rlabel polysilicon 968 -886 968 -886 0 3
rlabel polysilicon 975 -880 975 -880 0 1
rlabel polysilicon 975 -886 975 -886 0 3
rlabel polysilicon 982 -880 982 -880 0 1
rlabel polysilicon 982 -886 982 -886 0 3
rlabel polysilicon 989 -880 989 -880 0 1
rlabel polysilicon 992 -880 992 -880 0 2
rlabel polysilicon 989 -886 989 -886 0 3
rlabel polysilicon 992 -886 992 -886 0 4
rlabel polysilicon 996 -880 996 -880 0 1
rlabel polysilicon 996 -886 996 -886 0 3
rlabel polysilicon 1003 -880 1003 -880 0 1
rlabel polysilicon 1003 -886 1003 -886 0 3
rlabel polysilicon 1013 -880 1013 -880 0 2
rlabel polysilicon 1010 -886 1010 -886 0 3
rlabel polysilicon 1013 -886 1013 -886 0 4
rlabel polysilicon 1017 -880 1017 -880 0 1
rlabel polysilicon 1017 -886 1017 -886 0 3
rlabel polysilicon 1024 -880 1024 -880 0 1
rlabel polysilicon 1024 -886 1024 -886 0 3
rlabel polysilicon 1038 -880 1038 -880 0 1
rlabel polysilicon 1038 -886 1038 -886 0 3
rlabel polysilicon 1080 -880 1080 -880 0 1
rlabel polysilicon 1080 -886 1080 -886 0 3
rlabel polysilicon 12 -967 12 -967 0 4
rlabel polysilicon 16 -961 16 -961 0 1
rlabel polysilicon 16 -967 16 -967 0 3
rlabel polysilicon 23 -961 23 -961 0 1
rlabel polysilicon 23 -967 23 -967 0 3
rlabel polysilicon 30 -961 30 -961 0 1
rlabel polysilicon 30 -967 30 -967 0 3
rlabel polysilicon 37 -961 37 -961 0 1
rlabel polysilicon 37 -967 37 -967 0 3
rlabel polysilicon 44 -961 44 -961 0 1
rlabel polysilicon 44 -967 44 -967 0 3
rlabel polysilicon 51 -961 51 -961 0 1
rlabel polysilicon 51 -967 51 -967 0 3
rlabel polysilicon 58 -961 58 -961 0 1
rlabel polysilicon 58 -967 58 -967 0 3
rlabel polysilicon 65 -961 65 -961 0 1
rlabel polysilicon 65 -967 65 -967 0 3
rlabel polysilicon 72 -961 72 -961 0 1
rlabel polysilicon 72 -967 72 -967 0 3
rlabel polysilicon 79 -961 79 -961 0 1
rlabel polysilicon 79 -967 79 -967 0 3
rlabel polysilicon 86 -961 86 -961 0 1
rlabel polysilicon 86 -967 86 -967 0 3
rlabel polysilicon 93 -961 93 -961 0 1
rlabel polysilicon 93 -967 93 -967 0 3
rlabel polysilicon 100 -961 100 -961 0 1
rlabel polysilicon 100 -967 100 -967 0 3
rlabel polysilicon 107 -961 107 -961 0 1
rlabel polysilicon 107 -967 107 -967 0 3
rlabel polysilicon 114 -961 114 -961 0 1
rlabel polysilicon 114 -967 114 -967 0 3
rlabel polysilicon 121 -961 121 -961 0 1
rlabel polysilicon 121 -967 121 -967 0 3
rlabel polysilicon 128 -967 128 -967 0 3
rlabel polysilicon 131 -967 131 -967 0 4
rlabel polysilicon 135 -961 135 -961 0 1
rlabel polysilicon 135 -967 135 -967 0 3
rlabel polysilicon 142 -961 142 -961 0 1
rlabel polysilicon 142 -967 142 -967 0 3
rlabel polysilicon 149 -961 149 -961 0 1
rlabel polysilicon 149 -967 149 -967 0 3
rlabel polysilicon 156 -961 156 -961 0 1
rlabel polysilicon 156 -967 156 -967 0 3
rlabel polysilicon 163 -961 163 -961 0 1
rlabel polysilicon 163 -967 163 -967 0 3
rlabel polysilicon 170 -961 170 -961 0 1
rlabel polysilicon 170 -967 170 -967 0 3
rlabel polysilicon 180 -961 180 -961 0 2
rlabel polysilicon 177 -967 177 -967 0 3
rlabel polysilicon 180 -967 180 -967 0 4
rlabel polysilicon 184 -961 184 -961 0 1
rlabel polysilicon 184 -967 184 -967 0 3
rlabel polysilicon 191 -961 191 -961 0 1
rlabel polysilicon 191 -967 191 -967 0 3
rlabel polysilicon 198 -961 198 -961 0 1
rlabel polysilicon 198 -967 198 -967 0 3
rlabel polysilicon 205 -961 205 -961 0 1
rlabel polysilicon 205 -967 205 -967 0 3
rlabel polysilicon 212 -961 212 -961 0 1
rlabel polysilicon 215 -961 215 -961 0 2
rlabel polysilicon 219 -961 219 -961 0 1
rlabel polysilicon 222 -961 222 -961 0 2
rlabel polysilicon 222 -967 222 -967 0 4
rlabel polysilicon 226 -961 226 -961 0 1
rlabel polysilicon 226 -967 226 -967 0 3
rlabel polysilicon 233 -961 233 -961 0 1
rlabel polysilicon 236 -961 236 -961 0 2
rlabel polysilicon 240 -961 240 -961 0 1
rlabel polysilicon 240 -967 240 -967 0 3
rlabel polysilicon 243 -967 243 -967 0 4
rlabel polysilicon 247 -961 247 -961 0 1
rlabel polysilicon 247 -967 247 -967 0 3
rlabel polysilicon 254 -961 254 -961 0 1
rlabel polysilicon 254 -967 254 -967 0 3
rlabel polysilicon 261 -961 261 -961 0 1
rlabel polysilicon 261 -967 261 -967 0 3
rlabel polysilicon 268 -961 268 -961 0 1
rlabel polysilicon 268 -967 268 -967 0 3
rlabel polysilicon 275 -961 275 -961 0 1
rlabel polysilicon 278 -961 278 -961 0 2
rlabel polysilicon 282 -961 282 -961 0 1
rlabel polysilicon 285 -961 285 -961 0 2
rlabel polysilicon 285 -967 285 -967 0 4
rlabel polysilicon 289 -961 289 -961 0 1
rlabel polysilicon 289 -967 289 -967 0 3
rlabel polysilicon 296 -961 296 -961 0 1
rlabel polysilicon 296 -967 296 -967 0 3
rlabel polysilicon 303 -961 303 -961 0 1
rlabel polysilicon 303 -967 303 -967 0 3
rlabel polysilicon 310 -961 310 -961 0 1
rlabel polysilicon 310 -967 310 -967 0 3
rlabel polysilicon 317 -961 317 -961 0 1
rlabel polysilicon 317 -967 317 -967 0 3
rlabel polysilicon 324 -961 324 -961 0 1
rlabel polysilicon 324 -967 324 -967 0 3
rlabel polysilicon 327 -967 327 -967 0 4
rlabel polysilicon 331 -961 331 -961 0 1
rlabel polysilicon 331 -967 331 -967 0 3
rlabel polysilicon 338 -961 338 -961 0 1
rlabel polysilicon 338 -967 338 -967 0 3
rlabel polysilicon 345 -961 345 -961 0 1
rlabel polysilicon 345 -967 345 -967 0 3
rlabel polysilicon 352 -961 352 -961 0 1
rlabel polysilicon 352 -967 352 -967 0 3
rlabel polysilicon 359 -961 359 -961 0 1
rlabel polysilicon 359 -967 359 -967 0 3
rlabel polysilicon 362 -967 362 -967 0 4
rlabel polysilicon 366 -961 366 -961 0 1
rlabel polysilicon 366 -967 366 -967 0 3
rlabel polysilicon 373 -961 373 -961 0 1
rlabel polysilicon 373 -967 373 -967 0 3
rlabel polysilicon 380 -967 380 -967 0 3
rlabel polysilicon 383 -967 383 -967 0 4
rlabel polysilicon 387 -961 387 -961 0 1
rlabel polysilicon 387 -967 387 -967 0 3
rlabel polysilicon 397 -967 397 -967 0 4
rlabel polysilicon 401 -961 401 -961 0 1
rlabel polysilicon 401 -967 401 -967 0 3
rlabel polysilicon 408 -961 408 -961 0 1
rlabel polysilicon 408 -967 408 -967 0 3
rlabel polysilicon 415 -961 415 -961 0 1
rlabel polysilicon 418 -961 418 -961 0 2
rlabel polysilicon 418 -967 418 -967 0 4
rlabel polysilicon 422 -961 422 -961 0 1
rlabel polysilicon 422 -967 422 -967 0 3
rlabel polysilicon 429 -961 429 -961 0 1
rlabel polysilicon 429 -967 429 -967 0 3
rlabel polysilicon 439 -961 439 -961 0 2
rlabel polysilicon 436 -967 436 -967 0 3
rlabel polysilicon 439 -967 439 -967 0 4
rlabel polysilicon 443 -961 443 -961 0 1
rlabel polysilicon 443 -967 443 -967 0 3
rlabel polysilicon 450 -967 450 -967 0 3
rlabel polysilicon 453 -967 453 -967 0 4
rlabel polysilicon 457 -961 457 -961 0 1
rlabel polysilicon 457 -967 457 -967 0 3
rlabel polysilicon 464 -961 464 -961 0 1
rlabel polysilicon 464 -967 464 -967 0 3
rlabel polysilicon 471 -961 471 -961 0 1
rlabel polysilicon 474 -961 474 -961 0 2
rlabel polysilicon 471 -967 471 -967 0 3
rlabel polysilicon 474 -967 474 -967 0 4
rlabel polysilicon 478 -961 478 -961 0 1
rlabel polysilicon 478 -967 478 -967 0 3
rlabel polysilicon 481 -967 481 -967 0 4
rlabel polysilicon 485 -961 485 -961 0 1
rlabel polysilicon 485 -967 485 -967 0 3
rlabel polysilicon 492 -961 492 -961 0 1
rlabel polysilicon 492 -967 492 -967 0 3
rlabel polysilicon 495 -967 495 -967 0 4
rlabel polysilicon 499 -961 499 -961 0 1
rlabel polysilicon 499 -967 499 -967 0 3
rlabel polysilicon 506 -961 506 -961 0 1
rlabel polysilicon 506 -967 506 -967 0 3
rlabel polysilicon 513 -961 513 -961 0 1
rlabel polysilicon 520 -961 520 -961 0 1
rlabel polysilicon 520 -967 520 -967 0 3
rlabel polysilicon 530 -961 530 -961 0 2
rlabel polysilicon 530 -967 530 -967 0 4
rlabel polysilicon 534 -961 534 -961 0 1
rlabel polysilicon 534 -967 534 -967 0 3
rlabel polysilicon 541 -961 541 -961 0 1
rlabel polysilicon 541 -967 541 -967 0 3
rlabel polysilicon 548 -961 548 -961 0 1
rlabel polysilicon 548 -967 548 -967 0 3
rlabel polysilicon 555 -961 555 -961 0 1
rlabel polysilicon 555 -967 555 -967 0 3
rlabel polysilicon 562 -961 562 -961 0 1
rlabel polysilicon 562 -967 562 -967 0 3
rlabel polysilicon 565 -967 565 -967 0 4
rlabel polysilicon 569 -961 569 -961 0 1
rlabel polysilicon 569 -967 569 -967 0 3
rlabel polysilicon 576 -961 576 -961 0 1
rlabel polysilicon 576 -967 576 -967 0 3
rlabel polysilicon 583 -961 583 -961 0 1
rlabel polysilicon 583 -967 583 -967 0 3
rlabel polysilicon 590 -961 590 -961 0 1
rlabel polysilicon 590 -967 590 -967 0 3
rlabel polysilicon 597 -961 597 -961 0 1
rlabel polysilicon 600 -961 600 -961 0 2
rlabel polysilicon 597 -967 597 -967 0 3
rlabel polysilicon 600 -967 600 -967 0 4
rlabel polysilicon 604 -961 604 -961 0 1
rlabel polysilicon 604 -967 604 -967 0 3
rlabel polysilicon 607 -967 607 -967 0 4
rlabel polysilicon 611 -961 611 -961 0 1
rlabel polysilicon 611 -967 611 -967 0 3
rlabel polysilicon 618 -961 618 -961 0 1
rlabel polysilicon 618 -967 618 -967 0 3
rlabel polysilicon 628 -961 628 -961 0 2
rlabel polysilicon 625 -967 625 -967 0 3
rlabel polysilicon 635 -961 635 -961 0 2
rlabel polysilicon 632 -967 632 -967 0 3
rlabel polysilicon 635 -967 635 -967 0 4
rlabel polysilicon 639 -961 639 -961 0 1
rlabel polysilicon 639 -967 639 -967 0 3
rlabel polysilicon 646 -961 646 -961 0 1
rlabel polysilicon 646 -967 646 -967 0 3
rlabel polysilicon 656 -961 656 -961 0 2
rlabel polysilicon 653 -967 653 -967 0 3
rlabel polysilicon 660 -961 660 -961 0 1
rlabel polysilicon 660 -967 660 -967 0 3
rlabel polysilicon 667 -961 667 -961 0 1
rlabel polysilicon 667 -967 667 -967 0 3
rlabel polysilicon 674 -961 674 -961 0 1
rlabel polysilicon 674 -967 674 -967 0 3
rlabel polysilicon 681 -961 681 -961 0 1
rlabel polysilicon 681 -967 681 -967 0 3
rlabel polysilicon 688 -961 688 -961 0 1
rlabel polysilicon 688 -967 688 -967 0 3
rlabel polysilicon 695 -961 695 -961 0 1
rlabel polysilicon 695 -967 695 -967 0 3
rlabel polysilicon 698 -967 698 -967 0 4
rlabel polysilicon 702 -961 702 -961 0 1
rlabel polysilicon 702 -967 702 -967 0 3
rlabel polysilicon 709 -961 709 -961 0 1
rlabel polysilicon 709 -967 709 -967 0 3
rlabel polysilicon 716 -961 716 -961 0 1
rlabel polysilicon 716 -967 716 -967 0 3
rlabel polysilicon 723 -961 723 -961 0 1
rlabel polysilicon 723 -967 723 -967 0 3
rlabel polysilicon 730 -961 730 -961 0 1
rlabel polysilicon 730 -967 730 -967 0 3
rlabel polysilicon 737 -961 737 -961 0 1
rlabel polysilicon 737 -967 737 -967 0 3
rlabel polysilicon 744 -961 744 -961 0 1
rlabel polysilicon 744 -967 744 -967 0 3
rlabel polysilicon 751 -961 751 -961 0 1
rlabel polysilicon 751 -967 751 -967 0 3
rlabel polysilicon 758 -961 758 -961 0 1
rlabel polysilicon 758 -967 758 -967 0 3
rlabel polysilicon 765 -961 765 -961 0 1
rlabel polysilicon 765 -967 765 -967 0 3
rlabel polysilicon 772 -961 772 -961 0 1
rlabel polysilicon 772 -967 772 -967 0 3
rlabel polysilicon 779 -961 779 -961 0 1
rlabel polysilicon 779 -967 779 -967 0 3
rlabel polysilicon 786 -961 786 -961 0 1
rlabel polysilicon 786 -967 786 -967 0 3
rlabel polysilicon 793 -961 793 -961 0 1
rlabel polysilicon 793 -967 793 -967 0 3
rlabel polysilicon 800 -961 800 -961 0 1
rlabel polysilicon 800 -967 800 -967 0 3
rlabel polysilicon 807 -961 807 -961 0 1
rlabel polysilicon 807 -967 807 -967 0 3
rlabel polysilicon 814 -961 814 -961 0 1
rlabel polysilicon 814 -967 814 -967 0 3
rlabel polysilicon 821 -961 821 -961 0 1
rlabel polysilicon 821 -967 821 -967 0 3
rlabel polysilicon 828 -961 828 -961 0 1
rlabel polysilicon 828 -967 828 -967 0 3
rlabel polysilicon 835 -961 835 -961 0 1
rlabel polysilicon 835 -967 835 -967 0 3
rlabel polysilicon 842 -961 842 -961 0 1
rlabel polysilicon 842 -967 842 -967 0 3
rlabel polysilicon 849 -961 849 -961 0 1
rlabel polysilicon 849 -967 849 -967 0 3
rlabel polysilicon 856 -961 856 -961 0 1
rlabel polysilicon 856 -967 856 -967 0 3
rlabel polysilicon 863 -961 863 -961 0 1
rlabel polysilicon 863 -967 863 -967 0 3
rlabel polysilicon 870 -961 870 -961 0 1
rlabel polysilicon 870 -967 870 -967 0 3
rlabel polysilicon 877 -961 877 -961 0 1
rlabel polysilicon 877 -967 877 -967 0 3
rlabel polysilicon 884 -961 884 -961 0 1
rlabel polysilicon 884 -967 884 -967 0 3
rlabel polysilicon 891 -961 891 -961 0 1
rlabel polysilicon 891 -967 891 -967 0 3
rlabel polysilicon 898 -961 898 -961 0 1
rlabel polysilicon 898 -967 898 -967 0 3
rlabel polysilicon 905 -961 905 -961 0 1
rlabel polysilicon 905 -967 905 -967 0 3
rlabel polysilicon 912 -961 912 -961 0 1
rlabel polysilicon 915 -961 915 -961 0 2
rlabel polysilicon 915 -967 915 -967 0 4
rlabel polysilicon 922 -961 922 -961 0 2
rlabel polysilicon 919 -967 919 -967 0 3
rlabel polysilicon 922 -967 922 -967 0 4
rlabel polysilicon 929 -961 929 -961 0 2
rlabel polysilicon 926 -967 926 -967 0 3
rlabel polysilicon 929 -967 929 -967 0 4
rlabel polysilicon 933 -961 933 -961 0 1
rlabel polysilicon 933 -967 933 -967 0 3
rlabel polysilicon 943 -961 943 -961 0 2
rlabel polysilicon 943 -967 943 -967 0 4
rlabel polysilicon 947 -961 947 -961 0 1
rlabel polysilicon 947 -967 947 -967 0 3
rlabel polysilicon 954 -961 954 -961 0 1
rlabel polysilicon 954 -967 954 -967 0 3
rlabel polysilicon 961 -961 961 -961 0 1
rlabel polysilicon 961 -967 961 -967 0 3
rlabel polysilicon 968 -961 968 -961 0 1
rlabel polysilicon 968 -967 968 -967 0 3
rlabel polysilicon 982 -961 982 -961 0 1
rlabel polysilicon 982 -967 982 -967 0 3
rlabel polysilicon 1010 -961 1010 -961 0 1
rlabel polysilicon 1010 -967 1010 -967 0 3
rlabel polysilicon 1038 -961 1038 -961 0 1
rlabel polysilicon 1038 -967 1038 -967 0 3
rlabel polysilicon 1059 -961 1059 -961 0 1
rlabel polysilicon 1059 -967 1059 -967 0 3
rlabel polysilicon 1087 -961 1087 -961 0 1
rlabel polysilicon 1087 -967 1087 -967 0 3
rlabel polysilicon 9 -1054 9 -1054 0 1
rlabel polysilicon 9 -1060 9 -1060 0 3
rlabel polysilicon 16 -1054 16 -1054 0 1
rlabel polysilicon 16 -1060 16 -1060 0 3
rlabel polysilicon 23 -1054 23 -1054 0 1
rlabel polysilicon 23 -1060 23 -1060 0 3
rlabel polysilicon 30 -1054 30 -1054 0 1
rlabel polysilicon 30 -1060 30 -1060 0 3
rlabel polysilicon 40 -1054 40 -1054 0 2
rlabel polysilicon 44 -1054 44 -1054 0 1
rlabel polysilicon 44 -1060 44 -1060 0 3
rlabel polysilicon 51 -1054 51 -1054 0 1
rlabel polysilicon 51 -1060 51 -1060 0 3
rlabel polysilicon 61 -1054 61 -1054 0 2
rlabel polysilicon 58 -1060 58 -1060 0 3
rlabel polysilicon 65 -1054 65 -1054 0 1
rlabel polysilicon 65 -1060 65 -1060 0 3
rlabel polysilicon 72 -1054 72 -1054 0 1
rlabel polysilicon 72 -1060 72 -1060 0 3
rlabel polysilicon 79 -1054 79 -1054 0 1
rlabel polysilicon 79 -1060 79 -1060 0 3
rlabel polysilicon 86 -1054 86 -1054 0 1
rlabel polysilicon 86 -1060 86 -1060 0 3
rlabel polysilicon 93 -1054 93 -1054 0 1
rlabel polysilicon 93 -1060 93 -1060 0 3
rlabel polysilicon 100 -1054 100 -1054 0 1
rlabel polysilicon 100 -1060 100 -1060 0 3
rlabel polysilicon 107 -1054 107 -1054 0 1
rlabel polysilicon 107 -1060 107 -1060 0 3
rlabel polysilicon 114 -1054 114 -1054 0 1
rlabel polysilicon 114 -1060 114 -1060 0 3
rlabel polysilicon 121 -1054 121 -1054 0 1
rlabel polysilicon 121 -1060 121 -1060 0 3
rlabel polysilicon 131 -1054 131 -1054 0 2
rlabel polysilicon 135 -1054 135 -1054 0 1
rlabel polysilicon 135 -1060 135 -1060 0 3
rlabel polysilicon 142 -1054 142 -1054 0 1
rlabel polysilicon 145 -1054 145 -1054 0 2
rlabel polysilicon 142 -1060 142 -1060 0 3
rlabel polysilicon 149 -1054 149 -1054 0 1
rlabel polysilicon 149 -1060 149 -1060 0 3
rlabel polysilicon 156 -1054 156 -1054 0 1
rlabel polysilicon 156 -1060 156 -1060 0 3
rlabel polysilicon 163 -1054 163 -1054 0 1
rlabel polysilicon 166 -1060 166 -1060 0 4
rlabel polysilicon 170 -1060 170 -1060 0 3
rlabel polysilicon 173 -1060 173 -1060 0 4
rlabel polysilicon 180 -1054 180 -1054 0 2
rlabel polysilicon 180 -1060 180 -1060 0 4
rlabel polysilicon 184 -1054 184 -1054 0 1
rlabel polysilicon 184 -1060 184 -1060 0 3
rlabel polysilicon 191 -1054 191 -1054 0 1
rlabel polysilicon 191 -1060 191 -1060 0 3
rlabel polysilicon 198 -1054 198 -1054 0 1
rlabel polysilicon 198 -1060 198 -1060 0 3
rlabel polysilicon 205 -1054 205 -1054 0 1
rlabel polysilicon 208 -1054 208 -1054 0 2
rlabel polysilicon 205 -1060 205 -1060 0 3
rlabel polysilicon 212 -1054 212 -1054 0 1
rlabel polysilicon 219 -1054 219 -1054 0 1
rlabel polysilicon 222 -1060 222 -1060 0 4
rlabel polysilicon 226 -1054 226 -1054 0 1
rlabel polysilicon 226 -1060 226 -1060 0 3
rlabel polysilicon 233 -1054 233 -1054 0 1
rlabel polysilicon 233 -1060 233 -1060 0 3
rlabel polysilicon 240 -1054 240 -1054 0 1
rlabel polysilicon 240 -1060 240 -1060 0 3
rlabel polysilicon 247 -1054 247 -1054 0 1
rlabel polysilicon 247 -1060 247 -1060 0 3
rlabel polysilicon 257 -1054 257 -1054 0 2
rlabel polysilicon 261 -1054 261 -1054 0 1
rlabel polysilicon 261 -1060 261 -1060 0 3
rlabel polysilicon 268 -1054 268 -1054 0 1
rlabel polysilicon 268 -1060 268 -1060 0 3
rlabel polysilicon 275 -1054 275 -1054 0 1
rlabel polysilicon 275 -1060 275 -1060 0 3
rlabel polysilicon 282 -1054 282 -1054 0 1
rlabel polysilicon 282 -1060 282 -1060 0 3
rlabel polysilicon 289 -1054 289 -1054 0 1
rlabel polysilicon 289 -1060 289 -1060 0 3
rlabel polysilicon 296 -1054 296 -1054 0 1
rlabel polysilicon 299 -1054 299 -1054 0 2
rlabel polysilicon 299 -1060 299 -1060 0 4
rlabel polysilicon 303 -1054 303 -1054 0 1
rlabel polysilicon 303 -1060 303 -1060 0 3
rlabel polysilicon 310 -1054 310 -1054 0 1
rlabel polysilicon 310 -1060 310 -1060 0 3
rlabel polysilicon 317 -1054 317 -1054 0 1
rlabel polysilicon 317 -1060 317 -1060 0 3
rlabel polysilicon 324 -1054 324 -1054 0 1
rlabel polysilicon 324 -1060 324 -1060 0 3
rlabel polysilicon 331 -1054 331 -1054 0 1
rlabel polysilicon 331 -1060 331 -1060 0 3
rlabel polysilicon 338 -1054 338 -1054 0 1
rlabel polysilicon 338 -1060 338 -1060 0 3
rlabel polysilicon 345 -1054 345 -1054 0 1
rlabel polysilicon 345 -1060 345 -1060 0 3
rlabel polysilicon 352 -1054 352 -1054 0 1
rlabel polysilicon 355 -1054 355 -1054 0 2
rlabel polysilicon 352 -1060 352 -1060 0 3
rlabel polysilicon 355 -1060 355 -1060 0 4
rlabel polysilicon 359 -1054 359 -1054 0 1
rlabel polysilicon 359 -1060 359 -1060 0 3
rlabel polysilicon 366 -1054 366 -1054 0 1
rlabel polysilicon 366 -1060 366 -1060 0 3
rlabel polysilicon 373 -1054 373 -1054 0 1
rlabel polysilicon 373 -1060 373 -1060 0 3
rlabel polysilicon 380 -1054 380 -1054 0 1
rlabel polysilicon 380 -1060 380 -1060 0 3
rlabel polysilicon 387 -1054 387 -1054 0 1
rlabel polysilicon 387 -1060 387 -1060 0 3
rlabel polysilicon 394 -1054 394 -1054 0 1
rlabel polysilicon 394 -1060 394 -1060 0 3
rlabel polysilicon 401 -1054 401 -1054 0 1
rlabel polysilicon 401 -1060 401 -1060 0 3
rlabel polysilicon 411 -1054 411 -1054 0 2
rlabel polysilicon 408 -1060 408 -1060 0 3
rlabel polysilicon 411 -1060 411 -1060 0 4
rlabel polysilicon 415 -1054 415 -1054 0 1
rlabel polysilicon 415 -1060 415 -1060 0 3
rlabel polysilicon 422 -1054 422 -1054 0 1
rlabel polysilicon 422 -1060 422 -1060 0 3
rlabel polysilicon 429 -1054 429 -1054 0 1
rlabel polysilicon 432 -1054 432 -1054 0 2
rlabel polysilicon 429 -1060 429 -1060 0 3
rlabel polysilicon 436 -1054 436 -1054 0 1
rlabel polysilicon 436 -1060 436 -1060 0 3
rlabel polysilicon 443 -1054 443 -1054 0 1
rlabel polysilicon 446 -1054 446 -1054 0 2
rlabel polysilicon 443 -1060 443 -1060 0 3
rlabel polysilicon 446 -1060 446 -1060 0 4
rlabel polysilicon 450 -1054 450 -1054 0 1
rlabel polysilicon 453 -1054 453 -1054 0 2
rlabel polysilicon 453 -1060 453 -1060 0 4
rlabel polysilicon 457 -1054 457 -1054 0 1
rlabel polysilicon 457 -1060 457 -1060 0 3
rlabel polysilicon 464 -1054 464 -1054 0 1
rlabel polysilicon 464 -1060 464 -1060 0 3
rlabel polysilicon 471 -1054 471 -1054 0 1
rlabel polysilicon 474 -1054 474 -1054 0 2
rlabel polysilicon 478 -1054 478 -1054 0 1
rlabel polysilicon 478 -1060 478 -1060 0 3
rlabel polysilicon 488 -1054 488 -1054 0 2
rlabel polysilicon 485 -1060 485 -1060 0 3
rlabel polysilicon 492 -1054 492 -1054 0 1
rlabel polysilicon 492 -1060 492 -1060 0 3
rlabel polysilicon 495 -1060 495 -1060 0 4
rlabel polysilicon 499 -1054 499 -1054 0 1
rlabel polysilicon 499 -1060 499 -1060 0 3
rlabel polysilicon 506 -1054 506 -1054 0 1
rlabel polysilicon 506 -1060 506 -1060 0 3
rlabel polysilicon 516 -1054 516 -1054 0 2
rlabel polysilicon 513 -1060 513 -1060 0 3
rlabel polysilicon 520 -1054 520 -1054 0 1
rlabel polysilicon 520 -1060 520 -1060 0 3
rlabel polysilicon 527 -1054 527 -1054 0 1
rlabel polysilicon 527 -1060 527 -1060 0 3
rlabel polysilicon 537 -1054 537 -1054 0 2
rlabel polysilicon 534 -1060 534 -1060 0 3
rlabel polysilicon 537 -1060 537 -1060 0 4
rlabel polysilicon 541 -1054 541 -1054 0 1
rlabel polysilicon 541 -1060 541 -1060 0 3
rlabel polysilicon 548 -1054 548 -1054 0 1
rlabel polysilicon 551 -1054 551 -1054 0 2
rlabel polysilicon 551 -1060 551 -1060 0 4
rlabel polysilicon 555 -1054 555 -1054 0 1
rlabel polysilicon 555 -1060 555 -1060 0 3
rlabel polysilicon 562 -1054 562 -1054 0 1
rlabel polysilicon 562 -1060 562 -1060 0 3
rlabel polysilicon 569 -1054 569 -1054 0 1
rlabel polysilicon 569 -1060 569 -1060 0 3
rlabel polysilicon 572 -1060 572 -1060 0 4
rlabel polysilicon 576 -1054 576 -1054 0 1
rlabel polysilicon 576 -1060 576 -1060 0 3
rlabel polysilicon 579 -1060 579 -1060 0 4
rlabel polysilicon 583 -1054 583 -1054 0 1
rlabel polysilicon 586 -1054 586 -1054 0 2
rlabel polysilicon 583 -1060 583 -1060 0 3
rlabel polysilicon 590 -1054 590 -1054 0 1
rlabel polysilicon 590 -1060 590 -1060 0 3
rlabel polysilicon 597 -1054 597 -1054 0 1
rlabel polysilicon 597 -1060 597 -1060 0 3
rlabel polysilicon 604 -1054 604 -1054 0 1
rlabel polysilicon 607 -1054 607 -1054 0 2
rlabel polysilicon 611 -1054 611 -1054 0 1
rlabel polysilicon 611 -1060 611 -1060 0 3
rlabel polysilicon 618 -1054 618 -1054 0 1
rlabel polysilicon 618 -1060 618 -1060 0 3
rlabel polysilicon 628 -1054 628 -1054 0 2
rlabel polysilicon 628 -1060 628 -1060 0 4
rlabel polysilicon 632 -1054 632 -1054 0 1
rlabel polysilicon 632 -1060 632 -1060 0 3
rlabel polysilicon 639 -1054 639 -1054 0 1
rlabel polysilicon 639 -1060 639 -1060 0 3
rlabel polysilicon 646 -1054 646 -1054 0 1
rlabel polysilicon 649 -1054 649 -1054 0 2
rlabel polysilicon 646 -1060 646 -1060 0 3
rlabel polysilicon 649 -1060 649 -1060 0 4
rlabel polysilicon 653 -1054 653 -1054 0 1
rlabel polysilicon 653 -1060 653 -1060 0 3
rlabel polysilicon 660 -1054 660 -1054 0 1
rlabel polysilicon 660 -1060 660 -1060 0 3
rlabel polysilicon 667 -1054 667 -1054 0 1
rlabel polysilicon 667 -1060 667 -1060 0 3
rlabel polysilicon 674 -1054 674 -1054 0 1
rlabel polysilicon 674 -1060 674 -1060 0 3
rlabel polysilicon 681 -1054 681 -1054 0 1
rlabel polysilicon 681 -1060 681 -1060 0 3
rlabel polysilicon 691 -1054 691 -1054 0 2
rlabel polysilicon 688 -1060 688 -1060 0 3
rlabel polysilicon 695 -1054 695 -1054 0 1
rlabel polysilicon 695 -1060 695 -1060 0 3
rlabel polysilicon 702 -1054 702 -1054 0 1
rlabel polysilicon 702 -1060 702 -1060 0 3
rlabel polysilicon 709 -1054 709 -1054 0 1
rlabel polysilicon 709 -1060 709 -1060 0 3
rlabel polysilicon 716 -1054 716 -1054 0 1
rlabel polysilicon 716 -1060 716 -1060 0 3
rlabel polysilicon 723 -1054 723 -1054 0 1
rlabel polysilicon 723 -1060 723 -1060 0 3
rlabel polysilicon 730 -1054 730 -1054 0 1
rlabel polysilicon 733 -1054 733 -1054 0 2
rlabel polysilicon 730 -1060 730 -1060 0 3
rlabel polysilicon 737 -1054 737 -1054 0 1
rlabel polysilicon 737 -1060 737 -1060 0 3
rlabel polysilicon 744 -1054 744 -1054 0 1
rlabel polysilicon 744 -1060 744 -1060 0 3
rlabel polysilicon 751 -1054 751 -1054 0 1
rlabel polysilicon 751 -1060 751 -1060 0 3
rlabel polysilicon 758 -1054 758 -1054 0 1
rlabel polysilicon 758 -1060 758 -1060 0 3
rlabel polysilicon 765 -1054 765 -1054 0 1
rlabel polysilicon 765 -1060 765 -1060 0 3
rlabel polysilicon 772 -1054 772 -1054 0 1
rlabel polysilicon 772 -1060 772 -1060 0 3
rlabel polysilicon 779 -1054 779 -1054 0 1
rlabel polysilicon 779 -1060 779 -1060 0 3
rlabel polysilicon 786 -1054 786 -1054 0 1
rlabel polysilicon 786 -1060 786 -1060 0 3
rlabel polysilicon 793 -1054 793 -1054 0 1
rlabel polysilicon 793 -1060 793 -1060 0 3
rlabel polysilicon 800 -1054 800 -1054 0 1
rlabel polysilicon 800 -1060 800 -1060 0 3
rlabel polysilicon 807 -1054 807 -1054 0 1
rlabel polysilicon 807 -1060 807 -1060 0 3
rlabel polysilicon 814 -1054 814 -1054 0 1
rlabel polysilicon 814 -1060 814 -1060 0 3
rlabel polysilicon 821 -1054 821 -1054 0 1
rlabel polysilicon 821 -1060 821 -1060 0 3
rlabel polysilicon 828 -1054 828 -1054 0 1
rlabel polysilicon 828 -1060 828 -1060 0 3
rlabel polysilicon 835 -1054 835 -1054 0 1
rlabel polysilicon 835 -1060 835 -1060 0 3
rlabel polysilicon 842 -1054 842 -1054 0 1
rlabel polysilicon 842 -1060 842 -1060 0 3
rlabel polysilicon 849 -1054 849 -1054 0 1
rlabel polysilicon 849 -1060 849 -1060 0 3
rlabel polysilicon 856 -1054 856 -1054 0 1
rlabel polysilicon 856 -1060 856 -1060 0 3
rlabel polysilicon 863 -1054 863 -1054 0 1
rlabel polysilicon 863 -1060 863 -1060 0 3
rlabel polysilicon 870 -1054 870 -1054 0 1
rlabel polysilicon 870 -1060 870 -1060 0 3
rlabel polysilicon 877 -1054 877 -1054 0 1
rlabel polysilicon 877 -1060 877 -1060 0 3
rlabel polysilicon 884 -1054 884 -1054 0 1
rlabel polysilicon 884 -1060 884 -1060 0 3
rlabel polysilicon 891 -1054 891 -1054 0 1
rlabel polysilicon 891 -1060 891 -1060 0 3
rlabel polysilicon 898 -1054 898 -1054 0 1
rlabel polysilicon 898 -1060 898 -1060 0 3
rlabel polysilicon 905 -1054 905 -1054 0 1
rlabel polysilicon 905 -1060 905 -1060 0 3
rlabel polysilicon 912 -1054 912 -1054 0 1
rlabel polysilicon 912 -1060 912 -1060 0 3
rlabel polysilicon 919 -1054 919 -1054 0 1
rlabel polysilicon 919 -1060 919 -1060 0 3
rlabel polysilicon 926 -1054 926 -1054 0 1
rlabel polysilicon 926 -1060 926 -1060 0 3
rlabel polysilicon 933 -1054 933 -1054 0 1
rlabel polysilicon 933 -1060 933 -1060 0 3
rlabel polysilicon 940 -1054 940 -1054 0 1
rlabel polysilicon 940 -1060 940 -1060 0 3
rlabel polysilicon 947 -1054 947 -1054 0 1
rlabel polysilicon 947 -1060 947 -1060 0 3
rlabel polysilicon 954 -1054 954 -1054 0 1
rlabel polysilicon 954 -1060 954 -1060 0 3
rlabel polysilicon 961 -1054 961 -1054 0 1
rlabel polysilicon 961 -1060 961 -1060 0 3
rlabel polysilicon 968 -1054 968 -1054 0 1
rlabel polysilicon 968 -1060 968 -1060 0 3
rlabel polysilicon 975 -1054 975 -1054 0 1
rlabel polysilicon 975 -1060 975 -1060 0 3
rlabel polysilicon 982 -1054 982 -1054 0 1
rlabel polysilicon 982 -1060 982 -1060 0 3
rlabel polysilicon 989 -1054 989 -1054 0 1
rlabel polysilicon 989 -1060 989 -1060 0 3
rlabel polysilicon 996 -1054 996 -1054 0 1
rlabel polysilicon 996 -1060 996 -1060 0 3
rlabel polysilicon 1003 -1054 1003 -1054 0 1
rlabel polysilicon 1003 -1060 1003 -1060 0 3
rlabel polysilicon 1010 -1054 1010 -1054 0 1
rlabel polysilicon 1010 -1060 1010 -1060 0 3
rlabel polysilicon 1017 -1054 1017 -1054 0 1
rlabel polysilicon 1017 -1060 1017 -1060 0 3
rlabel polysilicon 1027 -1060 1027 -1060 0 4
rlabel polysilicon 1031 -1054 1031 -1054 0 1
rlabel polysilicon 1031 -1060 1031 -1060 0 3
rlabel polysilicon 1038 -1054 1038 -1054 0 1
rlabel polysilicon 1038 -1060 1038 -1060 0 3
rlabel polysilicon 1045 -1054 1045 -1054 0 1
rlabel polysilicon 1045 -1060 1045 -1060 0 3
rlabel polysilicon 1052 -1054 1052 -1054 0 1
rlabel polysilicon 1052 -1060 1052 -1060 0 3
rlabel polysilicon 1059 -1054 1059 -1054 0 1
rlabel polysilicon 1059 -1060 1059 -1060 0 3
rlabel polysilicon 1066 -1054 1066 -1054 0 1
rlabel polysilicon 1069 -1054 1069 -1054 0 2
rlabel polysilicon 1069 -1060 1069 -1060 0 4
rlabel polysilicon 1073 -1054 1073 -1054 0 1
rlabel polysilicon 1076 -1054 1076 -1054 0 2
rlabel polysilicon 1076 -1060 1076 -1060 0 4
rlabel polysilicon 1080 -1060 1080 -1060 0 3
rlabel polysilicon 1083 -1060 1083 -1060 0 4
rlabel polysilicon 1087 -1054 1087 -1054 0 1
rlabel polysilicon 1087 -1060 1087 -1060 0 3
rlabel polysilicon 1094 -1054 1094 -1054 0 1
rlabel polysilicon 1094 -1060 1094 -1060 0 3
rlabel polysilicon 1097 -1060 1097 -1060 0 4
rlabel polysilicon 1101 -1054 1101 -1054 0 1
rlabel polysilicon 1101 -1060 1101 -1060 0 3
rlabel polysilicon 2 -1153 2 -1153 0 1
rlabel polysilicon 2 -1159 2 -1159 0 3
rlabel polysilicon 9 -1159 9 -1159 0 3
rlabel polysilicon 19 -1153 19 -1153 0 2
rlabel polysilicon 23 -1153 23 -1153 0 1
rlabel polysilicon 23 -1159 23 -1159 0 3
rlabel polysilicon 30 -1159 30 -1159 0 3
rlabel polysilicon 33 -1159 33 -1159 0 4
rlabel polysilicon 37 -1153 37 -1153 0 1
rlabel polysilicon 37 -1159 37 -1159 0 3
rlabel polysilicon 44 -1153 44 -1153 0 1
rlabel polysilicon 44 -1159 44 -1159 0 3
rlabel polysilicon 51 -1153 51 -1153 0 1
rlabel polysilicon 51 -1159 51 -1159 0 3
rlabel polysilicon 58 -1153 58 -1153 0 1
rlabel polysilicon 58 -1159 58 -1159 0 3
rlabel polysilicon 65 -1153 65 -1153 0 1
rlabel polysilicon 65 -1159 65 -1159 0 3
rlabel polysilicon 72 -1153 72 -1153 0 1
rlabel polysilicon 72 -1159 72 -1159 0 3
rlabel polysilicon 79 -1159 79 -1159 0 3
rlabel polysilicon 82 -1159 82 -1159 0 4
rlabel polysilicon 86 -1153 86 -1153 0 1
rlabel polysilicon 86 -1159 86 -1159 0 3
rlabel polysilicon 93 -1153 93 -1153 0 1
rlabel polysilicon 93 -1159 93 -1159 0 3
rlabel polysilicon 100 -1153 100 -1153 0 1
rlabel polysilicon 100 -1159 100 -1159 0 3
rlabel polysilicon 107 -1153 107 -1153 0 1
rlabel polysilicon 107 -1159 107 -1159 0 3
rlabel polysilicon 114 -1153 114 -1153 0 1
rlabel polysilicon 114 -1159 114 -1159 0 3
rlabel polysilicon 121 -1153 121 -1153 0 1
rlabel polysilicon 121 -1159 121 -1159 0 3
rlabel polysilicon 128 -1153 128 -1153 0 1
rlabel polysilicon 131 -1153 131 -1153 0 2
rlabel polysilicon 128 -1159 128 -1159 0 3
rlabel polysilicon 135 -1153 135 -1153 0 1
rlabel polysilicon 135 -1159 135 -1159 0 3
rlabel polysilicon 145 -1153 145 -1153 0 2
rlabel polysilicon 142 -1159 142 -1159 0 3
rlabel polysilicon 149 -1153 149 -1153 0 1
rlabel polysilicon 149 -1159 149 -1159 0 3
rlabel polysilicon 156 -1153 156 -1153 0 1
rlabel polysilicon 156 -1159 156 -1159 0 3
rlabel polysilicon 163 -1153 163 -1153 0 1
rlabel polysilicon 163 -1159 163 -1159 0 3
rlabel polysilicon 170 -1153 170 -1153 0 1
rlabel polysilicon 170 -1159 170 -1159 0 3
rlabel polysilicon 177 -1153 177 -1153 0 1
rlabel polysilicon 177 -1159 177 -1159 0 3
rlabel polysilicon 187 -1153 187 -1153 0 2
rlabel polysilicon 184 -1159 184 -1159 0 3
rlabel polysilicon 187 -1159 187 -1159 0 4
rlabel polysilicon 191 -1153 191 -1153 0 1
rlabel polysilicon 191 -1159 191 -1159 0 3
rlabel polysilicon 198 -1153 198 -1153 0 1
rlabel polysilicon 198 -1159 198 -1159 0 3
rlabel polysilicon 205 -1153 205 -1153 0 1
rlabel polysilicon 205 -1159 205 -1159 0 3
rlabel polysilicon 212 -1159 212 -1159 0 3
rlabel polysilicon 219 -1153 219 -1153 0 1
rlabel polysilicon 219 -1159 219 -1159 0 3
rlabel polysilicon 226 -1153 226 -1153 0 1
rlabel polysilicon 229 -1153 229 -1153 0 2
rlabel polysilicon 226 -1159 226 -1159 0 3
rlabel polysilicon 229 -1159 229 -1159 0 4
rlabel polysilicon 236 -1153 236 -1153 0 2
rlabel polysilicon 233 -1159 233 -1159 0 3
rlabel polysilicon 236 -1159 236 -1159 0 4
rlabel polysilicon 240 -1153 240 -1153 0 1
rlabel polysilicon 243 -1153 243 -1153 0 2
rlabel polysilicon 240 -1159 240 -1159 0 3
rlabel polysilicon 243 -1159 243 -1159 0 4
rlabel polysilicon 247 -1153 247 -1153 0 1
rlabel polysilicon 247 -1159 247 -1159 0 3
rlabel polysilicon 254 -1153 254 -1153 0 1
rlabel polysilicon 254 -1159 254 -1159 0 3
rlabel polysilicon 261 -1153 261 -1153 0 1
rlabel polysilicon 264 -1153 264 -1153 0 2
rlabel polysilicon 264 -1159 264 -1159 0 4
rlabel polysilicon 268 -1153 268 -1153 0 1
rlabel polysilicon 268 -1159 268 -1159 0 3
rlabel polysilicon 275 -1153 275 -1153 0 1
rlabel polysilicon 275 -1159 275 -1159 0 3
rlabel polysilicon 282 -1153 282 -1153 0 1
rlabel polysilicon 282 -1159 282 -1159 0 3
rlabel polysilicon 289 -1153 289 -1153 0 1
rlabel polysilicon 289 -1159 289 -1159 0 3
rlabel polysilicon 296 -1153 296 -1153 0 1
rlabel polysilicon 296 -1159 296 -1159 0 3
rlabel polysilicon 306 -1159 306 -1159 0 4
rlabel polysilicon 310 -1153 310 -1153 0 1
rlabel polysilicon 310 -1159 310 -1159 0 3
rlabel polysilicon 317 -1153 317 -1153 0 1
rlabel polysilicon 317 -1159 317 -1159 0 3
rlabel polysilicon 324 -1153 324 -1153 0 1
rlabel polysilicon 324 -1159 324 -1159 0 3
rlabel polysilicon 334 -1153 334 -1153 0 2
rlabel polysilicon 331 -1159 331 -1159 0 3
rlabel polysilicon 338 -1153 338 -1153 0 1
rlabel polysilicon 338 -1159 338 -1159 0 3
rlabel polysilicon 345 -1153 345 -1153 0 1
rlabel polysilicon 345 -1159 345 -1159 0 3
rlabel polysilicon 355 -1159 355 -1159 0 4
rlabel polysilicon 359 -1153 359 -1153 0 1
rlabel polysilicon 359 -1159 359 -1159 0 3
rlabel polysilicon 366 -1153 366 -1153 0 1
rlabel polysilicon 369 -1153 369 -1153 0 2
rlabel polysilicon 366 -1159 366 -1159 0 3
rlabel polysilicon 373 -1153 373 -1153 0 1
rlabel polysilicon 373 -1159 373 -1159 0 3
rlabel polysilicon 380 -1153 380 -1153 0 1
rlabel polysilicon 380 -1159 380 -1159 0 3
rlabel polysilicon 387 -1153 387 -1153 0 1
rlabel polysilicon 387 -1159 387 -1159 0 3
rlabel polysilicon 394 -1153 394 -1153 0 1
rlabel polysilicon 394 -1159 394 -1159 0 3
rlabel polysilicon 401 -1153 401 -1153 0 1
rlabel polysilicon 401 -1159 401 -1159 0 3
rlabel polysilicon 408 -1153 408 -1153 0 1
rlabel polysilicon 408 -1159 408 -1159 0 3
rlabel polysilicon 415 -1153 415 -1153 0 1
rlabel polysilicon 415 -1159 415 -1159 0 3
rlabel polysilicon 422 -1153 422 -1153 0 1
rlabel polysilicon 422 -1159 422 -1159 0 3
rlabel polysilicon 429 -1153 429 -1153 0 1
rlabel polysilicon 429 -1159 429 -1159 0 3
rlabel polysilicon 436 -1153 436 -1153 0 1
rlabel polysilicon 439 -1153 439 -1153 0 2
rlabel polysilicon 436 -1159 436 -1159 0 3
rlabel polysilicon 439 -1159 439 -1159 0 4
rlabel polysilicon 443 -1153 443 -1153 0 1
rlabel polysilicon 446 -1153 446 -1153 0 2
rlabel polysilicon 443 -1159 443 -1159 0 3
rlabel polysilicon 446 -1159 446 -1159 0 4
rlabel polysilicon 450 -1153 450 -1153 0 1
rlabel polysilicon 450 -1159 450 -1159 0 3
rlabel polysilicon 457 -1153 457 -1153 0 1
rlabel polysilicon 457 -1159 457 -1159 0 3
rlabel polysilicon 467 -1153 467 -1153 0 2
rlabel polysilicon 464 -1159 464 -1159 0 3
rlabel polysilicon 467 -1159 467 -1159 0 4
rlabel polysilicon 474 -1153 474 -1153 0 2
rlabel polysilicon 471 -1159 471 -1159 0 3
rlabel polysilicon 474 -1159 474 -1159 0 4
rlabel polysilicon 478 -1153 478 -1153 0 1
rlabel polysilicon 478 -1159 478 -1159 0 3
rlabel polysilicon 485 -1153 485 -1153 0 1
rlabel polysilicon 485 -1159 485 -1159 0 3
rlabel polysilicon 492 -1153 492 -1153 0 1
rlabel polysilicon 495 -1153 495 -1153 0 2
rlabel polysilicon 495 -1159 495 -1159 0 4
rlabel polysilicon 499 -1153 499 -1153 0 1
rlabel polysilicon 499 -1159 499 -1159 0 3
rlabel polysilicon 506 -1153 506 -1153 0 1
rlabel polysilicon 509 -1153 509 -1153 0 2
rlabel polysilicon 509 -1159 509 -1159 0 4
rlabel polysilicon 513 -1153 513 -1153 0 1
rlabel polysilicon 513 -1159 513 -1159 0 3
rlabel polysilicon 520 -1153 520 -1153 0 1
rlabel polysilicon 520 -1159 520 -1159 0 3
rlabel polysilicon 530 -1153 530 -1153 0 2
rlabel polysilicon 530 -1159 530 -1159 0 4
rlabel polysilicon 534 -1153 534 -1153 0 1
rlabel polysilicon 534 -1159 534 -1159 0 3
rlabel polysilicon 541 -1153 541 -1153 0 1
rlabel polysilicon 541 -1159 541 -1159 0 3
rlabel polysilicon 548 -1153 548 -1153 0 1
rlabel polysilicon 548 -1159 548 -1159 0 3
rlabel polysilicon 555 -1153 555 -1153 0 1
rlabel polysilicon 555 -1159 555 -1159 0 3
rlabel polysilicon 562 -1153 562 -1153 0 1
rlabel polysilicon 562 -1159 562 -1159 0 3
rlabel polysilicon 569 -1153 569 -1153 0 1
rlabel polysilicon 569 -1159 569 -1159 0 3
rlabel polysilicon 576 -1153 576 -1153 0 1
rlabel polysilicon 576 -1159 576 -1159 0 3
rlabel polysilicon 583 -1153 583 -1153 0 1
rlabel polysilicon 586 -1153 586 -1153 0 2
rlabel polysilicon 583 -1159 583 -1159 0 3
rlabel polysilicon 586 -1159 586 -1159 0 4
rlabel polysilicon 590 -1153 590 -1153 0 1
rlabel polysilicon 593 -1153 593 -1153 0 2
rlabel polysilicon 590 -1159 590 -1159 0 3
rlabel polysilicon 593 -1159 593 -1159 0 4
rlabel polysilicon 597 -1153 597 -1153 0 1
rlabel polysilicon 600 -1153 600 -1153 0 2
rlabel polysilicon 597 -1159 597 -1159 0 3
rlabel polysilicon 600 -1159 600 -1159 0 4
rlabel polysilicon 604 -1153 604 -1153 0 1
rlabel polysilicon 607 -1153 607 -1153 0 2
rlabel polysilicon 604 -1159 604 -1159 0 3
rlabel polysilicon 611 -1153 611 -1153 0 1
rlabel polysilicon 611 -1159 611 -1159 0 3
rlabel polysilicon 621 -1153 621 -1153 0 2
rlabel polysilicon 618 -1159 618 -1159 0 3
rlabel polysilicon 621 -1159 621 -1159 0 4
rlabel polysilicon 628 -1153 628 -1153 0 2
rlabel polysilicon 625 -1159 625 -1159 0 3
rlabel polysilicon 628 -1159 628 -1159 0 4
rlabel polysilicon 632 -1153 632 -1153 0 1
rlabel polysilicon 632 -1159 632 -1159 0 3
rlabel polysilicon 642 -1153 642 -1153 0 2
rlabel polysilicon 639 -1159 639 -1159 0 3
rlabel polysilicon 642 -1159 642 -1159 0 4
rlabel polysilicon 646 -1153 646 -1153 0 1
rlabel polysilicon 646 -1159 646 -1159 0 3
rlabel polysilicon 653 -1153 653 -1153 0 1
rlabel polysilicon 653 -1159 653 -1159 0 3
rlabel polysilicon 660 -1153 660 -1153 0 1
rlabel polysilicon 660 -1159 660 -1159 0 3
rlabel polysilicon 663 -1159 663 -1159 0 4
rlabel polysilicon 667 -1153 667 -1153 0 1
rlabel polysilicon 667 -1159 667 -1159 0 3
rlabel polysilicon 674 -1153 674 -1153 0 1
rlabel polysilicon 677 -1153 677 -1153 0 2
rlabel polysilicon 677 -1159 677 -1159 0 4
rlabel polysilicon 681 -1153 681 -1153 0 1
rlabel polysilicon 681 -1159 681 -1159 0 3
rlabel polysilicon 688 -1153 688 -1153 0 1
rlabel polysilicon 691 -1159 691 -1159 0 4
rlabel polysilicon 695 -1153 695 -1153 0 1
rlabel polysilicon 695 -1159 695 -1159 0 3
rlabel polysilicon 702 -1153 702 -1153 0 1
rlabel polysilicon 702 -1159 702 -1159 0 3
rlabel polysilicon 709 -1153 709 -1153 0 1
rlabel polysilicon 709 -1159 709 -1159 0 3
rlabel polysilicon 716 -1153 716 -1153 0 1
rlabel polysilicon 716 -1159 716 -1159 0 3
rlabel polysilicon 723 -1153 723 -1153 0 1
rlabel polysilicon 726 -1153 726 -1153 0 2
rlabel polysilicon 723 -1159 723 -1159 0 3
rlabel polysilicon 730 -1153 730 -1153 0 1
rlabel polysilicon 733 -1159 733 -1159 0 4
rlabel polysilicon 737 -1153 737 -1153 0 1
rlabel polysilicon 737 -1159 737 -1159 0 3
rlabel polysilicon 744 -1153 744 -1153 0 1
rlabel polysilicon 744 -1159 744 -1159 0 3
rlabel polysilicon 751 -1153 751 -1153 0 1
rlabel polysilicon 751 -1159 751 -1159 0 3
rlabel polysilicon 758 -1153 758 -1153 0 1
rlabel polysilicon 758 -1159 758 -1159 0 3
rlabel polysilicon 765 -1153 765 -1153 0 1
rlabel polysilicon 765 -1159 765 -1159 0 3
rlabel polysilicon 772 -1153 772 -1153 0 1
rlabel polysilicon 772 -1159 772 -1159 0 3
rlabel polysilicon 779 -1153 779 -1153 0 1
rlabel polysilicon 779 -1159 779 -1159 0 3
rlabel polysilicon 786 -1153 786 -1153 0 1
rlabel polysilicon 786 -1159 786 -1159 0 3
rlabel polysilicon 793 -1153 793 -1153 0 1
rlabel polysilicon 793 -1159 793 -1159 0 3
rlabel polysilicon 800 -1153 800 -1153 0 1
rlabel polysilicon 800 -1159 800 -1159 0 3
rlabel polysilicon 807 -1153 807 -1153 0 1
rlabel polysilicon 807 -1159 807 -1159 0 3
rlabel polysilicon 814 -1153 814 -1153 0 1
rlabel polysilicon 814 -1159 814 -1159 0 3
rlabel polysilicon 821 -1153 821 -1153 0 1
rlabel polysilicon 821 -1159 821 -1159 0 3
rlabel polysilicon 828 -1153 828 -1153 0 1
rlabel polysilicon 828 -1159 828 -1159 0 3
rlabel polysilicon 835 -1153 835 -1153 0 1
rlabel polysilicon 835 -1159 835 -1159 0 3
rlabel polysilicon 842 -1153 842 -1153 0 1
rlabel polysilicon 842 -1159 842 -1159 0 3
rlabel polysilicon 849 -1153 849 -1153 0 1
rlabel polysilicon 849 -1159 849 -1159 0 3
rlabel polysilicon 856 -1153 856 -1153 0 1
rlabel polysilicon 856 -1159 856 -1159 0 3
rlabel polysilicon 863 -1153 863 -1153 0 1
rlabel polysilicon 863 -1159 863 -1159 0 3
rlabel polysilicon 870 -1153 870 -1153 0 1
rlabel polysilicon 870 -1159 870 -1159 0 3
rlabel polysilicon 877 -1153 877 -1153 0 1
rlabel polysilicon 877 -1159 877 -1159 0 3
rlabel polysilicon 884 -1153 884 -1153 0 1
rlabel polysilicon 884 -1159 884 -1159 0 3
rlabel polysilicon 891 -1153 891 -1153 0 1
rlabel polysilicon 891 -1159 891 -1159 0 3
rlabel polysilicon 898 -1153 898 -1153 0 1
rlabel polysilicon 898 -1159 898 -1159 0 3
rlabel polysilicon 905 -1153 905 -1153 0 1
rlabel polysilicon 905 -1159 905 -1159 0 3
rlabel polysilicon 912 -1153 912 -1153 0 1
rlabel polysilicon 912 -1159 912 -1159 0 3
rlabel polysilicon 919 -1153 919 -1153 0 1
rlabel polysilicon 919 -1159 919 -1159 0 3
rlabel polysilicon 926 -1153 926 -1153 0 1
rlabel polysilicon 926 -1159 926 -1159 0 3
rlabel polysilicon 933 -1153 933 -1153 0 1
rlabel polysilicon 933 -1159 933 -1159 0 3
rlabel polysilicon 940 -1153 940 -1153 0 1
rlabel polysilicon 940 -1159 940 -1159 0 3
rlabel polysilicon 947 -1153 947 -1153 0 1
rlabel polysilicon 947 -1159 947 -1159 0 3
rlabel polysilicon 954 -1153 954 -1153 0 1
rlabel polysilicon 954 -1159 954 -1159 0 3
rlabel polysilicon 961 -1153 961 -1153 0 1
rlabel polysilicon 961 -1159 961 -1159 0 3
rlabel polysilicon 968 -1153 968 -1153 0 1
rlabel polysilicon 968 -1159 968 -1159 0 3
rlabel polysilicon 975 -1153 975 -1153 0 1
rlabel polysilicon 975 -1159 975 -1159 0 3
rlabel polysilicon 982 -1153 982 -1153 0 1
rlabel polysilicon 982 -1159 982 -1159 0 3
rlabel polysilicon 989 -1153 989 -1153 0 1
rlabel polysilicon 989 -1159 989 -1159 0 3
rlabel polysilicon 996 -1153 996 -1153 0 1
rlabel polysilicon 996 -1159 996 -1159 0 3
rlabel polysilicon 1003 -1153 1003 -1153 0 1
rlabel polysilicon 1003 -1159 1003 -1159 0 3
rlabel polysilicon 1010 -1153 1010 -1153 0 1
rlabel polysilicon 1010 -1159 1010 -1159 0 3
rlabel polysilicon 1017 -1153 1017 -1153 0 1
rlabel polysilicon 1017 -1159 1017 -1159 0 3
rlabel polysilicon 1024 -1153 1024 -1153 0 1
rlabel polysilicon 1024 -1159 1024 -1159 0 3
rlabel polysilicon 1031 -1153 1031 -1153 0 1
rlabel polysilicon 1031 -1159 1031 -1159 0 3
rlabel polysilicon 1038 -1153 1038 -1153 0 1
rlabel polysilicon 1038 -1159 1038 -1159 0 3
rlabel polysilicon 1045 -1153 1045 -1153 0 1
rlabel polysilicon 1045 -1159 1045 -1159 0 3
rlabel polysilicon 1052 -1153 1052 -1153 0 1
rlabel polysilicon 1052 -1159 1052 -1159 0 3
rlabel polysilicon 1059 -1153 1059 -1153 0 1
rlabel polysilicon 1059 -1159 1059 -1159 0 3
rlabel polysilicon 1066 -1153 1066 -1153 0 1
rlabel polysilicon 1066 -1159 1066 -1159 0 3
rlabel polysilicon 1073 -1153 1073 -1153 0 1
rlabel polysilicon 1073 -1159 1073 -1159 0 3
rlabel polysilicon 1080 -1153 1080 -1153 0 1
rlabel polysilicon 1080 -1159 1080 -1159 0 3
rlabel polysilicon 1087 -1153 1087 -1153 0 1
rlabel polysilicon 1087 -1159 1087 -1159 0 3
rlabel polysilicon 1090 -1159 1090 -1159 0 4
rlabel polysilicon 1094 -1153 1094 -1153 0 1
rlabel polysilicon 1097 -1153 1097 -1153 0 2
rlabel polysilicon 1094 -1159 1094 -1159 0 3
rlabel polysilicon 1101 -1153 1101 -1153 0 1
rlabel polysilicon 1101 -1159 1101 -1159 0 3
rlabel polysilicon 2 -1256 2 -1256 0 1
rlabel polysilicon 2 -1262 2 -1262 0 3
rlabel polysilicon 9 -1256 9 -1256 0 1
rlabel polysilicon 9 -1262 9 -1262 0 3
rlabel polysilicon 16 -1256 16 -1256 0 1
rlabel polysilicon 23 -1256 23 -1256 0 1
rlabel polysilicon 26 -1256 26 -1256 0 2
rlabel polysilicon 23 -1262 23 -1262 0 3
rlabel polysilicon 30 -1256 30 -1256 0 1
rlabel polysilicon 30 -1262 30 -1262 0 3
rlabel polysilicon 37 -1256 37 -1256 0 1
rlabel polysilicon 37 -1262 37 -1262 0 3
rlabel polysilicon 44 -1256 44 -1256 0 1
rlabel polysilicon 44 -1262 44 -1262 0 3
rlabel polysilicon 51 -1256 51 -1256 0 1
rlabel polysilicon 51 -1262 51 -1262 0 3
rlabel polysilicon 54 -1262 54 -1262 0 4
rlabel polysilicon 58 -1256 58 -1256 0 1
rlabel polysilicon 58 -1262 58 -1262 0 3
rlabel polysilicon 65 -1256 65 -1256 0 1
rlabel polysilicon 65 -1262 65 -1262 0 3
rlabel polysilicon 72 -1256 72 -1256 0 1
rlabel polysilicon 72 -1262 72 -1262 0 3
rlabel polysilicon 79 -1256 79 -1256 0 1
rlabel polysilicon 82 -1256 82 -1256 0 2
rlabel polysilicon 86 -1256 86 -1256 0 1
rlabel polysilicon 86 -1262 86 -1262 0 3
rlabel polysilicon 93 -1256 93 -1256 0 1
rlabel polysilicon 93 -1262 93 -1262 0 3
rlabel polysilicon 100 -1256 100 -1256 0 1
rlabel polysilicon 100 -1262 100 -1262 0 3
rlabel polysilicon 107 -1256 107 -1256 0 1
rlabel polysilicon 107 -1262 107 -1262 0 3
rlabel polysilicon 114 -1256 114 -1256 0 1
rlabel polysilicon 117 -1256 117 -1256 0 2
rlabel polysilicon 114 -1262 114 -1262 0 3
rlabel polysilicon 117 -1262 117 -1262 0 4
rlabel polysilicon 121 -1256 121 -1256 0 1
rlabel polysilicon 121 -1262 121 -1262 0 3
rlabel polysilicon 128 -1256 128 -1256 0 1
rlabel polysilicon 128 -1262 128 -1262 0 3
rlabel polysilicon 135 -1256 135 -1256 0 1
rlabel polysilicon 135 -1262 135 -1262 0 3
rlabel polysilicon 142 -1256 142 -1256 0 1
rlabel polysilicon 142 -1262 142 -1262 0 3
rlabel polysilicon 149 -1256 149 -1256 0 1
rlabel polysilicon 149 -1262 149 -1262 0 3
rlabel polysilicon 156 -1256 156 -1256 0 1
rlabel polysilicon 156 -1262 156 -1262 0 3
rlabel polysilicon 163 -1256 163 -1256 0 1
rlabel polysilicon 166 -1256 166 -1256 0 2
rlabel polysilicon 163 -1262 163 -1262 0 3
rlabel polysilicon 166 -1262 166 -1262 0 4
rlabel polysilicon 170 -1256 170 -1256 0 1
rlabel polysilicon 170 -1262 170 -1262 0 3
rlabel polysilicon 177 -1256 177 -1256 0 1
rlabel polysilicon 177 -1262 177 -1262 0 3
rlabel polysilicon 184 -1256 184 -1256 0 1
rlabel polysilicon 187 -1256 187 -1256 0 2
rlabel polysilicon 184 -1262 184 -1262 0 3
rlabel polysilicon 187 -1262 187 -1262 0 4
rlabel polysilicon 191 -1256 191 -1256 0 1
rlabel polysilicon 194 -1256 194 -1256 0 2
rlabel polysilicon 194 -1262 194 -1262 0 4
rlabel polysilicon 198 -1256 198 -1256 0 1
rlabel polysilicon 201 -1262 201 -1262 0 4
rlabel polysilicon 205 -1256 205 -1256 0 1
rlabel polysilicon 205 -1262 205 -1262 0 3
rlabel polysilicon 215 -1256 215 -1256 0 2
rlabel polysilicon 212 -1262 212 -1262 0 3
rlabel polysilicon 215 -1262 215 -1262 0 4
rlabel polysilicon 219 -1256 219 -1256 0 1
rlabel polysilicon 219 -1262 219 -1262 0 3
rlabel polysilicon 222 -1262 222 -1262 0 4
rlabel polysilicon 226 -1256 226 -1256 0 1
rlabel polysilicon 226 -1262 226 -1262 0 3
rlabel polysilicon 233 -1256 233 -1256 0 1
rlabel polysilicon 233 -1262 233 -1262 0 3
rlabel polysilicon 240 -1256 240 -1256 0 1
rlabel polysilicon 240 -1262 240 -1262 0 3
rlabel polysilicon 247 -1256 247 -1256 0 1
rlabel polysilicon 247 -1262 247 -1262 0 3
rlabel polysilicon 254 -1256 254 -1256 0 1
rlabel polysilicon 254 -1262 254 -1262 0 3
rlabel polysilicon 261 -1256 261 -1256 0 1
rlabel polysilicon 261 -1262 261 -1262 0 3
rlabel polysilicon 268 -1256 268 -1256 0 1
rlabel polysilicon 268 -1262 268 -1262 0 3
rlabel polysilicon 275 -1256 275 -1256 0 1
rlabel polysilicon 275 -1262 275 -1262 0 3
rlabel polysilicon 282 -1256 282 -1256 0 1
rlabel polysilicon 282 -1262 282 -1262 0 3
rlabel polysilicon 289 -1256 289 -1256 0 1
rlabel polysilicon 292 -1256 292 -1256 0 2
rlabel polysilicon 289 -1262 289 -1262 0 3
rlabel polysilicon 292 -1262 292 -1262 0 4
rlabel polysilicon 296 -1256 296 -1256 0 1
rlabel polysilicon 296 -1262 296 -1262 0 3
rlabel polysilicon 303 -1256 303 -1256 0 1
rlabel polysilicon 303 -1262 303 -1262 0 3
rlabel polysilicon 310 -1256 310 -1256 0 1
rlabel polysilicon 310 -1262 310 -1262 0 3
rlabel polysilicon 317 -1256 317 -1256 0 1
rlabel polysilicon 317 -1262 317 -1262 0 3
rlabel polysilicon 324 -1256 324 -1256 0 1
rlabel polysilicon 324 -1262 324 -1262 0 3
rlabel polysilicon 331 -1256 331 -1256 0 1
rlabel polysilicon 331 -1262 331 -1262 0 3
rlabel polysilicon 338 -1256 338 -1256 0 1
rlabel polysilicon 338 -1262 338 -1262 0 3
rlabel polysilicon 345 -1256 345 -1256 0 1
rlabel polysilicon 345 -1262 345 -1262 0 3
rlabel polysilicon 352 -1256 352 -1256 0 1
rlabel polysilicon 352 -1262 352 -1262 0 3
rlabel polysilicon 359 -1256 359 -1256 0 1
rlabel polysilicon 359 -1262 359 -1262 0 3
rlabel polysilicon 366 -1256 366 -1256 0 1
rlabel polysilicon 366 -1262 366 -1262 0 3
rlabel polysilicon 373 -1256 373 -1256 0 1
rlabel polysilicon 373 -1262 373 -1262 0 3
rlabel polysilicon 380 -1256 380 -1256 0 1
rlabel polysilicon 380 -1262 380 -1262 0 3
rlabel polysilicon 387 -1256 387 -1256 0 1
rlabel polysilicon 387 -1262 387 -1262 0 3
rlabel polysilicon 394 -1256 394 -1256 0 1
rlabel polysilicon 394 -1262 394 -1262 0 3
rlabel polysilicon 401 -1256 401 -1256 0 1
rlabel polysilicon 401 -1262 401 -1262 0 3
rlabel polysilicon 408 -1256 408 -1256 0 1
rlabel polysilicon 408 -1262 408 -1262 0 3
rlabel polysilicon 415 -1256 415 -1256 0 1
rlabel polysilicon 415 -1262 415 -1262 0 3
rlabel polysilicon 422 -1256 422 -1256 0 1
rlabel polysilicon 422 -1262 422 -1262 0 3
rlabel polysilicon 425 -1262 425 -1262 0 4
rlabel polysilicon 429 -1256 429 -1256 0 1
rlabel polysilicon 432 -1262 432 -1262 0 4
rlabel polysilicon 436 -1256 436 -1256 0 1
rlabel polysilicon 436 -1262 436 -1262 0 3
rlabel polysilicon 443 -1256 443 -1256 0 1
rlabel polysilicon 443 -1262 443 -1262 0 3
rlabel polysilicon 450 -1256 450 -1256 0 1
rlabel polysilicon 450 -1262 450 -1262 0 3
rlabel polysilicon 457 -1256 457 -1256 0 1
rlabel polysilicon 460 -1256 460 -1256 0 2
rlabel polysilicon 457 -1262 457 -1262 0 3
rlabel polysilicon 464 -1256 464 -1256 0 1
rlabel polysilicon 464 -1262 464 -1262 0 3
rlabel polysilicon 471 -1256 471 -1256 0 1
rlabel polysilicon 474 -1256 474 -1256 0 2
rlabel polysilicon 471 -1262 471 -1262 0 3
rlabel polysilicon 478 -1256 478 -1256 0 1
rlabel polysilicon 478 -1262 478 -1262 0 3
rlabel polysilicon 485 -1256 485 -1256 0 1
rlabel polysilicon 485 -1262 485 -1262 0 3
rlabel polysilicon 492 -1256 492 -1256 0 1
rlabel polysilicon 495 -1256 495 -1256 0 2
rlabel polysilicon 492 -1262 492 -1262 0 3
rlabel polysilicon 495 -1262 495 -1262 0 4
rlabel polysilicon 499 -1256 499 -1256 0 1
rlabel polysilicon 502 -1256 502 -1256 0 2
rlabel polysilicon 499 -1262 499 -1262 0 3
rlabel polysilicon 502 -1262 502 -1262 0 4
rlabel polysilicon 506 -1256 506 -1256 0 1
rlabel polysilicon 506 -1262 506 -1262 0 3
rlabel polysilicon 513 -1256 513 -1256 0 1
rlabel polysilicon 516 -1256 516 -1256 0 2
rlabel polysilicon 513 -1262 513 -1262 0 3
rlabel polysilicon 516 -1262 516 -1262 0 4
rlabel polysilicon 523 -1256 523 -1256 0 2
rlabel polysilicon 520 -1262 520 -1262 0 3
rlabel polysilicon 527 -1256 527 -1256 0 1
rlabel polysilicon 527 -1262 527 -1262 0 3
rlabel polysilicon 537 -1262 537 -1262 0 4
rlabel polysilicon 541 -1256 541 -1256 0 1
rlabel polysilicon 544 -1256 544 -1256 0 2
rlabel polysilicon 541 -1262 541 -1262 0 3
rlabel polysilicon 544 -1262 544 -1262 0 4
rlabel polysilicon 548 -1256 548 -1256 0 1
rlabel polysilicon 551 -1256 551 -1256 0 2
rlabel polysilicon 548 -1262 548 -1262 0 3
rlabel polysilicon 555 -1256 555 -1256 0 1
rlabel polysilicon 555 -1262 555 -1262 0 3
rlabel polysilicon 562 -1256 562 -1256 0 1
rlabel polysilicon 565 -1256 565 -1256 0 2
rlabel polysilicon 562 -1262 562 -1262 0 3
rlabel polysilicon 565 -1262 565 -1262 0 4
rlabel polysilicon 569 -1256 569 -1256 0 1
rlabel polysilicon 569 -1262 569 -1262 0 3
rlabel polysilicon 576 -1256 576 -1256 0 1
rlabel polysilicon 576 -1262 576 -1262 0 3
rlabel polysilicon 586 -1256 586 -1256 0 2
rlabel polysilicon 583 -1262 583 -1262 0 3
rlabel polysilicon 586 -1262 586 -1262 0 4
rlabel polysilicon 590 -1256 590 -1256 0 1
rlabel polysilicon 597 -1256 597 -1256 0 1
rlabel polysilicon 597 -1262 597 -1262 0 3
rlabel polysilicon 604 -1256 604 -1256 0 1
rlabel polysilicon 607 -1256 607 -1256 0 2
rlabel polysilicon 604 -1262 604 -1262 0 3
rlabel polysilicon 607 -1262 607 -1262 0 4
rlabel polysilicon 611 -1256 611 -1256 0 1
rlabel polysilicon 611 -1262 611 -1262 0 3
rlabel polysilicon 618 -1256 618 -1256 0 1
rlabel polysilicon 618 -1262 618 -1262 0 3
rlabel polysilicon 625 -1256 625 -1256 0 1
rlabel polysilicon 625 -1262 625 -1262 0 3
rlabel polysilicon 632 -1256 632 -1256 0 1
rlabel polysilicon 632 -1262 632 -1262 0 3
rlabel polysilicon 639 -1256 639 -1256 0 1
rlabel polysilicon 639 -1262 639 -1262 0 3
rlabel polysilicon 646 -1256 646 -1256 0 1
rlabel polysilicon 646 -1262 646 -1262 0 3
rlabel polysilicon 656 -1256 656 -1256 0 2
rlabel polysilicon 653 -1262 653 -1262 0 3
rlabel polysilicon 656 -1262 656 -1262 0 4
rlabel polysilicon 660 -1256 660 -1256 0 1
rlabel polysilicon 660 -1262 660 -1262 0 3
rlabel polysilicon 667 -1256 667 -1256 0 1
rlabel polysilicon 667 -1262 667 -1262 0 3
rlabel polysilicon 674 -1256 674 -1256 0 1
rlabel polysilicon 674 -1262 674 -1262 0 3
rlabel polysilicon 681 -1256 681 -1256 0 1
rlabel polysilicon 684 -1256 684 -1256 0 2
rlabel polysilicon 688 -1256 688 -1256 0 1
rlabel polysilicon 688 -1262 688 -1262 0 3
rlabel polysilicon 695 -1256 695 -1256 0 1
rlabel polysilicon 695 -1262 695 -1262 0 3
rlabel polysilicon 702 -1256 702 -1256 0 1
rlabel polysilicon 702 -1262 702 -1262 0 3
rlabel polysilicon 709 -1256 709 -1256 0 1
rlabel polysilicon 709 -1262 709 -1262 0 3
rlabel polysilicon 716 -1256 716 -1256 0 1
rlabel polysilicon 719 -1256 719 -1256 0 2
rlabel polysilicon 716 -1262 716 -1262 0 3
rlabel polysilicon 723 -1256 723 -1256 0 1
rlabel polysilicon 723 -1262 723 -1262 0 3
rlabel polysilicon 730 -1256 730 -1256 0 1
rlabel polysilicon 730 -1262 730 -1262 0 3
rlabel polysilicon 737 -1256 737 -1256 0 1
rlabel polysilicon 737 -1262 737 -1262 0 3
rlabel polysilicon 744 -1256 744 -1256 0 1
rlabel polysilicon 744 -1262 744 -1262 0 3
rlabel polysilicon 751 -1256 751 -1256 0 1
rlabel polysilicon 751 -1262 751 -1262 0 3
rlabel polysilicon 758 -1256 758 -1256 0 1
rlabel polysilicon 758 -1262 758 -1262 0 3
rlabel polysilicon 765 -1256 765 -1256 0 1
rlabel polysilicon 765 -1262 765 -1262 0 3
rlabel polysilicon 772 -1256 772 -1256 0 1
rlabel polysilicon 772 -1262 772 -1262 0 3
rlabel polysilicon 779 -1256 779 -1256 0 1
rlabel polysilicon 782 -1256 782 -1256 0 2
rlabel polysilicon 786 -1256 786 -1256 0 1
rlabel polysilicon 786 -1262 786 -1262 0 3
rlabel polysilicon 793 -1256 793 -1256 0 1
rlabel polysilicon 793 -1262 793 -1262 0 3
rlabel polysilicon 800 -1256 800 -1256 0 1
rlabel polysilicon 800 -1262 800 -1262 0 3
rlabel polysilicon 807 -1256 807 -1256 0 1
rlabel polysilicon 807 -1262 807 -1262 0 3
rlabel polysilicon 814 -1256 814 -1256 0 1
rlabel polysilicon 817 -1262 817 -1262 0 4
rlabel polysilicon 821 -1256 821 -1256 0 1
rlabel polysilicon 821 -1262 821 -1262 0 3
rlabel polysilicon 828 -1256 828 -1256 0 1
rlabel polysilicon 828 -1262 828 -1262 0 3
rlabel polysilicon 835 -1256 835 -1256 0 1
rlabel polysilicon 835 -1262 835 -1262 0 3
rlabel polysilicon 842 -1256 842 -1256 0 1
rlabel polysilicon 842 -1262 842 -1262 0 3
rlabel polysilicon 849 -1256 849 -1256 0 1
rlabel polysilicon 849 -1262 849 -1262 0 3
rlabel polysilicon 856 -1256 856 -1256 0 1
rlabel polysilicon 856 -1262 856 -1262 0 3
rlabel polysilicon 863 -1256 863 -1256 0 1
rlabel polysilicon 863 -1262 863 -1262 0 3
rlabel polysilicon 870 -1256 870 -1256 0 1
rlabel polysilicon 870 -1262 870 -1262 0 3
rlabel polysilicon 877 -1256 877 -1256 0 1
rlabel polysilicon 877 -1262 877 -1262 0 3
rlabel polysilicon 884 -1256 884 -1256 0 1
rlabel polysilicon 884 -1262 884 -1262 0 3
rlabel polysilicon 891 -1256 891 -1256 0 1
rlabel polysilicon 891 -1262 891 -1262 0 3
rlabel polysilicon 898 -1256 898 -1256 0 1
rlabel polysilicon 898 -1262 898 -1262 0 3
rlabel polysilicon 905 -1256 905 -1256 0 1
rlabel polysilicon 905 -1262 905 -1262 0 3
rlabel polysilicon 912 -1256 912 -1256 0 1
rlabel polysilicon 912 -1262 912 -1262 0 3
rlabel polysilicon 919 -1256 919 -1256 0 1
rlabel polysilicon 919 -1262 919 -1262 0 3
rlabel polysilicon 926 -1256 926 -1256 0 1
rlabel polysilicon 933 -1256 933 -1256 0 1
rlabel polysilicon 933 -1262 933 -1262 0 3
rlabel polysilicon 940 -1256 940 -1256 0 1
rlabel polysilicon 940 -1262 940 -1262 0 3
rlabel polysilicon 947 -1256 947 -1256 0 1
rlabel polysilicon 947 -1262 947 -1262 0 3
rlabel polysilicon 954 -1256 954 -1256 0 1
rlabel polysilicon 954 -1262 954 -1262 0 3
rlabel polysilicon 961 -1256 961 -1256 0 1
rlabel polysilicon 961 -1262 961 -1262 0 3
rlabel polysilicon 968 -1256 968 -1256 0 1
rlabel polysilicon 968 -1262 968 -1262 0 3
rlabel polysilicon 975 -1256 975 -1256 0 1
rlabel polysilicon 975 -1262 975 -1262 0 3
rlabel polysilicon 982 -1256 982 -1256 0 1
rlabel polysilicon 982 -1262 982 -1262 0 3
rlabel polysilicon 989 -1256 989 -1256 0 1
rlabel polysilicon 989 -1262 989 -1262 0 3
rlabel polysilicon 996 -1256 996 -1256 0 1
rlabel polysilicon 996 -1262 996 -1262 0 3
rlabel polysilicon 1003 -1256 1003 -1256 0 1
rlabel polysilicon 1003 -1262 1003 -1262 0 3
rlabel polysilicon 1010 -1256 1010 -1256 0 1
rlabel polysilicon 1010 -1262 1010 -1262 0 3
rlabel polysilicon 1017 -1256 1017 -1256 0 1
rlabel polysilicon 1017 -1262 1017 -1262 0 3
rlabel polysilicon 1020 -1262 1020 -1262 0 4
rlabel polysilicon 1024 -1256 1024 -1256 0 1
rlabel polysilicon 1024 -1262 1024 -1262 0 3
rlabel polysilicon 1031 -1256 1031 -1256 0 1
rlabel polysilicon 1038 -1256 1038 -1256 0 1
rlabel polysilicon 1041 -1256 1041 -1256 0 2
rlabel polysilicon 1041 -1262 1041 -1262 0 4
rlabel polysilicon 1045 -1256 1045 -1256 0 1
rlabel polysilicon 1045 -1262 1045 -1262 0 3
rlabel polysilicon 1052 -1256 1052 -1256 0 1
rlabel polysilicon 1052 -1262 1052 -1262 0 3
rlabel polysilicon 1059 -1256 1059 -1256 0 1
rlabel polysilicon 1059 -1262 1059 -1262 0 3
rlabel polysilicon 1066 -1256 1066 -1256 0 1
rlabel polysilicon 1066 -1262 1066 -1262 0 3
rlabel polysilicon 1073 -1256 1073 -1256 0 1
rlabel polysilicon 1073 -1262 1073 -1262 0 3
rlabel polysilicon 9 -1335 9 -1335 0 1
rlabel polysilicon 9 -1341 9 -1341 0 3
rlabel polysilicon 16 -1335 16 -1335 0 1
rlabel polysilicon 16 -1341 16 -1341 0 3
rlabel polysilicon 23 -1335 23 -1335 0 1
rlabel polysilicon 23 -1341 23 -1341 0 3
rlabel polysilicon 30 -1335 30 -1335 0 1
rlabel polysilicon 30 -1341 30 -1341 0 3
rlabel polysilicon 37 -1335 37 -1335 0 1
rlabel polysilicon 37 -1341 37 -1341 0 3
rlabel polysilicon 44 -1335 44 -1335 0 1
rlabel polysilicon 44 -1341 44 -1341 0 3
rlabel polysilicon 51 -1335 51 -1335 0 1
rlabel polysilicon 51 -1341 51 -1341 0 3
rlabel polysilicon 58 -1335 58 -1335 0 1
rlabel polysilicon 58 -1341 58 -1341 0 3
rlabel polysilicon 65 -1335 65 -1335 0 1
rlabel polysilicon 65 -1341 65 -1341 0 3
rlabel polysilicon 72 -1335 72 -1335 0 1
rlabel polysilicon 72 -1341 72 -1341 0 3
rlabel polysilicon 79 -1341 79 -1341 0 3
rlabel polysilicon 86 -1335 86 -1335 0 1
rlabel polysilicon 86 -1341 86 -1341 0 3
rlabel polysilicon 93 -1335 93 -1335 0 1
rlabel polysilicon 93 -1341 93 -1341 0 3
rlabel polysilicon 100 -1335 100 -1335 0 1
rlabel polysilicon 100 -1341 100 -1341 0 3
rlabel polysilicon 107 -1335 107 -1335 0 1
rlabel polysilicon 107 -1341 107 -1341 0 3
rlabel polysilicon 117 -1335 117 -1335 0 2
rlabel polysilicon 121 -1335 121 -1335 0 1
rlabel polysilicon 121 -1341 121 -1341 0 3
rlabel polysilicon 131 -1335 131 -1335 0 2
rlabel polysilicon 128 -1341 128 -1341 0 3
rlabel polysilicon 138 -1335 138 -1335 0 2
rlabel polysilicon 138 -1341 138 -1341 0 4
rlabel polysilicon 142 -1335 142 -1335 0 1
rlabel polysilicon 142 -1341 142 -1341 0 3
rlabel polysilicon 149 -1335 149 -1335 0 1
rlabel polysilicon 149 -1341 149 -1341 0 3
rlabel polysilicon 159 -1335 159 -1335 0 2
rlabel polysilicon 159 -1341 159 -1341 0 4
rlabel polysilicon 163 -1335 163 -1335 0 1
rlabel polysilicon 163 -1341 163 -1341 0 3
rlabel polysilicon 170 -1335 170 -1335 0 1
rlabel polysilicon 173 -1335 173 -1335 0 2
rlabel polysilicon 173 -1341 173 -1341 0 4
rlabel polysilicon 177 -1341 177 -1341 0 3
rlabel polysilicon 180 -1341 180 -1341 0 4
rlabel polysilicon 184 -1335 184 -1335 0 1
rlabel polysilicon 184 -1341 184 -1341 0 3
rlabel polysilicon 191 -1335 191 -1335 0 1
rlabel polysilicon 194 -1335 194 -1335 0 2
rlabel polysilicon 194 -1341 194 -1341 0 4
rlabel polysilicon 198 -1335 198 -1335 0 1
rlabel polysilicon 198 -1341 198 -1341 0 3
rlabel polysilicon 205 -1335 205 -1335 0 1
rlabel polysilicon 205 -1341 205 -1341 0 3
rlabel polysilicon 212 -1335 212 -1335 0 1
rlabel polysilicon 212 -1341 212 -1341 0 3
rlabel polysilicon 219 -1335 219 -1335 0 1
rlabel polysilicon 222 -1335 222 -1335 0 2
rlabel polysilicon 219 -1341 219 -1341 0 3
rlabel polysilicon 222 -1341 222 -1341 0 4
rlabel polysilicon 226 -1335 226 -1335 0 1
rlabel polysilicon 226 -1341 226 -1341 0 3
rlabel polysilicon 233 -1335 233 -1335 0 1
rlabel polysilicon 233 -1341 233 -1341 0 3
rlabel polysilicon 240 -1335 240 -1335 0 1
rlabel polysilicon 240 -1341 240 -1341 0 3
rlabel polysilicon 247 -1335 247 -1335 0 1
rlabel polysilicon 247 -1341 247 -1341 0 3
rlabel polysilicon 254 -1335 254 -1335 0 1
rlabel polysilicon 254 -1341 254 -1341 0 3
rlabel polysilicon 261 -1335 261 -1335 0 1
rlabel polysilicon 261 -1341 261 -1341 0 3
rlabel polysilicon 268 -1335 268 -1335 0 1
rlabel polysilicon 268 -1341 268 -1341 0 3
rlabel polysilicon 275 -1335 275 -1335 0 1
rlabel polysilicon 275 -1341 275 -1341 0 3
rlabel polysilicon 282 -1335 282 -1335 0 1
rlabel polysilicon 282 -1341 282 -1341 0 3
rlabel polysilicon 292 -1335 292 -1335 0 2
rlabel polysilicon 292 -1341 292 -1341 0 4
rlabel polysilicon 296 -1335 296 -1335 0 1
rlabel polysilicon 296 -1341 296 -1341 0 3
rlabel polysilicon 303 -1335 303 -1335 0 1
rlabel polysilicon 303 -1341 303 -1341 0 3
rlabel polysilicon 310 -1335 310 -1335 0 1
rlabel polysilicon 310 -1341 310 -1341 0 3
rlabel polysilicon 317 -1335 317 -1335 0 1
rlabel polysilicon 320 -1335 320 -1335 0 2
rlabel polysilicon 317 -1341 317 -1341 0 3
rlabel polysilicon 327 -1335 327 -1335 0 2
rlabel polysilicon 324 -1341 324 -1341 0 3
rlabel polysilicon 327 -1341 327 -1341 0 4
rlabel polysilicon 331 -1335 331 -1335 0 1
rlabel polysilicon 331 -1341 331 -1341 0 3
rlabel polysilicon 338 -1335 338 -1335 0 1
rlabel polysilicon 338 -1341 338 -1341 0 3
rlabel polysilicon 345 -1335 345 -1335 0 1
rlabel polysilicon 345 -1341 345 -1341 0 3
rlabel polysilicon 352 -1335 352 -1335 0 1
rlabel polysilicon 355 -1335 355 -1335 0 2
rlabel polysilicon 352 -1341 352 -1341 0 3
rlabel polysilicon 355 -1341 355 -1341 0 4
rlabel polysilicon 359 -1335 359 -1335 0 1
rlabel polysilicon 359 -1341 359 -1341 0 3
rlabel polysilicon 366 -1335 366 -1335 0 1
rlabel polysilicon 369 -1335 369 -1335 0 2
rlabel polysilicon 369 -1341 369 -1341 0 4
rlabel polysilicon 373 -1335 373 -1335 0 1
rlabel polysilicon 373 -1341 373 -1341 0 3
rlabel polysilicon 380 -1335 380 -1335 0 1
rlabel polysilicon 380 -1341 380 -1341 0 3
rlabel polysilicon 387 -1335 387 -1335 0 1
rlabel polysilicon 387 -1341 387 -1341 0 3
rlabel polysilicon 394 -1335 394 -1335 0 1
rlabel polysilicon 394 -1341 394 -1341 0 3
rlabel polysilicon 401 -1335 401 -1335 0 1
rlabel polysilicon 401 -1341 401 -1341 0 3
rlabel polysilicon 408 -1335 408 -1335 0 1
rlabel polysilicon 408 -1341 408 -1341 0 3
rlabel polysilicon 415 -1335 415 -1335 0 1
rlabel polysilicon 415 -1341 415 -1341 0 3
rlabel polysilicon 422 -1335 422 -1335 0 1
rlabel polysilicon 422 -1341 422 -1341 0 3
rlabel polysilicon 432 -1335 432 -1335 0 2
rlabel polysilicon 429 -1341 429 -1341 0 3
rlabel polysilicon 432 -1341 432 -1341 0 4
rlabel polysilicon 436 -1335 436 -1335 0 1
rlabel polysilicon 436 -1341 436 -1341 0 3
rlabel polysilicon 443 -1335 443 -1335 0 1
rlabel polysilicon 443 -1341 443 -1341 0 3
rlabel polysilicon 450 -1335 450 -1335 0 1
rlabel polysilicon 450 -1341 450 -1341 0 3
rlabel polysilicon 457 -1335 457 -1335 0 1
rlabel polysilicon 460 -1335 460 -1335 0 2
rlabel polysilicon 460 -1341 460 -1341 0 4
rlabel polysilicon 464 -1335 464 -1335 0 1
rlabel polysilicon 464 -1341 464 -1341 0 3
rlabel polysilicon 474 -1335 474 -1335 0 2
rlabel polysilicon 471 -1341 471 -1341 0 3
rlabel polysilicon 478 -1335 478 -1335 0 1
rlabel polysilicon 478 -1341 478 -1341 0 3
rlabel polysilicon 485 -1335 485 -1335 0 1
rlabel polysilicon 485 -1341 485 -1341 0 3
rlabel polysilicon 492 -1335 492 -1335 0 1
rlabel polysilicon 492 -1341 492 -1341 0 3
rlabel polysilicon 495 -1341 495 -1341 0 4
rlabel polysilicon 499 -1335 499 -1335 0 1
rlabel polysilicon 499 -1341 499 -1341 0 3
rlabel polysilicon 509 -1335 509 -1335 0 2
rlabel polysilicon 506 -1341 506 -1341 0 3
rlabel polysilicon 513 -1335 513 -1335 0 1
rlabel polysilicon 513 -1341 513 -1341 0 3
rlabel polysilicon 520 -1335 520 -1335 0 1
rlabel polysilicon 520 -1341 520 -1341 0 3
rlabel polysilicon 527 -1335 527 -1335 0 1
rlabel polysilicon 527 -1341 527 -1341 0 3
rlabel polysilicon 534 -1335 534 -1335 0 1
rlabel polysilicon 537 -1335 537 -1335 0 2
rlabel polysilicon 541 -1335 541 -1335 0 1
rlabel polysilicon 541 -1341 541 -1341 0 3
rlabel polysilicon 548 -1335 548 -1335 0 1
rlabel polysilicon 548 -1341 548 -1341 0 3
rlabel polysilicon 555 -1335 555 -1335 0 1
rlabel polysilicon 555 -1341 555 -1341 0 3
rlabel polysilicon 562 -1335 562 -1335 0 1
rlabel polysilicon 562 -1341 562 -1341 0 3
rlabel polysilicon 569 -1335 569 -1335 0 1
rlabel polysilicon 569 -1341 569 -1341 0 3
rlabel polysilicon 576 -1335 576 -1335 0 1
rlabel polysilicon 579 -1335 579 -1335 0 2
rlabel polysilicon 576 -1341 576 -1341 0 3
rlabel polysilicon 579 -1341 579 -1341 0 4
rlabel polysilicon 583 -1335 583 -1335 0 1
rlabel polysilicon 583 -1341 583 -1341 0 3
rlabel polysilicon 590 -1335 590 -1335 0 1
rlabel polysilicon 590 -1341 590 -1341 0 3
rlabel polysilicon 597 -1335 597 -1335 0 1
rlabel polysilicon 597 -1341 597 -1341 0 3
rlabel polysilicon 600 -1341 600 -1341 0 4
rlabel polysilicon 604 -1335 604 -1335 0 1
rlabel polysilicon 604 -1341 604 -1341 0 3
rlabel polysilicon 611 -1335 611 -1335 0 1
rlabel polysilicon 611 -1341 611 -1341 0 3
rlabel polysilicon 621 -1335 621 -1335 0 2
rlabel polysilicon 618 -1341 618 -1341 0 3
rlabel polysilicon 625 -1335 625 -1335 0 1
rlabel polysilicon 625 -1341 625 -1341 0 3
rlabel polysilicon 632 -1335 632 -1335 0 1
rlabel polysilicon 632 -1341 632 -1341 0 3
rlabel polysilicon 639 -1335 639 -1335 0 1
rlabel polysilicon 639 -1341 639 -1341 0 3
rlabel polysilicon 646 -1335 646 -1335 0 1
rlabel polysilicon 646 -1341 646 -1341 0 3
rlabel polysilicon 649 -1341 649 -1341 0 4
rlabel polysilicon 653 -1335 653 -1335 0 1
rlabel polysilicon 653 -1341 653 -1341 0 3
rlabel polysilicon 660 -1335 660 -1335 0 1
rlabel polysilicon 660 -1341 660 -1341 0 3
rlabel polysilicon 667 -1335 667 -1335 0 1
rlabel polysilicon 667 -1341 667 -1341 0 3
rlabel polysilicon 677 -1335 677 -1335 0 2
rlabel polysilicon 674 -1341 674 -1341 0 3
rlabel polysilicon 677 -1341 677 -1341 0 4
rlabel polysilicon 681 -1335 681 -1335 0 1
rlabel polysilicon 681 -1341 681 -1341 0 3
rlabel polysilicon 688 -1335 688 -1335 0 1
rlabel polysilicon 688 -1341 688 -1341 0 3
rlabel polysilicon 695 -1335 695 -1335 0 1
rlabel polysilicon 695 -1341 695 -1341 0 3
rlabel polysilicon 702 -1341 702 -1341 0 3
rlabel polysilicon 705 -1341 705 -1341 0 4
rlabel polysilicon 709 -1335 709 -1335 0 1
rlabel polysilicon 709 -1341 709 -1341 0 3
rlabel polysilicon 716 -1335 716 -1335 0 1
rlabel polysilicon 716 -1341 716 -1341 0 3
rlabel polysilicon 723 -1335 723 -1335 0 1
rlabel polysilicon 723 -1341 723 -1341 0 3
rlabel polysilicon 730 -1335 730 -1335 0 1
rlabel polysilicon 730 -1341 730 -1341 0 3
rlabel polysilicon 737 -1341 737 -1341 0 3
rlabel polysilicon 744 -1335 744 -1335 0 1
rlabel polysilicon 744 -1341 744 -1341 0 3
rlabel polysilicon 751 -1335 751 -1335 0 1
rlabel polysilicon 751 -1341 751 -1341 0 3
rlabel polysilicon 758 -1335 758 -1335 0 1
rlabel polysilicon 761 -1335 761 -1335 0 2
rlabel polysilicon 758 -1341 758 -1341 0 3
rlabel polysilicon 765 -1335 765 -1335 0 1
rlabel polysilicon 765 -1341 765 -1341 0 3
rlabel polysilicon 772 -1335 772 -1335 0 1
rlabel polysilicon 772 -1341 772 -1341 0 3
rlabel polysilicon 779 -1335 779 -1335 0 1
rlabel polysilicon 779 -1341 779 -1341 0 3
rlabel polysilicon 786 -1335 786 -1335 0 1
rlabel polysilicon 786 -1341 786 -1341 0 3
rlabel polysilicon 793 -1335 793 -1335 0 1
rlabel polysilicon 793 -1341 793 -1341 0 3
rlabel polysilicon 800 -1335 800 -1335 0 1
rlabel polysilicon 800 -1341 800 -1341 0 3
rlabel polysilicon 807 -1335 807 -1335 0 1
rlabel polysilicon 807 -1341 807 -1341 0 3
rlabel polysilicon 814 -1335 814 -1335 0 1
rlabel polysilicon 814 -1341 814 -1341 0 3
rlabel polysilicon 821 -1335 821 -1335 0 1
rlabel polysilicon 821 -1341 821 -1341 0 3
rlabel polysilicon 828 -1335 828 -1335 0 1
rlabel polysilicon 828 -1341 828 -1341 0 3
rlabel polysilicon 835 -1335 835 -1335 0 1
rlabel polysilicon 835 -1341 835 -1341 0 3
rlabel polysilicon 842 -1335 842 -1335 0 1
rlabel polysilicon 842 -1341 842 -1341 0 3
rlabel polysilicon 849 -1335 849 -1335 0 1
rlabel polysilicon 849 -1341 849 -1341 0 3
rlabel polysilicon 856 -1335 856 -1335 0 1
rlabel polysilicon 856 -1341 856 -1341 0 3
rlabel polysilicon 863 -1335 863 -1335 0 1
rlabel polysilicon 863 -1341 863 -1341 0 3
rlabel polysilicon 870 -1335 870 -1335 0 1
rlabel polysilicon 870 -1341 870 -1341 0 3
rlabel polysilicon 877 -1335 877 -1335 0 1
rlabel polysilicon 877 -1341 877 -1341 0 3
rlabel polysilicon 884 -1335 884 -1335 0 1
rlabel polysilicon 884 -1341 884 -1341 0 3
rlabel polysilicon 891 -1335 891 -1335 0 1
rlabel polysilicon 891 -1341 891 -1341 0 3
rlabel polysilicon 898 -1335 898 -1335 0 1
rlabel polysilicon 898 -1341 898 -1341 0 3
rlabel polysilicon 905 -1335 905 -1335 0 1
rlabel polysilicon 905 -1341 905 -1341 0 3
rlabel polysilicon 912 -1335 912 -1335 0 1
rlabel polysilicon 912 -1341 912 -1341 0 3
rlabel polysilicon 919 -1335 919 -1335 0 1
rlabel polysilicon 919 -1341 919 -1341 0 3
rlabel polysilicon 926 -1341 926 -1341 0 3
rlabel polysilicon 933 -1335 933 -1335 0 1
rlabel polysilicon 933 -1341 933 -1341 0 3
rlabel polysilicon 940 -1335 940 -1335 0 1
rlabel polysilicon 940 -1341 940 -1341 0 3
rlabel polysilicon 947 -1335 947 -1335 0 1
rlabel polysilicon 947 -1341 947 -1341 0 3
rlabel polysilicon 954 -1335 954 -1335 0 1
rlabel polysilicon 954 -1341 954 -1341 0 3
rlabel polysilicon 961 -1335 961 -1335 0 1
rlabel polysilicon 961 -1341 961 -1341 0 3
rlabel polysilicon 968 -1335 968 -1335 0 1
rlabel polysilicon 968 -1341 968 -1341 0 3
rlabel polysilicon 975 -1335 975 -1335 0 1
rlabel polysilicon 975 -1341 975 -1341 0 3
rlabel polysilicon 982 -1335 982 -1335 0 1
rlabel polysilicon 982 -1341 982 -1341 0 3
rlabel polysilicon 989 -1335 989 -1335 0 1
rlabel polysilicon 989 -1341 989 -1341 0 3
rlabel polysilicon 996 -1335 996 -1335 0 1
rlabel polysilicon 996 -1341 996 -1341 0 3
rlabel polysilicon 1003 -1335 1003 -1335 0 1
rlabel polysilicon 1003 -1341 1003 -1341 0 3
rlabel polysilicon 1010 -1335 1010 -1335 0 1
rlabel polysilicon 1010 -1341 1010 -1341 0 3
rlabel polysilicon 1017 -1335 1017 -1335 0 1
rlabel polysilicon 1020 -1335 1020 -1335 0 2
rlabel polysilicon 1017 -1341 1017 -1341 0 3
rlabel polysilicon 1024 -1341 1024 -1341 0 3
rlabel polysilicon 1031 -1335 1031 -1335 0 1
rlabel polysilicon 1034 -1335 1034 -1335 0 2
rlabel polysilicon 1031 -1341 1031 -1341 0 3
rlabel polysilicon 1034 -1341 1034 -1341 0 4
rlabel polysilicon 1038 -1335 1038 -1335 0 1
rlabel polysilicon 1038 -1341 1038 -1341 0 3
rlabel polysilicon 1045 -1335 1045 -1335 0 1
rlabel polysilicon 1048 -1335 1048 -1335 0 2
rlabel polysilicon 1048 -1341 1048 -1341 0 4
rlabel polysilicon 1052 -1335 1052 -1335 0 1
rlabel polysilicon 1052 -1341 1052 -1341 0 3
rlabel polysilicon 1059 -1335 1059 -1335 0 1
rlabel polysilicon 1062 -1335 1062 -1335 0 2
rlabel polysilicon 1066 -1335 1066 -1335 0 1
rlabel polysilicon 1066 -1341 1066 -1341 0 3
rlabel polysilicon 1073 -1335 1073 -1335 0 1
rlabel polysilicon 1073 -1341 1073 -1341 0 3
rlabel polysilicon 1080 -1335 1080 -1335 0 1
rlabel polysilicon 1080 -1341 1080 -1341 0 3
rlabel polysilicon 16 -1412 16 -1412 0 1
rlabel polysilicon 16 -1418 16 -1418 0 3
rlabel polysilicon 23 -1412 23 -1412 0 1
rlabel polysilicon 23 -1418 23 -1418 0 3
rlabel polysilicon 30 -1412 30 -1412 0 1
rlabel polysilicon 30 -1418 30 -1418 0 3
rlabel polysilicon 37 -1412 37 -1412 0 1
rlabel polysilicon 37 -1418 37 -1418 0 3
rlabel polysilicon 44 -1412 44 -1412 0 1
rlabel polysilicon 44 -1418 44 -1418 0 3
rlabel polysilicon 54 -1412 54 -1412 0 2
rlabel polysilicon 51 -1418 51 -1418 0 3
rlabel polysilicon 61 -1412 61 -1412 0 2
rlabel polysilicon 65 -1412 65 -1412 0 1
rlabel polysilicon 65 -1418 65 -1418 0 3
rlabel polysilicon 72 -1412 72 -1412 0 1
rlabel polysilicon 72 -1418 72 -1418 0 3
rlabel polysilicon 79 -1412 79 -1412 0 1
rlabel polysilicon 79 -1418 79 -1418 0 3
rlabel polysilicon 86 -1412 86 -1412 0 1
rlabel polysilicon 89 -1412 89 -1412 0 2
rlabel polysilicon 86 -1418 86 -1418 0 3
rlabel polysilicon 89 -1418 89 -1418 0 4
rlabel polysilicon 93 -1412 93 -1412 0 1
rlabel polysilicon 93 -1418 93 -1418 0 3
rlabel polysilicon 100 -1412 100 -1412 0 1
rlabel polysilicon 100 -1418 100 -1418 0 3
rlabel polysilicon 107 -1412 107 -1412 0 1
rlabel polysilicon 107 -1418 107 -1418 0 3
rlabel polysilicon 114 -1412 114 -1412 0 1
rlabel polysilicon 114 -1418 114 -1418 0 3
rlabel polysilicon 121 -1412 121 -1412 0 1
rlabel polysilicon 121 -1418 121 -1418 0 3
rlabel polysilicon 128 -1412 128 -1412 0 1
rlabel polysilicon 128 -1418 128 -1418 0 3
rlabel polysilicon 135 -1412 135 -1412 0 1
rlabel polysilicon 138 -1418 138 -1418 0 4
rlabel polysilicon 145 -1412 145 -1412 0 2
rlabel polysilicon 142 -1418 142 -1418 0 3
rlabel polysilicon 149 -1412 149 -1412 0 1
rlabel polysilicon 149 -1418 149 -1418 0 3
rlabel polysilicon 156 -1412 156 -1412 0 1
rlabel polysilicon 159 -1418 159 -1418 0 4
rlabel polysilicon 163 -1412 163 -1412 0 1
rlabel polysilicon 163 -1418 163 -1418 0 3
rlabel polysilicon 166 -1418 166 -1418 0 4
rlabel polysilicon 170 -1412 170 -1412 0 1
rlabel polysilicon 170 -1418 170 -1418 0 3
rlabel polysilicon 177 -1412 177 -1412 0 1
rlabel polysilicon 177 -1418 177 -1418 0 3
rlabel polysilicon 184 -1412 184 -1412 0 1
rlabel polysilicon 184 -1418 184 -1418 0 3
rlabel polysilicon 191 -1412 191 -1412 0 1
rlabel polysilicon 191 -1418 191 -1418 0 3
rlabel polysilicon 198 -1412 198 -1412 0 1
rlabel polysilicon 198 -1418 198 -1418 0 3
rlabel polysilicon 205 -1412 205 -1412 0 1
rlabel polysilicon 208 -1412 208 -1412 0 2
rlabel polysilicon 205 -1418 205 -1418 0 3
rlabel polysilicon 212 -1412 212 -1412 0 1
rlabel polysilicon 212 -1418 212 -1418 0 3
rlabel polysilicon 222 -1412 222 -1412 0 2
rlabel polysilicon 219 -1418 219 -1418 0 3
rlabel polysilicon 222 -1418 222 -1418 0 4
rlabel polysilicon 226 -1412 226 -1412 0 1
rlabel polysilicon 226 -1418 226 -1418 0 3
rlabel polysilicon 233 -1412 233 -1412 0 1
rlabel polysilicon 233 -1418 233 -1418 0 3
rlabel polysilicon 240 -1418 240 -1418 0 3
rlabel polysilicon 243 -1418 243 -1418 0 4
rlabel polysilicon 247 -1412 247 -1412 0 1
rlabel polysilicon 247 -1418 247 -1418 0 3
rlabel polysilicon 254 -1412 254 -1412 0 1
rlabel polysilicon 254 -1418 254 -1418 0 3
rlabel polysilicon 261 -1412 261 -1412 0 1
rlabel polysilicon 261 -1418 261 -1418 0 3
rlabel polysilicon 268 -1412 268 -1412 0 1
rlabel polysilicon 268 -1418 268 -1418 0 3
rlabel polysilicon 275 -1412 275 -1412 0 1
rlabel polysilicon 275 -1418 275 -1418 0 3
rlabel polysilicon 282 -1412 282 -1412 0 1
rlabel polysilicon 282 -1418 282 -1418 0 3
rlabel polysilicon 289 -1412 289 -1412 0 1
rlabel polysilicon 289 -1418 289 -1418 0 3
rlabel polysilicon 296 -1412 296 -1412 0 1
rlabel polysilicon 296 -1418 296 -1418 0 3
rlabel polysilicon 303 -1412 303 -1412 0 1
rlabel polysilicon 303 -1418 303 -1418 0 3
rlabel polysilicon 306 -1418 306 -1418 0 4
rlabel polysilicon 310 -1412 310 -1412 0 1
rlabel polysilicon 310 -1418 310 -1418 0 3
rlabel polysilicon 317 -1412 317 -1412 0 1
rlabel polysilicon 317 -1418 317 -1418 0 3
rlabel polysilicon 324 -1412 324 -1412 0 1
rlabel polysilicon 324 -1418 324 -1418 0 3
rlabel polysilicon 331 -1412 331 -1412 0 1
rlabel polysilicon 331 -1418 331 -1418 0 3
rlabel polysilicon 338 -1412 338 -1412 0 1
rlabel polysilicon 338 -1418 338 -1418 0 3
rlabel polysilicon 345 -1412 345 -1412 0 1
rlabel polysilicon 345 -1418 345 -1418 0 3
rlabel polysilicon 352 -1412 352 -1412 0 1
rlabel polysilicon 355 -1412 355 -1412 0 2
rlabel polysilicon 355 -1418 355 -1418 0 4
rlabel polysilicon 359 -1412 359 -1412 0 1
rlabel polysilicon 362 -1418 362 -1418 0 4
rlabel polysilicon 366 -1412 366 -1412 0 1
rlabel polysilicon 366 -1418 366 -1418 0 3
rlabel polysilicon 373 -1412 373 -1412 0 1
rlabel polysilicon 373 -1418 373 -1418 0 3
rlabel polysilicon 380 -1412 380 -1412 0 1
rlabel polysilicon 380 -1418 380 -1418 0 3
rlabel polysilicon 387 -1412 387 -1412 0 1
rlabel polysilicon 390 -1418 390 -1418 0 4
rlabel polysilicon 394 -1412 394 -1412 0 1
rlabel polysilicon 394 -1418 394 -1418 0 3
rlabel polysilicon 401 -1412 401 -1412 0 1
rlabel polysilicon 401 -1418 401 -1418 0 3
rlabel polysilicon 408 -1412 408 -1412 0 1
rlabel polysilicon 411 -1412 411 -1412 0 2
rlabel polysilicon 408 -1418 408 -1418 0 3
rlabel polysilicon 411 -1418 411 -1418 0 4
rlabel polysilicon 415 -1412 415 -1412 0 1
rlabel polysilicon 415 -1418 415 -1418 0 3
rlabel polysilicon 422 -1412 422 -1412 0 1
rlabel polysilicon 422 -1418 422 -1418 0 3
rlabel polysilicon 429 -1412 429 -1412 0 1
rlabel polysilicon 429 -1418 429 -1418 0 3
rlabel polysilicon 436 -1412 436 -1412 0 1
rlabel polysilicon 436 -1418 436 -1418 0 3
rlabel polysilicon 443 -1412 443 -1412 0 1
rlabel polysilicon 443 -1418 443 -1418 0 3
rlabel polysilicon 450 -1412 450 -1412 0 1
rlabel polysilicon 450 -1418 450 -1418 0 3
rlabel polysilicon 457 -1412 457 -1412 0 1
rlabel polysilicon 457 -1418 457 -1418 0 3
rlabel polysilicon 464 -1412 464 -1412 0 1
rlabel polysilicon 464 -1418 464 -1418 0 3
rlabel polysilicon 471 -1412 471 -1412 0 1
rlabel polysilicon 471 -1418 471 -1418 0 3
rlabel polysilicon 478 -1412 478 -1412 0 1
rlabel polysilicon 478 -1418 478 -1418 0 3
rlabel polysilicon 485 -1412 485 -1412 0 1
rlabel polysilicon 485 -1418 485 -1418 0 3
rlabel polysilicon 492 -1412 492 -1412 0 1
rlabel polysilicon 492 -1418 492 -1418 0 3
rlabel polysilicon 499 -1412 499 -1412 0 1
rlabel polysilicon 499 -1418 499 -1418 0 3
rlabel polysilicon 506 -1412 506 -1412 0 1
rlabel polysilicon 509 -1412 509 -1412 0 2
rlabel polysilicon 506 -1418 506 -1418 0 3
rlabel polysilicon 516 -1412 516 -1412 0 2
rlabel polysilicon 513 -1418 513 -1418 0 3
rlabel polysilicon 516 -1418 516 -1418 0 4
rlabel polysilicon 520 -1412 520 -1412 0 1
rlabel polysilicon 523 -1412 523 -1412 0 2
rlabel polysilicon 523 -1418 523 -1418 0 4
rlabel polysilicon 527 -1412 527 -1412 0 1
rlabel polysilicon 527 -1418 527 -1418 0 3
rlabel polysilicon 534 -1412 534 -1412 0 1
rlabel polysilicon 534 -1418 534 -1418 0 3
rlabel polysilicon 541 -1412 541 -1412 0 1
rlabel polysilicon 541 -1418 541 -1418 0 3
rlabel polysilicon 548 -1412 548 -1412 0 1
rlabel polysilicon 548 -1418 548 -1418 0 3
rlabel polysilicon 555 -1412 555 -1412 0 1
rlabel polysilicon 555 -1418 555 -1418 0 3
rlabel polysilicon 565 -1412 565 -1412 0 2
rlabel polysilicon 562 -1418 562 -1418 0 3
rlabel polysilicon 569 -1412 569 -1412 0 1
rlabel polysilicon 572 -1412 572 -1412 0 2
rlabel polysilicon 569 -1418 569 -1418 0 3
rlabel polysilicon 576 -1412 576 -1412 0 1
rlabel polysilicon 579 -1412 579 -1412 0 2
rlabel polysilicon 576 -1418 576 -1418 0 3
rlabel polysilicon 583 -1412 583 -1412 0 1
rlabel polysilicon 586 -1412 586 -1412 0 2
rlabel polysilicon 583 -1418 583 -1418 0 3
rlabel polysilicon 586 -1418 586 -1418 0 4
rlabel polysilicon 590 -1412 590 -1412 0 1
rlabel polysilicon 590 -1418 590 -1418 0 3
rlabel polysilicon 597 -1412 597 -1412 0 1
rlabel polysilicon 597 -1418 597 -1418 0 3
rlabel polysilicon 604 -1412 604 -1412 0 1
rlabel polysilicon 604 -1418 604 -1418 0 3
rlabel polysilicon 611 -1412 611 -1412 0 1
rlabel polysilicon 611 -1418 611 -1418 0 3
rlabel polysilicon 618 -1412 618 -1412 0 1
rlabel polysilicon 618 -1418 618 -1418 0 3
rlabel polysilicon 625 -1412 625 -1412 0 1
rlabel polysilicon 625 -1418 625 -1418 0 3
rlabel polysilicon 632 -1412 632 -1412 0 1
rlabel polysilicon 632 -1418 632 -1418 0 3
rlabel polysilicon 639 -1412 639 -1412 0 1
rlabel polysilicon 639 -1418 639 -1418 0 3
rlabel polysilicon 646 -1412 646 -1412 0 1
rlabel polysilicon 646 -1418 646 -1418 0 3
rlabel polysilicon 653 -1412 653 -1412 0 1
rlabel polysilicon 653 -1418 653 -1418 0 3
rlabel polysilicon 660 -1412 660 -1412 0 1
rlabel polysilicon 663 -1412 663 -1412 0 2
rlabel polysilicon 660 -1418 660 -1418 0 3
rlabel polysilicon 663 -1418 663 -1418 0 4
rlabel polysilicon 667 -1412 667 -1412 0 1
rlabel polysilicon 667 -1418 667 -1418 0 3
rlabel polysilicon 674 -1412 674 -1412 0 1
rlabel polysilicon 674 -1418 674 -1418 0 3
rlabel polysilicon 681 -1412 681 -1412 0 1
rlabel polysilicon 684 -1412 684 -1412 0 2
rlabel polysilicon 681 -1418 681 -1418 0 3
rlabel polysilicon 688 -1412 688 -1412 0 1
rlabel polysilicon 688 -1418 688 -1418 0 3
rlabel polysilicon 695 -1412 695 -1412 0 1
rlabel polysilicon 695 -1418 695 -1418 0 3
rlabel polysilicon 705 -1412 705 -1412 0 2
rlabel polysilicon 702 -1418 702 -1418 0 3
rlabel polysilicon 709 -1412 709 -1412 0 1
rlabel polysilicon 709 -1418 709 -1418 0 3
rlabel polysilicon 712 -1418 712 -1418 0 4
rlabel polysilicon 716 -1412 716 -1412 0 1
rlabel polysilicon 716 -1418 716 -1418 0 3
rlabel polysilicon 723 -1412 723 -1412 0 1
rlabel polysilicon 723 -1418 723 -1418 0 3
rlabel polysilicon 730 -1412 730 -1412 0 1
rlabel polysilicon 730 -1418 730 -1418 0 3
rlabel polysilicon 737 -1412 737 -1412 0 1
rlabel polysilicon 744 -1412 744 -1412 0 1
rlabel polysilicon 744 -1418 744 -1418 0 3
rlabel polysilicon 751 -1412 751 -1412 0 1
rlabel polysilicon 751 -1418 751 -1418 0 3
rlabel polysilicon 758 -1412 758 -1412 0 1
rlabel polysilicon 758 -1418 758 -1418 0 3
rlabel polysilicon 765 -1418 765 -1418 0 3
rlabel polysilicon 768 -1418 768 -1418 0 4
rlabel polysilicon 772 -1412 772 -1412 0 1
rlabel polysilicon 772 -1418 772 -1418 0 3
rlabel polysilicon 779 -1412 779 -1412 0 1
rlabel polysilicon 779 -1418 779 -1418 0 3
rlabel polysilicon 786 -1412 786 -1412 0 1
rlabel polysilicon 786 -1418 786 -1418 0 3
rlabel polysilicon 793 -1412 793 -1412 0 1
rlabel polysilicon 793 -1418 793 -1418 0 3
rlabel polysilicon 800 -1412 800 -1412 0 1
rlabel polysilicon 800 -1418 800 -1418 0 3
rlabel polysilicon 807 -1412 807 -1412 0 1
rlabel polysilicon 807 -1418 807 -1418 0 3
rlabel polysilicon 814 -1412 814 -1412 0 1
rlabel polysilicon 814 -1418 814 -1418 0 3
rlabel polysilicon 821 -1412 821 -1412 0 1
rlabel polysilicon 821 -1418 821 -1418 0 3
rlabel polysilicon 828 -1412 828 -1412 0 1
rlabel polysilicon 828 -1418 828 -1418 0 3
rlabel polysilicon 835 -1412 835 -1412 0 1
rlabel polysilicon 835 -1418 835 -1418 0 3
rlabel polysilicon 842 -1412 842 -1412 0 1
rlabel polysilicon 842 -1418 842 -1418 0 3
rlabel polysilicon 849 -1412 849 -1412 0 1
rlabel polysilicon 849 -1418 849 -1418 0 3
rlabel polysilicon 856 -1412 856 -1412 0 1
rlabel polysilicon 856 -1418 856 -1418 0 3
rlabel polysilicon 863 -1412 863 -1412 0 1
rlabel polysilicon 863 -1418 863 -1418 0 3
rlabel polysilicon 870 -1412 870 -1412 0 1
rlabel polysilicon 870 -1418 870 -1418 0 3
rlabel polysilicon 877 -1412 877 -1412 0 1
rlabel polysilicon 877 -1418 877 -1418 0 3
rlabel polysilicon 884 -1412 884 -1412 0 1
rlabel polysilicon 884 -1418 884 -1418 0 3
rlabel polysilicon 891 -1412 891 -1412 0 1
rlabel polysilicon 891 -1418 891 -1418 0 3
rlabel polysilicon 898 -1412 898 -1412 0 1
rlabel polysilicon 898 -1418 898 -1418 0 3
rlabel polysilicon 905 -1412 905 -1412 0 1
rlabel polysilicon 905 -1418 905 -1418 0 3
rlabel polysilicon 912 -1412 912 -1412 0 1
rlabel polysilicon 912 -1418 912 -1418 0 3
rlabel polysilicon 919 -1412 919 -1412 0 1
rlabel polysilicon 919 -1418 919 -1418 0 3
rlabel polysilicon 926 -1418 926 -1418 0 3
rlabel polysilicon 929 -1418 929 -1418 0 4
rlabel polysilicon 933 -1412 933 -1412 0 1
rlabel polysilicon 933 -1418 933 -1418 0 3
rlabel polysilicon 940 -1412 940 -1412 0 1
rlabel polysilicon 940 -1418 940 -1418 0 3
rlabel polysilicon 950 -1412 950 -1412 0 2
rlabel polysilicon 947 -1418 947 -1418 0 3
rlabel polysilicon 950 -1418 950 -1418 0 4
rlabel polysilicon 954 -1412 954 -1412 0 1
rlabel polysilicon 954 -1418 954 -1418 0 3
rlabel polysilicon 961 -1412 961 -1412 0 1
rlabel polysilicon 961 -1418 961 -1418 0 3
rlabel polysilicon 971 -1412 971 -1412 0 2
rlabel polysilicon 968 -1418 968 -1418 0 3
rlabel polysilicon 971 -1418 971 -1418 0 4
rlabel polysilicon 975 -1412 975 -1412 0 1
rlabel polysilicon 975 -1418 975 -1418 0 3
rlabel polysilicon 982 -1412 982 -1412 0 1
rlabel polysilicon 982 -1418 982 -1418 0 3
rlabel polysilicon 989 -1412 989 -1412 0 1
rlabel polysilicon 989 -1418 989 -1418 0 3
rlabel polysilicon 996 -1412 996 -1412 0 1
rlabel polysilicon 996 -1418 996 -1418 0 3
rlabel polysilicon 1003 -1412 1003 -1412 0 1
rlabel polysilicon 1006 -1418 1006 -1418 0 4
rlabel polysilicon 1010 -1412 1010 -1412 0 1
rlabel polysilicon 1010 -1418 1010 -1418 0 3
rlabel polysilicon 1017 -1412 1017 -1412 0 1
rlabel polysilicon 1017 -1418 1017 -1418 0 3
rlabel polysilicon 1024 -1412 1024 -1412 0 1
rlabel polysilicon 1024 -1418 1024 -1418 0 3
rlabel polysilicon 1031 -1412 1031 -1412 0 1
rlabel polysilicon 1031 -1418 1031 -1418 0 3
rlabel polysilicon 1041 -1418 1041 -1418 0 4
rlabel polysilicon 1045 -1412 1045 -1412 0 1
rlabel polysilicon 1045 -1418 1045 -1418 0 3
rlabel polysilicon 1052 -1412 1052 -1412 0 1
rlabel polysilicon 1052 -1418 1052 -1418 0 3
rlabel polysilicon 1073 -1412 1073 -1412 0 1
rlabel polysilicon 1073 -1418 1073 -1418 0 3
rlabel polysilicon 26 -1493 26 -1493 0 2
rlabel polysilicon 30 -1493 30 -1493 0 1
rlabel polysilicon 30 -1499 30 -1499 0 3
rlabel polysilicon 37 -1493 37 -1493 0 1
rlabel polysilicon 37 -1499 37 -1499 0 3
rlabel polysilicon 44 -1493 44 -1493 0 1
rlabel polysilicon 44 -1499 44 -1499 0 3
rlabel polysilicon 51 -1493 51 -1493 0 1
rlabel polysilicon 54 -1493 54 -1493 0 2
rlabel polysilicon 58 -1493 58 -1493 0 1
rlabel polysilicon 58 -1499 58 -1499 0 3
rlabel polysilicon 65 -1493 65 -1493 0 1
rlabel polysilicon 65 -1499 65 -1499 0 3
rlabel polysilicon 72 -1493 72 -1493 0 1
rlabel polysilicon 75 -1493 75 -1493 0 2
rlabel polysilicon 75 -1499 75 -1499 0 4
rlabel polysilicon 79 -1493 79 -1493 0 1
rlabel polysilicon 79 -1499 79 -1499 0 3
rlabel polysilicon 86 -1493 86 -1493 0 1
rlabel polysilicon 86 -1499 86 -1499 0 3
rlabel polysilicon 93 -1493 93 -1493 0 1
rlabel polysilicon 93 -1499 93 -1499 0 3
rlabel polysilicon 100 -1493 100 -1493 0 1
rlabel polysilicon 100 -1499 100 -1499 0 3
rlabel polysilicon 107 -1493 107 -1493 0 1
rlabel polysilicon 107 -1499 107 -1499 0 3
rlabel polysilicon 114 -1493 114 -1493 0 1
rlabel polysilicon 114 -1499 114 -1499 0 3
rlabel polysilicon 121 -1493 121 -1493 0 1
rlabel polysilicon 124 -1493 124 -1493 0 2
rlabel polysilicon 121 -1499 121 -1499 0 3
rlabel polysilicon 128 -1493 128 -1493 0 1
rlabel polysilicon 131 -1499 131 -1499 0 4
rlabel polysilicon 135 -1493 135 -1493 0 1
rlabel polysilicon 135 -1499 135 -1499 0 3
rlabel polysilicon 142 -1493 142 -1493 0 1
rlabel polysilicon 142 -1499 142 -1499 0 3
rlabel polysilicon 149 -1493 149 -1493 0 1
rlabel polysilicon 149 -1499 149 -1499 0 3
rlabel polysilicon 156 -1493 156 -1493 0 1
rlabel polysilicon 156 -1499 156 -1499 0 3
rlabel polysilicon 163 -1493 163 -1493 0 1
rlabel polysilicon 163 -1499 163 -1499 0 3
rlabel polysilicon 170 -1493 170 -1493 0 1
rlabel polysilicon 170 -1499 170 -1499 0 3
rlabel polysilicon 177 -1493 177 -1493 0 1
rlabel polysilicon 180 -1499 180 -1499 0 4
rlabel polysilicon 184 -1493 184 -1493 0 1
rlabel polysilicon 187 -1493 187 -1493 0 2
rlabel polysilicon 187 -1499 187 -1499 0 4
rlabel polysilicon 191 -1493 191 -1493 0 1
rlabel polysilicon 191 -1499 191 -1499 0 3
rlabel polysilicon 198 -1493 198 -1493 0 1
rlabel polysilicon 198 -1499 198 -1499 0 3
rlabel polysilicon 205 -1493 205 -1493 0 1
rlabel polysilicon 205 -1499 205 -1499 0 3
rlabel polysilicon 212 -1493 212 -1493 0 1
rlabel polysilicon 212 -1499 212 -1499 0 3
rlabel polysilicon 219 -1493 219 -1493 0 1
rlabel polysilicon 219 -1499 219 -1499 0 3
rlabel polysilicon 226 -1493 226 -1493 0 1
rlabel polysilicon 226 -1499 226 -1499 0 3
rlabel polysilicon 233 -1493 233 -1493 0 1
rlabel polysilicon 233 -1499 233 -1499 0 3
rlabel polysilicon 243 -1493 243 -1493 0 2
rlabel polysilicon 240 -1499 240 -1499 0 3
rlabel polysilicon 243 -1499 243 -1499 0 4
rlabel polysilicon 247 -1493 247 -1493 0 1
rlabel polysilicon 247 -1499 247 -1499 0 3
rlabel polysilicon 254 -1493 254 -1493 0 1
rlabel polysilicon 254 -1499 254 -1499 0 3
rlabel polysilicon 261 -1493 261 -1493 0 1
rlabel polysilicon 261 -1499 261 -1499 0 3
rlabel polysilicon 268 -1493 268 -1493 0 1
rlabel polysilicon 268 -1499 268 -1499 0 3
rlabel polysilicon 275 -1493 275 -1493 0 1
rlabel polysilicon 275 -1499 275 -1499 0 3
rlabel polysilicon 282 -1493 282 -1493 0 1
rlabel polysilicon 282 -1499 282 -1499 0 3
rlabel polysilicon 289 -1493 289 -1493 0 1
rlabel polysilicon 292 -1493 292 -1493 0 2
rlabel polysilicon 292 -1499 292 -1499 0 4
rlabel polysilicon 296 -1493 296 -1493 0 1
rlabel polysilicon 296 -1499 296 -1499 0 3
rlabel polysilicon 306 -1493 306 -1493 0 2
rlabel polysilicon 303 -1499 303 -1499 0 3
rlabel polysilicon 306 -1499 306 -1499 0 4
rlabel polysilicon 310 -1493 310 -1493 0 1
rlabel polysilicon 310 -1499 310 -1499 0 3
rlabel polysilicon 313 -1499 313 -1499 0 4
rlabel polysilicon 317 -1493 317 -1493 0 1
rlabel polysilicon 320 -1493 320 -1493 0 2
rlabel polysilicon 317 -1499 317 -1499 0 3
rlabel polysilicon 324 -1493 324 -1493 0 1
rlabel polysilicon 324 -1499 324 -1499 0 3
rlabel polysilicon 331 -1493 331 -1493 0 1
rlabel polysilicon 331 -1499 331 -1499 0 3
rlabel polysilicon 338 -1493 338 -1493 0 1
rlabel polysilicon 338 -1499 338 -1499 0 3
rlabel polysilicon 345 -1493 345 -1493 0 1
rlabel polysilicon 345 -1499 345 -1499 0 3
rlabel polysilicon 352 -1493 352 -1493 0 1
rlabel polysilicon 352 -1499 352 -1499 0 3
rlabel polysilicon 359 -1493 359 -1493 0 1
rlabel polysilicon 359 -1499 359 -1499 0 3
rlabel polysilicon 366 -1493 366 -1493 0 1
rlabel polysilicon 366 -1499 366 -1499 0 3
rlabel polysilicon 373 -1493 373 -1493 0 1
rlabel polysilicon 373 -1499 373 -1499 0 3
rlabel polysilicon 380 -1493 380 -1493 0 1
rlabel polysilicon 380 -1499 380 -1499 0 3
rlabel polysilicon 387 -1493 387 -1493 0 1
rlabel polysilicon 387 -1499 387 -1499 0 3
rlabel polysilicon 394 -1493 394 -1493 0 1
rlabel polysilicon 397 -1493 397 -1493 0 2
rlabel polysilicon 394 -1499 394 -1499 0 3
rlabel polysilicon 397 -1499 397 -1499 0 4
rlabel polysilicon 401 -1493 401 -1493 0 1
rlabel polysilicon 401 -1499 401 -1499 0 3
rlabel polysilicon 408 -1493 408 -1493 0 1
rlabel polysilicon 408 -1499 408 -1499 0 3
rlabel polysilicon 415 -1493 415 -1493 0 1
rlabel polysilicon 418 -1493 418 -1493 0 2
rlabel polysilicon 415 -1499 415 -1499 0 3
rlabel polysilicon 418 -1499 418 -1499 0 4
rlabel polysilicon 422 -1493 422 -1493 0 1
rlabel polysilicon 422 -1499 422 -1499 0 3
rlabel polysilicon 429 -1493 429 -1493 0 1
rlabel polysilicon 429 -1499 429 -1499 0 3
rlabel polysilicon 436 -1493 436 -1493 0 1
rlabel polysilicon 439 -1499 439 -1499 0 4
rlabel polysilicon 443 -1493 443 -1493 0 1
rlabel polysilicon 443 -1499 443 -1499 0 3
rlabel polysilicon 450 -1493 450 -1493 0 1
rlabel polysilicon 450 -1499 450 -1499 0 3
rlabel polysilicon 457 -1493 457 -1493 0 1
rlabel polysilicon 457 -1499 457 -1499 0 3
rlabel polysilicon 464 -1493 464 -1493 0 1
rlabel polysilicon 464 -1499 464 -1499 0 3
rlabel polysilicon 471 -1493 471 -1493 0 1
rlabel polysilicon 471 -1499 471 -1499 0 3
rlabel polysilicon 478 -1493 478 -1493 0 1
rlabel polysilicon 478 -1499 478 -1499 0 3
rlabel polysilicon 485 -1493 485 -1493 0 1
rlabel polysilicon 485 -1499 485 -1499 0 3
rlabel polysilicon 492 -1493 492 -1493 0 1
rlabel polysilicon 492 -1499 492 -1499 0 3
rlabel polysilicon 499 -1493 499 -1493 0 1
rlabel polysilicon 499 -1499 499 -1499 0 3
rlabel polysilicon 506 -1493 506 -1493 0 1
rlabel polysilicon 506 -1499 506 -1499 0 3
rlabel polysilicon 513 -1493 513 -1493 0 1
rlabel polysilicon 513 -1499 513 -1499 0 3
rlabel polysilicon 520 -1493 520 -1493 0 1
rlabel polysilicon 520 -1499 520 -1499 0 3
rlabel polysilicon 527 -1493 527 -1493 0 1
rlabel polysilicon 527 -1499 527 -1499 0 3
rlabel polysilicon 537 -1493 537 -1493 0 2
rlabel polysilicon 534 -1499 534 -1499 0 3
rlabel polysilicon 537 -1499 537 -1499 0 4
rlabel polysilicon 544 -1493 544 -1493 0 2
rlabel polysilicon 544 -1499 544 -1499 0 4
rlabel polysilicon 548 -1493 548 -1493 0 1
rlabel polysilicon 548 -1499 548 -1499 0 3
rlabel polysilicon 555 -1493 555 -1493 0 1
rlabel polysilicon 558 -1493 558 -1493 0 2
rlabel polysilicon 558 -1499 558 -1499 0 4
rlabel polysilicon 562 -1493 562 -1493 0 1
rlabel polysilicon 565 -1493 565 -1493 0 2
rlabel polysilicon 562 -1499 562 -1499 0 3
rlabel polysilicon 565 -1499 565 -1499 0 4
rlabel polysilicon 569 -1493 569 -1493 0 1
rlabel polysilicon 569 -1499 569 -1499 0 3
rlabel polysilicon 579 -1493 579 -1493 0 2
rlabel polysilicon 576 -1499 576 -1499 0 3
rlabel polysilicon 579 -1499 579 -1499 0 4
rlabel polysilicon 583 -1493 583 -1493 0 1
rlabel polysilicon 583 -1499 583 -1499 0 3
rlabel polysilicon 590 -1493 590 -1493 0 1
rlabel polysilicon 590 -1499 590 -1499 0 3
rlabel polysilicon 597 -1493 597 -1493 0 1
rlabel polysilicon 597 -1499 597 -1499 0 3
rlabel polysilicon 604 -1493 604 -1493 0 1
rlabel polysilicon 604 -1499 604 -1499 0 3
rlabel polysilicon 611 -1493 611 -1493 0 1
rlabel polysilicon 611 -1499 611 -1499 0 3
rlabel polysilicon 618 -1493 618 -1493 0 1
rlabel polysilicon 618 -1499 618 -1499 0 3
rlabel polysilicon 625 -1493 625 -1493 0 1
rlabel polysilicon 625 -1499 625 -1499 0 3
rlabel polysilicon 635 -1493 635 -1493 0 2
rlabel polysilicon 639 -1493 639 -1493 0 1
rlabel polysilicon 639 -1499 639 -1499 0 3
rlabel polysilicon 646 -1493 646 -1493 0 1
rlabel polysilicon 646 -1499 646 -1499 0 3
rlabel polysilicon 656 -1493 656 -1493 0 2
rlabel polysilicon 653 -1499 653 -1499 0 3
rlabel polysilicon 656 -1499 656 -1499 0 4
rlabel polysilicon 660 -1493 660 -1493 0 1
rlabel polysilicon 660 -1499 660 -1499 0 3
rlabel polysilicon 667 -1493 667 -1493 0 1
rlabel polysilicon 667 -1499 667 -1499 0 3
rlabel polysilicon 674 -1493 674 -1493 0 1
rlabel polysilicon 674 -1499 674 -1499 0 3
rlabel polysilicon 681 -1493 681 -1493 0 1
rlabel polysilicon 684 -1493 684 -1493 0 2
rlabel polysilicon 681 -1499 681 -1499 0 3
rlabel polysilicon 684 -1499 684 -1499 0 4
rlabel polysilicon 688 -1493 688 -1493 0 1
rlabel polysilicon 688 -1499 688 -1499 0 3
rlabel polysilicon 695 -1493 695 -1493 0 1
rlabel polysilicon 695 -1499 695 -1499 0 3
rlabel polysilicon 702 -1493 702 -1493 0 1
rlabel polysilicon 702 -1499 702 -1499 0 3
rlabel polysilicon 709 -1493 709 -1493 0 1
rlabel polysilicon 709 -1499 709 -1499 0 3
rlabel polysilicon 716 -1493 716 -1493 0 1
rlabel polysilicon 716 -1499 716 -1499 0 3
rlabel polysilicon 726 -1493 726 -1493 0 2
rlabel polysilicon 723 -1499 723 -1499 0 3
rlabel polysilicon 726 -1499 726 -1499 0 4
rlabel polysilicon 730 -1493 730 -1493 0 1
rlabel polysilicon 730 -1499 730 -1499 0 3
rlabel polysilicon 737 -1493 737 -1493 0 1
rlabel polysilicon 737 -1499 737 -1499 0 3
rlabel polysilicon 744 -1493 744 -1493 0 1
rlabel polysilicon 744 -1499 744 -1499 0 3
rlabel polysilicon 751 -1493 751 -1493 0 1
rlabel polysilicon 751 -1499 751 -1499 0 3
rlabel polysilicon 758 -1493 758 -1493 0 1
rlabel polysilicon 758 -1499 758 -1499 0 3
rlabel polysilicon 765 -1493 765 -1493 0 1
rlabel polysilicon 765 -1499 765 -1499 0 3
rlabel polysilicon 772 -1493 772 -1493 0 1
rlabel polysilicon 772 -1499 772 -1499 0 3
rlabel polysilicon 779 -1493 779 -1493 0 1
rlabel polysilicon 779 -1499 779 -1499 0 3
rlabel polysilicon 786 -1493 786 -1493 0 1
rlabel polysilicon 786 -1499 786 -1499 0 3
rlabel polysilicon 793 -1493 793 -1493 0 1
rlabel polysilicon 793 -1499 793 -1499 0 3
rlabel polysilicon 800 -1499 800 -1499 0 3
rlabel polysilicon 803 -1499 803 -1499 0 4
rlabel polysilicon 807 -1493 807 -1493 0 1
rlabel polysilicon 807 -1499 807 -1499 0 3
rlabel polysilicon 814 -1493 814 -1493 0 1
rlabel polysilicon 814 -1499 814 -1499 0 3
rlabel polysilicon 821 -1493 821 -1493 0 1
rlabel polysilicon 821 -1499 821 -1499 0 3
rlabel polysilicon 828 -1493 828 -1493 0 1
rlabel polysilicon 828 -1499 828 -1499 0 3
rlabel polysilicon 835 -1493 835 -1493 0 1
rlabel polysilicon 835 -1499 835 -1499 0 3
rlabel polysilicon 842 -1493 842 -1493 0 1
rlabel polysilicon 842 -1499 842 -1499 0 3
rlabel polysilicon 849 -1493 849 -1493 0 1
rlabel polysilicon 849 -1499 849 -1499 0 3
rlabel polysilicon 856 -1493 856 -1493 0 1
rlabel polysilicon 856 -1499 856 -1499 0 3
rlabel polysilicon 863 -1493 863 -1493 0 1
rlabel polysilicon 863 -1499 863 -1499 0 3
rlabel polysilicon 870 -1493 870 -1493 0 1
rlabel polysilicon 870 -1499 870 -1499 0 3
rlabel polysilicon 877 -1493 877 -1493 0 1
rlabel polysilicon 877 -1499 877 -1499 0 3
rlabel polysilicon 884 -1493 884 -1493 0 1
rlabel polysilicon 884 -1499 884 -1499 0 3
rlabel polysilicon 891 -1493 891 -1493 0 1
rlabel polysilicon 891 -1499 891 -1499 0 3
rlabel polysilicon 898 -1493 898 -1493 0 1
rlabel polysilicon 898 -1499 898 -1499 0 3
rlabel polysilicon 905 -1493 905 -1493 0 1
rlabel polysilicon 905 -1499 905 -1499 0 3
rlabel polysilicon 912 -1493 912 -1493 0 1
rlabel polysilicon 912 -1499 912 -1499 0 3
rlabel polysilicon 919 -1493 919 -1493 0 1
rlabel polysilicon 922 -1493 922 -1493 0 2
rlabel polysilicon 922 -1499 922 -1499 0 4
rlabel polysilicon 926 -1493 926 -1493 0 1
rlabel polysilicon 926 -1499 926 -1499 0 3
rlabel polysilicon 933 -1493 933 -1493 0 1
rlabel polysilicon 933 -1499 933 -1499 0 3
rlabel polysilicon 940 -1493 940 -1493 0 1
rlabel polysilicon 943 -1493 943 -1493 0 2
rlabel polysilicon 947 -1493 947 -1493 0 1
rlabel polysilicon 947 -1499 947 -1499 0 3
rlabel polysilicon 954 -1493 954 -1493 0 1
rlabel polysilicon 954 -1499 954 -1499 0 3
rlabel polysilicon 964 -1499 964 -1499 0 4
rlabel polysilicon 971 -1493 971 -1493 0 2
rlabel polysilicon 971 -1499 971 -1499 0 4
rlabel polysilicon 975 -1493 975 -1493 0 1
rlabel polysilicon 975 -1499 975 -1499 0 3
rlabel polysilicon 982 -1493 982 -1493 0 1
rlabel polysilicon 982 -1499 982 -1499 0 3
rlabel polysilicon 989 -1493 989 -1493 0 1
rlabel polysilicon 989 -1499 989 -1499 0 3
rlabel polysilicon 996 -1493 996 -1493 0 1
rlabel polysilicon 996 -1499 996 -1499 0 3
rlabel polysilicon 1003 -1493 1003 -1493 0 1
rlabel polysilicon 1003 -1499 1003 -1499 0 3
rlabel polysilicon 1038 -1493 1038 -1493 0 1
rlabel polysilicon 1038 -1499 1038 -1499 0 3
rlabel polysilicon 1066 -1493 1066 -1493 0 1
rlabel polysilicon 2 -1590 2 -1590 0 1
rlabel polysilicon 2 -1596 2 -1596 0 3
rlabel polysilicon 9 -1590 9 -1590 0 1
rlabel polysilicon 9 -1596 9 -1596 0 3
rlabel polysilicon 16 -1590 16 -1590 0 1
rlabel polysilicon 16 -1596 16 -1596 0 3
rlabel polysilicon 23 -1590 23 -1590 0 1
rlabel polysilicon 23 -1596 23 -1596 0 3
rlabel polysilicon 30 -1590 30 -1590 0 1
rlabel polysilicon 30 -1596 30 -1596 0 3
rlabel polysilicon 37 -1590 37 -1590 0 1
rlabel polysilicon 37 -1596 37 -1596 0 3
rlabel polysilicon 47 -1596 47 -1596 0 4
rlabel polysilicon 51 -1590 51 -1590 0 1
rlabel polysilicon 51 -1596 51 -1596 0 3
rlabel polysilicon 58 -1590 58 -1590 0 1
rlabel polysilicon 58 -1596 58 -1596 0 3
rlabel polysilicon 65 -1590 65 -1590 0 1
rlabel polysilicon 65 -1596 65 -1596 0 3
rlabel polysilicon 72 -1590 72 -1590 0 1
rlabel polysilicon 72 -1596 72 -1596 0 3
rlabel polysilicon 75 -1596 75 -1596 0 4
rlabel polysilicon 79 -1590 79 -1590 0 1
rlabel polysilicon 82 -1590 82 -1590 0 2
rlabel polysilicon 82 -1596 82 -1596 0 4
rlabel polysilicon 86 -1590 86 -1590 0 1
rlabel polysilicon 86 -1596 86 -1596 0 3
rlabel polysilicon 93 -1590 93 -1590 0 1
rlabel polysilicon 93 -1596 93 -1596 0 3
rlabel polysilicon 100 -1590 100 -1590 0 1
rlabel polysilicon 100 -1596 100 -1596 0 3
rlabel polysilicon 107 -1590 107 -1590 0 1
rlabel polysilicon 107 -1596 107 -1596 0 3
rlabel polysilicon 114 -1590 114 -1590 0 1
rlabel polysilicon 114 -1596 114 -1596 0 3
rlabel polysilicon 124 -1590 124 -1590 0 2
rlabel polysilicon 121 -1596 121 -1596 0 3
rlabel polysilicon 124 -1596 124 -1596 0 4
rlabel polysilicon 128 -1590 128 -1590 0 1
rlabel polysilicon 128 -1596 128 -1596 0 3
rlabel polysilicon 135 -1590 135 -1590 0 1
rlabel polysilicon 135 -1596 135 -1596 0 3
rlabel polysilicon 142 -1590 142 -1590 0 1
rlabel polysilicon 142 -1596 142 -1596 0 3
rlabel polysilicon 149 -1590 149 -1590 0 1
rlabel polysilicon 149 -1596 149 -1596 0 3
rlabel polysilicon 156 -1590 156 -1590 0 1
rlabel polysilicon 156 -1596 156 -1596 0 3
rlabel polysilicon 163 -1590 163 -1590 0 1
rlabel polysilicon 163 -1596 163 -1596 0 3
rlabel polysilicon 170 -1590 170 -1590 0 1
rlabel polysilicon 170 -1596 170 -1596 0 3
rlabel polysilicon 177 -1590 177 -1590 0 1
rlabel polysilicon 177 -1596 177 -1596 0 3
rlabel polysilicon 184 -1590 184 -1590 0 1
rlabel polysilicon 184 -1596 184 -1596 0 3
rlabel polysilicon 194 -1590 194 -1590 0 2
rlabel polysilicon 194 -1596 194 -1596 0 4
rlabel polysilicon 198 -1590 198 -1590 0 1
rlabel polysilicon 198 -1596 198 -1596 0 3
rlabel polysilicon 205 -1590 205 -1590 0 1
rlabel polysilicon 205 -1596 205 -1596 0 3
rlabel polysilicon 212 -1590 212 -1590 0 1
rlabel polysilicon 212 -1596 212 -1596 0 3
rlabel polysilicon 222 -1590 222 -1590 0 2
rlabel polysilicon 222 -1596 222 -1596 0 4
rlabel polysilicon 226 -1590 226 -1590 0 1
rlabel polysilicon 229 -1590 229 -1590 0 2
rlabel polysilicon 226 -1596 226 -1596 0 3
rlabel polysilicon 233 -1590 233 -1590 0 1
rlabel polysilicon 233 -1596 233 -1596 0 3
rlabel polysilicon 240 -1590 240 -1590 0 1
rlabel polysilicon 243 -1590 243 -1590 0 2
rlabel polysilicon 243 -1596 243 -1596 0 4
rlabel polysilicon 247 -1590 247 -1590 0 1
rlabel polysilicon 247 -1596 247 -1596 0 3
rlabel polysilicon 250 -1596 250 -1596 0 4
rlabel polysilicon 254 -1590 254 -1590 0 1
rlabel polysilicon 254 -1596 254 -1596 0 3
rlabel polysilicon 261 -1590 261 -1590 0 1
rlabel polysilicon 261 -1596 261 -1596 0 3
rlabel polysilicon 268 -1590 268 -1590 0 1
rlabel polysilicon 268 -1596 268 -1596 0 3
rlabel polysilicon 275 -1590 275 -1590 0 1
rlabel polysilicon 275 -1596 275 -1596 0 3
rlabel polysilicon 282 -1590 282 -1590 0 1
rlabel polysilicon 282 -1596 282 -1596 0 3
rlabel polysilicon 289 -1590 289 -1590 0 1
rlabel polysilicon 289 -1596 289 -1596 0 3
rlabel polysilicon 296 -1590 296 -1590 0 1
rlabel polysilicon 296 -1596 296 -1596 0 3
rlabel polysilicon 303 -1590 303 -1590 0 1
rlabel polysilicon 303 -1596 303 -1596 0 3
rlabel polysilicon 310 -1590 310 -1590 0 1
rlabel polysilicon 310 -1596 310 -1596 0 3
rlabel polysilicon 317 -1590 317 -1590 0 1
rlabel polysilicon 317 -1596 317 -1596 0 3
rlabel polysilicon 324 -1590 324 -1590 0 1
rlabel polysilicon 327 -1590 327 -1590 0 2
rlabel polysilicon 331 -1590 331 -1590 0 1
rlabel polysilicon 331 -1596 331 -1596 0 3
rlabel polysilicon 338 -1590 338 -1590 0 1
rlabel polysilicon 341 -1590 341 -1590 0 2
rlabel polysilicon 338 -1596 338 -1596 0 3
rlabel polysilicon 341 -1596 341 -1596 0 4
rlabel polysilicon 345 -1590 345 -1590 0 1
rlabel polysilicon 345 -1596 345 -1596 0 3
rlabel polysilicon 352 -1590 352 -1590 0 1
rlabel polysilicon 355 -1590 355 -1590 0 2
rlabel polysilicon 355 -1596 355 -1596 0 4
rlabel polysilicon 359 -1590 359 -1590 0 1
rlabel polysilicon 362 -1590 362 -1590 0 2
rlabel polysilicon 362 -1596 362 -1596 0 4
rlabel polysilicon 366 -1590 366 -1590 0 1
rlabel polysilicon 366 -1596 366 -1596 0 3
rlabel polysilicon 373 -1590 373 -1590 0 1
rlabel polysilicon 376 -1590 376 -1590 0 2
rlabel polysilicon 373 -1596 373 -1596 0 3
rlabel polysilicon 376 -1596 376 -1596 0 4
rlabel polysilicon 380 -1590 380 -1590 0 1
rlabel polysilicon 380 -1596 380 -1596 0 3
rlabel polysilicon 387 -1590 387 -1590 0 1
rlabel polysilicon 387 -1596 387 -1596 0 3
rlabel polysilicon 394 -1590 394 -1590 0 1
rlabel polysilicon 397 -1590 397 -1590 0 2
rlabel polysilicon 394 -1596 394 -1596 0 3
rlabel polysilicon 401 -1590 401 -1590 0 1
rlabel polysilicon 401 -1596 401 -1596 0 3
rlabel polysilicon 408 -1590 408 -1590 0 1
rlabel polysilicon 408 -1596 408 -1596 0 3
rlabel polysilicon 418 -1590 418 -1590 0 2
rlabel polysilicon 422 -1590 422 -1590 0 1
rlabel polysilicon 422 -1596 422 -1596 0 3
rlabel polysilicon 429 -1590 429 -1590 0 1
rlabel polysilicon 429 -1596 429 -1596 0 3
rlabel polysilicon 436 -1590 436 -1590 0 1
rlabel polysilicon 439 -1590 439 -1590 0 2
rlabel polysilicon 436 -1596 436 -1596 0 3
rlabel polysilicon 443 -1590 443 -1590 0 1
rlabel polysilicon 443 -1596 443 -1596 0 3
rlabel polysilicon 450 -1590 450 -1590 0 1
rlabel polysilicon 450 -1596 450 -1596 0 3
rlabel polysilicon 453 -1596 453 -1596 0 4
rlabel polysilicon 457 -1590 457 -1590 0 1
rlabel polysilicon 460 -1590 460 -1590 0 2
rlabel polysilicon 457 -1596 457 -1596 0 3
rlabel polysilicon 460 -1596 460 -1596 0 4
rlabel polysilicon 464 -1590 464 -1590 0 1
rlabel polysilicon 464 -1596 464 -1596 0 3
rlabel polysilicon 471 -1590 471 -1590 0 1
rlabel polysilicon 474 -1590 474 -1590 0 2
rlabel polysilicon 471 -1596 471 -1596 0 3
rlabel polysilicon 474 -1596 474 -1596 0 4
rlabel polysilicon 478 -1590 478 -1590 0 1
rlabel polysilicon 478 -1596 478 -1596 0 3
rlabel polysilicon 485 -1590 485 -1590 0 1
rlabel polysilicon 485 -1596 485 -1596 0 3
rlabel polysilicon 495 -1590 495 -1590 0 2
rlabel polysilicon 492 -1596 492 -1596 0 3
rlabel polysilicon 499 -1590 499 -1590 0 1
rlabel polysilicon 499 -1596 499 -1596 0 3
rlabel polysilicon 506 -1590 506 -1590 0 1
rlabel polysilicon 506 -1596 506 -1596 0 3
rlabel polysilicon 513 -1590 513 -1590 0 1
rlabel polysilicon 516 -1590 516 -1590 0 2
rlabel polysilicon 513 -1596 513 -1596 0 3
rlabel polysilicon 520 -1590 520 -1590 0 1
rlabel polysilicon 520 -1596 520 -1596 0 3
rlabel polysilicon 527 -1590 527 -1590 0 1
rlabel polysilicon 527 -1596 527 -1596 0 3
rlabel polysilicon 534 -1590 534 -1590 0 1
rlabel polysilicon 537 -1596 537 -1596 0 4
rlabel polysilicon 544 -1590 544 -1590 0 2
rlabel polysilicon 544 -1596 544 -1596 0 4
rlabel polysilicon 548 -1590 548 -1590 0 1
rlabel polysilicon 548 -1596 548 -1596 0 3
rlabel polysilicon 555 -1590 555 -1590 0 1
rlabel polysilicon 555 -1596 555 -1596 0 3
rlabel polysilicon 562 -1590 562 -1590 0 1
rlabel polysilicon 562 -1596 562 -1596 0 3
rlabel polysilicon 569 -1590 569 -1590 0 1
rlabel polysilicon 569 -1596 569 -1596 0 3
rlabel polysilicon 576 -1590 576 -1590 0 1
rlabel polysilicon 576 -1596 576 -1596 0 3
rlabel polysilicon 583 -1590 583 -1590 0 1
rlabel polysilicon 583 -1596 583 -1596 0 3
rlabel polysilicon 590 -1590 590 -1590 0 1
rlabel polysilicon 590 -1596 590 -1596 0 3
rlabel polysilicon 597 -1590 597 -1590 0 1
rlabel polysilicon 597 -1596 597 -1596 0 3
rlabel polysilicon 604 -1590 604 -1590 0 1
rlabel polysilicon 604 -1596 604 -1596 0 3
rlabel polysilicon 611 -1590 611 -1590 0 1
rlabel polysilicon 611 -1596 611 -1596 0 3
rlabel polysilicon 618 -1590 618 -1590 0 1
rlabel polysilicon 618 -1596 618 -1596 0 3
rlabel polysilicon 625 -1590 625 -1590 0 1
rlabel polysilicon 625 -1596 625 -1596 0 3
rlabel polysilicon 632 -1590 632 -1590 0 1
rlabel polysilicon 632 -1596 632 -1596 0 3
rlabel polysilicon 639 -1590 639 -1590 0 1
rlabel polysilicon 639 -1596 639 -1596 0 3
rlabel polysilicon 646 -1590 646 -1590 0 1
rlabel polysilicon 646 -1596 646 -1596 0 3
rlabel polysilicon 653 -1590 653 -1590 0 1
rlabel polysilicon 653 -1596 653 -1596 0 3
rlabel polysilicon 660 -1590 660 -1590 0 1
rlabel polysilicon 663 -1590 663 -1590 0 2
rlabel polysilicon 663 -1596 663 -1596 0 4
rlabel polysilicon 667 -1590 667 -1590 0 1
rlabel polysilicon 667 -1596 667 -1596 0 3
rlabel polysilicon 674 -1590 674 -1590 0 1
rlabel polysilicon 674 -1596 674 -1596 0 3
rlabel polysilicon 681 -1590 681 -1590 0 1
rlabel polysilicon 684 -1590 684 -1590 0 2
rlabel polysilicon 684 -1596 684 -1596 0 4
rlabel polysilicon 688 -1590 688 -1590 0 1
rlabel polysilicon 688 -1596 688 -1596 0 3
rlabel polysilicon 695 -1590 695 -1590 0 1
rlabel polysilicon 695 -1596 695 -1596 0 3
rlabel polysilicon 702 -1590 702 -1590 0 1
rlabel polysilicon 702 -1596 702 -1596 0 3
rlabel polysilicon 709 -1590 709 -1590 0 1
rlabel polysilicon 712 -1590 712 -1590 0 2
rlabel polysilicon 709 -1596 709 -1596 0 3
rlabel polysilicon 716 -1590 716 -1590 0 1
rlabel polysilicon 716 -1596 716 -1596 0 3
rlabel polysilicon 723 -1590 723 -1590 0 1
rlabel polysilicon 723 -1596 723 -1596 0 3
rlabel polysilicon 733 -1590 733 -1590 0 2
rlabel polysilicon 730 -1596 730 -1596 0 3
rlabel polysilicon 733 -1596 733 -1596 0 4
rlabel polysilicon 737 -1590 737 -1590 0 1
rlabel polysilicon 737 -1596 737 -1596 0 3
rlabel polysilicon 744 -1590 744 -1590 0 1
rlabel polysilicon 744 -1596 744 -1596 0 3
rlabel polysilicon 751 -1590 751 -1590 0 1
rlabel polysilicon 751 -1596 751 -1596 0 3
rlabel polysilicon 758 -1590 758 -1590 0 1
rlabel polysilicon 758 -1596 758 -1596 0 3
rlabel polysilicon 765 -1590 765 -1590 0 1
rlabel polysilicon 765 -1596 765 -1596 0 3
rlabel polysilicon 772 -1590 772 -1590 0 1
rlabel polysilicon 772 -1596 772 -1596 0 3
rlabel polysilicon 779 -1590 779 -1590 0 1
rlabel polysilicon 779 -1596 779 -1596 0 3
rlabel polysilicon 786 -1590 786 -1590 0 1
rlabel polysilicon 786 -1596 786 -1596 0 3
rlabel polysilicon 793 -1590 793 -1590 0 1
rlabel polysilicon 793 -1596 793 -1596 0 3
rlabel polysilicon 800 -1590 800 -1590 0 1
rlabel polysilicon 803 -1590 803 -1590 0 2
rlabel polysilicon 803 -1596 803 -1596 0 4
rlabel polysilicon 807 -1590 807 -1590 0 1
rlabel polysilicon 807 -1596 807 -1596 0 3
rlabel polysilicon 814 -1590 814 -1590 0 1
rlabel polysilicon 814 -1596 814 -1596 0 3
rlabel polysilicon 821 -1590 821 -1590 0 1
rlabel polysilicon 821 -1596 821 -1596 0 3
rlabel polysilicon 828 -1590 828 -1590 0 1
rlabel polysilicon 828 -1596 828 -1596 0 3
rlabel polysilicon 835 -1590 835 -1590 0 1
rlabel polysilicon 835 -1596 835 -1596 0 3
rlabel polysilicon 842 -1590 842 -1590 0 1
rlabel polysilicon 842 -1596 842 -1596 0 3
rlabel polysilicon 849 -1590 849 -1590 0 1
rlabel polysilicon 849 -1596 849 -1596 0 3
rlabel polysilicon 856 -1590 856 -1590 0 1
rlabel polysilicon 856 -1596 856 -1596 0 3
rlabel polysilicon 863 -1590 863 -1590 0 1
rlabel polysilicon 863 -1596 863 -1596 0 3
rlabel polysilicon 870 -1590 870 -1590 0 1
rlabel polysilicon 870 -1596 870 -1596 0 3
rlabel polysilicon 877 -1590 877 -1590 0 1
rlabel polysilicon 877 -1596 877 -1596 0 3
rlabel polysilicon 884 -1590 884 -1590 0 1
rlabel polysilicon 884 -1596 884 -1596 0 3
rlabel polysilicon 891 -1590 891 -1590 0 1
rlabel polysilicon 891 -1596 891 -1596 0 3
rlabel polysilicon 898 -1590 898 -1590 0 1
rlabel polysilicon 898 -1596 898 -1596 0 3
rlabel polysilicon 905 -1590 905 -1590 0 1
rlabel polysilicon 905 -1596 905 -1596 0 3
rlabel polysilicon 912 -1590 912 -1590 0 1
rlabel polysilicon 912 -1596 912 -1596 0 3
rlabel polysilicon 919 -1590 919 -1590 0 1
rlabel polysilicon 919 -1596 919 -1596 0 3
rlabel polysilicon 926 -1590 926 -1590 0 1
rlabel polysilicon 926 -1596 926 -1596 0 3
rlabel polysilicon 933 -1590 933 -1590 0 1
rlabel polysilicon 933 -1596 933 -1596 0 3
rlabel polysilicon 940 -1590 940 -1590 0 1
rlabel polysilicon 940 -1596 940 -1596 0 3
rlabel polysilicon 947 -1590 947 -1590 0 1
rlabel polysilicon 947 -1596 947 -1596 0 3
rlabel polysilicon 954 -1590 954 -1590 0 1
rlabel polysilicon 954 -1596 954 -1596 0 3
rlabel polysilicon 961 -1590 961 -1590 0 1
rlabel polysilicon 961 -1596 961 -1596 0 3
rlabel polysilicon 968 -1590 968 -1590 0 1
rlabel polysilicon 968 -1596 968 -1596 0 3
rlabel polysilicon 975 -1590 975 -1590 0 1
rlabel polysilicon 975 -1596 975 -1596 0 3
rlabel polysilicon 982 -1590 982 -1590 0 1
rlabel polysilicon 982 -1596 982 -1596 0 3
rlabel polysilicon 989 -1590 989 -1590 0 1
rlabel polysilicon 989 -1596 989 -1596 0 3
rlabel polysilicon 996 -1590 996 -1590 0 1
rlabel polysilicon 996 -1596 996 -1596 0 3
rlabel polysilicon 1003 -1590 1003 -1590 0 1
rlabel polysilicon 1003 -1596 1003 -1596 0 3
rlabel polysilicon 1010 -1590 1010 -1590 0 1
rlabel polysilicon 1010 -1596 1010 -1596 0 3
rlabel polysilicon 1017 -1590 1017 -1590 0 1
rlabel polysilicon 1017 -1596 1017 -1596 0 3
rlabel polysilicon 1024 -1590 1024 -1590 0 1
rlabel polysilicon 1024 -1596 1024 -1596 0 3
rlabel polysilicon 1031 -1590 1031 -1590 0 1
rlabel polysilicon 1031 -1596 1031 -1596 0 3
rlabel polysilicon 1038 -1590 1038 -1590 0 1
rlabel polysilicon 1038 -1596 1038 -1596 0 3
rlabel polysilicon 1045 -1590 1045 -1590 0 1
rlabel polysilicon 1045 -1596 1045 -1596 0 3
rlabel polysilicon 1052 -1590 1052 -1590 0 1
rlabel polysilicon 1052 -1596 1052 -1596 0 3
rlabel polysilicon 1059 -1590 1059 -1590 0 1
rlabel polysilicon 1059 -1596 1059 -1596 0 3
rlabel polysilicon 1066 -1590 1066 -1590 0 1
rlabel polysilicon 1066 -1596 1066 -1596 0 3
rlabel polysilicon 1073 -1590 1073 -1590 0 1
rlabel polysilicon 1073 -1596 1073 -1596 0 3
rlabel polysilicon 1080 -1590 1080 -1590 0 1
rlabel polysilicon 1080 -1596 1080 -1596 0 3
rlabel polysilicon 1087 -1590 1087 -1590 0 1
rlabel polysilicon 1087 -1596 1087 -1596 0 3
rlabel polysilicon 1094 -1590 1094 -1590 0 1
rlabel polysilicon 1094 -1596 1094 -1596 0 3
rlabel polysilicon 1101 -1590 1101 -1590 0 1
rlabel polysilicon 1101 -1596 1101 -1596 0 3
rlabel polysilicon 1108 -1590 1108 -1590 0 1
rlabel polysilicon 1111 -1590 1111 -1590 0 2
rlabel polysilicon 1108 -1596 1108 -1596 0 3
rlabel polysilicon 2 -1677 2 -1677 0 1
rlabel polysilicon 2 -1683 2 -1683 0 3
rlabel polysilicon 9 -1677 9 -1677 0 1
rlabel polysilicon 9 -1683 9 -1683 0 3
rlabel polysilicon 16 -1677 16 -1677 0 1
rlabel polysilicon 16 -1683 16 -1683 0 3
rlabel polysilicon 23 -1677 23 -1677 0 1
rlabel polysilicon 23 -1683 23 -1683 0 3
rlabel polysilicon 30 -1677 30 -1677 0 1
rlabel polysilicon 30 -1683 30 -1683 0 3
rlabel polysilicon 37 -1677 37 -1677 0 1
rlabel polysilicon 37 -1683 37 -1683 0 3
rlabel polysilicon 44 -1677 44 -1677 0 1
rlabel polysilicon 44 -1683 44 -1683 0 3
rlabel polysilicon 51 -1677 51 -1677 0 1
rlabel polysilicon 51 -1683 51 -1683 0 3
rlabel polysilicon 61 -1677 61 -1677 0 2
rlabel polysilicon 65 -1677 65 -1677 0 1
rlabel polysilicon 65 -1683 65 -1683 0 3
rlabel polysilicon 72 -1677 72 -1677 0 1
rlabel polysilicon 72 -1683 72 -1683 0 3
rlabel polysilicon 79 -1677 79 -1677 0 1
rlabel polysilicon 86 -1677 86 -1677 0 1
rlabel polysilicon 86 -1683 86 -1683 0 3
rlabel polysilicon 96 -1683 96 -1683 0 4
rlabel polysilicon 100 -1677 100 -1677 0 1
rlabel polysilicon 100 -1683 100 -1683 0 3
rlabel polysilicon 107 -1677 107 -1677 0 1
rlabel polysilicon 107 -1683 107 -1683 0 3
rlabel polysilicon 114 -1677 114 -1677 0 1
rlabel polysilicon 114 -1683 114 -1683 0 3
rlabel polysilicon 121 -1677 121 -1677 0 1
rlabel polysilicon 121 -1683 121 -1683 0 3
rlabel polysilicon 128 -1677 128 -1677 0 1
rlabel polysilicon 128 -1683 128 -1683 0 3
rlabel polysilicon 135 -1677 135 -1677 0 1
rlabel polysilicon 138 -1677 138 -1677 0 2
rlabel polysilicon 138 -1683 138 -1683 0 4
rlabel polysilicon 142 -1677 142 -1677 0 1
rlabel polysilicon 142 -1683 142 -1683 0 3
rlabel polysilicon 149 -1677 149 -1677 0 1
rlabel polysilicon 149 -1683 149 -1683 0 3
rlabel polysilicon 152 -1683 152 -1683 0 4
rlabel polysilicon 159 -1677 159 -1677 0 2
rlabel polysilicon 156 -1683 156 -1683 0 3
rlabel polysilicon 163 -1677 163 -1677 0 1
rlabel polysilicon 163 -1683 163 -1683 0 3
rlabel polysilicon 170 -1677 170 -1677 0 1
rlabel polysilicon 170 -1683 170 -1683 0 3
rlabel polysilicon 177 -1677 177 -1677 0 1
rlabel polysilicon 177 -1683 177 -1683 0 3
rlabel polysilicon 184 -1677 184 -1677 0 1
rlabel polysilicon 184 -1683 184 -1683 0 3
rlabel polysilicon 194 -1677 194 -1677 0 2
rlabel polysilicon 191 -1683 191 -1683 0 3
rlabel polysilicon 194 -1683 194 -1683 0 4
rlabel polysilicon 198 -1677 198 -1677 0 1
rlabel polysilicon 198 -1683 198 -1683 0 3
rlabel polysilicon 201 -1683 201 -1683 0 4
rlabel polysilicon 205 -1677 205 -1677 0 1
rlabel polysilicon 205 -1683 205 -1683 0 3
rlabel polysilicon 212 -1677 212 -1677 0 1
rlabel polysilicon 215 -1683 215 -1683 0 4
rlabel polysilicon 222 -1677 222 -1677 0 2
rlabel polysilicon 222 -1683 222 -1683 0 4
rlabel polysilicon 226 -1677 226 -1677 0 1
rlabel polysilicon 226 -1683 226 -1683 0 3
rlabel polysilicon 229 -1683 229 -1683 0 4
rlabel polysilicon 233 -1677 233 -1677 0 1
rlabel polysilicon 236 -1677 236 -1677 0 2
rlabel polysilicon 240 -1677 240 -1677 0 1
rlabel polysilicon 240 -1683 240 -1683 0 3
rlabel polysilicon 247 -1677 247 -1677 0 1
rlabel polysilicon 247 -1683 247 -1683 0 3
rlabel polysilicon 254 -1677 254 -1677 0 1
rlabel polysilicon 254 -1683 254 -1683 0 3
rlabel polysilicon 261 -1677 261 -1677 0 1
rlabel polysilicon 261 -1683 261 -1683 0 3
rlabel polysilicon 268 -1677 268 -1677 0 1
rlabel polysilicon 268 -1683 268 -1683 0 3
rlabel polysilicon 275 -1677 275 -1677 0 1
rlabel polysilicon 275 -1683 275 -1683 0 3
rlabel polysilicon 282 -1677 282 -1677 0 1
rlabel polysilicon 285 -1683 285 -1683 0 4
rlabel polysilicon 289 -1677 289 -1677 0 1
rlabel polysilicon 289 -1683 289 -1683 0 3
rlabel polysilicon 292 -1683 292 -1683 0 4
rlabel polysilicon 296 -1677 296 -1677 0 1
rlabel polysilicon 299 -1677 299 -1677 0 2
rlabel polysilicon 299 -1683 299 -1683 0 4
rlabel polysilicon 303 -1677 303 -1677 0 1
rlabel polysilicon 303 -1683 303 -1683 0 3
rlabel polysilicon 310 -1677 310 -1677 0 1
rlabel polysilicon 310 -1683 310 -1683 0 3
rlabel polysilicon 317 -1677 317 -1677 0 1
rlabel polysilicon 317 -1683 317 -1683 0 3
rlabel polysilicon 324 -1677 324 -1677 0 1
rlabel polysilicon 324 -1683 324 -1683 0 3
rlabel polysilicon 331 -1677 331 -1677 0 1
rlabel polysilicon 331 -1683 331 -1683 0 3
rlabel polysilicon 338 -1677 338 -1677 0 1
rlabel polysilicon 338 -1683 338 -1683 0 3
rlabel polysilicon 345 -1677 345 -1677 0 1
rlabel polysilicon 345 -1683 345 -1683 0 3
rlabel polysilicon 348 -1683 348 -1683 0 4
rlabel polysilicon 352 -1677 352 -1677 0 1
rlabel polysilicon 352 -1683 352 -1683 0 3
rlabel polysilicon 359 -1677 359 -1677 0 1
rlabel polysilicon 359 -1683 359 -1683 0 3
rlabel polysilicon 366 -1677 366 -1677 0 1
rlabel polysilicon 366 -1683 366 -1683 0 3
rlabel polysilicon 369 -1683 369 -1683 0 4
rlabel polysilicon 373 -1677 373 -1677 0 1
rlabel polysilicon 373 -1683 373 -1683 0 3
rlabel polysilicon 380 -1683 380 -1683 0 3
rlabel polysilicon 383 -1683 383 -1683 0 4
rlabel polysilicon 387 -1677 387 -1677 0 1
rlabel polysilicon 390 -1677 390 -1677 0 2
rlabel polysilicon 394 -1677 394 -1677 0 1
rlabel polysilicon 394 -1683 394 -1683 0 3
rlabel polysilicon 401 -1677 401 -1677 0 1
rlabel polysilicon 401 -1683 401 -1683 0 3
rlabel polysilicon 408 -1677 408 -1677 0 1
rlabel polysilicon 408 -1683 408 -1683 0 3
rlabel polysilicon 415 -1677 415 -1677 0 1
rlabel polysilicon 415 -1683 415 -1683 0 3
rlabel polysilicon 422 -1677 422 -1677 0 1
rlabel polysilicon 422 -1683 422 -1683 0 3
rlabel polysilicon 429 -1677 429 -1677 0 1
rlabel polysilicon 429 -1683 429 -1683 0 3
rlabel polysilicon 436 -1677 436 -1677 0 1
rlabel polysilicon 436 -1683 436 -1683 0 3
rlabel polysilicon 443 -1677 443 -1677 0 1
rlabel polysilicon 443 -1683 443 -1683 0 3
rlabel polysilicon 450 -1677 450 -1677 0 1
rlabel polysilicon 453 -1677 453 -1677 0 2
rlabel polysilicon 450 -1683 450 -1683 0 3
rlabel polysilicon 453 -1683 453 -1683 0 4
rlabel polysilicon 457 -1677 457 -1677 0 1
rlabel polysilicon 457 -1683 457 -1683 0 3
rlabel polysilicon 464 -1677 464 -1677 0 1
rlabel polysilicon 467 -1677 467 -1677 0 2
rlabel polysilicon 464 -1683 464 -1683 0 3
rlabel polysilicon 467 -1683 467 -1683 0 4
rlabel polysilicon 474 -1677 474 -1677 0 2
rlabel polysilicon 471 -1683 471 -1683 0 3
rlabel polysilicon 474 -1683 474 -1683 0 4
rlabel polysilicon 478 -1677 478 -1677 0 1
rlabel polysilicon 481 -1677 481 -1677 0 2
rlabel polysilicon 478 -1683 478 -1683 0 3
rlabel polysilicon 481 -1683 481 -1683 0 4
rlabel polysilicon 488 -1677 488 -1677 0 2
rlabel polysilicon 485 -1683 485 -1683 0 3
rlabel polysilicon 488 -1683 488 -1683 0 4
rlabel polysilicon 492 -1677 492 -1677 0 1
rlabel polysilicon 492 -1683 492 -1683 0 3
rlabel polysilicon 495 -1683 495 -1683 0 4
rlabel polysilicon 499 -1677 499 -1677 0 1
rlabel polysilicon 499 -1683 499 -1683 0 3
rlabel polysilicon 506 -1677 506 -1677 0 1
rlabel polysilicon 506 -1683 506 -1683 0 3
rlabel polysilicon 513 -1677 513 -1677 0 1
rlabel polysilicon 513 -1683 513 -1683 0 3
rlabel polysilicon 520 -1677 520 -1677 0 1
rlabel polysilicon 520 -1683 520 -1683 0 3
rlabel polysilicon 527 -1677 527 -1677 0 1
rlabel polysilicon 527 -1683 527 -1683 0 3
rlabel polysilicon 534 -1677 534 -1677 0 1
rlabel polysilicon 537 -1677 537 -1677 0 2
rlabel polysilicon 541 -1677 541 -1677 0 1
rlabel polysilicon 541 -1683 541 -1683 0 3
rlabel polysilicon 548 -1677 548 -1677 0 1
rlabel polysilicon 548 -1683 548 -1683 0 3
rlabel polysilicon 551 -1683 551 -1683 0 4
rlabel polysilicon 555 -1677 555 -1677 0 1
rlabel polysilicon 558 -1677 558 -1677 0 2
rlabel polysilicon 558 -1683 558 -1683 0 4
rlabel polysilicon 565 -1677 565 -1677 0 2
rlabel polysilicon 562 -1683 562 -1683 0 3
rlabel polysilicon 565 -1683 565 -1683 0 4
rlabel polysilicon 569 -1677 569 -1677 0 1
rlabel polysilicon 569 -1683 569 -1683 0 3
rlabel polysilicon 576 -1677 576 -1677 0 1
rlabel polysilicon 576 -1683 576 -1683 0 3
rlabel polysilicon 583 -1677 583 -1677 0 1
rlabel polysilicon 583 -1683 583 -1683 0 3
rlabel polysilicon 590 -1677 590 -1677 0 1
rlabel polysilicon 590 -1683 590 -1683 0 3
rlabel polysilicon 597 -1677 597 -1677 0 1
rlabel polysilicon 597 -1683 597 -1683 0 3
rlabel polysilicon 604 -1677 604 -1677 0 1
rlabel polysilicon 604 -1683 604 -1683 0 3
rlabel polysilicon 611 -1677 611 -1677 0 1
rlabel polysilicon 611 -1683 611 -1683 0 3
rlabel polysilicon 618 -1677 618 -1677 0 1
rlabel polysilicon 618 -1683 618 -1683 0 3
rlabel polysilicon 625 -1677 625 -1677 0 1
rlabel polysilicon 625 -1683 625 -1683 0 3
rlabel polysilicon 632 -1677 632 -1677 0 1
rlabel polysilicon 632 -1683 632 -1683 0 3
rlabel polysilicon 639 -1677 639 -1677 0 1
rlabel polysilicon 639 -1683 639 -1683 0 3
rlabel polysilicon 646 -1677 646 -1677 0 1
rlabel polysilicon 646 -1683 646 -1683 0 3
rlabel polysilicon 653 -1677 653 -1677 0 1
rlabel polysilicon 653 -1683 653 -1683 0 3
rlabel polysilicon 660 -1677 660 -1677 0 1
rlabel polysilicon 660 -1683 660 -1683 0 3
rlabel polysilicon 667 -1677 667 -1677 0 1
rlabel polysilicon 667 -1683 667 -1683 0 3
rlabel polysilicon 674 -1677 674 -1677 0 1
rlabel polysilicon 674 -1683 674 -1683 0 3
rlabel polysilicon 681 -1677 681 -1677 0 1
rlabel polysilicon 681 -1683 681 -1683 0 3
rlabel polysilicon 688 -1677 688 -1677 0 1
rlabel polysilicon 688 -1683 688 -1683 0 3
rlabel polysilicon 695 -1677 695 -1677 0 1
rlabel polysilicon 695 -1683 695 -1683 0 3
rlabel polysilicon 702 -1677 702 -1677 0 1
rlabel polysilicon 702 -1683 702 -1683 0 3
rlabel polysilicon 709 -1677 709 -1677 0 1
rlabel polysilicon 709 -1683 709 -1683 0 3
rlabel polysilicon 716 -1677 716 -1677 0 1
rlabel polysilicon 716 -1683 716 -1683 0 3
rlabel polysilicon 723 -1677 723 -1677 0 1
rlabel polysilicon 723 -1683 723 -1683 0 3
rlabel polysilicon 730 -1683 730 -1683 0 3
rlabel polysilicon 733 -1683 733 -1683 0 4
rlabel polysilicon 737 -1677 737 -1677 0 1
rlabel polysilicon 737 -1683 737 -1683 0 3
rlabel polysilicon 744 -1677 744 -1677 0 1
rlabel polysilicon 744 -1683 744 -1683 0 3
rlabel polysilicon 751 -1677 751 -1677 0 1
rlabel polysilicon 751 -1683 751 -1683 0 3
rlabel polysilicon 758 -1677 758 -1677 0 1
rlabel polysilicon 758 -1683 758 -1683 0 3
rlabel polysilicon 765 -1677 765 -1677 0 1
rlabel polysilicon 765 -1683 765 -1683 0 3
rlabel polysilicon 772 -1677 772 -1677 0 1
rlabel polysilicon 772 -1683 772 -1683 0 3
rlabel polysilicon 779 -1677 779 -1677 0 1
rlabel polysilicon 779 -1683 779 -1683 0 3
rlabel polysilicon 786 -1677 786 -1677 0 1
rlabel polysilicon 786 -1683 786 -1683 0 3
rlabel polysilicon 793 -1677 793 -1677 0 1
rlabel polysilicon 793 -1683 793 -1683 0 3
rlabel polysilicon 800 -1677 800 -1677 0 1
rlabel polysilicon 800 -1683 800 -1683 0 3
rlabel polysilicon 807 -1677 807 -1677 0 1
rlabel polysilicon 807 -1683 807 -1683 0 3
rlabel polysilicon 814 -1677 814 -1677 0 1
rlabel polysilicon 814 -1683 814 -1683 0 3
rlabel polysilicon 821 -1677 821 -1677 0 1
rlabel polysilicon 824 -1677 824 -1677 0 2
rlabel polysilicon 821 -1683 821 -1683 0 3
rlabel polysilicon 828 -1677 828 -1677 0 1
rlabel polysilicon 828 -1683 828 -1683 0 3
rlabel polysilicon 835 -1677 835 -1677 0 1
rlabel polysilicon 835 -1683 835 -1683 0 3
rlabel polysilicon 842 -1677 842 -1677 0 1
rlabel polysilicon 842 -1683 842 -1683 0 3
rlabel polysilicon 849 -1677 849 -1677 0 1
rlabel polysilicon 849 -1683 849 -1683 0 3
rlabel polysilicon 856 -1677 856 -1677 0 1
rlabel polysilicon 856 -1683 856 -1683 0 3
rlabel polysilicon 863 -1677 863 -1677 0 1
rlabel polysilicon 863 -1683 863 -1683 0 3
rlabel polysilicon 870 -1677 870 -1677 0 1
rlabel polysilicon 870 -1683 870 -1683 0 3
rlabel polysilicon 877 -1677 877 -1677 0 1
rlabel polysilicon 877 -1683 877 -1683 0 3
rlabel polysilicon 887 -1677 887 -1677 0 2
rlabel polysilicon 884 -1683 884 -1683 0 3
rlabel polysilicon 887 -1683 887 -1683 0 4
rlabel polysilicon 891 -1677 891 -1677 0 1
rlabel polysilicon 894 -1677 894 -1677 0 2
rlabel polysilicon 891 -1683 891 -1683 0 3
rlabel polysilicon 894 -1683 894 -1683 0 4
rlabel polysilicon 898 -1677 898 -1677 0 1
rlabel polysilicon 898 -1683 898 -1683 0 3
rlabel polysilicon 905 -1677 905 -1677 0 1
rlabel polysilicon 905 -1683 905 -1683 0 3
rlabel polysilicon 915 -1677 915 -1677 0 2
rlabel polysilicon 912 -1683 912 -1683 0 3
rlabel polysilicon 919 -1677 919 -1677 0 1
rlabel polysilicon 919 -1683 919 -1683 0 3
rlabel polysilicon 926 -1677 926 -1677 0 1
rlabel polysilicon 926 -1683 926 -1683 0 3
rlabel polysilicon 933 -1677 933 -1677 0 1
rlabel polysilicon 933 -1683 933 -1683 0 3
rlabel polysilicon 940 -1677 940 -1677 0 1
rlabel polysilicon 940 -1683 940 -1683 0 3
rlabel polysilicon 947 -1677 947 -1677 0 1
rlabel polysilicon 947 -1683 947 -1683 0 3
rlabel polysilicon 954 -1677 954 -1677 0 1
rlabel polysilicon 954 -1683 954 -1683 0 3
rlabel polysilicon 961 -1677 961 -1677 0 1
rlabel polysilicon 961 -1683 961 -1683 0 3
rlabel polysilicon 975 -1677 975 -1677 0 1
rlabel polysilicon 975 -1683 975 -1683 0 3
rlabel polysilicon 982 -1677 982 -1677 0 1
rlabel polysilicon 982 -1683 982 -1683 0 3
rlabel polysilicon 1003 -1677 1003 -1677 0 1
rlabel polysilicon 1003 -1683 1003 -1683 0 3
rlabel polysilicon 1024 -1683 1024 -1683 0 3
rlabel polysilicon 1027 -1683 1027 -1683 0 4
rlabel polysilicon 1052 -1677 1052 -1677 0 1
rlabel polysilicon 1052 -1683 1052 -1683 0 3
rlabel polysilicon 2 -1772 2 -1772 0 1
rlabel polysilicon 2 -1778 2 -1778 0 3
rlabel polysilicon 9 -1778 9 -1778 0 3
rlabel polysilicon 16 -1772 16 -1772 0 1
rlabel polysilicon 23 -1772 23 -1772 0 1
rlabel polysilicon 23 -1778 23 -1778 0 3
rlabel polysilicon 30 -1772 30 -1772 0 1
rlabel polysilicon 30 -1778 30 -1778 0 3
rlabel polysilicon 37 -1772 37 -1772 0 1
rlabel polysilicon 37 -1778 37 -1778 0 3
rlabel polysilicon 44 -1772 44 -1772 0 1
rlabel polysilicon 44 -1778 44 -1778 0 3
rlabel polysilicon 51 -1772 51 -1772 0 1
rlabel polysilicon 54 -1772 54 -1772 0 2
rlabel polysilicon 51 -1778 51 -1778 0 3
rlabel polysilicon 54 -1778 54 -1778 0 4
rlabel polysilicon 61 -1772 61 -1772 0 2
rlabel polysilicon 65 -1772 65 -1772 0 1
rlabel polysilicon 65 -1778 65 -1778 0 3
rlabel polysilicon 72 -1772 72 -1772 0 1
rlabel polysilicon 72 -1778 72 -1778 0 3
rlabel polysilicon 79 -1772 79 -1772 0 1
rlabel polysilicon 79 -1778 79 -1778 0 3
rlabel polysilicon 86 -1772 86 -1772 0 1
rlabel polysilicon 86 -1778 86 -1778 0 3
rlabel polysilicon 93 -1772 93 -1772 0 1
rlabel polysilicon 93 -1778 93 -1778 0 3
rlabel polysilicon 100 -1772 100 -1772 0 1
rlabel polysilicon 103 -1772 103 -1772 0 2
rlabel polysilicon 100 -1778 100 -1778 0 3
rlabel polysilicon 103 -1778 103 -1778 0 4
rlabel polysilicon 107 -1772 107 -1772 0 1
rlabel polysilicon 110 -1772 110 -1772 0 2
rlabel polysilicon 110 -1778 110 -1778 0 4
rlabel polysilicon 114 -1772 114 -1772 0 1
rlabel polysilicon 114 -1778 114 -1778 0 3
rlabel polysilicon 121 -1772 121 -1772 0 1
rlabel polysilicon 121 -1778 121 -1778 0 3
rlabel polysilicon 128 -1772 128 -1772 0 1
rlabel polysilicon 128 -1778 128 -1778 0 3
rlabel polysilicon 135 -1772 135 -1772 0 1
rlabel polysilicon 135 -1778 135 -1778 0 3
rlabel polysilicon 142 -1772 142 -1772 0 1
rlabel polysilicon 142 -1778 142 -1778 0 3
rlabel polysilicon 149 -1772 149 -1772 0 1
rlabel polysilicon 149 -1778 149 -1778 0 3
rlabel polysilicon 156 -1772 156 -1772 0 1
rlabel polysilicon 156 -1778 156 -1778 0 3
rlabel polysilicon 163 -1772 163 -1772 0 1
rlabel polysilicon 166 -1772 166 -1772 0 2
rlabel polysilicon 170 -1772 170 -1772 0 1
rlabel polysilicon 170 -1778 170 -1778 0 3
rlabel polysilicon 177 -1772 177 -1772 0 1
rlabel polysilicon 180 -1772 180 -1772 0 2
rlabel polysilicon 177 -1778 177 -1778 0 3
rlabel polysilicon 187 -1772 187 -1772 0 2
rlabel polysilicon 187 -1778 187 -1778 0 4
rlabel polysilicon 191 -1772 191 -1772 0 1
rlabel polysilicon 191 -1778 191 -1778 0 3
rlabel polysilicon 198 -1772 198 -1772 0 1
rlabel polysilicon 198 -1778 198 -1778 0 3
rlabel polysilicon 205 -1772 205 -1772 0 1
rlabel polysilicon 205 -1778 205 -1778 0 3
rlabel polysilicon 215 -1778 215 -1778 0 4
rlabel polysilicon 222 -1772 222 -1772 0 2
rlabel polysilicon 219 -1778 219 -1778 0 3
rlabel polysilicon 226 -1772 226 -1772 0 1
rlabel polysilicon 226 -1778 226 -1778 0 3
rlabel polysilicon 233 -1772 233 -1772 0 1
rlabel polysilicon 233 -1778 233 -1778 0 3
rlabel polysilicon 240 -1772 240 -1772 0 1
rlabel polysilicon 243 -1772 243 -1772 0 2
rlabel polysilicon 240 -1778 240 -1778 0 3
rlabel polysilicon 243 -1778 243 -1778 0 4
rlabel polysilicon 247 -1772 247 -1772 0 1
rlabel polysilicon 247 -1778 247 -1778 0 3
rlabel polysilicon 254 -1772 254 -1772 0 1
rlabel polysilicon 254 -1778 254 -1778 0 3
rlabel polysilicon 261 -1772 261 -1772 0 1
rlabel polysilicon 261 -1778 261 -1778 0 3
rlabel polysilicon 268 -1772 268 -1772 0 1
rlabel polysilicon 268 -1778 268 -1778 0 3
rlabel polysilicon 275 -1772 275 -1772 0 1
rlabel polysilicon 275 -1778 275 -1778 0 3
rlabel polysilicon 282 -1772 282 -1772 0 1
rlabel polysilicon 282 -1778 282 -1778 0 3
rlabel polysilicon 289 -1772 289 -1772 0 1
rlabel polysilicon 289 -1778 289 -1778 0 3
rlabel polysilicon 296 -1772 296 -1772 0 1
rlabel polysilicon 296 -1778 296 -1778 0 3
rlabel polysilicon 303 -1772 303 -1772 0 1
rlabel polysilicon 303 -1778 303 -1778 0 3
rlabel polysilicon 313 -1772 313 -1772 0 2
rlabel polysilicon 310 -1778 310 -1778 0 3
rlabel polysilicon 313 -1778 313 -1778 0 4
rlabel polysilicon 317 -1772 317 -1772 0 1
rlabel polysilicon 317 -1778 317 -1778 0 3
rlabel polysilicon 324 -1772 324 -1772 0 1
rlabel polysilicon 324 -1778 324 -1778 0 3
rlabel polysilicon 327 -1778 327 -1778 0 4
rlabel polysilicon 331 -1772 331 -1772 0 1
rlabel polysilicon 331 -1778 331 -1778 0 3
rlabel polysilicon 338 -1772 338 -1772 0 1
rlabel polysilicon 338 -1778 338 -1778 0 3
rlabel polysilicon 345 -1772 345 -1772 0 1
rlabel polysilicon 345 -1778 345 -1778 0 3
rlabel polysilicon 352 -1772 352 -1772 0 1
rlabel polysilicon 352 -1778 352 -1778 0 3
rlabel polysilicon 359 -1772 359 -1772 0 1
rlabel polysilicon 359 -1778 359 -1778 0 3
rlabel polysilicon 366 -1772 366 -1772 0 1
rlabel polysilicon 369 -1772 369 -1772 0 2
rlabel polysilicon 366 -1778 366 -1778 0 3
rlabel polysilicon 369 -1778 369 -1778 0 4
rlabel polysilicon 373 -1772 373 -1772 0 1
rlabel polysilicon 376 -1772 376 -1772 0 2
rlabel polysilicon 373 -1778 373 -1778 0 3
rlabel polysilicon 376 -1778 376 -1778 0 4
rlabel polysilicon 383 -1772 383 -1772 0 2
rlabel polysilicon 380 -1778 380 -1778 0 3
rlabel polysilicon 387 -1772 387 -1772 0 1
rlabel polysilicon 387 -1778 387 -1778 0 3
rlabel polysilicon 394 -1772 394 -1772 0 1
rlabel polysilicon 394 -1778 394 -1778 0 3
rlabel polysilicon 401 -1772 401 -1772 0 1
rlabel polysilicon 404 -1772 404 -1772 0 2
rlabel polysilicon 401 -1778 401 -1778 0 3
rlabel polysilicon 408 -1772 408 -1772 0 1
rlabel polysilicon 411 -1772 411 -1772 0 2
rlabel polysilicon 408 -1778 408 -1778 0 3
rlabel polysilicon 415 -1772 415 -1772 0 1
rlabel polysilicon 415 -1778 415 -1778 0 3
rlabel polysilicon 422 -1772 422 -1772 0 1
rlabel polysilicon 425 -1772 425 -1772 0 2
rlabel polysilicon 429 -1772 429 -1772 0 1
rlabel polysilicon 429 -1778 429 -1778 0 3
rlabel polysilicon 436 -1772 436 -1772 0 1
rlabel polysilicon 436 -1778 436 -1778 0 3
rlabel polysilicon 443 -1772 443 -1772 0 1
rlabel polysilicon 443 -1778 443 -1778 0 3
rlabel polysilicon 450 -1772 450 -1772 0 1
rlabel polysilicon 450 -1778 450 -1778 0 3
rlabel polysilicon 457 -1772 457 -1772 0 1
rlabel polysilicon 457 -1778 457 -1778 0 3
rlabel polysilicon 464 -1772 464 -1772 0 1
rlabel polysilicon 467 -1772 467 -1772 0 2
rlabel polysilicon 464 -1778 464 -1778 0 3
rlabel polysilicon 467 -1778 467 -1778 0 4
rlabel polysilicon 471 -1772 471 -1772 0 1
rlabel polysilicon 471 -1778 471 -1778 0 3
rlabel polysilicon 478 -1772 478 -1772 0 1
rlabel polysilicon 481 -1772 481 -1772 0 2
rlabel polysilicon 485 -1772 485 -1772 0 1
rlabel polysilicon 485 -1778 485 -1778 0 3
rlabel polysilicon 492 -1772 492 -1772 0 1
rlabel polysilicon 492 -1778 492 -1778 0 3
rlabel polysilicon 499 -1772 499 -1772 0 1
rlabel polysilicon 499 -1778 499 -1778 0 3
rlabel polysilicon 506 -1772 506 -1772 0 1
rlabel polysilicon 506 -1778 506 -1778 0 3
rlabel polysilicon 513 -1772 513 -1772 0 1
rlabel polysilicon 516 -1772 516 -1772 0 2
rlabel polysilicon 516 -1778 516 -1778 0 4
rlabel polysilicon 520 -1772 520 -1772 0 1
rlabel polysilicon 520 -1778 520 -1778 0 3
rlabel polysilicon 527 -1772 527 -1772 0 1
rlabel polysilicon 527 -1778 527 -1778 0 3
rlabel polysilicon 534 -1772 534 -1772 0 1
rlabel polysilicon 534 -1778 534 -1778 0 3
rlabel polysilicon 541 -1772 541 -1772 0 1
rlabel polysilicon 541 -1778 541 -1778 0 3
rlabel polysilicon 548 -1772 548 -1772 0 1
rlabel polysilicon 548 -1778 548 -1778 0 3
rlabel polysilicon 555 -1772 555 -1772 0 1
rlabel polysilicon 555 -1778 555 -1778 0 3
rlabel polysilicon 562 -1772 562 -1772 0 1
rlabel polysilicon 562 -1778 562 -1778 0 3
rlabel polysilicon 569 -1772 569 -1772 0 1
rlabel polysilicon 569 -1778 569 -1778 0 3
rlabel polysilicon 576 -1772 576 -1772 0 1
rlabel polysilicon 576 -1778 576 -1778 0 3
rlabel polysilicon 583 -1772 583 -1772 0 1
rlabel polysilicon 583 -1778 583 -1778 0 3
rlabel polysilicon 593 -1772 593 -1772 0 2
rlabel polysilicon 590 -1778 590 -1778 0 3
rlabel polysilicon 593 -1778 593 -1778 0 4
rlabel polysilicon 597 -1772 597 -1772 0 1
rlabel polysilicon 597 -1778 597 -1778 0 3
rlabel polysilicon 604 -1772 604 -1772 0 1
rlabel polysilicon 604 -1778 604 -1778 0 3
rlabel polysilicon 614 -1772 614 -1772 0 2
rlabel polysilicon 611 -1778 611 -1778 0 3
rlabel polysilicon 618 -1772 618 -1772 0 1
rlabel polysilicon 621 -1772 621 -1772 0 2
rlabel polysilicon 618 -1778 618 -1778 0 3
rlabel polysilicon 621 -1778 621 -1778 0 4
rlabel polysilicon 625 -1772 625 -1772 0 1
rlabel polysilicon 625 -1778 625 -1778 0 3
rlabel polysilicon 632 -1778 632 -1778 0 3
rlabel polysilicon 635 -1778 635 -1778 0 4
rlabel polysilicon 639 -1772 639 -1772 0 1
rlabel polysilicon 639 -1778 639 -1778 0 3
rlabel polysilicon 646 -1772 646 -1772 0 1
rlabel polysilicon 649 -1772 649 -1772 0 2
rlabel polysilicon 646 -1778 646 -1778 0 3
rlabel polysilicon 653 -1772 653 -1772 0 1
rlabel polysilicon 653 -1778 653 -1778 0 3
rlabel polysilicon 656 -1778 656 -1778 0 4
rlabel polysilicon 660 -1772 660 -1772 0 1
rlabel polysilicon 660 -1778 660 -1778 0 3
rlabel polysilicon 667 -1772 667 -1772 0 1
rlabel polysilicon 667 -1778 667 -1778 0 3
rlabel polysilicon 674 -1772 674 -1772 0 1
rlabel polysilicon 677 -1772 677 -1772 0 2
rlabel polysilicon 674 -1778 674 -1778 0 3
rlabel polysilicon 677 -1778 677 -1778 0 4
rlabel polysilicon 681 -1772 681 -1772 0 1
rlabel polysilicon 681 -1778 681 -1778 0 3
rlabel polysilicon 688 -1772 688 -1772 0 1
rlabel polysilicon 688 -1778 688 -1778 0 3
rlabel polysilicon 695 -1772 695 -1772 0 1
rlabel polysilicon 695 -1778 695 -1778 0 3
rlabel polysilicon 702 -1772 702 -1772 0 1
rlabel polysilicon 702 -1778 702 -1778 0 3
rlabel polysilicon 709 -1772 709 -1772 0 1
rlabel polysilicon 709 -1778 709 -1778 0 3
rlabel polysilicon 716 -1772 716 -1772 0 1
rlabel polysilicon 716 -1778 716 -1778 0 3
rlabel polysilicon 723 -1772 723 -1772 0 1
rlabel polysilicon 723 -1778 723 -1778 0 3
rlabel polysilicon 730 -1772 730 -1772 0 1
rlabel polysilicon 730 -1778 730 -1778 0 3
rlabel polysilicon 737 -1772 737 -1772 0 1
rlabel polysilicon 737 -1778 737 -1778 0 3
rlabel polysilicon 744 -1772 744 -1772 0 1
rlabel polysilicon 744 -1778 744 -1778 0 3
rlabel polysilicon 751 -1772 751 -1772 0 1
rlabel polysilicon 751 -1778 751 -1778 0 3
rlabel polysilicon 758 -1772 758 -1772 0 1
rlabel polysilicon 758 -1778 758 -1778 0 3
rlabel polysilicon 765 -1772 765 -1772 0 1
rlabel polysilicon 765 -1778 765 -1778 0 3
rlabel polysilicon 772 -1772 772 -1772 0 1
rlabel polysilicon 772 -1778 772 -1778 0 3
rlabel polysilicon 779 -1772 779 -1772 0 1
rlabel polysilicon 779 -1778 779 -1778 0 3
rlabel polysilicon 786 -1772 786 -1772 0 1
rlabel polysilicon 786 -1778 786 -1778 0 3
rlabel polysilicon 793 -1772 793 -1772 0 1
rlabel polysilicon 793 -1778 793 -1778 0 3
rlabel polysilicon 803 -1772 803 -1772 0 2
rlabel polysilicon 807 -1772 807 -1772 0 1
rlabel polysilicon 807 -1778 807 -1778 0 3
rlabel polysilicon 814 -1772 814 -1772 0 1
rlabel polysilicon 814 -1778 814 -1778 0 3
rlabel polysilicon 821 -1772 821 -1772 0 1
rlabel polysilicon 821 -1778 821 -1778 0 3
rlabel polysilicon 828 -1772 828 -1772 0 1
rlabel polysilicon 828 -1778 828 -1778 0 3
rlabel polysilicon 835 -1772 835 -1772 0 1
rlabel polysilicon 835 -1778 835 -1778 0 3
rlabel polysilicon 842 -1772 842 -1772 0 1
rlabel polysilicon 842 -1778 842 -1778 0 3
rlabel polysilicon 849 -1772 849 -1772 0 1
rlabel polysilicon 849 -1778 849 -1778 0 3
rlabel polysilicon 856 -1772 856 -1772 0 1
rlabel polysilicon 856 -1778 856 -1778 0 3
rlabel polysilicon 863 -1772 863 -1772 0 1
rlabel polysilicon 863 -1778 863 -1778 0 3
rlabel polysilicon 870 -1772 870 -1772 0 1
rlabel polysilicon 870 -1778 870 -1778 0 3
rlabel polysilicon 877 -1772 877 -1772 0 1
rlabel polysilicon 877 -1778 877 -1778 0 3
rlabel polysilicon 884 -1772 884 -1772 0 1
rlabel polysilicon 884 -1778 884 -1778 0 3
rlabel polysilicon 891 -1772 891 -1772 0 1
rlabel polysilicon 891 -1778 891 -1778 0 3
rlabel polysilicon 898 -1772 898 -1772 0 1
rlabel polysilicon 898 -1778 898 -1778 0 3
rlabel polysilicon 905 -1772 905 -1772 0 1
rlabel polysilicon 905 -1778 905 -1778 0 3
rlabel polysilicon 912 -1772 912 -1772 0 1
rlabel polysilicon 912 -1778 912 -1778 0 3
rlabel polysilicon 919 -1772 919 -1772 0 1
rlabel polysilicon 919 -1778 919 -1778 0 3
rlabel polysilicon 926 -1772 926 -1772 0 1
rlabel polysilicon 926 -1778 926 -1778 0 3
rlabel polysilicon 933 -1772 933 -1772 0 1
rlabel polysilicon 933 -1778 933 -1778 0 3
rlabel polysilicon 940 -1772 940 -1772 0 1
rlabel polysilicon 940 -1778 940 -1778 0 3
rlabel polysilicon 947 -1772 947 -1772 0 1
rlabel polysilicon 947 -1778 947 -1778 0 3
rlabel polysilicon 954 -1772 954 -1772 0 1
rlabel polysilicon 954 -1778 954 -1778 0 3
rlabel polysilicon 961 -1772 961 -1772 0 1
rlabel polysilicon 961 -1778 961 -1778 0 3
rlabel polysilicon 968 -1772 968 -1772 0 1
rlabel polysilicon 968 -1778 968 -1778 0 3
rlabel polysilicon 975 -1772 975 -1772 0 1
rlabel polysilicon 975 -1778 975 -1778 0 3
rlabel polysilicon 982 -1772 982 -1772 0 1
rlabel polysilicon 982 -1778 982 -1778 0 3
rlabel polysilicon 989 -1772 989 -1772 0 1
rlabel polysilicon 989 -1778 989 -1778 0 3
rlabel polysilicon 996 -1778 996 -1778 0 3
rlabel polysilicon 999 -1778 999 -1778 0 4
rlabel polysilicon 1006 -1772 1006 -1772 0 2
rlabel polysilicon 1003 -1778 1003 -1778 0 3
rlabel polysilicon 1010 -1772 1010 -1772 0 1
rlabel polysilicon 1010 -1778 1010 -1778 0 3
rlabel polysilicon 1017 -1772 1017 -1772 0 1
rlabel polysilicon 1017 -1778 1017 -1778 0 3
rlabel polysilicon 1024 -1772 1024 -1772 0 1
rlabel polysilicon 1024 -1778 1024 -1778 0 3
rlabel polysilicon 51 -1863 51 -1863 0 1
rlabel polysilicon 51 -1869 51 -1869 0 3
rlabel polysilicon 58 -1863 58 -1863 0 1
rlabel polysilicon 58 -1869 58 -1869 0 3
rlabel polysilicon 65 -1863 65 -1863 0 1
rlabel polysilicon 65 -1869 65 -1869 0 3
rlabel polysilicon 72 -1863 72 -1863 0 1
rlabel polysilicon 72 -1869 72 -1869 0 3
rlabel polysilicon 79 -1863 79 -1863 0 1
rlabel polysilicon 79 -1869 79 -1869 0 3
rlabel polysilicon 86 -1863 86 -1863 0 1
rlabel polysilicon 86 -1869 86 -1869 0 3
rlabel polysilicon 93 -1863 93 -1863 0 1
rlabel polysilicon 93 -1869 93 -1869 0 3
rlabel polysilicon 100 -1863 100 -1863 0 1
rlabel polysilicon 100 -1869 100 -1869 0 3
rlabel polysilicon 107 -1863 107 -1863 0 1
rlabel polysilicon 107 -1869 107 -1869 0 3
rlabel polysilicon 114 -1863 114 -1863 0 1
rlabel polysilicon 114 -1869 114 -1869 0 3
rlabel polysilicon 121 -1863 121 -1863 0 1
rlabel polysilicon 121 -1869 121 -1869 0 3
rlabel polysilicon 128 -1863 128 -1863 0 1
rlabel polysilicon 131 -1869 131 -1869 0 4
rlabel polysilicon 135 -1863 135 -1863 0 1
rlabel polysilicon 135 -1869 135 -1869 0 3
rlabel polysilicon 142 -1863 142 -1863 0 1
rlabel polysilicon 142 -1869 142 -1869 0 3
rlabel polysilicon 149 -1863 149 -1863 0 1
rlabel polysilicon 149 -1869 149 -1869 0 3
rlabel polysilicon 156 -1863 156 -1863 0 1
rlabel polysilicon 156 -1869 156 -1869 0 3
rlabel polysilicon 163 -1863 163 -1863 0 1
rlabel polysilicon 163 -1869 163 -1869 0 3
rlabel polysilicon 166 -1869 166 -1869 0 4
rlabel polysilicon 170 -1863 170 -1863 0 1
rlabel polysilicon 170 -1869 170 -1869 0 3
rlabel polysilicon 177 -1863 177 -1863 0 1
rlabel polysilicon 177 -1869 177 -1869 0 3
rlabel polysilicon 184 -1863 184 -1863 0 1
rlabel polysilicon 184 -1869 184 -1869 0 3
rlabel polysilicon 194 -1863 194 -1863 0 2
rlabel polysilicon 191 -1869 191 -1869 0 3
rlabel polysilicon 201 -1863 201 -1863 0 2
rlabel polysilicon 198 -1869 198 -1869 0 3
rlabel polysilicon 205 -1869 205 -1869 0 3
rlabel polysilicon 212 -1863 212 -1863 0 1
rlabel polysilicon 215 -1863 215 -1863 0 2
rlabel polysilicon 212 -1869 212 -1869 0 3
rlabel polysilicon 215 -1869 215 -1869 0 4
rlabel polysilicon 219 -1863 219 -1863 0 1
rlabel polysilicon 219 -1869 219 -1869 0 3
rlabel polysilicon 226 -1863 226 -1863 0 1
rlabel polysilicon 229 -1863 229 -1863 0 2
rlabel polysilicon 229 -1869 229 -1869 0 4
rlabel polysilicon 233 -1863 233 -1863 0 1
rlabel polysilicon 233 -1869 233 -1869 0 3
rlabel polysilicon 240 -1869 240 -1869 0 3
rlabel polysilicon 243 -1869 243 -1869 0 4
rlabel polysilicon 247 -1863 247 -1863 0 1
rlabel polysilicon 247 -1869 247 -1869 0 3
rlabel polysilicon 254 -1863 254 -1863 0 1
rlabel polysilicon 254 -1869 254 -1869 0 3
rlabel polysilicon 261 -1863 261 -1863 0 1
rlabel polysilicon 261 -1869 261 -1869 0 3
rlabel polysilicon 268 -1863 268 -1863 0 1
rlabel polysilicon 268 -1869 268 -1869 0 3
rlabel polysilicon 275 -1863 275 -1863 0 1
rlabel polysilicon 275 -1869 275 -1869 0 3
rlabel polysilicon 282 -1863 282 -1863 0 1
rlabel polysilicon 282 -1869 282 -1869 0 3
rlabel polysilicon 289 -1863 289 -1863 0 1
rlabel polysilicon 289 -1869 289 -1869 0 3
rlabel polysilicon 296 -1863 296 -1863 0 1
rlabel polysilicon 296 -1869 296 -1869 0 3
rlabel polysilicon 303 -1863 303 -1863 0 1
rlabel polysilicon 303 -1869 303 -1869 0 3
rlabel polysilicon 310 -1863 310 -1863 0 1
rlabel polysilicon 310 -1869 310 -1869 0 3
rlabel polysilicon 317 -1863 317 -1863 0 1
rlabel polysilicon 317 -1869 317 -1869 0 3
rlabel polysilicon 324 -1863 324 -1863 0 1
rlabel polysilicon 324 -1869 324 -1869 0 3
rlabel polysilicon 331 -1863 331 -1863 0 1
rlabel polysilicon 331 -1869 331 -1869 0 3
rlabel polysilicon 338 -1863 338 -1863 0 1
rlabel polysilicon 338 -1869 338 -1869 0 3
rlabel polysilicon 345 -1863 345 -1863 0 1
rlabel polysilicon 348 -1863 348 -1863 0 2
rlabel polysilicon 345 -1869 345 -1869 0 3
rlabel polysilicon 348 -1869 348 -1869 0 4
rlabel polysilicon 352 -1863 352 -1863 0 1
rlabel polysilicon 352 -1869 352 -1869 0 3
rlabel polysilicon 362 -1869 362 -1869 0 4
rlabel polysilicon 369 -1863 369 -1863 0 2
rlabel polysilicon 373 -1863 373 -1863 0 1
rlabel polysilicon 373 -1869 373 -1869 0 3
rlabel polysilicon 380 -1863 380 -1863 0 1
rlabel polysilicon 380 -1869 380 -1869 0 3
rlabel polysilicon 387 -1863 387 -1863 0 1
rlabel polysilicon 387 -1869 387 -1869 0 3
rlabel polysilicon 394 -1863 394 -1863 0 1
rlabel polysilicon 394 -1869 394 -1869 0 3
rlabel polysilicon 401 -1863 401 -1863 0 1
rlabel polysilicon 401 -1869 401 -1869 0 3
rlabel polysilicon 408 -1863 408 -1863 0 1
rlabel polysilicon 408 -1869 408 -1869 0 3
rlabel polysilicon 411 -1869 411 -1869 0 4
rlabel polysilicon 415 -1863 415 -1863 0 1
rlabel polysilicon 418 -1863 418 -1863 0 2
rlabel polysilicon 415 -1869 415 -1869 0 3
rlabel polysilicon 418 -1869 418 -1869 0 4
rlabel polysilicon 422 -1863 422 -1863 0 1
rlabel polysilicon 425 -1863 425 -1863 0 2
rlabel polysilicon 422 -1869 422 -1869 0 3
rlabel polysilicon 429 -1863 429 -1863 0 1
rlabel polysilicon 429 -1869 429 -1869 0 3
rlabel polysilicon 436 -1863 436 -1863 0 1
rlabel polysilicon 436 -1869 436 -1869 0 3
rlabel polysilicon 443 -1863 443 -1863 0 1
rlabel polysilicon 443 -1869 443 -1869 0 3
rlabel polysilicon 450 -1863 450 -1863 0 1
rlabel polysilicon 450 -1869 450 -1869 0 3
rlabel polysilicon 457 -1863 457 -1863 0 1
rlabel polysilicon 460 -1863 460 -1863 0 2
rlabel polysilicon 457 -1869 457 -1869 0 3
rlabel polysilicon 464 -1863 464 -1863 0 1
rlabel polysilicon 464 -1869 464 -1869 0 3
rlabel polysilicon 471 -1863 471 -1863 0 1
rlabel polysilicon 471 -1869 471 -1869 0 3
rlabel polysilicon 478 -1863 478 -1863 0 1
rlabel polysilicon 478 -1869 478 -1869 0 3
rlabel polysilicon 485 -1863 485 -1863 0 1
rlabel polysilicon 485 -1869 485 -1869 0 3
rlabel polysilicon 492 -1863 492 -1863 0 1
rlabel polysilicon 492 -1869 492 -1869 0 3
rlabel polysilicon 499 -1863 499 -1863 0 1
rlabel polysilicon 499 -1869 499 -1869 0 3
rlabel polysilicon 506 -1863 506 -1863 0 1
rlabel polysilicon 506 -1869 506 -1869 0 3
rlabel polysilicon 509 -1869 509 -1869 0 4
rlabel polysilicon 513 -1863 513 -1863 0 1
rlabel polysilicon 513 -1869 513 -1869 0 3
rlabel polysilicon 520 -1863 520 -1863 0 1
rlabel polysilicon 523 -1863 523 -1863 0 2
rlabel polysilicon 523 -1869 523 -1869 0 4
rlabel polysilicon 527 -1863 527 -1863 0 1
rlabel polysilicon 530 -1869 530 -1869 0 4
rlabel polysilicon 534 -1863 534 -1863 0 1
rlabel polysilicon 534 -1869 534 -1869 0 3
rlabel polysilicon 541 -1863 541 -1863 0 1
rlabel polysilicon 541 -1869 541 -1869 0 3
rlabel polysilicon 548 -1863 548 -1863 0 1
rlabel polysilicon 551 -1863 551 -1863 0 2
rlabel polysilicon 548 -1869 548 -1869 0 3
rlabel polysilicon 551 -1869 551 -1869 0 4
rlabel polysilicon 555 -1863 555 -1863 0 1
rlabel polysilicon 555 -1869 555 -1869 0 3
rlabel polysilicon 562 -1863 562 -1863 0 1
rlabel polysilicon 565 -1863 565 -1863 0 2
rlabel polysilicon 562 -1869 562 -1869 0 3
rlabel polysilicon 569 -1863 569 -1863 0 1
rlabel polysilicon 569 -1869 569 -1869 0 3
rlabel polysilicon 576 -1863 576 -1863 0 1
rlabel polysilicon 576 -1869 576 -1869 0 3
rlabel polysilicon 583 -1863 583 -1863 0 1
rlabel polysilicon 583 -1869 583 -1869 0 3
rlabel polysilicon 590 -1863 590 -1863 0 1
rlabel polysilicon 590 -1869 590 -1869 0 3
rlabel polysilicon 597 -1863 597 -1863 0 1
rlabel polysilicon 597 -1869 597 -1869 0 3
rlabel polysilicon 604 -1863 604 -1863 0 1
rlabel polysilicon 604 -1869 604 -1869 0 3
rlabel polysilicon 611 -1863 611 -1863 0 1
rlabel polysilicon 611 -1869 611 -1869 0 3
rlabel polysilicon 618 -1863 618 -1863 0 1
rlabel polysilicon 618 -1869 618 -1869 0 3
rlabel polysilicon 628 -1863 628 -1863 0 2
rlabel polysilicon 625 -1869 625 -1869 0 3
rlabel polysilicon 628 -1869 628 -1869 0 4
rlabel polysilicon 632 -1869 632 -1869 0 3
rlabel polysilicon 642 -1863 642 -1863 0 2
rlabel polysilicon 642 -1869 642 -1869 0 4
rlabel polysilicon 646 -1863 646 -1863 0 1
rlabel polysilicon 646 -1869 646 -1869 0 3
rlabel polysilicon 653 -1863 653 -1863 0 1
rlabel polysilicon 653 -1869 653 -1869 0 3
rlabel polysilicon 660 -1863 660 -1863 0 1
rlabel polysilicon 660 -1869 660 -1869 0 3
rlabel polysilicon 663 -1869 663 -1869 0 4
rlabel polysilicon 667 -1863 667 -1863 0 1
rlabel polysilicon 667 -1869 667 -1869 0 3
rlabel polysilicon 674 -1863 674 -1863 0 1
rlabel polysilicon 674 -1869 674 -1869 0 3
rlabel polysilicon 681 -1863 681 -1863 0 1
rlabel polysilicon 681 -1869 681 -1869 0 3
rlabel polysilicon 688 -1863 688 -1863 0 1
rlabel polysilicon 688 -1869 688 -1869 0 3
rlabel polysilicon 695 -1863 695 -1863 0 1
rlabel polysilicon 695 -1869 695 -1869 0 3
rlabel polysilicon 702 -1863 702 -1863 0 1
rlabel polysilicon 702 -1869 702 -1869 0 3
rlabel polysilicon 709 -1863 709 -1863 0 1
rlabel polysilicon 709 -1869 709 -1869 0 3
rlabel polysilicon 716 -1863 716 -1863 0 1
rlabel polysilicon 716 -1869 716 -1869 0 3
rlabel polysilicon 726 -1863 726 -1863 0 2
rlabel polysilicon 723 -1869 723 -1869 0 3
rlabel polysilicon 726 -1869 726 -1869 0 4
rlabel polysilicon 730 -1863 730 -1863 0 1
rlabel polysilicon 730 -1869 730 -1869 0 3
rlabel polysilicon 737 -1863 737 -1863 0 1
rlabel polysilicon 737 -1869 737 -1869 0 3
rlabel polysilicon 744 -1863 744 -1863 0 1
rlabel polysilicon 744 -1869 744 -1869 0 3
rlabel polysilicon 751 -1863 751 -1863 0 1
rlabel polysilicon 751 -1869 751 -1869 0 3
rlabel polysilicon 758 -1863 758 -1863 0 1
rlabel polysilicon 758 -1869 758 -1869 0 3
rlabel polysilicon 765 -1863 765 -1863 0 1
rlabel polysilicon 765 -1869 765 -1869 0 3
rlabel polysilicon 772 -1863 772 -1863 0 1
rlabel polysilicon 772 -1869 772 -1869 0 3
rlabel polysilicon 779 -1863 779 -1863 0 1
rlabel polysilicon 779 -1869 779 -1869 0 3
rlabel polysilicon 786 -1863 786 -1863 0 1
rlabel polysilicon 786 -1869 786 -1869 0 3
rlabel polysilicon 793 -1863 793 -1863 0 1
rlabel polysilicon 793 -1869 793 -1869 0 3
rlabel polysilicon 800 -1863 800 -1863 0 1
rlabel polysilicon 800 -1869 800 -1869 0 3
rlabel polysilicon 807 -1863 807 -1863 0 1
rlabel polysilicon 807 -1869 807 -1869 0 3
rlabel polysilicon 814 -1863 814 -1863 0 1
rlabel polysilicon 814 -1869 814 -1869 0 3
rlabel polysilicon 817 -1869 817 -1869 0 4
rlabel polysilicon 821 -1863 821 -1863 0 1
rlabel polysilicon 821 -1869 821 -1869 0 3
rlabel polysilicon 828 -1863 828 -1863 0 1
rlabel polysilicon 828 -1869 828 -1869 0 3
rlabel polysilicon 835 -1863 835 -1863 0 1
rlabel polysilicon 838 -1863 838 -1863 0 2
rlabel polysilicon 842 -1863 842 -1863 0 1
rlabel polysilicon 845 -1863 845 -1863 0 2
rlabel polysilicon 845 -1869 845 -1869 0 4
rlabel polysilicon 849 -1863 849 -1863 0 1
rlabel polysilicon 852 -1863 852 -1863 0 2
rlabel polysilicon 856 -1863 856 -1863 0 1
rlabel polysilicon 856 -1869 856 -1869 0 3
rlabel polysilicon 863 -1863 863 -1863 0 1
rlabel polysilicon 863 -1869 863 -1869 0 3
rlabel polysilicon 870 -1863 870 -1863 0 1
rlabel polysilicon 870 -1869 870 -1869 0 3
rlabel polysilicon 877 -1863 877 -1863 0 1
rlabel polysilicon 877 -1869 877 -1869 0 3
rlabel polysilicon 898 -1863 898 -1863 0 1
rlabel polysilicon 898 -1869 898 -1869 0 3
rlabel polysilicon 915 -1863 915 -1863 0 2
rlabel polysilicon 947 -1863 947 -1863 0 1
rlabel polysilicon 950 -1863 950 -1863 0 2
rlabel polysilicon 16 -1934 16 -1934 0 1
rlabel polysilicon 16 -1940 16 -1940 0 3
rlabel polysilicon 23 -1934 23 -1934 0 1
rlabel polysilicon 23 -1940 23 -1940 0 3
rlabel polysilicon 33 -1940 33 -1940 0 4
rlabel polysilicon 37 -1940 37 -1940 0 3
rlabel polysilicon 40 -1940 40 -1940 0 4
rlabel polysilicon 44 -1934 44 -1934 0 1
rlabel polysilicon 47 -1940 47 -1940 0 4
rlabel polysilicon 51 -1934 51 -1934 0 1
rlabel polysilicon 51 -1940 51 -1940 0 3
rlabel polysilicon 58 -1934 58 -1934 0 1
rlabel polysilicon 58 -1940 58 -1940 0 3
rlabel polysilicon 65 -1934 65 -1934 0 1
rlabel polysilicon 65 -1940 65 -1940 0 3
rlabel polysilicon 72 -1934 72 -1934 0 1
rlabel polysilicon 72 -1940 72 -1940 0 3
rlabel polysilicon 79 -1934 79 -1934 0 1
rlabel polysilicon 79 -1940 79 -1940 0 3
rlabel polysilicon 86 -1934 86 -1934 0 1
rlabel polysilicon 86 -1940 86 -1940 0 3
rlabel polysilicon 93 -1934 93 -1934 0 1
rlabel polysilicon 93 -1940 93 -1940 0 3
rlabel polysilicon 100 -1934 100 -1934 0 1
rlabel polysilicon 100 -1940 100 -1940 0 3
rlabel polysilicon 107 -1934 107 -1934 0 1
rlabel polysilicon 107 -1940 107 -1940 0 3
rlabel polysilicon 114 -1934 114 -1934 0 1
rlabel polysilicon 114 -1940 114 -1940 0 3
rlabel polysilicon 121 -1934 121 -1934 0 1
rlabel polysilicon 124 -1934 124 -1934 0 2
rlabel polysilicon 128 -1934 128 -1934 0 1
rlabel polysilicon 128 -1940 128 -1940 0 3
rlabel polysilicon 135 -1934 135 -1934 0 1
rlabel polysilicon 135 -1940 135 -1940 0 3
rlabel polysilicon 142 -1934 142 -1934 0 1
rlabel polysilicon 145 -1934 145 -1934 0 2
rlabel polysilicon 142 -1940 142 -1940 0 3
rlabel polysilicon 149 -1934 149 -1934 0 1
rlabel polysilicon 149 -1940 149 -1940 0 3
rlabel polysilicon 156 -1934 156 -1934 0 1
rlabel polysilicon 159 -1934 159 -1934 0 2
rlabel polysilicon 159 -1940 159 -1940 0 4
rlabel polysilicon 163 -1934 163 -1934 0 1
rlabel polysilicon 163 -1940 163 -1940 0 3
rlabel polysilicon 170 -1934 170 -1934 0 1
rlabel polysilicon 170 -1940 170 -1940 0 3
rlabel polysilicon 177 -1934 177 -1934 0 1
rlabel polysilicon 177 -1940 177 -1940 0 3
rlabel polysilicon 180 -1940 180 -1940 0 4
rlabel polysilicon 184 -1934 184 -1934 0 1
rlabel polysilicon 184 -1940 184 -1940 0 3
rlabel polysilicon 191 -1934 191 -1934 0 1
rlabel polysilicon 194 -1934 194 -1934 0 2
rlabel polysilicon 191 -1940 191 -1940 0 3
rlabel polysilicon 194 -1940 194 -1940 0 4
rlabel polysilicon 198 -1934 198 -1934 0 1
rlabel polysilicon 198 -1940 198 -1940 0 3
rlabel polysilicon 205 -1934 205 -1934 0 1
rlabel polysilicon 205 -1940 205 -1940 0 3
rlabel polysilicon 212 -1934 212 -1934 0 1
rlabel polysilicon 212 -1940 212 -1940 0 3
rlabel polysilicon 219 -1940 219 -1940 0 3
rlabel polysilicon 222 -1940 222 -1940 0 4
rlabel polysilicon 229 -1934 229 -1934 0 2
rlabel polysilicon 226 -1940 226 -1940 0 3
rlabel polysilicon 229 -1940 229 -1940 0 4
rlabel polysilicon 233 -1940 233 -1940 0 3
rlabel polysilicon 236 -1940 236 -1940 0 4
rlabel polysilicon 240 -1934 240 -1934 0 1
rlabel polysilicon 243 -1934 243 -1934 0 2
rlabel polysilicon 240 -1940 240 -1940 0 3
rlabel polysilicon 243 -1940 243 -1940 0 4
rlabel polysilicon 247 -1934 247 -1934 0 1
rlabel polysilicon 247 -1940 247 -1940 0 3
rlabel polysilicon 254 -1934 254 -1934 0 1
rlabel polysilicon 254 -1940 254 -1940 0 3
rlabel polysilicon 261 -1934 261 -1934 0 1
rlabel polysilicon 261 -1940 261 -1940 0 3
rlabel polysilicon 268 -1934 268 -1934 0 1
rlabel polysilicon 268 -1940 268 -1940 0 3
rlabel polysilicon 275 -1934 275 -1934 0 1
rlabel polysilicon 275 -1940 275 -1940 0 3
rlabel polysilicon 282 -1934 282 -1934 0 1
rlabel polysilicon 285 -1934 285 -1934 0 2
rlabel polysilicon 282 -1940 282 -1940 0 3
rlabel polysilicon 289 -1934 289 -1934 0 1
rlabel polysilicon 289 -1940 289 -1940 0 3
rlabel polysilicon 296 -1934 296 -1934 0 1
rlabel polysilicon 296 -1940 296 -1940 0 3
rlabel polysilicon 303 -1934 303 -1934 0 1
rlabel polysilicon 303 -1940 303 -1940 0 3
rlabel polysilicon 310 -1934 310 -1934 0 1
rlabel polysilicon 310 -1940 310 -1940 0 3
rlabel polysilicon 317 -1934 317 -1934 0 1
rlabel polysilicon 317 -1940 317 -1940 0 3
rlabel polysilicon 320 -1940 320 -1940 0 4
rlabel polysilicon 324 -1934 324 -1934 0 1
rlabel polysilicon 324 -1940 324 -1940 0 3
rlabel polysilicon 331 -1934 331 -1934 0 1
rlabel polysilicon 334 -1934 334 -1934 0 2
rlabel polysilicon 331 -1940 331 -1940 0 3
rlabel polysilicon 334 -1940 334 -1940 0 4
rlabel polysilicon 338 -1934 338 -1934 0 1
rlabel polysilicon 338 -1940 338 -1940 0 3
rlabel polysilicon 345 -1934 345 -1934 0 1
rlabel polysilicon 345 -1940 345 -1940 0 3
rlabel polysilicon 352 -1934 352 -1934 0 1
rlabel polysilicon 352 -1940 352 -1940 0 3
rlabel polysilicon 359 -1934 359 -1934 0 1
rlabel polysilicon 359 -1940 359 -1940 0 3
rlabel polysilicon 366 -1934 366 -1934 0 1
rlabel polysilicon 366 -1940 366 -1940 0 3
rlabel polysilicon 373 -1934 373 -1934 0 1
rlabel polysilicon 373 -1940 373 -1940 0 3
rlabel polysilicon 380 -1934 380 -1934 0 1
rlabel polysilicon 380 -1940 380 -1940 0 3
rlabel polysilicon 387 -1934 387 -1934 0 1
rlabel polysilicon 387 -1940 387 -1940 0 3
rlabel polysilicon 394 -1934 394 -1934 0 1
rlabel polysilicon 394 -1940 394 -1940 0 3
rlabel polysilicon 401 -1934 401 -1934 0 1
rlabel polysilicon 401 -1940 401 -1940 0 3
rlabel polysilicon 408 -1934 408 -1934 0 1
rlabel polysilicon 411 -1934 411 -1934 0 2
rlabel polysilicon 408 -1940 408 -1940 0 3
rlabel polysilicon 411 -1940 411 -1940 0 4
rlabel polysilicon 418 -1934 418 -1934 0 2
rlabel polysilicon 415 -1940 415 -1940 0 3
rlabel polysilicon 418 -1940 418 -1940 0 4
rlabel polysilicon 422 -1934 422 -1934 0 1
rlabel polysilicon 422 -1940 422 -1940 0 3
rlabel polysilicon 429 -1934 429 -1934 0 1
rlabel polysilicon 429 -1940 429 -1940 0 3
rlabel polysilicon 436 -1934 436 -1934 0 1
rlabel polysilicon 439 -1934 439 -1934 0 2
rlabel polysilicon 436 -1940 436 -1940 0 3
rlabel polysilicon 439 -1940 439 -1940 0 4
rlabel polysilicon 443 -1934 443 -1934 0 1
rlabel polysilicon 443 -1940 443 -1940 0 3
rlabel polysilicon 450 -1934 450 -1934 0 1
rlabel polysilicon 453 -1934 453 -1934 0 2
rlabel polysilicon 450 -1940 450 -1940 0 3
rlabel polysilicon 453 -1940 453 -1940 0 4
rlabel polysilicon 457 -1934 457 -1934 0 1
rlabel polysilicon 460 -1934 460 -1934 0 2
rlabel polysilicon 457 -1940 457 -1940 0 3
rlabel polysilicon 460 -1940 460 -1940 0 4
rlabel polysilicon 464 -1934 464 -1934 0 1
rlabel polysilicon 464 -1940 464 -1940 0 3
rlabel polysilicon 471 -1934 471 -1934 0 1
rlabel polysilicon 474 -1940 474 -1940 0 4
rlabel polysilicon 478 -1934 478 -1934 0 1
rlabel polysilicon 478 -1940 478 -1940 0 3
rlabel polysilicon 485 -1934 485 -1934 0 1
rlabel polysilicon 485 -1940 485 -1940 0 3
rlabel polysilicon 492 -1934 492 -1934 0 1
rlabel polysilicon 492 -1940 492 -1940 0 3
rlabel polysilicon 499 -1934 499 -1934 0 1
rlabel polysilicon 499 -1940 499 -1940 0 3
rlabel polysilicon 502 -1940 502 -1940 0 4
rlabel polysilicon 506 -1934 506 -1934 0 1
rlabel polysilicon 506 -1940 506 -1940 0 3
rlabel polysilicon 513 -1934 513 -1934 0 1
rlabel polysilicon 513 -1940 513 -1940 0 3
rlabel polysilicon 520 -1934 520 -1934 0 1
rlabel polysilicon 520 -1940 520 -1940 0 3
rlabel polysilicon 527 -1934 527 -1934 0 1
rlabel polysilicon 527 -1940 527 -1940 0 3
rlabel polysilicon 534 -1934 534 -1934 0 1
rlabel polysilicon 534 -1940 534 -1940 0 3
rlabel polysilicon 541 -1934 541 -1934 0 1
rlabel polysilicon 541 -1940 541 -1940 0 3
rlabel polysilicon 548 -1934 548 -1934 0 1
rlabel polysilicon 548 -1940 548 -1940 0 3
rlabel polysilicon 555 -1934 555 -1934 0 1
rlabel polysilicon 555 -1940 555 -1940 0 3
rlabel polysilicon 562 -1934 562 -1934 0 1
rlabel polysilicon 562 -1940 562 -1940 0 3
rlabel polysilicon 569 -1934 569 -1934 0 1
rlabel polysilicon 569 -1940 569 -1940 0 3
rlabel polysilicon 576 -1934 576 -1934 0 1
rlabel polysilicon 576 -1940 576 -1940 0 3
rlabel polysilicon 579 -1940 579 -1940 0 4
rlabel polysilicon 583 -1934 583 -1934 0 1
rlabel polysilicon 583 -1940 583 -1940 0 3
rlabel polysilicon 590 -1940 590 -1940 0 3
rlabel polysilicon 593 -1940 593 -1940 0 4
rlabel polysilicon 597 -1934 597 -1934 0 1
rlabel polysilicon 597 -1940 597 -1940 0 3
rlabel polysilicon 604 -1934 604 -1934 0 1
rlabel polysilicon 604 -1940 604 -1940 0 3
rlabel polysilicon 611 -1934 611 -1934 0 1
rlabel polysilicon 611 -1940 611 -1940 0 3
rlabel polysilicon 618 -1934 618 -1934 0 1
rlabel polysilicon 618 -1940 618 -1940 0 3
rlabel polysilicon 625 -1934 625 -1934 0 1
rlabel polysilicon 625 -1940 625 -1940 0 3
rlabel polysilicon 632 -1934 632 -1934 0 1
rlabel polysilicon 632 -1940 632 -1940 0 3
rlabel polysilicon 639 -1934 639 -1934 0 1
rlabel polysilicon 639 -1940 639 -1940 0 3
rlabel polysilicon 646 -1934 646 -1934 0 1
rlabel polysilicon 646 -1940 646 -1940 0 3
rlabel polysilicon 653 -1934 653 -1934 0 1
rlabel polysilicon 653 -1940 653 -1940 0 3
rlabel polysilicon 660 -1934 660 -1934 0 1
rlabel polysilicon 660 -1940 660 -1940 0 3
rlabel polysilicon 667 -1934 667 -1934 0 1
rlabel polysilicon 667 -1940 667 -1940 0 3
rlabel polysilicon 674 -1934 674 -1934 0 1
rlabel polysilicon 674 -1940 674 -1940 0 3
rlabel polysilicon 681 -1934 681 -1934 0 1
rlabel polysilicon 681 -1940 681 -1940 0 3
rlabel polysilicon 684 -1940 684 -1940 0 4
rlabel polysilicon 688 -1934 688 -1934 0 1
rlabel polysilicon 688 -1940 688 -1940 0 3
rlabel polysilicon 695 -1934 695 -1934 0 1
rlabel polysilicon 695 -1940 695 -1940 0 3
rlabel polysilicon 702 -1934 702 -1934 0 1
rlabel polysilicon 702 -1940 702 -1940 0 3
rlabel polysilicon 709 -1934 709 -1934 0 1
rlabel polysilicon 709 -1940 709 -1940 0 3
rlabel polysilicon 716 -1934 716 -1934 0 1
rlabel polysilicon 716 -1940 716 -1940 0 3
rlabel polysilicon 723 -1934 723 -1934 0 1
rlabel polysilicon 723 -1940 723 -1940 0 3
rlabel polysilicon 730 -1934 730 -1934 0 1
rlabel polysilicon 730 -1940 730 -1940 0 3
rlabel polysilicon 737 -1934 737 -1934 0 1
rlabel polysilicon 737 -1940 737 -1940 0 3
rlabel polysilicon 744 -1934 744 -1934 0 1
rlabel polysilicon 744 -1940 744 -1940 0 3
rlabel polysilicon 751 -1934 751 -1934 0 1
rlabel polysilicon 751 -1940 751 -1940 0 3
rlabel polysilicon 758 -1934 758 -1934 0 1
rlabel polysilicon 761 -1934 761 -1934 0 2
rlabel polysilicon 758 -1940 758 -1940 0 3
rlabel polysilicon 765 -1934 765 -1934 0 1
rlabel polysilicon 765 -1940 765 -1940 0 3
rlabel polysilicon 772 -1934 772 -1934 0 1
rlabel polysilicon 772 -1940 772 -1940 0 3
rlabel polysilicon 782 -1934 782 -1934 0 2
rlabel polysilicon 779 -1940 779 -1940 0 3
rlabel polysilicon 782 -1940 782 -1940 0 4
rlabel polysilicon 786 -1934 786 -1934 0 1
rlabel polysilicon 786 -1940 786 -1940 0 3
rlabel polysilicon 793 -1934 793 -1934 0 1
rlabel polysilicon 793 -1940 793 -1940 0 3
rlabel polysilicon 814 -1934 814 -1934 0 1
rlabel polysilicon 814 -1940 814 -1940 0 3
rlabel polysilicon 821 -1934 821 -1934 0 1
rlabel polysilicon 821 -1940 821 -1940 0 3
rlabel polysilicon 37 -1993 37 -1993 0 1
rlabel polysilicon 37 -1999 37 -1999 0 3
rlabel polysilicon 44 -1993 44 -1993 0 1
rlabel polysilicon 44 -1999 44 -1999 0 3
rlabel polysilicon 51 -1993 51 -1993 0 1
rlabel polysilicon 51 -1999 51 -1999 0 3
rlabel polysilicon 58 -1993 58 -1993 0 1
rlabel polysilicon 58 -1999 58 -1999 0 3
rlabel polysilicon 65 -1993 65 -1993 0 1
rlabel polysilicon 65 -1999 65 -1999 0 3
rlabel polysilicon 72 -1993 72 -1993 0 1
rlabel polysilicon 72 -1999 72 -1999 0 3
rlabel polysilicon 79 -1993 79 -1993 0 1
rlabel polysilicon 79 -1999 79 -1999 0 3
rlabel polysilicon 86 -1993 86 -1993 0 1
rlabel polysilicon 86 -1999 86 -1999 0 3
rlabel polysilicon 93 -1993 93 -1993 0 1
rlabel polysilicon 93 -1999 93 -1999 0 3
rlabel polysilicon 100 -1993 100 -1993 0 1
rlabel polysilicon 100 -1999 100 -1999 0 3
rlabel polysilicon 107 -1993 107 -1993 0 1
rlabel polysilicon 107 -1999 107 -1999 0 3
rlabel polysilicon 114 -1993 114 -1993 0 1
rlabel polysilicon 114 -1999 114 -1999 0 3
rlabel polysilicon 121 -1993 121 -1993 0 1
rlabel polysilicon 121 -1999 121 -1999 0 3
rlabel polysilicon 128 -1993 128 -1993 0 1
rlabel polysilicon 128 -1999 128 -1999 0 3
rlabel polysilicon 135 -1993 135 -1993 0 1
rlabel polysilicon 138 -1993 138 -1993 0 2
rlabel polysilicon 135 -1999 135 -1999 0 3
rlabel polysilicon 142 -1993 142 -1993 0 1
rlabel polysilicon 142 -1999 142 -1999 0 3
rlabel polysilicon 149 -1993 149 -1993 0 1
rlabel polysilicon 149 -1999 149 -1999 0 3
rlabel polysilicon 156 -1993 156 -1993 0 1
rlabel polysilicon 159 -1993 159 -1993 0 2
rlabel polysilicon 163 -1993 163 -1993 0 1
rlabel polysilicon 163 -1999 163 -1999 0 3
rlabel polysilicon 170 -1993 170 -1993 0 1
rlabel polysilicon 170 -1999 170 -1999 0 3
rlabel polysilicon 177 -1993 177 -1993 0 1
rlabel polysilicon 177 -1999 177 -1999 0 3
rlabel polysilicon 184 -1993 184 -1993 0 1
rlabel polysilicon 184 -1999 184 -1999 0 3
rlabel polysilicon 191 -1993 191 -1993 0 1
rlabel polysilicon 191 -1999 191 -1999 0 3
rlabel polysilicon 198 -1993 198 -1993 0 1
rlabel polysilicon 198 -1999 198 -1999 0 3
rlabel polysilicon 201 -1999 201 -1999 0 4
rlabel polysilicon 205 -1993 205 -1993 0 1
rlabel polysilicon 205 -1999 205 -1999 0 3
rlabel polysilicon 212 -1993 212 -1993 0 1
rlabel polysilicon 212 -1999 212 -1999 0 3
rlabel polysilicon 219 -1993 219 -1993 0 1
rlabel polysilicon 219 -1999 219 -1999 0 3
rlabel polysilicon 229 -1993 229 -1993 0 2
rlabel polysilicon 229 -1999 229 -1999 0 4
rlabel polysilicon 233 -1993 233 -1993 0 1
rlabel polysilicon 233 -1999 233 -1999 0 3
rlabel polysilicon 240 -1999 240 -1999 0 3
rlabel polysilicon 243 -1999 243 -1999 0 4
rlabel polysilicon 247 -1993 247 -1993 0 1
rlabel polysilicon 247 -1999 247 -1999 0 3
rlabel polysilicon 254 -1993 254 -1993 0 1
rlabel polysilicon 254 -1999 254 -1999 0 3
rlabel polysilicon 261 -1993 261 -1993 0 1
rlabel polysilicon 264 -1993 264 -1993 0 2
rlabel polysilicon 261 -1999 261 -1999 0 3
rlabel polysilicon 264 -1999 264 -1999 0 4
rlabel polysilicon 268 -1993 268 -1993 0 1
rlabel polysilicon 271 -1993 271 -1993 0 2
rlabel polysilicon 271 -1999 271 -1999 0 4
rlabel polysilicon 275 -1993 275 -1993 0 1
rlabel polysilicon 275 -1999 275 -1999 0 3
rlabel polysilicon 282 -1993 282 -1993 0 1
rlabel polysilicon 282 -1999 282 -1999 0 3
rlabel polysilicon 289 -1999 289 -1999 0 3
rlabel polysilicon 292 -1999 292 -1999 0 4
rlabel polysilicon 296 -1993 296 -1993 0 1
rlabel polysilicon 296 -1999 296 -1999 0 3
rlabel polysilicon 303 -1993 303 -1993 0 1
rlabel polysilicon 303 -1999 303 -1999 0 3
rlabel polysilicon 313 -1999 313 -1999 0 4
rlabel polysilicon 317 -1993 317 -1993 0 1
rlabel polysilicon 317 -1999 317 -1999 0 3
rlabel polysilicon 324 -1993 324 -1993 0 1
rlabel polysilicon 324 -1999 324 -1999 0 3
rlabel polysilicon 331 -1993 331 -1993 0 1
rlabel polysilicon 331 -1999 331 -1999 0 3
rlabel polysilicon 338 -1993 338 -1993 0 1
rlabel polysilicon 338 -1999 338 -1999 0 3
rlabel polysilicon 345 -1993 345 -1993 0 1
rlabel polysilicon 345 -1999 345 -1999 0 3
rlabel polysilicon 352 -1993 352 -1993 0 1
rlabel polysilicon 352 -1999 352 -1999 0 3
rlabel polysilicon 359 -1993 359 -1993 0 1
rlabel polysilicon 359 -1999 359 -1999 0 3
rlabel polysilicon 369 -1993 369 -1993 0 2
rlabel polysilicon 373 -1993 373 -1993 0 1
rlabel polysilicon 373 -1999 373 -1999 0 3
rlabel polysilicon 380 -1993 380 -1993 0 1
rlabel polysilicon 380 -1999 380 -1999 0 3
rlabel polysilicon 387 -1993 387 -1993 0 1
rlabel polysilicon 387 -1999 387 -1999 0 3
rlabel polysilicon 394 -1993 394 -1993 0 1
rlabel polysilicon 394 -1999 394 -1999 0 3
rlabel polysilicon 401 -1993 401 -1993 0 1
rlabel polysilicon 401 -1999 401 -1999 0 3
rlabel polysilicon 408 -1993 408 -1993 0 1
rlabel polysilicon 408 -1999 408 -1999 0 3
rlabel polysilicon 415 -1993 415 -1993 0 1
rlabel polysilicon 415 -1999 415 -1999 0 3
rlabel polysilicon 422 -1993 422 -1993 0 1
rlabel polysilicon 422 -1999 422 -1999 0 3
rlabel polysilicon 432 -1993 432 -1993 0 2
rlabel polysilicon 429 -1999 429 -1999 0 3
rlabel polysilicon 432 -1999 432 -1999 0 4
rlabel polysilicon 436 -1993 436 -1993 0 1
rlabel polysilicon 439 -1993 439 -1993 0 2
rlabel polysilicon 446 -1993 446 -1993 0 2
rlabel polysilicon 443 -1999 443 -1999 0 3
rlabel polysilicon 446 -1999 446 -1999 0 4
rlabel polysilicon 450 -1993 450 -1993 0 1
rlabel polysilicon 450 -1999 450 -1999 0 3
rlabel polysilicon 457 -1993 457 -1993 0 1
rlabel polysilicon 457 -1999 457 -1999 0 3
rlabel polysilicon 464 -1993 464 -1993 0 1
rlabel polysilicon 464 -1999 464 -1999 0 3
rlabel polysilicon 471 -1993 471 -1993 0 1
rlabel polysilicon 471 -1999 471 -1999 0 3
rlabel polysilicon 478 -1993 478 -1993 0 1
rlabel polysilicon 478 -1999 478 -1999 0 3
rlabel polysilicon 485 -1993 485 -1993 0 1
rlabel polysilicon 485 -1999 485 -1999 0 3
rlabel polysilicon 492 -1993 492 -1993 0 1
rlabel polysilicon 495 -1993 495 -1993 0 2
rlabel polysilicon 492 -1999 492 -1999 0 3
rlabel polysilicon 499 -1993 499 -1993 0 1
rlabel polysilicon 499 -1999 499 -1999 0 3
rlabel polysilicon 506 -1993 506 -1993 0 1
rlabel polysilicon 506 -1999 506 -1999 0 3
rlabel polysilicon 516 -1993 516 -1993 0 2
rlabel polysilicon 513 -1999 513 -1999 0 3
rlabel polysilicon 520 -1993 520 -1993 0 1
rlabel polysilicon 520 -1999 520 -1999 0 3
rlabel polysilicon 527 -1993 527 -1993 0 1
rlabel polysilicon 527 -1999 527 -1999 0 3
rlabel polysilicon 534 -1993 534 -1993 0 1
rlabel polysilicon 534 -1999 534 -1999 0 3
rlabel polysilicon 541 -1993 541 -1993 0 1
rlabel polysilicon 541 -1999 541 -1999 0 3
rlabel polysilicon 548 -1993 548 -1993 0 1
rlabel polysilicon 548 -1999 548 -1999 0 3
rlabel polysilicon 555 -1993 555 -1993 0 1
rlabel polysilicon 555 -1999 555 -1999 0 3
rlabel polysilicon 562 -1993 562 -1993 0 1
rlabel polysilicon 562 -1999 562 -1999 0 3
rlabel polysilicon 569 -1993 569 -1993 0 1
rlabel polysilicon 569 -1999 569 -1999 0 3
rlabel polysilicon 576 -1993 576 -1993 0 1
rlabel polysilicon 576 -1999 576 -1999 0 3
rlabel polysilicon 583 -1999 583 -1999 0 3
rlabel polysilicon 586 -1999 586 -1999 0 4
rlabel polysilicon 593 -1993 593 -1993 0 2
rlabel polysilicon 590 -1999 590 -1999 0 3
rlabel polysilicon 593 -1999 593 -1999 0 4
rlabel polysilicon 597 -1993 597 -1993 0 1
rlabel polysilicon 597 -1999 597 -1999 0 3
rlabel polysilicon 600 -1999 600 -1999 0 4
rlabel polysilicon 604 -1993 604 -1993 0 1
rlabel polysilicon 604 -1999 604 -1999 0 3
rlabel polysilicon 611 -1993 611 -1993 0 1
rlabel polysilicon 611 -1999 611 -1999 0 3
rlabel polysilicon 618 -1993 618 -1993 0 1
rlabel polysilicon 618 -1999 618 -1999 0 3
rlabel polysilicon 625 -1993 625 -1993 0 1
rlabel polysilicon 625 -1999 625 -1999 0 3
rlabel polysilicon 632 -1993 632 -1993 0 1
rlabel polysilicon 632 -1999 632 -1999 0 3
rlabel polysilicon 639 -1993 639 -1993 0 1
rlabel polysilicon 639 -1999 639 -1999 0 3
rlabel polysilicon 646 -1993 646 -1993 0 1
rlabel polysilicon 646 -1999 646 -1999 0 3
rlabel polysilicon 653 -1993 653 -1993 0 1
rlabel polysilicon 653 -1999 653 -1999 0 3
rlabel polysilicon 660 -1999 660 -1999 0 3
rlabel polysilicon 663 -1999 663 -1999 0 4
rlabel polysilicon 667 -1993 667 -1993 0 1
rlabel polysilicon 667 -1999 667 -1999 0 3
rlabel polysilicon 674 -1993 674 -1993 0 1
rlabel polysilicon 677 -1993 677 -1993 0 2
rlabel polysilicon 674 -1999 674 -1999 0 3
rlabel polysilicon 677 -1999 677 -1999 0 4
rlabel polysilicon 681 -1993 681 -1993 0 1
rlabel polysilicon 681 -1999 681 -1999 0 3
rlabel polysilicon 688 -1993 688 -1993 0 1
rlabel polysilicon 691 -1999 691 -1999 0 4
rlabel polysilicon 695 -1993 695 -1993 0 1
rlabel polysilicon 695 -1999 695 -1999 0 3
rlabel polysilicon 702 -1993 702 -1993 0 1
rlabel polysilicon 702 -1999 702 -1999 0 3
rlabel polysilicon 709 -1993 709 -1993 0 1
rlabel polysilicon 709 -1999 709 -1999 0 3
rlabel polysilicon 716 -1993 716 -1993 0 1
rlabel polysilicon 716 -1999 716 -1999 0 3
rlabel polysilicon 723 -1993 723 -1993 0 1
rlabel polysilicon 726 -1993 726 -1993 0 2
rlabel polysilicon 730 -1993 730 -1993 0 1
rlabel polysilicon 730 -1999 730 -1999 0 3
rlabel polysilicon 737 -1993 737 -1993 0 1
rlabel polysilicon 737 -1999 737 -1999 0 3
rlabel polysilicon 744 -1993 744 -1993 0 1
rlabel polysilicon 744 -1999 744 -1999 0 3
rlabel polysilicon 751 -1993 751 -1993 0 1
rlabel polysilicon 751 -1999 751 -1999 0 3
rlabel polysilicon 758 -1993 758 -1993 0 1
rlabel polysilicon 758 -1999 758 -1999 0 3
rlabel polysilicon 765 -1993 765 -1993 0 1
rlabel polysilicon 765 -1999 765 -1999 0 3
rlabel polysilicon 772 -1993 772 -1993 0 1
rlabel polysilicon 772 -1999 772 -1999 0 3
rlabel polysilicon 779 -1993 779 -1993 0 1
rlabel polysilicon 786 -1993 786 -1993 0 1
rlabel polysilicon 786 -1999 786 -1999 0 3
rlabel polysilicon 793 -1999 793 -1999 0 3
rlabel polysilicon 796 -1999 796 -1999 0 4
rlabel polysilicon 800 -1993 800 -1993 0 1
rlabel polysilicon 800 -1999 800 -1999 0 3
rlabel polysilicon 807 -1993 807 -1993 0 1
rlabel polysilicon 807 -1999 807 -1999 0 3
rlabel polysilicon 814 -1993 814 -1993 0 1
rlabel polysilicon 814 -1999 814 -1999 0 3
rlabel polysilicon 16 -2056 16 -2056 0 1
rlabel polysilicon 16 -2062 16 -2062 0 3
rlabel polysilicon 23 -2056 23 -2056 0 1
rlabel polysilicon 23 -2062 23 -2062 0 3
rlabel polysilicon 30 -2056 30 -2056 0 1
rlabel polysilicon 30 -2062 30 -2062 0 3
rlabel polysilicon 37 -2056 37 -2056 0 1
rlabel polysilicon 37 -2062 37 -2062 0 3
rlabel polysilicon 44 -2056 44 -2056 0 1
rlabel polysilicon 44 -2062 44 -2062 0 3
rlabel polysilicon 51 -2056 51 -2056 0 1
rlabel polysilicon 51 -2062 51 -2062 0 3
rlabel polysilicon 58 -2056 58 -2056 0 1
rlabel polysilicon 58 -2062 58 -2062 0 3
rlabel polysilicon 65 -2056 65 -2056 0 1
rlabel polysilicon 65 -2062 65 -2062 0 3
rlabel polysilicon 72 -2056 72 -2056 0 1
rlabel polysilicon 72 -2062 72 -2062 0 3
rlabel polysilicon 79 -2056 79 -2056 0 1
rlabel polysilicon 79 -2062 79 -2062 0 3
rlabel polysilicon 86 -2056 86 -2056 0 1
rlabel polysilicon 86 -2062 86 -2062 0 3
rlabel polysilicon 93 -2056 93 -2056 0 1
rlabel polysilicon 93 -2062 93 -2062 0 3
rlabel polysilicon 100 -2056 100 -2056 0 1
rlabel polysilicon 100 -2062 100 -2062 0 3
rlabel polysilicon 107 -2056 107 -2056 0 1
rlabel polysilicon 107 -2062 107 -2062 0 3
rlabel polysilicon 114 -2056 114 -2056 0 1
rlabel polysilicon 114 -2062 114 -2062 0 3
rlabel polysilicon 121 -2056 121 -2056 0 1
rlabel polysilicon 124 -2062 124 -2062 0 4
rlabel polysilicon 128 -2056 128 -2056 0 1
rlabel polysilicon 128 -2062 128 -2062 0 3
rlabel polysilicon 131 -2062 131 -2062 0 4
rlabel polysilicon 135 -2056 135 -2056 0 1
rlabel polysilicon 135 -2062 135 -2062 0 3
rlabel polysilicon 142 -2056 142 -2056 0 1
rlabel polysilicon 142 -2062 142 -2062 0 3
rlabel polysilicon 145 -2062 145 -2062 0 4
rlabel polysilicon 149 -2056 149 -2056 0 1
rlabel polysilicon 149 -2062 149 -2062 0 3
rlabel polysilicon 156 -2056 156 -2056 0 1
rlabel polysilicon 156 -2062 156 -2062 0 3
rlabel polysilicon 166 -2056 166 -2056 0 2
rlabel polysilicon 163 -2062 163 -2062 0 3
rlabel polysilicon 170 -2056 170 -2056 0 1
rlabel polysilicon 170 -2062 170 -2062 0 3
rlabel polysilicon 177 -2062 177 -2062 0 3
rlabel polysilicon 180 -2062 180 -2062 0 4
rlabel polysilicon 184 -2056 184 -2056 0 1
rlabel polysilicon 187 -2056 187 -2056 0 2
rlabel polysilicon 184 -2062 184 -2062 0 3
rlabel polysilicon 187 -2062 187 -2062 0 4
rlabel polysilicon 191 -2056 191 -2056 0 1
rlabel polysilicon 191 -2062 191 -2062 0 3
rlabel polysilicon 198 -2056 198 -2056 0 1
rlabel polysilicon 198 -2062 198 -2062 0 3
rlabel polysilicon 205 -2056 205 -2056 0 1
rlabel polysilicon 205 -2062 205 -2062 0 3
rlabel polysilicon 212 -2056 212 -2056 0 1
rlabel polysilicon 212 -2062 212 -2062 0 3
rlabel polysilicon 219 -2056 219 -2056 0 1
rlabel polysilicon 219 -2062 219 -2062 0 3
rlabel polysilicon 226 -2056 226 -2056 0 1
rlabel polysilicon 229 -2056 229 -2056 0 2
rlabel polysilicon 229 -2062 229 -2062 0 4
rlabel polysilicon 233 -2056 233 -2056 0 1
rlabel polysilicon 236 -2056 236 -2056 0 2
rlabel polysilicon 233 -2062 233 -2062 0 3
rlabel polysilicon 236 -2062 236 -2062 0 4
rlabel polysilicon 243 -2056 243 -2056 0 2
rlabel polysilicon 240 -2062 240 -2062 0 3
rlabel polysilicon 243 -2062 243 -2062 0 4
rlabel polysilicon 247 -2056 247 -2056 0 1
rlabel polysilicon 247 -2062 247 -2062 0 3
rlabel polysilicon 254 -2056 254 -2056 0 1
rlabel polysilicon 257 -2056 257 -2056 0 2
rlabel polysilicon 254 -2062 254 -2062 0 3
rlabel polysilicon 257 -2062 257 -2062 0 4
rlabel polysilicon 261 -2056 261 -2056 0 1
rlabel polysilicon 261 -2062 261 -2062 0 3
rlabel polysilicon 268 -2056 268 -2056 0 1
rlabel polysilicon 268 -2062 268 -2062 0 3
rlabel polysilicon 275 -2056 275 -2056 0 1
rlabel polysilicon 275 -2062 275 -2062 0 3
rlabel polysilicon 282 -2056 282 -2056 0 1
rlabel polysilicon 282 -2062 282 -2062 0 3
rlabel polysilicon 289 -2056 289 -2056 0 1
rlabel polysilicon 289 -2062 289 -2062 0 3
rlabel polysilicon 296 -2056 296 -2056 0 1
rlabel polysilicon 296 -2062 296 -2062 0 3
rlabel polysilicon 303 -2056 303 -2056 0 1
rlabel polysilicon 303 -2062 303 -2062 0 3
rlabel polysilicon 310 -2056 310 -2056 0 1
rlabel polysilicon 310 -2062 310 -2062 0 3
rlabel polysilicon 317 -2056 317 -2056 0 1
rlabel polysilicon 317 -2062 317 -2062 0 3
rlabel polysilicon 324 -2056 324 -2056 0 1
rlabel polysilicon 324 -2062 324 -2062 0 3
rlabel polysilicon 331 -2056 331 -2056 0 1
rlabel polysilicon 331 -2062 331 -2062 0 3
rlabel polysilicon 338 -2056 338 -2056 0 1
rlabel polysilicon 338 -2062 338 -2062 0 3
rlabel polysilicon 345 -2056 345 -2056 0 1
rlabel polysilicon 348 -2056 348 -2056 0 2
rlabel polysilicon 345 -2062 345 -2062 0 3
rlabel polysilicon 352 -2056 352 -2056 0 1
rlabel polysilicon 352 -2062 352 -2062 0 3
rlabel polysilicon 359 -2056 359 -2056 0 1
rlabel polysilicon 359 -2062 359 -2062 0 3
rlabel polysilicon 366 -2056 366 -2056 0 1
rlabel polysilicon 366 -2062 366 -2062 0 3
rlabel polysilicon 373 -2056 373 -2056 0 1
rlabel polysilicon 373 -2062 373 -2062 0 3
rlabel polysilicon 380 -2056 380 -2056 0 1
rlabel polysilicon 380 -2062 380 -2062 0 3
rlabel polysilicon 387 -2056 387 -2056 0 1
rlabel polysilicon 387 -2062 387 -2062 0 3
rlabel polysilicon 394 -2056 394 -2056 0 1
rlabel polysilicon 397 -2056 397 -2056 0 2
rlabel polysilicon 394 -2062 394 -2062 0 3
rlabel polysilicon 397 -2062 397 -2062 0 4
rlabel polysilicon 401 -2056 401 -2056 0 1
rlabel polysilicon 404 -2056 404 -2056 0 2
rlabel polysilicon 408 -2056 408 -2056 0 1
rlabel polysilicon 408 -2062 408 -2062 0 3
rlabel polysilicon 415 -2056 415 -2056 0 1
rlabel polysilicon 418 -2056 418 -2056 0 2
rlabel polysilicon 415 -2062 415 -2062 0 3
rlabel polysilicon 418 -2062 418 -2062 0 4
rlabel polysilicon 422 -2056 422 -2056 0 1
rlabel polysilicon 422 -2062 422 -2062 0 3
rlabel polysilicon 432 -2056 432 -2056 0 2
rlabel polysilicon 432 -2062 432 -2062 0 4
rlabel polysilicon 436 -2056 436 -2056 0 1
rlabel polysilicon 436 -2062 436 -2062 0 3
rlabel polysilicon 443 -2056 443 -2056 0 1
rlabel polysilicon 443 -2062 443 -2062 0 3
rlabel polysilicon 450 -2056 450 -2056 0 1
rlabel polysilicon 450 -2062 450 -2062 0 3
rlabel polysilicon 457 -2056 457 -2056 0 1
rlabel polysilicon 460 -2056 460 -2056 0 2
rlabel polysilicon 457 -2062 457 -2062 0 3
rlabel polysilicon 460 -2062 460 -2062 0 4
rlabel polysilicon 464 -2056 464 -2056 0 1
rlabel polysilicon 464 -2062 464 -2062 0 3
rlabel polysilicon 474 -2056 474 -2056 0 2
rlabel polysilicon 471 -2062 471 -2062 0 3
rlabel polysilicon 474 -2062 474 -2062 0 4
rlabel polysilicon 478 -2056 478 -2056 0 1
rlabel polysilicon 478 -2062 478 -2062 0 3
rlabel polysilicon 488 -2056 488 -2056 0 2
rlabel polysilicon 485 -2062 485 -2062 0 3
rlabel polysilicon 488 -2062 488 -2062 0 4
rlabel polysilicon 492 -2056 492 -2056 0 1
rlabel polysilicon 492 -2062 492 -2062 0 3
rlabel polysilicon 499 -2056 499 -2056 0 1
rlabel polysilicon 499 -2062 499 -2062 0 3
rlabel polysilicon 506 -2062 506 -2062 0 3
rlabel polysilicon 509 -2062 509 -2062 0 4
rlabel polysilicon 513 -2056 513 -2056 0 1
rlabel polysilicon 513 -2062 513 -2062 0 3
rlabel polysilicon 516 -2062 516 -2062 0 4
rlabel polysilicon 520 -2056 520 -2056 0 1
rlabel polysilicon 520 -2062 520 -2062 0 3
rlabel polysilicon 527 -2056 527 -2056 0 1
rlabel polysilicon 527 -2062 527 -2062 0 3
rlabel polysilicon 534 -2056 534 -2056 0 1
rlabel polysilicon 534 -2062 534 -2062 0 3
rlabel polysilicon 541 -2056 541 -2056 0 1
rlabel polysilicon 541 -2062 541 -2062 0 3
rlabel polysilicon 548 -2056 548 -2056 0 1
rlabel polysilicon 548 -2062 548 -2062 0 3
rlabel polysilicon 555 -2056 555 -2056 0 1
rlabel polysilicon 555 -2062 555 -2062 0 3
rlabel polysilicon 565 -2056 565 -2056 0 2
rlabel polysilicon 562 -2062 562 -2062 0 3
rlabel polysilicon 569 -2056 569 -2056 0 1
rlabel polysilicon 569 -2062 569 -2062 0 3
rlabel polysilicon 576 -2056 576 -2056 0 1
rlabel polysilicon 576 -2062 576 -2062 0 3
rlabel polysilicon 583 -2056 583 -2056 0 1
rlabel polysilicon 583 -2062 583 -2062 0 3
rlabel polysilicon 590 -2056 590 -2056 0 1
rlabel polysilicon 590 -2062 590 -2062 0 3
rlabel polysilicon 597 -2056 597 -2056 0 1
rlabel polysilicon 597 -2062 597 -2062 0 3
rlabel polysilicon 604 -2056 604 -2056 0 1
rlabel polysilicon 604 -2062 604 -2062 0 3
rlabel polysilicon 611 -2056 611 -2056 0 1
rlabel polysilicon 611 -2062 611 -2062 0 3
rlabel polysilicon 618 -2056 618 -2056 0 1
rlabel polysilicon 618 -2062 618 -2062 0 3
rlabel polysilicon 625 -2056 625 -2056 0 1
rlabel polysilicon 625 -2062 625 -2062 0 3
rlabel polysilicon 632 -2056 632 -2056 0 1
rlabel polysilicon 632 -2062 632 -2062 0 3
rlabel polysilicon 639 -2056 639 -2056 0 1
rlabel polysilicon 639 -2062 639 -2062 0 3
rlabel polysilicon 646 -2056 646 -2056 0 1
rlabel polysilicon 646 -2062 646 -2062 0 3
rlabel polysilicon 653 -2056 653 -2056 0 1
rlabel polysilicon 660 -2056 660 -2056 0 1
rlabel polysilicon 660 -2062 660 -2062 0 3
rlabel polysilicon 667 -2056 667 -2056 0 1
rlabel polysilicon 670 -2056 670 -2056 0 2
rlabel polysilicon 670 -2062 670 -2062 0 4
rlabel polysilicon 674 -2056 674 -2056 0 1
rlabel polysilicon 674 -2062 674 -2062 0 3
rlabel polysilicon 681 -2056 681 -2056 0 1
rlabel polysilicon 681 -2062 681 -2062 0 3
rlabel polysilicon 688 -2056 688 -2056 0 1
rlabel polysilicon 688 -2062 688 -2062 0 3
rlabel polysilicon 695 -2056 695 -2056 0 1
rlabel polysilicon 695 -2062 695 -2062 0 3
rlabel polysilicon 702 -2056 702 -2056 0 1
rlabel polysilicon 702 -2062 702 -2062 0 3
rlabel polysilicon 709 -2056 709 -2056 0 1
rlabel polysilicon 709 -2062 709 -2062 0 3
rlabel polysilicon 716 -2056 716 -2056 0 1
rlabel polysilicon 716 -2062 716 -2062 0 3
rlabel polysilicon 726 -2056 726 -2056 0 2
rlabel polysilicon 723 -2062 723 -2062 0 3
rlabel polysilicon 726 -2062 726 -2062 0 4
rlabel polysilicon 730 -2056 730 -2056 0 1
rlabel polysilicon 730 -2062 730 -2062 0 3
rlabel polysilicon 737 -2056 737 -2056 0 1
rlabel polysilicon 737 -2062 737 -2062 0 3
rlabel polysilicon 744 -2056 744 -2056 0 1
rlabel polysilicon 744 -2062 744 -2062 0 3
rlabel polysilicon 751 -2056 751 -2056 0 1
rlabel polysilicon 751 -2062 751 -2062 0 3
rlabel polysilicon 758 -2056 758 -2056 0 1
rlabel polysilicon 758 -2062 758 -2062 0 3
rlabel polysilicon 765 -2056 765 -2056 0 1
rlabel polysilicon 765 -2062 765 -2062 0 3
rlabel polysilicon 772 -2056 772 -2056 0 1
rlabel polysilicon 772 -2062 772 -2062 0 3
rlabel polysilicon 779 -2056 779 -2056 0 1
rlabel polysilicon 779 -2062 779 -2062 0 3
rlabel polysilicon 786 -2056 786 -2056 0 1
rlabel polysilicon 786 -2062 786 -2062 0 3
rlabel polysilicon 16 -2121 16 -2121 0 1
rlabel polysilicon 16 -2127 16 -2127 0 3
rlabel polysilicon 23 -2121 23 -2121 0 1
rlabel polysilicon 23 -2127 23 -2127 0 3
rlabel polysilicon 30 -2121 30 -2121 0 1
rlabel polysilicon 30 -2127 30 -2127 0 3
rlabel polysilicon 40 -2127 40 -2127 0 4
rlabel polysilicon 44 -2121 44 -2121 0 1
rlabel polysilicon 44 -2127 44 -2127 0 3
rlabel polysilicon 51 -2121 51 -2121 0 1
rlabel polysilicon 51 -2127 51 -2127 0 3
rlabel polysilicon 58 -2121 58 -2121 0 1
rlabel polysilicon 58 -2127 58 -2127 0 3
rlabel polysilicon 65 -2121 65 -2121 0 1
rlabel polysilicon 65 -2127 65 -2127 0 3
rlabel polysilicon 72 -2121 72 -2121 0 1
rlabel polysilicon 72 -2127 72 -2127 0 3
rlabel polysilicon 79 -2121 79 -2121 0 1
rlabel polysilicon 79 -2127 79 -2127 0 3
rlabel polysilicon 86 -2121 86 -2121 0 1
rlabel polysilicon 86 -2127 86 -2127 0 3
rlabel polysilicon 93 -2121 93 -2121 0 1
rlabel polysilicon 96 -2121 96 -2121 0 2
rlabel polysilicon 103 -2121 103 -2121 0 2
rlabel polysilicon 100 -2127 100 -2127 0 3
rlabel polysilicon 107 -2121 107 -2121 0 1
rlabel polysilicon 107 -2127 107 -2127 0 3
rlabel polysilicon 114 -2121 114 -2121 0 1
rlabel polysilicon 114 -2127 114 -2127 0 3
rlabel polysilicon 121 -2121 121 -2121 0 1
rlabel polysilicon 121 -2127 121 -2127 0 3
rlabel polysilicon 128 -2121 128 -2121 0 1
rlabel polysilicon 128 -2127 128 -2127 0 3
rlabel polysilicon 135 -2121 135 -2121 0 1
rlabel polysilicon 138 -2121 138 -2121 0 2
rlabel polysilicon 135 -2127 135 -2127 0 3
rlabel polysilicon 142 -2121 142 -2121 0 1
rlabel polysilicon 142 -2127 142 -2127 0 3
rlabel polysilicon 149 -2121 149 -2121 0 1
rlabel polysilicon 149 -2127 149 -2127 0 3
rlabel polysilicon 156 -2121 156 -2121 0 1
rlabel polysilicon 156 -2127 156 -2127 0 3
rlabel polysilicon 159 -2127 159 -2127 0 4
rlabel polysilicon 163 -2121 163 -2121 0 1
rlabel polysilicon 163 -2127 163 -2127 0 3
rlabel polysilicon 173 -2121 173 -2121 0 2
rlabel polysilicon 170 -2127 170 -2127 0 3
rlabel polysilicon 173 -2127 173 -2127 0 4
rlabel polysilicon 177 -2121 177 -2121 0 1
rlabel polysilicon 180 -2121 180 -2121 0 2
rlabel polysilicon 177 -2127 177 -2127 0 3
rlabel polysilicon 180 -2127 180 -2127 0 4
rlabel polysilicon 184 -2121 184 -2121 0 1
rlabel polysilicon 191 -2121 191 -2121 0 1
rlabel polysilicon 191 -2127 191 -2127 0 3
rlabel polysilicon 198 -2121 198 -2121 0 1
rlabel polysilicon 198 -2127 198 -2127 0 3
rlabel polysilicon 201 -2127 201 -2127 0 4
rlabel polysilicon 205 -2121 205 -2121 0 1
rlabel polysilicon 205 -2127 205 -2127 0 3
rlabel polysilicon 208 -2127 208 -2127 0 4
rlabel polysilicon 212 -2121 212 -2121 0 1
rlabel polysilicon 212 -2127 212 -2127 0 3
rlabel polysilicon 219 -2121 219 -2121 0 1
rlabel polysilicon 219 -2127 219 -2127 0 3
rlabel polysilicon 222 -2127 222 -2127 0 4
rlabel polysilicon 229 -2121 229 -2121 0 2
rlabel polysilicon 226 -2127 226 -2127 0 3
rlabel polysilicon 233 -2121 233 -2121 0 1
rlabel polysilicon 233 -2127 233 -2127 0 3
rlabel polysilicon 240 -2121 240 -2121 0 1
rlabel polysilicon 240 -2127 240 -2127 0 3
rlabel polysilicon 247 -2121 247 -2121 0 1
rlabel polysilicon 250 -2127 250 -2127 0 4
rlabel polysilicon 254 -2121 254 -2121 0 1
rlabel polysilicon 254 -2127 254 -2127 0 3
rlabel polysilicon 261 -2121 261 -2121 0 1
rlabel polysilicon 261 -2127 261 -2127 0 3
rlabel polysilicon 268 -2121 268 -2121 0 1
rlabel polysilicon 268 -2127 268 -2127 0 3
rlabel polysilicon 275 -2121 275 -2121 0 1
rlabel polysilicon 275 -2127 275 -2127 0 3
rlabel polysilicon 282 -2121 282 -2121 0 1
rlabel polysilicon 282 -2127 282 -2127 0 3
rlabel polysilicon 289 -2121 289 -2121 0 1
rlabel polysilicon 292 -2121 292 -2121 0 2
rlabel polysilicon 296 -2121 296 -2121 0 1
rlabel polysilicon 296 -2127 296 -2127 0 3
rlabel polysilicon 303 -2121 303 -2121 0 1
rlabel polysilicon 303 -2127 303 -2127 0 3
rlabel polysilicon 310 -2121 310 -2121 0 1
rlabel polysilicon 310 -2127 310 -2127 0 3
rlabel polysilicon 317 -2121 317 -2121 0 1
rlabel polysilicon 320 -2121 320 -2121 0 2
rlabel polysilicon 320 -2127 320 -2127 0 4
rlabel polysilicon 324 -2121 324 -2121 0 1
rlabel polysilicon 324 -2127 324 -2127 0 3
rlabel polysilicon 331 -2121 331 -2121 0 1
rlabel polysilicon 331 -2127 331 -2127 0 3
rlabel polysilicon 338 -2121 338 -2121 0 1
rlabel polysilicon 338 -2127 338 -2127 0 3
rlabel polysilicon 348 -2121 348 -2121 0 2
rlabel polysilicon 345 -2127 345 -2127 0 3
rlabel polysilicon 348 -2127 348 -2127 0 4
rlabel polysilicon 352 -2121 352 -2121 0 1
rlabel polysilicon 352 -2127 352 -2127 0 3
rlabel polysilicon 362 -2121 362 -2121 0 2
rlabel polysilicon 362 -2127 362 -2127 0 4
rlabel polysilicon 366 -2121 366 -2121 0 1
rlabel polysilicon 366 -2127 366 -2127 0 3
rlabel polysilicon 373 -2121 373 -2121 0 1
rlabel polysilicon 373 -2127 373 -2127 0 3
rlabel polysilicon 383 -2121 383 -2121 0 2
rlabel polysilicon 380 -2127 380 -2127 0 3
rlabel polysilicon 387 -2121 387 -2121 0 1
rlabel polysilicon 387 -2127 387 -2127 0 3
rlabel polysilicon 394 -2121 394 -2121 0 1
rlabel polysilicon 394 -2127 394 -2127 0 3
rlabel polysilicon 401 -2121 401 -2121 0 1
rlabel polysilicon 401 -2127 401 -2127 0 3
rlabel polysilicon 411 -2121 411 -2121 0 2
rlabel polysilicon 408 -2127 408 -2127 0 3
rlabel polysilicon 411 -2127 411 -2127 0 4
rlabel polysilicon 415 -2121 415 -2121 0 1
rlabel polysilicon 415 -2127 415 -2127 0 3
rlabel polysilicon 422 -2121 422 -2121 0 1
rlabel polysilicon 422 -2127 422 -2127 0 3
rlabel polysilicon 429 -2121 429 -2121 0 1
rlabel polysilicon 429 -2127 429 -2127 0 3
rlabel polysilicon 439 -2121 439 -2121 0 2
rlabel polysilicon 439 -2127 439 -2127 0 4
rlabel polysilicon 443 -2121 443 -2121 0 1
rlabel polysilicon 443 -2127 443 -2127 0 3
rlabel polysilicon 450 -2121 450 -2121 0 1
rlabel polysilicon 450 -2127 450 -2127 0 3
rlabel polysilicon 457 -2121 457 -2121 0 1
rlabel polysilicon 460 -2121 460 -2121 0 2
rlabel polysilicon 464 -2121 464 -2121 0 1
rlabel polysilicon 464 -2127 464 -2127 0 3
rlabel polysilicon 467 -2127 467 -2127 0 4
rlabel polysilicon 474 -2121 474 -2121 0 2
rlabel polysilicon 471 -2127 471 -2127 0 3
rlabel polysilicon 474 -2127 474 -2127 0 4
rlabel polysilicon 478 -2121 478 -2121 0 1
rlabel polysilicon 478 -2127 478 -2127 0 3
rlabel polysilicon 485 -2121 485 -2121 0 1
rlabel polysilicon 485 -2127 485 -2127 0 3
rlabel polysilicon 492 -2121 492 -2121 0 1
rlabel polysilicon 492 -2127 492 -2127 0 3
rlabel polysilicon 499 -2121 499 -2121 0 1
rlabel polysilicon 499 -2127 499 -2127 0 3
rlabel polysilicon 506 -2121 506 -2121 0 1
rlabel polysilicon 506 -2127 506 -2127 0 3
rlabel polysilicon 509 -2127 509 -2127 0 4
rlabel polysilicon 513 -2121 513 -2121 0 1
rlabel polysilicon 513 -2127 513 -2127 0 3
rlabel polysilicon 520 -2121 520 -2121 0 1
rlabel polysilicon 520 -2127 520 -2127 0 3
rlabel polysilicon 527 -2121 527 -2121 0 1
rlabel polysilicon 527 -2127 527 -2127 0 3
rlabel polysilicon 534 -2121 534 -2121 0 1
rlabel polysilicon 534 -2127 534 -2127 0 3
rlabel polysilicon 541 -2121 541 -2121 0 1
rlabel polysilicon 541 -2127 541 -2127 0 3
rlabel polysilicon 548 -2121 548 -2121 0 1
rlabel polysilicon 548 -2127 548 -2127 0 3
rlabel polysilicon 555 -2121 555 -2121 0 1
rlabel polysilicon 555 -2127 555 -2127 0 3
rlabel polysilicon 562 -2121 562 -2121 0 1
rlabel polysilicon 562 -2127 562 -2127 0 3
rlabel polysilicon 569 -2121 569 -2121 0 1
rlabel polysilicon 569 -2127 569 -2127 0 3
rlabel polysilicon 576 -2121 576 -2121 0 1
rlabel polysilicon 576 -2127 576 -2127 0 3
rlabel polysilicon 583 -2121 583 -2121 0 1
rlabel polysilicon 583 -2127 583 -2127 0 3
rlabel polysilicon 593 -2121 593 -2121 0 2
rlabel polysilicon 593 -2127 593 -2127 0 4
rlabel polysilicon 597 -2121 597 -2121 0 1
rlabel polysilicon 597 -2127 597 -2127 0 3
rlabel polysilicon 604 -2121 604 -2121 0 1
rlabel polysilicon 604 -2127 604 -2127 0 3
rlabel polysilicon 611 -2121 611 -2121 0 1
rlabel polysilicon 611 -2127 611 -2127 0 3
rlabel polysilicon 618 -2121 618 -2121 0 1
rlabel polysilicon 618 -2127 618 -2127 0 3
rlabel polysilicon 625 -2121 625 -2121 0 1
rlabel polysilicon 625 -2127 625 -2127 0 3
rlabel polysilicon 632 -2121 632 -2121 0 1
rlabel polysilicon 632 -2127 632 -2127 0 3
rlabel polysilicon 639 -2121 639 -2121 0 1
rlabel polysilicon 639 -2127 639 -2127 0 3
rlabel polysilicon 646 -2121 646 -2121 0 1
rlabel polysilicon 646 -2127 646 -2127 0 3
rlabel polysilicon 653 -2121 653 -2121 0 1
rlabel polysilicon 653 -2127 653 -2127 0 3
rlabel polysilicon 660 -2121 660 -2121 0 1
rlabel polysilicon 660 -2127 660 -2127 0 3
rlabel polysilicon 667 -2121 667 -2121 0 1
rlabel polysilicon 667 -2127 667 -2127 0 3
rlabel polysilicon 674 -2121 674 -2121 0 1
rlabel polysilicon 674 -2127 674 -2127 0 3
rlabel polysilicon 681 -2121 681 -2121 0 1
rlabel polysilicon 681 -2127 681 -2127 0 3
rlabel polysilicon 688 -2121 688 -2121 0 1
rlabel polysilicon 688 -2127 688 -2127 0 3
rlabel polysilicon 695 -2121 695 -2121 0 1
rlabel polysilicon 695 -2127 695 -2127 0 3
rlabel polysilicon 702 -2121 702 -2121 0 1
rlabel polysilicon 702 -2127 702 -2127 0 3
rlabel polysilicon 709 -2121 709 -2121 0 1
rlabel polysilicon 709 -2127 709 -2127 0 3
rlabel polysilicon 716 -2121 716 -2121 0 1
rlabel polysilicon 716 -2127 716 -2127 0 3
rlabel polysilicon 723 -2121 723 -2121 0 1
rlabel polysilicon 723 -2127 723 -2127 0 3
rlabel polysilicon 730 -2127 730 -2127 0 3
rlabel polysilicon 737 -2121 737 -2121 0 1
rlabel polysilicon 737 -2127 737 -2127 0 3
rlabel polysilicon 86 -2172 86 -2172 0 1
rlabel polysilicon 86 -2178 86 -2178 0 3
rlabel polysilicon 100 -2172 100 -2172 0 1
rlabel polysilicon 100 -2178 100 -2178 0 3
rlabel polysilicon 107 -2172 107 -2172 0 1
rlabel polysilicon 107 -2178 107 -2178 0 3
rlabel polysilicon 114 -2172 114 -2172 0 1
rlabel polysilicon 114 -2178 114 -2178 0 3
rlabel polysilicon 121 -2172 121 -2172 0 1
rlabel polysilicon 121 -2178 121 -2178 0 3
rlabel polysilicon 128 -2172 128 -2172 0 1
rlabel polysilicon 128 -2178 128 -2178 0 3
rlabel polysilicon 131 -2178 131 -2178 0 4
rlabel polysilicon 135 -2172 135 -2172 0 1
rlabel polysilicon 142 -2172 142 -2172 0 1
rlabel polysilicon 142 -2178 142 -2178 0 3
rlabel polysilicon 152 -2172 152 -2172 0 2
rlabel polysilicon 152 -2178 152 -2178 0 4
rlabel polysilicon 156 -2172 156 -2172 0 1
rlabel polysilicon 159 -2172 159 -2172 0 2
rlabel polysilicon 156 -2178 156 -2178 0 3
rlabel polysilicon 163 -2172 163 -2172 0 1
rlabel polysilicon 163 -2178 163 -2178 0 3
rlabel polysilicon 170 -2172 170 -2172 0 1
rlabel polysilicon 170 -2178 170 -2178 0 3
rlabel polysilicon 177 -2172 177 -2172 0 1
rlabel polysilicon 177 -2178 177 -2178 0 3
rlabel polysilicon 184 -2172 184 -2172 0 1
rlabel polysilicon 184 -2178 184 -2178 0 3
rlabel polysilicon 191 -2172 191 -2172 0 1
rlabel polysilicon 191 -2178 191 -2178 0 3
rlabel polysilicon 198 -2172 198 -2172 0 1
rlabel polysilicon 198 -2178 198 -2178 0 3
rlabel polysilicon 205 -2172 205 -2172 0 1
rlabel polysilicon 205 -2178 205 -2178 0 3
rlabel polysilicon 212 -2172 212 -2172 0 1
rlabel polysilicon 212 -2178 212 -2178 0 3
rlabel polysilicon 219 -2172 219 -2172 0 1
rlabel polysilicon 222 -2172 222 -2172 0 2
rlabel polysilicon 219 -2178 219 -2178 0 3
rlabel polysilicon 222 -2178 222 -2178 0 4
rlabel polysilicon 226 -2172 226 -2172 0 1
rlabel polysilicon 229 -2172 229 -2172 0 2
rlabel polysilicon 233 -2172 233 -2172 0 1
rlabel polysilicon 233 -2178 233 -2178 0 3
rlabel polysilicon 240 -2178 240 -2178 0 3
rlabel polysilicon 243 -2178 243 -2178 0 4
rlabel polysilicon 247 -2172 247 -2172 0 1
rlabel polysilicon 247 -2178 247 -2178 0 3
rlabel polysilicon 254 -2172 254 -2172 0 1
rlabel polysilicon 254 -2178 254 -2178 0 3
rlabel polysilicon 261 -2172 261 -2172 0 1
rlabel polysilicon 261 -2178 261 -2178 0 3
rlabel polysilicon 268 -2172 268 -2172 0 1
rlabel polysilicon 268 -2178 268 -2178 0 3
rlabel polysilicon 275 -2172 275 -2172 0 1
rlabel polysilicon 275 -2178 275 -2178 0 3
rlabel polysilicon 282 -2172 282 -2172 0 1
rlabel polysilicon 285 -2172 285 -2172 0 2
rlabel polysilicon 282 -2178 282 -2178 0 3
rlabel polysilicon 285 -2178 285 -2178 0 4
rlabel polysilicon 289 -2172 289 -2172 0 1
rlabel polysilicon 289 -2178 289 -2178 0 3
rlabel polysilicon 296 -2172 296 -2172 0 1
rlabel polysilicon 299 -2178 299 -2178 0 4
rlabel polysilicon 303 -2172 303 -2172 0 1
rlabel polysilicon 303 -2178 303 -2178 0 3
rlabel polysilicon 310 -2172 310 -2172 0 1
rlabel polysilicon 313 -2172 313 -2172 0 2
rlabel polysilicon 310 -2178 310 -2178 0 3
rlabel polysilicon 317 -2172 317 -2172 0 1
rlabel polysilicon 317 -2178 317 -2178 0 3
rlabel polysilicon 324 -2172 324 -2172 0 1
rlabel polysilicon 324 -2178 324 -2178 0 3
rlabel polysilicon 331 -2172 331 -2172 0 1
rlabel polysilicon 334 -2172 334 -2172 0 2
rlabel polysilicon 331 -2178 331 -2178 0 3
rlabel polysilicon 338 -2172 338 -2172 0 1
rlabel polysilicon 338 -2178 338 -2178 0 3
rlabel polysilicon 345 -2172 345 -2172 0 1
rlabel polysilicon 345 -2178 345 -2178 0 3
rlabel polysilicon 352 -2172 352 -2172 0 1
rlabel polysilicon 352 -2178 352 -2178 0 3
rlabel polysilicon 359 -2172 359 -2172 0 1
rlabel polysilicon 359 -2178 359 -2178 0 3
rlabel polysilicon 366 -2172 366 -2172 0 1
rlabel polysilicon 366 -2178 366 -2178 0 3
rlabel polysilicon 373 -2172 373 -2172 0 1
rlabel polysilicon 373 -2178 373 -2178 0 3
rlabel polysilicon 380 -2172 380 -2172 0 1
rlabel polysilicon 380 -2178 380 -2178 0 3
rlabel polysilicon 387 -2172 387 -2172 0 1
rlabel polysilicon 390 -2172 390 -2172 0 2
rlabel polysilicon 390 -2178 390 -2178 0 4
rlabel polysilicon 394 -2172 394 -2172 0 1
rlabel polysilicon 394 -2178 394 -2178 0 3
rlabel polysilicon 401 -2172 401 -2172 0 1
rlabel polysilicon 401 -2178 401 -2178 0 3
rlabel polysilicon 408 -2172 408 -2172 0 1
rlabel polysilicon 411 -2178 411 -2178 0 4
rlabel polysilicon 415 -2172 415 -2172 0 1
rlabel polysilicon 415 -2178 415 -2178 0 3
rlabel polysilicon 422 -2172 422 -2172 0 1
rlabel polysilicon 422 -2178 422 -2178 0 3
rlabel polysilicon 429 -2172 429 -2172 0 1
rlabel polysilicon 429 -2178 429 -2178 0 3
rlabel polysilicon 432 -2178 432 -2178 0 4
rlabel polysilicon 436 -2172 436 -2172 0 1
rlabel polysilicon 436 -2178 436 -2178 0 3
rlabel polysilicon 443 -2172 443 -2172 0 1
rlabel polysilicon 443 -2178 443 -2178 0 3
rlabel polysilicon 453 -2172 453 -2172 0 2
rlabel polysilicon 450 -2178 450 -2178 0 3
rlabel polysilicon 457 -2172 457 -2172 0 1
rlabel polysilicon 460 -2178 460 -2178 0 4
rlabel polysilicon 464 -2172 464 -2172 0 1
rlabel polysilicon 464 -2178 464 -2178 0 3
rlabel polysilicon 471 -2172 471 -2172 0 1
rlabel polysilicon 471 -2178 471 -2178 0 3
rlabel polysilicon 478 -2172 478 -2172 0 1
rlabel polysilicon 478 -2178 478 -2178 0 3
rlabel polysilicon 485 -2172 485 -2172 0 1
rlabel polysilicon 485 -2178 485 -2178 0 3
rlabel polysilicon 492 -2178 492 -2178 0 3
rlabel polysilicon 499 -2172 499 -2172 0 1
rlabel polysilicon 499 -2178 499 -2178 0 3
rlabel polysilicon 509 -2172 509 -2172 0 2
rlabel polysilicon 509 -2178 509 -2178 0 4
rlabel polysilicon 513 -2172 513 -2172 0 1
rlabel polysilicon 513 -2178 513 -2178 0 3
rlabel polysilicon 520 -2172 520 -2172 0 1
rlabel polysilicon 520 -2178 520 -2178 0 3
rlabel polysilicon 527 -2172 527 -2172 0 1
rlabel polysilicon 527 -2178 527 -2178 0 3
rlabel polysilicon 534 -2172 534 -2172 0 1
rlabel polysilicon 534 -2178 534 -2178 0 3
rlabel polysilicon 541 -2172 541 -2172 0 1
rlabel polysilicon 541 -2178 541 -2178 0 3
rlabel polysilicon 548 -2172 548 -2172 0 1
rlabel polysilicon 548 -2178 548 -2178 0 3
rlabel polysilicon 555 -2172 555 -2172 0 1
rlabel polysilicon 558 -2172 558 -2172 0 2
rlabel polysilicon 555 -2178 555 -2178 0 3
rlabel polysilicon 558 -2178 558 -2178 0 4
rlabel polysilicon 562 -2172 562 -2172 0 1
rlabel polysilicon 562 -2178 562 -2178 0 3
rlabel polysilicon 569 -2172 569 -2172 0 1
rlabel polysilicon 569 -2178 569 -2178 0 3
rlabel polysilicon 576 -2172 576 -2172 0 1
rlabel polysilicon 579 -2172 579 -2172 0 2
rlabel polysilicon 576 -2178 576 -2178 0 3
rlabel polysilicon 583 -2178 583 -2178 0 3
rlabel polysilicon 586 -2178 586 -2178 0 4
rlabel polysilicon 590 -2172 590 -2172 0 1
rlabel polysilicon 590 -2178 590 -2178 0 3
rlabel polysilicon 597 -2172 597 -2172 0 1
rlabel polysilicon 597 -2178 597 -2178 0 3
rlabel polysilicon 604 -2172 604 -2172 0 1
rlabel polysilicon 604 -2178 604 -2178 0 3
rlabel polysilicon 611 -2172 611 -2172 0 1
rlabel polysilicon 611 -2178 611 -2178 0 3
rlabel polysilicon 618 -2172 618 -2172 0 1
rlabel polysilicon 618 -2178 618 -2178 0 3
rlabel polysilicon 625 -2172 625 -2172 0 1
rlabel polysilicon 625 -2178 625 -2178 0 3
rlabel polysilicon 632 -2172 632 -2172 0 1
rlabel polysilicon 632 -2178 632 -2178 0 3
rlabel polysilicon 639 -2172 639 -2172 0 1
rlabel polysilicon 639 -2178 639 -2178 0 3
rlabel polysilicon 646 -2172 646 -2172 0 1
rlabel polysilicon 646 -2178 646 -2178 0 3
rlabel polysilicon 653 -2172 653 -2172 0 1
rlabel polysilicon 653 -2178 653 -2178 0 3
rlabel polysilicon 660 -2172 660 -2172 0 1
rlabel polysilicon 660 -2178 660 -2178 0 3
rlabel polysilicon 667 -2172 667 -2172 0 1
rlabel polysilicon 667 -2178 667 -2178 0 3
rlabel polysilicon 670 -2178 670 -2178 0 4
rlabel polysilicon 674 -2172 674 -2172 0 1
rlabel polysilicon 674 -2178 674 -2178 0 3
rlabel polysilicon 681 -2178 681 -2178 0 3
rlabel polysilicon 688 -2172 688 -2172 0 1
rlabel polysilicon 688 -2178 688 -2178 0 3
rlabel polysilicon 695 -2172 695 -2172 0 1
rlabel polysilicon 698 -2172 698 -2172 0 2
rlabel polysilicon 702 -2172 702 -2172 0 1
rlabel polysilicon 702 -2178 702 -2178 0 3
rlabel polysilicon 709 -2172 709 -2172 0 1
rlabel polysilicon 709 -2178 709 -2178 0 3
rlabel polysilicon 716 -2172 716 -2172 0 1
rlabel polysilicon 716 -2178 716 -2178 0 3
rlabel polysilicon 723 -2172 723 -2172 0 1
rlabel polysilicon 723 -2178 723 -2178 0 3
rlabel polysilicon 89 -2225 89 -2225 0 2
rlabel polysilicon 107 -2225 107 -2225 0 1
rlabel polysilicon 107 -2231 107 -2231 0 3
rlabel polysilicon 114 -2225 114 -2225 0 1
rlabel polysilicon 114 -2231 114 -2231 0 3
rlabel polysilicon 124 -2225 124 -2225 0 2
rlabel polysilicon 124 -2231 124 -2231 0 4
rlabel polysilicon 131 -2225 131 -2225 0 2
rlabel polysilicon 128 -2231 128 -2231 0 3
rlabel polysilicon 138 -2231 138 -2231 0 4
rlabel polysilicon 142 -2225 142 -2225 0 1
rlabel polysilicon 142 -2231 142 -2231 0 3
rlabel polysilicon 149 -2225 149 -2225 0 1
rlabel polysilicon 149 -2231 149 -2231 0 3
rlabel polysilicon 156 -2225 156 -2225 0 1
rlabel polysilicon 156 -2231 156 -2231 0 3
rlabel polysilicon 163 -2231 163 -2231 0 3
rlabel polysilicon 166 -2231 166 -2231 0 4
rlabel polysilicon 170 -2225 170 -2225 0 1
rlabel polysilicon 173 -2231 173 -2231 0 4
rlabel polysilicon 177 -2225 177 -2225 0 1
rlabel polysilicon 177 -2231 177 -2231 0 3
rlabel polysilicon 180 -2231 180 -2231 0 4
rlabel polysilicon 184 -2225 184 -2225 0 1
rlabel polysilicon 184 -2231 184 -2231 0 3
rlabel polysilicon 191 -2225 191 -2225 0 1
rlabel polysilicon 191 -2231 191 -2231 0 3
rlabel polysilicon 201 -2231 201 -2231 0 4
rlabel polysilicon 205 -2225 205 -2225 0 1
rlabel polysilicon 208 -2231 208 -2231 0 4
rlabel polysilicon 212 -2225 212 -2225 0 1
rlabel polysilicon 212 -2231 212 -2231 0 3
rlabel polysilicon 219 -2225 219 -2225 0 1
rlabel polysilicon 219 -2231 219 -2231 0 3
rlabel polysilicon 226 -2231 226 -2231 0 3
rlabel polysilicon 229 -2231 229 -2231 0 4
rlabel polysilicon 233 -2225 233 -2225 0 1
rlabel polysilicon 233 -2231 233 -2231 0 3
rlabel polysilicon 240 -2225 240 -2225 0 1
rlabel polysilicon 240 -2231 240 -2231 0 3
rlabel polysilicon 247 -2225 247 -2225 0 1
rlabel polysilicon 247 -2231 247 -2231 0 3
rlabel polysilicon 254 -2225 254 -2225 0 1
rlabel polysilicon 254 -2231 254 -2231 0 3
rlabel polysilicon 261 -2225 261 -2225 0 1
rlabel polysilicon 261 -2231 261 -2231 0 3
rlabel polysilicon 268 -2225 268 -2225 0 1
rlabel polysilicon 268 -2231 268 -2231 0 3
rlabel polysilicon 275 -2225 275 -2225 0 1
rlabel polysilicon 275 -2231 275 -2231 0 3
rlabel polysilicon 285 -2225 285 -2225 0 2
rlabel polysilicon 282 -2231 282 -2231 0 3
rlabel polysilicon 289 -2225 289 -2225 0 1
rlabel polysilicon 289 -2231 289 -2231 0 3
rlabel polysilicon 296 -2225 296 -2225 0 1
rlabel polysilicon 296 -2231 296 -2231 0 3
rlabel polysilicon 306 -2225 306 -2225 0 2
rlabel polysilicon 303 -2231 303 -2231 0 3
rlabel polysilicon 306 -2231 306 -2231 0 4
rlabel polysilicon 310 -2225 310 -2225 0 1
rlabel polysilicon 310 -2231 310 -2231 0 3
rlabel polysilicon 317 -2225 317 -2225 0 1
rlabel polysilicon 317 -2231 317 -2231 0 3
rlabel polysilicon 324 -2225 324 -2225 0 1
rlabel polysilicon 324 -2231 324 -2231 0 3
rlabel polysilicon 331 -2225 331 -2225 0 1
rlabel polysilicon 331 -2231 331 -2231 0 3
rlabel polysilicon 338 -2225 338 -2225 0 1
rlabel polysilicon 338 -2231 338 -2231 0 3
rlabel polysilicon 345 -2225 345 -2225 0 1
rlabel polysilicon 345 -2231 345 -2231 0 3
rlabel polysilicon 352 -2225 352 -2225 0 1
rlabel polysilicon 352 -2231 352 -2231 0 3
rlabel polysilicon 359 -2231 359 -2231 0 3
rlabel polysilicon 366 -2225 366 -2225 0 1
rlabel polysilicon 366 -2231 366 -2231 0 3
rlabel polysilicon 373 -2231 373 -2231 0 3
rlabel polysilicon 376 -2231 376 -2231 0 4
rlabel polysilicon 380 -2225 380 -2225 0 1
rlabel polysilicon 380 -2231 380 -2231 0 3
rlabel polysilicon 387 -2225 387 -2225 0 1
rlabel polysilicon 390 -2225 390 -2225 0 2
rlabel polysilicon 390 -2231 390 -2231 0 4
rlabel polysilicon 394 -2225 394 -2225 0 1
rlabel polysilicon 394 -2231 394 -2231 0 3
rlabel polysilicon 401 -2225 401 -2225 0 1
rlabel polysilicon 401 -2231 401 -2231 0 3
rlabel polysilicon 408 -2225 408 -2225 0 1
rlabel polysilicon 408 -2231 408 -2231 0 3
rlabel polysilicon 415 -2225 415 -2225 0 1
rlabel polysilicon 415 -2231 415 -2231 0 3
rlabel polysilicon 425 -2225 425 -2225 0 2
rlabel polysilicon 425 -2231 425 -2231 0 4
rlabel polysilicon 429 -2225 429 -2225 0 1
rlabel polysilicon 429 -2231 429 -2231 0 3
rlabel polysilicon 436 -2225 436 -2225 0 1
rlabel polysilicon 436 -2231 436 -2231 0 3
rlabel polysilicon 443 -2231 443 -2231 0 3
rlabel polysilicon 446 -2231 446 -2231 0 4
rlabel polysilicon 450 -2225 450 -2225 0 1
rlabel polysilicon 450 -2231 450 -2231 0 3
rlabel polysilicon 457 -2225 457 -2225 0 1
rlabel polysilicon 457 -2231 457 -2231 0 3
rlabel polysilicon 464 -2225 464 -2225 0 1
rlabel polysilicon 464 -2231 464 -2231 0 3
rlabel polysilicon 467 -2231 467 -2231 0 4
rlabel polysilicon 471 -2225 471 -2225 0 1
rlabel polysilicon 471 -2231 471 -2231 0 3
rlabel polysilicon 478 -2225 478 -2225 0 1
rlabel polysilicon 478 -2231 478 -2231 0 3
rlabel polysilicon 485 -2225 485 -2225 0 1
rlabel polysilicon 485 -2231 485 -2231 0 3
rlabel polysilicon 492 -2225 492 -2225 0 1
rlabel polysilicon 492 -2231 492 -2231 0 3
rlabel polysilicon 499 -2225 499 -2225 0 1
rlabel polysilicon 499 -2231 499 -2231 0 3
rlabel polysilicon 506 -2225 506 -2225 0 1
rlabel polysilicon 506 -2231 506 -2231 0 3
rlabel polysilicon 513 -2225 513 -2225 0 1
rlabel polysilicon 513 -2231 513 -2231 0 3
rlabel polysilicon 520 -2225 520 -2225 0 1
rlabel polysilicon 520 -2231 520 -2231 0 3
rlabel polysilicon 527 -2225 527 -2225 0 1
rlabel polysilicon 527 -2231 527 -2231 0 3
rlabel polysilicon 534 -2225 534 -2225 0 1
rlabel polysilicon 534 -2231 534 -2231 0 3
rlabel polysilicon 541 -2225 541 -2225 0 1
rlabel polysilicon 541 -2231 541 -2231 0 3
rlabel polysilicon 548 -2225 548 -2225 0 1
rlabel polysilicon 548 -2231 548 -2231 0 3
rlabel polysilicon 555 -2225 555 -2225 0 1
rlabel polysilicon 555 -2231 555 -2231 0 3
rlabel polysilicon 562 -2225 562 -2225 0 1
rlabel polysilicon 565 -2231 565 -2231 0 4
rlabel polysilicon 569 -2225 569 -2225 0 1
rlabel polysilicon 569 -2231 569 -2231 0 3
rlabel polysilicon 579 -2225 579 -2225 0 2
rlabel polysilicon 576 -2231 576 -2231 0 3
rlabel polysilicon 579 -2231 579 -2231 0 4
rlabel polysilicon 583 -2225 583 -2225 0 1
rlabel polysilicon 583 -2231 583 -2231 0 3
rlabel polysilicon 590 -2225 590 -2225 0 1
rlabel polysilicon 590 -2231 590 -2231 0 3
rlabel polysilicon 597 -2225 597 -2225 0 1
rlabel polysilicon 597 -2231 597 -2231 0 3
rlabel polysilicon 604 -2225 604 -2225 0 1
rlabel polysilicon 607 -2231 607 -2231 0 4
rlabel polysilicon 614 -2225 614 -2225 0 2
rlabel polysilicon 611 -2231 611 -2231 0 3
rlabel polysilicon 618 -2225 618 -2225 0 1
rlabel polysilicon 621 -2225 621 -2225 0 2
rlabel polysilicon 625 -2225 625 -2225 0 1
rlabel polysilicon 632 -2225 632 -2225 0 1
rlabel polysilicon 632 -2231 632 -2231 0 3
rlabel polysilicon 639 -2225 639 -2225 0 1
rlabel polysilicon 639 -2231 639 -2231 0 3
rlabel polysilicon 660 -2225 660 -2225 0 1
rlabel polysilicon 660 -2231 660 -2231 0 3
rlabel polysilicon 114 -2262 114 -2262 0 1
rlabel polysilicon 114 -2268 114 -2268 0 3
rlabel polysilicon 121 -2262 121 -2262 0 1
rlabel polysilicon 124 -2262 124 -2262 0 2
rlabel polysilicon 124 -2268 124 -2268 0 4
rlabel polysilicon 131 -2262 131 -2262 0 2
rlabel polysilicon 131 -2268 131 -2268 0 4
rlabel polysilicon 135 -2262 135 -2262 0 1
rlabel polysilicon 135 -2268 135 -2268 0 3
rlabel polysilicon 145 -2262 145 -2262 0 2
rlabel polysilicon 142 -2268 142 -2268 0 3
rlabel polysilicon 145 -2268 145 -2268 0 4
rlabel polysilicon 149 -2262 149 -2262 0 1
rlabel polysilicon 156 -2262 156 -2262 0 1
rlabel polysilicon 156 -2268 156 -2268 0 3
rlabel polysilicon 163 -2262 163 -2262 0 1
rlabel polysilicon 163 -2268 163 -2268 0 3
rlabel polysilicon 170 -2262 170 -2262 0 1
rlabel polysilicon 170 -2268 170 -2268 0 3
rlabel polysilicon 177 -2262 177 -2262 0 1
rlabel polysilicon 177 -2268 177 -2268 0 3
rlabel polysilicon 184 -2262 184 -2262 0 1
rlabel polysilicon 184 -2268 184 -2268 0 3
rlabel polysilicon 191 -2262 191 -2262 0 1
rlabel polysilicon 194 -2262 194 -2262 0 2
rlabel polysilicon 198 -2262 198 -2262 0 1
rlabel polysilicon 198 -2268 198 -2268 0 3
rlabel polysilicon 205 -2262 205 -2262 0 1
rlabel polysilicon 205 -2268 205 -2268 0 3
rlabel polysilicon 212 -2262 212 -2262 0 1
rlabel polysilicon 212 -2268 212 -2268 0 3
rlabel polysilicon 215 -2268 215 -2268 0 4
rlabel polysilicon 219 -2262 219 -2262 0 1
rlabel polysilicon 219 -2268 219 -2268 0 3
rlabel polysilicon 226 -2262 226 -2262 0 1
rlabel polysilicon 226 -2268 226 -2268 0 3
rlabel polysilicon 236 -2262 236 -2262 0 2
rlabel polysilicon 233 -2268 233 -2268 0 3
rlabel polysilicon 240 -2262 240 -2262 0 1
rlabel polysilicon 243 -2268 243 -2268 0 4
rlabel polysilicon 247 -2262 247 -2262 0 1
rlabel polysilicon 247 -2268 247 -2268 0 3
rlabel polysilicon 254 -2262 254 -2262 0 1
rlabel polysilicon 254 -2268 254 -2268 0 3
rlabel polysilicon 261 -2262 261 -2262 0 1
rlabel polysilicon 261 -2268 261 -2268 0 3
rlabel polysilicon 268 -2262 268 -2262 0 1
rlabel polysilicon 268 -2268 268 -2268 0 3
rlabel polysilicon 275 -2262 275 -2262 0 1
rlabel polysilicon 275 -2268 275 -2268 0 3
rlabel polysilicon 282 -2262 282 -2262 0 1
rlabel polysilicon 282 -2268 282 -2268 0 3
rlabel polysilicon 289 -2262 289 -2262 0 1
rlabel polysilicon 289 -2268 289 -2268 0 3
rlabel polysilicon 296 -2262 296 -2262 0 1
rlabel polysilicon 296 -2268 296 -2268 0 3
rlabel polysilicon 303 -2262 303 -2262 0 1
rlabel polysilicon 306 -2262 306 -2262 0 2
rlabel polysilicon 303 -2268 303 -2268 0 3
rlabel polysilicon 306 -2268 306 -2268 0 4
rlabel polysilicon 313 -2262 313 -2262 0 2
rlabel polysilicon 313 -2268 313 -2268 0 4
rlabel polysilicon 317 -2262 317 -2262 0 1
rlabel polysilicon 317 -2268 317 -2268 0 3
rlabel polysilicon 324 -2262 324 -2262 0 1
rlabel polysilicon 327 -2262 327 -2262 0 2
rlabel polysilicon 331 -2262 331 -2262 0 1
rlabel polysilicon 331 -2268 331 -2268 0 3
rlabel polysilicon 338 -2262 338 -2262 0 1
rlabel polysilicon 338 -2268 338 -2268 0 3
rlabel polysilicon 345 -2262 345 -2262 0 1
rlabel polysilicon 345 -2268 345 -2268 0 3
rlabel polysilicon 352 -2262 352 -2262 0 1
rlabel polysilicon 352 -2268 352 -2268 0 3
rlabel polysilicon 359 -2262 359 -2262 0 1
rlabel polysilicon 362 -2262 362 -2262 0 2
rlabel polysilicon 359 -2268 359 -2268 0 3
rlabel polysilicon 362 -2268 362 -2268 0 4
rlabel polysilicon 366 -2262 366 -2262 0 1
rlabel polysilicon 366 -2268 366 -2268 0 3
rlabel polysilicon 373 -2262 373 -2262 0 1
rlabel polysilicon 373 -2268 373 -2268 0 3
rlabel polysilicon 380 -2262 380 -2262 0 1
rlabel polysilicon 380 -2268 380 -2268 0 3
rlabel polysilicon 390 -2262 390 -2262 0 2
rlabel polysilicon 387 -2268 387 -2268 0 3
rlabel polysilicon 394 -2262 394 -2262 0 1
rlabel polysilicon 397 -2262 397 -2262 0 2
rlabel polysilicon 401 -2262 401 -2262 0 1
rlabel polysilicon 401 -2268 401 -2268 0 3
rlabel polysilicon 408 -2262 408 -2262 0 1
rlabel polysilicon 408 -2268 408 -2268 0 3
rlabel polysilicon 415 -2262 415 -2262 0 1
rlabel polysilicon 415 -2268 415 -2268 0 3
rlabel polysilicon 422 -2262 422 -2262 0 1
rlabel polysilicon 422 -2268 422 -2268 0 3
rlabel polysilicon 432 -2262 432 -2262 0 2
rlabel polysilicon 429 -2268 429 -2268 0 3
rlabel polysilicon 432 -2268 432 -2268 0 4
rlabel polysilicon 436 -2262 436 -2262 0 1
rlabel polysilicon 436 -2268 436 -2268 0 3
rlabel polysilicon 443 -2262 443 -2262 0 1
rlabel polysilicon 443 -2268 443 -2268 0 3
rlabel polysilicon 450 -2262 450 -2262 0 1
rlabel polysilicon 450 -2268 450 -2268 0 3
rlabel polysilicon 457 -2262 457 -2262 0 1
rlabel polysilicon 457 -2268 457 -2268 0 3
rlabel polysilicon 464 -2262 464 -2262 0 1
rlabel polysilicon 464 -2268 464 -2268 0 3
rlabel polysilicon 471 -2268 471 -2268 0 3
rlabel polysilicon 474 -2268 474 -2268 0 4
rlabel polysilicon 478 -2262 478 -2262 0 1
rlabel polysilicon 478 -2268 478 -2268 0 3
rlabel polysilicon 485 -2262 485 -2262 0 1
rlabel polysilicon 485 -2268 485 -2268 0 3
rlabel polysilicon 492 -2262 492 -2262 0 1
rlabel polysilicon 492 -2268 492 -2268 0 3
rlabel polysilicon 499 -2262 499 -2262 0 1
rlabel polysilicon 499 -2268 499 -2268 0 3
rlabel polysilicon 506 -2262 506 -2262 0 1
rlabel polysilicon 506 -2268 506 -2268 0 3
rlabel polysilicon 513 -2262 513 -2262 0 1
rlabel polysilicon 513 -2268 513 -2268 0 3
rlabel polysilicon 520 -2262 520 -2262 0 1
rlabel polysilicon 520 -2268 520 -2268 0 3
rlabel polysilicon 527 -2262 527 -2262 0 1
rlabel polysilicon 527 -2268 527 -2268 0 3
rlabel polysilicon 534 -2262 534 -2262 0 1
rlabel polysilicon 534 -2268 534 -2268 0 3
rlabel polysilicon 541 -2262 541 -2262 0 1
rlabel polysilicon 541 -2268 541 -2268 0 3
rlabel polysilicon 548 -2262 548 -2262 0 1
rlabel polysilicon 548 -2268 548 -2268 0 3
rlabel polysilicon 555 -2262 555 -2262 0 1
rlabel polysilicon 555 -2268 555 -2268 0 3
rlabel polysilicon 562 -2262 562 -2262 0 1
rlabel polysilicon 565 -2262 565 -2262 0 2
rlabel polysilicon 569 -2268 569 -2268 0 3
rlabel polysilicon 576 -2262 576 -2262 0 1
rlabel polysilicon 576 -2268 576 -2268 0 3
rlabel polysilicon 583 -2262 583 -2262 0 1
rlabel polysilicon 583 -2268 583 -2268 0 3
rlabel polysilicon 639 -2262 639 -2262 0 1
rlabel polysilicon 639 -2268 639 -2268 0 3
rlabel polysilicon 121 -2289 121 -2289 0 1
rlabel polysilicon 177 -2289 177 -2289 0 1
rlabel polysilicon 177 -2295 177 -2295 0 3
rlabel polysilicon 212 -2289 212 -2289 0 1
rlabel polysilicon 212 -2295 212 -2295 0 3
rlabel polysilicon 222 -2289 222 -2289 0 2
rlabel polysilicon 226 -2289 226 -2289 0 1
rlabel polysilicon 226 -2295 226 -2295 0 3
rlabel polysilicon 233 -2289 233 -2289 0 1
rlabel polysilicon 233 -2295 233 -2295 0 3
rlabel polysilicon 240 -2289 240 -2289 0 1
rlabel polysilicon 243 -2295 243 -2295 0 4
rlabel polysilicon 250 -2289 250 -2289 0 2
rlabel polysilicon 254 -2289 254 -2289 0 1
rlabel polysilicon 254 -2295 254 -2295 0 3
rlabel polysilicon 268 -2289 268 -2289 0 1
rlabel polysilicon 268 -2295 268 -2295 0 3
rlabel polysilicon 275 -2289 275 -2289 0 1
rlabel polysilicon 275 -2295 275 -2295 0 3
rlabel polysilicon 282 -2289 282 -2289 0 1
rlabel polysilicon 282 -2295 282 -2295 0 3
rlabel polysilicon 289 -2289 289 -2289 0 1
rlabel polysilicon 289 -2295 289 -2295 0 3
rlabel polysilicon 296 -2289 296 -2289 0 1
rlabel polysilicon 296 -2295 296 -2295 0 3
rlabel polysilicon 303 -2289 303 -2289 0 1
rlabel polysilicon 306 -2295 306 -2295 0 4
rlabel polysilicon 310 -2289 310 -2289 0 1
rlabel polysilicon 310 -2295 310 -2295 0 3
rlabel polysilicon 317 -2289 317 -2289 0 1
rlabel polysilicon 317 -2295 317 -2295 0 3
rlabel polysilicon 327 -2295 327 -2295 0 4
rlabel polysilicon 331 -2289 331 -2289 0 1
rlabel polysilicon 331 -2295 331 -2295 0 3
rlabel polysilicon 338 -2295 338 -2295 0 3
rlabel polysilicon 345 -2289 345 -2289 0 1
rlabel polysilicon 345 -2295 345 -2295 0 3
rlabel polysilicon 366 -2289 366 -2289 0 1
rlabel polysilicon 366 -2295 366 -2295 0 3
rlabel polysilicon 380 -2289 380 -2289 0 1
rlabel polysilicon 380 -2295 380 -2295 0 3
rlabel polysilicon 404 -2289 404 -2289 0 2
rlabel polysilicon 415 -2289 415 -2289 0 1
rlabel polysilicon 415 -2295 415 -2295 0 3
rlabel polysilicon 422 -2289 422 -2289 0 1
rlabel polysilicon 422 -2295 422 -2295 0 3
rlabel polysilicon 432 -2295 432 -2295 0 4
rlabel polysilicon 439 -2289 439 -2289 0 2
rlabel polysilicon 439 -2295 439 -2295 0 4
rlabel polysilicon 443 -2295 443 -2295 0 3
rlabel polysilicon 446 -2295 446 -2295 0 4
rlabel polysilicon 450 -2289 450 -2289 0 1
rlabel polysilicon 450 -2295 450 -2295 0 3
rlabel polysilicon 457 -2289 457 -2289 0 1
rlabel polysilicon 457 -2295 457 -2295 0 3
rlabel polysilicon 464 -2289 464 -2289 0 1
rlabel polysilicon 464 -2295 464 -2295 0 3
rlabel polysilicon 474 -2289 474 -2289 0 2
rlabel polysilicon 478 -2289 478 -2289 0 1
rlabel polysilicon 502 -2289 502 -2289 0 2
rlabel polysilicon 502 -2295 502 -2295 0 4
rlabel polysilicon 506 -2289 506 -2289 0 1
rlabel polysilicon 506 -2295 506 -2295 0 3
rlabel polysilicon 513 -2289 513 -2289 0 1
rlabel polysilicon 513 -2295 513 -2295 0 3
rlabel polysilicon 520 -2289 520 -2289 0 1
rlabel polysilicon 520 -2295 520 -2295 0 3
rlabel polysilicon 527 -2289 527 -2289 0 1
rlabel polysilicon 530 -2289 530 -2289 0 2
rlabel polysilicon 534 -2289 534 -2289 0 1
rlabel polysilicon 534 -2295 534 -2295 0 3
rlabel polysilicon 541 -2289 541 -2289 0 1
rlabel polysilicon 541 -2295 541 -2295 0 3
rlabel polysilicon 548 -2289 548 -2289 0 1
rlabel polysilicon 572 -2289 572 -2289 0 2
rlabel polysilicon 569 -2295 569 -2295 0 3
rlabel polysilicon 576 -2289 576 -2289 0 1
rlabel polysilicon 576 -2295 576 -2295 0 3
rlabel polysilicon 639 -2289 639 -2289 0 1
rlabel polysilicon 639 -2295 639 -2295 0 3
rlabel polysilicon 170 -2312 170 -2312 0 3
rlabel polysilicon 177 -2306 177 -2306 0 1
rlabel polysilicon 177 -2312 177 -2312 0 3
rlabel polysilicon 215 -2306 215 -2306 0 2
rlabel polysilicon 226 -2306 226 -2306 0 1
rlabel polysilicon 226 -2312 226 -2312 0 3
rlabel polysilicon 233 -2306 233 -2306 0 1
rlabel polysilicon 233 -2312 233 -2312 0 3
rlabel polysilicon 240 -2312 240 -2312 0 3
rlabel polysilicon 247 -2306 247 -2306 0 1
rlabel polysilicon 247 -2312 247 -2312 0 3
rlabel polysilicon 254 -2306 254 -2306 0 1
rlabel polysilicon 254 -2312 254 -2312 0 3
rlabel polysilicon 264 -2306 264 -2306 0 2
rlabel polysilicon 268 -2312 268 -2312 0 3
rlabel polysilicon 275 -2312 275 -2312 0 3
rlabel polysilicon 278 -2312 278 -2312 0 4
rlabel polysilicon 285 -2306 285 -2306 0 2
rlabel polysilicon 282 -2312 282 -2312 0 3
rlabel polysilicon 289 -2306 289 -2306 0 1
rlabel polysilicon 296 -2306 296 -2306 0 1
rlabel polysilicon 296 -2312 296 -2312 0 3
rlabel polysilicon 306 -2312 306 -2312 0 4
rlabel polysilicon 313 -2306 313 -2306 0 2
rlabel polysilicon 317 -2306 317 -2306 0 1
rlabel polysilicon 317 -2312 317 -2312 0 3
rlabel polysilicon 369 -2306 369 -2306 0 2
rlabel polysilicon 380 -2306 380 -2306 0 1
rlabel polysilicon 380 -2312 380 -2312 0 3
rlabel polysilicon 387 -2312 387 -2312 0 3
rlabel polysilicon 404 -2312 404 -2312 0 4
rlabel polysilicon 408 -2306 408 -2306 0 1
rlabel polysilicon 408 -2312 408 -2312 0 3
rlabel polysilicon 509 -2306 509 -2306 0 2
rlabel polysilicon 527 -2306 527 -2306 0 1
rlabel polysilicon 527 -2312 527 -2312 0 3
rlabel polysilicon 534 -2312 534 -2312 0 3
rlabel polysilicon 597 -2306 597 -2306 0 1
rlabel polysilicon 597 -2312 597 -2312 0 3
rlabel polysilicon 604 -2306 604 -2306 0 1
rlabel polysilicon 614 -2306 614 -2306 0 2
rlabel polysilicon 611 -2312 611 -2312 0 3
rlabel polysilicon 639 -2306 639 -2306 0 1
rlabel polysilicon 642 -2312 642 -2312 0 4
rlabel polysilicon 646 -2306 646 -2306 0 1
rlabel polysilicon 646 -2312 646 -2312 0 3
rlabel metal2 177 1 177 1 0 net=3643
rlabel metal2 205 1 205 1 0 net=6163
rlabel metal2 257 1 257 1 0 net=2849
rlabel metal2 310 1 310 1 0 net=3565
rlabel metal2 359 1 359 1 0 net=5247
rlabel metal2 271 -1 271 -1 0 net=1385
rlabel metal2 177 -12 177 -12 0 net=3644
rlabel metal2 194 -12 194 -12 0 net=677
rlabel metal2 212 -12 212 -12 0 net=6165
rlabel metal2 233 -12 233 -12 0 net=3399
rlabel metal2 261 -12 261 -12 0 net=1387
rlabel metal2 282 -12 282 -12 0 net=2851
rlabel metal2 282 -12 282 -12 0 net=2851
rlabel metal2 303 -12 303 -12 0 net=3567
rlabel metal2 341 -12 341 -12 0 net=5329
rlabel metal2 184 -14 184 -14 0 net=1089
rlabel metal2 215 -14 215 -14 0 net=6603
rlabel metal2 348 -14 348 -14 0 net=4139
rlabel metal2 198 -16 198 -16 0 net=620
rlabel metal2 240 -16 240 -16 0 net=1403
rlabel metal2 366 -16 366 -16 0 net=5249
rlabel metal2 366 -18 366 -18 0 net=2435
rlabel metal2 156 -29 156 -29 0 net=5051
rlabel metal2 156 -29 156 -29 0 net=5051
rlabel metal2 166 -29 166 -29 0 net=2281
rlabel metal2 205 -29 205 -29 0 net=2319
rlabel metal2 282 -29 282 -29 0 net=2853
rlabel metal2 282 -29 282 -29 0 net=2853
rlabel metal2 289 -29 289 -29 0 net=5099
rlabel metal2 299 -29 299 -29 0 net=4179
rlabel metal2 387 -29 387 -29 0 net=4141
rlabel metal2 177 -31 177 -31 0 net=3823
rlabel metal2 215 -31 215 -31 0 net=6166
rlabel metal2 226 -31 226 -31 0 net=1405
rlabel metal2 247 -31 247 -31 0 net=1389
rlabel metal2 268 -31 268 -31 0 net=2865
rlabel metal2 345 -31 345 -31 0 net=2437
rlabel metal2 380 -31 380 -31 0 net=4371
rlabel metal2 394 -31 394 -31 0 net=5331
rlabel metal2 194 -33 194 -33 0 net=3531
rlabel metal2 296 -33 296 -33 0 net=4641
rlabel metal2 373 -33 373 -33 0 net=5251
rlabel metal2 411 -33 411 -33 0 net=5161
rlabel metal2 212 -35 212 -35 0 net=3400
rlabel metal2 254 -35 254 -35 0 net=6605
rlabel metal2 317 -35 317 -35 0 net=4907
rlabel metal2 366 -35 366 -35 0 net=3675
rlabel metal2 380 -35 380 -35 0 net=5447
rlabel metal2 219 -37 219 -37 0 net=1475
rlabel metal2 261 -37 261 -37 0 net=2977
rlabel metal2 233 -39 233 -39 0 net=2399
rlabel metal2 303 -39 303 -39 0 net=3569
rlabel metal2 86 -50 86 -50 0 net=2755
rlabel metal2 121 -50 121 -50 0 net=2253
rlabel metal2 142 -50 142 -50 0 net=5571
rlabel metal2 177 -50 177 -50 0 net=3824
rlabel metal2 191 -50 191 -50 0 net=1477
rlabel metal2 233 -50 233 -50 0 net=6606
rlabel metal2 317 -50 317 -50 0 net=4909
rlabel metal2 579 -50 579 -50 0 net=4065
rlabel metal2 93 -52 93 -52 0 net=4687
rlabel metal2 107 -52 107 -52 0 net=2187
rlabel metal2 177 -52 177 -52 0 net=1407
rlabel metal2 247 -52 247 -52 0 net=1391
rlabel metal2 303 -52 303 -52 0 net=4180
rlabel metal2 355 -52 355 -52 0 net=4115
rlabel metal2 436 -52 436 -52 0 net=6843
rlabel metal2 135 -54 135 -54 0 net=5655
rlabel metal2 247 -54 247 -54 0 net=2979
rlabel metal2 268 -54 268 -54 0 net=2867
rlabel metal2 268 -54 268 -54 0 net=2867
rlabel metal2 275 -54 275 -54 0 net=3533
rlabel metal2 394 -54 394 -54 0 net=5253
rlabel metal2 443 -54 443 -54 0 net=5321
rlabel metal2 149 -56 149 -56 0 net=3073
rlabel metal2 275 -56 275 -56 0 net=2043
rlabel metal2 376 -56 376 -56 0 net=4671
rlabel metal2 429 -56 429 -56 0 net=4143
rlabel metal2 450 -56 450 -56 0 net=5163
rlabel metal2 156 -58 156 -58 0 net=5052
rlabel metal2 156 -58 156 -58 0 net=5052
rlabel metal2 163 -58 163 -58 0 net=3445
rlabel metal2 240 -58 240 -58 0 net=2401
rlabel metal2 303 -58 303 -58 0 net=2439
rlabel metal2 348 -58 348 -58 0 net=5537
rlabel metal2 205 -60 205 -60 0 net=2321
rlabel metal2 331 -60 331 -60 0 net=4642
rlabel metal2 422 -60 422 -60 0 net=5333
rlabel metal2 198 -62 198 -62 0 net=2283
rlabel metal2 215 -62 215 -62 0 net=1663
rlabel metal2 324 -62 324 -62 0 net=3571
rlabel metal2 338 -62 338 -62 0 net=3099
rlabel metal2 387 -62 387 -62 0 net=4373
rlabel metal2 100 -64 100 -64 0 net=4077
rlabel metal2 289 -64 289 -64 0 net=5101
rlabel metal2 282 -66 282 -66 0 net=2855
rlabel metal2 310 -66 310 -66 0 net=2485
rlabel metal2 338 -66 338 -66 0 net=5448
rlabel metal2 282 -68 282 -68 0 net=1967
rlabel metal2 341 -70 341 -70 0 net=4309
rlabel metal2 362 -72 362 -72 0 net=5789
rlabel metal2 366 -74 366 -74 0 net=3677
rlabel metal2 401 -76 401 -76 0 net=3657
rlabel metal2 58 -87 58 -87 0 net=5657
rlabel metal2 149 -87 149 -87 0 net=3074
rlabel metal2 282 -87 282 -87 0 net=1969
rlabel metal2 313 -87 313 -87 0 net=3678
rlabel metal2 436 -87 436 -87 0 net=5255
rlabel metal2 562 -87 562 -87 0 net=1399
rlabel metal2 562 -87 562 -87 0 net=1399
rlabel metal2 565 -87 565 -87 0 net=3207
rlabel metal2 65 -89 65 -89 0 net=5573
rlabel metal2 177 -89 177 -89 0 net=1409
rlabel metal2 247 -89 247 -89 0 net=2981
rlabel metal2 436 -89 436 -89 0 net=6697
rlabel metal2 583 -89 583 -89 0 net=4067
rlabel metal2 72 -91 72 -91 0 net=4427
rlabel metal2 282 -91 282 -91 0 net=2856
rlabel metal2 324 -91 324 -91 0 net=2487
rlabel metal2 324 -91 324 -91 0 net=2487
rlabel metal2 345 -91 345 -91 0 net=3658
rlabel metal2 443 -91 443 -91 0 net=4145
rlabel metal2 443 -91 443 -91 0 net=4145
rlabel metal2 450 -91 450 -91 0 net=5335
rlabel metal2 79 -93 79 -93 0 net=3449
rlabel metal2 121 -93 121 -93 0 net=1479
rlabel metal2 205 -93 205 -93 0 net=2285
rlabel metal2 268 -93 268 -93 0 net=2869
rlabel metal2 457 -93 457 -93 0 net=5165
rlabel metal2 86 -95 86 -95 0 net=2756
rlabel metal2 128 -95 128 -95 0 net=2255
rlabel metal2 128 -95 128 -95 0 net=2255
rlabel metal2 180 -95 180 -95 0 net=6809
rlabel metal2 86 -97 86 -97 0 net=3447
rlabel metal2 184 -97 184 -97 0 net=1913
rlabel metal2 205 -97 205 -97 0 net=1665
rlabel metal2 247 -97 247 -97 0 net=1393
rlabel metal2 317 -97 317 -97 0 net=2323
rlabel metal2 348 -97 348 -97 0 net=4910
rlabel metal2 478 -97 478 -97 0 net=5539
rlabel metal2 93 -99 93 -99 0 net=4688
rlabel metal2 149 -99 149 -99 0 net=2863
rlabel metal2 187 -99 187 -99 0 net=449
rlabel metal2 268 -99 268 -99 0 net=2735
rlabel metal2 352 -99 352 -99 0 net=4310
rlabel metal2 485 -99 485 -99 0 net=6845
rlabel metal2 93 -101 93 -101 0 net=3223
rlabel metal2 163 -101 163 -101 0 net=2189
rlabel metal2 226 -101 226 -101 0 net=1150
rlabel metal2 331 -101 331 -101 0 net=3573
rlabel metal2 114 -103 114 -103 0 net=1939
rlabel metal2 275 -103 275 -103 0 net=2045
rlabel metal2 331 -103 331 -103 0 net=5489
rlabel metal2 170 -105 170 -105 0 net=1679
rlabel metal2 289 -105 289 -105 0 net=2441
rlabel metal2 355 -105 355 -105 0 net=5322
rlabel metal2 156 -107 156 -107 0 net=2347
rlabel metal2 306 -107 306 -107 0 net=3673
rlabel metal2 243 -109 243 -109 0 net=270
rlabel metal2 261 -111 261 -111 0 net=2403
rlabel metal2 359 -111 359 -111 0 net=5790
rlabel metal2 222 -113 222 -113 0 net=1755
rlabel metal2 362 -113 362 -113 0 net=330
rlabel metal2 387 -113 387 -113 0 net=5103
rlabel metal2 107 -115 107 -115 0 net=2903
rlabel metal2 366 -115 366 -115 0 net=5275
rlabel metal2 142 -117 142 -117 0 net=2451
rlabel metal2 369 -117 369 -117 0 net=3971
rlabel metal2 177 -119 177 -119 0 net=673
rlabel metal2 373 -119 373 -119 0 net=3535
rlabel metal2 100 -121 100 -121 0 net=4078
rlabel metal2 376 -121 376 -121 0 net=5169
rlabel metal2 100 -123 100 -123 0 net=4751
rlabel metal2 387 -123 387 -123 0 net=6767
rlabel metal2 394 -125 394 -125 0 net=4673
rlabel metal2 334 -127 334 -127 0 net=5871
rlabel metal2 408 -127 408 -127 0 net=4117
rlabel metal2 380 -129 380 -129 0 net=3101
rlabel metal2 422 -129 422 -129 0 net=4375
rlabel metal2 422 -131 422 -131 0 net=5823
rlabel metal2 51 -142 51 -142 0 net=575
rlabel metal2 208 -142 208 -142 0 net=1193
rlabel metal2 380 -142 380 -142 0 net=3674
rlabel metal2 485 -142 485 -142 0 net=4377
rlabel metal2 485 -142 485 -142 0 net=4377
rlabel metal2 544 -142 544 -142 0 net=579
rlabel metal2 618 -142 618 -142 0 net=3209
rlabel metal2 642 -142 642 -142 0 net=6861
rlabel metal2 65 -144 65 -144 0 net=5574
rlabel metal2 222 -144 222 -144 0 net=2286
rlabel metal2 282 -144 282 -144 0 net=3574
rlabel metal2 439 -144 439 -144 0 net=5490
rlabel metal2 65 -146 65 -146 0 net=2905
rlabel metal2 121 -146 121 -146 0 net=1480
rlabel metal2 236 -146 236 -146 0 net=2404
rlabel metal2 282 -146 282 -146 0 net=2047
rlabel metal2 320 -146 320 -146 0 net=2870
rlabel metal2 457 -146 457 -146 0 net=4675
rlabel metal2 506 -146 506 -146 0 net=6769
rlabel metal2 72 -148 72 -148 0 net=4428
rlabel metal2 387 -148 387 -148 0 net=5336
rlabel metal2 79 -150 79 -150 0 net=3450
rlabel metal2 180 -150 180 -150 0 net=231
rlabel metal2 366 -150 366 -150 0 net=5166
rlabel metal2 79 -152 79 -152 0 net=4753
rlabel metal2 138 -152 138 -152 0 net=2789
rlabel metal2 390 -152 390 -152 0 net=1400
rlabel metal2 86 -154 86 -154 0 net=3448
rlabel metal2 247 -154 247 -154 0 net=1395
rlabel metal2 285 -154 285 -154 0 net=2982
rlabel metal2 457 -154 457 -154 0 net=2539
rlabel metal2 86 -156 86 -156 0 net=6905
rlabel metal2 296 -156 296 -156 0 net=5104
rlabel metal2 100 -158 100 -158 0 net=2191
rlabel metal2 173 -158 173 -158 0 net=1237
rlabel metal2 296 -158 296 -158 0 net=3972
rlabel metal2 527 -158 527 -158 0 net=6811
rlabel metal2 107 -160 107 -160 0 net=2349
rlabel metal2 191 -160 191 -160 0 net=1495
rlabel metal2 317 -160 317 -160 0 net=2488
rlabel metal2 331 -160 331 -160 0 net=3536
rlabel metal2 527 -160 527 -160 0 net=5733
rlabel metal2 114 -162 114 -162 0 net=1941
rlabel metal2 341 -162 341 -162 0 net=2699
rlabel metal2 408 -162 408 -162 0 net=3103
rlabel metal2 464 -162 464 -162 0 net=4119
rlabel metal2 114 -164 114 -164 0 net=2257
rlabel metal2 135 -164 135 -164 0 net=661
rlabel metal2 324 -164 324 -164 0 net=4631
rlabel metal2 408 -164 408 -164 0 net=4643
rlabel metal2 443 -164 443 -164 0 net=4147
rlabel metal2 478 -164 478 -164 0 net=5825
rlabel metal2 121 -166 121 -166 0 net=1681
rlabel metal2 177 -166 177 -166 0 net=1281
rlabel metal2 345 -166 345 -166 0 net=2325
rlabel metal2 394 -166 394 -166 0 net=5873
rlabel metal2 492 -166 492 -166 0 net=5541
rlabel metal2 513 -166 513 -166 0 net=5171
rlabel metal2 128 -168 128 -168 0 net=1971
rlabel metal2 338 -168 338 -168 0 net=3727
rlabel metal2 352 -168 352 -168 0 net=5935
rlabel metal2 436 -168 436 -168 0 net=6699
rlabel metal2 149 -170 149 -170 0 net=2864
rlabel metal2 359 -170 359 -170 0 net=6846
rlabel metal2 149 -172 149 -172 0 net=4475
rlabel metal2 362 -172 362 -172 0 net=4059
rlabel metal2 450 -172 450 -172 0 net=5277
rlabel metal2 583 -172 583 -172 0 net=4069
rlabel metal2 156 -174 156 -174 0 net=1667
rlabel metal2 261 -174 261 -174 0 net=1757
rlabel metal2 355 -174 355 -174 0 net=2749
rlabel metal2 163 -176 163 -176 0 net=1263
rlabel metal2 355 -176 355 -176 0 net=5256
rlabel metal2 170 -178 170 -178 0 net=2736
rlabel metal2 275 -178 275 -178 0 net=2171
rlabel metal2 551 -178 551 -178 0 net=5409
rlabel metal2 205 -180 205 -180 0 net=5597
rlabel metal2 226 -182 226 -182 0 net=2129
rlabel metal2 289 -182 289 -182 0 net=2443
rlabel metal2 198 -184 198 -184 0 net=1915
rlabel metal2 233 -184 233 -184 0 net=1411
rlabel metal2 289 -184 289 -184 0 net=1963
rlabel metal2 93 -186 93 -186 0 net=3224
rlabel metal2 93 -188 93 -188 0 net=2453
rlabel metal2 198 -188 198 -188 0 net=1327
rlabel metal2 58 -190 58 -190 0 net=5658
rlabel metal2 215 -190 215 -190 0 net=2013
rlabel metal2 16 -201 16 -201 0 net=1669
rlabel metal2 187 -201 187 -201 0 net=2172
rlabel metal2 303 -201 303 -201 0 net=5701
rlabel metal2 646 -201 646 -201 0 net=6863
rlabel metal2 37 -203 37 -203 0 net=5287
rlabel metal2 198 -203 198 -203 0 net=1328
rlabel metal2 317 -203 317 -203 0 net=2661
rlabel metal2 317 -203 317 -203 0 net=2661
rlabel metal2 320 -203 320 -203 0 net=2750
rlabel metal2 460 -203 460 -203 0 net=6719
rlabel metal2 670 -203 670 -203 0 net=6299
rlabel metal2 44 -205 44 -205 0 net=4379
rlabel metal2 205 -205 205 -205 0 net=6700
rlabel metal2 520 -205 520 -205 0 net=5827
rlabel metal2 65 -207 65 -207 0 net=2906
rlabel metal2 212 -207 212 -207 0 net=2014
rlabel metal2 233 -207 233 -207 0 net=1979
rlabel metal2 411 -207 411 -207 0 net=1025
rlabel metal2 467 -207 467 -207 0 net=5683
rlabel metal2 618 -207 618 -207 0 net=3211
rlabel metal2 65 -209 65 -209 0 net=2101
rlabel metal2 233 -209 233 -209 0 net=1239
rlabel metal2 261 -209 261 -209 0 net=1413
rlabel metal2 289 -209 289 -209 0 net=1965
rlabel metal2 331 -209 331 -209 0 net=1942
rlabel metal2 513 -209 513 -209 0 net=4121
rlabel metal2 562 -209 562 -209 0 net=2541
rlabel metal2 79 -211 79 -211 0 net=4754
rlabel metal2 236 -211 236 -211 0 net=1609
rlabel metal2 355 -211 355 -211 0 net=4765
rlabel metal2 569 -211 569 -211 0 net=4070
rlabel metal2 590 -211 590 -211 0 net=5173
rlabel metal2 51 -213 51 -213 0 net=2199
rlabel metal2 86 -213 86 -213 0 net=6906
rlabel metal2 173 -213 173 -213 0 net=1521
rlabel metal2 359 -213 359 -213 0 net=2327
rlabel metal2 390 -213 390 -213 0 net=5874
rlabel metal2 520 -213 520 -213 0 net=5411
rlabel metal2 569 -213 569 -213 0 net=6629
rlabel metal2 86 -215 86 -215 0 net=4477
rlabel metal2 222 -215 222 -215 0 net=3299
rlabel metal2 397 -215 397 -215 0 net=4148
rlabel metal2 471 -215 471 -215 0 net=4677
rlabel metal2 576 -215 576 -215 0 net=6771
rlabel metal2 93 -217 93 -217 0 net=2455
rlabel metal2 268 -217 268 -217 0 net=2131
rlabel metal2 373 -217 373 -217 0 net=4847
rlabel metal2 93 -219 93 -219 0 net=3195
rlabel metal2 198 -219 198 -219 0 net=2035
rlabel metal2 282 -219 282 -219 0 net=2049
rlabel metal2 376 -219 376 -219 0 net=4378
rlabel metal2 492 -219 492 -219 0 net=5279
rlabel metal2 597 -219 597 -219 0 net=4903
rlabel metal2 100 -221 100 -221 0 net=2193
rlabel metal2 240 -221 240 -221 0 net=1397
rlabel metal2 299 -221 299 -221 0 net=3265
rlabel metal2 527 -221 527 -221 0 net=5735
rlabel metal2 30 -223 30 -223 0 net=5649
rlabel metal2 107 -223 107 -223 0 net=2350
rlabel metal2 226 -223 226 -223 0 net=1917
rlabel metal2 397 -223 397 -223 0 net=2711
rlabel metal2 464 -223 464 -223 0 net=6812
rlabel metal2 544 -223 544 -223 0 net=4857
rlabel metal2 23 -225 23 -225 0 net=6607
rlabel metal2 121 -225 121 -225 0 net=1683
rlabel metal2 177 -225 177 -225 0 net=1283
rlabel metal2 324 -225 324 -225 0 net=4633
rlabel metal2 58 -227 58 -227 0 net=4785
rlabel metal2 310 -227 310 -227 0 net=1759
rlabel metal2 404 -227 404 -227 0 net=750
rlabel metal2 509 -227 509 -227 0 net=4575
rlabel metal2 72 -229 72 -229 0 net=126
rlabel metal2 247 -229 247 -229 0 net=1497
rlabel metal2 408 -229 408 -229 0 net=4645
rlabel metal2 72 -231 72 -231 0 net=2259
rlabel metal2 121 -231 121 -231 0 net=2173
rlabel metal2 163 -231 163 -231 0 net=1265
rlabel metal2 408 -231 408 -231 0 net=5542
rlabel metal2 114 -233 114 -233 0 net=2575
rlabel metal2 415 -233 415 -233 0 net=3105
rlabel metal2 443 -233 443 -233 0 net=4061
rlabel metal2 128 -235 128 -235 0 net=1973
rlabel metal2 366 -235 366 -235 0 net=2791
rlabel metal2 485 -235 485 -235 0 net=3911
rlabel metal2 128 -237 128 -237 0 net=1813
rlabel metal2 208 -237 208 -237 0 net=5353
rlabel metal2 138 -239 138 -239 0 net=1887
rlabel metal2 338 -239 338 -239 0 net=2445
rlabel metal2 422 -239 422 -239 0 net=5599
rlabel metal2 163 -241 163 -241 0 net=2467
rlabel metal2 338 -241 338 -241 0 net=4071
rlabel metal2 345 -243 345 -243 0 net=3728
rlabel metal2 418 -243 418 -243 0 net=3035
rlabel metal2 429 -243 429 -243 0 net=5936
rlabel metal2 345 -245 345 -245 0 net=2701
rlabel metal2 394 -245 394 -245 0 net=3043
rlabel metal2 394 -247 394 -247 0 net=3519
rlabel metal2 23 -258 23 -258 0 net=6608
rlabel metal2 142 -258 142 -258 0 net=2457
rlabel metal2 299 -258 299 -258 0 net=602
rlabel metal2 439 -258 439 -258 0 net=5280
rlabel metal2 583 -258 583 -258 0 net=4859
rlabel metal2 583 -258 583 -258 0 net=4859
rlabel metal2 590 -258 590 -258 0 net=5601
rlabel metal2 597 -258 597 -258 0 net=4905
rlabel metal2 604 -258 604 -258 0 net=3520
rlabel metal2 674 -258 674 -258 0 net=6301
rlabel metal2 751 -258 751 -258 0 net=6631
rlabel metal2 856 -258 856 -258 0 net=6683
rlabel metal2 51 -260 51 -260 0 net=4787
rlabel metal2 65 -260 65 -260 0 net=2102
rlabel metal2 240 -260 240 -260 0 net=1398
rlabel metal2 334 -260 334 -260 0 net=6720
rlabel metal2 681 -260 681 -260 0 net=6773
rlabel metal2 16 -262 16 -262 0 net=1670
rlabel metal2 247 -262 247 -262 0 net=1266
rlabel metal2 401 -262 401 -262 0 net=1980
rlabel metal2 590 -262 590 -262 0 net=5703
rlabel metal2 646 -262 646 -262 0 net=5737
rlabel metal2 688 -262 688 -262 0 net=6865
rlabel metal2 58 -264 58 -264 0 net=2201
rlabel metal2 107 -264 107 -264 0 net=2174
rlabel metal2 128 -264 128 -264 0 net=1513
rlabel metal2 229 -264 229 -264 0 net=1918
rlabel metal2 261 -264 261 -264 0 net=1415
rlabel metal2 338 -264 338 -264 0 net=1974
rlabel metal2 359 -264 359 -264 0 net=2329
rlabel metal2 415 -264 415 -264 0 net=3037
rlabel metal2 443 -264 443 -264 0 net=2793
rlabel metal2 485 -264 485 -264 0 net=3913
rlabel metal2 485 -264 485 -264 0 net=3913
rlabel metal2 492 -264 492 -264 0 net=4063
rlabel metal2 492 -264 492 -264 0 net=4063
rlabel metal2 499 -264 499 -264 0 net=4073
rlabel metal2 534 -264 534 -264 0 net=4635
rlabel metal2 597 -264 597 -264 0 net=5685
rlabel metal2 618 -264 618 -264 0 net=3212
rlabel metal2 688 -264 688 -264 0 net=6085
rlabel metal2 44 -266 44 -266 0 net=4380
rlabel metal2 107 -266 107 -266 0 net=3085
rlabel metal2 191 -266 191 -266 0 net=2051
rlabel metal2 205 -266 205 -266 0 net=1297
rlabel metal2 268 -266 268 -266 0 net=6009
rlabel metal2 359 -266 359 -266 0 net=2207
rlabel metal2 446 -266 446 -266 0 net=5875
rlabel metal2 625 -266 625 -266 0 net=4849
rlabel metal2 68 -268 68 -268 0 net=867
rlabel metal2 114 -268 114 -268 0 net=2576
rlabel metal2 184 -268 184 -268 0 net=2195
rlabel metal2 275 -268 275 -268 0 net=1499
rlabel metal2 341 -268 341 -268 0 net=3165
rlabel metal2 460 -268 460 -268 0 net=6261
rlabel metal2 72 -270 72 -270 0 net=2260
rlabel metal2 149 -270 149 -270 0 net=1685
rlabel metal2 177 -270 177 -270 0 net=1889
rlabel metal2 205 -270 205 -270 0 net=1611
rlabel metal2 310 -270 310 -270 0 net=2663
rlabel metal2 373 -270 373 -270 0 net=2050
rlabel metal2 481 -270 481 -270 0 net=5693
rlabel metal2 37 -272 37 -272 0 net=5288
rlabel metal2 215 -272 215 -272 0 net=1141
rlabel metal2 499 -272 499 -272 0 net=4123
rlabel metal2 520 -272 520 -272 0 net=5413
rlabel metal2 632 -272 632 -272 0 net=5175
rlabel metal2 30 -274 30 -274 0 net=5650
rlabel metal2 222 -274 222 -274 0 net=1284
rlabel metal2 296 -274 296 -274 0 net=1966
rlabel metal2 317 -274 317 -274 0 net=1761
rlabel metal2 373 -274 373 -274 0 net=6901
rlabel metal2 30 -276 30 -276 0 net=4479
rlabel metal2 100 -276 100 -276 0 net=513
rlabel metal2 117 -276 117 -276 0 net=6757
rlabel metal2 639 -276 639 -276 0 net=5829
rlabel metal2 37 -278 37 -278 0 net=3197
rlabel metal2 121 -278 121 -278 0 net=2037
rlabel metal2 282 -278 282 -278 0 net=2133
rlabel metal2 380 -278 380 -278 0 net=3301
rlabel metal2 471 -278 471 -278 0 net=3267
rlabel metal2 541 -278 541 -278 0 net=5355
rlabel metal2 72 -280 72 -280 0 net=2469
rlabel metal2 180 -280 180 -280 0 net=2405
rlabel metal2 243 -280 243 -280 0 net=4335
rlabel metal2 390 -280 390 -280 0 net=66
rlabel metal2 555 -280 555 -280 0 net=4679
rlabel metal2 86 -282 86 -282 0 net=3493
rlabel metal2 394 -282 394 -282 0 net=4193
rlabel metal2 562 -282 562 -282 0 net=4767
rlabel metal2 600 -282 600 -282 0 net=1
rlabel metal2 93 -284 93 -284 0 net=3395
rlabel metal2 289 -284 289 -284 0 net=1523
rlabel metal2 324 -284 324 -284 0 net=2447
rlabel metal2 429 -284 429 -284 0 net=3045
rlabel metal2 527 -284 527 -284 0 net=4577
rlabel metal2 565 -284 565 -284 0 net=5891
rlabel metal2 149 -286 149 -286 0 net=1815
rlabel metal2 345 -286 345 -286 0 net=2703
rlabel metal2 411 -286 411 -286 0 net=4103
rlabel metal2 163 -288 163 -288 0 net=3305
rlabel metal2 170 -290 170 -290 0 net=1241
rlabel metal2 345 -290 345 -290 0 net=4647
rlabel metal2 387 -292 387 -292 0 net=4223
rlabel metal2 387 -294 387 -294 0 net=2543
rlabel metal2 429 -296 429 -296 0 net=3107
rlabel metal2 450 -296 450 -296 0 net=2712
rlabel metal2 422 -298 422 -298 0 net=3087
rlabel metal2 506 -298 506 -298 0 net=6551
rlabel metal2 338 -300 338 -300 0 net=4969
rlabel metal2 2 -311 2 -311 0 net=5949
rlabel metal2 107 -311 107 -311 0 net=3086
rlabel metal2 121 -311 121 -311 0 net=2038
rlabel metal2 128 -311 128 -311 0 net=1514
rlabel metal2 653 -311 653 -311 0 net=5603
rlabel metal2 849 -311 849 -311 0 net=6235
rlabel metal2 9 -313 9 -313 0 net=5691
rlabel metal2 72 -313 72 -313 0 net=2470
rlabel metal2 226 -313 226 -313 0 net=1299
rlabel metal2 226 -313 226 -313 0 net=1299
rlabel metal2 233 -313 233 -313 0 net=4648
rlabel metal2 352 -313 352 -313 0 net=6010
rlabel metal2 590 -313 590 -313 0 net=5705
rlabel metal2 674 -313 674 -313 0 net=6245
rlabel metal2 681 -313 681 -313 0 net=5739
rlabel metal2 726 -313 726 -313 0 net=6785
rlabel metal2 16 -315 16 -315 0 net=5887
rlabel metal2 114 -315 114 -315 0 net=3039
rlabel metal2 422 -315 422 -315 0 net=4064
rlabel metal2 534 -315 534 -315 0 net=4195
rlabel metal2 569 -315 569 -315 0 net=4637
rlabel metal2 695 -315 695 -315 0 net=6553
rlabel metal2 828 -315 828 -315 0 net=6633
rlabel metal2 23 -317 23 -317 0 net=4917
rlabel metal2 215 -317 215 -317 0 net=246
rlabel metal2 257 -317 257 -317 0 net=1416
rlabel metal2 275 -317 275 -317 0 net=1500
rlabel metal2 352 -317 352 -317 0 net=3915
rlabel metal2 513 -317 513 -317 0 net=4075
rlabel metal2 548 -317 548 -317 0 net=4225
rlabel metal2 597 -317 597 -317 0 net=5687
rlabel metal2 702 -317 702 -317 0 net=5893
rlabel metal2 852 -317 852 -317 0 net=6684
rlabel metal2 30 -319 30 -319 0 net=4481
rlabel metal2 96 -319 96 -319 0 net=3717
rlabel metal2 219 -319 219 -319 0 net=3341
rlabel metal2 359 -319 359 -319 0 net=2208
rlabel metal2 450 -319 450 -319 0 net=3089
rlabel metal2 513 -319 513 -319 0 net=3268
rlabel metal2 544 -319 544 -319 0 net=6609
rlabel metal2 709 -319 709 -319 0 net=4851
rlabel metal2 44 -321 44 -321 0 net=972
rlabel metal2 121 -321 121 -321 0 net=4265
rlabel metal2 401 -321 401 -321 0 net=4680
rlabel metal2 667 -321 667 -321 0 net=5695
rlabel metal2 716 -321 716 -321 0 net=6303
rlabel metal2 716 -321 716 -321 0 net=6303
rlabel metal2 730 -321 730 -321 0 net=6263
rlabel metal2 44 -323 44 -323 0 net=4863
rlabel metal2 240 -323 240 -323 0 net=3705
rlabel metal2 450 -323 450 -323 0 net=3047
rlabel metal2 520 -323 520 -323 0 net=4105
rlabel metal2 583 -323 583 -323 0 net=4861
rlabel metal2 618 -323 618 -323 0 net=5357
rlabel metal2 737 -323 737 -323 0 net=6775
rlabel metal2 51 -325 51 -325 0 net=4788
rlabel metal2 362 -325 362 -325 0 net=6229
rlabel metal2 51 -327 51 -327 0 net=1891
rlabel metal2 233 -327 233 -327 0 net=6217
rlabel metal2 37 -329 37 -329 0 net=3199
rlabel metal2 240 -329 240 -329 0 net=2135
rlabel metal2 289 -329 289 -329 0 net=5483
rlabel metal2 744 -329 744 -329 0 net=6867
rlabel metal2 58 -331 58 -331 0 net=2202
rlabel metal2 135 -331 135 -331 0 net=984
rlabel metal2 247 -331 247 -331 0 net=1763
rlabel metal2 334 -331 334 -331 0 net=2330
rlabel metal2 471 -331 471 -331 0 net=2794
rlabel metal2 499 -331 499 -331 0 net=4125
rlabel metal2 583 -331 583 -331 0 net=6758
rlabel metal2 639 -331 639 -331 0 net=5831
rlabel metal2 751 -331 751 -331 0 net=6903
rlabel metal2 58 -333 58 -333 0 net=1817
rlabel metal2 212 -333 212 -333 0 net=3013
rlabel metal2 474 -333 474 -333 0 net=5711
rlabel metal2 639 -333 639 -333 0 net=5481
rlabel metal2 65 -335 65 -335 0 net=2053
rlabel metal2 261 -335 261 -335 0 net=1525
rlabel metal2 310 -335 310 -335 0 net=2665
rlabel metal2 373 -335 373 -335 0 net=5937
rlabel metal2 75 -337 75 -337 0 net=472
rlabel metal2 170 -337 170 -337 0 net=1243
rlabel metal2 282 -337 282 -337 0 net=2449
rlabel metal2 380 -337 380 -337 0 net=4337
rlabel metal2 586 -337 586 -337 0 net=6449
rlabel metal2 86 -339 86 -339 0 net=3495
rlabel metal2 380 -339 380 -339 0 net=2545
rlabel metal2 394 -339 394 -339 0 net=3167
rlabel metal2 506 -339 506 -339 0 net=4971
rlabel metal2 646 -339 646 -339 0 net=5177
rlabel metal2 688 -339 688 -339 0 net=6087
rlabel metal2 86 -341 86 -341 0 net=2197
rlabel metal2 289 -341 289 -341 0 net=2495
rlabel metal2 401 -341 401 -341 0 net=566
rlabel metal2 436 -341 436 -341 0 net=5669
rlabel metal2 93 -343 93 -343 0 net=3397
rlabel metal2 429 -343 429 -343 0 net=3109
rlabel metal2 457 -343 457 -343 0 net=3303
rlabel metal2 516 -343 516 -343 0 net=5987
rlabel metal2 93 -345 93 -345 0 net=6353
rlabel metal2 100 -347 100 -347 0 net=1709
rlabel metal2 429 -347 429 -347 0 net=3955
rlabel metal2 604 -347 604 -347 0 net=5877
rlabel metal2 128 -349 128 -349 0 net=4227
rlabel metal2 254 -349 254 -349 0 net=2783
rlabel metal2 604 -349 604 -349 0 net=4906
rlabel metal2 625 -349 625 -349 0 net=5415
rlabel metal2 138 -351 138 -351 0 net=438
rlabel metal2 296 -351 296 -351 0 net=1873
rlabel metal2 576 -351 576 -351 0 net=4769
rlabel metal2 142 -353 142 -353 0 net=2458
rlabel metal2 555 -353 555 -353 0 net=4579
rlabel metal2 30 -355 30 -355 0 net=4975
rlabel metal2 145 -355 145 -355 0 net=3967
rlabel metal2 156 -357 156 -357 0 net=1687
rlabel metal2 156 -359 156 -359 0 net=3307
rlabel metal2 254 -359 254 -359 0 net=2617
rlabel metal2 331 -359 331 -359 0 net=4601
rlabel metal2 37 -361 37 -361 0 net=2953
rlabel metal2 334 -361 334 -361 0 net=4919
rlabel metal2 163 -363 163 -363 0 net=1613
rlabel metal2 268 -363 268 -363 0 net=1607
rlabel metal2 453 -363 453 -363 0 net=1
rlabel metal2 205 -365 205 -365 0 net=3699
rlabel metal2 299 -367 299 -367 0 net=4213
rlabel metal2 303 -369 303 -369 0 net=2705
rlabel metal2 366 -371 366 -371 0 net=6203
rlabel metal2 2 -382 2 -382 0 net=5950
rlabel metal2 205 -382 205 -382 0 net=6621
rlabel metal2 2 -384 2 -384 0 net=4707
rlabel metal2 226 -384 226 -384 0 net=1301
rlabel metal2 226 -384 226 -384 0 net=1301
rlabel metal2 261 -384 261 -384 0 net=1526
rlabel metal2 369 -384 369 -384 0 net=4076
rlabel metal2 621 -384 621 -384 0 net=5482
rlabel metal2 660 -384 660 -384 0 net=5359
rlabel metal2 660 -384 660 -384 0 net=5359
rlabel metal2 758 -384 758 -384 0 net=4853
rlabel metal2 758 -384 758 -384 0 net=4853
rlabel metal2 828 -384 828 -384 0 net=6265
rlabel metal2 16 -386 16 -386 0 net=5888
rlabel metal2 159 -386 159 -386 0 net=6373
rlabel metal2 16 -388 16 -388 0 net=4865
rlabel metal2 51 -388 51 -388 0 net=1892
rlabel metal2 261 -388 261 -388 0 net=2471
rlabel metal2 478 -388 478 -388 0 net=3090
rlabel metal2 516 -388 516 -388 0 net=5878
rlabel metal2 842 -388 842 -388 0 net=6355
rlabel metal2 23 -390 23 -390 0 net=4918
rlabel metal2 275 -390 275 -390 0 net=2351
rlabel metal2 436 -390 436 -390 0 net=3111
rlabel metal2 502 -390 502 -390 0 net=6776
rlabel metal2 852 -390 852 -390 0 net=6634
rlabel metal2 23 -392 23 -392 0 net=3719
rlabel metal2 282 -392 282 -392 0 net=2450
rlabel metal2 390 -392 390 -392 0 net=6554
rlabel metal2 807 -392 807 -392 0 net=6701
rlabel metal2 863 -392 863 -392 0 net=6236
rlabel metal2 37 -394 37 -394 0 net=2954
rlabel metal2 509 -394 509 -394 0 net=6803
rlabel metal2 37 -396 37 -396 0 net=3185
rlabel metal2 107 -396 107 -396 0 net=792
rlabel metal2 310 -396 310 -396 0 net=3398
rlabel metal2 359 -396 359 -396 0 net=5706
rlabel metal2 716 -396 716 -396 0 net=6305
rlabel metal2 44 -398 44 -398 0 net=2039
rlabel metal2 184 -398 184 -398 0 net=3201
rlabel metal2 303 -398 303 -398 0 net=2707
rlabel metal2 317 -398 317 -398 0 net=3497
rlabel metal2 495 -398 495 -398 0 net=6721
rlabel metal2 54 -400 54 -400 0 net=1114
rlabel metal2 145 -400 145 -400 0 net=5757
rlabel metal2 870 -400 870 -400 0 net=6787
rlabel metal2 75 -402 75 -402 0 net=1608
rlabel metal2 303 -402 303 -402 0 net=6904
rlabel metal2 79 -404 79 -404 0 net=4482
rlabel metal2 100 -404 100 -404 0 net=1711
rlabel metal2 201 -404 201 -404 0 net=4941
rlabel metal2 324 -404 324 -404 0 net=3169
rlabel metal2 401 -404 401 -404 0 net=3304
rlabel metal2 520 -404 520 -404 0 net=4107
rlabel metal2 604 -404 604 -404 0 net=5609
rlabel metal2 674 -404 674 -404 0 net=6247
rlabel metal2 9 -406 9 -406 0 net=5692
rlabel metal2 86 -406 86 -406 0 net=2198
rlabel metal2 240 -406 240 -406 0 net=2137
rlabel metal2 373 -406 373 -406 0 net=6405
rlabel metal2 9 -408 9 -408 0 net=4229
rlabel metal2 240 -408 240 -408 0 net=2341
rlabel metal2 331 -408 331 -408 0 net=3916
rlabel metal2 408 -408 408 -408 0 net=3014
rlabel metal2 520 -408 520 -408 0 net=6088
rlabel metal2 772 -408 772 -408 0 net=6205
rlabel metal2 72 -410 72 -410 0 net=1287
rlabel metal2 369 -410 369 -410 0 net=2957
rlabel metal2 415 -410 415 -410 0 net=3701
rlabel metal2 555 -410 555 -410 0 net=4603
rlabel metal2 695 -410 695 -410 0 net=5689
rlabel metal2 814 -410 814 -410 0 net=5895
rlabel metal2 72 -412 72 -412 0 net=1615
rlabel metal2 170 -412 170 -412 0 net=1689
rlabel metal2 212 -412 212 -412 0 net=5039
rlabel metal2 86 -414 86 -414 0 net=3309
rlabel metal2 163 -414 163 -414 0 net=4226
rlabel metal2 576 -414 576 -414 0 net=4581
rlabel metal2 625 -414 625 -414 0 net=4921
rlabel metal2 716 -414 716 -414 0 net=6231
rlabel metal2 93 -416 93 -416 0 net=1765
rlabel metal2 254 -416 254 -416 0 net=2619
rlabel metal2 422 -416 422 -416 0 net=6517
rlabel metal2 65 -418 65 -418 0 net=2055
rlabel metal2 289 -418 289 -418 0 net=2497
rlabel metal2 422 -418 422 -418 0 net=5485
rlabel metal2 730 -418 730 -418 0 net=5833
rlabel metal2 58 -420 58 -420 0 net=1819
rlabel metal2 107 -420 107 -420 0 net=731
rlabel metal2 425 -420 425 -420 0 net=4862
rlabel metal2 611 -420 611 -420 0 net=4771
rlabel metal2 646 -420 646 -420 0 net=5417
rlabel metal2 730 -420 730 -420 0 net=5939
rlabel metal2 58 -422 58 -422 0 net=1875
rlabel metal2 338 -422 338 -422 0 net=2667
rlabel metal2 110 -424 110 -424 0 net=2939
rlabel metal2 289 -424 289 -424 0 net=2547
rlabel metal2 436 -424 436 -424 0 net=5604
rlabel metal2 117 -426 117 -426 0 net=97
rlabel metal2 450 -426 450 -426 0 net=3048
rlabel metal2 471 -426 471 -426 0 net=6281
rlabel metal2 835 -426 835 -426 0 net=6451
rlabel metal2 114 -428 114 -428 0 net=3041
rlabel metal2 485 -428 485 -428 0 net=3969
rlabel metal2 590 -428 590 -428 0 net=4639
rlabel metal2 688 -428 688 -428 0 net=5671
rlabel metal2 114 -430 114 -430 0 net=4271
rlabel metal2 632 -430 632 -430 0 net=4973
rlabel metal2 121 -432 121 -432 0 net=4267
rlabel metal2 418 -432 418 -432 0 net=3459
rlabel metal2 523 -432 523 -432 0 net=6737
rlabel metal2 121 -434 121 -434 0 net=2971
rlabel metal2 156 -434 156 -434 0 net=1088
rlabel metal2 345 -434 345 -434 0 net=3343
rlabel metal2 527 -434 527 -434 0 net=4127
rlabel metal2 646 -434 646 -434 0 net=5179
rlabel metal2 688 -434 688 -434 0 net=5697
rlabel metal2 751 -434 751 -434 0 net=6869
rlabel metal2 30 -436 30 -436 0 net=4976
rlabel metal2 212 -436 212 -436 0 net=6731
rlabel metal2 30 -438 30 -438 0 net=3543
rlabel metal2 135 -438 135 -438 0 net=1859
rlabel metal2 366 -438 366 -438 0 net=4507
rlabel metal2 618 -438 618 -438 0 net=5713
rlabel metal2 128 -440 128 -440 0 net=1245
rlabel metal2 233 -440 233 -440 0 net=1927
rlabel metal2 548 -440 548 -440 0 net=4339
rlabel metal2 667 -440 667 -440 0 net=5989
rlabel metal2 142 -442 142 -442 0 net=2737
rlabel metal2 191 -442 191 -442 0 net=1995
rlabel metal2 404 -442 404 -442 0 net=3551
rlabel metal2 555 -442 555 -442 0 net=4197
rlabel metal2 611 -442 611 -442 0 net=5743
rlabel metal2 702 -442 702 -442 0 net=6611
rlabel metal2 142 -444 142 -444 0 net=2583
rlabel metal2 443 -444 443 -444 0 net=3707
rlabel metal2 702 -444 702 -444 0 net=6219
rlabel metal2 152 -446 152 -446 0 net=1435
rlabel metal2 296 -448 296 -448 0 net=6193
rlabel metal2 331 -450 331 -450 0 net=2311
rlabel metal2 541 -450 541 -450 0 net=4215
rlabel metal2 723 -450 723 -450 0 net=5741
rlabel metal2 299 -452 299 -452 0 net=5079
rlabel metal2 387 -454 387 -454 0 net=2785
rlabel metal2 499 -454 499 -454 0 net=3957
rlabel metal2 278 -456 278 -456 0 net=950
rlabel metal2 387 -458 387 -458 0 net=2408
rlabel metal2 415 -460 415 -460 0 net=1863
rlabel metal2 2 -471 2 -471 0 net=4708
rlabel metal2 268 -471 268 -471 0 net=4942
rlabel metal2 429 -471 429 -471 0 net=5834
rlabel metal2 2 -473 2 -473 0 net=6555
rlabel metal2 243 -473 243 -473 0 net=3344
rlabel metal2 544 -473 544 -473 0 net=6306
rlabel metal2 9 -475 9 -475 0 net=4230
rlabel metal2 607 -475 607 -475 0 net=6189
rlabel metal2 716 -475 716 -475 0 net=6233
rlabel metal2 716 -475 716 -475 0 net=6233
rlabel metal2 726 -475 726 -475 0 net=5896
rlabel metal2 9 -477 9 -477 0 net=6691
rlabel metal2 51 -477 51 -477 0 net=496
rlabel metal2 170 -477 170 -477 0 net=2739
rlabel metal2 170 -477 170 -477 0 net=2739
rlabel metal2 180 -477 180 -477 0 net=1093
rlabel metal2 212 -477 212 -477 0 net=6622
rlabel metal2 30 -479 30 -479 0 net=3545
rlabel metal2 54 -479 54 -479 0 net=4922
rlabel metal2 807 -479 807 -479 0 net=6703
rlabel metal2 807 -479 807 -479 0 net=6703
rlabel metal2 814 -479 814 -479 0 net=6739
rlabel metal2 30 -481 30 -481 0 net=3187
rlabel metal2 58 -481 58 -481 0 net=1876
rlabel metal2 313 -481 313 -481 0 net=2668
rlabel metal2 37 -483 37 -483 0 net=3795
rlabel metal2 394 -483 394 -483 0 net=2498
rlabel metal2 439 -483 439 -483 0 net=817
rlabel metal2 58 -485 58 -485 0 net=1861
rlabel metal2 184 -485 184 -485 0 net=1713
rlabel metal2 243 -485 243 -485 0 net=3202
rlabel metal2 303 -485 303 -485 0 net=2343
rlabel metal2 320 -485 320 -485 0 net=3708
rlabel metal2 695 -485 695 -485 0 net=6221
rlabel metal2 79 -487 79 -487 0 net=333
rlabel metal2 100 -487 100 -487 0 net=4604
rlabel metal2 660 -487 660 -487 0 net=5361
rlabel metal2 23 -489 23 -489 0 net=3721
rlabel metal2 86 -489 86 -489 0 net=3310
rlabel metal2 324 -489 324 -489 0 net=3171
rlabel metal2 401 -489 401 -489 0 net=4269
rlabel metal2 86 -491 86 -491 0 net=2941
rlabel metal2 352 -491 352 -491 0 net=1288
rlabel metal2 443 -491 443 -491 0 net=2787
rlabel metal2 443 -491 443 -491 0 net=2787
rlabel metal2 460 -491 460 -491 0 net=5672
rlabel metal2 100 -493 100 -493 0 net=1527
rlabel metal2 114 -493 114 -493 0 net=2669
rlabel metal2 408 -493 408 -493 0 net=2959
rlabel metal2 464 -493 464 -493 0 net=1864
rlabel metal2 541 -493 541 -493 0 net=3959
rlabel metal2 639 -493 639 -493 0 net=5611
rlabel metal2 765 -493 765 -493 0 net=6453
rlabel metal2 82 -495 82 -495 0 net=1491
rlabel metal2 117 -495 117 -495 0 net=4640
rlabel metal2 835 -495 835 -495 0 net=6519
rlabel metal2 121 -497 121 -497 0 net=2973
rlabel metal2 415 -497 415 -497 0 net=5742
rlabel metal2 121 -499 121 -499 0 net=2477
rlabel metal2 359 -499 359 -499 0 net=2138
rlabel metal2 373 -499 373 -499 0 net=2621
rlabel metal2 415 -499 415 -499 0 net=3970
rlabel metal2 639 -499 639 -499 0 net=5991
rlabel metal2 674 -499 674 -499 0 net=5699
rlabel metal2 128 -501 128 -501 0 net=1246
rlabel metal2 324 -501 324 -501 0 net=4017
rlabel metal2 576 -501 576 -501 0 net=4583
rlabel metal2 646 -501 646 -501 0 net=5181
rlabel metal2 667 -501 667 -501 0 net=4527
rlabel metal2 16 -503 16 -503 0 net=4867
rlabel metal2 135 -503 135 -503 0 net=2709
rlabel metal2 366 -503 366 -503 0 net=3042
rlabel metal2 485 -503 485 -503 0 net=5040
rlabel metal2 16 -505 16 -505 0 net=6505
rlabel metal2 166 -505 166 -505 0 net=6391
rlabel metal2 488 -505 488 -505 0 net=6248
rlabel metal2 142 -507 142 -507 0 net=2585
rlabel metal2 373 -507 373 -507 0 net=3703
rlabel metal2 646 -507 646 -507 0 net=6206
rlabel metal2 149 -509 149 -509 0 net=662
rlabel metal2 177 -509 177 -509 0 net=2041
rlabel metal2 296 -509 296 -509 0 net=1211
rlabel metal2 338 -509 338 -509 0 net=1997
rlabel metal2 380 -509 380 -509 0 net=4340
rlabel metal2 688 -509 688 -509 0 net=6195
rlabel metal2 779 -509 779 -509 0 net=6723
rlabel metal2 65 -511 65 -511 0 net=1821
rlabel metal2 156 -511 156 -511 0 net=6313
rlabel metal2 502 -511 502 -511 0 net=6356
rlabel metal2 65 -513 65 -513 0 net=3807
rlabel metal2 464 -513 464 -513 0 net=4799
rlabel metal2 506 -513 506 -513 0 net=5714
rlabel metal2 163 -515 163 -515 0 net=5486
rlabel metal2 509 -515 509 -515 0 net=4974
rlabel metal2 184 -517 184 -517 0 net=1303
rlabel metal2 247 -517 247 -517 0 net=2365
rlabel metal2 422 -517 422 -517 0 net=4108
rlabel metal2 632 -517 632 -517 0 net=5419
rlabel metal2 709 -517 709 -517 0 net=6613
rlabel metal2 786 -517 786 -517 0 net=6805
rlabel metal2 191 -519 191 -519 0 net=5690
rlabel metal2 856 -519 856 -519 0 net=6789
rlabel metal2 93 -521 93 -521 0 net=1767
rlabel metal2 194 -521 194 -521 0 net=794
rlabel metal2 254 -521 254 -521 0 net=2057
rlabel metal2 387 -521 387 -521 0 net=4128
rlabel metal2 709 -521 709 -521 0 net=6283
rlabel metal2 93 -523 93 -523 0 net=1094
rlabel metal2 341 -523 341 -523 0 net=5207
rlabel metal2 569 -523 569 -523 0 net=4273
rlabel metal2 590 -523 590 -523 0 net=4509
rlabel metal2 751 -523 751 -523 0 net=6871
rlabel metal2 800 -523 800 -523 0 net=6733
rlabel metal2 198 -525 198 -525 0 net=1929
rlabel metal2 240 -525 240 -525 0 net=6374
rlabel metal2 226 -527 226 -527 0 net=3499
rlabel metal2 513 -527 513 -527 0 net=3553
rlabel metal2 597 -527 597 -527 0 net=4773
rlabel metal2 233 -529 233 -529 0 net=1733
rlabel metal2 520 -529 520 -529 0 net=1436
rlabel metal2 254 -531 254 -531 0 net=2353
rlabel metal2 289 -531 289 -531 0 net=2549
rlabel metal2 436 -531 436 -531 0 net=4951
rlabel metal2 611 -531 611 -531 0 net=5745
rlabel metal2 744 -531 744 -531 0 net=4855
rlabel metal2 205 -533 205 -533 0 net=1691
rlabel metal2 289 -533 289 -533 0 net=2313
rlabel metal2 453 -533 453 -533 0 net=4777
rlabel metal2 730 -533 730 -533 0 net=5941
rlabel metal2 72 -535 72 -535 0 net=1616
rlabel metal2 268 -535 268 -535 0 net=2021
rlabel metal2 457 -535 457 -535 0 net=6877
rlabel metal2 730 -535 730 -535 0 net=6407
rlabel metal2 72 -537 72 -537 0 net=3461
rlabel metal2 457 -537 457 -537 0 net=3113
rlabel metal2 499 -537 499 -537 0 net=5758
rlabel metal2 450 -539 450 -539 0 net=896
rlabel metal2 527 -539 527 -539 0 net=4217
rlabel metal2 478 -541 478 -541 0 net=5080
rlabel metal2 555 -543 555 -543 0 net=4199
rlabel metal2 723 -543 723 -543 0 net=6266
rlabel metal2 261 -545 261 -545 0 net=2473
rlabel metal2 261 -547 261 -547 0 net=2745
rlabel metal2 2 -558 2 -558 0 net=6556
rlabel metal2 502 -558 502 -558 0 net=4584
rlabel metal2 583 -558 583 -558 0 net=4275
rlabel metal2 607 -558 607 -558 0 net=5746
rlabel metal2 681 -558 681 -558 0 net=6879
rlabel metal2 2 -560 2 -560 0 net=3189
rlabel metal2 37 -560 37 -560 0 net=3796
rlabel metal2 107 -560 107 -560 0 net=1493
rlabel metal2 107 -560 107 -560 0 net=1493
rlabel metal2 131 -560 131 -560 0 net=2361
rlabel metal2 177 -560 177 -560 0 net=730
rlabel metal2 345 -560 345 -560 0 net=2058
rlabel metal2 373 -560 373 -560 0 net=3704
rlabel metal2 506 -560 506 -560 0 net=4743
rlabel metal2 541 -560 541 -560 0 net=6645
rlabel metal2 835 -560 835 -560 0 net=6521
rlabel metal2 9 -562 9 -562 0 net=6692
rlabel metal2 135 -562 135 -562 0 net=2710
rlabel metal2 373 -562 373 -562 0 net=2623
rlabel metal2 404 -562 404 -562 0 net=6847
rlabel metal2 9 -564 9 -564 0 net=2943
rlabel metal2 156 -564 156 -564 0 net=4555
rlabel metal2 254 -564 254 -564 0 net=2355
rlabel metal2 254 -564 254 -564 0 net=2355
rlabel metal2 317 -564 317 -564 0 net=1919
rlabel metal2 544 -564 544 -564 0 net=2921
rlabel metal2 23 -566 23 -566 0 net=500
rlabel metal2 191 -566 191 -566 0 net=1768
rlabel metal2 401 -566 401 -566 0 net=3151
rlabel metal2 520 -566 520 -566 0 net=4445
rlabel metal2 646 -566 646 -566 0 net=6655
rlabel metal2 23 -568 23 -568 0 net=3547
rlabel metal2 58 -568 58 -568 0 net=1862
rlabel metal2 415 -568 415 -568 0 net=2559
rlabel metal2 453 -568 453 -568 0 net=4218
rlabel metal2 555 -568 555 -568 0 net=2474
rlabel metal2 744 -568 744 -568 0 net=4856
rlabel metal2 754 -568 754 -568 0 net=3679
rlabel metal2 30 -570 30 -570 0 net=2533
rlabel metal2 436 -570 436 -570 0 net=2746
rlabel metal2 562 -570 562 -570 0 net=4201
rlabel metal2 583 -570 583 -570 0 net=4775
rlabel metal2 660 -570 660 -570 0 net=5613
rlabel metal2 695 -570 695 -570 0 net=6223
rlabel metal2 765 -570 765 -570 0 net=6455
rlabel metal2 40 -572 40 -572 0 net=215
rlabel metal2 429 -572 429 -572 0 net=2961
rlabel metal2 457 -572 457 -572 0 net=3115
rlabel metal2 597 -572 597 -572 0 net=6196
rlabel metal2 723 -572 723 -572 0 net=5393
rlabel metal2 44 -574 44 -574 0 net=4023
rlabel metal2 103 -574 103 -574 0 net=1319
rlabel metal2 348 -574 348 -574 0 net=3819
rlabel metal2 457 -574 457 -574 0 net=3555
rlabel metal2 548 -574 548 -574 0 net=3961
rlabel metal2 618 -574 618 -574 0 net=6191
rlabel metal2 744 -574 744 -574 0 net=5943
rlabel metal2 772 -574 772 -574 0 net=6873
rlabel metal2 51 -576 51 -576 0 net=2479
rlabel metal2 128 -576 128 -576 0 net=4869
rlabel metal2 653 -576 653 -576 0 net=5183
rlabel metal2 698 -576 698 -576 0 net=6307
rlabel metal2 786 -576 786 -576 0 net=6807
rlabel metal2 65 -578 65 -578 0 net=3809
rlabel metal2 79 -578 79 -578 0 net=3722
rlabel metal2 474 -578 474 -578 0 net=5420
rlabel metal2 702 -578 702 -578 0 net=5363
rlabel metal2 793 -578 793 -578 0 net=6790
rlabel metal2 65 -580 65 -580 0 net=1553
rlabel metal2 338 -580 338 -580 0 net=6357
rlabel metal2 800 -580 800 -580 0 net=6735
rlabel metal2 79 -582 79 -582 0 net=1305
rlabel metal2 191 -582 191 -582 0 net=2713
rlabel metal2 485 -582 485 -582 0 net=6393
rlabel metal2 779 -582 779 -582 0 net=6725
rlabel metal2 93 -584 93 -584 0 net=6429
rlabel metal2 800 -584 800 -584 0 net=6705
rlabel metal2 814 -584 814 -584 0 net=6741
rlabel metal2 93 -586 93 -586 0 net=1529
rlabel metal2 135 -586 135 -586 0 net=5951
rlabel metal2 730 -586 730 -586 0 net=6409
rlabel metal2 159 -588 159 -588 0 net=102
rlabel metal2 264 -588 264 -588 0 net=5623
rlabel metal2 737 -588 737 -588 0 net=6615
rlabel metal2 166 -590 166 -590 0 net=4803
rlabel metal2 173 -592 173 -592 0 net=2165
rlabel metal2 184 -592 184 -592 0 net=1931
rlabel metal2 205 -592 205 -592 0 net=6751
rlabel metal2 198 -594 198 -594 0 net=1213
rlabel metal2 313 -594 313 -594 0 net=2788
rlabel metal2 471 -594 471 -594 0 net=6315
rlabel metal2 205 -596 205 -596 0 net=1715
rlabel metal2 226 -596 226 -596 0 net=3501
rlabel metal2 534 -596 534 -596 0 net=5209
rlabel metal2 212 -598 212 -598 0 net=2042
rlabel metal2 289 -598 289 -598 0 net=2315
rlabel metal2 471 -598 471 -598 0 net=4510
rlabel metal2 632 -598 632 -598 0 net=4529
rlabel metal2 16 -600 16 -600 0 net=6506
rlabel metal2 215 -600 215 -600 0 net=357
rlabel metal2 359 -600 359 -600 0 net=4615
rlabel metal2 513 -600 513 -600 0 net=3117
rlabel metal2 569 -600 569 -600 0 net=4953
rlabel metal2 16 -602 16 -602 0 net=3921
rlabel metal2 219 -602 219 -602 0 net=1735
rlabel metal2 236 -602 236 -602 0 net=754
rlabel metal2 425 -602 425 -602 0 net=3621
rlabel metal2 114 -604 114 -604 0 net=2671
rlabel metal2 590 -604 590 -604 0 net=5700
rlabel metal2 114 -606 114 -606 0 net=2741
rlabel metal2 226 -606 226 -606 0 net=2022
rlabel metal2 275 -606 275 -606 0 net=1693
rlabel metal2 359 -606 359 -606 0 net=1999
rlabel metal2 380 -606 380 -606 0 net=2551
rlabel metal2 639 -606 639 -606 0 net=5993
rlabel metal2 149 -608 149 -608 0 net=1822
rlabel metal2 247 -608 247 -608 0 net=2367
rlabel metal2 275 -608 275 -608 0 net=2759
rlabel metal2 611 -608 611 -608 0 net=4779
rlabel metal2 149 -610 149 -610 0 net=4019
rlabel metal2 338 -610 338 -610 0 net=2499
rlabel metal2 467 -610 467 -610 0 net=4083
rlabel metal2 611 -610 611 -610 0 net=6234
rlabel metal2 145 -612 145 -612 0 net=2381
rlabel metal2 366 -612 366 -612 0 net=3173
rlabel metal2 492 -612 492 -612 0 net=5553
rlabel metal2 709 -612 709 -612 0 net=6285
rlabel metal2 247 -614 247 -614 0 net=1485
rlabel metal2 450 -614 450 -614 0 net=5119
rlabel metal2 72 -616 72 -616 0 net=3463
rlabel metal2 72 -618 72 -618 0 net=3067
rlabel metal2 334 -618 334 -618 0 net=3311
rlabel metal2 282 -620 282 -620 0 net=2345
rlabel metal2 352 -620 352 -620 0 net=2587
rlabel metal2 289 -622 289 -622 0 net=2975
rlabel metal2 352 -626 352 -626 0 net=4801
rlabel metal2 464 -628 464 -628 0 net=4270
rlabel metal2 593 -630 593 -630 0 net=5631
rlabel metal2 2 -641 2 -641 0 net=3190
rlabel metal2 61 -641 61 -641 0 net=451
rlabel metal2 138 -641 138 -641 0 net=170
rlabel metal2 464 -641 464 -641 0 net=6192
rlabel metal2 821 -641 821 -641 0 net=5633
rlabel metal2 2 -643 2 -643 0 net=4557
rlabel metal2 173 -643 173 -643 0 net=2346
rlabel metal2 289 -643 289 -643 0 net=2976
rlabel metal2 331 -643 331 -643 0 net=2552
rlabel metal2 590 -643 590 -643 0 net=6736
rlabel metal2 947 -643 947 -643 0 net=5395
rlabel metal2 16 -645 16 -645 0 net=3922
rlabel metal2 93 -645 93 -645 0 net=1530
rlabel metal2 184 -645 184 -645 0 net=1932
rlabel metal2 436 -645 436 -645 0 net=2963
rlabel metal2 488 -645 488 -645 0 net=4776
rlabel metal2 593 -645 593 -645 0 net=2922
rlabel metal2 16 -647 16 -647 0 net=4021
rlabel metal2 184 -647 184 -647 0 net=2369
rlabel metal2 289 -647 289 -647 0 net=2589
rlabel metal2 404 -647 404 -647 0 net=3116
rlabel metal2 562 -647 562 -647 0 net=3963
rlabel metal2 583 -647 583 -647 0 net=4531
rlabel metal2 660 -647 660 -647 0 net=5185
rlabel metal2 793 -647 793 -647 0 net=6431
rlabel metal2 891 -647 891 -647 0 net=6875
rlabel metal2 37 -649 37 -649 0 net=3741
rlabel metal2 338 -649 338 -649 0 net=3174
rlabel metal2 387 -649 387 -649 0 net=3465
rlabel metal2 481 -649 481 -649 0 net=753
rlabel metal2 604 -649 604 -649 0 net=4277
rlabel metal2 621 -649 621 -649 0 net=5364
rlabel metal2 786 -649 786 -649 0 net=6359
rlabel metal2 814 -649 814 -649 0 net=6617
rlabel metal2 51 -651 51 -651 0 net=2480
rlabel metal2 502 -651 502 -651 0 net=6410
rlabel metal2 828 -651 828 -651 0 net=6647
rlabel metal2 30 -653 30 -653 0 net=2534
rlabel metal2 513 -653 513 -653 0 net=3119
rlabel metal2 537 -653 537 -653 0 net=6394
rlabel metal2 779 -653 779 -653 0 net=6317
rlabel metal2 51 -655 51 -655 0 net=3153
rlabel metal2 520 -655 520 -655 0 net=6808
rlabel metal2 58 -657 58 -657 0 net=2167
rlabel metal2 198 -657 198 -657 0 net=1215
rlabel metal2 338 -657 338 -657 0 net=1575
rlabel metal2 506 -657 506 -657 0 net=4745
rlabel metal2 523 -657 523 -657 0 net=585
rlabel metal2 611 -657 611 -657 0 net=6539
rlabel metal2 912 -657 912 -657 0 net=3681
rlabel metal2 65 -659 65 -659 0 net=1555
rlabel metal2 177 -659 177 -659 0 net=2761
rlabel metal2 341 -659 341 -659 0 net=2624
rlabel metal2 436 -659 436 -659 0 net=2643
rlabel metal2 551 -659 551 -659 0 net=5994
rlabel metal2 716 -659 716 -659 0 net=6287
rlabel metal2 65 -661 65 -661 0 net=4097
rlabel metal2 149 -661 149 -661 0 net=2715
rlabel metal2 198 -661 198 -661 0 net=1737
rlabel metal2 233 -661 233 -661 0 net=1921
rlabel metal2 345 -661 345 -661 0 net=3502
rlabel metal2 541 -661 541 -661 0 net=5120
rlabel metal2 730 -661 730 -661 0 net=5625
rlabel metal2 72 -663 72 -663 0 net=3069
rlabel metal2 359 -663 359 -663 0 net=2000
rlabel metal2 408 -663 408 -663 0 net=3811
rlabel metal2 541 -663 541 -663 0 net=6726
rlabel metal2 72 -665 72 -665 0 net=2317
rlabel metal2 474 -665 474 -665 0 net=6665
rlabel metal2 79 -667 79 -667 0 net=1306
rlabel metal2 247 -667 247 -667 0 net=1487
rlabel metal2 366 -667 366 -667 0 net=1285
rlabel metal2 443 -667 443 -667 0 net=2685
rlabel metal2 499 -667 499 -667 0 net=4085
rlabel metal2 555 -667 555 -667 0 net=4954
rlabel metal2 765 -667 765 -667 0 net=6657
rlabel metal2 9 -669 9 -669 0 net=2944
rlabel metal2 250 -669 250 -669 0 net=2356
rlabel metal2 275 -669 275 -669 0 net=2560
rlabel metal2 478 -669 478 -669 0 net=5093
rlabel metal2 9 -671 9 -671 0 net=4025
rlabel metal2 79 -671 79 -671 0 net=2501
rlabel metal2 390 -671 390 -671 0 net=6475
rlabel metal2 23 -673 23 -673 0 net=3549
rlabel metal2 86 -673 86 -673 0 net=6587
rlabel metal2 93 -675 93 -675 0 net=1957
rlabel metal2 170 -675 170 -675 0 net=1233
rlabel metal2 205 -675 205 -675 0 net=1717
rlabel metal2 324 -675 324 -675 0 net=2383
rlabel metal2 562 -675 562 -675 0 net=6456
rlabel metal2 100 -677 100 -677 0 net=4870
rlabel metal2 576 -677 576 -677 0 net=4203
rlabel metal2 614 -677 614 -677 0 net=1072
rlabel metal2 103 -679 103 -679 0 net=4209
rlabel metal2 625 -679 625 -679 0 net=4447
rlabel metal2 639 -679 639 -679 0 net=4781
rlabel metal2 667 -679 667 -679 0 net=3623
rlabel metal2 100 -681 100 -681 0 net=5889
rlabel metal2 674 -681 674 -681 0 net=5555
rlabel metal2 730 -681 730 -681 0 net=6707
rlabel metal2 842 -681 842 -681 0 net=6523
rlabel metal2 103 -683 103 -683 0 net=685
rlabel metal2 170 -683 170 -683 0 net=1321
rlabel metal2 324 -683 324 -683 0 net=3821
rlabel metal2 576 -683 576 -683 0 net=4053
rlabel metal2 639 -683 639 -683 0 net=4469
rlabel metal2 107 -685 107 -685 0 net=1494
rlabel metal2 205 -685 205 -685 0 net=1877
rlabel metal2 261 -685 261 -685 0 net=1247
rlabel metal2 352 -685 352 -685 0 net=4802
rlabel metal2 422 -685 422 -685 0 net=2673
rlabel metal2 646 -685 646 -685 0 net=4805
rlabel metal2 688 -685 688 -685 0 net=5953
rlabel metal2 772 -685 772 -685 0 net=6309
rlabel metal2 842 -685 842 -685 0 net=6753
rlabel metal2 114 -687 114 -687 0 net=2743
rlabel metal2 352 -687 352 -687 0 net=2523
rlabel metal2 653 -687 653 -687 0 net=5211
rlabel metal2 751 -687 751 -687 0 net=6225
rlabel metal2 877 -687 877 -687 0 net=6881
rlabel metal2 89 -689 89 -689 0 net=1325
rlabel metal2 121 -689 121 -689 0 net=2363
rlabel metal2 212 -689 212 -689 0 net=5421
rlabel metal2 744 -689 744 -689 0 net=5945
rlabel metal2 863 -689 863 -689 0 net=6743
rlabel metal2 135 -691 135 -691 0 net=1617
rlabel metal2 219 -691 219 -691 0 net=1695
rlabel metal2 380 -691 380 -691 0 net=3557
rlabel metal2 485 -691 485 -691 0 net=4617
rlabel metal2 681 -691 681 -691 0 net=5615
rlabel metal2 863 -691 863 -691 0 net=6849
rlabel metal2 145 -693 145 -693 0 net=5381
rlabel metal2 163 -695 163 -695 0 net=1839
rlabel metal2 226 -697 226 -697 0 net=347
rlabel metal2 422 -697 422 -697 0 net=2103
rlabel metal2 558 -697 558 -697 0 net=4999
rlabel metal2 229 -699 229 -699 0 net=3503
rlabel metal2 485 -699 485 -699 0 net=5457
rlabel metal2 236 -701 236 -701 0 net=5429
rlabel metal2 240 -703 240 -703 0 net=2331
rlabel metal2 492 -703 492 -703 0 net=3313
rlabel metal2 240 -705 240 -705 0 net=6433
rlabel metal2 296 -707 296 -707 0 net=2807
rlabel metal2 348 -709 348 -709 0 net=3033
rlabel metal2 16 -720 16 -720 0 net=4022
rlabel metal2 135 -720 135 -720 0 net=1618
rlabel metal2 415 -720 415 -720 0 net=6658
rlabel metal2 849 -720 849 -720 0 net=6525
rlabel metal2 908 -720 908 -720 0 net=3682
rlabel metal2 926 -720 926 -720 0 net=5627
rlabel metal2 1006 -720 1006 -720 0 net=6333
rlabel metal2 1031 -720 1031 -720 0 net=5397
rlabel metal2 23 -722 23 -722 0 net=5673
rlabel metal2 135 -722 135 -722 0 net=2717
rlabel metal2 170 -722 170 -722 0 net=1322
rlabel metal2 478 -722 478 -722 0 net=309
rlabel metal2 551 -722 551 -722 0 net=6588
rlabel metal2 912 -722 912 -722 0 net=2071
rlabel metal2 26 -724 26 -724 0 net=1158
rlabel metal2 33 -724 33 -724 0 net=284
rlabel metal2 716 -724 716 -724 0 net=5459
rlabel metal2 793 -724 793 -724 0 net=6361
rlabel metal2 954 -724 954 -724 0 net=5635
rlabel metal2 30 -726 30 -726 0 net=1841
rlabel metal2 170 -726 170 -726 0 net=1701
rlabel metal2 229 -726 229 -726 0 net=2744
rlabel metal2 317 -726 317 -726 0 net=3070
rlabel metal2 464 -726 464 -726 0 net=2965
rlabel metal2 481 -726 481 -726 0 net=4532
rlabel metal2 590 -726 590 -726 0 net=5879
rlabel metal2 744 -726 744 -726 0 net=5617
rlabel metal2 807 -726 807 -726 0 net=6435
rlabel metal2 44 -728 44 -728 0 net=3550
rlabel metal2 128 -728 128 -728 0 net=626
rlabel metal2 436 -728 436 -728 0 net=2645
rlabel metal2 488 -728 488 -728 0 net=3120
rlabel metal2 555 -728 555 -728 0 net=6476
rlabel metal2 2 -730 2 -730 0 net=4559
rlabel metal2 58 -730 58 -730 0 net=2168
rlabel metal2 240 -730 240 -730 0 net=556
rlabel metal2 558 -730 558 -730 0 net=6648
rlabel metal2 58 -732 58 -732 0 net=1235
rlabel metal2 205 -732 205 -732 0 net=1923
rlabel metal2 247 -732 247 -732 0 net=1577
rlabel metal2 348 -732 348 -732 0 net=3034
rlabel metal2 516 -732 516 -732 0 net=3314
rlabel metal2 674 -732 674 -732 0 net=4807
rlabel metal2 779 -732 779 -732 0 net=6289
rlabel metal2 891 -732 891 -732 0 net=404
rlabel metal2 86 -734 86 -734 0 net=5422
rlabel metal2 621 -734 621 -734 0 net=6876
rlabel metal2 86 -736 86 -736 0 net=1489
rlabel metal2 317 -736 317 -736 0 net=1867
rlabel metal2 506 -736 506 -736 0 net=4087
rlabel metal2 625 -736 625 -736 0 net=6744
rlabel metal2 51 -738 51 -738 0 net=3155
rlabel metal2 527 -738 527 -738 0 net=3813
rlabel metal2 565 -738 565 -738 0 net=6310
rlabel metal2 898 -738 898 -738 0 net=3625
rlabel metal2 65 -740 65 -740 0 net=4099
rlabel metal2 541 -740 541 -740 0 net=6255
rlabel metal2 723 -740 723 -740 0 net=5557
rlabel metal2 814 -740 814 -740 0 net=6541
rlabel metal2 89 -742 89 -742 0 net=5890
rlabel metal2 688 -742 688 -742 0 net=5383
rlabel metal2 737 -742 737 -742 0 net=5095
rlabel metal2 93 -744 93 -744 0 net=1958
rlabel metal2 254 -744 254 -744 0 net=1878
rlabel metal2 373 -744 373 -744 0 net=6432
rlabel metal2 51 -746 51 -746 0 net=3385
rlabel metal2 128 -746 128 -746 0 net=1729
rlabel metal2 569 -746 569 -746 0 net=3965
rlabel metal2 625 -746 625 -746 0 net=4471
rlabel metal2 667 -746 667 -746 0 net=6708
rlabel metal2 758 -746 758 -746 0 net=5955
rlabel metal2 821 -746 821 -746 0 net=6667
rlabel metal2 72 -748 72 -748 0 net=2318
rlabel metal2 394 -748 394 -748 0 net=4611
rlabel metal2 569 -748 569 -748 0 net=4055
rlabel metal2 579 -748 579 -748 0 net=6226
rlabel metal2 142 -750 142 -750 0 net=1696
rlabel metal2 261 -750 261 -750 0 net=1248
rlabel metal2 268 -750 268 -750 0 net=1217
rlabel metal2 331 -750 331 -750 0 net=2675
rlabel metal2 436 -750 436 -750 0 net=3505
rlabel metal2 485 -750 485 -750 0 net=5575
rlabel metal2 660 -750 660 -750 0 net=4783
rlabel metal2 9 -752 9 -752 0 net=4027
rlabel metal2 527 -752 527 -752 0 net=6831
rlabel metal2 107 -754 107 -754 0 net=1721
rlabel metal2 296 -754 296 -754 0 net=2809
rlabel metal2 576 -754 576 -754 0 net=5469
rlabel metal2 107 -756 107 -756 0 net=1326
rlabel metal2 142 -756 142 -756 0 net=2525
rlabel metal2 380 -756 380 -756 0 net=3559
rlabel metal2 583 -756 583 -756 0 net=4205
rlabel metal2 628 -756 628 -756 0 net=6618
rlabel metal2 100 -758 100 -758 0 net=564
rlabel metal2 145 -758 145 -758 0 net=2579
rlabel metal2 156 -758 156 -758 0 net=1557
rlabel metal2 191 -758 191 -758 0 net=4533
rlabel metal2 254 -758 254 -758 0 net=3833
rlabel metal2 296 -758 296 -758 0 net=1465
rlabel metal2 359 -758 359 -758 0 net=2333
rlabel metal2 394 -758 394 -758 0 net=2385
rlabel metal2 415 -758 415 -758 0 net=6641
rlabel metal2 842 -758 842 -758 0 net=6755
rlabel metal2 100 -760 100 -760 0 net=2725
rlabel metal2 639 -760 639 -760 0 net=4619
rlabel metal2 688 -760 688 -760 0 net=5947
rlabel metal2 786 -760 786 -760 0 net=6319
rlabel metal2 156 -762 156 -762 0 net=1739
rlabel metal2 212 -762 212 -762 0 net=1789
rlabel metal2 236 -762 236 -762 0 net=4733
rlabel metal2 702 -762 702 -762 0 net=5213
rlabel metal2 751 -762 751 -762 0 net=6883
rlabel metal2 37 -764 37 -764 0 net=3742
rlabel metal2 243 -764 243 -764 0 net=3601
rlabel metal2 408 -764 408 -764 0 net=2687
rlabel metal2 450 -764 450 -764 0 net=3467
rlabel metal2 681 -764 681 -764 0 net=5001
rlabel metal2 709 -764 709 -764 0 net=5431
rlabel metal2 863 -764 863 -764 0 net=6851
rlabel metal2 37 -766 37 -766 0 net=6619
rlabel metal2 520 -766 520 -766 0 net=4747
rlabel metal2 695 -766 695 -766 0 net=5187
rlabel metal2 177 -768 177 -768 0 net=2763
rlabel metal2 275 -768 275 -768 0 net=1130
rlabel metal2 404 -768 404 -768 0 net=2795
rlabel metal2 450 -768 450 -768 0 net=2209
rlabel metal2 611 -768 611 -768 0 net=4211
rlabel metal2 79 -770 79 -770 0 net=2503
rlabel metal2 289 -770 289 -770 0 net=2591
rlabel metal2 562 -770 562 -770 0 net=4319
rlabel metal2 632 -770 632 -770 0 net=4449
rlabel metal2 79 -772 79 -772 0 net=3393
rlabel metal2 492 -772 492 -772 0 net=6677
rlabel metal2 177 -774 177 -774 0 net=2371
rlabel metal2 289 -774 289 -774 0 net=1719
rlabel metal2 324 -774 324 -774 0 net=3822
rlabel metal2 513 -774 513 -774 0 net=4789
rlabel metal2 618 -774 618 -774 0 net=4279
rlabel metal2 121 -776 121 -776 0 net=2364
rlabel metal2 310 -776 310 -776 0 net=4159
rlabel metal2 338 -776 338 -776 0 net=1286
rlabel metal2 471 -776 471 -776 0 net=2871
rlabel metal2 110 -778 110 -778 0 net=2945
rlabel metal2 131 -778 131 -778 0 net=3061
rlabel metal2 345 -778 345 -778 0 net=1259
rlabel metal2 366 -780 366 -780 0 net=2105
rlabel metal2 16 -791 16 -791 0 net=5535
rlabel metal2 68 -791 68 -791 0 net=1137
rlabel metal2 114 -791 114 -791 0 net=63
rlabel metal2 310 -791 310 -791 0 net=1843
rlabel metal2 387 -791 387 -791 0 net=6759
rlabel metal2 961 -791 961 -791 0 net=2072
rlabel metal2 1017 -791 1017 -791 0 net=6335
rlabel metal2 1066 -791 1066 -791 0 net=5399
rlabel metal2 23 -793 23 -793 0 net=5674
rlabel metal2 79 -793 79 -793 0 net=3394
rlabel metal2 233 -793 233 -793 0 net=3062
rlabel metal2 338 -793 338 -793 0 net=2211
rlabel metal2 492 -793 492 -793 0 net=4808
rlabel metal2 814 -793 814 -793 0 net=6643
rlabel metal2 975 -793 975 -793 0 net=5629
rlabel metal2 23 -795 23 -795 0 net=2581
rlabel metal2 173 -795 173 -795 0 net=354
rlabel metal2 411 -795 411 -795 0 net=2592
rlabel metal2 523 -795 523 -795 0 net=6362
rlabel metal2 863 -795 863 -795 0 net=6679
rlabel metal2 989 -795 989 -795 0 net=765
rlabel metal2 1010 -795 1010 -795 0 net=5637
rlabel metal2 30 -797 30 -797 0 net=1842
rlabel metal2 380 -797 380 -797 0 net=2334
rlabel metal2 530 -797 530 -797 0 net=4620
rlabel metal2 653 -797 653 -797 0 net=5577
rlabel metal2 877 -797 877 -797 0 net=6853
rlabel metal2 37 -799 37 -799 0 net=6620
rlabel metal2 233 -799 233 -799 0 net=1467
rlabel metal2 380 -799 380 -799 0 net=2149
rlabel metal2 551 -799 551 -799 0 net=4489
rlabel metal2 695 -799 695 -799 0 net=4212
rlabel metal2 915 -799 915 -799 0 net=1401
rlabel metal2 37 -801 37 -801 0 net=3513
rlabel metal2 240 -801 240 -801 0 net=1720
rlabel metal2 296 -801 296 -801 0 net=1697
rlabel metal2 618 -801 618 -801 0 net=4450
rlabel metal2 817 -801 817 -801 0 net=6055
rlabel metal2 44 -803 44 -803 0 net=4560
rlabel metal2 254 -803 254 -803 0 net=3835
rlabel metal2 621 -803 621 -803 0 net=3626
rlabel metal2 919 -803 919 -803 0 net=6543
rlabel metal2 919 -803 919 -803 0 net=6543
rlabel metal2 47 -805 47 -805 0 net=729
rlabel metal2 268 -805 268 -805 0 net=1723
rlabel metal2 422 -805 422 -805 0 net=6777
rlabel metal2 51 -807 51 -807 0 net=2475
rlabel metal2 254 -807 254 -807 0 net=1869
rlabel metal2 422 -807 422 -807 0 net=2811
rlabel metal2 439 -807 439 -807 0 net=6443
rlabel metal2 30 -809 30 -809 0 net=2415
rlabel metal2 261 -809 261 -809 0 net=1453
rlabel metal2 537 -809 537 -809 0 net=6884
rlabel metal2 800 -809 800 -809 0 net=5957
rlabel metal2 58 -811 58 -811 0 net=1236
rlabel metal2 429 -811 429 -811 0 net=5215
rlabel metal2 751 -811 751 -811 0 net=5365
rlabel metal2 12 -813 12 -813 0 net=2377
rlabel metal2 72 -813 72 -813 0 net=2527
rlabel metal2 149 -813 149 -813 0 net=1791
rlabel metal2 282 -813 282 -813 0 net=1218
rlabel metal2 450 -813 450 -813 0 net=2967
rlabel metal2 485 -813 485 -813 0 net=3561
rlabel metal2 544 -813 544 -813 0 net=5217
rlabel metal2 639 -813 639 -813 0 net=4257
rlabel metal2 79 -815 79 -815 0 net=2489
rlabel metal2 471 -815 471 -815 0 net=2873
rlabel metal2 492 -815 492 -815 0 net=5121
rlabel metal2 821 -815 821 -815 0 net=6669
rlabel metal2 86 -817 86 -817 0 net=1490
rlabel metal2 443 -817 443 -817 0 net=2797
rlabel metal2 478 -817 478 -817 0 net=3255
rlabel metal2 681 -817 681 -817 0 net=4749
rlabel metal2 765 -817 765 -817 0 net=5461
rlabel metal2 828 -817 828 -817 0 net=6833
rlabel metal2 86 -819 86 -819 0 net=3387
rlabel metal2 114 -819 114 -819 0 net=2688
rlabel metal2 499 -819 499 -819 0 net=4101
rlabel metal2 695 -819 695 -819 0 net=2517
rlabel metal2 828 -819 828 -819 0 net=6527
rlabel metal2 891 -819 891 -819 0 net=6589
rlabel metal2 891 -819 891 -819 0 net=6589
rlabel metal2 93 -821 93 -821 0 net=1559
rlabel metal2 184 -821 184 -821 0 net=1261
rlabel metal2 506 -821 506 -821 0 net=3157
rlabel metal2 506 -821 506 -821 0 net=3157
rlabel metal2 513 -821 513 -821 0 net=3966
rlabel metal2 667 -821 667 -821 0 net=5948
rlabel metal2 709 -821 709 -821 0 net=5189
rlabel metal2 709 -821 709 -821 0 net=5189
rlabel metal2 716 -821 716 -821 0 net=5881
rlabel metal2 121 -823 121 -823 0 net=2947
rlabel metal2 513 -823 513 -823 0 net=4473
rlabel metal2 723 -823 723 -823 0 net=5385
rlabel metal2 835 -823 835 -823 0 net=5097
rlabel metal2 121 -825 121 -825 0 net=2719
rlabel metal2 138 -825 138 -825 0 net=4534
rlabel metal2 205 -825 205 -825 0 net=1925
rlabel metal2 289 -825 289 -825 0 net=2107
rlabel metal2 373 -825 373 -825 0 net=5047
rlabel metal2 730 -825 730 -825 0 net=4784
rlabel metal2 2 -827 2 -827 0 net=3733
rlabel metal2 219 -827 219 -827 0 net=6256
rlabel metal2 772 -827 772 -827 0 net=5471
rlabel metal2 128 -829 128 -829 0 net=1731
rlabel metal2 345 -829 345 -829 0 net=2119
rlabel metal2 516 -829 516 -829 0 net=4280
rlabel metal2 660 -829 660 -829 0 net=4735
rlabel metal2 772 -829 772 -829 0 net=6291
rlabel metal2 110 -831 110 -831 0 net=4627
rlabel metal2 670 -831 670 -831 0 net=5113
rlabel metal2 758 -831 758 -831 0 net=5433
rlabel metal2 117 -833 117 -833 0 net=4433
rlabel metal2 702 -833 702 -833 0 net=5003
rlabel metal2 131 -835 131 -835 0 net=6436
rlabel metal2 135 -837 135 -837 0 net=5901
rlabel metal2 142 -839 142 -839 0 net=2765
rlabel metal2 240 -839 240 -839 0 net=3987
rlabel metal2 534 -839 534 -839 0 net=4613
rlabel metal2 163 -841 163 -841 0 net=1703
rlabel metal2 191 -841 191 -841 0 net=1579
rlabel metal2 268 -841 268 -841 0 net=3427
rlabel metal2 415 -841 415 -841 0 net=4088
rlabel metal2 604 -841 604 -841 0 net=4791
rlabel metal2 156 -843 156 -843 0 net=1741
rlabel metal2 324 -843 324 -843 0 net=4161
rlabel metal2 611 -843 611 -843 0 net=4321
rlabel metal2 100 -845 100 -845 0 net=2727
rlabel metal2 355 -845 355 -845 0 net=4887
rlabel metal2 100 -847 100 -847 0 net=2677
rlabel metal2 355 -847 355 -847 0 net=6756
rlabel metal2 156 -849 156 -849 0 net=2553
rlabel metal2 331 -849 331 -849 0 net=2387
rlabel metal2 457 -849 457 -849 0 net=4029
rlabel metal2 793 -849 793 -849 0 net=5619
rlabel metal2 170 -851 170 -851 0 net=2372
rlabel metal2 198 -851 198 -851 0 net=2217
rlabel metal2 275 -851 275 -851 0 net=2505
rlabel metal2 457 -851 457 -851 0 net=2647
rlabel metal2 548 -851 548 -851 0 net=3815
rlabel metal2 177 -853 177 -853 0 net=2247
rlabel metal2 464 -853 464 -853 0 net=6623
rlabel metal2 212 -855 212 -855 0 net=5135
rlabel metal2 366 -857 366 -857 0 net=1044
rlabel metal2 579 -857 579 -857 0 net=6479
rlabel metal2 373 -859 373 -859 0 net=2141
rlabel metal2 548 -859 548 -859 0 net=2493
rlabel metal2 555 -861 555 -861 0 net=5663
rlabel metal2 359 -863 359 -863 0 net=3603
rlabel metal2 562 -863 562 -863 0 net=6133
rlabel metal2 275 -865 275 -865 0 net=4535
rlabel metal2 565 -865 565 -865 0 net=5117
rlabel metal2 565 -867 565 -867 0 net=6320
rlabel metal2 583 -869 583 -869 0 net=4207
rlabel metal2 779 -869 779 -869 0 net=5559
rlabel metal2 436 -871 436 -871 0 net=3507
rlabel metal2 436 -873 436 -873 0 net=3468
rlabel metal2 562 -875 562 -875 0 net=1501
rlabel metal2 569 -877 569 -877 0 net=4057
rlabel metal2 16 -888 16 -888 0 net=5536
rlabel metal2 121 -888 121 -888 0 net=2721
rlabel metal2 121 -888 121 -888 0 net=2721
rlabel metal2 135 -888 135 -888 0 net=2389
rlabel metal2 359 -888 359 -888 0 net=3508
rlabel metal2 600 -888 600 -888 0 net=5620
rlabel metal2 915 -888 915 -888 0 net=6544
rlabel metal2 947 -888 947 -888 0 net=6761
rlabel metal2 947 -888 947 -888 0 net=6761
rlabel metal2 954 -888 954 -888 0 net=6644
rlabel metal2 1013 -888 1013 -888 0 net=6336
rlabel metal2 1038 -888 1038 -888 0 net=5639
rlabel metal2 1080 -888 1080 -888 0 net=5401
rlabel metal2 16 -890 16 -890 0 net=5137
rlabel metal2 184 -890 184 -890 0 net=1262
rlabel metal2 366 -890 366 -890 0 net=4102
rlabel metal2 807 -890 807 -890 0 net=5435
rlabel metal2 807 -890 807 -890 0 net=5435
rlabel metal2 814 -890 814 -890 0 net=5463
rlabel metal2 870 -890 870 -890 0 net=6855
rlabel metal2 1010 -890 1010 -890 0 net=6457
rlabel metal2 23 -892 23 -892 0 net=2582
rlabel metal2 243 -892 243 -892 0 net=4536
rlabel metal2 289 -892 289 -892 0 net=2109
rlabel metal2 366 -892 366 -892 0 net=2813
rlabel metal2 429 -892 429 -892 0 net=5216
rlabel metal2 534 -892 534 -892 0 net=1502
rlabel metal2 817 -892 817 -892 0 net=6528
rlabel metal2 961 -892 961 -892 0 net=6057
rlabel metal2 2 -894 2 -894 0 net=3735
rlabel metal2 51 -894 51 -894 0 net=2476
rlabel metal2 422 -894 422 -894 0 net=2263
rlabel metal2 534 -894 534 -894 0 net=3605
rlabel metal2 569 -894 569 -894 0 net=5958
rlabel metal2 961 -894 961 -894 0 net=6779
rlabel metal2 989 -894 989 -894 0 net=5630
rlabel metal2 51 -896 51 -896 0 net=1793
rlabel metal2 156 -896 156 -896 0 net=2555
rlabel metal2 205 -896 205 -896 0 net=1417
rlabel metal2 289 -896 289 -896 0 net=1219
rlabel metal2 369 -896 369 -896 0 net=4474
rlabel metal2 520 -896 520 -896 0 net=5118
rlabel metal2 828 -896 828 -896 0 net=5579
rlabel metal2 891 -896 891 -896 0 net=6591
rlabel metal2 968 -896 968 -896 0 net=6835
rlabel metal2 58 -898 58 -898 0 net=2378
rlabel metal2 219 -898 219 -898 0 net=4750
rlabel metal2 765 -898 765 -898 0 net=5387
rlabel metal2 849 -898 849 -898 0 net=6135
rlabel metal2 891 -898 891 -898 0 net=6625
rlabel metal2 58 -900 58 -900 0 net=2249
rlabel metal2 408 -900 408 -900 0 net=2968
rlabel metal2 464 -900 464 -900 0 net=2799
rlabel metal2 474 -900 474 -900 0 net=3816
rlabel metal2 884 -900 884 -900 0 net=6681
rlabel metal2 65 -902 65 -902 0 net=2213
rlabel metal2 352 -902 352 -902 0 net=2143
rlabel metal2 387 -902 387 -902 0 net=2507
rlabel metal2 408 -902 408 -902 0 net=3837
rlabel metal2 628 -902 628 -902 0 net=5136
rlabel metal2 933 -902 933 -902 0 net=5098
rlabel metal2 72 -904 72 -904 0 net=2528
rlabel metal2 278 -904 278 -904 0 net=3063
rlabel metal2 527 -904 527 -904 0 net=3563
rlabel metal2 730 -904 730 -904 0 net=5115
rlabel metal2 72 -906 72 -906 0 net=1845
rlabel metal2 317 -906 317 -906 0 net=1732
rlabel metal2 499 -906 499 -906 0 net=4614
rlabel metal2 737 -906 737 -906 0 net=5123
rlabel metal2 751 -906 751 -906 0 net=5367
rlabel metal2 800 -906 800 -906 0 net=5561
rlabel metal2 93 -908 93 -908 0 net=1560
rlabel metal2 261 -908 261 -908 0 net=1455
rlabel metal2 324 -908 324 -908 0 net=2729
rlabel metal2 345 -908 345 -908 0 net=2120
rlabel metal2 499 -908 499 -908 0 net=3159
rlabel metal2 537 -908 537 -908 0 net=3743
rlabel metal2 548 -908 548 -908 0 net=6670
rlabel metal2 93 -910 93 -910 0 net=4031
rlabel metal2 635 -910 635 -910 0 net=4829
rlabel metal2 765 -910 765 -910 0 net=5473
rlabel metal2 842 -910 842 -910 0 net=5665
rlabel metal2 905 -910 905 -910 0 net=6481
rlabel metal2 107 -912 107 -912 0 net=2494
rlabel metal2 688 -912 688 -912 0 net=4793
rlabel metal2 723 -912 723 -912 0 net=5049
rlabel metal2 779 -912 779 -912 0 net=5273
rlabel metal2 107 -914 107 -914 0 net=2593
rlabel metal2 261 -914 261 -914 0 net=1725
rlabel metal2 310 -914 310 -914 0 net=2391
rlabel metal2 597 -914 597 -914 0 net=4365
rlabel metal2 702 -914 702 -914 0 net=4889
rlabel metal2 856 -914 856 -914 0 net=5883
rlabel metal2 905 -914 905 -914 0 net=6445
rlabel metal2 110 -916 110 -916 0 net=1870
rlabel metal2 285 -916 285 -916 0 net=3437
rlabel metal2 373 -916 373 -916 0 net=4011
rlabel metal2 604 -916 604 -916 0 net=4163
rlabel metal2 653 -916 653 -916 0 net=4491
rlabel metal2 709 -916 709 -916 0 net=5191
rlabel metal2 863 -916 863 -916 0 net=5903
rlabel metal2 912 -916 912 -916 0 net=365
rlabel metal2 114 -918 114 -918 0 net=1581
rlabel metal2 198 -918 198 -918 0 net=2219
rlabel metal2 411 -918 411 -918 0 net=4511
rlabel metal2 149 -920 149 -920 0 net=1705
rlabel metal2 170 -920 170 -920 0 net=2059
rlabel metal2 429 -920 429 -920 0 net=2649
rlabel metal2 467 -920 467 -920 0 net=4058
rlabel metal2 660 -920 660 -920 0 net=4629
rlabel metal2 30 -922 30 -922 0 net=2417
rlabel metal2 180 -922 180 -922 0 net=989
rlabel metal2 436 -922 436 -922 0 net=3345
rlabel metal2 551 -922 551 -922 0 net=4208
rlabel metal2 639 -922 639 -922 0 net=4259
rlabel metal2 660 -922 660 -922 0 net=4737
rlabel metal2 30 -924 30 -924 0 net=6013
rlabel metal2 439 -924 439 -924 0 net=517
rlabel metal2 86 -926 86 -926 0 net=3388
rlabel metal2 191 -926 191 -926 0 net=1469
rlabel metal2 439 -926 439 -926 0 net=4347
rlabel metal2 513 -926 513 -926 0 net=4035
rlabel metal2 625 -926 625 -926 0 net=4323
rlabel metal2 86 -928 86 -928 0 net=2767
rlabel metal2 156 -928 156 -928 0 net=3429
rlabel metal2 443 -928 443 -928 0 net=3989
rlabel metal2 632 -928 632 -928 0 net=4435
rlabel metal2 37 -930 37 -930 0 net=3515
rlabel metal2 457 -930 457 -930 0 net=2875
rlabel metal2 502 -930 502 -930 0 net=4381
rlabel metal2 37 -932 37 -932 0 net=4181
rlabel metal2 142 -932 142 -932 0 net=1699
rlabel metal2 471 -932 471 -932 0 net=3779
rlabel metal2 173 -934 173 -934 0 net=2425
rlabel metal2 478 -934 478 -934 0 net=3257
rlabel metal2 555 -934 555 -934 0 net=2519
rlabel metal2 198 -936 198 -936 0 net=3121
rlabel metal2 695 -936 695 -936 0 net=1402
rlabel metal2 208 -938 208 -938 0 net=1926
rlabel metal2 478 -938 478 -938 0 net=6105
rlabel metal2 44 -940 44 -940 0 net=812
rlabel metal2 562 -940 562 -940 0 net=5659
rlabel metal2 44 -942 44 -942 0 net=2949
rlabel metal2 212 -944 212 -944 0 net=838
rlabel metal2 233 -944 233 -944 0 net=1742
rlabel metal2 268 -944 268 -944 0 net=2151
rlabel metal2 401 -944 401 -944 0 net=2083
rlabel metal2 100 -946 100 -946 0 net=2679
rlabel metal2 79 -948 79 -948 0 net=2491
rlabel metal2 222 -948 222 -948 0 net=1503
rlabel metal2 79 -950 79 -950 0 net=1567
rlabel metal2 415 -952 415 -952 0 net=5004
rlabel metal2 758 -954 758 -954 0 net=6293
rlabel metal2 618 -956 618 -956 0 net=5219
rlabel metal2 618 -958 618 -958 0 net=3711
rlabel metal2 9 -969 9 -969 0 net=4013
rlabel metal2 380 -969 380 -969 0 net=3346
rlabel metal2 565 -969 565 -969 0 net=5116
rlabel metal2 835 -969 835 -969 0 net=5661
rlabel metal2 947 -969 947 -969 0 net=6763
rlabel metal2 1010 -969 1010 -969 0 net=6059
rlabel metal2 1038 -969 1038 -969 0 net=6458
rlabel metal2 1087 -969 1087 -969 0 net=5403
rlabel metal2 16 -971 16 -971 0 net=5138
rlabel metal2 474 -971 474 -971 0 net=372
rlabel metal2 16 -973 16 -973 0 net=2815
rlabel metal2 373 -973 373 -973 0 net=2085
rlabel metal2 408 -973 408 -973 0 net=3838
rlabel metal2 453 -973 453 -973 0 net=2800
rlabel metal2 481 -973 481 -973 0 net=4324
rlabel metal2 698 -973 698 -973 0 net=6856
rlabel metal2 891 -973 891 -973 0 net=6627
rlabel metal2 1059 -973 1059 -973 0 net=5641
rlabel metal2 37 -975 37 -975 0 net=4182
rlabel metal2 226 -975 226 -975 0 net=176
rlabel metal2 600 -975 600 -975 0 net=4830
rlabel metal2 751 -975 751 -975 0 net=5193
rlabel metal2 842 -975 842 -975 0 net=5667
rlabel metal2 954 -975 954 -975 0 net=3713
rlabel metal2 58 -977 58 -977 0 net=2250
rlabel metal2 488 -977 488 -977 0 net=3564
rlabel metal2 607 -977 607 -977 0 net=5562
rlabel metal2 828 -977 828 -977 0 net=5581
rlabel metal2 863 -977 863 -977 0 net=5905
rlabel metal2 898 -977 898 -977 0 net=6593
rlabel metal2 30 -979 30 -979 0 net=6014
rlabel metal2 635 -979 635 -979 0 net=6311
rlabel metal2 30 -981 30 -981 0 net=3123
rlabel metal2 240 -981 240 -981 0 net=439
rlabel metal2 639 -981 639 -981 0 net=4437
rlabel metal2 681 -981 681 -981 0 net=4383
rlabel metal2 758 -981 758 -981 0 net=6295
rlabel metal2 919 -981 919 -981 0 net=6836
rlabel metal2 982 -981 982 -981 0 net=6482
rlabel metal2 61 -983 61 -983 0 net=3973
rlabel metal2 653 -983 653 -983 0 net=6682
rlabel metal2 905 -983 905 -983 0 net=6447
rlabel metal2 93 -985 93 -985 0 net=4032
rlabel metal2 247 -985 247 -985 0 net=2681
rlabel metal2 471 -985 471 -985 0 net=5725
rlabel metal2 100 -987 100 -987 0 net=2492
rlabel metal2 338 -987 338 -987 0 net=2730
rlabel metal2 418 -987 418 -987 0 net=511
rlabel metal2 737 -987 737 -987 0 net=5125
rlabel metal2 856 -987 856 -987 0 net=5885
rlabel metal2 100 -989 100 -989 0 net=2409
rlabel metal2 247 -989 247 -989 0 net=1505
rlabel metal2 366 -989 366 -989 0 net=2877
rlabel metal2 492 -989 492 -989 0 net=4630
rlabel metal2 716 -989 716 -989 0 net=4795
rlabel metal2 765 -989 765 -989 0 net=5475
rlabel metal2 905 -989 905 -989 0 net=5569
rlabel metal2 929 -989 929 -989 0 net=6780
rlabel metal2 93 -991 93 -991 0 net=3269
rlabel metal2 495 -991 495 -991 0 net=6895
rlabel metal2 114 -993 114 -993 0 net=1583
rlabel metal2 261 -993 261 -993 0 net=1727
rlabel metal2 380 -993 380 -993 0 net=3259
rlabel metal2 506 -993 506 -993 0 net=4349
rlabel metal2 730 -993 730 -993 0 net=5857
rlabel metal2 933 -993 933 -993 0 net=6545
rlabel metal2 114 -995 114 -995 0 net=1707
rlabel metal2 177 -995 177 -995 0 net=897
rlabel metal2 383 -995 383 -995 0 net=2155
rlabel metal2 436 -995 436 -995 0 net=4995
rlabel metal2 793 -995 793 -995 0 net=5369
rlabel metal2 814 -995 814 -995 0 net=5465
rlabel metal2 943 -995 943 -995 0 net=6653
rlabel metal2 121 -997 121 -997 0 net=2722
rlabel metal2 131 -997 131 -997 0 net=6367
rlabel metal2 72 -999 72 -999 0 net=1847
rlabel metal2 131 -999 131 -999 0 net=3213
rlabel metal2 261 -999 261 -999 0 net=2265
rlabel metal2 457 -999 457 -999 0 net=3745
rlabel metal2 548 -999 548 -999 0 net=5427
rlabel metal2 65 -1001 65 -1001 0 net=2215
rlabel metal2 506 -1001 506 -1001 0 net=2625
rlabel metal2 660 -1001 660 -1001 0 net=4739
rlabel metal2 786 -1001 786 -1001 0 net=5389
rlabel metal2 814 -1001 814 -1001 0 net=4729
rlabel metal2 65 -1003 65 -1003 0 net=3431
rlabel metal2 180 -1003 180 -1003 0 net=1645
rlabel metal2 282 -1003 282 -1003 0 net=1437
rlabel metal2 576 -1003 576 -1003 0 net=6639
rlabel metal2 72 -1005 72 -1005 0 net=2221
rlabel metal2 285 -1005 285 -1005 0 net=5274
rlabel metal2 135 -1007 135 -1007 0 net=2390
rlabel metal2 450 -1007 450 -1007 0 net=5281
rlabel metal2 135 -1009 135 -1009 0 net=1601
rlabel metal2 142 -1011 142 -1011 0 net=1700
rlabel metal2 537 -1011 537 -1011 0 net=6136
rlabel metal2 44 -1013 44 -1013 0 net=2950
rlabel metal2 145 -1013 145 -1013 0 net=6857
rlabel metal2 149 -1015 149 -1015 0 net=2419
rlabel metal2 180 -1015 180 -1015 0 net=3521
rlabel metal2 296 -1015 296 -1015 0 net=2427
rlabel metal2 450 -1015 450 -1015 0 net=6321
rlabel metal2 23 -1017 23 -1017 0 net=3736
rlabel metal2 191 -1017 191 -1017 0 net=1471
rlabel metal2 299 -1017 299 -1017 0 net=3064
rlabel metal2 527 -1017 527 -1017 0 net=4367
rlabel metal2 723 -1017 723 -1017 0 net=4891
rlabel metal2 849 -1017 849 -1017 0 net=6107
rlabel metal2 23 -1019 23 -1019 0 net=3861
rlabel metal2 303 -1019 303 -1019 0 net=3439
rlabel metal2 597 -1019 597 -1019 0 net=6015
rlabel metal2 40 -1021 40 -1021 0 net=1429
rlabel metal2 198 -1021 198 -1021 0 net=1419
rlabel metal2 257 -1021 257 -1021 0 net=3391
rlabel metal2 604 -1021 604 -1021 0 net=5543
rlabel metal2 51 -1023 51 -1023 0 net=1794
rlabel metal2 303 -1023 303 -1023 0 net=2651
rlabel metal2 443 -1023 443 -1023 0 net=3517
rlabel metal2 702 -1023 702 -1023 0 net=4493
rlabel metal2 807 -1023 807 -1023 0 net=5437
rlabel metal2 51 -1025 51 -1025 0 net=2769
rlabel metal2 156 -1025 156 -1025 0 net=1329
rlabel metal2 310 -1025 310 -1025 0 net=2392
rlabel metal2 499 -1025 499 -1025 0 net=3161
rlabel metal2 541 -1025 541 -1025 0 net=4037
rlabel metal2 604 -1025 604 -1025 0 net=5651
rlabel metal2 44 -1027 44 -1027 0 net=2997
rlabel metal2 499 -1027 499 -1027 0 net=2601
rlabel metal2 79 -1029 79 -1029 0 net=1569
rlabel metal2 317 -1029 317 -1029 0 net=1457
rlabel metal2 387 -1029 387 -1029 0 net=2509
rlabel metal2 397 -1029 397 -1029 0 net=1383
rlabel metal2 443 -1029 443 -1029 0 net=5050
rlabel metal2 79 -1031 79 -1031 0 net=1885
rlabel metal2 516 -1031 516 -1031 0 net=5220
rlabel metal2 268 -1033 268 -1033 0 net=2153
rlabel metal2 324 -1033 324 -1033 0 net=2373
rlabel metal2 429 -1033 429 -1033 0 net=4819
rlabel metal2 107 -1035 107 -1035 0 net=2595
rlabel metal2 331 -1035 331 -1035 0 net=2111
rlabel metal2 534 -1035 534 -1035 0 net=3607
rlabel metal2 611 -1035 611 -1035 0 net=4165
rlabel metal2 702 -1035 702 -1035 0 net=4513
rlabel metal2 107 -1037 107 -1037 0 net=2061
rlabel metal2 184 -1037 184 -1037 0 net=2557
rlabel metal2 331 -1037 331 -1037 0 net=2145
rlabel metal2 551 -1037 551 -1037 0 net=5585
rlabel metal2 12 -1039 12 -1039 0 net=793
rlabel metal2 555 -1039 555 -1039 0 net=2521
rlabel metal2 646 -1039 646 -1039 0 net=4261
rlabel metal2 691 -1039 691 -1039 0 net=4521
rlabel metal2 184 -1041 184 -1041 0 net=1221
rlabel metal2 453 -1041 453 -1041 0 net=3289
rlabel metal2 569 -1041 569 -1041 0 net=3991
rlabel metal2 618 -1041 618 -1041 0 net=4653
rlabel metal2 289 -1043 289 -1043 0 net=1975
rlabel metal2 446 -1043 446 -1043 0 net=4875
rlabel metal2 625 -1043 625 -1043 0 net=6363
rlabel metal2 569 -1045 569 -1045 0 net=427
rlabel metal2 583 -1047 583 -1047 0 net=3781
rlabel metal2 86 -1049 86 -1049 0 net=1905
rlabel metal2 628 -1049 628 -1049 0 net=4109
rlabel metal2 646 -1051 646 -1051 0 net=4429
rlabel metal2 16 -1062 16 -1062 0 net=2817
rlabel metal2 478 -1062 478 -1062 0 net=5126
rlabel metal2 961 -1062 961 -1062 0 net=6365
rlabel metal2 1027 -1062 1027 -1062 0 net=6640
rlabel metal2 1059 -1062 1059 -1062 0 net=6654
rlabel metal2 1094 -1062 1094 -1062 0 net=5405
rlabel metal2 19 -1064 19 -1064 0 net=27
rlabel metal2 338 -1064 338 -1064 0 net=1458
rlabel metal2 464 -1064 464 -1064 0 net=2683
rlabel metal2 495 -1064 495 -1064 0 net=5438
rlabel metal2 989 -1064 989 -1064 0 net=6595
rlabel metal2 1094 -1064 1094 -1064 0 net=5643
rlabel metal2 30 -1066 30 -1066 0 net=3125
rlabel metal2 51 -1066 51 -1066 0 net=2770
rlabel metal2 65 -1066 65 -1066 0 net=3432
rlabel metal2 156 -1066 156 -1066 0 net=1330
rlabel metal2 191 -1066 191 -1066 0 net=1431
rlabel metal2 205 -1066 205 -1066 0 net=1355
rlabel metal2 205 -1066 205 -1066 0 net=1355
rlabel metal2 219 -1066 219 -1066 0 net=1675
rlabel metal2 275 -1066 275 -1066 0 net=3523
rlabel metal2 569 -1066 569 -1066 0 net=5544
rlabel metal2 996 -1066 996 -1066 0 net=6765
rlabel metal2 51 -1068 51 -1068 0 net=2571
rlabel metal2 142 -1068 142 -1068 0 net=25
rlabel metal2 282 -1068 282 -1068 0 net=1438
rlabel metal2 513 -1068 513 -1068 0 net=587
rlabel metal2 579 -1068 579 -1068 0 net=5428
rlabel metal2 1017 -1068 1017 -1068 0 net=6897
rlabel metal2 58 -1070 58 -1070 0 net=1747
rlabel metal2 369 -1070 369 -1070 0 net=5652
rlabel metal2 65 -1072 65 -1072 0 net=2267
rlabel metal2 296 -1072 296 -1072 0 net=2087
rlabel metal2 387 -1072 387 -1072 0 net=2375
rlabel metal2 576 -1072 576 -1072 0 net=3509
rlabel metal2 604 -1072 604 -1072 0 net=5041
rlabel metal2 926 -1072 926 -1072 0 net=6323
rlabel metal2 2 -1074 2 -1074 0 net=3295
rlabel metal2 303 -1074 303 -1074 0 net=2652
rlabel metal2 583 -1074 583 -1074 0 net=6628
rlabel metal2 79 -1076 79 -1076 0 net=1886
rlabel metal2 191 -1076 191 -1076 0 net=1585
rlabel metal2 222 -1076 222 -1076 0 net=1728
rlabel metal2 352 -1076 352 -1076 0 net=5662
rlabel metal2 86 -1078 86 -1078 0 net=1907
rlabel metal2 86 -1078 86 -1078 0 net=1907
rlabel metal2 114 -1078 114 -1078 0 net=1708
rlabel metal2 177 -1078 177 -1078 0 net=1421
rlabel metal2 233 -1078 233 -1078 0 net=1473
rlabel metal2 310 -1078 310 -1078 0 net=1570
rlabel metal2 569 -1078 569 -1078 0 net=3843
rlabel metal2 586 -1078 586 -1078 0 net=6296
rlabel metal2 940 -1078 940 -1078 0 net=3715
rlabel metal2 1097 -1078 1097 -1078 0 net=1
rlabel metal2 93 -1080 93 -1080 0 net=3271
rlabel metal2 121 -1080 121 -1080 0 net=1849
rlabel metal2 317 -1080 317 -1080 0 net=2154
rlabel metal2 572 -1080 572 -1080 0 net=6403
rlabel metal2 44 -1082 44 -1082 0 net=2999
rlabel metal2 156 -1082 156 -1082 0 net=1977
rlabel metal2 324 -1082 324 -1082 0 net=2558
rlabel metal2 593 -1082 593 -1082 0 net=5726
rlabel metal2 44 -1084 44 -1084 0 net=2757
rlabel metal2 597 -1084 597 -1084 0 net=3392
rlabel metal2 621 -1084 621 -1084 0 net=6563
rlabel metal2 93 -1086 93 -1086 0 net=1651
rlabel metal2 247 -1086 247 -1086 0 net=1507
rlabel metal2 289 -1086 289 -1086 0 net=2147
rlabel metal2 338 -1086 338 -1086 0 net=2429
rlabel metal2 439 -1086 439 -1086 0 net=4038
rlabel metal2 628 -1086 628 -1086 0 net=5194
rlabel metal2 863 -1086 863 -1086 0 net=5859
rlabel metal2 135 -1088 135 -1088 0 net=1603
rlabel metal2 345 -1088 345 -1088 0 net=3609
rlabel metal2 628 -1088 628 -1088 0 net=5668
rlabel metal2 107 -1090 107 -1090 0 net=2063
rlabel metal2 163 -1090 163 -1090 0 net=3737
rlabel metal2 509 -1090 509 -1090 0 net=6019
rlabel metal2 107 -1092 107 -1092 0 net=3617
rlabel metal2 184 -1092 184 -1092 0 net=1223
rlabel metal2 359 -1092 359 -1092 0 net=2113
rlabel metal2 387 -1092 387 -1092 0 net=2157
rlabel metal2 408 -1092 408 -1092 0 net=5067
rlabel metal2 912 -1092 912 -1092 0 net=6547
rlabel metal2 100 -1094 100 -1094 0 net=2411
rlabel metal2 198 -1094 198 -1094 0 net=3261
rlabel metal2 394 -1094 394 -1094 0 net=2511
rlabel metal2 411 -1094 411 -1094 0 net=131
rlabel metal2 541 -1094 541 -1094 0 net=3075
rlabel metal2 9 -1096 9 -1096 0 net=4015
rlabel metal2 166 -1096 166 -1096 0 net=6257
rlabel metal2 240 -1098 240 -1098 0 net=1647
rlabel metal2 359 -1098 359 -1098 0 net=1531
rlabel metal2 590 -1098 590 -1098 0 net=5466
rlabel metal2 919 -1098 919 -1098 0 net=6017
rlabel metal2 247 -1100 247 -1100 0 net=3401
rlabel metal2 646 -1100 646 -1100 0 net=691
rlabel metal2 688 -1100 688 -1100 0 net=5570
rlabel metal2 919 -1100 919 -1100 0 net=6131
rlabel metal2 380 -1102 380 -1102 0 net=2627
rlabel metal2 649 -1102 649 -1102 0 net=5886
rlabel metal2 1003 -1102 1003 -1102 0 net=6859
rlabel metal2 72 -1104 72 -1104 0 net=2222
rlabel metal2 688 -1104 688 -1104 0 net=6167
rlabel metal2 23 -1106 23 -1106 0 net=3863
rlabel metal2 394 -1106 394 -1106 0 net=3441
rlabel metal2 723 -1106 723 -1106 0 net=4495
rlabel metal2 849 -1106 849 -1106 0 net=6109
rlabel metal2 23 -1108 23 -1108 0 net=2969
rlabel metal2 401 -1108 401 -1108 0 net=2297
rlabel metal2 555 -1108 555 -1108 0 net=3291
rlabel metal2 639 -1108 639 -1108 0 net=2522
rlabel metal2 726 -1108 726 -1108 0 net=6139
rlabel metal2 422 -1110 422 -1110 0 net=2216
rlabel metal2 555 -1110 555 -1110 0 net=3993
rlabel metal2 730 -1110 730 -1110 0 net=6173
rlabel metal2 268 -1112 268 -1112 0 net=2597
rlabel metal2 429 -1112 429 -1112 0 net=3518
rlabel metal2 730 -1112 730 -1112 0 net=6448
rlabel metal2 429 -1114 429 -1114 0 net=4369
rlabel metal2 611 -1114 611 -1114 0 net=3975
rlabel metal2 667 -1114 667 -1114 0 net=4385
rlabel metal2 765 -1114 765 -1114 0 net=4997
rlabel metal2 856 -1114 856 -1114 0 net=5587
rlabel metal2 1038 -1114 1038 -1114 0 net=6375
rlabel metal2 436 -1116 436 -1116 0 net=6791
rlabel metal2 457 -1118 457 -1118 0 net=3747
rlabel metal2 779 -1118 779 -1118 0 net=5283
rlabel metal2 457 -1120 457 -1120 0 net=2603
rlabel metal2 520 -1120 520 -1120 0 net=3163
rlabel metal2 618 -1120 618 -1120 0 net=4877
rlabel metal2 786 -1120 786 -1120 0 net=4893
rlabel metal2 226 -1122 226 -1122 0 net=3215
rlabel metal2 520 -1122 520 -1122 0 net=4263
rlabel metal2 716 -1122 716 -1122 0 net=4655
rlabel metal2 800 -1122 800 -1122 0 net=5371
rlabel metal2 226 -1124 226 -1124 0 net=2821
rlabel metal2 530 -1124 530 -1124 0 net=4537
rlabel metal2 800 -1124 800 -1124 0 net=4731
rlabel metal2 821 -1124 821 -1124 0 net=5477
rlabel metal2 632 -1126 632 -1126 0 net=4741
rlabel metal2 758 -1126 758 -1126 0 net=4797
rlabel metal2 653 -1128 653 -1128 0 net=4167
rlabel metal2 807 -1128 807 -1128 0 net=4111
rlabel metal2 653 -1130 653 -1130 0 net=3783
rlabel metal2 772 -1130 772 -1130 0 net=4821
rlabel metal2 240 -1132 240 -1132 0 net=4457
rlabel metal2 807 -1132 807 -1132 0 net=5907
rlabel metal2 660 -1134 660 -1134 0 net=6312
rlabel metal2 681 -1136 681 -1136 0 net=4351
rlabel metal2 793 -1136 793 -1136 0 net=5391
rlabel metal2 1010 -1136 1010 -1136 0 net=6061
rlabel metal2 299 -1138 299 -1138 0 net=5037
rlabel metal2 695 -1138 695 -1138 0 net=4431
rlabel metal2 842 -1138 842 -1138 0 net=5583
rlabel metal2 492 -1140 492 -1140 0 net=4755
rlabel metal2 842 -1140 842 -1140 0 net=6369
rlabel metal2 485 -1142 485 -1142 0 net=6483
rlabel metal2 366 -1144 366 -1144 0 net=2879
rlabel metal2 674 -1144 674 -1144 0 net=4439
rlabel metal2 702 -1144 702 -1144 0 net=4515
rlabel metal2 366 -1146 366 -1146 0 net=1384
rlabel metal2 642 -1146 642 -1146 0 net=4695
rlabel metal2 709 -1146 709 -1146 0 net=4523
rlabel metal2 149 -1148 149 -1148 0 net=2421
rlabel metal2 674 -1148 674 -1148 0 net=5751
rlabel metal2 149 -1150 149 -1150 0 net=3613
rlabel metal2 709 -1150 709 -1150 0 net=3175
rlabel metal2 30 -1161 30 -1161 0 net=1192
rlabel metal2 590 -1161 590 -1161 0 net=524
rlabel metal2 639 -1161 639 -1161 0 net=5392
rlabel metal2 1090 -1161 1090 -1161 0 net=5406
rlabel metal2 30 -1163 30 -1163 0 net=3615
rlabel metal2 156 -1163 156 -1163 0 net=1978
rlabel metal2 243 -1163 243 -1163 0 net=1648
rlabel metal2 331 -1163 331 -1163 0 net=6132
rlabel metal2 33 -1165 33 -1165 0 net=1652
rlabel metal2 121 -1165 121 -1165 0 net=3001
rlabel metal2 156 -1165 156 -1165 0 net=1879
rlabel metal2 429 -1165 429 -1165 0 net=4370
rlabel metal2 464 -1165 464 -1165 0 net=6860
rlabel metal2 51 -1167 51 -1167 0 net=2573
rlabel metal2 436 -1167 436 -1167 0 net=157
rlabel metal2 58 -1169 58 -1169 0 net=1748
rlabel metal2 93 -1169 93 -1169 0 net=3739
rlabel metal2 194 -1169 194 -1169 0 net=884
rlabel metal2 247 -1169 247 -1169 0 net=3403
rlabel metal2 471 -1169 471 -1169 0 net=6366
rlabel metal2 58 -1171 58 -1171 0 net=1909
rlabel metal2 114 -1171 114 -1171 0 net=3273
rlabel metal2 128 -1171 128 -1171 0 net=2158
rlabel metal2 439 -1171 439 -1171 0 net=2684
rlabel metal2 495 -1171 495 -1171 0 net=4998
rlabel metal2 891 -1171 891 -1171 0 net=6565
rlabel metal2 51 -1173 51 -1173 0 net=4935
rlabel metal2 114 -1173 114 -1173 0 net=5038
rlabel metal2 684 -1173 684 -1173 0 net=4894
rlabel metal2 65 -1175 65 -1175 0 net=2269
rlabel metal2 65 -1175 65 -1175 0 net=2269
rlabel metal2 82 -1175 82 -1175 0 net=4016
rlabel metal2 128 -1175 128 -1175 0 net=2065
rlabel metal2 163 -1175 163 -1175 0 net=6018
rlabel metal2 135 -1177 135 -1177 0 net=1433
rlabel metal2 226 -1177 226 -1177 0 net=1183
rlabel metal2 639 -1177 639 -1177 0 net=4517
rlabel metal2 842 -1177 842 -1177 0 net=6371
rlabel metal2 117 -1179 117 -1179 0 net=4045
rlabel metal2 642 -1179 642 -1179 0 net=4432
rlabel metal2 772 -1179 772 -1179 0 net=5043
rlabel metal2 842 -1179 842 -1179 0 net=5439
rlabel metal2 170 -1181 170 -1181 0 net=2413
rlabel metal2 247 -1181 247 -1181 0 net=3443
rlabel metal2 446 -1181 446 -1181 0 net=3164
rlabel metal2 544 -1181 544 -1181 0 net=4732
rlabel metal2 919 -1181 919 -1181 0 net=6175
rlabel metal2 184 -1183 184 -1183 0 net=6331
rlabel metal2 37 -1185 37 -1185 0 net=3126
rlabel metal2 198 -1185 198 -1185 0 net=3263
rlabel metal2 495 -1185 495 -1185 0 net=4168
rlabel metal2 954 -1185 954 -1185 0 net=6793
rlabel metal2 37 -1187 37 -1187 0 net=5523
rlabel metal2 226 -1187 226 -1187 0 net=1225
rlabel metal2 331 -1187 331 -1187 0 net=3611
rlabel metal2 352 -1187 352 -1187 0 net=2115
rlabel metal2 380 -1187 380 -1187 0 net=2629
rlabel metal2 450 -1187 450 -1187 0 net=2819
rlabel metal2 548 -1187 548 -1187 0 net=3524
rlabel metal2 590 -1187 590 -1187 0 net=6351
rlabel metal2 79 -1189 79 -1189 0 net=2093
rlabel metal2 380 -1189 380 -1189 0 net=2299
rlabel metal2 450 -1189 450 -1189 0 net=2881
rlabel metal2 509 -1189 509 -1189 0 net=6324
rlabel metal2 79 -1191 79 -1191 0 net=3751
rlabel metal2 513 -1191 513 -1191 0 net=2376
rlabel metal2 597 -1191 597 -1191 0 net=5584
rlabel metal2 44 -1193 44 -1193 0 net=2758
rlabel metal2 516 -1193 516 -1193 0 net=5995
rlabel metal2 1010 -1193 1010 -1193 0 net=6063
rlabel metal2 44 -1195 44 -1195 0 net=1823
rlabel metal2 229 -1195 229 -1195 0 net=1474
rlabel metal2 282 -1195 282 -1195 0 net=1508
rlabel metal2 600 -1195 600 -1195 0 net=3716
rlabel metal2 72 -1197 72 -1197 0 net=3865
rlabel metal2 604 -1197 604 -1197 0 net=4352
rlabel metal2 723 -1197 723 -1197 0 net=6766
rlabel metal2 26 -1199 26 -1199 0 net=269
rlabel metal2 611 -1199 611 -1199 0 net=3977
rlabel metal2 611 -1199 611 -1199 0 net=3977
rlabel metal2 618 -1199 618 -1199 0 net=3748
rlabel metal2 660 -1199 660 -1199 0 net=6273
rlabel metal2 835 -1199 835 -1199 0 net=4497
rlabel metal2 72 -1201 72 -1201 0 net=1605
rlabel metal2 387 -1201 387 -1201 0 net=3845
rlabel metal2 618 -1201 618 -1201 0 net=4353
rlabel metal2 660 -1201 660 -1201 0 net=4441
rlabel metal2 716 -1201 716 -1201 0 net=5372
rlabel metal2 912 -1201 912 -1201 0 net=6549
rlabel metal2 107 -1203 107 -1203 0 net=3619
rlabel metal2 394 -1203 394 -1203 0 net=2423
rlabel metal2 485 -1203 485 -1203 0 net=3177
rlabel metal2 723 -1203 723 -1203 0 net=4823
rlabel metal2 884 -1203 884 -1203 0 net=6169
rlabel metal2 107 -1205 107 -1205 0 net=3477
rlabel metal2 233 -1205 233 -1205 0 net=75
rlabel metal2 310 -1205 310 -1205 0 net=3077
rlabel metal2 555 -1205 555 -1205 0 net=3995
rlabel metal2 667 -1205 667 -1205 0 net=4387
rlabel metal2 691 -1205 691 -1205 0 net=6663
rlabel metal2 219 -1207 219 -1207 0 net=1677
rlabel metal2 254 -1207 254 -1207 0 net=1851
rlabel metal2 401 -1207 401 -1207 0 net=2513
rlabel metal2 492 -1207 492 -1207 0 net=5293
rlabel metal2 677 -1207 677 -1207 0 net=6404
rlabel metal2 16 -1209 16 -1209 0 net=3997
rlabel metal2 261 -1209 261 -1209 0 net=1443
rlabel metal2 555 -1209 555 -1209 0 net=3511
rlabel metal2 586 -1209 586 -1209 0 net=6207
rlabel metal2 1045 -1209 1045 -1209 0 net=6899
rlabel metal2 177 -1211 177 -1211 0 net=1422
rlabel metal2 264 -1211 264 -1211 0 net=4137
rlabel metal2 695 -1211 695 -1211 0 net=4539
rlabel metal2 814 -1211 814 -1211 0 net=6376
rlabel metal2 1073 -1211 1073 -1211 0 net=5645
rlabel metal2 177 -1213 177 -1213 0 net=4389
rlabel metal2 541 -1213 541 -1213 0 net=1124
rlabel metal2 1038 -1213 1038 -1213 0 net=5155
rlabel metal2 268 -1215 268 -1215 0 net=2823
rlabel metal2 502 -1215 502 -1215 0 net=5961
rlabel metal2 856 -1215 856 -1215 0 net=4113
rlabel metal2 268 -1217 268 -1217 0 net=3627
rlabel metal2 520 -1217 520 -1217 0 net=4264
rlabel metal2 562 -1217 562 -1217 0 net=3293
rlabel metal2 653 -1217 653 -1217 0 net=3785
rlabel metal2 807 -1217 807 -1217 0 net=5909
rlabel metal2 275 -1219 275 -1219 0 net=1533
rlabel metal2 408 -1219 408 -1219 0 net=2529
rlabel metal2 562 -1219 562 -1219 0 net=4798
rlabel metal2 282 -1221 282 -1221 0 net=2857
rlabel metal2 709 -1221 709 -1221 0 net=5777
rlabel metal2 730 -1221 730 -1221 0 net=5479
rlabel metal2 142 -1223 142 -1223 0 net=6157
rlabel metal2 2 -1225 2 -1225 0 net=3297
rlabel metal2 289 -1225 289 -1225 0 net=2148
rlabel metal2 457 -1225 457 -1225 0 net=2604
rlabel metal2 569 -1225 569 -1225 0 net=4657
rlabel metal2 807 -1225 807 -1225 0 net=5589
rlabel metal2 2 -1227 2 -1227 0 net=1357
rlabel metal2 292 -1227 292 -1227 0 net=229
rlabel metal2 737 -1227 737 -1227 0 net=4459
rlabel metal2 758 -1227 758 -1227 0 net=4525
rlabel metal2 821 -1227 821 -1227 0 net=5285
rlabel metal2 9 -1229 9 -1229 0 net=741
rlabel metal2 296 -1229 296 -1229 0 net=2089
rlabel metal2 663 -1229 663 -1229 0 net=6395
rlabel metal2 9 -1231 9 -1231 0 net=3873
rlabel metal2 296 -1231 296 -1231 0 net=3217
rlabel metal2 702 -1231 702 -1231 0 net=4697
rlabel metal2 751 -1231 751 -1231 0 net=4879
rlabel metal2 779 -1231 779 -1231 0 net=6411
rlabel metal2 23 -1233 23 -1233 0 net=2970
rlabel metal2 499 -1233 499 -1233 0 net=4742
rlabel metal2 681 -1233 681 -1233 0 net=4605
rlabel metal2 751 -1233 751 -1233 0 net=4809
rlabel metal2 870 -1233 870 -1233 0 net=6021
rlabel metal2 23 -1235 23 -1235 0 net=5752
rlabel metal2 947 -1235 947 -1235 0 net=6485
rlabel metal2 191 -1237 191 -1237 0 net=1587
rlabel metal2 303 -1237 303 -1237 0 net=1769
rlabel metal2 933 -1237 933 -1237 0 net=6597
rlabel metal2 100 -1239 100 -1239 0 net=3451
rlabel metal2 338 -1239 338 -1239 0 net=2431
rlabel metal2 422 -1239 422 -1239 0 net=2599
rlabel metal2 793 -1239 793 -1239 0 net=4757
rlabel metal2 338 -1241 338 -1241 0 net=2223
rlabel metal2 961 -1241 961 -1241 0 net=6259
rlabel metal2 355 -1243 355 -1243 0 net=1068
rlabel metal2 443 -1243 443 -1243 0 net=5923
rlabel metal2 961 -1243 961 -1243 0 net=6111
rlabel metal2 443 -1245 443 -1245 0 net=3797
rlabel metal2 898 -1245 898 -1245 0 net=6141
rlabel metal2 863 -1247 863 -1247 0 net=5069
rlabel metal2 863 -1249 863 -1249 0 net=5861
rlabel metal2 187 -1251 187 -1251 0 net=6337
rlabel metal2 187 -1253 187 -1253 0 net=5675
rlabel metal2 2 -1264 2 -1264 0 net=1358
rlabel metal2 520 -1264 520 -1264 0 net=4526
rlabel metal2 814 -1264 814 -1264 0 net=5441
rlabel metal2 863 -1264 863 -1264 0 net=5863
rlabel metal2 863 -1264 863 -1264 0 net=5863
rlabel metal2 870 -1264 870 -1264 0 net=6023
rlabel metal2 898 -1264 898 -1264 0 net=5071
rlabel metal2 898 -1264 898 -1264 0 net=5071
rlabel metal2 982 -1264 982 -1264 0 net=4114
rlabel metal2 1066 -1264 1066 -1264 0 net=5157
rlabel metal2 9 -1266 9 -1266 0 net=3875
rlabel metal2 30 -1266 30 -1266 0 net=3616
rlabel metal2 170 -1266 170 -1266 0 net=2414
rlabel metal2 254 -1266 254 -1266 0 net=3998
rlabel metal2 513 -1266 513 -1266 0 net=5286
rlabel metal2 870 -1266 870 -1266 0 net=6339
rlabel metal2 947 -1266 947 -1266 0 net=6487
rlabel metal2 1017 -1266 1017 -1266 0 net=6065
rlabel metal2 1045 -1266 1045 -1266 0 net=6900
rlabel metal2 1045 -1266 1045 -1266 0 net=6900
rlabel metal2 1073 -1266 1073 -1266 0 net=5647
rlabel metal2 1073 -1266 1073 -1266 0 net=5647
rlabel metal2 9 -1268 9 -1268 0 net=1911
rlabel metal2 86 -1268 86 -1268 0 net=4937
rlabel metal2 604 -1268 604 -1268 0 net=5127
rlabel metal2 912 -1268 912 -1268 0 net=6209
rlabel metal2 1017 -1268 1017 -1268 0 net=4499
rlabel metal2 30 -1270 30 -1270 0 net=2073
rlabel metal2 93 -1270 93 -1270 0 net=3740
rlabel metal2 219 -1270 219 -1270 0 net=1678
rlabel metal2 240 -1270 240 -1270 0 net=1445
rlabel metal2 317 -1270 317 -1270 0 net=1852
rlabel metal2 331 -1270 331 -1270 0 net=3612
rlabel metal2 464 -1270 464 -1270 0 net=3405
rlabel metal2 541 -1270 541 -1270 0 net=6372
rlabel metal2 1020 -1270 1020 -1270 0 net=1
rlabel metal2 51 -1272 51 -1272 0 net=3218
rlabel metal2 320 -1272 320 -1272 0 net=3264
rlabel metal2 548 -1272 548 -1272 0 net=5480
rlabel metal2 744 -1272 744 -1272 0 net=4699
rlabel metal2 744 -1272 744 -1272 0 net=4699
rlabel metal2 751 -1272 751 -1272 0 net=4811
rlabel metal2 51 -1274 51 -1274 0 net=3003
rlabel metal2 159 -1274 159 -1274 0 net=627
rlabel metal2 478 -1274 478 -1274 0 net=4541
rlabel metal2 761 -1274 761 -1274 0 net=5491
rlabel metal2 884 -1274 884 -1274 0 net=6171
rlabel metal2 1003 -1274 1003 -1274 0 net=6577
rlabel metal2 54 -1276 54 -1276 0 net=3078
rlabel metal2 366 -1276 366 -1276 0 net=2574
rlabel metal2 576 -1276 576 -1276 0 net=3294
rlabel metal2 586 -1276 586 -1276 0 net=4388
rlabel metal2 884 -1276 884 -1276 0 net=6567
rlabel metal2 58 -1278 58 -1278 0 net=2859
rlabel metal2 292 -1278 292 -1278 0 net=4943
rlabel metal2 835 -1278 835 -1278 0 net=5963
rlabel metal2 65 -1280 65 -1280 0 net=2271
rlabel metal2 170 -1280 170 -1280 0 net=4138
rlabel metal2 677 -1280 677 -1280 0 net=6550
rlabel metal2 65 -1282 65 -1282 0 net=2225
rlabel metal2 369 -1282 369 -1282 0 net=2820
rlabel metal2 555 -1282 555 -1282 0 net=3512
rlabel metal2 583 -1282 583 -1282 0 net=2600
rlabel metal2 639 -1282 639 -1282 0 net=4519
rlabel metal2 817 -1282 817 -1282 0 net=5839
rlabel metal2 954 -1282 954 -1282 0 net=6795
rlabel metal2 93 -1284 93 -1284 0 net=3453
rlabel metal2 114 -1284 114 -1284 0 net=601
rlabel metal2 135 -1284 135 -1284 0 net=1434
rlabel metal2 331 -1284 331 -1284 0 net=3203
rlabel metal2 422 -1284 422 -1284 0 net=3917
rlabel metal2 565 -1284 565 -1284 0 net=4977
rlabel metal2 653 -1284 653 -1284 0 net=6112
rlabel metal2 100 -1286 100 -1286 0 net=3275
rlabel metal2 142 -1286 142 -1286 0 net=3298
rlabel metal2 292 -1286 292 -1286 0 net=3620
rlabel metal2 338 -1286 338 -1286 0 net=2117
rlabel metal2 425 -1286 425 -1286 0 net=2630
rlabel metal2 443 -1286 443 -1286 0 net=3799
rlabel metal2 604 -1286 604 -1286 0 net=3979
rlabel metal2 625 -1286 625 -1286 0 net=4047
rlabel metal2 653 -1286 653 -1286 0 net=4759
rlabel metal2 23 -1288 23 -1288 0 net=4325
rlabel metal2 142 -1288 142 -1288 0 net=1227
rlabel metal2 261 -1288 261 -1288 0 net=1535
rlabel metal2 282 -1288 282 -1288 0 net=2433
rlabel metal2 415 -1288 415 -1288 0 net=2825
rlabel metal2 443 -1288 443 -1288 0 net=4405
rlabel metal2 527 -1288 527 -1288 0 net=3893
rlabel metal2 537 -1288 537 -1288 0 net=4361
rlabel metal2 607 -1288 607 -1288 0 net=5910
rlabel metal2 940 -1288 940 -1288 0 net=6413
rlabel metal2 23 -1290 23 -1290 0 net=3479
rlabel metal2 117 -1290 117 -1290 0 net=4460
rlabel metal2 751 -1290 751 -1290 0 net=4593
rlabel metal2 72 -1292 72 -1292 0 net=1606
rlabel metal2 359 -1292 359 -1292 0 net=3787
rlabel metal2 793 -1292 793 -1292 0 net=5925
rlabel metal2 919 -1292 919 -1292 0 net=6177
rlabel metal2 72 -1294 72 -1294 0 net=3847
rlabel metal2 464 -1294 464 -1294 0 net=3753
rlabel metal2 537 -1294 537 -1294 0 net=3996
rlabel metal2 656 -1294 656 -1294 0 net=6332
rlabel metal2 107 -1296 107 -1296 0 net=1795
rlabel metal2 163 -1296 163 -1296 0 net=4585
rlabel metal2 660 -1296 660 -1296 0 net=4443
rlabel metal2 849 -1296 849 -1296 0 net=5997
rlabel metal2 968 -1296 968 -1296 0 net=6143
rlabel metal2 117 -1298 117 -1298 0 net=5753
rlabel metal2 373 -1298 373 -1298 0 net=2091
rlabel metal2 611 -1298 611 -1298 0 net=4355
rlabel metal2 660 -1298 660 -1298 0 net=4607
rlabel metal2 716 -1298 716 -1298 0 net=5019
rlabel metal2 793 -1298 793 -1298 0 net=4249
rlabel metal2 128 -1300 128 -1300 0 net=2067
rlabel metal2 173 -1300 173 -1300 0 net=6664
rlabel metal2 187 -1302 187 -1302 0 net=6352
rlabel metal2 191 -1304 191 -1304 0 net=6260
rlabel metal2 996 -1304 996 -1304 0 net=1745
rlabel metal2 194 -1306 194 -1306 0 net=3444
rlabel metal2 268 -1306 268 -1306 0 net=3628
rlabel metal2 667 -1306 667 -1306 0 net=5295
rlabel metal2 807 -1306 807 -1306 0 net=5591
rlabel metal2 194 -1308 194 -1308 0 net=2121
rlabel metal2 268 -1308 268 -1308 0 net=2095
rlabel metal2 373 -1308 373 -1308 0 net=3179
rlabel metal2 667 -1308 667 -1308 0 net=4649
rlabel metal2 198 -1310 198 -1310 0 net=2179
rlabel metal2 247 -1310 247 -1310 0 net=2883
rlabel metal2 485 -1310 485 -1310 0 net=3929
rlabel metal2 681 -1310 681 -1310 0 net=5045
rlabel metal2 786 -1310 786 -1310 0 net=5677
rlabel metal2 905 -1310 905 -1310 0 net=6397
rlabel metal2 184 -1312 184 -1312 0 net=810
rlabel metal2 275 -1312 275 -1312 0 net=2983
rlabel metal2 562 -1312 562 -1312 0 net=5787
rlabel metal2 933 -1312 933 -1312 0 net=6599
rlabel metal2 44 -1314 44 -1314 0 net=1825
rlabel metal2 201 -1314 201 -1314 0 net=2424
rlabel metal2 432 -1314 432 -1314 0 net=3017
rlabel metal2 509 -1314 509 -1314 0 net=1749
rlabel metal2 688 -1314 688 -1314 0 net=5779
rlabel metal2 716 -1314 716 -1314 0 net=4881
rlabel metal2 877 -1314 877 -1314 0 net=6159
rlabel metal2 44 -1316 44 -1316 0 net=4391
rlabel metal2 205 -1316 205 -1316 0 net=1589
rlabel metal2 296 -1316 296 -1316 0 net=2955
rlabel metal2 709 -1316 709 -1316 0 net=4825
rlabel metal2 758 -1316 758 -1316 0 net=6093
rlabel metal2 156 -1318 156 -1318 0 net=1881
rlabel metal2 212 -1318 212 -1318 0 net=3539
rlabel metal2 345 -1318 345 -1318 0 net=3057
rlabel metal2 499 -1318 499 -1318 0 net=3235
rlabel metal2 212 -1320 212 -1320 0 net=1771
rlabel metal2 355 -1320 355 -1320 0 net=5223
rlabel metal2 828 -1320 828 -1320 0 net=6275
rlabel metal2 37 -1322 37 -1322 0 net=5525
rlabel metal2 380 -1322 380 -1322 0 net=2301
rlabel metal2 432 -1322 432 -1322 0 net=3389
rlabel metal2 597 -1322 597 -1322 0 net=3867
rlabel metal2 37 -1324 37 -1324 0 net=2019
rlabel metal2 380 -1324 380 -1324 0 net=2515
rlabel metal2 422 -1324 422 -1324 0 net=2535
rlabel metal2 401 -1326 401 -1326 0 net=2531
rlabel metal2 457 -1326 457 -1326 0 net=5843
rlabel metal2 408 -1328 408 -1328 0 net=4659
rlabel metal2 492 -1330 492 -1330 0 net=5511
rlabel metal2 415 -1332 415 -1332 0 net=3415
rlabel metal2 569 -1332 569 -1332 0 net=3825
rlabel metal2 16 -1343 16 -1343 0 net=3876
rlabel metal2 89 -1343 89 -1343 0 net=2956
rlabel metal2 303 -1343 303 -1343 0 net=5526
rlabel metal2 352 -1343 352 -1343 0 net=2516
rlabel metal2 387 -1343 387 -1343 0 net=2092
rlabel metal2 471 -1343 471 -1343 0 net=4048
rlabel metal2 646 -1343 646 -1343 0 net=6094
rlabel metal2 919 -1343 919 -1343 0 net=5999
rlabel metal2 919 -1343 919 -1343 0 net=5999
rlabel metal2 950 -1343 950 -1343 0 net=1746
rlabel metal2 1031 -1343 1031 -1343 0 net=6066
rlabel metal2 16 -1345 16 -1345 0 net=5377
rlabel metal2 222 -1345 222 -1345 0 net=2434
rlabel metal2 292 -1345 292 -1345 0 net=4235
rlabel metal2 576 -1345 576 -1345 0 net=4444
rlabel metal2 891 -1345 891 -1345 0 net=5965
rlabel metal2 1024 -1345 1024 -1345 0 net=6137
rlabel metal2 1038 -1345 1038 -1345 0 net=5648
rlabel metal2 23 -1347 23 -1347 0 net=3480
rlabel metal2 107 -1347 107 -1347 0 net=1797
rlabel metal2 222 -1347 222 -1347 0 net=5754
rlabel metal2 338 -1347 338 -1347 0 net=2118
rlabel metal2 366 -1347 366 -1347 0 net=3019
rlabel metal2 471 -1347 471 -1347 0 net=4939
rlabel metal2 597 -1347 597 -1347 0 net=6172
rlabel metal2 971 -1347 971 -1347 0 net=6389
rlabel metal2 1045 -1347 1045 -1347 0 net=4003
rlabel metal2 1073 -1347 1073 -1347 0 net=5159
rlabel metal2 9 -1349 9 -1349 0 net=1912
rlabel metal2 107 -1349 107 -1349 0 net=3205
rlabel metal2 338 -1349 338 -1349 0 net=3755
rlabel metal2 495 -1349 495 -1349 0 net=3868
rlabel metal2 737 -1349 737 -1349 0 net=6340
rlabel metal2 30 -1351 30 -1351 0 net=2074
rlabel metal2 65 -1351 65 -1351 0 net=2227
rlabel metal2 79 -1351 79 -1351 0 net=3419
rlabel metal2 380 -1351 380 -1351 0 net=2303
rlabel metal2 411 -1351 411 -1351 0 net=1750
rlabel metal2 576 -1351 576 -1351 0 net=5046
rlabel metal2 705 -1351 705 -1351 0 net=4700
rlabel metal2 758 -1351 758 -1351 0 net=6600
rlabel metal2 30 -1353 30 -1353 0 net=3277
rlabel metal2 114 -1353 114 -1353 0 net=1983
rlabel metal2 254 -1353 254 -1353 0 net=2123
rlabel metal2 331 -1353 331 -1353 0 net=3919
rlabel metal2 579 -1353 579 -1353 0 net=6178
rlabel metal2 961 -1353 961 -1353 0 net=6415
rlabel metal2 37 -1355 37 -1355 0 net=2020
rlabel metal2 138 -1355 138 -1355 0 net=2532
rlabel metal2 415 -1355 415 -1355 0 net=3417
rlabel metal2 506 -1355 506 -1355 0 net=5780
rlabel metal2 705 -1355 705 -1355 0 net=4500
rlabel metal2 37 -1357 37 -1357 0 net=4393
rlabel metal2 51 -1357 51 -1357 0 net=3004
rlabel metal2 254 -1357 254 -1357 0 net=1267
rlabel metal2 509 -1357 509 -1357 0 net=4520
rlabel metal2 723 -1357 723 -1357 0 net=5225
rlabel metal2 821 -1357 821 -1357 0 net=5493
rlabel metal2 821 -1357 821 -1357 0 net=5493
rlabel metal2 835 -1357 835 -1357 0 net=5841
rlabel metal2 44 -1359 44 -1359 0 net=3059
rlabel metal2 401 -1359 401 -1359 0 net=3826
rlabel metal2 590 -1359 590 -1359 0 net=3981
rlabel metal2 618 -1359 618 -1359 0 net=6398
rlabel metal2 54 -1361 54 -1361 0 net=847
rlabel metal2 611 -1361 611 -1361 0 net=4357
rlabel metal2 632 -1361 632 -1361 0 net=4595
rlabel metal2 758 -1361 758 -1361 0 net=5129
rlabel metal2 835 -1361 835 -1361 0 net=5927
rlabel metal2 863 -1361 863 -1361 0 net=5865
rlabel metal2 65 -1363 65 -1363 0 net=3455
rlabel metal2 100 -1363 100 -1363 0 net=2537
rlabel metal2 429 -1363 429 -1363 0 net=6507
rlabel metal2 93 -1365 93 -1365 0 net=4543
rlabel metal2 523 -1365 523 -1365 0 net=5621
rlabel metal2 611 -1365 611 -1365 0 net=2465
rlabel metal2 684 -1365 684 -1365 0 net=6099
rlabel metal2 121 -1367 121 -1367 0 net=4326
rlabel metal2 247 -1367 247 -1367 0 net=2885
rlabel metal2 355 -1367 355 -1367 0 net=3729
rlabel metal2 429 -1367 429 -1367 0 net=3487
rlabel metal2 548 -1367 548 -1367 0 net=3591
rlabel metal2 688 -1367 688 -1367 0 net=4957
rlabel metal2 709 -1367 709 -1367 0 net=4827
rlabel metal2 842 -1367 842 -1367 0 net=5073
rlabel metal2 58 -1369 58 -1369 0 net=2861
rlabel metal2 128 -1369 128 -1369 0 net=3390
rlabel metal2 572 -1369 572 -1369 0 net=5139
rlabel metal2 765 -1369 765 -1369 0 net=5021
rlabel metal2 128 -1371 128 -1371 0 net=3239
rlabel metal2 268 -1371 268 -1371 0 net=2097
rlabel metal2 303 -1371 303 -1371 0 net=265
rlabel metal2 730 -1371 730 -1371 0 net=4945
rlabel metal2 779 -1371 779 -1371 0 net=5297
rlabel metal2 849 -1371 849 -1371 0 net=5845
rlabel metal2 145 -1373 145 -1373 0 net=623
rlabel metal2 159 -1373 159 -1373 0 net=3800
rlabel metal2 579 -1373 579 -1373 0 net=5835
rlabel metal2 870 -1373 870 -1373 0 net=6277
rlabel metal2 884 -1373 884 -1373 0 net=6569
rlabel metal2 149 -1375 149 -1375 0 net=2273
rlabel metal2 275 -1375 275 -1375 0 net=2985
rlabel metal2 415 -1375 415 -1375 0 net=2731
rlabel metal2 674 -1375 674 -1375 0 net=4883
rlabel metal2 737 -1375 737 -1375 0 net=5788
rlabel metal2 800 -1375 800 -1375 0 net=5679
rlabel metal2 884 -1375 884 -1375 0 net=6489
rlabel metal2 149 -1377 149 -1377 0 net=3869
rlabel metal2 184 -1377 184 -1377 0 net=1827
rlabel metal2 261 -1377 261 -1377 0 net=1537
rlabel metal2 282 -1377 282 -1377 0 net=2653
rlabel metal2 450 -1377 450 -1377 0 net=3237
rlabel metal2 583 -1377 583 -1377 0 net=5729
rlabel metal2 982 -1377 982 -1377 0 net=6145
rlabel metal2 163 -1379 163 -1379 0 net=2069
rlabel metal2 205 -1379 205 -1379 0 net=1883
rlabel metal2 324 -1379 324 -1379 0 net=1629
rlabel metal2 492 -1379 492 -1379 0 net=5057
rlabel metal2 23 -1381 23 -1381 0 net=3083
rlabel metal2 324 -1381 324 -1381 0 net=3181
rlabel metal2 443 -1381 443 -1381 0 net=4407
rlabel metal2 583 -1381 583 -1381 0 net=5592
rlabel metal2 443 -1383 443 -1383 0 net=3931
rlabel metal2 492 -1383 492 -1383 0 net=3407
rlabel metal2 586 -1383 586 -1383 0 net=6469
rlabel metal2 163 -1385 163 -1385 0 net=3631
rlabel metal2 359 -1385 359 -1385 0 net=3789
rlabel metal2 772 -1385 772 -1385 0 net=5513
rlabel metal2 947 -1385 947 -1385 0 net=6211
rlabel metal2 177 -1387 177 -1387 0 net=2181
rlabel metal2 359 -1387 359 -1387 0 net=2826
rlabel metal2 464 -1387 464 -1387 0 net=3135
rlabel metal2 597 -1387 597 -1387 0 net=4813
rlabel metal2 184 -1389 184 -1389 0 net=2481
rlabel metal2 369 -1389 369 -1389 0 net=5545
rlabel metal2 198 -1391 198 -1391 0 net=1591
rlabel metal2 317 -1391 317 -1391 0 net=1853
rlabel metal2 485 -1391 485 -1391 0 net=4363
rlabel metal2 565 -1391 565 -1391 0 net=5307
rlabel metal2 72 -1393 72 -1393 0 net=3849
rlabel metal2 646 -1393 646 -1393 0 net=4761
rlabel metal2 660 -1393 660 -1393 0 net=4609
rlabel metal2 72 -1395 72 -1395 0 net=3541
rlabel metal2 408 -1395 408 -1395 0 net=4660
rlabel metal2 653 -1395 653 -1395 0 net=5373
rlabel metal2 142 -1397 142 -1397 0 net=1229
rlabel metal2 408 -1397 408 -1397 0 net=1333
rlabel metal2 660 -1397 660 -1397 0 net=6796
rlabel metal2 212 -1399 212 -1399 0 net=1773
rlabel metal2 436 -1399 436 -1399 0 net=3895
rlabel metal2 681 -1399 681 -1399 0 net=5819
rlabel metal2 1003 -1399 1003 -1399 0 net=6579
rlabel metal2 212 -1401 212 -1401 0 net=1447
rlabel metal2 527 -1401 527 -1401 0 net=4587
rlabel metal2 695 -1401 695 -1401 0 net=5443
rlabel metal2 1003 -1401 1003 -1401 0 net=6713
rlabel metal2 625 -1403 625 -1403 0 net=4651
rlabel metal2 814 -1403 814 -1403 0 net=6161
rlabel metal2 639 -1405 639 -1405 0 net=4979
rlabel metal2 926 -1405 926 -1405 0 net=6025
rlabel metal2 639 -1407 639 -1407 0 net=4251
rlabel metal2 649 -1409 649 -1409 0 net=5563
rlabel metal2 16 -1420 16 -1420 0 net=5378
rlabel metal2 135 -1420 135 -1420 0 net=2099
rlabel metal2 310 -1420 310 -1420 0 net=2125
rlabel metal2 380 -1420 380 -1420 0 net=2305
rlabel metal2 380 -1420 380 -1420 0 net=2305
rlabel metal2 390 -1420 390 -1420 0 net=3238
rlabel metal2 471 -1420 471 -1420 0 net=4940
rlabel metal2 569 -1420 569 -1420 0 net=4884
rlabel metal2 681 -1420 681 -1420 0 net=5680
rlabel metal2 828 -1420 828 -1420 0 net=5309
rlabel metal2 842 -1420 842 -1420 0 net=5074
rlabel metal2 971 -1420 971 -1420 0 net=6138
rlabel metal2 1066 -1420 1066 -1420 0 net=5160
rlabel metal2 23 -1422 23 -1422 0 net=3084
rlabel metal2 268 -1422 268 -1422 0 net=2274
rlabel metal2 310 -1422 310 -1422 0 net=5005
rlabel metal2 758 -1422 758 -1422 0 net=5131
rlabel metal2 758 -1422 758 -1422 0 net=5131
rlabel metal2 793 -1422 793 -1422 0 net=5564
rlabel metal2 975 -1422 975 -1422 0 net=6417
rlabel metal2 1010 -1422 1010 -1422 0 net=6581
rlabel metal2 30 -1424 30 -1424 0 net=3278
rlabel metal2 163 -1424 163 -1424 0 net=321
rlabel metal2 338 -1424 338 -1424 0 net=3756
rlabel metal2 579 -1424 579 -1424 0 net=4828
rlabel metal2 793 -1424 793 -1424 0 net=5495
rlabel metal2 828 -1424 828 -1424 0 net=5547
rlabel metal2 877 -1424 877 -1424 0 net=5820
rlabel metal2 1024 -1424 1024 -1424 0 net=6390
rlabel metal2 30 -1426 30 -1426 0 net=5815
rlabel metal2 54 -1426 54 -1426 0 net=3240
rlabel metal2 138 -1426 138 -1426 0 net=947
rlabel metal2 163 -1426 163 -1426 0 net=1449
rlabel metal2 219 -1426 219 -1426 0 net=5374
rlabel metal2 663 -1426 663 -1426 0 net=5298
rlabel metal2 821 -1426 821 -1426 0 net=5967
rlabel metal2 929 -1426 929 -1426 0 net=5866
rlabel metal2 44 -1428 44 -1428 0 net=3060
rlabel metal2 142 -1428 142 -1428 0 net=1799
rlabel metal2 205 -1428 205 -1428 0 net=5842
rlabel metal2 44 -1430 44 -1430 0 net=3247
rlabel metal2 205 -1430 205 -1430 0 net=2005
rlabel metal2 289 -1430 289 -1430 0 net=3633
rlabel metal2 499 -1430 499 -1430 0 net=4408
rlabel metal2 516 -1430 516 -1430 0 net=4610
rlabel metal2 744 -1430 744 -1430 0 net=4947
rlabel metal2 58 -1432 58 -1432 0 net=5791
rlabel metal2 688 -1432 688 -1432 0 net=4959
rlabel metal2 723 -1432 723 -1432 0 net=5227
rlabel metal2 772 -1432 772 -1432 0 net=5515
rlabel metal2 835 -1432 835 -1432 0 net=5929
rlabel metal2 877 -1432 877 -1432 0 net=6183
rlabel metal2 65 -1434 65 -1434 0 net=3457
rlabel metal2 65 -1434 65 -1434 0 net=3457
rlabel metal2 72 -1434 72 -1434 0 net=3542
rlabel metal2 408 -1434 408 -1434 0 net=2723
rlabel metal2 523 -1434 523 -1434 0 net=4652
rlabel metal2 635 -1434 635 -1434 0 net=5058
rlabel metal2 835 -1434 835 -1434 0 net=6279
rlabel metal2 884 -1434 884 -1434 0 net=6490
rlabel metal2 926 -1434 926 -1434 0 net=6213
rlabel metal2 37 -1436 37 -1436 0 net=4394
rlabel metal2 75 -1436 75 -1436 0 net=4451
rlabel metal2 338 -1436 338 -1436 0 net=3827
rlabel metal2 597 -1436 597 -1436 0 net=4815
rlabel metal2 712 -1436 712 -1436 0 net=6162
rlabel metal2 842 -1436 842 -1436 0 net=6101
rlabel metal2 954 -1436 954 -1436 0 net=6715
rlabel metal2 37 -1438 37 -1438 0 net=3871
rlabel metal2 170 -1438 170 -1438 0 net=2183
rlabel metal2 212 -1438 212 -1438 0 net=1855
rlabel metal2 345 -1438 345 -1438 0 net=2887
rlabel metal2 394 -1438 394 -1438 0 net=2987
rlabel metal2 411 -1438 411 -1438 0 net=4364
rlabel metal2 513 -1438 513 -1438 0 net=3801
rlabel metal2 765 -1438 765 -1438 0 net=6601
rlabel metal2 86 -1440 86 -1440 0 net=5299
rlabel metal2 807 -1440 807 -1440 0 net=5731
rlabel metal2 870 -1440 870 -1440 0 net=6471
rlabel metal2 26 -1442 26 -1442 0 net=191
rlabel metal2 89 -1442 89 -1442 0 net=5265
rlabel metal2 814 -1442 814 -1442 0 net=5837
rlabel metal2 947 -1442 947 -1442 0 net=5533
rlabel metal2 93 -1444 93 -1444 0 net=4544
rlabel metal2 555 -1444 555 -1444 0 net=3851
rlabel metal2 583 -1444 583 -1444 0 net=4358
rlabel metal2 639 -1444 639 -1444 0 net=4253
rlabel metal2 681 -1444 681 -1444 0 net=6570
rlabel metal2 912 -1444 912 -1444 0 net=5847
rlabel metal2 93 -1446 93 -1446 0 net=1593
rlabel metal2 219 -1446 219 -1446 0 net=1884
rlabel metal2 292 -1446 292 -1446 0 net=2293
rlabel metal2 352 -1446 352 -1446 0 net=1335
rlabel metal2 555 -1446 555 -1446 0 net=2466
rlabel metal2 632 -1446 632 -1446 0 net=4597
rlabel metal2 646 -1446 646 -1446 0 net=4763
rlabel metal2 726 -1446 726 -1446 0 net=6341
rlabel metal2 100 -1448 100 -1448 0 net=2538
rlabel metal2 604 -1448 604 -1448 0 net=5622
rlabel metal2 79 -1450 79 -1450 0 net=3421
rlabel metal2 107 -1450 107 -1450 0 net=3206
rlabel metal2 660 -1450 660 -1450 0 net=5959
rlabel metal2 79 -1452 79 -1452 0 net=3183
rlabel metal2 362 -1452 362 -1452 0 net=4241
rlabel metal2 611 -1452 611 -1452 0 net=3791
rlabel metal2 751 -1452 751 -1452 0 net=5141
rlabel metal2 856 -1452 856 -1452 0 net=6001
rlabel metal2 107 -1454 107 -1454 0 net=2605
rlabel metal2 667 -1454 667 -1454 0 net=4981
rlabel metal2 863 -1454 863 -1454 0 net=6027
rlabel metal2 121 -1456 121 -1456 0 net=2862
rlabel metal2 247 -1456 247 -1456 0 net=1829
rlabel metal2 397 -1456 397 -1456 0 net=5022
rlabel metal2 121 -1458 121 -1458 0 net=3859
rlabel metal2 317 -1458 317 -1458 0 net=2732
rlabel metal2 418 -1458 418 -1458 0 net=3418
rlabel metal2 478 -1458 478 -1458 0 net=1631
rlabel metal2 702 -1458 702 -1458 0 net=5239
rlabel metal2 919 -1458 919 -1458 0 net=4004
rlabel metal2 149 -1460 149 -1460 0 net=3489
rlabel metal2 450 -1460 450 -1460 0 net=3137
rlabel metal2 478 -1460 478 -1460 0 net=3983
rlabel metal2 695 -1460 695 -1460 0 net=5445
rlabel metal2 933 -1460 933 -1460 0 net=6509
rlabel metal2 166 -1462 166 -1462 0 net=4621
rlabel metal2 590 -1462 590 -1462 0 net=4089
rlabel metal2 177 -1464 177 -1464 0 net=2070
rlabel metal2 198 -1464 198 -1464 0 net=3639
rlabel metal2 401 -1464 401 -1464 0 net=1289
rlabel metal2 562 -1464 562 -1464 0 net=4719
rlabel metal2 695 -1464 695 -1464 0 net=3877
rlabel metal2 982 -1464 982 -1464 0 net=6147
rlabel metal2 184 -1466 184 -1466 0 net=2483
rlabel metal2 366 -1466 366 -1466 0 net=3021
rlabel metal2 457 -1466 457 -1466 0 net=4237
rlabel metal2 618 -1466 618 -1466 0 net=5053
rlabel metal2 184 -1468 184 -1468 0 net=3920
rlabel metal2 366 -1468 366 -1468 0 net=2229
rlabel metal2 415 -1468 415 -1468 0 net=4009
rlabel metal2 191 -1470 191 -1470 0 net=1275
rlabel metal2 527 -1470 527 -1470 0 net=4589
rlabel metal2 243 -1472 243 -1472 0 net=4661
rlabel metal2 247 -1474 247 -1474 0 net=2275
rlabel metal2 320 -1474 320 -1474 0 net=3763
rlabel metal2 355 -1474 355 -1474 0 net=3903
rlabel metal2 443 -1474 443 -1474 0 net=3933
rlabel metal2 51 -1476 51 -1476 0 net=3347
rlabel metal2 464 -1476 464 -1476 0 net=3409
rlabel metal2 506 -1476 506 -1476 0 net=3593
rlabel metal2 254 -1478 254 -1478 0 net=1268
rlabel metal2 422 -1478 422 -1478 0 net=3731
rlabel metal2 548 -1478 548 -1478 0 net=3645
rlabel metal2 233 -1480 233 -1480 0 net=1775
rlabel metal2 422 -1480 422 -1480 0 net=3897
rlabel metal2 485 -1480 485 -1480 0 net=4689
rlabel metal2 114 -1482 114 -1482 0 net=1985
rlabel metal2 436 -1482 436 -1482 0 net=6399
rlabel metal2 114 -1484 114 -1484 0 net=2655
rlabel metal2 275 -1486 275 -1486 0 net=1539
rlabel metal2 226 -1488 226 -1488 0 net=1231
rlabel metal2 156 -1490 156 -1490 0 net=1459
rlabel metal2 9 -1501 9 -1501 0 net=1291
rlabel metal2 418 -1501 418 -1501 0 net=3732
rlabel metal2 506 -1501 506 -1501 0 net=3594
rlabel metal2 558 -1501 558 -1501 0 net=5142
rlabel metal2 800 -1501 800 -1501 0 net=6280
rlabel metal2 856 -1501 856 -1501 0 net=6003
rlabel metal2 996 -1501 996 -1501 0 net=6149
rlabel metal2 996 -1501 996 -1501 0 net=6149
rlabel metal2 1038 -1501 1038 -1501 0 net=6583
rlabel metal2 16 -1503 16 -1503 0 net=3491
rlabel metal2 194 -1503 194 -1503 0 net=625
rlabel metal2 506 -1503 506 -1503 0 net=906
rlabel metal2 726 -1503 726 -1503 0 net=5732
rlabel metal2 835 -1503 835 -1503 0 net=5313
rlabel metal2 23 -1505 23 -1505 0 net=1451
rlabel metal2 226 -1505 226 -1505 0 net=2126
rlabel metal2 366 -1505 366 -1505 0 net=2231
rlabel metal2 366 -1505 366 -1505 0 net=2231
rlabel metal2 380 -1505 380 -1505 0 net=2307
rlabel metal2 380 -1505 380 -1505 0 net=2307
rlabel metal2 394 -1505 394 -1505 0 net=6745
rlabel metal2 30 -1507 30 -1507 0 net=5816
rlabel metal2 268 -1507 268 -1507 0 net=3860
rlabel metal2 327 -1507 327 -1507 0 net=4010
rlabel metal2 667 -1507 667 -1507 0 net=4721
rlabel metal2 870 -1507 870 -1507 0 net=6473
rlabel metal2 30 -1509 30 -1509 0 net=1801
rlabel metal2 149 -1509 149 -1509 0 net=1359
rlabel metal2 418 -1509 418 -1509 0 net=2724
rlabel metal2 534 -1509 534 -1509 0 net=4931
rlabel metal2 870 -1509 870 -1509 0 net=5055
rlabel metal2 1003 -1509 1003 -1509 0 net=6419
rlabel metal2 37 -1511 37 -1511 0 net=3872
rlabel metal2 268 -1511 268 -1511 0 net=1831
rlabel metal2 341 -1511 341 -1511 0 net=5548
rlabel metal2 842 -1511 842 -1511 0 net=6103
rlabel metal2 37 -1513 37 -1513 0 net=4033
rlabel metal2 681 -1513 681 -1513 0 net=6602
rlabel metal2 891 -1513 891 -1513 0 net=5960
rlabel metal2 51 -1515 51 -1515 0 net=3423
rlabel metal2 121 -1515 121 -1515 0 net=5527
rlabel metal2 947 -1515 947 -1515 0 net=5848
rlabel metal2 58 -1517 58 -1517 0 net=5792
rlabel metal2 128 -1517 128 -1517 0 net=1461
rlabel metal2 163 -1517 163 -1517 0 net=1857
rlabel metal2 229 -1517 229 -1517 0 net=2484
rlabel metal2 275 -1517 275 -1517 0 net=1232
rlabel metal2 317 -1517 317 -1517 0 net=3985
rlabel metal2 513 -1517 513 -1517 0 net=3803
rlabel metal2 562 -1517 562 -1517 0 net=5446
rlabel metal2 733 -1517 733 -1517 0 net=6709
rlabel metal2 58 -1519 58 -1519 0 net=4283
rlabel metal2 422 -1519 422 -1519 0 net=3899
rlabel metal2 646 -1519 646 -1519 0 net=4591
rlabel metal2 65 -1521 65 -1521 0 net=3458
rlabel metal2 93 -1521 93 -1521 0 net=1594
rlabel metal2 352 -1521 352 -1521 0 net=1336
rlabel metal2 450 -1521 450 -1521 0 net=3138
rlabel metal2 520 -1521 520 -1521 0 net=3433
rlabel metal2 562 -1521 562 -1521 0 net=4243
rlabel metal2 618 -1521 618 -1521 0 net=4955
rlabel metal2 877 -1521 877 -1521 0 net=6185
rlabel metal2 44 -1523 44 -1523 0 net=3249
rlabel metal2 72 -1523 72 -1523 0 net=4231
rlabel metal2 877 -1523 877 -1523 0 net=6511
rlabel metal2 954 -1523 954 -1523 0 net=6717
rlabel metal2 79 -1525 79 -1525 0 net=3184
rlabel metal2 565 -1525 565 -1525 0 net=5838
rlabel metal2 898 -1525 898 -1525 0 net=6343
rlabel metal2 79 -1527 79 -1527 0 net=3646
rlabel metal2 618 -1527 618 -1527 0 net=3879
rlabel metal2 702 -1527 702 -1527 0 net=4983
rlabel metal2 744 -1527 744 -1527 0 net=5229
rlabel metal2 898 -1527 898 -1527 0 net=4949
rlabel metal2 82 -1529 82 -1529 0 net=3145
rlabel metal2 534 -1529 534 -1529 0 net=6649
rlabel metal2 86 -1531 86 -1531 0 net=2185
rlabel metal2 177 -1531 177 -1531 0 net=1987
rlabel metal2 247 -1531 247 -1531 0 net=2277
rlabel metal2 282 -1531 282 -1531 0 net=1540
rlabel metal2 359 -1531 359 -1531 0 net=3065
rlabel metal2 646 -1531 646 -1531 0 net=4005
rlabel metal2 863 -1531 863 -1531 0 net=6029
rlabel metal2 93 -1533 93 -1533 0 net=1201
rlabel metal2 436 -1533 436 -1533 0 net=19
rlabel metal2 905 -1533 905 -1533 0 net=6401
rlabel metal2 100 -1535 100 -1535 0 net=3525
rlabel metal2 254 -1535 254 -1535 0 net=1777
rlabel metal2 306 -1535 306 -1535 0 net=5291
rlabel metal2 912 -1535 912 -1535 0 net=5311
rlabel metal2 922 -1535 922 -1535 0 net=3749
rlabel metal2 964 -1535 964 -1535 0 net=5534
rlabel metal2 135 -1537 135 -1537 0 net=2100
rlabel metal2 464 -1537 464 -1537 0 net=3411
rlabel metal2 548 -1537 548 -1537 0 net=3793
rlabel metal2 653 -1537 653 -1537 0 net=5605
rlabel metal2 135 -1539 135 -1539 0 net=4239
rlabel metal2 474 -1539 474 -1539 0 net=4764
rlabel metal2 716 -1539 716 -1539 0 net=4961
rlabel metal2 926 -1539 926 -1539 0 net=6215
rlabel metal2 142 -1541 142 -1541 0 net=2295
rlabel metal2 362 -1541 362 -1541 0 net=5719
rlabel metal2 156 -1543 156 -1543 0 net=3023
rlabel metal2 569 -1543 569 -1543 0 net=3853
rlabel metal2 674 -1543 674 -1543 0 net=4255
rlabel metal2 180 -1545 180 -1545 0 net=2923
rlabel metal2 219 -1545 219 -1545 0 net=2831
rlabel metal2 289 -1545 289 -1545 0 net=3049
rlabel metal2 590 -1545 590 -1545 0 net=4091
rlabel metal2 660 -1545 660 -1545 0 net=4663
rlabel metal2 681 -1545 681 -1545 0 net=5968
rlabel metal2 184 -1547 184 -1547 0 net=2357
rlabel metal2 331 -1547 331 -1547 0 net=3765
rlabel metal2 604 -1547 604 -1547 0 net=1633
rlabel metal2 751 -1547 751 -1547 0 net=5241
rlabel metal2 107 -1549 107 -1549 0 net=2607
rlabel metal2 338 -1549 338 -1549 0 net=3829
rlabel metal2 590 -1549 590 -1549 0 net=4817
rlabel metal2 695 -1549 695 -1549 0 net=5007
rlabel metal2 758 -1549 758 -1549 0 net=5133
rlabel metal2 107 -1551 107 -1551 0 net=2657
rlabel metal2 170 -1551 170 -1551 0 net=2075
rlabel metal2 345 -1551 345 -1551 0 net=3349
rlabel metal2 460 -1551 460 -1551 0 net=4409
rlabel metal2 758 -1551 758 -1551 0 net=5339
rlabel metal2 114 -1553 114 -1553 0 net=3225
rlabel metal2 485 -1553 485 -1553 0 net=4691
rlabel metal2 772 -1553 772 -1553 0 net=5267
rlabel metal2 187 -1555 187 -1555 0 net=420
rlabel metal2 471 -1555 471 -1555 0 net=3635
rlabel metal2 663 -1555 663 -1555 0 net=4303
rlabel metal2 709 -1555 709 -1555 0 net=6239
rlabel metal2 222 -1557 222 -1557 0 net=40
rlabel metal2 684 -1557 684 -1557 0 net=6197
rlabel metal2 233 -1559 233 -1559 0 net=1986
rlabel metal2 723 -1559 723 -1559 0 net=6043
rlabel metal2 786 -1559 786 -1559 0 net=5517
rlabel metal2 233 -1561 233 -1561 0 net=4299
rlabel metal2 723 -1561 723 -1561 0 net=5301
rlabel metal2 793 -1561 793 -1561 0 net=5497
rlabel metal2 131 -1563 131 -1563 0 net=4625
rlabel metal2 803 -1563 803 -1563 0 net=6529
rlabel metal2 243 -1565 243 -1565 0 net=3697
rlabel metal2 583 -1565 583 -1565 0 net=4623
rlabel metal2 821 -1565 821 -1565 0 net=5931
rlabel metal2 247 -1567 247 -1567 0 net=297
rlabel metal2 254 -1569 254 -1569 0 net=3071
rlabel metal2 296 -1569 296 -1569 0 net=4453
rlabel metal2 639 -1569 639 -1569 0 net=4599
rlabel metal2 198 -1571 198 -1571 0 net=3641
rlabel metal2 310 -1571 310 -1571 0 net=4545
rlabel metal2 75 -1573 75 -1573 0 net=4081
rlabel metal2 373 -1573 373 -1573 0 net=3905
rlabel metal2 527 -1573 527 -1573 0 net=3935
rlabel metal2 2 -1575 2 -1575 0 net=3629
rlabel metal2 387 -1575 387 -1575 0 net=2889
rlabel metal2 495 -1575 495 -1575 0 net=3687
rlabel metal2 579 -1575 579 -1575 0 net=4157
rlabel metal2 198 -1577 198 -1577 0 net=2007
rlabel metal2 261 -1577 261 -1577 0 net=2001
rlabel metal2 191 -1579 191 -1579 0 net=1277
rlabel metal2 387 -1579 387 -1579 0 net=1619
rlabel metal2 397 -1581 397 -1581 0 net=3079
rlabel metal2 401 -1583 401 -1583 0 net=3709
rlabel metal2 408 -1585 408 -1585 0 net=2989
rlabel metal2 355 -1587 355 -1587 0 net=2841
rlabel metal2 2 -1598 2 -1598 0 net=3630
rlabel metal2 303 -1598 303 -1598 0 net=1779
rlabel metal2 355 -1598 355 -1598 0 net=4624
rlabel metal2 803 -1598 803 -1598 0 net=6216
rlabel metal2 2 -1600 2 -1600 0 net=6011
rlabel metal2 163 -1600 163 -1600 0 net=1858
rlabel metal2 359 -1600 359 -1600 0 net=2991
rlabel metal2 453 -1600 453 -1600 0 net=4592
rlabel metal2 23 -1602 23 -1602 0 net=1452
rlabel metal2 261 -1602 261 -1602 0 net=2003
rlabel metal2 373 -1602 373 -1602 0 net=3710
rlabel metal2 660 -1602 660 -1602 0 net=4305
rlabel metal2 709 -1602 709 -1602 0 net=6718
rlabel metal2 23 -1604 23 -1604 0 net=2659
rlabel metal2 114 -1604 114 -1604 0 net=3227
rlabel metal2 114 -1604 114 -1604 0 net=3227
rlabel metal2 121 -1604 121 -1604 0 net=4626
rlabel metal2 824 -1604 824 -1604 0 net=5312
rlabel metal2 982 -1604 982 -1604 0 net=6711
rlabel metal2 30 -1606 30 -1606 0 net=1802
rlabel metal2 236 -1606 236 -1606 0 net=3072
rlabel metal2 282 -1606 282 -1606 0 net=2833
rlabel metal2 429 -1606 429 -1606 0 net=3689
rlabel metal2 548 -1606 548 -1606 0 net=3794
rlabel metal2 548 -1606 548 -1606 0 net=3794
rlabel metal2 555 -1606 555 -1606 0 net=3805
rlabel metal2 723 -1606 723 -1606 0 net=5303
rlabel metal2 849 -1606 849 -1606 0 net=4158
rlabel metal2 919 -1606 919 -1606 0 net=6005
rlabel metal2 30 -1608 30 -1608 0 net=3637
rlabel metal2 492 -1608 492 -1608 0 net=4818
rlabel metal2 663 -1608 663 -1608 0 net=4256
rlabel metal2 37 -1610 37 -1610 0 net=4034
rlabel metal2 61 -1610 61 -1610 0 net=534
rlabel metal2 453 -1610 453 -1610 0 net=4950
rlabel metal2 37 -1612 37 -1612 0 net=1463
rlabel metal2 135 -1612 135 -1612 0 net=4240
rlabel metal2 376 -1612 376 -1612 0 net=2308
rlabel metal2 390 -1612 390 -1612 0 net=3698
rlabel metal2 583 -1612 583 -1612 0 net=3855
rlabel metal2 681 -1612 681 -1612 0 net=4411
rlabel metal2 758 -1612 758 -1612 0 net=5134
rlabel metal2 72 -1614 72 -1614 0 net=4232
rlabel metal2 891 -1614 891 -1614 0 net=3750
rlabel metal2 72 -1616 72 -1616 0 net=3081
rlabel metal2 457 -1616 457 -1616 0 net=4600
rlabel metal2 786 -1616 786 -1616 0 net=5315
rlabel metal2 947 -1616 947 -1616 0 net=5607
rlabel metal2 75 -1618 75 -1618 0 net=2937
rlabel metal2 289 -1618 289 -1618 0 net=3051
rlabel metal2 460 -1618 460 -1618 0 net=4341
rlabel metal2 555 -1618 555 -1618 0 net=6104
rlabel metal2 79 -1620 79 -1620 0 net=3066
rlabel metal2 688 -1620 688 -1620 0 net=4985
rlabel metal2 716 -1620 716 -1620 0 net=1635
rlabel metal2 996 -1620 996 -1620 0 net=6151
rlabel metal2 58 -1622 58 -1622 0 net=4285
rlabel metal2 674 -1622 674 -1622 0 net=4665
rlabel metal2 723 -1622 723 -1622 0 net=4723
rlabel metal2 772 -1622 772 -1622 0 net=6045
rlabel metal2 877 -1622 877 -1622 0 net=6513
rlabel metal2 82 -1624 82 -1624 0 net=3766
rlabel metal2 611 -1624 611 -1624 0 net=3937
rlabel metal2 695 -1624 695 -1624 0 net=5009
rlabel metal2 765 -1624 765 -1624 0 net=5231
rlabel metal2 877 -1624 877 -1624 0 net=6031
rlabel metal2 86 -1626 86 -1626 0 net=2186
rlabel metal2 289 -1626 289 -1626 0 net=4082
rlabel metal2 317 -1626 317 -1626 0 net=3986
rlabel metal2 562 -1626 562 -1626 0 net=4245
rlabel metal2 590 -1626 590 -1626 0 net=3881
rlabel metal2 639 -1626 639 -1626 0 net=5721
rlabel metal2 975 -1626 975 -1626 0 net=6421
rlabel metal2 107 -1628 107 -1628 0 net=2393
rlabel metal2 467 -1628 467 -1628 0 net=6402
rlabel metal2 121 -1630 121 -1630 0 net=1439
rlabel metal2 205 -1630 205 -1630 0 net=1279
rlabel metal2 268 -1630 268 -1630 0 net=1833
rlabel metal2 471 -1630 471 -1630 0 net=4483
rlabel metal2 702 -1630 702 -1630 0 net=4547
rlabel metal2 751 -1630 751 -1630 0 net=4693
rlabel metal2 1052 -1630 1052 -1630 0 net=6585
rlabel metal2 9 -1632 9 -1632 0 net=1293
rlabel metal2 212 -1632 212 -1632 0 net=2925
rlabel metal2 303 -1632 303 -1632 0 net=2843
rlabel metal2 474 -1632 474 -1632 0 net=363
rlabel metal2 9 -1634 9 -1634 0 net=5971
rlabel metal2 138 -1634 138 -1634 0 net=2733
rlabel metal2 310 -1634 310 -1634 0 net=1621
rlabel metal2 408 -1634 408 -1634 0 net=4007
rlabel metal2 730 -1634 730 -1634 0 net=6186
rlabel metal2 128 -1636 128 -1636 0 net=2359
rlabel metal2 212 -1636 212 -1636 0 net=4956
rlabel metal2 856 -1636 856 -1636 0 net=5499
rlabel metal2 142 -1638 142 -1638 0 net=2296
rlabel metal2 474 -1638 474 -1638 0 net=5289
rlabel metal2 744 -1638 744 -1638 0 net=4963
rlabel metal2 835 -1638 835 -1638 0 net=5519
rlabel metal2 65 -1640 65 -1640 0 net=3251
rlabel metal2 481 -1640 481 -1640 0 net=5292
rlabel metal2 926 -1640 926 -1640 0 net=6531
rlabel metal2 65 -1642 65 -1642 0 net=2309
rlabel metal2 142 -1642 142 -1642 0 net=1989
rlabel metal2 222 -1642 222 -1642 0 net=3642
rlabel metal2 317 -1642 317 -1642 0 net=1743
rlabel metal2 492 -1642 492 -1642 0 net=5449
rlabel metal2 842 -1642 842 -1642 0 net=5529
rlabel metal2 149 -1644 149 -1644 0 net=1361
rlabel metal2 194 -1644 194 -1644 0 net=1595
rlabel metal2 499 -1644 499 -1644 0 net=3413
rlabel metal2 537 -1644 537 -1644 0 net=6650
rlabel metal2 44 -1646 44 -1646 0 net=3015
rlabel metal2 156 -1646 156 -1646 0 net=3025
rlabel metal2 478 -1646 478 -1646 0 net=3147
rlabel metal2 513 -1646 513 -1646 0 net=6746
rlabel metal2 170 -1648 170 -1648 0 net=2076
rlabel metal2 544 -1648 544 -1648 0 net=5197
rlabel metal2 684 -1648 684 -1648 0 net=6459
rlabel metal2 170 -1650 170 -1650 0 net=2009
rlabel metal2 222 -1650 222 -1650 0 net=2278
rlabel metal2 296 -1650 296 -1650 0 net=666
rlabel metal2 513 -1650 513 -1650 0 net=3339
rlabel metal2 905 -1650 905 -1650 0 net=6241
rlabel metal2 86 -1652 86 -1652 0 net=5081
rlabel metal2 226 -1652 226 -1652 0 net=5056
rlabel metal2 933 -1652 933 -1652 0 net=6345
rlabel metal2 16 -1654 16 -1654 0 net=3492
rlabel metal2 233 -1654 233 -1654 0 net=267
rlabel metal2 366 -1654 366 -1654 0 net=2233
rlabel metal2 520 -1654 520 -1654 0 net=3435
rlabel metal2 772 -1654 772 -1654 0 net=5257
rlabel metal2 16 -1656 16 -1656 0 net=3425
rlabel metal2 163 -1656 163 -1656 0 net=1571
rlabel metal2 387 -1656 387 -1656 0 net=540
rlabel metal2 565 -1656 565 -1656 0 net=6474
rlabel metal2 51 -1658 51 -1658 0 net=3831
rlabel metal2 597 -1658 597 -1658 0 net=3901
rlabel metal2 779 -1658 779 -1658 0 net=5269
rlabel metal2 177 -1660 177 -1660 0 net=2891
rlabel metal2 558 -1660 558 -1660 0 net=4561
rlabel metal2 604 -1660 604 -1660 0 net=4455
rlabel metal2 793 -1660 793 -1660 0 net=5243
rlabel metal2 100 -1662 100 -1662 0 net=3527
rlabel metal2 464 -1662 464 -1662 0 net=3907
rlabel metal2 625 -1662 625 -1662 0 net=4093
rlabel metal2 814 -1662 814 -1662 0 net=5341
rlabel metal2 100 -1664 100 -1664 0 net=3127
rlabel metal2 275 -1664 275 -1664 0 net=4933
rlabel metal2 821 -1664 821 -1664 0 net=5933
rlabel metal2 93 -1666 93 -1666 0 net=1203
rlabel metal2 345 -1666 345 -1666 0 net=3351
rlabel metal2 653 -1666 653 -1666 0 net=4301
rlabel metal2 733 -1666 733 -1666 0 net=5487
rlabel metal2 863 -1666 863 -1666 0 net=6199
rlabel metal2 345 -1668 345 -1668 0 net=5349
rlabel metal2 478 -1668 478 -1668 0 net=364
rlabel metal2 394 -1670 394 -1670 0 net=4291
rlabel metal2 331 -1672 331 -1672 0 net=2609
rlabel metal2 488 -1672 488 -1672 0 net=4327
rlabel metal2 331 -1674 331 -1674 0 net=1803
rlabel metal2 2 -1685 2 -1685 0 net=6012
rlabel metal2 443 -1685 443 -1685 0 net=3026
rlabel metal2 593 -1685 593 -1685 0 net=4233
rlabel metal2 1024 -1685 1024 -1685 0 net=5167
rlabel metal2 1024 -1685 1024 -1685 0 net=5167
rlabel metal2 1027 -1685 1027 -1685 0 net=6586
rlabel metal2 2 -1687 2 -1687 0 net=1565
rlabel metal2 110 -1687 110 -1687 0 net=2360
rlabel metal2 152 -1687 152 -1687 0 net=4934
rlabel metal2 282 -1687 282 -1687 0 net=2611
rlabel metal2 429 -1687 429 -1687 0 net=3691
rlabel metal2 621 -1687 621 -1687 0 net=4666
rlabel metal2 730 -1687 730 -1687 0 net=5934
rlabel metal2 887 -1687 887 -1687 0 net=5608
rlabel metal2 1003 -1687 1003 -1687 0 net=6153
rlabel metal2 9 -1689 9 -1689 0 net=5972
rlabel metal2 198 -1689 198 -1689 0 net=3902
rlabel metal2 649 -1689 649 -1689 0 net=5500
rlabel metal2 891 -1689 891 -1689 0 net=6712
rlabel metal2 16 -1691 16 -1691 0 net=3426
rlabel metal2 233 -1691 233 -1691 0 net=1597
rlabel metal2 443 -1691 443 -1691 0 net=3923
rlabel metal2 716 -1691 716 -1691 0 net=4725
rlabel metal2 730 -1691 730 -1691 0 net=5011
rlabel metal2 779 -1691 779 -1691 0 net=5271
rlabel metal2 803 -1691 803 -1691 0 net=5488
rlabel metal2 821 -1691 821 -1691 0 net=6747
rlabel metal2 23 -1693 23 -1693 0 net=2660
rlabel metal2 198 -1693 198 -1693 0 net=2927
rlabel metal2 275 -1693 275 -1693 0 net=2771
rlabel metal2 779 -1693 779 -1693 0 net=5343
rlabel metal2 835 -1693 835 -1693 0 net=5521
rlabel metal2 912 -1693 912 -1693 0 net=6422
rlabel metal2 23 -1695 23 -1695 0 net=2933
rlabel metal2 240 -1695 240 -1695 0 net=2938
rlabel metal2 415 -1695 415 -1695 0 net=2835
rlabel metal2 457 -1695 457 -1695 0 net=5351
rlabel metal2 898 -1695 898 -1695 0 net=1637
rlabel metal2 30 -1697 30 -1697 0 net=3638
rlabel metal2 471 -1697 471 -1697 0 net=4456
rlabel metal2 793 -1697 793 -1697 0 net=5245
rlabel metal2 835 -1697 835 -1697 0 net=6461
rlabel metal2 30 -1699 30 -1699 0 net=5221
rlabel metal2 348 -1699 348 -1699 0 net=2163
rlabel metal2 394 -1699 394 -1699 0 net=2235
rlabel metal2 548 -1699 548 -1699 0 net=5801
rlabel metal2 849 -1699 849 -1699 0 net=6047
rlabel metal2 849 -1699 849 -1699 0 net=6047
rlabel metal2 898 -1699 898 -1699 0 net=6007
rlabel metal2 926 -1699 926 -1699 0 net=6533
rlabel metal2 37 -1701 37 -1701 0 net=1464
rlabel metal2 184 -1701 184 -1701 0 net=1363
rlabel metal2 205 -1701 205 -1701 0 net=1295
rlabel metal2 205 -1701 205 -1701 0 net=1295
rlabel metal2 222 -1701 222 -1701 0 net=1280
rlabel metal2 285 -1701 285 -1701 0 net=4008
rlabel metal2 467 -1701 467 -1701 0 net=5290
rlabel metal2 793 -1701 793 -1701 0 net=5451
rlabel metal2 863 -1701 863 -1701 0 net=6201
rlabel metal2 940 -1701 940 -1701 0 net=6693
rlabel metal2 37 -1703 37 -1703 0 net=4359
rlabel metal2 299 -1703 299 -1703 0 net=479
rlabel metal2 555 -1703 555 -1703 0 net=5199
rlabel metal2 639 -1703 639 -1703 0 net=5723
rlabel metal2 44 -1705 44 -1705 0 net=3016
rlabel metal2 65 -1705 65 -1705 0 net=2310
rlabel metal2 170 -1705 170 -1705 0 net=2011
rlabel metal2 317 -1705 317 -1705 0 net=1744
rlabel metal2 464 -1705 464 -1705 0 net=4079
rlabel metal2 688 -1705 688 -1705 0 net=4987
rlabel metal2 16 -1707 16 -1707 0 net=872
rlabel metal2 471 -1707 471 -1707 0 net=3939
rlabel metal2 569 -1707 569 -1707 0 net=4563
rlabel metal2 723 -1707 723 -1707 0 net=4965
rlabel metal2 44 -1709 44 -1709 0 net=3321
rlabel metal2 408 -1709 408 -1709 0 net=3806
rlabel metal2 51 -1711 51 -1711 0 net=3832
rlabel metal2 478 -1711 478 -1711 0 net=3315
rlabel metal2 548 -1711 548 -1711 0 net=4247
rlabel metal2 597 -1711 597 -1711 0 net=4287
rlabel metal2 51 -1713 51 -1713 0 net=1257
rlabel metal2 128 -1713 128 -1713 0 net=2279
rlabel metal2 485 -1713 485 -1713 0 net=6537
rlabel metal2 54 -1715 54 -1715 0 net=4155
rlabel metal2 261 -1715 261 -1715 0 net=1781
rlabel metal2 338 -1715 338 -1715 0 net=1835
rlabel metal2 352 -1715 352 -1715 0 net=2004
rlabel metal2 481 -1715 481 -1715 0 net=3938
rlabel metal2 614 -1715 614 -1715 0 net=4667
rlabel metal2 65 -1717 65 -1717 0 net=2127
rlabel metal2 243 -1717 243 -1717 0 net=2734
rlabel metal2 289 -1717 289 -1717 0 net=3340
rlabel metal2 516 -1717 516 -1717 0 net=5061
rlabel metal2 72 -1719 72 -1719 0 net=3082
rlabel metal2 488 -1719 488 -1719 0 net=3414
rlabel metal2 576 -1719 576 -1719 0 net=3883
rlabel metal2 618 -1719 618 -1719 0 net=5089
rlabel metal2 72 -1721 72 -1721 0 net=1573
rlabel metal2 177 -1721 177 -1721 0 net=2893
rlabel metal2 450 -1721 450 -1721 0 net=4307
rlabel metal2 79 -1723 79 -1723 0 net=1441
rlabel metal2 135 -1723 135 -1723 0 net=4133
rlabel metal2 492 -1723 492 -1723 0 net=4694
rlabel metal2 86 -1725 86 -1725 0 net=5083
rlabel metal2 947 -1725 947 -1725 0 net=6515
rlabel metal2 86 -1727 86 -1727 0 net=3659
rlabel metal2 121 -1727 121 -1727 0 net=1991
rlabel metal2 149 -1727 149 -1727 0 net=470
rlabel metal2 401 -1727 401 -1727 0 net=3253
rlabel metal2 541 -1727 541 -1727 0 net=4343
rlabel metal2 905 -1727 905 -1727 0 net=6243
rlabel metal2 138 -1729 138 -1729 0 net=5653
rlabel metal2 142 -1731 142 -1731 0 net=2845
rlabel metal2 317 -1731 317 -1731 0 net=1641
rlabel metal2 492 -1731 492 -1731 0 net=3031
rlabel metal2 149 -1733 149 -1733 0 net=762
rlabel metal2 247 -1733 247 -1733 0 net=1204
rlabel metal2 156 -1735 156 -1735 0 net=421
rlabel metal2 268 -1735 268 -1735 0 net=1649
rlabel metal2 331 -1735 331 -1735 0 net=1805
rlabel metal2 352 -1735 352 -1735 0 net=1893
rlabel metal2 495 -1735 495 -1735 0 net=3436
rlabel metal2 156 -1737 156 -1737 0 net=4149
rlabel metal2 289 -1737 289 -1737 0 net=2993
rlabel metal2 366 -1737 366 -1737 0 net=4302
rlabel metal2 674 -1737 674 -1737 0 net=6032
rlabel metal2 100 -1739 100 -1739 0 net=3129
rlabel metal2 366 -1739 366 -1739 0 net=6535
rlabel metal2 100 -1741 100 -1741 0 net=1351
rlabel metal2 177 -1741 177 -1741 0 net=2077
rlabel metal2 303 -1741 303 -1741 0 net=1623
rlabel metal2 369 -1741 369 -1741 0 net=3352
rlabel metal2 541 -1741 541 -1741 0 net=6089
rlabel metal2 114 -1743 114 -1743 0 net=3229
rlabel metal2 842 -1743 842 -1743 0 net=5531
rlabel metal2 107 -1745 107 -1745 0 net=2395
rlabel metal2 163 -1745 163 -1745 0 net=694
rlabel metal2 331 -1745 331 -1745 0 net=3323
rlabel metal2 373 -1745 373 -1745 0 net=3053
rlabel metal2 485 -1745 485 -1745 0 net=3005
rlabel metal2 786 -1745 786 -1745 0 net=5317
rlabel metal2 107 -1747 107 -1747 0 net=5849
rlabel metal2 187 -1749 187 -1749 0 net=6067
rlabel metal2 226 -1751 226 -1751 0 net=4095
rlabel metal2 786 -1751 786 -1751 0 net=6347
rlabel metal2 401 -1753 401 -1753 0 net=2897
rlabel metal2 499 -1753 499 -1753 0 net=3149
rlabel metal2 513 -1753 513 -1753 0 net=3856
rlabel metal2 625 -1753 625 -1753 0 net=4329
rlabel metal2 884 -1753 884 -1753 0 net=5681
rlabel metal2 373 -1755 373 -1755 0 net=2567
rlabel metal2 583 -1755 583 -1755 0 net=4549
rlabel metal2 800 -1755 800 -1755 0 net=5305
rlabel metal2 604 -1757 604 -1757 0 net=3909
rlabel metal2 604 -1759 604 -1759 0 net=4293
rlabel metal2 667 -1759 667 -1759 0 net=4413
rlabel metal2 569 -1761 569 -1761 0 net=4171
rlabel metal2 681 -1761 681 -1761 0 net=4485
rlabel metal2 695 -1763 695 -1763 0 net=5233
rlabel metal2 765 -1765 765 -1765 0 net=5259
rlabel metal2 422 -1767 422 -1767 0 net=3529
rlabel metal2 422 -1769 422 -1769 0 net=6659
rlabel metal2 2 -1780 2 -1780 0 net=1566
rlabel metal2 205 -1780 205 -1780 0 net=1296
rlabel metal2 565 -1780 565 -1780 0 net=6244
rlabel metal2 975 -1780 975 -1780 0 net=1638
rlabel metal2 9 -1782 9 -1782 0 net=5222
rlabel metal2 37 -1782 37 -1782 0 net=4360
rlabel metal2 313 -1782 313 -1782 0 net=2568
rlabel metal2 506 -1782 506 -1782 0 net=3150
rlabel metal2 583 -1782 583 -1782 0 net=4551
rlabel metal2 583 -1782 583 -1782 0 net=4551
rlabel metal2 590 -1782 590 -1782 0 net=6534
rlabel metal2 996 -1782 996 -1782 0 net=6154
rlabel metal2 23 -1784 23 -1784 0 net=2934
rlabel metal2 215 -1784 215 -1784 0 net=2012
rlabel metal2 310 -1784 310 -1784 0 net=2899
rlabel metal2 460 -1784 460 -1784 0 net=6202
rlabel metal2 947 -1784 947 -1784 0 net=5168
rlabel metal2 44 -1786 44 -1786 0 net=3322
rlabel metal2 369 -1786 369 -1786 0 net=2236
rlabel metal2 422 -1786 422 -1786 0 net=3910
rlabel metal2 726 -1786 726 -1786 0 net=6516
rlabel metal2 51 -1788 51 -1788 0 net=5724
rlabel metal2 915 -1788 915 -1788 0 net=5682
rlabel metal2 51 -1790 51 -1790 0 net=5323
rlabel metal2 369 -1790 369 -1790 0 net=2164
rlabel metal2 450 -1790 450 -1790 0 net=4308
rlabel metal2 590 -1790 590 -1790 0 net=4295
rlabel metal2 611 -1790 611 -1790 0 net=5352
rlabel metal2 54 -1792 54 -1792 0 net=1574
rlabel metal2 79 -1792 79 -1792 0 net=1442
rlabel metal2 107 -1792 107 -1792 0 net=1365
rlabel metal2 215 -1792 215 -1792 0 net=603
rlabel metal2 674 -1792 674 -1792 0 net=5246
rlabel metal2 842 -1792 842 -1792 0 net=5318
rlabel metal2 58 -1794 58 -1794 0 net=1993
rlabel metal2 128 -1794 128 -1794 0 net=2280
rlabel metal2 177 -1794 177 -1794 0 net=105
rlabel metal2 240 -1794 240 -1794 0 net=3254
rlabel metal2 541 -1794 541 -1794 0 net=4461
rlabel metal2 632 -1794 632 -1794 0 net=5654
rlabel metal2 65 -1796 65 -1796 0 net=2128
rlabel metal2 380 -1796 380 -1796 0 net=4080
rlabel metal2 642 -1796 642 -1796 0 net=6538
rlabel metal2 65 -1798 65 -1798 0 net=2847
rlabel metal2 149 -1798 149 -1798 0 net=4151
rlabel metal2 170 -1798 170 -1798 0 net=1353
rlabel metal2 226 -1798 226 -1798 0 net=4096
rlabel metal2 415 -1798 415 -1798 0 net=3055
rlabel metal2 464 -1798 464 -1798 0 net=4248
rlabel metal2 604 -1798 604 -1798 0 net=5085
rlabel metal2 814 -1798 814 -1798 0 net=6008
rlabel metal2 72 -1800 72 -1800 0 net=6181
rlabel metal2 464 -1800 464 -1800 0 net=3693
rlabel metal2 611 -1800 611 -1800 0 net=5261
rlabel metal2 898 -1800 898 -1800 0 net=5817
rlabel metal2 79 -1802 79 -1802 0 net=2251
rlabel metal2 618 -1802 618 -1802 0 net=4988
rlabel metal2 93 -1804 93 -1804 0 net=1258
rlabel metal2 135 -1804 135 -1804 0 net=4135
rlabel metal2 226 -1804 226 -1804 0 net=278
rlabel metal2 618 -1804 618 -1804 0 net=4967
rlabel metal2 751 -1804 751 -1804 0 net=6049
rlabel metal2 93 -1806 93 -1806 0 net=2397
rlabel metal2 121 -1806 121 -1806 0 net=3581
rlabel metal2 467 -1806 467 -1806 0 net=4701
rlabel metal2 527 -1806 527 -1806 0 net=6536
rlabel metal2 100 -1808 100 -1808 0 net=2751
rlabel metal2 478 -1808 478 -1808 0 net=3317
rlabel metal2 548 -1808 548 -1808 0 net=5897
rlabel metal2 100 -1810 100 -1810 0 net=2929
rlabel metal2 243 -1810 243 -1810 0 net=1249
rlabel metal2 499 -1810 499 -1810 0 net=4331
rlabel metal2 635 -1810 635 -1810 0 net=5272
rlabel metal2 110 -1812 110 -1812 0 net=3032
rlabel metal2 506 -1812 506 -1812 0 net=3530
rlabel metal2 828 -1812 828 -1812 0 net=6463
rlabel metal2 86 -1814 86 -1814 0 net=3661
rlabel metal2 534 -1814 534 -1814 0 net=5201
rlabel metal2 576 -1814 576 -1814 0 net=3884
rlabel metal2 86 -1816 86 -1816 0 net=2169
rlabel metal2 254 -1816 254 -1816 0 net=4156
rlabel metal2 576 -1816 576 -1816 0 net=4289
rlabel metal2 621 -1816 621 -1816 0 net=6113
rlabel metal2 114 -1818 114 -1818 0 net=3925
rlabel metal2 555 -1818 555 -1818 0 net=4415
rlabel metal2 674 -1818 674 -1818 0 net=4727
rlabel metal2 135 -1820 135 -1820 0 net=4911
rlabel metal2 170 -1820 170 -1820 0 net=3595
rlabel metal2 646 -1820 646 -1820 0 net=3999
rlabel metal2 142 -1822 142 -1822 0 net=1625
rlabel metal2 380 -1822 380 -1822 0 net=3231
rlabel metal2 653 -1822 653 -1822 0 net=5522
rlabel metal2 156 -1824 156 -1824 0 net=1205
rlabel metal2 247 -1824 247 -1824 0 net=2079
rlabel metal2 418 -1824 418 -1824 0 net=6571
rlabel metal2 653 -1824 653 -1824 0 net=5013
rlabel metal2 194 -1826 194 -1826 0 net=525
rlabel metal2 247 -1826 247 -1826 0 net=2773
rlabel metal2 282 -1826 282 -1826 0 net=2613
rlabel metal2 443 -1826 443 -1826 0 net=4565
rlabel metal2 702 -1826 702 -1826 0 net=4234
rlabel metal2 254 -1828 254 -1828 0 net=2287
rlabel metal2 520 -1828 520 -1828 0 net=5532
rlabel metal2 268 -1830 268 -1830 0 net=1650
rlabel metal2 660 -1830 660 -1830 0 net=4345
rlabel metal2 786 -1830 786 -1830 0 net=6349
rlabel metal2 261 -1832 261 -1832 0 net=1783
rlabel metal2 275 -1832 275 -1832 0 net=2177
rlabel metal2 681 -1832 681 -1832 0 net=4487
rlabel metal2 233 -1834 233 -1834 0 net=1599
rlabel metal2 282 -1834 282 -1834 0 net=1807
rlabel metal2 373 -1834 373 -1834 0 net=6671
rlabel metal2 597 -1834 597 -1834 0 net=2561
rlabel metal2 667 -1834 667 -1834 0 net=6695
rlabel metal2 233 -1836 233 -1836 0 net=1895
rlabel metal2 408 -1836 408 -1836 0 net=450
rlabel metal2 289 -1838 289 -1838 0 net=2995
rlabel metal2 681 -1838 681 -1838 0 net=5235
rlabel metal2 709 -1838 709 -1838 0 net=4669
rlabel metal2 289 -1840 289 -1840 0 net=3325
rlabel metal2 338 -1840 338 -1840 0 net=3007
rlabel metal2 688 -1840 688 -1840 0 net=5345
rlabel metal2 786 -1840 786 -1840 0 net=6069
rlabel metal2 296 -1842 296 -1842 0 net=1751
rlabel metal2 695 -1842 695 -1842 0 net=5453
rlabel metal2 838 -1842 838 -1842 0 net=4401
rlabel metal2 317 -1844 317 -1844 0 net=1643
rlabel metal2 709 -1844 709 -1844 0 net=5091
rlabel metal2 793 -1844 793 -1844 0 net=1871
rlabel metal2 317 -1846 317 -1846 0 net=1837
rlabel metal2 716 -1846 716 -1846 0 net=5803
rlabel metal2 324 -1848 324 -1848 0 net=2837
rlabel metal2 730 -1848 730 -1848 0 net=5851
rlabel metal2 331 -1850 331 -1850 0 net=4173
rlabel metal2 737 -1850 737 -1850 0 net=5063
rlabel metal2 807 -1850 807 -1850 0 net=6749
rlabel metal2 345 -1852 345 -1852 0 net=1156
rlabel metal2 429 -1854 429 -1854 0 net=2895
rlabel metal2 569 -1854 569 -1854 0 net=5306
rlabel metal2 429 -1856 429 -1856 0 net=3941
rlabel metal2 737 -1856 737 -1856 0 net=6661
rlabel metal2 359 -1858 359 -1858 0 net=3131
rlabel metal2 758 -1858 758 -1858 0 net=6121
rlabel metal2 821 -1860 821 -1860 0 net=6091
rlabel metal2 16 -1871 16 -1871 0 net=5325
rlabel metal2 58 -1871 58 -1871 0 net=1994
rlabel metal2 184 -1871 184 -1871 0 net=4136
rlabel metal2 219 -1871 219 -1871 0 net=1600
rlabel metal2 285 -1871 285 -1871 0 net=4670
rlabel metal2 23 -1873 23 -1873 0 net=6071
rlabel metal2 194 -1873 194 -1873 0 net=3095
rlabel metal2 229 -1873 229 -1873 0 net=805
rlabel metal2 243 -1873 243 -1873 0 net=1838
rlabel metal2 324 -1873 324 -1873 0 net=2838
rlabel metal2 415 -1873 415 -1873 0 net=3056
rlabel metal2 464 -1873 464 -1873 0 net=3694
rlabel metal2 509 -1873 509 -1873 0 net=6662
rlabel metal2 744 -1873 744 -1873 0 net=6115
rlabel metal2 744 -1873 744 -1873 0 net=6115
rlabel metal2 765 -1873 765 -1873 0 net=5899
rlabel metal2 765 -1873 765 -1873 0 net=5899
rlabel metal2 782 -1873 782 -1873 0 net=6350
rlabel metal2 51 -1875 51 -1875 0 net=5407
rlabel metal2 247 -1875 247 -1875 0 net=2775
rlabel metal2 334 -1875 334 -1875 0 net=5092
rlabel metal2 845 -1875 845 -1875 0 net=5818
rlabel metal2 58 -1877 58 -1877 0 net=1753
rlabel metal2 345 -1877 345 -1877 0 net=2459
rlabel metal2 345 -1877 345 -1877 0 net=2459
rlabel metal2 348 -1877 348 -1877 0 net=2996
rlabel metal2 359 -1877 359 -1877 0 net=4709
rlabel metal2 443 -1877 443 -1877 0 net=4567
rlabel metal2 702 -1877 702 -1877 0 net=6092
rlabel metal2 65 -1879 65 -1879 0 net=2848
rlabel metal2 177 -1879 177 -1879 0 net=1354
rlabel metal2 247 -1879 247 -1879 0 net=1251
rlabel metal2 411 -1879 411 -1879 0 net=1042
rlabel metal2 464 -1879 464 -1879 0 net=3319
rlabel metal2 520 -1879 520 -1879 0 net=4553
rlabel metal2 618 -1879 618 -1879 0 net=4968
rlabel metal2 702 -1879 702 -1879 0 net=6123
rlabel metal2 821 -1879 821 -1879 0 net=4403
rlabel metal2 65 -1881 65 -1881 0 net=5143
rlabel metal2 128 -1881 128 -1881 0 net=4153
rlabel metal2 177 -1881 177 -1881 0 net=312
rlabel metal2 471 -1881 471 -1881 0 net=3133
rlabel metal2 758 -1881 758 -1881 0 net=1872
rlabel metal2 72 -1883 72 -1883 0 net=6182
rlabel metal2 296 -1883 296 -1883 0 net=2753
rlabel metal2 418 -1883 418 -1883 0 net=6837
rlabel metal2 628 -1883 628 -1883 0 net=4728
rlabel metal2 709 -1883 709 -1883 0 net=1561
rlabel metal2 793 -1883 793 -1883 0 net=4001
rlabel metal2 72 -1885 72 -1885 0 net=5149
rlabel metal2 191 -1885 191 -1885 0 net=2178
rlabel metal2 338 -1885 338 -1885 0 net=3009
rlabel metal2 362 -1885 362 -1885 0 net=1644
rlabel metal2 527 -1885 527 -1885 0 net=4895
rlabel metal2 79 -1887 79 -1887 0 net=2252
rlabel metal2 289 -1887 289 -1887 0 net=3327
rlabel metal2 366 -1887 366 -1887 0 net=3651
rlabel metal2 530 -1887 530 -1887 0 net=2562
rlabel metal2 632 -1887 632 -1887 0 net=6070
rlabel metal2 814 -1887 814 -1887 0 net=6465
rlabel metal2 79 -1889 79 -1889 0 net=1809
rlabel metal2 289 -1889 289 -1889 0 net=3353
rlabel metal2 373 -1889 373 -1889 0 net=6673
rlabel metal2 674 -1889 674 -1889 0 net=5805
rlabel metal2 751 -1889 751 -1889 0 net=6051
rlabel metal2 44 -1891 44 -1891 0 net=394
rlabel metal2 310 -1891 310 -1891 0 net=2901
rlabel metal2 387 -1891 387 -1891 0 net=3857
rlabel metal2 471 -1891 471 -1891 0 net=4346
rlabel metal2 100 -1893 100 -1893 0 net=2931
rlabel metal2 394 -1893 394 -1893 0 net=2615
rlabel metal2 408 -1893 408 -1893 0 net=5919
rlabel metal2 646 -1893 646 -1893 0 net=6573
rlabel metal2 751 -1893 751 -1893 0 net=5065
rlabel metal2 100 -1895 100 -1895 0 net=3927
rlabel metal2 121 -1895 121 -1895 0 net=3583
rlabel metal2 215 -1895 215 -1895 0 net=115
rlabel metal2 422 -1895 422 -1895 0 net=99
rlabel metal2 646 -1895 646 -1895 0 net=5347
rlabel metal2 86 -1897 86 -1897 0 net=2170
rlabel metal2 142 -1897 142 -1897 0 net=1627
rlabel metal2 408 -1897 408 -1897 0 net=6696
rlabel metal2 681 -1897 681 -1897 0 net=5237
rlabel metal2 86 -1899 86 -1899 0 net=1897
rlabel metal2 380 -1899 380 -1899 0 net=3233
rlabel metal2 681 -1899 681 -1899 0 net=6237
rlabel metal2 93 -1901 93 -1901 0 net=2398
rlabel metal2 212 -1901 212 -1901 0 net=5715
rlabel metal2 422 -1901 422 -1901 0 net=3241
rlabel metal2 93 -1903 93 -1903 0 net=4175
rlabel metal2 429 -1903 429 -1903 0 net=3943
rlabel metal2 478 -1903 478 -1903 0 net=3663
rlabel metal2 548 -1903 548 -1903 0 net=747
rlabel metal2 107 -1905 107 -1905 0 net=1366
rlabel metal2 212 -1905 212 -1905 0 net=1785
rlabel metal2 310 -1905 310 -1905 0 net=3469
rlabel metal2 429 -1905 429 -1905 0 net=4703
rlabel metal2 548 -1905 548 -1905 0 net=5087
rlabel metal2 625 -1905 625 -1905 0 net=6635
rlabel metal2 107 -1907 107 -1907 0 net=4913
rlabel metal2 166 -1907 166 -1907 0 net=1381
rlabel metal2 268 -1907 268 -1907 0 net=2081
rlabel metal2 436 -1907 436 -1907 0 net=2896
rlabel metal2 436 -1907 436 -1907 0 net=2896
rlabel metal2 457 -1907 457 -1907 0 net=4831
rlabel metal2 551 -1907 551 -1907 0 net=4488
rlabel metal2 114 -1909 114 -1909 0 net=1207
rlabel metal2 254 -1909 254 -1909 0 net=2289
rlabel metal2 485 -1909 485 -1909 0 net=3771
rlabel metal2 583 -1909 583 -1909 0 net=5023
rlabel metal2 135 -1911 135 -1911 0 net=3597
rlabel metal2 254 -1911 254 -1911 0 net=2203
rlabel metal2 604 -1911 604 -1911 0 net=6750
rlabel metal2 131 -1913 131 -1913 0 net=2913
rlabel metal2 492 -1913 492 -1913 0 net=4333
rlabel metal2 506 -1913 506 -1913 0 net=4463
rlabel metal2 562 -1913 562 -1913 0 net=6033
rlabel metal2 149 -1915 149 -1915 0 net=2379
rlabel metal2 394 -1915 394 -1915 0 net=4501
rlabel metal2 625 -1915 625 -1915 0 net=5455
rlabel metal2 499 -1917 499 -1917 0 net=4290
rlabel metal2 653 -1917 653 -1917 0 net=5015
rlabel metal2 611 -1919 611 -1919 0 net=5263
rlabel metal2 453 -1921 453 -1921 0 net=6823
rlabel metal2 534 -1923 534 -1923 0 net=5203
rlabel metal2 534 -1925 534 -1925 0 net=4297
rlabel metal2 541 -1927 541 -1927 0 net=4417
rlabel metal2 555 -1929 555 -1929 0 net=5853
rlabel metal2 730 -1931 730 -1931 0 net=2261
rlabel metal2 33 -1942 33 -1942 0 net=806
rlabel metal2 40 -1942 40 -1942 0 net=54
rlabel metal2 51 -1942 51 -1942 0 net=5408
rlabel metal2 418 -1942 418 -1942 0 net=3234
rlabel metal2 677 -1942 677 -1942 0 net=5238
rlabel metal2 695 -1942 695 -1942 0 net=5017
rlabel metal2 814 -1942 814 -1942 0 net=6467
rlabel metal2 814 -1942 814 -1942 0 net=6467
rlabel metal2 37 -1944 37 -1944 0 net=1209
rlabel metal2 121 -1944 121 -1944 0 net=1933
rlabel metal2 191 -1944 191 -1944 0 net=5088
rlabel metal2 576 -1944 576 -1944 0 net=2262
rlabel metal2 782 -1944 782 -1944 0 net=4404
rlabel metal2 44 -1946 44 -1946 0 net=3599
rlabel metal2 138 -1946 138 -1946 0 net=1022
rlabel metal2 275 -1946 275 -1946 0 net=1628
rlabel metal2 373 -1946 373 -1946 0 net=2902
rlabel metal2 446 -1946 446 -1946 0 net=4334
rlabel metal2 495 -1946 495 -1946 0 net=4418
rlabel metal2 593 -1946 593 -1946 0 net=5456
rlabel metal2 653 -1946 653 -1946 0 net=5264
rlabel metal2 786 -1946 786 -1946 0 net=6053
rlabel metal2 58 -1948 58 -1948 0 net=1754
rlabel metal2 243 -1948 243 -1948 0 net=3858
rlabel metal2 394 -1948 394 -1948 0 net=2689
rlabel metal2 72 -1950 72 -1950 0 net=5151
rlabel metal2 93 -1950 93 -1950 0 net=4176
rlabel metal2 439 -1950 439 -1950 0 net=5769
rlabel metal2 653 -1950 653 -1950 0 net=5807
rlabel metal2 684 -1950 684 -1950 0 net=5066
rlabel metal2 772 -1950 772 -1950 0 net=6238
rlabel metal2 72 -1952 72 -1952 0 net=4915
rlabel metal2 114 -1952 114 -1952 0 net=5707
rlabel metal2 170 -1952 170 -1952 0 net=2915
rlabel metal2 219 -1952 219 -1952 0 net=3354
rlabel metal2 296 -1952 296 -1952 0 net=2754
rlabel metal2 611 -1952 611 -1952 0 net=6825
rlabel metal2 128 -1954 128 -1954 0 net=4154
rlabel metal2 229 -1954 229 -1954 0 net=2932
rlabel metal2 275 -1954 275 -1954 0 net=1423
rlabel metal2 352 -1954 352 -1954 0 net=3011
rlabel metal2 439 -1954 439 -1954 0 net=3320
rlabel metal2 499 -1954 499 -1954 0 net=6249
rlabel metal2 709 -1954 709 -1954 0 net=1563
rlabel metal2 51 -1956 51 -1956 0 net=5423
rlabel metal2 233 -1956 233 -1956 0 net=2082
rlabel metal2 296 -1956 296 -1956 0 net=2563
rlabel metal2 478 -1956 478 -1956 0 net=3665
rlabel metal2 506 -1956 506 -1956 0 net=4465
rlabel metal2 583 -1956 583 -1956 0 net=5025
rlabel metal2 618 -1956 618 -1956 0 net=6839
rlabel metal2 58 -1958 58 -1958 0 net=2139
rlabel metal2 142 -1958 142 -1958 0 net=1653
rlabel metal2 205 -1958 205 -1958 0 net=1382
rlabel metal2 317 -1958 317 -1958 0 net=5911
rlabel metal2 506 -1958 506 -1958 0 net=4833
rlabel metal2 516 -1958 516 -1958 0 net=6885
rlabel metal2 86 -1960 86 -1960 0 net=1899
rlabel metal2 254 -1960 254 -1960 0 net=2205
rlabel metal2 352 -1960 352 -1960 0 net=1943
rlabel metal2 415 -1960 415 -1960 0 net=6437
rlabel metal2 86 -1962 86 -1962 0 net=2337
rlabel metal2 317 -1962 317 -1962 0 net=2461
rlabel metal2 359 -1962 359 -1962 0 net=4711
rlabel metal2 408 -1962 408 -1962 0 net=3243
rlabel metal2 450 -1962 450 -1962 0 net=5854
rlabel metal2 579 -1962 579 -1962 0 net=5501
rlabel metal2 660 -1962 660 -1962 0 net=6035
rlabel metal2 688 -1962 688 -1962 0 net=5900
rlabel metal2 93 -1964 93 -1964 0 net=5867
rlabel metal2 184 -1964 184 -1964 0 net=3471
rlabel metal2 320 -1964 320 -1964 0 net=2616
rlabel metal2 415 -1964 415 -1964 0 net=2907
rlabel metal2 527 -1964 527 -1964 0 net=4897
rlabel metal2 555 -1964 555 -1964 0 net=4503
rlabel metal2 593 -1964 593 -1964 0 net=6797
rlabel metal2 744 -1964 744 -1964 0 net=6117
rlabel metal2 100 -1966 100 -1966 0 net=3928
rlabel metal2 163 -1966 163 -1966 0 net=3585
rlabel metal2 205 -1966 205 -1966 0 net=1371
rlabel metal2 247 -1966 247 -1966 0 net=1253
rlabel metal2 271 -1966 271 -1966 0 net=3279
rlabel metal2 453 -1966 453 -1966 0 net=3134
rlabel metal2 100 -1968 100 -1968 0 net=3381
rlabel metal2 149 -1968 149 -1968 0 net=2380
rlabel metal2 282 -1968 282 -1968 0 net=1551
rlabel metal2 527 -1968 527 -1968 0 net=4129
rlabel metal2 149 -1970 149 -1970 0 net=389
rlabel metal2 303 -1970 303 -1970 0 net=2291
rlabel metal2 366 -1970 366 -1970 0 net=3653
rlabel metal2 534 -1970 534 -1970 0 net=4298
rlabel metal2 597 -1970 597 -1970 0 net=5921
rlabel metal2 723 -1970 723 -1970 0 net=6637
rlabel metal2 159 -1972 159 -1972 0 net=4395
rlabel metal2 324 -1972 324 -1972 0 net=2777
rlabel metal2 369 -1972 369 -1972 0 net=4177
rlabel metal2 562 -1972 562 -1972 0 net=4569
rlabel metal2 723 -1972 723 -1972 0 net=4002
rlabel metal2 79 -1974 79 -1974 0 net=1811
rlabel metal2 401 -1974 401 -1974 0 net=3773
rlabel metal2 576 -1974 576 -1974 0 net=5593
rlabel metal2 65 -1976 65 -1976 0 net=5145
rlabel metal2 159 -1976 159 -1976 0 net=3355
rlabel metal2 198 -1976 198 -1976 0 net=3097
rlabel metal2 422 -1976 422 -1976 0 net=2577
rlabel metal2 597 -1976 597 -1976 0 net=5348
rlabel metal2 16 -1978 16 -1978 0 net=5327
rlabel metal2 191 -1978 191 -1978 0 net=2015
rlabel metal2 212 -1978 212 -1978 0 net=1787
rlabel metal2 443 -1978 443 -1978 0 net=3945
rlabel metal2 632 -1978 632 -1978 0 net=6675
rlabel metal2 646 -1978 646 -1978 0 net=5821
rlabel metal2 212 -1980 212 -1980 0 net=1269
rlabel metal2 457 -1980 457 -1980 0 net=4554
rlabel metal2 569 -1980 569 -1980 0 net=5205
rlabel metal2 338 -1982 338 -1982 0 net=3329
rlabel metal2 520 -1982 520 -1982 0 net=3191
rlabel metal2 338 -1984 338 -1984 0 net=5717
rlabel metal2 429 -1984 429 -1984 0 net=4705
rlabel metal2 681 -1984 681 -1984 0 net=6125
rlabel metal2 380 -1986 380 -1986 0 net=5747
rlabel metal2 702 -1986 702 -1986 0 net=6575
rlabel metal2 436 -1988 436 -1988 0 net=6491
rlabel metal2 23 -1990 23 -1990 0 net=6072
rlabel metal2 16 -2001 16 -2001 0 net=5869
rlabel metal2 156 -2001 156 -2001 0 net=1959
rlabel metal2 201 -2001 201 -2001 0 net=37
rlabel metal2 229 -2001 229 -2001 0 net=5718
rlabel metal2 387 -2001 387 -2001 0 net=3012
rlabel metal2 432 -2001 432 -2001 0 net=4706
rlabel metal2 576 -2001 576 -2001 0 net=5595
rlabel metal2 576 -2001 576 -2001 0 net=5595
rlabel metal2 586 -2001 586 -2001 0 net=6676
rlabel metal2 646 -2001 646 -2001 0 net=5822
rlabel metal2 670 -2001 670 -2001 0 net=1564
rlabel metal2 796 -2001 796 -2001 0 net=6468
rlabel metal2 30 -2003 30 -2003 0 net=5147
rlabel metal2 177 -2003 177 -2003 0 net=2917
rlabel metal2 313 -2003 313 -2003 0 net=1812
rlabel metal2 331 -2003 331 -2003 0 net=2206
rlabel metal2 488 -2003 488 -2003 0 net=263
rlabel metal2 548 -2003 548 -2003 0 net=4467
rlabel metal2 37 -2005 37 -2005 0 net=1210
rlabel metal2 229 -2005 229 -2005 0 net=1945
rlabel metal2 271 -2005 271 -2005 0 net=2292
rlabel metal2 387 -2005 387 -2005 0 net=1509
rlabel metal2 513 -2005 513 -2005 0 net=5206
rlabel metal2 639 -2005 639 -2005 0 net=6251
rlabel metal2 744 -2005 744 -2005 0 net=6054
rlabel metal2 37 -2007 37 -2007 0 net=3473
rlabel metal2 233 -2007 233 -2007 0 net=1788
rlabel metal2 247 -2007 247 -2007 0 net=3098
rlabel metal2 492 -2007 492 -2007 0 net=4505
rlabel metal2 569 -2007 569 -2007 0 net=187
rlabel metal2 44 -2009 44 -2009 0 net=3600
rlabel metal2 236 -2009 236 -2009 0 net=4871
rlabel metal2 555 -2009 555 -2009 0 net=5503
rlabel metal2 625 -2009 625 -2009 0 net=5771
rlabel metal2 625 -2009 625 -2009 0 net=5771
rlabel metal2 660 -2009 660 -2009 0 net=6576
rlabel metal2 744 -2009 744 -2009 0 net=6827
rlabel metal2 758 -2009 758 -2009 0 net=6841
rlabel metal2 44 -2011 44 -2011 0 net=5153
rlabel metal2 149 -2011 149 -2011 0 net=3587
rlabel metal2 191 -2011 191 -2011 0 net=2017
rlabel metal2 247 -2011 247 -2011 0 net=1255
rlabel metal2 264 -2011 264 -2011 0 net=5969
rlabel metal2 653 -2011 653 -2011 0 net=5809
rlabel metal2 674 -2011 674 -2011 0 net=5973
rlabel metal2 751 -2011 751 -2011 0 net=6887
rlabel metal2 51 -2013 51 -2013 0 net=5424
rlabel metal2 170 -2013 170 -2013 0 net=1367
rlabel metal2 275 -2013 275 -2013 0 net=1425
rlabel metal2 275 -2013 275 -2013 0 net=1425
rlabel metal2 289 -2013 289 -2013 0 net=1944
rlabel metal2 359 -2013 359 -2013 0 net=4713
rlabel metal2 380 -2013 380 -2013 0 net=3245
rlabel metal2 464 -2013 464 -2013 0 net=5913
rlabel metal2 688 -2013 688 -2013 0 net=6799
rlabel metal2 758 -2013 758 -2013 0 net=6119
rlabel metal2 51 -2015 51 -2015 0 net=5727
rlabel metal2 593 -2015 593 -2015 0 net=5018
rlabel metal2 58 -2017 58 -2017 0 net=2140
rlabel metal2 289 -2017 289 -2017 0 net=1337
rlabel metal2 352 -2017 352 -2017 0 net=2578
rlabel metal2 464 -2017 464 -2017 0 net=3655
rlabel metal2 562 -2017 562 -2017 0 net=4571
rlabel metal2 691 -2017 691 -2017 0 net=6638
rlabel metal2 58 -2019 58 -2019 0 net=5709
rlabel metal2 191 -2019 191 -2019 0 net=1271
rlabel metal2 243 -2019 243 -2019 0 net=1552
rlabel metal2 292 -2019 292 -2019 0 net=568
rlabel metal2 471 -2019 471 -2019 0 net=5749
rlabel metal2 716 -2019 716 -2019 0 net=6493
rlabel metal2 65 -2021 65 -2021 0 net=5328
rlabel metal2 296 -2021 296 -2021 0 net=2565
rlabel metal2 373 -2021 373 -2021 0 net=3281
rlabel metal2 565 -2021 565 -2021 0 net=6557
rlabel metal2 65 -2023 65 -2023 0 net=4281
rlabel metal2 583 -2023 583 -2023 0 net=710
rlabel metal2 709 -2023 709 -2023 0 net=6439
rlabel metal2 72 -2025 72 -2025 0 net=4916
rlabel metal2 163 -2025 163 -2025 0 net=3357
rlabel metal2 303 -2025 303 -2025 0 net=4397
rlabel metal2 450 -2025 450 -2025 0 net=3363
rlabel metal2 681 -2025 681 -2025 0 net=6127
rlabel metal2 72 -2027 72 -2027 0 net=3383
rlabel metal2 107 -2027 107 -2027 0 net=2827
rlabel metal2 303 -2027 303 -2027 0 net=2023
rlabel metal2 541 -2027 541 -2027 0 net=4899
rlabel metal2 667 -2027 667 -2027 0 net=6037
rlabel metal2 79 -2029 79 -2029 0 net=2463
rlabel metal2 324 -2029 324 -2029 0 net=2691
rlabel metal2 401 -2029 401 -2029 0 net=3775
rlabel metal2 86 -2031 86 -2031 0 net=2339
rlabel metal2 219 -2031 219 -2031 0 net=1901
rlabel metal2 317 -2031 317 -2031 0 net=3331
rlabel metal2 527 -2031 527 -2031 0 net=4131
rlabel metal2 583 -2031 583 -2031 0 net=5027
rlabel metal2 646 -2031 646 -2031 0 net=6377
rlabel metal2 86 -2033 86 -2033 0 net=3193
rlabel metal2 590 -2033 590 -2033 0 net=3575
rlabel metal2 100 -2035 100 -2035 0 net=1935
rlabel metal2 128 -2035 128 -2035 0 net=3367
rlabel metal2 261 -2035 261 -2035 0 net=6813
rlabel metal2 611 -2035 611 -2035 0 net=5075
rlabel metal2 23 -2037 23 -2037 0 net=5425
rlabel metal2 205 -2037 205 -2037 0 net=1373
rlabel metal2 261 -2037 261 -2037 0 net=2779
rlabel metal2 394 -2037 394 -2037 0 net=6907
rlabel metal2 114 -2039 114 -2039 0 net=1655
rlabel metal2 205 -2039 205 -2039 0 net=3139
rlabel metal2 457 -2039 457 -2039 0 net=5922
rlabel metal2 93 -2041 93 -2041 0 net=1661
rlabel metal2 331 -2041 331 -2041 0 net=2635
rlabel metal2 408 -2041 408 -2041 0 net=2909
rlabel metal2 418 -2041 418 -2041 0 net=4925
rlabel metal2 121 -2043 121 -2043 0 net=1146
rlabel metal2 338 -2043 338 -2043 0 net=2829
rlabel metal2 345 -2045 345 -2045 0 net=1121
rlabel metal2 506 -2045 506 -2045 0 net=4835
rlabel metal2 415 -2047 415 -2047 0 net=4178
rlabel metal2 422 -2049 422 -2049 0 net=3667
rlabel metal2 429 -2051 429 -2051 0 net=4183
rlabel metal2 478 -2051 478 -2051 0 net=3029
rlabel metal2 485 -2053 485 -2053 0 net=3947
rlabel metal2 23 -2064 23 -2064 0 net=5426
rlabel metal2 411 -2064 411 -2064 0 net=380
rlabel metal2 534 -2064 534 -2064 0 net=3949
rlabel metal2 541 -2064 541 -2064 0 net=4132
rlabel metal2 611 -2064 611 -2064 0 net=5077
rlabel metal2 611 -2064 611 -2064 0 net=5077
rlabel metal2 653 -2064 653 -2064 0 net=6559
rlabel metal2 23 -2066 23 -2066 0 net=1331
rlabel metal2 254 -2066 254 -2066 0 net=1902
rlabel metal2 292 -2066 292 -2066 0 net=2566
rlabel metal2 373 -2066 373 -2066 0 net=3283
rlabel metal2 418 -2066 418 -2066 0 net=3030
rlabel metal2 534 -2066 534 -2066 0 net=5505
rlabel metal2 569 -2066 569 -2066 0 net=5970
rlabel metal2 667 -2066 667 -2066 0 net=6039
rlabel metal2 723 -2066 723 -2066 0 net=6120
rlabel metal2 30 -2068 30 -2068 0 net=5148
rlabel metal2 184 -2068 184 -2068 0 net=322
rlabel metal2 240 -2068 240 -2068 0 net=1427
rlabel metal2 345 -2068 345 -2068 0 net=3668
rlabel metal2 436 -2068 436 -2068 0 net=4399
rlabel metal2 569 -2068 569 -2068 0 net=5029
rlabel metal2 632 -2068 632 -2068 0 net=6379
rlabel metal2 670 -2068 670 -2068 0 net=6842
rlabel metal2 30 -2070 30 -2070 0 net=6187
rlabel metal2 474 -2070 474 -2070 0 net=4572
rlabel metal2 646 -2070 646 -2070 0 net=6495
rlabel metal2 37 -2072 37 -2072 0 net=3474
rlabel metal2 257 -2072 257 -2072 0 net=4681
rlabel metal2 443 -2072 443 -2072 0 net=4185
rlabel metal2 443 -2072 443 -2072 0 net=4185
rlabel metal2 457 -2072 457 -2072 0 net=4468
rlabel metal2 44 -2074 44 -2074 0 net=5154
rlabel metal2 212 -2074 212 -2074 0 net=3369
rlabel metal2 296 -2074 296 -2074 0 net=3359
rlabel metal2 457 -2074 457 -2074 0 net=5793
rlabel metal2 618 -2074 618 -2074 0 net=5811
rlabel metal2 681 -2074 681 -2074 0 net=6909
rlabel metal2 44 -2076 44 -2076 0 net=1369
rlabel metal2 212 -2076 212 -2076 0 net=1307
rlabel metal2 352 -2076 352 -2076 0 net=70
rlabel metal2 660 -2076 660 -2076 0 net=5915
rlabel metal2 709 -2076 709 -2076 0 net=6129
rlabel metal2 726 -2076 726 -2076 0 net=3475
rlabel metal2 51 -2078 51 -2078 0 net=5728
rlabel metal2 135 -2078 135 -2078 0 net=2340
rlabel metal2 219 -2078 219 -2078 0 net=1375
rlabel metal2 275 -2078 275 -2078 0 net=2919
rlabel metal2 324 -2078 324 -2078 0 net=2693
rlabel metal2 373 -2078 373 -2078 0 net=2631
rlabel metal2 488 -2078 488 -2078 0 net=4506
rlabel metal2 499 -2078 499 -2078 0 net=3577
rlabel metal2 709 -2078 709 -2078 0 net=6889
rlabel metal2 51 -2080 51 -2080 0 net=3589
rlabel metal2 268 -2080 268 -2080 0 net=1947
rlabel metal2 317 -2080 317 -2080 0 net=3333
rlabel metal2 359 -2080 359 -2080 0 net=4715
rlabel metal2 492 -2080 492 -2080 0 net=4873
rlabel metal2 562 -2080 562 -2080 0 net=4901
rlabel metal2 58 -2082 58 -2082 0 net=5710
rlabel metal2 135 -2082 135 -2082 0 net=2830
rlabel metal2 380 -2082 380 -2082 0 net=3246
rlabel metal2 464 -2082 464 -2082 0 net=3656
rlabel metal2 527 -2082 527 -2082 0 net=6815
rlabel metal2 58 -2084 58 -2084 0 net=3817
rlabel metal2 142 -2084 142 -2084 0 net=644
rlabel metal2 366 -2084 366 -2084 0 net=3839
rlabel metal2 474 -2084 474 -2084 0 net=5596
rlabel metal2 65 -2086 65 -2086 0 net=4282
rlabel metal2 142 -2086 142 -2086 0 net=1961
rlabel metal2 233 -2086 233 -2086 0 net=5565
rlabel metal2 296 -2086 296 -2086 0 net=2637
rlabel metal2 338 -2086 338 -2086 0 net=3723
rlabel metal2 478 -2086 478 -2086 0 net=5750
rlabel metal2 65 -2088 65 -2088 0 net=2569
rlabel metal2 317 -2088 317 -2088 0 net=5755
rlabel metal2 688 -2088 688 -2088 0 net=6801
rlabel metal2 72 -2090 72 -2090 0 net=3384
rlabel metal2 107 -2090 107 -2090 0 net=2828
rlabel metal2 233 -2090 233 -2090 0 net=1339
rlabel metal2 331 -2090 331 -2090 0 net=1511
rlabel metal2 415 -2090 415 -2090 0 net=3365
rlabel metal2 460 -2090 460 -2090 0 net=3776
rlabel metal2 72 -2092 72 -2092 0 net=2781
rlabel metal2 320 -2092 320 -2092 0 net=4573
rlabel metal2 478 -2092 478 -2092 0 net=4419
rlabel metal2 520 -2092 520 -2092 0 net=4837
rlabel metal2 576 -2092 576 -2092 0 net=5773
rlabel metal2 688 -2092 688 -2092 0 net=6441
rlabel metal2 79 -2094 79 -2094 0 net=2464
rlabel metal2 506 -2094 506 -2094 0 net=5763
rlabel metal2 625 -2094 625 -2094 0 net=6253
rlabel metal2 716 -2094 716 -2094 0 net=6829
rlabel metal2 79 -2096 79 -2096 0 net=3537
rlabel metal2 247 -2096 247 -2096 0 net=1256
rlabel metal2 387 -2096 387 -2096 0 net=2805
rlabel metal2 520 -2096 520 -2096 0 net=4927
rlabel metal2 86 -2098 86 -2098 0 net=3194
rlabel metal2 261 -2098 261 -2098 0 net=1981
rlabel metal2 604 -2098 604 -2098 0 net=5975
rlabel metal2 86 -2100 86 -2100 0 net=2159
rlabel metal2 100 -2100 100 -2100 0 net=1937
rlabel metal2 114 -2100 114 -2100 0 net=1657
rlabel metal2 114 -2100 114 -2100 0 net=1657
rlabel metal2 121 -2100 121 -2100 0 net=2025
rlabel metal2 394 -2100 394 -2100 0 net=6685
rlabel metal2 93 -2102 93 -2102 0 net=1662
rlabel metal2 303 -2102 303 -2102 0 net=1515
rlabel metal2 394 -2102 394 -2102 0 net=2911
rlabel metal2 16 -2104 16 -2104 0 net=5870
rlabel metal2 128 -2104 128 -2104 0 net=5059
rlabel metal2 149 -2106 149 -2106 0 net=1273
rlabel metal2 163 -2108 163 -2108 0 net=221
rlabel metal2 156 -2110 156 -2110 0 net=2175
rlabel metal2 180 -2110 180 -2110 0 net=6651
rlabel metal2 180 -2112 180 -2112 0 net=2018
rlabel metal2 191 -2114 191 -2114 0 net=3141
rlabel metal2 16 -2116 16 -2116 0 net=6329
rlabel metal2 198 -2118 198 -2118 0 net=705
rlabel metal2 16 -2129 16 -2129 0 net=6330
rlabel metal2 506 -2129 506 -2129 0 net=6254
rlabel metal2 632 -2129 632 -2129 0 net=6381
rlabel metal2 632 -2129 632 -2129 0 net=6381
rlabel metal2 688 -2129 688 -2129 0 net=6442
rlabel metal2 40 -2131 40 -2131 0 net=444
rlabel metal2 163 -2131 163 -2131 0 net=2176
rlabel metal2 184 -2131 184 -2131 0 net=1377
rlabel metal2 261 -2131 261 -2131 0 net=1982
rlabel metal2 457 -2131 457 -2131 0 net=3891
rlabel metal2 695 -2131 695 -2131 0 net=6652
rlabel metal2 44 -2133 44 -2133 0 net=1370
rlabel metal2 254 -2133 254 -2133 0 net=3725
rlabel metal2 345 -2133 345 -2133 0 net=5756
rlabel metal2 625 -2133 625 -2133 0 net=6891
rlabel metal2 51 -2135 51 -2135 0 net=3590
rlabel metal2 226 -2135 226 -2135 0 net=1428
rlabel metal2 261 -2135 261 -2135 0 net=2695
rlabel metal2 359 -2135 359 -2135 0 net=4683
rlabel metal2 436 -2135 436 -2135 0 net=3767
rlabel metal2 509 -2135 509 -2135 0 net=5060
rlabel metal2 558 -2135 558 -2135 0 net=6830
rlabel metal2 58 -2137 58 -2137 0 net=3818
rlabel metal2 121 -2137 121 -2137 0 net=2027
rlabel metal2 268 -2137 268 -2137 0 net=5567
rlabel metal2 348 -2137 348 -2137 0 net=216
rlabel metal2 439 -2137 439 -2137 0 net=5078
rlabel metal2 660 -2137 660 -2137 0 net=5917
rlabel metal2 65 -2139 65 -2139 0 net=2570
rlabel metal2 324 -2139 324 -2139 0 net=3335
rlabel metal2 380 -2139 380 -2139 0 net=2912
rlabel metal2 408 -2139 408 -2139 0 net=4400
rlabel metal2 534 -2139 534 -2139 0 net=5507
rlabel metal2 72 -2141 72 -2141 0 net=2782
rlabel metal2 362 -2141 362 -2141 0 net=6155
rlabel metal2 390 -2141 390 -2141 0 net=4874
rlabel metal2 513 -2141 513 -2141 0 net=4929
rlabel metal2 541 -2141 541 -2141 0 net=5765
rlabel metal2 579 -2141 579 -2141 0 net=6802
rlabel metal2 86 -2143 86 -2143 0 net=2161
rlabel metal2 86 -2143 86 -2143 0 net=2161
rlabel metal2 100 -2143 100 -2143 0 net=1659
rlabel metal2 128 -2143 128 -2143 0 net=465
rlabel metal2 170 -2143 170 -2143 0 net=3366
rlabel metal2 464 -2143 464 -2143 0 net=4902
rlabel metal2 583 -2143 583 -2143 0 net=5795
rlabel metal2 593 -2143 593 -2143 0 net=471
rlabel metal2 30 -2145 30 -2145 0 net=6188
rlabel metal2 135 -2145 135 -2145 0 net=1541
rlabel metal2 198 -2145 198 -2145 0 net=4574
rlabel metal2 464 -2145 464 -2145 0 net=3579
rlabel metal2 520 -2145 520 -2145 0 net=4839
rlabel metal2 548 -2145 548 -2145 0 net=5031
rlabel metal2 597 -2145 597 -2145 0 net=5977
rlabel metal2 611 -2145 611 -2145 0 net=6561
rlabel metal2 107 -2147 107 -2147 0 net=1938
rlabel metal2 142 -2147 142 -2147 0 net=1962
rlabel metal2 198 -2147 198 -2147 0 net=3757
rlabel metal2 226 -2147 226 -2147 0 net=3091
rlabel metal2 282 -2147 282 -2147 0 net=3371
rlabel metal2 296 -2147 296 -2147 0 net=2639
rlabel metal2 373 -2147 373 -2147 0 net=2633
rlabel metal2 408 -2147 408 -2147 0 net=5195
rlabel metal2 555 -2147 555 -2147 0 net=3951
rlabel metal2 23 -2149 23 -2149 0 net=1332
rlabel metal2 170 -2149 170 -2149 0 net=2237
rlabel metal2 604 -2149 604 -2149 0 net=5813
rlabel metal2 639 -2149 639 -2149 0 net=6687
rlabel metal2 107 -2151 107 -2151 0 net=3669
rlabel metal2 201 -2151 201 -2151 0 net=2920
rlabel metal2 282 -2151 282 -2151 0 net=4039
rlabel metal2 331 -2151 331 -2151 0 net=1512
rlabel metal2 471 -2151 471 -2151 0 net=5379
rlabel metal2 639 -2151 639 -2151 0 net=6911
rlabel metal2 114 -2153 114 -2153 0 net=1865
rlabel metal2 296 -2153 296 -2153 0 net=2806
rlabel metal2 443 -2153 443 -2153 0 net=4187
rlabel metal2 485 -2153 485 -2153 0 net=4717
rlabel metal2 646 -2153 646 -2153 0 net=6497
rlabel metal2 121 -2155 121 -2155 0 net=4989
rlabel metal2 443 -2155 443 -2155 0 net=4421
rlabel metal2 499 -2155 499 -2155 0 net=6077
rlabel metal2 646 -2155 646 -2155 0 net=6817
rlabel metal2 142 -2157 142 -2157 0 net=1341
rlabel metal2 275 -2157 275 -2157 0 net=1517
rlabel metal2 313 -2157 313 -2157 0 net=3476
rlabel metal2 149 -2159 149 -2159 0 net=1274
rlabel metal2 212 -2159 212 -2159 0 net=1309
rlabel metal2 303 -2159 303 -2159 0 net=1949
rlabel metal2 331 -2159 331 -2159 0 net=5549
rlabel metal2 667 -2159 667 -2159 0 net=6041
rlabel metal2 79 -2161 79 -2161 0 net=3538
rlabel metal2 219 -2161 219 -2161 0 net=5781
rlabel metal2 478 -2161 478 -2161 0 net=4311
rlabel metal2 667 -2161 667 -2161 0 net=6130
rlabel metal2 156 -2163 156 -2163 0 net=605
rlabel metal2 366 -2163 366 -2163 0 net=3841
rlabel metal2 576 -2163 576 -2163 0 net=5775
rlabel metal2 177 -2165 177 -2165 0 net=2801
rlabel metal2 191 -2165 191 -2165 0 net=3143
rlabel metal2 222 -2165 222 -2165 0 net=3481
rlabel metal2 366 -2165 366 -2165 0 net=3361
rlabel metal2 191 -2167 191 -2167 0 net=1481
rlabel metal2 373 -2167 373 -2167 0 net=3285
rlabel metal2 422 -2167 422 -2167 0 net=6325
rlabel metal2 250 -2169 250 -2169 0 net=5337
rlabel metal2 86 -2180 86 -2180 0 net=2162
rlabel metal2 107 -2180 107 -2180 0 net=3671
rlabel metal2 107 -2180 107 -2180 0 net=3671
rlabel metal2 114 -2180 114 -2180 0 net=1866
rlabel metal2 380 -2180 380 -2180 0 net=6156
rlabel metal2 506 -2180 506 -2180 0 net=5551
rlabel metal2 534 -2180 534 -2180 0 net=5196
rlabel metal2 674 -2180 674 -2180 0 net=6042
rlabel metal2 114 -2182 114 -2182 0 net=1379
rlabel metal2 191 -2182 191 -2182 0 net=1483
rlabel metal2 191 -2182 191 -2182 0 net=1483
rlabel metal2 205 -2182 205 -2182 0 net=3144
rlabel metal2 222 -2182 222 -2182 0 net=224
rlabel metal2 579 -2182 579 -2182 0 net=5776
rlabel metal2 121 -2184 121 -2184 0 net=4991
rlabel metal2 163 -2184 163 -2184 0 net=1543
rlabel metal2 205 -2184 205 -2184 0 net=790
rlabel metal2 324 -2184 324 -2184 0 net=4041
rlabel metal2 401 -2184 401 -2184 0 net=5338
rlabel metal2 492 -2184 492 -2184 0 net=6073
rlabel metal2 569 -2184 569 -2184 0 net=5918
rlabel metal2 124 -2186 124 -2186 0 net=3726
rlabel metal2 275 -2186 275 -2186 0 net=1519
rlabel metal2 275 -2186 275 -2186 0 net=1519
rlabel metal2 282 -2186 282 -2186 0 net=3362
rlabel metal2 401 -2186 401 -2186 0 net=6327
rlabel metal2 425 -2186 425 -2186 0 net=5380
rlabel metal2 583 -2186 583 -2186 0 net=3892
rlabel metal2 128 -2188 128 -2188 0 net=1106
rlabel metal2 429 -2188 429 -2188 0 net=4718
rlabel metal2 639 -2188 639 -2188 0 net=6912
rlabel metal2 142 -2190 142 -2190 0 net=1343
rlabel metal2 233 -2190 233 -2190 0 net=1311
rlabel metal2 233 -2190 233 -2190 0 net=1311
rlabel metal2 240 -2190 240 -2190 0 net=4930
rlabel metal2 555 -2190 555 -2190 0 net=6562
rlabel metal2 170 -2192 170 -2192 0 net=2239
rlabel metal2 243 -2192 243 -2192 0 net=3219
rlabel metal2 285 -2192 285 -2192 0 net=680
rlabel metal2 394 -2192 394 -2192 0 net=2634
rlabel metal2 569 -2192 569 -2192 0 net=6781
rlabel metal2 142 -2194 142 -2194 0 net=3647
rlabel metal2 198 -2194 198 -2194 0 net=3759
rlabel metal2 408 -2194 408 -2194 0 net=4423
rlabel metal2 450 -2194 450 -2194 0 net=3580
rlabel metal2 499 -2194 499 -2194 0 net=6079
rlabel metal2 555 -2194 555 -2194 0 net=6383
rlabel metal2 212 -2196 212 -2196 0 net=5568
rlabel metal2 366 -2196 366 -2196 0 net=3287
rlabel metal2 387 -2196 387 -2196 0 net=721
rlabel metal2 513 -2196 513 -2196 0 net=5033
rlabel metal2 583 -2196 583 -2196 0 net=6499
rlabel metal2 152 -2198 152 -2198 0 net=4923
rlabel metal2 285 -2198 285 -2198 0 net=5105
rlabel metal2 548 -2198 548 -2198 0 net=5797
rlabel metal2 597 -2198 597 -2198 0 net=5979
rlabel metal2 296 -2200 296 -2200 0 net=1671
rlabel metal2 632 -2200 632 -2200 0 net=3953
rlabel metal2 317 -2202 317 -2202 0 net=3483
rlabel metal2 415 -2202 415 -2202 0 net=5783
rlabel metal2 586 -2202 586 -2202 0 net=5814
rlabel metal2 317 -2204 317 -2204 0 net=4189
rlabel metal2 509 -2204 509 -2204 0 net=983
rlabel metal2 324 -2206 324 -2206 0 net=3337
rlabel metal2 359 -2206 359 -2206 0 net=4685
rlabel metal2 429 -2206 429 -2206 0 net=4313
rlabel metal2 590 -2206 590 -2206 0 net=6893
rlabel metal2 268 -2208 268 -2208 0 net=3093
rlabel metal2 432 -2208 432 -2208 0 net=6267
rlabel metal2 478 -2208 478 -2208 0 net=6297
rlabel metal2 268 -2210 268 -2210 0 net=2935
rlabel metal2 331 -2210 331 -2210 0 net=6179
rlabel metal2 485 -2210 485 -2210 0 net=3842
rlabel metal2 261 -2212 261 -2212 0 net=2697
rlabel metal2 436 -2212 436 -2212 0 net=3769
rlabel metal2 597 -2212 597 -2212 0 net=6819
rlabel metal2 261 -2214 261 -2214 0 net=2641
rlabel metal2 390 -2214 390 -2214 0 net=5319
rlabel metal2 485 -2214 485 -2214 0 net=4841
rlabel metal2 156 -2216 156 -2216 0 net=1639
rlabel metal2 520 -2216 520 -2216 0 net=5767
rlabel metal2 156 -2218 156 -2218 0 net=2803
rlabel metal2 289 -2218 289 -2218 0 net=3373
rlabel metal2 541 -2218 541 -2218 0 net=6689
rlabel metal2 131 -2220 131 -2220 0 net=145
rlabel metal2 247 -2220 247 -2220 0 net=2029
rlabel metal2 660 -2220 660 -2220 0 net=5509
rlabel metal2 100 -2222 100 -2222 0 net=1660
rlabel metal2 247 -2222 247 -2222 0 net=1951
rlabel metal2 107 -2233 107 -2233 0 net=3672
rlabel metal2 275 -2233 275 -2233 0 net=1520
rlabel metal2 289 -2233 289 -2233 0 net=2031
rlabel metal2 289 -2233 289 -2233 0 net=2031
rlabel metal2 306 -2233 306 -2233 0 net=6298
rlabel metal2 499 -2233 499 -2233 0 net=5785
rlabel metal2 499 -2233 499 -2233 0 net=5785
rlabel metal2 534 -2233 534 -2233 0 net=3770
rlabel metal2 639 -2233 639 -2233 0 net=5981
rlabel metal2 639 -2233 639 -2233 0 net=5981
rlabel metal2 114 -2235 114 -2235 0 net=1380
rlabel metal2 198 -2235 198 -2235 0 net=2335
rlabel metal2 254 -2235 254 -2235 0 net=3221
rlabel metal2 313 -2235 313 -2235 0 net=6328
rlabel metal2 415 -2235 415 -2235 0 net=4686
rlabel metal2 443 -2235 443 -2235 0 net=3695
rlabel metal2 527 -2235 527 -2235 0 net=6081
rlabel metal2 548 -2235 548 -2235 0 net=5799
rlabel metal2 548 -2235 548 -2235 0 net=5799
rlabel metal2 562 -2235 562 -2235 0 net=6894
rlabel metal2 607 -2235 607 -2235 0 net=5510
rlabel metal2 114 -2237 114 -2237 0 net=3649
rlabel metal2 149 -2237 149 -2237 0 net=4993
rlabel metal2 173 -2237 173 -2237 0 net=1484
rlabel metal2 201 -2237 201 -2237 0 net=4924
rlabel metal2 219 -2237 219 -2237 0 net=1345
rlabel metal2 317 -2237 317 -2237 0 net=4191
rlabel metal2 317 -2237 317 -2237 0 net=4191
rlabel metal2 324 -2237 324 -2237 0 net=3338
rlabel metal2 366 -2237 366 -2237 0 net=3288
rlabel metal2 390 -2237 390 -2237 0 net=4885
rlabel metal2 422 -2237 422 -2237 0 net=4315
rlabel metal2 446 -2237 446 -2237 0 net=6690
rlabel metal2 565 -2237 565 -2237 0 net=3954
rlabel metal2 121 -2239 121 -2239 0 net=586
rlabel metal2 128 -2239 128 -2239 0 net=520
rlabel metal2 149 -2239 149 -2239 0 net=1100
rlabel metal2 212 -2239 212 -2239 0 net=3683
rlabel metal2 261 -2239 261 -2239 0 net=2642
rlabel metal2 327 -2239 327 -2239 0 net=434
rlabel metal2 366 -2239 366 -2239 0 net=4043
rlabel metal2 397 -2239 397 -2239 0 net=6180
rlabel metal2 513 -2239 513 -2239 0 net=5035
rlabel metal2 583 -2239 583 -2239 0 net=6501
rlabel metal2 583 -2239 583 -2239 0 net=6501
rlabel metal2 124 -2241 124 -2241 0 net=798
rlabel metal2 156 -2241 156 -2241 0 net=2804
rlabel metal2 205 -2241 205 -2241 0 net=6727
rlabel metal2 331 -2241 331 -2241 0 net=2698
rlabel metal2 401 -2241 401 -2241 0 net=4425
rlabel metal2 457 -2241 457 -2241 0 net=6269
rlabel metal2 457 -2241 457 -2241 0 net=6269
rlabel metal2 464 -2241 464 -2241 0 net=5768
rlabel metal2 527 -2241 527 -2241 0 net=6385
rlabel metal2 131 -2243 131 -2243 0 net=2747
rlabel metal2 156 -2243 156 -2243 0 net=5375
rlabel metal2 261 -2243 261 -2243 0 net=4219
rlabel metal2 467 -2243 467 -2243 0 net=5552
rlabel metal2 513 -2243 513 -2243 0 net=6423
rlabel metal2 163 -2245 163 -2245 0 net=2936
rlabel metal2 296 -2245 296 -2245 0 net=1673
rlabel metal2 338 -2245 338 -2245 0 net=1640
rlabel metal2 576 -2245 576 -2245 0 net=6821
rlabel metal2 163 -2247 163 -2247 0 net=4169
rlabel metal2 247 -2247 247 -2247 0 net=1953
rlabel metal2 310 -2247 310 -2247 0 net=3375
rlabel metal2 345 -2247 345 -2247 0 net=3485
rlabel metal2 492 -2247 492 -2247 0 net=6075
rlabel metal2 555 -2247 555 -2247 0 net=6783
rlabel metal2 166 -2249 166 -2249 0 net=433
rlabel metal2 485 -2249 485 -2249 0 net=4843
rlabel metal2 506 -2249 506 -2249 0 net=2951
rlabel metal2 177 -2251 177 -2251 0 net=1545
rlabel metal2 240 -2251 240 -2251 0 net=2241
rlabel metal2 268 -2251 268 -2251 0 net=4049
rlabel metal2 303 -2251 303 -2251 0 net=5759
rlabel metal2 359 -2251 359 -2251 0 net=6095
rlabel metal2 184 -2253 184 -2253 0 net=3027
rlabel metal2 373 -2253 373 -2253 0 net=5320
rlabel metal2 352 -2255 352 -2255 0 net=3094
rlabel metal2 394 -2255 394 -2255 0 net=3761
rlabel metal2 226 -2257 226 -2257 0 net=6227
rlabel metal2 380 -2257 380 -2257 0 net=3885
rlabel metal2 436 -2257 436 -2257 0 net=5107
rlabel metal2 226 -2259 226 -2259 0 net=1313
rlabel metal2 303 -2259 303 -2259 0 net=1903
rlabel metal2 114 -2270 114 -2270 0 net=3650
rlabel metal2 135 -2270 135 -2270 0 net=2748
rlabel metal2 163 -2270 163 -2270 0 net=4170
rlabel metal2 317 -2270 317 -2270 0 net=4192
rlabel metal2 380 -2270 380 -2270 0 net=3887
rlabel metal2 380 -2270 380 -2270 0 net=3887
rlabel metal2 401 -2270 401 -2270 0 net=4426
rlabel metal2 450 -2270 450 -2270 0 net=1904
rlabel metal2 639 -2270 639 -2270 0 net=5983
rlabel metal2 639 -2270 639 -2270 0 net=5983
rlabel metal2 121 -2272 121 -2272 0 net=971
rlabel metal2 142 -2272 142 -2272 0 net=5376
rlabel metal2 170 -2272 170 -2272 0 net=4994
rlabel metal2 215 -2272 215 -2272 0 net=901
rlabel metal2 240 -2272 240 -2272 0 net=1135
rlabel metal2 254 -2272 254 -2272 0 net=1347
rlabel metal2 254 -2272 254 -2272 0 net=1347
rlabel metal2 275 -2272 275 -2272 0 net=3222
rlabel metal2 289 -2272 289 -2272 0 net=2033
rlabel metal2 345 -2272 345 -2272 0 net=5761
rlabel metal2 345 -2272 345 -2272 0 net=5761
rlabel metal2 352 -2272 352 -2272 0 net=6228
rlabel metal2 404 -2272 404 -2272 0 net=4886
rlabel metal2 422 -2272 422 -2272 0 net=4317
rlabel metal2 422 -2272 422 -2272 0 net=4317
rlabel metal2 429 -2272 429 -2272 0 net=940
rlabel metal2 541 -2272 541 -2272 0 net=5036
rlabel metal2 177 -2274 177 -2274 0 net=1547
rlabel metal2 177 -2274 177 -2274 0 net=1547
rlabel metal2 184 -2274 184 -2274 0 net=3028
rlabel metal2 243 -2274 243 -2274 0 net=3696
rlabel metal2 485 -2274 485 -2274 0 net=3762
rlabel metal2 534 -2274 534 -2274 0 net=6083
rlabel metal2 548 -2274 548 -2274 0 net=5800
rlabel metal2 548 -2274 548 -2274 0 net=5800
rlabel metal2 198 -2276 198 -2276 0 net=2336
rlabel metal2 359 -2276 359 -2276 0 net=3486
rlabel metal2 471 -2276 471 -2276 0 net=5786
rlabel metal2 534 -2276 534 -2276 0 net=6784
rlabel metal2 212 -2278 212 -2278 0 net=3685
rlabel metal2 226 -2278 226 -2278 0 net=1315
rlabel metal2 261 -2278 261 -2278 0 net=4221
rlabel metal2 289 -2278 289 -2278 0 net=2839
rlabel metal2 408 -2278 408 -2278 0 net=6076
rlabel metal2 205 -2280 205 -2280 0 net=6729
rlabel metal2 268 -2280 268 -2280 0 net=4051
rlabel metal2 296 -2280 296 -2280 0 net=1955
rlabel metal2 296 -2280 296 -2280 0 net=1955
rlabel metal2 303 -2280 303 -2280 0 net=1674
rlabel metal2 415 -2280 415 -2280 0 net=5109
rlabel metal2 457 -2280 457 -2280 0 net=6271
rlabel metal2 474 -2280 474 -2280 0 net=1172
rlabel metal2 513 -2280 513 -2280 0 net=6425
rlabel metal2 247 -2282 247 -2282 0 net=2243
rlabel metal2 303 -2282 303 -2282 0 net=4044
rlabel metal2 432 -2282 432 -2282 0 net=2952
rlabel metal2 513 -2282 513 -2282 0 net=6387
rlabel metal2 331 -2284 331 -2284 0 net=3377
rlabel metal2 362 -2284 362 -2284 0 net=1323
rlabel metal2 443 -2284 443 -2284 0 net=6097
rlabel metal2 492 -2284 492 -2284 0 net=4845
rlabel metal2 527 -2284 527 -2284 0 net=6822
rlabel metal2 450 -2286 450 -2286 0 net=6477
rlabel metal2 576 -2286 576 -2286 0 net=6503
rlabel metal2 177 -2297 177 -2297 0 net=1549
rlabel metal2 177 -2297 177 -2297 0 net=1549
rlabel metal2 212 -2297 212 -2297 0 net=3686
rlabel metal2 226 -2297 226 -2297 0 net=6730
rlabel metal2 247 -2297 247 -2297 0 net=1349
rlabel metal2 275 -2297 275 -2297 0 net=4222
rlabel metal2 338 -2297 338 -2297 0 net=5762
rlabel metal2 366 -2297 366 -2297 0 net=1324
rlabel metal2 380 -2297 380 -2297 0 net=3889
rlabel metal2 380 -2297 380 -2297 0 net=3889
rlabel metal2 408 -2297 408 -2297 0 net=5111
rlabel metal2 422 -2297 422 -2297 0 net=4318
rlabel metal2 443 -2297 443 -2297 0 net=6272
rlabel metal2 502 -2297 502 -2297 0 net=6388
rlabel metal2 520 -2297 520 -2297 0 net=6427
rlabel metal2 534 -2297 534 -2297 0 net=6084
rlabel metal2 569 -2297 569 -2297 0 net=6504
rlabel metal2 597 -2297 597 -2297 0 net=5467
rlabel metal2 639 -2297 639 -2297 0 net=5985
rlabel metal2 226 -2299 226 -2299 0 net=5855
rlabel metal2 282 -2299 282 -2299 0 net=4052
rlabel metal2 296 -2299 296 -2299 0 net=1956
rlabel metal2 313 -2299 313 -2299 0 net=2840
rlabel metal2 432 -2299 432 -2299 0 net=6098
rlabel metal2 506 -2299 506 -2299 0 net=4846
rlabel metal2 614 -2299 614 -2299 0 net=915
rlabel metal2 233 -2301 233 -2301 0 net=1317
rlabel metal2 233 -2301 233 -2301 0 net=1317
rlabel metal2 254 -2301 254 -2301 0 net=3777
rlabel metal2 289 -2301 289 -2301 0 net=2034
rlabel metal2 317 -2301 317 -2301 0 net=3379
rlabel metal2 446 -2301 446 -2301 0 net=6478
rlabel metal2 268 -2303 268 -2303 0 net=2245
rlabel metal2 170 -2314 170 -2314 0 net=1550
rlabel metal2 226 -2314 226 -2314 0 net=5856
rlabel metal2 296 -2314 296 -2314 0 net=2246
rlabel metal2 380 -2314 380 -2314 0 net=3890
rlabel metal2 404 -2314 404 -2314 0 net=5112
rlabel metal2 527 -2314 527 -2314 0 net=6428
rlabel metal2 597 -2314 597 -2314 0 net=5468
rlabel metal2 642 -2314 642 -2314 0 net=5986
rlabel metal2 233 -2316 233 -2316 0 net=1318
rlabel metal2 247 -2316 247 -2316 0 net=1350
rlabel metal2 278 -2316 278 -2316 0 net=3380
rlabel metal2 254 -2318 254 -2318 0 net=3778
<< end >>
