magic
tech scmos
timestamp 1555018107 
<< pdiffusion >>
rect 1 -20 7 -14
rect 8 -20 14 -14
rect 15 -20 21 -14
rect 22 -20 28 -14
rect 29 -20 35 -14
rect 36 -20 42 -14
rect 43 -20 49 -14
rect 50 -20 56 -14
rect 57 -20 63 -14
rect 64 -20 70 -14
rect 71 -20 77 -14
rect 78 -20 84 -14
rect 85 -20 91 -14
rect 92 -20 98 -14
rect 99 -20 105 -14
rect 106 -20 112 -14
rect 113 -20 119 -14
rect 120 -20 126 -14
rect 127 -20 133 -14
rect 134 -20 140 -14
rect 232 -20 235 -14
rect 344 -20 347 -14
rect 351 -20 357 -14
rect 358 -20 361 -14
rect 379 -20 382 -14
rect 400 -20 403 -14
rect 407 -20 410 -14
rect 414 -20 417 -14
rect 421 -20 424 -14
rect 428 -20 434 -14
rect 435 -20 441 -14
rect 442 -20 445 -14
rect 449 -20 455 -14
rect 456 -20 462 -14
rect 463 -20 469 -14
rect 470 -20 473 -14
rect 505 -20 511 -14
rect 526 -20 529 -14
rect 533 -20 539 -14
rect 547 -20 553 -14
rect 554 -20 557 -14
rect 603 -20 606 -14
rect 610 -20 616 -14
rect 652 -20 655 -14
rect 666 -20 672 -14
rect 673 -20 679 -14
rect 687 -20 690 -14
rect 715 -20 721 -14
rect 750 -20 756 -14
rect 799 -20 802 -14
rect 876 -20 882 -14
rect 953 -20 956 -14
rect 1 -57 7 -51
rect 8 -57 14 -51
rect 15 -57 21 -51
rect 22 -57 28 -51
rect 29 -57 35 -51
rect 36 -57 42 -51
rect 43 -57 49 -51
rect 50 -57 56 -51
rect 57 -57 63 -51
rect 64 -57 70 -51
rect 71 -57 77 -51
rect 78 -57 84 -51
rect 85 -57 91 -51
rect 92 -57 98 -51
rect 141 -57 147 -51
rect 148 -57 151 -51
rect 155 -57 158 -51
rect 225 -57 228 -51
rect 232 -57 238 -51
rect 260 -57 263 -51
rect 281 -57 284 -51
rect 302 -57 308 -51
rect 323 -57 326 -51
rect 330 -57 333 -51
rect 337 -57 340 -51
rect 372 -57 375 -51
rect 379 -57 382 -51
rect 386 -57 392 -51
rect 393 -57 396 -51
rect 400 -57 403 -51
rect 407 -57 413 -51
rect 414 -57 420 -51
rect 421 -57 427 -51
rect 428 -57 431 -51
rect 435 -57 438 -51
rect 442 -57 448 -51
rect 449 -57 452 -51
rect 456 -57 462 -51
rect 463 -57 466 -51
rect 470 -57 473 -51
rect 477 -57 480 -51
rect 491 -57 497 -51
rect 498 -57 501 -51
rect 505 -57 508 -51
rect 512 -57 518 -51
rect 519 -57 525 -51
rect 526 -57 532 -51
rect 533 -57 536 -51
rect 540 -57 543 -51
rect 547 -57 550 -51
rect 554 -57 557 -51
rect 561 -57 564 -51
rect 568 -57 574 -51
rect 575 -57 578 -51
rect 582 -57 585 -51
rect 589 -57 595 -51
rect 596 -57 599 -51
rect 603 -57 606 -51
rect 610 -57 613 -51
rect 617 -57 620 -51
rect 624 -57 627 -51
rect 631 -57 637 -51
rect 638 -57 641 -51
rect 645 -57 648 -51
rect 652 -57 655 -51
rect 659 -57 662 -51
rect 666 -57 669 -51
rect 673 -57 679 -51
rect 680 -57 683 -51
rect 687 -57 690 -51
rect 701 -57 704 -51
rect 708 -57 714 -51
rect 715 -57 718 -51
rect 729 -57 732 -51
rect 743 -57 746 -51
rect 757 -57 763 -51
rect 771 -57 774 -51
rect 813 -57 816 -51
rect 820 -57 823 -51
rect 827 -57 830 -51
rect 841 -57 844 -51
rect 883 -57 889 -51
rect 897 -57 900 -51
rect 932 -57 938 -51
rect 988 -57 991 -51
rect 995 -57 998 -51
rect 1 -104 7 -98
rect 8 -104 14 -98
rect 15 -104 21 -98
rect 22 -104 28 -98
rect 29 -104 35 -98
rect 36 -104 42 -98
rect 43 -104 49 -98
rect 50 -104 56 -98
rect 57 -104 63 -98
rect 64 -104 70 -98
rect 71 -104 77 -98
rect 78 -104 84 -98
rect 85 -104 91 -98
rect 92 -104 98 -98
rect 99 -104 105 -98
rect 106 -104 112 -98
rect 127 -104 130 -98
rect 148 -104 151 -98
rect 190 -104 193 -98
rect 197 -104 203 -98
rect 204 -104 207 -98
rect 218 -104 221 -98
rect 246 -104 252 -98
rect 253 -104 256 -98
rect 260 -104 263 -98
rect 267 -104 270 -98
rect 274 -104 277 -98
rect 281 -104 284 -98
rect 288 -104 294 -98
rect 295 -104 298 -98
rect 302 -104 305 -98
rect 309 -104 312 -98
rect 316 -104 319 -98
rect 323 -104 326 -98
rect 330 -104 336 -98
rect 337 -104 340 -98
rect 344 -104 347 -98
rect 351 -104 354 -98
rect 358 -104 361 -98
rect 365 -104 368 -98
rect 372 -104 378 -98
rect 379 -104 382 -98
rect 386 -104 389 -98
rect 393 -104 396 -98
rect 400 -104 403 -98
rect 407 -104 413 -98
rect 414 -104 417 -98
rect 421 -104 424 -98
rect 428 -104 434 -98
rect 435 -104 438 -98
rect 442 -104 445 -98
rect 449 -104 452 -98
rect 456 -104 462 -98
rect 463 -104 466 -98
rect 470 -104 476 -98
rect 477 -104 480 -98
rect 484 -104 490 -98
rect 491 -104 494 -98
rect 498 -104 501 -98
rect 505 -104 508 -98
rect 512 -104 515 -98
rect 519 -104 522 -98
rect 526 -104 532 -98
rect 533 -104 539 -98
rect 540 -104 543 -98
rect 547 -104 553 -98
rect 554 -104 557 -98
rect 561 -104 564 -98
rect 568 -104 571 -98
rect 575 -104 578 -98
rect 582 -104 585 -98
rect 589 -104 592 -98
rect 596 -104 599 -98
rect 603 -104 606 -98
rect 610 -104 613 -98
rect 617 -104 620 -98
rect 624 -104 627 -98
rect 631 -104 634 -98
rect 638 -104 641 -98
rect 645 -104 651 -98
rect 652 -104 655 -98
rect 659 -104 662 -98
rect 666 -104 669 -98
rect 673 -104 676 -98
rect 680 -104 683 -98
rect 687 -104 690 -98
rect 694 -104 697 -98
rect 701 -104 704 -98
rect 708 -104 711 -98
rect 715 -104 718 -98
rect 722 -104 725 -98
rect 729 -104 732 -98
rect 736 -104 739 -98
rect 743 -104 746 -98
rect 750 -104 753 -98
rect 778 -104 781 -98
rect 785 -104 788 -98
rect 792 -104 798 -98
rect 799 -104 802 -98
rect 806 -104 812 -98
rect 813 -104 819 -98
rect 820 -104 826 -98
rect 827 -104 830 -98
rect 834 -104 837 -98
rect 841 -104 844 -98
rect 855 -104 858 -98
rect 862 -104 865 -98
rect 869 -104 872 -98
rect 883 -104 889 -98
rect 890 -104 893 -98
rect 939 -104 942 -98
rect 946 -104 949 -98
rect 953 -104 956 -98
rect 1009 -104 1012 -98
rect 1086 -104 1089 -98
rect 1 -173 7 -167
rect 8 -173 14 -167
rect 15 -173 21 -167
rect 22 -173 28 -167
rect 29 -173 35 -167
rect 36 -173 42 -167
rect 43 -173 49 -167
rect 50 -173 56 -167
rect 57 -173 63 -167
rect 64 -173 70 -167
rect 71 -173 77 -167
rect 78 -173 84 -167
rect 92 -173 95 -167
rect 113 -173 116 -167
rect 134 -173 137 -167
rect 141 -173 144 -167
rect 148 -173 151 -167
rect 155 -173 158 -167
rect 162 -173 165 -167
rect 169 -173 172 -167
rect 176 -173 179 -167
rect 183 -173 186 -167
rect 190 -173 193 -167
rect 197 -173 200 -167
rect 204 -173 210 -167
rect 211 -173 217 -167
rect 218 -173 221 -167
rect 225 -173 228 -167
rect 232 -173 238 -167
rect 239 -173 245 -167
rect 246 -173 249 -167
rect 253 -173 256 -167
rect 260 -173 263 -167
rect 267 -173 270 -167
rect 274 -173 277 -167
rect 281 -173 284 -167
rect 288 -173 291 -167
rect 295 -173 298 -167
rect 302 -173 305 -167
rect 309 -173 312 -167
rect 316 -173 319 -167
rect 323 -173 326 -167
rect 330 -173 333 -167
rect 337 -173 340 -167
rect 344 -173 347 -167
rect 351 -173 357 -167
rect 358 -173 364 -167
rect 365 -173 368 -167
rect 372 -173 375 -167
rect 379 -173 382 -167
rect 386 -173 389 -167
rect 393 -173 396 -167
rect 400 -173 403 -167
rect 407 -173 410 -167
rect 414 -173 417 -167
rect 421 -173 424 -167
rect 428 -173 434 -167
rect 435 -173 438 -167
rect 442 -173 445 -167
rect 449 -173 452 -167
rect 456 -173 459 -167
rect 463 -173 469 -167
rect 470 -173 473 -167
rect 477 -173 483 -167
rect 484 -173 487 -167
rect 491 -173 494 -167
rect 498 -173 504 -167
rect 505 -173 511 -167
rect 512 -173 518 -167
rect 519 -173 525 -167
rect 526 -173 529 -167
rect 533 -173 536 -167
rect 540 -173 546 -167
rect 547 -173 550 -167
rect 554 -173 557 -167
rect 561 -173 564 -167
rect 568 -173 571 -167
rect 575 -173 578 -167
rect 582 -173 585 -167
rect 589 -173 592 -167
rect 596 -173 599 -167
rect 603 -173 606 -167
rect 610 -173 616 -167
rect 617 -173 620 -167
rect 624 -173 627 -167
rect 631 -173 634 -167
rect 638 -173 641 -167
rect 645 -173 648 -167
rect 652 -173 658 -167
rect 659 -173 662 -167
rect 666 -173 669 -167
rect 673 -173 676 -167
rect 680 -173 683 -167
rect 687 -173 690 -167
rect 694 -173 700 -167
rect 701 -173 704 -167
rect 708 -173 711 -167
rect 715 -173 718 -167
rect 722 -173 725 -167
rect 729 -173 732 -167
rect 736 -173 739 -167
rect 743 -173 746 -167
rect 750 -173 753 -167
rect 757 -173 760 -167
rect 764 -173 770 -167
rect 771 -173 774 -167
rect 778 -173 781 -167
rect 785 -173 788 -167
rect 792 -173 798 -167
rect 799 -173 802 -167
rect 806 -173 809 -167
rect 813 -173 816 -167
rect 820 -173 826 -167
rect 827 -173 830 -167
rect 834 -173 837 -167
rect 841 -173 844 -167
rect 848 -173 851 -167
rect 855 -173 858 -167
rect 862 -173 865 -167
rect 869 -173 872 -167
rect 876 -173 882 -167
rect 883 -173 889 -167
rect 890 -173 893 -167
rect 897 -173 900 -167
rect 904 -173 907 -167
rect 911 -173 914 -167
rect 918 -173 921 -167
rect 925 -173 928 -167
rect 932 -173 935 -167
rect 939 -173 942 -167
rect 946 -173 949 -167
rect 953 -173 956 -167
rect 960 -173 963 -167
rect 967 -173 970 -167
rect 974 -173 977 -167
rect 981 -173 984 -167
rect 995 -173 998 -167
rect 1009 -173 1012 -167
rect 1037 -173 1040 -167
rect 1128 -173 1131 -167
rect 1135 -173 1138 -167
rect 1191 -173 1197 -167
rect 1219 -173 1222 -167
rect 1 -260 7 -254
rect 8 -260 14 -254
rect 15 -260 21 -254
rect 22 -260 28 -254
rect 29 -260 35 -254
rect 36 -260 42 -254
rect 50 -260 53 -254
rect 57 -260 60 -254
rect 64 -260 67 -254
rect 71 -260 74 -254
rect 78 -260 81 -254
rect 85 -260 88 -254
rect 92 -260 95 -254
rect 99 -260 102 -254
rect 106 -260 109 -254
rect 113 -260 119 -254
rect 120 -260 123 -254
rect 127 -260 130 -254
rect 134 -260 137 -254
rect 141 -260 144 -254
rect 148 -260 151 -254
rect 155 -260 158 -254
rect 162 -260 165 -254
rect 169 -260 175 -254
rect 176 -260 179 -254
rect 183 -260 186 -254
rect 190 -260 196 -254
rect 197 -260 203 -254
rect 204 -260 207 -254
rect 211 -260 217 -254
rect 218 -260 221 -254
rect 225 -260 228 -254
rect 232 -260 238 -254
rect 239 -260 245 -254
rect 246 -260 249 -254
rect 253 -260 256 -254
rect 260 -260 263 -254
rect 267 -260 270 -254
rect 274 -260 277 -254
rect 281 -260 284 -254
rect 288 -260 294 -254
rect 295 -260 298 -254
rect 302 -260 305 -254
rect 309 -260 312 -254
rect 316 -260 319 -254
rect 323 -260 326 -254
rect 330 -260 333 -254
rect 337 -260 340 -254
rect 344 -260 347 -254
rect 351 -260 354 -254
rect 358 -260 361 -254
rect 365 -260 368 -254
rect 372 -260 375 -254
rect 379 -260 385 -254
rect 386 -260 389 -254
rect 393 -260 396 -254
rect 400 -260 403 -254
rect 407 -260 410 -254
rect 414 -260 417 -254
rect 421 -260 424 -254
rect 428 -260 431 -254
rect 435 -260 438 -254
rect 442 -260 448 -254
rect 449 -260 452 -254
rect 456 -260 462 -254
rect 463 -260 469 -254
rect 470 -260 476 -254
rect 477 -260 480 -254
rect 484 -260 487 -254
rect 491 -260 497 -254
rect 498 -260 501 -254
rect 505 -260 511 -254
rect 512 -260 515 -254
rect 519 -260 522 -254
rect 526 -260 532 -254
rect 533 -260 536 -254
rect 540 -260 546 -254
rect 547 -260 550 -254
rect 554 -260 557 -254
rect 561 -260 564 -254
rect 568 -260 574 -254
rect 575 -260 581 -254
rect 582 -260 585 -254
rect 589 -260 595 -254
rect 596 -260 599 -254
rect 603 -260 606 -254
rect 610 -260 616 -254
rect 617 -260 620 -254
rect 624 -260 627 -254
rect 631 -260 634 -254
rect 638 -260 641 -254
rect 645 -260 648 -254
rect 652 -260 655 -254
rect 659 -260 662 -254
rect 666 -260 669 -254
rect 673 -260 676 -254
rect 680 -260 683 -254
rect 687 -260 690 -254
rect 694 -260 697 -254
rect 701 -260 704 -254
rect 708 -260 711 -254
rect 715 -260 721 -254
rect 722 -260 725 -254
rect 729 -260 732 -254
rect 736 -260 739 -254
rect 743 -260 746 -254
rect 750 -260 753 -254
rect 757 -260 760 -254
rect 764 -260 767 -254
rect 771 -260 777 -254
rect 778 -260 781 -254
rect 785 -260 791 -254
rect 792 -260 795 -254
rect 799 -260 802 -254
rect 806 -260 809 -254
rect 813 -260 816 -254
rect 820 -260 823 -254
rect 827 -260 833 -254
rect 834 -260 837 -254
rect 841 -260 844 -254
rect 848 -260 851 -254
rect 855 -260 858 -254
rect 862 -260 865 -254
rect 869 -260 872 -254
rect 876 -260 879 -254
rect 883 -260 886 -254
rect 890 -260 893 -254
rect 897 -260 900 -254
rect 904 -260 907 -254
rect 911 -260 914 -254
rect 918 -260 921 -254
rect 925 -260 928 -254
rect 932 -260 935 -254
rect 939 -260 942 -254
rect 946 -260 949 -254
rect 953 -260 956 -254
rect 960 -260 963 -254
rect 967 -260 970 -254
rect 974 -260 977 -254
rect 981 -260 984 -254
rect 988 -260 991 -254
rect 995 -260 1001 -254
rect 1002 -260 1005 -254
rect 1009 -260 1012 -254
rect 1016 -260 1019 -254
rect 1023 -260 1026 -254
rect 1030 -260 1033 -254
rect 1037 -260 1040 -254
rect 1044 -260 1047 -254
rect 1051 -260 1054 -254
rect 1058 -260 1061 -254
rect 1065 -260 1068 -254
rect 1072 -260 1075 -254
rect 1079 -260 1082 -254
rect 1086 -260 1089 -254
rect 1093 -260 1099 -254
rect 1100 -260 1103 -254
rect 1107 -260 1110 -254
rect 1114 -260 1120 -254
rect 1121 -260 1127 -254
rect 1128 -260 1131 -254
rect 1135 -260 1138 -254
rect 1142 -260 1145 -254
rect 1149 -260 1152 -254
rect 1156 -260 1159 -254
rect 1163 -260 1166 -254
rect 1170 -260 1173 -254
rect 1226 -260 1229 -254
rect 1254 -260 1257 -254
rect 1282 -260 1285 -254
rect 1 -391 7 -385
rect 8 -391 14 -385
rect 15 -391 21 -385
rect 22 -391 28 -385
rect 29 -391 35 -385
rect 36 -391 42 -385
rect 43 -391 46 -385
rect 50 -391 53 -385
rect 57 -391 63 -385
rect 64 -391 67 -385
rect 71 -391 74 -385
rect 78 -391 81 -385
rect 85 -391 88 -385
rect 92 -391 98 -385
rect 99 -391 102 -385
rect 106 -391 109 -385
rect 113 -391 119 -385
rect 120 -391 126 -385
rect 127 -391 130 -385
rect 134 -391 140 -385
rect 141 -391 144 -385
rect 148 -391 151 -385
rect 155 -391 158 -385
rect 162 -391 165 -385
rect 169 -391 172 -385
rect 176 -391 179 -385
rect 183 -391 186 -385
rect 190 -391 193 -385
rect 197 -391 203 -385
rect 204 -391 210 -385
rect 211 -391 217 -385
rect 218 -391 221 -385
rect 225 -391 228 -385
rect 232 -391 238 -385
rect 239 -391 242 -385
rect 246 -391 252 -385
rect 253 -391 256 -385
rect 260 -391 263 -385
rect 267 -391 270 -385
rect 274 -391 277 -385
rect 281 -391 287 -385
rect 288 -391 291 -385
rect 295 -391 298 -385
rect 302 -391 305 -385
rect 309 -391 312 -385
rect 316 -391 322 -385
rect 323 -391 326 -385
rect 330 -391 333 -385
rect 337 -391 343 -385
rect 344 -391 347 -385
rect 351 -391 354 -385
rect 358 -391 361 -385
rect 365 -391 368 -385
rect 372 -391 375 -385
rect 379 -391 382 -385
rect 386 -391 389 -385
rect 393 -391 396 -385
rect 400 -391 403 -385
rect 407 -391 413 -385
rect 414 -391 417 -385
rect 421 -391 424 -385
rect 428 -391 431 -385
rect 435 -391 441 -385
rect 442 -391 445 -385
rect 449 -391 455 -385
rect 456 -391 459 -385
rect 463 -391 466 -385
rect 470 -391 476 -385
rect 477 -391 480 -385
rect 484 -391 487 -385
rect 491 -391 494 -385
rect 498 -391 501 -385
rect 505 -391 511 -385
rect 512 -391 515 -385
rect 519 -391 522 -385
rect 526 -391 529 -385
rect 533 -391 536 -385
rect 540 -391 543 -385
rect 547 -391 550 -385
rect 554 -391 557 -385
rect 561 -391 564 -385
rect 568 -391 574 -385
rect 575 -391 578 -385
rect 582 -391 585 -385
rect 589 -391 592 -385
rect 596 -391 599 -385
rect 603 -391 609 -385
rect 610 -391 616 -385
rect 617 -391 620 -385
rect 624 -391 627 -385
rect 631 -391 634 -385
rect 638 -391 641 -385
rect 645 -391 648 -385
rect 652 -391 655 -385
rect 659 -391 662 -385
rect 666 -391 672 -385
rect 673 -391 676 -385
rect 680 -391 683 -385
rect 687 -391 690 -385
rect 694 -391 697 -385
rect 701 -391 707 -385
rect 708 -391 714 -385
rect 715 -391 718 -385
rect 722 -391 725 -385
rect 729 -391 735 -385
rect 736 -391 739 -385
rect 743 -391 749 -385
rect 750 -391 756 -385
rect 757 -391 760 -385
rect 764 -391 767 -385
rect 771 -391 774 -385
rect 778 -391 781 -385
rect 785 -391 788 -385
rect 792 -391 795 -385
rect 799 -391 802 -385
rect 806 -391 809 -385
rect 813 -391 816 -385
rect 820 -391 823 -385
rect 827 -391 830 -385
rect 834 -391 837 -385
rect 841 -391 844 -385
rect 848 -391 851 -385
rect 855 -391 858 -385
rect 862 -391 865 -385
rect 869 -391 872 -385
rect 876 -391 879 -385
rect 883 -391 886 -385
rect 890 -391 893 -385
rect 897 -391 900 -385
rect 904 -391 907 -385
rect 911 -391 914 -385
rect 918 -391 921 -385
rect 925 -391 928 -385
rect 932 -391 935 -385
rect 939 -391 942 -385
rect 946 -391 949 -385
rect 953 -391 956 -385
rect 960 -391 963 -385
rect 967 -391 970 -385
rect 974 -391 977 -385
rect 981 -391 984 -385
rect 988 -391 991 -385
rect 995 -391 998 -385
rect 1002 -391 1005 -385
rect 1009 -391 1012 -385
rect 1016 -391 1019 -385
rect 1023 -391 1026 -385
rect 1030 -391 1033 -385
rect 1037 -391 1040 -385
rect 1044 -391 1047 -385
rect 1051 -391 1054 -385
rect 1058 -391 1061 -385
rect 1065 -391 1068 -385
rect 1072 -391 1075 -385
rect 1079 -391 1082 -385
rect 1086 -391 1089 -385
rect 1093 -391 1096 -385
rect 1100 -391 1103 -385
rect 1107 -391 1110 -385
rect 1114 -391 1117 -385
rect 1121 -391 1124 -385
rect 1128 -391 1131 -385
rect 1135 -391 1138 -385
rect 1142 -391 1145 -385
rect 1149 -391 1152 -385
rect 1156 -391 1159 -385
rect 1163 -391 1166 -385
rect 1170 -391 1173 -385
rect 1177 -391 1180 -385
rect 1184 -391 1187 -385
rect 1191 -391 1194 -385
rect 1198 -391 1204 -385
rect 1205 -391 1208 -385
rect 1212 -391 1215 -385
rect 1219 -391 1222 -385
rect 1226 -391 1229 -385
rect 1233 -391 1236 -385
rect 1240 -391 1243 -385
rect 1247 -391 1250 -385
rect 1254 -391 1257 -385
rect 1261 -391 1264 -385
rect 1268 -391 1271 -385
rect 1275 -391 1278 -385
rect 1282 -391 1285 -385
rect 1289 -391 1292 -385
rect 1296 -391 1299 -385
rect 1303 -391 1306 -385
rect 1310 -391 1313 -385
rect 1317 -391 1320 -385
rect 1324 -391 1327 -385
rect 1331 -391 1334 -385
rect 1338 -391 1341 -385
rect 1345 -391 1348 -385
rect 1352 -391 1355 -385
rect 1359 -391 1362 -385
rect 1366 -391 1369 -385
rect 1373 -391 1376 -385
rect 1380 -391 1383 -385
rect 1387 -391 1390 -385
rect 1394 -391 1400 -385
rect 1590 -391 1593 -385
rect 1 -502 7 -496
rect 8 -502 14 -496
rect 15 -502 21 -496
rect 22 -502 28 -496
rect 29 -502 32 -496
rect 36 -502 39 -496
rect 43 -502 46 -496
rect 50 -502 53 -496
rect 57 -502 60 -496
rect 64 -502 67 -496
rect 71 -502 74 -496
rect 78 -502 84 -496
rect 85 -502 91 -496
rect 92 -502 95 -496
rect 99 -502 105 -496
rect 106 -502 112 -496
rect 113 -502 116 -496
rect 120 -502 123 -496
rect 127 -502 130 -496
rect 134 -502 140 -496
rect 141 -502 144 -496
rect 148 -502 151 -496
rect 155 -502 158 -496
rect 162 -502 165 -496
rect 169 -502 172 -496
rect 176 -502 182 -496
rect 183 -502 189 -496
rect 190 -502 196 -496
rect 197 -502 200 -496
rect 204 -502 207 -496
rect 211 -502 214 -496
rect 218 -502 224 -496
rect 225 -502 228 -496
rect 232 -502 235 -496
rect 239 -502 242 -496
rect 246 -502 249 -496
rect 253 -502 256 -496
rect 260 -502 263 -496
rect 267 -502 270 -496
rect 274 -502 277 -496
rect 281 -502 284 -496
rect 288 -502 291 -496
rect 295 -502 301 -496
rect 302 -502 305 -496
rect 309 -502 312 -496
rect 316 -502 319 -496
rect 323 -502 326 -496
rect 330 -502 333 -496
rect 337 -502 340 -496
rect 344 -502 347 -496
rect 351 -502 354 -496
rect 358 -502 364 -496
rect 365 -502 368 -496
rect 372 -502 375 -496
rect 379 -502 382 -496
rect 386 -502 389 -496
rect 393 -502 396 -496
rect 400 -502 403 -496
rect 407 -502 410 -496
rect 414 -502 420 -496
rect 421 -502 424 -496
rect 428 -502 431 -496
rect 435 -502 438 -496
rect 442 -502 445 -496
rect 449 -502 455 -496
rect 456 -502 459 -496
rect 463 -502 466 -496
rect 470 -502 476 -496
rect 477 -502 483 -496
rect 484 -502 487 -496
rect 491 -502 497 -496
rect 498 -502 501 -496
rect 505 -502 508 -496
rect 512 -502 518 -496
rect 519 -502 525 -496
rect 526 -502 532 -496
rect 533 -502 539 -496
rect 540 -502 543 -496
rect 547 -502 550 -496
rect 554 -502 557 -496
rect 561 -502 564 -496
rect 568 -502 571 -496
rect 575 -502 578 -496
rect 582 -502 585 -496
rect 589 -502 595 -496
rect 596 -502 602 -496
rect 603 -502 606 -496
rect 610 -502 613 -496
rect 617 -502 620 -496
rect 624 -502 627 -496
rect 631 -502 637 -496
rect 638 -502 641 -496
rect 645 -502 651 -496
rect 652 -502 655 -496
rect 659 -502 662 -496
rect 666 -502 669 -496
rect 673 -502 676 -496
rect 680 -502 683 -496
rect 687 -502 690 -496
rect 694 -502 700 -496
rect 701 -502 704 -496
rect 708 -502 714 -496
rect 715 -502 718 -496
rect 722 -502 725 -496
rect 729 -502 732 -496
rect 736 -502 739 -496
rect 743 -502 746 -496
rect 750 -502 753 -496
rect 757 -502 763 -496
rect 764 -502 767 -496
rect 771 -502 774 -496
rect 778 -502 781 -496
rect 785 -502 788 -496
rect 792 -502 795 -496
rect 799 -502 802 -496
rect 806 -502 809 -496
rect 813 -502 816 -496
rect 820 -502 823 -496
rect 827 -502 833 -496
rect 834 -502 837 -496
rect 841 -502 844 -496
rect 848 -502 851 -496
rect 855 -502 858 -496
rect 862 -502 865 -496
rect 869 -502 872 -496
rect 876 -502 879 -496
rect 883 -502 886 -496
rect 890 -502 893 -496
rect 897 -502 903 -496
rect 904 -502 907 -496
rect 911 -502 914 -496
rect 918 -502 921 -496
rect 925 -502 928 -496
rect 932 -502 935 -496
rect 939 -502 942 -496
rect 946 -502 949 -496
rect 953 -502 956 -496
rect 960 -502 963 -496
rect 967 -502 970 -496
rect 974 -502 977 -496
rect 981 -502 984 -496
rect 988 -502 991 -496
rect 995 -502 998 -496
rect 1002 -502 1005 -496
rect 1009 -502 1012 -496
rect 1016 -502 1019 -496
rect 1023 -502 1026 -496
rect 1030 -502 1033 -496
rect 1037 -502 1040 -496
rect 1044 -502 1047 -496
rect 1051 -502 1054 -496
rect 1058 -502 1061 -496
rect 1065 -502 1068 -496
rect 1072 -502 1075 -496
rect 1079 -502 1082 -496
rect 1086 -502 1089 -496
rect 1093 -502 1096 -496
rect 1100 -502 1103 -496
rect 1107 -502 1110 -496
rect 1114 -502 1117 -496
rect 1121 -502 1124 -496
rect 1128 -502 1131 -496
rect 1135 -502 1138 -496
rect 1142 -502 1145 -496
rect 1149 -502 1152 -496
rect 1156 -502 1159 -496
rect 1163 -502 1166 -496
rect 1170 -502 1173 -496
rect 1177 -502 1180 -496
rect 1184 -502 1187 -496
rect 1191 -502 1197 -496
rect 1198 -502 1201 -496
rect 1205 -502 1208 -496
rect 1212 -502 1215 -496
rect 1219 -502 1222 -496
rect 1226 -502 1229 -496
rect 1233 -502 1236 -496
rect 1240 -502 1243 -496
rect 1247 -502 1250 -496
rect 1254 -502 1257 -496
rect 1261 -502 1264 -496
rect 1268 -502 1271 -496
rect 1275 -502 1278 -496
rect 1282 -502 1285 -496
rect 1289 -502 1292 -496
rect 1296 -502 1299 -496
rect 1303 -502 1306 -496
rect 1310 -502 1313 -496
rect 1317 -502 1320 -496
rect 1324 -502 1327 -496
rect 1331 -502 1334 -496
rect 1338 -502 1341 -496
rect 1345 -502 1348 -496
rect 1352 -502 1355 -496
rect 1359 -502 1362 -496
rect 1366 -502 1369 -496
rect 1373 -502 1376 -496
rect 1380 -502 1383 -496
rect 1387 -502 1390 -496
rect 1394 -502 1397 -496
rect 1401 -502 1404 -496
rect 1408 -502 1411 -496
rect 1415 -502 1418 -496
rect 1422 -502 1425 -496
rect 1429 -502 1432 -496
rect 1436 -502 1439 -496
rect 1443 -502 1446 -496
rect 1450 -502 1453 -496
rect 1457 -502 1460 -496
rect 1464 -502 1467 -496
rect 1471 -502 1474 -496
rect 1478 -502 1481 -496
rect 1485 -502 1488 -496
rect 1492 -502 1495 -496
rect 1499 -502 1502 -496
rect 1506 -502 1509 -496
rect 1513 -502 1516 -496
rect 1520 -502 1526 -496
rect 1527 -502 1530 -496
rect 1709 -502 1712 -496
rect 1 -609 7 -603
rect 8 -609 11 -603
rect 15 -609 21 -603
rect 22 -609 25 -603
rect 29 -609 35 -603
rect 36 -609 42 -603
rect 43 -609 46 -603
rect 50 -609 53 -603
rect 57 -609 63 -603
rect 64 -609 67 -603
rect 71 -609 74 -603
rect 78 -609 81 -603
rect 85 -609 88 -603
rect 92 -609 95 -603
rect 99 -609 105 -603
rect 106 -609 109 -603
rect 113 -609 116 -603
rect 120 -609 123 -603
rect 127 -609 130 -603
rect 134 -609 137 -603
rect 141 -609 144 -603
rect 148 -609 154 -603
rect 155 -609 158 -603
rect 162 -609 165 -603
rect 169 -609 172 -603
rect 176 -609 179 -603
rect 183 -609 189 -603
rect 190 -609 193 -603
rect 197 -609 200 -603
rect 204 -609 207 -603
rect 211 -609 214 -603
rect 218 -609 221 -603
rect 225 -609 228 -603
rect 232 -609 238 -603
rect 239 -609 245 -603
rect 246 -609 249 -603
rect 253 -609 256 -603
rect 260 -609 263 -603
rect 267 -609 270 -603
rect 274 -609 277 -603
rect 281 -609 284 -603
rect 288 -609 291 -603
rect 295 -609 298 -603
rect 302 -609 305 -603
rect 309 -609 312 -603
rect 316 -609 322 -603
rect 323 -609 326 -603
rect 330 -609 333 -603
rect 337 -609 343 -603
rect 344 -609 347 -603
rect 351 -609 354 -603
rect 358 -609 361 -603
rect 365 -609 368 -603
rect 372 -609 375 -603
rect 379 -609 385 -603
rect 386 -609 389 -603
rect 393 -609 396 -603
rect 400 -609 403 -603
rect 407 -609 410 -603
rect 414 -609 417 -603
rect 421 -609 424 -603
rect 428 -609 434 -603
rect 435 -609 438 -603
rect 442 -609 445 -603
rect 449 -609 455 -603
rect 456 -609 462 -603
rect 463 -609 466 -603
rect 470 -609 473 -603
rect 477 -609 480 -603
rect 484 -609 487 -603
rect 491 -609 494 -603
rect 498 -609 501 -603
rect 505 -609 508 -603
rect 512 -609 518 -603
rect 519 -609 522 -603
rect 526 -609 532 -603
rect 533 -609 536 -603
rect 540 -609 543 -603
rect 547 -609 550 -603
rect 554 -609 557 -603
rect 561 -609 564 -603
rect 568 -609 571 -603
rect 575 -609 581 -603
rect 582 -609 588 -603
rect 589 -609 595 -603
rect 596 -609 599 -603
rect 603 -609 606 -603
rect 610 -609 613 -603
rect 617 -609 620 -603
rect 624 -609 627 -603
rect 631 -609 637 -603
rect 638 -609 641 -603
rect 645 -609 648 -603
rect 652 -609 655 -603
rect 659 -609 662 -603
rect 666 -609 669 -603
rect 673 -609 679 -603
rect 680 -609 683 -603
rect 687 -609 690 -603
rect 694 -609 700 -603
rect 701 -609 704 -603
rect 708 -609 711 -603
rect 715 -609 718 -603
rect 722 -609 725 -603
rect 729 -609 732 -603
rect 736 -609 739 -603
rect 743 -609 746 -603
rect 750 -609 753 -603
rect 757 -609 760 -603
rect 764 -609 767 -603
rect 771 -609 774 -603
rect 778 -609 784 -603
rect 785 -609 788 -603
rect 792 -609 795 -603
rect 799 -609 802 -603
rect 806 -609 809 -603
rect 813 -609 816 -603
rect 820 -609 826 -603
rect 827 -609 830 -603
rect 834 -609 837 -603
rect 841 -609 847 -603
rect 848 -609 854 -603
rect 855 -609 858 -603
rect 862 -609 868 -603
rect 869 -609 875 -603
rect 876 -609 879 -603
rect 883 -609 886 -603
rect 890 -609 896 -603
rect 897 -609 900 -603
rect 904 -609 907 -603
rect 911 -609 917 -603
rect 918 -609 921 -603
rect 925 -609 928 -603
rect 932 -609 938 -603
rect 939 -609 942 -603
rect 946 -609 949 -603
rect 953 -609 956 -603
rect 960 -609 963 -603
rect 967 -609 970 -603
rect 974 -609 977 -603
rect 981 -609 984 -603
rect 988 -609 991 -603
rect 995 -609 998 -603
rect 1002 -609 1005 -603
rect 1009 -609 1012 -603
rect 1016 -609 1019 -603
rect 1023 -609 1026 -603
rect 1030 -609 1033 -603
rect 1037 -609 1040 -603
rect 1044 -609 1047 -603
rect 1051 -609 1057 -603
rect 1058 -609 1061 -603
rect 1065 -609 1068 -603
rect 1072 -609 1075 -603
rect 1079 -609 1082 -603
rect 1086 -609 1089 -603
rect 1093 -609 1096 -603
rect 1100 -609 1103 -603
rect 1107 -609 1110 -603
rect 1114 -609 1117 -603
rect 1121 -609 1124 -603
rect 1128 -609 1131 -603
rect 1135 -609 1138 -603
rect 1142 -609 1145 -603
rect 1149 -609 1152 -603
rect 1156 -609 1159 -603
rect 1163 -609 1166 -603
rect 1170 -609 1173 -603
rect 1177 -609 1180 -603
rect 1184 -609 1187 -603
rect 1191 -609 1194 -603
rect 1198 -609 1201 -603
rect 1205 -609 1208 -603
rect 1212 -609 1215 -603
rect 1219 -609 1222 -603
rect 1226 -609 1229 -603
rect 1233 -609 1236 -603
rect 1240 -609 1243 -603
rect 1247 -609 1250 -603
rect 1254 -609 1257 -603
rect 1261 -609 1264 -603
rect 1268 -609 1271 -603
rect 1275 -609 1278 -603
rect 1282 -609 1285 -603
rect 1289 -609 1292 -603
rect 1296 -609 1299 -603
rect 1303 -609 1306 -603
rect 1310 -609 1313 -603
rect 1317 -609 1320 -603
rect 1324 -609 1327 -603
rect 1331 -609 1334 -603
rect 1338 -609 1341 -603
rect 1345 -609 1348 -603
rect 1352 -609 1355 -603
rect 1359 -609 1362 -603
rect 1366 -609 1369 -603
rect 1373 -609 1376 -603
rect 1380 -609 1383 -603
rect 1387 -609 1390 -603
rect 1394 -609 1397 -603
rect 1401 -609 1404 -603
rect 1408 -609 1411 -603
rect 1415 -609 1418 -603
rect 1422 -609 1425 -603
rect 1429 -609 1432 -603
rect 1436 -609 1439 -603
rect 1443 -609 1446 -603
rect 1450 -609 1453 -603
rect 1457 -609 1460 -603
rect 1464 -609 1470 -603
rect 1471 -609 1474 -603
rect 1478 -609 1481 -603
rect 1485 -609 1488 -603
rect 1492 -609 1495 -603
rect 1499 -609 1502 -603
rect 1506 -609 1509 -603
rect 1513 -609 1516 -603
rect 1520 -609 1523 -603
rect 1534 -609 1537 -603
rect 1555 -609 1558 -603
rect 1737 -609 1740 -603
rect 1758 -609 1761 -603
rect 1765 -609 1768 -603
rect 1 -718 7 -712
rect 8 -718 11 -712
rect 15 -718 18 -712
rect 22 -718 25 -712
rect 29 -718 32 -712
rect 36 -718 39 -712
rect 43 -718 46 -712
rect 50 -718 53 -712
rect 57 -718 60 -712
rect 64 -718 67 -712
rect 71 -718 74 -712
rect 78 -718 81 -712
rect 85 -718 88 -712
rect 92 -718 98 -712
rect 99 -718 102 -712
rect 106 -718 109 -712
rect 113 -718 119 -712
rect 120 -718 123 -712
rect 127 -718 130 -712
rect 134 -718 140 -712
rect 141 -718 147 -712
rect 148 -718 151 -712
rect 155 -718 158 -712
rect 162 -718 165 -712
rect 169 -718 175 -712
rect 176 -718 179 -712
rect 183 -718 189 -712
rect 190 -718 193 -712
rect 197 -718 200 -712
rect 204 -718 207 -712
rect 211 -718 214 -712
rect 218 -718 221 -712
rect 225 -718 228 -712
rect 232 -718 238 -712
rect 239 -718 242 -712
rect 246 -718 249 -712
rect 253 -718 256 -712
rect 260 -718 263 -712
rect 267 -718 270 -712
rect 274 -718 277 -712
rect 281 -718 284 -712
rect 288 -718 291 -712
rect 295 -718 298 -712
rect 302 -718 305 -712
rect 309 -718 312 -712
rect 316 -718 319 -712
rect 323 -718 326 -712
rect 330 -718 333 -712
rect 337 -718 340 -712
rect 344 -718 347 -712
rect 351 -718 354 -712
rect 358 -718 364 -712
rect 365 -718 368 -712
rect 372 -718 375 -712
rect 379 -718 382 -712
rect 386 -718 389 -712
rect 393 -718 396 -712
rect 400 -718 403 -712
rect 407 -718 410 -712
rect 414 -718 417 -712
rect 421 -718 424 -712
rect 428 -718 431 -712
rect 435 -718 438 -712
rect 442 -718 445 -712
rect 449 -718 452 -712
rect 456 -718 459 -712
rect 463 -718 469 -712
rect 470 -718 473 -712
rect 477 -718 483 -712
rect 484 -718 487 -712
rect 491 -718 494 -712
rect 498 -718 501 -712
rect 505 -718 511 -712
rect 512 -718 515 -712
rect 519 -718 522 -712
rect 526 -718 529 -712
rect 533 -718 536 -712
rect 540 -718 546 -712
rect 547 -718 550 -712
rect 554 -718 560 -712
rect 561 -718 564 -712
rect 568 -718 571 -712
rect 575 -718 578 -712
rect 582 -718 585 -712
rect 589 -718 592 -712
rect 596 -718 602 -712
rect 603 -718 606 -712
rect 610 -718 613 -712
rect 617 -718 623 -712
rect 624 -718 627 -712
rect 631 -718 634 -712
rect 638 -718 641 -712
rect 645 -718 651 -712
rect 652 -718 655 -712
rect 659 -718 662 -712
rect 666 -718 669 -712
rect 673 -718 676 -712
rect 680 -718 683 -712
rect 687 -718 693 -712
rect 694 -718 697 -712
rect 701 -718 704 -712
rect 708 -718 714 -712
rect 715 -718 721 -712
rect 722 -718 725 -712
rect 729 -718 732 -712
rect 736 -718 742 -712
rect 743 -718 746 -712
rect 750 -718 753 -712
rect 757 -718 763 -712
rect 764 -718 767 -712
rect 771 -718 774 -712
rect 778 -718 784 -712
rect 785 -718 788 -712
rect 792 -718 798 -712
rect 799 -718 802 -712
rect 806 -718 809 -712
rect 813 -718 816 -712
rect 820 -718 823 -712
rect 827 -718 833 -712
rect 834 -718 837 -712
rect 841 -718 847 -712
rect 848 -718 851 -712
rect 855 -718 858 -712
rect 862 -718 865 -712
rect 869 -718 872 -712
rect 876 -718 879 -712
rect 883 -718 886 -712
rect 890 -718 893 -712
rect 897 -718 903 -712
rect 904 -718 910 -712
rect 911 -718 914 -712
rect 918 -718 924 -712
rect 925 -718 928 -712
rect 932 -718 935 -712
rect 939 -718 942 -712
rect 946 -718 949 -712
rect 953 -718 956 -712
rect 960 -718 963 -712
rect 967 -718 973 -712
rect 974 -718 977 -712
rect 981 -718 984 -712
rect 988 -718 991 -712
rect 995 -718 1001 -712
rect 1002 -718 1005 -712
rect 1009 -718 1012 -712
rect 1016 -718 1022 -712
rect 1023 -718 1026 -712
rect 1030 -718 1033 -712
rect 1037 -718 1040 -712
rect 1044 -718 1047 -712
rect 1051 -718 1054 -712
rect 1058 -718 1061 -712
rect 1065 -718 1068 -712
rect 1072 -718 1075 -712
rect 1079 -718 1082 -712
rect 1086 -718 1089 -712
rect 1093 -718 1096 -712
rect 1100 -718 1103 -712
rect 1107 -718 1110 -712
rect 1114 -718 1117 -712
rect 1121 -718 1127 -712
rect 1128 -718 1131 -712
rect 1135 -718 1138 -712
rect 1142 -718 1145 -712
rect 1149 -718 1152 -712
rect 1156 -718 1159 -712
rect 1163 -718 1166 -712
rect 1170 -718 1173 -712
rect 1177 -718 1180 -712
rect 1184 -718 1187 -712
rect 1191 -718 1194 -712
rect 1198 -718 1201 -712
rect 1205 -718 1208 -712
rect 1212 -718 1215 -712
rect 1219 -718 1222 -712
rect 1226 -718 1229 -712
rect 1233 -718 1236 -712
rect 1240 -718 1243 -712
rect 1247 -718 1250 -712
rect 1254 -718 1257 -712
rect 1261 -718 1264 -712
rect 1268 -718 1271 -712
rect 1275 -718 1278 -712
rect 1282 -718 1285 -712
rect 1289 -718 1292 -712
rect 1296 -718 1299 -712
rect 1303 -718 1306 -712
rect 1310 -718 1313 -712
rect 1317 -718 1320 -712
rect 1324 -718 1327 -712
rect 1331 -718 1334 -712
rect 1338 -718 1341 -712
rect 1345 -718 1348 -712
rect 1352 -718 1355 -712
rect 1359 -718 1362 -712
rect 1366 -718 1369 -712
rect 1373 -718 1376 -712
rect 1380 -718 1383 -712
rect 1387 -718 1390 -712
rect 1394 -718 1397 -712
rect 1401 -718 1404 -712
rect 1408 -718 1411 -712
rect 1415 -718 1418 -712
rect 1422 -718 1425 -712
rect 1429 -718 1432 -712
rect 1436 -718 1439 -712
rect 1443 -718 1446 -712
rect 1450 -718 1453 -712
rect 1457 -718 1460 -712
rect 1464 -718 1467 -712
rect 1471 -718 1474 -712
rect 1478 -718 1481 -712
rect 1485 -718 1488 -712
rect 1492 -718 1495 -712
rect 1499 -718 1502 -712
rect 1506 -718 1509 -712
rect 1513 -718 1516 -712
rect 1520 -718 1523 -712
rect 1527 -718 1530 -712
rect 1534 -718 1537 -712
rect 1541 -718 1544 -712
rect 1548 -718 1551 -712
rect 1555 -718 1558 -712
rect 1562 -718 1565 -712
rect 1569 -718 1572 -712
rect 1576 -718 1579 -712
rect 1583 -718 1586 -712
rect 1590 -718 1593 -712
rect 1597 -718 1600 -712
rect 1604 -718 1607 -712
rect 1611 -718 1614 -712
rect 1618 -718 1621 -712
rect 1625 -718 1628 -712
rect 1632 -718 1635 -712
rect 1639 -718 1642 -712
rect 1646 -718 1649 -712
rect 1653 -718 1659 -712
rect 1660 -718 1663 -712
rect 1667 -718 1673 -712
rect 1786 -718 1789 -712
rect 1793 -718 1796 -712
rect 1800 -718 1803 -712
rect 1821 -718 1824 -712
rect 1856 -718 1859 -712
rect 1 -863 7 -857
rect 8 -863 11 -857
rect 15 -863 21 -857
rect 22 -863 25 -857
rect 29 -863 32 -857
rect 36 -863 39 -857
rect 43 -863 49 -857
rect 50 -863 56 -857
rect 57 -863 60 -857
rect 64 -863 67 -857
rect 71 -863 74 -857
rect 78 -863 84 -857
rect 85 -863 88 -857
rect 92 -863 95 -857
rect 99 -863 102 -857
rect 106 -863 109 -857
rect 113 -863 116 -857
rect 120 -863 126 -857
rect 127 -863 130 -857
rect 134 -863 137 -857
rect 141 -863 144 -857
rect 148 -863 151 -857
rect 155 -863 158 -857
rect 162 -863 168 -857
rect 169 -863 172 -857
rect 176 -863 182 -857
rect 183 -863 186 -857
rect 190 -863 196 -857
rect 197 -863 203 -857
rect 204 -863 207 -857
rect 211 -863 214 -857
rect 218 -863 221 -857
rect 225 -863 228 -857
rect 232 -863 235 -857
rect 239 -863 242 -857
rect 246 -863 249 -857
rect 253 -863 256 -857
rect 260 -863 263 -857
rect 267 -863 270 -857
rect 274 -863 277 -857
rect 281 -863 284 -857
rect 288 -863 291 -857
rect 295 -863 298 -857
rect 302 -863 305 -857
rect 309 -863 312 -857
rect 316 -863 319 -857
rect 323 -863 326 -857
rect 330 -863 333 -857
rect 337 -863 340 -857
rect 344 -863 347 -857
rect 351 -863 354 -857
rect 358 -863 361 -857
rect 365 -863 368 -857
rect 372 -863 375 -857
rect 379 -863 382 -857
rect 386 -863 389 -857
rect 393 -863 396 -857
rect 400 -863 403 -857
rect 407 -863 410 -857
rect 414 -863 417 -857
rect 421 -863 424 -857
rect 428 -863 431 -857
rect 435 -863 441 -857
rect 442 -863 445 -857
rect 449 -863 452 -857
rect 456 -863 459 -857
rect 463 -863 466 -857
rect 470 -863 473 -857
rect 477 -863 480 -857
rect 484 -863 487 -857
rect 491 -863 497 -857
rect 498 -863 501 -857
rect 505 -863 508 -857
rect 512 -863 518 -857
rect 519 -863 522 -857
rect 526 -863 529 -857
rect 533 -863 536 -857
rect 540 -863 543 -857
rect 547 -863 553 -857
rect 554 -863 560 -857
rect 561 -863 564 -857
rect 568 -863 574 -857
rect 575 -863 581 -857
rect 582 -863 588 -857
rect 589 -863 592 -857
rect 596 -863 602 -857
rect 603 -863 606 -857
rect 610 -863 616 -857
rect 617 -863 623 -857
rect 624 -863 630 -857
rect 631 -863 634 -857
rect 638 -863 641 -857
rect 645 -863 648 -857
rect 652 -863 655 -857
rect 659 -863 662 -857
rect 666 -863 669 -857
rect 673 -863 676 -857
rect 680 -863 683 -857
rect 687 -863 693 -857
rect 694 -863 697 -857
rect 701 -863 707 -857
rect 708 -863 711 -857
rect 715 -863 718 -857
rect 722 -863 725 -857
rect 729 -863 732 -857
rect 736 -863 739 -857
rect 743 -863 746 -857
rect 750 -863 753 -857
rect 757 -863 763 -857
rect 764 -863 767 -857
rect 771 -863 774 -857
rect 778 -863 784 -857
rect 785 -863 791 -857
rect 792 -863 795 -857
rect 799 -863 802 -857
rect 806 -863 809 -857
rect 813 -863 816 -857
rect 820 -863 826 -857
rect 827 -863 833 -857
rect 834 -863 837 -857
rect 841 -863 844 -857
rect 848 -863 851 -857
rect 855 -863 858 -857
rect 862 -863 865 -857
rect 869 -863 872 -857
rect 876 -863 879 -857
rect 883 -863 886 -857
rect 890 -863 893 -857
rect 897 -863 900 -857
rect 904 -863 907 -857
rect 911 -863 914 -857
rect 918 -863 924 -857
rect 925 -863 928 -857
rect 932 -863 935 -857
rect 939 -863 942 -857
rect 946 -863 949 -857
rect 953 -863 956 -857
rect 960 -863 963 -857
rect 967 -863 970 -857
rect 974 -863 980 -857
rect 981 -863 984 -857
rect 988 -863 991 -857
rect 995 -863 998 -857
rect 1002 -863 1005 -857
rect 1009 -863 1012 -857
rect 1016 -863 1019 -857
rect 1023 -863 1026 -857
rect 1030 -863 1036 -857
rect 1037 -863 1040 -857
rect 1044 -863 1047 -857
rect 1051 -863 1054 -857
rect 1058 -863 1061 -857
rect 1065 -863 1068 -857
rect 1072 -863 1075 -857
rect 1079 -863 1082 -857
rect 1086 -863 1089 -857
rect 1093 -863 1096 -857
rect 1100 -863 1103 -857
rect 1107 -863 1110 -857
rect 1114 -863 1117 -857
rect 1121 -863 1124 -857
rect 1128 -863 1131 -857
rect 1135 -863 1138 -857
rect 1142 -863 1145 -857
rect 1149 -863 1152 -857
rect 1156 -863 1159 -857
rect 1163 -863 1166 -857
rect 1170 -863 1173 -857
rect 1177 -863 1180 -857
rect 1184 -863 1187 -857
rect 1191 -863 1197 -857
rect 1198 -863 1201 -857
rect 1205 -863 1208 -857
rect 1212 -863 1215 -857
rect 1219 -863 1222 -857
rect 1226 -863 1229 -857
rect 1233 -863 1236 -857
rect 1240 -863 1243 -857
rect 1247 -863 1250 -857
rect 1254 -863 1257 -857
rect 1261 -863 1264 -857
rect 1268 -863 1271 -857
rect 1275 -863 1278 -857
rect 1282 -863 1285 -857
rect 1289 -863 1292 -857
rect 1296 -863 1299 -857
rect 1303 -863 1306 -857
rect 1310 -863 1313 -857
rect 1317 -863 1320 -857
rect 1324 -863 1327 -857
rect 1331 -863 1334 -857
rect 1338 -863 1341 -857
rect 1345 -863 1348 -857
rect 1352 -863 1355 -857
rect 1359 -863 1362 -857
rect 1366 -863 1369 -857
rect 1373 -863 1376 -857
rect 1380 -863 1383 -857
rect 1387 -863 1390 -857
rect 1394 -863 1397 -857
rect 1401 -863 1404 -857
rect 1408 -863 1411 -857
rect 1415 -863 1418 -857
rect 1422 -863 1425 -857
rect 1429 -863 1432 -857
rect 1436 -863 1439 -857
rect 1443 -863 1446 -857
rect 1450 -863 1453 -857
rect 1457 -863 1460 -857
rect 1464 -863 1467 -857
rect 1471 -863 1474 -857
rect 1478 -863 1481 -857
rect 1485 -863 1488 -857
rect 1492 -863 1495 -857
rect 1499 -863 1502 -857
rect 1506 -863 1509 -857
rect 1513 -863 1516 -857
rect 1520 -863 1523 -857
rect 1527 -863 1530 -857
rect 1534 -863 1537 -857
rect 1541 -863 1544 -857
rect 1548 -863 1551 -857
rect 1555 -863 1558 -857
rect 1562 -863 1565 -857
rect 1569 -863 1572 -857
rect 1576 -863 1579 -857
rect 1583 -863 1586 -857
rect 1590 -863 1593 -857
rect 1597 -863 1600 -857
rect 1604 -863 1607 -857
rect 1611 -863 1614 -857
rect 1618 -863 1621 -857
rect 1625 -863 1628 -857
rect 1632 -863 1635 -857
rect 1639 -863 1642 -857
rect 1646 -863 1649 -857
rect 1653 -863 1656 -857
rect 1660 -863 1663 -857
rect 1667 -863 1670 -857
rect 1674 -863 1677 -857
rect 1681 -863 1684 -857
rect 1688 -863 1691 -857
rect 1695 -863 1698 -857
rect 1702 -863 1705 -857
rect 1709 -863 1712 -857
rect 1716 -863 1719 -857
rect 1723 -863 1726 -857
rect 1730 -863 1733 -857
rect 1737 -863 1740 -857
rect 1744 -863 1747 -857
rect 1751 -863 1754 -857
rect 1758 -863 1761 -857
rect 1765 -863 1768 -857
rect 1772 -863 1775 -857
rect 1779 -863 1785 -857
rect 1786 -863 1789 -857
rect 1793 -863 1796 -857
rect 1800 -863 1803 -857
rect 1807 -863 1810 -857
rect 1814 -863 1820 -857
rect 1821 -863 1824 -857
rect 1828 -863 1831 -857
rect 1835 -863 1838 -857
rect 1842 -863 1845 -857
rect 1849 -863 1852 -857
rect 1856 -863 1859 -857
rect 1884 -863 1887 -857
rect 1891 -863 1894 -857
rect 1 -984 4 -978
rect 8 -984 11 -978
rect 15 -984 18 -978
rect 22 -984 25 -978
rect 29 -984 32 -978
rect 36 -984 39 -978
rect 43 -984 46 -978
rect 50 -984 53 -978
rect 57 -984 60 -978
rect 64 -984 70 -978
rect 71 -984 74 -978
rect 78 -984 81 -978
rect 85 -984 88 -978
rect 92 -984 98 -978
rect 99 -984 102 -978
rect 106 -984 112 -978
rect 113 -984 116 -978
rect 120 -984 123 -978
rect 127 -984 130 -978
rect 134 -984 137 -978
rect 141 -984 147 -978
rect 148 -984 151 -978
rect 155 -984 161 -978
rect 162 -984 165 -978
rect 169 -984 172 -978
rect 176 -984 179 -978
rect 183 -984 189 -978
rect 190 -984 193 -978
rect 197 -984 200 -978
rect 204 -984 207 -978
rect 211 -984 214 -978
rect 218 -984 221 -978
rect 225 -984 228 -978
rect 232 -984 238 -978
rect 239 -984 242 -978
rect 246 -984 249 -978
rect 253 -984 256 -978
rect 260 -984 263 -978
rect 267 -984 270 -978
rect 274 -984 277 -978
rect 281 -984 284 -978
rect 288 -984 291 -978
rect 295 -984 298 -978
rect 302 -984 305 -978
rect 309 -984 312 -978
rect 316 -984 319 -978
rect 323 -984 326 -978
rect 330 -984 333 -978
rect 337 -984 340 -978
rect 344 -984 347 -978
rect 351 -984 354 -978
rect 358 -984 361 -978
rect 365 -984 368 -978
rect 372 -984 375 -978
rect 379 -984 382 -978
rect 386 -984 392 -978
rect 393 -984 396 -978
rect 400 -984 403 -978
rect 407 -984 410 -978
rect 414 -984 417 -978
rect 421 -984 424 -978
rect 428 -984 431 -978
rect 435 -984 438 -978
rect 442 -984 445 -978
rect 449 -984 452 -978
rect 456 -984 462 -978
rect 463 -984 466 -978
rect 470 -984 473 -978
rect 477 -984 480 -978
rect 484 -984 487 -978
rect 491 -984 494 -978
rect 498 -984 501 -978
rect 505 -984 508 -978
rect 512 -984 515 -978
rect 519 -984 522 -978
rect 526 -984 529 -978
rect 533 -984 539 -978
rect 540 -984 546 -978
rect 547 -984 550 -978
rect 554 -984 557 -978
rect 561 -984 564 -978
rect 568 -984 571 -978
rect 575 -984 578 -978
rect 582 -984 585 -978
rect 589 -984 592 -978
rect 596 -984 599 -978
rect 603 -984 609 -978
rect 610 -984 613 -978
rect 617 -984 620 -978
rect 624 -984 627 -978
rect 631 -984 634 -978
rect 638 -984 641 -978
rect 645 -984 648 -978
rect 652 -984 655 -978
rect 659 -984 662 -978
rect 666 -984 669 -978
rect 673 -984 676 -978
rect 680 -984 686 -978
rect 687 -984 690 -978
rect 694 -984 697 -978
rect 701 -984 704 -978
rect 708 -984 711 -978
rect 715 -984 718 -978
rect 722 -984 728 -978
rect 729 -984 732 -978
rect 736 -984 742 -978
rect 743 -984 749 -978
rect 750 -984 756 -978
rect 757 -984 760 -978
rect 764 -984 767 -978
rect 771 -984 777 -978
rect 778 -984 781 -978
rect 785 -984 788 -978
rect 792 -984 795 -978
rect 799 -984 802 -978
rect 806 -984 809 -978
rect 813 -984 816 -978
rect 820 -984 823 -978
rect 827 -984 830 -978
rect 834 -984 837 -978
rect 841 -984 844 -978
rect 848 -984 851 -978
rect 855 -984 858 -978
rect 862 -984 865 -978
rect 869 -984 872 -978
rect 876 -984 879 -978
rect 883 -984 886 -978
rect 890 -984 893 -978
rect 897 -984 900 -978
rect 904 -984 907 -978
rect 911 -984 917 -978
rect 918 -984 924 -978
rect 925 -984 928 -978
rect 932 -984 935 -978
rect 939 -984 945 -978
rect 946 -984 949 -978
rect 953 -984 956 -978
rect 960 -984 963 -978
rect 967 -984 970 -978
rect 974 -984 977 -978
rect 981 -984 987 -978
rect 988 -984 991 -978
rect 995 -984 998 -978
rect 1002 -984 1008 -978
rect 1009 -984 1015 -978
rect 1016 -984 1019 -978
rect 1023 -984 1026 -978
rect 1030 -984 1036 -978
rect 1037 -984 1043 -978
rect 1044 -984 1047 -978
rect 1051 -984 1054 -978
rect 1058 -984 1064 -978
rect 1065 -984 1068 -978
rect 1072 -984 1075 -978
rect 1079 -984 1085 -978
rect 1086 -984 1089 -978
rect 1093 -984 1096 -978
rect 1100 -984 1103 -978
rect 1107 -984 1110 -978
rect 1114 -984 1117 -978
rect 1121 -984 1124 -978
rect 1128 -984 1131 -978
rect 1135 -984 1138 -978
rect 1142 -984 1145 -978
rect 1149 -984 1155 -978
rect 1156 -984 1162 -978
rect 1163 -984 1166 -978
rect 1170 -984 1173 -978
rect 1177 -984 1180 -978
rect 1184 -984 1187 -978
rect 1191 -984 1194 -978
rect 1198 -984 1201 -978
rect 1205 -984 1208 -978
rect 1212 -984 1215 -978
rect 1219 -984 1222 -978
rect 1226 -984 1232 -978
rect 1233 -984 1236 -978
rect 1240 -984 1243 -978
rect 1247 -984 1250 -978
rect 1254 -984 1257 -978
rect 1261 -984 1264 -978
rect 1268 -984 1271 -978
rect 1275 -984 1278 -978
rect 1282 -984 1285 -978
rect 1289 -984 1292 -978
rect 1296 -984 1299 -978
rect 1303 -984 1306 -978
rect 1310 -984 1313 -978
rect 1317 -984 1320 -978
rect 1324 -984 1327 -978
rect 1331 -984 1334 -978
rect 1338 -984 1341 -978
rect 1345 -984 1348 -978
rect 1352 -984 1355 -978
rect 1359 -984 1362 -978
rect 1366 -984 1369 -978
rect 1373 -984 1376 -978
rect 1380 -984 1383 -978
rect 1387 -984 1390 -978
rect 1394 -984 1397 -978
rect 1401 -984 1404 -978
rect 1408 -984 1411 -978
rect 1415 -984 1418 -978
rect 1422 -984 1425 -978
rect 1429 -984 1432 -978
rect 1436 -984 1439 -978
rect 1443 -984 1446 -978
rect 1450 -984 1453 -978
rect 1457 -984 1460 -978
rect 1464 -984 1467 -978
rect 1471 -984 1474 -978
rect 1478 -984 1481 -978
rect 1485 -984 1488 -978
rect 1492 -984 1495 -978
rect 1499 -984 1502 -978
rect 1506 -984 1509 -978
rect 1513 -984 1516 -978
rect 1520 -984 1523 -978
rect 1527 -984 1530 -978
rect 1534 -984 1537 -978
rect 1541 -984 1544 -978
rect 1548 -984 1551 -978
rect 1555 -984 1558 -978
rect 1562 -984 1565 -978
rect 1569 -984 1572 -978
rect 1576 -984 1579 -978
rect 1583 -984 1586 -978
rect 1590 -984 1593 -978
rect 1597 -984 1600 -978
rect 1604 -984 1607 -978
rect 1611 -984 1614 -978
rect 1618 -984 1621 -978
rect 1625 -984 1628 -978
rect 1632 -984 1635 -978
rect 1639 -984 1642 -978
rect 1646 -984 1649 -978
rect 1653 -984 1656 -978
rect 1660 -984 1663 -978
rect 1667 -984 1670 -978
rect 1674 -984 1677 -978
rect 1681 -984 1684 -978
rect 1688 -984 1691 -978
rect 1695 -984 1698 -978
rect 1702 -984 1705 -978
rect 1709 -984 1712 -978
rect 1716 -984 1719 -978
rect 1723 -984 1726 -978
rect 1730 -984 1733 -978
rect 1737 -984 1740 -978
rect 1744 -984 1747 -978
rect 1751 -984 1754 -978
rect 1758 -984 1761 -978
rect 1765 -984 1768 -978
rect 1772 -984 1775 -978
rect 1779 -984 1782 -978
rect 1786 -984 1789 -978
rect 1793 -984 1796 -978
rect 1800 -984 1803 -978
rect 1807 -984 1810 -978
rect 1814 -984 1817 -978
rect 1821 -984 1824 -978
rect 1828 -984 1831 -978
rect 1835 -984 1838 -978
rect 1842 -984 1845 -978
rect 1849 -984 1852 -978
rect 1856 -984 1859 -978
rect 1863 -984 1866 -978
rect 1870 -984 1873 -978
rect 1877 -984 1883 -978
rect 1884 -984 1887 -978
rect 1891 -984 1894 -978
rect 1898 -984 1904 -978
rect 1905 -984 1908 -978
rect 1912 -984 1918 -978
rect 1919 -984 1925 -978
rect 1926 -984 1929 -978
rect 1933 -984 1936 -978
rect 1940 -984 1943 -978
rect 1947 -984 1950 -978
rect 1954 -984 1957 -978
rect 1 -1115 7 -1109
rect 8 -1115 11 -1109
rect 15 -1115 18 -1109
rect 22 -1115 25 -1109
rect 29 -1115 32 -1109
rect 36 -1115 39 -1109
rect 43 -1115 49 -1109
rect 50 -1115 53 -1109
rect 57 -1115 60 -1109
rect 64 -1115 70 -1109
rect 71 -1115 74 -1109
rect 78 -1115 84 -1109
rect 85 -1115 88 -1109
rect 92 -1115 95 -1109
rect 99 -1115 102 -1109
rect 106 -1115 109 -1109
rect 113 -1115 116 -1109
rect 120 -1115 123 -1109
rect 127 -1115 133 -1109
rect 134 -1115 137 -1109
rect 141 -1115 144 -1109
rect 148 -1115 151 -1109
rect 155 -1115 158 -1109
rect 162 -1115 165 -1109
rect 169 -1115 172 -1109
rect 176 -1115 179 -1109
rect 183 -1115 186 -1109
rect 190 -1115 193 -1109
rect 197 -1115 200 -1109
rect 204 -1115 207 -1109
rect 211 -1115 217 -1109
rect 218 -1115 224 -1109
rect 225 -1115 228 -1109
rect 232 -1115 235 -1109
rect 239 -1115 242 -1109
rect 246 -1115 249 -1109
rect 253 -1115 256 -1109
rect 260 -1115 263 -1109
rect 267 -1115 270 -1109
rect 274 -1115 277 -1109
rect 281 -1115 284 -1109
rect 288 -1115 291 -1109
rect 295 -1115 298 -1109
rect 302 -1115 305 -1109
rect 309 -1115 315 -1109
rect 316 -1115 319 -1109
rect 323 -1115 326 -1109
rect 330 -1115 333 -1109
rect 337 -1115 340 -1109
rect 344 -1115 347 -1109
rect 351 -1115 354 -1109
rect 358 -1115 361 -1109
rect 365 -1115 368 -1109
rect 372 -1115 375 -1109
rect 379 -1115 382 -1109
rect 386 -1115 389 -1109
rect 393 -1115 399 -1109
rect 400 -1115 403 -1109
rect 407 -1115 410 -1109
rect 414 -1115 417 -1109
rect 421 -1115 424 -1109
rect 428 -1115 431 -1109
rect 435 -1115 438 -1109
rect 442 -1115 445 -1109
rect 449 -1115 455 -1109
rect 456 -1115 459 -1109
rect 463 -1115 466 -1109
rect 470 -1115 473 -1109
rect 477 -1115 480 -1109
rect 484 -1115 487 -1109
rect 491 -1115 494 -1109
rect 498 -1115 501 -1109
rect 505 -1115 508 -1109
rect 512 -1115 515 -1109
rect 519 -1115 525 -1109
rect 526 -1115 529 -1109
rect 533 -1115 536 -1109
rect 540 -1115 543 -1109
rect 547 -1115 550 -1109
rect 554 -1115 557 -1109
rect 561 -1115 567 -1109
rect 568 -1115 574 -1109
rect 575 -1115 581 -1109
rect 582 -1115 585 -1109
rect 589 -1115 592 -1109
rect 596 -1115 599 -1109
rect 603 -1115 606 -1109
rect 610 -1115 613 -1109
rect 617 -1115 620 -1109
rect 624 -1115 630 -1109
rect 631 -1115 637 -1109
rect 638 -1115 641 -1109
rect 645 -1115 651 -1109
rect 652 -1115 658 -1109
rect 659 -1115 662 -1109
rect 666 -1115 669 -1109
rect 673 -1115 676 -1109
rect 680 -1115 686 -1109
rect 687 -1115 690 -1109
rect 694 -1115 697 -1109
rect 701 -1115 704 -1109
rect 708 -1115 711 -1109
rect 715 -1115 718 -1109
rect 722 -1115 725 -1109
rect 729 -1115 735 -1109
rect 736 -1115 742 -1109
rect 743 -1115 746 -1109
rect 750 -1115 756 -1109
rect 757 -1115 763 -1109
rect 764 -1115 767 -1109
rect 771 -1115 774 -1109
rect 778 -1115 784 -1109
rect 785 -1115 791 -1109
rect 792 -1115 795 -1109
rect 799 -1115 802 -1109
rect 806 -1115 809 -1109
rect 813 -1115 816 -1109
rect 820 -1115 823 -1109
rect 827 -1115 830 -1109
rect 834 -1115 837 -1109
rect 841 -1115 844 -1109
rect 848 -1115 854 -1109
rect 855 -1115 858 -1109
rect 862 -1115 868 -1109
rect 869 -1115 872 -1109
rect 876 -1115 879 -1109
rect 883 -1115 886 -1109
rect 890 -1115 896 -1109
rect 897 -1115 900 -1109
rect 904 -1115 907 -1109
rect 911 -1115 914 -1109
rect 918 -1115 921 -1109
rect 925 -1115 928 -1109
rect 932 -1115 935 -1109
rect 939 -1115 942 -1109
rect 946 -1115 949 -1109
rect 953 -1115 959 -1109
rect 960 -1115 963 -1109
rect 967 -1115 970 -1109
rect 974 -1115 977 -1109
rect 981 -1115 984 -1109
rect 988 -1115 991 -1109
rect 995 -1115 998 -1109
rect 1002 -1115 1005 -1109
rect 1009 -1115 1012 -1109
rect 1016 -1115 1022 -1109
rect 1023 -1115 1026 -1109
rect 1030 -1115 1033 -1109
rect 1037 -1115 1040 -1109
rect 1044 -1115 1050 -1109
rect 1051 -1115 1054 -1109
rect 1058 -1115 1061 -1109
rect 1065 -1115 1068 -1109
rect 1072 -1115 1075 -1109
rect 1079 -1115 1082 -1109
rect 1086 -1115 1089 -1109
rect 1093 -1115 1096 -1109
rect 1100 -1115 1103 -1109
rect 1107 -1115 1110 -1109
rect 1114 -1115 1117 -1109
rect 1121 -1115 1124 -1109
rect 1128 -1115 1131 -1109
rect 1135 -1115 1141 -1109
rect 1142 -1115 1145 -1109
rect 1149 -1115 1155 -1109
rect 1156 -1115 1159 -1109
rect 1163 -1115 1166 -1109
rect 1170 -1115 1173 -1109
rect 1177 -1115 1180 -1109
rect 1184 -1115 1187 -1109
rect 1191 -1115 1194 -1109
rect 1198 -1115 1201 -1109
rect 1205 -1115 1208 -1109
rect 1212 -1115 1215 -1109
rect 1219 -1115 1222 -1109
rect 1226 -1115 1232 -1109
rect 1233 -1115 1236 -1109
rect 1240 -1115 1243 -1109
rect 1247 -1115 1250 -1109
rect 1254 -1115 1257 -1109
rect 1261 -1115 1264 -1109
rect 1268 -1115 1271 -1109
rect 1275 -1115 1278 -1109
rect 1282 -1115 1285 -1109
rect 1289 -1115 1292 -1109
rect 1296 -1115 1299 -1109
rect 1303 -1115 1306 -1109
rect 1310 -1115 1313 -1109
rect 1317 -1115 1320 -1109
rect 1324 -1115 1327 -1109
rect 1331 -1115 1334 -1109
rect 1338 -1115 1341 -1109
rect 1345 -1115 1348 -1109
rect 1352 -1115 1355 -1109
rect 1359 -1115 1362 -1109
rect 1366 -1115 1369 -1109
rect 1373 -1115 1376 -1109
rect 1380 -1115 1383 -1109
rect 1387 -1115 1390 -1109
rect 1394 -1115 1397 -1109
rect 1401 -1115 1404 -1109
rect 1408 -1115 1411 -1109
rect 1415 -1115 1418 -1109
rect 1422 -1115 1425 -1109
rect 1429 -1115 1432 -1109
rect 1436 -1115 1439 -1109
rect 1443 -1115 1446 -1109
rect 1450 -1115 1453 -1109
rect 1457 -1115 1460 -1109
rect 1464 -1115 1467 -1109
rect 1471 -1115 1474 -1109
rect 1478 -1115 1481 -1109
rect 1485 -1115 1488 -1109
rect 1492 -1115 1495 -1109
rect 1499 -1115 1502 -1109
rect 1506 -1115 1509 -1109
rect 1513 -1115 1516 -1109
rect 1520 -1115 1523 -1109
rect 1527 -1115 1530 -1109
rect 1534 -1115 1537 -1109
rect 1541 -1115 1544 -1109
rect 1548 -1115 1551 -1109
rect 1555 -1115 1558 -1109
rect 1562 -1115 1565 -1109
rect 1569 -1115 1572 -1109
rect 1576 -1115 1579 -1109
rect 1583 -1115 1586 -1109
rect 1590 -1115 1593 -1109
rect 1597 -1115 1600 -1109
rect 1604 -1115 1607 -1109
rect 1611 -1115 1614 -1109
rect 1618 -1115 1621 -1109
rect 1625 -1115 1628 -1109
rect 1632 -1115 1635 -1109
rect 1639 -1115 1642 -1109
rect 1646 -1115 1649 -1109
rect 1653 -1115 1656 -1109
rect 1660 -1115 1663 -1109
rect 1667 -1115 1670 -1109
rect 1674 -1115 1677 -1109
rect 1681 -1115 1684 -1109
rect 1688 -1115 1691 -1109
rect 1695 -1115 1698 -1109
rect 1702 -1115 1705 -1109
rect 1709 -1115 1712 -1109
rect 1716 -1115 1719 -1109
rect 1723 -1115 1726 -1109
rect 1730 -1115 1733 -1109
rect 1737 -1115 1740 -1109
rect 1744 -1115 1747 -1109
rect 1751 -1115 1754 -1109
rect 1758 -1115 1761 -1109
rect 1765 -1115 1768 -1109
rect 1772 -1115 1775 -1109
rect 1779 -1115 1782 -1109
rect 1786 -1115 1789 -1109
rect 1793 -1115 1796 -1109
rect 1800 -1115 1803 -1109
rect 1807 -1115 1810 -1109
rect 1814 -1115 1817 -1109
rect 1821 -1115 1824 -1109
rect 1828 -1115 1831 -1109
rect 1835 -1115 1838 -1109
rect 1842 -1115 1845 -1109
rect 1849 -1115 1852 -1109
rect 1856 -1115 1859 -1109
rect 1863 -1115 1869 -1109
rect 1870 -1115 1873 -1109
rect 1877 -1115 1880 -1109
rect 1926 -1115 1929 -1109
rect 1947 -1115 1950 -1109
rect 1961 -1115 1964 -1109
rect 1968 -1115 1971 -1109
rect 1975 -1115 1978 -1109
rect 1 -1250 4 -1244
rect 8 -1250 11 -1244
rect 15 -1250 18 -1244
rect 22 -1250 28 -1244
rect 29 -1250 32 -1244
rect 36 -1250 42 -1244
rect 43 -1250 46 -1244
rect 50 -1250 53 -1244
rect 57 -1250 63 -1244
rect 64 -1250 67 -1244
rect 71 -1250 74 -1244
rect 78 -1250 84 -1244
rect 85 -1250 88 -1244
rect 92 -1250 95 -1244
rect 99 -1250 102 -1244
rect 106 -1250 109 -1244
rect 113 -1250 116 -1244
rect 120 -1250 126 -1244
rect 127 -1250 130 -1244
rect 134 -1250 137 -1244
rect 141 -1250 144 -1244
rect 148 -1250 151 -1244
rect 155 -1250 161 -1244
rect 162 -1250 165 -1244
rect 169 -1250 175 -1244
rect 176 -1250 182 -1244
rect 183 -1250 186 -1244
rect 190 -1250 193 -1244
rect 197 -1250 200 -1244
rect 204 -1250 207 -1244
rect 211 -1250 214 -1244
rect 218 -1250 221 -1244
rect 225 -1250 231 -1244
rect 232 -1250 235 -1244
rect 239 -1250 242 -1244
rect 246 -1250 249 -1244
rect 253 -1250 256 -1244
rect 260 -1250 266 -1244
rect 267 -1250 270 -1244
rect 274 -1250 277 -1244
rect 281 -1250 284 -1244
rect 288 -1250 294 -1244
rect 295 -1250 298 -1244
rect 302 -1250 305 -1244
rect 309 -1250 312 -1244
rect 316 -1250 319 -1244
rect 323 -1250 326 -1244
rect 330 -1250 333 -1244
rect 337 -1250 340 -1244
rect 344 -1250 347 -1244
rect 351 -1250 354 -1244
rect 358 -1250 361 -1244
rect 365 -1250 368 -1244
rect 372 -1250 375 -1244
rect 379 -1250 382 -1244
rect 386 -1250 389 -1244
rect 393 -1250 396 -1244
rect 400 -1250 403 -1244
rect 407 -1250 410 -1244
rect 414 -1250 417 -1244
rect 421 -1250 427 -1244
rect 428 -1250 431 -1244
rect 435 -1250 438 -1244
rect 442 -1250 448 -1244
rect 449 -1250 455 -1244
rect 456 -1250 459 -1244
rect 463 -1250 466 -1244
rect 470 -1250 476 -1244
rect 477 -1250 480 -1244
rect 484 -1250 487 -1244
rect 491 -1250 494 -1244
rect 498 -1250 501 -1244
rect 505 -1250 508 -1244
rect 512 -1250 518 -1244
rect 519 -1250 522 -1244
rect 526 -1250 529 -1244
rect 533 -1250 536 -1244
rect 540 -1250 543 -1244
rect 547 -1250 550 -1244
rect 554 -1250 557 -1244
rect 561 -1250 567 -1244
rect 568 -1250 571 -1244
rect 575 -1250 578 -1244
rect 582 -1250 588 -1244
rect 589 -1250 592 -1244
rect 596 -1250 599 -1244
rect 603 -1250 606 -1244
rect 610 -1250 613 -1244
rect 617 -1250 620 -1244
rect 624 -1250 627 -1244
rect 631 -1250 634 -1244
rect 638 -1250 641 -1244
rect 645 -1250 648 -1244
rect 652 -1250 655 -1244
rect 659 -1250 662 -1244
rect 666 -1250 672 -1244
rect 673 -1250 676 -1244
rect 680 -1250 683 -1244
rect 687 -1250 690 -1244
rect 694 -1250 697 -1244
rect 701 -1250 704 -1244
rect 708 -1250 711 -1244
rect 715 -1250 718 -1244
rect 722 -1250 725 -1244
rect 729 -1250 732 -1244
rect 736 -1250 739 -1244
rect 743 -1250 746 -1244
rect 750 -1250 753 -1244
rect 757 -1250 760 -1244
rect 764 -1250 767 -1244
rect 771 -1250 777 -1244
rect 778 -1250 784 -1244
rect 785 -1250 788 -1244
rect 792 -1250 798 -1244
rect 799 -1250 802 -1244
rect 806 -1250 812 -1244
rect 813 -1250 816 -1244
rect 820 -1250 826 -1244
rect 827 -1250 830 -1244
rect 834 -1250 837 -1244
rect 841 -1250 844 -1244
rect 848 -1250 851 -1244
rect 855 -1250 861 -1244
rect 862 -1250 865 -1244
rect 869 -1250 875 -1244
rect 876 -1250 882 -1244
rect 883 -1250 886 -1244
rect 890 -1250 893 -1244
rect 897 -1250 900 -1244
rect 904 -1250 910 -1244
rect 911 -1250 914 -1244
rect 918 -1250 921 -1244
rect 925 -1250 931 -1244
rect 932 -1250 935 -1244
rect 939 -1250 942 -1244
rect 946 -1250 949 -1244
rect 953 -1250 956 -1244
rect 960 -1250 966 -1244
rect 967 -1250 970 -1244
rect 974 -1250 977 -1244
rect 981 -1250 984 -1244
rect 988 -1250 991 -1244
rect 995 -1250 998 -1244
rect 1002 -1250 1005 -1244
rect 1009 -1250 1012 -1244
rect 1016 -1250 1022 -1244
rect 1023 -1250 1026 -1244
rect 1030 -1250 1033 -1244
rect 1037 -1250 1040 -1244
rect 1044 -1250 1050 -1244
rect 1051 -1250 1054 -1244
rect 1058 -1250 1061 -1244
rect 1065 -1250 1068 -1244
rect 1072 -1250 1075 -1244
rect 1079 -1250 1082 -1244
rect 1086 -1250 1089 -1244
rect 1093 -1250 1096 -1244
rect 1100 -1250 1103 -1244
rect 1107 -1250 1110 -1244
rect 1114 -1250 1117 -1244
rect 1121 -1250 1124 -1244
rect 1128 -1250 1134 -1244
rect 1135 -1250 1138 -1244
rect 1142 -1250 1145 -1244
rect 1149 -1250 1152 -1244
rect 1156 -1250 1162 -1244
rect 1163 -1250 1166 -1244
rect 1170 -1250 1173 -1244
rect 1177 -1250 1183 -1244
rect 1184 -1250 1187 -1244
rect 1191 -1250 1194 -1244
rect 1198 -1250 1201 -1244
rect 1205 -1250 1208 -1244
rect 1212 -1250 1215 -1244
rect 1219 -1250 1222 -1244
rect 1226 -1250 1229 -1244
rect 1233 -1250 1236 -1244
rect 1240 -1250 1243 -1244
rect 1247 -1250 1250 -1244
rect 1254 -1250 1257 -1244
rect 1261 -1250 1264 -1244
rect 1268 -1250 1271 -1244
rect 1275 -1250 1278 -1244
rect 1282 -1250 1285 -1244
rect 1289 -1250 1292 -1244
rect 1296 -1250 1299 -1244
rect 1303 -1250 1306 -1244
rect 1310 -1250 1313 -1244
rect 1317 -1250 1320 -1244
rect 1324 -1250 1327 -1244
rect 1331 -1250 1334 -1244
rect 1338 -1250 1341 -1244
rect 1345 -1250 1348 -1244
rect 1352 -1250 1355 -1244
rect 1359 -1250 1362 -1244
rect 1366 -1250 1369 -1244
rect 1373 -1250 1376 -1244
rect 1380 -1250 1383 -1244
rect 1387 -1250 1390 -1244
rect 1394 -1250 1397 -1244
rect 1401 -1250 1404 -1244
rect 1408 -1250 1411 -1244
rect 1415 -1250 1418 -1244
rect 1422 -1250 1425 -1244
rect 1429 -1250 1432 -1244
rect 1436 -1250 1439 -1244
rect 1443 -1250 1446 -1244
rect 1450 -1250 1453 -1244
rect 1457 -1250 1460 -1244
rect 1464 -1250 1467 -1244
rect 1471 -1250 1474 -1244
rect 1478 -1250 1481 -1244
rect 1485 -1250 1488 -1244
rect 1492 -1250 1495 -1244
rect 1499 -1250 1502 -1244
rect 1506 -1250 1509 -1244
rect 1513 -1250 1516 -1244
rect 1520 -1250 1523 -1244
rect 1527 -1250 1530 -1244
rect 1534 -1250 1537 -1244
rect 1541 -1250 1544 -1244
rect 1548 -1250 1551 -1244
rect 1555 -1250 1558 -1244
rect 1562 -1250 1565 -1244
rect 1569 -1250 1572 -1244
rect 1576 -1250 1579 -1244
rect 1583 -1250 1586 -1244
rect 1590 -1250 1593 -1244
rect 1597 -1250 1600 -1244
rect 1604 -1250 1607 -1244
rect 1611 -1250 1614 -1244
rect 1618 -1250 1621 -1244
rect 1625 -1250 1628 -1244
rect 1632 -1250 1635 -1244
rect 1639 -1250 1642 -1244
rect 1646 -1250 1649 -1244
rect 1653 -1250 1656 -1244
rect 1660 -1250 1663 -1244
rect 1667 -1250 1670 -1244
rect 1674 -1250 1677 -1244
rect 1681 -1250 1684 -1244
rect 1688 -1250 1691 -1244
rect 1695 -1250 1698 -1244
rect 1702 -1250 1705 -1244
rect 1709 -1250 1712 -1244
rect 1716 -1250 1719 -1244
rect 1723 -1250 1726 -1244
rect 1730 -1250 1733 -1244
rect 1737 -1250 1740 -1244
rect 1744 -1250 1747 -1244
rect 1751 -1250 1754 -1244
rect 1758 -1250 1761 -1244
rect 1765 -1250 1768 -1244
rect 1772 -1250 1775 -1244
rect 1779 -1250 1782 -1244
rect 1786 -1250 1789 -1244
rect 1793 -1250 1796 -1244
rect 1800 -1250 1803 -1244
rect 1807 -1250 1810 -1244
rect 1814 -1250 1817 -1244
rect 1821 -1250 1824 -1244
rect 1828 -1250 1831 -1244
rect 1835 -1250 1838 -1244
rect 1842 -1250 1845 -1244
rect 1849 -1250 1852 -1244
rect 1856 -1250 1859 -1244
rect 1863 -1250 1866 -1244
rect 1870 -1250 1873 -1244
rect 1877 -1250 1880 -1244
rect 1884 -1250 1887 -1244
rect 1891 -1250 1894 -1244
rect 1898 -1250 1901 -1244
rect 1905 -1250 1908 -1244
rect 1912 -1250 1915 -1244
rect 1919 -1250 1922 -1244
rect 1926 -1250 1929 -1244
rect 1954 -1250 1957 -1244
rect 1961 -1250 1964 -1244
rect 1968 -1250 1971 -1244
rect 1975 -1250 1978 -1244
rect 1989 -1250 1992 -1244
rect 1 -1393 7 -1387
rect 8 -1393 11 -1387
rect 15 -1393 18 -1387
rect 22 -1393 25 -1387
rect 29 -1393 32 -1387
rect 36 -1393 39 -1387
rect 43 -1393 46 -1387
rect 50 -1393 56 -1387
rect 57 -1393 63 -1387
rect 64 -1393 67 -1387
rect 71 -1393 77 -1387
rect 78 -1393 81 -1387
rect 85 -1393 88 -1387
rect 92 -1393 95 -1387
rect 99 -1393 102 -1387
rect 106 -1393 112 -1387
rect 113 -1393 116 -1387
rect 120 -1393 123 -1387
rect 127 -1393 133 -1387
rect 134 -1393 137 -1387
rect 141 -1393 147 -1387
rect 148 -1393 154 -1387
rect 155 -1393 158 -1387
rect 162 -1393 168 -1387
rect 169 -1393 172 -1387
rect 176 -1393 179 -1387
rect 183 -1393 186 -1387
rect 190 -1393 193 -1387
rect 197 -1393 200 -1387
rect 204 -1393 210 -1387
rect 211 -1393 214 -1387
rect 218 -1393 221 -1387
rect 225 -1393 228 -1387
rect 232 -1393 235 -1387
rect 239 -1393 242 -1387
rect 246 -1393 249 -1387
rect 253 -1393 256 -1387
rect 260 -1393 263 -1387
rect 267 -1393 270 -1387
rect 274 -1393 277 -1387
rect 281 -1393 284 -1387
rect 288 -1393 291 -1387
rect 295 -1393 298 -1387
rect 302 -1393 305 -1387
rect 309 -1393 312 -1387
rect 316 -1393 319 -1387
rect 323 -1393 326 -1387
rect 330 -1393 333 -1387
rect 337 -1393 340 -1387
rect 344 -1393 347 -1387
rect 351 -1393 354 -1387
rect 358 -1393 361 -1387
rect 365 -1393 368 -1387
rect 372 -1393 375 -1387
rect 379 -1393 382 -1387
rect 386 -1393 389 -1387
rect 393 -1393 396 -1387
rect 400 -1393 403 -1387
rect 407 -1393 410 -1387
rect 414 -1393 417 -1387
rect 421 -1393 424 -1387
rect 428 -1393 434 -1387
rect 435 -1393 438 -1387
rect 442 -1393 445 -1387
rect 449 -1393 452 -1387
rect 456 -1393 459 -1387
rect 463 -1393 466 -1387
rect 470 -1393 473 -1387
rect 477 -1393 480 -1387
rect 484 -1393 487 -1387
rect 491 -1393 494 -1387
rect 498 -1393 501 -1387
rect 505 -1393 508 -1387
rect 512 -1393 515 -1387
rect 519 -1393 522 -1387
rect 526 -1393 532 -1387
rect 533 -1393 536 -1387
rect 540 -1393 543 -1387
rect 547 -1393 550 -1387
rect 554 -1393 557 -1387
rect 561 -1393 564 -1387
rect 568 -1393 571 -1387
rect 575 -1393 581 -1387
rect 582 -1393 585 -1387
rect 589 -1393 592 -1387
rect 596 -1393 599 -1387
rect 603 -1393 606 -1387
rect 610 -1393 613 -1387
rect 617 -1393 620 -1387
rect 624 -1393 630 -1387
rect 631 -1393 634 -1387
rect 638 -1393 641 -1387
rect 645 -1393 648 -1387
rect 652 -1393 658 -1387
rect 659 -1393 662 -1387
rect 666 -1393 672 -1387
rect 673 -1393 679 -1387
rect 680 -1393 683 -1387
rect 687 -1393 690 -1387
rect 694 -1393 697 -1387
rect 701 -1393 704 -1387
rect 708 -1393 714 -1387
rect 715 -1393 718 -1387
rect 722 -1393 725 -1387
rect 729 -1393 732 -1387
rect 736 -1393 739 -1387
rect 743 -1393 746 -1387
rect 750 -1393 753 -1387
rect 757 -1393 760 -1387
rect 764 -1393 767 -1387
rect 771 -1393 774 -1387
rect 778 -1393 781 -1387
rect 785 -1393 788 -1387
rect 792 -1393 795 -1387
rect 799 -1393 802 -1387
rect 806 -1393 809 -1387
rect 813 -1393 816 -1387
rect 820 -1393 823 -1387
rect 827 -1393 830 -1387
rect 834 -1393 840 -1387
rect 841 -1393 844 -1387
rect 848 -1393 851 -1387
rect 855 -1393 861 -1387
rect 862 -1393 865 -1387
rect 869 -1393 872 -1387
rect 876 -1393 879 -1387
rect 883 -1393 886 -1387
rect 890 -1393 893 -1387
rect 897 -1393 900 -1387
rect 904 -1393 907 -1387
rect 911 -1393 914 -1387
rect 918 -1393 924 -1387
rect 925 -1393 931 -1387
rect 932 -1393 935 -1387
rect 939 -1393 945 -1387
rect 946 -1393 949 -1387
rect 953 -1393 956 -1387
rect 960 -1393 963 -1387
rect 967 -1393 973 -1387
rect 974 -1393 977 -1387
rect 981 -1393 984 -1387
rect 988 -1393 991 -1387
rect 995 -1393 1001 -1387
rect 1002 -1393 1005 -1387
rect 1009 -1393 1012 -1387
rect 1016 -1393 1019 -1387
rect 1023 -1393 1026 -1387
rect 1030 -1393 1036 -1387
rect 1037 -1393 1040 -1387
rect 1044 -1393 1047 -1387
rect 1051 -1393 1057 -1387
rect 1058 -1393 1061 -1387
rect 1065 -1393 1071 -1387
rect 1072 -1393 1078 -1387
rect 1079 -1393 1082 -1387
rect 1086 -1393 1089 -1387
rect 1093 -1393 1096 -1387
rect 1100 -1393 1103 -1387
rect 1107 -1393 1113 -1387
rect 1114 -1393 1117 -1387
rect 1121 -1393 1124 -1387
rect 1128 -1393 1131 -1387
rect 1135 -1393 1138 -1387
rect 1142 -1393 1145 -1387
rect 1149 -1393 1152 -1387
rect 1156 -1393 1159 -1387
rect 1163 -1393 1166 -1387
rect 1170 -1393 1176 -1387
rect 1177 -1393 1180 -1387
rect 1184 -1393 1190 -1387
rect 1191 -1393 1194 -1387
rect 1198 -1393 1201 -1387
rect 1205 -1393 1208 -1387
rect 1212 -1393 1215 -1387
rect 1219 -1393 1222 -1387
rect 1226 -1393 1229 -1387
rect 1233 -1393 1236 -1387
rect 1240 -1393 1246 -1387
rect 1247 -1393 1250 -1387
rect 1254 -1393 1257 -1387
rect 1261 -1393 1264 -1387
rect 1268 -1393 1271 -1387
rect 1275 -1393 1278 -1387
rect 1282 -1393 1288 -1387
rect 1289 -1393 1292 -1387
rect 1296 -1393 1299 -1387
rect 1303 -1393 1306 -1387
rect 1310 -1393 1313 -1387
rect 1317 -1393 1320 -1387
rect 1324 -1393 1327 -1387
rect 1331 -1393 1334 -1387
rect 1338 -1393 1341 -1387
rect 1345 -1393 1348 -1387
rect 1352 -1393 1355 -1387
rect 1359 -1393 1362 -1387
rect 1366 -1393 1369 -1387
rect 1373 -1393 1376 -1387
rect 1380 -1393 1383 -1387
rect 1387 -1393 1390 -1387
rect 1394 -1393 1397 -1387
rect 1401 -1393 1404 -1387
rect 1408 -1393 1411 -1387
rect 1415 -1393 1418 -1387
rect 1422 -1393 1425 -1387
rect 1429 -1393 1432 -1387
rect 1436 -1393 1439 -1387
rect 1443 -1393 1446 -1387
rect 1450 -1393 1453 -1387
rect 1457 -1393 1460 -1387
rect 1464 -1393 1467 -1387
rect 1471 -1393 1474 -1387
rect 1478 -1393 1481 -1387
rect 1485 -1393 1488 -1387
rect 1492 -1393 1495 -1387
rect 1499 -1393 1502 -1387
rect 1506 -1393 1509 -1387
rect 1513 -1393 1516 -1387
rect 1520 -1393 1523 -1387
rect 1527 -1393 1530 -1387
rect 1534 -1393 1537 -1387
rect 1541 -1393 1544 -1387
rect 1548 -1393 1551 -1387
rect 1555 -1393 1558 -1387
rect 1562 -1393 1565 -1387
rect 1569 -1393 1572 -1387
rect 1576 -1393 1579 -1387
rect 1583 -1393 1586 -1387
rect 1590 -1393 1593 -1387
rect 1597 -1393 1600 -1387
rect 1604 -1393 1607 -1387
rect 1611 -1393 1614 -1387
rect 1618 -1393 1621 -1387
rect 1625 -1393 1628 -1387
rect 1632 -1393 1635 -1387
rect 1639 -1393 1642 -1387
rect 1646 -1393 1649 -1387
rect 1653 -1393 1656 -1387
rect 1660 -1393 1663 -1387
rect 1667 -1393 1670 -1387
rect 1674 -1393 1677 -1387
rect 1681 -1393 1684 -1387
rect 1688 -1393 1691 -1387
rect 1695 -1393 1698 -1387
rect 1702 -1393 1705 -1387
rect 1709 -1393 1712 -1387
rect 1716 -1393 1719 -1387
rect 1723 -1393 1726 -1387
rect 1730 -1393 1733 -1387
rect 1737 -1393 1740 -1387
rect 1744 -1393 1747 -1387
rect 1751 -1393 1754 -1387
rect 1758 -1393 1761 -1387
rect 1765 -1393 1768 -1387
rect 1772 -1393 1775 -1387
rect 1779 -1393 1782 -1387
rect 1786 -1393 1789 -1387
rect 1793 -1393 1796 -1387
rect 1800 -1393 1803 -1387
rect 1807 -1393 1810 -1387
rect 1814 -1393 1817 -1387
rect 1821 -1393 1824 -1387
rect 1828 -1393 1831 -1387
rect 1835 -1393 1838 -1387
rect 1842 -1393 1845 -1387
rect 1849 -1393 1852 -1387
rect 1856 -1393 1859 -1387
rect 1863 -1393 1866 -1387
rect 1870 -1393 1873 -1387
rect 1877 -1393 1880 -1387
rect 1884 -1393 1887 -1387
rect 1891 -1393 1894 -1387
rect 1898 -1393 1901 -1387
rect 1905 -1393 1908 -1387
rect 1912 -1393 1918 -1387
rect 1919 -1393 1922 -1387
rect 1926 -1393 1929 -1387
rect 1933 -1393 1936 -1387
rect 1940 -1393 1943 -1387
rect 1947 -1393 1950 -1387
rect 1968 -1393 1971 -1387
rect 1975 -1393 1978 -1387
rect 1982 -1393 1985 -1387
rect 1989 -1393 1992 -1387
rect 1996 -1393 1999 -1387
rect 1 -1524 4 -1518
rect 8 -1524 11 -1518
rect 15 -1524 18 -1518
rect 22 -1524 25 -1518
rect 29 -1524 32 -1518
rect 36 -1524 39 -1518
rect 43 -1524 49 -1518
rect 50 -1524 53 -1518
rect 57 -1524 63 -1518
rect 64 -1524 67 -1518
rect 71 -1524 74 -1518
rect 78 -1524 84 -1518
rect 85 -1524 88 -1518
rect 92 -1524 95 -1518
rect 99 -1524 102 -1518
rect 106 -1524 109 -1518
rect 113 -1524 116 -1518
rect 120 -1524 123 -1518
rect 127 -1524 130 -1518
rect 134 -1524 137 -1518
rect 141 -1524 147 -1518
rect 148 -1524 151 -1518
rect 155 -1524 158 -1518
rect 162 -1524 165 -1518
rect 169 -1524 172 -1518
rect 176 -1524 179 -1518
rect 183 -1524 186 -1518
rect 190 -1524 196 -1518
rect 197 -1524 200 -1518
rect 204 -1524 207 -1518
rect 211 -1524 217 -1518
rect 218 -1524 221 -1518
rect 225 -1524 228 -1518
rect 232 -1524 238 -1518
rect 239 -1524 245 -1518
rect 246 -1524 249 -1518
rect 253 -1524 256 -1518
rect 260 -1524 263 -1518
rect 267 -1524 270 -1518
rect 274 -1524 277 -1518
rect 281 -1524 284 -1518
rect 288 -1524 291 -1518
rect 295 -1524 298 -1518
rect 302 -1524 305 -1518
rect 309 -1524 312 -1518
rect 316 -1524 319 -1518
rect 323 -1524 326 -1518
rect 330 -1524 333 -1518
rect 337 -1524 340 -1518
rect 344 -1524 347 -1518
rect 351 -1524 354 -1518
rect 358 -1524 361 -1518
rect 365 -1524 368 -1518
rect 372 -1524 375 -1518
rect 379 -1524 382 -1518
rect 386 -1524 389 -1518
rect 393 -1524 396 -1518
rect 400 -1524 403 -1518
rect 407 -1524 410 -1518
rect 414 -1524 417 -1518
rect 421 -1524 424 -1518
rect 428 -1524 431 -1518
rect 435 -1524 438 -1518
rect 442 -1524 445 -1518
rect 449 -1524 452 -1518
rect 456 -1524 459 -1518
rect 463 -1524 466 -1518
rect 470 -1524 473 -1518
rect 477 -1524 480 -1518
rect 484 -1524 487 -1518
rect 491 -1524 494 -1518
rect 498 -1524 504 -1518
rect 505 -1524 508 -1518
rect 512 -1524 515 -1518
rect 519 -1524 522 -1518
rect 526 -1524 529 -1518
rect 533 -1524 536 -1518
rect 540 -1524 543 -1518
rect 547 -1524 550 -1518
rect 554 -1524 557 -1518
rect 561 -1524 564 -1518
rect 568 -1524 571 -1518
rect 575 -1524 578 -1518
rect 582 -1524 585 -1518
rect 589 -1524 595 -1518
rect 596 -1524 599 -1518
rect 603 -1524 606 -1518
rect 610 -1524 613 -1518
rect 617 -1524 620 -1518
rect 624 -1524 630 -1518
rect 631 -1524 634 -1518
rect 638 -1524 641 -1518
rect 645 -1524 648 -1518
rect 652 -1524 655 -1518
rect 659 -1524 665 -1518
rect 666 -1524 672 -1518
rect 673 -1524 676 -1518
rect 680 -1524 683 -1518
rect 687 -1524 690 -1518
rect 694 -1524 697 -1518
rect 701 -1524 704 -1518
rect 708 -1524 714 -1518
rect 715 -1524 718 -1518
rect 722 -1524 725 -1518
rect 729 -1524 732 -1518
rect 736 -1524 739 -1518
rect 743 -1524 746 -1518
rect 750 -1524 756 -1518
rect 757 -1524 760 -1518
rect 764 -1524 767 -1518
rect 771 -1524 774 -1518
rect 778 -1524 781 -1518
rect 785 -1524 788 -1518
rect 792 -1524 795 -1518
rect 799 -1524 802 -1518
rect 806 -1524 809 -1518
rect 813 -1524 816 -1518
rect 820 -1524 823 -1518
rect 827 -1524 830 -1518
rect 834 -1524 837 -1518
rect 841 -1524 844 -1518
rect 848 -1524 851 -1518
rect 855 -1524 858 -1518
rect 862 -1524 865 -1518
rect 869 -1524 872 -1518
rect 876 -1524 879 -1518
rect 883 -1524 886 -1518
rect 890 -1524 893 -1518
rect 897 -1524 900 -1518
rect 904 -1524 907 -1518
rect 911 -1524 914 -1518
rect 918 -1524 924 -1518
rect 925 -1524 928 -1518
rect 932 -1524 935 -1518
rect 939 -1524 942 -1518
rect 946 -1524 952 -1518
rect 953 -1524 959 -1518
rect 960 -1524 966 -1518
rect 967 -1524 970 -1518
rect 974 -1524 977 -1518
rect 981 -1524 987 -1518
rect 988 -1524 991 -1518
rect 995 -1524 998 -1518
rect 1002 -1524 1008 -1518
rect 1009 -1524 1012 -1518
rect 1016 -1524 1019 -1518
rect 1023 -1524 1026 -1518
rect 1030 -1524 1033 -1518
rect 1037 -1524 1040 -1518
rect 1044 -1524 1047 -1518
rect 1051 -1524 1054 -1518
rect 1058 -1524 1061 -1518
rect 1065 -1524 1071 -1518
rect 1072 -1524 1075 -1518
rect 1079 -1524 1082 -1518
rect 1086 -1524 1089 -1518
rect 1093 -1524 1096 -1518
rect 1100 -1524 1106 -1518
rect 1107 -1524 1113 -1518
rect 1114 -1524 1120 -1518
rect 1121 -1524 1124 -1518
rect 1128 -1524 1134 -1518
rect 1135 -1524 1138 -1518
rect 1142 -1524 1145 -1518
rect 1149 -1524 1152 -1518
rect 1156 -1524 1162 -1518
rect 1163 -1524 1166 -1518
rect 1170 -1524 1173 -1518
rect 1177 -1524 1180 -1518
rect 1184 -1524 1187 -1518
rect 1191 -1524 1197 -1518
rect 1198 -1524 1201 -1518
rect 1205 -1524 1208 -1518
rect 1212 -1524 1215 -1518
rect 1219 -1524 1222 -1518
rect 1226 -1524 1229 -1518
rect 1233 -1524 1236 -1518
rect 1240 -1524 1243 -1518
rect 1247 -1524 1250 -1518
rect 1254 -1524 1257 -1518
rect 1261 -1524 1267 -1518
rect 1268 -1524 1271 -1518
rect 1275 -1524 1278 -1518
rect 1282 -1524 1285 -1518
rect 1289 -1524 1292 -1518
rect 1296 -1524 1299 -1518
rect 1303 -1524 1309 -1518
rect 1310 -1524 1313 -1518
rect 1317 -1524 1320 -1518
rect 1324 -1524 1327 -1518
rect 1331 -1524 1337 -1518
rect 1338 -1524 1341 -1518
rect 1345 -1524 1348 -1518
rect 1352 -1524 1355 -1518
rect 1359 -1524 1362 -1518
rect 1366 -1524 1369 -1518
rect 1373 -1524 1376 -1518
rect 1380 -1524 1383 -1518
rect 1387 -1524 1390 -1518
rect 1394 -1524 1397 -1518
rect 1401 -1524 1404 -1518
rect 1408 -1524 1411 -1518
rect 1415 -1524 1418 -1518
rect 1422 -1524 1425 -1518
rect 1429 -1524 1432 -1518
rect 1436 -1524 1439 -1518
rect 1443 -1524 1446 -1518
rect 1450 -1524 1453 -1518
rect 1457 -1524 1460 -1518
rect 1464 -1524 1467 -1518
rect 1471 -1524 1474 -1518
rect 1478 -1524 1481 -1518
rect 1485 -1524 1488 -1518
rect 1492 -1524 1495 -1518
rect 1499 -1524 1502 -1518
rect 1506 -1524 1509 -1518
rect 1513 -1524 1516 -1518
rect 1520 -1524 1523 -1518
rect 1527 -1524 1530 -1518
rect 1534 -1524 1537 -1518
rect 1541 -1524 1544 -1518
rect 1548 -1524 1551 -1518
rect 1555 -1524 1558 -1518
rect 1562 -1524 1565 -1518
rect 1569 -1524 1572 -1518
rect 1576 -1524 1579 -1518
rect 1583 -1524 1586 -1518
rect 1590 -1524 1593 -1518
rect 1597 -1524 1600 -1518
rect 1604 -1524 1607 -1518
rect 1611 -1524 1614 -1518
rect 1618 -1524 1621 -1518
rect 1625 -1524 1628 -1518
rect 1632 -1524 1635 -1518
rect 1639 -1524 1642 -1518
rect 1646 -1524 1649 -1518
rect 1653 -1524 1656 -1518
rect 1660 -1524 1663 -1518
rect 1667 -1524 1670 -1518
rect 1674 -1524 1677 -1518
rect 1681 -1524 1684 -1518
rect 1688 -1524 1691 -1518
rect 1695 -1524 1698 -1518
rect 1702 -1524 1705 -1518
rect 1709 -1524 1712 -1518
rect 1716 -1524 1719 -1518
rect 1723 -1524 1726 -1518
rect 1730 -1524 1733 -1518
rect 1737 -1524 1740 -1518
rect 1744 -1524 1747 -1518
rect 1751 -1524 1754 -1518
rect 1758 -1524 1761 -1518
rect 1765 -1524 1768 -1518
rect 1772 -1524 1775 -1518
rect 1779 -1524 1782 -1518
rect 1786 -1524 1789 -1518
rect 1793 -1524 1796 -1518
rect 1800 -1524 1803 -1518
rect 1807 -1524 1810 -1518
rect 1814 -1524 1817 -1518
rect 1821 -1524 1824 -1518
rect 1828 -1524 1831 -1518
rect 1835 -1524 1838 -1518
rect 1842 -1524 1845 -1518
rect 1849 -1524 1852 -1518
rect 1856 -1524 1859 -1518
rect 1863 -1524 1866 -1518
rect 1870 -1524 1873 -1518
rect 1877 -1524 1880 -1518
rect 1884 -1524 1887 -1518
rect 1891 -1524 1894 -1518
rect 1898 -1524 1901 -1518
rect 1905 -1524 1908 -1518
rect 1912 -1524 1915 -1518
rect 1919 -1524 1922 -1518
rect 1926 -1524 1929 -1518
rect 1933 -1524 1936 -1518
rect 1940 -1524 1943 -1518
rect 1947 -1524 1950 -1518
rect 1954 -1524 1957 -1518
rect 1961 -1524 1964 -1518
rect 1968 -1524 1974 -1518
rect 1975 -1524 1981 -1518
rect 1982 -1524 1985 -1518
rect 1989 -1524 1992 -1518
rect 1996 -1524 2002 -1518
rect 2003 -1524 2009 -1518
rect 2010 -1524 2013 -1518
rect 2017 -1524 2020 -1518
rect 2024 -1524 2027 -1518
rect 1 -1651 4 -1645
rect 8 -1651 11 -1645
rect 15 -1651 18 -1645
rect 22 -1651 25 -1645
rect 29 -1651 32 -1645
rect 36 -1651 39 -1645
rect 43 -1651 46 -1645
rect 50 -1651 53 -1645
rect 57 -1651 60 -1645
rect 64 -1651 70 -1645
rect 71 -1651 74 -1645
rect 78 -1651 84 -1645
rect 85 -1651 91 -1645
rect 92 -1651 95 -1645
rect 99 -1651 102 -1645
rect 106 -1651 109 -1645
rect 113 -1651 119 -1645
rect 120 -1651 123 -1645
rect 127 -1651 130 -1645
rect 134 -1651 137 -1645
rect 141 -1651 147 -1645
rect 148 -1651 151 -1645
rect 155 -1651 158 -1645
rect 162 -1651 165 -1645
rect 169 -1651 175 -1645
rect 176 -1651 182 -1645
rect 183 -1651 186 -1645
rect 190 -1651 193 -1645
rect 197 -1651 200 -1645
rect 204 -1651 207 -1645
rect 211 -1651 214 -1645
rect 218 -1651 221 -1645
rect 225 -1651 228 -1645
rect 232 -1651 235 -1645
rect 239 -1651 242 -1645
rect 246 -1651 249 -1645
rect 253 -1651 256 -1645
rect 260 -1651 263 -1645
rect 267 -1651 270 -1645
rect 274 -1651 277 -1645
rect 281 -1651 284 -1645
rect 288 -1651 291 -1645
rect 295 -1651 298 -1645
rect 302 -1651 305 -1645
rect 309 -1651 312 -1645
rect 316 -1651 319 -1645
rect 323 -1651 326 -1645
rect 330 -1651 333 -1645
rect 337 -1651 340 -1645
rect 344 -1651 347 -1645
rect 351 -1651 354 -1645
rect 358 -1651 361 -1645
rect 365 -1651 368 -1645
rect 372 -1651 375 -1645
rect 379 -1651 382 -1645
rect 386 -1651 389 -1645
rect 393 -1651 399 -1645
rect 400 -1651 403 -1645
rect 407 -1651 410 -1645
rect 414 -1651 420 -1645
rect 421 -1651 424 -1645
rect 428 -1651 431 -1645
rect 435 -1651 438 -1645
rect 442 -1651 445 -1645
rect 449 -1651 452 -1645
rect 456 -1651 459 -1645
rect 463 -1651 466 -1645
rect 470 -1651 473 -1645
rect 477 -1651 480 -1645
rect 484 -1651 487 -1645
rect 491 -1651 494 -1645
rect 498 -1651 501 -1645
rect 505 -1651 508 -1645
rect 512 -1651 515 -1645
rect 519 -1651 522 -1645
rect 526 -1651 529 -1645
rect 533 -1651 536 -1645
rect 540 -1651 546 -1645
rect 547 -1651 550 -1645
rect 554 -1651 557 -1645
rect 561 -1651 564 -1645
rect 568 -1651 571 -1645
rect 575 -1651 578 -1645
rect 582 -1651 585 -1645
rect 589 -1651 592 -1645
rect 596 -1651 599 -1645
rect 603 -1651 606 -1645
rect 610 -1651 613 -1645
rect 617 -1651 620 -1645
rect 624 -1651 627 -1645
rect 631 -1651 634 -1645
rect 638 -1651 641 -1645
rect 645 -1651 648 -1645
rect 652 -1651 655 -1645
rect 659 -1651 665 -1645
rect 666 -1651 672 -1645
rect 673 -1651 676 -1645
rect 680 -1651 683 -1645
rect 687 -1651 690 -1645
rect 694 -1651 700 -1645
rect 701 -1651 704 -1645
rect 708 -1651 714 -1645
rect 715 -1651 718 -1645
rect 722 -1651 725 -1645
rect 729 -1651 732 -1645
rect 736 -1651 742 -1645
rect 743 -1651 746 -1645
rect 750 -1651 753 -1645
rect 757 -1651 760 -1645
rect 764 -1651 770 -1645
rect 771 -1651 774 -1645
rect 778 -1651 781 -1645
rect 785 -1651 788 -1645
rect 792 -1651 795 -1645
rect 799 -1651 802 -1645
rect 806 -1651 809 -1645
rect 813 -1651 819 -1645
rect 820 -1651 823 -1645
rect 827 -1651 833 -1645
rect 834 -1651 837 -1645
rect 841 -1651 844 -1645
rect 848 -1651 851 -1645
rect 855 -1651 858 -1645
rect 862 -1651 865 -1645
rect 869 -1651 872 -1645
rect 876 -1651 879 -1645
rect 883 -1651 886 -1645
rect 890 -1651 893 -1645
rect 897 -1651 900 -1645
rect 904 -1651 907 -1645
rect 911 -1651 914 -1645
rect 918 -1651 924 -1645
rect 925 -1651 928 -1645
rect 932 -1651 935 -1645
rect 939 -1651 945 -1645
rect 946 -1651 949 -1645
rect 953 -1651 956 -1645
rect 960 -1651 963 -1645
rect 967 -1651 973 -1645
rect 974 -1651 977 -1645
rect 981 -1651 984 -1645
rect 988 -1651 991 -1645
rect 995 -1651 998 -1645
rect 1002 -1651 1005 -1645
rect 1009 -1651 1012 -1645
rect 1016 -1651 1019 -1645
rect 1023 -1651 1026 -1645
rect 1030 -1651 1033 -1645
rect 1037 -1651 1043 -1645
rect 1044 -1651 1047 -1645
rect 1051 -1651 1057 -1645
rect 1058 -1651 1061 -1645
rect 1065 -1651 1068 -1645
rect 1072 -1651 1075 -1645
rect 1079 -1651 1082 -1645
rect 1086 -1651 1092 -1645
rect 1093 -1651 1096 -1645
rect 1100 -1651 1103 -1645
rect 1107 -1651 1110 -1645
rect 1114 -1651 1117 -1645
rect 1121 -1651 1124 -1645
rect 1128 -1651 1134 -1645
rect 1135 -1651 1138 -1645
rect 1142 -1651 1145 -1645
rect 1149 -1651 1152 -1645
rect 1156 -1651 1159 -1645
rect 1163 -1651 1166 -1645
rect 1170 -1651 1173 -1645
rect 1177 -1651 1180 -1645
rect 1184 -1651 1187 -1645
rect 1191 -1651 1194 -1645
rect 1198 -1651 1201 -1645
rect 1205 -1651 1211 -1645
rect 1212 -1651 1215 -1645
rect 1219 -1651 1222 -1645
rect 1226 -1651 1229 -1645
rect 1233 -1651 1236 -1645
rect 1240 -1651 1246 -1645
rect 1247 -1651 1250 -1645
rect 1254 -1651 1257 -1645
rect 1261 -1651 1264 -1645
rect 1268 -1651 1271 -1645
rect 1275 -1651 1278 -1645
rect 1282 -1651 1288 -1645
rect 1289 -1651 1292 -1645
rect 1296 -1651 1299 -1645
rect 1303 -1651 1309 -1645
rect 1310 -1651 1313 -1645
rect 1317 -1651 1320 -1645
rect 1324 -1651 1327 -1645
rect 1331 -1651 1337 -1645
rect 1338 -1651 1341 -1645
rect 1345 -1651 1348 -1645
rect 1352 -1651 1358 -1645
rect 1359 -1651 1362 -1645
rect 1366 -1651 1369 -1645
rect 1373 -1651 1376 -1645
rect 1380 -1651 1383 -1645
rect 1387 -1651 1390 -1645
rect 1394 -1651 1397 -1645
rect 1401 -1651 1404 -1645
rect 1408 -1651 1411 -1645
rect 1415 -1651 1418 -1645
rect 1422 -1651 1425 -1645
rect 1429 -1651 1432 -1645
rect 1436 -1651 1439 -1645
rect 1443 -1651 1446 -1645
rect 1450 -1651 1453 -1645
rect 1457 -1651 1460 -1645
rect 1464 -1651 1470 -1645
rect 1471 -1651 1474 -1645
rect 1478 -1651 1481 -1645
rect 1485 -1651 1488 -1645
rect 1492 -1651 1495 -1645
rect 1499 -1651 1505 -1645
rect 1506 -1651 1509 -1645
rect 1513 -1651 1516 -1645
rect 1520 -1651 1523 -1645
rect 1527 -1651 1530 -1645
rect 1534 -1651 1537 -1645
rect 1541 -1651 1544 -1645
rect 1548 -1651 1551 -1645
rect 1555 -1651 1558 -1645
rect 1562 -1651 1565 -1645
rect 1569 -1651 1572 -1645
rect 1576 -1651 1579 -1645
rect 1583 -1651 1586 -1645
rect 1590 -1651 1593 -1645
rect 1597 -1651 1600 -1645
rect 1604 -1651 1607 -1645
rect 1611 -1651 1614 -1645
rect 1618 -1651 1621 -1645
rect 1625 -1651 1628 -1645
rect 1632 -1651 1635 -1645
rect 1639 -1651 1642 -1645
rect 1646 -1651 1649 -1645
rect 1653 -1651 1656 -1645
rect 1660 -1651 1663 -1645
rect 1667 -1651 1670 -1645
rect 1674 -1651 1677 -1645
rect 1681 -1651 1684 -1645
rect 1688 -1651 1691 -1645
rect 1695 -1651 1698 -1645
rect 1702 -1651 1705 -1645
rect 1709 -1651 1712 -1645
rect 1716 -1651 1719 -1645
rect 1723 -1651 1726 -1645
rect 1730 -1651 1733 -1645
rect 1737 -1651 1740 -1645
rect 1744 -1651 1747 -1645
rect 1751 -1651 1754 -1645
rect 1758 -1651 1761 -1645
rect 1765 -1651 1768 -1645
rect 1772 -1651 1775 -1645
rect 1779 -1651 1782 -1645
rect 1786 -1651 1789 -1645
rect 1793 -1651 1796 -1645
rect 1800 -1651 1803 -1645
rect 1807 -1651 1810 -1645
rect 1814 -1651 1817 -1645
rect 1821 -1651 1824 -1645
rect 1828 -1651 1831 -1645
rect 1835 -1651 1838 -1645
rect 1842 -1651 1848 -1645
rect 1849 -1651 1852 -1645
rect 1856 -1651 1859 -1645
rect 1863 -1651 1866 -1645
rect 1870 -1651 1873 -1645
rect 1877 -1651 1883 -1645
rect 1884 -1651 1887 -1645
rect 1891 -1651 1894 -1645
rect 1898 -1651 1901 -1645
rect 1905 -1651 1908 -1645
rect 1912 -1651 1915 -1645
rect 1919 -1651 1922 -1645
rect 1926 -1651 1929 -1645
rect 1933 -1651 1936 -1645
rect 1940 -1651 1943 -1645
rect 1947 -1651 1950 -1645
rect 1975 -1651 1978 -1645
rect 2017 -1651 2020 -1645
rect 8 -1780 11 -1774
rect 15 -1780 18 -1774
rect 22 -1780 25 -1774
rect 29 -1780 32 -1774
rect 36 -1780 39 -1774
rect 43 -1780 46 -1774
rect 50 -1780 53 -1774
rect 57 -1780 60 -1774
rect 64 -1780 70 -1774
rect 71 -1780 74 -1774
rect 78 -1780 81 -1774
rect 85 -1780 88 -1774
rect 92 -1780 95 -1774
rect 99 -1780 102 -1774
rect 106 -1780 109 -1774
rect 113 -1780 116 -1774
rect 120 -1780 123 -1774
rect 127 -1780 133 -1774
rect 134 -1780 137 -1774
rect 141 -1780 144 -1774
rect 148 -1780 151 -1774
rect 155 -1780 158 -1774
rect 162 -1780 165 -1774
rect 169 -1780 172 -1774
rect 176 -1780 179 -1774
rect 183 -1780 189 -1774
rect 190 -1780 196 -1774
rect 197 -1780 203 -1774
rect 204 -1780 207 -1774
rect 211 -1780 214 -1774
rect 218 -1780 221 -1774
rect 225 -1780 228 -1774
rect 232 -1780 235 -1774
rect 239 -1780 242 -1774
rect 246 -1780 249 -1774
rect 253 -1780 256 -1774
rect 260 -1780 263 -1774
rect 267 -1780 270 -1774
rect 274 -1780 277 -1774
rect 281 -1780 284 -1774
rect 288 -1780 291 -1774
rect 295 -1780 298 -1774
rect 302 -1780 305 -1774
rect 309 -1780 312 -1774
rect 316 -1780 319 -1774
rect 323 -1780 326 -1774
rect 330 -1780 333 -1774
rect 337 -1780 340 -1774
rect 344 -1780 347 -1774
rect 351 -1780 354 -1774
rect 358 -1780 361 -1774
rect 365 -1780 368 -1774
rect 372 -1780 375 -1774
rect 379 -1780 382 -1774
rect 386 -1780 389 -1774
rect 393 -1780 399 -1774
rect 400 -1780 403 -1774
rect 407 -1780 410 -1774
rect 414 -1780 420 -1774
rect 421 -1780 424 -1774
rect 428 -1780 431 -1774
rect 435 -1780 438 -1774
rect 442 -1780 445 -1774
rect 449 -1780 452 -1774
rect 456 -1780 459 -1774
rect 463 -1780 466 -1774
rect 470 -1780 473 -1774
rect 477 -1780 483 -1774
rect 484 -1780 487 -1774
rect 491 -1780 494 -1774
rect 498 -1780 501 -1774
rect 505 -1780 508 -1774
rect 512 -1780 518 -1774
rect 519 -1780 525 -1774
rect 526 -1780 529 -1774
rect 533 -1780 536 -1774
rect 540 -1780 543 -1774
rect 547 -1780 550 -1774
rect 554 -1780 560 -1774
rect 561 -1780 567 -1774
rect 568 -1780 571 -1774
rect 575 -1780 578 -1774
rect 582 -1780 585 -1774
rect 589 -1780 592 -1774
rect 596 -1780 602 -1774
rect 603 -1780 606 -1774
rect 610 -1780 613 -1774
rect 617 -1780 620 -1774
rect 624 -1780 627 -1774
rect 631 -1780 634 -1774
rect 638 -1780 641 -1774
rect 645 -1780 651 -1774
rect 652 -1780 655 -1774
rect 659 -1780 662 -1774
rect 666 -1780 669 -1774
rect 673 -1780 676 -1774
rect 680 -1780 686 -1774
rect 687 -1780 690 -1774
rect 694 -1780 700 -1774
rect 701 -1780 704 -1774
rect 708 -1780 711 -1774
rect 715 -1780 718 -1774
rect 722 -1780 725 -1774
rect 729 -1780 732 -1774
rect 736 -1780 742 -1774
rect 743 -1780 746 -1774
rect 750 -1780 753 -1774
rect 757 -1780 760 -1774
rect 764 -1780 767 -1774
rect 771 -1780 774 -1774
rect 778 -1780 781 -1774
rect 785 -1780 788 -1774
rect 792 -1780 795 -1774
rect 799 -1780 802 -1774
rect 806 -1780 812 -1774
rect 813 -1780 816 -1774
rect 820 -1780 823 -1774
rect 827 -1780 833 -1774
rect 834 -1780 837 -1774
rect 841 -1780 844 -1774
rect 848 -1780 851 -1774
rect 855 -1780 858 -1774
rect 862 -1780 865 -1774
rect 869 -1780 872 -1774
rect 876 -1780 879 -1774
rect 883 -1780 889 -1774
rect 890 -1780 893 -1774
rect 897 -1780 903 -1774
rect 904 -1780 907 -1774
rect 911 -1780 914 -1774
rect 918 -1780 921 -1774
rect 925 -1780 928 -1774
rect 932 -1780 935 -1774
rect 939 -1780 945 -1774
rect 946 -1780 949 -1774
rect 953 -1780 956 -1774
rect 960 -1780 963 -1774
rect 967 -1780 970 -1774
rect 974 -1780 977 -1774
rect 981 -1780 987 -1774
rect 988 -1780 991 -1774
rect 995 -1780 998 -1774
rect 1002 -1780 1005 -1774
rect 1009 -1780 1012 -1774
rect 1016 -1780 1019 -1774
rect 1023 -1780 1026 -1774
rect 1030 -1780 1033 -1774
rect 1037 -1780 1040 -1774
rect 1044 -1780 1047 -1774
rect 1051 -1780 1054 -1774
rect 1058 -1780 1061 -1774
rect 1065 -1780 1068 -1774
rect 1072 -1780 1078 -1774
rect 1079 -1780 1085 -1774
rect 1086 -1780 1089 -1774
rect 1093 -1780 1096 -1774
rect 1100 -1780 1106 -1774
rect 1107 -1780 1113 -1774
rect 1114 -1780 1117 -1774
rect 1121 -1780 1124 -1774
rect 1128 -1780 1131 -1774
rect 1135 -1780 1138 -1774
rect 1142 -1780 1145 -1774
rect 1149 -1780 1152 -1774
rect 1156 -1780 1159 -1774
rect 1163 -1780 1166 -1774
rect 1170 -1780 1173 -1774
rect 1177 -1780 1180 -1774
rect 1184 -1780 1187 -1774
rect 1191 -1780 1194 -1774
rect 1198 -1780 1201 -1774
rect 1205 -1780 1208 -1774
rect 1212 -1780 1215 -1774
rect 1219 -1780 1222 -1774
rect 1226 -1780 1229 -1774
rect 1233 -1780 1236 -1774
rect 1240 -1780 1246 -1774
rect 1247 -1780 1250 -1774
rect 1254 -1780 1257 -1774
rect 1261 -1780 1264 -1774
rect 1268 -1780 1271 -1774
rect 1275 -1780 1278 -1774
rect 1282 -1780 1285 -1774
rect 1289 -1780 1292 -1774
rect 1296 -1780 1299 -1774
rect 1303 -1780 1309 -1774
rect 1310 -1780 1313 -1774
rect 1317 -1780 1323 -1774
rect 1324 -1780 1327 -1774
rect 1331 -1780 1334 -1774
rect 1338 -1780 1341 -1774
rect 1345 -1780 1348 -1774
rect 1352 -1780 1358 -1774
rect 1359 -1780 1365 -1774
rect 1366 -1780 1369 -1774
rect 1373 -1780 1376 -1774
rect 1380 -1780 1383 -1774
rect 1387 -1780 1390 -1774
rect 1394 -1780 1397 -1774
rect 1401 -1780 1404 -1774
rect 1408 -1780 1411 -1774
rect 1415 -1780 1418 -1774
rect 1422 -1780 1425 -1774
rect 1429 -1780 1432 -1774
rect 1436 -1780 1439 -1774
rect 1443 -1780 1446 -1774
rect 1450 -1780 1453 -1774
rect 1457 -1780 1460 -1774
rect 1464 -1780 1470 -1774
rect 1471 -1780 1474 -1774
rect 1478 -1780 1481 -1774
rect 1485 -1780 1488 -1774
rect 1492 -1780 1495 -1774
rect 1499 -1780 1502 -1774
rect 1506 -1780 1509 -1774
rect 1513 -1780 1516 -1774
rect 1520 -1780 1523 -1774
rect 1527 -1780 1530 -1774
rect 1534 -1780 1537 -1774
rect 1541 -1780 1544 -1774
rect 1548 -1780 1551 -1774
rect 1555 -1780 1558 -1774
rect 1562 -1780 1565 -1774
rect 1569 -1780 1572 -1774
rect 1576 -1780 1579 -1774
rect 1583 -1780 1586 -1774
rect 1590 -1780 1593 -1774
rect 1597 -1780 1600 -1774
rect 1604 -1780 1607 -1774
rect 1611 -1780 1614 -1774
rect 1618 -1780 1621 -1774
rect 1625 -1780 1628 -1774
rect 1632 -1780 1635 -1774
rect 1639 -1780 1642 -1774
rect 1646 -1780 1649 -1774
rect 1653 -1780 1656 -1774
rect 1660 -1780 1663 -1774
rect 1667 -1780 1670 -1774
rect 1674 -1780 1677 -1774
rect 1681 -1780 1684 -1774
rect 1688 -1780 1691 -1774
rect 1695 -1780 1698 -1774
rect 1702 -1780 1705 -1774
rect 1709 -1780 1712 -1774
rect 1716 -1780 1719 -1774
rect 1723 -1780 1726 -1774
rect 1730 -1780 1733 -1774
rect 1737 -1780 1740 -1774
rect 1744 -1780 1747 -1774
rect 1751 -1780 1754 -1774
rect 1758 -1780 1761 -1774
rect 1765 -1780 1768 -1774
rect 1772 -1780 1775 -1774
rect 1779 -1780 1782 -1774
rect 1786 -1780 1789 -1774
rect 1793 -1780 1796 -1774
rect 1800 -1780 1803 -1774
rect 1807 -1780 1810 -1774
rect 1814 -1780 1817 -1774
rect 1821 -1780 1824 -1774
rect 1828 -1780 1831 -1774
rect 1835 -1780 1838 -1774
rect 1842 -1780 1845 -1774
rect 1849 -1780 1852 -1774
rect 1856 -1780 1859 -1774
rect 1863 -1780 1866 -1774
rect 1870 -1780 1873 -1774
rect 1877 -1780 1880 -1774
rect 1884 -1780 1887 -1774
rect 1891 -1780 1894 -1774
rect 1898 -1780 1901 -1774
rect 1905 -1780 1908 -1774
rect 1912 -1780 1915 -1774
rect 1919 -1780 1922 -1774
rect 1926 -1780 1929 -1774
rect 1933 -1780 1939 -1774
rect 1940 -1780 1946 -1774
rect 1947 -1780 1950 -1774
rect 1954 -1780 1957 -1774
rect 1961 -1780 1964 -1774
rect 1968 -1780 1971 -1774
rect 2017 -1780 2020 -1774
rect 1 -1905 7 -1899
rect 8 -1905 14 -1899
rect 15 -1905 18 -1899
rect 22 -1905 25 -1899
rect 29 -1905 32 -1899
rect 36 -1905 39 -1899
rect 43 -1905 46 -1899
rect 50 -1905 53 -1899
rect 57 -1905 63 -1899
rect 64 -1905 67 -1899
rect 71 -1905 74 -1899
rect 78 -1905 81 -1899
rect 85 -1905 88 -1899
rect 92 -1905 95 -1899
rect 99 -1905 105 -1899
rect 106 -1905 109 -1899
rect 113 -1905 116 -1899
rect 120 -1905 123 -1899
rect 127 -1905 130 -1899
rect 134 -1905 140 -1899
rect 141 -1905 147 -1899
rect 148 -1905 151 -1899
rect 155 -1905 158 -1899
rect 162 -1905 165 -1899
rect 169 -1905 172 -1899
rect 176 -1905 179 -1899
rect 183 -1905 186 -1899
rect 190 -1905 193 -1899
rect 197 -1905 203 -1899
rect 204 -1905 207 -1899
rect 211 -1905 214 -1899
rect 218 -1905 221 -1899
rect 225 -1905 228 -1899
rect 232 -1905 235 -1899
rect 239 -1905 242 -1899
rect 246 -1905 249 -1899
rect 253 -1905 256 -1899
rect 260 -1905 263 -1899
rect 267 -1905 270 -1899
rect 274 -1905 277 -1899
rect 281 -1905 284 -1899
rect 288 -1905 291 -1899
rect 295 -1905 298 -1899
rect 302 -1905 305 -1899
rect 309 -1905 312 -1899
rect 316 -1905 319 -1899
rect 323 -1905 326 -1899
rect 330 -1905 333 -1899
rect 337 -1905 340 -1899
rect 344 -1905 347 -1899
rect 351 -1905 354 -1899
rect 358 -1905 361 -1899
rect 365 -1905 368 -1899
rect 372 -1905 375 -1899
rect 379 -1905 382 -1899
rect 386 -1905 389 -1899
rect 393 -1905 396 -1899
rect 400 -1905 406 -1899
rect 407 -1905 410 -1899
rect 414 -1905 417 -1899
rect 421 -1905 424 -1899
rect 428 -1905 431 -1899
rect 435 -1905 438 -1899
rect 442 -1905 445 -1899
rect 449 -1905 452 -1899
rect 456 -1905 459 -1899
rect 463 -1905 466 -1899
rect 470 -1905 473 -1899
rect 477 -1905 483 -1899
rect 484 -1905 490 -1899
rect 491 -1905 494 -1899
rect 498 -1905 501 -1899
rect 505 -1905 511 -1899
rect 512 -1905 515 -1899
rect 519 -1905 522 -1899
rect 526 -1905 529 -1899
rect 533 -1905 536 -1899
rect 540 -1905 543 -1899
rect 547 -1905 550 -1899
rect 554 -1905 557 -1899
rect 561 -1905 564 -1899
rect 568 -1905 571 -1899
rect 575 -1905 581 -1899
rect 582 -1905 585 -1899
rect 589 -1905 592 -1899
rect 596 -1905 599 -1899
rect 603 -1905 606 -1899
rect 610 -1905 616 -1899
rect 617 -1905 623 -1899
rect 624 -1905 627 -1899
rect 631 -1905 634 -1899
rect 638 -1905 641 -1899
rect 645 -1905 648 -1899
rect 652 -1905 655 -1899
rect 659 -1905 662 -1899
rect 666 -1905 669 -1899
rect 673 -1905 676 -1899
rect 680 -1905 683 -1899
rect 687 -1905 693 -1899
rect 694 -1905 697 -1899
rect 701 -1905 704 -1899
rect 708 -1905 711 -1899
rect 715 -1905 721 -1899
rect 722 -1905 728 -1899
rect 729 -1905 732 -1899
rect 736 -1905 739 -1899
rect 743 -1905 746 -1899
rect 750 -1905 753 -1899
rect 757 -1905 760 -1899
rect 764 -1905 770 -1899
rect 771 -1905 777 -1899
rect 778 -1905 781 -1899
rect 785 -1905 788 -1899
rect 792 -1905 795 -1899
rect 799 -1905 802 -1899
rect 806 -1905 809 -1899
rect 813 -1905 816 -1899
rect 820 -1905 823 -1899
rect 827 -1905 830 -1899
rect 834 -1905 837 -1899
rect 841 -1905 844 -1899
rect 848 -1905 851 -1899
rect 855 -1905 858 -1899
rect 862 -1905 865 -1899
rect 869 -1905 872 -1899
rect 876 -1905 879 -1899
rect 883 -1905 889 -1899
rect 890 -1905 893 -1899
rect 897 -1905 900 -1899
rect 904 -1905 910 -1899
rect 911 -1905 914 -1899
rect 918 -1905 921 -1899
rect 925 -1905 928 -1899
rect 932 -1905 938 -1899
rect 939 -1905 942 -1899
rect 946 -1905 949 -1899
rect 953 -1905 956 -1899
rect 960 -1905 963 -1899
rect 967 -1905 970 -1899
rect 974 -1905 977 -1899
rect 981 -1905 987 -1899
rect 988 -1905 991 -1899
rect 995 -1905 998 -1899
rect 1002 -1905 1005 -1899
rect 1009 -1905 1012 -1899
rect 1016 -1905 1019 -1899
rect 1023 -1905 1029 -1899
rect 1030 -1905 1033 -1899
rect 1037 -1905 1040 -1899
rect 1044 -1905 1047 -1899
rect 1051 -1905 1054 -1899
rect 1058 -1905 1064 -1899
rect 1065 -1905 1068 -1899
rect 1072 -1905 1075 -1899
rect 1079 -1905 1082 -1899
rect 1086 -1905 1092 -1899
rect 1093 -1905 1096 -1899
rect 1100 -1905 1106 -1899
rect 1107 -1905 1113 -1899
rect 1114 -1905 1117 -1899
rect 1121 -1905 1127 -1899
rect 1128 -1905 1131 -1899
rect 1135 -1905 1138 -1899
rect 1142 -1905 1145 -1899
rect 1149 -1905 1155 -1899
rect 1156 -1905 1159 -1899
rect 1163 -1905 1166 -1899
rect 1170 -1905 1173 -1899
rect 1177 -1905 1180 -1899
rect 1184 -1905 1187 -1899
rect 1191 -1905 1194 -1899
rect 1198 -1905 1201 -1899
rect 1205 -1905 1211 -1899
rect 1212 -1905 1215 -1899
rect 1219 -1905 1225 -1899
rect 1226 -1905 1229 -1899
rect 1233 -1905 1236 -1899
rect 1240 -1905 1243 -1899
rect 1247 -1905 1250 -1899
rect 1254 -1905 1257 -1899
rect 1261 -1905 1264 -1899
rect 1268 -1905 1271 -1899
rect 1275 -1905 1281 -1899
rect 1282 -1905 1285 -1899
rect 1289 -1905 1292 -1899
rect 1296 -1905 1299 -1899
rect 1303 -1905 1306 -1899
rect 1310 -1905 1313 -1899
rect 1317 -1905 1320 -1899
rect 1324 -1905 1327 -1899
rect 1331 -1905 1334 -1899
rect 1338 -1905 1341 -1899
rect 1345 -1905 1348 -1899
rect 1352 -1905 1355 -1899
rect 1359 -1905 1362 -1899
rect 1366 -1905 1369 -1899
rect 1373 -1905 1376 -1899
rect 1380 -1905 1383 -1899
rect 1387 -1905 1390 -1899
rect 1394 -1905 1397 -1899
rect 1401 -1905 1404 -1899
rect 1408 -1905 1411 -1899
rect 1415 -1905 1418 -1899
rect 1422 -1905 1425 -1899
rect 1429 -1905 1432 -1899
rect 1436 -1905 1439 -1899
rect 1443 -1905 1446 -1899
rect 1450 -1905 1453 -1899
rect 1457 -1905 1460 -1899
rect 1464 -1905 1467 -1899
rect 1471 -1905 1474 -1899
rect 1478 -1905 1481 -1899
rect 1485 -1905 1488 -1899
rect 1492 -1905 1495 -1899
rect 1499 -1905 1502 -1899
rect 1506 -1905 1509 -1899
rect 1513 -1905 1516 -1899
rect 1520 -1905 1523 -1899
rect 1527 -1905 1530 -1899
rect 1534 -1905 1537 -1899
rect 1541 -1905 1544 -1899
rect 1548 -1905 1551 -1899
rect 1555 -1905 1558 -1899
rect 1562 -1905 1568 -1899
rect 1569 -1905 1572 -1899
rect 1576 -1905 1579 -1899
rect 1583 -1905 1586 -1899
rect 1590 -1905 1593 -1899
rect 1597 -1905 1600 -1899
rect 1604 -1905 1607 -1899
rect 1611 -1905 1614 -1899
rect 1618 -1905 1621 -1899
rect 1625 -1905 1628 -1899
rect 1632 -1905 1635 -1899
rect 1639 -1905 1642 -1899
rect 1646 -1905 1649 -1899
rect 1653 -1905 1656 -1899
rect 1660 -1905 1663 -1899
rect 1667 -1905 1670 -1899
rect 1674 -1905 1677 -1899
rect 1681 -1905 1684 -1899
rect 1688 -1905 1691 -1899
rect 1695 -1905 1698 -1899
rect 1702 -1905 1705 -1899
rect 1709 -1905 1712 -1899
rect 1716 -1905 1719 -1899
rect 1723 -1905 1726 -1899
rect 1730 -1905 1733 -1899
rect 1737 -1905 1740 -1899
rect 1744 -1905 1747 -1899
rect 1751 -1905 1754 -1899
rect 1758 -1905 1761 -1899
rect 1765 -1905 1768 -1899
rect 1772 -1905 1775 -1899
rect 1779 -1905 1782 -1899
rect 1786 -1905 1789 -1899
rect 1793 -1905 1796 -1899
rect 1800 -1905 1803 -1899
rect 1807 -1905 1810 -1899
rect 1814 -1905 1817 -1899
rect 1821 -1905 1824 -1899
rect 1828 -1905 1831 -1899
rect 1835 -1905 1838 -1899
rect 1842 -1905 1845 -1899
rect 1849 -1905 1852 -1899
rect 1856 -1905 1859 -1899
rect 1863 -1905 1866 -1899
rect 1870 -1905 1873 -1899
rect 1877 -1905 1880 -1899
rect 1884 -1905 1887 -1899
rect 1891 -1905 1894 -1899
rect 1898 -1905 1901 -1899
rect 1905 -1905 1908 -1899
rect 1912 -1905 1915 -1899
rect 1919 -1905 1922 -1899
rect 1926 -1905 1929 -1899
rect 1933 -1905 1936 -1899
rect 1940 -1905 1943 -1899
rect 1947 -1905 1950 -1899
rect 1954 -1905 1957 -1899
rect 1961 -1905 1964 -1899
rect 1968 -1905 1971 -1899
rect 1975 -1905 1978 -1899
rect 1982 -1905 1985 -1899
rect 1989 -1905 1992 -1899
rect 1996 -1905 1999 -1899
rect 2003 -1905 2006 -1899
rect 2010 -1905 2016 -1899
rect 2017 -1905 2020 -1899
rect 2024 -1905 2027 -1899
rect 1 -2052 4 -2046
rect 8 -2052 11 -2046
rect 15 -2052 21 -2046
rect 22 -2052 25 -2046
rect 29 -2052 32 -2046
rect 36 -2052 39 -2046
rect 43 -2052 46 -2046
rect 50 -2052 53 -2046
rect 57 -2052 60 -2046
rect 64 -2052 70 -2046
rect 71 -2052 74 -2046
rect 78 -2052 81 -2046
rect 85 -2052 88 -2046
rect 92 -2052 95 -2046
rect 99 -2052 102 -2046
rect 106 -2052 109 -2046
rect 113 -2052 119 -2046
rect 120 -2052 123 -2046
rect 127 -2052 130 -2046
rect 134 -2052 137 -2046
rect 141 -2052 147 -2046
rect 148 -2052 151 -2046
rect 155 -2052 158 -2046
rect 162 -2052 165 -2046
rect 169 -2052 172 -2046
rect 176 -2052 179 -2046
rect 183 -2052 186 -2046
rect 190 -2052 193 -2046
rect 197 -2052 200 -2046
rect 204 -2052 207 -2046
rect 211 -2052 214 -2046
rect 218 -2052 224 -2046
rect 225 -2052 228 -2046
rect 232 -2052 235 -2046
rect 239 -2052 245 -2046
rect 246 -2052 249 -2046
rect 253 -2052 256 -2046
rect 260 -2052 263 -2046
rect 267 -2052 270 -2046
rect 274 -2052 277 -2046
rect 281 -2052 284 -2046
rect 288 -2052 291 -2046
rect 295 -2052 298 -2046
rect 302 -2052 305 -2046
rect 309 -2052 315 -2046
rect 316 -2052 319 -2046
rect 323 -2052 326 -2046
rect 330 -2052 333 -2046
rect 337 -2052 343 -2046
rect 344 -2052 347 -2046
rect 351 -2052 354 -2046
rect 358 -2052 361 -2046
rect 365 -2052 368 -2046
rect 372 -2052 375 -2046
rect 379 -2052 382 -2046
rect 386 -2052 389 -2046
rect 393 -2052 396 -2046
rect 400 -2052 403 -2046
rect 407 -2052 410 -2046
rect 414 -2052 417 -2046
rect 421 -2052 424 -2046
rect 428 -2052 431 -2046
rect 435 -2052 438 -2046
rect 442 -2052 445 -2046
rect 449 -2052 455 -2046
rect 456 -2052 459 -2046
rect 463 -2052 466 -2046
rect 470 -2052 473 -2046
rect 477 -2052 480 -2046
rect 484 -2052 487 -2046
rect 491 -2052 494 -2046
rect 498 -2052 501 -2046
rect 505 -2052 508 -2046
rect 512 -2052 515 -2046
rect 519 -2052 522 -2046
rect 526 -2052 532 -2046
rect 533 -2052 539 -2046
rect 540 -2052 543 -2046
rect 547 -2052 550 -2046
rect 554 -2052 557 -2046
rect 561 -2052 564 -2046
rect 568 -2052 571 -2046
rect 575 -2052 578 -2046
rect 582 -2052 585 -2046
rect 589 -2052 592 -2046
rect 596 -2052 599 -2046
rect 603 -2052 606 -2046
rect 610 -2052 613 -2046
rect 617 -2052 620 -2046
rect 624 -2052 627 -2046
rect 631 -2052 634 -2046
rect 638 -2052 641 -2046
rect 645 -2052 648 -2046
rect 652 -2052 655 -2046
rect 659 -2052 662 -2046
rect 666 -2052 669 -2046
rect 673 -2052 676 -2046
rect 680 -2052 683 -2046
rect 687 -2052 690 -2046
rect 694 -2052 700 -2046
rect 701 -2052 704 -2046
rect 708 -2052 711 -2046
rect 715 -2052 718 -2046
rect 722 -2052 728 -2046
rect 729 -2052 735 -2046
rect 736 -2052 739 -2046
rect 743 -2052 746 -2046
rect 750 -2052 756 -2046
rect 757 -2052 763 -2046
rect 764 -2052 767 -2046
rect 771 -2052 777 -2046
rect 778 -2052 781 -2046
rect 785 -2052 788 -2046
rect 792 -2052 795 -2046
rect 799 -2052 802 -2046
rect 806 -2052 809 -2046
rect 813 -2052 819 -2046
rect 820 -2052 823 -2046
rect 827 -2052 830 -2046
rect 834 -2052 837 -2046
rect 841 -2052 847 -2046
rect 848 -2052 854 -2046
rect 855 -2052 858 -2046
rect 862 -2052 868 -2046
rect 869 -2052 872 -2046
rect 876 -2052 882 -2046
rect 883 -2052 886 -2046
rect 890 -2052 896 -2046
rect 897 -2052 900 -2046
rect 904 -2052 907 -2046
rect 911 -2052 914 -2046
rect 918 -2052 924 -2046
rect 925 -2052 928 -2046
rect 932 -2052 935 -2046
rect 939 -2052 942 -2046
rect 946 -2052 949 -2046
rect 953 -2052 956 -2046
rect 960 -2052 966 -2046
rect 967 -2052 973 -2046
rect 974 -2052 977 -2046
rect 981 -2052 984 -2046
rect 988 -2052 991 -2046
rect 995 -2052 998 -2046
rect 1002 -2052 1005 -2046
rect 1009 -2052 1012 -2046
rect 1016 -2052 1019 -2046
rect 1023 -2052 1026 -2046
rect 1030 -2052 1033 -2046
rect 1037 -2052 1040 -2046
rect 1044 -2052 1047 -2046
rect 1051 -2052 1054 -2046
rect 1058 -2052 1061 -2046
rect 1065 -2052 1068 -2046
rect 1072 -2052 1075 -2046
rect 1079 -2052 1082 -2046
rect 1086 -2052 1092 -2046
rect 1093 -2052 1096 -2046
rect 1100 -2052 1103 -2046
rect 1107 -2052 1113 -2046
rect 1114 -2052 1117 -2046
rect 1121 -2052 1124 -2046
rect 1128 -2052 1131 -2046
rect 1135 -2052 1138 -2046
rect 1142 -2052 1145 -2046
rect 1149 -2052 1152 -2046
rect 1156 -2052 1159 -2046
rect 1163 -2052 1166 -2046
rect 1170 -2052 1173 -2046
rect 1177 -2052 1180 -2046
rect 1184 -2052 1187 -2046
rect 1191 -2052 1197 -2046
rect 1198 -2052 1201 -2046
rect 1205 -2052 1208 -2046
rect 1212 -2052 1215 -2046
rect 1219 -2052 1222 -2046
rect 1226 -2052 1229 -2046
rect 1233 -2052 1239 -2046
rect 1240 -2052 1243 -2046
rect 1247 -2052 1250 -2046
rect 1254 -2052 1260 -2046
rect 1261 -2052 1267 -2046
rect 1268 -2052 1271 -2046
rect 1275 -2052 1278 -2046
rect 1282 -2052 1285 -2046
rect 1289 -2052 1295 -2046
rect 1296 -2052 1299 -2046
rect 1303 -2052 1306 -2046
rect 1310 -2052 1313 -2046
rect 1317 -2052 1320 -2046
rect 1324 -2052 1327 -2046
rect 1331 -2052 1334 -2046
rect 1338 -2052 1341 -2046
rect 1345 -2052 1348 -2046
rect 1352 -2052 1355 -2046
rect 1359 -2052 1362 -2046
rect 1366 -2052 1369 -2046
rect 1373 -2052 1376 -2046
rect 1380 -2052 1383 -2046
rect 1387 -2052 1390 -2046
rect 1394 -2052 1397 -2046
rect 1401 -2052 1404 -2046
rect 1408 -2052 1411 -2046
rect 1415 -2052 1418 -2046
rect 1422 -2052 1425 -2046
rect 1429 -2052 1432 -2046
rect 1436 -2052 1439 -2046
rect 1443 -2052 1446 -2046
rect 1450 -2052 1456 -2046
rect 1457 -2052 1460 -2046
rect 1464 -2052 1467 -2046
rect 1471 -2052 1474 -2046
rect 1478 -2052 1481 -2046
rect 1485 -2052 1488 -2046
rect 1492 -2052 1495 -2046
rect 1499 -2052 1502 -2046
rect 1506 -2052 1509 -2046
rect 1513 -2052 1516 -2046
rect 1520 -2052 1523 -2046
rect 1527 -2052 1530 -2046
rect 1534 -2052 1537 -2046
rect 1541 -2052 1544 -2046
rect 1548 -2052 1551 -2046
rect 1555 -2052 1558 -2046
rect 1562 -2052 1565 -2046
rect 1569 -2052 1572 -2046
rect 1576 -2052 1579 -2046
rect 1583 -2052 1586 -2046
rect 1590 -2052 1593 -2046
rect 1597 -2052 1600 -2046
rect 1604 -2052 1607 -2046
rect 1611 -2052 1614 -2046
rect 1618 -2052 1621 -2046
rect 1625 -2052 1628 -2046
rect 1632 -2052 1635 -2046
rect 1639 -2052 1642 -2046
rect 1646 -2052 1649 -2046
rect 1653 -2052 1656 -2046
rect 1660 -2052 1663 -2046
rect 1667 -2052 1670 -2046
rect 1674 -2052 1677 -2046
rect 1681 -2052 1684 -2046
rect 1688 -2052 1691 -2046
rect 1695 -2052 1698 -2046
rect 1702 -2052 1705 -2046
rect 1709 -2052 1712 -2046
rect 1716 -2052 1719 -2046
rect 1723 -2052 1726 -2046
rect 1730 -2052 1733 -2046
rect 1737 -2052 1740 -2046
rect 1744 -2052 1747 -2046
rect 1751 -2052 1754 -2046
rect 1758 -2052 1761 -2046
rect 1765 -2052 1768 -2046
rect 1772 -2052 1775 -2046
rect 1779 -2052 1782 -2046
rect 1786 -2052 1789 -2046
rect 1793 -2052 1796 -2046
rect 1800 -2052 1803 -2046
rect 1807 -2052 1810 -2046
rect 1814 -2052 1817 -2046
rect 1821 -2052 1824 -2046
rect 1828 -2052 1831 -2046
rect 1835 -2052 1838 -2046
rect 1842 -2052 1845 -2046
rect 1849 -2052 1852 -2046
rect 1856 -2052 1859 -2046
rect 1863 -2052 1866 -2046
rect 1870 -2052 1873 -2046
rect 1877 -2052 1880 -2046
rect 1884 -2052 1887 -2046
rect 1891 -2052 1894 -2046
rect 1898 -2052 1901 -2046
rect 1905 -2052 1908 -2046
rect 1912 -2052 1915 -2046
rect 1919 -2052 1925 -2046
rect 1926 -2052 1929 -2046
rect 1933 -2052 1936 -2046
rect 1940 -2052 1943 -2046
rect 1947 -2052 1950 -2046
rect 1954 -2052 1957 -2046
rect 1961 -2052 1964 -2046
rect 1968 -2052 1971 -2046
rect 1975 -2052 1978 -2046
rect 1982 -2052 1985 -2046
rect 1989 -2052 1992 -2046
rect 1 -2193 4 -2187
rect 8 -2193 14 -2187
rect 15 -2193 18 -2187
rect 22 -2193 25 -2187
rect 29 -2193 35 -2187
rect 36 -2193 42 -2187
rect 43 -2193 46 -2187
rect 50 -2193 53 -2187
rect 57 -2193 60 -2187
rect 64 -2193 67 -2187
rect 71 -2193 74 -2187
rect 78 -2193 81 -2187
rect 85 -2193 91 -2187
rect 92 -2193 98 -2187
rect 99 -2193 102 -2187
rect 106 -2193 112 -2187
rect 113 -2193 119 -2187
rect 120 -2193 123 -2187
rect 127 -2193 130 -2187
rect 134 -2193 137 -2187
rect 141 -2193 144 -2187
rect 148 -2193 151 -2187
rect 155 -2193 158 -2187
rect 162 -2193 165 -2187
rect 169 -2193 172 -2187
rect 176 -2193 179 -2187
rect 183 -2193 186 -2187
rect 190 -2193 193 -2187
rect 197 -2193 200 -2187
rect 204 -2193 207 -2187
rect 211 -2193 214 -2187
rect 218 -2193 221 -2187
rect 225 -2193 228 -2187
rect 232 -2193 238 -2187
rect 239 -2193 242 -2187
rect 246 -2193 249 -2187
rect 253 -2193 256 -2187
rect 260 -2193 263 -2187
rect 267 -2193 270 -2187
rect 274 -2193 277 -2187
rect 281 -2193 284 -2187
rect 288 -2193 291 -2187
rect 295 -2193 298 -2187
rect 302 -2193 305 -2187
rect 309 -2193 312 -2187
rect 316 -2193 319 -2187
rect 323 -2193 326 -2187
rect 330 -2193 333 -2187
rect 337 -2193 343 -2187
rect 344 -2193 347 -2187
rect 351 -2193 354 -2187
rect 358 -2193 361 -2187
rect 365 -2193 368 -2187
rect 372 -2193 375 -2187
rect 379 -2193 382 -2187
rect 386 -2193 392 -2187
rect 393 -2193 396 -2187
rect 400 -2193 406 -2187
rect 407 -2193 410 -2187
rect 414 -2193 417 -2187
rect 421 -2193 424 -2187
rect 428 -2193 431 -2187
rect 435 -2193 441 -2187
rect 442 -2193 445 -2187
rect 449 -2193 452 -2187
rect 456 -2193 459 -2187
rect 463 -2193 469 -2187
rect 470 -2193 473 -2187
rect 477 -2193 480 -2187
rect 484 -2193 487 -2187
rect 491 -2193 494 -2187
rect 498 -2193 501 -2187
rect 505 -2193 511 -2187
rect 512 -2193 515 -2187
rect 519 -2193 522 -2187
rect 526 -2193 529 -2187
rect 533 -2193 536 -2187
rect 540 -2193 546 -2187
rect 547 -2193 550 -2187
rect 554 -2193 557 -2187
rect 561 -2193 564 -2187
rect 568 -2193 571 -2187
rect 575 -2193 578 -2187
rect 582 -2193 585 -2187
rect 589 -2193 595 -2187
rect 596 -2193 599 -2187
rect 603 -2193 606 -2187
rect 610 -2193 613 -2187
rect 617 -2193 620 -2187
rect 624 -2193 630 -2187
rect 631 -2193 634 -2187
rect 638 -2193 641 -2187
rect 645 -2193 651 -2187
rect 652 -2193 655 -2187
rect 659 -2193 662 -2187
rect 666 -2193 669 -2187
rect 673 -2193 676 -2187
rect 680 -2193 683 -2187
rect 687 -2193 690 -2187
rect 694 -2193 697 -2187
rect 701 -2193 704 -2187
rect 708 -2193 711 -2187
rect 715 -2193 718 -2187
rect 722 -2193 725 -2187
rect 729 -2193 732 -2187
rect 736 -2193 739 -2187
rect 743 -2193 746 -2187
rect 750 -2193 753 -2187
rect 757 -2193 760 -2187
rect 764 -2193 767 -2187
rect 771 -2193 774 -2187
rect 778 -2193 781 -2187
rect 785 -2193 788 -2187
rect 792 -2193 795 -2187
rect 799 -2193 802 -2187
rect 806 -2193 809 -2187
rect 813 -2193 816 -2187
rect 820 -2193 823 -2187
rect 827 -2193 830 -2187
rect 834 -2193 840 -2187
rect 841 -2193 844 -2187
rect 848 -2193 851 -2187
rect 855 -2193 858 -2187
rect 862 -2193 865 -2187
rect 869 -2193 872 -2187
rect 876 -2193 882 -2187
rect 883 -2193 886 -2187
rect 890 -2193 893 -2187
rect 897 -2193 900 -2187
rect 904 -2193 907 -2187
rect 911 -2193 914 -2187
rect 918 -2193 921 -2187
rect 925 -2193 928 -2187
rect 932 -2193 935 -2187
rect 939 -2193 942 -2187
rect 946 -2193 949 -2187
rect 953 -2193 956 -2187
rect 960 -2193 963 -2187
rect 967 -2193 973 -2187
rect 974 -2193 980 -2187
rect 981 -2193 984 -2187
rect 988 -2193 991 -2187
rect 995 -2193 998 -2187
rect 1002 -2193 1005 -2187
rect 1009 -2193 1012 -2187
rect 1016 -2193 1019 -2187
rect 1023 -2193 1026 -2187
rect 1030 -2193 1033 -2187
rect 1037 -2193 1040 -2187
rect 1044 -2193 1047 -2187
rect 1051 -2193 1057 -2187
rect 1058 -2193 1061 -2187
rect 1065 -2193 1071 -2187
rect 1072 -2193 1075 -2187
rect 1079 -2193 1085 -2187
rect 1086 -2193 1089 -2187
rect 1093 -2193 1096 -2187
rect 1100 -2193 1103 -2187
rect 1107 -2193 1113 -2187
rect 1114 -2193 1117 -2187
rect 1121 -2193 1124 -2187
rect 1128 -2193 1131 -2187
rect 1135 -2193 1141 -2187
rect 1142 -2193 1145 -2187
rect 1149 -2193 1152 -2187
rect 1156 -2193 1162 -2187
rect 1163 -2193 1166 -2187
rect 1170 -2193 1173 -2187
rect 1177 -2193 1180 -2187
rect 1184 -2193 1187 -2187
rect 1191 -2193 1194 -2187
rect 1198 -2193 1201 -2187
rect 1205 -2193 1208 -2187
rect 1212 -2193 1215 -2187
rect 1219 -2193 1222 -2187
rect 1226 -2193 1229 -2187
rect 1233 -2193 1236 -2187
rect 1240 -2193 1243 -2187
rect 1247 -2193 1250 -2187
rect 1254 -2193 1257 -2187
rect 1261 -2193 1264 -2187
rect 1268 -2193 1271 -2187
rect 1275 -2193 1281 -2187
rect 1282 -2193 1285 -2187
rect 1289 -2193 1292 -2187
rect 1296 -2193 1299 -2187
rect 1303 -2193 1306 -2187
rect 1310 -2193 1313 -2187
rect 1317 -2193 1320 -2187
rect 1324 -2193 1327 -2187
rect 1331 -2193 1334 -2187
rect 1338 -2193 1341 -2187
rect 1345 -2193 1348 -2187
rect 1352 -2193 1355 -2187
rect 1359 -2193 1365 -2187
rect 1366 -2193 1369 -2187
rect 1373 -2193 1379 -2187
rect 1380 -2193 1383 -2187
rect 1387 -2193 1390 -2187
rect 1394 -2193 1400 -2187
rect 1401 -2193 1407 -2187
rect 1408 -2193 1411 -2187
rect 1415 -2193 1418 -2187
rect 1422 -2193 1425 -2187
rect 1429 -2193 1432 -2187
rect 1436 -2193 1439 -2187
rect 1443 -2193 1446 -2187
rect 1450 -2193 1456 -2187
rect 1457 -2193 1460 -2187
rect 1464 -2193 1467 -2187
rect 1471 -2193 1477 -2187
rect 1478 -2193 1481 -2187
rect 1485 -2193 1488 -2187
rect 1492 -2193 1495 -2187
rect 1499 -2193 1502 -2187
rect 1506 -2193 1509 -2187
rect 1513 -2193 1516 -2187
rect 1520 -2193 1523 -2187
rect 1527 -2193 1530 -2187
rect 1534 -2193 1537 -2187
rect 1541 -2193 1544 -2187
rect 1548 -2193 1551 -2187
rect 1555 -2193 1558 -2187
rect 1562 -2193 1565 -2187
rect 1569 -2193 1572 -2187
rect 1576 -2193 1579 -2187
rect 1583 -2193 1586 -2187
rect 1590 -2193 1593 -2187
rect 1597 -2193 1600 -2187
rect 1604 -2193 1607 -2187
rect 1611 -2193 1614 -2187
rect 1618 -2193 1621 -2187
rect 1625 -2193 1628 -2187
rect 1632 -2193 1635 -2187
rect 1639 -2193 1642 -2187
rect 1646 -2193 1649 -2187
rect 1653 -2193 1656 -2187
rect 1660 -2193 1663 -2187
rect 1667 -2193 1670 -2187
rect 1674 -2193 1677 -2187
rect 1681 -2193 1684 -2187
rect 1688 -2193 1691 -2187
rect 1695 -2193 1698 -2187
rect 1702 -2193 1705 -2187
rect 1709 -2193 1712 -2187
rect 1716 -2193 1719 -2187
rect 1723 -2193 1726 -2187
rect 1730 -2193 1733 -2187
rect 1737 -2193 1740 -2187
rect 1744 -2193 1747 -2187
rect 1751 -2193 1754 -2187
rect 1758 -2193 1761 -2187
rect 1765 -2193 1768 -2187
rect 1772 -2193 1775 -2187
rect 1779 -2193 1782 -2187
rect 1786 -2193 1789 -2187
rect 1793 -2193 1796 -2187
rect 1800 -2193 1803 -2187
rect 1807 -2193 1810 -2187
rect 1814 -2193 1817 -2187
rect 1821 -2193 1824 -2187
rect 1828 -2193 1831 -2187
rect 1835 -2193 1838 -2187
rect 1842 -2193 1845 -2187
rect 1849 -2193 1852 -2187
rect 1856 -2193 1859 -2187
rect 1863 -2193 1866 -2187
rect 1870 -2193 1873 -2187
rect 1877 -2193 1880 -2187
rect 1884 -2193 1887 -2187
rect 1891 -2193 1894 -2187
rect 1898 -2193 1901 -2187
rect 1905 -2193 1908 -2187
rect 1912 -2193 1915 -2187
rect 1 -2322 7 -2316
rect 8 -2322 11 -2316
rect 15 -2322 21 -2316
rect 22 -2322 25 -2316
rect 29 -2322 32 -2316
rect 36 -2322 39 -2316
rect 43 -2322 46 -2316
rect 50 -2322 53 -2316
rect 57 -2322 60 -2316
rect 64 -2322 70 -2316
rect 71 -2322 74 -2316
rect 78 -2322 81 -2316
rect 85 -2322 88 -2316
rect 92 -2322 95 -2316
rect 99 -2322 102 -2316
rect 106 -2322 109 -2316
rect 113 -2322 119 -2316
rect 120 -2322 126 -2316
rect 127 -2322 130 -2316
rect 134 -2322 137 -2316
rect 141 -2322 144 -2316
rect 148 -2322 151 -2316
rect 155 -2322 161 -2316
rect 162 -2322 165 -2316
rect 169 -2322 175 -2316
rect 176 -2322 179 -2316
rect 183 -2322 186 -2316
rect 190 -2322 193 -2316
rect 197 -2322 200 -2316
rect 204 -2322 210 -2316
rect 211 -2322 217 -2316
rect 218 -2322 224 -2316
rect 225 -2322 228 -2316
rect 232 -2322 238 -2316
rect 239 -2322 245 -2316
rect 246 -2322 249 -2316
rect 253 -2322 256 -2316
rect 260 -2322 263 -2316
rect 267 -2322 270 -2316
rect 274 -2322 277 -2316
rect 281 -2322 284 -2316
rect 288 -2322 291 -2316
rect 295 -2322 298 -2316
rect 302 -2322 305 -2316
rect 309 -2322 312 -2316
rect 316 -2322 319 -2316
rect 323 -2322 326 -2316
rect 330 -2322 333 -2316
rect 337 -2322 340 -2316
rect 344 -2322 347 -2316
rect 351 -2322 354 -2316
rect 358 -2322 361 -2316
rect 365 -2322 368 -2316
rect 372 -2322 375 -2316
rect 379 -2322 382 -2316
rect 386 -2322 389 -2316
rect 393 -2322 396 -2316
rect 400 -2322 403 -2316
rect 407 -2322 410 -2316
rect 414 -2322 417 -2316
rect 421 -2322 424 -2316
rect 428 -2322 431 -2316
rect 435 -2322 438 -2316
rect 442 -2322 445 -2316
rect 449 -2322 452 -2316
rect 456 -2322 459 -2316
rect 463 -2322 469 -2316
rect 470 -2322 473 -2316
rect 477 -2322 480 -2316
rect 484 -2322 487 -2316
rect 491 -2322 494 -2316
rect 498 -2322 501 -2316
rect 505 -2322 508 -2316
rect 512 -2322 515 -2316
rect 519 -2322 522 -2316
rect 526 -2322 529 -2316
rect 533 -2322 536 -2316
rect 540 -2322 543 -2316
rect 547 -2322 550 -2316
rect 554 -2322 557 -2316
rect 561 -2322 564 -2316
rect 568 -2322 574 -2316
rect 575 -2322 578 -2316
rect 582 -2322 585 -2316
rect 589 -2322 592 -2316
rect 596 -2322 599 -2316
rect 603 -2322 606 -2316
rect 610 -2322 613 -2316
rect 617 -2322 620 -2316
rect 624 -2322 630 -2316
rect 631 -2322 634 -2316
rect 638 -2322 641 -2316
rect 645 -2322 648 -2316
rect 652 -2322 658 -2316
rect 659 -2322 662 -2316
rect 666 -2322 672 -2316
rect 673 -2322 679 -2316
rect 680 -2322 683 -2316
rect 687 -2322 690 -2316
rect 694 -2322 697 -2316
rect 701 -2322 704 -2316
rect 708 -2322 711 -2316
rect 715 -2322 718 -2316
rect 722 -2322 725 -2316
rect 729 -2322 732 -2316
rect 736 -2322 739 -2316
rect 743 -2322 746 -2316
rect 750 -2322 753 -2316
rect 757 -2322 763 -2316
rect 764 -2322 767 -2316
rect 771 -2322 774 -2316
rect 778 -2322 781 -2316
rect 785 -2322 788 -2316
rect 792 -2322 798 -2316
rect 799 -2322 802 -2316
rect 806 -2322 809 -2316
rect 813 -2322 819 -2316
rect 820 -2322 826 -2316
rect 827 -2322 830 -2316
rect 834 -2322 837 -2316
rect 841 -2322 844 -2316
rect 848 -2322 851 -2316
rect 855 -2322 858 -2316
rect 862 -2322 865 -2316
rect 869 -2322 872 -2316
rect 876 -2322 879 -2316
rect 883 -2322 889 -2316
rect 890 -2322 893 -2316
rect 897 -2322 900 -2316
rect 904 -2322 907 -2316
rect 911 -2322 914 -2316
rect 918 -2322 921 -2316
rect 925 -2322 928 -2316
rect 932 -2322 935 -2316
rect 939 -2322 942 -2316
rect 946 -2322 952 -2316
rect 953 -2322 956 -2316
rect 960 -2322 963 -2316
rect 967 -2322 970 -2316
rect 974 -2322 977 -2316
rect 981 -2322 984 -2316
rect 988 -2322 991 -2316
rect 995 -2322 1001 -2316
rect 1002 -2322 1005 -2316
rect 1009 -2322 1012 -2316
rect 1016 -2322 1019 -2316
rect 1023 -2322 1026 -2316
rect 1030 -2322 1033 -2316
rect 1037 -2322 1040 -2316
rect 1044 -2322 1047 -2316
rect 1051 -2322 1054 -2316
rect 1058 -2322 1061 -2316
rect 1065 -2322 1071 -2316
rect 1072 -2322 1075 -2316
rect 1079 -2322 1082 -2316
rect 1086 -2322 1089 -2316
rect 1093 -2322 1096 -2316
rect 1100 -2322 1103 -2316
rect 1107 -2322 1110 -2316
rect 1114 -2322 1120 -2316
rect 1121 -2322 1127 -2316
rect 1128 -2322 1131 -2316
rect 1135 -2322 1138 -2316
rect 1142 -2322 1145 -2316
rect 1149 -2322 1152 -2316
rect 1156 -2322 1159 -2316
rect 1163 -2322 1166 -2316
rect 1170 -2322 1173 -2316
rect 1177 -2322 1180 -2316
rect 1184 -2322 1190 -2316
rect 1191 -2322 1194 -2316
rect 1198 -2322 1201 -2316
rect 1205 -2322 1208 -2316
rect 1212 -2322 1215 -2316
rect 1219 -2322 1222 -2316
rect 1226 -2322 1229 -2316
rect 1233 -2322 1236 -2316
rect 1240 -2322 1243 -2316
rect 1247 -2322 1250 -2316
rect 1254 -2322 1257 -2316
rect 1261 -2322 1264 -2316
rect 1268 -2322 1271 -2316
rect 1275 -2322 1278 -2316
rect 1282 -2322 1285 -2316
rect 1289 -2322 1295 -2316
rect 1296 -2322 1299 -2316
rect 1303 -2322 1309 -2316
rect 1310 -2322 1313 -2316
rect 1317 -2322 1320 -2316
rect 1324 -2322 1327 -2316
rect 1331 -2322 1334 -2316
rect 1338 -2322 1341 -2316
rect 1345 -2322 1348 -2316
rect 1352 -2322 1355 -2316
rect 1359 -2322 1362 -2316
rect 1366 -2322 1372 -2316
rect 1373 -2322 1376 -2316
rect 1380 -2322 1383 -2316
rect 1387 -2322 1390 -2316
rect 1394 -2322 1397 -2316
rect 1401 -2322 1404 -2316
rect 1408 -2322 1411 -2316
rect 1415 -2322 1418 -2316
rect 1422 -2322 1425 -2316
rect 1429 -2322 1432 -2316
rect 1436 -2322 1439 -2316
rect 1443 -2322 1446 -2316
rect 1450 -2322 1453 -2316
rect 1457 -2322 1460 -2316
rect 1464 -2322 1467 -2316
rect 1471 -2322 1474 -2316
rect 1478 -2322 1481 -2316
rect 1485 -2322 1488 -2316
rect 1492 -2322 1495 -2316
rect 1499 -2322 1502 -2316
rect 1506 -2322 1509 -2316
rect 1513 -2322 1516 -2316
rect 1520 -2322 1523 -2316
rect 1527 -2322 1530 -2316
rect 1534 -2322 1537 -2316
rect 1541 -2322 1544 -2316
rect 1548 -2322 1551 -2316
rect 1555 -2322 1558 -2316
rect 1562 -2322 1565 -2316
rect 1569 -2322 1572 -2316
rect 1576 -2322 1579 -2316
rect 1583 -2322 1586 -2316
rect 1590 -2322 1593 -2316
rect 1597 -2322 1600 -2316
rect 1604 -2322 1607 -2316
rect 1611 -2322 1614 -2316
rect 1618 -2322 1621 -2316
rect 1625 -2322 1628 -2316
rect 1632 -2322 1635 -2316
rect 1639 -2322 1642 -2316
rect 1646 -2322 1649 -2316
rect 1653 -2322 1656 -2316
rect 1660 -2322 1663 -2316
rect 1667 -2322 1670 -2316
rect 1674 -2322 1677 -2316
rect 1681 -2322 1684 -2316
rect 1688 -2322 1691 -2316
rect 1695 -2322 1698 -2316
rect 1702 -2322 1705 -2316
rect 1709 -2322 1715 -2316
rect 1716 -2322 1719 -2316
rect 1723 -2322 1729 -2316
rect 1730 -2322 1733 -2316
rect 1737 -2322 1740 -2316
rect 1744 -2322 1750 -2316
rect 1751 -2322 1754 -2316
rect 1758 -2322 1761 -2316
rect 1765 -2322 1768 -2316
rect 1772 -2322 1775 -2316
rect 1779 -2322 1782 -2316
rect 1786 -2322 1789 -2316
rect 1793 -2322 1796 -2316
rect 1821 -2322 1824 -2316
rect 1828 -2322 1831 -2316
rect 1 -2447 7 -2441
rect 8 -2447 11 -2441
rect 15 -2447 18 -2441
rect 22 -2447 28 -2441
rect 29 -2447 32 -2441
rect 36 -2447 39 -2441
rect 43 -2447 46 -2441
rect 50 -2447 53 -2441
rect 57 -2447 60 -2441
rect 64 -2447 67 -2441
rect 71 -2447 74 -2441
rect 78 -2447 84 -2441
rect 85 -2447 88 -2441
rect 92 -2447 98 -2441
rect 99 -2447 102 -2441
rect 106 -2447 112 -2441
rect 113 -2447 116 -2441
rect 120 -2447 123 -2441
rect 127 -2447 133 -2441
rect 134 -2447 137 -2441
rect 141 -2447 144 -2441
rect 148 -2447 151 -2441
rect 155 -2447 158 -2441
rect 162 -2447 165 -2441
rect 169 -2447 172 -2441
rect 176 -2447 179 -2441
rect 183 -2447 186 -2441
rect 190 -2447 196 -2441
rect 197 -2447 200 -2441
rect 204 -2447 207 -2441
rect 211 -2447 214 -2441
rect 218 -2447 221 -2441
rect 225 -2447 228 -2441
rect 232 -2447 235 -2441
rect 239 -2447 242 -2441
rect 246 -2447 249 -2441
rect 253 -2447 256 -2441
rect 260 -2447 263 -2441
rect 267 -2447 270 -2441
rect 274 -2447 277 -2441
rect 281 -2447 284 -2441
rect 288 -2447 291 -2441
rect 295 -2447 298 -2441
rect 302 -2447 305 -2441
rect 309 -2447 312 -2441
rect 316 -2447 319 -2441
rect 323 -2447 326 -2441
rect 330 -2447 333 -2441
rect 337 -2447 343 -2441
rect 344 -2447 347 -2441
rect 351 -2447 354 -2441
rect 358 -2447 361 -2441
rect 365 -2447 368 -2441
rect 372 -2447 375 -2441
rect 379 -2447 382 -2441
rect 386 -2447 392 -2441
rect 393 -2447 396 -2441
rect 400 -2447 406 -2441
rect 407 -2447 410 -2441
rect 414 -2447 417 -2441
rect 421 -2447 424 -2441
rect 428 -2447 434 -2441
rect 435 -2447 441 -2441
rect 442 -2447 448 -2441
rect 449 -2447 452 -2441
rect 456 -2447 462 -2441
rect 463 -2447 466 -2441
rect 470 -2447 473 -2441
rect 477 -2447 480 -2441
rect 484 -2447 487 -2441
rect 491 -2447 494 -2441
rect 498 -2447 501 -2441
rect 505 -2447 508 -2441
rect 512 -2447 518 -2441
rect 519 -2447 522 -2441
rect 526 -2447 532 -2441
rect 533 -2447 536 -2441
rect 540 -2447 546 -2441
rect 547 -2447 550 -2441
rect 554 -2447 557 -2441
rect 561 -2447 564 -2441
rect 568 -2447 571 -2441
rect 575 -2447 578 -2441
rect 582 -2447 585 -2441
rect 589 -2447 592 -2441
rect 596 -2447 602 -2441
rect 603 -2447 606 -2441
rect 610 -2447 613 -2441
rect 617 -2447 620 -2441
rect 624 -2447 627 -2441
rect 631 -2447 634 -2441
rect 638 -2447 641 -2441
rect 645 -2447 648 -2441
rect 652 -2447 655 -2441
rect 659 -2447 662 -2441
rect 666 -2447 669 -2441
rect 673 -2447 679 -2441
rect 680 -2447 683 -2441
rect 687 -2447 690 -2441
rect 694 -2447 700 -2441
rect 701 -2447 704 -2441
rect 708 -2447 711 -2441
rect 715 -2447 721 -2441
rect 722 -2447 725 -2441
rect 729 -2447 735 -2441
rect 736 -2447 739 -2441
rect 743 -2447 746 -2441
rect 750 -2447 753 -2441
rect 757 -2447 760 -2441
rect 764 -2447 767 -2441
rect 771 -2447 774 -2441
rect 778 -2447 781 -2441
rect 785 -2447 791 -2441
rect 792 -2447 795 -2441
rect 799 -2447 802 -2441
rect 806 -2447 809 -2441
rect 813 -2447 816 -2441
rect 820 -2447 823 -2441
rect 827 -2447 833 -2441
rect 834 -2447 837 -2441
rect 841 -2447 844 -2441
rect 848 -2447 851 -2441
rect 855 -2447 858 -2441
rect 862 -2447 865 -2441
rect 869 -2447 872 -2441
rect 876 -2447 879 -2441
rect 883 -2447 889 -2441
rect 890 -2447 893 -2441
rect 897 -2447 900 -2441
rect 904 -2447 907 -2441
rect 911 -2447 914 -2441
rect 918 -2447 921 -2441
rect 925 -2447 928 -2441
rect 932 -2447 935 -2441
rect 939 -2447 942 -2441
rect 946 -2447 949 -2441
rect 953 -2447 956 -2441
rect 960 -2447 963 -2441
rect 967 -2447 970 -2441
rect 974 -2447 977 -2441
rect 981 -2447 984 -2441
rect 988 -2447 991 -2441
rect 995 -2447 998 -2441
rect 1002 -2447 1005 -2441
rect 1009 -2447 1012 -2441
rect 1016 -2447 1022 -2441
rect 1023 -2447 1026 -2441
rect 1030 -2447 1033 -2441
rect 1037 -2447 1040 -2441
rect 1044 -2447 1047 -2441
rect 1051 -2447 1057 -2441
rect 1058 -2447 1061 -2441
rect 1065 -2447 1068 -2441
rect 1072 -2447 1075 -2441
rect 1079 -2447 1085 -2441
rect 1086 -2447 1089 -2441
rect 1093 -2447 1096 -2441
rect 1100 -2447 1103 -2441
rect 1107 -2447 1110 -2441
rect 1114 -2447 1117 -2441
rect 1121 -2447 1124 -2441
rect 1128 -2447 1131 -2441
rect 1135 -2447 1138 -2441
rect 1142 -2447 1145 -2441
rect 1149 -2447 1152 -2441
rect 1156 -2447 1159 -2441
rect 1163 -2447 1169 -2441
rect 1170 -2447 1173 -2441
rect 1177 -2447 1180 -2441
rect 1184 -2447 1187 -2441
rect 1191 -2447 1194 -2441
rect 1198 -2447 1201 -2441
rect 1205 -2447 1208 -2441
rect 1212 -2447 1218 -2441
rect 1219 -2447 1222 -2441
rect 1226 -2447 1229 -2441
rect 1233 -2447 1236 -2441
rect 1240 -2447 1243 -2441
rect 1247 -2447 1250 -2441
rect 1254 -2447 1257 -2441
rect 1261 -2447 1264 -2441
rect 1268 -2447 1271 -2441
rect 1275 -2447 1278 -2441
rect 1282 -2447 1285 -2441
rect 1289 -2447 1292 -2441
rect 1296 -2447 1299 -2441
rect 1303 -2447 1306 -2441
rect 1310 -2447 1313 -2441
rect 1317 -2447 1323 -2441
rect 1324 -2447 1327 -2441
rect 1331 -2447 1334 -2441
rect 1338 -2447 1344 -2441
rect 1345 -2447 1348 -2441
rect 1352 -2447 1355 -2441
rect 1359 -2447 1362 -2441
rect 1366 -2447 1369 -2441
rect 1373 -2447 1376 -2441
rect 1380 -2447 1383 -2441
rect 1387 -2447 1393 -2441
rect 1394 -2447 1397 -2441
rect 1401 -2447 1404 -2441
rect 1408 -2447 1411 -2441
rect 1415 -2447 1418 -2441
rect 1422 -2447 1425 -2441
rect 1429 -2447 1432 -2441
rect 1436 -2447 1439 -2441
rect 1443 -2447 1446 -2441
rect 1450 -2447 1453 -2441
rect 1457 -2447 1460 -2441
rect 1464 -2447 1467 -2441
rect 1471 -2447 1474 -2441
rect 1478 -2447 1481 -2441
rect 1485 -2447 1488 -2441
rect 1492 -2447 1495 -2441
rect 1499 -2447 1502 -2441
rect 1506 -2447 1509 -2441
rect 1513 -2447 1516 -2441
rect 1520 -2447 1523 -2441
rect 1527 -2447 1530 -2441
rect 1534 -2447 1537 -2441
rect 1541 -2447 1544 -2441
rect 1548 -2447 1551 -2441
rect 1555 -2447 1558 -2441
rect 1562 -2447 1565 -2441
rect 1569 -2447 1572 -2441
rect 1576 -2447 1579 -2441
rect 1583 -2447 1586 -2441
rect 1590 -2447 1593 -2441
rect 1597 -2447 1600 -2441
rect 1604 -2447 1607 -2441
rect 1611 -2447 1614 -2441
rect 1618 -2447 1621 -2441
rect 1625 -2447 1628 -2441
rect 1632 -2447 1635 -2441
rect 1639 -2447 1642 -2441
rect 1646 -2447 1649 -2441
rect 1653 -2447 1656 -2441
rect 1660 -2447 1663 -2441
rect 1667 -2447 1670 -2441
rect 1674 -2447 1677 -2441
rect 1681 -2447 1684 -2441
rect 1688 -2447 1691 -2441
rect 1695 -2447 1698 -2441
rect 1702 -2447 1705 -2441
rect 1709 -2447 1712 -2441
rect 1716 -2447 1719 -2441
rect 1723 -2447 1726 -2441
rect 1730 -2447 1733 -2441
rect 1737 -2447 1740 -2441
rect 1744 -2447 1747 -2441
rect 1751 -2447 1757 -2441
rect 1758 -2447 1761 -2441
rect 1765 -2447 1768 -2441
rect 1772 -2447 1775 -2441
rect 1779 -2447 1782 -2441
rect 1786 -2447 1789 -2441
rect 1793 -2447 1799 -2441
rect 1800 -2447 1803 -2441
rect 1807 -2447 1810 -2441
rect 1 -2582 7 -2576
rect 8 -2582 14 -2576
rect 15 -2582 18 -2576
rect 22 -2582 25 -2576
rect 29 -2582 32 -2576
rect 36 -2582 39 -2576
rect 43 -2582 46 -2576
rect 50 -2582 53 -2576
rect 57 -2582 60 -2576
rect 64 -2582 67 -2576
rect 71 -2582 74 -2576
rect 78 -2582 81 -2576
rect 85 -2582 88 -2576
rect 92 -2582 95 -2576
rect 99 -2582 105 -2576
rect 106 -2582 112 -2576
rect 113 -2582 116 -2576
rect 120 -2582 123 -2576
rect 127 -2582 130 -2576
rect 134 -2582 137 -2576
rect 141 -2582 144 -2576
rect 148 -2582 154 -2576
rect 155 -2582 161 -2576
rect 162 -2582 165 -2576
rect 169 -2582 175 -2576
rect 176 -2582 179 -2576
rect 183 -2582 186 -2576
rect 190 -2582 193 -2576
rect 197 -2582 200 -2576
rect 204 -2582 207 -2576
rect 211 -2582 214 -2576
rect 218 -2582 221 -2576
rect 225 -2582 228 -2576
rect 232 -2582 235 -2576
rect 239 -2582 245 -2576
rect 246 -2582 249 -2576
rect 253 -2582 256 -2576
rect 260 -2582 263 -2576
rect 267 -2582 270 -2576
rect 274 -2582 277 -2576
rect 281 -2582 284 -2576
rect 288 -2582 291 -2576
rect 295 -2582 298 -2576
rect 302 -2582 305 -2576
rect 309 -2582 312 -2576
rect 316 -2582 319 -2576
rect 323 -2582 326 -2576
rect 330 -2582 333 -2576
rect 337 -2582 340 -2576
rect 344 -2582 347 -2576
rect 351 -2582 354 -2576
rect 358 -2582 361 -2576
rect 365 -2582 368 -2576
rect 372 -2582 375 -2576
rect 379 -2582 382 -2576
rect 386 -2582 389 -2576
rect 393 -2582 396 -2576
rect 400 -2582 403 -2576
rect 407 -2582 410 -2576
rect 414 -2582 417 -2576
rect 421 -2582 424 -2576
rect 428 -2582 431 -2576
rect 435 -2582 438 -2576
rect 442 -2582 445 -2576
rect 449 -2582 455 -2576
rect 456 -2582 459 -2576
rect 463 -2582 466 -2576
rect 470 -2582 473 -2576
rect 477 -2582 480 -2576
rect 484 -2582 487 -2576
rect 491 -2582 494 -2576
rect 498 -2582 501 -2576
rect 505 -2582 508 -2576
rect 512 -2582 515 -2576
rect 519 -2582 522 -2576
rect 526 -2582 529 -2576
rect 533 -2582 536 -2576
rect 540 -2582 543 -2576
rect 547 -2582 550 -2576
rect 554 -2582 560 -2576
rect 561 -2582 564 -2576
rect 568 -2582 571 -2576
rect 575 -2582 578 -2576
rect 582 -2582 585 -2576
rect 589 -2582 592 -2576
rect 596 -2582 602 -2576
rect 603 -2582 606 -2576
rect 610 -2582 613 -2576
rect 617 -2582 620 -2576
rect 624 -2582 630 -2576
rect 631 -2582 634 -2576
rect 638 -2582 644 -2576
rect 645 -2582 648 -2576
rect 652 -2582 655 -2576
rect 659 -2582 662 -2576
rect 666 -2582 672 -2576
rect 673 -2582 676 -2576
rect 680 -2582 683 -2576
rect 687 -2582 690 -2576
rect 694 -2582 697 -2576
rect 701 -2582 704 -2576
rect 708 -2582 714 -2576
rect 715 -2582 718 -2576
rect 722 -2582 728 -2576
rect 729 -2582 732 -2576
rect 736 -2582 742 -2576
rect 743 -2582 746 -2576
rect 750 -2582 753 -2576
rect 757 -2582 760 -2576
rect 764 -2582 767 -2576
rect 771 -2582 774 -2576
rect 778 -2582 781 -2576
rect 785 -2582 788 -2576
rect 792 -2582 795 -2576
rect 799 -2582 802 -2576
rect 806 -2582 809 -2576
rect 813 -2582 816 -2576
rect 820 -2582 823 -2576
rect 827 -2582 830 -2576
rect 834 -2582 837 -2576
rect 841 -2582 844 -2576
rect 848 -2582 854 -2576
rect 855 -2582 858 -2576
rect 862 -2582 865 -2576
rect 869 -2582 872 -2576
rect 876 -2582 879 -2576
rect 883 -2582 886 -2576
rect 890 -2582 893 -2576
rect 897 -2582 900 -2576
rect 904 -2582 907 -2576
rect 911 -2582 914 -2576
rect 918 -2582 921 -2576
rect 925 -2582 928 -2576
rect 932 -2582 935 -2576
rect 939 -2582 942 -2576
rect 946 -2582 952 -2576
rect 953 -2582 956 -2576
rect 960 -2582 963 -2576
rect 967 -2582 973 -2576
rect 974 -2582 977 -2576
rect 981 -2582 984 -2576
rect 988 -2582 994 -2576
rect 995 -2582 998 -2576
rect 1002 -2582 1005 -2576
rect 1009 -2582 1012 -2576
rect 1016 -2582 1022 -2576
rect 1023 -2582 1026 -2576
rect 1030 -2582 1033 -2576
rect 1037 -2582 1040 -2576
rect 1044 -2582 1050 -2576
rect 1051 -2582 1057 -2576
rect 1058 -2582 1061 -2576
rect 1065 -2582 1068 -2576
rect 1072 -2582 1078 -2576
rect 1079 -2582 1082 -2576
rect 1086 -2582 1089 -2576
rect 1093 -2582 1096 -2576
rect 1100 -2582 1103 -2576
rect 1107 -2582 1110 -2576
rect 1114 -2582 1120 -2576
rect 1121 -2582 1124 -2576
rect 1128 -2582 1134 -2576
rect 1135 -2582 1141 -2576
rect 1142 -2582 1145 -2576
rect 1149 -2582 1152 -2576
rect 1156 -2582 1162 -2576
rect 1163 -2582 1166 -2576
rect 1170 -2582 1176 -2576
rect 1177 -2582 1180 -2576
rect 1184 -2582 1187 -2576
rect 1191 -2582 1197 -2576
rect 1198 -2582 1201 -2576
rect 1205 -2582 1208 -2576
rect 1212 -2582 1215 -2576
rect 1219 -2582 1222 -2576
rect 1226 -2582 1229 -2576
rect 1233 -2582 1236 -2576
rect 1240 -2582 1243 -2576
rect 1247 -2582 1250 -2576
rect 1254 -2582 1257 -2576
rect 1261 -2582 1264 -2576
rect 1268 -2582 1271 -2576
rect 1275 -2582 1278 -2576
rect 1282 -2582 1285 -2576
rect 1289 -2582 1292 -2576
rect 1296 -2582 1299 -2576
rect 1303 -2582 1306 -2576
rect 1310 -2582 1313 -2576
rect 1317 -2582 1320 -2576
rect 1324 -2582 1327 -2576
rect 1331 -2582 1334 -2576
rect 1338 -2582 1341 -2576
rect 1345 -2582 1348 -2576
rect 1352 -2582 1355 -2576
rect 1359 -2582 1362 -2576
rect 1366 -2582 1369 -2576
rect 1373 -2582 1376 -2576
rect 1380 -2582 1383 -2576
rect 1387 -2582 1390 -2576
rect 1394 -2582 1397 -2576
rect 1401 -2582 1404 -2576
rect 1408 -2582 1411 -2576
rect 1415 -2582 1418 -2576
rect 1422 -2582 1425 -2576
rect 1429 -2582 1432 -2576
rect 1436 -2582 1439 -2576
rect 1443 -2582 1446 -2576
rect 1450 -2582 1453 -2576
rect 1457 -2582 1460 -2576
rect 1464 -2582 1467 -2576
rect 1471 -2582 1474 -2576
rect 1478 -2582 1481 -2576
rect 1485 -2582 1488 -2576
rect 1492 -2582 1495 -2576
rect 1499 -2582 1502 -2576
rect 1506 -2582 1512 -2576
rect 1513 -2582 1516 -2576
rect 1520 -2582 1523 -2576
rect 1527 -2582 1530 -2576
rect 1534 -2582 1537 -2576
rect 1541 -2582 1544 -2576
rect 1548 -2582 1551 -2576
rect 1555 -2582 1558 -2576
rect 1562 -2582 1565 -2576
rect 1569 -2582 1572 -2576
rect 1576 -2582 1579 -2576
rect 1583 -2582 1586 -2576
rect 1590 -2582 1593 -2576
rect 1597 -2582 1600 -2576
rect 1604 -2582 1607 -2576
rect 1611 -2582 1614 -2576
rect 1618 -2582 1621 -2576
rect 1625 -2582 1628 -2576
rect 1632 -2582 1635 -2576
rect 1639 -2582 1642 -2576
rect 1646 -2582 1649 -2576
rect 1653 -2582 1656 -2576
rect 1660 -2582 1663 -2576
rect 1667 -2582 1670 -2576
rect 1674 -2582 1677 -2576
rect 1681 -2582 1684 -2576
rect 1688 -2582 1691 -2576
rect 1695 -2582 1701 -2576
rect 1702 -2582 1705 -2576
rect 1709 -2582 1712 -2576
rect 1716 -2582 1719 -2576
rect 1723 -2582 1726 -2576
rect 1730 -2582 1733 -2576
rect 1737 -2582 1743 -2576
rect 1744 -2582 1747 -2576
rect 1751 -2582 1754 -2576
rect 1758 -2582 1761 -2576
rect 1765 -2582 1768 -2576
rect 1772 -2582 1775 -2576
rect 1779 -2582 1782 -2576
rect 1786 -2582 1789 -2576
rect 1793 -2582 1799 -2576
rect 1800 -2582 1803 -2576
rect 1807 -2582 1810 -2576
rect 1814 -2582 1817 -2576
rect 1 -2715 7 -2709
rect 8 -2715 11 -2709
rect 15 -2715 21 -2709
rect 22 -2715 28 -2709
rect 29 -2715 32 -2709
rect 36 -2715 39 -2709
rect 43 -2715 46 -2709
rect 50 -2715 53 -2709
rect 57 -2715 63 -2709
rect 64 -2715 70 -2709
rect 71 -2715 74 -2709
rect 78 -2715 81 -2709
rect 85 -2715 88 -2709
rect 92 -2715 95 -2709
rect 99 -2715 102 -2709
rect 106 -2715 109 -2709
rect 113 -2715 116 -2709
rect 120 -2715 123 -2709
rect 127 -2715 130 -2709
rect 134 -2715 137 -2709
rect 141 -2715 144 -2709
rect 148 -2715 151 -2709
rect 155 -2715 158 -2709
rect 162 -2715 165 -2709
rect 169 -2715 172 -2709
rect 176 -2715 179 -2709
rect 183 -2715 186 -2709
rect 190 -2715 193 -2709
rect 197 -2715 203 -2709
rect 204 -2715 210 -2709
rect 211 -2715 214 -2709
rect 218 -2715 221 -2709
rect 225 -2715 228 -2709
rect 232 -2715 235 -2709
rect 239 -2715 242 -2709
rect 246 -2715 249 -2709
rect 253 -2715 256 -2709
rect 260 -2715 263 -2709
rect 267 -2715 270 -2709
rect 274 -2715 277 -2709
rect 281 -2715 284 -2709
rect 288 -2715 294 -2709
rect 295 -2715 298 -2709
rect 302 -2715 305 -2709
rect 309 -2715 312 -2709
rect 316 -2715 319 -2709
rect 323 -2715 326 -2709
rect 330 -2715 333 -2709
rect 337 -2715 340 -2709
rect 344 -2715 347 -2709
rect 351 -2715 354 -2709
rect 358 -2715 361 -2709
rect 365 -2715 368 -2709
rect 372 -2715 375 -2709
rect 379 -2715 382 -2709
rect 386 -2715 389 -2709
rect 393 -2715 396 -2709
rect 400 -2715 403 -2709
rect 407 -2715 410 -2709
rect 414 -2715 417 -2709
rect 421 -2715 427 -2709
rect 428 -2715 431 -2709
rect 435 -2715 438 -2709
rect 442 -2715 445 -2709
rect 449 -2715 452 -2709
rect 456 -2715 459 -2709
rect 463 -2715 466 -2709
rect 470 -2715 473 -2709
rect 477 -2715 480 -2709
rect 484 -2715 487 -2709
rect 491 -2715 494 -2709
rect 498 -2715 501 -2709
rect 505 -2715 508 -2709
rect 512 -2715 515 -2709
rect 519 -2715 525 -2709
rect 526 -2715 529 -2709
rect 533 -2715 536 -2709
rect 540 -2715 543 -2709
rect 547 -2715 550 -2709
rect 554 -2715 557 -2709
rect 561 -2715 564 -2709
rect 568 -2715 571 -2709
rect 575 -2715 578 -2709
rect 582 -2715 588 -2709
rect 589 -2715 592 -2709
rect 596 -2715 599 -2709
rect 603 -2715 609 -2709
rect 610 -2715 613 -2709
rect 617 -2715 620 -2709
rect 624 -2715 627 -2709
rect 631 -2715 637 -2709
rect 638 -2715 644 -2709
rect 645 -2715 648 -2709
rect 652 -2715 655 -2709
rect 659 -2715 662 -2709
rect 666 -2715 669 -2709
rect 673 -2715 676 -2709
rect 680 -2715 683 -2709
rect 687 -2715 690 -2709
rect 694 -2715 697 -2709
rect 701 -2715 704 -2709
rect 708 -2715 714 -2709
rect 715 -2715 718 -2709
rect 722 -2715 725 -2709
rect 729 -2715 732 -2709
rect 736 -2715 739 -2709
rect 743 -2715 746 -2709
rect 750 -2715 753 -2709
rect 757 -2715 760 -2709
rect 764 -2715 767 -2709
rect 771 -2715 777 -2709
rect 778 -2715 781 -2709
rect 785 -2715 788 -2709
rect 792 -2715 795 -2709
rect 799 -2715 802 -2709
rect 806 -2715 809 -2709
rect 813 -2715 816 -2709
rect 820 -2715 823 -2709
rect 827 -2715 830 -2709
rect 834 -2715 837 -2709
rect 841 -2715 847 -2709
rect 848 -2715 854 -2709
rect 855 -2715 858 -2709
rect 862 -2715 868 -2709
rect 869 -2715 872 -2709
rect 876 -2715 879 -2709
rect 883 -2715 889 -2709
rect 890 -2715 893 -2709
rect 897 -2715 900 -2709
rect 904 -2715 907 -2709
rect 911 -2715 917 -2709
rect 918 -2715 924 -2709
rect 925 -2715 928 -2709
rect 932 -2715 935 -2709
rect 939 -2715 942 -2709
rect 946 -2715 949 -2709
rect 953 -2715 956 -2709
rect 960 -2715 963 -2709
rect 967 -2715 970 -2709
rect 974 -2715 980 -2709
rect 981 -2715 984 -2709
rect 988 -2715 991 -2709
rect 995 -2715 998 -2709
rect 1002 -2715 1005 -2709
rect 1009 -2715 1012 -2709
rect 1016 -2715 1022 -2709
rect 1023 -2715 1026 -2709
rect 1030 -2715 1033 -2709
rect 1037 -2715 1040 -2709
rect 1044 -2715 1047 -2709
rect 1051 -2715 1057 -2709
rect 1058 -2715 1064 -2709
rect 1065 -2715 1068 -2709
rect 1072 -2715 1075 -2709
rect 1079 -2715 1082 -2709
rect 1086 -2715 1089 -2709
rect 1093 -2715 1096 -2709
rect 1100 -2715 1103 -2709
rect 1107 -2715 1110 -2709
rect 1114 -2715 1117 -2709
rect 1121 -2715 1124 -2709
rect 1128 -2715 1131 -2709
rect 1135 -2715 1138 -2709
rect 1142 -2715 1145 -2709
rect 1149 -2715 1155 -2709
rect 1156 -2715 1159 -2709
rect 1163 -2715 1166 -2709
rect 1170 -2715 1173 -2709
rect 1177 -2715 1180 -2709
rect 1184 -2715 1187 -2709
rect 1191 -2715 1197 -2709
rect 1198 -2715 1201 -2709
rect 1205 -2715 1208 -2709
rect 1212 -2715 1215 -2709
rect 1219 -2715 1222 -2709
rect 1226 -2715 1229 -2709
rect 1233 -2715 1236 -2709
rect 1240 -2715 1246 -2709
rect 1247 -2715 1250 -2709
rect 1254 -2715 1257 -2709
rect 1261 -2715 1264 -2709
rect 1268 -2715 1271 -2709
rect 1275 -2715 1278 -2709
rect 1282 -2715 1285 -2709
rect 1289 -2715 1295 -2709
rect 1296 -2715 1299 -2709
rect 1303 -2715 1306 -2709
rect 1310 -2715 1313 -2709
rect 1317 -2715 1323 -2709
rect 1324 -2715 1330 -2709
rect 1331 -2715 1334 -2709
rect 1338 -2715 1341 -2709
rect 1345 -2715 1348 -2709
rect 1352 -2715 1355 -2709
rect 1359 -2715 1362 -2709
rect 1366 -2715 1369 -2709
rect 1373 -2715 1376 -2709
rect 1380 -2715 1383 -2709
rect 1387 -2715 1390 -2709
rect 1394 -2715 1397 -2709
rect 1401 -2715 1404 -2709
rect 1408 -2715 1411 -2709
rect 1415 -2715 1418 -2709
rect 1422 -2715 1425 -2709
rect 1429 -2715 1432 -2709
rect 1436 -2715 1439 -2709
rect 1443 -2715 1446 -2709
rect 1450 -2715 1453 -2709
rect 1457 -2715 1460 -2709
rect 1464 -2715 1467 -2709
rect 1471 -2715 1474 -2709
rect 1478 -2715 1481 -2709
rect 1485 -2715 1488 -2709
rect 1492 -2715 1495 -2709
rect 1499 -2715 1502 -2709
rect 1506 -2715 1509 -2709
rect 1513 -2715 1516 -2709
rect 1520 -2715 1523 -2709
rect 1527 -2715 1530 -2709
rect 1534 -2715 1537 -2709
rect 1541 -2715 1544 -2709
rect 1548 -2715 1551 -2709
rect 1555 -2715 1558 -2709
rect 1562 -2715 1565 -2709
rect 1569 -2715 1572 -2709
rect 1576 -2715 1579 -2709
rect 1583 -2715 1586 -2709
rect 1590 -2715 1593 -2709
rect 1597 -2715 1600 -2709
rect 1604 -2715 1607 -2709
rect 1611 -2715 1614 -2709
rect 1618 -2715 1621 -2709
rect 1625 -2715 1628 -2709
rect 1632 -2715 1635 -2709
rect 1639 -2715 1642 -2709
rect 1646 -2715 1649 -2709
rect 1653 -2715 1656 -2709
rect 1660 -2715 1663 -2709
rect 1667 -2715 1670 -2709
rect 1674 -2715 1677 -2709
rect 1681 -2715 1684 -2709
rect 1688 -2715 1691 -2709
rect 1695 -2715 1698 -2709
rect 1702 -2715 1705 -2709
rect 1709 -2715 1712 -2709
rect 1716 -2715 1719 -2709
rect 1723 -2715 1726 -2709
rect 1730 -2715 1733 -2709
rect 1737 -2715 1740 -2709
rect 1744 -2715 1747 -2709
rect 1751 -2715 1754 -2709
rect 1758 -2715 1761 -2709
rect 1765 -2715 1771 -2709
rect 1772 -2715 1778 -2709
rect 1779 -2715 1785 -2709
rect 1786 -2715 1789 -2709
rect 1793 -2715 1796 -2709
rect 1800 -2715 1803 -2709
rect 1807 -2715 1810 -2709
rect 1 -2836 7 -2830
rect 8 -2836 14 -2830
rect 15 -2836 21 -2830
rect 36 -2836 39 -2830
rect 43 -2836 46 -2830
rect 50 -2836 53 -2830
rect 57 -2836 60 -2830
rect 64 -2836 67 -2830
rect 71 -2836 74 -2830
rect 78 -2836 81 -2830
rect 85 -2836 88 -2830
rect 92 -2836 98 -2830
rect 99 -2836 102 -2830
rect 106 -2836 109 -2830
rect 113 -2836 116 -2830
rect 120 -2836 123 -2830
rect 127 -2836 130 -2830
rect 134 -2836 137 -2830
rect 141 -2836 144 -2830
rect 148 -2836 151 -2830
rect 155 -2836 158 -2830
rect 162 -2836 165 -2830
rect 169 -2836 172 -2830
rect 176 -2836 179 -2830
rect 183 -2836 186 -2830
rect 190 -2836 193 -2830
rect 197 -2836 200 -2830
rect 204 -2836 207 -2830
rect 211 -2836 214 -2830
rect 218 -2836 221 -2830
rect 225 -2836 228 -2830
rect 232 -2836 235 -2830
rect 239 -2836 242 -2830
rect 246 -2836 249 -2830
rect 253 -2836 256 -2830
rect 260 -2836 263 -2830
rect 267 -2836 270 -2830
rect 274 -2836 277 -2830
rect 281 -2836 284 -2830
rect 288 -2836 291 -2830
rect 295 -2836 298 -2830
rect 302 -2836 305 -2830
rect 309 -2836 312 -2830
rect 316 -2836 319 -2830
rect 323 -2836 326 -2830
rect 330 -2836 333 -2830
rect 337 -2836 340 -2830
rect 344 -2836 347 -2830
rect 351 -2836 357 -2830
rect 358 -2836 361 -2830
rect 365 -2836 368 -2830
rect 372 -2836 375 -2830
rect 379 -2836 382 -2830
rect 386 -2836 389 -2830
rect 393 -2836 396 -2830
rect 400 -2836 403 -2830
rect 407 -2836 410 -2830
rect 414 -2836 417 -2830
rect 421 -2836 424 -2830
rect 428 -2836 431 -2830
rect 435 -2836 438 -2830
rect 442 -2836 445 -2830
rect 449 -2836 452 -2830
rect 456 -2836 459 -2830
rect 463 -2836 466 -2830
rect 470 -2836 473 -2830
rect 477 -2836 483 -2830
rect 484 -2836 487 -2830
rect 491 -2836 494 -2830
rect 498 -2836 501 -2830
rect 505 -2836 508 -2830
rect 512 -2836 515 -2830
rect 519 -2836 522 -2830
rect 526 -2836 529 -2830
rect 533 -2836 536 -2830
rect 540 -2836 543 -2830
rect 547 -2836 550 -2830
rect 554 -2836 560 -2830
rect 561 -2836 567 -2830
rect 568 -2836 571 -2830
rect 575 -2836 578 -2830
rect 582 -2836 588 -2830
rect 589 -2836 592 -2830
rect 596 -2836 599 -2830
rect 603 -2836 606 -2830
rect 610 -2836 613 -2830
rect 617 -2836 623 -2830
rect 624 -2836 627 -2830
rect 631 -2836 634 -2830
rect 638 -2836 641 -2830
rect 645 -2836 648 -2830
rect 652 -2836 655 -2830
rect 659 -2836 665 -2830
rect 666 -2836 669 -2830
rect 673 -2836 676 -2830
rect 680 -2836 683 -2830
rect 687 -2836 690 -2830
rect 694 -2836 697 -2830
rect 701 -2836 707 -2830
rect 708 -2836 714 -2830
rect 715 -2836 718 -2830
rect 722 -2836 725 -2830
rect 729 -2836 735 -2830
rect 736 -2836 739 -2830
rect 743 -2836 746 -2830
rect 750 -2836 753 -2830
rect 757 -2836 760 -2830
rect 764 -2836 767 -2830
rect 771 -2836 774 -2830
rect 778 -2836 781 -2830
rect 785 -2836 788 -2830
rect 792 -2836 795 -2830
rect 799 -2836 802 -2830
rect 806 -2836 809 -2830
rect 813 -2836 816 -2830
rect 820 -2836 823 -2830
rect 827 -2836 833 -2830
rect 834 -2836 837 -2830
rect 841 -2836 844 -2830
rect 848 -2836 854 -2830
rect 855 -2836 861 -2830
rect 862 -2836 865 -2830
rect 869 -2836 875 -2830
rect 876 -2836 879 -2830
rect 883 -2836 886 -2830
rect 890 -2836 893 -2830
rect 897 -2836 900 -2830
rect 904 -2836 907 -2830
rect 911 -2836 914 -2830
rect 918 -2836 921 -2830
rect 925 -2836 928 -2830
rect 932 -2836 935 -2830
rect 939 -2836 942 -2830
rect 946 -2836 949 -2830
rect 953 -2836 956 -2830
rect 960 -2836 963 -2830
rect 967 -2836 970 -2830
rect 974 -2836 977 -2830
rect 981 -2836 984 -2830
rect 988 -2836 991 -2830
rect 995 -2836 1001 -2830
rect 1002 -2836 1005 -2830
rect 1009 -2836 1015 -2830
rect 1016 -2836 1022 -2830
rect 1023 -2836 1026 -2830
rect 1030 -2836 1033 -2830
rect 1037 -2836 1040 -2830
rect 1044 -2836 1047 -2830
rect 1051 -2836 1054 -2830
rect 1058 -2836 1061 -2830
rect 1065 -2836 1071 -2830
rect 1072 -2836 1075 -2830
rect 1079 -2836 1082 -2830
rect 1086 -2836 1089 -2830
rect 1093 -2836 1096 -2830
rect 1100 -2836 1103 -2830
rect 1107 -2836 1110 -2830
rect 1114 -2836 1120 -2830
rect 1121 -2836 1127 -2830
rect 1128 -2836 1134 -2830
rect 1135 -2836 1138 -2830
rect 1142 -2836 1145 -2830
rect 1149 -2836 1152 -2830
rect 1156 -2836 1159 -2830
rect 1163 -2836 1166 -2830
rect 1170 -2836 1173 -2830
rect 1177 -2836 1183 -2830
rect 1184 -2836 1187 -2830
rect 1191 -2836 1194 -2830
rect 1198 -2836 1204 -2830
rect 1205 -2836 1208 -2830
rect 1212 -2836 1215 -2830
rect 1219 -2836 1222 -2830
rect 1226 -2836 1229 -2830
rect 1233 -2836 1239 -2830
rect 1240 -2836 1243 -2830
rect 1247 -2836 1250 -2830
rect 1254 -2836 1257 -2830
rect 1261 -2836 1264 -2830
rect 1268 -2836 1271 -2830
rect 1275 -2836 1278 -2830
rect 1282 -2836 1288 -2830
rect 1289 -2836 1292 -2830
rect 1296 -2836 1299 -2830
rect 1303 -2836 1306 -2830
rect 1310 -2836 1313 -2830
rect 1317 -2836 1320 -2830
rect 1324 -2836 1327 -2830
rect 1331 -2836 1334 -2830
rect 1338 -2836 1344 -2830
rect 1345 -2836 1348 -2830
rect 1352 -2836 1358 -2830
rect 1359 -2836 1362 -2830
rect 1366 -2836 1369 -2830
rect 1373 -2836 1376 -2830
rect 1380 -2836 1383 -2830
rect 1387 -2836 1390 -2830
rect 1394 -2836 1397 -2830
rect 1401 -2836 1404 -2830
rect 1408 -2836 1411 -2830
rect 1415 -2836 1418 -2830
rect 1422 -2836 1425 -2830
rect 1429 -2836 1435 -2830
rect 1436 -2836 1439 -2830
rect 1443 -2836 1446 -2830
rect 1450 -2836 1453 -2830
rect 1457 -2836 1460 -2830
rect 1464 -2836 1467 -2830
rect 1471 -2836 1474 -2830
rect 1478 -2836 1481 -2830
rect 1485 -2836 1488 -2830
rect 1492 -2836 1495 -2830
rect 1499 -2836 1502 -2830
rect 1506 -2836 1509 -2830
rect 1513 -2836 1516 -2830
rect 1520 -2836 1523 -2830
rect 1527 -2836 1530 -2830
rect 1534 -2836 1537 -2830
rect 1541 -2836 1544 -2830
rect 1548 -2836 1551 -2830
rect 1555 -2836 1558 -2830
rect 1562 -2836 1565 -2830
rect 1569 -2836 1572 -2830
rect 1576 -2836 1579 -2830
rect 1583 -2836 1586 -2830
rect 1590 -2836 1593 -2830
rect 1597 -2836 1600 -2830
rect 1604 -2836 1607 -2830
rect 1611 -2836 1614 -2830
rect 1618 -2836 1621 -2830
rect 1625 -2836 1628 -2830
rect 1632 -2836 1635 -2830
rect 1639 -2836 1642 -2830
rect 1646 -2836 1649 -2830
rect 1653 -2836 1656 -2830
rect 1660 -2836 1663 -2830
rect 1667 -2836 1670 -2830
rect 1674 -2836 1677 -2830
rect 1681 -2836 1684 -2830
rect 1688 -2836 1691 -2830
rect 1695 -2836 1698 -2830
rect 1702 -2836 1705 -2830
rect 1709 -2836 1715 -2830
rect 1716 -2836 1722 -2830
rect 1723 -2836 1729 -2830
rect 1730 -2836 1733 -2830
rect 1737 -2836 1740 -2830
rect 1744 -2836 1747 -2830
rect 1751 -2836 1754 -2830
rect 1758 -2836 1761 -2830
rect 1765 -2836 1768 -2830
rect 1772 -2836 1775 -2830
rect 1 -2955 7 -2949
rect 8 -2955 14 -2949
rect 15 -2955 21 -2949
rect 22 -2955 25 -2949
rect 29 -2955 35 -2949
rect 36 -2955 42 -2949
rect 43 -2955 49 -2949
rect 50 -2955 53 -2949
rect 57 -2955 60 -2949
rect 64 -2955 67 -2949
rect 71 -2955 74 -2949
rect 78 -2955 84 -2949
rect 85 -2955 88 -2949
rect 92 -2955 95 -2949
rect 99 -2955 102 -2949
rect 106 -2955 112 -2949
rect 113 -2955 116 -2949
rect 120 -2955 123 -2949
rect 127 -2955 130 -2949
rect 134 -2955 140 -2949
rect 141 -2955 147 -2949
rect 148 -2955 151 -2949
rect 155 -2955 158 -2949
rect 162 -2955 168 -2949
rect 169 -2955 172 -2949
rect 176 -2955 179 -2949
rect 183 -2955 186 -2949
rect 190 -2955 193 -2949
rect 197 -2955 200 -2949
rect 204 -2955 210 -2949
rect 211 -2955 214 -2949
rect 218 -2955 224 -2949
rect 225 -2955 231 -2949
rect 232 -2955 235 -2949
rect 239 -2955 242 -2949
rect 246 -2955 249 -2949
rect 253 -2955 256 -2949
rect 260 -2955 263 -2949
rect 267 -2955 270 -2949
rect 274 -2955 277 -2949
rect 281 -2955 284 -2949
rect 288 -2955 291 -2949
rect 295 -2955 298 -2949
rect 302 -2955 305 -2949
rect 309 -2955 312 -2949
rect 316 -2955 319 -2949
rect 323 -2955 326 -2949
rect 330 -2955 333 -2949
rect 337 -2955 340 -2949
rect 344 -2955 347 -2949
rect 351 -2955 354 -2949
rect 358 -2955 361 -2949
rect 365 -2955 368 -2949
rect 372 -2955 375 -2949
rect 379 -2955 382 -2949
rect 386 -2955 389 -2949
rect 393 -2955 396 -2949
rect 400 -2955 403 -2949
rect 407 -2955 413 -2949
rect 414 -2955 417 -2949
rect 421 -2955 424 -2949
rect 428 -2955 431 -2949
rect 435 -2955 441 -2949
rect 442 -2955 445 -2949
rect 449 -2955 452 -2949
rect 456 -2955 459 -2949
rect 463 -2955 469 -2949
rect 470 -2955 473 -2949
rect 477 -2955 480 -2949
rect 484 -2955 487 -2949
rect 491 -2955 494 -2949
rect 498 -2955 501 -2949
rect 505 -2955 508 -2949
rect 512 -2955 515 -2949
rect 519 -2955 522 -2949
rect 526 -2955 529 -2949
rect 533 -2955 539 -2949
rect 540 -2955 543 -2949
rect 547 -2955 550 -2949
rect 554 -2955 557 -2949
rect 561 -2955 564 -2949
rect 568 -2955 571 -2949
rect 575 -2955 578 -2949
rect 582 -2955 585 -2949
rect 589 -2955 592 -2949
rect 596 -2955 599 -2949
rect 603 -2955 606 -2949
rect 610 -2955 613 -2949
rect 617 -2955 620 -2949
rect 624 -2955 627 -2949
rect 631 -2955 634 -2949
rect 638 -2955 641 -2949
rect 645 -2955 648 -2949
rect 652 -2955 658 -2949
rect 659 -2955 665 -2949
rect 666 -2955 669 -2949
rect 673 -2955 676 -2949
rect 680 -2955 683 -2949
rect 687 -2955 690 -2949
rect 694 -2955 697 -2949
rect 701 -2955 704 -2949
rect 708 -2955 711 -2949
rect 715 -2955 718 -2949
rect 722 -2955 725 -2949
rect 729 -2955 732 -2949
rect 736 -2955 739 -2949
rect 743 -2955 746 -2949
rect 750 -2955 753 -2949
rect 757 -2955 760 -2949
rect 764 -2955 767 -2949
rect 771 -2955 774 -2949
rect 778 -2955 784 -2949
rect 785 -2955 788 -2949
rect 792 -2955 795 -2949
rect 799 -2955 802 -2949
rect 806 -2955 809 -2949
rect 813 -2955 816 -2949
rect 820 -2955 826 -2949
rect 827 -2955 830 -2949
rect 834 -2955 837 -2949
rect 841 -2955 844 -2949
rect 848 -2955 854 -2949
rect 855 -2955 858 -2949
rect 862 -2955 868 -2949
rect 869 -2955 872 -2949
rect 876 -2955 879 -2949
rect 883 -2955 886 -2949
rect 890 -2955 893 -2949
rect 897 -2955 900 -2949
rect 904 -2955 907 -2949
rect 911 -2955 917 -2949
rect 918 -2955 921 -2949
rect 925 -2955 928 -2949
rect 932 -2955 935 -2949
rect 939 -2955 945 -2949
rect 946 -2955 949 -2949
rect 953 -2955 956 -2949
rect 960 -2955 963 -2949
rect 967 -2955 973 -2949
rect 974 -2955 977 -2949
rect 981 -2955 984 -2949
rect 988 -2955 991 -2949
rect 995 -2955 998 -2949
rect 1002 -2955 1005 -2949
rect 1009 -2955 1012 -2949
rect 1016 -2955 1019 -2949
rect 1023 -2955 1029 -2949
rect 1030 -2955 1036 -2949
rect 1037 -2955 1040 -2949
rect 1044 -2955 1047 -2949
rect 1051 -2955 1057 -2949
rect 1058 -2955 1061 -2949
rect 1065 -2955 1068 -2949
rect 1072 -2955 1075 -2949
rect 1079 -2955 1082 -2949
rect 1086 -2955 1089 -2949
rect 1093 -2955 1099 -2949
rect 1100 -2955 1103 -2949
rect 1107 -2955 1110 -2949
rect 1114 -2955 1117 -2949
rect 1121 -2955 1124 -2949
rect 1128 -2955 1131 -2949
rect 1135 -2955 1138 -2949
rect 1142 -2955 1145 -2949
rect 1149 -2955 1152 -2949
rect 1156 -2955 1159 -2949
rect 1163 -2955 1166 -2949
rect 1170 -2955 1173 -2949
rect 1177 -2955 1180 -2949
rect 1184 -2955 1187 -2949
rect 1191 -2955 1194 -2949
rect 1198 -2955 1204 -2949
rect 1205 -2955 1208 -2949
rect 1212 -2955 1215 -2949
rect 1219 -2955 1222 -2949
rect 1226 -2955 1229 -2949
rect 1233 -2955 1236 -2949
rect 1240 -2955 1243 -2949
rect 1247 -2955 1250 -2949
rect 1254 -2955 1257 -2949
rect 1261 -2955 1264 -2949
rect 1268 -2955 1271 -2949
rect 1275 -2955 1278 -2949
rect 1282 -2955 1285 -2949
rect 1289 -2955 1292 -2949
rect 1296 -2955 1299 -2949
rect 1303 -2955 1306 -2949
rect 1310 -2955 1313 -2949
rect 1317 -2955 1320 -2949
rect 1324 -2955 1327 -2949
rect 1331 -2955 1337 -2949
rect 1338 -2955 1341 -2949
rect 1345 -2955 1348 -2949
rect 1352 -2955 1355 -2949
rect 1359 -2955 1362 -2949
rect 1366 -2955 1369 -2949
rect 1373 -2955 1376 -2949
rect 1380 -2955 1383 -2949
rect 1387 -2955 1390 -2949
rect 1394 -2955 1397 -2949
rect 1401 -2955 1404 -2949
rect 1408 -2955 1411 -2949
rect 1415 -2955 1418 -2949
rect 1422 -2955 1425 -2949
rect 1429 -2955 1432 -2949
rect 1436 -2955 1439 -2949
rect 1443 -2955 1446 -2949
rect 1450 -2955 1453 -2949
rect 1457 -2955 1460 -2949
rect 1464 -2955 1467 -2949
rect 1471 -2955 1474 -2949
rect 1478 -2955 1481 -2949
rect 1485 -2955 1488 -2949
rect 1492 -2955 1495 -2949
rect 1499 -2955 1502 -2949
rect 1506 -2955 1509 -2949
rect 1513 -2955 1516 -2949
rect 1520 -2955 1523 -2949
rect 1527 -2955 1530 -2949
rect 1534 -2955 1537 -2949
rect 1541 -2955 1544 -2949
rect 1548 -2955 1551 -2949
rect 1555 -2955 1558 -2949
rect 1562 -2955 1565 -2949
rect 1569 -2955 1572 -2949
rect 1576 -2955 1579 -2949
rect 1583 -2955 1586 -2949
rect 1590 -2955 1593 -2949
rect 1597 -2955 1600 -2949
rect 1604 -2955 1607 -2949
rect 1611 -2955 1614 -2949
rect 1618 -2955 1621 -2949
rect 1625 -2955 1628 -2949
rect 1632 -2955 1635 -2949
rect 1639 -2955 1645 -2949
rect 1646 -2955 1649 -2949
rect 1653 -2955 1656 -2949
rect 1660 -2955 1663 -2949
rect 1667 -2955 1670 -2949
rect 1674 -2955 1677 -2949
rect 1681 -2955 1684 -2949
rect 1688 -2955 1691 -2949
rect 1695 -2955 1698 -2949
rect 1702 -2955 1708 -2949
rect 1 -3082 7 -3076
rect 8 -3082 14 -3076
rect 15 -3082 21 -3076
rect 22 -3082 28 -3076
rect 29 -3082 32 -3076
rect 36 -3082 39 -3076
rect 43 -3082 46 -3076
rect 50 -3082 53 -3076
rect 57 -3082 63 -3076
rect 64 -3082 67 -3076
rect 71 -3082 74 -3076
rect 78 -3082 84 -3076
rect 85 -3082 91 -3076
rect 92 -3082 95 -3076
rect 99 -3082 102 -3076
rect 106 -3082 109 -3076
rect 113 -3082 116 -3076
rect 120 -3082 123 -3076
rect 127 -3082 130 -3076
rect 134 -3082 140 -3076
rect 141 -3082 147 -3076
rect 148 -3082 154 -3076
rect 155 -3082 158 -3076
rect 162 -3082 165 -3076
rect 169 -3082 172 -3076
rect 176 -3082 179 -3076
rect 183 -3082 189 -3076
rect 190 -3082 193 -3076
rect 197 -3082 203 -3076
rect 204 -3082 210 -3076
rect 211 -3082 217 -3076
rect 218 -3082 221 -3076
rect 225 -3082 228 -3076
rect 232 -3082 235 -3076
rect 239 -3082 242 -3076
rect 246 -3082 249 -3076
rect 253 -3082 256 -3076
rect 260 -3082 263 -3076
rect 267 -3082 270 -3076
rect 274 -3082 277 -3076
rect 281 -3082 284 -3076
rect 288 -3082 291 -3076
rect 295 -3082 298 -3076
rect 302 -3082 305 -3076
rect 309 -3082 312 -3076
rect 316 -3082 319 -3076
rect 323 -3082 326 -3076
rect 330 -3082 333 -3076
rect 337 -3082 340 -3076
rect 344 -3082 350 -3076
rect 351 -3082 354 -3076
rect 358 -3082 361 -3076
rect 365 -3082 371 -3076
rect 372 -3082 375 -3076
rect 379 -3082 382 -3076
rect 386 -3082 389 -3076
rect 393 -3082 399 -3076
rect 400 -3082 403 -3076
rect 407 -3082 410 -3076
rect 414 -3082 417 -3076
rect 421 -3082 424 -3076
rect 428 -3082 431 -3076
rect 435 -3082 438 -3076
rect 442 -3082 445 -3076
rect 449 -3082 455 -3076
rect 456 -3082 459 -3076
rect 463 -3082 466 -3076
rect 470 -3082 473 -3076
rect 477 -3082 480 -3076
rect 484 -3082 487 -3076
rect 491 -3082 494 -3076
rect 498 -3082 501 -3076
rect 505 -3082 508 -3076
rect 512 -3082 515 -3076
rect 519 -3082 522 -3076
rect 526 -3082 529 -3076
rect 533 -3082 536 -3076
rect 540 -3082 543 -3076
rect 547 -3082 550 -3076
rect 554 -3082 557 -3076
rect 561 -3082 564 -3076
rect 568 -3082 571 -3076
rect 575 -3082 578 -3076
rect 582 -3082 585 -3076
rect 589 -3082 592 -3076
rect 596 -3082 599 -3076
rect 603 -3082 606 -3076
rect 610 -3082 613 -3076
rect 617 -3082 623 -3076
rect 624 -3082 627 -3076
rect 631 -3082 637 -3076
rect 638 -3082 641 -3076
rect 645 -3082 648 -3076
rect 652 -3082 655 -3076
rect 659 -3082 662 -3076
rect 666 -3082 669 -3076
rect 673 -3082 676 -3076
rect 680 -3082 683 -3076
rect 687 -3082 693 -3076
rect 694 -3082 697 -3076
rect 701 -3082 704 -3076
rect 708 -3082 711 -3076
rect 715 -3082 718 -3076
rect 722 -3082 725 -3076
rect 729 -3082 732 -3076
rect 736 -3082 742 -3076
rect 743 -3082 746 -3076
rect 750 -3082 753 -3076
rect 757 -3082 763 -3076
rect 764 -3082 767 -3076
rect 771 -3082 774 -3076
rect 778 -3082 781 -3076
rect 785 -3082 791 -3076
rect 792 -3082 795 -3076
rect 799 -3082 805 -3076
rect 806 -3082 809 -3076
rect 813 -3082 816 -3076
rect 820 -3082 823 -3076
rect 827 -3082 833 -3076
rect 834 -3082 840 -3076
rect 841 -3082 844 -3076
rect 848 -3082 851 -3076
rect 855 -3082 858 -3076
rect 862 -3082 865 -3076
rect 869 -3082 872 -3076
rect 876 -3082 882 -3076
rect 883 -3082 886 -3076
rect 890 -3082 893 -3076
rect 897 -3082 903 -3076
rect 904 -3082 907 -3076
rect 911 -3082 917 -3076
rect 918 -3082 921 -3076
rect 925 -3082 928 -3076
rect 932 -3082 935 -3076
rect 939 -3082 942 -3076
rect 946 -3082 952 -3076
rect 953 -3082 956 -3076
rect 960 -3082 963 -3076
rect 967 -3082 970 -3076
rect 974 -3082 980 -3076
rect 981 -3082 984 -3076
rect 988 -3082 991 -3076
rect 995 -3082 998 -3076
rect 1002 -3082 1005 -3076
rect 1009 -3082 1012 -3076
rect 1016 -3082 1022 -3076
rect 1023 -3082 1026 -3076
rect 1030 -3082 1033 -3076
rect 1037 -3082 1040 -3076
rect 1044 -3082 1047 -3076
rect 1051 -3082 1054 -3076
rect 1058 -3082 1061 -3076
rect 1065 -3082 1068 -3076
rect 1072 -3082 1075 -3076
rect 1079 -3082 1085 -3076
rect 1086 -3082 1092 -3076
rect 1093 -3082 1096 -3076
rect 1100 -3082 1103 -3076
rect 1107 -3082 1110 -3076
rect 1114 -3082 1117 -3076
rect 1121 -3082 1124 -3076
rect 1128 -3082 1131 -3076
rect 1135 -3082 1138 -3076
rect 1142 -3082 1145 -3076
rect 1149 -3082 1152 -3076
rect 1156 -3082 1159 -3076
rect 1163 -3082 1166 -3076
rect 1170 -3082 1173 -3076
rect 1177 -3082 1180 -3076
rect 1184 -3082 1187 -3076
rect 1191 -3082 1194 -3076
rect 1198 -3082 1201 -3076
rect 1205 -3082 1208 -3076
rect 1212 -3082 1215 -3076
rect 1219 -3082 1222 -3076
rect 1226 -3082 1229 -3076
rect 1233 -3082 1236 -3076
rect 1240 -3082 1243 -3076
rect 1247 -3082 1250 -3076
rect 1254 -3082 1257 -3076
rect 1261 -3082 1264 -3076
rect 1268 -3082 1271 -3076
rect 1275 -3082 1278 -3076
rect 1282 -3082 1285 -3076
rect 1289 -3082 1292 -3076
rect 1296 -3082 1299 -3076
rect 1303 -3082 1306 -3076
rect 1310 -3082 1313 -3076
rect 1317 -3082 1320 -3076
rect 1324 -3082 1327 -3076
rect 1331 -3082 1334 -3076
rect 1338 -3082 1341 -3076
rect 1345 -3082 1348 -3076
rect 1352 -3082 1355 -3076
rect 1359 -3082 1362 -3076
rect 1366 -3082 1369 -3076
rect 1373 -3082 1376 -3076
rect 1380 -3082 1383 -3076
rect 1387 -3082 1390 -3076
rect 1394 -3082 1397 -3076
rect 1401 -3082 1404 -3076
rect 1408 -3082 1411 -3076
rect 1415 -3082 1418 -3076
rect 1422 -3082 1425 -3076
rect 1429 -3082 1432 -3076
rect 1436 -3082 1439 -3076
rect 1443 -3082 1446 -3076
rect 1450 -3082 1453 -3076
rect 1457 -3082 1460 -3076
rect 1464 -3082 1467 -3076
rect 1471 -3082 1474 -3076
rect 1478 -3082 1481 -3076
rect 1485 -3082 1488 -3076
rect 1492 -3082 1495 -3076
rect 1499 -3082 1502 -3076
rect 1506 -3082 1509 -3076
rect 1513 -3082 1516 -3076
rect 1520 -3082 1523 -3076
rect 1527 -3082 1530 -3076
rect 1534 -3082 1537 -3076
rect 1541 -3082 1544 -3076
rect 1548 -3082 1551 -3076
rect 1555 -3082 1558 -3076
rect 1562 -3082 1565 -3076
rect 1569 -3082 1572 -3076
rect 1576 -3082 1579 -3076
rect 1583 -3082 1586 -3076
rect 1590 -3082 1593 -3076
rect 1597 -3082 1600 -3076
rect 1604 -3082 1607 -3076
rect 1611 -3082 1614 -3076
rect 1618 -3082 1621 -3076
rect 1625 -3082 1628 -3076
rect 1632 -3082 1635 -3076
rect 1639 -3082 1642 -3076
rect 1646 -3082 1649 -3076
rect 1653 -3082 1656 -3076
rect 1 -3221 7 -3215
rect 8 -3221 14 -3215
rect 15 -3221 21 -3215
rect 22 -3221 28 -3215
rect 64 -3221 70 -3215
rect 71 -3221 74 -3215
rect 78 -3221 81 -3215
rect 85 -3221 88 -3215
rect 92 -3221 95 -3215
rect 99 -3221 102 -3215
rect 106 -3221 109 -3215
rect 113 -3221 119 -3215
rect 120 -3221 123 -3215
rect 127 -3221 133 -3215
rect 134 -3221 137 -3215
rect 141 -3221 144 -3215
rect 148 -3221 154 -3215
rect 155 -3221 158 -3215
rect 162 -3221 165 -3215
rect 169 -3221 172 -3215
rect 176 -3221 179 -3215
rect 183 -3221 186 -3215
rect 190 -3221 193 -3215
rect 197 -3221 200 -3215
rect 204 -3221 207 -3215
rect 211 -3221 214 -3215
rect 218 -3221 221 -3215
rect 225 -3221 228 -3215
rect 232 -3221 235 -3215
rect 239 -3221 245 -3215
rect 246 -3221 249 -3215
rect 253 -3221 256 -3215
rect 260 -3221 263 -3215
rect 267 -3221 270 -3215
rect 274 -3221 277 -3215
rect 281 -3221 284 -3215
rect 288 -3221 291 -3215
rect 295 -3221 298 -3215
rect 302 -3221 305 -3215
rect 309 -3221 312 -3215
rect 316 -3221 319 -3215
rect 323 -3221 326 -3215
rect 330 -3221 333 -3215
rect 337 -3221 340 -3215
rect 344 -3221 347 -3215
rect 351 -3221 354 -3215
rect 358 -3221 361 -3215
rect 365 -3221 368 -3215
rect 372 -3221 375 -3215
rect 379 -3221 382 -3215
rect 386 -3221 389 -3215
rect 393 -3221 396 -3215
rect 400 -3221 406 -3215
rect 407 -3221 410 -3215
rect 414 -3221 417 -3215
rect 421 -3221 424 -3215
rect 428 -3221 434 -3215
rect 435 -3221 438 -3215
rect 442 -3221 445 -3215
rect 449 -3221 452 -3215
rect 456 -3221 459 -3215
rect 463 -3221 466 -3215
rect 470 -3221 476 -3215
rect 477 -3221 480 -3215
rect 484 -3221 487 -3215
rect 491 -3221 497 -3215
rect 498 -3221 504 -3215
rect 505 -3221 508 -3215
rect 512 -3221 515 -3215
rect 519 -3221 522 -3215
rect 526 -3221 529 -3215
rect 533 -3221 539 -3215
rect 540 -3221 546 -3215
rect 547 -3221 550 -3215
rect 554 -3221 557 -3215
rect 561 -3221 564 -3215
rect 568 -3221 571 -3215
rect 575 -3221 581 -3215
rect 582 -3221 585 -3215
rect 589 -3221 595 -3215
rect 596 -3221 599 -3215
rect 603 -3221 606 -3215
rect 610 -3221 613 -3215
rect 617 -3221 620 -3215
rect 624 -3221 627 -3215
rect 631 -3221 634 -3215
rect 638 -3221 641 -3215
rect 645 -3221 648 -3215
rect 652 -3221 658 -3215
rect 659 -3221 662 -3215
rect 666 -3221 669 -3215
rect 673 -3221 676 -3215
rect 680 -3221 686 -3215
rect 687 -3221 690 -3215
rect 694 -3221 697 -3215
rect 701 -3221 704 -3215
rect 708 -3221 711 -3215
rect 715 -3221 718 -3215
rect 722 -3221 725 -3215
rect 729 -3221 732 -3215
rect 736 -3221 739 -3215
rect 743 -3221 746 -3215
rect 750 -3221 753 -3215
rect 757 -3221 760 -3215
rect 764 -3221 767 -3215
rect 771 -3221 774 -3215
rect 778 -3221 784 -3215
rect 785 -3221 788 -3215
rect 792 -3221 798 -3215
rect 799 -3221 802 -3215
rect 806 -3221 809 -3215
rect 813 -3221 816 -3215
rect 820 -3221 826 -3215
rect 827 -3221 830 -3215
rect 834 -3221 840 -3215
rect 841 -3221 844 -3215
rect 848 -3221 851 -3215
rect 855 -3221 858 -3215
rect 862 -3221 865 -3215
rect 869 -3221 872 -3215
rect 876 -3221 879 -3215
rect 883 -3221 886 -3215
rect 890 -3221 896 -3215
rect 897 -3221 900 -3215
rect 904 -3221 907 -3215
rect 911 -3221 914 -3215
rect 918 -3221 921 -3215
rect 925 -3221 928 -3215
rect 932 -3221 935 -3215
rect 939 -3221 942 -3215
rect 946 -3221 952 -3215
rect 953 -3221 956 -3215
rect 960 -3221 963 -3215
rect 967 -3221 970 -3215
rect 974 -3221 977 -3215
rect 981 -3221 984 -3215
rect 988 -3221 991 -3215
rect 995 -3221 1001 -3215
rect 1002 -3221 1005 -3215
rect 1009 -3221 1015 -3215
rect 1016 -3221 1019 -3215
rect 1023 -3221 1026 -3215
rect 1030 -3221 1033 -3215
rect 1037 -3221 1040 -3215
rect 1044 -3221 1047 -3215
rect 1051 -3221 1054 -3215
rect 1058 -3221 1064 -3215
rect 1065 -3221 1068 -3215
rect 1072 -3221 1075 -3215
rect 1079 -3221 1082 -3215
rect 1086 -3221 1092 -3215
rect 1093 -3221 1096 -3215
rect 1100 -3221 1103 -3215
rect 1107 -3221 1110 -3215
rect 1114 -3221 1117 -3215
rect 1121 -3221 1124 -3215
rect 1128 -3221 1131 -3215
rect 1135 -3221 1138 -3215
rect 1142 -3221 1145 -3215
rect 1149 -3221 1152 -3215
rect 1156 -3221 1159 -3215
rect 1163 -3221 1166 -3215
rect 1170 -3221 1173 -3215
rect 1177 -3221 1180 -3215
rect 1184 -3221 1187 -3215
rect 1191 -3221 1194 -3215
rect 1198 -3221 1201 -3215
rect 1205 -3221 1208 -3215
rect 1212 -3221 1215 -3215
rect 1219 -3221 1222 -3215
rect 1226 -3221 1229 -3215
rect 1233 -3221 1236 -3215
rect 1240 -3221 1243 -3215
rect 1247 -3221 1250 -3215
rect 1254 -3221 1257 -3215
rect 1261 -3221 1264 -3215
rect 1268 -3221 1271 -3215
rect 1275 -3221 1278 -3215
rect 1282 -3221 1285 -3215
rect 1289 -3221 1292 -3215
rect 1296 -3221 1302 -3215
rect 1303 -3221 1306 -3215
rect 1310 -3221 1313 -3215
rect 1317 -3221 1320 -3215
rect 1324 -3221 1327 -3215
rect 1331 -3221 1334 -3215
rect 1338 -3221 1341 -3215
rect 1345 -3221 1351 -3215
rect 1352 -3221 1358 -3215
rect 1359 -3221 1362 -3215
rect 1366 -3221 1369 -3215
rect 1373 -3221 1376 -3215
rect 1380 -3221 1383 -3215
rect 1387 -3221 1390 -3215
rect 1394 -3221 1397 -3215
rect 1401 -3221 1404 -3215
rect 1408 -3221 1414 -3215
rect 1415 -3221 1418 -3215
rect 1422 -3221 1425 -3215
rect 1429 -3221 1432 -3215
rect 1436 -3221 1439 -3215
rect 1443 -3221 1446 -3215
rect 1450 -3221 1453 -3215
rect 1457 -3221 1460 -3215
rect 1464 -3221 1467 -3215
rect 1471 -3221 1477 -3215
rect 1478 -3221 1481 -3215
rect 1485 -3221 1488 -3215
rect 1492 -3221 1495 -3215
rect 1499 -3221 1502 -3215
rect 1506 -3221 1509 -3215
rect 1513 -3221 1516 -3215
rect 1520 -3221 1523 -3215
rect 1604 -3221 1607 -3215
rect 1 -3314 7 -3308
rect 8 -3314 14 -3308
rect 15 -3314 21 -3308
rect 22 -3314 28 -3308
rect 127 -3314 133 -3308
rect 134 -3314 137 -3308
rect 162 -3314 165 -3308
rect 169 -3314 172 -3308
rect 176 -3314 179 -3308
rect 183 -3314 186 -3308
rect 190 -3314 193 -3308
rect 197 -3314 200 -3308
rect 204 -3314 207 -3308
rect 211 -3314 214 -3308
rect 218 -3314 221 -3308
rect 225 -3314 228 -3308
rect 232 -3314 235 -3308
rect 239 -3314 242 -3308
rect 246 -3314 249 -3308
rect 253 -3314 256 -3308
rect 260 -3314 263 -3308
rect 267 -3314 270 -3308
rect 274 -3314 277 -3308
rect 281 -3314 284 -3308
rect 288 -3314 291 -3308
rect 295 -3314 298 -3308
rect 302 -3314 305 -3308
rect 309 -3314 312 -3308
rect 316 -3314 319 -3308
rect 323 -3314 326 -3308
rect 330 -3314 333 -3308
rect 337 -3314 340 -3308
rect 344 -3314 350 -3308
rect 351 -3314 354 -3308
rect 358 -3314 361 -3308
rect 365 -3314 368 -3308
rect 372 -3314 375 -3308
rect 379 -3314 382 -3308
rect 386 -3314 389 -3308
rect 393 -3314 396 -3308
rect 400 -3314 406 -3308
rect 407 -3314 410 -3308
rect 414 -3314 417 -3308
rect 421 -3314 424 -3308
rect 428 -3314 431 -3308
rect 435 -3314 441 -3308
rect 442 -3314 448 -3308
rect 449 -3314 452 -3308
rect 456 -3314 459 -3308
rect 463 -3314 466 -3308
rect 470 -3314 473 -3308
rect 477 -3314 480 -3308
rect 484 -3314 487 -3308
rect 491 -3314 497 -3308
rect 498 -3314 501 -3308
rect 505 -3314 508 -3308
rect 512 -3314 515 -3308
rect 519 -3314 522 -3308
rect 526 -3314 532 -3308
rect 533 -3314 536 -3308
rect 540 -3314 546 -3308
rect 547 -3314 550 -3308
rect 554 -3314 557 -3308
rect 561 -3314 564 -3308
rect 568 -3314 571 -3308
rect 575 -3314 578 -3308
rect 582 -3314 585 -3308
rect 589 -3314 592 -3308
rect 596 -3314 599 -3308
rect 603 -3314 606 -3308
rect 610 -3314 613 -3308
rect 617 -3314 623 -3308
rect 624 -3314 627 -3308
rect 631 -3314 634 -3308
rect 638 -3314 641 -3308
rect 645 -3314 648 -3308
rect 652 -3314 655 -3308
rect 659 -3314 662 -3308
rect 666 -3314 669 -3308
rect 673 -3314 679 -3308
rect 680 -3314 683 -3308
rect 687 -3314 693 -3308
rect 694 -3314 697 -3308
rect 701 -3314 707 -3308
rect 708 -3314 711 -3308
rect 715 -3314 718 -3308
rect 722 -3314 725 -3308
rect 729 -3314 732 -3308
rect 736 -3314 739 -3308
rect 743 -3314 746 -3308
rect 750 -3314 753 -3308
rect 757 -3314 760 -3308
rect 764 -3314 767 -3308
rect 771 -3314 774 -3308
rect 778 -3314 781 -3308
rect 785 -3314 791 -3308
rect 792 -3314 795 -3308
rect 799 -3314 802 -3308
rect 806 -3314 809 -3308
rect 813 -3314 816 -3308
rect 820 -3314 823 -3308
rect 827 -3314 830 -3308
rect 834 -3314 837 -3308
rect 841 -3314 844 -3308
rect 848 -3314 851 -3308
rect 855 -3314 858 -3308
rect 862 -3314 865 -3308
rect 869 -3314 875 -3308
rect 876 -3314 882 -3308
rect 883 -3314 886 -3308
rect 890 -3314 893 -3308
rect 897 -3314 903 -3308
rect 904 -3314 910 -3308
rect 911 -3314 917 -3308
rect 918 -3314 921 -3308
rect 925 -3314 928 -3308
rect 932 -3314 935 -3308
rect 939 -3314 942 -3308
rect 946 -3314 949 -3308
rect 953 -3314 956 -3308
rect 960 -3314 963 -3308
rect 967 -3314 970 -3308
rect 974 -3314 977 -3308
rect 981 -3314 987 -3308
rect 988 -3314 991 -3308
rect 995 -3314 998 -3308
rect 1002 -3314 1005 -3308
rect 1009 -3314 1012 -3308
rect 1016 -3314 1022 -3308
rect 1023 -3314 1026 -3308
rect 1030 -3314 1033 -3308
rect 1037 -3314 1040 -3308
rect 1044 -3314 1047 -3308
rect 1051 -3314 1054 -3308
rect 1058 -3314 1061 -3308
rect 1065 -3314 1068 -3308
rect 1072 -3314 1075 -3308
rect 1079 -3314 1082 -3308
rect 1086 -3314 1089 -3308
rect 1093 -3314 1096 -3308
rect 1100 -3314 1103 -3308
rect 1107 -3314 1113 -3308
rect 1114 -3314 1117 -3308
rect 1121 -3314 1124 -3308
rect 1128 -3314 1134 -3308
rect 1135 -3314 1138 -3308
rect 1142 -3314 1145 -3308
rect 1149 -3314 1152 -3308
rect 1156 -3314 1159 -3308
rect 1163 -3314 1166 -3308
rect 1170 -3314 1173 -3308
rect 1177 -3314 1183 -3308
rect 1184 -3314 1190 -3308
rect 1191 -3314 1194 -3308
rect 1198 -3314 1201 -3308
rect 1205 -3314 1211 -3308
rect 1212 -3314 1218 -3308
rect 1219 -3314 1222 -3308
rect 1226 -3314 1229 -3308
rect 1233 -3314 1236 -3308
rect 1240 -3314 1243 -3308
rect 1247 -3314 1253 -3308
rect 1254 -3314 1260 -3308
rect 1261 -3314 1267 -3308
rect 1268 -3314 1271 -3308
rect 1275 -3314 1278 -3308
rect 1282 -3314 1285 -3308
rect 1289 -3314 1292 -3308
rect 1296 -3314 1299 -3308
rect 1303 -3314 1306 -3308
rect 1310 -3314 1313 -3308
rect 1317 -3314 1320 -3308
rect 1324 -3314 1327 -3308
rect 1331 -3314 1334 -3308
rect 1338 -3314 1341 -3308
rect 1345 -3314 1348 -3308
rect 1352 -3314 1355 -3308
rect 1359 -3314 1362 -3308
rect 1380 -3314 1383 -3308
rect 1387 -3314 1390 -3308
rect 1527 -3314 1533 -3308
rect 1583 -3314 1586 -3308
rect 1 -3411 7 -3405
rect 8 -3411 14 -3405
rect 15 -3411 21 -3405
rect 22 -3411 28 -3405
rect 29 -3411 35 -3405
rect 36 -3411 42 -3405
rect 43 -3411 49 -3405
rect 50 -3411 56 -3405
rect 57 -3411 63 -3405
rect 239 -3411 242 -3405
rect 246 -3411 249 -3405
rect 267 -3411 270 -3405
rect 281 -3411 284 -3405
rect 288 -3411 294 -3405
rect 295 -3411 301 -3405
rect 302 -3411 305 -3405
rect 309 -3411 312 -3405
rect 316 -3411 319 -3405
rect 323 -3411 326 -3405
rect 330 -3411 333 -3405
rect 337 -3411 340 -3405
rect 344 -3411 347 -3405
rect 351 -3411 354 -3405
rect 358 -3411 361 -3405
rect 365 -3411 368 -3405
rect 372 -3411 378 -3405
rect 379 -3411 382 -3405
rect 386 -3411 389 -3405
rect 393 -3411 396 -3405
rect 400 -3411 403 -3405
rect 407 -3411 410 -3405
rect 414 -3411 417 -3405
rect 421 -3411 424 -3405
rect 428 -3411 431 -3405
rect 435 -3411 438 -3405
rect 442 -3411 445 -3405
rect 449 -3411 452 -3405
rect 456 -3411 459 -3405
rect 463 -3411 466 -3405
rect 470 -3411 473 -3405
rect 477 -3411 480 -3405
rect 484 -3411 487 -3405
rect 491 -3411 494 -3405
rect 498 -3411 504 -3405
rect 505 -3411 508 -3405
rect 512 -3411 515 -3405
rect 519 -3411 525 -3405
rect 526 -3411 529 -3405
rect 533 -3411 536 -3405
rect 540 -3411 543 -3405
rect 547 -3411 550 -3405
rect 554 -3411 557 -3405
rect 561 -3411 564 -3405
rect 568 -3411 571 -3405
rect 575 -3411 581 -3405
rect 582 -3411 585 -3405
rect 589 -3411 592 -3405
rect 596 -3411 599 -3405
rect 603 -3411 606 -3405
rect 610 -3411 616 -3405
rect 617 -3411 620 -3405
rect 624 -3411 627 -3405
rect 631 -3411 634 -3405
rect 638 -3411 641 -3405
rect 645 -3411 648 -3405
rect 652 -3411 655 -3405
rect 659 -3411 662 -3405
rect 666 -3411 669 -3405
rect 673 -3411 676 -3405
rect 680 -3411 683 -3405
rect 687 -3411 690 -3405
rect 694 -3411 697 -3405
rect 701 -3411 704 -3405
rect 708 -3411 711 -3405
rect 715 -3411 718 -3405
rect 722 -3411 725 -3405
rect 729 -3411 735 -3405
rect 736 -3411 739 -3405
rect 743 -3411 746 -3405
rect 750 -3411 753 -3405
rect 757 -3411 760 -3405
rect 764 -3411 767 -3405
rect 771 -3411 774 -3405
rect 778 -3411 781 -3405
rect 785 -3411 788 -3405
rect 792 -3411 795 -3405
rect 799 -3411 805 -3405
rect 806 -3411 809 -3405
rect 813 -3411 816 -3405
rect 820 -3411 823 -3405
rect 827 -3411 830 -3405
rect 834 -3411 837 -3405
rect 841 -3411 844 -3405
rect 848 -3411 851 -3405
rect 855 -3411 858 -3405
rect 862 -3411 865 -3405
rect 869 -3411 872 -3405
rect 876 -3411 882 -3405
rect 883 -3411 886 -3405
rect 890 -3411 896 -3405
rect 897 -3411 900 -3405
rect 904 -3411 907 -3405
rect 911 -3411 914 -3405
rect 918 -3411 921 -3405
rect 925 -3411 928 -3405
rect 932 -3411 935 -3405
rect 939 -3411 942 -3405
rect 946 -3411 952 -3405
rect 953 -3411 956 -3405
rect 960 -3411 963 -3405
rect 967 -3411 970 -3405
rect 974 -3411 977 -3405
rect 981 -3411 984 -3405
rect 988 -3411 991 -3405
rect 995 -3411 998 -3405
rect 1002 -3411 1005 -3405
rect 1009 -3411 1015 -3405
rect 1016 -3411 1022 -3405
rect 1023 -3411 1029 -3405
rect 1030 -3411 1033 -3405
rect 1037 -3411 1043 -3405
rect 1044 -3411 1047 -3405
rect 1051 -3411 1057 -3405
rect 1058 -3411 1064 -3405
rect 1065 -3411 1068 -3405
rect 1072 -3411 1075 -3405
rect 1079 -3411 1082 -3405
rect 1086 -3411 1089 -3405
rect 1093 -3411 1096 -3405
rect 1100 -3411 1103 -3405
rect 1107 -3411 1113 -3405
rect 1114 -3411 1117 -3405
rect 1121 -3411 1124 -3405
rect 1128 -3411 1131 -3405
rect 1135 -3411 1138 -3405
rect 1142 -3411 1145 -3405
rect 1149 -3411 1155 -3405
rect 1156 -3411 1162 -3405
rect 1163 -3411 1169 -3405
rect 1170 -3411 1173 -3405
rect 1184 -3411 1187 -3405
rect 1191 -3411 1194 -3405
rect 1198 -3411 1201 -3405
rect 1205 -3411 1208 -3405
rect 1212 -3411 1218 -3405
rect 1233 -3411 1236 -3405
rect 1240 -3411 1243 -3405
rect 1247 -3411 1250 -3405
rect 1261 -3411 1267 -3405
rect 1310 -3411 1313 -3405
rect 1317 -3411 1320 -3405
rect 1331 -3411 1334 -3405
rect 1373 -3411 1376 -3405
rect 1380 -3411 1383 -3405
rect 1387 -3411 1390 -3405
rect 1576 -3411 1579 -3405
rect 1 -3458 7 -3452
rect 8 -3458 14 -3452
rect 15 -3458 21 -3452
rect 22 -3458 28 -3452
rect 29 -3458 35 -3452
rect 36 -3458 42 -3452
rect 43 -3458 49 -3452
rect 50 -3458 56 -3452
rect 57 -3458 63 -3452
rect 64 -3458 70 -3452
rect 71 -3458 77 -3452
rect 78 -3458 84 -3452
rect 85 -3458 91 -3452
rect 92 -3458 98 -3452
rect 99 -3458 105 -3452
rect 260 -3458 263 -3452
rect 309 -3458 312 -3452
rect 316 -3458 319 -3452
rect 337 -3458 340 -3452
rect 344 -3458 347 -3452
rect 351 -3458 357 -3452
rect 358 -3458 361 -3452
rect 365 -3458 368 -3452
rect 372 -3458 375 -3452
rect 379 -3458 382 -3452
rect 386 -3458 389 -3452
rect 393 -3458 396 -3452
rect 400 -3458 403 -3452
rect 407 -3458 413 -3452
rect 414 -3458 417 -3452
rect 421 -3458 424 -3452
rect 428 -3458 431 -3452
rect 435 -3458 438 -3452
rect 442 -3458 445 -3452
rect 449 -3458 452 -3452
rect 456 -3458 459 -3452
rect 463 -3458 466 -3452
rect 470 -3458 476 -3452
rect 477 -3458 480 -3452
rect 484 -3458 487 -3452
rect 491 -3458 494 -3452
rect 498 -3458 501 -3452
rect 505 -3458 511 -3452
rect 512 -3458 515 -3452
rect 519 -3458 522 -3452
rect 526 -3458 529 -3452
rect 533 -3458 536 -3452
rect 540 -3458 543 -3452
rect 547 -3458 550 -3452
rect 554 -3458 557 -3452
rect 561 -3458 564 -3452
rect 568 -3458 571 -3452
rect 575 -3458 578 -3452
rect 582 -3458 588 -3452
rect 589 -3458 595 -3452
rect 596 -3458 599 -3452
rect 603 -3458 609 -3452
rect 610 -3458 613 -3452
rect 617 -3458 623 -3452
rect 624 -3458 627 -3452
rect 631 -3458 634 -3452
rect 638 -3458 641 -3452
rect 645 -3458 648 -3452
rect 652 -3458 658 -3452
rect 659 -3458 665 -3452
rect 666 -3458 669 -3452
rect 673 -3458 676 -3452
rect 680 -3458 683 -3452
rect 687 -3458 690 -3452
rect 694 -3458 697 -3452
rect 701 -3458 704 -3452
rect 708 -3458 711 -3452
rect 715 -3458 721 -3452
rect 722 -3458 725 -3452
rect 729 -3458 732 -3452
rect 736 -3458 739 -3452
rect 743 -3458 746 -3452
rect 750 -3458 753 -3452
rect 757 -3458 760 -3452
rect 764 -3458 767 -3452
rect 771 -3458 774 -3452
rect 778 -3458 781 -3452
rect 785 -3458 788 -3452
rect 792 -3458 795 -3452
rect 799 -3458 802 -3452
rect 806 -3458 812 -3452
rect 813 -3458 816 -3452
rect 820 -3458 826 -3452
rect 827 -3458 830 -3452
rect 834 -3458 837 -3452
rect 841 -3458 844 -3452
rect 848 -3458 854 -3452
rect 855 -3458 858 -3452
rect 862 -3458 865 -3452
rect 869 -3458 872 -3452
rect 876 -3458 879 -3452
rect 883 -3458 886 -3452
rect 890 -3458 893 -3452
rect 897 -3458 900 -3452
rect 904 -3458 907 -3452
rect 911 -3458 914 -3452
rect 918 -3458 921 -3452
rect 925 -3458 928 -3452
rect 932 -3458 935 -3452
rect 939 -3458 942 -3452
rect 946 -3458 949 -3452
rect 953 -3458 956 -3452
rect 960 -3458 963 -3452
rect 967 -3458 973 -3452
rect 974 -3458 977 -3452
rect 981 -3458 984 -3452
rect 988 -3458 991 -3452
rect 995 -3458 1001 -3452
rect 1002 -3458 1005 -3452
rect 1009 -3458 1012 -3452
rect 1016 -3458 1019 -3452
rect 1023 -3458 1026 -3452
rect 1030 -3458 1033 -3452
rect 1051 -3458 1054 -3452
rect 1072 -3458 1075 -3452
rect 1079 -3458 1082 -3452
rect 1100 -3458 1103 -3452
rect 1114 -3458 1117 -3452
rect 1121 -3458 1124 -3452
rect 1128 -3458 1131 -3452
rect 1135 -3458 1138 -3452
rect 1142 -3458 1145 -3452
rect 1191 -3458 1194 -3452
rect 1198 -3458 1201 -3452
rect 1205 -3458 1208 -3452
rect 1212 -3458 1215 -3452
rect 1268 -3458 1271 -3452
rect 1296 -3458 1302 -3452
rect 1303 -3458 1306 -3452
rect 1317 -3458 1320 -3452
rect 1345 -3458 1348 -3452
rect 1380 -3458 1383 -3452
rect 1387 -3458 1390 -3452
rect 1394 -3458 1397 -3452
rect 1576 -3458 1579 -3452
rect 1 -3499 7 -3493
rect 8 -3499 14 -3493
rect 15 -3499 21 -3493
rect 22 -3499 28 -3493
rect 29 -3499 35 -3493
rect 36 -3499 42 -3493
rect 43 -3499 49 -3493
rect 50 -3499 56 -3493
rect 57 -3499 63 -3493
rect 64 -3499 70 -3493
rect 71 -3499 77 -3493
rect 78 -3499 84 -3493
rect 85 -3499 91 -3493
rect 92 -3499 98 -3493
rect 99 -3499 105 -3493
rect 106 -3499 112 -3493
rect 113 -3499 119 -3493
rect 120 -3499 126 -3493
rect 267 -3499 270 -3493
rect 281 -3499 287 -3493
rect 295 -3499 298 -3493
rect 365 -3499 368 -3493
rect 372 -3499 375 -3493
rect 379 -3499 382 -3493
rect 386 -3499 392 -3493
rect 407 -3499 410 -3493
rect 421 -3499 427 -3493
rect 428 -3499 431 -3493
rect 435 -3499 441 -3493
rect 442 -3499 445 -3493
rect 449 -3499 452 -3493
rect 456 -3499 459 -3493
rect 470 -3499 473 -3493
rect 477 -3499 480 -3493
rect 484 -3499 487 -3493
rect 491 -3499 494 -3493
rect 498 -3499 501 -3493
rect 505 -3499 508 -3493
rect 512 -3499 515 -3493
rect 526 -3499 529 -3493
rect 533 -3499 536 -3493
rect 540 -3499 543 -3493
rect 547 -3499 550 -3493
rect 554 -3499 557 -3493
rect 561 -3499 564 -3493
rect 568 -3499 571 -3493
rect 575 -3499 578 -3493
rect 582 -3499 585 -3493
rect 589 -3499 592 -3493
rect 603 -3499 606 -3493
rect 617 -3499 620 -3493
rect 631 -3499 634 -3493
rect 638 -3499 641 -3493
rect 645 -3499 648 -3493
rect 652 -3499 658 -3493
rect 687 -3499 690 -3493
rect 694 -3499 697 -3493
rect 701 -3499 704 -3493
rect 708 -3499 711 -3493
rect 715 -3499 718 -3493
rect 722 -3499 728 -3493
rect 729 -3499 735 -3493
rect 736 -3499 739 -3493
rect 743 -3499 746 -3493
rect 750 -3499 756 -3493
rect 757 -3499 760 -3493
rect 764 -3499 767 -3493
rect 771 -3499 774 -3493
rect 785 -3499 788 -3493
rect 792 -3499 795 -3493
rect 799 -3499 802 -3493
rect 806 -3499 809 -3493
rect 813 -3499 816 -3493
rect 820 -3499 823 -3493
rect 827 -3499 830 -3493
rect 876 -3499 879 -3493
rect 883 -3499 886 -3493
rect 890 -3499 893 -3493
rect 897 -3499 900 -3493
rect 904 -3499 907 -3493
rect 911 -3499 917 -3493
rect 918 -3499 921 -3493
rect 925 -3499 928 -3493
rect 932 -3499 935 -3493
rect 939 -3499 942 -3493
rect 946 -3499 949 -3493
rect 953 -3499 956 -3493
rect 960 -3499 963 -3493
rect 974 -3499 977 -3493
rect 995 -3499 998 -3493
rect 1002 -3499 1008 -3493
rect 1009 -3499 1012 -3493
rect 1023 -3499 1026 -3493
rect 1037 -3499 1040 -3493
rect 1044 -3499 1047 -3493
rect 1051 -3499 1054 -3493
rect 1058 -3499 1061 -3493
rect 1065 -3499 1068 -3493
rect 1072 -3499 1075 -3493
rect 1079 -3499 1082 -3493
rect 1086 -3499 1092 -3493
rect 1114 -3499 1117 -3493
rect 1121 -3499 1124 -3493
rect 1135 -3499 1138 -3493
rect 1156 -3499 1159 -3493
rect 1177 -3499 1183 -3493
rect 1184 -3499 1187 -3493
rect 1191 -3499 1194 -3493
rect 1233 -3499 1236 -3493
rect 1247 -3499 1250 -3493
rect 1268 -3499 1271 -3493
rect 1275 -3499 1278 -3493
rect 1373 -3499 1376 -3493
rect 1380 -3499 1386 -3493
rect 1387 -3499 1390 -3493
rect 1394 -3499 1397 -3493
rect 1415 -3499 1418 -3493
rect 1576 -3499 1579 -3493
rect 1 -3530 7 -3524
rect 8 -3530 14 -3524
rect 15 -3530 21 -3524
rect 22 -3530 28 -3524
rect 29 -3530 35 -3524
rect 36 -3530 42 -3524
rect 43 -3530 49 -3524
rect 50 -3530 56 -3524
rect 57 -3530 63 -3524
rect 64 -3530 70 -3524
rect 71 -3530 77 -3524
rect 78 -3530 84 -3524
rect 85 -3530 91 -3524
rect 92 -3530 98 -3524
rect 379 -3530 382 -3524
rect 386 -3530 389 -3524
rect 393 -3530 396 -3524
rect 400 -3530 403 -3524
rect 428 -3530 431 -3524
rect 442 -3530 445 -3524
rect 449 -3530 452 -3524
rect 463 -3530 466 -3524
rect 477 -3530 483 -3524
rect 484 -3530 487 -3524
rect 491 -3530 494 -3524
rect 498 -3530 501 -3524
rect 505 -3530 508 -3524
rect 512 -3530 515 -3524
rect 519 -3530 525 -3524
rect 526 -3530 529 -3524
rect 533 -3530 536 -3524
rect 540 -3530 543 -3524
rect 547 -3530 550 -3524
rect 554 -3530 560 -3524
rect 561 -3530 567 -3524
rect 568 -3530 571 -3524
rect 575 -3530 578 -3524
rect 582 -3530 585 -3524
rect 589 -3530 592 -3524
rect 596 -3530 599 -3524
rect 603 -3530 606 -3524
rect 645 -3530 648 -3524
rect 652 -3530 655 -3524
rect 673 -3530 676 -3524
rect 694 -3530 697 -3524
rect 701 -3530 704 -3524
rect 708 -3530 711 -3524
rect 729 -3530 732 -3524
rect 757 -3530 760 -3524
rect 764 -3530 767 -3524
rect 771 -3530 774 -3524
rect 778 -3530 781 -3524
rect 785 -3530 788 -3524
rect 792 -3530 795 -3524
rect 799 -3530 802 -3524
rect 806 -3530 809 -3524
rect 813 -3530 816 -3524
rect 820 -3530 826 -3524
rect 841 -3530 844 -3524
rect 862 -3530 865 -3524
rect 876 -3530 879 -3524
rect 883 -3530 886 -3524
rect 890 -3530 896 -3524
rect 897 -3530 900 -3524
rect 904 -3530 907 -3524
rect 918 -3530 921 -3524
rect 925 -3530 928 -3524
rect 932 -3530 935 -3524
rect 939 -3530 942 -3524
rect 946 -3530 952 -3524
rect 953 -3530 959 -3524
rect 960 -3530 966 -3524
rect 967 -3530 970 -3524
rect 1002 -3530 1008 -3524
rect 1016 -3530 1022 -3524
rect 1030 -3530 1036 -3524
rect 1037 -3530 1043 -3524
rect 1044 -3530 1047 -3524
rect 1051 -3530 1054 -3524
rect 1058 -3530 1064 -3524
rect 1072 -3530 1075 -3524
rect 1114 -3530 1117 -3524
rect 1128 -3530 1131 -3524
rect 1135 -3530 1138 -3524
rect 1142 -3530 1145 -3524
rect 1156 -3530 1162 -3524
rect 1163 -3530 1166 -3524
rect 1177 -3530 1180 -3524
rect 1191 -3530 1194 -3524
rect 1261 -3530 1264 -3524
rect 1275 -3530 1281 -3524
rect 1338 -3530 1341 -3524
rect 1380 -3530 1383 -3524
rect 1394 -3530 1397 -3524
rect 1499 -3530 1502 -3524
rect 1576 -3530 1582 -3524
rect 1 -3559 7 -3553
rect 8 -3559 14 -3553
rect 15 -3559 21 -3553
rect 22 -3559 28 -3553
rect 29 -3559 35 -3553
rect 36 -3559 42 -3553
rect 43 -3559 49 -3553
rect 50 -3559 56 -3553
rect 57 -3559 63 -3553
rect 64 -3559 70 -3553
rect 71 -3559 77 -3553
rect 78 -3559 84 -3553
rect 85 -3559 91 -3553
rect 92 -3559 98 -3553
rect 99 -3559 105 -3553
rect 106 -3559 112 -3553
rect 113 -3559 119 -3553
rect 379 -3559 382 -3553
rect 386 -3559 389 -3553
rect 393 -3559 396 -3553
rect 400 -3559 403 -3553
rect 407 -3559 410 -3553
rect 449 -3559 452 -3553
rect 456 -3559 459 -3553
rect 470 -3559 476 -3553
rect 477 -3559 480 -3553
rect 491 -3559 494 -3553
rect 498 -3559 504 -3553
rect 505 -3559 508 -3553
rect 512 -3559 515 -3553
rect 526 -3559 532 -3553
rect 533 -3559 536 -3553
rect 540 -3559 543 -3553
rect 547 -3559 550 -3553
rect 554 -3559 557 -3553
rect 561 -3559 567 -3553
rect 568 -3559 571 -3553
rect 575 -3559 581 -3553
rect 582 -3559 585 -3553
rect 589 -3559 592 -3553
rect 596 -3559 599 -3553
rect 603 -3559 609 -3553
rect 659 -3559 665 -3553
rect 666 -3559 669 -3553
rect 701 -3559 707 -3553
rect 708 -3559 711 -3553
rect 736 -3559 739 -3553
rect 757 -3559 760 -3553
rect 764 -3559 770 -3553
rect 771 -3559 774 -3553
rect 778 -3559 781 -3553
rect 785 -3559 788 -3553
rect 792 -3559 798 -3553
rect 799 -3559 802 -3553
rect 806 -3559 809 -3553
rect 813 -3559 816 -3553
rect 876 -3559 879 -3553
rect 883 -3559 886 -3553
rect 897 -3559 900 -3553
rect 904 -3559 907 -3553
rect 925 -3559 928 -3553
rect 932 -3559 938 -3553
rect 939 -3559 942 -3553
rect 946 -3559 952 -3553
rect 1107 -3559 1113 -3553
rect 1114 -3559 1117 -3553
rect 1128 -3559 1131 -3553
rect 1135 -3559 1138 -3553
rect 1163 -3559 1166 -3553
rect 1177 -3559 1180 -3553
rect 1191 -3559 1194 -3553
rect 1359 -3559 1362 -3553
rect 1387 -3559 1390 -3553
rect 1394 -3559 1397 -3553
rect 1 -3574 7 -3568
rect 8 -3574 14 -3568
rect 15 -3574 21 -3568
rect 22 -3574 28 -3568
rect 29 -3574 35 -3568
rect 36 -3574 42 -3568
rect 43 -3574 49 -3568
rect 50 -3574 56 -3568
rect 57 -3574 63 -3568
rect 64 -3574 70 -3568
rect 71 -3574 77 -3568
rect 78 -3574 84 -3568
rect 85 -3574 91 -3568
rect 92 -3574 98 -3568
rect 99 -3574 105 -3568
rect 386 -3574 389 -3568
rect 393 -3574 399 -3568
rect 400 -3574 406 -3568
rect 407 -3574 410 -3568
rect 456 -3574 462 -3568
rect 463 -3574 466 -3568
rect 491 -3574 494 -3568
rect 498 -3574 504 -3568
rect 561 -3574 564 -3568
rect 575 -3574 581 -3568
rect 589 -3574 592 -3568
rect 596 -3574 602 -3568
rect 631 -3574 634 -3568
rect 743 -3574 749 -3568
rect 757 -3574 760 -3568
rect 799 -3574 802 -3568
rect 806 -3574 812 -3568
rect 883 -3574 886 -3568
rect 890 -3574 896 -3568
rect 897 -3574 903 -3568
rect 1128 -3574 1134 -3568
rect 1135 -3574 1138 -3568
rect 1170 -3574 1173 -3568
rect 1177 -3574 1183 -3568
rect 1184 -3574 1187 -3568
rect 1191 -3574 1197 -3568
rect 1198 -3574 1201 -3568
rect 1387 -3574 1393 -3568
rect 1394 -3574 1397 -3568
<< polysilicon >>
rect 233 -15 234 -13
rect 233 -21 234 -19
rect 345 -15 346 -13
rect 345 -21 346 -19
rect 352 -15 353 -13
rect 359 -15 360 -13
rect 359 -21 360 -19
rect 380 -15 381 -13
rect 380 -21 381 -19
rect 401 -15 402 -13
rect 401 -21 402 -19
rect 408 -15 409 -13
rect 408 -21 409 -19
rect 415 -15 416 -13
rect 415 -21 416 -19
rect 422 -15 423 -13
rect 422 -21 423 -19
rect 432 -15 433 -13
rect 432 -21 433 -19
rect 436 -15 437 -13
rect 436 -21 437 -19
rect 443 -15 444 -13
rect 443 -21 444 -19
rect 450 -15 451 -13
rect 453 -15 454 -13
rect 457 -15 458 -13
rect 460 -15 461 -13
rect 460 -21 461 -19
rect 467 -15 468 -13
rect 464 -21 465 -19
rect 471 -15 472 -13
rect 471 -21 472 -19
rect 506 -15 507 -13
rect 509 -21 510 -19
rect 527 -15 528 -13
rect 527 -21 528 -19
rect 534 -15 535 -13
rect 534 -21 535 -19
rect 537 -21 538 -19
rect 548 -15 549 -13
rect 551 -21 552 -19
rect 555 -15 556 -13
rect 555 -21 556 -19
rect 604 -15 605 -13
rect 604 -21 605 -19
rect 614 -15 615 -13
rect 653 -15 654 -13
rect 653 -21 654 -19
rect 670 -15 671 -13
rect 670 -21 671 -19
rect 677 -15 678 -13
rect 677 -21 678 -19
rect 688 -15 689 -13
rect 688 -21 689 -19
rect 716 -15 717 -13
rect 719 -21 720 -19
rect 754 -15 755 -13
rect 751 -21 752 -19
rect 754 -21 755 -19
rect 800 -15 801 -13
rect 800 -21 801 -19
rect 877 -15 878 -13
rect 880 -21 881 -19
rect 954 -15 955 -13
rect 954 -21 955 -19
rect 145 -52 146 -50
rect 149 -52 150 -50
rect 149 -58 150 -56
rect 156 -52 157 -50
rect 156 -58 157 -56
rect 226 -52 227 -50
rect 226 -58 227 -56
rect 236 -52 237 -50
rect 261 -52 262 -50
rect 261 -58 262 -56
rect 282 -52 283 -50
rect 282 -58 283 -56
rect 306 -52 307 -50
rect 306 -58 307 -56
rect 324 -52 325 -50
rect 324 -58 325 -56
rect 331 -52 332 -50
rect 331 -58 332 -56
rect 338 -52 339 -50
rect 338 -58 339 -56
rect 373 -52 374 -50
rect 373 -58 374 -56
rect 380 -52 381 -50
rect 380 -58 381 -56
rect 390 -52 391 -50
rect 387 -58 388 -56
rect 394 -52 395 -50
rect 394 -58 395 -56
rect 401 -52 402 -50
rect 401 -58 402 -56
rect 408 -52 409 -50
rect 408 -58 409 -56
rect 415 -58 416 -56
rect 425 -52 426 -50
rect 422 -58 423 -56
rect 429 -52 430 -50
rect 429 -58 430 -56
rect 436 -52 437 -50
rect 436 -58 437 -56
rect 443 -52 444 -50
rect 450 -52 451 -50
rect 450 -58 451 -56
rect 460 -52 461 -50
rect 457 -58 458 -56
rect 460 -58 461 -56
rect 464 -52 465 -50
rect 464 -58 465 -56
rect 471 -52 472 -50
rect 471 -58 472 -56
rect 478 -52 479 -50
rect 478 -58 479 -56
rect 492 -52 493 -50
rect 495 -52 496 -50
rect 499 -52 500 -50
rect 499 -58 500 -56
rect 506 -52 507 -50
rect 506 -58 507 -56
rect 513 -52 514 -50
rect 516 -52 517 -50
rect 516 -58 517 -56
rect 520 -52 521 -50
rect 523 -52 524 -50
rect 523 -58 524 -56
rect 527 -52 528 -50
rect 530 -52 531 -50
rect 534 -52 535 -50
rect 534 -58 535 -56
rect 541 -52 542 -50
rect 541 -58 542 -56
rect 548 -52 549 -50
rect 548 -58 549 -56
rect 555 -52 556 -50
rect 555 -58 556 -56
rect 562 -52 563 -50
rect 562 -58 563 -56
rect 569 -58 570 -56
rect 576 -52 577 -50
rect 576 -58 577 -56
rect 583 -52 584 -50
rect 583 -58 584 -56
rect 590 -52 591 -50
rect 590 -58 591 -56
rect 593 -58 594 -56
rect 597 -52 598 -50
rect 597 -58 598 -56
rect 604 -52 605 -50
rect 604 -58 605 -56
rect 611 -52 612 -50
rect 611 -58 612 -56
rect 618 -52 619 -50
rect 618 -58 619 -56
rect 625 -52 626 -50
rect 625 -58 626 -56
rect 632 -52 633 -50
rect 639 -52 640 -50
rect 639 -58 640 -56
rect 646 -52 647 -50
rect 646 -58 647 -56
rect 653 -52 654 -50
rect 653 -58 654 -56
rect 660 -52 661 -50
rect 660 -58 661 -56
rect 667 -52 668 -50
rect 667 -58 668 -56
rect 677 -52 678 -50
rect 677 -58 678 -56
rect 681 -52 682 -50
rect 681 -58 682 -56
rect 688 -52 689 -50
rect 688 -58 689 -56
rect 702 -52 703 -50
rect 702 -58 703 -56
rect 712 -52 713 -50
rect 709 -58 710 -56
rect 712 -58 713 -56
rect 716 -52 717 -50
rect 716 -58 717 -56
rect 730 -52 731 -50
rect 730 -58 731 -56
rect 744 -52 745 -50
rect 744 -58 745 -56
rect 758 -52 759 -50
rect 758 -58 759 -56
rect 772 -52 773 -50
rect 772 -58 773 -56
rect 814 -52 815 -50
rect 814 -58 815 -56
rect 821 -52 822 -50
rect 821 -58 822 -56
rect 828 -52 829 -50
rect 828 -58 829 -56
rect 842 -52 843 -50
rect 842 -58 843 -56
rect 884 -52 885 -50
rect 884 -58 885 -56
rect 898 -52 899 -50
rect 898 -58 899 -56
rect 936 -58 937 -56
rect 989 -52 990 -50
rect 989 -58 990 -56
rect 996 -52 997 -50
rect 996 -58 997 -56
rect 89 -105 90 -103
rect 128 -99 129 -97
rect 128 -105 129 -103
rect 149 -99 150 -97
rect 149 -105 150 -103
rect 191 -99 192 -97
rect 191 -105 192 -103
rect 198 -99 199 -97
rect 205 -99 206 -97
rect 205 -105 206 -103
rect 219 -99 220 -97
rect 219 -105 220 -103
rect 247 -99 248 -97
rect 247 -105 248 -103
rect 250 -105 251 -103
rect 254 -99 255 -97
rect 254 -105 255 -103
rect 261 -99 262 -97
rect 261 -105 262 -103
rect 268 -99 269 -97
rect 268 -105 269 -103
rect 275 -99 276 -97
rect 275 -105 276 -103
rect 282 -99 283 -97
rect 282 -105 283 -103
rect 289 -99 290 -97
rect 292 -105 293 -103
rect 296 -99 297 -97
rect 296 -105 297 -103
rect 303 -99 304 -97
rect 303 -105 304 -103
rect 310 -99 311 -97
rect 310 -105 311 -103
rect 317 -99 318 -97
rect 317 -105 318 -103
rect 324 -99 325 -97
rect 324 -105 325 -103
rect 331 -99 332 -97
rect 334 -99 335 -97
rect 331 -105 332 -103
rect 338 -99 339 -97
rect 338 -105 339 -103
rect 345 -99 346 -97
rect 345 -105 346 -103
rect 352 -99 353 -97
rect 352 -105 353 -103
rect 359 -99 360 -97
rect 359 -105 360 -103
rect 366 -99 367 -97
rect 366 -105 367 -103
rect 373 -99 374 -97
rect 376 -99 377 -97
rect 373 -105 374 -103
rect 376 -105 377 -103
rect 380 -99 381 -97
rect 380 -105 381 -103
rect 387 -99 388 -97
rect 387 -105 388 -103
rect 394 -99 395 -97
rect 394 -105 395 -103
rect 401 -99 402 -97
rect 401 -105 402 -103
rect 411 -99 412 -97
rect 408 -105 409 -103
rect 415 -99 416 -97
rect 415 -105 416 -103
rect 422 -99 423 -97
rect 422 -105 423 -103
rect 432 -99 433 -97
rect 432 -105 433 -103
rect 436 -99 437 -97
rect 436 -105 437 -103
rect 443 -99 444 -97
rect 443 -105 444 -103
rect 450 -99 451 -97
rect 450 -105 451 -103
rect 457 -105 458 -103
rect 460 -105 461 -103
rect 464 -99 465 -97
rect 464 -105 465 -103
rect 474 -99 475 -97
rect 471 -105 472 -103
rect 474 -105 475 -103
rect 478 -99 479 -97
rect 478 -105 479 -103
rect 488 -99 489 -97
rect 485 -105 486 -103
rect 488 -105 489 -103
rect 492 -99 493 -97
rect 492 -105 493 -103
rect 499 -99 500 -97
rect 499 -105 500 -103
rect 506 -99 507 -97
rect 506 -105 507 -103
rect 513 -99 514 -97
rect 513 -105 514 -103
rect 520 -99 521 -97
rect 520 -105 521 -103
rect 530 -99 531 -97
rect 527 -105 528 -103
rect 530 -105 531 -103
rect 534 -99 535 -97
rect 534 -105 535 -103
rect 537 -105 538 -103
rect 541 -99 542 -97
rect 541 -105 542 -103
rect 551 -99 552 -97
rect 548 -105 549 -103
rect 551 -105 552 -103
rect 555 -99 556 -97
rect 555 -105 556 -103
rect 562 -99 563 -97
rect 562 -105 563 -103
rect 569 -99 570 -97
rect 569 -105 570 -103
rect 576 -99 577 -97
rect 576 -105 577 -103
rect 583 -99 584 -97
rect 583 -105 584 -103
rect 590 -99 591 -97
rect 590 -105 591 -103
rect 597 -99 598 -97
rect 597 -105 598 -103
rect 604 -99 605 -97
rect 604 -105 605 -103
rect 611 -99 612 -97
rect 611 -105 612 -103
rect 618 -99 619 -97
rect 618 -105 619 -103
rect 625 -99 626 -97
rect 625 -105 626 -103
rect 632 -99 633 -97
rect 632 -105 633 -103
rect 639 -99 640 -97
rect 639 -105 640 -103
rect 649 -99 650 -97
rect 646 -105 647 -103
rect 649 -105 650 -103
rect 653 -99 654 -97
rect 653 -105 654 -103
rect 660 -99 661 -97
rect 660 -105 661 -103
rect 667 -99 668 -97
rect 667 -105 668 -103
rect 674 -99 675 -97
rect 674 -105 675 -103
rect 681 -99 682 -97
rect 681 -105 682 -103
rect 688 -99 689 -97
rect 688 -105 689 -103
rect 695 -99 696 -97
rect 695 -105 696 -103
rect 702 -99 703 -97
rect 702 -105 703 -103
rect 709 -99 710 -97
rect 709 -105 710 -103
rect 716 -99 717 -97
rect 716 -105 717 -103
rect 723 -99 724 -97
rect 723 -105 724 -103
rect 730 -99 731 -97
rect 730 -105 731 -103
rect 737 -99 738 -97
rect 737 -105 738 -103
rect 744 -99 745 -97
rect 744 -105 745 -103
rect 751 -99 752 -97
rect 751 -105 752 -103
rect 779 -99 780 -97
rect 779 -105 780 -103
rect 786 -99 787 -97
rect 786 -105 787 -103
rect 793 -99 794 -97
rect 796 -99 797 -97
rect 793 -105 794 -103
rect 796 -105 797 -103
rect 800 -99 801 -97
rect 800 -105 801 -103
rect 807 -99 808 -97
rect 810 -99 811 -97
rect 810 -105 811 -103
rect 817 -99 818 -97
rect 814 -105 815 -103
rect 817 -105 818 -103
rect 821 -99 822 -97
rect 824 -105 825 -103
rect 828 -99 829 -97
rect 828 -105 829 -103
rect 835 -99 836 -97
rect 835 -105 836 -103
rect 842 -99 843 -97
rect 842 -105 843 -103
rect 856 -99 857 -97
rect 856 -105 857 -103
rect 863 -99 864 -97
rect 863 -105 864 -103
rect 870 -99 871 -97
rect 870 -105 871 -103
rect 884 -99 885 -97
rect 887 -99 888 -97
rect 884 -105 885 -103
rect 891 -99 892 -97
rect 891 -105 892 -103
rect 940 -99 941 -97
rect 940 -105 941 -103
rect 947 -99 948 -97
rect 947 -105 948 -103
rect 954 -99 955 -97
rect 954 -105 955 -103
rect 1010 -99 1011 -97
rect 1010 -105 1011 -103
rect 1087 -99 1088 -97
rect 1087 -105 1088 -103
rect 93 -168 94 -166
rect 93 -174 94 -172
rect 114 -168 115 -166
rect 114 -174 115 -172
rect 135 -168 136 -166
rect 135 -174 136 -172
rect 142 -168 143 -166
rect 142 -174 143 -172
rect 149 -168 150 -166
rect 149 -174 150 -172
rect 156 -168 157 -166
rect 156 -174 157 -172
rect 163 -168 164 -166
rect 163 -174 164 -172
rect 170 -168 171 -166
rect 170 -174 171 -172
rect 177 -168 178 -166
rect 177 -174 178 -172
rect 184 -168 185 -166
rect 184 -174 185 -172
rect 191 -168 192 -166
rect 191 -174 192 -172
rect 198 -168 199 -166
rect 198 -174 199 -172
rect 208 -168 209 -166
rect 208 -174 209 -172
rect 215 -174 216 -172
rect 219 -168 220 -166
rect 219 -174 220 -172
rect 226 -168 227 -166
rect 226 -174 227 -172
rect 233 -174 234 -172
rect 236 -174 237 -172
rect 243 -168 244 -166
rect 240 -174 241 -172
rect 243 -174 244 -172
rect 247 -168 248 -166
rect 247 -174 248 -172
rect 254 -168 255 -166
rect 254 -174 255 -172
rect 261 -168 262 -166
rect 261 -174 262 -172
rect 268 -168 269 -166
rect 268 -174 269 -172
rect 275 -168 276 -166
rect 275 -174 276 -172
rect 282 -168 283 -166
rect 282 -174 283 -172
rect 289 -168 290 -166
rect 289 -174 290 -172
rect 296 -168 297 -166
rect 296 -174 297 -172
rect 303 -168 304 -166
rect 303 -174 304 -172
rect 310 -168 311 -166
rect 310 -174 311 -172
rect 317 -168 318 -166
rect 317 -174 318 -172
rect 324 -168 325 -166
rect 324 -174 325 -172
rect 331 -168 332 -166
rect 331 -174 332 -172
rect 338 -168 339 -166
rect 338 -174 339 -172
rect 345 -168 346 -166
rect 345 -174 346 -172
rect 352 -168 353 -166
rect 355 -168 356 -166
rect 352 -174 353 -172
rect 359 -168 360 -166
rect 362 -168 363 -166
rect 359 -174 360 -172
rect 362 -174 363 -172
rect 366 -168 367 -166
rect 366 -174 367 -172
rect 373 -168 374 -166
rect 373 -174 374 -172
rect 380 -168 381 -166
rect 380 -174 381 -172
rect 387 -168 388 -166
rect 387 -174 388 -172
rect 394 -168 395 -166
rect 394 -174 395 -172
rect 401 -168 402 -166
rect 401 -174 402 -172
rect 408 -168 409 -166
rect 408 -174 409 -172
rect 415 -168 416 -166
rect 415 -174 416 -172
rect 422 -168 423 -166
rect 422 -174 423 -172
rect 429 -168 430 -166
rect 432 -168 433 -166
rect 432 -174 433 -172
rect 436 -168 437 -166
rect 436 -174 437 -172
rect 443 -168 444 -166
rect 443 -174 444 -172
rect 450 -168 451 -166
rect 450 -174 451 -172
rect 457 -168 458 -166
rect 457 -174 458 -172
rect 464 -168 465 -166
rect 467 -168 468 -166
rect 464 -174 465 -172
rect 471 -168 472 -166
rect 471 -174 472 -172
rect 478 -168 479 -166
rect 481 -168 482 -166
rect 481 -174 482 -172
rect 485 -168 486 -166
rect 485 -174 486 -172
rect 492 -168 493 -166
rect 492 -174 493 -172
rect 499 -168 500 -166
rect 502 -168 503 -166
rect 499 -174 500 -172
rect 502 -174 503 -172
rect 506 -168 507 -166
rect 509 -168 510 -166
rect 509 -174 510 -172
rect 513 -168 514 -166
rect 513 -174 514 -172
rect 516 -174 517 -172
rect 520 -168 521 -166
rect 520 -174 521 -172
rect 523 -174 524 -172
rect 527 -168 528 -166
rect 527 -174 528 -172
rect 534 -168 535 -166
rect 534 -174 535 -172
rect 541 -168 542 -166
rect 541 -174 542 -172
rect 544 -174 545 -172
rect 548 -168 549 -166
rect 548 -174 549 -172
rect 555 -168 556 -166
rect 555 -174 556 -172
rect 562 -168 563 -166
rect 562 -174 563 -172
rect 569 -168 570 -166
rect 569 -174 570 -172
rect 576 -168 577 -166
rect 576 -174 577 -172
rect 583 -168 584 -166
rect 583 -174 584 -172
rect 590 -168 591 -166
rect 590 -174 591 -172
rect 597 -168 598 -166
rect 597 -174 598 -172
rect 604 -168 605 -166
rect 604 -174 605 -172
rect 611 -168 612 -166
rect 611 -174 612 -172
rect 614 -174 615 -172
rect 618 -168 619 -166
rect 618 -174 619 -172
rect 625 -168 626 -166
rect 625 -174 626 -172
rect 632 -168 633 -166
rect 632 -174 633 -172
rect 639 -168 640 -166
rect 639 -174 640 -172
rect 646 -168 647 -166
rect 646 -174 647 -172
rect 653 -168 654 -166
rect 656 -168 657 -166
rect 653 -174 654 -172
rect 656 -174 657 -172
rect 660 -168 661 -166
rect 660 -174 661 -172
rect 667 -168 668 -166
rect 667 -174 668 -172
rect 674 -168 675 -166
rect 674 -174 675 -172
rect 681 -168 682 -166
rect 681 -174 682 -172
rect 688 -168 689 -166
rect 688 -174 689 -172
rect 698 -168 699 -166
rect 695 -174 696 -172
rect 698 -174 699 -172
rect 702 -168 703 -166
rect 702 -174 703 -172
rect 709 -168 710 -166
rect 709 -174 710 -172
rect 716 -168 717 -166
rect 716 -174 717 -172
rect 723 -168 724 -166
rect 723 -174 724 -172
rect 730 -168 731 -166
rect 730 -174 731 -172
rect 737 -168 738 -166
rect 737 -174 738 -172
rect 744 -168 745 -166
rect 744 -174 745 -172
rect 751 -168 752 -166
rect 751 -174 752 -172
rect 758 -168 759 -166
rect 758 -174 759 -172
rect 768 -168 769 -166
rect 765 -174 766 -172
rect 768 -174 769 -172
rect 772 -168 773 -166
rect 772 -174 773 -172
rect 779 -168 780 -166
rect 779 -174 780 -172
rect 786 -168 787 -166
rect 786 -174 787 -172
rect 793 -168 794 -166
rect 793 -174 794 -172
rect 796 -174 797 -172
rect 800 -168 801 -166
rect 800 -174 801 -172
rect 807 -168 808 -166
rect 807 -174 808 -172
rect 814 -168 815 -166
rect 814 -174 815 -172
rect 821 -168 822 -166
rect 828 -168 829 -166
rect 828 -174 829 -172
rect 835 -168 836 -166
rect 835 -174 836 -172
rect 842 -168 843 -166
rect 842 -174 843 -172
rect 849 -168 850 -166
rect 849 -174 850 -172
rect 856 -168 857 -166
rect 856 -174 857 -172
rect 863 -168 864 -166
rect 863 -174 864 -172
rect 870 -168 871 -166
rect 870 -174 871 -172
rect 877 -168 878 -166
rect 880 -168 881 -166
rect 880 -174 881 -172
rect 887 -168 888 -166
rect 887 -174 888 -172
rect 891 -168 892 -166
rect 891 -174 892 -172
rect 898 -168 899 -166
rect 898 -174 899 -172
rect 905 -168 906 -166
rect 905 -174 906 -172
rect 912 -168 913 -166
rect 912 -174 913 -172
rect 919 -168 920 -166
rect 919 -174 920 -172
rect 926 -168 927 -166
rect 926 -174 927 -172
rect 933 -168 934 -166
rect 933 -174 934 -172
rect 940 -168 941 -166
rect 940 -174 941 -172
rect 947 -168 948 -166
rect 947 -174 948 -172
rect 954 -168 955 -166
rect 954 -174 955 -172
rect 961 -168 962 -166
rect 961 -174 962 -172
rect 968 -168 969 -166
rect 968 -174 969 -172
rect 975 -168 976 -166
rect 975 -174 976 -172
rect 982 -168 983 -166
rect 982 -174 983 -172
rect 996 -168 997 -166
rect 996 -174 997 -172
rect 1010 -168 1011 -166
rect 1010 -174 1011 -172
rect 1038 -168 1039 -166
rect 1038 -174 1039 -172
rect 1129 -168 1130 -166
rect 1129 -174 1130 -172
rect 1136 -168 1137 -166
rect 1136 -174 1137 -172
rect 1195 -168 1196 -166
rect 1195 -174 1196 -172
rect 1220 -168 1221 -166
rect 1220 -174 1221 -172
rect 51 -255 52 -253
rect 51 -261 52 -259
rect 58 -255 59 -253
rect 58 -261 59 -259
rect 65 -255 66 -253
rect 65 -261 66 -259
rect 72 -255 73 -253
rect 72 -261 73 -259
rect 79 -255 80 -253
rect 79 -261 80 -259
rect 86 -255 87 -253
rect 86 -261 87 -259
rect 93 -255 94 -253
rect 93 -261 94 -259
rect 100 -255 101 -253
rect 100 -261 101 -259
rect 107 -255 108 -253
rect 107 -261 108 -259
rect 117 -255 118 -253
rect 117 -261 118 -259
rect 121 -255 122 -253
rect 121 -261 122 -259
rect 128 -255 129 -253
rect 128 -261 129 -259
rect 135 -255 136 -253
rect 135 -261 136 -259
rect 142 -255 143 -253
rect 142 -261 143 -259
rect 149 -255 150 -253
rect 149 -261 150 -259
rect 156 -255 157 -253
rect 156 -261 157 -259
rect 163 -255 164 -253
rect 163 -261 164 -259
rect 170 -255 171 -253
rect 173 -261 174 -259
rect 177 -255 178 -253
rect 177 -261 178 -259
rect 184 -255 185 -253
rect 184 -261 185 -259
rect 191 -255 192 -253
rect 191 -261 192 -259
rect 194 -261 195 -259
rect 201 -255 202 -253
rect 198 -261 199 -259
rect 205 -255 206 -253
rect 205 -261 206 -259
rect 212 -255 213 -253
rect 215 -261 216 -259
rect 219 -255 220 -253
rect 219 -261 220 -259
rect 226 -255 227 -253
rect 226 -261 227 -259
rect 233 -255 234 -253
rect 236 -255 237 -253
rect 233 -261 234 -259
rect 236 -261 237 -259
rect 243 -255 244 -253
rect 243 -261 244 -259
rect 247 -255 248 -253
rect 247 -261 248 -259
rect 254 -255 255 -253
rect 254 -261 255 -259
rect 261 -255 262 -253
rect 261 -261 262 -259
rect 268 -255 269 -253
rect 268 -261 269 -259
rect 275 -255 276 -253
rect 275 -261 276 -259
rect 282 -255 283 -253
rect 282 -261 283 -259
rect 289 -255 290 -253
rect 292 -255 293 -253
rect 289 -261 290 -259
rect 296 -255 297 -253
rect 296 -261 297 -259
rect 303 -255 304 -253
rect 303 -261 304 -259
rect 310 -255 311 -253
rect 310 -261 311 -259
rect 317 -255 318 -253
rect 317 -261 318 -259
rect 324 -255 325 -253
rect 324 -261 325 -259
rect 331 -255 332 -253
rect 331 -261 332 -259
rect 338 -255 339 -253
rect 338 -261 339 -259
rect 345 -255 346 -253
rect 345 -261 346 -259
rect 352 -255 353 -253
rect 352 -261 353 -259
rect 359 -255 360 -253
rect 359 -261 360 -259
rect 366 -255 367 -253
rect 366 -261 367 -259
rect 373 -255 374 -253
rect 373 -261 374 -259
rect 380 -255 381 -253
rect 383 -255 384 -253
rect 383 -261 384 -259
rect 387 -255 388 -253
rect 387 -261 388 -259
rect 394 -255 395 -253
rect 394 -261 395 -259
rect 401 -255 402 -253
rect 401 -261 402 -259
rect 408 -255 409 -253
rect 408 -261 409 -259
rect 415 -255 416 -253
rect 415 -261 416 -259
rect 422 -255 423 -253
rect 422 -261 423 -259
rect 429 -255 430 -253
rect 429 -261 430 -259
rect 436 -255 437 -253
rect 436 -261 437 -259
rect 443 -255 444 -253
rect 446 -255 447 -253
rect 443 -261 444 -259
rect 450 -255 451 -253
rect 450 -261 451 -259
rect 457 -255 458 -253
rect 460 -255 461 -253
rect 457 -261 458 -259
rect 460 -261 461 -259
rect 467 -255 468 -253
rect 467 -261 468 -259
rect 471 -255 472 -253
rect 474 -255 475 -253
rect 471 -261 472 -259
rect 474 -261 475 -259
rect 478 -255 479 -253
rect 478 -261 479 -259
rect 485 -255 486 -253
rect 485 -261 486 -259
rect 495 -255 496 -253
rect 492 -261 493 -259
rect 495 -261 496 -259
rect 499 -255 500 -253
rect 499 -261 500 -259
rect 506 -255 507 -253
rect 509 -255 510 -253
rect 506 -261 507 -259
rect 509 -261 510 -259
rect 513 -255 514 -253
rect 513 -261 514 -259
rect 520 -255 521 -253
rect 520 -261 521 -259
rect 530 -255 531 -253
rect 527 -261 528 -259
rect 530 -261 531 -259
rect 534 -255 535 -253
rect 534 -261 535 -259
rect 541 -255 542 -253
rect 544 -255 545 -253
rect 544 -261 545 -259
rect 548 -255 549 -253
rect 548 -261 549 -259
rect 555 -255 556 -253
rect 555 -261 556 -259
rect 562 -255 563 -253
rect 562 -261 563 -259
rect 569 -255 570 -253
rect 572 -255 573 -253
rect 569 -261 570 -259
rect 572 -261 573 -259
rect 579 -255 580 -253
rect 576 -261 577 -259
rect 579 -261 580 -259
rect 583 -255 584 -253
rect 583 -261 584 -259
rect 590 -255 591 -253
rect 593 -255 594 -253
rect 593 -261 594 -259
rect 597 -255 598 -253
rect 597 -261 598 -259
rect 604 -255 605 -253
rect 604 -261 605 -259
rect 611 -255 612 -253
rect 614 -255 615 -253
rect 611 -261 612 -259
rect 614 -261 615 -259
rect 618 -255 619 -253
rect 618 -261 619 -259
rect 625 -255 626 -253
rect 625 -261 626 -259
rect 632 -255 633 -253
rect 632 -261 633 -259
rect 639 -255 640 -253
rect 639 -261 640 -259
rect 646 -255 647 -253
rect 646 -261 647 -259
rect 653 -255 654 -253
rect 653 -261 654 -259
rect 660 -255 661 -253
rect 660 -261 661 -259
rect 667 -255 668 -253
rect 667 -261 668 -259
rect 674 -255 675 -253
rect 674 -261 675 -259
rect 681 -255 682 -253
rect 681 -261 682 -259
rect 688 -255 689 -253
rect 688 -261 689 -259
rect 695 -255 696 -253
rect 695 -261 696 -259
rect 702 -255 703 -253
rect 702 -261 703 -259
rect 709 -255 710 -253
rect 709 -261 710 -259
rect 719 -255 720 -253
rect 716 -261 717 -259
rect 723 -255 724 -253
rect 723 -261 724 -259
rect 730 -255 731 -253
rect 730 -261 731 -259
rect 737 -255 738 -253
rect 737 -261 738 -259
rect 744 -255 745 -253
rect 744 -261 745 -259
rect 751 -255 752 -253
rect 751 -261 752 -259
rect 758 -255 759 -253
rect 758 -261 759 -259
rect 765 -255 766 -253
rect 765 -261 766 -259
rect 772 -255 773 -253
rect 779 -255 780 -253
rect 779 -261 780 -259
rect 789 -255 790 -253
rect 786 -261 787 -259
rect 789 -261 790 -259
rect 793 -255 794 -253
rect 793 -261 794 -259
rect 800 -255 801 -253
rect 800 -261 801 -259
rect 807 -255 808 -253
rect 807 -261 808 -259
rect 814 -255 815 -253
rect 814 -261 815 -259
rect 821 -255 822 -253
rect 821 -261 822 -259
rect 831 -255 832 -253
rect 828 -261 829 -259
rect 835 -255 836 -253
rect 835 -261 836 -259
rect 842 -255 843 -253
rect 842 -261 843 -259
rect 849 -255 850 -253
rect 849 -261 850 -259
rect 856 -255 857 -253
rect 856 -261 857 -259
rect 863 -255 864 -253
rect 863 -261 864 -259
rect 870 -255 871 -253
rect 870 -261 871 -259
rect 877 -255 878 -253
rect 877 -261 878 -259
rect 884 -255 885 -253
rect 884 -261 885 -259
rect 891 -255 892 -253
rect 891 -261 892 -259
rect 898 -255 899 -253
rect 898 -261 899 -259
rect 905 -255 906 -253
rect 905 -261 906 -259
rect 912 -255 913 -253
rect 912 -261 913 -259
rect 919 -255 920 -253
rect 919 -261 920 -259
rect 926 -255 927 -253
rect 926 -261 927 -259
rect 933 -255 934 -253
rect 933 -261 934 -259
rect 940 -255 941 -253
rect 940 -261 941 -259
rect 947 -255 948 -253
rect 947 -261 948 -259
rect 954 -255 955 -253
rect 954 -261 955 -259
rect 961 -255 962 -253
rect 961 -261 962 -259
rect 968 -255 969 -253
rect 968 -261 969 -259
rect 975 -255 976 -253
rect 975 -261 976 -259
rect 982 -255 983 -253
rect 982 -261 983 -259
rect 989 -255 990 -253
rect 989 -261 990 -259
rect 996 -255 997 -253
rect 999 -255 1000 -253
rect 999 -261 1000 -259
rect 1003 -255 1004 -253
rect 1003 -261 1004 -259
rect 1010 -255 1011 -253
rect 1010 -261 1011 -259
rect 1017 -255 1018 -253
rect 1017 -261 1018 -259
rect 1024 -255 1025 -253
rect 1024 -261 1025 -259
rect 1031 -255 1032 -253
rect 1031 -261 1032 -259
rect 1038 -255 1039 -253
rect 1038 -261 1039 -259
rect 1045 -255 1046 -253
rect 1045 -261 1046 -259
rect 1052 -255 1053 -253
rect 1052 -261 1053 -259
rect 1059 -255 1060 -253
rect 1059 -261 1060 -259
rect 1066 -255 1067 -253
rect 1066 -261 1067 -259
rect 1073 -255 1074 -253
rect 1073 -261 1074 -259
rect 1080 -255 1081 -253
rect 1080 -261 1081 -259
rect 1087 -255 1088 -253
rect 1087 -261 1088 -259
rect 1097 -255 1098 -253
rect 1094 -261 1095 -259
rect 1097 -261 1098 -259
rect 1101 -255 1102 -253
rect 1101 -261 1102 -259
rect 1108 -255 1109 -253
rect 1108 -261 1109 -259
rect 1118 -255 1119 -253
rect 1115 -261 1116 -259
rect 1118 -261 1119 -259
rect 1125 -255 1126 -253
rect 1122 -261 1123 -259
rect 1129 -255 1130 -253
rect 1129 -261 1130 -259
rect 1136 -255 1137 -253
rect 1136 -261 1137 -259
rect 1143 -255 1144 -253
rect 1143 -261 1144 -259
rect 1150 -255 1151 -253
rect 1150 -261 1151 -259
rect 1157 -255 1158 -253
rect 1157 -261 1158 -259
rect 1164 -255 1165 -253
rect 1164 -261 1165 -259
rect 1171 -255 1172 -253
rect 1171 -261 1172 -259
rect 1227 -255 1228 -253
rect 1227 -261 1228 -259
rect 1255 -255 1256 -253
rect 1255 -261 1256 -259
rect 1283 -255 1284 -253
rect 1283 -261 1284 -259
rect 44 -386 45 -384
rect 44 -392 45 -390
rect 51 -386 52 -384
rect 51 -392 52 -390
rect 58 -386 59 -384
rect 61 -386 62 -384
rect 65 -386 66 -384
rect 65 -392 66 -390
rect 72 -386 73 -384
rect 72 -392 73 -390
rect 79 -386 80 -384
rect 79 -392 80 -390
rect 86 -386 87 -384
rect 86 -392 87 -390
rect 93 -386 94 -384
rect 96 -386 97 -384
rect 96 -392 97 -390
rect 100 -386 101 -384
rect 100 -392 101 -390
rect 107 -386 108 -384
rect 107 -392 108 -390
rect 114 -386 115 -384
rect 117 -386 118 -384
rect 117 -392 118 -390
rect 121 -386 122 -384
rect 121 -392 122 -390
rect 124 -392 125 -390
rect 128 -386 129 -384
rect 128 -392 129 -390
rect 138 -386 139 -384
rect 135 -392 136 -390
rect 138 -392 139 -390
rect 142 -386 143 -384
rect 142 -392 143 -390
rect 149 -386 150 -384
rect 149 -392 150 -390
rect 156 -386 157 -384
rect 156 -392 157 -390
rect 163 -386 164 -384
rect 163 -392 164 -390
rect 170 -386 171 -384
rect 170 -392 171 -390
rect 177 -386 178 -384
rect 177 -392 178 -390
rect 184 -386 185 -384
rect 184 -392 185 -390
rect 191 -386 192 -384
rect 191 -392 192 -390
rect 198 -386 199 -384
rect 201 -386 202 -384
rect 198 -392 199 -390
rect 205 -386 206 -384
rect 208 -386 209 -384
rect 205 -392 206 -390
rect 212 -392 213 -390
rect 215 -392 216 -390
rect 219 -386 220 -384
rect 219 -392 220 -390
rect 226 -386 227 -384
rect 226 -392 227 -390
rect 240 -386 241 -384
rect 240 -392 241 -390
rect 254 -386 255 -384
rect 254 -392 255 -390
rect 261 -386 262 -384
rect 261 -392 262 -390
rect 268 -386 269 -384
rect 268 -392 269 -390
rect 275 -386 276 -384
rect 275 -392 276 -390
rect 282 -386 283 -384
rect 285 -386 286 -384
rect 282 -392 283 -390
rect 285 -392 286 -390
rect 289 -386 290 -384
rect 289 -392 290 -390
rect 296 -386 297 -384
rect 296 -392 297 -390
rect 303 -386 304 -384
rect 303 -392 304 -390
rect 310 -386 311 -384
rect 310 -392 311 -390
rect 320 -392 321 -390
rect 324 -386 325 -384
rect 324 -392 325 -390
rect 331 -386 332 -384
rect 331 -392 332 -390
rect 338 -386 339 -384
rect 341 -386 342 -384
rect 338 -392 339 -390
rect 345 -386 346 -384
rect 345 -392 346 -390
rect 352 -386 353 -384
rect 352 -392 353 -390
rect 359 -386 360 -384
rect 359 -392 360 -390
rect 366 -386 367 -384
rect 366 -392 367 -390
rect 373 -386 374 -384
rect 373 -392 374 -390
rect 380 -386 381 -384
rect 380 -392 381 -390
rect 387 -386 388 -384
rect 387 -392 388 -390
rect 394 -386 395 -384
rect 394 -392 395 -390
rect 401 -386 402 -384
rect 401 -392 402 -390
rect 408 -386 409 -384
rect 411 -386 412 -384
rect 408 -392 409 -390
rect 415 -386 416 -384
rect 415 -392 416 -390
rect 422 -386 423 -384
rect 422 -392 423 -390
rect 429 -386 430 -384
rect 429 -392 430 -390
rect 436 -386 437 -384
rect 439 -386 440 -384
rect 436 -392 437 -390
rect 439 -392 440 -390
rect 443 -386 444 -384
rect 443 -392 444 -390
rect 450 -386 451 -384
rect 453 -386 454 -384
rect 450 -392 451 -390
rect 457 -386 458 -384
rect 457 -392 458 -390
rect 464 -386 465 -384
rect 464 -392 465 -390
rect 471 -386 472 -384
rect 474 -386 475 -384
rect 474 -392 475 -390
rect 478 -386 479 -384
rect 478 -392 479 -390
rect 485 -386 486 -384
rect 485 -392 486 -390
rect 492 -386 493 -384
rect 492 -392 493 -390
rect 499 -386 500 -384
rect 499 -392 500 -390
rect 506 -386 507 -384
rect 509 -386 510 -384
rect 506 -392 507 -390
rect 509 -392 510 -390
rect 513 -386 514 -384
rect 513 -392 514 -390
rect 520 -386 521 -384
rect 520 -392 521 -390
rect 527 -386 528 -384
rect 527 -392 528 -390
rect 534 -386 535 -384
rect 534 -392 535 -390
rect 541 -386 542 -384
rect 541 -392 542 -390
rect 548 -386 549 -384
rect 548 -392 549 -390
rect 555 -386 556 -384
rect 555 -392 556 -390
rect 562 -386 563 -384
rect 562 -392 563 -390
rect 569 -386 570 -384
rect 569 -392 570 -390
rect 576 -386 577 -384
rect 576 -392 577 -390
rect 583 -386 584 -384
rect 583 -392 584 -390
rect 590 -386 591 -384
rect 590 -392 591 -390
rect 597 -386 598 -384
rect 597 -392 598 -390
rect 604 -386 605 -384
rect 607 -386 608 -384
rect 604 -392 605 -390
rect 607 -392 608 -390
rect 611 -386 612 -384
rect 614 -386 615 -384
rect 611 -392 612 -390
rect 614 -392 615 -390
rect 618 -386 619 -384
rect 618 -392 619 -390
rect 625 -386 626 -384
rect 625 -392 626 -390
rect 632 -386 633 -384
rect 632 -392 633 -390
rect 639 -386 640 -384
rect 639 -392 640 -390
rect 646 -386 647 -384
rect 646 -392 647 -390
rect 653 -386 654 -384
rect 653 -392 654 -390
rect 660 -386 661 -384
rect 660 -392 661 -390
rect 667 -386 668 -384
rect 670 -386 671 -384
rect 670 -392 671 -390
rect 674 -386 675 -384
rect 674 -392 675 -390
rect 681 -386 682 -384
rect 681 -392 682 -390
rect 688 -386 689 -384
rect 688 -392 689 -390
rect 695 -386 696 -384
rect 695 -392 696 -390
rect 702 -386 703 -384
rect 705 -386 706 -384
rect 702 -392 703 -390
rect 709 -386 710 -384
rect 712 -386 713 -384
rect 712 -392 713 -390
rect 716 -386 717 -384
rect 716 -392 717 -390
rect 723 -386 724 -384
rect 723 -392 724 -390
rect 730 -386 731 -384
rect 733 -386 734 -384
rect 730 -392 731 -390
rect 733 -392 734 -390
rect 737 -386 738 -384
rect 737 -392 738 -390
rect 747 -386 748 -384
rect 744 -392 745 -390
rect 747 -392 748 -390
rect 751 -386 752 -384
rect 754 -386 755 -384
rect 751 -392 752 -390
rect 758 -386 759 -384
rect 758 -392 759 -390
rect 765 -386 766 -384
rect 765 -392 766 -390
rect 772 -386 773 -384
rect 772 -392 773 -390
rect 779 -386 780 -384
rect 779 -392 780 -390
rect 786 -386 787 -384
rect 786 -392 787 -390
rect 793 -386 794 -384
rect 793 -392 794 -390
rect 800 -386 801 -384
rect 800 -392 801 -390
rect 807 -386 808 -384
rect 807 -392 808 -390
rect 814 -386 815 -384
rect 814 -392 815 -390
rect 821 -386 822 -384
rect 821 -392 822 -390
rect 828 -386 829 -384
rect 828 -392 829 -390
rect 835 -386 836 -384
rect 835 -392 836 -390
rect 842 -386 843 -384
rect 842 -392 843 -390
rect 849 -386 850 -384
rect 849 -392 850 -390
rect 856 -386 857 -384
rect 856 -392 857 -390
rect 863 -386 864 -384
rect 863 -392 864 -390
rect 870 -386 871 -384
rect 870 -392 871 -390
rect 877 -386 878 -384
rect 877 -392 878 -390
rect 884 -386 885 -384
rect 884 -392 885 -390
rect 891 -386 892 -384
rect 891 -392 892 -390
rect 898 -386 899 -384
rect 898 -392 899 -390
rect 905 -386 906 -384
rect 905 -392 906 -390
rect 912 -386 913 -384
rect 912 -392 913 -390
rect 919 -386 920 -384
rect 919 -392 920 -390
rect 926 -386 927 -384
rect 926 -392 927 -390
rect 933 -386 934 -384
rect 933 -392 934 -390
rect 940 -386 941 -384
rect 940 -392 941 -390
rect 947 -386 948 -384
rect 947 -392 948 -390
rect 954 -386 955 -384
rect 954 -392 955 -390
rect 961 -386 962 -384
rect 961 -392 962 -390
rect 968 -386 969 -384
rect 968 -392 969 -390
rect 975 -386 976 -384
rect 975 -392 976 -390
rect 982 -386 983 -384
rect 982 -392 983 -390
rect 989 -386 990 -384
rect 989 -392 990 -390
rect 996 -386 997 -384
rect 996 -392 997 -390
rect 1003 -386 1004 -384
rect 1003 -392 1004 -390
rect 1010 -386 1011 -384
rect 1010 -392 1011 -390
rect 1017 -386 1018 -384
rect 1017 -392 1018 -390
rect 1024 -386 1025 -384
rect 1024 -392 1025 -390
rect 1031 -386 1032 -384
rect 1031 -392 1032 -390
rect 1038 -386 1039 -384
rect 1038 -392 1039 -390
rect 1045 -386 1046 -384
rect 1045 -392 1046 -390
rect 1052 -386 1053 -384
rect 1052 -392 1053 -390
rect 1059 -386 1060 -384
rect 1059 -392 1060 -390
rect 1066 -386 1067 -384
rect 1066 -392 1067 -390
rect 1073 -386 1074 -384
rect 1073 -392 1074 -390
rect 1080 -386 1081 -384
rect 1080 -392 1081 -390
rect 1087 -386 1088 -384
rect 1087 -392 1088 -390
rect 1094 -386 1095 -384
rect 1094 -392 1095 -390
rect 1101 -386 1102 -384
rect 1101 -392 1102 -390
rect 1108 -386 1109 -384
rect 1108 -392 1109 -390
rect 1115 -386 1116 -384
rect 1115 -392 1116 -390
rect 1122 -386 1123 -384
rect 1122 -392 1123 -390
rect 1129 -386 1130 -384
rect 1129 -392 1130 -390
rect 1136 -386 1137 -384
rect 1136 -392 1137 -390
rect 1143 -386 1144 -384
rect 1143 -392 1144 -390
rect 1150 -386 1151 -384
rect 1150 -392 1151 -390
rect 1157 -386 1158 -384
rect 1157 -392 1158 -390
rect 1164 -386 1165 -384
rect 1164 -392 1165 -390
rect 1171 -386 1172 -384
rect 1171 -392 1172 -390
rect 1178 -386 1179 -384
rect 1178 -392 1179 -390
rect 1185 -386 1186 -384
rect 1185 -392 1186 -390
rect 1192 -386 1193 -384
rect 1192 -392 1193 -390
rect 1202 -386 1203 -384
rect 1199 -392 1200 -390
rect 1206 -386 1207 -384
rect 1206 -392 1207 -390
rect 1213 -386 1214 -384
rect 1213 -392 1214 -390
rect 1220 -386 1221 -384
rect 1220 -392 1221 -390
rect 1227 -386 1228 -384
rect 1227 -392 1228 -390
rect 1234 -386 1235 -384
rect 1234 -392 1235 -390
rect 1241 -386 1242 -384
rect 1241 -392 1242 -390
rect 1248 -386 1249 -384
rect 1248 -392 1249 -390
rect 1255 -386 1256 -384
rect 1255 -392 1256 -390
rect 1262 -386 1263 -384
rect 1262 -392 1263 -390
rect 1269 -386 1270 -384
rect 1269 -392 1270 -390
rect 1276 -386 1277 -384
rect 1276 -392 1277 -390
rect 1283 -386 1284 -384
rect 1283 -392 1284 -390
rect 1290 -386 1291 -384
rect 1290 -392 1291 -390
rect 1297 -386 1298 -384
rect 1297 -392 1298 -390
rect 1304 -386 1305 -384
rect 1304 -392 1305 -390
rect 1311 -386 1312 -384
rect 1311 -392 1312 -390
rect 1318 -386 1319 -384
rect 1318 -392 1319 -390
rect 1325 -386 1326 -384
rect 1325 -392 1326 -390
rect 1332 -386 1333 -384
rect 1332 -392 1333 -390
rect 1339 -386 1340 -384
rect 1339 -392 1340 -390
rect 1346 -386 1347 -384
rect 1346 -392 1347 -390
rect 1353 -386 1354 -384
rect 1353 -392 1354 -390
rect 1360 -386 1361 -384
rect 1360 -392 1361 -390
rect 1367 -386 1368 -384
rect 1367 -392 1368 -390
rect 1374 -386 1375 -384
rect 1374 -392 1375 -390
rect 1381 -386 1382 -384
rect 1381 -392 1382 -390
rect 1388 -386 1389 -384
rect 1388 -392 1389 -390
rect 1395 -386 1396 -384
rect 1395 -392 1396 -390
rect 1398 -392 1399 -390
rect 1591 -386 1592 -384
rect 1591 -392 1592 -390
rect 23 -497 24 -495
rect 26 -497 27 -495
rect 30 -497 31 -495
rect 30 -503 31 -501
rect 37 -497 38 -495
rect 37 -503 38 -501
rect 44 -497 45 -495
rect 44 -503 45 -501
rect 51 -497 52 -495
rect 51 -503 52 -501
rect 58 -497 59 -495
rect 58 -503 59 -501
rect 65 -497 66 -495
rect 65 -503 66 -501
rect 72 -497 73 -495
rect 72 -503 73 -501
rect 79 -497 80 -495
rect 82 -497 83 -495
rect 79 -503 80 -501
rect 86 -497 87 -495
rect 89 -497 90 -495
rect 86 -503 87 -501
rect 93 -497 94 -495
rect 93 -503 94 -501
rect 100 -497 101 -495
rect 103 -497 104 -495
rect 100 -503 101 -501
rect 103 -503 104 -501
rect 107 -497 108 -495
rect 110 -497 111 -495
rect 110 -503 111 -501
rect 114 -497 115 -495
rect 114 -503 115 -501
rect 121 -497 122 -495
rect 121 -503 122 -501
rect 128 -497 129 -495
rect 128 -503 129 -501
rect 135 -497 136 -495
rect 138 -497 139 -495
rect 135 -503 136 -501
rect 138 -503 139 -501
rect 142 -497 143 -495
rect 142 -503 143 -501
rect 149 -497 150 -495
rect 149 -503 150 -501
rect 156 -497 157 -495
rect 156 -503 157 -501
rect 163 -497 164 -495
rect 163 -503 164 -501
rect 170 -497 171 -495
rect 170 -503 171 -501
rect 177 -497 178 -495
rect 180 -497 181 -495
rect 180 -503 181 -501
rect 187 -497 188 -495
rect 187 -503 188 -501
rect 191 -497 192 -495
rect 194 -497 195 -495
rect 194 -503 195 -501
rect 198 -497 199 -495
rect 198 -503 199 -501
rect 205 -497 206 -495
rect 205 -503 206 -501
rect 212 -497 213 -495
rect 212 -503 213 -501
rect 219 -497 220 -495
rect 222 -503 223 -501
rect 226 -497 227 -495
rect 226 -503 227 -501
rect 233 -497 234 -495
rect 233 -503 234 -501
rect 240 -497 241 -495
rect 240 -503 241 -501
rect 247 -497 248 -495
rect 247 -503 248 -501
rect 254 -497 255 -495
rect 254 -503 255 -501
rect 261 -497 262 -495
rect 261 -503 262 -501
rect 268 -497 269 -495
rect 268 -503 269 -501
rect 275 -497 276 -495
rect 275 -503 276 -501
rect 282 -497 283 -495
rect 282 -503 283 -501
rect 289 -497 290 -495
rect 289 -503 290 -501
rect 299 -497 300 -495
rect 299 -503 300 -501
rect 303 -497 304 -495
rect 303 -503 304 -501
rect 310 -497 311 -495
rect 310 -503 311 -501
rect 317 -497 318 -495
rect 317 -503 318 -501
rect 324 -497 325 -495
rect 324 -503 325 -501
rect 331 -497 332 -495
rect 331 -503 332 -501
rect 338 -497 339 -495
rect 338 -503 339 -501
rect 345 -497 346 -495
rect 345 -503 346 -501
rect 352 -497 353 -495
rect 352 -503 353 -501
rect 359 -497 360 -495
rect 362 -497 363 -495
rect 359 -503 360 -501
rect 362 -503 363 -501
rect 366 -497 367 -495
rect 366 -503 367 -501
rect 373 -497 374 -495
rect 373 -503 374 -501
rect 380 -497 381 -495
rect 380 -503 381 -501
rect 387 -497 388 -495
rect 387 -503 388 -501
rect 394 -497 395 -495
rect 394 -503 395 -501
rect 401 -497 402 -495
rect 401 -503 402 -501
rect 408 -497 409 -495
rect 408 -503 409 -501
rect 418 -497 419 -495
rect 418 -503 419 -501
rect 422 -497 423 -495
rect 422 -503 423 -501
rect 429 -497 430 -495
rect 429 -503 430 -501
rect 436 -497 437 -495
rect 436 -503 437 -501
rect 443 -497 444 -495
rect 443 -503 444 -501
rect 453 -497 454 -495
rect 450 -503 451 -501
rect 453 -503 454 -501
rect 457 -497 458 -495
rect 457 -503 458 -501
rect 464 -497 465 -495
rect 464 -503 465 -501
rect 471 -497 472 -495
rect 474 -497 475 -495
rect 474 -503 475 -501
rect 478 -497 479 -495
rect 481 -497 482 -495
rect 478 -503 479 -501
rect 481 -503 482 -501
rect 485 -497 486 -495
rect 485 -503 486 -501
rect 492 -497 493 -495
rect 495 -497 496 -495
rect 492 -503 493 -501
rect 495 -503 496 -501
rect 499 -497 500 -495
rect 499 -503 500 -501
rect 506 -497 507 -495
rect 506 -503 507 -501
rect 513 -497 514 -495
rect 516 -503 517 -501
rect 520 -497 521 -495
rect 523 -497 524 -495
rect 520 -503 521 -501
rect 523 -503 524 -501
rect 527 -497 528 -495
rect 530 -497 531 -495
rect 527 -503 528 -501
rect 530 -503 531 -501
rect 534 -497 535 -495
rect 534 -503 535 -501
rect 537 -503 538 -501
rect 541 -497 542 -495
rect 541 -503 542 -501
rect 548 -497 549 -495
rect 548 -503 549 -501
rect 555 -497 556 -495
rect 555 -503 556 -501
rect 562 -497 563 -495
rect 562 -503 563 -501
rect 569 -497 570 -495
rect 569 -503 570 -501
rect 576 -497 577 -495
rect 576 -503 577 -501
rect 583 -497 584 -495
rect 583 -503 584 -501
rect 590 -497 591 -495
rect 593 -497 594 -495
rect 593 -503 594 -501
rect 597 -497 598 -495
rect 597 -503 598 -501
rect 600 -503 601 -501
rect 604 -497 605 -495
rect 604 -503 605 -501
rect 611 -497 612 -495
rect 611 -503 612 -501
rect 618 -497 619 -495
rect 618 -503 619 -501
rect 625 -497 626 -495
rect 625 -503 626 -501
rect 632 -497 633 -495
rect 635 -497 636 -495
rect 635 -503 636 -501
rect 639 -497 640 -495
rect 639 -503 640 -501
rect 646 -497 647 -495
rect 649 -497 650 -495
rect 649 -503 650 -501
rect 653 -497 654 -495
rect 653 -503 654 -501
rect 660 -497 661 -495
rect 660 -503 661 -501
rect 667 -497 668 -495
rect 667 -503 668 -501
rect 674 -497 675 -495
rect 674 -503 675 -501
rect 681 -497 682 -495
rect 681 -503 682 -501
rect 688 -497 689 -495
rect 688 -503 689 -501
rect 695 -497 696 -495
rect 695 -503 696 -501
rect 698 -503 699 -501
rect 702 -497 703 -495
rect 702 -503 703 -501
rect 709 -497 710 -495
rect 709 -503 710 -501
rect 712 -503 713 -501
rect 716 -497 717 -495
rect 716 -503 717 -501
rect 723 -497 724 -495
rect 723 -503 724 -501
rect 730 -497 731 -495
rect 730 -503 731 -501
rect 737 -497 738 -495
rect 737 -503 738 -501
rect 744 -497 745 -495
rect 744 -503 745 -501
rect 751 -497 752 -495
rect 751 -503 752 -501
rect 758 -497 759 -495
rect 758 -503 759 -501
rect 761 -503 762 -501
rect 765 -497 766 -495
rect 765 -503 766 -501
rect 772 -497 773 -495
rect 772 -503 773 -501
rect 779 -497 780 -495
rect 779 -503 780 -501
rect 786 -497 787 -495
rect 786 -503 787 -501
rect 793 -497 794 -495
rect 793 -503 794 -501
rect 800 -497 801 -495
rect 800 -503 801 -501
rect 807 -497 808 -495
rect 807 -503 808 -501
rect 814 -497 815 -495
rect 814 -503 815 -501
rect 821 -497 822 -495
rect 821 -503 822 -501
rect 828 -497 829 -495
rect 828 -503 829 -501
rect 831 -503 832 -501
rect 835 -497 836 -495
rect 835 -503 836 -501
rect 842 -497 843 -495
rect 842 -503 843 -501
rect 849 -497 850 -495
rect 849 -503 850 -501
rect 856 -497 857 -495
rect 856 -503 857 -501
rect 863 -497 864 -495
rect 863 -503 864 -501
rect 870 -497 871 -495
rect 870 -503 871 -501
rect 877 -497 878 -495
rect 877 -503 878 -501
rect 884 -497 885 -495
rect 884 -503 885 -501
rect 891 -497 892 -495
rect 891 -503 892 -501
rect 898 -497 899 -495
rect 901 -503 902 -501
rect 905 -497 906 -495
rect 905 -503 906 -501
rect 912 -497 913 -495
rect 912 -503 913 -501
rect 919 -497 920 -495
rect 919 -503 920 -501
rect 926 -497 927 -495
rect 926 -503 927 -501
rect 933 -497 934 -495
rect 933 -503 934 -501
rect 940 -497 941 -495
rect 940 -503 941 -501
rect 947 -497 948 -495
rect 947 -503 948 -501
rect 954 -497 955 -495
rect 954 -503 955 -501
rect 961 -497 962 -495
rect 961 -503 962 -501
rect 968 -497 969 -495
rect 968 -503 969 -501
rect 975 -497 976 -495
rect 975 -503 976 -501
rect 982 -497 983 -495
rect 982 -503 983 -501
rect 989 -497 990 -495
rect 996 -497 997 -495
rect 996 -503 997 -501
rect 1003 -497 1004 -495
rect 1003 -503 1004 -501
rect 1010 -497 1011 -495
rect 1010 -503 1011 -501
rect 1017 -497 1018 -495
rect 1017 -503 1018 -501
rect 1024 -497 1025 -495
rect 1024 -503 1025 -501
rect 1031 -497 1032 -495
rect 1031 -503 1032 -501
rect 1038 -497 1039 -495
rect 1038 -503 1039 -501
rect 1045 -497 1046 -495
rect 1045 -503 1046 -501
rect 1052 -497 1053 -495
rect 1052 -503 1053 -501
rect 1059 -497 1060 -495
rect 1059 -503 1060 -501
rect 1066 -497 1067 -495
rect 1066 -503 1067 -501
rect 1073 -497 1074 -495
rect 1073 -503 1074 -501
rect 1080 -497 1081 -495
rect 1080 -503 1081 -501
rect 1087 -497 1088 -495
rect 1087 -503 1088 -501
rect 1094 -497 1095 -495
rect 1094 -503 1095 -501
rect 1101 -497 1102 -495
rect 1101 -503 1102 -501
rect 1108 -497 1109 -495
rect 1108 -503 1109 -501
rect 1115 -497 1116 -495
rect 1115 -503 1116 -501
rect 1122 -497 1123 -495
rect 1122 -503 1123 -501
rect 1129 -497 1130 -495
rect 1129 -503 1130 -501
rect 1136 -497 1137 -495
rect 1136 -503 1137 -501
rect 1143 -497 1144 -495
rect 1143 -503 1144 -501
rect 1150 -497 1151 -495
rect 1150 -503 1151 -501
rect 1157 -497 1158 -495
rect 1157 -503 1158 -501
rect 1164 -497 1165 -495
rect 1164 -503 1165 -501
rect 1171 -497 1172 -495
rect 1171 -503 1172 -501
rect 1178 -497 1179 -495
rect 1178 -503 1179 -501
rect 1185 -497 1186 -495
rect 1185 -503 1186 -501
rect 1195 -503 1196 -501
rect 1199 -497 1200 -495
rect 1199 -503 1200 -501
rect 1206 -497 1207 -495
rect 1206 -503 1207 -501
rect 1213 -497 1214 -495
rect 1213 -503 1214 -501
rect 1220 -497 1221 -495
rect 1220 -503 1221 -501
rect 1227 -497 1228 -495
rect 1227 -503 1228 -501
rect 1234 -497 1235 -495
rect 1234 -503 1235 -501
rect 1241 -497 1242 -495
rect 1241 -503 1242 -501
rect 1248 -497 1249 -495
rect 1248 -503 1249 -501
rect 1255 -497 1256 -495
rect 1255 -503 1256 -501
rect 1262 -497 1263 -495
rect 1262 -503 1263 -501
rect 1269 -497 1270 -495
rect 1269 -503 1270 -501
rect 1272 -503 1273 -501
rect 1276 -497 1277 -495
rect 1276 -503 1277 -501
rect 1283 -497 1284 -495
rect 1283 -503 1284 -501
rect 1290 -497 1291 -495
rect 1290 -503 1291 -501
rect 1297 -497 1298 -495
rect 1297 -503 1298 -501
rect 1304 -497 1305 -495
rect 1304 -503 1305 -501
rect 1311 -497 1312 -495
rect 1311 -503 1312 -501
rect 1318 -497 1319 -495
rect 1318 -503 1319 -501
rect 1325 -497 1326 -495
rect 1325 -503 1326 -501
rect 1332 -497 1333 -495
rect 1332 -503 1333 -501
rect 1339 -497 1340 -495
rect 1339 -503 1340 -501
rect 1346 -497 1347 -495
rect 1346 -503 1347 -501
rect 1353 -497 1354 -495
rect 1353 -503 1354 -501
rect 1360 -497 1361 -495
rect 1360 -503 1361 -501
rect 1367 -497 1368 -495
rect 1367 -503 1368 -501
rect 1374 -497 1375 -495
rect 1374 -503 1375 -501
rect 1381 -497 1382 -495
rect 1381 -503 1382 -501
rect 1388 -497 1389 -495
rect 1388 -503 1389 -501
rect 1395 -497 1396 -495
rect 1395 -503 1396 -501
rect 1402 -497 1403 -495
rect 1402 -503 1403 -501
rect 1409 -497 1410 -495
rect 1409 -503 1410 -501
rect 1416 -497 1417 -495
rect 1416 -503 1417 -501
rect 1423 -497 1424 -495
rect 1423 -503 1424 -501
rect 1430 -497 1431 -495
rect 1430 -503 1431 -501
rect 1437 -497 1438 -495
rect 1437 -503 1438 -501
rect 1444 -497 1445 -495
rect 1444 -503 1445 -501
rect 1451 -497 1452 -495
rect 1451 -503 1452 -501
rect 1458 -497 1459 -495
rect 1458 -503 1459 -501
rect 1465 -497 1466 -495
rect 1465 -503 1466 -501
rect 1472 -497 1473 -495
rect 1472 -503 1473 -501
rect 1479 -497 1480 -495
rect 1479 -503 1480 -501
rect 1486 -497 1487 -495
rect 1486 -503 1487 -501
rect 1493 -497 1494 -495
rect 1493 -503 1494 -501
rect 1500 -497 1501 -495
rect 1500 -503 1501 -501
rect 1503 -503 1504 -501
rect 1507 -497 1508 -495
rect 1507 -503 1508 -501
rect 1514 -497 1515 -495
rect 1514 -503 1515 -501
rect 1524 -497 1525 -495
rect 1528 -497 1529 -495
rect 1528 -503 1529 -501
rect 1710 -497 1711 -495
rect 1710 -503 1711 -501
rect 9 -604 10 -602
rect 9 -610 10 -608
rect 23 -604 24 -602
rect 23 -610 24 -608
rect 30 -604 31 -602
rect 30 -610 31 -608
rect 44 -604 45 -602
rect 44 -610 45 -608
rect 51 -604 52 -602
rect 51 -610 52 -608
rect 61 -604 62 -602
rect 58 -610 59 -608
rect 61 -610 62 -608
rect 65 -604 66 -602
rect 65 -610 66 -608
rect 72 -604 73 -602
rect 72 -610 73 -608
rect 79 -604 80 -602
rect 79 -610 80 -608
rect 86 -604 87 -602
rect 86 -610 87 -608
rect 93 -604 94 -602
rect 93 -610 94 -608
rect 103 -604 104 -602
rect 100 -610 101 -608
rect 103 -610 104 -608
rect 107 -604 108 -602
rect 114 -604 115 -602
rect 114 -610 115 -608
rect 121 -604 122 -602
rect 121 -610 122 -608
rect 128 -604 129 -602
rect 128 -610 129 -608
rect 135 -604 136 -602
rect 135 -610 136 -608
rect 142 -604 143 -602
rect 142 -610 143 -608
rect 149 -604 150 -602
rect 152 -604 153 -602
rect 149 -610 150 -608
rect 152 -610 153 -608
rect 156 -604 157 -602
rect 156 -610 157 -608
rect 163 -604 164 -602
rect 163 -610 164 -608
rect 170 -604 171 -602
rect 170 -610 171 -608
rect 177 -604 178 -602
rect 177 -610 178 -608
rect 184 -604 185 -602
rect 184 -610 185 -608
rect 187 -610 188 -608
rect 191 -604 192 -602
rect 191 -610 192 -608
rect 198 -604 199 -602
rect 198 -610 199 -608
rect 205 -604 206 -602
rect 205 -610 206 -608
rect 212 -604 213 -602
rect 212 -610 213 -608
rect 219 -604 220 -602
rect 219 -610 220 -608
rect 226 -604 227 -602
rect 226 -610 227 -608
rect 233 -610 234 -608
rect 236 -610 237 -608
rect 240 -604 241 -602
rect 243 -604 244 -602
rect 240 -610 241 -608
rect 243 -610 244 -608
rect 247 -604 248 -602
rect 247 -610 248 -608
rect 254 -604 255 -602
rect 254 -610 255 -608
rect 261 -604 262 -602
rect 261 -610 262 -608
rect 268 -604 269 -602
rect 268 -610 269 -608
rect 275 -604 276 -602
rect 275 -610 276 -608
rect 282 -604 283 -602
rect 282 -610 283 -608
rect 289 -604 290 -602
rect 289 -610 290 -608
rect 296 -604 297 -602
rect 296 -610 297 -608
rect 303 -604 304 -602
rect 303 -610 304 -608
rect 310 -604 311 -602
rect 310 -610 311 -608
rect 317 -604 318 -602
rect 320 -610 321 -608
rect 324 -604 325 -602
rect 324 -610 325 -608
rect 331 -604 332 -602
rect 331 -610 332 -608
rect 338 -604 339 -602
rect 341 -604 342 -602
rect 338 -610 339 -608
rect 345 -604 346 -602
rect 345 -610 346 -608
rect 352 -604 353 -602
rect 352 -610 353 -608
rect 359 -604 360 -602
rect 359 -610 360 -608
rect 366 -604 367 -602
rect 366 -610 367 -608
rect 373 -604 374 -602
rect 373 -610 374 -608
rect 383 -610 384 -608
rect 387 -604 388 -602
rect 387 -610 388 -608
rect 394 -604 395 -602
rect 394 -610 395 -608
rect 401 -604 402 -602
rect 401 -610 402 -608
rect 408 -604 409 -602
rect 408 -610 409 -608
rect 415 -604 416 -602
rect 415 -610 416 -608
rect 422 -604 423 -602
rect 422 -610 423 -608
rect 429 -610 430 -608
rect 432 -610 433 -608
rect 436 -604 437 -602
rect 436 -610 437 -608
rect 443 -604 444 -602
rect 443 -610 444 -608
rect 450 -604 451 -602
rect 453 -604 454 -602
rect 450 -610 451 -608
rect 453 -610 454 -608
rect 457 -604 458 -602
rect 460 -604 461 -602
rect 457 -610 458 -608
rect 464 -604 465 -602
rect 464 -610 465 -608
rect 471 -604 472 -602
rect 471 -610 472 -608
rect 478 -604 479 -602
rect 478 -610 479 -608
rect 485 -604 486 -602
rect 485 -610 486 -608
rect 492 -604 493 -602
rect 492 -610 493 -608
rect 499 -604 500 -602
rect 499 -610 500 -608
rect 506 -604 507 -602
rect 506 -610 507 -608
rect 513 -604 514 -602
rect 516 -604 517 -602
rect 513 -610 514 -608
rect 520 -604 521 -602
rect 520 -610 521 -608
rect 527 -604 528 -602
rect 530 -604 531 -602
rect 527 -610 528 -608
rect 530 -610 531 -608
rect 534 -604 535 -602
rect 534 -610 535 -608
rect 541 -604 542 -602
rect 541 -610 542 -608
rect 548 -604 549 -602
rect 548 -610 549 -608
rect 555 -604 556 -602
rect 555 -610 556 -608
rect 562 -604 563 -602
rect 562 -610 563 -608
rect 569 -604 570 -602
rect 569 -610 570 -608
rect 576 -604 577 -602
rect 579 -604 580 -602
rect 576 -610 577 -608
rect 583 -604 584 -602
rect 586 -604 587 -602
rect 586 -610 587 -608
rect 590 -604 591 -602
rect 593 -604 594 -602
rect 590 -610 591 -608
rect 593 -610 594 -608
rect 597 -604 598 -602
rect 597 -610 598 -608
rect 604 -604 605 -602
rect 604 -610 605 -608
rect 611 -604 612 -602
rect 611 -610 612 -608
rect 618 -604 619 -602
rect 618 -610 619 -608
rect 625 -604 626 -602
rect 625 -610 626 -608
rect 632 -604 633 -602
rect 635 -604 636 -602
rect 635 -610 636 -608
rect 639 -604 640 -602
rect 639 -610 640 -608
rect 646 -604 647 -602
rect 646 -610 647 -608
rect 653 -604 654 -602
rect 653 -610 654 -608
rect 656 -610 657 -608
rect 660 -604 661 -602
rect 660 -610 661 -608
rect 667 -604 668 -602
rect 667 -610 668 -608
rect 674 -604 675 -602
rect 677 -604 678 -602
rect 677 -610 678 -608
rect 681 -604 682 -602
rect 681 -610 682 -608
rect 688 -604 689 -602
rect 688 -610 689 -608
rect 698 -604 699 -602
rect 695 -610 696 -608
rect 698 -610 699 -608
rect 702 -604 703 -602
rect 702 -610 703 -608
rect 709 -604 710 -602
rect 709 -610 710 -608
rect 716 -604 717 -602
rect 716 -610 717 -608
rect 723 -604 724 -602
rect 723 -610 724 -608
rect 730 -604 731 -602
rect 730 -610 731 -608
rect 737 -604 738 -602
rect 737 -610 738 -608
rect 744 -604 745 -602
rect 744 -610 745 -608
rect 751 -604 752 -602
rect 751 -610 752 -608
rect 758 -604 759 -602
rect 758 -610 759 -608
rect 765 -604 766 -602
rect 765 -610 766 -608
rect 772 -604 773 -602
rect 772 -610 773 -608
rect 779 -604 780 -602
rect 779 -610 780 -608
rect 786 -604 787 -602
rect 786 -610 787 -608
rect 793 -604 794 -602
rect 793 -610 794 -608
rect 800 -604 801 -602
rect 800 -610 801 -608
rect 807 -604 808 -602
rect 807 -610 808 -608
rect 814 -604 815 -602
rect 814 -610 815 -608
rect 821 -604 822 -602
rect 824 -604 825 -602
rect 821 -610 822 -608
rect 824 -610 825 -608
rect 828 -604 829 -602
rect 828 -610 829 -608
rect 835 -604 836 -602
rect 835 -610 836 -608
rect 842 -604 843 -602
rect 845 -604 846 -602
rect 842 -610 843 -608
rect 849 -604 850 -602
rect 852 -604 853 -602
rect 849 -610 850 -608
rect 852 -610 853 -608
rect 856 -604 857 -602
rect 856 -610 857 -608
rect 866 -604 867 -602
rect 863 -610 864 -608
rect 866 -610 867 -608
rect 873 -604 874 -602
rect 870 -610 871 -608
rect 873 -610 874 -608
rect 877 -604 878 -602
rect 877 -610 878 -608
rect 884 -604 885 -602
rect 884 -610 885 -608
rect 891 -604 892 -602
rect 894 -604 895 -602
rect 894 -610 895 -608
rect 898 -610 899 -608
rect 905 -604 906 -602
rect 905 -610 906 -608
rect 912 -604 913 -602
rect 915 -604 916 -602
rect 915 -610 916 -608
rect 919 -604 920 -602
rect 919 -610 920 -608
rect 926 -604 927 -602
rect 926 -610 927 -608
rect 933 -610 934 -608
rect 940 -604 941 -602
rect 940 -610 941 -608
rect 947 -604 948 -602
rect 947 -610 948 -608
rect 954 -604 955 -602
rect 954 -610 955 -608
rect 961 -604 962 -602
rect 961 -610 962 -608
rect 968 -604 969 -602
rect 968 -610 969 -608
rect 975 -604 976 -602
rect 975 -610 976 -608
rect 982 -604 983 -602
rect 982 -610 983 -608
rect 989 -610 990 -608
rect 996 -604 997 -602
rect 996 -610 997 -608
rect 1003 -604 1004 -602
rect 1003 -610 1004 -608
rect 1010 -604 1011 -602
rect 1010 -610 1011 -608
rect 1017 -604 1018 -602
rect 1017 -610 1018 -608
rect 1024 -604 1025 -602
rect 1024 -610 1025 -608
rect 1031 -604 1032 -602
rect 1031 -610 1032 -608
rect 1038 -604 1039 -602
rect 1038 -610 1039 -608
rect 1045 -604 1046 -602
rect 1045 -610 1046 -608
rect 1052 -604 1053 -602
rect 1055 -604 1056 -602
rect 1059 -604 1060 -602
rect 1059 -610 1060 -608
rect 1066 -604 1067 -602
rect 1066 -610 1067 -608
rect 1073 -604 1074 -602
rect 1073 -610 1074 -608
rect 1080 -604 1081 -602
rect 1080 -610 1081 -608
rect 1087 -604 1088 -602
rect 1087 -610 1088 -608
rect 1094 -604 1095 -602
rect 1094 -610 1095 -608
rect 1101 -604 1102 -602
rect 1101 -610 1102 -608
rect 1108 -604 1109 -602
rect 1108 -610 1109 -608
rect 1115 -604 1116 -602
rect 1115 -610 1116 -608
rect 1122 -604 1123 -602
rect 1122 -610 1123 -608
rect 1129 -604 1130 -602
rect 1129 -610 1130 -608
rect 1136 -604 1137 -602
rect 1136 -610 1137 -608
rect 1143 -604 1144 -602
rect 1143 -610 1144 -608
rect 1150 -604 1151 -602
rect 1150 -610 1151 -608
rect 1157 -604 1158 -602
rect 1157 -610 1158 -608
rect 1164 -604 1165 -602
rect 1164 -610 1165 -608
rect 1171 -604 1172 -602
rect 1171 -610 1172 -608
rect 1178 -604 1179 -602
rect 1178 -610 1179 -608
rect 1185 -604 1186 -602
rect 1185 -610 1186 -608
rect 1192 -604 1193 -602
rect 1192 -610 1193 -608
rect 1199 -604 1200 -602
rect 1199 -610 1200 -608
rect 1206 -604 1207 -602
rect 1206 -610 1207 -608
rect 1213 -604 1214 -602
rect 1213 -610 1214 -608
rect 1220 -604 1221 -602
rect 1220 -610 1221 -608
rect 1227 -604 1228 -602
rect 1227 -610 1228 -608
rect 1234 -604 1235 -602
rect 1234 -610 1235 -608
rect 1241 -604 1242 -602
rect 1241 -610 1242 -608
rect 1248 -604 1249 -602
rect 1248 -610 1249 -608
rect 1255 -604 1256 -602
rect 1255 -610 1256 -608
rect 1262 -604 1263 -602
rect 1262 -610 1263 -608
rect 1269 -604 1270 -602
rect 1272 -604 1273 -602
rect 1269 -610 1270 -608
rect 1276 -604 1277 -602
rect 1276 -610 1277 -608
rect 1283 -604 1284 -602
rect 1283 -610 1284 -608
rect 1290 -604 1291 -602
rect 1290 -610 1291 -608
rect 1297 -604 1298 -602
rect 1297 -610 1298 -608
rect 1304 -604 1305 -602
rect 1304 -610 1305 -608
rect 1311 -604 1312 -602
rect 1311 -610 1312 -608
rect 1318 -604 1319 -602
rect 1318 -610 1319 -608
rect 1325 -604 1326 -602
rect 1325 -610 1326 -608
rect 1332 -604 1333 -602
rect 1332 -610 1333 -608
rect 1339 -604 1340 -602
rect 1339 -610 1340 -608
rect 1346 -604 1347 -602
rect 1346 -610 1347 -608
rect 1353 -604 1354 -602
rect 1353 -610 1354 -608
rect 1360 -604 1361 -602
rect 1360 -610 1361 -608
rect 1367 -604 1368 -602
rect 1367 -610 1368 -608
rect 1374 -604 1375 -602
rect 1374 -610 1375 -608
rect 1381 -604 1382 -602
rect 1381 -610 1382 -608
rect 1388 -604 1389 -602
rect 1388 -610 1389 -608
rect 1395 -604 1396 -602
rect 1395 -610 1396 -608
rect 1402 -604 1403 -602
rect 1402 -610 1403 -608
rect 1409 -604 1410 -602
rect 1409 -610 1410 -608
rect 1416 -604 1417 -602
rect 1416 -610 1417 -608
rect 1423 -604 1424 -602
rect 1423 -610 1424 -608
rect 1430 -604 1431 -602
rect 1430 -610 1431 -608
rect 1437 -604 1438 -602
rect 1437 -610 1438 -608
rect 1444 -604 1445 -602
rect 1444 -610 1445 -608
rect 1451 -604 1452 -602
rect 1451 -610 1452 -608
rect 1458 -604 1459 -602
rect 1458 -610 1459 -608
rect 1468 -604 1469 -602
rect 1465 -610 1466 -608
rect 1468 -610 1469 -608
rect 1472 -604 1473 -602
rect 1472 -610 1473 -608
rect 1479 -604 1480 -602
rect 1479 -610 1480 -608
rect 1486 -604 1487 -602
rect 1486 -610 1487 -608
rect 1493 -604 1494 -602
rect 1493 -610 1494 -608
rect 1500 -604 1501 -602
rect 1503 -604 1504 -602
rect 1500 -610 1501 -608
rect 1507 -604 1508 -602
rect 1507 -610 1508 -608
rect 1514 -604 1515 -602
rect 1514 -610 1515 -608
rect 1521 -604 1522 -602
rect 1521 -610 1522 -608
rect 1535 -604 1536 -602
rect 1535 -610 1536 -608
rect 1556 -604 1557 -602
rect 1556 -610 1557 -608
rect 1738 -604 1739 -602
rect 1738 -610 1739 -608
rect 1759 -604 1760 -602
rect 1759 -610 1760 -608
rect 1766 -604 1767 -602
rect 1766 -610 1767 -608
rect 9 -713 10 -711
rect 9 -719 10 -717
rect 16 -713 17 -711
rect 16 -719 17 -717
rect 23 -713 24 -711
rect 23 -719 24 -717
rect 30 -713 31 -711
rect 30 -719 31 -717
rect 37 -713 38 -711
rect 37 -719 38 -717
rect 44 -713 45 -711
rect 44 -719 45 -717
rect 51 -713 52 -711
rect 51 -719 52 -717
rect 58 -713 59 -711
rect 58 -719 59 -717
rect 65 -713 66 -711
rect 65 -719 66 -717
rect 72 -713 73 -711
rect 72 -719 73 -717
rect 79 -713 80 -711
rect 79 -719 80 -717
rect 86 -713 87 -711
rect 86 -719 87 -717
rect 96 -713 97 -711
rect 93 -719 94 -717
rect 96 -719 97 -717
rect 100 -713 101 -711
rect 100 -719 101 -717
rect 107 -719 108 -717
rect 114 -713 115 -711
rect 117 -713 118 -711
rect 114 -719 115 -717
rect 117 -719 118 -717
rect 121 -713 122 -711
rect 121 -719 122 -717
rect 128 -713 129 -711
rect 128 -719 129 -717
rect 135 -713 136 -711
rect 135 -719 136 -717
rect 138 -719 139 -717
rect 142 -713 143 -711
rect 145 -713 146 -711
rect 142 -719 143 -717
rect 145 -719 146 -717
rect 149 -713 150 -711
rect 149 -719 150 -717
rect 156 -713 157 -711
rect 156 -719 157 -717
rect 163 -713 164 -711
rect 163 -719 164 -717
rect 170 -713 171 -711
rect 173 -713 174 -711
rect 170 -719 171 -717
rect 173 -719 174 -717
rect 177 -713 178 -711
rect 177 -719 178 -717
rect 184 -719 185 -717
rect 187 -719 188 -717
rect 191 -713 192 -711
rect 191 -719 192 -717
rect 198 -713 199 -711
rect 198 -719 199 -717
rect 205 -713 206 -711
rect 205 -719 206 -717
rect 212 -713 213 -711
rect 212 -719 213 -717
rect 219 -713 220 -711
rect 219 -719 220 -717
rect 226 -713 227 -711
rect 226 -719 227 -717
rect 236 -713 237 -711
rect 233 -719 234 -717
rect 240 -713 241 -711
rect 240 -719 241 -717
rect 247 -713 248 -711
rect 247 -719 248 -717
rect 254 -713 255 -711
rect 254 -719 255 -717
rect 261 -713 262 -711
rect 261 -719 262 -717
rect 268 -713 269 -711
rect 268 -719 269 -717
rect 275 -713 276 -711
rect 275 -719 276 -717
rect 282 -713 283 -711
rect 282 -719 283 -717
rect 289 -713 290 -711
rect 289 -719 290 -717
rect 296 -713 297 -711
rect 296 -719 297 -717
rect 303 -713 304 -711
rect 303 -719 304 -717
rect 310 -713 311 -711
rect 310 -719 311 -717
rect 317 -713 318 -711
rect 324 -713 325 -711
rect 324 -719 325 -717
rect 331 -713 332 -711
rect 331 -719 332 -717
rect 338 -713 339 -711
rect 338 -719 339 -717
rect 345 -713 346 -711
rect 345 -719 346 -717
rect 352 -713 353 -711
rect 352 -719 353 -717
rect 359 -713 360 -711
rect 362 -713 363 -711
rect 359 -719 360 -717
rect 366 -713 367 -711
rect 366 -719 367 -717
rect 373 -713 374 -711
rect 373 -719 374 -717
rect 380 -713 381 -711
rect 380 -719 381 -717
rect 387 -713 388 -711
rect 387 -719 388 -717
rect 394 -713 395 -711
rect 394 -719 395 -717
rect 401 -713 402 -711
rect 401 -719 402 -717
rect 408 -713 409 -711
rect 408 -719 409 -717
rect 415 -713 416 -711
rect 415 -719 416 -717
rect 422 -713 423 -711
rect 422 -719 423 -717
rect 429 -713 430 -711
rect 429 -719 430 -717
rect 436 -713 437 -711
rect 436 -719 437 -717
rect 443 -713 444 -711
rect 443 -719 444 -717
rect 450 -713 451 -711
rect 450 -719 451 -717
rect 457 -713 458 -711
rect 457 -719 458 -717
rect 464 -713 465 -711
rect 467 -713 468 -711
rect 464 -719 465 -717
rect 467 -719 468 -717
rect 471 -713 472 -711
rect 471 -719 472 -717
rect 478 -713 479 -711
rect 481 -713 482 -711
rect 478 -719 479 -717
rect 485 -713 486 -711
rect 485 -719 486 -717
rect 492 -713 493 -711
rect 492 -719 493 -717
rect 499 -713 500 -711
rect 499 -719 500 -717
rect 506 -713 507 -711
rect 509 -713 510 -711
rect 509 -719 510 -717
rect 513 -713 514 -711
rect 513 -719 514 -717
rect 520 -713 521 -711
rect 520 -719 521 -717
rect 527 -713 528 -711
rect 527 -719 528 -717
rect 534 -713 535 -711
rect 534 -719 535 -717
rect 541 -713 542 -711
rect 544 -713 545 -711
rect 544 -719 545 -717
rect 548 -713 549 -711
rect 548 -719 549 -717
rect 555 -719 556 -717
rect 558 -719 559 -717
rect 562 -713 563 -711
rect 562 -719 563 -717
rect 569 -713 570 -711
rect 569 -719 570 -717
rect 576 -713 577 -711
rect 576 -719 577 -717
rect 583 -713 584 -711
rect 583 -719 584 -717
rect 590 -713 591 -711
rect 590 -719 591 -717
rect 597 -713 598 -711
rect 600 -713 601 -711
rect 600 -719 601 -717
rect 604 -713 605 -711
rect 604 -719 605 -717
rect 611 -713 612 -711
rect 611 -719 612 -717
rect 618 -713 619 -711
rect 621 -713 622 -711
rect 618 -719 619 -717
rect 621 -719 622 -717
rect 625 -713 626 -711
rect 625 -719 626 -717
rect 632 -713 633 -711
rect 632 -719 633 -717
rect 639 -713 640 -711
rect 639 -719 640 -717
rect 646 -713 647 -711
rect 649 -713 650 -711
rect 646 -719 647 -717
rect 649 -719 650 -717
rect 653 -713 654 -711
rect 656 -713 657 -711
rect 653 -719 654 -717
rect 660 -713 661 -711
rect 660 -719 661 -717
rect 667 -713 668 -711
rect 667 -719 668 -717
rect 674 -713 675 -711
rect 674 -719 675 -717
rect 681 -713 682 -711
rect 681 -719 682 -717
rect 691 -713 692 -711
rect 688 -719 689 -717
rect 695 -713 696 -711
rect 695 -719 696 -717
rect 702 -713 703 -711
rect 702 -719 703 -717
rect 709 -713 710 -711
rect 712 -713 713 -711
rect 709 -719 710 -717
rect 712 -719 713 -717
rect 719 -713 720 -711
rect 716 -719 717 -717
rect 719 -719 720 -717
rect 723 -713 724 -711
rect 723 -719 724 -717
rect 730 -713 731 -711
rect 730 -719 731 -717
rect 737 -713 738 -711
rect 740 -713 741 -711
rect 737 -719 738 -717
rect 740 -719 741 -717
rect 744 -713 745 -711
rect 744 -719 745 -717
rect 751 -713 752 -711
rect 751 -719 752 -717
rect 758 -713 759 -711
rect 761 -713 762 -711
rect 758 -719 759 -717
rect 761 -719 762 -717
rect 765 -713 766 -711
rect 765 -719 766 -717
rect 772 -713 773 -711
rect 772 -719 773 -717
rect 779 -713 780 -711
rect 782 -713 783 -711
rect 779 -719 780 -717
rect 782 -719 783 -717
rect 786 -713 787 -711
rect 786 -719 787 -717
rect 793 -713 794 -711
rect 796 -713 797 -711
rect 793 -719 794 -717
rect 800 -713 801 -711
rect 800 -719 801 -717
rect 803 -719 804 -717
rect 807 -713 808 -711
rect 807 -719 808 -717
rect 814 -713 815 -711
rect 814 -719 815 -717
rect 821 -713 822 -711
rect 821 -719 822 -717
rect 828 -713 829 -711
rect 831 -713 832 -711
rect 828 -719 829 -717
rect 835 -713 836 -711
rect 835 -719 836 -717
rect 842 -713 843 -711
rect 845 -713 846 -711
rect 842 -719 843 -717
rect 845 -719 846 -717
rect 849 -713 850 -711
rect 849 -719 850 -717
rect 856 -713 857 -711
rect 856 -719 857 -717
rect 863 -713 864 -711
rect 863 -719 864 -717
rect 870 -713 871 -711
rect 870 -719 871 -717
rect 877 -713 878 -711
rect 877 -719 878 -717
rect 884 -713 885 -711
rect 884 -719 885 -717
rect 891 -713 892 -711
rect 891 -719 892 -717
rect 898 -713 899 -711
rect 901 -713 902 -711
rect 898 -719 899 -717
rect 901 -719 902 -717
rect 908 -713 909 -711
rect 908 -719 909 -717
rect 912 -713 913 -711
rect 912 -719 913 -717
rect 922 -713 923 -711
rect 919 -719 920 -717
rect 922 -719 923 -717
rect 926 -713 927 -711
rect 926 -719 927 -717
rect 933 -713 934 -711
rect 933 -719 934 -717
rect 940 -713 941 -711
rect 940 -719 941 -717
rect 947 -713 948 -711
rect 947 -719 948 -717
rect 954 -713 955 -711
rect 954 -719 955 -717
rect 961 -713 962 -711
rect 961 -719 962 -717
rect 971 -713 972 -711
rect 968 -719 969 -717
rect 971 -719 972 -717
rect 975 -713 976 -711
rect 975 -719 976 -717
rect 982 -713 983 -711
rect 982 -719 983 -717
rect 989 -713 990 -711
rect 989 -719 990 -717
rect 999 -713 1000 -711
rect 999 -719 1000 -717
rect 1003 -713 1004 -711
rect 1003 -719 1004 -717
rect 1010 -713 1011 -711
rect 1010 -719 1011 -717
rect 1020 -713 1021 -711
rect 1017 -719 1018 -717
rect 1020 -719 1021 -717
rect 1024 -713 1025 -711
rect 1024 -719 1025 -717
rect 1031 -713 1032 -711
rect 1031 -719 1032 -717
rect 1038 -713 1039 -711
rect 1038 -719 1039 -717
rect 1045 -713 1046 -711
rect 1045 -719 1046 -717
rect 1052 -713 1053 -711
rect 1052 -719 1053 -717
rect 1059 -713 1060 -711
rect 1059 -719 1060 -717
rect 1066 -713 1067 -711
rect 1066 -719 1067 -717
rect 1073 -713 1074 -711
rect 1073 -719 1074 -717
rect 1080 -713 1081 -711
rect 1080 -719 1081 -717
rect 1087 -713 1088 -711
rect 1087 -719 1088 -717
rect 1094 -713 1095 -711
rect 1094 -719 1095 -717
rect 1101 -713 1102 -711
rect 1101 -719 1102 -717
rect 1108 -713 1109 -711
rect 1108 -719 1109 -717
rect 1115 -713 1116 -711
rect 1115 -719 1116 -717
rect 1122 -713 1123 -711
rect 1122 -719 1123 -717
rect 1129 -713 1130 -711
rect 1129 -719 1130 -717
rect 1136 -713 1137 -711
rect 1136 -719 1137 -717
rect 1143 -713 1144 -711
rect 1143 -719 1144 -717
rect 1150 -713 1151 -711
rect 1150 -719 1151 -717
rect 1157 -713 1158 -711
rect 1157 -719 1158 -717
rect 1164 -713 1165 -711
rect 1164 -719 1165 -717
rect 1171 -713 1172 -711
rect 1171 -719 1172 -717
rect 1178 -713 1179 -711
rect 1178 -719 1179 -717
rect 1185 -713 1186 -711
rect 1185 -719 1186 -717
rect 1192 -713 1193 -711
rect 1192 -719 1193 -717
rect 1199 -713 1200 -711
rect 1199 -719 1200 -717
rect 1206 -713 1207 -711
rect 1206 -719 1207 -717
rect 1213 -713 1214 -711
rect 1213 -719 1214 -717
rect 1220 -713 1221 -711
rect 1220 -719 1221 -717
rect 1227 -713 1228 -711
rect 1227 -719 1228 -717
rect 1234 -713 1235 -711
rect 1234 -719 1235 -717
rect 1241 -713 1242 -711
rect 1241 -719 1242 -717
rect 1248 -713 1249 -711
rect 1248 -719 1249 -717
rect 1255 -713 1256 -711
rect 1255 -719 1256 -717
rect 1262 -713 1263 -711
rect 1262 -719 1263 -717
rect 1269 -713 1270 -711
rect 1269 -719 1270 -717
rect 1276 -713 1277 -711
rect 1276 -719 1277 -717
rect 1283 -713 1284 -711
rect 1283 -719 1284 -717
rect 1290 -713 1291 -711
rect 1290 -719 1291 -717
rect 1297 -713 1298 -711
rect 1297 -719 1298 -717
rect 1304 -713 1305 -711
rect 1304 -719 1305 -717
rect 1311 -713 1312 -711
rect 1311 -719 1312 -717
rect 1318 -713 1319 -711
rect 1318 -719 1319 -717
rect 1325 -713 1326 -711
rect 1325 -719 1326 -717
rect 1332 -713 1333 -711
rect 1332 -719 1333 -717
rect 1339 -713 1340 -711
rect 1339 -719 1340 -717
rect 1346 -713 1347 -711
rect 1346 -719 1347 -717
rect 1353 -713 1354 -711
rect 1353 -719 1354 -717
rect 1360 -713 1361 -711
rect 1360 -719 1361 -717
rect 1367 -713 1368 -711
rect 1367 -719 1368 -717
rect 1374 -713 1375 -711
rect 1374 -719 1375 -717
rect 1381 -713 1382 -711
rect 1381 -719 1382 -717
rect 1388 -713 1389 -711
rect 1388 -719 1389 -717
rect 1395 -713 1396 -711
rect 1395 -719 1396 -717
rect 1402 -713 1403 -711
rect 1402 -719 1403 -717
rect 1409 -713 1410 -711
rect 1409 -719 1410 -717
rect 1416 -713 1417 -711
rect 1416 -719 1417 -717
rect 1423 -713 1424 -711
rect 1423 -719 1424 -717
rect 1430 -713 1431 -711
rect 1430 -719 1431 -717
rect 1437 -713 1438 -711
rect 1437 -719 1438 -717
rect 1444 -713 1445 -711
rect 1444 -719 1445 -717
rect 1451 -713 1452 -711
rect 1451 -719 1452 -717
rect 1458 -713 1459 -711
rect 1458 -719 1459 -717
rect 1465 -713 1466 -711
rect 1465 -719 1466 -717
rect 1472 -713 1473 -711
rect 1472 -719 1473 -717
rect 1479 -713 1480 -711
rect 1479 -719 1480 -717
rect 1486 -713 1487 -711
rect 1486 -719 1487 -717
rect 1493 -713 1494 -711
rect 1493 -719 1494 -717
rect 1500 -713 1501 -711
rect 1500 -719 1501 -717
rect 1507 -713 1508 -711
rect 1507 -719 1508 -717
rect 1514 -713 1515 -711
rect 1514 -719 1515 -717
rect 1521 -713 1522 -711
rect 1521 -719 1522 -717
rect 1528 -713 1529 -711
rect 1528 -719 1529 -717
rect 1535 -713 1536 -711
rect 1535 -719 1536 -717
rect 1542 -713 1543 -711
rect 1542 -719 1543 -717
rect 1549 -713 1550 -711
rect 1549 -719 1550 -717
rect 1556 -713 1557 -711
rect 1556 -719 1557 -717
rect 1563 -713 1564 -711
rect 1563 -719 1564 -717
rect 1570 -713 1571 -711
rect 1570 -719 1571 -717
rect 1577 -713 1578 -711
rect 1577 -719 1578 -717
rect 1584 -713 1585 -711
rect 1584 -719 1585 -717
rect 1591 -713 1592 -711
rect 1591 -719 1592 -717
rect 1598 -713 1599 -711
rect 1598 -719 1599 -717
rect 1605 -713 1606 -711
rect 1605 -719 1606 -717
rect 1612 -713 1613 -711
rect 1612 -719 1613 -717
rect 1619 -713 1620 -711
rect 1619 -719 1620 -717
rect 1626 -713 1627 -711
rect 1626 -719 1627 -717
rect 1633 -713 1634 -711
rect 1633 -719 1634 -717
rect 1640 -713 1641 -711
rect 1640 -719 1641 -717
rect 1647 -713 1648 -711
rect 1647 -719 1648 -717
rect 1657 -713 1658 -711
rect 1654 -719 1655 -717
rect 1661 -713 1662 -711
rect 1661 -719 1662 -717
rect 1668 -713 1669 -711
rect 1671 -713 1672 -711
rect 1671 -719 1672 -717
rect 1787 -713 1788 -711
rect 1787 -719 1788 -717
rect 1794 -713 1795 -711
rect 1794 -719 1795 -717
rect 1801 -713 1802 -711
rect 1801 -719 1802 -717
rect 1822 -713 1823 -711
rect 1822 -719 1823 -717
rect 1857 -713 1858 -711
rect 1857 -719 1858 -717
rect 9 -858 10 -856
rect 9 -864 10 -862
rect 16 -864 17 -862
rect 23 -858 24 -856
rect 23 -864 24 -862
rect 30 -858 31 -856
rect 30 -864 31 -862
rect 37 -858 38 -856
rect 37 -864 38 -862
rect 44 -858 45 -856
rect 47 -864 48 -862
rect 54 -858 55 -856
rect 51 -864 52 -862
rect 54 -864 55 -862
rect 58 -858 59 -856
rect 58 -864 59 -862
rect 65 -858 66 -856
rect 65 -864 66 -862
rect 72 -858 73 -856
rect 72 -864 73 -862
rect 79 -858 80 -856
rect 82 -858 83 -856
rect 79 -864 80 -862
rect 86 -858 87 -856
rect 86 -864 87 -862
rect 93 -858 94 -856
rect 93 -864 94 -862
rect 100 -858 101 -856
rect 100 -864 101 -862
rect 107 -858 108 -856
rect 107 -864 108 -862
rect 114 -858 115 -856
rect 114 -864 115 -862
rect 121 -858 122 -856
rect 124 -858 125 -856
rect 121 -864 122 -862
rect 128 -858 129 -856
rect 128 -864 129 -862
rect 135 -858 136 -856
rect 135 -864 136 -862
rect 142 -858 143 -856
rect 142 -864 143 -862
rect 149 -858 150 -856
rect 149 -864 150 -862
rect 156 -858 157 -856
rect 156 -864 157 -862
rect 163 -858 164 -856
rect 166 -858 167 -856
rect 163 -864 164 -862
rect 166 -864 167 -862
rect 170 -858 171 -856
rect 170 -864 171 -862
rect 177 -858 178 -856
rect 180 -858 181 -856
rect 177 -864 178 -862
rect 180 -864 181 -862
rect 184 -858 185 -856
rect 184 -864 185 -862
rect 191 -858 192 -856
rect 194 -864 195 -862
rect 198 -858 199 -856
rect 201 -858 202 -856
rect 198 -864 199 -862
rect 201 -864 202 -862
rect 205 -858 206 -856
rect 205 -864 206 -862
rect 212 -858 213 -856
rect 212 -864 213 -862
rect 219 -858 220 -856
rect 226 -858 227 -856
rect 226 -864 227 -862
rect 233 -858 234 -856
rect 233 -864 234 -862
rect 240 -858 241 -856
rect 240 -864 241 -862
rect 247 -858 248 -856
rect 247 -864 248 -862
rect 254 -858 255 -856
rect 254 -864 255 -862
rect 261 -858 262 -856
rect 261 -864 262 -862
rect 268 -858 269 -856
rect 268 -864 269 -862
rect 275 -858 276 -856
rect 275 -864 276 -862
rect 282 -858 283 -856
rect 282 -864 283 -862
rect 289 -858 290 -856
rect 289 -864 290 -862
rect 296 -858 297 -856
rect 296 -864 297 -862
rect 303 -858 304 -856
rect 310 -858 311 -856
rect 310 -864 311 -862
rect 317 -864 318 -862
rect 324 -858 325 -856
rect 324 -864 325 -862
rect 331 -858 332 -856
rect 331 -864 332 -862
rect 338 -858 339 -856
rect 338 -864 339 -862
rect 345 -858 346 -856
rect 345 -864 346 -862
rect 352 -858 353 -856
rect 352 -864 353 -862
rect 359 -858 360 -856
rect 359 -864 360 -862
rect 366 -858 367 -856
rect 366 -864 367 -862
rect 373 -858 374 -856
rect 373 -864 374 -862
rect 380 -858 381 -856
rect 380 -864 381 -862
rect 387 -858 388 -856
rect 387 -864 388 -862
rect 394 -858 395 -856
rect 394 -864 395 -862
rect 401 -858 402 -856
rect 401 -864 402 -862
rect 408 -858 409 -856
rect 408 -864 409 -862
rect 415 -858 416 -856
rect 415 -864 416 -862
rect 422 -858 423 -856
rect 422 -864 423 -862
rect 429 -858 430 -856
rect 429 -864 430 -862
rect 439 -858 440 -856
rect 436 -864 437 -862
rect 439 -864 440 -862
rect 443 -858 444 -856
rect 443 -864 444 -862
rect 450 -858 451 -856
rect 450 -864 451 -862
rect 457 -858 458 -856
rect 457 -864 458 -862
rect 464 -858 465 -856
rect 464 -864 465 -862
rect 471 -858 472 -856
rect 471 -864 472 -862
rect 478 -858 479 -856
rect 478 -864 479 -862
rect 485 -858 486 -856
rect 485 -864 486 -862
rect 492 -858 493 -856
rect 495 -858 496 -856
rect 492 -864 493 -862
rect 495 -864 496 -862
rect 499 -858 500 -856
rect 499 -864 500 -862
rect 506 -858 507 -856
rect 506 -864 507 -862
rect 513 -858 514 -856
rect 516 -858 517 -856
rect 513 -864 514 -862
rect 516 -864 517 -862
rect 520 -858 521 -856
rect 520 -864 521 -862
rect 527 -858 528 -856
rect 527 -864 528 -862
rect 534 -858 535 -856
rect 534 -864 535 -862
rect 541 -858 542 -856
rect 541 -864 542 -862
rect 548 -858 549 -856
rect 548 -864 549 -862
rect 555 -858 556 -856
rect 558 -858 559 -856
rect 558 -864 559 -862
rect 562 -858 563 -856
rect 562 -864 563 -862
rect 572 -858 573 -856
rect 569 -864 570 -862
rect 572 -864 573 -862
rect 576 -858 577 -856
rect 579 -858 580 -856
rect 576 -864 577 -862
rect 583 -858 584 -856
rect 586 -858 587 -856
rect 583 -864 584 -862
rect 586 -864 587 -862
rect 590 -858 591 -856
rect 590 -864 591 -862
rect 597 -858 598 -856
rect 597 -864 598 -862
rect 600 -864 601 -862
rect 604 -858 605 -856
rect 604 -864 605 -862
rect 611 -858 612 -856
rect 614 -858 615 -856
rect 611 -864 612 -862
rect 618 -858 619 -856
rect 621 -858 622 -856
rect 618 -864 619 -862
rect 621 -864 622 -862
rect 625 -858 626 -856
rect 628 -858 629 -856
rect 625 -864 626 -862
rect 628 -864 629 -862
rect 632 -858 633 -856
rect 632 -864 633 -862
rect 639 -858 640 -856
rect 639 -864 640 -862
rect 646 -858 647 -856
rect 646 -864 647 -862
rect 653 -858 654 -856
rect 653 -864 654 -862
rect 660 -858 661 -856
rect 660 -864 661 -862
rect 667 -858 668 -856
rect 667 -864 668 -862
rect 674 -858 675 -856
rect 674 -864 675 -862
rect 681 -858 682 -856
rect 681 -864 682 -862
rect 691 -858 692 -856
rect 688 -864 689 -862
rect 691 -864 692 -862
rect 695 -858 696 -856
rect 695 -864 696 -862
rect 702 -864 703 -862
rect 705 -864 706 -862
rect 709 -858 710 -856
rect 709 -864 710 -862
rect 716 -858 717 -856
rect 716 -864 717 -862
rect 723 -858 724 -856
rect 723 -864 724 -862
rect 730 -858 731 -856
rect 730 -864 731 -862
rect 737 -858 738 -856
rect 737 -864 738 -862
rect 744 -858 745 -856
rect 744 -864 745 -862
rect 751 -858 752 -856
rect 751 -864 752 -862
rect 761 -858 762 -856
rect 758 -864 759 -862
rect 761 -864 762 -862
rect 765 -858 766 -856
rect 765 -864 766 -862
rect 772 -858 773 -856
rect 772 -864 773 -862
rect 779 -858 780 -856
rect 782 -858 783 -856
rect 779 -864 780 -862
rect 782 -864 783 -862
rect 786 -858 787 -856
rect 789 -858 790 -856
rect 786 -864 787 -862
rect 789 -864 790 -862
rect 793 -858 794 -856
rect 793 -864 794 -862
rect 800 -858 801 -856
rect 803 -858 804 -856
rect 800 -864 801 -862
rect 807 -858 808 -856
rect 807 -864 808 -862
rect 814 -858 815 -856
rect 814 -864 815 -862
rect 821 -858 822 -856
rect 824 -858 825 -856
rect 821 -864 822 -862
rect 824 -864 825 -862
rect 828 -858 829 -856
rect 831 -858 832 -856
rect 828 -864 829 -862
rect 831 -864 832 -862
rect 835 -858 836 -856
rect 835 -864 836 -862
rect 842 -858 843 -856
rect 842 -864 843 -862
rect 849 -858 850 -856
rect 849 -864 850 -862
rect 856 -858 857 -856
rect 856 -864 857 -862
rect 863 -858 864 -856
rect 863 -864 864 -862
rect 870 -858 871 -856
rect 870 -864 871 -862
rect 877 -858 878 -856
rect 877 -864 878 -862
rect 884 -858 885 -856
rect 884 -864 885 -862
rect 891 -858 892 -856
rect 891 -864 892 -862
rect 898 -858 899 -856
rect 898 -864 899 -862
rect 905 -858 906 -856
rect 905 -864 906 -862
rect 912 -858 913 -856
rect 912 -864 913 -862
rect 919 -858 920 -856
rect 919 -864 920 -862
rect 922 -864 923 -862
rect 926 -858 927 -856
rect 926 -864 927 -862
rect 933 -858 934 -856
rect 933 -864 934 -862
rect 940 -858 941 -856
rect 940 -864 941 -862
rect 947 -858 948 -856
rect 947 -864 948 -862
rect 954 -858 955 -856
rect 954 -864 955 -862
rect 961 -858 962 -856
rect 961 -864 962 -862
rect 968 -858 969 -856
rect 968 -864 969 -862
rect 975 -864 976 -862
rect 982 -858 983 -856
rect 982 -864 983 -862
rect 989 -858 990 -856
rect 989 -864 990 -862
rect 996 -858 997 -856
rect 996 -864 997 -862
rect 1003 -858 1004 -856
rect 1003 -864 1004 -862
rect 1010 -858 1011 -856
rect 1010 -864 1011 -862
rect 1017 -858 1018 -856
rect 1017 -864 1018 -862
rect 1024 -858 1025 -856
rect 1024 -864 1025 -862
rect 1031 -858 1032 -856
rect 1034 -858 1035 -856
rect 1031 -864 1032 -862
rect 1034 -864 1035 -862
rect 1038 -858 1039 -856
rect 1038 -864 1039 -862
rect 1045 -858 1046 -856
rect 1045 -864 1046 -862
rect 1052 -858 1053 -856
rect 1052 -864 1053 -862
rect 1059 -858 1060 -856
rect 1059 -864 1060 -862
rect 1066 -858 1067 -856
rect 1066 -864 1067 -862
rect 1073 -858 1074 -856
rect 1073 -864 1074 -862
rect 1080 -858 1081 -856
rect 1080 -864 1081 -862
rect 1087 -858 1088 -856
rect 1087 -864 1088 -862
rect 1094 -858 1095 -856
rect 1094 -864 1095 -862
rect 1101 -858 1102 -856
rect 1101 -864 1102 -862
rect 1108 -858 1109 -856
rect 1108 -864 1109 -862
rect 1111 -864 1112 -862
rect 1115 -858 1116 -856
rect 1115 -864 1116 -862
rect 1122 -858 1123 -856
rect 1122 -864 1123 -862
rect 1129 -858 1130 -856
rect 1129 -864 1130 -862
rect 1136 -858 1137 -856
rect 1136 -864 1137 -862
rect 1143 -858 1144 -856
rect 1143 -864 1144 -862
rect 1150 -858 1151 -856
rect 1150 -864 1151 -862
rect 1157 -858 1158 -856
rect 1157 -864 1158 -862
rect 1164 -858 1165 -856
rect 1164 -864 1165 -862
rect 1171 -858 1172 -856
rect 1171 -864 1172 -862
rect 1178 -858 1179 -856
rect 1178 -864 1179 -862
rect 1185 -858 1186 -856
rect 1185 -864 1186 -862
rect 1192 -858 1193 -856
rect 1195 -858 1196 -856
rect 1192 -864 1193 -862
rect 1199 -858 1200 -856
rect 1199 -864 1200 -862
rect 1206 -858 1207 -856
rect 1206 -864 1207 -862
rect 1213 -858 1214 -856
rect 1213 -864 1214 -862
rect 1220 -858 1221 -856
rect 1220 -864 1221 -862
rect 1227 -858 1228 -856
rect 1227 -864 1228 -862
rect 1234 -858 1235 -856
rect 1234 -864 1235 -862
rect 1241 -858 1242 -856
rect 1241 -864 1242 -862
rect 1248 -858 1249 -856
rect 1248 -864 1249 -862
rect 1255 -858 1256 -856
rect 1255 -864 1256 -862
rect 1262 -858 1263 -856
rect 1262 -864 1263 -862
rect 1269 -858 1270 -856
rect 1269 -864 1270 -862
rect 1276 -858 1277 -856
rect 1276 -864 1277 -862
rect 1283 -858 1284 -856
rect 1283 -864 1284 -862
rect 1290 -858 1291 -856
rect 1290 -864 1291 -862
rect 1297 -858 1298 -856
rect 1297 -864 1298 -862
rect 1304 -858 1305 -856
rect 1304 -864 1305 -862
rect 1311 -858 1312 -856
rect 1311 -864 1312 -862
rect 1318 -858 1319 -856
rect 1318 -864 1319 -862
rect 1325 -858 1326 -856
rect 1325 -864 1326 -862
rect 1332 -858 1333 -856
rect 1332 -864 1333 -862
rect 1339 -858 1340 -856
rect 1339 -864 1340 -862
rect 1346 -858 1347 -856
rect 1346 -864 1347 -862
rect 1353 -858 1354 -856
rect 1353 -864 1354 -862
rect 1360 -858 1361 -856
rect 1360 -864 1361 -862
rect 1367 -858 1368 -856
rect 1367 -864 1368 -862
rect 1374 -858 1375 -856
rect 1374 -864 1375 -862
rect 1381 -858 1382 -856
rect 1381 -864 1382 -862
rect 1388 -858 1389 -856
rect 1388 -864 1389 -862
rect 1395 -858 1396 -856
rect 1395 -864 1396 -862
rect 1402 -858 1403 -856
rect 1402 -864 1403 -862
rect 1409 -858 1410 -856
rect 1409 -864 1410 -862
rect 1416 -858 1417 -856
rect 1416 -864 1417 -862
rect 1423 -858 1424 -856
rect 1423 -864 1424 -862
rect 1430 -858 1431 -856
rect 1430 -864 1431 -862
rect 1437 -858 1438 -856
rect 1437 -864 1438 -862
rect 1444 -858 1445 -856
rect 1444 -864 1445 -862
rect 1451 -858 1452 -856
rect 1451 -864 1452 -862
rect 1458 -858 1459 -856
rect 1458 -864 1459 -862
rect 1465 -858 1466 -856
rect 1465 -864 1466 -862
rect 1472 -858 1473 -856
rect 1472 -864 1473 -862
rect 1479 -858 1480 -856
rect 1479 -864 1480 -862
rect 1486 -858 1487 -856
rect 1486 -864 1487 -862
rect 1493 -858 1494 -856
rect 1493 -864 1494 -862
rect 1500 -858 1501 -856
rect 1500 -864 1501 -862
rect 1507 -858 1508 -856
rect 1507 -864 1508 -862
rect 1514 -858 1515 -856
rect 1514 -864 1515 -862
rect 1521 -858 1522 -856
rect 1521 -864 1522 -862
rect 1528 -858 1529 -856
rect 1528 -864 1529 -862
rect 1535 -858 1536 -856
rect 1535 -864 1536 -862
rect 1542 -858 1543 -856
rect 1542 -864 1543 -862
rect 1549 -858 1550 -856
rect 1549 -864 1550 -862
rect 1556 -858 1557 -856
rect 1556 -864 1557 -862
rect 1563 -858 1564 -856
rect 1563 -864 1564 -862
rect 1570 -858 1571 -856
rect 1570 -864 1571 -862
rect 1577 -858 1578 -856
rect 1577 -864 1578 -862
rect 1584 -858 1585 -856
rect 1584 -864 1585 -862
rect 1591 -858 1592 -856
rect 1591 -864 1592 -862
rect 1594 -864 1595 -862
rect 1598 -858 1599 -856
rect 1598 -864 1599 -862
rect 1605 -858 1606 -856
rect 1605 -864 1606 -862
rect 1612 -858 1613 -856
rect 1612 -864 1613 -862
rect 1619 -858 1620 -856
rect 1619 -864 1620 -862
rect 1626 -858 1627 -856
rect 1626 -864 1627 -862
rect 1633 -858 1634 -856
rect 1633 -864 1634 -862
rect 1640 -858 1641 -856
rect 1640 -864 1641 -862
rect 1647 -858 1648 -856
rect 1647 -864 1648 -862
rect 1654 -858 1655 -856
rect 1654 -864 1655 -862
rect 1661 -858 1662 -856
rect 1661 -864 1662 -862
rect 1668 -858 1669 -856
rect 1668 -864 1669 -862
rect 1675 -858 1676 -856
rect 1675 -864 1676 -862
rect 1682 -858 1683 -856
rect 1682 -864 1683 -862
rect 1689 -858 1690 -856
rect 1689 -864 1690 -862
rect 1696 -858 1697 -856
rect 1696 -864 1697 -862
rect 1703 -858 1704 -856
rect 1703 -864 1704 -862
rect 1710 -858 1711 -856
rect 1710 -864 1711 -862
rect 1717 -858 1718 -856
rect 1717 -864 1718 -862
rect 1724 -858 1725 -856
rect 1724 -864 1725 -862
rect 1731 -858 1732 -856
rect 1731 -864 1732 -862
rect 1738 -858 1739 -856
rect 1738 -864 1739 -862
rect 1745 -858 1746 -856
rect 1745 -864 1746 -862
rect 1752 -858 1753 -856
rect 1752 -864 1753 -862
rect 1759 -858 1760 -856
rect 1759 -864 1760 -862
rect 1766 -858 1767 -856
rect 1766 -864 1767 -862
rect 1773 -858 1774 -856
rect 1773 -864 1774 -862
rect 1780 -858 1781 -856
rect 1783 -858 1784 -856
rect 1780 -864 1781 -862
rect 1783 -864 1784 -862
rect 1787 -858 1788 -856
rect 1787 -864 1788 -862
rect 1794 -858 1795 -856
rect 1794 -864 1795 -862
rect 1801 -858 1802 -856
rect 1801 -864 1802 -862
rect 1808 -858 1809 -856
rect 1808 -864 1809 -862
rect 1818 -864 1819 -862
rect 1822 -858 1823 -856
rect 1822 -864 1823 -862
rect 1829 -858 1830 -856
rect 1829 -864 1830 -862
rect 1836 -858 1837 -856
rect 1836 -864 1837 -862
rect 1843 -858 1844 -856
rect 1843 -864 1844 -862
rect 1850 -858 1851 -856
rect 1850 -864 1851 -862
rect 1857 -858 1858 -856
rect 1857 -864 1858 -862
rect 1885 -858 1886 -856
rect 1885 -864 1886 -862
rect 1892 -858 1893 -856
rect 1892 -864 1893 -862
rect 2 -979 3 -977
rect 2 -985 3 -983
rect 9 -979 10 -977
rect 9 -985 10 -983
rect 16 -979 17 -977
rect 16 -985 17 -983
rect 23 -979 24 -977
rect 23 -985 24 -983
rect 30 -979 31 -977
rect 30 -985 31 -983
rect 37 -979 38 -977
rect 37 -985 38 -983
rect 44 -979 45 -977
rect 44 -985 45 -983
rect 51 -979 52 -977
rect 51 -985 52 -983
rect 58 -979 59 -977
rect 58 -985 59 -983
rect 65 -979 66 -977
rect 68 -979 69 -977
rect 65 -985 66 -983
rect 68 -985 69 -983
rect 72 -979 73 -977
rect 72 -985 73 -983
rect 79 -979 80 -977
rect 79 -985 80 -983
rect 86 -979 87 -977
rect 86 -985 87 -983
rect 93 -979 94 -977
rect 96 -985 97 -983
rect 100 -979 101 -977
rect 100 -985 101 -983
rect 107 -979 108 -977
rect 110 -979 111 -977
rect 110 -985 111 -983
rect 114 -979 115 -977
rect 114 -985 115 -983
rect 121 -979 122 -977
rect 121 -985 122 -983
rect 128 -979 129 -977
rect 128 -985 129 -983
rect 135 -979 136 -977
rect 135 -985 136 -983
rect 142 -979 143 -977
rect 142 -985 143 -983
rect 145 -985 146 -983
rect 149 -979 150 -977
rect 149 -985 150 -983
rect 156 -979 157 -977
rect 156 -985 157 -983
rect 159 -985 160 -983
rect 163 -979 164 -977
rect 163 -985 164 -983
rect 170 -979 171 -977
rect 170 -985 171 -983
rect 177 -979 178 -977
rect 177 -985 178 -983
rect 184 -979 185 -977
rect 187 -979 188 -977
rect 184 -985 185 -983
rect 191 -979 192 -977
rect 191 -985 192 -983
rect 198 -979 199 -977
rect 198 -985 199 -983
rect 205 -979 206 -977
rect 205 -985 206 -983
rect 212 -979 213 -977
rect 212 -985 213 -983
rect 219 -985 220 -983
rect 226 -979 227 -977
rect 226 -985 227 -983
rect 233 -979 234 -977
rect 236 -979 237 -977
rect 236 -985 237 -983
rect 240 -979 241 -977
rect 240 -985 241 -983
rect 247 -979 248 -977
rect 247 -985 248 -983
rect 254 -979 255 -977
rect 254 -985 255 -983
rect 261 -979 262 -977
rect 261 -985 262 -983
rect 268 -979 269 -977
rect 268 -985 269 -983
rect 275 -979 276 -977
rect 275 -985 276 -983
rect 282 -979 283 -977
rect 282 -985 283 -983
rect 289 -979 290 -977
rect 289 -985 290 -983
rect 296 -979 297 -977
rect 296 -985 297 -983
rect 303 -985 304 -983
rect 310 -979 311 -977
rect 310 -985 311 -983
rect 317 -979 318 -977
rect 317 -985 318 -983
rect 324 -979 325 -977
rect 324 -985 325 -983
rect 331 -979 332 -977
rect 331 -985 332 -983
rect 338 -979 339 -977
rect 338 -985 339 -983
rect 345 -979 346 -977
rect 345 -985 346 -983
rect 352 -979 353 -977
rect 352 -985 353 -983
rect 359 -979 360 -977
rect 359 -985 360 -983
rect 366 -979 367 -977
rect 366 -985 367 -983
rect 373 -979 374 -977
rect 373 -985 374 -983
rect 380 -979 381 -977
rect 380 -985 381 -983
rect 390 -979 391 -977
rect 387 -985 388 -983
rect 390 -985 391 -983
rect 394 -979 395 -977
rect 394 -985 395 -983
rect 401 -979 402 -977
rect 401 -985 402 -983
rect 408 -979 409 -977
rect 408 -985 409 -983
rect 415 -979 416 -977
rect 415 -985 416 -983
rect 422 -979 423 -977
rect 422 -985 423 -983
rect 429 -979 430 -977
rect 429 -985 430 -983
rect 436 -979 437 -977
rect 436 -985 437 -983
rect 443 -979 444 -977
rect 443 -985 444 -983
rect 450 -979 451 -977
rect 450 -985 451 -983
rect 457 -979 458 -977
rect 460 -979 461 -977
rect 457 -985 458 -983
rect 464 -979 465 -977
rect 464 -985 465 -983
rect 471 -979 472 -977
rect 471 -985 472 -983
rect 478 -979 479 -977
rect 478 -985 479 -983
rect 485 -979 486 -977
rect 485 -985 486 -983
rect 492 -979 493 -977
rect 492 -985 493 -983
rect 499 -979 500 -977
rect 499 -985 500 -983
rect 506 -979 507 -977
rect 506 -985 507 -983
rect 513 -979 514 -977
rect 513 -985 514 -983
rect 520 -979 521 -977
rect 520 -985 521 -983
rect 527 -979 528 -977
rect 527 -985 528 -983
rect 534 -979 535 -977
rect 537 -979 538 -977
rect 534 -985 535 -983
rect 537 -985 538 -983
rect 541 -979 542 -977
rect 544 -979 545 -977
rect 548 -979 549 -977
rect 548 -985 549 -983
rect 555 -979 556 -977
rect 555 -985 556 -983
rect 562 -979 563 -977
rect 562 -985 563 -983
rect 569 -979 570 -977
rect 569 -985 570 -983
rect 576 -979 577 -977
rect 576 -985 577 -983
rect 583 -979 584 -977
rect 583 -985 584 -983
rect 590 -979 591 -977
rect 590 -985 591 -983
rect 597 -979 598 -977
rect 597 -985 598 -983
rect 604 -979 605 -977
rect 604 -985 605 -983
rect 607 -985 608 -983
rect 611 -979 612 -977
rect 611 -985 612 -983
rect 618 -979 619 -977
rect 618 -985 619 -983
rect 625 -979 626 -977
rect 625 -985 626 -983
rect 632 -979 633 -977
rect 632 -985 633 -983
rect 639 -979 640 -977
rect 639 -985 640 -983
rect 646 -979 647 -977
rect 646 -985 647 -983
rect 653 -979 654 -977
rect 653 -985 654 -983
rect 660 -979 661 -977
rect 660 -985 661 -983
rect 667 -979 668 -977
rect 667 -985 668 -983
rect 674 -979 675 -977
rect 674 -985 675 -983
rect 684 -979 685 -977
rect 681 -985 682 -983
rect 684 -985 685 -983
rect 688 -979 689 -977
rect 688 -985 689 -983
rect 695 -979 696 -977
rect 695 -985 696 -983
rect 702 -979 703 -977
rect 702 -985 703 -983
rect 709 -979 710 -977
rect 709 -985 710 -983
rect 716 -979 717 -977
rect 716 -985 717 -983
rect 726 -979 727 -977
rect 723 -985 724 -983
rect 726 -985 727 -983
rect 730 -979 731 -977
rect 730 -985 731 -983
rect 740 -979 741 -977
rect 737 -985 738 -983
rect 740 -985 741 -983
rect 744 -979 745 -977
rect 747 -979 748 -977
rect 744 -985 745 -983
rect 747 -985 748 -983
rect 754 -979 755 -977
rect 751 -985 752 -983
rect 754 -985 755 -983
rect 758 -979 759 -977
rect 758 -985 759 -983
rect 765 -979 766 -977
rect 765 -985 766 -983
rect 772 -979 773 -977
rect 775 -979 776 -977
rect 772 -985 773 -983
rect 775 -985 776 -983
rect 779 -979 780 -977
rect 779 -985 780 -983
rect 786 -979 787 -977
rect 786 -985 787 -983
rect 793 -979 794 -977
rect 793 -985 794 -983
rect 800 -979 801 -977
rect 800 -985 801 -983
rect 807 -979 808 -977
rect 807 -985 808 -983
rect 814 -979 815 -977
rect 814 -985 815 -983
rect 821 -979 822 -977
rect 821 -985 822 -983
rect 828 -979 829 -977
rect 828 -985 829 -983
rect 835 -979 836 -977
rect 835 -985 836 -983
rect 842 -979 843 -977
rect 842 -985 843 -983
rect 849 -979 850 -977
rect 849 -985 850 -983
rect 856 -979 857 -977
rect 856 -985 857 -983
rect 863 -979 864 -977
rect 863 -985 864 -983
rect 870 -979 871 -977
rect 870 -985 871 -983
rect 877 -979 878 -977
rect 877 -985 878 -983
rect 884 -979 885 -977
rect 884 -985 885 -983
rect 891 -979 892 -977
rect 891 -985 892 -983
rect 898 -979 899 -977
rect 898 -985 899 -983
rect 905 -979 906 -977
rect 905 -985 906 -983
rect 915 -979 916 -977
rect 912 -985 913 -983
rect 915 -985 916 -983
rect 922 -979 923 -977
rect 919 -985 920 -983
rect 922 -985 923 -983
rect 926 -979 927 -977
rect 926 -985 927 -983
rect 933 -979 934 -977
rect 933 -985 934 -983
rect 940 -979 941 -977
rect 943 -979 944 -977
rect 940 -985 941 -983
rect 943 -985 944 -983
rect 947 -979 948 -977
rect 947 -985 948 -983
rect 954 -979 955 -977
rect 954 -985 955 -983
rect 961 -979 962 -977
rect 961 -985 962 -983
rect 968 -979 969 -977
rect 968 -985 969 -983
rect 975 -979 976 -977
rect 975 -985 976 -983
rect 982 -979 983 -977
rect 985 -979 986 -977
rect 982 -985 983 -983
rect 985 -985 986 -983
rect 989 -979 990 -977
rect 989 -985 990 -983
rect 996 -979 997 -977
rect 996 -985 997 -983
rect 1003 -979 1004 -977
rect 1006 -979 1007 -977
rect 1003 -985 1004 -983
rect 1006 -985 1007 -983
rect 1010 -979 1011 -977
rect 1013 -979 1014 -977
rect 1010 -985 1011 -983
rect 1013 -985 1014 -983
rect 1017 -979 1018 -977
rect 1017 -985 1018 -983
rect 1024 -979 1025 -977
rect 1024 -985 1025 -983
rect 1031 -979 1032 -977
rect 1034 -979 1035 -977
rect 1031 -985 1032 -983
rect 1034 -985 1035 -983
rect 1038 -979 1039 -977
rect 1041 -979 1042 -977
rect 1038 -985 1039 -983
rect 1041 -985 1042 -983
rect 1045 -979 1046 -977
rect 1045 -985 1046 -983
rect 1052 -979 1053 -977
rect 1052 -985 1053 -983
rect 1059 -979 1060 -977
rect 1062 -979 1063 -977
rect 1059 -985 1060 -983
rect 1062 -985 1063 -983
rect 1066 -979 1067 -977
rect 1066 -985 1067 -983
rect 1073 -979 1074 -977
rect 1073 -985 1074 -983
rect 1080 -979 1081 -977
rect 1083 -979 1084 -977
rect 1080 -985 1081 -983
rect 1083 -985 1084 -983
rect 1087 -979 1088 -977
rect 1087 -985 1088 -983
rect 1094 -979 1095 -977
rect 1094 -985 1095 -983
rect 1101 -979 1102 -977
rect 1101 -985 1102 -983
rect 1108 -979 1109 -977
rect 1111 -979 1112 -977
rect 1108 -985 1109 -983
rect 1115 -979 1116 -977
rect 1115 -985 1116 -983
rect 1122 -979 1123 -977
rect 1122 -985 1123 -983
rect 1129 -979 1130 -977
rect 1129 -985 1130 -983
rect 1136 -979 1137 -977
rect 1136 -985 1137 -983
rect 1143 -979 1144 -977
rect 1143 -985 1144 -983
rect 1153 -979 1154 -977
rect 1150 -985 1151 -983
rect 1153 -985 1154 -983
rect 1157 -979 1158 -977
rect 1160 -979 1161 -977
rect 1160 -985 1161 -983
rect 1164 -979 1165 -977
rect 1164 -985 1165 -983
rect 1171 -979 1172 -977
rect 1171 -985 1172 -983
rect 1178 -979 1179 -977
rect 1178 -985 1179 -983
rect 1185 -979 1186 -977
rect 1185 -985 1186 -983
rect 1192 -979 1193 -977
rect 1192 -985 1193 -983
rect 1199 -979 1200 -977
rect 1199 -985 1200 -983
rect 1206 -979 1207 -977
rect 1206 -985 1207 -983
rect 1213 -979 1214 -977
rect 1213 -985 1214 -983
rect 1220 -979 1221 -977
rect 1220 -985 1221 -983
rect 1227 -985 1228 -983
rect 1230 -985 1231 -983
rect 1234 -979 1235 -977
rect 1234 -985 1235 -983
rect 1241 -979 1242 -977
rect 1241 -985 1242 -983
rect 1248 -979 1249 -977
rect 1248 -985 1249 -983
rect 1255 -979 1256 -977
rect 1255 -985 1256 -983
rect 1262 -979 1263 -977
rect 1262 -985 1263 -983
rect 1269 -979 1270 -977
rect 1269 -985 1270 -983
rect 1276 -979 1277 -977
rect 1276 -985 1277 -983
rect 1283 -979 1284 -977
rect 1283 -985 1284 -983
rect 1290 -979 1291 -977
rect 1290 -985 1291 -983
rect 1297 -979 1298 -977
rect 1297 -985 1298 -983
rect 1304 -979 1305 -977
rect 1304 -985 1305 -983
rect 1311 -979 1312 -977
rect 1311 -985 1312 -983
rect 1318 -979 1319 -977
rect 1318 -985 1319 -983
rect 1325 -979 1326 -977
rect 1325 -985 1326 -983
rect 1332 -979 1333 -977
rect 1332 -985 1333 -983
rect 1339 -979 1340 -977
rect 1339 -985 1340 -983
rect 1346 -979 1347 -977
rect 1346 -985 1347 -983
rect 1353 -979 1354 -977
rect 1353 -985 1354 -983
rect 1360 -979 1361 -977
rect 1360 -985 1361 -983
rect 1367 -979 1368 -977
rect 1367 -985 1368 -983
rect 1374 -979 1375 -977
rect 1374 -985 1375 -983
rect 1381 -979 1382 -977
rect 1381 -985 1382 -983
rect 1388 -979 1389 -977
rect 1388 -985 1389 -983
rect 1395 -979 1396 -977
rect 1395 -985 1396 -983
rect 1402 -979 1403 -977
rect 1402 -985 1403 -983
rect 1409 -979 1410 -977
rect 1409 -985 1410 -983
rect 1416 -979 1417 -977
rect 1416 -985 1417 -983
rect 1423 -979 1424 -977
rect 1423 -985 1424 -983
rect 1430 -979 1431 -977
rect 1430 -985 1431 -983
rect 1437 -979 1438 -977
rect 1437 -985 1438 -983
rect 1444 -979 1445 -977
rect 1444 -985 1445 -983
rect 1451 -979 1452 -977
rect 1451 -985 1452 -983
rect 1458 -979 1459 -977
rect 1458 -985 1459 -983
rect 1465 -979 1466 -977
rect 1465 -985 1466 -983
rect 1472 -979 1473 -977
rect 1472 -985 1473 -983
rect 1479 -979 1480 -977
rect 1479 -985 1480 -983
rect 1486 -979 1487 -977
rect 1486 -985 1487 -983
rect 1493 -979 1494 -977
rect 1493 -985 1494 -983
rect 1500 -979 1501 -977
rect 1500 -985 1501 -983
rect 1507 -979 1508 -977
rect 1507 -985 1508 -983
rect 1514 -979 1515 -977
rect 1514 -985 1515 -983
rect 1521 -979 1522 -977
rect 1521 -985 1522 -983
rect 1528 -979 1529 -977
rect 1528 -985 1529 -983
rect 1535 -979 1536 -977
rect 1535 -985 1536 -983
rect 1542 -979 1543 -977
rect 1542 -985 1543 -983
rect 1549 -979 1550 -977
rect 1549 -985 1550 -983
rect 1556 -979 1557 -977
rect 1556 -985 1557 -983
rect 1563 -979 1564 -977
rect 1563 -985 1564 -983
rect 1570 -979 1571 -977
rect 1570 -985 1571 -983
rect 1577 -979 1578 -977
rect 1577 -985 1578 -983
rect 1584 -979 1585 -977
rect 1584 -985 1585 -983
rect 1591 -979 1592 -977
rect 1594 -979 1595 -977
rect 1591 -985 1592 -983
rect 1598 -979 1599 -977
rect 1598 -985 1599 -983
rect 1605 -979 1606 -977
rect 1605 -985 1606 -983
rect 1612 -979 1613 -977
rect 1612 -985 1613 -983
rect 1619 -979 1620 -977
rect 1619 -985 1620 -983
rect 1626 -979 1627 -977
rect 1626 -985 1627 -983
rect 1633 -979 1634 -977
rect 1633 -985 1634 -983
rect 1640 -979 1641 -977
rect 1640 -985 1641 -983
rect 1647 -979 1648 -977
rect 1647 -985 1648 -983
rect 1654 -979 1655 -977
rect 1654 -985 1655 -983
rect 1661 -979 1662 -977
rect 1661 -985 1662 -983
rect 1668 -979 1669 -977
rect 1668 -985 1669 -983
rect 1675 -979 1676 -977
rect 1675 -985 1676 -983
rect 1682 -979 1683 -977
rect 1682 -985 1683 -983
rect 1689 -979 1690 -977
rect 1689 -985 1690 -983
rect 1696 -979 1697 -977
rect 1696 -985 1697 -983
rect 1703 -979 1704 -977
rect 1703 -985 1704 -983
rect 1710 -979 1711 -977
rect 1710 -985 1711 -983
rect 1717 -979 1718 -977
rect 1717 -985 1718 -983
rect 1724 -979 1725 -977
rect 1724 -985 1725 -983
rect 1731 -979 1732 -977
rect 1731 -985 1732 -983
rect 1738 -979 1739 -977
rect 1738 -985 1739 -983
rect 1745 -979 1746 -977
rect 1745 -985 1746 -983
rect 1752 -979 1753 -977
rect 1752 -985 1753 -983
rect 1759 -979 1760 -977
rect 1759 -985 1760 -983
rect 1766 -979 1767 -977
rect 1766 -985 1767 -983
rect 1773 -979 1774 -977
rect 1773 -985 1774 -983
rect 1780 -979 1781 -977
rect 1780 -985 1781 -983
rect 1787 -979 1788 -977
rect 1787 -985 1788 -983
rect 1794 -979 1795 -977
rect 1794 -985 1795 -983
rect 1801 -979 1802 -977
rect 1801 -985 1802 -983
rect 1808 -979 1809 -977
rect 1808 -985 1809 -983
rect 1815 -979 1816 -977
rect 1815 -985 1816 -983
rect 1822 -979 1823 -977
rect 1822 -985 1823 -983
rect 1829 -979 1830 -977
rect 1829 -985 1830 -983
rect 1836 -979 1837 -977
rect 1836 -985 1837 -983
rect 1843 -979 1844 -977
rect 1843 -985 1844 -983
rect 1850 -979 1851 -977
rect 1850 -985 1851 -983
rect 1857 -979 1858 -977
rect 1857 -985 1858 -983
rect 1864 -979 1865 -977
rect 1864 -985 1865 -983
rect 1871 -979 1872 -977
rect 1871 -985 1872 -983
rect 1878 -979 1879 -977
rect 1881 -979 1882 -977
rect 1878 -985 1879 -983
rect 1881 -985 1882 -983
rect 1885 -979 1886 -977
rect 1885 -985 1886 -983
rect 1892 -979 1893 -977
rect 1892 -985 1893 -983
rect 1899 -979 1900 -977
rect 1899 -985 1900 -983
rect 1902 -985 1903 -983
rect 1906 -979 1907 -977
rect 1906 -985 1907 -983
rect 1913 -979 1914 -977
rect 1916 -979 1917 -977
rect 1920 -979 1921 -977
rect 1920 -985 1921 -983
rect 1927 -979 1928 -977
rect 1927 -985 1928 -983
rect 1934 -979 1935 -977
rect 1934 -985 1935 -983
rect 1941 -979 1942 -977
rect 1941 -985 1942 -983
rect 1948 -979 1949 -977
rect 1948 -985 1949 -983
rect 1955 -979 1956 -977
rect 1955 -985 1956 -983
rect 9 -1110 10 -1108
rect 9 -1116 10 -1114
rect 16 -1110 17 -1108
rect 16 -1116 17 -1114
rect 23 -1110 24 -1108
rect 23 -1116 24 -1114
rect 30 -1110 31 -1108
rect 30 -1116 31 -1114
rect 37 -1110 38 -1108
rect 37 -1116 38 -1114
rect 47 -1110 48 -1108
rect 44 -1116 45 -1114
rect 47 -1116 48 -1114
rect 51 -1110 52 -1108
rect 51 -1116 52 -1114
rect 58 -1110 59 -1108
rect 58 -1116 59 -1114
rect 65 -1110 66 -1108
rect 68 -1110 69 -1108
rect 65 -1116 66 -1114
rect 72 -1110 73 -1108
rect 72 -1116 73 -1114
rect 79 -1110 80 -1108
rect 82 -1110 83 -1108
rect 82 -1116 83 -1114
rect 86 -1110 87 -1108
rect 86 -1116 87 -1114
rect 93 -1110 94 -1108
rect 93 -1116 94 -1114
rect 100 -1110 101 -1108
rect 100 -1116 101 -1114
rect 107 -1110 108 -1108
rect 107 -1116 108 -1114
rect 114 -1110 115 -1108
rect 114 -1116 115 -1114
rect 121 -1110 122 -1108
rect 121 -1116 122 -1114
rect 128 -1110 129 -1108
rect 128 -1116 129 -1114
rect 131 -1116 132 -1114
rect 135 -1110 136 -1108
rect 135 -1116 136 -1114
rect 142 -1110 143 -1108
rect 142 -1116 143 -1114
rect 149 -1110 150 -1108
rect 149 -1116 150 -1114
rect 156 -1110 157 -1108
rect 156 -1116 157 -1114
rect 163 -1110 164 -1108
rect 163 -1116 164 -1114
rect 170 -1110 171 -1108
rect 170 -1116 171 -1114
rect 177 -1110 178 -1108
rect 177 -1116 178 -1114
rect 184 -1110 185 -1108
rect 184 -1116 185 -1114
rect 191 -1110 192 -1108
rect 191 -1116 192 -1114
rect 198 -1110 199 -1108
rect 198 -1116 199 -1114
rect 205 -1110 206 -1108
rect 205 -1116 206 -1114
rect 212 -1110 213 -1108
rect 215 -1110 216 -1108
rect 212 -1116 213 -1114
rect 219 -1110 220 -1108
rect 222 -1116 223 -1114
rect 226 -1110 227 -1108
rect 226 -1116 227 -1114
rect 233 -1110 234 -1108
rect 233 -1116 234 -1114
rect 240 -1110 241 -1108
rect 240 -1116 241 -1114
rect 247 -1110 248 -1108
rect 247 -1116 248 -1114
rect 254 -1110 255 -1108
rect 254 -1116 255 -1114
rect 261 -1110 262 -1108
rect 261 -1116 262 -1114
rect 268 -1110 269 -1108
rect 268 -1116 269 -1114
rect 275 -1110 276 -1108
rect 275 -1116 276 -1114
rect 282 -1110 283 -1108
rect 282 -1116 283 -1114
rect 289 -1110 290 -1108
rect 289 -1116 290 -1114
rect 296 -1110 297 -1108
rect 296 -1116 297 -1114
rect 303 -1110 304 -1108
rect 303 -1116 304 -1114
rect 310 -1110 311 -1108
rect 313 -1116 314 -1114
rect 317 -1110 318 -1108
rect 317 -1116 318 -1114
rect 324 -1110 325 -1108
rect 324 -1116 325 -1114
rect 331 -1110 332 -1108
rect 331 -1116 332 -1114
rect 338 -1110 339 -1108
rect 338 -1116 339 -1114
rect 345 -1110 346 -1108
rect 345 -1116 346 -1114
rect 352 -1110 353 -1108
rect 352 -1116 353 -1114
rect 359 -1110 360 -1108
rect 359 -1116 360 -1114
rect 366 -1110 367 -1108
rect 366 -1116 367 -1114
rect 373 -1110 374 -1108
rect 373 -1116 374 -1114
rect 380 -1110 381 -1108
rect 380 -1116 381 -1114
rect 387 -1110 388 -1108
rect 394 -1110 395 -1108
rect 397 -1110 398 -1108
rect 394 -1116 395 -1114
rect 401 -1110 402 -1108
rect 401 -1116 402 -1114
rect 408 -1110 409 -1108
rect 408 -1116 409 -1114
rect 415 -1110 416 -1108
rect 415 -1116 416 -1114
rect 422 -1110 423 -1108
rect 422 -1116 423 -1114
rect 429 -1110 430 -1108
rect 429 -1116 430 -1114
rect 436 -1110 437 -1108
rect 436 -1116 437 -1114
rect 443 -1110 444 -1108
rect 443 -1116 444 -1114
rect 450 -1110 451 -1108
rect 453 -1110 454 -1108
rect 450 -1116 451 -1114
rect 453 -1116 454 -1114
rect 457 -1110 458 -1108
rect 457 -1116 458 -1114
rect 464 -1110 465 -1108
rect 464 -1116 465 -1114
rect 471 -1110 472 -1108
rect 471 -1116 472 -1114
rect 478 -1110 479 -1108
rect 478 -1116 479 -1114
rect 485 -1110 486 -1108
rect 485 -1116 486 -1114
rect 492 -1110 493 -1108
rect 492 -1116 493 -1114
rect 499 -1110 500 -1108
rect 499 -1116 500 -1114
rect 506 -1110 507 -1108
rect 506 -1116 507 -1114
rect 513 -1110 514 -1108
rect 513 -1116 514 -1114
rect 520 -1110 521 -1108
rect 520 -1116 521 -1114
rect 523 -1116 524 -1114
rect 527 -1110 528 -1108
rect 527 -1116 528 -1114
rect 534 -1110 535 -1108
rect 534 -1116 535 -1114
rect 541 -1110 542 -1108
rect 541 -1116 542 -1114
rect 548 -1110 549 -1108
rect 548 -1116 549 -1114
rect 555 -1110 556 -1108
rect 555 -1116 556 -1114
rect 565 -1110 566 -1108
rect 562 -1116 563 -1114
rect 565 -1116 566 -1114
rect 569 -1110 570 -1108
rect 572 -1110 573 -1108
rect 569 -1116 570 -1114
rect 572 -1116 573 -1114
rect 576 -1110 577 -1108
rect 579 -1110 580 -1108
rect 576 -1116 577 -1114
rect 579 -1116 580 -1114
rect 583 -1110 584 -1108
rect 583 -1116 584 -1114
rect 590 -1110 591 -1108
rect 590 -1116 591 -1114
rect 597 -1110 598 -1108
rect 597 -1116 598 -1114
rect 604 -1110 605 -1108
rect 604 -1116 605 -1114
rect 611 -1110 612 -1108
rect 611 -1116 612 -1114
rect 618 -1110 619 -1108
rect 618 -1116 619 -1114
rect 625 -1110 626 -1108
rect 628 -1110 629 -1108
rect 625 -1116 626 -1114
rect 628 -1116 629 -1114
rect 632 -1110 633 -1108
rect 635 -1110 636 -1108
rect 632 -1116 633 -1114
rect 639 -1110 640 -1108
rect 639 -1116 640 -1114
rect 646 -1110 647 -1108
rect 649 -1110 650 -1108
rect 646 -1116 647 -1114
rect 653 -1110 654 -1108
rect 656 -1110 657 -1108
rect 653 -1116 654 -1114
rect 656 -1116 657 -1114
rect 660 -1110 661 -1108
rect 660 -1116 661 -1114
rect 667 -1110 668 -1108
rect 667 -1116 668 -1114
rect 674 -1110 675 -1108
rect 674 -1116 675 -1114
rect 681 -1110 682 -1108
rect 684 -1110 685 -1108
rect 681 -1116 682 -1114
rect 684 -1116 685 -1114
rect 688 -1110 689 -1108
rect 688 -1116 689 -1114
rect 695 -1110 696 -1108
rect 695 -1116 696 -1114
rect 702 -1110 703 -1108
rect 702 -1116 703 -1114
rect 709 -1110 710 -1108
rect 709 -1116 710 -1114
rect 716 -1110 717 -1108
rect 716 -1116 717 -1114
rect 723 -1110 724 -1108
rect 723 -1116 724 -1114
rect 730 -1110 731 -1108
rect 733 -1110 734 -1108
rect 730 -1116 731 -1114
rect 733 -1116 734 -1114
rect 737 -1110 738 -1108
rect 740 -1110 741 -1108
rect 737 -1116 738 -1114
rect 740 -1116 741 -1114
rect 744 -1110 745 -1108
rect 744 -1116 745 -1114
rect 747 -1116 748 -1114
rect 751 -1110 752 -1108
rect 751 -1116 752 -1114
rect 754 -1116 755 -1114
rect 758 -1110 759 -1108
rect 761 -1110 762 -1108
rect 761 -1116 762 -1114
rect 765 -1110 766 -1108
rect 765 -1116 766 -1114
rect 772 -1110 773 -1108
rect 772 -1116 773 -1114
rect 779 -1110 780 -1108
rect 782 -1110 783 -1108
rect 779 -1116 780 -1114
rect 782 -1116 783 -1114
rect 786 -1110 787 -1108
rect 789 -1110 790 -1108
rect 789 -1116 790 -1114
rect 793 -1110 794 -1108
rect 793 -1116 794 -1114
rect 800 -1110 801 -1108
rect 800 -1116 801 -1114
rect 807 -1110 808 -1108
rect 807 -1116 808 -1114
rect 814 -1110 815 -1108
rect 814 -1116 815 -1114
rect 821 -1110 822 -1108
rect 821 -1116 822 -1114
rect 828 -1110 829 -1108
rect 828 -1116 829 -1114
rect 835 -1110 836 -1108
rect 835 -1116 836 -1114
rect 842 -1110 843 -1108
rect 842 -1116 843 -1114
rect 849 -1110 850 -1108
rect 849 -1116 850 -1114
rect 852 -1116 853 -1114
rect 856 -1110 857 -1108
rect 856 -1116 857 -1114
rect 863 -1110 864 -1108
rect 866 -1110 867 -1108
rect 863 -1116 864 -1114
rect 866 -1116 867 -1114
rect 870 -1110 871 -1108
rect 870 -1116 871 -1114
rect 877 -1110 878 -1108
rect 877 -1116 878 -1114
rect 884 -1110 885 -1108
rect 884 -1116 885 -1114
rect 891 -1110 892 -1108
rect 894 -1110 895 -1108
rect 891 -1116 892 -1114
rect 894 -1116 895 -1114
rect 898 -1110 899 -1108
rect 898 -1116 899 -1114
rect 905 -1110 906 -1108
rect 905 -1116 906 -1114
rect 912 -1110 913 -1108
rect 912 -1116 913 -1114
rect 919 -1110 920 -1108
rect 919 -1116 920 -1114
rect 926 -1110 927 -1108
rect 926 -1116 927 -1114
rect 933 -1110 934 -1108
rect 933 -1116 934 -1114
rect 940 -1110 941 -1108
rect 940 -1116 941 -1114
rect 947 -1110 948 -1108
rect 947 -1116 948 -1114
rect 954 -1110 955 -1108
rect 957 -1110 958 -1108
rect 954 -1116 955 -1114
rect 957 -1116 958 -1114
rect 961 -1110 962 -1108
rect 961 -1116 962 -1114
rect 968 -1110 969 -1108
rect 968 -1116 969 -1114
rect 975 -1110 976 -1108
rect 975 -1116 976 -1114
rect 982 -1110 983 -1108
rect 982 -1116 983 -1114
rect 989 -1110 990 -1108
rect 989 -1116 990 -1114
rect 996 -1110 997 -1108
rect 996 -1116 997 -1114
rect 1003 -1110 1004 -1108
rect 1003 -1116 1004 -1114
rect 1010 -1110 1011 -1108
rect 1010 -1116 1011 -1114
rect 1017 -1110 1018 -1108
rect 1020 -1110 1021 -1108
rect 1017 -1116 1018 -1114
rect 1020 -1116 1021 -1114
rect 1024 -1110 1025 -1108
rect 1024 -1116 1025 -1114
rect 1031 -1110 1032 -1108
rect 1031 -1116 1032 -1114
rect 1038 -1110 1039 -1108
rect 1038 -1116 1039 -1114
rect 1045 -1110 1046 -1108
rect 1048 -1110 1049 -1108
rect 1045 -1116 1046 -1114
rect 1048 -1116 1049 -1114
rect 1052 -1110 1053 -1108
rect 1052 -1116 1053 -1114
rect 1059 -1110 1060 -1108
rect 1059 -1116 1060 -1114
rect 1066 -1110 1067 -1108
rect 1066 -1116 1067 -1114
rect 1073 -1110 1074 -1108
rect 1073 -1116 1074 -1114
rect 1080 -1110 1081 -1108
rect 1080 -1116 1081 -1114
rect 1087 -1110 1088 -1108
rect 1087 -1116 1088 -1114
rect 1094 -1110 1095 -1108
rect 1094 -1116 1095 -1114
rect 1101 -1110 1102 -1108
rect 1101 -1116 1102 -1114
rect 1108 -1110 1109 -1108
rect 1108 -1116 1109 -1114
rect 1115 -1110 1116 -1108
rect 1115 -1116 1116 -1114
rect 1122 -1110 1123 -1108
rect 1122 -1116 1123 -1114
rect 1129 -1110 1130 -1108
rect 1129 -1116 1130 -1114
rect 1136 -1110 1137 -1108
rect 1139 -1110 1140 -1108
rect 1136 -1116 1137 -1114
rect 1139 -1116 1140 -1114
rect 1143 -1110 1144 -1108
rect 1143 -1116 1144 -1114
rect 1150 -1110 1151 -1108
rect 1153 -1110 1154 -1108
rect 1153 -1116 1154 -1114
rect 1157 -1110 1158 -1108
rect 1157 -1116 1158 -1114
rect 1164 -1110 1165 -1108
rect 1164 -1116 1165 -1114
rect 1171 -1110 1172 -1108
rect 1171 -1116 1172 -1114
rect 1178 -1110 1179 -1108
rect 1178 -1116 1179 -1114
rect 1185 -1110 1186 -1108
rect 1185 -1116 1186 -1114
rect 1192 -1110 1193 -1108
rect 1192 -1116 1193 -1114
rect 1199 -1110 1200 -1108
rect 1199 -1116 1200 -1114
rect 1206 -1110 1207 -1108
rect 1206 -1116 1207 -1114
rect 1213 -1110 1214 -1108
rect 1213 -1116 1214 -1114
rect 1220 -1110 1221 -1108
rect 1220 -1116 1221 -1114
rect 1227 -1110 1228 -1108
rect 1230 -1110 1231 -1108
rect 1230 -1116 1231 -1114
rect 1234 -1110 1235 -1108
rect 1234 -1116 1235 -1114
rect 1241 -1110 1242 -1108
rect 1241 -1116 1242 -1114
rect 1248 -1110 1249 -1108
rect 1248 -1116 1249 -1114
rect 1255 -1110 1256 -1108
rect 1255 -1116 1256 -1114
rect 1262 -1110 1263 -1108
rect 1262 -1116 1263 -1114
rect 1269 -1110 1270 -1108
rect 1269 -1116 1270 -1114
rect 1276 -1110 1277 -1108
rect 1276 -1116 1277 -1114
rect 1283 -1110 1284 -1108
rect 1283 -1116 1284 -1114
rect 1290 -1110 1291 -1108
rect 1290 -1116 1291 -1114
rect 1297 -1110 1298 -1108
rect 1297 -1116 1298 -1114
rect 1304 -1110 1305 -1108
rect 1304 -1116 1305 -1114
rect 1311 -1110 1312 -1108
rect 1311 -1116 1312 -1114
rect 1318 -1110 1319 -1108
rect 1318 -1116 1319 -1114
rect 1325 -1110 1326 -1108
rect 1325 -1116 1326 -1114
rect 1332 -1110 1333 -1108
rect 1332 -1116 1333 -1114
rect 1339 -1110 1340 -1108
rect 1339 -1116 1340 -1114
rect 1346 -1110 1347 -1108
rect 1346 -1116 1347 -1114
rect 1353 -1110 1354 -1108
rect 1353 -1116 1354 -1114
rect 1360 -1110 1361 -1108
rect 1360 -1116 1361 -1114
rect 1367 -1110 1368 -1108
rect 1367 -1116 1368 -1114
rect 1374 -1110 1375 -1108
rect 1374 -1116 1375 -1114
rect 1381 -1110 1382 -1108
rect 1381 -1116 1382 -1114
rect 1388 -1110 1389 -1108
rect 1388 -1116 1389 -1114
rect 1395 -1110 1396 -1108
rect 1395 -1116 1396 -1114
rect 1402 -1110 1403 -1108
rect 1402 -1116 1403 -1114
rect 1409 -1110 1410 -1108
rect 1409 -1116 1410 -1114
rect 1416 -1110 1417 -1108
rect 1416 -1116 1417 -1114
rect 1423 -1110 1424 -1108
rect 1423 -1116 1424 -1114
rect 1430 -1110 1431 -1108
rect 1430 -1116 1431 -1114
rect 1437 -1110 1438 -1108
rect 1437 -1116 1438 -1114
rect 1444 -1110 1445 -1108
rect 1444 -1116 1445 -1114
rect 1451 -1110 1452 -1108
rect 1451 -1116 1452 -1114
rect 1458 -1110 1459 -1108
rect 1458 -1116 1459 -1114
rect 1465 -1110 1466 -1108
rect 1465 -1116 1466 -1114
rect 1472 -1110 1473 -1108
rect 1472 -1116 1473 -1114
rect 1479 -1110 1480 -1108
rect 1479 -1116 1480 -1114
rect 1486 -1110 1487 -1108
rect 1486 -1116 1487 -1114
rect 1493 -1110 1494 -1108
rect 1493 -1116 1494 -1114
rect 1500 -1110 1501 -1108
rect 1500 -1116 1501 -1114
rect 1507 -1110 1508 -1108
rect 1507 -1116 1508 -1114
rect 1514 -1110 1515 -1108
rect 1514 -1116 1515 -1114
rect 1521 -1110 1522 -1108
rect 1521 -1116 1522 -1114
rect 1528 -1110 1529 -1108
rect 1528 -1116 1529 -1114
rect 1535 -1110 1536 -1108
rect 1535 -1116 1536 -1114
rect 1542 -1110 1543 -1108
rect 1542 -1116 1543 -1114
rect 1549 -1110 1550 -1108
rect 1549 -1116 1550 -1114
rect 1556 -1110 1557 -1108
rect 1556 -1116 1557 -1114
rect 1563 -1110 1564 -1108
rect 1563 -1116 1564 -1114
rect 1570 -1110 1571 -1108
rect 1570 -1116 1571 -1114
rect 1577 -1110 1578 -1108
rect 1577 -1116 1578 -1114
rect 1584 -1110 1585 -1108
rect 1584 -1116 1585 -1114
rect 1591 -1110 1592 -1108
rect 1591 -1116 1592 -1114
rect 1598 -1110 1599 -1108
rect 1598 -1116 1599 -1114
rect 1605 -1110 1606 -1108
rect 1605 -1116 1606 -1114
rect 1612 -1110 1613 -1108
rect 1612 -1116 1613 -1114
rect 1619 -1110 1620 -1108
rect 1619 -1116 1620 -1114
rect 1626 -1110 1627 -1108
rect 1626 -1116 1627 -1114
rect 1633 -1110 1634 -1108
rect 1633 -1116 1634 -1114
rect 1640 -1110 1641 -1108
rect 1640 -1116 1641 -1114
rect 1647 -1110 1648 -1108
rect 1647 -1116 1648 -1114
rect 1654 -1110 1655 -1108
rect 1654 -1116 1655 -1114
rect 1661 -1110 1662 -1108
rect 1661 -1116 1662 -1114
rect 1668 -1110 1669 -1108
rect 1668 -1116 1669 -1114
rect 1675 -1110 1676 -1108
rect 1675 -1116 1676 -1114
rect 1682 -1110 1683 -1108
rect 1682 -1116 1683 -1114
rect 1689 -1110 1690 -1108
rect 1689 -1116 1690 -1114
rect 1696 -1110 1697 -1108
rect 1696 -1116 1697 -1114
rect 1703 -1110 1704 -1108
rect 1703 -1116 1704 -1114
rect 1710 -1110 1711 -1108
rect 1710 -1116 1711 -1114
rect 1717 -1110 1718 -1108
rect 1717 -1116 1718 -1114
rect 1724 -1110 1725 -1108
rect 1724 -1116 1725 -1114
rect 1731 -1110 1732 -1108
rect 1731 -1116 1732 -1114
rect 1738 -1110 1739 -1108
rect 1738 -1116 1739 -1114
rect 1745 -1110 1746 -1108
rect 1745 -1116 1746 -1114
rect 1752 -1110 1753 -1108
rect 1752 -1116 1753 -1114
rect 1759 -1110 1760 -1108
rect 1759 -1116 1760 -1114
rect 1766 -1110 1767 -1108
rect 1766 -1116 1767 -1114
rect 1773 -1110 1774 -1108
rect 1773 -1116 1774 -1114
rect 1780 -1110 1781 -1108
rect 1780 -1116 1781 -1114
rect 1787 -1110 1788 -1108
rect 1787 -1116 1788 -1114
rect 1794 -1110 1795 -1108
rect 1794 -1116 1795 -1114
rect 1801 -1110 1802 -1108
rect 1801 -1116 1802 -1114
rect 1808 -1110 1809 -1108
rect 1808 -1116 1809 -1114
rect 1815 -1110 1816 -1108
rect 1815 -1116 1816 -1114
rect 1822 -1110 1823 -1108
rect 1822 -1116 1823 -1114
rect 1829 -1110 1830 -1108
rect 1829 -1116 1830 -1114
rect 1836 -1110 1837 -1108
rect 1836 -1116 1837 -1114
rect 1843 -1110 1844 -1108
rect 1843 -1116 1844 -1114
rect 1850 -1110 1851 -1108
rect 1850 -1116 1851 -1114
rect 1857 -1110 1858 -1108
rect 1857 -1116 1858 -1114
rect 1867 -1110 1868 -1108
rect 1864 -1116 1865 -1114
rect 1867 -1116 1868 -1114
rect 1871 -1110 1872 -1108
rect 1871 -1116 1872 -1114
rect 1878 -1110 1879 -1108
rect 1878 -1116 1879 -1114
rect 1927 -1110 1928 -1108
rect 1927 -1116 1928 -1114
rect 1948 -1110 1949 -1108
rect 1948 -1116 1949 -1114
rect 1962 -1110 1963 -1108
rect 1962 -1116 1963 -1114
rect 1969 -1110 1970 -1108
rect 1969 -1116 1970 -1114
rect 1976 -1110 1977 -1108
rect 1976 -1116 1977 -1114
rect 2 -1245 3 -1243
rect 2 -1251 3 -1249
rect 9 -1245 10 -1243
rect 9 -1251 10 -1249
rect 16 -1245 17 -1243
rect 16 -1251 17 -1249
rect 30 -1245 31 -1243
rect 30 -1251 31 -1249
rect 37 -1245 38 -1243
rect 40 -1245 41 -1243
rect 40 -1251 41 -1249
rect 44 -1245 45 -1243
rect 44 -1251 45 -1249
rect 51 -1245 52 -1243
rect 51 -1251 52 -1249
rect 58 -1245 59 -1243
rect 61 -1245 62 -1243
rect 58 -1251 59 -1249
rect 61 -1251 62 -1249
rect 65 -1245 66 -1243
rect 65 -1251 66 -1249
rect 72 -1245 73 -1243
rect 72 -1251 73 -1249
rect 79 -1245 80 -1243
rect 82 -1245 83 -1243
rect 79 -1251 80 -1249
rect 82 -1251 83 -1249
rect 86 -1245 87 -1243
rect 86 -1251 87 -1249
rect 93 -1245 94 -1243
rect 93 -1251 94 -1249
rect 100 -1245 101 -1243
rect 100 -1251 101 -1249
rect 107 -1245 108 -1243
rect 107 -1251 108 -1249
rect 114 -1245 115 -1243
rect 114 -1251 115 -1249
rect 121 -1245 122 -1243
rect 124 -1245 125 -1243
rect 124 -1251 125 -1249
rect 128 -1245 129 -1243
rect 128 -1251 129 -1249
rect 135 -1245 136 -1243
rect 135 -1251 136 -1249
rect 142 -1245 143 -1243
rect 142 -1251 143 -1249
rect 149 -1245 150 -1243
rect 149 -1251 150 -1249
rect 159 -1245 160 -1243
rect 156 -1251 157 -1249
rect 159 -1251 160 -1249
rect 163 -1245 164 -1243
rect 163 -1251 164 -1249
rect 170 -1245 171 -1243
rect 170 -1251 171 -1249
rect 173 -1251 174 -1249
rect 177 -1245 178 -1243
rect 180 -1245 181 -1243
rect 177 -1251 178 -1249
rect 180 -1251 181 -1249
rect 184 -1245 185 -1243
rect 184 -1251 185 -1249
rect 191 -1245 192 -1243
rect 191 -1251 192 -1249
rect 198 -1245 199 -1243
rect 198 -1251 199 -1249
rect 205 -1245 206 -1243
rect 205 -1251 206 -1249
rect 212 -1245 213 -1243
rect 212 -1251 213 -1249
rect 219 -1245 220 -1243
rect 219 -1251 220 -1249
rect 229 -1245 230 -1243
rect 226 -1251 227 -1249
rect 229 -1251 230 -1249
rect 233 -1245 234 -1243
rect 233 -1251 234 -1249
rect 240 -1245 241 -1243
rect 240 -1251 241 -1249
rect 247 -1245 248 -1243
rect 247 -1251 248 -1249
rect 254 -1245 255 -1243
rect 254 -1251 255 -1249
rect 261 -1251 262 -1249
rect 264 -1251 265 -1249
rect 268 -1245 269 -1243
rect 268 -1251 269 -1249
rect 275 -1245 276 -1243
rect 275 -1251 276 -1249
rect 282 -1245 283 -1243
rect 282 -1251 283 -1249
rect 289 -1245 290 -1243
rect 292 -1245 293 -1243
rect 296 -1245 297 -1243
rect 296 -1251 297 -1249
rect 303 -1245 304 -1243
rect 303 -1251 304 -1249
rect 310 -1245 311 -1243
rect 310 -1251 311 -1249
rect 317 -1245 318 -1243
rect 317 -1251 318 -1249
rect 324 -1245 325 -1243
rect 324 -1251 325 -1249
rect 331 -1245 332 -1243
rect 338 -1245 339 -1243
rect 338 -1251 339 -1249
rect 345 -1245 346 -1243
rect 345 -1251 346 -1249
rect 352 -1245 353 -1243
rect 352 -1251 353 -1249
rect 359 -1245 360 -1243
rect 359 -1251 360 -1249
rect 366 -1245 367 -1243
rect 366 -1251 367 -1249
rect 373 -1245 374 -1243
rect 373 -1251 374 -1249
rect 380 -1245 381 -1243
rect 380 -1251 381 -1249
rect 387 -1251 388 -1249
rect 394 -1245 395 -1243
rect 394 -1251 395 -1249
rect 401 -1245 402 -1243
rect 401 -1251 402 -1249
rect 408 -1245 409 -1243
rect 408 -1251 409 -1249
rect 415 -1245 416 -1243
rect 415 -1251 416 -1249
rect 422 -1245 423 -1243
rect 425 -1245 426 -1243
rect 422 -1251 423 -1249
rect 425 -1251 426 -1249
rect 429 -1245 430 -1243
rect 429 -1251 430 -1249
rect 436 -1245 437 -1243
rect 436 -1251 437 -1249
rect 443 -1245 444 -1243
rect 446 -1245 447 -1243
rect 443 -1251 444 -1249
rect 446 -1251 447 -1249
rect 450 -1245 451 -1243
rect 453 -1245 454 -1243
rect 450 -1251 451 -1249
rect 453 -1251 454 -1249
rect 457 -1245 458 -1243
rect 457 -1251 458 -1249
rect 464 -1245 465 -1243
rect 464 -1251 465 -1249
rect 471 -1245 472 -1243
rect 474 -1245 475 -1243
rect 474 -1251 475 -1249
rect 478 -1245 479 -1243
rect 478 -1251 479 -1249
rect 485 -1245 486 -1243
rect 485 -1251 486 -1249
rect 492 -1245 493 -1243
rect 492 -1251 493 -1249
rect 499 -1245 500 -1243
rect 499 -1251 500 -1249
rect 506 -1245 507 -1243
rect 506 -1251 507 -1249
rect 516 -1245 517 -1243
rect 513 -1251 514 -1249
rect 516 -1251 517 -1249
rect 520 -1245 521 -1243
rect 520 -1251 521 -1249
rect 527 -1245 528 -1243
rect 527 -1251 528 -1249
rect 534 -1245 535 -1243
rect 534 -1251 535 -1249
rect 541 -1245 542 -1243
rect 541 -1251 542 -1249
rect 548 -1245 549 -1243
rect 548 -1251 549 -1249
rect 555 -1245 556 -1243
rect 555 -1251 556 -1249
rect 562 -1245 563 -1243
rect 562 -1251 563 -1249
rect 565 -1251 566 -1249
rect 569 -1245 570 -1243
rect 569 -1251 570 -1249
rect 576 -1245 577 -1243
rect 576 -1251 577 -1249
rect 583 -1245 584 -1243
rect 586 -1245 587 -1243
rect 583 -1251 584 -1249
rect 586 -1251 587 -1249
rect 590 -1245 591 -1243
rect 590 -1251 591 -1249
rect 597 -1245 598 -1243
rect 597 -1251 598 -1249
rect 604 -1245 605 -1243
rect 604 -1251 605 -1249
rect 611 -1245 612 -1243
rect 611 -1251 612 -1249
rect 618 -1245 619 -1243
rect 618 -1251 619 -1249
rect 625 -1245 626 -1243
rect 625 -1251 626 -1249
rect 632 -1245 633 -1243
rect 632 -1251 633 -1249
rect 639 -1245 640 -1243
rect 639 -1251 640 -1249
rect 646 -1245 647 -1243
rect 646 -1251 647 -1249
rect 653 -1245 654 -1243
rect 653 -1251 654 -1249
rect 660 -1245 661 -1243
rect 660 -1251 661 -1249
rect 667 -1245 668 -1243
rect 670 -1245 671 -1243
rect 667 -1251 668 -1249
rect 670 -1251 671 -1249
rect 674 -1245 675 -1243
rect 674 -1251 675 -1249
rect 681 -1245 682 -1243
rect 681 -1251 682 -1249
rect 688 -1245 689 -1243
rect 688 -1251 689 -1249
rect 695 -1245 696 -1243
rect 695 -1251 696 -1249
rect 702 -1245 703 -1243
rect 702 -1251 703 -1249
rect 709 -1245 710 -1243
rect 709 -1251 710 -1249
rect 716 -1245 717 -1243
rect 716 -1251 717 -1249
rect 723 -1245 724 -1243
rect 723 -1251 724 -1249
rect 730 -1245 731 -1243
rect 730 -1251 731 -1249
rect 737 -1245 738 -1243
rect 737 -1251 738 -1249
rect 744 -1245 745 -1243
rect 747 -1245 748 -1243
rect 744 -1251 745 -1249
rect 751 -1245 752 -1243
rect 751 -1251 752 -1249
rect 758 -1245 759 -1243
rect 758 -1251 759 -1249
rect 765 -1245 766 -1243
rect 765 -1251 766 -1249
rect 772 -1245 773 -1243
rect 775 -1245 776 -1243
rect 772 -1251 773 -1249
rect 775 -1251 776 -1249
rect 779 -1245 780 -1243
rect 782 -1245 783 -1243
rect 779 -1251 780 -1249
rect 786 -1245 787 -1243
rect 786 -1251 787 -1249
rect 793 -1245 794 -1243
rect 793 -1251 794 -1249
rect 800 -1245 801 -1243
rect 800 -1251 801 -1249
rect 807 -1245 808 -1243
rect 810 -1245 811 -1243
rect 807 -1251 808 -1249
rect 810 -1251 811 -1249
rect 814 -1245 815 -1243
rect 814 -1251 815 -1249
rect 821 -1245 822 -1243
rect 821 -1251 822 -1249
rect 824 -1251 825 -1249
rect 828 -1245 829 -1243
rect 828 -1251 829 -1249
rect 835 -1245 836 -1243
rect 835 -1251 836 -1249
rect 842 -1245 843 -1243
rect 842 -1251 843 -1249
rect 849 -1245 850 -1243
rect 849 -1251 850 -1249
rect 856 -1245 857 -1243
rect 859 -1245 860 -1243
rect 856 -1251 857 -1249
rect 859 -1251 860 -1249
rect 863 -1245 864 -1243
rect 863 -1251 864 -1249
rect 870 -1245 871 -1243
rect 873 -1245 874 -1243
rect 873 -1251 874 -1249
rect 877 -1245 878 -1243
rect 880 -1245 881 -1243
rect 877 -1251 878 -1249
rect 884 -1245 885 -1243
rect 884 -1251 885 -1249
rect 891 -1245 892 -1243
rect 891 -1251 892 -1249
rect 898 -1245 899 -1243
rect 898 -1251 899 -1249
rect 905 -1245 906 -1243
rect 908 -1245 909 -1243
rect 905 -1251 906 -1249
rect 908 -1251 909 -1249
rect 912 -1245 913 -1243
rect 912 -1251 913 -1249
rect 919 -1245 920 -1243
rect 919 -1251 920 -1249
rect 926 -1245 927 -1243
rect 929 -1245 930 -1243
rect 926 -1251 927 -1249
rect 929 -1251 930 -1249
rect 933 -1245 934 -1243
rect 933 -1251 934 -1249
rect 940 -1245 941 -1243
rect 940 -1251 941 -1249
rect 947 -1245 948 -1243
rect 947 -1251 948 -1249
rect 954 -1245 955 -1243
rect 954 -1251 955 -1249
rect 964 -1245 965 -1243
rect 961 -1251 962 -1249
rect 964 -1251 965 -1249
rect 968 -1245 969 -1243
rect 968 -1251 969 -1249
rect 975 -1245 976 -1243
rect 975 -1251 976 -1249
rect 982 -1245 983 -1243
rect 982 -1251 983 -1249
rect 989 -1245 990 -1243
rect 989 -1251 990 -1249
rect 996 -1245 997 -1243
rect 996 -1251 997 -1249
rect 1003 -1245 1004 -1243
rect 1003 -1251 1004 -1249
rect 1010 -1245 1011 -1243
rect 1010 -1251 1011 -1249
rect 1017 -1245 1018 -1243
rect 1017 -1251 1018 -1249
rect 1020 -1251 1021 -1249
rect 1024 -1245 1025 -1243
rect 1024 -1251 1025 -1249
rect 1031 -1245 1032 -1243
rect 1031 -1251 1032 -1249
rect 1038 -1245 1039 -1243
rect 1038 -1251 1039 -1249
rect 1045 -1245 1046 -1243
rect 1048 -1245 1049 -1243
rect 1052 -1245 1053 -1243
rect 1052 -1251 1053 -1249
rect 1059 -1245 1060 -1243
rect 1059 -1251 1060 -1249
rect 1066 -1245 1067 -1243
rect 1066 -1251 1067 -1249
rect 1073 -1245 1074 -1243
rect 1073 -1251 1074 -1249
rect 1080 -1245 1081 -1243
rect 1080 -1251 1081 -1249
rect 1087 -1245 1088 -1243
rect 1087 -1251 1088 -1249
rect 1094 -1245 1095 -1243
rect 1094 -1251 1095 -1249
rect 1101 -1245 1102 -1243
rect 1101 -1251 1102 -1249
rect 1108 -1245 1109 -1243
rect 1108 -1251 1109 -1249
rect 1115 -1245 1116 -1243
rect 1115 -1251 1116 -1249
rect 1122 -1245 1123 -1243
rect 1122 -1251 1123 -1249
rect 1129 -1245 1130 -1243
rect 1132 -1245 1133 -1243
rect 1129 -1251 1130 -1249
rect 1132 -1251 1133 -1249
rect 1136 -1245 1137 -1243
rect 1136 -1251 1137 -1249
rect 1143 -1245 1144 -1243
rect 1143 -1251 1144 -1249
rect 1150 -1245 1151 -1243
rect 1150 -1251 1151 -1249
rect 1157 -1245 1158 -1243
rect 1160 -1245 1161 -1243
rect 1164 -1245 1165 -1243
rect 1164 -1251 1165 -1249
rect 1171 -1245 1172 -1243
rect 1171 -1251 1172 -1249
rect 1178 -1245 1179 -1243
rect 1181 -1245 1182 -1243
rect 1178 -1251 1179 -1249
rect 1181 -1251 1182 -1249
rect 1185 -1245 1186 -1243
rect 1185 -1251 1186 -1249
rect 1192 -1245 1193 -1243
rect 1192 -1251 1193 -1249
rect 1199 -1245 1200 -1243
rect 1199 -1251 1200 -1249
rect 1206 -1245 1207 -1243
rect 1206 -1251 1207 -1249
rect 1213 -1245 1214 -1243
rect 1213 -1251 1214 -1249
rect 1220 -1245 1221 -1243
rect 1220 -1251 1221 -1249
rect 1227 -1245 1228 -1243
rect 1227 -1251 1228 -1249
rect 1234 -1245 1235 -1243
rect 1234 -1251 1235 -1249
rect 1241 -1245 1242 -1243
rect 1241 -1251 1242 -1249
rect 1248 -1245 1249 -1243
rect 1248 -1251 1249 -1249
rect 1255 -1245 1256 -1243
rect 1255 -1251 1256 -1249
rect 1262 -1245 1263 -1243
rect 1262 -1251 1263 -1249
rect 1269 -1245 1270 -1243
rect 1269 -1251 1270 -1249
rect 1276 -1245 1277 -1243
rect 1276 -1251 1277 -1249
rect 1283 -1245 1284 -1243
rect 1283 -1251 1284 -1249
rect 1290 -1245 1291 -1243
rect 1290 -1251 1291 -1249
rect 1297 -1245 1298 -1243
rect 1297 -1251 1298 -1249
rect 1304 -1245 1305 -1243
rect 1304 -1251 1305 -1249
rect 1311 -1245 1312 -1243
rect 1311 -1251 1312 -1249
rect 1318 -1245 1319 -1243
rect 1318 -1251 1319 -1249
rect 1325 -1245 1326 -1243
rect 1325 -1251 1326 -1249
rect 1332 -1245 1333 -1243
rect 1332 -1251 1333 -1249
rect 1339 -1245 1340 -1243
rect 1339 -1251 1340 -1249
rect 1346 -1245 1347 -1243
rect 1346 -1251 1347 -1249
rect 1353 -1245 1354 -1243
rect 1353 -1251 1354 -1249
rect 1360 -1245 1361 -1243
rect 1360 -1251 1361 -1249
rect 1367 -1245 1368 -1243
rect 1367 -1251 1368 -1249
rect 1374 -1245 1375 -1243
rect 1374 -1251 1375 -1249
rect 1381 -1245 1382 -1243
rect 1381 -1251 1382 -1249
rect 1388 -1245 1389 -1243
rect 1388 -1251 1389 -1249
rect 1391 -1251 1392 -1249
rect 1395 -1245 1396 -1243
rect 1395 -1251 1396 -1249
rect 1402 -1245 1403 -1243
rect 1402 -1251 1403 -1249
rect 1409 -1245 1410 -1243
rect 1409 -1251 1410 -1249
rect 1416 -1245 1417 -1243
rect 1416 -1251 1417 -1249
rect 1423 -1245 1424 -1243
rect 1423 -1251 1424 -1249
rect 1430 -1245 1431 -1243
rect 1430 -1251 1431 -1249
rect 1437 -1245 1438 -1243
rect 1437 -1251 1438 -1249
rect 1444 -1245 1445 -1243
rect 1444 -1251 1445 -1249
rect 1451 -1245 1452 -1243
rect 1451 -1251 1452 -1249
rect 1458 -1245 1459 -1243
rect 1458 -1251 1459 -1249
rect 1465 -1245 1466 -1243
rect 1465 -1251 1466 -1249
rect 1472 -1245 1473 -1243
rect 1472 -1251 1473 -1249
rect 1479 -1245 1480 -1243
rect 1479 -1251 1480 -1249
rect 1486 -1245 1487 -1243
rect 1486 -1251 1487 -1249
rect 1493 -1245 1494 -1243
rect 1493 -1251 1494 -1249
rect 1500 -1245 1501 -1243
rect 1500 -1251 1501 -1249
rect 1507 -1245 1508 -1243
rect 1507 -1251 1508 -1249
rect 1514 -1245 1515 -1243
rect 1514 -1251 1515 -1249
rect 1521 -1245 1522 -1243
rect 1521 -1251 1522 -1249
rect 1528 -1245 1529 -1243
rect 1528 -1251 1529 -1249
rect 1535 -1245 1536 -1243
rect 1535 -1251 1536 -1249
rect 1542 -1245 1543 -1243
rect 1542 -1251 1543 -1249
rect 1549 -1245 1550 -1243
rect 1549 -1251 1550 -1249
rect 1556 -1245 1557 -1243
rect 1556 -1251 1557 -1249
rect 1563 -1245 1564 -1243
rect 1563 -1251 1564 -1249
rect 1570 -1245 1571 -1243
rect 1570 -1251 1571 -1249
rect 1577 -1245 1578 -1243
rect 1577 -1251 1578 -1249
rect 1584 -1245 1585 -1243
rect 1584 -1251 1585 -1249
rect 1591 -1245 1592 -1243
rect 1591 -1251 1592 -1249
rect 1598 -1245 1599 -1243
rect 1598 -1251 1599 -1249
rect 1605 -1245 1606 -1243
rect 1605 -1251 1606 -1249
rect 1612 -1245 1613 -1243
rect 1612 -1251 1613 -1249
rect 1619 -1245 1620 -1243
rect 1619 -1251 1620 -1249
rect 1626 -1245 1627 -1243
rect 1626 -1251 1627 -1249
rect 1633 -1245 1634 -1243
rect 1633 -1251 1634 -1249
rect 1640 -1245 1641 -1243
rect 1640 -1251 1641 -1249
rect 1647 -1245 1648 -1243
rect 1647 -1251 1648 -1249
rect 1654 -1245 1655 -1243
rect 1654 -1251 1655 -1249
rect 1661 -1245 1662 -1243
rect 1661 -1251 1662 -1249
rect 1668 -1245 1669 -1243
rect 1668 -1251 1669 -1249
rect 1675 -1245 1676 -1243
rect 1675 -1251 1676 -1249
rect 1682 -1245 1683 -1243
rect 1682 -1251 1683 -1249
rect 1689 -1245 1690 -1243
rect 1689 -1251 1690 -1249
rect 1696 -1245 1697 -1243
rect 1696 -1251 1697 -1249
rect 1703 -1245 1704 -1243
rect 1703 -1251 1704 -1249
rect 1710 -1245 1711 -1243
rect 1710 -1251 1711 -1249
rect 1717 -1245 1718 -1243
rect 1717 -1251 1718 -1249
rect 1724 -1245 1725 -1243
rect 1724 -1251 1725 -1249
rect 1731 -1245 1732 -1243
rect 1731 -1251 1732 -1249
rect 1738 -1245 1739 -1243
rect 1738 -1251 1739 -1249
rect 1745 -1245 1746 -1243
rect 1745 -1251 1746 -1249
rect 1752 -1245 1753 -1243
rect 1752 -1251 1753 -1249
rect 1759 -1245 1760 -1243
rect 1759 -1251 1760 -1249
rect 1766 -1245 1767 -1243
rect 1766 -1251 1767 -1249
rect 1773 -1245 1774 -1243
rect 1773 -1251 1774 -1249
rect 1780 -1245 1781 -1243
rect 1780 -1251 1781 -1249
rect 1787 -1245 1788 -1243
rect 1787 -1251 1788 -1249
rect 1794 -1245 1795 -1243
rect 1794 -1251 1795 -1249
rect 1801 -1245 1802 -1243
rect 1801 -1251 1802 -1249
rect 1808 -1245 1809 -1243
rect 1808 -1251 1809 -1249
rect 1815 -1245 1816 -1243
rect 1815 -1251 1816 -1249
rect 1822 -1245 1823 -1243
rect 1822 -1251 1823 -1249
rect 1829 -1245 1830 -1243
rect 1829 -1251 1830 -1249
rect 1836 -1245 1837 -1243
rect 1836 -1251 1837 -1249
rect 1843 -1245 1844 -1243
rect 1843 -1251 1844 -1249
rect 1850 -1245 1851 -1243
rect 1850 -1251 1851 -1249
rect 1857 -1245 1858 -1243
rect 1857 -1251 1858 -1249
rect 1864 -1245 1865 -1243
rect 1864 -1251 1865 -1249
rect 1871 -1245 1872 -1243
rect 1871 -1251 1872 -1249
rect 1878 -1245 1879 -1243
rect 1878 -1251 1879 -1249
rect 1885 -1245 1886 -1243
rect 1885 -1251 1886 -1249
rect 1892 -1245 1893 -1243
rect 1892 -1251 1893 -1249
rect 1899 -1245 1900 -1243
rect 1899 -1251 1900 -1249
rect 1906 -1245 1907 -1243
rect 1906 -1251 1907 -1249
rect 1913 -1245 1914 -1243
rect 1913 -1251 1914 -1249
rect 1920 -1245 1921 -1243
rect 1920 -1251 1921 -1249
rect 1927 -1245 1928 -1243
rect 1927 -1251 1928 -1249
rect 1955 -1245 1956 -1243
rect 1955 -1251 1956 -1249
rect 1962 -1245 1963 -1243
rect 1962 -1251 1963 -1249
rect 1969 -1245 1970 -1243
rect 1969 -1251 1970 -1249
rect 1976 -1245 1977 -1243
rect 1976 -1251 1977 -1249
rect 1990 -1245 1991 -1243
rect 1990 -1251 1991 -1249
rect 9 -1388 10 -1386
rect 9 -1394 10 -1392
rect 16 -1388 17 -1386
rect 16 -1394 17 -1392
rect 23 -1388 24 -1386
rect 23 -1394 24 -1392
rect 30 -1388 31 -1386
rect 30 -1394 31 -1392
rect 37 -1388 38 -1386
rect 37 -1394 38 -1392
rect 44 -1388 45 -1386
rect 44 -1394 45 -1392
rect 51 -1388 52 -1386
rect 54 -1388 55 -1386
rect 51 -1394 52 -1392
rect 58 -1388 59 -1386
rect 58 -1394 59 -1392
rect 61 -1394 62 -1392
rect 65 -1388 66 -1386
rect 65 -1394 66 -1392
rect 72 -1388 73 -1386
rect 75 -1388 76 -1386
rect 75 -1394 76 -1392
rect 79 -1388 80 -1386
rect 79 -1394 80 -1392
rect 86 -1388 87 -1386
rect 86 -1394 87 -1392
rect 93 -1388 94 -1386
rect 93 -1394 94 -1392
rect 100 -1388 101 -1386
rect 100 -1394 101 -1392
rect 107 -1388 108 -1386
rect 110 -1388 111 -1386
rect 110 -1394 111 -1392
rect 114 -1388 115 -1386
rect 114 -1394 115 -1392
rect 121 -1388 122 -1386
rect 121 -1394 122 -1392
rect 128 -1388 129 -1386
rect 128 -1394 129 -1392
rect 131 -1394 132 -1392
rect 135 -1388 136 -1386
rect 135 -1394 136 -1392
rect 142 -1388 143 -1386
rect 145 -1388 146 -1386
rect 145 -1394 146 -1392
rect 152 -1388 153 -1386
rect 149 -1394 150 -1392
rect 152 -1394 153 -1392
rect 156 -1388 157 -1386
rect 156 -1394 157 -1392
rect 163 -1388 164 -1386
rect 163 -1394 164 -1392
rect 166 -1394 167 -1392
rect 170 -1388 171 -1386
rect 170 -1394 171 -1392
rect 177 -1388 178 -1386
rect 177 -1394 178 -1392
rect 184 -1388 185 -1386
rect 184 -1394 185 -1392
rect 191 -1388 192 -1386
rect 191 -1394 192 -1392
rect 198 -1388 199 -1386
rect 198 -1394 199 -1392
rect 205 -1388 206 -1386
rect 208 -1388 209 -1386
rect 208 -1394 209 -1392
rect 212 -1388 213 -1386
rect 212 -1394 213 -1392
rect 219 -1388 220 -1386
rect 219 -1394 220 -1392
rect 226 -1388 227 -1386
rect 226 -1394 227 -1392
rect 233 -1388 234 -1386
rect 233 -1394 234 -1392
rect 240 -1388 241 -1386
rect 240 -1394 241 -1392
rect 247 -1388 248 -1386
rect 247 -1394 248 -1392
rect 254 -1388 255 -1386
rect 254 -1394 255 -1392
rect 261 -1388 262 -1386
rect 261 -1394 262 -1392
rect 268 -1388 269 -1386
rect 268 -1394 269 -1392
rect 275 -1388 276 -1386
rect 275 -1394 276 -1392
rect 282 -1388 283 -1386
rect 282 -1394 283 -1392
rect 289 -1388 290 -1386
rect 289 -1394 290 -1392
rect 296 -1388 297 -1386
rect 296 -1394 297 -1392
rect 303 -1388 304 -1386
rect 303 -1394 304 -1392
rect 310 -1388 311 -1386
rect 310 -1394 311 -1392
rect 317 -1388 318 -1386
rect 317 -1394 318 -1392
rect 324 -1388 325 -1386
rect 324 -1394 325 -1392
rect 331 -1394 332 -1392
rect 338 -1388 339 -1386
rect 338 -1394 339 -1392
rect 345 -1388 346 -1386
rect 345 -1394 346 -1392
rect 352 -1388 353 -1386
rect 352 -1394 353 -1392
rect 359 -1388 360 -1386
rect 359 -1394 360 -1392
rect 366 -1388 367 -1386
rect 366 -1394 367 -1392
rect 373 -1388 374 -1386
rect 373 -1394 374 -1392
rect 380 -1388 381 -1386
rect 380 -1394 381 -1392
rect 387 -1388 388 -1386
rect 387 -1394 388 -1392
rect 394 -1388 395 -1386
rect 394 -1394 395 -1392
rect 401 -1388 402 -1386
rect 401 -1394 402 -1392
rect 408 -1388 409 -1386
rect 408 -1394 409 -1392
rect 415 -1388 416 -1386
rect 415 -1394 416 -1392
rect 422 -1388 423 -1386
rect 422 -1394 423 -1392
rect 429 -1388 430 -1386
rect 432 -1388 433 -1386
rect 429 -1394 430 -1392
rect 432 -1394 433 -1392
rect 436 -1388 437 -1386
rect 436 -1394 437 -1392
rect 443 -1388 444 -1386
rect 443 -1394 444 -1392
rect 450 -1388 451 -1386
rect 450 -1394 451 -1392
rect 457 -1388 458 -1386
rect 457 -1394 458 -1392
rect 464 -1388 465 -1386
rect 464 -1394 465 -1392
rect 471 -1388 472 -1386
rect 471 -1394 472 -1392
rect 478 -1388 479 -1386
rect 478 -1394 479 -1392
rect 485 -1388 486 -1386
rect 485 -1394 486 -1392
rect 492 -1388 493 -1386
rect 492 -1394 493 -1392
rect 499 -1388 500 -1386
rect 499 -1394 500 -1392
rect 506 -1388 507 -1386
rect 506 -1394 507 -1392
rect 513 -1388 514 -1386
rect 513 -1394 514 -1392
rect 520 -1388 521 -1386
rect 520 -1394 521 -1392
rect 527 -1388 528 -1386
rect 530 -1388 531 -1386
rect 527 -1394 528 -1392
rect 530 -1394 531 -1392
rect 534 -1388 535 -1386
rect 534 -1394 535 -1392
rect 541 -1388 542 -1386
rect 541 -1394 542 -1392
rect 548 -1388 549 -1386
rect 548 -1394 549 -1392
rect 555 -1388 556 -1386
rect 555 -1394 556 -1392
rect 562 -1388 563 -1386
rect 562 -1394 563 -1392
rect 569 -1388 570 -1386
rect 569 -1394 570 -1392
rect 579 -1388 580 -1386
rect 576 -1394 577 -1392
rect 579 -1394 580 -1392
rect 583 -1388 584 -1386
rect 583 -1394 584 -1392
rect 590 -1388 591 -1386
rect 590 -1394 591 -1392
rect 597 -1388 598 -1386
rect 597 -1394 598 -1392
rect 604 -1388 605 -1386
rect 604 -1394 605 -1392
rect 611 -1388 612 -1386
rect 611 -1394 612 -1392
rect 618 -1388 619 -1386
rect 618 -1394 619 -1392
rect 625 -1388 626 -1386
rect 628 -1388 629 -1386
rect 625 -1394 626 -1392
rect 628 -1394 629 -1392
rect 632 -1388 633 -1386
rect 632 -1394 633 -1392
rect 639 -1388 640 -1386
rect 639 -1394 640 -1392
rect 646 -1388 647 -1386
rect 646 -1394 647 -1392
rect 653 -1388 654 -1386
rect 656 -1388 657 -1386
rect 653 -1394 654 -1392
rect 656 -1394 657 -1392
rect 660 -1388 661 -1386
rect 660 -1394 661 -1392
rect 667 -1388 668 -1386
rect 670 -1388 671 -1386
rect 667 -1394 668 -1392
rect 674 -1388 675 -1386
rect 677 -1388 678 -1386
rect 677 -1394 678 -1392
rect 681 -1388 682 -1386
rect 681 -1394 682 -1392
rect 688 -1388 689 -1386
rect 688 -1394 689 -1392
rect 695 -1388 696 -1386
rect 695 -1394 696 -1392
rect 702 -1388 703 -1386
rect 702 -1394 703 -1392
rect 709 -1388 710 -1386
rect 712 -1388 713 -1386
rect 709 -1394 710 -1392
rect 712 -1394 713 -1392
rect 716 -1388 717 -1386
rect 716 -1394 717 -1392
rect 723 -1388 724 -1386
rect 723 -1394 724 -1392
rect 730 -1388 731 -1386
rect 730 -1394 731 -1392
rect 737 -1388 738 -1386
rect 737 -1394 738 -1392
rect 744 -1388 745 -1386
rect 744 -1394 745 -1392
rect 751 -1388 752 -1386
rect 751 -1394 752 -1392
rect 758 -1388 759 -1386
rect 758 -1394 759 -1392
rect 765 -1388 766 -1386
rect 765 -1394 766 -1392
rect 772 -1388 773 -1386
rect 772 -1394 773 -1392
rect 779 -1388 780 -1386
rect 779 -1394 780 -1392
rect 786 -1388 787 -1386
rect 786 -1394 787 -1392
rect 793 -1388 794 -1386
rect 793 -1394 794 -1392
rect 800 -1388 801 -1386
rect 800 -1394 801 -1392
rect 807 -1388 808 -1386
rect 807 -1394 808 -1392
rect 814 -1388 815 -1386
rect 814 -1394 815 -1392
rect 821 -1388 822 -1386
rect 821 -1394 822 -1392
rect 828 -1388 829 -1386
rect 828 -1394 829 -1392
rect 835 -1388 836 -1386
rect 838 -1388 839 -1386
rect 835 -1394 836 -1392
rect 842 -1388 843 -1386
rect 842 -1394 843 -1392
rect 849 -1388 850 -1386
rect 849 -1394 850 -1392
rect 856 -1388 857 -1386
rect 859 -1388 860 -1386
rect 856 -1394 857 -1392
rect 859 -1394 860 -1392
rect 863 -1388 864 -1386
rect 863 -1394 864 -1392
rect 870 -1388 871 -1386
rect 870 -1394 871 -1392
rect 877 -1388 878 -1386
rect 877 -1394 878 -1392
rect 884 -1388 885 -1386
rect 884 -1394 885 -1392
rect 891 -1388 892 -1386
rect 891 -1394 892 -1392
rect 898 -1388 899 -1386
rect 898 -1394 899 -1392
rect 905 -1388 906 -1386
rect 905 -1394 906 -1392
rect 912 -1388 913 -1386
rect 912 -1394 913 -1392
rect 919 -1388 920 -1386
rect 922 -1388 923 -1386
rect 919 -1394 920 -1392
rect 922 -1394 923 -1392
rect 929 -1388 930 -1386
rect 926 -1394 927 -1392
rect 929 -1394 930 -1392
rect 933 -1388 934 -1386
rect 933 -1394 934 -1392
rect 943 -1388 944 -1386
rect 940 -1394 941 -1392
rect 943 -1394 944 -1392
rect 947 -1388 948 -1386
rect 947 -1394 948 -1392
rect 954 -1388 955 -1386
rect 954 -1394 955 -1392
rect 961 -1388 962 -1386
rect 961 -1394 962 -1392
rect 968 -1388 969 -1386
rect 968 -1394 969 -1392
rect 975 -1388 976 -1386
rect 975 -1394 976 -1392
rect 982 -1388 983 -1386
rect 982 -1394 983 -1392
rect 989 -1388 990 -1386
rect 989 -1394 990 -1392
rect 996 -1388 997 -1386
rect 999 -1388 1000 -1386
rect 996 -1394 997 -1392
rect 999 -1394 1000 -1392
rect 1003 -1388 1004 -1386
rect 1003 -1394 1004 -1392
rect 1010 -1388 1011 -1386
rect 1010 -1394 1011 -1392
rect 1017 -1388 1018 -1386
rect 1017 -1394 1018 -1392
rect 1024 -1388 1025 -1386
rect 1024 -1394 1025 -1392
rect 1031 -1388 1032 -1386
rect 1031 -1394 1032 -1392
rect 1034 -1394 1035 -1392
rect 1038 -1388 1039 -1386
rect 1038 -1394 1039 -1392
rect 1045 -1388 1046 -1386
rect 1052 -1388 1053 -1386
rect 1055 -1388 1056 -1386
rect 1052 -1394 1053 -1392
rect 1055 -1394 1056 -1392
rect 1059 -1388 1060 -1386
rect 1059 -1394 1060 -1392
rect 1066 -1388 1067 -1386
rect 1069 -1388 1070 -1386
rect 1066 -1394 1067 -1392
rect 1069 -1394 1070 -1392
rect 1073 -1388 1074 -1386
rect 1076 -1388 1077 -1386
rect 1076 -1394 1077 -1392
rect 1080 -1388 1081 -1386
rect 1080 -1394 1081 -1392
rect 1087 -1388 1088 -1386
rect 1087 -1394 1088 -1392
rect 1094 -1388 1095 -1386
rect 1094 -1394 1095 -1392
rect 1101 -1388 1102 -1386
rect 1101 -1394 1102 -1392
rect 1108 -1388 1109 -1386
rect 1111 -1388 1112 -1386
rect 1108 -1394 1109 -1392
rect 1111 -1394 1112 -1392
rect 1115 -1388 1116 -1386
rect 1115 -1394 1116 -1392
rect 1122 -1388 1123 -1386
rect 1122 -1394 1123 -1392
rect 1129 -1388 1130 -1386
rect 1129 -1394 1130 -1392
rect 1136 -1388 1137 -1386
rect 1136 -1394 1137 -1392
rect 1143 -1388 1144 -1386
rect 1143 -1394 1144 -1392
rect 1150 -1388 1151 -1386
rect 1150 -1394 1151 -1392
rect 1157 -1388 1158 -1386
rect 1157 -1394 1158 -1392
rect 1164 -1388 1165 -1386
rect 1164 -1394 1165 -1392
rect 1171 -1388 1172 -1386
rect 1171 -1394 1172 -1392
rect 1178 -1388 1179 -1386
rect 1178 -1394 1179 -1392
rect 1185 -1388 1186 -1386
rect 1185 -1394 1186 -1392
rect 1192 -1388 1193 -1386
rect 1192 -1394 1193 -1392
rect 1199 -1388 1200 -1386
rect 1199 -1394 1200 -1392
rect 1206 -1388 1207 -1386
rect 1206 -1394 1207 -1392
rect 1213 -1388 1214 -1386
rect 1213 -1394 1214 -1392
rect 1220 -1388 1221 -1386
rect 1220 -1394 1221 -1392
rect 1227 -1388 1228 -1386
rect 1227 -1394 1228 -1392
rect 1234 -1388 1235 -1386
rect 1234 -1394 1235 -1392
rect 1241 -1388 1242 -1386
rect 1244 -1388 1245 -1386
rect 1241 -1394 1242 -1392
rect 1244 -1394 1245 -1392
rect 1248 -1388 1249 -1386
rect 1248 -1394 1249 -1392
rect 1255 -1388 1256 -1386
rect 1255 -1394 1256 -1392
rect 1262 -1388 1263 -1386
rect 1262 -1394 1263 -1392
rect 1269 -1388 1270 -1386
rect 1269 -1394 1270 -1392
rect 1276 -1388 1277 -1386
rect 1276 -1394 1277 -1392
rect 1283 -1388 1284 -1386
rect 1283 -1394 1284 -1392
rect 1286 -1394 1287 -1392
rect 1290 -1388 1291 -1386
rect 1290 -1394 1291 -1392
rect 1297 -1388 1298 -1386
rect 1297 -1394 1298 -1392
rect 1304 -1388 1305 -1386
rect 1304 -1394 1305 -1392
rect 1311 -1388 1312 -1386
rect 1311 -1394 1312 -1392
rect 1318 -1388 1319 -1386
rect 1318 -1394 1319 -1392
rect 1325 -1388 1326 -1386
rect 1325 -1394 1326 -1392
rect 1332 -1388 1333 -1386
rect 1332 -1394 1333 -1392
rect 1339 -1388 1340 -1386
rect 1339 -1394 1340 -1392
rect 1346 -1388 1347 -1386
rect 1346 -1394 1347 -1392
rect 1353 -1388 1354 -1386
rect 1353 -1394 1354 -1392
rect 1360 -1388 1361 -1386
rect 1360 -1394 1361 -1392
rect 1367 -1388 1368 -1386
rect 1367 -1394 1368 -1392
rect 1374 -1388 1375 -1386
rect 1374 -1394 1375 -1392
rect 1381 -1388 1382 -1386
rect 1381 -1394 1382 -1392
rect 1388 -1388 1389 -1386
rect 1391 -1388 1392 -1386
rect 1388 -1394 1389 -1392
rect 1395 -1388 1396 -1386
rect 1395 -1394 1396 -1392
rect 1402 -1388 1403 -1386
rect 1402 -1394 1403 -1392
rect 1409 -1388 1410 -1386
rect 1409 -1394 1410 -1392
rect 1416 -1388 1417 -1386
rect 1416 -1394 1417 -1392
rect 1423 -1388 1424 -1386
rect 1423 -1394 1424 -1392
rect 1430 -1388 1431 -1386
rect 1430 -1394 1431 -1392
rect 1437 -1388 1438 -1386
rect 1437 -1394 1438 -1392
rect 1444 -1388 1445 -1386
rect 1444 -1394 1445 -1392
rect 1451 -1388 1452 -1386
rect 1451 -1394 1452 -1392
rect 1458 -1388 1459 -1386
rect 1458 -1394 1459 -1392
rect 1465 -1388 1466 -1386
rect 1465 -1394 1466 -1392
rect 1472 -1388 1473 -1386
rect 1472 -1394 1473 -1392
rect 1479 -1388 1480 -1386
rect 1479 -1394 1480 -1392
rect 1486 -1388 1487 -1386
rect 1486 -1394 1487 -1392
rect 1493 -1388 1494 -1386
rect 1493 -1394 1494 -1392
rect 1500 -1388 1501 -1386
rect 1500 -1394 1501 -1392
rect 1507 -1388 1508 -1386
rect 1507 -1394 1508 -1392
rect 1514 -1388 1515 -1386
rect 1514 -1394 1515 -1392
rect 1521 -1388 1522 -1386
rect 1521 -1394 1522 -1392
rect 1528 -1388 1529 -1386
rect 1528 -1394 1529 -1392
rect 1535 -1388 1536 -1386
rect 1535 -1394 1536 -1392
rect 1542 -1388 1543 -1386
rect 1542 -1394 1543 -1392
rect 1549 -1388 1550 -1386
rect 1549 -1394 1550 -1392
rect 1556 -1388 1557 -1386
rect 1556 -1394 1557 -1392
rect 1563 -1388 1564 -1386
rect 1563 -1394 1564 -1392
rect 1570 -1388 1571 -1386
rect 1570 -1394 1571 -1392
rect 1577 -1388 1578 -1386
rect 1577 -1394 1578 -1392
rect 1584 -1388 1585 -1386
rect 1584 -1394 1585 -1392
rect 1591 -1388 1592 -1386
rect 1591 -1394 1592 -1392
rect 1598 -1388 1599 -1386
rect 1598 -1394 1599 -1392
rect 1605 -1388 1606 -1386
rect 1605 -1394 1606 -1392
rect 1612 -1388 1613 -1386
rect 1612 -1394 1613 -1392
rect 1619 -1388 1620 -1386
rect 1619 -1394 1620 -1392
rect 1626 -1388 1627 -1386
rect 1626 -1394 1627 -1392
rect 1633 -1388 1634 -1386
rect 1633 -1394 1634 -1392
rect 1640 -1388 1641 -1386
rect 1640 -1394 1641 -1392
rect 1647 -1388 1648 -1386
rect 1647 -1394 1648 -1392
rect 1654 -1388 1655 -1386
rect 1654 -1394 1655 -1392
rect 1661 -1388 1662 -1386
rect 1661 -1394 1662 -1392
rect 1668 -1388 1669 -1386
rect 1668 -1394 1669 -1392
rect 1675 -1388 1676 -1386
rect 1675 -1394 1676 -1392
rect 1682 -1388 1683 -1386
rect 1682 -1394 1683 -1392
rect 1689 -1388 1690 -1386
rect 1689 -1394 1690 -1392
rect 1696 -1388 1697 -1386
rect 1696 -1394 1697 -1392
rect 1703 -1388 1704 -1386
rect 1703 -1394 1704 -1392
rect 1710 -1388 1711 -1386
rect 1710 -1394 1711 -1392
rect 1717 -1388 1718 -1386
rect 1717 -1394 1718 -1392
rect 1724 -1388 1725 -1386
rect 1724 -1394 1725 -1392
rect 1731 -1388 1732 -1386
rect 1731 -1394 1732 -1392
rect 1738 -1388 1739 -1386
rect 1738 -1394 1739 -1392
rect 1745 -1388 1746 -1386
rect 1745 -1394 1746 -1392
rect 1752 -1388 1753 -1386
rect 1752 -1394 1753 -1392
rect 1759 -1388 1760 -1386
rect 1759 -1394 1760 -1392
rect 1766 -1388 1767 -1386
rect 1766 -1394 1767 -1392
rect 1773 -1388 1774 -1386
rect 1773 -1394 1774 -1392
rect 1780 -1388 1781 -1386
rect 1780 -1394 1781 -1392
rect 1787 -1388 1788 -1386
rect 1787 -1394 1788 -1392
rect 1794 -1388 1795 -1386
rect 1794 -1394 1795 -1392
rect 1801 -1388 1802 -1386
rect 1801 -1394 1802 -1392
rect 1808 -1388 1809 -1386
rect 1808 -1394 1809 -1392
rect 1815 -1388 1816 -1386
rect 1815 -1394 1816 -1392
rect 1822 -1388 1823 -1386
rect 1822 -1394 1823 -1392
rect 1829 -1388 1830 -1386
rect 1829 -1394 1830 -1392
rect 1836 -1388 1837 -1386
rect 1836 -1394 1837 -1392
rect 1843 -1388 1844 -1386
rect 1843 -1394 1844 -1392
rect 1850 -1388 1851 -1386
rect 1850 -1394 1851 -1392
rect 1857 -1388 1858 -1386
rect 1857 -1394 1858 -1392
rect 1864 -1388 1865 -1386
rect 1864 -1394 1865 -1392
rect 1871 -1388 1872 -1386
rect 1871 -1394 1872 -1392
rect 1878 -1388 1879 -1386
rect 1878 -1394 1879 -1392
rect 1885 -1388 1886 -1386
rect 1885 -1394 1886 -1392
rect 1892 -1388 1893 -1386
rect 1892 -1394 1893 -1392
rect 1899 -1388 1900 -1386
rect 1899 -1394 1900 -1392
rect 1906 -1388 1907 -1386
rect 1906 -1394 1907 -1392
rect 1913 -1388 1914 -1386
rect 1916 -1388 1917 -1386
rect 1913 -1394 1914 -1392
rect 1916 -1394 1917 -1392
rect 1920 -1388 1921 -1386
rect 1920 -1394 1921 -1392
rect 1927 -1388 1928 -1386
rect 1927 -1394 1928 -1392
rect 1934 -1388 1935 -1386
rect 1934 -1394 1935 -1392
rect 1941 -1388 1942 -1386
rect 1941 -1394 1942 -1392
rect 1948 -1388 1949 -1386
rect 1948 -1394 1949 -1392
rect 1969 -1388 1970 -1386
rect 1969 -1394 1970 -1392
rect 1976 -1388 1977 -1386
rect 1976 -1394 1977 -1392
rect 1983 -1388 1984 -1386
rect 1983 -1394 1984 -1392
rect 1986 -1394 1987 -1392
rect 1990 -1388 1991 -1386
rect 1990 -1394 1991 -1392
rect 1997 -1388 1998 -1386
rect 1997 -1394 1998 -1392
rect 2 -1519 3 -1517
rect 2 -1525 3 -1523
rect 9 -1519 10 -1517
rect 9 -1525 10 -1523
rect 16 -1519 17 -1517
rect 16 -1525 17 -1523
rect 23 -1519 24 -1517
rect 23 -1525 24 -1523
rect 30 -1519 31 -1517
rect 30 -1525 31 -1523
rect 37 -1519 38 -1517
rect 37 -1525 38 -1523
rect 44 -1519 45 -1517
rect 47 -1519 48 -1517
rect 44 -1525 45 -1523
rect 47 -1525 48 -1523
rect 51 -1519 52 -1517
rect 51 -1525 52 -1523
rect 58 -1519 59 -1517
rect 61 -1519 62 -1517
rect 58 -1525 59 -1523
rect 65 -1519 66 -1517
rect 65 -1525 66 -1523
rect 72 -1519 73 -1517
rect 72 -1525 73 -1523
rect 79 -1519 80 -1517
rect 82 -1519 83 -1517
rect 79 -1525 80 -1523
rect 82 -1525 83 -1523
rect 86 -1519 87 -1517
rect 86 -1525 87 -1523
rect 93 -1519 94 -1517
rect 93 -1525 94 -1523
rect 100 -1519 101 -1517
rect 100 -1525 101 -1523
rect 107 -1519 108 -1517
rect 107 -1525 108 -1523
rect 114 -1519 115 -1517
rect 114 -1525 115 -1523
rect 121 -1519 122 -1517
rect 121 -1525 122 -1523
rect 128 -1519 129 -1517
rect 128 -1525 129 -1523
rect 135 -1519 136 -1517
rect 135 -1525 136 -1523
rect 142 -1519 143 -1517
rect 145 -1519 146 -1517
rect 142 -1525 143 -1523
rect 145 -1525 146 -1523
rect 149 -1519 150 -1517
rect 149 -1525 150 -1523
rect 156 -1519 157 -1517
rect 156 -1525 157 -1523
rect 163 -1519 164 -1517
rect 163 -1525 164 -1523
rect 170 -1519 171 -1517
rect 170 -1525 171 -1523
rect 177 -1519 178 -1517
rect 177 -1525 178 -1523
rect 184 -1519 185 -1517
rect 184 -1525 185 -1523
rect 191 -1519 192 -1517
rect 194 -1519 195 -1517
rect 191 -1525 192 -1523
rect 194 -1525 195 -1523
rect 198 -1519 199 -1517
rect 198 -1525 199 -1523
rect 205 -1519 206 -1517
rect 205 -1525 206 -1523
rect 212 -1519 213 -1517
rect 215 -1519 216 -1517
rect 212 -1525 213 -1523
rect 219 -1519 220 -1517
rect 219 -1525 220 -1523
rect 226 -1519 227 -1517
rect 226 -1525 227 -1523
rect 233 -1519 234 -1517
rect 233 -1525 234 -1523
rect 240 -1519 241 -1517
rect 243 -1519 244 -1517
rect 240 -1525 241 -1523
rect 247 -1519 248 -1517
rect 247 -1525 248 -1523
rect 254 -1519 255 -1517
rect 254 -1525 255 -1523
rect 261 -1519 262 -1517
rect 261 -1525 262 -1523
rect 268 -1519 269 -1517
rect 268 -1525 269 -1523
rect 275 -1519 276 -1517
rect 275 -1525 276 -1523
rect 282 -1519 283 -1517
rect 282 -1525 283 -1523
rect 289 -1519 290 -1517
rect 289 -1525 290 -1523
rect 296 -1519 297 -1517
rect 296 -1525 297 -1523
rect 303 -1519 304 -1517
rect 303 -1525 304 -1523
rect 310 -1519 311 -1517
rect 310 -1525 311 -1523
rect 317 -1519 318 -1517
rect 317 -1525 318 -1523
rect 324 -1519 325 -1517
rect 324 -1525 325 -1523
rect 331 -1519 332 -1517
rect 331 -1525 332 -1523
rect 338 -1519 339 -1517
rect 338 -1525 339 -1523
rect 345 -1519 346 -1517
rect 345 -1525 346 -1523
rect 352 -1519 353 -1517
rect 352 -1525 353 -1523
rect 359 -1519 360 -1517
rect 359 -1525 360 -1523
rect 366 -1519 367 -1517
rect 366 -1525 367 -1523
rect 373 -1519 374 -1517
rect 373 -1525 374 -1523
rect 380 -1519 381 -1517
rect 380 -1525 381 -1523
rect 387 -1519 388 -1517
rect 387 -1525 388 -1523
rect 394 -1519 395 -1517
rect 394 -1525 395 -1523
rect 401 -1519 402 -1517
rect 401 -1525 402 -1523
rect 408 -1519 409 -1517
rect 408 -1525 409 -1523
rect 415 -1519 416 -1517
rect 415 -1525 416 -1523
rect 422 -1519 423 -1517
rect 422 -1525 423 -1523
rect 429 -1519 430 -1517
rect 429 -1525 430 -1523
rect 436 -1519 437 -1517
rect 436 -1525 437 -1523
rect 443 -1519 444 -1517
rect 443 -1525 444 -1523
rect 450 -1519 451 -1517
rect 450 -1525 451 -1523
rect 457 -1519 458 -1517
rect 457 -1525 458 -1523
rect 464 -1519 465 -1517
rect 464 -1525 465 -1523
rect 471 -1519 472 -1517
rect 471 -1525 472 -1523
rect 478 -1519 479 -1517
rect 478 -1525 479 -1523
rect 485 -1519 486 -1517
rect 485 -1525 486 -1523
rect 492 -1519 493 -1517
rect 492 -1525 493 -1523
rect 502 -1519 503 -1517
rect 499 -1525 500 -1523
rect 502 -1525 503 -1523
rect 506 -1519 507 -1517
rect 506 -1525 507 -1523
rect 513 -1519 514 -1517
rect 513 -1525 514 -1523
rect 520 -1519 521 -1517
rect 520 -1525 521 -1523
rect 527 -1519 528 -1517
rect 527 -1525 528 -1523
rect 534 -1519 535 -1517
rect 534 -1525 535 -1523
rect 541 -1519 542 -1517
rect 541 -1525 542 -1523
rect 548 -1519 549 -1517
rect 548 -1525 549 -1523
rect 555 -1519 556 -1517
rect 555 -1525 556 -1523
rect 562 -1519 563 -1517
rect 562 -1525 563 -1523
rect 569 -1519 570 -1517
rect 569 -1525 570 -1523
rect 576 -1519 577 -1517
rect 576 -1525 577 -1523
rect 583 -1519 584 -1517
rect 583 -1525 584 -1523
rect 590 -1519 591 -1517
rect 590 -1525 591 -1523
rect 593 -1525 594 -1523
rect 597 -1519 598 -1517
rect 597 -1525 598 -1523
rect 604 -1519 605 -1517
rect 604 -1525 605 -1523
rect 611 -1519 612 -1517
rect 611 -1525 612 -1523
rect 618 -1519 619 -1517
rect 618 -1525 619 -1523
rect 625 -1519 626 -1517
rect 628 -1519 629 -1517
rect 625 -1525 626 -1523
rect 628 -1525 629 -1523
rect 632 -1519 633 -1517
rect 632 -1525 633 -1523
rect 639 -1519 640 -1517
rect 639 -1525 640 -1523
rect 646 -1519 647 -1517
rect 646 -1525 647 -1523
rect 653 -1519 654 -1517
rect 653 -1525 654 -1523
rect 660 -1519 661 -1517
rect 663 -1519 664 -1517
rect 660 -1525 661 -1523
rect 663 -1525 664 -1523
rect 667 -1519 668 -1517
rect 670 -1519 671 -1517
rect 667 -1525 668 -1523
rect 670 -1525 671 -1523
rect 674 -1519 675 -1517
rect 674 -1525 675 -1523
rect 681 -1519 682 -1517
rect 681 -1525 682 -1523
rect 688 -1519 689 -1517
rect 688 -1525 689 -1523
rect 695 -1519 696 -1517
rect 695 -1525 696 -1523
rect 702 -1519 703 -1517
rect 702 -1525 703 -1523
rect 709 -1519 710 -1517
rect 712 -1519 713 -1517
rect 709 -1525 710 -1523
rect 712 -1525 713 -1523
rect 716 -1519 717 -1517
rect 716 -1525 717 -1523
rect 723 -1519 724 -1517
rect 723 -1525 724 -1523
rect 730 -1519 731 -1517
rect 730 -1525 731 -1523
rect 737 -1519 738 -1517
rect 737 -1525 738 -1523
rect 744 -1519 745 -1517
rect 744 -1525 745 -1523
rect 751 -1519 752 -1517
rect 754 -1519 755 -1517
rect 751 -1525 752 -1523
rect 754 -1525 755 -1523
rect 758 -1519 759 -1517
rect 758 -1525 759 -1523
rect 765 -1519 766 -1517
rect 765 -1525 766 -1523
rect 772 -1519 773 -1517
rect 772 -1525 773 -1523
rect 779 -1519 780 -1517
rect 779 -1525 780 -1523
rect 786 -1519 787 -1517
rect 786 -1525 787 -1523
rect 793 -1519 794 -1517
rect 793 -1525 794 -1523
rect 800 -1519 801 -1517
rect 800 -1525 801 -1523
rect 807 -1519 808 -1517
rect 807 -1525 808 -1523
rect 814 -1519 815 -1517
rect 814 -1525 815 -1523
rect 821 -1519 822 -1517
rect 821 -1525 822 -1523
rect 828 -1519 829 -1517
rect 828 -1525 829 -1523
rect 835 -1519 836 -1517
rect 835 -1525 836 -1523
rect 842 -1519 843 -1517
rect 842 -1525 843 -1523
rect 849 -1519 850 -1517
rect 849 -1525 850 -1523
rect 856 -1519 857 -1517
rect 856 -1525 857 -1523
rect 863 -1519 864 -1517
rect 863 -1525 864 -1523
rect 870 -1519 871 -1517
rect 870 -1525 871 -1523
rect 877 -1519 878 -1517
rect 877 -1525 878 -1523
rect 884 -1519 885 -1517
rect 884 -1525 885 -1523
rect 891 -1519 892 -1517
rect 891 -1525 892 -1523
rect 898 -1519 899 -1517
rect 898 -1525 899 -1523
rect 905 -1519 906 -1517
rect 905 -1525 906 -1523
rect 912 -1519 913 -1517
rect 912 -1525 913 -1523
rect 922 -1519 923 -1517
rect 919 -1525 920 -1523
rect 922 -1525 923 -1523
rect 926 -1519 927 -1517
rect 926 -1525 927 -1523
rect 933 -1519 934 -1517
rect 933 -1525 934 -1523
rect 940 -1519 941 -1517
rect 940 -1525 941 -1523
rect 947 -1519 948 -1517
rect 950 -1519 951 -1517
rect 950 -1525 951 -1523
rect 954 -1519 955 -1517
rect 957 -1519 958 -1517
rect 954 -1525 955 -1523
rect 957 -1525 958 -1523
rect 961 -1519 962 -1517
rect 968 -1519 969 -1517
rect 968 -1525 969 -1523
rect 975 -1519 976 -1517
rect 975 -1525 976 -1523
rect 982 -1519 983 -1517
rect 985 -1519 986 -1517
rect 982 -1525 983 -1523
rect 985 -1525 986 -1523
rect 989 -1519 990 -1517
rect 989 -1525 990 -1523
rect 996 -1519 997 -1517
rect 996 -1525 997 -1523
rect 1003 -1519 1004 -1517
rect 1006 -1519 1007 -1517
rect 1003 -1525 1004 -1523
rect 1006 -1525 1007 -1523
rect 1010 -1519 1011 -1517
rect 1010 -1525 1011 -1523
rect 1017 -1519 1018 -1517
rect 1017 -1525 1018 -1523
rect 1024 -1519 1025 -1517
rect 1024 -1525 1025 -1523
rect 1031 -1519 1032 -1517
rect 1031 -1525 1032 -1523
rect 1038 -1519 1039 -1517
rect 1038 -1525 1039 -1523
rect 1045 -1525 1046 -1523
rect 1052 -1519 1053 -1517
rect 1052 -1525 1053 -1523
rect 1059 -1519 1060 -1517
rect 1059 -1525 1060 -1523
rect 1069 -1519 1070 -1517
rect 1066 -1525 1067 -1523
rect 1069 -1525 1070 -1523
rect 1073 -1519 1074 -1517
rect 1073 -1525 1074 -1523
rect 1080 -1519 1081 -1517
rect 1080 -1525 1081 -1523
rect 1087 -1519 1088 -1517
rect 1087 -1525 1088 -1523
rect 1094 -1519 1095 -1517
rect 1094 -1525 1095 -1523
rect 1101 -1519 1102 -1517
rect 1104 -1519 1105 -1517
rect 1101 -1525 1102 -1523
rect 1104 -1525 1105 -1523
rect 1108 -1519 1109 -1517
rect 1111 -1519 1112 -1517
rect 1108 -1525 1109 -1523
rect 1111 -1525 1112 -1523
rect 1115 -1519 1116 -1517
rect 1118 -1519 1119 -1517
rect 1115 -1525 1116 -1523
rect 1118 -1525 1119 -1523
rect 1122 -1519 1123 -1517
rect 1122 -1525 1123 -1523
rect 1129 -1519 1130 -1517
rect 1132 -1519 1133 -1517
rect 1129 -1525 1130 -1523
rect 1132 -1525 1133 -1523
rect 1136 -1519 1137 -1517
rect 1136 -1525 1137 -1523
rect 1143 -1519 1144 -1517
rect 1143 -1525 1144 -1523
rect 1150 -1519 1151 -1517
rect 1150 -1525 1151 -1523
rect 1157 -1519 1158 -1517
rect 1160 -1519 1161 -1517
rect 1157 -1525 1158 -1523
rect 1160 -1525 1161 -1523
rect 1164 -1519 1165 -1517
rect 1164 -1525 1165 -1523
rect 1171 -1519 1172 -1517
rect 1171 -1525 1172 -1523
rect 1178 -1519 1179 -1517
rect 1178 -1525 1179 -1523
rect 1185 -1519 1186 -1517
rect 1185 -1525 1186 -1523
rect 1192 -1519 1193 -1517
rect 1192 -1525 1193 -1523
rect 1195 -1525 1196 -1523
rect 1199 -1519 1200 -1517
rect 1199 -1525 1200 -1523
rect 1206 -1519 1207 -1517
rect 1206 -1525 1207 -1523
rect 1213 -1519 1214 -1517
rect 1213 -1525 1214 -1523
rect 1220 -1519 1221 -1517
rect 1220 -1525 1221 -1523
rect 1227 -1519 1228 -1517
rect 1227 -1525 1228 -1523
rect 1234 -1519 1235 -1517
rect 1234 -1525 1235 -1523
rect 1241 -1519 1242 -1517
rect 1241 -1525 1242 -1523
rect 1248 -1519 1249 -1517
rect 1248 -1525 1249 -1523
rect 1255 -1519 1256 -1517
rect 1255 -1525 1256 -1523
rect 1262 -1519 1263 -1517
rect 1265 -1519 1266 -1517
rect 1262 -1525 1263 -1523
rect 1265 -1525 1266 -1523
rect 1269 -1519 1270 -1517
rect 1269 -1525 1270 -1523
rect 1276 -1519 1277 -1517
rect 1276 -1525 1277 -1523
rect 1283 -1519 1284 -1517
rect 1283 -1525 1284 -1523
rect 1290 -1519 1291 -1517
rect 1290 -1525 1291 -1523
rect 1297 -1519 1298 -1517
rect 1297 -1525 1298 -1523
rect 1304 -1519 1305 -1517
rect 1307 -1519 1308 -1517
rect 1307 -1525 1308 -1523
rect 1311 -1519 1312 -1517
rect 1311 -1525 1312 -1523
rect 1318 -1519 1319 -1517
rect 1318 -1525 1319 -1523
rect 1325 -1519 1326 -1517
rect 1325 -1525 1326 -1523
rect 1332 -1519 1333 -1517
rect 1335 -1519 1336 -1517
rect 1332 -1525 1333 -1523
rect 1335 -1525 1336 -1523
rect 1339 -1519 1340 -1517
rect 1339 -1525 1340 -1523
rect 1346 -1519 1347 -1517
rect 1346 -1525 1347 -1523
rect 1353 -1519 1354 -1517
rect 1353 -1525 1354 -1523
rect 1360 -1519 1361 -1517
rect 1360 -1525 1361 -1523
rect 1367 -1519 1368 -1517
rect 1367 -1525 1368 -1523
rect 1374 -1519 1375 -1517
rect 1374 -1525 1375 -1523
rect 1381 -1519 1382 -1517
rect 1381 -1525 1382 -1523
rect 1388 -1519 1389 -1517
rect 1388 -1525 1389 -1523
rect 1395 -1519 1396 -1517
rect 1395 -1525 1396 -1523
rect 1402 -1519 1403 -1517
rect 1402 -1525 1403 -1523
rect 1409 -1519 1410 -1517
rect 1409 -1525 1410 -1523
rect 1416 -1519 1417 -1517
rect 1416 -1525 1417 -1523
rect 1423 -1519 1424 -1517
rect 1423 -1525 1424 -1523
rect 1430 -1519 1431 -1517
rect 1430 -1525 1431 -1523
rect 1437 -1519 1438 -1517
rect 1437 -1525 1438 -1523
rect 1444 -1519 1445 -1517
rect 1444 -1525 1445 -1523
rect 1451 -1519 1452 -1517
rect 1451 -1525 1452 -1523
rect 1458 -1519 1459 -1517
rect 1458 -1525 1459 -1523
rect 1465 -1519 1466 -1517
rect 1465 -1525 1466 -1523
rect 1472 -1519 1473 -1517
rect 1472 -1525 1473 -1523
rect 1479 -1519 1480 -1517
rect 1479 -1525 1480 -1523
rect 1486 -1519 1487 -1517
rect 1486 -1525 1487 -1523
rect 1493 -1519 1494 -1517
rect 1493 -1525 1494 -1523
rect 1500 -1519 1501 -1517
rect 1500 -1525 1501 -1523
rect 1507 -1519 1508 -1517
rect 1507 -1525 1508 -1523
rect 1514 -1519 1515 -1517
rect 1514 -1525 1515 -1523
rect 1521 -1519 1522 -1517
rect 1521 -1525 1522 -1523
rect 1528 -1519 1529 -1517
rect 1528 -1525 1529 -1523
rect 1535 -1519 1536 -1517
rect 1535 -1525 1536 -1523
rect 1542 -1519 1543 -1517
rect 1542 -1525 1543 -1523
rect 1549 -1519 1550 -1517
rect 1549 -1525 1550 -1523
rect 1556 -1519 1557 -1517
rect 1556 -1525 1557 -1523
rect 1563 -1519 1564 -1517
rect 1563 -1525 1564 -1523
rect 1570 -1519 1571 -1517
rect 1570 -1525 1571 -1523
rect 1577 -1519 1578 -1517
rect 1577 -1525 1578 -1523
rect 1584 -1519 1585 -1517
rect 1584 -1525 1585 -1523
rect 1591 -1519 1592 -1517
rect 1591 -1525 1592 -1523
rect 1598 -1519 1599 -1517
rect 1598 -1525 1599 -1523
rect 1605 -1519 1606 -1517
rect 1605 -1525 1606 -1523
rect 1612 -1519 1613 -1517
rect 1612 -1525 1613 -1523
rect 1619 -1519 1620 -1517
rect 1619 -1525 1620 -1523
rect 1626 -1519 1627 -1517
rect 1626 -1525 1627 -1523
rect 1633 -1519 1634 -1517
rect 1633 -1525 1634 -1523
rect 1640 -1519 1641 -1517
rect 1640 -1525 1641 -1523
rect 1647 -1519 1648 -1517
rect 1647 -1525 1648 -1523
rect 1654 -1519 1655 -1517
rect 1654 -1525 1655 -1523
rect 1661 -1519 1662 -1517
rect 1661 -1525 1662 -1523
rect 1668 -1519 1669 -1517
rect 1668 -1525 1669 -1523
rect 1675 -1519 1676 -1517
rect 1675 -1525 1676 -1523
rect 1682 -1519 1683 -1517
rect 1682 -1525 1683 -1523
rect 1689 -1519 1690 -1517
rect 1689 -1525 1690 -1523
rect 1696 -1519 1697 -1517
rect 1696 -1525 1697 -1523
rect 1703 -1519 1704 -1517
rect 1703 -1525 1704 -1523
rect 1710 -1519 1711 -1517
rect 1710 -1525 1711 -1523
rect 1717 -1519 1718 -1517
rect 1717 -1525 1718 -1523
rect 1724 -1519 1725 -1517
rect 1724 -1525 1725 -1523
rect 1731 -1519 1732 -1517
rect 1731 -1525 1732 -1523
rect 1738 -1519 1739 -1517
rect 1738 -1525 1739 -1523
rect 1745 -1519 1746 -1517
rect 1745 -1525 1746 -1523
rect 1752 -1519 1753 -1517
rect 1752 -1525 1753 -1523
rect 1759 -1519 1760 -1517
rect 1759 -1525 1760 -1523
rect 1766 -1519 1767 -1517
rect 1766 -1525 1767 -1523
rect 1773 -1519 1774 -1517
rect 1773 -1525 1774 -1523
rect 1780 -1519 1781 -1517
rect 1780 -1525 1781 -1523
rect 1787 -1519 1788 -1517
rect 1787 -1525 1788 -1523
rect 1794 -1519 1795 -1517
rect 1794 -1525 1795 -1523
rect 1801 -1519 1802 -1517
rect 1801 -1525 1802 -1523
rect 1808 -1519 1809 -1517
rect 1808 -1525 1809 -1523
rect 1815 -1519 1816 -1517
rect 1815 -1525 1816 -1523
rect 1822 -1519 1823 -1517
rect 1822 -1525 1823 -1523
rect 1829 -1519 1830 -1517
rect 1829 -1525 1830 -1523
rect 1836 -1519 1837 -1517
rect 1836 -1525 1837 -1523
rect 1843 -1519 1844 -1517
rect 1843 -1525 1844 -1523
rect 1850 -1519 1851 -1517
rect 1850 -1525 1851 -1523
rect 1857 -1519 1858 -1517
rect 1857 -1525 1858 -1523
rect 1864 -1519 1865 -1517
rect 1864 -1525 1865 -1523
rect 1871 -1519 1872 -1517
rect 1871 -1525 1872 -1523
rect 1878 -1519 1879 -1517
rect 1878 -1525 1879 -1523
rect 1885 -1519 1886 -1517
rect 1885 -1525 1886 -1523
rect 1892 -1519 1893 -1517
rect 1892 -1525 1893 -1523
rect 1899 -1519 1900 -1517
rect 1899 -1525 1900 -1523
rect 1906 -1519 1907 -1517
rect 1906 -1525 1907 -1523
rect 1913 -1519 1914 -1517
rect 1913 -1525 1914 -1523
rect 1920 -1519 1921 -1517
rect 1920 -1525 1921 -1523
rect 1927 -1519 1928 -1517
rect 1927 -1525 1928 -1523
rect 1934 -1519 1935 -1517
rect 1934 -1525 1935 -1523
rect 1941 -1519 1942 -1517
rect 1941 -1525 1942 -1523
rect 1948 -1519 1949 -1517
rect 1948 -1525 1949 -1523
rect 1955 -1519 1956 -1517
rect 1955 -1525 1956 -1523
rect 1962 -1519 1963 -1517
rect 1962 -1525 1963 -1523
rect 1969 -1519 1970 -1517
rect 1969 -1525 1970 -1523
rect 1972 -1525 1973 -1523
rect 1976 -1525 1977 -1523
rect 1979 -1525 1980 -1523
rect 1983 -1519 1984 -1517
rect 1986 -1519 1987 -1517
rect 1983 -1525 1984 -1523
rect 1990 -1519 1991 -1517
rect 1990 -1525 1991 -1523
rect 1997 -1519 1998 -1517
rect 2000 -1525 2001 -1523
rect 2007 -1519 2008 -1517
rect 2004 -1525 2005 -1523
rect 2007 -1525 2008 -1523
rect 2011 -1519 2012 -1517
rect 2011 -1525 2012 -1523
rect 2018 -1519 2019 -1517
rect 2018 -1525 2019 -1523
rect 2025 -1519 2026 -1517
rect 2025 -1525 2026 -1523
rect 2 -1646 3 -1644
rect 2 -1652 3 -1650
rect 9 -1646 10 -1644
rect 9 -1652 10 -1650
rect 16 -1646 17 -1644
rect 16 -1652 17 -1650
rect 23 -1646 24 -1644
rect 23 -1652 24 -1650
rect 30 -1646 31 -1644
rect 30 -1652 31 -1650
rect 37 -1646 38 -1644
rect 37 -1652 38 -1650
rect 44 -1646 45 -1644
rect 44 -1652 45 -1650
rect 51 -1646 52 -1644
rect 51 -1652 52 -1650
rect 58 -1646 59 -1644
rect 58 -1652 59 -1650
rect 65 -1646 66 -1644
rect 68 -1646 69 -1644
rect 65 -1652 66 -1650
rect 72 -1646 73 -1644
rect 72 -1652 73 -1650
rect 79 -1646 80 -1644
rect 82 -1646 83 -1644
rect 82 -1652 83 -1650
rect 86 -1646 87 -1644
rect 89 -1646 90 -1644
rect 89 -1652 90 -1650
rect 93 -1646 94 -1644
rect 93 -1652 94 -1650
rect 100 -1646 101 -1644
rect 100 -1652 101 -1650
rect 107 -1646 108 -1644
rect 107 -1652 108 -1650
rect 114 -1646 115 -1644
rect 117 -1646 118 -1644
rect 114 -1652 115 -1650
rect 117 -1652 118 -1650
rect 121 -1646 122 -1644
rect 121 -1652 122 -1650
rect 128 -1646 129 -1644
rect 128 -1652 129 -1650
rect 135 -1646 136 -1644
rect 135 -1652 136 -1650
rect 142 -1646 143 -1644
rect 145 -1646 146 -1644
rect 142 -1652 143 -1650
rect 149 -1646 150 -1644
rect 149 -1652 150 -1650
rect 156 -1646 157 -1644
rect 156 -1652 157 -1650
rect 163 -1646 164 -1644
rect 163 -1652 164 -1650
rect 170 -1646 171 -1644
rect 173 -1646 174 -1644
rect 170 -1652 171 -1650
rect 177 -1646 178 -1644
rect 180 -1646 181 -1644
rect 180 -1652 181 -1650
rect 184 -1646 185 -1644
rect 184 -1652 185 -1650
rect 191 -1646 192 -1644
rect 191 -1652 192 -1650
rect 198 -1646 199 -1644
rect 198 -1652 199 -1650
rect 205 -1646 206 -1644
rect 205 -1652 206 -1650
rect 212 -1646 213 -1644
rect 212 -1652 213 -1650
rect 219 -1646 220 -1644
rect 219 -1652 220 -1650
rect 226 -1646 227 -1644
rect 226 -1652 227 -1650
rect 233 -1646 234 -1644
rect 233 -1652 234 -1650
rect 240 -1646 241 -1644
rect 240 -1652 241 -1650
rect 247 -1646 248 -1644
rect 247 -1652 248 -1650
rect 254 -1646 255 -1644
rect 254 -1652 255 -1650
rect 261 -1646 262 -1644
rect 261 -1652 262 -1650
rect 268 -1646 269 -1644
rect 268 -1652 269 -1650
rect 275 -1646 276 -1644
rect 275 -1652 276 -1650
rect 282 -1646 283 -1644
rect 282 -1652 283 -1650
rect 289 -1646 290 -1644
rect 289 -1652 290 -1650
rect 296 -1646 297 -1644
rect 296 -1652 297 -1650
rect 303 -1646 304 -1644
rect 303 -1652 304 -1650
rect 310 -1646 311 -1644
rect 310 -1652 311 -1650
rect 317 -1646 318 -1644
rect 317 -1652 318 -1650
rect 324 -1646 325 -1644
rect 324 -1652 325 -1650
rect 331 -1646 332 -1644
rect 331 -1652 332 -1650
rect 338 -1646 339 -1644
rect 338 -1652 339 -1650
rect 345 -1646 346 -1644
rect 345 -1652 346 -1650
rect 352 -1646 353 -1644
rect 352 -1652 353 -1650
rect 359 -1646 360 -1644
rect 359 -1652 360 -1650
rect 366 -1646 367 -1644
rect 366 -1652 367 -1650
rect 373 -1646 374 -1644
rect 373 -1652 374 -1650
rect 380 -1646 381 -1644
rect 380 -1652 381 -1650
rect 387 -1646 388 -1644
rect 387 -1652 388 -1650
rect 394 -1646 395 -1644
rect 397 -1646 398 -1644
rect 394 -1652 395 -1650
rect 397 -1652 398 -1650
rect 401 -1646 402 -1644
rect 401 -1652 402 -1650
rect 408 -1646 409 -1644
rect 408 -1652 409 -1650
rect 418 -1646 419 -1644
rect 418 -1652 419 -1650
rect 422 -1646 423 -1644
rect 422 -1652 423 -1650
rect 429 -1646 430 -1644
rect 429 -1652 430 -1650
rect 436 -1646 437 -1644
rect 436 -1652 437 -1650
rect 443 -1646 444 -1644
rect 443 -1652 444 -1650
rect 450 -1646 451 -1644
rect 450 -1652 451 -1650
rect 457 -1646 458 -1644
rect 457 -1652 458 -1650
rect 464 -1646 465 -1644
rect 464 -1652 465 -1650
rect 471 -1646 472 -1644
rect 471 -1652 472 -1650
rect 478 -1646 479 -1644
rect 478 -1652 479 -1650
rect 485 -1646 486 -1644
rect 485 -1652 486 -1650
rect 492 -1646 493 -1644
rect 492 -1652 493 -1650
rect 499 -1646 500 -1644
rect 499 -1652 500 -1650
rect 506 -1646 507 -1644
rect 506 -1652 507 -1650
rect 513 -1646 514 -1644
rect 513 -1652 514 -1650
rect 520 -1646 521 -1644
rect 520 -1652 521 -1650
rect 527 -1646 528 -1644
rect 527 -1652 528 -1650
rect 534 -1646 535 -1644
rect 534 -1652 535 -1650
rect 541 -1646 542 -1644
rect 544 -1646 545 -1644
rect 541 -1652 542 -1650
rect 544 -1652 545 -1650
rect 548 -1646 549 -1644
rect 548 -1652 549 -1650
rect 555 -1646 556 -1644
rect 555 -1652 556 -1650
rect 562 -1646 563 -1644
rect 562 -1652 563 -1650
rect 569 -1646 570 -1644
rect 569 -1652 570 -1650
rect 576 -1646 577 -1644
rect 576 -1652 577 -1650
rect 583 -1646 584 -1644
rect 583 -1652 584 -1650
rect 590 -1646 591 -1644
rect 590 -1652 591 -1650
rect 597 -1646 598 -1644
rect 597 -1652 598 -1650
rect 604 -1646 605 -1644
rect 604 -1652 605 -1650
rect 611 -1646 612 -1644
rect 611 -1652 612 -1650
rect 618 -1646 619 -1644
rect 618 -1652 619 -1650
rect 625 -1646 626 -1644
rect 625 -1652 626 -1650
rect 632 -1646 633 -1644
rect 632 -1652 633 -1650
rect 639 -1646 640 -1644
rect 639 -1652 640 -1650
rect 646 -1646 647 -1644
rect 646 -1652 647 -1650
rect 653 -1646 654 -1644
rect 653 -1652 654 -1650
rect 660 -1646 661 -1644
rect 663 -1646 664 -1644
rect 660 -1652 661 -1650
rect 663 -1652 664 -1650
rect 667 -1646 668 -1644
rect 670 -1646 671 -1644
rect 667 -1652 668 -1650
rect 670 -1652 671 -1650
rect 674 -1646 675 -1644
rect 674 -1652 675 -1650
rect 681 -1646 682 -1644
rect 681 -1652 682 -1650
rect 688 -1646 689 -1644
rect 688 -1652 689 -1650
rect 698 -1646 699 -1644
rect 695 -1652 696 -1650
rect 702 -1646 703 -1644
rect 702 -1652 703 -1650
rect 712 -1646 713 -1644
rect 709 -1652 710 -1650
rect 712 -1652 713 -1650
rect 716 -1646 717 -1644
rect 716 -1652 717 -1650
rect 723 -1646 724 -1644
rect 723 -1652 724 -1650
rect 730 -1646 731 -1644
rect 730 -1652 731 -1650
rect 737 -1646 738 -1644
rect 740 -1646 741 -1644
rect 737 -1652 738 -1650
rect 740 -1652 741 -1650
rect 744 -1646 745 -1644
rect 744 -1652 745 -1650
rect 751 -1646 752 -1644
rect 751 -1652 752 -1650
rect 758 -1646 759 -1644
rect 758 -1652 759 -1650
rect 768 -1646 769 -1644
rect 768 -1652 769 -1650
rect 772 -1646 773 -1644
rect 772 -1652 773 -1650
rect 779 -1646 780 -1644
rect 779 -1652 780 -1650
rect 786 -1646 787 -1644
rect 786 -1652 787 -1650
rect 793 -1646 794 -1644
rect 793 -1652 794 -1650
rect 800 -1646 801 -1644
rect 800 -1652 801 -1650
rect 807 -1646 808 -1644
rect 807 -1652 808 -1650
rect 814 -1646 815 -1644
rect 817 -1646 818 -1644
rect 814 -1652 815 -1650
rect 821 -1646 822 -1644
rect 821 -1652 822 -1650
rect 828 -1646 829 -1644
rect 831 -1646 832 -1644
rect 828 -1652 829 -1650
rect 831 -1652 832 -1650
rect 835 -1646 836 -1644
rect 835 -1652 836 -1650
rect 842 -1646 843 -1644
rect 842 -1652 843 -1650
rect 849 -1646 850 -1644
rect 849 -1652 850 -1650
rect 856 -1646 857 -1644
rect 856 -1652 857 -1650
rect 863 -1646 864 -1644
rect 863 -1652 864 -1650
rect 870 -1646 871 -1644
rect 870 -1652 871 -1650
rect 877 -1646 878 -1644
rect 877 -1652 878 -1650
rect 884 -1646 885 -1644
rect 884 -1652 885 -1650
rect 891 -1646 892 -1644
rect 891 -1652 892 -1650
rect 898 -1646 899 -1644
rect 898 -1652 899 -1650
rect 905 -1646 906 -1644
rect 905 -1652 906 -1650
rect 912 -1646 913 -1644
rect 912 -1652 913 -1650
rect 919 -1646 920 -1644
rect 922 -1646 923 -1644
rect 919 -1652 920 -1650
rect 922 -1652 923 -1650
rect 926 -1646 927 -1644
rect 926 -1652 927 -1650
rect 933 -1646 934 -1644
rect 933 -1652 934 -1650
rect 940 -1646 941 -1644
rect 940 -1652 941 -1650
rect 943 -1652 944 -1650
rect 947 -1646 948 -1644
rect 947 -1652 948 -1650
rect 954 -1646 955 -1644
rect 954 -1652 955 -1650
rect 961 -1646 962 -1644
rect 961 -1652 962 -1650
rect 968 -1646 969 -1644
rect 971 -1646 972 -1644
rect 968 -1652 969 -1650
rect 971 -1652 972 -1650
rect 975 -1646 976 -1644
rect 975 -1652 976 -1650
rect 982 -1646 983 -1644
rect 982 -1652 983 -1650
rect 989 -1646 990 -1644
rect 989 -1652 990 -1650
rect 996 -1646 997 -1644
rect 996 -1652 997 -1650
rect 1003 -1646 1004 -1644
rect 1003 -1652 1004 -1650
rect 1010 -1646 1011 -1644
rect 1010 -1652 1011 -1650
rect 1017 -1646 1018 -1644
rect 1017 -1652 1018 -1650
rect 1024 -1646 1025 -1644
rect 1024 -1652 1025 -1650
rect 1031 -1646 1032 -1644
rect 1031 -1652 1032 -1650
rect 1038 -1646 1039 -1644
rect 1038 -1652 1039 -1650
rect 1041 -1652 1042 -1650
rect 1045 -1646 1046 -1644
rect 1045 -1652 1046 -1650
rect 1052 -1646 1053 -1644
rect 1055 -1646 1056 -1644
rect 1052 -1652 1053 -1650
rect 1055 -1652 1056 -1650
rect 1059 -1646 1060 -1644
rect 1059 -1652 1060 -1650
rect 1066 -1646 1067 -1644
rect 1066 -1652 1067 -1650
rect 1073 -1646 1074 -1644
rect 1073 -1652 1074 -1650
rect 1080 -1646 1081 -1644
rect 1080 -1652 1081 -1650
rect 1087 -1646 1088 -1644
rect 1090 -1646 1091 -1644
rect 1087 -1652 1088 -1650
rect 1094 -1646 1095 -1644
rect 1094 -1652 1095 -1650
rect 1101 -1646 1102 -1644
rect 1101 -1652 1102 -1650
rect 1108 -1646 1109 -1644
rect 1108 -1652 1109 -1650
rect 1115 -1646 1116 -1644
rect 1115 -1652 1116 -1650
rect 1122 -1646 1123 -1644
rect 1122 -1652 1123 -1650
rect 1129 -1646 1130 -1644
rect 1132 -1646 1133 -1644
rect 1129 -1652 1130 -1650
rect 1132 -1652 1133 -1650
rect 1136 -1646 1137 -1644
rect 1136 -1652 1137 -1650
rect 1143 -1646 1144 -1644
rect 1143 -1652 1144 -1650
rect 1150 -1646 1151 -1644
rect 1150 -1652 1151 -1650
rect 1157 -1646 1158 -1644
rect 1157 -1652 1158 -1650
rect 1164 -1646 1165 -1644
rect 1164 -1652 1165 -1650
rect 1171 -1646 1172 -1644
rect 1171 -1652 1172 -1650
rect 1178 -1646 1179 -1644
rect 1178 -1652 1179 -1650
rect 1185 -1646 1186 -1644
rect 1185 -1652 1186 -1650
rect 1192 -1646 1193 -1644
rect 1192 -1652 1193 -1650
rect 1199 -1646 1200 -1644
rect 1199 -1652 1200 -1650
rect 1206 -1646 1207 -1644
rect 1209 -1646 1210 -1644
rect 1206 -1652 1207 -1650
rect 1209 -1652 1210 -1650
rect 1213 -1646 1214 -1644
rect 1213 -1652 1214 -1650
rect 1220 -1646 1221 -1644
rect 1220 -1652 1221 -1650
rect 1227 -1646 1228 -1644
rect 1227 -1652 1228 -1650
rect 1234 -1646 1235 -1644
rect 1234 -1652 1235 -1650
rect 1241 -1646 1242 -1644
rect 1244 -1646 1245 -1644
rect 1241 -1652 1242 -1650
rect 1244 -1652 1245 -1650
rect 1248 -1646 1249 -1644
rect 1248 -1652 1249 -1650
rect 1255 -1646 1256 -1644
rect 1255 -1652 1256 -1650
rect 1262 -1646 1263 -1644
rect 1262 -1652 1263 -1650
rect 1269 -1646 1270 -1644
rect 1269 -1652 1270 -1650
rect 1276 -1646 1277 -1644
rect 1276 -1652 1277 -1650
rect 1283 -1646 1284 -1644
rect 1286 -1646 1287 -1644
rect 1283 -1652 1284 -1650
rect 1286 -1652 1287 -1650
rect 1290 -1646 1291 -1644
rect 1290 -1652 1291 -1650
rect 1297 -1646 1298 -1644
rect 1297 -1652 1298 -1650
rect 1304 -1646 1305 -1644
rect 1307 -1646 1308 -1644
rect 1304 -1652 1305 -1650
rect 1307 -1652 1308 -1650
rect 1311 -1646 1312 -1644
rect 1311 -1652 1312 -1650
rect 1318 -1646 1319 -1644
rect 1318 -1652 1319 -1650
rect 1325 -1646 1326 -1644
rect 1325 -1652 1326 -1650
rect 1332 -1646 1333 -1644
rect 1335 -1646 1336 -1644
rect 1332 -1652 1333 -1650
rect 1335 -1652 1336 -1650
rect 1339 -1646 1340 -1644
rect 1339 -1652 1340 -1650
rect 1346 -1646 1347 -1644
rect 1346 -1652 1347 -1650
rect 1353 -1646 1354 -1644
rect 1356 -1646 1357 -1644
rect 1353 -1652 1354 -1650
rect 1356 -1652 1357 -1650
rect 1360 -1646 1361 -1644
rect 1360 -1652 1361 -1650
rect 1367 -1646 1368 -1644
rect 1367 -1652 1368 -1650
rect 1374 -1646 1375 -1644
rect 1374 -1652 1375 -1650
rect 1381 -1646 1382 -1644
rect 1381 -1652 1382 -1650
rect 1388 -1646 1389 -1644
rect 1388 -1652 1389 -1650
rect 1395 -1646 1396 -1644
rect 1395 -1652 1396 -1650
rect 1402 -1646 1403 -1644
rect 1402 -1652 1403 -1650
rect 1409 -1646 1410 -1644
rect 1409 -1652 1410 -1650
rect 1416 -1646 1417 -1644
rect 1416 -1652 1417 -1650
rect 1423 -1646 1424 -1644
rect 1423 -1652 1424 -1650
rect 1430 -1646 1431 -1644
rect 1430 -1652 1431 -1650
rect 1437 -1646 1438 -1644
rect 1437 -1652 1438 -1650
rect 1444 -1646 1445 -1644
rect 1444 -1652 1445 -1650
rect 1451 -1646 1452 -1644
rect 1451 -1652 1452 -1650
rect 1458 -1646 1459 -1644
rect 1458 -1652 1459 -1650
rect 1465 -1646 1466 -1644
rect 1465 -1652 1466 -1650
rect 1468 -1652 1469 -1650
rect 1472 -1646 1473 -1644
rect 1472 -1652 1473 -1650
rect 1479 -1646 1480 -1644
rect 1479 -1652 1480 -1650
rect 1486 -1646 1487 -1644
rect 1486 -1652 1487 -1650
rect 1493 -1646 1494 -1644
rect 1493 -1652 1494 -1650
rect 1500 -1646 1501 -1644
rect 1503 -1646 1504 -1644
rect 1500 -1652 1501 -1650
rect 1507 -1646 1508 -1644
rect 1507 -1652 1508 -1650
rect 1514 -1646 1515 -1644
rect 1514 -1652 1515 -1650
rect 1521 -1646 1522 -1644
rect 1521 -1652 1522 -1650
rect 1528 -1646 1529 -1644
rect 1528 -1652 1529 -1650
rect 1535 -1646 1536 -1644
rect 1535 -1652 1536 -1650
rect 1542 -1646 1543 -1644
rect 1542 -1652 1543 -1650
rect 1549 -1646 1550 -1644
rect 1549 -1652 1550 -1650
rect 1556 -1646 1557 -1644
rect 1556 -1652 1557 -1650
rect 1563 -1646 1564 -1644
rect 1563 -1652 1564 -1650
rect 1570 -1646 1571 -1644
rect 1570 -1652 1571 -1650
rect 1577 -1646 1578 -1644
rect 1577 -1652 1578 -1650
rect 1584 -1646 1585 -1644
rect 1584 -1652 1585 -1650
rect 1591 -1646 1592 -1644
rect 1591 -1652 1592 -1650
rect 1598 -1646 1599 -1644
rect 1598 -1652 1599 -1650
rect 1605 -1646 1606 -1644
rect 1605 -1652 1606 -1650
rect 1612 -1646 1613 -1644
rect 1612 -1652 1613 -1650
rect 1619 -1646 1620 -1644
rect 1619 -1652 1620 -1650
rect 1626 -1646 1627 -1644
rect 1626 -1652 1627 -1650
rect 1633 -1646 1634 -1644
rect 1633 -1652 1634 -1650
rect 1640 -1646 1641 -1644
rect 1640 -1652 1641 -1650
rect 1647 -1646 1648 -1644
rect 1647 -1652 1648 -1650
rect 1654 -1646 1655 -1644
rect 1654 -1652 1655 -1650
rect 1661 -1646 1662 -1644
rect 1661 -1652 1662 -1650
rect 1668 -1646 1669 -1644
rect 1668 -1652 1669 -1650
rect 1675 -1646 1676 -1644
rect 1675 -1652 1676 -1650
rect 1682 -1646 1683 -1644
rect 1682 -1652 1683 -1650
rect 1689 -1646 1690 -1644
rect 1689 -1652 1690 -1650
rect 1696 -1646 1697 -1644
rect 1696 -1652 1697 -1650
rect 1703 -1646 1704 -1644
rect 1703 -1652 1704 -1650
rect 1710 -1646 1711 -1644
rect 1710 -1652 1711 -1650
rect 1717 -1646 1718 -1644
rect 1717 -1652 1718 -1650
rect 1724 -1646 1725 -1644
rect 1724 -1652 1725 -1650
rect 1731 -1646 1732 -1644
rect 1731 -1652 1732 -1650
rect 1738 -1646 1739 -1644
rect 1738 -1652 1739 -1650
rect 1745 -1646 1746 -1644
rect 1745 -1652 1746 -1650
rect 1752 -1646 1753 -1644
rect 1752 -1652 1753 -1650
rect 1759 -1646 1760 -1644
rect 1759 -1652 1760 -1650
rect 1766 -1646 1767 -1644
rect 1766 -1652 1767 -1650
rect 1773 -1646 1774 -1644
rect 1773 -1652 1774 -1650
rect 1780 -1646 1781 -1644
rect 1780 -1652 1781 -1650
rect 1787 -1646 1788 -1644
rect 1787 -1652 1788 -1650
rect 1794 -1646 1795 -1644
rect 1794 -1652 1795 -1650
rect 1801 -1646 1802 -1644
rect 1801 -1652 1802 -1650
rect 1808 -1646 1809 -1644
rect 1808 -1652 1809 -1650
rect 1815 -1646 1816 -1644
rect 1815 -1652 1816 -1650
rect 1822 -1646 1823 -1644
rect 1822 -1652 1823 -1650
rect 1829 -1646 1830 -1644
rect 1829 -1652 1830 -1650
rect 1836 -1646 1837 -1644
rect 1836 -1652 1837 -1650
rect 1843 -1646 1844 -1644
rect 1843 -1652 1844 -1650
rect 1846 -1652 1847 -1650
rect 1850 -1646 1851 -1644
rect 1850 -1652 1851 -1650
rect 1857 -1646 1858 -1644
rect 1857 -1652 1858 -1650
rect 1864 -1646 1865 -1644
rect 1864 -1652 1865 -1650
rect 1871 -1646 1872 -1644
rect 1871 -1652 1872 -1650
rect 1878 -1646 1879 -1644
rect 1881 -1646 1882 -1644
rect 1878 -1652 1879 -1650
rect 1885 -1646 1886 -1644
rect 1885 -1652 1886 -1650
rect 1892 -1646 1893 -1644
rect 1892 -1652 1893 -1650
rect 1899 -1646 1900 -1644
rect 1899 -1652 1900 -1650
rect 1906 -1646 1907 -1644
rect 1906 -1652 1907 -1650
rect 1913 -1646 1914 -1644
rect 1913 -1652 1914 -1650
rect 1920 -1646 1921 -1644
rect 1920 -1652 1921 -1650
rect 1927 -1646 1928 -1644
rect 1927 -1652 1928 -1650
rect 1934 -1646 1935 -1644
rect 1934 -1652 1935 -1650
rect 1941 -1646 1942 -1644
rect 1941 -1652 1942 -1650
rect 1948 -1646 1949 -1644
rect 1948 -1652 1949 -1650
rect 1976 -1646 1977 -1644
rect 1976 -1652 1977 -1650
rect 2018 -1646 2019 -1644
rect 2018 -1652 2019 -1650
rect 9 -1775 10 -1773
rect 9 -1781 10 -1779
rect 16 -1775 17 -1773
rect 16 -1781 17 -1779
rect 23 -1775 24 -1773
rect 23 -1781 24 -1779
rect 30 -1775 31 -1773
rect 30 -1781 31 -1779
rect 37 -1775 38 -1773
rect 37 -1781 38 -1779
rect 44 -1775 45 -1773
rect 44 -1781 45 -1779
rect 51 -1775 52 -1773
rect 51 -1781 52 -1779
rect 58 -1775 59 -1773
rect 58 -1781 59 -1779
rect 68 -1775 69 -1773
rect 65 -1781 66 -1779
rect 68 -1781 69 -1779
rect 72 -1775 73 -1773
rect 72 -1781 73 -1779
rect 79 -1775 80 -1773
rect 79 -1781 80 -1779
rect 86 -1775 87 -1773
rect 86 -1781 87 -1779
rect 93 -1775 94 -1773
rect 93 -1781 94 -1779
rect 100 -1775 101 -1773
rect 100 -1781 101 -1779
rect 107 -1775 108 -1773
rect 107 -1781 108 -1779
rect 114 -1775 115 -1773
rect 114 -1781 115 -1779
rect 121 -1775 122 -1773
rect 121 -1781 122 -1779
rect 128 -1775 129 -1773
rect 131 -1775 132 -1773
rect 131 -1781 132 -1779
rect 135 -1775 136 -1773
rect 135 -1781 136 -1779
rect 142 -1775 143 -1773
rect 142 -1781 143 -1779
rect 149 -1775 150 -1773
rect 149 -1781 150 -1779
rect 156 -1775 157 -1773
rect 156 -1781 157 -1779
rect 163 -1775 164 -1773
rect 163 -1781 164 -1779
rect 170 -1775 171 -1773
rect 170 -1781 171 -1779
rect 177 -1775 178 -1773
rect 177 -1781 178 -1779
rect 184 -1775 185 -1773
rect 187 -1775 188 -1773
rect 184 -1781 185 -1779
rect 187 -1781 188 -1779
rect 191 -1775 192 -1773
rect 194 -1775 195 -1773
rect 191 -1781 192 -1779
rect 198 -1775 199 -1773
rect 201 -1775 202 -1773
rect 198 -1781 199 -1779
rect 205 -1775 206 -1773
rect 205 -1781 206 -1779
rect 212 -1775 213 -1773
rect 212 -1781 213 -1779
rect 219 -1775 220 -1773
rect 219 -1781 220 -1779
rect 226 -1775 227 -1773
rect 226 -1781 227 -1779
rect 233 -1775 234 -1773
rect 233 -1781 234 -1779
rect 240 -1775 241 -1773
rect 240 -1781 241 -1779
rect 247 -1775 248 -1773
rect 247 -1781 248 -1779
rect 254 -1775 255 -1773
rect 254 -1781 255 -1779
rect 261 -1775 262 -1773
rect 261 -1781 262 -1779
rect 268 -1775 269 -1773
rect 268 -1781 269 -1779
rect 275 -1775 276 -1773
rect 275 -1781 276 -1779
rect 282 -1775 283 -1773
rect 282 -1781 283 -1779
rect 289 -1775 290 -1773
rect 289 -1781 290 -1779
rect 296 -1775 297 -1773
rect 296 -1781 297 -1779
rect 303 -1775 304 -1773
rect 303 -1781 304 -1779
rect 310 -1775 311 -1773
rect 310 -1781 311 -1779
rect 317 -1775 318 -1773
rect 317 -1781 318 -1779
rect 324 -1775 325 -1773
rect 324 -1781 325 -1779
rect 331 -1775 332 -1773
rect 331 -1781 332 -1779
rect 338 -1775 339 -1773
rect 345 -1775 346 -1773
rect 345 -1781 346 -1779
rect 352 -1775 353 -1773
rect 352 -1781 353 -1779
rect 359 -1775 360 -1773
rect 359 -1781 360 -1779
rect 366 -1775 367 -1773
rect 366 -1781 367 -1779
rect 373 -1775 374 -1773
rect 373 -1781 374 -1779
rect 380 -1775 381 -1773
rect 380 -1781 381 -1779
rect 387 -1775 388 -1773
rect 387 -1781 388 -1779
rect 394 -1775 395 -1773
rect 397 -1775 398 -1773
rect 394 -1781 395 -1779
rect 397 -1781 398 -1779
rect 401 -1775 402 -1773
rect 401 -1781 402 -1779
rect 408 -1775 409 -1773
rect 408 -1781 409 -1779
rect 415 -1775 416 -1773
rect 418 -1775 419 -1773
rect 415 -1781 416 -1779
rect 418 -1781 419 -1779
rect 422 -1775 423 -1773
rect 422 -1781 423 -1779
rect 429 -1775 430 -1773
rect 429 -1781 430 -1779
rect 436 -1775 437 -1773
rect 436 -1781 437 -1779
rect 443 -1775 444 -1773
rect 443 -1781 444 -1779
rect 450 -1775 451 -1773
rect 450 -1781 451 -1779
rect 457 -1775 458 -1773
rect 457 -1781 458 -1779
rect 464 -1775 465 -1773
rect 464 -1781 465 -1779
rect 471 -1775 472 -1773
rect 471 -1781 472 -1779
rect 481 -1775 482 -1773
rect 478 -1781 479 -1779
rect 481 -1781 482 -1779
rect 485 -1775 486 -1773
rect 485 -1781 486 -1779
rect 492 -1775 493 -1773
rect 492 -1781 493 -1779
rect 499 -1775 500 -1773
rect 499 -1781 500 -1779
rect 506 -1775 507 -1773
rect 506 -1781 507 -1779
rect 513 -1775 514 -1773
rect 516 -1775 517 -1773
rect 513 -1781 514 -1779
rect 516 -1781 517 -1779
rect 523 -1775 524 -1773
rect 520 -1781 521 -1779
rect 523 -1781 524 -1779
rect 527 -1775 528 -1773
rect 527 -1781 528 -1779
rect 530 -1781 531 -1779
rect 534 -1775 535 -1773
rect 534 -1781 535 -1779
rect 541 -1775 542 -1773
rect 541 -1781 542 -1779
rect 548 -1775 549 -1773
rect 548 -1781 549 -1779
rect 555 -1775 556 -1773
rect 558 -1775 559 -1773
rect 555 -1781 556 -1779
rect 558 -1781 559 -1779
rect 565 -1775 566 -1773
rect 562 -1781 563 -1779
rect 565 -1781 566 -1779
rect 569 -1775 570 -1773
rect 569 -1781 570 -1779
rect 576 -1775 577 -1773
rect 576 -1781 577 -1779
rect 583 -1775 584 -1773
rect 583 -1781 584 -1779
rect 590 -1775 591 -1773
rect 590 -1781 591 -1779
rect 597 -1775 598 -1773
rect 600 -1775 601 -1773
rect 597 -1781 598 -1779
rect 600 -1781 601 -1779
rect 604 -1775 605 -1773
rect 604 -1781 605 -1779
rect 611 -1775 612 -1773
rect 611 -1781 612 -1779
rect 618 -1775 619 -1773
rect 618 -1781 619 -1779
rect 625 -1775 626 -1773
rect 625 -1781 626 -1779
rect 632 -1775 633 -1773
rect 632 -1781 633 -1779
rect 639 -1775 640 -1773
rect 639 -1781 640 -1779
rect 646 -1775 647 -1773
rect 649 -1775 650 -1773
rect 646 -1781 647 -1779
rect 649 -1781 650 -1779
rect 653 -1775 654 -1773
rect 653 -1781 654 -1779
rect 660 -1775 661 -1773
rect 660 -1781 661 -1779
rect 667 -1775 668 -1773
rect 667 -1781 668 -1779
rect 674 -1775 675 -1773
rect 674 -1781 675 -1779
rect 681 -1775 682 -1773
rect 684 -1775 685 -1773
rect 681 -1781 682 -1779
rect 684 -1781 685 -1779
rect 688 -1775 689 -1773
rect 688 -1781 689 -1779
rect 695 -1775 696 -1773
rect 698 -1775 699 -1773
rect 695 -1781 696 -1779
rect 702 -1775 703 -1773
rect 702 -1781 703 -1779
rect 709 -1775 710 -1773
rect 709 -1781 710 -1779
rect 716 -1775 717 -1773
rect 716 -1781 717 -1779
rect 723 -1775 724 -1773
rect 723 -1781 724 -1779
rect 730 -1775 731 -1773
rect 730 -1781 731 -1779
rect 737 -1775 738 -1773
rect 740 -1775 741 -1773
rect 737 -1781 738 -1779
rect 744 -1775 745 -1773
rect 744 -1781 745 -1779
rect 751 -1775 752 -1773
rect 751 -1781 752 -1779
rect 758 -1775 759 -1773
rect 758 -1781 759 -1779
rect 765 -1775 766 -1773
rect 765 -1781 766 -1779
rect 772 -1775 773 -1773
rect 772 -1781 773 -1779
rect 779 -1775 780 -1773
rect 779 -1781 780 -1779
rect 786 -1775 787 -1773
rect 786 -1781 787 -1779
rect 793 -1775 794 -1773
rect 793 -1781 794 -1779
rect 800 -1775 801 -1773
rect 800 -1781 801 -1779
rect 810 -1775 811 -1773
rect 810 -1781 811 -1779
rect 814 -1775 815 -1773
rect 814 -1781 815 -1779
rect 821 -1775 822 -1773
rect 821 -1781 822 -1779
rect 831 -1775 832 -1773
rect 828 -1781 829 -1779
rect 831 -1781 832 -1779
rect 835 -1775 836 -1773
rect 835 -1781 836 -1779
rect 842 -1775 843 -1773
rect 842 -1781 843 -1779
rect 849 -1775 850 -1773
rect 849 -1781 850 -1779
rect 856 -1775 857 -1773
rect 856 -1781 857 -1779
rect 863 -1775 864 -1773
rect 863 -1781 864 -1779
rect 870 -1775 871 -1773
rect 870 -1781 871 -1779
rect 877 -1775 878 -1773
rect 877 -1781 878 -1779
rect 887 -1775 888 -1773
rect 884 -1781 885 -1779
rect 887 -1781 888 -1779
rect 891 -1775 892 -1773
rect 891 -1781 892 -1779
rect 898 -1775 899 -1773
rect 901 -1775 902 -1773
rect 905 -1775 906 -1773
rect 905 -1781 906 -1779
rect 912 -1775 913 -1773
rect 912 -1781 913 -1779
rect 919 -1775 920 -1773
rect 919 -1781 920 -1779
rect 926 -1775 927 -1773
rect 926 -1781 927 -1779
rect 933 -1775 934 -1773
rect 933 -1781 934 -1779
rect 943 -1775 944 -1773
rect 940 -1781 941 -1779
rect 943 -1781 944 -1779
rect 947 -1775 948 -1773
rect 947 -1781 948 -1779
rect 954 -1775 955 -1773
rect 954 -1781 955 -1779
rect 961 -1775 962 -1773
rect 961 -1781 962 -1779
rect 968 -1775 969 -1773
rect 968 -1781 969 -1779
rect 975 -1775 976 -1773
rect 975 -1781 976 -1779
rect 982 -1775 983 -1773
rect 985 -1775 986 -1773
rect 989 -1775 990 -1773
rect 989 -1781 990 -1779
rect 996 -1775 997 -1773
rect 996 -1781 997 -1779
rect 1003 -1775 1004 -1773
rect 1003 -1781 1004 -1779
rect 1010 -1775 1011 -1773
rect 1010 -1781 1011 -1779
rect 1017 -1775 1018 -1773
rect 1017 -1781 1018 -1779
rect 1024 -1775 1025 -1773
rect 1024 -1781 1025 -1779
rect 1031 -1775 1032 -1773
rect 1031 -1781 1032 -1779
rect 1038 -1775 1039 -1773
rect 1038 -1781 1039 -1779
rect 1045 -1775 1046 -1773
rect 1045 -1781 1046 -1779
rect 1052 -1775 1053 -1773
rect 1052 -1781 1053 -1779
rect 1059 -1775 1060 -1773
rect 1059 -1781 1060 -1779
rect 1066 -1775 1067 -1773
rect 1066 -1781 1067 -1779
rect 1073 -1775 1074 -1773
rect 1076 -1775 1077 -1773
rect 1073 -1781 1074 -1779
rect 1076 -1781 1077 -1779
rect 1080 -1775 1081 -1773
rect 1083 -1775 1084 -1773
rect 1080 -1781 1081 -1779
rect 1083 -1781 1084 -1779
rect 1087 -1775 1088 -1773
rect 1087 -1781 1088 -1779
rect 1094 -1775 1095 -1773
rect 1094 -1781 1095 -1779
rect 1101 -1775 1102 -1773
rect 1104 -1775 1105 -1773
rect 1104 -1781 1105 -1779
rect 1111 -1775 1112 -1773
rect 1108 -1781 1109 -1779
rect 1111 -1781 1112 -1779
rect 1115 -1775 1116 -1773
rect 1115 -1781 1116 -1779
rect 1122 -1775 1123 -1773
rect 1122 -1781 1123 -1779
rect 1129 -1775 1130 -1773
rect 1129 -1781 1130 -1779
rect 1136 -1775 1137 -1773
rect 1136 -1781 1137 -1779
rect 1143 -1775 1144 -1773
rect 1143 -1781 1144 -1779
rect 1150 -1775 1151 -1773
rect 1150 -1781 1151 -1779
rect 1157 -1775 1158 -1773
rect 1157 -1781 1158 -1779
rect 1164 -1775 1165 -1773
rect 1164 -1781 1165 -1779
rect 1171 -1775 1172 -1773
rect 1171 -1781 1172 -1779
rect 1178 -1775 1179 -1773
rect 1178 -1781 1179 -1779
rect 1185 -1775 1186 -1773
rect 1185 -1781 1186 -1779
rect 1192 -1775 1193 -1773
rect 1192 -1781 1193 -1779
rect 1199 -1775 1200 -1773
rect 1199 -1781 1200 -1779
rect 1206 -1775 1207 -1773
rect 1206 -1781 1207 -1779
rect 1213 -1775 1214 -1773
rect 1213 -1781 1214 -1779
rect 1220 -1775 1221 -1773
rect 1220 -1781 1221 -1779
rect 1227 -1775 1228 -1773
rect 1227 -1781 1228 -1779
rect 1234 -1775 1235 -1773
rect 1234 -1781 1235 -1779
rect 1241 -1775 1242 -1773
rect 1244 -1775 1245 -1773
rect 1241 -1781 1242 -1779
rect 1244 -1781 1245 -1779
rect 1248 -1775 1249 -1773
rect 1248 -1781 1249 -1779
rect 1255 -1775 1256 -1773
rect 1255 -1781 1256 -1779
rect 1262 -1775 1263 -1773
rect 1262 -1781 1263 -1779
rect 1269 -1775 1270 -1773
rect 1269 -1781 1270 -1779
rect 1276 -1775 1277 -1773
rect 1276 -1781 1277 -1779
rect 1283 -1775 1284 -1773
rect 1283 -1781 1284 -1779
rect 1290 -1775 1291 -1773
rect 1290 -1781 1291 -1779
rect 1297 -1775 1298 -1773
rect 1297 -1781 1298 -1779
rect 1304 -1775 1305 -1773
rect 1307 -1775 1308 -1773
rect 1304 -1781 1305 -1779
rect 1307 -1781 1308 -1779
rect 1311 -1775 1312 -1773
rect 1311 -1781 1312 -1779
rect 1318 -1775 1319 -1773
rect 1318 -1781 1319 -1779
rect 1321 -1781 1322 -1779
rect 1325 -1775 1326 -1773
rect 1325 -1781 1326 -1779
rect 1332 -1775 1333 -1773
rect 1332 -1781 1333 -1779
rect 1339 -1775 1340 -1773
rect 1339 -1781 1340 -1779
rect 1346 -1775 1347 -1773
rect 1346 -1781 1347 -1779
rect 1353 -1775 1354 -1773
rect 1356 -1775 1357 -1773
rect 1360 -1775 1361 -1773
rect 1363 -1775 1364 -1773
rect 1360 -1781 1361 -1779
rect 1363 -1781 1364 -1779
rect 1367 -1775 1368 -1773
rect 1367 -1781 1368 -1779
rect 1374 -1775 1375 -1773
rect 1374 -1781 1375 -1779
rect 1381 -1775 1382 -1773
rect 1381 -1781 1382 -1779
rect 1388 -1775 1389 -1773
rect 1388 -1781 1389 -1779
rect 1395 -1775 1396 -1773
rect 1395 -1781 1396 -1779
rect 1402 -1775 1403 -1773
rect 1402 -1781 1403 -1779
rect 1409 -1775 1410 -1773
rect 1409 -1781 1410 -1779
rect 1416 -1775 1417 -1773
rect 1416 -1781 1417 -1779
rect 1423 -1775 1424 -1773
rect 1423 -1781 1424 -1779
rect 1430 -1775 1431 -1773
rect 1430 -1781 1431 -1779
rect 1437 -1775 1438 -1773
rect 1437 -1781 1438 -1779
rect 1444 -1775 1445 -1773
rect 1444 -1781 1445 -1779
rect 1451 -1775 1452 -1773
rect 1451 -1781 1452 -1779
rect 1458 -1775 1459 -1773
rect 1458 -1781 1459 -1779
rect 1465 -1775 1466 -1773
rect 1468 -1775 1469 -1773
rect 1465 -1781 1466 -1779
rect 1468 -1781 1469 -1779
rect 1472 -1775 1473 -1773
rect 1472 -1781 1473 -1779
rect 1479 -1775 1480 -1773
rect 1479 -1781 1480 -1779
rect 1486 -1775 1487 -1773
rect 1486 -1781 1487 -1779
rect 1493 -1775 1494 -1773
rect 1493 -1781 1494 -1779
rect 1500 -1775 1501 -1773
rect 1500 -1781 1501 -1779
rect 1507 -1775 1508 -1773
rect 1507 -1781 1508 -1779
rect 1514 -1775 1515 -1773
rect 1514 -1781 1515 -1779
rect 1521 -1775 1522 -1773
rect 1521 -1781 1522 -1779
rect 1528 -1775 1529 -1773
rect 1528 -1781 1529 -1779
rect 1535 -1775 1536 -1773
rect 1535 -1781 1536 -1779
rect 1542 -1775 1543 -1773
rect 1542 -1781 1543 -1779
rect 1549 -1775 1550 -1773
rect 1549 -1781 1550 -1779
rect 1556 -1775 1557 -1773
rect 1556 -1781 1557 -1779
rect 1563 -1775 1564 -1773
rect 1563 -1781 1564 -1779
rect 1570 -1775 1571 -1773
rect 1570 -1781 1571 -1779
rect 1577 -1775 1578 -1773
rect 1577 -1781 1578 -1779
rect 1584 -1775 1585 -1773
rect 1584 -1781 1585 -1779
rect 1591 -1775 1592 -1773
rect 1591 -1781 1592 -1779
rect 1598 -1775 1599 -1773
rect 1598 -1781 1599 -1779
rect 1605 -1775 1606 -1773
rect 1605 -1781 1606 -1779
rect 1612 -1775 1613 -1773
rect 1612 -1781 1613 -1779
rect 1619 -1775 1620 -1773
rect 1619 -1781 1620 -1779
rect 1626 -1775 1627 -1773
rect 1626 -1781 1627 -1779
rect 1633 -1775 1634 -1773
rect 1633 -1781 1634 -1779
rect 1640 -1775 1641 -1773
rect 1640 -1781 1641 -1779
rect 1647 -1775 1648 -1773
rect 1647 -1781 1648 -1779
rect 1654 -1775 1655 -1773
rect 1654 -1781 1655 -1779
rect 1661 -1775 1662 -1773
rect 1661 -1781 1662 -1779
rect 1668 -1775 1669 -1773
rect 1668 -1781 1669 -1779
rect 1675 -1775 1676 -1773
rect 1675 -1781 1676 -1779
rect 1682 -1775 1683 -1773
rect 1682 -1781 1683 -1779
rect 1689 -1775 1690 -1773
rect 1689 -1781 1690 -1779
rect 1696 -1775 1697 -1773
rect 1696 -1781 1697 -1779
rect 1703 -1775 1704 -1773
rect 1703 -1781 1704 -1779
rect 1710 -1775 1711 -1773
rect 1710 -1781 1711 -1779
rect 1717 -1775 1718 -1773
rect 1717 -1781 1718 -1779
rect 1724 -1775 1725 -1773
rect 1724 -1781 1725 -1779
rect 1731 -1775 1732 -1773
rect 1731 -1781 1732 -1779
rect 1738 -1775 1739 -1773
rect 1738 -1781 1739 -1779
rect 1745 -1775 1746 -1773
rect 1745 -1781 1746 -1779
rect 1752 -1775 1753 -1773
rect 1752 -1781 1753 -1779
rect 1759 -1775 1760 -1773
rect 1759 -1781 1760 -1779
rect 1766 -1775 1767 -1773
rect 1766 -1781 1767 -1779
rect 1773 -1775 1774 -1773
rect 1773 -1781 1774 -1779
rect 1780 -1775 1781 -1773
rect 1780 -1781 1781 -1779
rect 1787 -1775 1788 -1773
rect 1787 -1781 1788 -1779
rect 1794 -1775 1795 -1773
rect 1794 -1781 1795 -1779
rect 1801 -1775 1802 -1773
rect 1801 -1781 1802 -1779
rect 1808 -1775 1809 -1773
rect 1808 -1781 1809 -1779
rect 1815 -1775 1816 -1773
rect 1815 -1781 1816 -1779
rect 1822 -1775 1823 -1773
rect 1822 -1781 1823 -1779
rect 1829 -1775 1830 -1773
rect 1829 -1781 1830 -1779
rect 1836 -1775 1837 -1773
rect 1836 -1781 1837 -1779
rect 1843 -1775 1844 -1773
rect 1843 -1781 1844 -1779
rect 1850 -1775 1851 -1773
rect 1850 -1781 1851 -1779
rect 1857 -1775 1858 -1773
rect 1857 -1781 1858 -1779
rect 1864 -1775 1865 -1773
rect 1864 -1781 1865 -1779
rect 1871 -1775 1872 -1773
rect 1871 -1781 1872 -1779
rect 1878 -1775 1879 -1773
rect 1878 -1781 1879 -1779
rect 1885 -1775 1886 -1773
rect 1885 -1781 1886 -1779
rect 1892 -1775 1893 -1773
rect 1892 -1781 1893 -1779
rect 1899 -1775 1900 -1773
rect 1899 -1781 1900 -1779
rect 1906 -1775 1907 -1773
rect 1906 -1781 1907 -1779
rect 1913 -1775 1914 -1773
rect 1913 -1781 1914 -1779
rect 1920 -1775 1921 -1773
rect 1920 -1781 1921 -1779
rect 1927 -1775 1928 -1773
rect 1927 -1781 1928 -1779
rect 1934 -1775 1935 -1773
rect 1937 -1775 1938 -1773
rect 1934 -1781 1935 -1779
rect 1941 -1775 1942 -1773
rect 1944 -1775 1945 -1773
rect 1941 -1781 1942 -1779
rect 1944 -1781 1945 -1779
rect 1948 -1775 1949 -1773
rect 1948 -1781 1949 -1779
rect 1955 -1775 1956 -1773
rect 1955 -1781 1956 -1779
rect 1962 -1775 1963 -1773
rect 1962 -1781 1963 -1779
rect 1969 -1775 1970 -1773
rect 1969 -1781 1970 -1779
rect 2018 -1775 2019 -1773
rect 2018 -1781 2019 -1779
rect 5 -1906 6 -1904
rect 16 -1900 17 -1898
rect 16 -1906 17 -1904
rect 23 -1900 24 -1898
rect 23 -1906 24 -1904
rect 30 -1900 31 -1898
rect 30 -1906 31 -1904
rect 37 -1900 38 -1898
rect 37 -1906 38 -1904
rect 44 -1900 45 -1898
rect 44 -1906 45 -1904
rect 51 -1900 52 -1898
rect 51 -1906 52 -1904
rect 58 -1900 59 -1898
rect 61 -1900 62 -1898
rect 61 -1906 62 -1904
rect 65 -1900 66 -1898
rect 65 -1906 66 -1904
rect 72 -1900 73 -1898
rect 72 -1906 73 -1904
rect 79 -1900 80 -1898
rect 79 -1906 80 -1904
rect 86 -1900 87 -1898
rect 86 -1906 87 -1904
rect 93 -1900 94 -1898
rect 93 -1906 94 -1904
rect 103 -1900 104 -1898
rect 100 -1906 101 -1904
rect 103 -1906 104 -1904
rect 107 -1900 108 -1898
rect 107 -1906 108 -1904
rect 114 -1900 115 -1898
rect 114 -1906 115 -1904
rect 121 -1900 122 -1898
rect 121 -1906 122 -1904
rect 128 -1900 129 -1898
rect 128 -1906 129 -1904
rect 135 -1900 136 -1898
rect 138 -1900 139 -1898
rect 135 -1906 136 -1904
rect 138 -1906 139 -1904
rect 142 -1900 143 -1898
rect 145 -1900 146 -1898
rect 142 -1906 143 -1904
rect 145 -1906 146 -1904
rect 149 -1900 150 -1898
rect 149 -1906 150 -1904
rect 156 -1900 157 -1898
rect 156 -1906 157 -1904
rect 163 -1900 164 -1898
rect 163 -1906 164 -1904
rect 170 -1900 171 -1898
rect 170 -1906 171 -1904
rect 177 -1900 178 -1898
rect 177 -1906 178 -1904
rect 184 -1900 185 -1898
rect 184 -1906 185 -1904
rect 191 -1900 192 -1898
rect 191 -1906 192 -1904
rect 198 -1900 199 -1898
rect 201 -1900 202 -1898
rect 198 -1906 199 -1904
rect 205 -1900 206 -1898
rect 205 -1906 206 -1904
rect 212 -1900 213 -1898
rect 212 -1906 213 -1904
rect 219 -1900 220 -1898
rect 219 -1906 220 -1904
rect 226 -1900 227 -1898
rect 226 -1906 227 -1904
rect 233 -1900 234 -1898
rect 233 -1906 234 -1904
rect 240 -1900 241 -1898
rect 240 -1906 241 -1904
rect 247 -1900 248 -1898
rect 247 -1906 248 -1904
rect 254 -1900 255 -1898
rect 254 -1906 255 -1904
rect 261 -1900 262 -1898
rect 261 -1906 262 -1904
rect 268 -1900 269 -1898
rect 268 -1906 269 -1904
rect 275 -1900 276 -1898
rect 275 -1906 276 -1904
rect 282 -1900 283 -1898
rect 282 -1906 283 -1904
rect 289 -1900 290 -1898
rect 289 -1906 290 -1904
rect 296 -1900 297 -1898
rect 296 -1906 297 -1904
rect 303 -1900 304 -1898
rect 303 -1906 304 -1904
rect 310 -1900 311 -1898
rect 310 -1906 311 -1904
rect 317 -1900 318 -1898
rect 317 -1906 318 -1904
rect 324 -1900 325 -1898
rect 324 -1906 325 -1904
rect 331 -1900 332 -1898
rect 331 -1906 332 -1904
rect 338 -1906 339 -1904
rect 345 -1900 346 -1898
rect 345 -1906 346 -1904
rect 352 -1900 353 -1898
rect 352 -1906 353 -1904
rect 359 -1900 360 -1898
rect 359 -1906 360 -1904
rect 366 -1900 367 -1898
rect 366 -1906 367 -1904
rect 373 -1900 374 -1898
rect 373 -1906 374 -1904
rect 380 -1900 381 -1898
rect 380 -1906 381 -1904
rect 387 -1900 388 -1898
rect 387 -1906 388 -1904
rect 394 -1900 395 -1898
rect 394 -1906 395 -1904
rect 401 -1900 402 -1898
rect 404 -1900 405 -1898
rect 408 -1900 409 -1898
rect 408 -1906 409 -1904
rect 415 -1900 416 -1898
rect 415 -1906 416 -1904
rect 422 -1900 423 -1898
rect 422 -1906 423 -1904
rect 429 -1900 430 -1898
rect 429 -1906 430 -1904
rect 436 -1900 437 -1898
rect 436 -1906 437 -1904
rect 443 -1900 444 -1898
rect 443 -1906 444 -1904
rect 450 -1900 451 -1898
rect 450 -1906 451 -1904
rect 457 -1900 458 -1898
rect 457 -1906 458 -1904
rect 464 -1900 465 -1898
rect 464 -1906 465 -1904
rect 471 -1900 472 -1898
rect 471 -1906 472 -1904
rect 478 -1900 479 -1898
rect 481 -1906 482 -1904
rect 485 -1900 486 -1898
rect 488 -1900 489 -1898
rect 485 -1906 486 -1904
rect 488 -1906 489 -1904
rect 492 -1900 493 -1898
rect 492 -1906 493 -1904
rect 499 -1900 500 -1898
rect 499 -1906 500 -1904
rect 509 -1900 510 -1898
rect 506 -1906 507 -1904
rect 509 -1906 510 -1904
rect 513 -1900 514 -1898
rect 513 -1906 514 -1904
rect 520 -1900 521 -1898
rect 520 -1906 521 -1904
rect 527 -1900 528 -1898
rect 530 -1900 531 -1898
rect 527 -1906 528 -1904
rect 534 -1900 535 -1898
rect 534 -1906 535 -1904
rect 541 -1900 542 -1898
rect 541 -1906 542 -1904
rect 548 -1900 549 -1898
rect 548 -1906 549 -1904
rect 555 -1900 556 -1898
rect 555 -1906 556 -1904
rect 562 -1900 563 -1898
rect 562 -1906 563 -1904
rect 569 -1900 570 -1898
rect 569 -1906 570 -1904
rect 579 -1900 580 -1898
rect 579 -1906 580 -1904
rect 583 -1900 584 -1898
rect 583 -1906 584 -1904
rect 590 -1900 591 -1898
rect 590 -1906 591 -1904
rect 597 -1900 598 -1898
rect 597 -1906 598 -1904
rect 604 -1900 605 -1898
rect 604 -1906 605 -1904
rect 611 -1900 612 -1898
rect 614 -1900 615 -1898
rect 611 -1906 612 -1904
rect 614 -1906 615 -1904
rect 618 -1900 619 -1898
rect 618 -1906 619 -1904
rect 625 -1900 626 -1898
rect 625 -1906 626 -1904
rect 632 -1900 633 -1898
rect 632 -1906 633 -1904
rect 639 -1900 640 -1898
rect 639 -1906 640 -1904
rect 646 -1900 647 -1898
rect 646 -1906 647 -1904
rect 653 -1900 654 -1898
rect 653 -1906 654 -1904
rect 660 -1900 661 -1898
rect 660 -1906 661 -1904
rect 667 -1900 668 -1898
rect 674 -1900 675 -1898
rect 674 -1906 675 -1904
rect 681 -1900 682 -1898
rect 681 -1906 682 -1904
rect 691 -1900 692 -1898
rect 688 -1906 689 -1904
rect 691 -1906 692 -1904
rect 695 -1900 696 -1898
rect 695 -1906 696 -1904
rect 702 -1900 703 -1898
rect 702 -1906 703 -1904
rect 709 -1900 710 -1898
rect 709 -1906 710 -1904
rect 716 -1900 717 -1898
rect 719 -1900 720 -1898
rect 716 -1906 717 -1904
rect 719 -1906 720 -1904
rect 723 -1900 724 -1898
rect 723 -1906 724 -1904
rect 726 -1906 727 -1904
rect 730 -1900 731 -1898
rect 730 -1906 731 -1904
rect 737 -1900 738 -1898
rect 737 -1906 738 -1904
rect 744 -1900 745 -1898
rect 744 -1906 745 -1904
rect 751 -1900 752 -1898
rect 751 -1906 752 -1904
rect 758 -1900 759 -1898
rect 758 -1906 759 -1904
rect 765 -1900 766 -1898
rect 768 -1900 769 -1898
rect 765 -1906 766 -1904
rect 768 -1906 769 -1904
rect 772 -1900 773 -1898
rect 772 -1906 773 -1904
rect 775 -1906 776 -1904
rect 779 -1900 780 -1898
rect 779 -1906 780 -1904
rect 786 -1900 787 -1898
rect 786 -1906 787 -1904
rect 793 -1900 794 -1898
rect 793 -1906 794 -1904
rect 800 -1900 801 -1898
rect 800 -1906 801 -1904
rect 807 -1900 808 -1898
rect 807 -1906 808 -1904
rect 814 -1900 815 -1898
rect 814 -1906 815 -1904
rect 821 -1900 822 -1898
rect 821 -1906 822 -1904
rect 828 -1900 829 -1898
rect 828 -1906 829 -1904
rect 835 -1900 836 -1898
rect 835 -1906 836 -1904
rect 842 -1900 843 -1898
rect 842 -1906 843 -1904
rect 849 -1900 850 -1898
rect 849 -1906 850 -1904
rect 856 -1900 857 -1898
rect 856 -1906 857 -1904
rect 863 -1900 864 -1898
rect 863 -1906 864 -1904
rect 870 -1900 871 -1898
rect 870 -1906 871 -1904
rect 877 -1900 878 -1898
rect 877 -1906 878 -1904
rect 884 -1900 885 -1898
rect 887 -1900 888 -1898
rect 884 -1906 885 -1904
rect 887 -1906 888 -1904
rect 891 -1900 892 -1898
rect 891 -1906 892 -1904
rect 898 -1900 899 -1898
rect 898 -1906 899 -1904
rect 905 -1900 906 -1898
rect 908 -1900 909 -1898
rect 905 -1906 906 -1904
rect 908 -1906 909 -1904
rect 912 -1900 913 -1898
rect 912 -1906 913 -1904
rect 919 -1900 920 -1898
rect 919 -1906 920 -1904
rect 926 -1900 927 -1898
rect 926 -1906 927 -1904
rect 933 -1900 934 -1898
rect 936 -1900 937 -1898
rect 933 -1906 934 -1904
rect 936 -1906 937 -1904
rect 940 -1900 941 -1898
rect 940 -1906 941 -1904
rect 947 -1900 948 -1898
rect 947 -1906 948 -1904
rect 954 -1900 955 -1898
rect 954 -1906 955 -1904
rect 961 -1900 962 -1898
rect 961 -1906 962 -1904
rect 968 -1900 969 -1898
rect 968 -1906 969 -1904
rect 975 -1900 976 -1898
rect 975 -1906 976 -1904
rect 982 -1900 983 -1898
rect 985 -1900 986 -1898
rect 982 -1906 983 -1904
rect 985 -1906 986 -1904
rect 989 -1900 990 -1898
rect 989 -1906 990 -1904
rect 996 -1900 997 -1898
rect 996 -1906 997 -1904
rect 1003 -1900 1004 -1898
rect 1003 -1906 1004 -1904
rect 1010 -1900 1011 -1898
rect 1010 -1906 1011 -1904
rect 1017 -1900 1018 -1898
rect 1017 -1906 1018 -1904
rect 1024 -1900 1025 -1898
rect 1024 -1906 1025 -1904
rect 1027 -1906 1028 -1904
rect 1031 -1900 1032 -1898
rect 1031 -1906 1032 -1904
rect 1038 -1900 1039 -1898
rect 1038 -1906 1039 -1904
rect 1045 -1900 1046 -1898
rect 1045 -1906 1046 -1904
rect 1052 -1900 1053 -1898
rect 1052 -1906 1053 -1904
rect 1059 -1900 1060 -1898
rect 1059 -1906 1060 -1904
rect 1066 -1900 1067 -1898
rect 1066 -1906 1067 -1904
rect 1073 -1900 1074 -1898
rect 1073 -1906 1074 -1904
rect 1080 -1900 1081 -1898
rect 1080 -1906 1081 -1904
rect 1090 -1900 1091 -1898
rect 1087 -1906 1088 -1904
rect 1090 -1906 1091 -1904
rect 1094 -1900 1095 -1898
rect 1094 -1906 1095 -1904
rect 1101 -1900 1102 -1898
rect 1104 -1900 1105 -1898
rect 1104 -1906 1105 -1904
rect 1108 -1900 1109 -1898
rect 1111 -1900 1112 -1898
rect 1108 -1906 1109 -1904
rect 1111 -1906 1112 -1904
rect 1115 -1900 1116 -1898
rect 1115 -1906 1116 -1904
rect 1122 -1900 1123 -1898
rect 1125 -1900 1126 -1898
rect 1122 -1906 1123 -1904
rect 1129 -1900 1130 -1898
rect 1129 -1906 1130 -1904
rect 1136 -1900 1137 -1898
rect 1136 -1906 1137 -1904
rect 1143 -1900 1144 -1898
rect 1143 -1906 1144 -1904
rect 1150 -1900 1151 -1898
rect 1153 -1900 1154 -1898
rect 1150 -1906 1151 -1904
rect 1153 -1906 1154 -1904
rect 1157 -1900 1158 -1898
rect 1157 -1906 1158 -1904
rect 1164 -1900 1165 -1898
rect 1164 -1906 1165 -1904
rect 1171 -1900 1172 -1898
rect 1171 -1906 1172 -1904
rect 1178 -1900 1179 -1898
rect 1178 -1906 1179 -1904
rect 1185 -1900 1186 -1898
rect 1185 -1906 1186 -1904
rect 1192 -1900 1193 -1898
rect 1192 -1906 1193 -1904
rect 1199 -1900 1200 -1898
rect 1199 -1906 1200 -1904
rect 1209 -1900 1210 -1898
rect 1206 -1906 1207 -1904
rect 1209 -1906 1210 -1904
rect 1213 -1900 1214 -1898
rect 1213 -1906 1214 -1904
rect 1216 -1906 1217 -1904
rect 1220 -1900 1221 -1898
rect 1223 -1900 1224 -1898
rect 1220 -1906 1221 -1904
rect 1223 -1906 1224 -1904
rect 1227 -1900 1228 -1898
rect 1227 -1906 1228 -1904
rect 1234 -1900 1235 -1898
rect 1234 -1906 1235 -1904
rect 1241 -1900 1242 -1898
rect 1241 -1906 1242 -1904
rect 1248 -1900 1249 -1898
rect 1248 -1906 1249 -1904
rect 1255 -1900 1256 -1898
rect 1255 -1906 1256 -1904
rect 1262 -1900 1263 -1898
rect 1262 -1906 1263 -1904
rect 1269 -1900 1270 -1898
rect 1269 -1906 1270 -1904
rect 1276 -1906 1277 -1904
rect 1279 -1906 1280 -1904
rect 1283 -1900 1284 -1898
rect 1283 -1906 1284 -1904
rect 1290 -1900 1291 -1898
rect 1290 -1906 1291 -1904
rect 1297 -1900 1298 -1898
rect 1297 -1906 1298 -1904
rect 1304 -1900 1305 -1898
rect 1304 -1906 1305 -1904
rect 1311 -1900 1312 -1898
rect 1311 -1906 1312 -1904
rect 1318 -1900 1319 -1898
rect 1318 -1906 1319 -1904
rect 1325 -1900 1326 -1898
rect 1325 -1906 1326 -1904
rect 1332 -1900 1333 -1898
rect 1332 -1906 1333 -1904
rect 1339 -1900 1340 -1898
rect 1339 -1906 1340 -1904
rect 1346 -1900 1347 -1898
rect 1346 -1906 1347 -1904
rect 1353 -1900 1354 -1898
rect 1353 -1906 1354 -1904
rect 1360 -1900 1361 -1898
rect 1360 -1906 1361 -1904
rect 1367 -1900 1368 -1898
rect 1367 -1906 1368 -1904
rect 1374 -1900 1375 -1898
rect 1374 -1906 1375 -1904
rect 1381 -1900 1382 -1898
rect 1381 -1906 1382 -1904
rect 1388 -1900 1389 -1898
rect 1388 -1906 1389 -1904
rect 1395 -1900 1396 -1898
rect 1395 -1906 1396 -1904
rect 1402 -1900 1403 -1898
rect 1402 -1906 1403 -1904
rect 1409 -1900 1410 -1898
rect 1409 -1906 1410 -1904
rect 1416 -1900 1417 -1898
rect 1416 -1906 1417 -1904
rect 1423 -1900 1424 -1898
rect 1423 -1906 1424 -1904
rect 1430 -1900 1431 -1898
rect 1430 -1906 1431 -1904
rect 1437 -1900 1438 -1898
rect 1437 -1906 1438 -1904
rect 1444 -1900 1445 -1898
rect 1444 -1906 1445 -1904
rect 1451 -1900 1452 -1898
rect 1451 -1906 1452 -1904
rect 1458 -1900 1459 -1898
rect 1458 -1906 1459 -1904
rect 1465 -1900 1466 -1898
rect 1465 -1906 1466 -1904
rect 1472 -1900 1473 -1898
rect 1472 -1906 1473 -1904
rect 1479 -1900 1480 -1898
rect 1479 -1906 1480 -1904
rect 1486 -1900 1487 -1898
rect 1486 -1906 1487 -1904
rect 1493 -1900 1494 -1898
rect 1493 -1906 1494 -1904
rect 1500 -1900 1501 -1898
rect 1500 -1906 1501 -1904
rect 1507 -1900 1508 -1898
rect 1507 -1906 1508 -1904
rect 1514 -1900 1515 -1898
rect 1514 -1906 1515 -1904
rect 1521 -1900 1522 -1898
rect 1521 -1906 1522 -1904
rect 1528 -1900 1529 -1898
rect 1528 -1906 1529 -1904
rect 1535 -1900 1536 -1898
rect 1535 -1906 1536 -1904
rect 1542 -1900 1543 -1898
rect 1542 -1906 1543 -1904
rect 1549 -1900 1550 -1898
rect 1549 -1906 1550 -1904
rect 1556 -1900 1557 -1898
rect 1556 -1906 1557 -1904
rect 1563 -1900 1564 -1898
rect 1566 -1900 1567 -1898
rect 1566 -1906 1567 -1904
rect 1570 -1900 1571 -1898
rect 1570 -1906 1571 -1904
rect 1577 -1900 1578 -1898
rect 1577 -1906 1578 -1904
rect 1584 -1900 1585 -1898
rect 1584 -1906 1585 -1904
rect 1591 -1900 1592 -1898
rect 1591 -1906 1592 -1904
rect 1598 -1900 1599 -1898
rect 1598 -1906 1599 -1904
rect 1605 -1900 1606 -1898
rect 1605 -1906 1606 -1904
rect 1612 -1900 1613 -1898
rect 1612 -1906 1613 -1904
rect 1619 -1900 1620 -1898
rect 1619 -1906 1620 -1904
rect 1626 -1900 1627 -1898
rect 1626 -1906 1627 -1904
rect 1633 -1900 1634 -1898
rect 1633 -1906 1634 -1904
rect 1640 -1900 1641 -1898
rect 1640 -1906 1641 -1904
rect 1647 -1900 1648 -1898
rect 1647 -1906 1648 -1904
rect 1654 -1900 1655 -1898
rect 1654 -1906 1655 -1904
rect 1661 -1900 1662 -1898
rect 1661 -1906 1662 -1904
rect 1668 -1900 1669 -1898
rect 1668 -1906 1669 -1904
rect 1675 -1900 1676 -1898
rect 1675 -1906 1676 -1904
rect 1682 -1900 1683 -1898
rect 1682 -1906 1683 -1904
rect 1689 -1900 1690 -1898
rect 1689 -1906 1690 -1904
rect 1696 -1900 1697 -1898
rect 1696 -1906 1697 -1904
rect 1703 -1900 1704 -1898
rect 1703 -1906 1704 -1904
rect 1710 -1900 1711 -1898
rect 1710 -1906 1711 -1904
rect 1717 -1900 1718 -1898
rect 1717 -1906 1718 -1904
rect 1724 -1900 1725 -1898
rect 1724 -1906 1725 -1904
rect 1731 -1900 1732 -1898
rect 1731 -1906 1732 -1904
rect 1738 -1900 1739 -1898
rect 1738 -1906 1739 -1904
rect 1745 -1900 1746 -1898
rect 1745 -1906 1746 -1904
rect 1752 -1900 1753 -1898
rect 1752 -1906 1753 -1904
rect 1759 -1900 1760 -1898
rect 1759 -1906 1760 -1904
rect 1766 -1900 1767 -1898
rect 1766 -1906 1767 -1904
rect 1773 -1900 1774 -1898
rect 1773 -1906 1774 -1904
rect 1780 -1900 1781 -1898
rect 1780 -1906 1781 -1904
rect 1787 -1900 1788 -1898
rect 1787 -1906 1788 -1904
rect 1794 -1900 1795 -1898
rect 1794 -1906 1795 -1904
rect 1801 -1900 1802 -1898
rect 1801 -1906 1802 -1904
rect 1808 -1900 1809 -1898
rect 1808 -1906 1809 -1904
rect 1815 -1900 1816 -1898
rect 1815 -1906 1816 -1904
rect 1822 -1900 1823 -1898
rect 1822 -1906 1823 -1904
rect 1829 -1900 1830 -1898
rect 1829 -1906 1830 -1904
rect 1836 -1900 1837 -1898
rect 1836 -1906 1837 -1904
rect 1843 -1900 1844 -1898
rect 1843 -1906 1844 -1904
rect 1850 -1900 1851 -1898
rect 1850 -1906 1851 -1904
rect 1857 -1900 1858 -1898
rect 1857 -1906 1858 -1904
rect 1864 -1900 1865 -1898
rect 1864 -1906 1865 -1904
rect 1871 -1900 1872 -1898
rect 1871 -1906 1872 -1904
rect 1878 -1900 1879 -1898
rect 1878 -1906 1879 -1904
rect 1885 -1900 1886 -1898
rect 1885 -1906 1886 -1904
rect 1892 -1900 1893 -1898
rect 1892 -1906 1893 -1904
rect 1899 -1900 1900 -1898
rect 1899 -1906 1900 -1904
rect 1906 -1900 1907 -1898
rect 1906 -1906 1907 -1904
rect 1913 -1900 1914 -1898
rect 1913 -1906 1914 -1904
rect 1920 -1900 1921 -1898
rect 1920 -1906 1921 -1904
rect 1927 -1900 1928 -1898
rect 1927 -1906 1928 -1904
rect 1934 -1900 1935 -1898
rect 1934 -1906 1935 -1904
rect 1941 -1900 1942 -1898
rect 1941 -1906 1942 -1904
rect 1948 -1900 1949 -1898
rect 1948 -1906 1949 -1904
rect 1955 -1900 1956 -1898
rect 1955 -1906 1956 -1904
rect 1962 -1900 1963 -1898
rect 1962 -1906 1963 -1904
rect 1969 -1900 1970 -1898
rect 1969 -1906 1970 -1904
rect 1976 -1900 1977 -1898
rect 1976 -1906 1977 -1904
rect 1983 -1900 1984 -1898
rect 1983 -1906 1984 -1904
rect 1990 -1900 1991 -1898
rect 1990 -1906 1991 -1904
rect 1997 -1900 1998 -1898
rect 1997 -1906 1998 -1904
rect 2004 -1900 2005 -1898
rect 2004 -1906 2005 -1904
rect 2011 -1900 2012 -1898
rect 2014 -1900 2015 -1898
rect 2011 -1906 2012 -1904
rect 2018 -1900 2019 -1898
rect 2018 -1906 2019 -1904
rect 2025 -1900 2026 -1898
rect 2025 -1906 2026 -1904
rect 2 -2047 3 -2045
rect 2 -2053 3 -2051
rect 9 -2047 10 -2045
rect 9 -2053 10 -2051
rect 16 -2047 17 -2045
rect 16 -2053 17 -2051
rect 23 -2047 24 -2045
rect 23 -2053 24 -2051
rect 30 -2047 31 -2045
rect 30 -2053 31 -2051
rect 37 -2047 38 -2045
rect 37 -2053 38 -2051
rect 44 -2047 45 -2045
rect 44 -2053 45 -2051
rect 51 -2047 52 -2045
rect 51 -2053 52 -2051
rect 58 -2047 59 -2045
rect 58 -2053 59 -2051
rect 68 -2047 69 -2045
rect 65 -2053 66 -2051
rect 68 -2053 69 -2051
rect 72 -2047 73 -2045
rect 72 -2053 73 -2051
rect 79 -2047 80 -2045
rect 79 -2053 80 -2051
rect 86 -2047 87 -2045
rect 86 -2053 87 -2051
rect 93 -2047 94 -2045
rect 93 -2053 94 -2051
rect 100 -2047 101 -2045
rect 100 -2053 101 -2051
rect 107 -2047 108 -2045
rect 107 -2053 108 -2051
rect 114 -2047 115 -2045
rect 114 -2053 115 -2051
rect 117 -2053 118 -2051
rect 121 -2047 122 -2045
rect 121 -2053 122 -2051
rect 128 -2047 129 -2045
rect 128 -2053 129 -2051
rect 135 -2047 136 -2045
rect 135 -2053 136 -2051
rect 142 -2047 143 -2045
rect 145 -2047 146 -2045
rect 142 -2053 143 -2051
rect 145 -2053 146 -2051
rect 149 -2047 150 -2045
rect 149 -2053 150 -2051
rect 156 -2047 157 -2045
rect 156 -2053 157 -2051
rect 163 -2047 164 -2045
rect 163 -2053 164 -2051
rect 170 -2047 171 -2045
rect 170 -2053 171 -2051
rect 177 -2047 178 -2045
rect 177 -2053 178 -2051
rect 184 -2047 185 -2045
rect 184 -2053 185 -2051
rect 191 -2047 192 -2045
rect 191 -2053 192 -2051
rect 198 -2047 199 -2045
rect 198 -2053 199 -2051
rect 205 -2047 206 -2045
rect 205 -2053 206 -2051
rect 212 -2047 213 -2045
rect 212 -2053 213 -2051
rect 219 -2047 220 -2045
rect 222 -2047 223 -2045
rect 219 -2053 220 -2051
rect 222 -2053 223 -2051
rect 226 -2047 227 -2045
rect 226 -2053 227 -2051
rect 233 -2047 234 -2045
rect 233 -2053 234 -2051
rect 243 -2047 244 -2045
rect 243 -2053 244 -2051
rect 247 -2047 248 -2045
rect 247 -2053 248 -2051
rect 254 -2047 255 -2045
rect 254 -2053 255 -2051
rect 261 -2047 262 -2045
rect 261 -2053 262 -2051
rect 268 -2047 269 -2045
rect 268 -2053 269 -2051
rect 275 -2047 276 -2045
rect 275 -2053 276 -2051
rect 282 -2047 283 -2045
rect 282 -2053 283 -2051
rect 289 -2047 290 -2045
rect 289 -2053 290 -2051
rect 296 -2047 297 -2045
rect 296 -2053 297 -2051
rect 303 -2047 304 -2045
rect 303 -2053 304 -2051
rect 310 -2047 311 -2045
rect 313 -2047 314 -2045
rect 310 -2053 311 -2051
rect 313 -2053 314 -2051
rect 317 -2047 318 -2045
rect 317 -2053 318 -2051
rect 324 -2047 325 -2045
rect 324 -2053 325 -2051
rect 331 -2047 332 -2045
rect 331 -2053 332 -2051
rect 341 -2047 342 -2045
rect 338 -2053 339 -2051
rect 345 -2047 346 -2045
rect 345 -2053 346 -2051
rect 352 -2047 353 -2045
rect 352 -2053 353 -2051
rect 359 -2047 360 -2045
rect 359 -2053 360 -2051
rect 366 -2047 367 -2045
rect 366 -2053 367 -2051
rect 373 -2047 374 -2045
rect 373 -2053 374 -2051
rect 380 -2047 381 -2045
rect 380 -2053 381 -2051
rect 387 -2047 388 -2045
rect 387 -2053 388 -2051
rect 394 -2047 395 -2045
rect 394 -2053 395 -2051
rect 401 -2047 402 -2045
rect 401 -2053 402 -2051
rect 408 -2047 409 -2045
rect 408 -2053 409 -2051
rect 415 -2047 416 -2045
rect 415 -2053 416 -2051
rect 422 -2047 423 -2045
rect 422 -2053 423 -2051
rect 429 -2047 430 -2045
rect 429 -2053 430 -2051
rect 436 -2047 437 -2045
rect 436 -2053 437 -2051
rect 443 -2047 444 -2045
rect 443 -2053 444 -2051
rect 450 -2053 451 -2051
rect 453 -2053 454 -2051
rect 457 -2047 458 -2045
rect 457 -2053 458 -2051
rect 464 -2047 465 -2045
rect 464 -2053 465 -2051
rect 471 -2047 472 -2045
rect 471 -2053 472 -2051
rect 478 -2047 479 -2045
rect 478 -2053 479 -2051
rect 485 -2047 486 -2045
rect 485 -2053 486 -2051
rect 492 -2047 493 -2045
rect 492 -2053 493 -2051
rect 499 -2047 500 -2045
rect 499 -2053 500 -2051
rect 506 -2047 507 -2045
rect 506 -2053 507 -2051
rect 513 -2047 514 -2045
rect 513 -2053 514 -2051
rect 520 -2047 521 -2045
rect 520 -2053 521 -2051
rect 527 -2047 528 -2045
rect 530 -2047 531 -2045
rect 527 -2053 528 -2051
rect 530 -2053 531 -2051
rect 534 -2047 535 -2045
rect 537 -2047 538 -2045
rect 534 -2053 535 -2051
rect 537 -2053 538 -2051
rect 541 -2047 542 -2045
rect 541 -2053 542 -2051
rect 548 -2047 549 -2045
rect 548 -2053 549 -2051
rect 555 -2047 556 -2045
rect 555 -2053 556 -2051
rect 562 -2047 563 -2045
rect 562 -2053 563 -2051
rect 569 -2047 570 -2045
rect 569 -2053 570 -2051
rect 576 -2047 577 -2045
rect 576 -2053 577 -2051
rect 583 -2047 584 -2045
rect 583 -2053 584 -2051
rect 590 -2047 591 -2045
rect 590 -2053 591 -2051
rect 597 -2047 598 -2045
rect 597 -2053 598 -2051
rect 604 -2047 605 -2045
rect 604 -2053 605 -2051
rect 611 -2047 612 -2045
rect 611 -2053 612 -2051
rect 618 -2047 619 -2045
rect 618 -2053 619 -2051
rect 625 -2047 626 -2045
rect 625 -2053 626 -2051
rect 632 -2047 633 -2045
rect 632 -2053 633 -2051
rect 639 -2047 640 -2045
rect 639 -2053 640 -2051
rect 646 -2047 647 -2045
rect 646 -2053 647 -2051
rect 653 -2047 654 -2045
rect 653 -2053 654 -2051
rect 660 -2047 661 -2045
rect 660 -2053 661 -2051
rect 667 -2053 668 -2051
rect 674 -2047 675 -2045
rect 674 -2053 675 -2051
rect 681 -2047 682 -2045
rect 681 -2053 682 -2051
rect 688 -2047 689 -2045
rect 688 -2053 689 -2051
rect 698 -2047 699 -2045
rect 695 -2053 696 -2051
rect 698 -2053 699 -2051
rect 702 -2047 703 -2045
rect 702 -2053 703 -2051
rect 709 -2047 710 -2045
rect 709 -2053 710 -2051
rect 716 -2047 717 -2045
rect 716 -2053 717 -2051
rect 723 -2047 724 -2045
rect 723 -2053 724 -2051
rect 726 -2053 727 -2051
rect 730 -2047 731 -2045
rect 733 -2047 734 -2045
rect 730 -2053 731 -2051
rect 733 -2053 734 -2051
rect 737 -2047 738 -2045
rect 737 -2053 738 -2051
rect 744 -2047 745 -2045
rect 744 -2053 745 -2051
rect 751 -2047 752 -2045
rect 754 -2047 755 -2045
rect 751 -2053 752 -2051
rect 754 -2053 755 -2051
rect 758 -2047 759 -2045
rect 761 -2047 762 -2045
rect 758 -2053 759 -2051
rect 761 -2053 762 -2051
rect 765 -2047 766 -2045
rect 765 -2053 766 -2051
rect 772 -2047 773 -2045
rect 775 -2047 776 -2045
rect 772 -2053 773 -2051
rect 779 -2047 780 -2045
rect 779 -2053 780 -2051
rect 786 -2047 787 -2045
rect 786 -2053 787 -2051
rect 793 -2047 794 -2045
rect 793 -2053 794 -2051
rect 800 -2047 801 -2045
rect 800 -2053 801 -2051
rect 807 -2047 808 -2045
rect 807 -2053 808 -2051
rect 814 -2047 815 -2045
rect 817 -2047 818 -2045
rect 814 -2053 815 -2051
rect 817 -2053 818 -2051
rect 821 -2047 822 -2045
rect 821 -2053 822 -2051
rect 828 -2047 829 -2045
rect 828 -2053 829 -2051
rect 835 -2047 836 -2045
rect 835 -2053 836 -2051
rect 842 -2047 843 -2045
rect 845 -2047 846 -2045
rect 842 -2053 843 -2051
rect 845 -2053 846 -2051
rect 849 -2047 850 -2045
rect 849 -2053 850 -2051
rect 852 -2053 853 -2051
rect 856 -2047 857 -2045
rect 856 -2053 857 -2051
rect 863 -2047 864 -2045
rect 866 -2047 867 -2045
rect 863 -2053 864 -2051
rect 866 -2053 867 -2051
rect 870 -2047 871 -2045
rect 870 -2053 871 -2051
rect 877 -2047 878 -2045
rect 880 -2047 881 -2045
rect 877 -2053 878 -2051
rect 880 -2053 881 -2051
rect 884 -2047 885 -2045
rect 884 -2053 885 -2051
rect 891 -2047 892 -2045
rect 894 -2047 895 -2045
rect 891 -2053 892 -2051
rect 894 -2053 895 -2051
rect 898 -2047 899 -2045
rect 898 -2053 899 -2051
rect 905 -2047 906 -2045
rect 905 -2053 906 -2051
rect 912 -2047 913 -2045
rect 912 -2053 913 -2051
rect 919 -2047 920 -2045
rect 922 -2047 923 -2045
rect 919 -2053 920 -2051
rect 922 -2053 923 -2051
rect 926 -2047 927 -2045
rect 926 -2053 927 -2051
rect 933 -2047 934 -2045
rect 933 -2053 934 -2051
rect 940 -2047 941 -2045
rect 940 -2053 941 -2051
rect 947 -2047 948 -2045
rect 947 -2053 948 -2051
rect 954 -2047 955 -2045
rect 954 -2053 955 -2051
rect 961 -2047 962 -2045
rect 964 -2047 965 -2045
rect 961 -2053 962 -2051
rect 964 -2053 965 -2051
rect 968 -2047 969 -2045
rect 968 -2053 969 -2051
rect 971 -2053 972 -2051
rect 975 -2047 976 -2045
rect 975 -2053 976 -2051
rect 982 -2047 983 -2045
rect 982 -2053 983 -2051
rect 989 -2047 990 -2045
rect 989 -2053 990 -2051
rect 996 -2047 997 -2045
rect 996 -2053 997 -2051
rect 1003 -2047 1004 -2045
rect 1003 -2053 1004 -2051
rect 1010 -2047 1011 -2045
rect 1010 -2053 1011 -2051
rect 1017 -2047 1018 -2045
rect 1017 -2053 1018 -2051
rect 1024 -2047 1025 -2045
rect 1024 -2053 1025 -2051
rect 1031 -2047 1032 -2045
rect 1031 -2053 1032 -2051
rect 1038 -2047 1039 -2045
rect 1038 -2053 1039 -2051
rect 1045 -2047 1046 -2045
rect 1045 -2053 1046 -2051
rect 1052 -2047 1053 -2045
rect 1052 -2053 1053 -2051
rect 1059 -2047 1060 -2045
rect 1059 -2053 1060 -2051
rect 1066 -2047 1067 -2045
rect 1066 -2053 1067 -2051
rect 1073 -2047 1074 -2045
rect 1073 -2053 1074 -2051
rect 1080 -2047 1081 -2045
rect 1080 -2053 1081 -2051
rect 1087 -2047 1088 -2045
rect 1087 -2053 1088 -2051
rect 1090 -2053 1091 -2051
rect 1094 -2047 1095 -2045
rect 1094 -2053 1095 -2051
rect 1101 -2047 1102 -2045
rect 1101 -2053 1102 -2051
rect 1108 -2047 1109 -2045
rect 1111 -2047 1112 -2045
rect 1108 -2053 1109 -2051
rect 1111 -2053 1112 -2051
rect 1115 -2047 1116 -2045
rect 1115 -2053 1116 -2051
rect 1122 -2047 1123 -2045
rect 1122 -2053 1123 -2051
rect 1129 -2047 1130 -2045
rect 1129 -2053 1130 -2051
rect 1136 -2047 1137 -2045
rect 1136 -2053 1137 -2051
rect 1143 -2047 1144 -2045
rect 1143 -2053 1144 -2051
rect 1150 -2047 1151 -2045
rect 1150 -2053 1151 -2051
rect 1157 -2047 1158 -2045
rect 1157 -2053 1158 -2051
rect 1164 -2047 1165 -2045
rect 1164 -2053 1165 -2051
rect 1171 -2047 1172 -2045
rect 1171 -2053 1172 -2051
rect 1178 -2047 1179 -2045
rect 1178 -2053 1179 -2051
rect 1185 -2047 1186 -2045
rect 1185 -2053 1186 -2051
rect 1192 -2047 1193 -2045
rect 1192 -2053 1193 -2051
rect 1199 -2047 1200 -2045
rect 1199 -2053 1200 -2051
rect 1206 -2047 1207 -2045
rect 1206 -2053 1207 -2051
rect 1213 -2047 1214 -2045
rect 1216 -2047 1217 -2045
rect 1213 -2053 1214 -2051
rect 1220 -2047 1221 -2045
rect 1220 -2053 1221 -2051
rect 1227 -2047 1228 -2045
rect 1227 -2053 1228 -2051
rect 1237 -2047 1238 -2045
rect 1237 -2053 1238 -2051
rect 1241 -2047 1242 -2045
rect 1241 -2053 1242 -2051
rect 1248 -2047 1249 -2045
rect 1248 -2053 1249 -2051
rect 1255 -2047 1256 -2045
rect 1255 -2053 1256 -2051
rect 1262 -2047 1263 -2045
rect 1265 -2047 1266 -2045
rect 1262 -2053 1263 -2051
rect 1265 -2053 1266 -2051
rect 1269 -2047 1270 -2045
rect 1269 -2053 1270 -2051
rect 1276 -2047 1277 -2045
rect 1276 -2053 1277 -2051
rect 1283 -2047 1284 -2045
rect 1283 -2053 1284 -2051
rect 1290 -2047 1291 -2045
rect 1293 -2047 1294 -2045
rect 1293 -2053 1294 -2051
rect 1297 -2047 1298 -2045
rect 1297 -2053 1298 -2051
rect 1304 -2047 1305 -2045
rect 1304 -2053 1305 -2051
rect 1311 -2047 1312 -2045
rect 1311 -2053 1312 -2051
rect 1318 -2047 1319 -2045
rect 1318 -2053 1319 -2051
rect 1325 -2047 1326 -2045
rect 1325 -2053 1326 -2051
rect 1332 -2047 1333 -2045
rect 1332 -2053 1333 -2051
rect 1339 -2047 1340 -2045
rect 1339 -2053 1340 -2051
rect 1346 -2047 1347 -2045
rect 1346 -2053 1347 -2051
rect 1353 -2047 1354 -2045
rect 1353 -2053 1354 -2051
rect 1360 -2047 1361 -2045
rect 1360 -2053 1361 -2051
rect 1367 -2047 1368 -2045
rect 1367 -2053 1368 -2051
rect 1374 -2047 1375 -2045
rect 1374 -2053 1375 -2051
rect 1381 -2047 1382 -2045
rect 1381 -2053 1382 -2051
rect 1388 -2047 1389 -2045
rect 1388 -2053 1389 -2051
rect 1395 -2047 1396 -2045
rect 1395 -2053 1396 -2051
rect 1402 -2047 1403 -2045
rect 1402 -2053 1403 -2051
rect 1409 -2047 1410 -2045
rect 1409 -2053 1410 -2051
rect 1416 -2047 1417 -2045
rect 1416 -2053 1417 -2051
rect 1423 -2047 1424 -2045
rect 1423 -2053 1424 -2051
rect 1430 -2047 1431 -2045
rect 1430 -2053 1431 -2051
rect 1437 -2047 1438 -2045
rect 1437 -2053 1438 -2051
rect 1444 -2047 1445 -2045
rect 1444 -2053 1445 -2051
rect 1451 -2047 1452 -2045
rect 1454 -2047 1455 -2045
rect 1451 -2053 1452 -2051
rect 1458 -2047 1459 -2045
rect 1458 -2053 1459 -2051
rect 1465 -2047 1466 -2045
rect 1465 -2053 1466 -2051
rect 1472 -2047 1473 -2045
rect 1472 -2053 1473 -2051
rect 1479 -2047 1480 -2045
rect 1479 -2053 1480 -2051
rect 1486 -2047 1487 -2045
rect 1486 -2053 1487 -2051
rect 1493 -2047 1494 -2045
rect 1493 -2053 1494 -2051
rect 1500 -2047 1501 -2045
rect 1500 -2053 1501 -2051
rect 1507 -2047 1508 -2045
rect 1507 -2053 1508 -2051
rect 1514 -2047 1515 -2045
rect 1514 -2053 1515 -2051
rect 1521 -2047 1522 -2045
rect 1521 -2053 1522 -2051
rect 1528 -2047 1529 -2045
rect 1528 -2053 1529 -2051
rect 1535 -2047 1536 -2045
rect 1535 -2053 1536 -2051
rect 1542 -2047 1543 -2045
rect 1542 -2053 1543 -2051
rect 1549 -2047 1550 -2045
rect 1549 -2053 1550 -2051
rect 1556 -2047 1557 -2045
rect 1556 -2053 1557 -2051
rect 1563 -2047 1564 -2045
rect 1563 -2053 1564 -2051
rect 1570 -2047 1571 -2045
rect 1570 -2053 1571 -2051
rect 1577 -2047 1578 -2045
rect 1577 -2053 1578 -2051
rect 1584 -2047 1585 -2045
rect 1584 -2053 1585 -2051
rect 1591 -2047 1592 -2045
rect 1591 -2053 1592 -2051
rect 1598 -2047 1599 -2045
rect 1598 -2053 1599 -2051
rect 1605 -2047 1606 -2045
rect 1605 -2053 1606 -2051
rect 1612 -2047 1613 -2045
rect 1612 -2053 1613 -2051
rect 1619 -2047 1620 -2045
rect 1619 -2053 1620 -2051
rect 1626 -2047 1627 -2045
rect 1626 -2053 1627 -2051
rect 1633 -2047 1634 -2045
rect 1633 -2053 1634 -2051
rect 1640 -2047 1641 -2045
rect 1640 -2053 1641 -2051
rect 1647 -2047 1648 -2045
rect 1647 -2053 1648 -2051
rect 1654 -2047 1655 -2045
rect 1654 -2053 1655 -2051
rect 1661 -2047 1662 -2045
rect 1661 -2053 1662 -2051
rect 1668 -2047 1669 -2045
rect 1668 -2053 1669 -2051
rect 1675 -2047 1676 -2045
rect 1675 -2053 1676 -2051
rect 1682 -2047 1683 -2045
rect 1682 -2053 1683 -2051
rect 1689 -2047 1690 -2045
rect 1689 -2053 1690 -2051
rect 1696 -2047 1697 -2045
rect 1696 -2053 1697 -2051
rect 1703 -2047 1704 -2045
rect 1703 -2053 1704 -2051
rect 1710 -2047 1711 -2045
rect 1710 -2053 1711 -2051
rect 1717 -2047 1718 -2045
rect 1717 -2053 1718 -2051
rect 1724 -2047 1725 -2045
rect 1724 -2053 1725 -2051
rect 1731 -2047 1732 -2045
rect 1731 -2053 1732 -2051
rect 1738 -2047 1739 -2045
rect 1738 -2053 1739 -2051
rect 1745 -2047 1746 -2045
rect 1745 -2053 1746 -2051
rect 1752 -2047 1753 -2045
rect 1752 -2053 1753 -2051
rect 1759 -2047 1760 -2045
rect 1759 -2053 1760 -2051
rect 1766 -2047 1767 -2045
rect 1766 -2053 1767 -2051
rect 1773 -2047 1774 -2045
rect 1773 -2053 1774 -2051
rect 1780 -2047 1781 -2045
rect 1780 -2053 1781 -2051
rect 1787 -2047 1788 -2045
rect 1787 -2053 1788 -2051
rect 1794 -2047 1795 -2045
rect 1794 -2053 1795 -2051
rect 1801 -2047 1802 -2045
rect 1801 -2053 1802 -2051
rect 1808 -2047 1809 -2045
rect 1808 -2053 1809 -2051
rect 1815 -2047 1816 -2045
rect 1815 -2053 1816 -2051
rect 1822 -2047 1823 -2045
rect 1822 -2053 1823 -2051
rect 1829 -2047 1830 -2045
rect 1829 -2053 1830 -2051
rect 1836 -2047 1837 -2045
rect 1836 -2053 1837 -2051
rect 1843 -2047 1844 -2045
rect 1843 -2053 1844 -2051
rect 1850 -2047 1851 -2045
rect 1850 -2053 1851 -2051
rect 1857 -2047 1858 -2045
rect 1857 -2053 1858 -2051
rect 1864 -2047 1865 -2045
rect 1864 -2053 1865 -2051
rect 1871 -2047 1872 -2045
rect 1871 -2053 1872 -2051
rect 1878 -2047 1879 -2045
rect 1878 -2053 1879 -2051
rect 1885 -2047 1886 -2045
rect 1885 -2053 1886 -2051
rect 1892 -2047 1893 -2045
rect 1892 -2053 1893 -2051
rect 1899 -2047 1900 -2045
rect 1899 -2053 1900 -2051
rect 1906 -2047 1907 -2045
rect 1906 -2053 1907 -2051
rect 1913 -2047 1914 -2045
rect 1913 -2053 1914 -2051
rect 1920 -2047 1921 -2045
rect 1920 -2053 1921 -2051
rect 1923 -2053 1924 -2051
rect 1927 -2047 1928 -2045
rect 1927 -2053 1928 -2051
rect 1934 -2047 1935 -2045
rect 1934 -2053 1935 -2051
rect 1941 -2047 1942 -2045
rect 1941 -2053 1942 -2051
rect 1948 -2047 1949 -2045
rect 1948 -2053 1949 -2051
rect 1955 -2047 1956 -2045
rect 1955 -2053 1956 -2051
rect 1962 -2047 1963 -2045
rect 1962 -2053 1963 -2051
rect 1969 -2047 1970 -2045
rect 1969 -2053 1970 -2051
rect 1976 -2047 1977 -2045
rect 1976 -2053 1977 -2051
rect 1983 -2047 1984 -2045
rect 1983 -2053 1984 -2051
rect 1990 -2047 1991 -2045
rect 1990 -2053 1991 -2051
rect 2 -2188 3 -2186
rect 2 -2194 3 -2192
rect 12 -2194 13 -2192
rect 16 -2188 17 -2186
rect 16 -2194 17 -2192
rect 23 -2188 24 -2186
rect 23 -2194 24 -2192
rect 30 -2188 31 -2186
rect 33 -2188 34 -2186
rect 30 -2194 31 -2192
rect 33 -2194 34 -2192
rect 40 -2188 41 -2186
rect 37 -2194 38 -2192
rect 40 -2194 41 -2192
rect 44 -2188 45 -2186
rect 44 -2194 45 -2192
rect 51 -2188 52 -2186
rect 51 -2194 52 -2192
rect 58 -2188 59 -2186
rect 58 -2194 59 -2192
rect 65 -2188 66 -2186
rect 65 -2194 66 -2192
rect 72 -2188 73 -2186
rect 72 -2194 73 -2192
rect 79 -2188 80 -2186
rect 79 -2194 80 -2192
rect 86 -2188 87 -2186
rect 89 -2188 90 -2186
rect 86 -2194 87 -2192
rect 89 -2194 90 -2192
rect 93 -2188 94 -2186
rect 96 -2188 97 -2186
rect 93 -2194 94 -2192
rect 100 -2188 101 -2186
rect 100 -2194 101 -2192
rect 110 -2188 111 -2186
rect 107 -2194 108 -2192
rect 110 -2194 111 -2192
rect 121 -2188 122 -2186
rect 121 -2194 122 -2192
rect 128 -2188 129 -2186
rect 128 -2194 129 -2192
rect 135 -2188 136 -2186
rect 135 -2194 136 -2192
rect 142 -2188 143 -2186
rect 142 -2194 143 -2192
rect 149 -2188 150 -2186
rect 149 -2194 150 -2192
rect 156 -2188 157 -2186
rect 156 -2194 157 -2192
rect 163 -2188 164 -2186
rect 163 -2194 164 -2192
rect 170 -2188 171 -2186
rect 170 -2194 171 -2192
rect 177 -2188 178 -2186
rect 177 -2194 178 -2192
rect 184 -2188 185 -2186
rect 184 -2194 185 -2192
rect 191 -2188 192 -2186
rect 191 -2194 192 -2192
rect 198 -2188 199 -2186
rect 198 -2194 199 -2192
rect 205 -2188 206 -2186
rect 205 -2194 206 -2192
rect 212 -2188 213 -2186
rect 212 -2194 213 -2192
rect 219 -2188 220 -2186
rect 219 -2194 220 -2192
rect 226 -2188 227 -2186
rect 226 -2194 227 -2192
rect 233 -2188 234 -2186
rect 236 -2188 237 -2186
rect 240 -2188 241 -2186
rect 240 -2194 241 -2192
rect 247 -2188 248 -2186
rect 247 -2194 248 -2192
rect 254 -2188 255 -2186
rect 254 -2194 255 -2192
rect 261 -2188 262 -2186
rect 261 -2194 262 -2192
rect 268 -2188 269 -2186
rect 268 -2194 269 -2192
rect 275 -2188 276 -2186
rect 275 -2194 276 -2192
rect 282 -2188 283 -2186
rect 282 -2194 283 -2192
rect 289 -2188 290 -2186
rect 289 -2194 290 -2192
rect 296 -2188 297 -2186
rect 296 -2194 297 -2192
rect 303 -2188 304 -2186
rect 303 -2194 304 -2192
rect 310 -2188 311 -2186
rect 310 -2194 311 -2192
rect 317 -2188 318 -2186
rect 317 -2194 318 -2192
rect 324 -2188 325 -2186
rect 324 -2194 325 -2192
rect 331 -2188 332 -2186
rect 331 -2194 332 -2192
rect 341 -2188 342 -2186
rect 341 -2194 342 -2192
rect 345 -2188 346 -2186
rect 345 -2194 346 -2192
rect 352 -2188 353 -2186
rect 352 -2194 353 -2192
rect 359 -2188 360 -2186
rect 359 -2194 360 -2192
rect 366 -2188 367 -2186
rect 366 -2194 367 -2192
rect 373 -2188 374 -2186
rect 373 -2194 374 -2192
rect 380 -2188 381 -2186
rect 380 -2194 381 -2192
rect 387 -2188 388 -2186
rect 390 -2188 391 -2186
rect 387 -2194 388 -2192
rect 390 -2194 391 -2192
rect 394 -2188 395 -2186
rect 394 -2194 395 -2192
rect 401 -2188 402 -2186
rect 404 -2188 405 -2186
rect 401 -2194 402 -2192
rect 408 -2188 409 -2186
rect 408 -2194 409 -2192
rect 415 -2188 416 -2186
rect 415 -2194 416 -2192
rect 422 -2188 423 -2186
rect 422 -2194 423 -2192
rect 429 -2188 430 -2186
rect 429 -2194 430 -2192
rect 436 -2188 437 -2186
rect 439 -2188 440 -2186
rect 436 -2194 437 -2192
rect 443 -2188 444 -2186
rect 443 -2194 444 -2192
rect 450 -2188 451 -2186
rect 450 -2194 451 -2192
rect 457 -2188 458 -2186
rect 457 -2194 458 -2192
rect 464 -2188 465 -2186
rect 467 -2188 468 -2186
rect 464 -2194 465 -2192
rect 471 -2188 472 -2186
rect 471 -2194 472 -2192
rect 478 -2188 479 -2186
rect 478 -2194 479 -2192
rect 485 -2188 486 -2186
rect 485 -2194 486 -2192
rect 492 -2188 493 -2186
rect 492 -2194 493 -2192
rect 499 -2188 500 -2186
rect 499 -2194 500 -2192
rect 506 -2188 507 -2186
rect 509 -2188 510 -2186
rect 506 -2194 507 -2192
rect 509 -2194 510 -2192
rect 513 -2188 514 -2186
rect 513 -2194 514 -2192
rect 520 -2188 521 -2186
rect 520 -2194 521 -2192
rect 527 -2188 528 -2186
rect 527 -2194 528 -2192
rect 534 -2188 535 -2186
rect 534 -2194 535 -2192
rect 541 -2194 542 -2192
rect 544 -2194 545 -2192
rect 548 -2188 549 -2186
rect 548 -2194 549 -2192
rect 555 -2188 556 -2186
rect 555 -2194 556 -2192
rect 562 -2188 563 -2186
rect 562 -2194 563 -2192
rect 569 -2188 570 -2186
rect 569 -2194 570 -2192
rect 576 -2188 577 -2186
rect 576 -2194 577 -2192
rect 583 -2188 584 -2186
rect 583 -2194 584 -2192
rect 590 -2188 591 -2186
rect 593 -2188 594 -2186
rect 590 -2194 591 -2192
rect 597 -2188 598 -2186
rect 597 -2194 598 -2192
rect 604 -2188 605 -2186
rect 604 -2194 605 -2192
rect 611 -2188 612 -2186
rect 611 -2194 612 -2192
rect 618 -2188 619 -2186
rect 618 -2194 619 -2192
rect 625 -2188 626 -2186
rect 628 -2188 629 -2186
rect 632 -2188 633 -2186
rect 632 -2194 633 -2192
rect 639 -2188 640 -2186
rect 639 -2194 640 -2192
rect 646 -2188 647 -2186
rect 649 -2188 650 -2186
rect 649 -2194 650 -2192
rect 653 -2188 654 -2186
rect 653 -2194 654 -2192
rect 660 -2188 661 -2186
rect 660 -2194 661 -2192
rect 667 -2188 668 -2186
rect 667 -2194 668 -2192
rect 674 -2188 675 -2186
rect 674 -2194 675 -2192
rect 681 -2188 682 -2186
rect 681 -2194 682 -2192
rect 688 -2188 689 -2186
rect 688 -2194 689 -2192
rect 695 -2188 696 -2186
rect 695 -2194 696 -2192
rect 702 -2188 703 -2186
rect 702 -2194 703 -2192
rect 709 -2188 710 -2186
rect 709 -2194 710 -2192
rect 716 -2188 717 -2186
rect 716 -2194 717 -2192
rect 723 -2188 724 -2186
rect 723 -2194 724 -2192
rect 730 -2188 731 -2186
rect 730 -2194 731 -2192
rect 737 -2188 738 -2186
rect 737 -2194 738 -2192
rect 744 -2188 745 -2186
rect 744 -2194 745 -2192
rect 751 -2188 752 -2186
rect 751 -2194 752 -2192
rect 758 -2188 759 -2186
rect 758 -2194 759 -2192
rect 765 -2188 766 -2186
rect 765 -2194 766 -2192
rect 772 -2188 773 -2186
rect 772 -2194 773 -2192
rect 779 -2188 780 -2186
rect 779 -2194 780 -2192
rect 786 -2188 787 -2186
rect 786 -2194 787 -2192
rect 793 -2188 794 -2186
rect 793 -2194 794 -2192
rect 800 -2188 801 -2186
rect 800 -2194 801 -2192
rect 807 -2188 808 -2186
rect 807 -2194 808 -2192
rect 814 -2188 815 -2186
rect 814 -2194 815 -2192
rect 821 -2188 822 -2186
rect 821 -2194 822 -2192
rect 828 -2188 829 -2186
rect 828 -2194 829 -2192
rect 835 -2188 836 -2186
rect 838 -2188 839 -2186
rect 835 -2194 836 -2192
rect 842 -2188 843 -2186
rect 842 -2194 843 -2192
rect 849 -2188 850 -2186
rect 849 -2194 850 -2192
rect 856 -2188 857 -2186
rect 856 -2194 857 -2192
rect 863 -2188 864 -2186
rect 863 -2194 864 -2192
rect 870 -2188 871 -2186
rect 870 -2194 871 -2192
rect 877 -2188 878 -2186
rect 880 -2188 881 -2186
rect 877 -2194 878 -2192
rect 880 -2194 881 -2192
rect 884 -2188 885 -2186
rect 884 -2194 885 -2192
rect 891 -2188 892 -2186
rect 891 -2194 892 -2192
rect 898 -2188 899 -2186
rect 898 -2194 899 -2192
rect 905 -2188 906 -2186
rect 905 -2194 906 -2192
rect 912 -2188 913 -2186
rect 912 -2194 913 -2192
rect 919 -2188 920 -2186
rect 919 -2194 920 -2192
rect 926 -2188 927 -2186
rect 926 -2194 927 -2192
rect 933 -2188 934 -2186
rect 933 -2194 934 -2192
rect 940 -2188 941 -2186
rect 940 -2194 941 -2192
rect 947 -2188 948 -2186
rect 947 -2194 948 -2192
rect 954 -2188 955 -2186
rect 954 -2194 955 -2192
rect 961 -2188 962 -2186
rect 961 -2194 962 -2192
rect 968 -2188 969 -2186
rect 971 -2188 972 -2186
rect 968 -2194 969 -2192
rect 971 -2194 972 -2192
rect 975 -2188 976 -2186
rect 978 -2188 979 -2186
rect 975 -2194 976 -2192
rect 978 -2194 979 -2192
rect 982 -2188 983 -2186
rect 982 -2194 983 -2192
rect 989 -2188 990 -2186
rect 989 -2194 990 -2192
rect 996 -2188 997 -2186
rect 996 -2194 997 -2192
rect 1003 -2188 1004 -2186
rect 1003 -2194 1004 -2192
rect 1010 -2188 1011 -2186
rect 1010 -2194 1011 -2192
rect 1017 -2188 1018 -2186
rect 1017 -2194 1018 -2192
rect 1024 -2188 1025 -2186
rect 1024 -2194 1025 -2192
rect 1031 -2188 1032 -2186
rect 1031 -2194 1032 -2192
rect 1038 -2188 1039 -2186
rect 1038 -2194 1039 -2192
rect 1045 -2188 1046 -2186
rect 1045 -2194 1046 -2192
rect 1052 -2188 1053 -2186
rect 1052 -2194 1053 -2192
rect 1055 -2194 1056 -2192
rect 1059 -2188 1060 -2186
rect 1059 -2194 1060 -2192
rect 1066 -2188 1067 -2186
rect 1069 -2188 1070 -2186
rect 1066 -2194 1067 -2192
rect 1069 -2194 1070 -2192
rect 1073 -2188 1074 -2186
rect 1073 -2194 1074 -2192
rect 1080 -2188 1081 -2186
rect 1083 -2188 1084 -2186
rect 1083 -2194 1084 -2192
rect 1087 -2188 1088 -2186
rect 1087 -2194 1088 -2192
rect 1094 -2188 1095 -2186
rect 1094 -2194 1095 -2192
rect 1101 -2188 1102 -2186
rect 1101 -2194 1102 -2192
rect 1108 -2188 1109 -2186
rect 1111 -2188 1112 -2186
rect 1108 -2194 1109 -2192
rect 1111 -2194 1112 -2192
rect 1115 -2188 1116 -2186
rect 1115 -2194 1116 -2192
rect 1122 -2188 1123 -2186
rect 1122 -2194 1123 -2192
rect 1129 -2188 1130 -2186
rect 1129 -2194 1130 -2192
rect 1139 -2188 1140 -2186
rect 1139 -2194 1140 -2192
rect 1143 -2188 1144 -2186
rect 1143 -2194 1144 -2192
rect 1150 -2188 1151 -2186
rect 1150 -2194 1151 -2192
rect 1157 -2188 1158 -2186
rect 1160 -2188 1161 -2186
rect 1157 -2194 1158 -2192
rect 1160 -2194 1161 -2192
rect 1164 -2188 1165 -2186
rect 1164 -2194 1165 -2192
rect 1171 -2188 1172 -2186
rect 1171 -2194 1172 -2192
rect 1178 -2188 1179 -2186
rect 1178 -2194 1179 -2192
rect 1185 -2188 1186 -2186
rect 1185 -2194 1186 -2192
rect 1192 -2188 1193 -2186
rect 1192 -2194 1193 -2192
rect 1199 -2188 1200 -2186
rect 1199 -2194 1200 -2192
rect 1206 -2188 1207 -2186
rect 1206 -2194 1207 -2192
rect 1213 -2188 1214 -2186
rect 1213 -2194 1214 -2192
rect 1220 -2188 1221 -2186
rect 1220 -2194 1221 -2192
rect 1227 -2188 1228 -2186
rect 1227 -2194 1228 -2192
rect 1234 -2188 1235 -2186
rect 1234 -2194 1235 -2192
rect 1241 -2188 1242 -2186
rect 1241 -2194 1242 -2192
rect 1248 -2188 1249 -2186
rect 1248 -2194 1249 -2192
rect 1255 -2188 1256 -2186
rect 1255 -2194 1256 -2192
rect 1262 -2188 1263 -2186
rect 1262 -2194 1263 -2192
rect 1269 -2188 1270 -2186
rect 1269 -2194 1270 -2192
rect 1276 -2188 1277 -2186
rect 1276 -2194 1277 -2192
rect 1279 -2194 1280 -2192
rect 1283 -2188 1284 -2186
rect 1283 -2194 1284 -2192
rect 1290 -2188 1291 -2186
rect 1290 -2194 1291 -2192
rect 1297 -2188 1298 -2186
rect 1297 -2194 1298 -2192
rect 1304 -2188 1305 -2186
rect 1304 -2194 1305 -2192
rect 1311 -2188 1312 -2186
rect 1311 -2194 1312 -2192
rect 1318 -2188 1319 -2186
rect 1318 -2194 1319 -2192
rect 1325 -2188 1326 -2186
rect 1325 -2194 1326 -2192
rect 1332 -2188 1333 -2186
rect 1332 -2194 1333 -2192
rect 1339 -2188 1340 -2186
rect 1339 -2194 1340 -2192
rect 1346 -2188 1347 -2186
rect 1346 -2194 1347 -2192
rect 1353 -2188 1354 -2186
rect 1353 -2194 1354 -2192
rect 1360 -2188 1361 -2186
rect 1363 -2188 1364 -2186
rect 1360 -2194 1361 -2192
rect 1367 -2188 1368 -2186
rect 1367 -2194 1368 -2192
rect 1374 -2188 1375 -2186
rect 1377 -2188 1378 -2186
rect 1374 -2194 1375 -2192
rect 1381 -2188 1382 -2186
rect 1381 -2194 1382 -2192
rect 1388 -2188 1389 -2186
rect 1388 -2194 1389 -2192
rect 1395 -2188 1396 -2186
rect 1398 -2188 1399 -2186
rect 1395 -2194 1396 -2192
rect 1398 -2194 1399 -2192
rect 1402 -2188 1403 -2186
rect 1402 -2194 1403 -2192
rect 1409 -2188 1410 -2186
rect 1409 -2194 1410 -2192
rect 1416 -2188 1417 -2186
rect 1416 -2194 1417 -2192
rect 1423 -2188 1424 -2186
rect 1423 -2194 1424 -2192
rect 1430 -2188 1431 -2186
rect 1430 -2194 1431 -2192
rect 1437 -2188 1438 -2186
rect 1437 -2194 1438 -2192
rect 1444 -2188 1445 -2186
rect 1444 -2194 1445 -2192
rect 1451 -2188 1452 -2186
rect 1454 -2188 1455 -2186
rect 1454 -2194 1455 -2192
rect 1458 -2188 1459 -2186
rect 1458 -2194 1459 -2192
rect 1465 -2188 1466 -2186
rect 1465 -2194 1466 -2192
rect 1475 -2188 1476 -2186
rect 1472 -2194 1473 -2192
rect 1475 -2194 1476 -2192
rect 1479 -2188 1480 -2186
rect 1479 -2194 1480 -2192
rect 1486 -2188 1487 -2186
rect 1486 -2194 1487 -2192
rect 1493 -2188 1494 -2186
rect 1493 -2194 1494 -2192
rect 1500 -2188 1501 -2186
rect 1500 -2194 1501 -2192
rect 1507 -2188 1508 -2186
rect 1507 -2194 1508 -2192
rect 1514 -2188 1515 -2186
rect 1514 -2194 1515 -2192
rect 1521 -2188 1522 -2186
rect 1521 -2194 1522 -2192
rect 1528 -2188 1529 -2186
rect 1528 -2194 1529 -2192
rect 1535 -2188 1536 -2186
rect 1535 -2194 1536 -2192
rect 1542 -2188 1543 -2186
rect 1542 -2194 1543 -2192
rect 1549 -2188 1550 -2186
rect 1549 -2194 1550 -2192
rect 1556 -2188 1557 -2186
rect 1556 -2194 1557 -2192
rect 1563 -2188 1564 -2186
rect 1563 -2194 1564 -2192
rect 1570 -2188 1571 -2186
rect 1570 -2194 1571 -2192
rect 1577 -2188 1578 -2186
rect 1577 -2194 1578 -2192
rect 1584 -2188 1585 -2186
rect 1584 -2194 1585 -2192
rect 1591 -2188 1592 -2186
rect 1591 -2194 1592 -2192
rect 1598 -2188 1599 -2186
rect 1598 -2194 1599 -2192
rect 1605 -2188 1606 -2186
rect 1605 -2194 1606 -2192
rect 1612 -2188 1613 -2186
rect 1612 -2194 1613 -2192
rect 1619 -2188 1620 -2186
rect 1619 -2194 1620 -2192
rect 1626 -2188 1627 -2186
rect 1626 -2194 1627 -2192
rect 1633 -2188 1634 -2186
rect 1633 -2194 1634 -2192
rect 1640 -2188 1641 -2186
rect 1640 -2194 1641 -2192
rect 1647 -2188 1648 -2186
rect 1647 -2194 1648 -2192
rect 1654 -2188 1655 -2186
rect 1654 -2194 1655 -2192
rect 1661 -2188 1662 -2186
rect 1661 -2194 1662 -2192
rect 1668 -2188 1669 -2186
rect 1668 -2194 1669 -2192
rect 1675 -2188 1676 -2186
rect 1675 -2194 1676 -2192
rect 1682 -2188 1683 -2186
rect 1682 -2194 1683 -2192
rect 1689 -2188 1690 -2186
rect 1689 -2194 1690 -2192
rect 1696 -2188 1697 -2186
rect 1696 -2194 1697 -2192
rect 1703 -2188 1704 -2186
rect 1703 -2194 1704 -2192
rect 1710 -2188 1711 -2186
rect 1710 -2194 1711 -2192
rect 1717 -2188 1718 -2186
rect 1717 -2194 1718 -2192
rect 1724 -2188 1725 -2186
rect 1724 -2194 1725 -2192
rect 1731 -2188 1732 -2186
rect 1731 -2194 1732 -2192
rect 1738 -2188 1739 -2186
rect 1738 -2194 1739 -2192
rect 1745 -2188 1746 -2186
rect 1745 -2194 1746 -2192
rect 1752 -2188 1753 -2186
rect 1752 -2194 1753 -2192
rect 1759 -2188 1760 -2186
rect 1759 -2194 1760 -2192
rect 1766 -2188 1767 -2186
rect 1766 -2194 1767 -2192
rect 1773 -2188 1774 -2186
rect 1773 -2194 1774 -2192
rect 1780 -2188 1781 -2186
rect 1780 -2194 1781 -2192
rect 1787 -2188 1788 -2186
rect 1787 -2194 1788 -2192
rect 1794 -2188 1795 -2186
rect 1794 -2194 1795 -2192
rect 1801 -2188 1802 -2186
rect 1801 -2194 1802 -2192
rect 1808 -2188 1809 -2186
rect 1808 -2194 1809 -2192
rect 1815 -2188 1816 -2186
rect 1815 -2194 1816 -2192
rect 1822 -2188 1823 -2186
rect 1822 -2194 1823 -2192
rect 1829 -2188 1830 -2186
rect 1829 -2194 1830 -2192
rect 1836 -2188 1837 -2186
rect 1836 -2194 1837 -2192
rect 1843 -2188 1844 -2186
rect 1843 -2194 1844 -2192
rect 1850 -2188 1851 -2186
rect 1850 -2194 1851 -2192
rect 1857 -2188 1858 -2186
rect 1857 -2194 1858 -2192
rect 1864 -2188 1865 -2186
rect 1864 -2194 1865 -2192
rect 1871 -2188 1872 -2186
rect 1871 -2194 1872 -2192
rect 1878 -2188 1879 -2186
rect 1878 -2194 1879 -2192
rect 1885 -2188 1886 -2186
rect 1885 -2194 1886 -2192
rect 1892 -2188 1893 -2186
rect 1892 -2194 1893 -2192
rect 1899 -2188 1900 -2186
rect 1899 -2194 1900 -2192
rect 1906 -2188 1907 -2186
rect 1906 -2194 1907 -2192
rect 1913 -2188 1914 -2186
rect 1913 -2194 1914 -2192
rect 9 -2317 10 -2315
rect 9 -2323 10 -2321
rect 16 -2317 17 -2315
rect 16 -2323 17 -2321
rect 23 -2317 24 -2315
rect 23 -2323 24 -2321
rect 30 -2317 31 -2315
rect 30 -2323 31 -2321
rect 37 -2317 38 -2315
rect 37 -2323 38 -2321
rect 44 -2317 45 -2315
rect 44 -2323 45 -2321
rect 51 -2317 52 -2315
rect 51 -2323 52 -2321
rect 58 -2317 59 -2315
rect 58 -2323 59 -2321
rect 65 -2317 66 -2315
rect 68 -2317 69 -2315
rect 72 -2317 73 -2315
rect 72 -2323 73 -2321
rect 79 -2317 80 -2315
rect 79 -2323 80 -2321
rect 86 -2317 87 -2315
rect 86 -2323 87 -2321
rect 93 -2317 94 -2315
rect 93 -2323 94 -2321
rect 100 -2317 101 -2315
rect 100 -2323 101 -2321
rect 107 -2317 108 -2315
rect 107 -2323 108 -2321
rect 117 -2317 118 -2315
rect 114 -2323 115 -2321
rect 117 -2323 118 -2321
rect 121 -2317 122 -2315
rect 124 -2317 125 -2315
rect 124 -2323 125 -2321
rect 128 -2317 129 -2315
rect 128 -2323 129 -2321
rect 135 -2317 136 -2315
rect 135 -2323 136 -2321
rect 142 -2317 143 -2315
rect 142 -2323 143 -2321
rect 149 -2317 150 -2315
rect 149 -2323 150 -2321
rect 156 -2317 157 -2315
rect 159 -2317 160 -2315
rect 156 -2323 157 -2321
rect 159 -2323 160 -2321
rect 163 -2317 164 -2315
rect 163 -2323 164 -2321
rect 170 -2317 171 -2315
rect 173 -2317 174 -2315
rect 170 -2323 171 -2321
rect 177 -2317 178 -2315
rect 177 -2323 178 -2321
rect 184 -2317 185 -2315
rect 184 -2323 185 -2321
rect 191 -2317 192 -2315
rect 191 -2323 192 -2321
rect 198 -2317 199 -2315
rect 198 -2323 199 -2321
rect 205 -2317 206 -2315
rect 208 -2317 209 -2315
rect 205 -2323 206 -2321
rect 212 -2317 213 -2315
rect 215 -2317 216 -2315
rect 212 -2323 213 -2321
rect 215 -2323 216 -2321
rect 219 -2317 220 -2315
rect 222 -2317 223 -2315
rect 219 -2323 220 -2321
rect 226 -2317 227 -2315
rect 226 -2323 227 -2321
rect 236 -2317 237 -2315
rect 236 -2323 237 -2321
rect 240 -2317 241 -2315
rect 240 -2323 241 -2321
rect 243 -2323 244 -2321
rect 247 -2317 248 -2315
rect 247 -2323 248 -2321
rect 254 -2317 255 -2315
rect 254 -2323 255 -2321
rect 261 -2317 262 -2315
rect 261 -2323 262 -2321
rect 268 -2317 269 -2315
rect 268 -2323 269 -2321
rect 275 -2317 276 -2315
rect 275 -2323 276 -2321
rect 282 -2317 283 -2315
rect 282 -2323 283 -2321
rect 289 -2317 290 -2315
rect 289 -2323 290 -2321
rect 296 -2317 297 -2315
rect 296 -2323 297 -2321
rect 303 -2317 304 -2315
rect 303 -2323 304 -2321
rect 310 -2317 311 -2315
rect 310 -2323 311 -2321
rect 317 -2317 318 -2315
rect 317 -2323 318 -2321
rect 324 -2317 325 -2315
rect 324 -2323 325 -2321
rect 331 -2317 332 -2315
rect 331 -2323 332 -2321
rect 338 -2317 339 -2315
rect 338 -2323 339 -2321
rect 345 -2317 346 -2315
rect 345 -2323 346 -2321
rect 352 -2317 353 -2315
rect 352 -2323 353 -2321
rect 359 -2317 360 -2315
rect 359 -2323 360 -2321
rect 366 -2317 367 -2315
rect 366 -2323 367 -2321
rect 373 -2317 374 -2315
rect 373 -2323 374 -2321
rect 380 -2317 381 -2315
rect 380 -2323 381 -2321
rect 387 -2317 388 -2315
rect 387 -2323 388 -2321
rect 394 -2317 395 -2315
rect 394 -2323 395 -2321
rect 401 -2317 402 -2315
rect 401 -2323 402 -2321
rect 408 -2317 409 -2315
rect 408 -2323 409 -2321
rect 415 -2317 416 -2315
rect 415 -2323 416 -2321
rect 422 -2317 423 -2315
rect 422 -2323 423 -2321
rect 429 -2317 430 -2315
rect 429 -2323 430 -2321
rect 436 -2317 437 -2315
rect 436 -2323 437 -2321
rect 443 -2317 444 -2315
rect 443 -2323 444 -2321
rect 450 -2317 451 -2315
rect 450 -2323 451 -2321
rect 457 -2317 458 -2315
rect 457 -2323 458 -2321
rect 467 -2317 468 -2315
rect 464 -2323 465 -2321
rect 467 -2323 468 -2321
rect 471 -2317 472 -2315
rect 471 -2323 472 -2321
rect 478 -2317 479 -2315
rect 478 -2323 479 -2321
rect 485 -2317 486 -2315
rect 485 -2323 486 -2321
rect 492 -2317 493 -2315
rect 492 -2323 493 -2321
rect 499 -2317 500 -2315
rect 499 -2323 500 -2321
rect 506 -2317 507 -2315
rect 506 -2323 507 -2321
rect 513 -2317 514 -2315
rect 513 -2323 514 -2321
rect 520 -2317 521 -2315
rect 520 -2323 521 -2321
rect 527 -2317 528 -2315
rect 527 -2323 528 -2321
rect 534 -2317 535 -2315
rect 534 -2323 535 -2321
rect 541 -2317 542 -2315
rect 541 -2323 542 -2321
rect 548 -2317 549 -2315
rect 548 -2323 549 -2321
rect 555 -2317 556 -2315
rect 555 -2323 556 -2321
rect 562 -2317 563 -2315
rect 562 -2323 563 -2321
rect 569 -2317 570 -2315
rect 572 -2317 573 -2315
rect 569 -2323 570 -2321
rect 572 -2323 573 -2321
rect 576 -2317 577 -2315
rect 576 -2323 577 -2321
rect 583 -2317 584 -2315
rect 583 -2323 584 -2321
rect 590 -2317 591 -2315
rect 590 -2323 591 -2321
rect 597 -2317 598 -2315
rect 597 -2323 598 -2321
rect 604 -2317 605 -2315
rect 604 -2323 605 -2321
rect 611 -2317 612 -2315
rect 611 -2323 612 -2321
rect 618 -2317 619 -2315
rect 618 -2323 619 -2321
rect 625 -2317 626 -2315
rect 628 -2317 629 -2315
rect 625 -2323 626 -2321
rect 632 -2317 633 -2315
rect 632 -2323 633 -2321
rect 639 -2317 640 -2315
rect 639 -2323 640 -2321
rect 646 -2317 647 -2315
rect 646 -2323 647 -2321
rect 653 -2317 654 -2315
rect 656 -2317 657 -2315
rect 656 -2323 657 -2321
rect 660 -2317 661 -2315
rect 660 -2323 661 -2321
rect 670 -2317 671 -2315
rect 667 -2323 668 -2321
rect 674 -2317 675 -2315
rect 677 -2317 678 -2315
rect 674 -2323 675 -2321
rect 677 -2323 678 -2321
rect 681 -2317 682 -2315
rect 681 -2323 682 -2321
rect 688 -2317 689 -2315
rect 688 -2323 689 -2321
rect 695 -2317 696 -2315
rect 695 -2323 696 -2321
rect 702 -2317 703 -2315
rect 702 -2323 703 -2321
rect 709 -2317 710 -2315
rect 709 -2323 710 -2321
rect 716 -2317 717 -2315
rect 716 -2323 717 -2321
rect 723 -2317 724 -2315
rect 723 -2323 724 -2321
rect 730 -2317 731 -2315
rect 730 -2323 731 -2321
rect 737 -2317 738 -2315
rect 737 -2323 738 -2321
rect 744 -2317 745 -2315
rect 744 -2323 745 -2321
rect 751 -2317 752 -2315
rect 751 -2323 752 -2321
rect 758 -2317 759 -2315
rect 761 -2317 762 -2315
rect 758 -2323 759 -2321
rect 765 -2317 766 -2315
rect 765 -2323 766 -2321
rect 772 -2317 773 -2315
rect 772 -2323 773 -2321
rect 779 -2317 780 -2315
rect 779 -2323 780 -2321
rect 786 -2317 787 -2315
rect 786 -2323 787 -2321
rect 793 -2317 794 -2315
rect 796 -2317 797 -2315
rect 796 -2323 797 -2321
rect 800 -2317 801 -2315
rect 800 -2323 801 -2321
rect 807 -2317 808 -2315
rect 807 -2323 808 -2321
rect 817 -2317 818 -2315
rect 817 -2323 818 -2321
rect 821 -2317 822 -2315
rect 824 -2317 825 -2315
rect 821 -2323 822 -2321
rect 824 -2323 825 -2321
rect 828 -2317 829 -2315
rect 828 -2323 829 -2321
rect 835 -2317 836 -2315
rect 835 -2323 836 -2321
rect 842 -2317 843 -2315
rect 842 -2323 843 -2321
rect 849 -2317 850 -2315
rect 849 -2323 850 -2321
rect 856 -2317 857 -2315
rect 856 -2323 857 -2321
rect 863 -2317 864 -2315
rect 863 -2323 864 -2321
rect 870 -2317 871 -2315
rect 870 -2323 871 -2321
rect 877 -2317 878 -2315
rect 877 -2323 878 -2321
rect 887 -2317 888 -2315
rect 884 -2323 885 -2321
rect 887 -2323 888 -2321
rect 891 -2317 892 -2315
rect 891 -2323 892 -2321
rect 898 -2317 899 -2315
rect 898 -2323 899 -2321
rect 905 -2317 906 -2315
rect 905 -2323 906 -2321
rect 912 -2317 913 -2315
rect 912 -2323 913 -2321
rect 919 -2317 920 -2315
rect 919 -2323 920 -2321
rect 926 -2317 927 -2315
rect 926 -2323 927 -2321
rect 933 -2317 934 -2315
rect 933 -2323 934 -2321
rect 940 -2317 941 -2315
rect 940 -2323 941 -2321
rect 947 -2317 948 -2315
rect 950 -2317 951 -2315
rect 947 -2323 948 -2321
rect 950 -2323 951 -2321
rect 954 -2317 955 -2315
rect 954 -2323 955 -2321
rect 961 -2317 962 -2315
rect 961 -2323 962 -2321
rect 968 -2317 969 -2315
rect 968 -2323 969 -2321
rect 975 -2317 976 -2315
rect 975 -2323 976 -2321
rect 982 -2317 983 -2315
rect 982 -2323 983 -2321
rect 989 -2317 990 -2315
rect 989 -2323 990 -2321
rect 996 -2317 997 -2315
rect 999 -2317 1000 -2315
rect 996 -2323 997 -2321
rect 999 -2323 1000 -2321
rect 1003 -2317 1004 -2315
rect 1003 -2323 1004 -2321
rect 1010 -2317 1011 -2315
rect 1010 -2323 1011 -2321
rect 1017 -2317 1018 -2315
rect 1017 -2323 1018 -2321
rect 1024 -2317 1025 -2315
rect 1024 -2323 1025 -2321
rect 1031 -2317 1032 -2315
rect 1031 -2323 1032 -2321
rect 1038 -2317 1039 -2315
rect 1038 -2323 1039 -2321
rect 1045 -2317 1046 -2315
rect 1045 -2323 1046 -2321
rect 1052 -2317 1053 -2315
rect 1052 -2323 1053 -2321
rect 1059 -2317 1060 -2315
rect 1059 -2323 1060 -2321
rect 1069 -2317 1070 -2315
rect 1066 -2323 1067 -2321
rect 1069 -2323 1070 -2321
rect 1073 -2317 1074 -2315
rect 1073 -2323 1074 -2321
rect 1080 -2317 1081 -2315
rect 1080 -2323 1081 -2321
rect 1087 -2317 1088 -2315
rect 1087 -2323 1088 -2321
rect 1094 -2317 1095 -2315
rect 1094 -2323 1095 -2321
rect 1101 -2317 1102 -2315
rect 1101 -2323 1102 -2321
rect 1108 -2317 1109 -2315
rect 1108 -2323 1109 -2321
rect 1115 -2317 1116 -2315
rect 1115 -2323 1116 -2321
rect 1118 -2323 1119 -2321
rect 1122 -2317 1123 -2315
rect 1125 -2317 1126 -2315
rect 1122 -2323 1123 -2321
rect 1129 -2317 1130 -2315
rect 1129 -2323 1130 -2321
rect 1136 -2317 1137 -2315
rect 1136 -2323 1137 -2321
rect 1143 -2317 1144 -2315
rect 1143 -2323 1144 -2321
rect 1150 -2317 1151 -2315
rect 1150 -2323 1151 -2321
rect 1157 -2317 1158 -2315
rect 1157 -2323 1158 -2321
rect 1164 -2317 1165 -2315
rect 1164 -2323 1165 -2321
rect 1171 -2317 1172 -2315
rect 1171 -2323 1172 -2321
rect 1178 -2317 1179 -2315
rect 1178 -2323 1179 -2321
rect 1185 -2317 1186 -2315
rect 1188 -2317 1189 -2315
rect 1185 -2323 1186 -2321
rect 1188 -2323 1189 -2321
rect 1192 -2317 1193 -2315
rect 1192 -2323 1193 -2321
rect 1199 -2317 1200 -2315
rect 1199 -2323 1200 -2321
rect 1206 -2317 1207 -2315
rect 1206 -2323 1207 -2321
rect 1213 -2317 1214 -2315
rect 1213 -2323 1214 -2321
rect 1220 -2317 1221 -2315
rect 1220 -2323 1221 -2321
rect 1227 -2317 1228 -2315
rect 1227 -2323 1228 -2321
rect 1234 -2317 1235 -2315
rect 1234 -2323 1235 -2321
rect 1241 -2317 1242 -2315
rect 1241 -2323 1242 -2321
rect 1248 -2317 1249 -2315
rect 1248 -2323 1249 -2321
rect 1255 -2317 1256 -2315
rect 1255 -2323 1256 -2321
rect 1262 -2317 1263 -2315
rect 1262 -2323 1263 -2321
rect 1269 -2317 1270 -2315
rect 1269 -2323 1270 -2321
rect 1276 -2317 1277 -2315
rect 1276 -2323 1277 -2321
rect 1283 -2317 1284 -2315
rect 1283 -2323 1284 -2321
rect 1290 -2317 1291 -2315
rect 1293 -2317 1294 -2315
rect 1290 -2323 1291 -2321
rect 1293 -2323 1294 -2321
rect 1297 -2317 1298 -2315
rect 1297 -2323 1298 -2321
rect 1304 -2317 1305 -2315
rect 1304 -2323 1305 -2321
rect 1307 -2323 1308 -2321
rect 1311 -2317 1312 -2315
rect 1311 -2323 1312 -2321
rect 1318 -2317 1319 -2315
rect 1318 -2323 1319 -2321
rect 1325 -2317 1326 -2315
rect 1325 -2323 1326 -2321
rect 1332 -2317 1333 -2315
rect 1332 -2323 1333 -2321
rect 1339 -2317 1340 -2315
rect 1339 -2323 1340 -2321
rect 1346 -2317 1347 -2315
rect 1346 -2323 1347 -2321
rect 1353 -2317 1354 -2315
rect 1353 -2323 1354 -2321
rect 1360 -2317 1361 -2315
rect 1360 -2323 1361 -2321
rect 1367 -2317 1368 -2315
rect 1367 -2323 1368 -2321
rect 1370 -2323 1371 -2321
rect 1374 -2317 1375 -2315
rect 1374 -2323 1375 -2321
rect 1381 -2317 1382 -2315
rect 1381 -2323 1382 -2321
rect 1388 -2317 1389 -2315
rect 1388 -2323 1389 -2321
rect 1395 -2317 1396 -2315
rect 1395 -2323 1396 -2321
rect 1402 -2317 1403 -2315
rect 1402 -2323 1403 -2321
rect 1409 -2317 1410 -2315
rect 1409 -2323 1410 -2321
rect 1416 -2317 1417 -2315
rect 1416 -2323 1417 -2321
rect 1423 -2317 1424 -2315
rect 1423 -2323 1424 -2321
rect 1430 -2317 1431 -2315
rect 1430 -2323 1431 -2321
rect 1437 -2317 1438 -2315
rect 1437 -2323 1438 -2321
rect 1444 -2317 1445 -2315
rect 1444 -2323 1445 -2321
rect 1451 -2317 1452 -2315
rect 1451 -2323 1452 -2321
rect 1458 -2317 1459 -2315
rect 1458 -2323 1459 -2321
rect 1465 -2317 1466 -2315
rect 1465 -2323 1466 -2321
rect 1472 -2317 1473 -2315
rect 1472 -2323 1473 -2321
rect 1479 -2317 1480 -2315
rect 1479 -2323 1480 -2321
rect 1486 -2317 1487 -2315
rect 1486 -2323 1487 -2321
rect 1493 -2317 1494 -2315
rect 1493 -2323 1494 -2321
rect 1500 -2317 1501 -2315
rect 1500 -2323 1501 -2321
rect 1507 -2317 1508 -2315
rect 1507 -2323 1508 -2321
rect 1514 -2317 1515 -2315
rect 1514 -2323 1515 -2321
rect 1521 -2317 1522 -2315
rect 1521 -2323 1522 -2321
rect 1528 -2317 1529 -2315
rect 1528 -2323 1529 -2321
rect 1535 -2317 1536 -2315
rect 1535 -2323 1536 -2321
rect 1542 -2317 1543 -2315
rect 1542 -2323 1543 -2321
rect 1549 -2317 1550 -2315
rect 1549 -2323 1550 -2321
rect 1556 -2317 1557 -2315
rect 1556 -2323 1557 -2321
rect 1563 -2317 1564 -2315
rect 1563 -2323 1564 -2321
rect 1570 -2317 1571 -2315
rect 1570 -2323 1571 -2321
rect 1577 -2317 1578 -2315
rect 1577 -2323 1578 -2321
rect 1584 -2317 1585 -2315
rect 1584 -2323 1585 -2321
rect 1591 -2317 1592 -2315
rect 1591 -2323 1592 -2321
rect 1598 -2317 1599 -2315
rect 1598 -2323 1599 -2321
rect 1605 -2317 1606 -2315
rect 1605 -2323 1606 -2321
rect 1612 -2317 1613 -2315
rect 1612 -2323 1613 -2321
rect 1619 -2317 1620 -2315
rect 1619 -2323 1620 -2321
rect 1626 -2317 1627 -2315
rect 1626 -2323 1627 -2321
rect 1633 -2317 1634 -2315
rect 1633 -2323 1634 -2321
rect 1640 -2317 1641 -2315
rect 1640 -2323 1641 -2321
rect 1647 -2317 1648 -2315
rect 1647 -2323 1648 -2321
rect 1654 -2317 1655 -2315
rect 1654 -2323 1655 -2321
rect 1661 -2317 1662 -2315
rect 1661 -2323 1662 -2321
rect 1668 -2317 1669 -2315
rect 1668 -2323 1669 -2321
rect 1675 -2317 1676 -2315
rect 1675 -2323 1676 -2321
rect 1682 -2317 1683 -2315
rect 1682 -2323 1683 -2321
rect 1689 -2317 1690 -2315
rect 1689 -2323 1690 -2321
rect 1696 -2317 1697 -2315
rect 1696 -2323 1697 -2321
rect 1703 -2317 1704 -2315
rect 1703 -2323 1704 -2321
rect 1710 -2317 1711 -2315
rect 1713 -2317 1714 -2315
rect 1713 -2323 1714 -2321
rect 1717 -2317 1718 -2315
rect 1717 -2323 1718 -2321
rect 1727 -2317 1728 -2315
rect 1727 -2323 1728 -2321
rect 1731 -2317 1732 -2315
rect 1731 -2323 1732 -2321
rect 1738 -2317 1739 -2315
rect 1738 -2323 1739 -2321
rect 1745 -2317 1746 -2315
rect 1748 -2323 1749 -2321
rect 1752 -2317 1753 -2315
rect 1752 -2323 1753 -2321
rect 1759 -2317 1760 -2315
rect 1759 -2323 1760 -2321
rect 1766 -2317 1767 -2315
rect 1766 -2323 1767 -2321
rect 1773 -2317 1774 -2315
rect 1773 -2323 1774 -2321
rect 1780 -2317 1781 -2315
rect 1780 -2323 1781 -2321
rect 1787 -2317 1788 -2315
rect 1787 -2323 1788 -2321
rect 1794 -2317 1795 -2315
rect 1794 -2323 1795 -2321
rect 1822 -2317 1823 -2315
rect 1822 -2323 1823 -2321
rect 1829 -2317 1830 -2315
rect 1829 -2323 1830 -2321
rect 9 -2442 10 -2440
rect 9 -2448 10 -2446
rect 16 -2442 17 -2440
rect 16 -2448 17 -2446
rect 30 -2442 31 -2440
rect 30 -2448 31 -2446
rect 37 -2442 38 -2440
rect 37 -2448 38 -2446
rect 44 -2442 45 -2440
rect 44 -2448 45 -2446
rect 51 -2442 52 -2440
rect 51 -2448 52 -2446
rect 58 -2442 59 -2440
rect 58 -2448 59 -2446
rect 65 -2442 66 -2440
rect 65 -2448 66 -2446
rect 72 -2442 73 -2440
rect 72 -2448 73 -2446
rect 82 -2442 83 -2440
rect 79 -2448 80 -2446
rect 82 -2448 83 -2446
rect 86 -2442 87 -2440
rect 86 -2448 87 -2446
rect 93 -2442 94 -2440
rect 96 -2442 97 -2440
rect 93 -2448 94 -2446
rect 96 -2448 97 -2446
rect 100 -2442 101 -2440
rect 100 -2448 101 -2446
rect 107 -2442 108 -2440
rect 110 -2442 111 -2440
rect 107 -2448 108 -2446
rect 110 -2448 111 -2446
rect 114 -2442 115 -2440
rect 114 -2448 115 -2446
rect 121 -2442 122 -2440
rect 121 -2448 122 -2446
rect 128 -2442 129 -2440
rect 131 -2442 132 -2440
rect 128 -2448 129 -2446
rect 131 -2448 132 -2446
rect 135 -2442 136 -2440
rect 135 -2448 136 -2446
rect 142 -2442 143 -2440
rect 142 -2448 143 -2446
rect 149 -2442 150 -2440
rect 149 -2448 150 -2446
rect 156 -2442 157 -2440
rect 156 -2448 157 -2446
rect 163 -2442 164 -2440
rect 163 -2448 164 -2446
rect 170 -2442 171 -2440
rect 170 -2448 171 -2446
rect 177 -2442 178 -2440
rect 177 -2448 178 -2446
rect 184 -2442 185 -2440
rect 184 -2448 185 -2446
rect 191 -2442 192 -2440
rect 191 -2448 192 -2446
rect 194 -2448 195 -2446
rect 198 -2442 199 -2440
rect 198 -2448 199 -2446
rect 205 -2442 206 -2440
rect 205 -2448 206 -2446
rect 212 -2442 213 -2440
rect 212 -2448 213 -2446
rect 219 -2442 220 -2440
rect 219 -2448 220 -2446
rect 226 -2442 227 -2440
rect 226 -2448 227 -2446
rect 233 -2442 234 -2440
rect 233 -2448 234 -2446
rect 240 -2442 241 -2440
rect 240 -2448 241 -2446
rect 247 -2442 248 -2440
rect 247 -2448 248 -2446
rect 254 -2442 255 -2440
rect 254 -2448 255 -2446
rect 261 -2442 262 -2440
rect 261 -2448 262 -2446
rect 268 -2442 269 -2440
rect 268 -2448 269 -2446
rect 275 -2442 276 -2440
rect 275 -2448 276 -2446
rect 282 -2442 283 -2440
rect 282 -2448 283 -2446
rect 289 -2442 290 -2440
rect 289 -2448 290 -2446
rect 296 -2442 297 -2440
rect 296 -2448 297 -2446
rect 303 -2442 304 -2440
rect 303 -2448 304 -2446
rect 310 -2442 311 -2440
rect 310 -2448 311 -2446
rect 317 -2442 318 -2440
rect 317 -2448 318 -2446
rect 324 -2442 325 -2440
rect 324 -2448 325 -2446
rect 331 -2442 332 -2440
rect 331 -2448 332 -2446
rect 338 -2442 339 -2440
rect 341 -2442 342 -2440
rect 338 -2448 339 -2446
rect 341 -2448 342 -2446
rect 345 -2442 346 -2440
rect 345 -2448 346 -2446
rect 352 -2442 353 -2440
rect 352 -2448 353 -2446
rect 359 -2442 360 -2440
rect 359 -2448 360 -2446
rect 366 -2442 367 -2440
rect 366 -2448 367 -2446
rect 373 -2442 374 -2440
rect 373 -2448 374 -2446
rect 380 -2442 381 -2440
rect 380 -2448 381 -2446
rect 387 -2442 388 -2440
rect 390 -2442 391 -2440
rect 387 -2448 388 -2446
rect 390 -2448 391 -2446
rect 394 -2442 395 -2440
rect 394 -2448 395 -2446
rect 401 -2442 402 -2440
rect 404 -2442 405 -2440
rect 401 -2448 402 -2446
rect 404 -2448 405 -2446
rect 408 -2442 409 -2440
rect 408 -2448 409 -2446
rect 415 -2442 416 -2440
rect 415 -2448 416 -2446
rect 422 -2442 423 -2440
rect 422 -2448 423 -2446
rect 429 -2442 430 -2440
rect 432 -2442 433 -2440
rect 432 -2448 433 -2446
rect 436 -2442 437 -2440
rect 439 -2442 440 -2440
rect 436 -2448 437 -2446
rect 439 -2448 440 -2446
rect 443 -2442 444 -2440
rect 446 -2442 447 -2440
rect 443 -2448 444 -2446
rect 450 -2442 451 -2440
rect 450 -2448 451 -2446
rect 457 -2442 458 -2440
rect 460 -2442 461 -2440
rect 457 -2448 458 -2446
rect 460 -2448 461 -2446
rect 464 -2442 465 -2440
rect 464 -2448 465 -2446
rect 471 -2442 472 -2440
rect 471 -2448 472 -2446
rect 478 -2442 479 -2440
rect 478 -2448 479 -2446
rect 485 -2442 486 -2440
rect 485 -2448 486 -2446
rect 492 -2442 493 -2440
rect 492 -2448 493 -2446
rect 499 -2442 500 -2440
rect 499 -2448 500 -2446
rect 506 -2442 507 -2440
rect 506 -2448 507 -2446
rect 513 -2442 514 -2440
rect 513 -2448 514 -2446
rect 516 -2448 517 -2446
rect 520 -2442 521 -2440
rect 520 -2448 521 -2446
rect 527 -2442 528 -2440
rect 530 -2442 531 -2440
rect 527 -2448 528 -2446
rect 530 -2448 531 -2446
rect 534 -2442 535 -2440
rect 534 -2448 535 -2446
rect 541 -2442 542 -2440
rect 544 -2442 545 -2440
rect 544 -2448 545 -2446
rect 548 -2442 549 -2440
rect 548 -2448 549 -2446
rect 555 -2442 556 -2440
rect 555 -2448 556 -2446
rect 562 -2442 563 -2440
rect 562 -2448 563 -2446
rect 569 -2442 570 -2440
rect 569 -2448 570 -2446
rect 576 -2442 577 -2440
rect 576 -2448 577 -2446
rect 583 -2442 584 -2440
rect 583 -2448 584 -2446
rect 590 -2442 591 -2440
rect 590 -2448 591 -2446
rect 597 -2442 598 -2440
rect 597 -2448 598 -2446
rect 600 -2448 601 -2446
rect 604 -2442 605 -2440
rect 604 -2448 605 -2446
rect 611 -2442 612 -2440
rect 611 -2448 612 -2446
rect 618 -2442 619 -2440
rect 618 -2448 619 -2446
rect 625 -2442 626 -2440
rect 625 -2448 626 -2446
rect 632 -2442 633 -2440
rect 632 -2448 633 -2446
rect 639 -2442 640 -2440
rect 639 -2448 640 -2446
rect 646 -2442 647 -2440
rect 646 -2448 647 -2446
rect 653 -2442 654 -2440
rect 653 -2448 654 -2446
rect 660 -2442 661 -2440
rect 660 -2448 661 -2446
rect 667 -2442 668 -2440
rect 667 -2448 668 -2446
rect 674 -2442 675 -2440
rect 677 -2442 678 -2440
rect 674 -2448 675 -2446
rect 677 -2448 678 -2446
rect 681 -2442 682 -2440
rect 681 -2448 682 -2446
rect 688 -2442 689 -2440
rect 688 -2448 689 -2446
rect 695 -2442 696 -2440
rect 698 -2442 699 -2440
rect 695 -2448 696 -2446
rect 702 -2442 703 -2440
rect 702 -2448 703 -2446
rect 709 -2442 710 -2440
rect 709 -2448 710 -2446
rect 716 -2448 717 -2446
rect 719 -2448 720 -2446
rect 723 -2442 724 -2440
rect 723 -2448 724 -2446
rect 730 -2442 731 -2440
rect 733 -2442 734 -2440
rect 730 -2448 731 -2446
rect 737 -2442 738 -2440
rect 737 -2448 738 -2446
rect 744 -2442 745 -2440
rect 744 -2448 745 -2446
rect 751 -2442 752 -2440
rect 751 -2448 752 -2446
rect 758 -2442 759 -2440
rect 758 -2448 759 -2446
rect 765 -2442 766 -2440
rect 765 -2448 766 -2446
rect 772 -2442 773 -2440
rect 772 -2448 773 -2446
rect 779 -2442 780 -2440
rect 779 -2448 780 -2446
rect 786 -2442 787 -2440
rect 786 -2448 787 -2446
rect 789 -2448 790 -2446
rect 793 -2442 794 -2440
rect 793 -2448 794 -2446
rect 800 -2442 801 -2440
rect 800 -2448 801 -2446
rect 807 -2442 808 -2440
rect 807 -2448 808 -2446
rect 814 -2442 815 -2440
rect 814 -2448 815 -2446
rect 821 -2442 822 -2440
rect 821 -2448 822 -2446
rect 828 -2442 829 -2440
rect 831 -2442 832 -2440
rect 828 -2448 829 -2446
rect 831 -2448 832 -2446
rect 835 -2442 836 -2440
rect 835 -2448 836 -2446
rect 842 -2442 843 -2440
rect 842 -2448 843 -2446
rect 849 -2442 850 -2440
rect 849 -2448 850 -2446
rect 856 -2442 857 -2440
rect 856 -2448 857 -2446
rect 863 -2442 864 -2440
rect 863 -2448 864 -2446
rect 870 -2442 871 -2440
rect 870 -2448 871 -2446
rect 877 -2442 878 -2440
rect 877 -2448 878 -2446
rect 884 -2442 885 -2440
rect 887 -2442 888 -2440
rect 884 -2448 885 -2446
rect 887 -2448 888 -2446
rect 891 -2442 892 -2440
rect 891 -2448 892 -2446
rect 898 -2442 899 -2440
rect 898 -2448 899 -2446
rect 905 -2442 906 -2440
rect 905 -2448 906 -2446
rect 912 -2442 913 -2440
rect 912 -2448 913 -2446
rect 919 -2442 920 -2440
rect 919 -2448 920 -2446
rect 926 -2442 927 -2440
rect 926 -2448 927 -2446
rect 933 -2442 934 -2440
rect 933 -2448 934 -2446
rect 940 -2442 941 -2440
rect 940 -2448 941 -2446
rect 947 -2442 948 -2440
rect 947 -2448 948 -2446
rect 954 -2442 955 -2440
rect 954 -2448 955 -2446
rect 961 -2442 962 -2440
rect 961 -2448 962 -2446
rect 968 -2442 969 -2440
rect 968 -2448 969 -2446
rect 975 -2442 976 -2440
rect 975 -2448 976 -2446
rect 982 -2442 983 -2440
rect 982 -2448 983 -2446
rect 989 -2442 990 -2440
rect 989 -2448 990 -2446
rect 996 -2442 997 -2440
rect 996 -2448 997 -2446
rect 1003 -2442 1004 -2440
rect 1003 -2448 1004 -2446
rect 1010 -2442 1011 -2440
rect 1010 -2448 1011 -2446
rect 1017 -2442 1018 -2440
rect 1020 -2442 1021 -2440
rect 1017 -2448 1018 -2446
rect 1020 -2448 1021 -2446
rect 1024 -2442 1025 -2440
rect 1024 -2448 1025 -2446
rect 1031 -2442 1032 -2440
rect 1031 -2448 1032 -2446
rect 1038 -2442 1039 -2440
rect 1038 -2448 1039 -2446
rect 1045 -2442 1046 -2440
rect 1045 -2448 1046 -2446
rect 1052 -2442 1053 -2440
rect 1055 -2442 1056 -2440
rect 1059 -2442 1060 -2440
rect 1059 -2448 1060 -2446
rect 1066 -2442 1067 -2440
rect 1066 -2448 1067 -2446
rect 1073 -2442 1074 -2440
rect 1073 -2448 1074 -2446
rect 1080 -2442 1081 -2440
rect 1083 -2442 1084 -2440
rect 1080 -2448 1081 -2446
rect 1087 -2442 1088 -2440
rect 1087 -2448 1088 -2446
rect 1094 -2442 1095 -2440
rect 1094 -2448 1095 -2446
rect 1101 -2442 1102 -2440
rect 1101 -2448 1102 -2446
rect 1108 -2442 1109 -2440
rect 1108 -2448 1109 -2446
rect 1115 -2442 1116 -2440
rect 1115 -2448 1116 -2446
rect 1122 -2442 1123 -2440
rect 1122 -2448 1123 -2446
rect 1129 -2442 1130 -2440
rect 1129 -2448 1130 -2446
rect 1136 -2442 1137 -2440
rect 1136 -2448 1137 -2446
rect 1143 -2442 1144 -2440
rect 1143 -2448 1144 -2446
rect 1150 -2442 1151 -2440
rect 1150 -2448 1151 -2446
rect 1157 -2442 1158 -2440
rect 1157 -2448 1158 -2446
rect 1164 -2442 1165 -2440
rect 1167 -2442 1168 -2440
rect 1164 -2448 1165 -2446
rect 1167 -2448 1168 -2446
rect 1171 -2442 1172 -2440
rect 1171 -2448 1172 -2446
rect 1178 -2442 1179 -2440
rect 1178 -2448 1179 -2446
rect 1185 -2442 1186 -2440
rect 1185 -2448 1186 -2446
rect 1192 -2442 1193 -2440
rect 1192 -2448 1193 -2446
rect 1199 -2442 1200 -2440
rect 1199 -2448 1200 -2446
rect 1206 -2442 1207 -2440
rect 1206 -2448 1207 -2446
rect 1213 -2442 1214 -2440
rect 1216 -2442 1217 -2440
rect 1213 -2448 1214 -2446
rect 1220 -2442 1221 -2440
rect 1220 -2448 1221 -2446
rect 1227 -2442 1228 -2440
rect 1227 -2448 1228 -2446
rect 1234 -2442 1235 -2440
rect 1234 -2448 1235 -2446
rect 1241 -2442 1242 -2440
rect 1241 -2448 1242 -2446
rect 1248 -2442 1249 -2440
rect 1248 -2448 1249 -2446
rect 1255 -2442 1256 -2440
rect 1255 -2448 1256 -2446
rect 1262 -2442 1263 -2440
rect 1262 -2448 1263 -2446
rect 1269 -2442 1270 -2440
rect 1269 -2448 1270 -2446
rect 1276 -2442 1277 -2440
rect 1276 -2448 1277 -2446
rect 1283 -2442 1284 -2440
rect 1283 -2448 1284 -2446
rect 1290 -2442 1291 -2440
rect 1290 -2448 1291 -2446
rect 1297 -2442 1298 -2440
rect 1297 -2448 1298 -2446
rect 1304 -2442 1305 -2440
rect 1304 -2448 1305 -2446
rect 1311 -2442 1312 -2440
rect 1311 -2448 1312 -2446
rect 1321 -2442 1322 -2440
rect 1318 -2448 1319 -2446
rect 1321 -2448 1322 -2446
rect 1325 -2442 1326 -2440
rect 1325 -2448 1326 -2446
rect 1332 -2442 1333 -2440
rect 1332 -2448 1333 -2446
rect 1339 -2442 1340 -2440
rect 1342 -2442 1343 -2440
rect 1346 -2442 1347 -2440
rect 1346 -2448 1347 -2446
rect 1353 -2442 1354 -2440
rect 1353 -2448 1354 -2446
rect 1360 -2442 1361 -2440
rect 1360 -2448 1361 -2446
rect 1367 -2442 1368 -2440
rect 1367 -2448 1368 -2446
rect 1374 -2442 1375 -2440
rect 1374 -2448 1375 -2446
rect 1381 -2442 1382 -2440
rect 1381 -2448 1382 -2446
rect 1388 -2442 1389 -2440
rect 1391 -2442 1392 -2440
rect 1388 -2448 1389 -2446
rect 1395 -2442 1396 -2440
rect 1395 -2448 1396 -2446
rect 1402 -2442 1403 -2440
rect 1402 -2448 1403 -2446
rect 1409 -2442 1410 -2440
rect 1409 -2448 1410 -2446
rect 1416 -2442 1417 -2440
rect 1416 -2448 1417 -2446
rect 1423 -2442 1424 -2440
rect 1423 -2448 1424 -2446
rect 1430 -2442 1431 -2440
rect 1430 -2448 1431 -2446
rect 1437 -2442 1438 -2440
rect 1437 -2448 1438 -2446
rect 1444 -2442 1445 -2440
rect 1444 -2448 1445 -2446
rect 1451 -2442 1452 -2440
rect 1451 -2448 1452 -2446
rect 1458 -2442 1459 -2440
rect 1458 -2448 1459 -2446
rect 1465 -2442 1466 -2440
rect 1465 -2448 1466 -2446
rect 1472 -2442 1473 -2440
rect 1472 -2448 1473 -2446
rect 1479 -2442 1480 -2440
rect 1479 -2448 1480 -2446
rect 1486 -2442 1487 -2440
rect 1486 -2448 1487 -2446
rect 1493 -2442 1494 -2440
rect 1493 -2448 1494 -2446
rect 1500 -2442 1501 -2440
rect 1500 -2448 1501 -2446
rect 1507 -2442 1508 -2440
rect 1507 -2448 1508 -2446
rect 1514 -2442 1515 -2440
rect 1514 -2448 1515 -2446
rect 1521 -2442 1522 -2440
rect 1521 -2448 1522 -2446
rect 1528 -2442 1529 -2440
rect 1528 -2448 1529 -2446
rect 1535 -2442 1536 -2440
rect 1535 -2448 1536 -2446
rect 1542 -2442 1543 -2440
rect 1542 -2448 1543 -2446
rect 1549 -2442 1550 -2440
rect 1549 -2448 1550 -2446
rect 1556 -2442 1557 -2440
rect 1556 -2448 1557 -2446
rect 1563 -2442 1564 -2440
rect 1563 -2448 1564 -2446
rect 1570 -2442 1571 -2440
rect 1570 -2448 1571 -2446
rect 1577 -2442 1578 -2440
rect 1577 -2448 1578 -2446
rect 1584 -2442 1585 -2440
rect 1584 -2448 1585 -2446
rect 1591 -2442 1592 -2440
rect 1591 -2448 1592 -2446
rect 1598 -2442 1599 -2440
rect 1598 -2448 1599 -2446
rect 1605 -2442 1606 -2440
rect 1605 -2448 1606 -2446
rect 1612 -2442 1613 -2440
rect 1612 -2448 1613 -2446
rect 1619 -2442 1620 -2440
rect 1619 -2448 1620 -2446
rect 1626 -2442 1627 -2440
rect 1626 -2448 1627 -2446
rect 1633 -2442 1634 -2440
rect 1633 -2448 1634 -2446
rect 1640 -2442 1641 -2440
rect 1640 -2448 1641 -2446
rect 1647 -2442 1648 -2440
rect 1647 -2448 1648 -2446
rect 1654 -2442 1655 -2440
rect 1654 -2448 1655 -2446
rect 1661 -2442 1662 -2440
rect 1661 -2448 1662 -2446
rect 1668 -2442 1669 -2440
rect 1668 -2448 1669 -2446
rect 1675 -2442 1676 -2440
rect 1675 -2448 1676 -2446
rect 1682 -2442 1683 -2440
rect 1682 -2448 1683 -2446
rect 1689 -2442 1690 -2440
rect 1689 -2448 1690 -2446
rect 1696 -2442 1697 -2440
rect 1696 -2448 1697 -2446
rect 1703 -2442 1704 -2440
rect 1703 -2448 1704 -2446
rect 1710 -2442 1711 -2440
rect 1710 -2448 1711 -2446
rect 1717 -2442 1718 -2440
rect 1717 -2448 1718 -2446
rect 1724 -2442 1725 -2440
rect 1724 -2448 1725 -2446
rect 1731 -2442 1732 -2440
rect 1731 -2448 1732 -2446
rect 1738 -2442 1739 -2440
rect 1738 -2448 1739 -2446
rect 1745 -2442 1746 -2440
rect 1745 -2448 1746 -2446
rect 1752 -2442 1753 -2440
rect 1755 -2442 1756 -2440
rect 1759 -2442 1760 -2440
rect 1759 -2448 1760 -2446
rect 1766 -2442 1767 -2440
rect 1766 -2448 1767 -2446
rect 1773 -2442 1774 -2440
rect 1773 -2448 1774 -2446
rect 1780 -2442 1781 -2440
rect 1780 -2448 1781 -2446
rect 1787 -2442 1788 -2440
rect 1787 -2448 1788 -2446
rect 1794 -2442 1795 -2440
rect 1797 -2442 1798 -2440
rect 1794 -2448 1795 -2446
rect 1801 -2442 1802 -2440
rect 1801 -2448 1802 -2446
rect 1808 -2442 1809 -2440
rect 1808 -2448 1809 -2446
rect 16 -2577 17 -2575
rect 16 -2583 17 -2581
rect 23 -2577 24 -2575
rect 23 -2583 24 -2581
rect 30 -2577 31 -2575
rect 30 -2583 31 -2581
rect 37 -2577 38 -2575
rect 37 -2583 38 -2581
rect 44 -2577 45 -2575
rect 44 -2583 45 -2581
rect 51 -2577 52 -2575
rect 51 -2583 52 -2581
rect 58 -2577 59 -2575
rect 58 -2583 59 -2581
rect 65 -2577 66 -2575
rect 65 -2583 66 -2581
rect 72 -2577 73 -2575
rect 72 -2583 73 -2581
rect 79 -2577 80 -2575
rect 79 -2583 80 -2581
rect 86 -2577 87 -2575
rect 86 -2583 87 -2581
rect 93 -2577 94 -2575
rect 93 -2583 94 -2581
rect 100 -2577 101 -2575
rect 103 -2577 104 -2575
rect 100 -2583 101 -2581
rect 103 -2583 104 -2581
rect 107 -2577 108 -2575
rect 110 -2577 111 -2575
rect 107 -2583 108 -2581
rect 110 -2583 111 -2581
rect 114 -2577 115 -2575
rect 114 -2583 115 -2581
rect 121 -2577 122 -2575
rect 121 -2583 122 -2581
rect 128 -2577 129 -2575
rect 128 -2583 129 -2581
rect 135 -2577 136 -2575
rect 135 -2583 136 -2581
rect 142 -2577 143 -2575
rect 142 -2583 143 -2581
rect 149 -2577 150 -2575
rect 152 -2577 153 -2575
rect 149 -2583 150 -2581
rect 152 -2583 153 -2581
rect 156 -2577 157 -2575
rect 159 -2577 160 -2575
rect 156 -2583 157 -2581
rect 159 -2583 160 -2581
rect 163 -2577 164 -2575
rect 163 -2583 164 -2581
rect 170 -2577 171 -2575
rect 173 -2577 174 -2575
rect 170 -2583 171 -2581
rect 173 -2583 174 -2581
rect 177 -2577 178 -2575
rect 177 -2583 178 -2581
rect 184 -2577 185 -2575
rect 184 -2583 185 -2581
rect 191 -2577 192 -2575
rect 191 -2583 192 -2581
rect 198 -2577 199 -2575
rect 198 -2583 199 -2581
rect 205 -2577 206 -2575
rect 205 -2583 206 -2581
rect 212 -2577 213 -2575
rect 212 -2583 213 -2581
rect 219 -2577 220 -2575
rect 219 -2583 220 -2581
rect 226 -2577 227 -2575
rect 226 -2583 227 -2581
rect 233 -2577 234 -2575
rect 233 -2583 234 -2581
rect 243 -2577 244 -2575
rect 243 -2583 244 -2581
rect 247 -2577 248 -2575
rect 247 -2583 248 -2581
rect 254 -2577 255 -2575
rect 254 -2583 255 -2581
rect 261 -2577 262 -2575
rect 261 -2583 262 -2581
rect 268 -2577 269 -2575
rect 268 -2583 269 -2581
rect 275 -2577 276 -2575
rect 275 -2583 276 -2581
rect 282 -2577 283 -2575
rect 282 -2583 283 -2581
rect 289 -2577 290 -2575
rect 289 -2583 290 -2581
rect 296 -2577 297 -2575
rect 296 -2583 297 -2581
rect 303 -2577 304 -2575
rect 303 -2583 304 -2581
rect 310 -2577 311 -2575
rect 310 -2583 311 -2581
rect 317 -2577 318 -2575
rect 317 -2583 318 -2581
rect 324 -2577 325 -2575
rect 324 -2583 325 -2581
rect 331 -2577 332 -2575
rect 331 -2583 332 -2581
rect 338 -2577 339 -2575
rect 338 -2583 339 -2581
rect 345 -2577 346 -2575
rect 345 -2583 346 -2581
rect 352 -2577 353 -2575
rect 352 -2583 353 -2581
rect 359 -2577 360 -2575
rect 359 -2583 360 -2581
rect 366 -2577 367 -2575
rect 366 -2583 367 -2581
rect 373 -2577 374 -2575
rect 373 -2583 374 -2581
rect 380 -2577 381 -2575
rect 380 -2583 381 -2581
rect 387 -2577 388 -2575
rect 387 -2583 388 -2581
rect 394 -2577 395 -2575
rect 394 -2583 395 -2581
rect 401 -2577 402 -2575
rect 401 -2583 402 -2581
rect 408 -2577 409 -2575
rect 408 -2583 409 -2581
rect 415 -2577 416 -2575
rect 415 -2583 416 -2581
rect 422 -2577 423 -2575
rect 422 -2583 423 -2581
rect 429 -2577 430 -2575
rect 429 -2583 430 -2581
rect 436 -2577 437 -2575
rect 436 -2583 437 -2581
rect 443 -2577 444 -2575
rect 443 -2583 444 -2581
rect 450 -2577 451 -2575
rect 453 -2577 454 -2575
rect 450 -2583 451 -2581
rect 453 -2583 454 -2581
rect 457 -2577 458 -2575
rect 457 -2583 458 -2581
rect 464 -2577 465 -2575
rect 464 -2583 465 -2581
rect 471 -2577 472 -2575
rect 471 -2583 472 -2581
rect 478 -2577 479 -2575
rect 478 -2583 479 -2581
rect 485 -2577 486 -2575
rect 485 -2583 486 -2581
rect 492 -2577 493 -2575
rect 492 -2583 493 -2581
rect 499 -2577 500 -2575
rect 499 -2583 500 -2581
rect 506 -2577 507 -2575
rect 506 -2583 507 -2581
rect 513 -2577 514 -2575
rect 513 -2583 514 -2581
rect 520 -2577 521 -2575
rect 520 -2583 521 -2581
rect 527 -2577 528 -2575
rect 527 -2583 528 -2581
rect 534 -2577 535 -2575
rect 534 -2583 535 -2581
rect 541 -2577 542 -2575
rect 541 -2583 542 -2581
rect 548 -2577 549 -2575
rect 548 -2583 549 -2581
rect 555 -2577 556 -2575
rect 558 -2577 559 -2575
rect 555 -2583 556 -2581
rect 558 -2583 559 -2581
rect 562 -2577 563 -2575
rect 562 -2583 563 -2581
rect 569 -2577 570 -2575
rect 569 -2583 570 -2581
rect 576 -2577 577 -2575
rect 576 -2583 577 -2581
rect 583 -2577 584 -2575
rect 583 -2583 584 -2581
rect 590 -2577 591 -2575
rect 590 -2583 591 -2581
rect 597 -2577 598 -2575
rect 600 -2577 601 -2575
rect 597 -2583 598 -2581
rect 604 -2577 605 -2575
rect 604 -2583 605 -2581
rect 611 -2577 612 -2575
rect 611 -2583 612 -2581
rect 618 -2577 619 -2575
rect 618 -2583 619 -2581
rect 625 -2577 626 -2575
rect 628 -2577 629 -2575
rect 625 -2583 626 -2581
rect 628 -2583 629 -2581
rect 632 -2577 633 -2575
rect 632 -2583 633 -2581
rect 639 -2577 640 -2575
rect 639 -2583 640 -2581
rect 646 -2577 647 -2575
rect 646 -2583 647 -2581
rect 653 -2577 654 -2575
rect 653 -2583 654 -2581
rect 660 -2577 661 -2575
rect 660 -2583 661 -2581
rect 670 -2577 671 -2575
rect 667 -2583 668 -2581
rect 670 -2583 671 -2581
rect 674 -2577 675 -2575
rect 674 -2583 675 -2581
rect 681 -2577 682 -2575
rect 681 -2583 682 -2581
rect 688 -2577 689 -2575
rect 688 -2583 689 -2581
rect 695 -2577 696 -2575
rect 695 -2583 696 -2581
rect 702 -2577 703 -2575
rect 702 -2583 703 -2581
rect 709 -2577 710 -2575
rect 712 -2577 713 -2575
rect 709 -2583 710 -2581
rect 712 -2583 713 -2581
rect 716 -2577 717 -2575
rect 716 -2583 717 -2581
rect 723 -2577 724 -2575
rect 726 -2577 727 -2575
rect 723 -2583 724 -2581
rect 726 -2583 727 -2581
rect 730 -2577 731 -2575
rect 730 -2583 731 -2581
rect 737 -2577 738 -2575
rect 740 -2577 741 -2575
rect 737 -2583 738 -2581
rect 740 -2583 741 -2581
rect 744 -2577 745 -2575
rect 744 -2583 745 -2581
rect 751 -2577 752 -2575
rect 751 -2583 752 -2581
rect 758 -2577 759 -2575
rect 758 -2583 759 -2581
rect 765 -2577 766 -2575
rect 765 -2583 766 -2581
rect 772 -2577 773 -2575
rect 772 -2583 773 -2581
rect 779 -2577 780 -2575
rect 779 -2583 780 -2581
rect 786 -2577 787 -2575
rect 786 -2583 787 -2581
rect 793 -2577 794 -2575
rect 793 -2583 794 -2581
rect 800 -2577 801 -2575
rect 800 -2583 801 -2581
rect 807 -2577 808 -2575
rect 807 -2583 808 -2581
rect 814 -2577 815 -2575
rect 814 -2583 815 -2581
rect 821 -2577 822 -2575
rect 821 -2583 822 -2581
rect 828 -2577 829 -2575
rect 828 -2583 829 -2581
rect 835 -2577 836 -2575
rect 835 -2583 836 -2581
rect 842 -2577 843 -2575
rect 842 -2583 843 -2581
rect 849 -2577 850 -2575
rect 852 -2577 853 -2575
rect 849 -2583 850 -2581
rect 852 -2583 853 -2581
rect 856 -2577 857 -2575
rect 856 -2583 857 -2581
rect 863 -2577 864 -2575
rect 863 -2583 864 -2581
rect 870 -2577 871 -2575
rect 870 -2583 871 -2581
rect 877 -2577 878 -2575
rect 877 -2583 878 -2581
rect 884 -2577 885 -2575
rect 884 -2583 885 -2581
rect 891 -2577 892 -2575
rect 891 -2583 892 -2581
rect 898 -2577 899 -2575
rect 898 -2583 899 -2581
rect 905 -2577 906 -2575
rect 905 -2583 906 -2581
rect 912 -2577 913 -2575
rect 912 -2583 913 -2581
rect 919 -2577 920 -2575
rect 919 -2583 920 -2581
rect 926 -2577 927 -2575
rect 926 -2583 927 -2581
rect 933 -2577 934 -2575
rect 933 -2583 934 -2581
rect 940 -2577 941 -2575
rect 940 -2583 941 -2581
rect 947 -2577 948 -2575
rect 950 -2577 951 -2575
rect 950 -2583 951 -2581
rect 954 -2577 955 -2575
rect 954 -2583 955 -2581
rect 961 -2577 962 -2575
rect 961 -2583 962 -2581
rect 968 -2577 969 -2575
rect 971 -2577 972 -2575
rect 968 -2583 969 -2581
rect 971 -2583 972 -2581
rect 975 -2577 976 -2575
rect 975 -2583 976 -2581
rect 982 -2577 983 -2575
rect 982 -2583 983 -2581
rect 989 -2577 990 -2575
rect 992 -2577 993 -2575
rect 989 -2583 990 -2581
rect 996 -2577 997 -2575
rect 996 -2583 997 -2581
rect 1003 -2577 1004 -2575
rect 1003 -2583 1004 -2581
rect 1010 -2577 1011 -2575
rect 1010 -2583 1011 -2581
rect 1017 -2577 1018 -2575
rect 1020 -2577 1021 -2575
rect 1017 -2583 1018 -2581
rect 1020 -2583 1021 -2581
rect 1024 -2577 1025 -2575
rect 1024 -2583 1025 -2581
rect 1031 -2577 1032 -2575
rect 1031 -2583 1032 -2581
rect 1038 -2577 1039 -2575
rect 1038 -2583 1039 -2581
rect 1045 -2577 1046 -2575
rect 1048 -2577 1049 -2575
rect 1045 -2583 1046 -2581
rect 1048 -2583 1049 -2581
rect 1052 -2577 1053 -2575
rect 1055 -2577 1056 -2575
rect 1052 -2583 1053 -2581
rect 1055 -2583 1056 -2581
rect 1059 -2577 1060 -2575
rect 1059 -2583 1060 -2581
rect 1066 -2577 1067 -2575
rect 1066 -2583 1067 -2581
rect 1076 -2577 1077 -2575
rect 1076 -2583 1077 -2581
rect 1080 -2577 1081 -2575
rect 1080 -2583 1081 -2581
rect 1087 -2577 1088 -2575
rect 1087 -2583 1088 -2581
rect 1094 -2577 1095 -2575
rect 1094 -2583 1095 -2581
rect 1101 -2577 1102 -2575
rect 1101 -2583 1102 -2581
rect 1108 -2577 1109 -2575
rect 1108 -2583 1109 -2581
rect 1115 -2577 1116 -2575
rect 1118 -2577 1119 -2575
rect 1118 -2583 1119 -2581
rect 1122 -2577 1123 -2575
rect 1122 -2583 1123 -2581
rect 1129 -2577 1130 -2575
rect 1132 -2577 1133 -2575
rect 1129 -2583 1130 -2581
rect 1132 -2583 1133 -2581
rect 1136 -2583 1137 -2581
rect 1139 -2583 1140 -2581
rect 1143 -2577 1144 -2575
rect 1143 -2583 1144 -2581
rect 1150 -2577 1151 -2575
rect 1150 -2583 1151 -2581
rect 1157 -2577 1158 -2575
rect 1160 -2577 1161 -2575
rect 1160 -2583 1161 -2581
rect 1164 -2577 1165 -2575
rect 1164 -2583 1165 -2581
rect 1171 -2577 1172 -2575
rect 1174 -2577 1175 -2575
rect 1171 -2583 1172 -2581
rect 1174 -2583 1175 -2581
rect 1178 -2577 1179 -2575
rect 1178 -2583 1179 -2581
rect 1185 -2577 1186 -2575
rect 1185 -2583 1186 -2581
rect 1192 -2577 1193 -2575
rect 1195 -2577 1196 -2575
rect 1192 -2583 1193 -2581
rect 1195 -2583 1196 -2581
rect 1199 -2577 1200 -2575
rect 1199 -2583 1200 -2581
rect 1206 -2577 1207 -2575
rect 1206 -2583 1207 -2581
rect 1213 -2577 1214 -2575
rect 1213 -2583 1214 -2581
rect 1220 -2577 1221 -2575
rect 1220 -2583 1221 -2581
rect 1227 -2577 1228 -2575
rect 1227 -2583 1228 -2581
rect 1234 -2577 1235 -2575
rect 1234 -2583 1235 -2581
rect 1241 -2577 1242 -2575
rect 1241 -2583 1242 -2581
rect 1248 -2577 1249 -2575
rect 1248 -2583 1249 -2581
rect 1255 -2577 1256 -2575
rect 1255 -2583 1256 -2581
rect 1262 -2577 1263 -2575
rect 1262 -2583 1263 -2581
rect 1269 -2577 1270 -2575
rect 1269 -2583 1270 -2581
rect 1276 -2577 1277 -2575
rect 1276 -2583 1277 -2581
rect 1283 -2577 1284 -2575
rect 1283 -2583 1284 -2581
rect 1290 -2577 1291 -2575
rect 1290 -2583 1291 -2581
rect 1297 -2577 1298 -2575
rect 1297 -2583 1298 -2581
rect 1304 -2577 1305 -2575
rect 1304 -2583 1305 -2581
rect 1311 -2577 1312 -2575
rect 1311 -2583 1312 -2581
rect 1318 -2577 1319 -2575
rect 1318 -2583 1319 -2581
rect 1325 -2577 1326 -2575
rect 1325 -2583 1326 -2581
rect 1332 -2577 1333 -2575
rect 1332 -2583 1333 -2581
rect 1339 -2577 1340 -2575
rect 1339 -2583 1340 -2581
rect 1346 -2577 1347 -2575
rect 1346 -2583 1347 -2581
rect 1353 -2577 1354 -2575
rect 1353 -2583 1354 -2581
rect 1360 -2577 1361 -2575
rect 1360 -2583 1361 -2581
rect 1367 -2577 1368 -2575
rect 1367 -2583 1368 -2581
rect 1374 -2577 1375 -2575
rect 1374 -2583 1375 -2581
rect 1381 -2577 1382 -2575
rect 1381 -2583 1382 -2581
rect 1388 -2577 1389 -2575
rect 1388 -2583 1389 -2581
rect 1395 -2577 1396 -2575
rect 1395 -2583 1396 -2581
rect 1402 -2577 1403 -2575
rect 1402 -2583 1403 -2581
rect 1409 -2577 1410 -2575
rect 1409 -2583 1410 -2581
rect 1416 -2577 1417 -2575
rect 1416 -2583 1417 -2581
rect 1423 -2577 1424 -2575
rect 1423 -2583 1424 -2581
rect 1430 -2577 1431 -2575
rect 1430 -2583 1431 -2581
rect 1437 -2577 1438 -2575
rect 1437 -2583 1438 -2581
rect 1444 -2577 1445 -2575
rect 1444 -2583 1445 -2581
rect 1451 -2577 1452 -2575
rect 1451 -2583 1452 -2581
rect 1458 -2577 1459 -2575
rect 1458 -2583 1459 -2581
rect 1465 -2577 1466 -2575
rect 1465 -2583 1466 -2581
rect 1472 -2577 1473 -2575
rect 1472 -2583 1473 -2581
rect 1479 -2577 1480 -2575
rect 1479 -2583 1480 -2581
rect 1486 -2577 1487 -2575
rect 1486 -2583 1487 -2581
rect 1493 -2577 1494 -2575
rect 1493 -2583 1494 -2581
rect 1500 -2577 1501 -2575
rect 1500 -2583 1501 -2581
rect 1507 -2583 1508 -2581
rect 1510 -2583 1511 -2581
rect 1514 -2577 1515 -2575
rect 1514 -2583 1515 -2581
rect 1521 -2577 1522 -2575
rect 1521 -2583 1522 -2581
rect 1528 -2577 1529 -2575
rect 1528 -2583 1529 -2581
rect 1535 -2577 1536 -2575
rect 1535 -2583 1536 -2581
rect 1542 -2577 1543 -2575
rect 1542 -2583 1543 -2581
rect 1549 -2577 1550 -2575
rect 1549 -2583 1550 -2581
rect 1556 -2577 1557 -2575
rect 1556 -2583 1557 -2581
rect 1563 -2577 1564 -2575
rect 1563 -2583 1564 -2581
rect 1570 -2577 1571 -2575
rect 1570 -2583 1571 -2581
rect 1577 -2577 1578 -2575
rect 1577 -2583 1578 -2581
rect 1584 -2577 1585 -2575
rect 1584 -2583 1585 -2581
rect 1591 -2577 1592 -2575
rect 1591 -2583 1592 -2581
rect 1598 -2577 1599 -2575
rect 1598 -2583 1599 -2581
rect 1605 -2577 1606 -2575
rect 1605 -2583 1606 -2581
rect 1612 -2577 1613 -2575
rect 1612 -2583 1613 -2581
rect 1619 -2577 1620 -2575
rect 1619 -2583 1620 -2581
rect 1626 -2577 1627 -2575
rect 1626 -2583 1627 -2581
rect 1633 -2577 1634 -2575
rect 1633 -2583 1634 -2581
rect 1640 -2577 1641 -2575
rect 1640 -2583 1641 -2581
rect 1647 -2577 1648 -2575
rect 1647 -2583 1648 -2581
rect 1654 -2577 1655 -2575
rect 1654 -2583 1655 -2581
rect 1661 -2577 1662 -2575
rect 1661 -2583 1662 -2581
rect 1668 -2577 1669 -2575
rect 1668 -2583 1669 -2581
rect 1675 -2577 1676 -2575
rect 1675 -2583 1676 -2581
rect 1682 -2577 1683 -2575
rect 1682 -2583 1683 -2581
rect 1689 -2577 1690 -2575
rect 1689 -2583 1690 -2581
rect 1696 -2577 1697 -2575
rect 1699 -2577 1700 -2575
rect 1696 -2583 1697 -2581
rect 1699 -2583 1700 -2581
rect 1703 -2577 1704 -2575
rect 1703 -2583 1704 -2581
rect 1710 -2577 1711 -2575
rect 1710 -2583 1711 -2581
rect 1717 -2577 1718 -2575
rect 1717 -2583 1718 -2581
rect 1724 -2577 1725 -2575
rect 1724 -2583 1725 -2581
rect 1731 -2577 1732 -2575
rect 1731 -2583 1732 -2581
rect 1738 -2577 1739 -2575
rect 1741 -2577 1742 -2575
rect 1738 -2583 1739 -2581
rect 1741 -2583 1742 -2581
rect 1745 -2577 1746 -2575
rect 1745 -2583 1746 -2581
rect 1752 -2577 1753 -2575
rect 1752 -2583 1753 -2581
rect 1759 -2577 1760 -2575
rect 1759 -2583 1760 -2581
rect 1766 -2577 1767 -2575
rect 1766 -2583 1767 -2581
rect 1773 -2577 1774 -2575
rect 1773 -2583 1774 -2581
rect 1780 -2577 1781 -2575
rect 1780 -2583 1781 -2581
rect 1787 -2577 1788 -2575
rect 1787 -2583 1788 -2581
rect 1794 -2583 1795 -2581
rect 1801 -2577 1802 -2575
rect 1801 -2583 1802 -2581
rect 1808 -2577 1809 -2575
rect 1808 -2583 1809 -2581
rect 1815 -2577 1816 -2575
rect 1815 -2583 1816 -2581
rect 9 -2710 10 -2708
rect 9 -2716 10 -2714
rect 16 -2710 17 -2708
rect 30 -2710 31 -2708
rect 30 -2716 31 -2714
rect 37 -2710 38 -2708
rect 37 -2716 38 -2714
rect 44 -2710 45 -2708
rect 44 -2716 45 -2714
rect 51 -2710 52 -2708
rect 51 -2716 52 -2714
rect 58 -2710 59 -2708
rect 58 -2716 59 -2714
rect 61 -2716 62 -2714
rect 68 -2710 69 -2708
rect 68 -2716 69 -2714
rect 72 -2710 73 -2708
rect 72 -2716 73 -2714
rect 79 -2710 80 -2708
rect 79 -2716 80 -2714
rect 86 -2710 87 -2708
rect 86 -2716 87 -2714
rect 93 -2710 94 -2708
rect 93 -2716 94 -2714
rect 100 -2710 101 -2708
rect 100 -2716 101 -2714
rect 107 -2710 108 -2708
rect 107 -2716 108 -2714
rect 114 -2710 115 -2708
rect 114 -2716 115 -2714
rect 121 -2710 122 -2708
rect 121 -2716 122 -2714
rect 128 -2710 129 -2708
rect 128 -2716 129 -2714
rect 135 -2710 136 -2708
rect 135 -2716 136 -2714
rect 142 -2710 143 -2708
rect 142 -2716 143 -2714
rect 149 -2710 150 -2708
rect 149 -2716 150 -2714
rect 156 -2710 157 -2708
rect 156 -2716 157 -2714
rect 163 -2710 164 -2708
rect 163 -2716 164 -2714
rect 170 -2710 171 -2708
rect 170 -2716 171 -2714
rect 177 -2710 178 -2708
rect 177 -2716 178 -2714
rect 184 -2710 185 -2708
rect 184 -2716 185 -2714
rect 191 -2710 192 -2708
rect 191 -2716 192 -2714
rect 198 -2710 199 -2708
rect 201 -2710 202 -2708
rect 198 -2716 199 -2714
rect 201 -2716 202 -2714
rect 205 -2710 206 -2708
rect 208 -2710 209 -2708
rect 208 -2716 209 -2714
rect 212 -2710 213 -2708
rect 212 -2716 213 -2714
rect 219 -2710 220 -2708
rect 219 -2716 220 -2714
rect 226 -2710 227 -2708
rect 226 -2716 227 -2714
rect 233 -2710 234 -2708
rect 233 -2716 234 -2714
rect 240 -2710 241 -2708
rect 240 -2716 241 -2714
rect 247 -2710 248 -2708
rect 247 -2716 248 -2714
rect 254 -2710 255 -2708
rect 254 -2716 255 -2714
rect 261 -2710 262 -2708
rect 261 -2716 262 -2714
rect 268 -2710 269 -2708
rect 268 -2716 269 -2714
rect 275 -2710 276 -2708
rect 275 -2716 276 -2714
rect 282 -2710 283 -2708
rect 282 -2716 283 -2714
rect 289 -2710 290 -2708
rect 292 -2710 293 -2708
rect 292 -2716 293 -2714
rect 296 -2710 297 -2708
rect 296 -2716 297 -2714
rect 303 -2710 304 -2708
rect 303 -2716 304 -2714
rect 310 -2710 311 -2708
rect 310 -2716 311 -2714
rect 317 -2710 318 -2708
rect 317 -2716 318 -2714
rect 324 -2710 325 -2708
rect 324 -2716 325 -2714
rect 331 -2710 332 -2708
rect 331 -2716 332 -2714
rect 338 -2710 339 -2708
rect 338 -2716 339 -2714
rect 345 -2710 346 -2708
rect 345 -2716 346 -2714
rect 352 -2710 353 -2708
rect 352 -2716 353 -2714
rect 359 -2710 360 -2708
rect 359 -2716 360 -2714
rect 366 -2710 367 -2708
rect 366 -2716 367 -2714
rect 373 -2710 374 -2708
rect 373 -2716 374 -2714
rect 380 -2710 381 -2708
rect 380 -2716 381 -2714
rect 387 -2710 388 -2708
rect 387 -2716 388 -2714
rect 394 -2710 395 -2708
rect 394 -2716 395 -2714
rect 401 -2710 402 -2708
rect 401 -2716 402 -2714
rect 408 -2710 409 -2708
rect 408 -2716 409 -2714
rect 415 -2710 416 -2708
rect 415 -2716 416 -2714
rect 422 -2710 423 -2708
rect 425 -2710 426 -2708
rect 422 -2716 423 -2714
rect 425 -2716 426 -2714
rect 429 -2710 430 -2708
rect 429 -2716 430 -2714
rect 436 -2710 437 -2708
rect 436 -2716 437 -2714
rect 443 -2710 444 -2708
rect 443 -2716 444 -2714
rect 450 -2710 451 -2708
rect 450 -2716 451 -2714
rect 457 -2710 458 -2708
rect 457 -2716 458 -2714
rect 464 -2710 465 -2708
rect 464 -2716 465 -2714
rect 471 -2710 472 -2708
rect 471 -2716 472 -2714
rect 478 -2710 479 -2708
rect 478 -2716 479 -2714
rect 485 -2710 486 -2708
rect 485 -2716 486 -2714
rect 492 -2710 493 -2708
rect 492 -2716 493 -2714
rect 499 -2710 500 -2708
rect 499 -2716 500 -2714
rect 506 -2710 507 -2708
rect 506 -2716 507 -2714
rect 513 -2710 514 -2708
rect 513 -2716 514 -2714
rect 520 -2710 521 -2708
rect 523 -2710 524 -2708
rect 520 -2716 521 -2714
rect 523 -2716 524 -2714
rect 527 -2710 528 -2708
rect 527 -2716 528 -2714
rect 534 -2710 535 -2708
rect 534 -2716 535 -2714
rect 541 -2710 542 -2708
rect 541 -2716 542 -2714
rect 548 -2710 549 -2708
rect 548 -2716 549 -2714
rect 555 -2710 556 -2708
rect 555 -2716 556 -2714
rect 562 -2710 563 -2708
rect 562 -2716 563 -2714
rect 569 -2710 570 -2708
rect 569 -2716 570 -2714
rect 576 -2710 577 -2708
rect 576 -2716 577 -2714
rect 583 -2710 584 -2708
rect 586 -2710 587 -2708
rect 583 -2716 584 -2714
rect 590 -2710 591 -2708
rect 590 -2716 591 -2714
rect 597 -2710 598 -2708
rect 597 -2716 598 -2714
rect 604 -2710 605 -2708
rect 607 -2716 608 -2714
rect 611 -2710 612 -2708
rect 611 -2716 612 -2714
rect 618 -2710 619 -2708
rect 618 -2716 619 -2714
rect 625 -2710 626 -2708
rect 625 -2716 626 -2714
rect 632 -2710 633 -2708
rect 635 -2710 636 -2708
rect 632 -2716 633 -2714
rect 635 -2716 636 -2714
rect 642 -2710 643 -2708
rect 639 -2716 640 -2714
rect 642 -2716 643 -2714
rect 646 -2710 647 -2708
rect 646 -2716 647 -2714
rect 653 -2710 654 -2708
rect 653 -2716 654 -2714
rect 660 -2710 661 -2708
rect 660 -2716 661 -2714
rect 667 -2710 668 -2708
rect 667 -2716 668 -2714
rect 674 -2710 675 -2708
rect 674 -2716 675 -2714
rect 681 -2710 682 -2708
rect 681 -2716 682 -2714
rect 688 -2710 689 -2708
rect 688 -2716 689 -2714
rect 695 -2710 696 -2708
rect 695 -2716 696 -2714
rect 702 -2710 703 -2708
rect 702 -2716 703 -2714
rect 709 -2710 710 -2708
rect 712 -2710 713 -2708
rect 709 -2716 710 -2714
rect 712 -2716 713 -2714
rect 716 -2710 717 -2708
rect 716 -2716 717 -2714
rect 723 -2710 724 -2708
rect 723 -2716 724 -2714
rect 730 -2710 731 -2708
rect 730 -2716 731 -2714
rect 737 -2710 738 -2708
rect 737 -2716 738 -2714
rect 744 -2710 745 -2708
rect 744 -2716 745 -2714
rect 751 -2710 752 -2708
rect 751 -2716 752 -2714
rect 758 -2710 759 -2708
rect 758 -2716 759 -2714
rect 765 -2710 766 -2708
rect 765 -2716 766 -2714
rect 772 -2710 773 -2708
rect 775 -2710 776 -2708
rect 775 -2716 776 -2714
rect 779 -2710 780 -2708
rect 779 -2716 780 -2714
rect 786 -2710 787 -2708
rect 786 -2716 787 -2714
rect 793 -2710 794 -2708
rect 793 -2716 794 -2714
rect 800 -2710 801 -2708
rect 800 -2716 801 -2714
rect 807 -2710 808 -2708
rect 807 -2716 808 -2714
rect 814 -2710 815 -2708
rect 814 -2716 815 -2714
rect 821 -2710 822 -2708
rect 821 -2716 822 -2714
rect 828 -2710 829 -2708
rect 828 -2716 829 -2714
rect 835 -2710 836 -2708
rect 835 -2716 836 -2714
rect 842 -2710 843 -2708
rect 845 -2710 846 -2708
rect 842 -2716 843 -2714
rect 845 -2716 846 -2714
rect 849 -2710 850 -2708
rect 852 -2710 853 -2708
rect 856 -2710 857 -2708
rect 856 -2716 857 -2714
rect 866 -2710 867 -2708
rect 863 -2716 864 -2714
rect 866 -2716 867 -2714
rect 870 -2710 871 -2708
rect 870 -2716 871 -2714
rect 877 -2710 878 -2708
rect 877 -2716 878 -2714
rect 884 -2716 885 -2714
rect 887 -2716 888 -2714
rect 891 -2710 892 -2708
rect 891 -2716 892 -2714
rect 898 -2710 899 -2708
rect 898 -2716 899 -2714
rect 905 -2710 906 -2708
rect 905 -2716 906 -2714
rect 912 -2710 913 -2708
rect 915 -2710 916 -2708
rect 912 -2716 913 -2714
rect 915 -2716 916 -2714
rect 919 -2716 920 -2714
rect 926 -2710 927 -2708
rect 926 -2716 927 -2714
rect 933 -2710 934 -2708
rect 933 -2716 934 -2714
rect 940 -2710 941 -2708
rect 940 -2716 941 -2714
rect 947 -2710 948 -2708
rect 947 -2716 948 -2714
rect 954 -2710 955 -2708
rect 954 -2716 955 -2714
rect 961 -2710 962 -2708
rect 961 -2716 962 -2714
rect 968 -2710 969 -2708
rect 968 -2716 969 -2714
rect 975 -2710 976 -2708
rect 978 -2710 979 -2708
rect 975 -2716 976 -2714
rect 978 -2716 979 -2714
rect 982 -2710 983 -2708
rect 982 -2716 983 -2714
rect 989 -2710 990 -2708
rect 989 -2716 990 -2714
rect 996 -2710 997 -2708
rect 996 -2716 997 -2714
rect 1003 -2710 1004 -2708
rect 1003 -2716 1004 -2714
rect 1010 -2710 1011 -2708
rect 1010 -2716 1011 -2714
rect 1017 -2710 1018 -2708
rect 1020 -2710 1021 -2708
rect 1020 -2716 1021 -2714
rect 1024 -2710 1025 -2708
rect 1024 -2716 1025 -2714
rect 1031 -2710 1032 -2708
rect 1031 -2716 1032 -2714
rect 1038 -2710 1039 -2708
rect 1038 -2716 1039 -2714
rect 1045 -2710 1046 -2708
rect 1045 -2716 1046 -2714
rect 1052 -2710 1053 -2708
rect 1055 -2710 1056 -2708
rect 1052 -2716 1053 -2714
rect 1059 -2710 1060 -2708
rect 1062 -2710 1063 -2708
rect 1059 -2716 1060 -2714
rect 1062 -2716 1063 -2714
rect 1066 -2710 1067 -2708
rect 1066 -2716 1067 -2714
rect 1073 -2710 1074 -2708
rect 1073 -2716 1074 -2714
rect 1080 -2710 1081 -2708
rect 1080 -2716 1081 -2714
rect 1087 -2710 1088 -2708
rect 1087 -2716 1088 -2714
rect 1094 -2710 1095 -2708
rect 1094 -2716 1095 -2714
rect 1101 -2710 1102 -2708
rect 1101 -2716 1102 -2714
rect 1108 -2710 1109 -2708
rect 1108 -2716 1109 -2714
rect 1115 -2710 1116 -2708
rect 1115 -2716 1116 -2714
rect 1122 -2710 1123 -2708
rect 1122 -2716 1123 -2714
rect 1129 -2710 1130 -2708
rect 1129 -2716 1130 -2714
rect 1136 -2710 1137 -2708
rect 1136 -2716 1137 -2714
rect 1143 -2710 1144 -2708
rect 1143 -2716 1144 -2714
rect 1150 -2710 1151 -2708
rect 1150 -2716 1151 -2714
rect 1153 -2716 1154 -2714
rect 1157 -2710 1158 -2708
rect 1157 -2716 1158 -2714
rect 1164 -2710 1165 -2708
rect 1164 -2716 1165 -2714
rect 1171 -2710 1172 -2708
rect 1171 -2716 1172 -2714
rect 1178 -2710 1179 -2708
rect 1178 -2716 1179 -2714
rect 1185 -2710 1186 -2708
rect 1185 -2716 1186 -2714
rect 1192 -2710 1193 -2708
rect 1195 -2710 1196 -2708
rect 1192 -2716 1193 -2714
rect 1195 -2716 1196 -2714
rect 1199 -2710 1200 -2708
rect 1199 -2716 1200 -2714
rect 1206 -2710 1207 -2708
rect 1206 -2716 1207 -2714
rect 1213 -2710 1214 -2708
rect 1213 -2716 1214 -2714
rect 1220 -2710 1221 -2708
rect 1220 -2716 1221 -2714
rect 1227 -2710 1228 -2708
rect 1227 -2716 1228 -2714
rect 1234 -2710 1235 -2708
rect 1234 -2716 1235 -2714
rect 1241 -2710 1242 -2708
rect 1244 -2710 1245 -2708
rect 1241 -2716 1242 -2714
rect 1244 -2716 1245 -2714
rect 1248 -2710 1249 -2708
rect 1248 -2716 1249 -2714
rect 1255 -2710 1256 -2708
rect 1255 -2716 1256 -2714
rect 1262 -2710 1263 -2708
rect 1262 -2716 1263 -2714
rect 1269 -2710 1270 -2708
rect 1269 -2716 1270 -2714
rect 1276 -2710 1277 -2708
rect 1276 -2716 1277 -2714
rect 1283 -2710 1284 -2708
rect 1283 -2716 1284 -2714
rect 1293 -2710 1294 -2708
rect 1297 -2710 1298 -2708
rect 1297 -2716 1298 -2714
rect 1304 -2710 1305 -2708
rect 1304 -2716 1305 -2714
rect 1311 -2710 1312 -2708
rect 1311 -2716 1312 -2714
rect 1318 -2710 1319 -2708
rect 1321 -2710 1322 -2708
rect 1318 -2716 1319 -2714
rect 1321 -2716 1322 -2714
rect 1325 -2710 1326 -2708
rect 1325 -2716 1326 -2714
rect 1328 -2716 1329 -2714
rect 1332 -2710 1333 -2708
rect 1332 -2716 1333 -2714
rect 1339 -2710 1340 -2708
rect 1339 -2716 1340 -2714
rect 1346 -2710 1347 -2708
rect 1346 -2716 1347 -2714
rect 1353 -2710 1354 -2708
rect 1353 -2716 1354 -2714
rect 1360 -2710 1361 -2708
rect 1360 -2716 1361 -2714
rect 1367 -2710 1368 -2708
rect 1367 -2716 1368 -2714
rect 1374 -2710 1375 -2708
rect 1374 -2716 1375 -2714
rect 1381 -2710 1382 -2708
rect 1381 -2716 1382 -2714
rect 1388 -2710 1389 -2708
rect 1388 -2716 1389 -2714
rect 1395 -2710 1396 -2708
rect 1395 -2716 1396 -2714
rect 1402 -2710 1403 -2708
rect 1402 -2716 1403 -2714
rect 1409 -2710 1410 -2708
rect 1409 -2716 1410 -2714
rect 1416 -2710 1417 -2708
rect 1416 -2716 1417 -2714
rect 1423 -2710 1424 -2708
rect 1423 -2716 1424 -2714
rect 1430 -2710 1431 -2708
rect 1430 -2716 1431 -2714
rect 1437 -2710 1438 -2708
rect 1437 -2716 1438 -2714
rect 1444 -2710 1445 -2708
rect 1444 -2716 1445 -2714
rect 1451 -2710 1452 -2708
rect 1451 -2716 1452 -2714
rect 1458 -2710 1459 -2708
rect 1458 -2716 1459 -2714
rect 1465 -2710 1466 -2708
rect 1465 -2716 1466 -2714
rect 1472 -2710 1473 -2708
rect 1472 -2716 1473 -2714
rect 1479 -2710 1480 -2708
rect 1479 -2716 1480 -2714
rect 1486 -2710 1487 -2708
rect 1486 -2716 1487 -2714
rect 1493 -2710 1494 -2708
rect 1493 -2716 1494 -2714
rect 1500 -2710 1501 -2708
rect 1500 -2716 1501 -2714
rect 1507 -2710 1508 -2708
rect 1507 -2716 1508 -2714
rect 1514 -2710 1515 -2708
rect 1514 -2716 1515 -2714
rect 1521 -2710 1522 -2708
rect 1521 -2716 1522 -2714
rect 1528 -2710 1529 -2708
rect 1528 -2716 1529 -2714
rect 1535 -2710 1536 -2708
rect 1535 -2716 1536 -2714
rect 1542 -2710 1543 -2708
rect 1542 -2716 1543 -2714
rect 1549 -2710 1550 -2708
rect 1549 -2716 1550 -2714
rect 1556 -2710 1557 -2708
rect 1556 -2716 1557 -2714
rect 1563 -2710 1564 -2708
rect 1563 -2716 1564 -2714
rect 1570 -2710 1571 -2708
rect 1570 -2716 1571 -2714
rect 1577 -2710 1578 -2708
rect 1577 -2716 1578 -2714
rect 1584 -2710 1585 -2708
rect 1584 -2716 1585 -2714
rect 1591 -2710 1592 -2708
rect 1591 -2716 1592 -2714
rect 1598 -2710 1599 -2708
rect 1598 -2716 1599 -2714
rect 1605 -2710 1606 -2708
rect 1605 -2716 1606 -2714
rect 1612 -2710 1613 -2708
rect 1612 -2716 1613 -2714
rect 1619 -2710 1620 -2708
rect 1619 -2716 1620 -2714
rect 1626 -2710 1627 -2708
rect 1626 -2716 1627 -2714
rect 1633 -2710 1634 -2708
rect 1633 -2716 1634 -2714
rect 1640 -2710 1641 -2708
rect 1640 -2716 1641 -2714
rect 1647 -2710 1648 -2708
rect 1647 -2716 1648 -2714
rect 1654 -2710 1655 -2708
rect 1654 -2716 1655 -2714
rect 1661 -2710 1662 -2708
rect 1661 -2716 1662 -2714
rect 1668 -2710 1669 -2708
rect 1668 -2716 1669 -2714
rect 1675 -2710 1676 -2708
rect 1675 -2716 1676 -2714
rect 1682 -2710 1683 -2708
rect 1682 -2716 1683 -2714
rect 1689 -2710 1690 -2708
rect 1689 -2716 1690 -2714
rect 1696 -2710 1697 -2708
rect 1696 -2716 1697 -2714
rect 1703 -2710 1704 -2708
rect 1703 -2716 1704 -2714
rect 1710 -2710 1711 -2708
rect 1710 -2716 1711 -2714
rect 1717 -2710 1718 -2708
rect 1717 -2716 1718 -2714
rect 1724 -2710 1725 -2708
rect 1724 -2716 1725 -2714
rect 1731 -2710 1732 -2708
rect 1731 -2716 1732 -2714
rect 1738 -2710 1739 -2708
rect 1738 -2716 1739 -2714
rect 1745 -2710 1746 -2708
rect 1745 -2716 1746 -2714
rect 1752 -2710 1753 -2708
rect 1752 -2716 1753 -2714
rect 1759 -2710 1760 -2708
rect 1759 -2716 1760 -2714
rect 1766 -2710 1767 -2708
rect 1769 -2710 1770 -2708
rect 1766 -2716 1767 -2714
rect 1769 -2716 1770 -2714
rect 1773 -2710 1774 -2708
rect 1776 -2710 1777 -2708
rect 1773 -2716 1774 -2714
rect 1776 -2716 1777 -2714
rect 1783 -2710 1784 -2708
rect 1780 -2716 1781 -2714
rect 1783 -2716 1784 -2714
rect 1787 -2710 1788 -2708
rect 1787 -2716 1788 -2714
rect 1794 -2710 1795 -2708
rect 1794 -2716 1795 -2714
rect 1801 -2710 1802 -2708
rect 1801 -2716 1802 -2714
rect 1808 -2710 1809 -2708
rect 1808 -2716 1809 -2714
rect 37 -2831 38 -2829
rect 37 -2837 38 -2835
rect 44 -2831 45 -2829
rect 44 -2837 45 -2835
rect 51 -2831 52 -2829
rect 51 -2837 52 -2835
rect 58 -2831 59 -2829
rect 58 -2837 59 -2835
rect 65 -2831 66 -2829
rect 65 -2837 66 -2835
rect 72 -2831 73 -2829
rect 72 -2837 73 -2835
rect 79 -2831 80 -2829
rect 79 -2837 80 -2835
rect 86 -2831 87 -2829
rect 86 -2837 87 -2835
rect 93 -2831 94 -2829
rect 96 -2831 97 -2829
rect 93 -2837 94 -2835
rect 96 -2837 97 -2835
rect 100 -2831 101 -2829
rect 100 -2837 101 -2835
rect 107 -2831 108 -2829
rect 107 -2837 108 -2835
rect 114 -2831 115 -2829
rect 114 -2837 115 -2835
rect 121 -2831 122 -2829
rect 121 -2837 122 -2835
rect 128 -2831 129 -2829
rect 128 -2837 129 -2835
rect 135 -2831 136 -2829
rect 135 -2837 136 -2835
rect 142 -2831 143 -2829
rect 142 -2837 143 -2835
rect 149 -2831 150 -2829
rect 149 -2837 150 -2835
rect 156 -2831 157 -2829
rect 156 -2837 157 -2835
rect 163 -2831 164 -2829
rect 163 -2837 164 -2835
rect 170 -2831 171 -2829
rect 170 -2837 171 -2835
rect 177 -2831 178 -2829
rect 177 -2837 178 -2835
rect 184 -2831 185 -2829
rect 184 -2837 185 -2835
rect 191 -2831 192 -2829
rect 191 -2837 192 -2835
rect 198 -2831 199 -2829
rect 198 -2837 199 -2835
rect 205 -2831 206 -2829
rect 205 -2837 206 -2835
rect 212 -2831 213 -2829
rect 212 -2837 213 -2835
rect 219 -2831 220 -2829
rect 219 -2837 220 -2835
rect 226 -2831 227 -2829
rect 226 -2837 227 -2835
rect 233 -2831 234 -2829
rect 233 -2837 234 -2835
rect 240 -2831 241 -2829
rect 240 -2837 241 -2835
rect 247 -2831 248 -2829
rect 247 -2837 248 -2835
rect 254 -2831 255 -2829
rect 254 -2837 255 -2835
rect 261 -2831 262 -2829
rect 261 -2837 262 -2835
rect 268 -2831 269 -2829
rect 268 -2837 269 -2835
rect 275 -2831 276 -2829
rect 275 -2837 276 -2835
rect 282 -2831 283 -2829
rect 282 -2837 283 -2835
rect 289 -2831 290 -2829
rect 289 -2837 290 -2835
rect 296 -2831 297 -2829
rect 296 -2837 297 -2835
rect 303 -2831 304 -2829
rect 303 -2837 304 -2835
rect 310 -2831 311 -2829
rect 310 -2837 311 -2835
rect 317 -2831 318 -2829
rect 317 -2837 318 -2835
rect 324 -2831 325 -2829
rect 324 -2837 325 -2835
rect 331 -2831 332 -2829
rect 331 -2837 332 -2835
rect 338 -2831 339 -2829
rect 338 -2837 339 -2835
rect 345 -2831 346 -2829
rect 345 -2837 346 -2835
rect 355 -2831 356 -2829
rect 355 -2837 356 -2835
rect 359 -2831 360 -2829
rect 359 -2837 360 -2835
rect 366 -2831 367 -2829
rect 366 -2837 367 -2835
rect 373 -2831 374 -2829
rect 373 -2837 374 -2835
rect 380 -2831 381 -2829
rect 380 -2837 381 -2835
rect 387 -2831 388 -2829
rect 387 -2837 388 -2835
rect 394 -2831 395 -2829
rect 394 -2837 395 -2835
rect 401 -2831 402 -2829
rect 401 -2837 402 -2835
rect 408 -2831 409 -2829
rect 408 -2837 409 -2835
rect 415 -2831 416 -2829
rect 415 -2837 416 -2835
rect 422 -2831 423 -2829
rect 422 -2837 423 -2835
rect 429 -2831 430 -2829
rect 429 -2837 430 -2835
rect 436 -2831 437 -2829
rect 436 -2837 437 -2835
rect 443 -2831 444 -2829
rect 443 -2837 444 -2835
rect 450 -2831 451 -2829
rect 450 -2837 451 -2835
rect 457 -2831 458 -2829
rect 457 -2837 458 -2835
rect 464 -2831 465 -2829
rect 464 -2837 465 -2835
rect 471 -2831 472 -2829
rect 471 -2837 472 -2835
rect 478 -2831 479 -2829
rect 481 -2831 482 -2829
rect 478 -2837 479 -2835
rect 481 -2837 482 -2835
rect 485 -2831 486 -2829
rect 485 -2837 486 -2835
rect 492 -2831 493 -2829
rect 492 -2837 493 -2835
rect 499 -2831 500 -2829
rect 499 -2837 500 -2835
rect 506 -2831 507 -2829
rect 506 -2837 507 -2835
rect 513 -2831 514 -2829
rect 513 -2837 514 -2835
rect 520 -2831 521 -2829
rect 520 -2837 521 -2835
rect 527 -2831 528 -2829
rect 527 -2837 528 -2835
rect 534 -2831 535 -2829
rect 534 -2837 535 -2835
rect 541 -2831 542 -2829
rect 541 -2837 542 -2835
rect 548 -2831 549 -2829
rect 548 -2837 549 -2835
rect 555 -2831 556 -2829
rect 555 -2837 556 -2835
rect 558 -2837 559 -2835
rect 562 -2831 563 -2829
rect 565 -2831 566 -2829
rect 562 -2837 563 -2835
rect 565 -2837 566 -2835
rect 569 -2831 570 -2829
rect 569 -2837 570 -2835
rect 576 -2831 577 -2829
rect 576 -2837 577 -2835
rect 583 -2831 584 -2829
rect 583 -2837 584 -2835
rect 586 -2837 587 -2835
rect 590 -2831 591 -2829
rect 590 -2837 591 -2835
rect 597 -2831 598 -2829
rect 597 -2837 598 -2835
rect 604 -2831 605 -2829
rect 604 -2837 605 -2835
rect 611 -2831 612 -2829
rect 611 -2837 612 -2835
rect 618 -2831 619 -2829
rect 621 -2831 622 -2829
rect 618 -2837 619 -2835
rect 621 -2837 622 -2835
rect 625 -2831 626 -2829
rect 625 -2837 626 -2835
rect 632 -2831 633 -2829
rect 632 -2837 633 -2835
rect 639 -2831 640 -2829
rect 639 -2837 640 -2835
rect 646 -2831 647 -2829
rect 646 -2837 647 -2835
rect 653 -2831 654 -2829
rect 653 -2837 654 -2835
rect 660 -2831 661 -2829
rect 663 -2831 664 -2829
rect 660 -2837 661 -2835
rect 663 -2837 664 -2835
rect 667 -2831 668 -2829
rect 667 -2837 668 -2835
rect 674 -2831 675 -2829
rect 674 -2837 675 -2835
rect 681 -2831 682 -2829
rect 681 -2837 682 -2835
rect 688 -2831 689 -2829
rect 688 -2837 689 -2835
rect 695 -2831 696 -2829
rect 695 -2837 696 -2835
rect 702 -2831 703 -2829
rect 705 -2831 706 -2829
rect 705 -2837 706 -2835
rect 709 -2831 710 -2829
rect 712 -2831 713 -2829
rect 712 -2837 713 -2835
rect 716 -2831 717 -2829
rect 716 -2837 717 -2835
rect 723 -2831 724 -2829
rect 723 -2837 724 -2835
rect 730 -2831 731 -2829
rect 733 -2831 734 -2829
rect 733 -2837 734 -2835
rect 737 -2831 738 -2829
rect 737 -2837 738 -2835
rect 744 -2831 745 -2829
rect 744 -2837 745 -2835
rect 751 -2831 752 -2829
rect 751 -2837 752 -2835
rect 758 -2831 759 -2829
rect 758 -2837 759 -2835
rect 765 -2831 766 -2829
rect 765 -2837 766 -2835
rect 772 -2831 773 -2829
rect 772 -2837 773 -2835
rect 779 -2831 780 -2829
rect 779 -2837 780 -2835
rect 786 -2831 787 -2829
rect 786 -2837 787 -2835
rect 793 -2831 794 -2829
rect 793 -2837 794 -2835
rect 800 -2831 801 -2829
rect 800 -2837 801 -2835
rect 807 -2831 808 -2829
rect 807 -2837 808 -2835
rect 814 -2831 815 -2829
rect 814 -2837 815 -2835
rect 821 -2831 822 -2829
rect 821 -2837 822 -2835
rect 831 -2831 832 -2829
rect 828 -2837 829 -2835
rect 835 -2831 836 -2829
rect 835 -2837 836 -2835
rect 842 -2831 843 -2829
rect 842 -2837 843 -2835
rect 849 -2831 850 -2829
rect 852 -2831 853 -2829
rect 849 -2837 850 -2835
rect 852 -2837 853 -2835
rect 856 -2831 857 -2829
rect 859 -2831 860 -2829
rect 856 -2837 857 -2835
rect 859 -2837 860 -2835
rect 863 -2831 864 -2829
rect 863 -2837 864 -2835
rect 870 -2837 871 -2835
rect 873 -2837 874 -2835
rect 877 -2831 878 -2829
rect 877 -2837 878 -2835
rect 884 -2831 885 -2829
rect 884 -2837 885 -2835
rect 891 -2831 892 -2829
rect 891 -2837 892 -2835
rect 898 -2831 899 -2829
rect 898 -2837 899 -2835
rect 905 -2831 906 -2829
rect 905 -2837 906 -2835
rect 912 -2831 913 -2829
rect 912 -2837 913 -2835
rect 919 -2831 920 -2829
rect 919 -2837 920 -2835
rect 926 -2831 927 -2829
rect 926 -2837 927 -2835
rect 933 -2831 934 -2829
rect 933 -2837 934 -2835
rect 940 -2831 941 -2829
rect 940 -2837 941 -2835
rect 947 -2831 948 -2829
rect 947 -2837 948 -2835
rect 954 -2831 955 -2829
rect 954 -2837 955 -2835
rect 961 -2831 962 -2829
rect 961 -2837 962 -2835
rect 968 -2831 969 -2829
rect 968 -2837 969 -2835
rect 975 -2831 976 -2829
rect 975 -2837 976 -2835
rect 982 -2831 983 -2829
rect 982 -2837 983 -2835
rect 989 -2831 990 -2829
rect 989 -2837 990 -2835
rect 996 -2831 997 -2829
rect 999 -2837 1000 -2835
rect 1003 -2831 1004 -2829
rect 1003 -2837 1004 -2835
rect 1010 -2831 1011 -2829
rect 1013 -2831 1014 -2829
rect 1010 -2837 1011 -2835
rect 1013 -2837 1014 -2835
rect 1017 -2831 1018 -2829
rect 1020 -2831 1021 -2829
rect 1020 -2837 1021 -2835
rect 1024 -2831 1025 -2829
rect 1024 -2837 1025 -2835
rect 1031 -2831 1032 -2829
rect 1031 -2837 1032 -2835
rect 1038 -2831 1039 -2829
rect 1038 -2837 1039 -2835
rect 1045 -2831 1046 -2829
rect 1045 -2837 1046 -2835
rect 1052 -2831 1053 -2829
rect 1052 -2837 1053 -2835
rect 1059 -2831 1060 -2829
rect 1059 -2837 1060 -2835
rect 1066 -2831 1067 -2829
rect 1069 -2831 1070 -2829
rect 1066 -2837 1067 -2835
rect 1069 -2837 1070 -2835
rect 1073 -2831 1074 -2829
rect 1073 -2837 1074 -2835
rect 1080 -2831 1081 -2829
rect 1080 -2837 1081 -2835
rect 1087 -2831 1088 -2829
rect 1087 -2837 1088 -2835
rect 1094 -2831 1095 -2829
rect 1094 -2837 1095 -2835
rect 1101 -2831 1102 -2829
rect 1101 -2837 1102 -2835
rect 1108 -2831 1109 -2829
rect 1108 -2837 1109 -2835
rect 1115 -2831 1116 -2829
rect 1118 -2831 1119 -2829
rect 1115 -2837 1116 -2835
rect 1125 -2831 1126 -2829
rect 1122 -2837 1123 -2835
rect 1125 -2837 1126 -2835
rect 1129 -2831 1130 -2829
rect 1129 -2837 1130 -2835
rect 1136 -2831 1137 -2829
rect 1136 -2837 1137 -2835
rect 1143 -2831 1144 -2829
rect 1143 -2837 1144 -2835
rect 1150 -2831 1151 -2829
rect 1150 -2837 1151 -2835
rect 1157 -2831 1158 -2829
rect 1157 -2837 1158 -2835
rect 1164 -2831 1165 -2829
rect 1164 -2837 1165 -2835
rect 1171 -2831 1172 -2829
rect 1171 -2837 1172 -2835
rect 1178 -2831 1179 -2829
rect 1181 -2831 1182 -2829
rect 1178 -2837 1179 -2835
rect 1185 -2831 1186 -2829
rect 1185 -2837 1186 -2835
rect 1192 -2831 1193 -2829
rect 1192 -2837 1193 -2835
rect 1199 -2831 1200 -2829
rect 1202 -2831 1203 -2829
rect 1199 -2837 1200 -2835
rect 1202 -2837 1203 -2835
rect 1206 -2831 1207 -2829
rect 1206 -2837 1207 -2835
rect 1213 -2831 1214 -2829
rect 1213 -2837 1214 -2835
rect 1220 -2831 1221 -2829
rect 1220 -2837 1221 -2835
rect 1227 -2831 1228 -2829
rect 1227 -2837 1228 -2835
rect 1237 -2831 1238 -2829
rect 1234 -2837 1235 -2835
rect 1237 -2837 1238 -2835
rect 1241 -2831 1242 -2829
rect 1241 -2837 1242 -2835
rect 1248 -2831 1249 -2829
rect 1248 -2837 1249 -2835
rect 1255 -2831 1256 -2829
rect 1255 -2837 1256 -2835
rect 1262 -2831 1263 -2829
rect 1262 -2837 1263 -2835
rect 1269 -2831 1270 -2829
rect 1269 -2837 1270 -2835
rect 1276 -2831 1277 -2829
rect 1276 -2837 1277 -2835
rect 1283 -2831 1284 -2829
rect 1283 -2837 1284 -2835
rect 1286 -2837 1287 -2835
rect 1290 -2831 1291 -2829
rect 1290 -2837 1291 -2835
rect 1297 -2831 1298 -2829
rect 1297 -2837 1298 -2835
rect 1304 -2831 1305 -2829
rect 1304 -2837 1305 -2835
rect 1311 -2831 1312 -2829
rect 1311 -2837 1312 -2835
rect 1318 -2831 1319 -2829
rect 1318 -2837 1319 -2835
rect 1325 -2831 1326 -2829
rect 1325 -2837 1326 -2835
rect 1332 -2831 1333 -2829
rect 1332 -2837 1333 -2835
rect 1342 -2831 1343 -2829
rect 1342 -2837 1343 -2835
rect 1346 -2831 1347 -2829
rect 1346 -2837 1347 -2835
rect 1353 -2831 1354 -2829
rect 1353 -2837 1354 -2835
rect 1356 -2837 1357 -2835
rect 1360 -2831 1361 -2829
rect 1360 -2837 1361 -2835
rect 1367 -2831 1368 -2829
rect 1367 -2837 1368 -2835
rect 1374 -2831 1375 -2829
rect 1374 -2837 1375 -2835
rect 1381 -2831 1382 -2829
rect 1381 -2837 1382 -2835
rect 1388 -2831 1389 -2829
rect 1388 -2837 1389 -2835
rect 1395 -2831 1396 -2829
rect 1395 -2837 1396 -2835
rect 1402 -2831 1403 -2829
rect 1402 -2837 1403 -2835
rect 1409 -2831 1410 -2829
rect 1409 -2837 1410 -2835
rect 1416 -2831 1417 -2829
rect 1416 -2837 1417 -2835
rect 1423 -2831 1424 -2829
rect 1423 -2837 1424 -2835
rect 1430 -2831 1431 -2829
rect 1433 -2831 1434 -2829
rect 1430 -2837 1431 -2835
rect 1433 -2837 1434 -2835
rect 1437 -2831 1438 -2829
rect 1437 -2837 1438 -2835
rect 1444 -2831 1445 -2829
rect 1444 -2837 1445 -2835
rect 1451 -2831 1452 -2829
rect 1451 -2837 1452 -2835
rect 1458 -2831 1459 -2829
rect 1458 -2837 1459 -2835
rect 1465 -2831 1466 -2829
rect 1465 -2837 1466 -2835
rect 1472 -2831 1473 -2829
rect 1472 -2837 1473 -2835
rect 1479 -2831 1480 -2829
rect 1479 -2837 1480 -2835
rect 1486 -2831 1487 -2829
rect 1486 -2837 1487 -2835
rect 1493 -2831 1494 -2829
rect 1493 -2837 1494 -2835
rect 1500 -2831 1501 -2829
rect 1500 -2837 1501 -2835
rect 1507 -2831 1508 -2829
rect 1507 -2837 1508 -2835
rect 1514 -2831 1515 -2829
rect 1514 -2837 1515 -2835
rect 1521 -2831 1522 -2829
rect 1521 -2837 1522 -2835
rect 1528 -2831 1529 -2829
rect 1528 -2837 1529 -2835
rect 1535 -2831 1536 -2829
rect 1535 -2837 1536 -2835
rect 1542 -2831 1543 -2829
rect 1542 -2837 1543 -2835
rect 1549 -2831 1550 -2829
rect 1549 -2837 1550 -2835
rect 1556 -2831 1557 -2829
rect 1556 -2837 1557 -2835
rect 1563 -2831 1564 -2829
rect 1563 -2837 1564 -2835
rect 1570 -2831 1571 -2829
rect 1570 -2837 1571 -2835
rect 1577 -2831 1578 -2829
rect 1577 -2837 1578 -2835
rect 1584 -2831 1585 -2829
rect 1584 -2837 1585 -2835
rect 1591 -2831 1592 -2829
rect 1591 -2837 1592 -2835
rect 1598 -2831 1599 -2829
rect 1598 -2837 1599 -2835
rect 1605 -2831 1606 -2829
rect 1605 -2837 1606 -2835
rect 1612 -2831 1613 -2829
rect 1612 -2837 1613 -2835
rect 1619 -2831 1620 -2829
rect 1619 -2837 1620 -2835
rect 1626 -2831 1627 -2829
rect 1626 -2837 1627 -2835
rect 1633 -2831 1634 -2829
rect 1633 -2837 1634 -2835
rect 1640 -2831 1641 -2829
rect 1640 -2837 1641 -2835
rect 1647 -2831 1648 -2829
rect 1647 -2837 1648 -2835
rect 1654 -2831 1655 -2829
rect 1654 -2837 1655 -2835
rect 1661 -2831 1662 -2829
rect 1661 -2837 1662 -2835
rect 1668 -2831 1669 -2829
rect 1668 -2837 1669 -2835
rect 1675 -2831 1676 -2829
rect 1675 -2837 1676 -2835
rect 1682 -2831 1683 -2829
rect 1682 -2837 1683 -2835
rect 1689 -2831 1690 -2829
rect 1689 -2837 1690 -2835
rect 1696 -2831 1697 -2829
rect 1696 -2837 1697 -2835
rect 1703 -2831 1704 -2829
rect 1703 -2837 1704 -2835
rect 1710 -2831 1711 -2829
rect 1713 -2831 1714 -2829
rect 1710 -2837 1711 -2835
rect 1713 -2837 1714 -2835
rect 1717 -2831 1718 -2829
rect 1720 -2831 1721 -2829
rect 1717 -2837 1718 -2835
rect 1720 -2837 1721 -2835
rect 1724 -2831 1725 -2829
rect 1724 -2837 1725 -2835
rect 1727 -2837 1728 -2835
rect 1731 -2831 1732 -2829
rect 1731 -2837 1732 -2835
rect 1738 -2831 1739 -2829
rect 1738 -2837 1739 -2835
rect 1745 -2831 1746 -2829
rect 1745 -2837 1746 -2835
rect 1752 -2831 1753 -2829
rect 1752 -2837 1753 -2835
rect 1759 -2831 1760 -2829
rect 1759 -2837 1760 -2835
rect 1766 -2831 1767 -2829
rect 1766 -2837 1767 -2835
rect 1773 -2831 1774 -2829
rect 1773 -2837 1774 -2835
rect 23 -2950 24 -2948
rect 23 -2956 24 -2954
rect 51 -2950 52 -2948
rect 51 -2956 52 -2954
rect 58 -2950 59 -2948
rect 58 -2956 59 -2954
rect 65 -2950 66 -2948
rect 65 -2956 66 -2954
rect 72 -2950 73 -2948
rect 72 -2956 73 -2954
rect 82 -2950 83 -2948
rect 79 -2956 80 -2954
rect 82 -2956 83 -2954
rect 86 -2950 87 -2948
rect 86 -2956 87 -2954
rect 93 -2950 94 -2948
rect 93 -2956 94 -2954
rect 100 -2950 101 -2948
rect 100 -2956 101 -2954
rect 107 -2950 108 -2948
rect 110 -2950 111 -2948
rect 107 -2956 108 -2954
rect 110 -2956 111 -2954
rect 114 -2950 115 -2948
rect 114 -2956 115 -2954
rect 121 -2950 122 -2948
rect 121 -2956 122 -2954
rect 128 -2950 129 -2948
rect 128 -2956 129 -2954
rect 135 -2956 136 -2954
rect 138 -2956 139 -2954
rect 142 -2950 143 -2948
rect 145 -2950 146 -2948
rect 142 -2956 143 -2954
rect 149 -2950 150 -2948
rect 149 -2956 150 -2954
rect 156 -2950 157 -2948
rect 156 -2956 157 -2954
rect 163 -2950 164 -2948
rect 166 -2950 167 -2948
rect 163 -2956 164 -2954
rect 170 -2950 171 -2948
rect 170 -2956 171 -2954
rect 177 -2950 178 -2948
rect 177 -2956 178 -2954
rect 184 -2950 185 -2948
rect 184 -2956 185 -2954
rect 191 -2950 192 -2948
rect 191 -2956 192 -2954
rect 198 -2950 199 -2948
rect 198 -2956 199 -2954
rect 205 -2950 206 -2948
rect 208 -2950 209 -2948
rect 205 -2956 206 -2954
rect 212 -2950 213 -2948
rect 212 -2956 213 -2954
rect 219 -2950 220 -2948
rect 219 -2956 220 -2954
rect 226 -2950 227 -2948
rect 229 -2950 230 -2948
rect 226 -2956 227 -2954
rect 233 -2950 234 -2948
rect 233 -2956 234 -2954
rect 240 -2950 241 -2948
rect 240 -2956 241 -2954
rect 247 -2950 248 -2948
rect 247 -2956 248 -2954
rect 254 -2950 255 -2948
rect 254 -2956 255 -2954
rect 261 -2950 262 -2948
rect 261 -2956 262 -2954
rect 268 -2950 269 -2948
rect 268 -2956 269 -2954
rect 275 -2950 276 -2948
rect 275 -2956 276 -2954
rect 282 -2950 283 -2948
rect 282 -2956 283 -2954
rect 289 -2950 290 -2948
rect 289 -2956 290 -2954
rect 296 -2950 297 -2948
rect 296 -2956 297 -2954
rect 303 -2950 304 -2948
rect 303 -2956 304 -2954
rect 310 -2950 311 -2948
rect 310 -2956 311 -2954
rect 317 -2950 318 -2948
rect 317 -2956 318 -2954
rect 324 -2950 325 -2948
rect 324 -2956 325 -2954
rect 331 -2950 332 -2948
rect 331 -2956 332 -2954
rect 338 -2950 339 -2948
rect 338 -2956 339 -2954
rect 345 -2950 346 -2948
rect 345 -2956 346 -2954
rect 352 -2950 353 -2948
rect 352 -2956 353 -2954
rect 359 -2950 360 -2948
rect 359 -2956 360 -2954
rect 366 -2950 367 -2948
rect 366 -2956 367 -2954
rect 373 -2950 374 -2948
rect 373 -2956 374 -2954
rect 380 -2950 381 -2948
rect 380 -2956 381 -2954
rect 387 -2950 388 -2948
rect 387 -2956 388 -2954
rect 394 -2950 395 -2948
rect 394 -2956 395 -2954
rect 401 -2950 402 -2948
rect 401 -2956 402 -2954
rect 411 -2950 412 -2948
rect 408 -2956 409 -2954
rect 411 -2956 412 -2954
rect 415 -2950 416 -2948
rect 415 -2956 416 -2954
rect 422 -2950 423 -2948
rect 422 -2956 423 -2954
rect 429 -2950 430 -2948
rect 429 -2956 430 -2954
rect 436 -2950 437 -2948
rect 439 -2950 440 -2948
rect 439 -2956 440 -2954
rect 443 -2950 444 -2948
rect 443 -2956 444 -2954
rect 450 -2950 451 -2948
rect 450 -2956 451 -2954
rect 457 -2950 458 -2948
rect 457 -2956 458 -2954
rect 464 -2950 465 -2948
rect 467 -2950 468 -2948
rect 464 -2956 465 -2954
rect 471 -2950 472 -2948
rect 471 -2956 472 -2954
rect 478 -2950 479 -2948
rect 478 -2956 479 -2954
rect 485 -2950 486 -2948
rect 485 -2956 486 -2954
rect 492 -2950 493 -2948
rect 492 -2956 493 -2954
rect 499 -2950 500 -2948
rect 499 -2956 500 -2954
rect 506 -2950 507 -2948
rect 506 -2956 507 -2954
rect 513 -2950 514 -2948
rect 513 -2956 514 -2954
rect 520 -2950 521 -2948
rect 520 -2956 521 -2954
rect 527 -2950 528 -2948
rect 527 -2956 528 -2954
rect 534 -2950 535 -2948
rect 537 -2950 538 -2948
rect 534 -2956 535 -2954
rect 537 -2956 538 -2954
rect 541 -2950 542 -2948
rect 541 -2956 542 -2954
rect 548 -2950 549 -2948
rect 548 -2956 549 -2954
rect 555 -2950 556 -2948
rect 555 -2956 556 -2954
rect 562 -2950 563 -2948
rect 562 -2956 563 -2954
rect 569 -2950 570 -2948
rect 569 -2956 570 -2954
rect 576 -2950 577 -2948
rect 576 -2956 577 -2954
rect 583 -2950 584 -2948
rect 583 -2956 584 -2954
rect 590 -2950 591 -2948
rect 590 -2956 591 -2954
rect 597 -2950 598 -2948
rect 597 -2956 598 -2954
rect 604 -2950 605 -2948
rect 604 -2956 605 -2954
rect 611 -2950 612 -2948
rect 611 -2956 612 -2954
rect 618 -2950 619 -2948
rect 618 -2956 619 -2954
rect 625 -2950 626 -2948
rect 625 -2956 626 -2954
rect 632 -2950 633 -2948
rect 632 -2956 633 -2954
rect 639 -2950 640 -2948
rect 639 -2956 640 -2954
rect 646 -2950 647 -2948
rect 646 -2956 647 -2954
rect 653 -2950 654 -2948
rect 656 -2950 657 -2948
rect 653 -2956 654 -2954
rect 656 -2956 657 -2954
rect 660 -2950 661 -2948
rect 663 -2950 664 -2948
rect 660 -2956 661 -2954
rect 663 -2956 664 -2954
rect 667 -2950 668 -2948
rect 667 -2956 668 -2954
rect 674 -2950 675 -2948
rect 674 -2956 675 -2954
rect 681 -2950 682 -2948
rect 681 -2956 682 -2954
rect 688 -2950 689 -2948
rect 688 -2956 689 -2954
rect 695 -2950 696 -2948
rect 695 -2956 696 -2954
rect 702 -2950 703 -2948
rect 702 -2956 703 -2954
rect 709 -2950 710 -2948
rect 709 -2956 710 -2954
rect 716 -2950 717 -2948
rect 716 -2956 717 -2954
rect 723 -2950 724 -2948
rect 723 -2956 724 -2954
rect 730 -2950 731 -2948
rect 730 -2956 731 -2954
rect 737 -2950 738 -2948
rect 737 -2956 738 -2954
rect 744 -2950 745 -2948
rect 744 -2956 745 -2954
rect 751 -2950 752 -2948
rect 751 -2956 752 -2954
rect 758 -2950 759 -2948
rect 758 -2956 759 -2954
rect 765 -2950 766 -2948
rect 765 -2956 766 -2954
rect 772 -2950 773 -2948
rect 772 -2956 773 -2954
rect 782 -2950 783 -2948
rect 779 -2956 780 -2954
rect 782 -2956 783 -2954
rect 786 -2950 787 -2948
rect 786 -2956 787 -2954
rect 793 -2950 794 -2948
rect 793 -2956 794 -2954
rect 800 -2950 801 -2948
rect 800 -2956 801 -2954
rect 807 -2950 808 -2948
rect 807 -2956 808 -2954
rect 814 -2950 815 -2948
rect 814 -2956 815 -2954
rect 824 -2950 825 -2948
rect 828 -2950 829 -2948
rect 828 -2956 829 -2954
rect 835 -2950 836 -2948
rect 835 -2956 836 -2954
rect 842 -2950 843 -2948
rect 842 -2956 843 -2954
rect 849 -2950 850 -2948
rect 852 -2950 853 -2948
rect 849 -2956 850 -2954
rect 852 -2956 853 -2954
rect 856 -2950 857 -2948
rect 856 -2956 857 -2954
rect 863 -2950 864 -2948
rect 866 -2950 867 -2948
rect 863 -2956 864 -2954
rect 866 -2956 867 -2954
rect 870 -2950 871 -2948
rect 870 -2956 871 -2954
rect 877 -2950 878 -2948
rect 877 -2956 878 -2954
rect 884 -2950 885 -2948
rect 884 -2956 885 -2954
rect 891 -2950 892 -2948
rect 891 -2956 892 -2954
rect 898 -2950 899 -2948
rect 898 -2956 899 -2954
rect 905 -2950 906 -2948
rect 905 -2956 906 -2954
rect 912 -2950 913 -2948
rect 915 -2950 916 -2948
rect 912 -2956 913 -2954
rect 915 -2956 916 -2954
rect 919 -2950 920 -2948
rect 919 -2956 920 -2954
rect 926 -2950 927 -2948
rect 926 -2956 927 -2954
rect 933 -2950 934 -2948
rect 933 -2956 934 -2954
rect 943 -2950 944 -2948
rect 940 -2956 941 -2954
rect 943 -2956 944 -2954
rect 947 -2950 948 -2948
rect 947 -2956 948 -2954
rect 954 -2950 955 -2948
rect 954 -2956 955 -2954
rect 961 -2950 962 -2948
rect 961 -2956 962 -2954
rect 968 -2950 969 -2948
rect 971 -2950 972 -2948
rect 968 -2956 969 -2954
rect 975 -2950 976 -2948
rect 975 -2956 976 -2954
rect 982 -2950 983 -2948
rect 982 -2956 983 -2954
rect 989 -2950 990 -2948
rect 989 -2956 990 -2954
rect 996 -2950 997 -2948
rect 996 -2956 997 -2954
rect 1003 -2950 1004 -2948
rect 1003 -2956 1004 -2954
rect 1010 -2950 1011 -2948
rect 1010 -2956 1011 -2954
rect 1017 -2950 1018 -2948
rect 1017 -2956 1018 -2954
rect 1024 -2950 1025 -2948
rect 1027 -2950 1028 -2948
rect 1024 -2956 1025 -2954
rect 1027 -2956 1028 -2954
rect 1031 -2950 1032 -2948
rect 1031 -2956 1032 -2954
rect 1034 -2956 1035 -2954
rect 1038 -2950 1039 -2948
rect 1038 -2956 1039 -2954
rect 1045 -2950 1046 -2948
rect 1045 -2956 1046 -2954
rect 1052 -2950 1053 -2948
rect 1055 -2950 1056 -2948
rect 1055 -2956 1056 -2954
rect 1059 -2950 1060 -2948
rect 1059 -2956 1060 -2954
rect 1066 -2950 1067 -2948
rect 1066 -2956 1067 -2954
rect 1073 -2950 1074 -2948
rect 1073 -2956 1074 -2954
rect 1080 -2950 1081 -2948
rect 1080 -2956 1081 -2954
rect 1087 -2950 1088 -2948
rect 1087 -2956 1088 -2954
rect 1097 -2950 1098 -2948
rect 1097 -2956 1098 -2954
rect 1101 -2950 1102 -2948
rect 1101 -2956 1102 -2954
rect 1108 -2950 1109 -2948
rect 1108 -2956 1109 -2954
rect 1115 -2950 1116 -2948
rect 1115 -2956 1116 -2954
rect 1122 -2950 1123 -2948
rect 1122 -2956 1123 -2954
rect 1129 -2950 1130 -2948
rect 1129 -2956 1130 -2954
rect 1136 -2950 1137 -2948
rect 1136 -2956 1137 -2954
rect 1143 -2950 1144 -2948
rect 1143 -2956 1144 -2954
rect 1150 -2950 1151 -2948
rect 1150 -2956 1151 -2954
rect 1157 -2950 1158 -2948
rect 1157 -2956 1158 -2954
rect 1164 -2950 1165 -2948
rect 1164 -2956 1165 -2954
rect 1171 -2950 1172 -2948
rect 1171 -2956 1172 -2954
rect 1178 -2950 1179 -2948
rect 1178 -2956 1179 -2954
rect 1185 -2950 1186 -2948
rect 1185 -2956 1186 -2954
rect 1192 -2950 1193 -2948
rect 1192 -2956 1193 -2954
rect 1202 -2950 1203 -2948
rect 1199 -2956 1200 -2954
rect 1202 -2956 1203 -2954
rect 1206 -2950 1207 -2948
rect 1206 -2956 1207 -2954
rect 1213 -2950 1214 -2948
rect 1213 -2956 1214 -2954
rect 1220 -2950 1221 -2948
rect 1220 -2956 1221 -2954
rect 1227 -2950 1228 -2948
rect 1227 -2956 1228 -2954
rect 1234 -2950 1235 -2948
rect 1234 -2956 1235 -2954
rect 1241 -2950 1242 -2948
rect 1241 -2956 1242 -2954
rect 1248 -2950 1249 -2948
rect 1248 -2956 1249 -2954
rect 1255 -2950 1256 -2948
rect 1255 -2956 1256 -2954
rect 1262 -2950 1263 -2948
rect 1262 -2956 1263 -2954
rect 1269 -2950 1270 -2948
rect 1269 -2956 1270 -2954
rect 1276 -2950 1277 -2948
rect 1276 -2956 1277 -2954
rect 1283 -2950 1284 -2948
rect 1283 -2956 1284 -2954
rect 1290 -2950 1291 -2948
rect 1290 -2956 1291 -2954
rect 1297 -2950 1298 -2948
rect 1297 -2956 1298 -2954
rect 1304 -2950 1305 -2948
rect 1304 -2956 1305 -2954
rect 1311 -2950 1312 -2948
rect 1311 -2956 1312 -2954
rect 1318 -2950 1319 -2948
rect 1318 -2956 1319 -2954
rect 1325 -2950 1326 -2948
rect 1325 -2956 1326 -2954
rect 1332 -2956 1333 -2954
rect 1335 -2956 1336 -2954
rect 1339 -2950 1340 -2948
rect 1339 -2956 1340 -2954
rect 1346 -2950 1347 -2948
rect 1346 -2956 1347 -2954
rect 1353 -2950 1354 -2948
rect 1353 -2956 1354 -2954
rect 1360 -2950 1361 -2948
rect 1360 -2956 1361 -2954
rect 1367 -2950 1368 -2948
rect 1367 -2956 1368 -2954
rect 1374 -2950 1375 -2948
rect 1374 -2956 1375 -2954
rect 1381 -2950 1382 -2948
rect 1381 -2956 1382 -2954
rect 1388 -2950 1389 -2948
rect 1388 -2956 1389 -2954
rect 1395 -2950 1396 -2948
rect 1395 -2956 1396 -2954
rect 1402 -2950 1403 -2948
rect 1402 -2956 1403 -2954
rect 1409 -2950 1410 -2948
rect 1409 -2956 1410 -2954
rect 1416 -2950 1417 -2948
rect 1416 -2956 1417 -2954
rect 1423 -2950 1424 -2948
rect 1423 -2956 1424 -2954
rect 1430 -2950 1431 -2948
rect 1430 -2956 1431 -2954
rect 1437 -2950 1438 -2948
rect 1437 -2956 1438 -2954
rect 1444 -2950 1445 -2948
rect 1444 -2956 1445 -2954
rect 1451 -2950 1452 -2948
rect 1451 -2956 1452 -2954
rect 1458 -2950 1459 -2948
rect 1458 -2956 1459 -2954
rect 1465 -2950 1466 -2948
rect 1465 -2956 1466 -2954
rect 1472 -2950 1473 -2948
rect 1472 -2956 1473 -2954
rect 1479 -2950 1480 -2948
rect 1479 -2956 1480 -2954
rect 1486 -2950 1487 -2948
rect 1486 -2956 1487 -2954
rect 1493 -2950 1494 -2948
rect 1493 -2956 1494 -2954
rect 1500 -2950 1501 -2948
rect 1500 -2956 1501 -2954
rect 1507 -2950 1508 -2948
rect 1507 -2956 1508 -2954
rect 1514 -2950 1515 -2948
rect 1514 -2956 1515 -2954
rect 1521 -2950 1522 -2948
rect 1521 -2956 1522 -2954
rect 1528 -2950 1529 -2948
rect 1528 -2956 1529 -2954
rect 1535 -2950 1536 -2948
rect 1535 -2956 1536 -2954
rect 1542 -2950 1543 -2948
rect 1542 -2956 1543 -2954
rect 1549 -2950 1550 -2948
rect 1549 -2956 1550 -2954
rect 1556 -2950 1557 -2948
rect 1556 -2956 1557 -2954
rect 1563 -2950 1564 -2948
rect 1563 -2956 1564 -2954
rect 1570 -2950 1571 -2948
rect 1570 -2956 1571 -2954
rect 1577 -2950 1578 -2948
rect 1577 -2956 1578 -2954
rect 1584 -2950 1585 -2948
rect 1584 -2956 1585 -2954
rect 1591 -2950 1592 -2948
rect 1591 -2956 1592 -2954
rect 1598 -2950 1599 -2948
rect 1598 -2956 1599 -2954
rect 1605 -2950 1606 -2948
rect 1605 -2956 1606 -2954
rect 1612 -2950 1613 -2948
rect 1612 -2956 1613 -2954
rect 1619 -2950 1620 -2948
rect 1619 -2956 1620 -2954
rect 1626 -2950 1627 -2948
rect 1626 -2956 1627 -2954
rect 1633 -2950 1634 -2948
rect 1633 -2956 1634 -2954
rect 1640 -2950 1641 -2948
rect 1640 -2956 1641 -2954
rect 1647 -2950 1648 -2948
rect 1647 -2956 1648 -2954
rect 1654 -2950 1655 -2948
rect 1654 -2956 1655 -2954
rect 1661 -2950 1662 -2948
rect 1661 -2956 1662 -2954
rect 1668 -2950 1669 -2948
rect 1668 -2956 1669 -2954
rect 1675 -2950 1676 -2948
rect 1675 -2956 1676 -2954
rect 1682 -2950 1683 -2948
rect 1682 -2956 1683 -2954
rect 1689 -2950 1690 -2948
rect 1689 -2956 1690 -2954
rect 1696 -2950 1697 -2948
rect 1696 -2956 1697 -2954
rect 1703 -2950 1704 -2948
rect 1703 -2956 1704 -2954
rect 1706 -2956 1707 -2954
rect 30 -3077 31 -3075
rect 30 -3083 31 -3081
rect 37 -3077 38 -3075
rect 37 -3083 38 -3081
rect 44 -3077 45 -3075
rect 44 -3083 45 -3081
rect 51 -3077 52 -3075
rect 51 -3083 52 -3081
rect 58 -3077 59 -3075
rect 61 -3077 62 -3075
rect 61 -3083 62 -3081
rect 65 -3077 66 -3075
rect 65 -3083 66 -3081
rect 72 -3077 73 -3075
rect 72 -3083 73 -3081
rect 79 -3077 80 -3075
rect 82 -3077 83 -3075
rect 79 -3083 80 -3081
rect 82 -3083 83 -3081
rect 86 -3077 87 -3075
rect 89 -3077 90 -3075
rect 86 -3083 87 -3081
rect 89 -3083 90 -3081
rect 93 -3077 94 -3075
rect 93 -3083 94 -3081
rect 100 -3077 101 -3075
rect 100 -3083 101 -3081
rect 107 -3077 108 -3075
rect 107 -3083 108 -3081
rect 114 -3077 115 -3075
rect 114 -3083 115 -3081
rect 121 -3077 122 -3075
rect 121 -3083 122 -3081
rect 128 -3077 129 -3075
rect 128 -3083 129 -3081
rect 135 -3083 136 -3081
rect 145 -3077 146 -3075
rect 142 -3083 143 -3081
rect 145 -3083 146 -3081
rect 149 -3077 150 -3075
rect 152 -3077 153 -3075
rect 149 -3083 150 -3081
rect 152 -3083 153 -3081
rect 156 -3077 157 -3075
rect 156 -3083 157 -3081
rect 163 -3077 164 -3075
rect 163 -3083 164 -3081
rect 170 -3077 171 -3075
rect 170 -3083 171 -3081
rect 177 -3077 178 -3075
rect 177 -3083 178 -3081
rect 184 -3077 185 -3075
rect 187 -3077 188 -3075
rect 184 -3083 185 -3081
rect 191 -3077 192 -3075
rect 191 -3083 192 -3081
rect 198 -3083 199 -3081
rect 201 -3083 202 -3081
rect 205 -3077 206 -3075
rect 208 -3077 209 -3075
rect 215 -3083 216 -3081
rect 219 -3077 220 -3075
rect 219 -3083 220 -3081
rect 226 -3077 227 -3075
rect 226 -3083 227 -3081
rect 233 -3077 234 -3075
rect 233 -3083 234 -3081
rect 240 -3077 241 -3075
rect 240 -3083 241 -3081
rect 247 -3077 248 -3075
rect 247 -3083 248 -3081
rect 254 -3077 255 -3075
rect 254 -3083 255 -3081
rect 261 -3077 262 -3075
rect 261 -3083 262 -3081
rect 268 -3077 269 -3075
rect 268 -3083 269 -3081
rect 275 -3077 276 -3075
rect 275 -3083 276 -3081
rect 282 -3077 283 -3075
rect 282 -3083 283 -3081
rect 289 -3077 290 -3075
rect 289 -3083 290 -3081
rect 296 -3077 297 -3075
rect 296 -3083 297 -3081
rect 303 -3077 304 -3075
rect 303 -3083 304 -3081
rect 310 -3077 311 -3075
rect 310 -3083 311 -3081
rect 317 -3077 318 -3075
rect 317 -3083 318 -3081
rect 324 -3077 325 -3075
rect 324 -3083 325 -3081
rect 331 -3077 332 -3075
rect 331 -3083 332 -3081
rect 338 -3077 339 -3075
rect 338 -3083 339 -3081
rect 345 -3077 346 -3075
rect 348 -3083 349 -3081
rect 352 -3077 353 -3075
rect 352 -3083 353 -3081
rect 359 -3077 360 -3075
rect 359 -3083 360 -3081
rect 366 -3077 367 -3075
rect 369 -3077 370 -3075
rect 366 -3083 367 -3081
rect 369 -3083 370 -3081
rect 373 -3077 374 -3075
rect 373 -3083 374 -3081
rect 380 -3077 381 -3075
rect 380 -3083 381 -3081
rect 387 -3077 388 -3075
rect 387 -3083 388 -3081
rect 394 -3077 395 -3075
rect 394 -3083 395 -3081
rect 401 -3077 402 -3075
rect 401 -3083 402 -3081
rect 408 -3077 409 -3075
rect 408 -3083 409 -3081
rect 415 -3077 416 -3075
rect 415 -3083 416 -3081
rect 422 -3077 423 -3075
rect 422 -3083 423 -3081
rect 429 -3077 430 -3075
rect 429 -3083 430 -3081
rect 436 -3077 437 -3075
rect 436 -3083 437 -3081
rect 443 -3077 444 -3075
rect 443 -3083 444 -3081
rect 450 -3077 451 -3075
rect 453 -3077 454 -3075
rect 450 -3083 451 -3081
rect 453 -3083 454 -3081
rect 457 -3077 458 -3075
rect 457 -3083 458 -3081
rect 464 -3077 465 -3075
rect 464 -3083 465 -3081
rect 471 -3077 472 -3075
rect 471 -3083 472 -3081
rect 478 -3077 479 -3075
rect 478 -3083 479 -3081
rect 485 -3077 486 -3075
rect 485 -3083 486 -3081
rect 492 -3077 493 -3075
rect 492 -3083 493 -3081
rect 499 -3077 500 -3075
rect 499 -3083 500 -3081
rect 506 -3077 507 -3075
rect 506 -3083 507 -3081
rect 513 -3077 514 -3075
rect 513 -3083 514 -3081
rect 520 -3077 521 -3075
rect 520 -3083 521 -3081
rect 527 -3077 528 -3075
rect 527 -3083 528 -3081
rect 534 -3077 535 -3075
rect 534 -3083 535 -3081
rect 541 -3077 542 -3075
rect 541 -3083 542 -3081
rect 548 -3077 549 -3075
rect 548 -3083 549 -3081
rect 555 -3077 556 -3075
rect 555 -3083 556 -3081
rect 562 -3077 563 -3075
rect 562 -3083 563 -3081
rect 569 -3077 570 -3075
rect 569 -3083 570 -3081
rect 576 -3077 577 -3075
rect 576 -3083 577 -3081
rect 583 -3077 584 -3075
rect 583 -3083 584 -3081
rect 590 -3077 591 -3075
rect 590 -3083 591 -3081
rect 597 -3077 598 -3075
rect 597 -3083 598 -3081
rect 604 -3077 605 -3075
rect 604 -3083 605 -3081
rect 611 -3077 612 -3075
rect 611 -3083 612 -3081
rect 618 -3077 619 -3075
rect 621 -3077 622 -3075
rect 621 -3083 622 -3081
rect 625 -3077 626 -3075
rect 625 -3083 626 -3081
rect 632 -3077 633 -3075
rect 635 -3077 636 -3075
rect 632 -3083 633 -3081
rect 635 -3083 636 -3081
rect 639 -3077 640 -3075
rect 639 -3083 640 -3081
rect 646 -3077 647 -3075
rect 646 -3083 647 -3081
rect 653 -3077 654 -3075
rect 653 -3083 654 -3081
rect 660 -3077 661 -3075
rect 660 -3083 661 -3081
rect 667 -3077 668 -3075
rect 667 -3083 668 -3081
rect 674 -3077 675 -3075
rect 674 -3083 675 -3081
rect 681 -3077 682 -3075
rect 681 -3083 682 -3081
rect 688 -3077 689 -3075
rect 691 -3077 692 -3075
rect 688 -3083 689 -3081
rect 691 -3083 692 -3081
rect 695 -3077 696 -3075
rect 695 -3083 696 -3081
rect 702 -3077 703 -3075
rect 702 -3083 703 -3081
rect 709 -3077 710 -3075
rect 709 -3083 710 -3081
rect 716 -3077 717 -3075
rect 716 -3083 717 -3081
rect 723 -3077 724 -3075
rect 723 -3083 724 -3081
rect 730 -3077 731 -3075
rect 730 -3083 731 -3081
rect 737 -3077 738 -3075
rect 740 -3077 741 -3075
rect 737 -3083 738 -3081
rect 740 -3083 741 -3081
rect 744 -3077 745 -3075
rect 744 -3083 745 -3081
rect 751 -3077 752 -3075
rect 751 -3083 752 -3081
rect 758 -3077 759 -3075
rect 761 -3083 762 -3081
rect 765 -3077 766 -3075
rect 765 -3083 766 -3081
rect 772 -3077 773 -3075
rect 772 -3083 773 -3081
rect 779 -3077 780 -3075
rect 779 -3083 780 -3081
rect 786 -3077 787 -3075
rect 789 -3077 790 -3075
rect 786 -3083 787 -3081
rect 789 -3083 790 -3081
rect 793 -3077 794 -3075
rect 793 -3083 794 -3081
rect 800 -3077 801 -3075
rect 800 -3083 801 -3081
rect 803 -3083 804 -3081
rect 807 -3077 808 -3075
rect 807 -3083 808 -3081
rect 814 -3077 815 -3075
rect 814 -3083 815 -3081
rect 821 -3077 822 -3075
rect 821 -3083 822 -3081
rect 828 -3077 829 -3075
rect 831 -3077 832 -3075
rect 828 -3083 829 -3081
rect 835 -3077 836 -3075
rect 835 -3083 836 -3081
rect 838 -3083 839 -3081
rect 842 -3077 843 -3075
rect 842 -3083 843 -3081
rect 849 -3077 850 -3075
rect 849 -3083 850 -3081
rect 856 -3077 857 -3075
rect 856 -3083 857 -3081
rect 863 -3077 864 -3075
rect 863 -3083 864 -3081
rect 870 -3077 871 -3075
rect 870 -3083 871 -3081
rect 877 -3077 878 -3075
rect 880 -3077 881 -3075
rect 877 -3083 878 -3081
rect 884 -3077 885 -3075
rect 884 -3083 885 -3081
rect 891 -3077 892 -3075
rect 891 -3083 892 -3081
rect 898 -3077 899 -3075
rect 901 -3077 902 -3075
rect 898 -3083 899 -3081
rect 905 -3077 906 -3075
rect 905 -3083 906 -3081
rect 915 -3077 916 -3075
rect 912 -3083 913 -3081
rect 915 -3083 916 -3081
rect 919 -3077 920 -3075
rect 919 -3083 920 -3081
rect 926 -3077 927 -3075
rect 926 -3083 927 -3081
rect 933 -3077 934 -3075
rect 933 -3083 934 -3081
rect 940 -3077 941 -3075
rect 940 -3083 941 -3081
rect 947 -3077 948 -3075
rect 947 -3083 948 -3081
rect 950 -3083 951 -3081
rect 954 -3077 955 -3075
rect 954 -3083 955 -3081
rect 961 -3077 962 -3075
rect 961 -3083 962 -3081
rect 968 -3077 969 -3075
rect 968 -3083 969 -3081
rect 978 -3077 979 -3075
rect 975 -3083 976 -3081
rect 978 -3083 979 -3081
rect 982 -3077 983 -3075
rect 982 -3083 983 -3081
rect 989 -3077 990 -3075
rect 989 -3083 990 -3081
rect 996 -3077 997 -3075
rect 996 -3083 997 -3081
rect 1003 -3077 1004 -3075
rect 1003 -3083 1004 -3081
rect 1010 -3077 1011 -3075
rect 1010 -3083 1011 -3081
rect 1017 -3077 1018 -3075
rect 1020 -3077 1021 -3075
rect 1017 -3083 1018 -3081
rect 1020 -3083 1021 -3081
rect 1024 -3077 1025 -3075
rect 1024 -3083 1025 -3081
rect 1031 -3077 1032 -3075
rect 1031 -3083 1032 -3081
rect 1038 -3077 1039 -3075
rect 1038 -3083 1039 -3081
rect 1045 -3077 1046 -3075
rect 1045 -3083 1046 -3081
rect 1052 -3077 1053 -3075
rect 1052 -3083 1053 -3081
rect 1059 -3077 1060 -3075
rect 1059 -3083 1060 -3081
rect 1066 -3077 1067 -3075
rect 1066 -3083 1067 -3081
rect 1073 -3077 1074 -3075
rect 1073 -3083 1074 -3081
rect 1080 -3077 1081 -3075
rect 1080 -3083 1081 -3081
rect 1083 -3083 1084 -3081
rect 1087 -3083 1088 -3081
rect 1090 -3083 1091 -3081
rect 1094 -3077 1095 -3075
rect 1094 -3083 1095 -3081
rect 1101 -3077 1102 -3075
rect 1101 -3083 1102 -3081
rect 1108 -3077 1109 -3075
rect 1108 -3083 1109 -3081
rect 1115 -3077 1116 -3075
rect 1115 -3083 1116 -3081
rect 1122 -3077 1123 -3075
rect 1122 -3083 1123 -3081
rect 1129 -3077 1130 -3075
rect 1129 -3083 1130 -3081
rect 1136 -3077 1137 -3075
rect 1136 -3083 1137 -3081
rect 1143 -3077 1144 -3075
rect 1143 -3083 1144 -3081
rect 1150 -3077 1151 -3075
rect 1150 -3083 1151 -3081
rect 1157 -3077 1158 -3075
rect 1157 -3083 1158 -3081
rect 1164 -3077 1165 -3075
rect 1164 -3083 1165 -3081
rect 1171 -3077 1172 -3075
rect 1171 -3083 1172 -3081
rect 1178 -3077 1179 -3075
rect 1178 -3083 1179 -3081
rect 1185 -3077 1186 -3075
rect 1185 -3083 1186 -3081
rect 1192 -3077 1193 -3075
rect 1192 -3083 1193 -3081
rect 1199 -3077 1200 -3075
rect 1199 -3083 1200 -3081
rect 1206 -3077 1207 -3075
rect 1206 -3083 1207 -3081
rect 1213 -3077 1214 -3075
rect 1213 -3083 1214 -3081
rect 1220 -3077 1221 -3075
rect 1220 -3083 1221 -3081
rect 1227 -3077 1228 -3075
rect 1227 -3083 1228 -3081
rect 1234 -3077 1235 -3075
rect 1234 -3083 1235 -3081
rect 1241 -3077 1242 -3075
rect 1241 -3083 1242 -3081
rect 1248 -3077 1249 -3075
rect 1248 -3083 1249 -3081
rect 1255 -3077 1256 -3075
rect 1255 -3083 1256 -3081
rect 1262 -3077 1263 -3075
rect 1262 -3083 1263 -3081
rect 1269 -3077 1270 -3075
rect 1269 -3083 1270 -3081
rect 1276 -3077 1277 -3075
rect 1276 -3083 1277 -3081
rect 1283 -3077 1284 -3075
rect 1283 -3083 1284 -3081
rect 1290 -3077 1291 -3075
rect 1290 -3083 1291 -3081
rect 1297 -3077 1298 -3075
rect 1297 -3083 1298 -3081
rect 1304 -3077 1305 -3075
rect 1304 -3083 1305 -3081
rect 1311 -3077 1312 -3075
rect 1311 -3083 1312 -3081
rect 1318 -3077 1319 -3075
rect 1318 -3083 1319 -3081
rect 1325 -3077 1326 -3075
rect 1325 -3083 1326 -3081
rect 1332 -3077 1333 -3075
rect 1332 -3083 1333 -3081
rect 1339 -3077 1340 -3075
rect 1339 -3083 1340 -3081
rect 1346 -3077 1347 -3075
rect 1346 -3083 1347 -3081
rect 1353 -3077 1354 -3075
rect 1353 -3083 1354 -3081
rect 1360 -3077 1361 -3075
rect 1360 -3083 1361 -3081
rect 1367 -3077 1368 -3075
rect 1367 -3083 1368 -3081
rect 1374 -3077 1375 -3075
rect 1374 -3083 1375 -3081
rect 1381 -3077 1382 -3075
rect 1381 -3083 1382 -3081
rect 1388 -3077 1389 -3075
rect 1388 -3083 1389 -3081
rect 1395 -3077 1396 -3075
rect 1395 -3083 1396 -3081
rect 1402 -3077 1403 -3075
rect 1402 -3083 1403 -3081
rect 1409 -3077 1410 -3075
rect 1409 -3083 1410 -3081
rect 1416 -3077 1417 -3075
rect 1416 -3083 1417 -3081
rect 1423 -3077 1424 -3075
rect 1423 -3083 1424 -3081
rect 1430 -3077 1431 -3075
rect 1430 -3083 1431 -3081
rect 1437 -3077 1438 -3075
rect 1437 -3083 1438 -3081
rect 1444 -3077 1445 -3075
rect 1444 -3083 1445 -3081
rect 1451 -3077 1452 -3075
rect 1451 -3083 1452 -3081
rect 1458 -3077 1459 -3075
rect 1458 -3083 1459 -3081
rect 1465 -3077 1466 -3075
rect 1465 -3083 1466 -3081
rect 1472 -3077 1473 -3075
rect 1472 -3083 1473 -3081
rect 1479 -3077 1480 -3075
rect 1479 -3083 1480 -3081
rect 1486 -3077 1487 -3075
rect 1486 -3083 1487 -3081
rect 1493 -3077 1494 -3075
rect 1493 -3083 1494 -3081
rect 1500 -3077 1501 -3075
rect 1500 -3083 1501 -3081
rect 1507 -3077 1508 -3075
rect 1507 -3083 1508 -3081
rect 1514 -3077 1515 -3075
rect 1514 -3083 1515 -3081
rect 1521 -3077 1522 -3075
rect 1521 -3083 1522 -3081
rect 1528 -3077 1529 -3075
rect 1528 -3083 1529 -3081
rect 1535 -3077 1536 -3075
rect 1535 -3083 1536 -3081
rect 1542 -3077 1543 -3075
rect 1542 -3083 1543 -3081
rect 1549 -3077 1550 -3075
rect 1549 -3083 1550 -3081
rect 1556 -3077 1557 -3075
rect 1556 -3083 1557 -3081
rect 1563 -3077 1564 -3075
rect 1563 -3083 1564 -3081
rect 1570 -3077 1571 -3075
rect 1570 -3083 1571 -3081
rect 1577 -3077 1578 -3075
rect 1577 -3083 1578 -3081
rect 1584 -3077 1585 -3075
rect 1584 -3083 1585 -3081
rect 1591 -3077 1592 -3075
rect 1591 -3083 1592 -3081
rect 1598 -3077 1599 -3075
rect 1598 -3083 1599 -3081
rect 1605 -3077 1606 -3075
rect 1605 -3083 1606 -3081
rect 1612 -3077 1613 -3075
rect 1612 -3083 1613 -3081
rect 1619 -3077 1620 -3075
rect 1619 -3083 1620 -3081
rect 1626 -3077 1627 -3075
rect 1626 -3083 1627 -3081
rect 1633 -3077 1634 -3075
rect 1633 -3083 1634 -3081
rect 1640 -3077 1641 -3075
rect 1640 -3083 1641 -3081
rect 1647 -3077 1648 -3075
rect 1647 -3083 1648 -3081
rect 1654 -3077 1655 -3075
rect 1654 -3083 1655 -3081
rect 65 -3222 66 -3220
rect 72 -3216 73 -3214
rect 72 -3222 73 -3220
rect 79 -3216 80 -3214
rect 79 -3222 80 -3220
rect 86 -3216 87 -3214
rect 86 -3222 87 -3220
rect 93 -3216 94 -3214
rect 93 -3222 94 -3220
rect 100 -3216 101 -3214
rect 100 -3222 101 -3220
rect 107 -3216 108 -3214
rect 107 -3222 108 -3220
rect 114 -3216 115 -3214
rect 117 -3216 118 -3214
rect 114 -3222 115 -3220
rect 121 -3216 122 -3214
rect 121 -3222 122 -3220
rect 128 -3216 129 -3214
rect 131 -3216 132 -3214
rect 128 -3222 129 -3220
rect 135 -3216 136 -3214
rect 135 -3222 136 -3220
rect 142 -3216 143 -3214
rect 142 -3222 143 -3220
rect 149 -3216 150 -3214
rect 152 -3216 153 -3214
rect 149 -3222 150 -3220
rect 152 -3222 153 -3220
rect 156 -3216 157 -3214
rect 156 -3222 157 -3220
rect 163 -3216 164 -3214
rect 163 -3222 164 -3220
rect 170 -3216 171 -3214
rect 170 -3222 171 -3220
rect 177 -3216 178 -3214
rect 177 -3222 178 -3220
rect 184 -3216 185 -3214
rect 184 -3222 185 -3220
rect 191 -3216 192 -3214
rect 191 -3222 192 -3220
rect 198 -3216 199 -3214
rect 198 -3222 199 -3220
rect 205 -3216 206 -3214
rect 205 -3222 206 -3220
rect 212 -3216 213 -3214
rect 212 -3222 213 -3220
rect 219 -3216 220 -3214
rect 219 -3222 220 -3220
rect 226 -3216 227 -3214
rect 226 -3222 227 -3220
rect 233 -3216 234 -3214
rect 233 -3222 234 -3220
rect 243 -3222 244 -3220
rect 247 -3216 248 -3214
rect 247 -3222 248 -3220
rect 254 -3216 255 -3214
rect 254 -3222 255 -3220
rect 261 -3216 262 -3214
rect 261 -3222 262 -3220
rect 268 -3216 269 -3214
rect 268 -3222 269 -3220
rect 275 -3216 276 -3214
rect 275 -3222 276 -3220
rect 282 -3216 283 -3214
rect 282 -3222 283 -3220
rect 289 -3216 290 -3214
rect 289 -3222 290 -3220
rect 296 -3216 297 -3214
rect 296 -3222 297 -3220
rect 303 -3216 304 -3214
rect 303 -3222 304 -3220
rect 310 -3216 311 -3214
rect 310 -3222 311 -3220
rect 317 -3216 318 -3214
rect 317 -3222 318 -3220
rect 324 -3216 325 -3214
rect 324 -3222 325 -3220
rect 331 -3216 332 -3214
rect 331 -3222 332 -3220
rect 338 -3216 339 -3214
rect 338 -3222 339 -3220
rect 345 -3216 346 -3214
rect 345 -3222 346 -3220
rect 352 -3216 353 -3214
rect 352 -3222 353 -3220
rect 359 -3216 360 -3214
rect 359 -3222 360 -3220
rect 366 -3216 367 -3214
rect 366 -3222 367 -3220
rect 373 -3216 374 -3214
rect 373 -3222 374 -3220
rect 380 -3216 381 -3214
rect 380 -3222 381 -3220
rect 387 -3216 388 -3214
rect 387 -3222 388 -3220
rect 394 -3216 395 -3214
rect 394 -3222 395 -3220
rect 401 -3216 402 -3214
rect 404 -3216 405 -3214
rect 401 -3222 402 -3220
rect 404 -3222 405 -3220
rect 408 -3216 409 -3214
rect 408 -3222 409 -3220
rect 415 -3216 416 -3214
rect 415 -3222 416 -3220
rect 422 -3216 423 -3214
rect 422 -3222 423 -3220
rect 429 -3216 430 -3214
rect 432 -3216 433 -3214
rect 429 -3222 430 -3220
rect 436 -3216 437 -3214
rect 436 -3222 437 -3220
rect 443 -3216 444 -3214
rect 443 -3222 444 -3220
rect 450 -3216 451 -3214
rect 450 -3222 451 -3220
rect 457 -3216 458 -3214
rect 457 -3222 458 -3220
rect 464 -3216 465 -3214
rect 464 -3222 465 -3220
rect 471 -3216 472 -3214
rect 474 -3216 475 -3214
rect 471 -3222 472 -3220
rect 478 -3216 479 -3214
rect 478 -3222 479 -3220
rect 485 -3216 486 -3214
rect 485 -3222 486 -3220
rect 492 -3216 493 -3214
rect 492 -3222 493 -3220
rect 495 -3222 496 -3220
rect 499 -3216 500 -3214
rect 502 -3216 503 -3214
rect 499 -3222 500 -3220
rect 502 -3222 503 -3220
rect 506 -3216 507 -3214
rect 506 -3222 507 -3220
rect 513 -3216 514 -3214
rect 513 -3222 514 -3220
rect 520 -3216 521 -3214
rect 520 -3222 521 -3220
rect 527 -3216 528 -3214
rect 527 -3222 528 -3220
rect 534 -3216 535 -3214
rect 537 -3216 538 -3214
rect 534 -3222 535 -3220
rect 541 -3222 542 -3220
rect 544 -3222 545 -3220
rect 548 -3216 549 -3214
rect 548 -3222 549 -3220
rect 555 -3216 556 -3214
rect 555 -3222 556 -3220
rect 562 -3216 563 -3214
rect 562 -3222 563 -3220
rect 569 -3216 570 -3214
rect 569 -3222 570 -3220
rect 576 -3216 577 -3214
rect 579 -3216 580 -3214
rect 576 -3222 577 -3220
rect 579 -3222 580 -3220
rect 583 -3216 584 -3214
rect 583 -3222 584 -3220
rect 590 -3216 591 -3214
rect 593 -3216 594 -3214
rect 593 -3222 594 -3220
rect 597 -3216 598 -3214
rect 597 -3222 598 -3220
rect 604 -3216 605 -3214
rect 604 -3222 605 -3220
rect 611 -3216 612 -3214
rect 611 -3222 612 -3220
rect 618 -3216 619 -3214
rect 618 -3222 619 -3220
rect 625 -3216 626 -3214
rect 625 -3222 626 -3220
rect 632 -3216 633 -3214
rect 632 -3222 633 -3220
rect 639 -3216 640 -3214
rect 639 -3222 640 -3220
rect 646 -3216 647 -3214
rect 653 -3216 654 -3214
rect 656 -3216 657 -3214
rect 656 -3222 657 -3220
rect 660 -3216 661 -3214
rect 660 -3222 661 -3220
rect 667 -3216 668 -3214
rect 667 -3222 668 -3220
rect 674 -3216 675 -3214
rect 674 -3222 675 -3220
rect 681 -3216 682 -3214
rect 684 -3216 685 -3214
rect 681 -3222 682 -3220
rect 684 -3222 685 -3220
rect 688 -3216 689 -3214
rect 688 -3222 689 -3220
rect 695 -3216 696 -3214
rect 695 -3222 696 -3220
rect 702 -3216 703 -3214
rect 702 -3222 703 -3220
rect 709 -3216 710 -3214
rect 709 -3222 710 -3220
rect 716 -3216 717 -3214
rect 716 -3222 717 -3220
rect 723 -3216 724 -3214
rect 723 -3222 724 -3220
rect 730 -3216 731 -3214
rect 730 -3222 731 -3220
rect 737 -3216 738 -3214
rect 737 -3222 738 -3220
rect 744 -3216 745 -3214
rect 744 -3222 745 -3220
rect 751 -3216 752 -3214
rect 751 -3222 752 -3220
rect 758 -3216 759 -3214
rect 758 -3222 759 -3220
rect 765 -3216 766 -3214
rect 765 -3222 766 -3220
rect 772 -3216 773 -3214
rect 772 -3222 773 -3220
rect 779 -3216 780 -3214
rect 782 -3216 783 -3214
rect 779 -3222 780 -3220
rect 786 -3216 787 -3214
rect 786 -3222 787 -3220
rect 793 -3216 794 -3214
rect 796 -3216 797 -3214
rect 793 -3222 794 -3220
rect 796 -3222 797 -3220
rect 800 -3216 801 -3214
rect 800 -3222 801 -3220
rect 807 -3216 808 -3214
rect 807 -3222 808 -3220
rect 814 -3216 815 -3214
rect 814 -3222 815 -3220
rect 821 -3216 822 -3214
rect 824 -3216 825 -3214
rect 821 -3222 822 -3220
rect 824 -3222 825 -3220
rect 828 -3216 829 -3214
rect 828 -3222 829 -3220
rect 835 -3216 836 -3214
rect 838 -3216 839 -3214
rect 835 -3222 836 -3220
rect 838 -3222 839 -3220
rect 842 -3216 843 -3214
rect 842 -3222 843 -3220
rect 849 -3216 850 -3214
rect 849 -3222 850 -3220
rect 856 -3216 857 -3214
rect 856 -3222 857 -3220
rect 863 -3216 864 -3214
rect 863 -3222 864 -3220
rect 870 -3216 871 -3214
rect 870 -3222 871 -3220
rect 877 -3216 878 -3214
rect 877 -3222 878 -3220
rect 884 -3216 885 -3214
rect 884 -3222 885 -3220
rect 891 -3222 892 -3220
rect 894 -3222 895 -3220
rect 898 -3216 899 -3214
rect 898 -3222 899 -3220
rect 905 -3216 906 -3214
rect 905 -3222 906 -3220
rect 912 -3216 913 -3214
rect 912 -3222 913 -3220
rect 919 -3216 920 -3214
rect 919 -3222 920 -3220
rect 926 -3216 927 -3214
rect 926 -3222 927 -3220
rect 933 -3216 934 -3214
rect 933 -3222 934 -3220
rect 940 -3216 941 -3214
rect 940 -3222 941 -3220
rect 947 -3216 948 -3214
rect 947 -3222 948 -3220
rect 950 -3222 951 -3220
rect 954 -3216 955 -3214
rect 954 -3222 955 -3220
rect 961 -3216 962 -3214
rect 961 -3222 962 -3220
rect 968 -3216 969 -3214
rect 968 -3222 969 -3220
rect 975 -3216 976 -3214
rect 975 -3222 976 -3220
rect 982 -3216 983 -3214
rect 982 -3222 983 -3220
rect 989 -3216 990 -3214
rect 989 -3222 990 -3220
rect 996 -3216 997 -3214
rect 999 -3216 1000 -3214
rect 996 -3222 997 -3220
rect 999 -3222 1000 -3220
rect 1003 -3216 1004 -3214
rect 1003 -3222 1004 -3220
rect 1013 -3216 1014 -3214
rect 1010 -3222 1011 -3220
rect 1013 -3222 1014 -3220
rect 1017 -3216 1018 -3214
rect 1017 -3222 1018 -3220
rect 1024 -3216 1025 -3214
rect 1024 -3222 1025 -3220
rect 1031 -3216 1032 -3214
rect 1031 -3222 1032 -3220
rect 1038 -3216 1039 -3214
rect 1038 -3222 1039 -3220
rect 1045 -3216 1046 -3214
rect 1045 -3222 1046 -3220
rect 1052 -3216 1053 -3214
rect 1052 -3222 1053 -3220
rect 1059 -3216 1060 -3214
rect 1062 -3216 1063 -3214
rect 1066 -3216 1067 -3214
rect 1066 -3222 1067 -3220
rect 1073 -3216 1074 -3214
rect 1073 -3222 1074 -3220
rect 1080 -3216 1081 -3214
rect 1080 -3222 1081 -3220
rect 1087 -3216 1088 -3214
rect 1090 -3216 1091 -3214
rect 1090 -3222 1091 -3220
rect 1094 -3216 1095 -3214
rect 1094 -3222 1095 -3220
rect 1101 -3216 1102 -3214
rect 1101 -3222 1102 -3220
rect 1108 -3216 1109 -3214
rect 1108 -3222 1109 -3220
rect 1115 -3216 1116 -3214
rect 1115 -3222 1116 -3220
rect 1122 -3216 1123 -3214
rect 1122 -3222 1123 -3220
rect 1129 -3216 1130 -3214
rect 1129 -3222 1130 -3220
rect 1136 -3216 1137 -3214
rect 1136 -3222 1137 -3220
rect 1143 -3216 1144 -3214
rect 1143 -3222 1144 -3220
rect 1150 -3216 1151 -3214
rect 1150 -3222 1151 -3220
rect 1157 -3216 1158 -3214
rect 1157 -3222 1158 -3220
rect 1164 -3216 1165 -3214
rect 1164 -3222 1165 -3220
rect 1171 -3216 1172 -3214
rect 1171 -3222 1172 -3220
rect 1178 -3216 1179 -3214
rect 1178 -3222 1179 -3220
rect 1185 -3216 1186 -3214
rect 1185 -3222 1186 -3220
rect 1192 -3216 1193 -3214
rect 1192 -3222 1193 -3220
rect 1199 -3216 1200 -3214
rect 1199 -3222 1200 -3220
rect 1206 -3216 1207 -3214
rect 1206 -3222 1207 -3220
rect 1213 -3216 1214 -3214
rect 1213 -3222 1214 -3220
rect 1220 -3216 1221 -3214
rect 1220 -3222 1221 -3220
rect 1227 -3216 1228 -3214
rect 1227 -3222 1228 -3220
rect 1234 -3216 1235 -3214
rect 1234 -3222 1235 -3220
rect 1241 -3216 1242 -3214
rect 1241 -3222 1242 -3220
rect 1248 -3216 1249 -3214
rect 1248 -3222 1249 -3220
rect 1255 -3216 1256 -3214
rect 1255 -3222 1256 -3220
rect 1262 -3216 1263 -3214
rect 1262 -3222 1263 -3220
rect 1269 -3216 1270 -3214
rect 1269 -3222 1270 -3220
rect 1276 -3216 1277 -3214
rect 1276 -3222 1277 -3220
rect 1283 -3216 1284 -3214
rect 1283 -3222 1284 -3220
rect 1290 -3216 1291 -3214
rect 1290 -3222 1291 -3220
rect 1297 -3216 1298 -3214
rect 1300 -3222 1301 -3220
rect 1304 -3216 1305 -3214
rect 1304 -3222 1305 -3220
rect 1311 -3216 1312 -3214
rect 1311 -3222 1312 -3220
rect 1318 -3216 1319 -3214
rect 1318 -3222 1319 -3220
rect 1325 -3216 1326 -3214
rect 1325 -3222 1326 -3220
rect 1328 -3222 1329 -3220
rect 1332 -3216 1333 -3214
rect 1332 -3222 1333 -3220
rect 1339 -3216 1340 -3214
rect 1339 -3222 1340 -3220
rect 1346 -3216 1347 -3214
rect 1346 -3222 1347 -3220
rect 1349 -3222 1350 -3220
rect 1353 -3222 1354 -3220
rect 1356 -3222 1357 -3220
rect 1360 -3216 1361 -3214
rect 1360 -3222 1361 -3220
rect 1367 -3216 1368 -3214
rect 1367 -3222 1368 -3220
rect 1374 -3216 1375 -3214
rect 1374 -3222 1375 -3220
rect 1381 -3216 1382 -3214
rect 1381 -3222 1382 -3220
rect 1388 -3216 1389 -3214
rect 1388 -3222 1389 -3220
rect 1395 -3216 1396 -3214
rect 1395 -3222 1396 -3220
rect 1402 -3216 1403 -3214
rect 1402 -3222 1403 -3220
rect 1409 -3216 1410 -3214
rect 1412 -3216 1413 -3214
rect 1409 -3222 1410 -3220
rect 1416 -3216 1417 -3214
rect 1416 -3222 1417 -3220
rect 1423 -3216 1424 -3214
rect 1423 -3222 1424 -3220
rect 1430 -3216 1431 -3214
rect 1430 -3222 1431 -3220
rect 1437 -3216 1438 -3214
rect 1437 -3222 1438 -3220
rect 1444 -3216 1445 -3214
rect 1444 -3222 1445 -3220
rect 1451 -3216 1452 -3214
rect 1451 -3222 1452 -3220
rect 1458 -3216 1459 -3214
rect 1458 -3222 1459 -3220
rect 1465 -3216 1466 -3214
rect 1465 -3222 1466 -3220
rect 1475 -3216 1476 -3214
rect 1475 -3222 1476 -3220
rect 1479 -3216 1480 -3214
rect 1479 -3222 1480 -3220
rect 1486 -3216 1487 -3214
rect 1486 -3222 1487 -3220
rect 1493 -3216 1494 -3214
rect 1493 -3222 1494 -3220
rect 1500 -3216 1501 -3214
rect 1500 -3222 1501 -3220
rect 1507 -3216 1508 -3214
rect 1507 -3222 1508 -3220
rect 1514 -3216 1515 -3214
rect 1514 -3222 1515 -3220
rect 1521 -3216 1522 -3214
rect 1521 -3222 1522 -3220
rect 1605 -3216 1606 -3214
rect 1605 -3222 1606 -3220
rect 131 -3315 132 -3313
rect 135 -3309 136 -3307
rect 135 -3315 136 -3313
rect 163 -3309 164 -3307
rect 163 -3315 164 -3313
rect 170 -3309 171 -3307
rect 170 -3315 171 -3313
rect 177 -3309 178 -3307
rect 177 -3315 178 -3313
rect 184 -3309 185 -3307
rect 184 -3315 185 -3313
rect 191 -3309 192 -3307
rect 191 -3315 192 -3313
rect 198 -3309 199 -3307
rect 198 -3315 199 -3313
rect 205 -3309 206 -3307
rect 205 -3315 206 -3313
rect 212 -3309 213 -3307
rect 212 -3315 213 -3313
rect 219 -3309 220 -3307
rect 219 -3315 220 -3313
rect 226 -3309 227 -3307
rect 226 -3315 227 -3313
rect 233 -3309 234 -3307
rect 233 -3315 234 -3313
rect 240 -3309 241 -3307
rect 240 -3315 241 -3313
rect 247 -3309 248 -3307
rect 247 -3315 248 -3313
rect 254 -3309 255 -3307
rect 254 -3315 255 -3313
rect 261 -3309 262 -3307
rect 261 -3315 262 -3313
rect 268 -3309 269 -3307
rect 268 -3315 269 -3313
rect 275 -3309 276 -3307
rect 275 -3315 276 -3313
rect 282 -3309 283 -3307
rect 282 -3315 283 -3313
rect 289 -3309 290 -3307
rect 289 -3315 290 -3313
rect 296 -3309 297 -3307
rect 296 -3315 297 -3313
rect 303 -3309 304 -3307
rect 303 -3315 304 -3313
rect 310 -3309 311 -3307
rect 310 -3315 311 -3313
rect 317 -3309 318 -3307
rect 317 -3315 318 -3313
rect 324 -3309 325 -3307
rect 324 -3315 325 -3313
rect 331 -3309 332 -3307
rect 331 -3315 332 -3313
rect 338 -3309 339 -3307
rect 338 -3315 339 -3313
rect 345 -3309 346 -3307
rect 348 -3309 349 -3307
rect 345 -3315 346 -3313
rect 352 -3309 353 -3307
rect 352 -3315 353 -3313
rect 359 -3309 360 -3307
rect 359 -3315 360 -3313
rect 366 -3309 367 -3307
rect 366 -3315 367 -3313
rect 373 -3309 374 -3307
rect 373 -3315 374 -3313
rect 380 -3309 381 -3307
rect 380 -3315 381 -3313
rect 387 -3309 388 -3307
rect 387 -3315 388 -3313
rect 394 -3309 395 -3307
rect 394 -3315 395 -3313
rect 401 -3315 402 -3313
rect 408 -3309 409 -3307
rect 408 -3315 409 -3313
rect 415 -3309 416 -3307
rect 415 -3315 416 -3313
rect 422 -3309 423 -3307
rect 422 -3315 423 -3313
rect 429 -3309 430 -3307
rect 429 -3315 430 -3313
rect 436 -3309 437 -3307
rect 439 -3309 440 -3307
rect 443 -3309 444 -3307
rect 443 -3315 444 -3313
rect 446 -3315 447 -3313
rect 450 -3309 451 -3307
rect 450 -3315 451 -3313
rect 457 -3309 458 -3307
rect 457 -3315 458 -3313
rect 464 -3309 465 -3307
rect 464 -3315 465 -3313
rect 471 -3309 472 -3307
rect 471 -3315 472 -3313
rect 478 -3309 479 -3307
rect 478 -3315 479 -3313
rect 485 -3309 486 -3307
rect 485 -3315 486 -3313
rect 492 -3309 493 -3307
rect 499 -3309 500 -3307
rect 499 -3315 500 -3313
rect 506 -3309 507 -3307
rect 506 -3315 507 -3313
rect 513 -3309 514 -3307
rect 513 -3315 514 -3313
rect 520 -3309 521 -3307
rect 520 -3315 521 -3313
rect 527 -3309 528 -3307
rect 530 -3309 531 -3307
rect 527 -3315 528 -3313
rect 530 -3315 531 -3313
rect 534 -3309 535 -3307
rect 534 -3315 535 -3313
rect 541 -3309 542 -3307
rect 544 -3309 545 -3307
rect 544 -3315 545 -3313
rect 548 -3309 549 -3307
rect 548 -3315 549 -3313
rect 555 -3309 556 -3307
rect 555 -3315 556 -3313
rect 562 -3309 563 -3307
rect 562 -3315 563 -3313
rect 569 -3309 570 -3307
rect 569 -3315 570 -3313
rect 576 -3309 577 -3307
rect 576 -3315 577 -3313
rect 583 -3309 584 -3307
rect 583 -3315 584 -3313
rect 590 -3309 591 -3307
rect 590 -3315 591 -3313
rect 597 -3309 598 -3307
rect 597 -3315 598 -3313
rect 604 -3309 605 -3307
rect 604 -3315 605 -3313
rect 611 -3309 612 -3307
rect 611 -3315 612 -3313
rect 618 -3309 619 -3307
rect 618 -3315 619 -3313
rect 621 -3315 622 -3313
rect 625 -3309 626 -3307
rect 625 -3315 626 -3313
rect 632 -3309 633 -3307
rect 632 -3315 633 -3313
rect 639 -3309 640 -3307
rect 639 -3315 640 -3313
rect 646 -3315 647 -3313
rect 653 -3309 654 -3307
rect 653 -3315 654 -3313
rect 660 -3309 661 -3307
rect 660 -3315 661 -3313
rect 667 -3309 668 -3307
rect 667 -3315 668 -3313
rect 677 -3309 678 -3307
rect 674 -3315 675 -3313
rect 681 -3309 682 -3307
rect 681 -3315 682 -3313
rect 688 -3315 689 -3313
rect 691 -3315 692 -3313
rect 695 -3309 696 -3307
rect 695 -3315 696 -3313
rect 702 -3309 703 -3307
rect 705 -3309 706 -3307
rect 702 -3315 703 -3313
rect 705 -3315 706 -3313
rect 709 -3309 710 -3307
rect 709 -3315 710 -3313
rect 716 -3309 717 -3307
rect 716 -3315 717 -3313
rect 723 -3309 724 -3307
rect 723 -3315 724 -3313
rect 730 -3309 731 -3307
rect 730 -3315 731 -3313
rect 737 -3309 738 -3307
rect 737 -3315 738 -3313
rect 744 -3309 745 -3307
rect 744 -3315 745 -3313
rect 751 -3309 752 -3307
rect 751 -3315 752 -3313
rect 758 -3309 759 -3307
rect 758 -3315 759 -3313
rect 765 -3309 766 -3307
rect 765 -3315 766 -3313
rect 772 -3309 773 -3307
rect 772 -3315 773 -3313
rect 779 -3309 780 -3307
rect 779 -3315 780 -3313
rect 789 -3309 790 -3307
rect 786 -3315 787 -3313
rect 789 -3315 790 -3313
rect 793 -3309 794 -3307
rect 793 -3315 794 -3313
rect 800 -3309 801 -3307
rect 800 -3315 801 -3313
rect 807 -3309 808 -3307
rect 807 -3315 808 -3313
rect 814 -3309 815 -3307
rect 814 -3315 815 -3313
rect 821 -3309 822 -3307
rect 821 -3315 822 -3313
rect 828 -3309 829 -3307
rect 828 -3315 829 -3313
rect 835 -3309 836 -3307
rect 835 -3315 836 -3313
rect 842 -3309 843 -3307
rect 842 -3315 843 -3313
rect 849 -3309 850 -3307
rect 849 -3315 850 -3313
rect 856 -3309 857 -3307
rect 856 -3315 857 -3313
rect 863 -3309 864 -3307
rect 863 -3315 864 -3313
rect 870 -3315 871 -3313
rect 873 -3315 874 -3313
rect 877 -3309 878 -3307
rect 880 -3309 881 -3307
rect 877 -3315 878 -3313
rect 880 -3315 881 -3313
rect 884 -3309 885 -3307
rect 884 -3315 885 -3313
rect 891 -3309 892 -3307
rect 891 -3315 892 -3313
rect 901 -3309 902 -3307
rect 898 -3315 899 -3313
rect 901 -3315 902 -3313
rect 905 -3309 906 -3307
rect 905 -3315 906 -3313
rect 908 -3315 909 -3313
rect 912 -3309 913 -3307
rect 915 -3309 916 -3307
rect 912 -3315 913 -3313
rect 915 -3315 916 -3313
rect 919 -3309 920 -3307
rect 919 -3315 920 -3313
rect 926 -3309 927 -3307
rect 926 -3315 927 -3313
rect 933 -3309 934 -3307
rect 933 -3315 934 -3313
rect 940 -3309 941 -3307
rect 940 -3315 941 -3313
rect 947 -3309 948 -3307
rect 947 -3315 948 -3313
rect 954 -3309 955 -3307
rect 954 -3315 955 -3313
rect 961 -3309 962 -3307
rect 961 -3315 962 -3313
rect 968 -3309 969 -3307
rect 968 -3315 969 -3313
rect 975 -3309 976 -3307
rect 975 -3315 976 -3313
rect 982 -3309 983 -3307
rect 985 -3309 986 -3307
rect 982 -3315 983 -3313
rect 985 -3315 986 -3313
rect 989 -3309 990 -3307
rect 989 -3315 990 -3313
rect 996 -3309 997 -3307
rect 996 -3315 997 -3313
rect 1003 -3309 1004 -3307
rect 1003 -3315 1004 -3313
rect 1010 -3309 1011 -3307
rect 1010 -3315 1011 -3313
rect 1020 -3309 1021 -3307
rect 1020 -3315 1021 -3313
rect 1024 -3309 1025 -3307
rect 1024 -3315 1025 -3313
rect 1031 -3309 1032 -3307
rect 1031 -3315 1032 -3313
rect 1038 -3309 1039 -3307
rect 1038 -3315 1039 -3313
rect 1045 -3309 1046 -3307
rect 1045 -3315 1046 -3313
rect 1052 -3309 1053 -3307
rect 1052 -3315 1053 -3313
rect 1059 -3309 1060 -3307
rect 1059 -3315 1060 -3313
rect 1066 -3309 1067 -3307
rect 1066 -3315 1067 -3313
rect 1073 -3309 1074 -3307
rect 1073 -3315 1074 -3313
rect 1080 -3309 1081 -3307
rect 1080 -3315 1081 -3313
rect 1087 -3309 1088 -3307
rect 1087 -3315 1088 -3313
rect 1094 -3309 1095 -3307
rect 1094 -3315 1095 -3313
rect 1101 -3309 1102 -3307
rect 1101 -3315 1102 -3313
rect 1108 -3309 1109 -3307
rect 1108 -3315 1109 -3313
rect 1111 -3315 1112 -3313
rect 1115 -3309 1116 -3307
rect 1115 -3315 1116 -3313
rect 1122 -3309 1123 -3307
rect 1122 -3315 1123 -3313
rect 1129 -3309 1130 -3307
rect 1129 -3315 1130 -3313
rect 1136 -3309 1137 -3307
rect 1136 -3315 1137 -3313
rect 1143 -3309 1144 -3307
rect 1143 -3315 1144 -3313
rect 1150 -3309 1151 -3307
rect 1150 -3315 1151 -3313
rect 1157 -3309 1158 -3307
rect 1157 -3315 1158 -3313
rect 1164 -3309 1165 -3307
rect 1164 -3315 1165 -3313
rect 1171 -3309 1172 -3307
rect 1171 -3315 1172 -3313
rect 1178 -3309 1179 -3307
rect 1178 -3315 1179 -3313
rect 1188 -3309 1189 -3307
rect 1185 -3315 1186 -3313
rect 1192 -3309 1193 -3307
rect 1192 -3315 1193 -3313
rect 1199 -3309 1200 -3307
rect 1199 -3315 1200 -3313
rect 1209 -3309 1210 -3307
rect 1206 -3315 1207 -3313
rect 1209 -3315 1210 -3313
rect 1213 -3309 1214 -3307
rect 1213 -3315 1214 -3313
rect 1216 -3315 1217 -3313
rect 1220 -3309 1221 -3307
rect 1220 -3315 1221 -3313
rect 1227 -3309 1228 -3307
rect 1227 -3315 1228 -3313
rect 1234 -3309 1235 -3307
rect 1234 -3315 1235 -3313
rect 1241 -3309 1242 -3307
rect 1241 -3315 1242 -3313
rect 1248 -3315 1249 -3313
rect 1251 -3315 1252 -3313
rect 1255 -3309 1256 -3307
rect 1258 -3309 1259 -3307
rect 1262 -3309 1263 -3307
rect 1265 -3309 1266 -3307
rect 1262 -3315 1263 -3313
rect 1265 -3315 1266 -3313
rect 1269 -3309 1270 -3307
rect 1269 -3315 1270 -3313
rect 1276 -3309 1277 -3307
rect 1276 -3315 1277 -3313
rect 1283 -3309 1284 -3307
rect 1283 -3315 1284 -3313
rect 1290 -3309 1291 -3307
rect 1290 -3315 1291 -3313
rect 1297 -3309 1298 -3307
rect 1297 -3315 1298 -3313
rect 1304 -3309 1305 -3307
rect 1304 -3315 1305 -3313
rect 1311 -3309 1312 -3307
rect 1311 -3315 1312 -3313
rect 1318 -3309 1319 -3307
rect 1318 -3315 1319 -3313
rect 1325 -3309 1326 -3307
rect 1328 -3309 1329 -3307
rect 1325 -3315 1326 -3313
rect 1332 -3309 1333 -3307
rect 1332 -3315 1333 -3313
rect 1339 -3309 1340 -3307
rect 1339 -3315 1340 -3313
rect 1346 -3309 1347 -3307
rect 1346 -3315 1347 -3313
rect 1353 -3309 1354 -3307
rect 1353 -3315 1354 -3313
rect 1360 -3309 1361 -3307
rect 1360 -3315 1361 -3313
rect 1381 -3309 1382 -3307
rect 1381 -3315 1382 -3313
rect 1388 -3309 1389 -3307
rect 1388 -3315 1389 -3313
rect 1531 -3309 1532 -3307
rect 1528 -3315 1529 -3313
rect 1584 -3309 1585 -3307
rect 1584 -3315 1585 -3313
rect 240 -3406 241 -3404
rect 240 -3412 241 -3410
rect 247 -3406 248 -3404
rect 247 -3412 248 -3410
rect 268 -3406 269 -3404
rect 268 -3412 269 -3410
rect 282 -3406 283 -3404
rect 282 -3412 283 -3410
rect 289 -3406 290 -3404
rect 289 -3412 290 -3410
rect 292 -3412 293 -3410
rect 296 -3406 297 -3404
rect 299 -3412 300 -3410
rect 303 -3406 304 -3404
rect 303 -3412 304 -3410
rect 310 -3406 311 -3404
rect 310 -3412 311 -3410
rect 317 -3406 318 -3404
rect 317 -3412 318 -3410
rect 324 -3406 325 -3404
rect 324 -3412 325 -3410
rect 331 -3406 332 -3404
rect 331 -3412 332 -3410
rect 338 -3406 339 -3404
rect 338 -3412 339 -3410
rect 345 -3406 346 -3404
rect 345 -3412 346 -3410
rect 352 -3406 353 -3404
rect 352 -3412 353 -3410
rect 359 -3406 360 -3404
rect 359 -3412 360 -3410
rect 366 -3406 367 -3404
rect 366 -3412 367 -3410
rect 373 -3406 374 -3404
rect 376 -3412 377 -3410
rect 380 -3406 381 -3404
rect 380 -3412 381 -3410
rect 387 -3406 388 -3404
rect 387 -3412 388 -3410
rect 394 -3406 395 -3404
rect 394 -3412 395 -3410
rect 401 -3406 402 -3404
rect 401 -3412 402 -3410
rect 408 -3406 409 -3404
rect 408 -3412 409 -3410
rect 415 -3406 416 -3404
rect 415 -3412 416 -3410
rect 422 -3406 423 -3404
rect 422 -3412 423 -3410
rect 429 -3406 430 -3404
rect 429 -3412 430 -3410
rect 436 -3406 437 -3404
rect 436 -3412 437 -3410
rect 443 -3406 444 -3404
rect 443 -3412 444 -3410
rect 450 -3406 451 -3404
rect 450 -3412 451 -3410
rect 457 -3406 458 -3404
rect 457 -3412 458 -3410
rect 464 -3406 465 -3404
rect 464 -3412 465 -3410
rect 471 -3406 472 -3404
rect 471 -3412 472 -3410
rect 478 -3406 479 -3404
rect 478 -3412 479 -3410
rect 485 -3406 486 -3404
rect 485 -3412 486 -3410
rect 492 -3406 493 -3404
rect 492 -3412 493 -3410
rect 499 -3406 500 -3404
rect 499 -3412 500 -3410
rect 506 -3406 507 -3404
rect 506 -3412 507 -3410
rect 513 -3406 514 -3404
rect 513 -3412 514 -3410
rect 523 -3406 524 -3404
rect 520 -3412 521 -3410
rect 523 -3412 524 -3410
rect 527 -3406 528 -3404
rect 527 -3412 528 -3410
rect 534 -3406 535 -3404
rect 534 -3412 535 -3410
rect 541 -3406 542 -3404
rect 541 -3412 542 -3410
rect 548 -3406 549 -3404
rect 548 -3412 549 -3410
rect 555 -3406 556 -3404
rect 555 -3412 556 -3410
rect 562 -3406 563 -3404
rect 562 -3412 563 -3410
rect 569 -3406 570 -3404
rect 569 -3412 570 -3410
rect 576 -3406 577 -3404
rect 579 -3406 580 -3404
rect 579 -3412 580 -3410
rect 583 -3406 584 -3404
rect 583 -3412 584 -3410
rect 590 -3406 591 -3404
rect 590 -3412 591 -3410
rect 597 -3406 598 -3404
rect 597 -3412 598 -3410
rect 604 -3406 605 -3404
rect 604 -3412 605 -3410
rect 611 -3406 612 -3404
rect 614 -3406 615 -3404
rect 614 -3412 615 -3410
rect 618 -3406 619 -3404
rect 618 -3412 619 -3410
rect 625 -3406 626 -3404
rect 625 -3412 626 -3410
rect 632 -3406 633 -3404
rect 632 -3412 633 -3410
rect 639 -3406 640 -3404
rect 639 -3412 640 -3410
rect 646 -3406 647 -3404
rect 646 -3412 647 -3410
rect 653 -3406 654 -3404
rect 653 -3412 654 -3410
rect 660 -3406 661 -3404
rect 660 -3412 661 -3410
rect 667 -3406 668 -3404
rect 667 -3412 668 -3410
rect 674 -3406 675 -3404
rect 674 -3412 675 -3410
rect 681 -3406 682 -3404
rect 681 -3412 682 -3410
rect 688 -3406 689 -3404
rect 688 -3412 689 -3410
rect 695 -3406 696 -3404
rect 695 -3412 696 -3410
rect 702 -3406 703 -3404
rect 702 -3412 703 -3410
rect 709 -3406 710 -3404
rect 709 -3412 710 -3410
rect 716 -3406 717 -3404
rect 716 -3412 717 -3410
rect 723 -3406 724 -3404
rect 723 -3412 724 -3410
rect 730 -3412 731 -3410
rect 733 -3412 734 -3410
rect 737 -3406 738 -3404
rect 737 -3412 738 -3410
rect 744 -3406 745 -3404
rect 744 -3412 745 -3410
rect 751 -3406 752 -3404
rect 751 -3412 752 -3410
rect 758 -3406 759 -3404
rect 758 -3412 759 -3410
rect 765 -3406 766 -3404
rect 765 -3412 766 -3410
rect 772 -3406 773 -3404
rect 772 -3412 773 -3410
rect 779 -3406 780 -3404
rect 779 -3412 780 -3410
rect 786 -3406 787 -3404
rect 786 -3412 787 -3410
rect 793 -3406 794 -3404
rect 793 -3412 794 -3410
rect 800 -3406 801 -3404
rect 803 -3406 804 -3404
rect 803 -3412 804 -3410
rect 807 -3406 808 -3404
rect 807 -3412 808 -3410
rect 814 -3406 815 -3404
rect 814 -3412 815 -3410
rect 821 -3406 822 -3404
rect 821 -3412 822 -3410
rect 828 -3406 829 -3404
rect 828 -3412 829 -3410
rect 835 -3406 836 -3404
rect 835 -3412 836 -3410
rect 842 -3406 843 -3404
rect 842 -3412 843 -3410
rect 849 -3406 850 -3404
rect 849 -3412 850 -3410
rect 856 -3406 857 -3404
rect 856 -3412 857 -3410
rect 863 -3406 864 -3404
rect 863 -3412 864 -3410
rect 870 -3406 871 -3404
rect 870 -3412 871 -3410
rect 877 -3406 878 -3404
rect 877 -3412 878 -3410
rect 884 -3406 885 -3404
rect 884 -3412 885 -3410
rect 894 -3406 895 -3404
rect 891 -3412 892 -3410
rect 894 -3412 895 -3410
rect 898 -3406 899 -3404
rect 898 -3412 899 -3410
rect 905 -3406 906 -3404
rect 905 -3412 906 -3410
rect 912 -3406 913 -3404
rect 912 -3412 913 -3410
rect 919 -3406 920 -3404
rect 919 -3412 920 -3410
rect 926 -3406 927 -3404
rect 926 -3412 927 -3410
rect 933 -3406 934 -3404
rect 933 -3412 934 -3410
rect 940 -3406 941 -3404
rect 940 -3412 941 -3410
rect 947 -3406 948 -3404
rect 950 -3406 951 -3404
rect 947 -3412 948 -3410
rect 954 -3406 955 -3404
rect 954 -3412 955 -3410
rect 961 -3406 962 -3404
rect 961 -3412 962 -3410
rect 968 -3406 969 -3404
rect 968 -3412 969 -3410
rect 975 -3406 976 -3404
rect 975 -3412 976 -3410
rect 982 -3406 983 -3404
rect 982 -3412 983 -3410
rect 989 -3406 990 -3404
rect 989 -3412 990 -3410
rect 996 -3406 997 -3404
rect 996 -3412 997 -3410
rect 1003 -3406 1004 -3404
rect 1003 -3412 1004 -3410
rect 1013 -3406 1014 -3404
rect 1010 -3412 1011 -3410
rect 1017 -3406 1018 -3404
rect 1020 -3406 1021 -3404
rect 1017 -3412 1018 -3410
rect 1020 -3412 1021 -3410
rect 1024 -3406 1025 -3404
rect 1024 -3412 1025 -3410
rect 1031 -3406 1032 -3404
rect 1031 -3412 1032 -3410
rect 1038 -3406 1039 -3404
rect 1038 -3412 1039 -3410
rect 1041 -3412 1042 -3410
rect 1045 -3406 1046 -3404
rect 1045 -3412 1046 -3410
rect 1055 -3412 1056 -3410
rect 1059 -3406 1060 -3404
rect 1062 -3406 1063 -3404
rect 1066 -3406 1067 -3404
rect 1066 -3412 1067 -3410
rect 1073 -3406 1074 -3404
rect 1073 -3412 1074 -3410
rect 1080 -3406 1081 -3404
rect 1080 -3412 1081 -3410
rect 1087 -3406 1088 -3404
rect 1087 -3412 1088 -3410
rect 1094 -3406 1095 -3404
rect 1094 -3412 1095 -3410
rect 1101 -3406 1102 -3404
rect 1101 -3412 1102 -3410
rect 1108 -3406 1109 -3404
rect 1111 -3412 1112 -3410
rect 1115 -3406 1116 -3404
rect 1115 -3412 1116 -3410
rect 1122 -3406 1123 -3404
rect 1122 -3412 1123 -3410
rect 1129 -3406 1130 -3404
rect 1129 -3412 1130 -3410
rect 1136 -3406 1137 -3404
rect 1136 -3412 1137 -3410
rect 1143 -3406 1144 -3404
rect 1153 -3406 1154 -3404
rect 1150 -3412 1151 -3410
rect 1153 -3412 1154 -3410
rect 1157 -3406 1158 -3404
rect 1157 -3412 1158 -3410
rect 1160 -3412 1161 -3410
rect 1164 -3406 1165 -3404
rect 1167 -3406 1168 -3404
rect 1167 -3412 1168 -3410
rect 1171 -3406 1172 -3404
rect 1171 -3412 1172 -3410
rect 1185 -3406 1186 -3404
rect 1185 -3412 1186 -3410
rect 1192 -3406 1193 -3404
rect 1192 -3412 1193 -3410
rect 1199 -3406 1200 -3404
rect 1199 -3412 1200 -3410
rect 1206 -3406 1207 -3404
rect 1206 -3412 1207 -3410
rect 1213 -3406 1214 -3404
rect 1213 -3412 1214 -3410
rect 1216 -3412 1217 -3410
rect 1234 -3406 1235 -3404
rect 1234 -3412 1235 -3410
rect 1241 -3406 1242 -3404
rect 1241 -3412 1242 -3410
rect 1248 -3406 1249 -3404
rect 1248 -3412 1249 -3410
rect 1265 -3406 1266 -3404
rect 1265 -3412 1266 -3410
rect 1311 -3406 1312 -3404
rect 1311 -3412 1312 -3410
rect 1318 -3406 1319 -3404
rect 1318 -3412 1319 -3410
rect 1332 -3406 1333 -3404
rect 1332 -3412 1333 -3410
rect 1374 -3406 1375 -3404
rect 1374 -3412 1375 -3410
rect 1381 -3406 1382 -3404
rect 1381 -3412 1382 -3410
rect 1384 -3412 1385 -3410
rect 1388 -3406 1389 -3404
rect 1388 -3412 1389 -3410
rect 1577 -3406 1578 -3404
rect 1577 -3412 1578 -3410
rect 261 -3453 262 -3451
rect 261 -3459 262 -3457
rect 310 -3453 311 -3451
rect 310 -3459 311 -3457
rect 317 -3453 318 -3451
rect 317 -3459 318 -3457
rect 338 -3453 339 -3451
rect 338 -3459 339 -3457
rect 345 -3453 346 -3451
rect 345 -3459 346 -3457
rect 352 -3453 353 -3451
rect 355 -3453 356 -3451
rect 355 -3459 356 -3457
rect 359 -3453 360 -3451
rect 359 -3459 360 -3457
rect 366 -3453 367 -3451
rect 366 -3459 367 -3457
rect 373 -3453 374 -3451
rect 373 -3459 374 -3457
rect 380 -3453 381 -3451
rect 380 -3459 381 -3457
rect 387 -3453 388 -3451
rect 387 -3459 388 -3457
rect 394 -3453 395 -3451
rect 394 -3459 395 -3457
rect 401 -3453 402 -3451
rect 401 -3459 402 -3457
rect 411 -3459 412 -3457
rect 415 -3453 416 -3451
rect 415 -3459 416 -3457
rect 422 -3453 423 -3451
rect 422 -3459 423 -3457
rect 429 -3453 430 -3451
rect 429 -3459 430 -3457
rect 436 -3453 437 -3451
rect 436 -3459 437 -3457
rect 443 -3453 444 -3451
rect 443 -3459 444 -3457
rect 450 -3453 451 -3451
rect 450 -3459 451 -3457
rect 457 -3453 458 -3451
rect 457 -3459 458 -3457
rect 464 -3453 465 -3451
rect 464 -3459 465 -3457
rect 471 -3453 472 -3451
rect 474 -3453 475 -3451
rect 478 -3453 479 -3451
rect 478 -3459 479 -3457
rect 485 -3453 486 -3451
rect 485 -3459 486 -3457
rect 492 -3453 493 -3451
rect 492 -3459 493 -3457
rect 499 -3453 500 -3451
rect 499 -3459 500 -3457
rect 506 -3453 507 -3451
rect 509 -3453 510 -3451
rect 506 -3459 507 -3457
rect 513 -3453 514 -3451
rect 513 -3459 514 -3457
rect 520 -3453 521 -3451
rect 520 -3459 521 -3457
rect 527 -3453 528 -3451
rect 527 -3459 528 -3457
rect 534 -3453 535 -3451
rect 534 -3459 535 -3457
rect 541 -3453 542 -3451
rect 541 -3459 542 -3457
rect 548 -3453 549 -3451
rect 548 -3459 549 -3457
rect 555 -3453 556 -3451
rect 555 -3459 556 -3457
rect 562 -3453 563 -3451
rect 562 -3459 563 -3457
rect 569 -3453 570 -3451
rect 569 -3459 570 -3457
rect 576 -3453 577 -3451
rect 576 -3459 577 -3457
rect 583 -3453 584 -3451
rect 586 -3453 587 -3451
rect 583 -3459 584 -3457
rect 586 -3459 587 -3457
rect 590 -3459 591 -3457
rect 593 -3459 594 -3457
rect 597 -3453 598 -3451
rect 597 -3459 598 -3457
rect 604 -3453 605 -3451
rect 604 -3459 605 -3457
rect 607 -3459 608 -3457
rect 611 -3453 612 -3451
rect 611 -3459 612 -3457
rect 621 -3453 622 -3451
rect 618 -3459 619 -3457
rect 621 -3459 622 -3457
rect 625 -3453 626 -3451
rect 625 -3459 626 -3457
rect 632 -3453 633 -3451
rect 632 -3459 633 -3457
rect 639 -3453 640 -3451
rect 639 -3459 640 -3457
rect 646 -3453 647 -3451
rect 646 -3459 647 -3457
rect 656 -3453 657 -3451
rect 653 -3459 654 -3457
rect 660 -3453 661 -3451
rect 663 -3453 664 -3451
rect 660 -3459 661 -3457
rect 663 -3459 664 -3457
rect 667 -3453 668 -3451
rect 667 -3459 668 -3457
rect 674 -3453 675 -3451
rect 674 -3459 675 -3457
rect 681 -3453 682 -3451
rect 681 -3459 682 -3457
rect 688 -3453 689 -3451
rect 688 -3459 689 -3457
rect 695 -3453 696 -3451
rect 695 -3459 696 -3457
rect 702 -3453 703 -3451
rect 702 -3459 703 -3457
rect 709 -3453 710 -3451
rect 709 -3459 710 -3457
rect 716 -3453 717 -3451
rect 719 -3459 720 -3457
rect 723 -3453 724 -3451
rect 723 -3459 724 -3457
rect 730 -3453 731 -3451
rect 730 -3459 731 -3457
rect 737 -3453 738 -3451
rect 737 -3459 738 -3457
rect 744 -3453 745 -3451
rect 744 -3459 745 -3457
rect 751 -3453 752 -3451
rect 751 -3459 752 -3457
rect 758 -3453 759 -3451
rect 758 -3459 759 -3457
rect 765 -3453 766 -3451
rect 765 -3459 766 -3457
rect 772 -3453 773 -3451
rect 772 -3459 773 -3457
rect 779 -3453 780 -3451
rect 779 -3459 780 -3457
rect 786 -3453 787 -3451
rect 786 -3459 787 -3457
rect 793 -3453 794 -3451
rect 793 -3459 794 -3457
rect 800 -3453 801 -3451
rect 800 -3459 801 -3457
rect 807 -3453 808 -3451
rect 810 -3453 811 -3451
rect 807 -3459 808 -3457
rect 814 -3453 815 -3451
rect 814 -3459 815 -3457
rect 821 -3453 822 -3451
rect 824 -3453 825 -3451
rect 821 -3459 822 -3457
rect 828 -3453 829 -3451
rect 828 -3459 829 -3457
rect 835 -3453 836 -3451
rect 835 -3459 836 -3457
rect 842 -3453 843 -3451
rect 842 -3459 843 -3457
rect 849 -3453 850 -3451
rect 852 -3453 853 -3451
rect 852 -3459 853 -3457
rect 856 -3453 857 -3451
rect 856 -3459 857 -3457
rect 863 -3453 864 -3451
rect 863 -3459 864 -3457
rect 870 -3453 871 -3451
rect 870 -3459 871 -3457
rect 877 -3453 878 -3451
rect 877 -3459 878 -3457
rect 884 -3453 885 -3451
rect 884 -3459 885 -3457
rect 891 -3453 892 -3451
rect 891 -3459 892 -3457
rect 898 -3453 899 -3451
rect 898 -3459 899 -3457
rect 905 -3453 906 -3451
rect 905 -3459 906 -3457
rect 912 -3453 913 -3451
rect 912 -3459 913 -3457
rect 919 -3453 920 -3451
rect 919 -3459 920 -3457
rect 926 -3453 927 -3451
rect 926 -3459 927 -3457
rect 933 -3453 934 -3451
rect 933 -3459 934 -3457
rect 940 -3453 941 -3451
rect 940 -3459 941 -3457
rect 947 -3453 948 -3451
rect 947 -3459 948 -3457
rect 954 -3453 955 -3451
rect 961 -3453 962 -3451
rect 961 -3459 962 -3457
rect 968 -3459 969 -3457
rect 975 -3453 976 -3451
rect 975 -3459 976 -3457
rect 982 -3453 983 -3451
rect 982 -3459 983 -3457
rect 989 -3453 990 -3451
rect 989 -3459 990 -3457
rect 996 -3453 997 -3451
rect 999 -3453 1000 -3451
rect 996 -3459 997 -3457
rect 1003 -3453 1004 -3451
rect 1003 -3459 1004 -3457
rect 1010 -3453 1011 -3451
rect 1010 -3459 1011 -3457
rect 1017 -3453 1018 -3451
rect 1017 -3459 1018 -3457
rect 1024 -3453 1025 -3451
rect 1024 -3459 1025 -3457
rect 1031 -3453 1032 -3451
rect 1031 -3459 1032 -3457
rect 1052 -3453 1053 -3451
rect 1052 -3459 1053 -3457
rect 1073 -3453 1074 -3451
rect 1073 -3459 1074 -3457
rect 1080 -3453 1081 -3451
rect 1080 -3459 1081 -3457
rect 1101 -3453 1102 -3451
rect 1101 -3459 1102 -3457
rect 1115 -3453 1116 -3451
rect 1115 -3459 1116 -3457
rect 1118 -3459 1119 -3457
rect 1122 -3453 1123 -3451
rect 1122 -3459 1123 -3457
rect 1129 -3453 1130 -3451
rect 1129 -3459 1130 -3457
rect 1136 -3453 1137 -3451
rect 1136 -3459 1137 -3457
rect 1143 -3459 1144 -3457
rect 1192 -3453 1193 -3451
rect 1192 -3459 1193 -3457
rect 1199 -3453 1200 -3451
rect 1199 -3459 1200 -3457
rect 1206 -3453 1207 -3451
rect 1206 -3459 1207 -3457
rect 1213 -3453 1214 -3451
rect 1213 -3459 1214 -3457
rect 1269 -3453 1270 -3451
rect 1269 -3459 1270 -3457
rect 1300 -3453 1301 -3451
rect 1297 -3459 1298 -3457
rect 1300 -3459 1301 -3457
rect 1304 -3453 1305 -3451
rect 1304 -3459 1305 -3457
rect 1318 -3453 1319 -3451
rect 1318 -3459 1319 -3457
rect 1346 -3453 1347 -3451
rect 1346 -3459 1347 -3457
rect 1381 -3453 1382 -3451
rect 1384 -3453 1385 -3451
rect 1381 -3459 1382 -3457
rect 1388 -3453 1389 -3451
rect 1388 -3459 1389 -3457
rect 1395 -3453 1396 -3451
rect 1395 -3459 1396 -3457
rect 1577 -3453 1578 -3451
rect 1577 -3459 1578 -3457
rect 268 -3494 269 -3492
rect 268 -3500 269 -3498
rect 282 -3500 283 -3498
rect 285 -3500 286 -3498
rect 296 -3494 297 -3492
rect 296 -3500 297 -3498
rect 366 -3494 367 -3492
rect 366 -3500 367 -3498
rect 373 -3494 374 -3492
rect 373 -3500 374 -3498
rect 380 -3494 381 -3492
rect 380 -3500 381 -3498
rect 390 -3494 391 -3492
rect 390 -3500 391 -3498
rect 408 -3494 409 -3492
rect 408 -3500 409 -3498
rect 422 -3494 423 -3492
rect 425 -3494 426 -3492
rect 429 -3494 430 -3492
rect 429 -3500 430 -3498
rect 439 -3494 440 -3492
rect 439 -3500 440 -3498
rect 443 -3494 444 -3492
rect 443 -3500 444 -3498
rect 450 -3494 451 -3492
rect 450 -3500 451 -3498
rect 457 -3494 458 -3492
rect 457 -3500 458 -3498
rect 471 -3494 472 -3492
rect 471 -3500 472 -3498
rect 478 -3494 479 -3492
rect 478 -3500 479 -3498
rect 485 -3494 486 -3492
rect 485 -3500 486 -3498
rect 492 -3494 493 -3492
rect 492 -3500 493 -3498
rect 499 -3494 500 -3492
rect 499 -3500 500 -3498
rect 506 -3494 507 -3492
rect 506 -3500 507 -3498
rect 513 -3494 514 -3492
rect 513 -3500 514 -3498
rect 527 -3494 528 -3492
rect 527 -3500 528 -3498
rect 534 -3494 535 -3492
rect 534 -3500 535 -3498
rect 541 -3494 542 -3492
rect 541 -3500 542 -3498
rect 548 -3494 549 -3492
rect 548 -3500 549 -3498
rect 555 -3494 556 -3492
rect 555 -3500 556 -3498
rect 562 -3494 563 -3492
rect 562 -3500 563 -3498
rect 569 -3494 570 -3492
rect 569 -3500 570 -3498
rect 576 -3494 577 -3492
rect 576 -3500 577 -3498
rect 583 -3494 584 -3492
rect 583 -3500 584 -3498
rect 590 -3494 591 -3492
rect 590 -3500 591 -3498
rect 604 -3494 605 -3492
rect 604 -3500 605 -3498
rect 618 -3494 619 -3492
rect 618 -3500 619 -3498
rect 632 -3494 633 -3492
rect 632 -3500 633 -3498
rect 639 -3494 640 -3492
rect 639 -3500 640 -3498
rect 646 -3494 647 -3492
rect 646 -3500 647 -3498
rect 653 -3494 654 -3492
rect 656 -3494 657 -3492
rect 656 -3500 657 -3498
rect 688 -3494 689 -3492
rect 688 -3500 689 -3498
rect 695 -3494 696 -3492
rect 695 -3500 696 -3498
rect 702 -3494 703 -3492
rect 702 -3500 703 -3498
rect 709 -3494 710 -3492
rect 709 -3500 710 -3498
rect 716 -3494 717 -3492
rect 716 -3500 717 -3498
rect 723 -3494 724 -3492
rect 726 -3500 727 -3498
rect 730 -3494 731 -3492
rect 733 -3494 734 -3492
rect 730 -3500 731 -3498
rect 733 -3500 734 -3498
rect 737 -3494 738 -3492
rect 737 -3500 738 -3498
rect 744 -3494 745 -3492
rect 744 -3500 745 -3498
rect 754 -3494 755 -3492
rect 754 -3500 755 -3498
rect 758 -3494 759 -3492
rect 758 -3500 759 -3498
rect 765 -3494 766 -3492
rect 765 -3500 766 -3498
rect 772 -3494 773 -3492
rect 772 -3500 773 -3498
rect 786 -3494 787 -3492
rect 786 -3500 787 -3498
rect 793 -3494 794 -3492
rect 800 -3494 801 -3492
rect 800 -3500 801 -3498
rect 807 -3494 808 -3492
rect 807 -3500 808 -3498
rect 814 -3494 815 -3492
rect 814 -3500 815 -3498
rect 821 -3494 822 -3492
rect 821 -3500 822 -3498
rect 828 -3494 829 -3492
rect 828 -3500 829 -3498
rect 877 -3494 878 -3492
rect 877 -3500 878 -3498
rect 884 -3494 885 -3492
rect 884 -3500 885 -3498
rect 891 -3494 892 -3492
rect 891 -3500 892 -3498
rect 898 -3494 899 -3492
rect 898 -3500 899 -3498
rect 905 -3494 906 -3492
rect 905 -3500 906 -3498
rect 912 -3494 913 -3492
rect 915 -3494 916 -3492
rect 912 -3500 913 -3498
rect 919 -3494 920 -3492
rect 919 -3500 920 -3498
rect 926 -3494 927 -3492
rect 926 -3500 927 -3498
rect 933 -3494 934 -3492
rect 933 -3500 934 -3498
rect 940 -3494 941 -3492
rect 940 -3500 941 -3498
rect 947 -3494 948 -3492
rect 947 -3500 948 -3498
rect 954 -3500 955 -3498
rect 961 -3494 962 -3492
rect 961 -3500 962 -3498
rect 975 -3494 976 -3492
rect 975 -3500 976 -3498
rect 996 -3494 997 -3492
rect 996 -3500 997 -3498
rect 1003 -3494 1004 -3492
rect 1006 -3494 1007 -3492
rect 1003 -3500 1004 -3498
rect 1010 -3494 1011 -3492
rect 1010 -3500 1011 -3498
rect 1024 -3494 1025 -3492
rect 1024 -3500 1025 -3498
rect 1038 -3494 1039 -3492
rect 1038 -3500 1039 -3498
rect 1045 -3494 1046 -3492
rect 1045 -3500 1046 -3498
rect 1048 -3500 1049 -3498
rect 1052 -3494 1053 -3492
rect 1052 -3500 1053 -3498
rect 1059 -3494 1060 -3492
rect 1059 -3500 1060 -3498
rect 1066 -3494 1067 -3492
rect 1066 -3500 1067 -3498
rect 1073 -3494 1074 -3492
rect 1073 -3500 1074 -3498
rect 1080 -3494 1081 -3492
rect 1080 -3500 1081 -3498
rect 1087 -3494 1088 -3492
rect 1090 -3494 1091 -3492
rect 1090 -3500 1091 -3498
rect 1115 -3494 1116 -3492
rect 1118 -3494 1119 -3492
rect 1115 -3500 1116 -3498
rect 1122 -3494 1123 -3492
rect 1122 -3500 1123 -3498
rect 1136 -3494 1137 -3492
rect 1136 -3500 1137 -3498
rect 1157 -3494 1158 -3492
rect 1157 -3500 1158 -3498
rect 1178 -3494 1179 -3492
rect 1181 -3494 1182 -3492
rect 1181 -3500 1182 -3498
rect 1185 -3494 1186 -3492
rect 1185 -3500 1186 -3498
rect 1192 -3494 1193 -3492
rect 1192 -3500 1193 -3498
rect 1234 -3494 1235 -3492
rect 1234 -3500 1235 -3498
rect 1248 -3494 1249 -3492
rect 1248 -3500 1249 -3498
rect 1269 -3494 1270 -3492
rect 1269 -3500 1270 -3498
rect 1276 -3494 1277 -3492
rect 1276 -3500 1277 -3498
rect 1374 -3494 1375 -3492
rect 1374 -3500 1375 -3498
rect 1381 -3494 1382 -3492
rect 1384 -3500 1385 -3498
rect 1388 -3494 1389 -3492
rect 1388 -3500 1389 -3498
rect 1395 -3494 1396 -3492
rect 1395 -3500 1396 -3498
rect 1416 -3494 1417 -3492
rect 1416 -3500 1417 -3498
rect 1577 -3494 1578 -3492
rect 1577 -3500 1578 -3498
rect 380 -3525 381 -3523
rect 380 -3531 381 -3529
rect 387 -3525 388 -3523
rect 387 -3531 388 -3529
rect 394 -3525 395 -3523
rect 394 -3531 395 -3529
rect 401 -3525 402 -3523
rect 401 -3531 402 -3529
rect 429 -3525 430 -3523
rect 429 -3531 430 -3529
rect 443 -3525 444 -3523
rect 443 -3531 444 -3529
rect 450 -3525 451 -3523
rect 450 -3531 451 -3529
rect 464 -3525 465 -3523
rect 464 -3531 465 -3529
rect 478 -3525 479 -3523
rect 481 -3525 482 -3523
rect 478 -3531 479 -3529
rect 485 -3525 486 -3523
rect 485 -3531 486 -3529
rect 492 -3525 493 -3523
rect 492 -3531 493 -3529
rect 499 -3525 500 -3523
rect 499 -3531 500 -3529
rect 506 -3525 507 -3523
rect 506 -3531 507 -3529
rect 513 -3525 514 -3523
rect 513 -3531 514 -3529
rect 520 -3525 521 -3523
rect 520 -3531 521 -3529
rect 527 -3525 528 -3523
rect 527 -3531 528 -3529
rect 534 -3525 535 -3523
rect 534 -3531 535 -3529
rect 541 -3525 542 -3523
rect 541 -3531 542 -3529
rect 548 -3525 549 -3523
rect 548 -3531 549 -3529
rect 558 -3525 559 -3523
rect 555 -3531 556 -3529
rect 558 -3531 559 -3529
rect 565 -3525 566 -3523
rect 562 -3531 563 -3529
rect 565 -3531 566 -3529
rect 569 -3525 570 -3523
rect 569 -3531 570 -3529
rect 576 -3525 577 -3523
rect 576 -3531 577 -3529
rect 583 -3525 584 -3523
rect 583 -3531 584 -3529
rect 590 -3525 591 -3523
rect 590 -3531 591 -3529
rect 597 -3525 598 -3523
rect 597 -3531 598 -3529
rect 604 -3525 605 -3523
rect 604 -3531 605 -3529
rect 646 -3525 647 -3523
rect 646 -3531 647 -3529
rect 653 -3525 654 -3523
rect 653 -3531 654 -3529
rect 674 -3525 675 -3523
rect 674 -3531 675 -3529
rect 695 -3525 696 -3523
rect 695 -3531 696 -3529
rect 702 -3525 703 -3523
rect 702 -3531 703 -3529
rect 709 -3525 710 -3523
rect 709 -3531 710 -3529
rect 730 -3525 731 -3523
rect 730 -3531 731 -3529
rect 758 -3525 759 -3523
rect 758 -3531 759 -3529
rect 765 -3525 766 -3523
rect 765 -3531 766 -3529
rect 772 -3525 773 -3523
rect 772 -3531 773 -3529
rect 779 -3525 780 -3523
rect 779 -3531 780 -3529
rect 786 -3525 787 -3523
rect 786 -3531 787 -3529
rect 793 -3531 794 -3529
rect 800 -3525 801 -3523
rect 800 -3531 801 -3529
rect 807 -3525 808 -3523
rect 807 -3531 808 -3529
rect 814 -3525 815 -3523
rect 814 -3531 815 -3529
rect 821 -3525 822 -3523
rect 824 -3531 825 -3529
rect 842 -3525 843 -3523
rect 842 -3531 843 -3529
rect 863 -3525 864 -3523
rect 863 -3531 864 -3529
rect 877 -3525 878 -3523
rect 877 -3531 878 -3529
rect 884 -3525 885 -3523
rect 884 -3531 885 -3529
rect 891 -3531 892 -3529
rect 898 -3525 899 -3523
rect 898 -3531 899 -3529
rect 905 -3525 906 -3523
rect 905 -3531 906 -3529
rect 919 -3525 920 -3523
rect 919 -3531 920 -3529
rect 926 -3525 927 -3523
rect 926 -3531 927 -3529
rect 933 -3525 934 -3523
rect 933 -3531 934 -3529
rect 940 -3525 941 -3523
rect 940 -3531 941 -3529
rect 947 -3525 948 -3523
rect 950 -3531 951 -3529
rect 954 -3525 955 -3523
rect 957 -3525 958 -3523
rect 957 -3531 958 -3529
rect 961 -3525 962 -3523
rect 964 -3525 965 -3523
rect 968 -3525 969 -3523
rect 968 -3531 969 -3529
rect 1003 -3525 1004 -3523
rect 1017 -3525 1018 -3523
rect 1020 -3525 1021 -3523
rect 1031 -3525 1032 -3523
rect 1034 -3525 1035 -3523
rect 1038 -3525 1039 -3523
rect 1041 -3525 1042 -3523
rect 1038 -3531 1039 -3529
rect 1045 -3525 1046 -3523
rect 1048 -3525 1049 -3523
rect 1045 -3531 1046 -3529
rect 1052 -3525 1053 -3523
rect 1052 -3531 1053 -3529
rect 1062 -3525 1063 -3523
rect 1059 -3531 1060 -3529
rect 1073 -3525 1074 -3523
rect 1073 -3531 1074 -3529
rect 1115 -3525 1116 -3523
rect 1115 -3531 1116 -3529
rect 1129 -3525 1130 -3523
rect 1129 -3531 1130 -3529
rect 1136 -3525 1137 -3523
rect 1136 -3531 1137 -3529
rect 1143 -3525 1144 -3523
rect 1143 -3531 1144 -3529
rect 1157 -3531 1158 -3529
rect 1164 -3525 1165 -3523
rect 1164 -3531 1165 -3529
rect 1178 -3525 1179 -3523
rect 1178 -3531 1179 -3529
rect 1192 -3525 1193 -3523
rect 1192 -3531 1193 -3529
rect 1262 -3525 1263 -3523
rect 1262 -3531 1263 -3529
rect 1276 -3525 1277 -3523
rect 1279 -3525 1280 -3523
rect 1279 -3531 1280 -3529
rect 1339 -3525 1340 -3523
rect 1339 -3531 1340 -3529
rect 1381 -3525 1382 -3523
rect 1381 -3531 1382 -3529
rect 1395 -3525 1396 -3523
rect 1395 -3531 1396 -3529
rect 1500 -3525 1501 -3523
rect 1500 -3531 1501 -3529
rect 1577 -3525 1578 -3523
rect 1580 -3531 1581 -3529
rect 380 -3554 381 -3552
rect 380 -3560 381 -3558
rect 387 -3554 388 -3552
rect 387 -3560 388 -3558
rect 394 -3554 395 -3552
rect 394 -3560 395 -3558
rect 401 -3554 402 -3552
rect 401 -3560 402 -3558
rect 408 -3554 409 -3552
rect 408 -3560 409 -3558
rect 450 -3554 451 -3552
rect 450 -3560 451 -3558
rect 457 -3554 458 -3552
rect 457 -3560 458 -3558
rect 474 -3554 475 -3552
rect 474 -3560 475 -3558
rect 478 -3554 479 -3552
rect 478 -3560 479 -3558
rect 492 -3554 493 -3552
rect 492 -3560 493 -3558
rect 499 -3554 500 -3552
rect 502 -3560 503 -3558
rect 506 -3554 507 -3552
rect 506 -3560 507 -3558
rect 513 -3554 514 -3552
rect 513 -3560 514 -3558
rect 527 -3554 528 -3552
rect 527 -3560 528 -3558
rect 530 -3560 531 -3558
rect 534 -3554 535 -3552
rect 534 -3560 535 -3558
rect 541 -3554 542 -3552
rect 541 -3560 542 -3558
rect 548 -3554 549 -3552
rect 548 -3560 549 -3558
rect 555 -3554 556 -3552
rect 555 -3560 556 -3558
rect 565 -3554 566 -3552
rect 562 -3560 563 -3558
rect 569 -3554 570 -3552
rect 569 -3560 570 -3558
rect 576 -3554 577 -3552
rect 576 -3560 577 -3558
rect 579 -3560 580 -3558
rect 583 -3554 584 -3552
rect 583 -3560 584 -3558
rect 590 -3554 591 -3552
rect 590 -3560 591 -3558
rect 597 -3554 598 -3552
rect 597 -3560 598 -3558
rect 607 -3554 608 -3552
rect 660 -3554 661 -3552
rect 663 -3554 664 -3552
rect 667 -3554 668 -3552
rect 667 -3560 668 -3558
rect 702 -3554 703 -3552
rect 705 -3554 706 -3552
rect 702 -3560 703 -3558
rect 709 -3554 710 -3552
rect 709 -3560 710 -3558
rect 737 -3554 738 -3552
rect 737 -3560 738 -3558
rect 758 -3554 759 -3552
rect 758 -3560 759 -3558
rect 765 -3560 766 -3558
rect 768 -3560 769 -3558
rect 772 -3554 773 -3552
rect 772 -3560 773 -3558
rect 779 -3554 780 -3552
rect 779 -3560 780 -3558
rect 786 -3554 787 -3552
rect 786 -3560 787 -3558
rect 796 -3554 797 -3552
rect 793 -3560 794 -3558
rect 796 -3560 797 -3558
rect 800 -3554 801 -3552
rect 800 -3560 801 -3558
rect 807 -3554 808 -3552
rect 807 -3560 808 -3558
rect 814 -3554 815 -3552
rect 814 -3560 815 -3558
rect 877 -3554 878 -3552
rect 877 -3560 878 -3558
rect 884 -3554 885 -3552
rect 884 -3560 885 -3558
rect 898 -3554 899 -3552
rect 898 -3560 899 -3558
rect 905 -3554 906 -3552
rect 905 -3560 906 -3558
rect 926 -3554 927 -3552
rect 926 -3560 927 -3558
rect 936 -3554 937 -3552
rect 933 -3560 934 -3558
rect 940 -3554 941 -3552
rect 940 -3560 941 -3558
rect 950 -3560 951 -3558
rect 1108 -3554 1109 -3552
rect 1111 -3554 1112 -3552
rect 1111 -3560 1112 -3558
rect 1115 -3554 1116 -3552
rect 1115 -3560 1116 -3558
rect 1129 -3554 1130 -3552
rect 1129 -3560 1130 -3558
rect 1136 -3554 1137 -3552
rect 1136 -3560 1137 -3558
rect 1164 -3554 1165 -3552
rect 1164 -3560 1165 -3558
rect 1178 -3554 1179 -3552
rect 1178 -3560 1179 -3558
rect 1192 -3554 1193 -3552
rect 1192 -3560 1193 -3558
rect 1360 -3554 1361 -3552
rect 1360 -3560 1361 -3558
rect 1388 -3554 1389 -3552
rect 1388 -3560 1389 -3558
rect 1395 -3554 1396 -3552
rect 1395 -3560 1396 -3558
rect 387 -3569 388 -3567
rect 387 -3575 388 -3573
rect 394 -3569 395 -3567
rect 397 -3575 398 -3573
rect 401 -3569 402 -3567
rect 404 -3569 405 -3567
rect 401 -3575 402 -3573
rect 408 -3569 409 -3567
rect 408 -3575 409 -3573
rect 457 -3569 458 -3567
rect 457 -3575 458 -3573
rect 464 -3569 465 -3567
rect 464 -3575 465 -3573
rect 492 -3569 493 -3567
rect 492 -3575 493 -3573
rect 499 -3569 500 -3567
rect 502 -3575 503 -3573
rect 562 -3569 563 -3567
rect 562 -3575 563 -3573
rect 576 -3569 577 -3567
rect 579 -3575 580 -3573
rect 590 -3569 591 -3567
rect 590 -3575 591 -3573
rect 597 -3575 598 -3573
rect 600 -3575 601 -3573
rect 632 -3569 633 -3567
rect 632 -3575 633 -3573
rect 747 -3569 748 -3567
rect 747 -3575 748 -3573
rect 758 -3569 759 -3567
rect 758 -3575 759 -3573
rect 800 -3569 801 -3567
rect 800 -3575 801 -3573
rect 807 -3569 808 -3567
rect 810 -3575 811 -3573
rect 884 -3569 885 -3567
rect 884 -3575 885 -3573
rect 891 -3569 892 -3567
rect 894 -3569 895 -3567
rect 901 -3569 902 -3567
rect 898 -3575 899 -3573
rect 1132 -3569 1133 -3567
rect 1129 -3575 1130 -3573
rect 1136 -3569 1137 -3567
rect 1136 -3575 1137 -3573
rect 1171 -3569 1172 -3567
rect 1171 -3575 1172 -3573
rect 1178 -3575 1179 -3573
rect 1181 -3575 1182 -3573
rect 1185 -3569 1186 -3567
rect 1185 -3575 1186 -3573
rect 1195 -3575 1196 -3573
rect 1199 -3569 1200 -3567
rect 1199 -3575 1200 -3573
rect 1388 -3569 1389 -3567
rect 1391 -3569 1392 -3567
rect 1388 -3575 1389 -3573
rect 1395 -3569 1396 -3567
rect 1395 -3575 1396 -3573
<< metal1 >>
rect 233 0 437 1
rect 443 0 458 1
rect 527 0 549 1
rect 555 0 755 1
rect 877 0 955 1
rect 345 -2 353 -1
rect 359 -2 468 -1
rect 604 -2 615 -1
rect 653 -2 678 -1
rect 716 -2 801 -1
rect 380 -4 535 -3
rect 670 -4 689 -3
rect 401 -6 461 -5
rect 408 -8 433 -7
rect 453 -8 472 -7
rect 415 -10 507 -9
rect 422 -12 451 -11
rect 145 -23 150 -22
rect 156 -23 234 -22
rect 261 -23 307 -22
rect 324 -23 360 -22
rect 373 -23 409 -22
rect 425 -23 444 -22
rect 450 -23 556 -22
rect 590 -23 822 -22
rect 842 -23 885 -22
rect 954 -23 990 -22
rect 226 -25 237 -24
rect 282 -25 391 -24
rect 394 -25 416 -24
rect 429 -25 444 -24
rect 460 -25 556 -24
rect 618 -25 633 -24
rect 653 -25 668 -24
rect 677 -25 682 -24
rect 688 -25 703 -24
rect 712 -25 773 -24
rect 800 -25 829 -24
rect 331 -27 381 -26
rect 408 -27 563 -26
rect 653 -27 671 -26
rect 677 -27 731 -26
rect 751 -27 997 -26
rect 338 -29 346 -28
rect 380 -29 402 -28
rect 436 -29 661 -28
rect 688 -29 720 -28
rect 758 -29 899 -28
rect 401 -31 423 -30
rect 432 -31 437 -30
rect 460 -31 745 -30
rect 814 -31 881 -30
rect 464 -33 598 -32
rect 716 -33 755 -32
rect 471 -35 479 -34
rect 492 -35 507 -34
rect 509 -35 612 -34
rect 471 -37 517 -36
rect 520 -37 640 -36
rect 495 -39 500 -38
rect 513 -39 626 -38
rect 523 -41 542 -40
rect 551 -41 577 -40
rect 530 -43 549 -42
rect 534 -45 647 -44
rect 527 -47 535 -46
rect 537 -47 584 -46
rect 464 -49 528 -48
rect 128 -60 157 -59
rect 191 -60 199 -59
rect 205 -60 227 -59
rect 254 -60 433 -59
rect 474 -60 738 -59
rect 744 -60 871 -59
rect 884 -60 941 -59
rect 989 -60 1011 -59
rect 219 -62 283 -61
rect 289 -62 325 -61
rect 345 -62 423 -61
rect 478 -62 489 -61
rect 492 -62 710 -61
rect 716 -62 745 -61
rect 751 -62 888 -61
rect 898 -62 955 -61
rect 996 -62 1088 -61
rect 261 -64 269 -63
rect 275 -64 458 -63
rect 478 -64 591 -63
rect 625 -64 696 -63
rect 730 -64 787 -63
rect 796 -64 864 -63
rect 936 -64 948 -63
rect 247 -66 262 -65
rect 282 -66 461 -65
rect 506 -66 521 -65
rect 551 -66 678 -65
rect 688 -66 717 -65
rect 772 -66 836 -65
rect 296 -68 409 -67
rect 422 -68 437 -67
rect 506 -68 594 -67
rect 625 -68 811 -67
rect 817 -68 857 -67
rect 303 -70 339 -69
rect 352 -70 416 -69
rect 555 -70 675 -69
rect 702 -70 731 -69
rect 779 -70 885 -69
rect 306 -72 360 -71
rect 366 -72 402 -71
rect 415 -72 517 -71
rect 555 -72 577 -71
rect 583 -72 689 -71
rect 800 -72 829 -71
rect 310 -74 451 -73
rect 530 -74 584 -73
rect 590 -74 619 -73
rect 646 -74 710 -73
rect 807 -74 843 -73
rect 317 -76 332 -75
rect 338 -76 465 -75
rect 541 -76 577 -75
rect 597 -76 703 -75
rect 712 -76 843 -75
rect 324 -78 374 -77
rect 376 -78 381 -77
rect 387 -78 437 -77
rect 464 -78 472 -77
rect 499 -78 542 -77
rect 604 -78 619 -77
rect 649 -78 794 -77
rect 814 -78 829 -77
rect 331 -80 444 -79
rect 534 -80 598 -79
rect 660 -80 724 -79
rect 821 -80 892 -79
rect 334 -82 500 -81
rect 513 -82 535 -81
rect 569 -82 605 -81
rect 611 -82 661 -81
rect 373 -84 381 -83
rect 387 -84 524 -83
rect 548 -84 570 -83
rect 632 -84 822 -83
rect 401 -86 430 -85
rect 562 -86 612 -85
rect 411 -88 451 -87
rect 562 -88 654 -87
rect 653 -90 668 -89
rect 667 -92 682 -91
rect 639 -94 682 -93
rect 639 -96 759 -95
rect 89 -107 94 -106
rect 114 -107 129 -106
rect 135 -107 220 -106
rect 226 -107 293 -106
rect 345 -107 363 -106
rect 373 -107 395 -106
rect 408 -107 468 -106
rect 471 -107 489 -106
rect 513 -107 549 -106
rect 611 -107 647 -106
rect 656 -107 745 -106
rect 793 -107 822 -106
rect 828 -107 913 -106
rect 940 -107 997 -106
rect 1010 -107 1039 -106
rect 1087 -107 1130 -106
rect 1195 -107 1221 -106
rect 142 -109 255 -108
rect 261 -109 472 -108
rect 481 -109 552 -108
rect 646 -109 717 -108
rect 723 -109 850 -108
rect 856 -109 899 -108
rect 947 -109 969 -108
rect 156 -111 332 -110
rect 380 -111 384 -110
rect 394 -111 640 -110
rect 674 -111 759 -110
rect 810 -111 941 -110
rect 954 -111 983 -110
rect 163 -113 206 -112
rect 219 -113 304 -112
rect 310 -113 374 -112
rect 380 -113 444 -112
rect 450 -113 458 -112
rect 485 -113 510 -112
rect 513 -113 934 -112
rect 170 -115 356 -114
rect 376 -115 486 -114
rect 530 -115 549 -114
rect 576 -115 640 -114
rect 681 -115 724 -114
rect 744 -115 801 -114
rect 817 -115 829 -114
rect 835 -115 920 -114
rect 177 -117 339 -116
rect 352 -117 458 -116
rect 537 -117 626 -116
rect 660 -117 801 -116
rect 824 -117 1011 -116
rect 184 -119 192 -118
rect 198 -119 248 -118
rect 250 -119 311 -118
rect 317 -119 332 -118
rect 338 -119 633 -118
rect 698 -119 906 -118
rect 191 -121 276 -120
rect 289 -121 430 -120
rect 450 -121 503 -120
rect 576 -121 654 -120
rect 709 -121 808 -120
rect 842 -121 962 -120
rect 208 -123 318 -122
rect 383 -123 444 -122
rect 460 -123 633 -122
rect 716 -123 769 -122
rect 779 -123 836 -122
rect 856 -123 878 -122
rect 880 -123 927 -122
rect 243 -125 346 -124
rect 408 -125 423 -124
rect 590 -125 675 -124
rect 796 -125 843 -124
rect 863 -125 955 -124
rect 247 -127 521 -126
rect 569 -127 591 -126
rect 597 -127 682 -126
rect 814 -127 864 -126
rect 870 -127 976 -126
rect 254 -129 283 -128
rect 296 -129 423 -128
rect 432 -129 598 -128
rect 611 -129 661 -128
rect 737 -129 815 -128
rect 884 -129 1137 -128
rect 261 -131 475 -130
rect 520 -131 948 -130
rect 268 -133 304 -132
rect 432 -133 465 -132
rect 618 -133 710 -132
rect 786 -133 871 -132
rect 268 -135 367 -134
rect 415 -135 465 -134
rect 618 -135 752 -134
rect 275 -137 563 -136
rect 625 -137 668 -136
rect 688 -137 752 -136
rect 282 -139 388 -138
rect 401 -139 416 -138
rect 534 -139 563 -138
rect 649 -139 780 -138
rect 296 -141 479 -140
rect 534 -141 556 -140
rect 667 -141 794 -140
rect 366 -143 654 -142
rect 702 -143 738 -142
rect 352 -145 703 -144
rect 730 -145 787 -144
rect 387 -147 437 -146
rect 478 -147 570 -146
rect 695 -147 731 -146
rect 401 -149 528 -148
rect 359 -151 528 -150
rect 359 -153 773 -152
rect 436 -155 542 -154
rect 492 -157 556 -156
rect 492 -159 507 -158
rect 541 -159 605 -158
rect 499 -161 605 -160
rect 499 -163 888 -162
rect 506 -165 689 -164
rect 51 -176 164 -175
rect 177 -176 507 -175
rect 516 -176 1158 -175
rect 1220 -176 1228 -175
rect 58 -178 262 -177
rect 296 -178 500 -177
rect 530 -178 829 -177
rect 849 -178 885 -177
rect 887 -178 1088 -177
rect 1097 -178 1151 -177
rect 65 -180 451 -179
rect 457 -180 482 -179
rect 544 -180 724 -179
rect 737 -180 1032 -179
rect 1038 -180 1109 -179
rect 1118 -180 1196 -179
rect 72 -182 157 -181
rect 163 -182 433 -181
rect 443 -182 500 -181
rect 541 -182 738 -181
rect 772 -182 1025 -181
rect 1129 -182 1172 -181
rect 79 -184 465 -183
rect 474 -184 1284 -183
rect 86 -186 241 -185
rect 261 -186 353 -185
rect 366 -186 496 -185
rect 548 -186 724 -185
rect 772 -186 822 -185
rect 863 -186 1039 -185
rect 1125 -186 1130 -185
rect 1136 -186 1256 -185
rect 93 -188 101 -187
rect 107 -188 115 -187
rect 121 -188 514 -187
rect 548 -188 615 -187
rect 653 -188 836 -187
rect 870 -188 1053 -187
rect 93 -190 171 -189
rect 177 -190 192 -189
rect 212 -190 304 -189
rect 317 -190 353 -189
rect 380 -190 510 -189
rect 614 -190 759 -189
rect 789 -190 843 -189
rect 877 -190 892 -189
rect 905 -190 1018 -189
rect 117 -192 171 -191
rect 184 -192 202 -191
rect 219 -192 360 -191
rect 380 -192 528 -191
rect 569 -192 843 -191
rect 880 -192 899 -191
rect 905 -192 969 -191
rect 975 -192 1081 -191
rect 128 -194 269 -193
rect 292 -194 367 -193
rect 383 -194 514 -193
rect 656 -194 976 -193
rect 996 -194 1102 -193
rect 142 -196 216 -195
rect 219 -196 283 -195
rect 296 -196 584 -195
rect 688 -196 836 -195
rect 898 -196 941 -195
rect 954 -196 1074 -195
rect 142 -198 150 -197
rect 156 -198 594 -197
rect 688 -198 857 -197
rect 933 -198 1144 -197
rect 149 -200 409 -199
rect 415 -200 447 -199
rect 457 -200 633 -199
rect 681 -200 857 -199
rect 940 -200 962 -199
rect 968 -200 983 -199
rect 996 -200 1060 -199
rect 184 -202 199 -201
rect 254 -202 283 -201
rect 303 -202 521 -201
rect 632 -202 675 -201
rect 681 -202 920 -201
rect 999 -202 1067 -201
rect 191 -204 206 -203
rect 254 -204 325 -203
rect 345 -204 409 -203
rect 429 -204 535 -203
rect 562 -204 675 -203
rect 698 -204 1004 -203
rect 1010 -204 1137 -203
rect 268 -206 388 -205
rect 394 -206 451 -205
rect 492 -206 584 -205
rect 709 -206 864 -205
rect 947 -206 1011 -205
rect 275 -208 416 -207
rect 509 -208 654 -207
rect 716 -208 1046 -207
rect 208 -210 276 -209
rect 289 -210 325 -209
rect 345 -210 363 -209
rect 387 -210 524 -209
rect 534 -210 731 -209
rect 744 -210 871 -209
rect 243 -212 290 -211
rect 310 -212 395 -211
rect 422 -212 731 -211
rect 751 -212 983 -211
rect 135 -214 244 -213
rect 310 -214 332 -213
rect 359 -214 832 -213
rect 135 -216 234 -215
rect 317 -216 339 -215
rect 422 -216 570 -215
rect 604 -216 710 -215
rect 765 -216 892 -215
rect 233 -218 759 -217
rect 765 -218 927 -217
rect 247 -220 339 -219
rect 471 -220 927 -219
rect 247 -222 545 -221
rect 562 -222 591 -221
rect 604 -222 626 -221
rect 660 -222 752 -221
rect 768 -222 920 -221
rect 331 -224 580 -223
rect 702 -224 745 -223
rect 779 -224 934 -223
rect 436 -226 472 -225
rect 478 -226 591 -225
rect 611 -226 780 -225
rect 793 -226 962 -225
rect 236 -228 437 -227
rect 520 -228 577 -227
rect 611 -228 948 -227
rect 226 -230 237 -229
rect 541 -230 626 -229
rect 793 -230 913 -229
rect 226 -232 374 -231
rect 555 -232 661 -231
rect 719 -232 913 -231
rect 373 -234 444 -233
rect 555 -234 696 -233
rect 796 -234 1165 -233
rect 572 -236 696 -235
rect 800 -236 850 -235
rect 502 -238 801 -237
rect 807 -238 990 -237
rect 618 -240 703 -239
rect 786 -240 808 -239
rect 814 -240 955 -239
rect 460 -242 619 -241
rect 597 -244 815 -243
rect 597 -246 668 -245
rect 485 -248 668 -247
rect 401 -250 486 -249
rect 401 -252 468 -251
rect 44 -263 297 -262
rect 383 -263 542 -262
rect 548 -263 591 -262
rect 593 -263 948 -262
rect 989 -263 1382 -262
rect 51 -265 237 -264
rect 285 -265 1151 -264
rect 1164 -265 1347 -264
rect 51 -267 430 -266
rect 460 -267 668 -266
rect 681 -267 948 -266
rect 996 -267 1158 -266
rect 1202 -267 1354 -266
rect 58 -269 342 -268
rect 415 -269 465 -268
rect 471 -269 752 -268
rect 772 -269 822 -268
rect 828 -269 1214 -268
rect 1255 -269 1375 -268
rect 61 -271 73 -270
rect 86 -271 472 -270
rect 474 -271 836 -270
rect 842 -271 1291 -270
rect 72 -273 94 -272
rect 96 -273 122 -272
rect 142 -273 416 -272
rect 474 -273 1326 -272
rect 65 -275 143 -274
rect 156 -275 234 -274
rect 338 -275 430 -274
rect 506 -275 1235 -274
rect 1283 -275 1592 -274
rect 65 -277 454 -276
rect 509 -277 857 -276
rect 863 -277 1340 -276
rect 86 -279 139 -278
rect 163 -279 468 -278
rect 513 -279 1389 -278
rect 107 -281 297 -280
rect 387 -281 514 -280
rect 527 -281 1361 -280
rect 107 -283 458 -282
rect 527 -283 584 -282
rect 614 -283 983 -282
rect 1024 -283 1207 -282
rect 93 -285 458 -284
rect 499 -285 584 -284
rect 632 -285 836 -284
rect 863 -285 1095 -284
rect 1101 -285 1368 -284
rect 121 -287 157 -286
rect 163 -287 206 -286
rect 215 -287 1263 -286
rect 170 -289 283 -288
rect 352 -289 388 -288
rect 450 -289 507 -288
rect 509 -289 633 -288
rect 667 -289 1277 -288
rect 198 -291 549 -290
rect 576 -291 829 -290
rect 891 -291 895 -290
rect 905 -291 990 -290
rect 1038 -291 1284 -290
rect 135 -293 577 -292
rect 579 -293 640 -292
rect 681 -293 717 -292
rect 723 -293 843 -292
rect 891 -293 899 -292
rect 912 -293 1242 -292
rect 201 -295 381 -294
rect 408 -295 451 -294
rect 478 -295 640 -294
rect 688 -295 822 -294
rect 894 -295 899 -294
rect 933 -295 1095 -294
rect 1101 -295 1144 -294
rect 1171 -295 1256 -294
rect 114 -297 934 -296
rect 1045 -297 1298 -296
rect 205 -299 531 -298
rect 544 -299 717 -298
rect 744 -299 983 -298
rect 1052 -299 1305 -298
rect 282 -301 346 -300
rect 359 -301 479 -300
rect 499 -301 1396 -300
rect 275 -303 346 -302
rect 359 -303 374 -302
rect 443 -303 1172 -302
rect 198 -305 444 -304
rect 611 -305 1039 -304
rect 1059 -305 1151 -304
rect 317 -307 353 -306
rect 373 -307 423 -306
rect 611 -307 1032 -306
rect 1073 -307 1333 -306
rect 58 -309 1032 -308
rect 1073 -309 1098 -308
rect 1108 -309 1319 -308
rect 324 -311 409 -310
rect 422 -311 556 -310
rect 614 -311 724 -310
rect 747 -311 1004 -310
rect 1017 -311 1109 -310
rect 1115 -311 1130 -310
rect 1136 -311 1312 -310
rect 173 -313 1116 -312
rect 1118 -313 1249 -312
rect 324 -315 734 -314
rect 751 -315 1186 -314
rect 492 -317 1130 -316
rect 226 -319 493 -318
rect 555 -319 794 -318
rect 800 -319 906 -318
rect 968 -319 1060 -318
rect 1066 -319 1137 -318
rect 149 -321 227 -320
rect 495 -321 801 -320
rect 814 -321 1025 -320
rect 1080 -321 1165 -320
rect 149 -323 244 -322
rect 618 -323 689 -322
rect 695 -323 913 -322
rect 919 -323 969 -322
rect 975 -323 1046 -322
rect 1087 -323 1221 -322
rect 607 -325 619 -324
rect 625 -325 696 -324
rect 705 -325 1179 -324
rect 520 -327 626 -326
rect 670 -327 1053 -326
rect 1122 -327 1193 -326
rect 520 -329 535 -328
rect 674 -329 794 -328
rect 870 -329 1004 -328
rect 366 -331 535 -330
rect 562 -331 871 -330
rect 926 -331 1088 -330
rect 191 -333 563 -332
rect 653 -333 675 -332
rect 709 -333 815 -332
rect 884 -333 927 -332
rect 961 -333 1123 -332
rect 79 -335 710 -334
rect 712 -335 1270 -334
rect 79 -337 332 -336
rect 439 -337 654 -336
rect 730 -337 920 -336
rect 975 -337 1011 -336
rect 177 -339 192 -338
rect 254 -339 367 -338
rect 730 -339 1018 -338
rect 177 -341 248 -340
rect 331 -341 573 -340
rect 754 -341 885 -340
rect 999 -341 1081 -340
rect 208 -343 255 -342
rect 758 -343 1067 -342
rect 646 -345 759 -344
rect 779 -345 857 -344
rect 877 -345 962 -344
rect 194 -347 647 -346
rect 660 -347 780 -346
rect 786 -347 1144 -346
rect 117 -349 787 -348
rect 789 -349 955 -348
rect 117 -351 241 -350
rect 569 -351 878 -350
rect 940 -351 955 -350
rect 569 -353 1158 -352
rect 604 -355 661 -354
rect 737 -355 941 -354
rect 485 -357 738 -356
rect 849 -357 1011 -356
rect 401 -359 486 -358
rect 597 -359 605 -358
rect 765 -359 850 -358
rect 289 -361 598 -360
rect 702 -361 766 -360
rect 275 -363 703 -362
rect 289 -365 304 -364
rect 338 -365 402 -364
rect 303 -367 395 -366
rect 268 -369 395 -368
rect 268 -371 311 -370
rect 261 -373 311 -372
rect 219 -375 262 -374
rect 219 -377 437 -376
rect 128 -379 437 -378
rect 100 -381 129 -380
rect 100 -383 412 -382
rect 23 -394 234 -393
rect 247 -394 454 -393
rect 506 -394 1291 -393
rect 1297 -394 1445 -393
rect 1591 -394 1711 -393
rect 30 -396 444 -395
rect 450 -396 1487 -395
rect 37 -398 101 -397
rect 107 -398 363 -397
rect 408 -398 584 -397
rect 597 -398 731 -397
rect 1143 -398 1452 -397
rect 58 -400 276 -399
rect 317 -400 388 -399
rect 429 -400 524 -399
rect 530 -400 745 -399
rect 1031 -400 1144 -399
rect 1164 -400 1466 -399
rect 82 -402 577 -401
rect 607 -402 1340 -401
rect 1346 -402 1501 -401
rect 86 -404 409 -403
rect 429 -404 759 -403
rect 933 -404 1032 -403
rect 1052 -404 1165 -403
rect 1171 -404 1340 -403
rect 1353 -404 1480 -403
rect 86 -406 584 -405
rect 611 -406 794 -405
rect 807 -406 1053 -405
rect 1066 -406 1172 -405
rect 1178 -406 1298 -405
rect 1304 -406 1410 -405
rect 89 -408 129 -407
rect 135 -408 934 -407
rect 982 -408 1067 -407
rect 1073 -408 1179 -407
rect 1220 -408 1494 -407
rect 93 -410 104 -409
rect 110 -410 920 -409
rect 982 -410 1081 -409
rect 1094 -410 1221 -409
rect 1227 -410 1291 -409
rect 1311 -410 1417 -409
rect 96 -412 682 -411
rect 695 -412 794 -411
rect 905 -412 1095 -411
rect 1115 -412 1228 -411
rect 1269 -412 1424 -411
rect 100 -414 1249 -413
rect 1269 -414 1399 -413
rect 114 -416 262 -415
rect 268 -416 286 -415
rect 324 -416 475 -415
rect 481 -416 1074 -415
rect 1136 -416 1347 -415
rect 1353 -416 1525 -415
rect 65 -418 269 -417
rect 324 -418 570 -417
rect 576 -418 689 -417
rect 695 -418 738 -417
rect 747 -418 1312 -417
rect 1318 -418 1431 -417
rect 65 -420 360 -419
rect 366 -420 388 -419
rect 436 -420 528 -419
rect 534 -420 594 -419
rect 618 -420 731 -419
rect 733 -420 1305 -419
rect 1325 -420 1473 -419
rect 79 -422 367 -421
rect 401 -422 437 -421
rect 439 -422 745 -421
rect 758 -422 843 -421
rect 884 -422 1326 -421
rect 1332 -422 1459 -421
rect 79 -424 360 -423
rect 474 -424 1137 -423
rect 1192 -424 1333 -423
rect 1374 -424 1508 -423
rect 121 -426 300 -425
rect 331 -426 402 -425
rect 485 -426 507 -425
rect 534 -426 1319 -425
rect 121 -428 500 -427
rect 541 -428 570 -427
rect 639 -428 752 -427
rect 842 -428 1123 -427
rect 1206 -428 1375 -427
rect 124 -430 1130 -429
rect 1276 -430 1403 -429
rect 128 -432 136 -431
rect 163 -432 167 -431
rect 170 -432 419 -431
rect 464 -432 486 -431
rect 492 -432 542 -431
rect 653 -432 752 -431
rect 856 -432 885 -431
rect 919 -432 927 -431
rect 954 -432 1249 -431
rect 1283 -432 1438 -431
rect 51 -434 654 -433
rect 660 -434 668 -433
rect 670 -434 1389 -433
rect 51 -436 304 -435
rect 331 -436 472 -435
rect 478 -436 500 -435
rect 509 -436 857 -435
rect 898 -436 955 -435
rect 968 -436 1130 -435
rect 1255 -436 1389 -435
rect 163 -438 290 -437
rect 303 -438 395 -437
rect 443 -438 493 -437
rect 604 -438 927 -437
rect 989 -438 1116 -437
rect 1150 -438 1256 -437
rect 1283 -438 1368 -437
rect 166 -440 290 -439
rect 352 -440 528 -439
rect 562 -440 605 -439
rect 625 -440 661 -439
rect 674 -440 682 -439
rect 702 -440 1382 -439
rect 26 -442 563 -441
rect 632 -442 675 -441
rect 712 -442 1277 -441
rect 142 -444 626 -443
rect 632 -444 1515 -443
rect 142 -446 297 -445
rect 352 -446 556 -445
rect 716 -446 808 -445
rect 863 -446 969 -445
rect 1010 -446 1123 -445
rect 1213 -446 1368 -445
rect 117 -448 717 -447
rect 800 -448 864 -447
rect 877 -448 990 -447
rect 1017 -448 1207 -447
rect 1241 -448 1382 -447
rect 170 -450 423 -449
rect 464 -450 591 -449
rect 649 -450 878 -449
rect 891 -450 1011 -449
rect 1017 -450 1102 -449
rect 1108 -450 1214 -449
rect 180 -452 703 -451
rect 709 -452 1242 -451
rect 187 -454 423 -453
rect 478 -454 1361 -453
rect 194 -456 612 -455
rect 779 -456 892 -455
rect 898 -456 1529 -455
rect 198 -458 906 -457
rect 996 -458 1109 -457
rect 1199 -458 1361 -457
rect 184 -460 199 -459
rect 205 -460 262 -459
rect 282 -460 738 -459
rect 870 -460 997 -459
rect 1003 -460 1102 -459
rect 1185 -460 1200 -459
rect 205 -462 514 -461
rect 520 -462 556 -461
rect 590 -462 822 -461
rect 870 -462 948 -461
rect 1003 -462 1396 -461
rect 44 -464 822 -463
rect 849 -464 948 -463
rect 1038 -464 1151 -463
rect 1262 -464 1396 -463
rect 44 -466 227 -465
rect 254 -466 276 -465
rect 282 -466 496 -465
rect 520 -466 1025 -465
rect 1045 -466 1081 -465
rect 1087 -466 1186 -465
rect 191 -468 227 -467
rect 254 -468 615 -467
rect 635 -468 1263 -467
rect 191 -470 514 -469
rect 723 -470 780 -469
rect 786 -470 850 -469
rect 940 -470 1046 -469
rect 1087 -470 1158 -469
rect 138 -472 787 -471
rect 961 -472 1039 -471
rect 1059 -472 1158 -471
rect 138 -474 619 -473
rect 723 -474 815 -473
rect 828 -474 1060 -473
rect 215 -476 689 -475
rect 828 -476 1235 -475
rect 107 -478 1235 -477
rect 219 -480 640 -479
rect 835 -480 962 -479
rect 975 -480 1025 -479
rect 338 -482 815 -481
rect 912 -482 976 -481
rect 338 -484 346 -483
rect 380 -484 395 -483
rect 548 -484 913 -483
rect 149 -486 381 -485
rect 457 -486 549 -485
rect 597 -486 941 -485
rect 149 -488 178 -487
rect 310 -488 346 -487
rect 457 -488 647 -487
rect 765 -488 836 -487
rect 177 -490 213 -489
rect 310 -490 416 -489
rect 646 -490 801 -489
rect 212 -492 241 -491
rect 373 -492 766 -491
rect 219 -494 241 -493
rect 320 -494 374 -493
rect 9 -505 283 -504
rect 317 -505 416 -504
rect 450 -505 864 -504
rect 873 -505 983 -504
rect 1136 -505 1193 -504
rect 1269 -505 1273 -504
rect 1468 -505 1557 -504
rect 1710 -505 1760 -504
rect 23 -507 52 -506
rect 58 -507 101 -506
rect 103 -507 325 -506
rect 359 -507 409 -506
rect 450 -507 570 -506
rect 583 -507 608 -506
rect 618 -507 983 -506
rect 1129 -507 1137 -506
rect 1269 -507 1305 -506
rect 1486 -507 1522 -506
rect 1528 -507 1767 -506
rect 37 -509 185 -508
rect 194 -509 1165 -508
rect 1500 -509 1504 -508
rect 1514 -509 1739 -508
rect 61 -511 1263 -510
rect 1458 -511 1515 -510
rect 79 -513 325 -512
rect 362 -513 752 -512
rect 758 -513 1361 -512
rect 1451 -513 1459 -512
rect 1500 -513 1508 -512
rect 72 -515 80 -514
rect 103 -515 409 -514
rect 453 -515 598 -514
rect 618 -515 1074 -514
rect 1122 -515 1130 -514
rect 1150 -515 1165 -514
rect 1325 -515 1361 -514
rect 1430 -515 1452 -514
rect 72 -517 115 -516
rect 128 -517 220 -516
rect 222 -517 689 -516
rect 709 -517 1221 -516
rect 1402 -517 1431 -516
rect 107 -519 122 -518
rect 128 -519 395 -518
rect 401 -519 475 -518
rect 481 -519 801 -518
rect 824 -519 1249 -518
rect 114 -521 538 -520
rect 548 -521 570 -520
rect 583 -521 962 -520
rect 1052 -521 1123 -520
rect 1185 -521 1221 -520
rect 121 -523 339 -522
rect 341 -523 549 -522
rect 590 -523 829 -522
rect 831 -523 1151 -522
rect 1199 -523 1326 -522
rect 138 -525 1445 -524
rect 152 -527 587 -526
rect 593 -527 1074 -526
rect 1080 -527 1403 -526
rect 1416 -527 1445 -526
rect 156 -529 188 -528
rect 243 -529 360 -528
rect 373 -529 535 -528
rect 593 -529 1200 -528
rect 1213 -529 1249 -528
rect 1395 -529 1417 -528
rect 44 -531 535 -530
rect 597 -531 815 -530
rect 828 -531 836 -530
rect 842 -531 1263 -530
rect 1367 -531 1396 -530
rect 44 -533 902 -532
rect 947 -533 951 -532
rect 961 -533 1067 -532
rect 1178 -533 1214 -532
rect 1332 -533 1368 -532
rect 93 -535 157 -534
rect 177 -535 199 -534
rect 268 -535 297 -534
rect 317 -535 766 -534
rect 779 -535 801 -534
rect 842 -535 1438 -534
rect 93 -537 143 -536
rect 180 -537 206 -536
rect 268 -537 521 -536
rect 530 -537 731 -536
rect 761 -537 1186 -536
rect 1318 -537 1333 -536
rect 1409 -537 1438 -536
rect 65 -539 521 -538
rect 530 -539 647 -538
rect 667 -539 713 -538
rect 716 -539 759 -538
rect 765 -539 1340 -538
rect 1388 -539 1410 -538
rect 65 -541 136 -540
rect 142 -541 458 -540
rect 460 -541 1424 -540
rect 135 -543 150 -542
rect 191 -543 458 -542
rect 464 -543 650 -542
rect 653 -543 668 -542
rect 677 -543 717 -542
rect 723 -543 815 -542
rect 915 -543 1389 -542
rect 149 -545 311 -544
rect 352 -545 654 -544
rect 681 -545 724 -544
rect 730 -545 794 -544
rect 947 -545 990 -544
rect 1017 -545 1081 -544
rect 1157 -545 1179 -544
rect 1297 -545 1319 -544
rect 1339 -545 1382 -544
rect 198 -547 255 -546
rect 275 -547 283 -546
rect 310 -547 507 -546
rect 516 -547 710 -546
rect 779 -547 1473 -546
rect 30 -549 507 -548
rect 516 -549 1158 -548
rect 1297 -549 1347 -548
rect 1472 -549 1480 -548
rect 163 -551 276 -550
rect 366 -551 374 -550
rect 380 -551 402 -550
rect 464 -551 696 -550
rect 786 -551 836 -550
rect 954 -551 1018 -550
rect 1038 -551 1067 -550
rect 1283 -551 1480 -550
rect 163 -553 262 -552
rect 366 -553 486 -552
rect 492 -553 892 -552
rect 919 -553 1039 -552
rect 1052 -553 1312 -552
rect 1346 -553 1466 -552
rect 205 -555 248 -554
rect 254 -555 577 -554
rect 625 -555 853 -554
rect 891 -555 1536 -554
rect 30 -557 248 -556
rect 261 -557 479 -556
rect 485 -557 612 -556
rect 625 -557 738 -556
rect 786 -557 1004 -556
rect 1241 -557 1284 -556
rect 1290 -557 1312 -556
rect 170 -559 612 -558
rect 632 -559 997 -558
rect 1087 -559 1291 -558
rect 170 -561 430 -560
rect 436 -561 479 -560
rect 492 -561 857 -560
rect 919 -561 1060 -560
rect 1087 -561 1228 -560
rect 226 -563 353 -562
rect 387 -563 395 -562
rect 418 -563 1242 -562
rect 226 -565 444 -564
rect 471 -565 563 -564
rect 576 -565 1109 -564
rect 1195 -565 1228 -564
rect 233 -567 444 -566
rect 495 -567 969 -566
rect 1055 -567 1109 -566
rect 303 -569 388 -568
rect 523 -569 1382 -568
rect 240 -571 304 -570
rect 331 -571 437 -570
rect 527 -571 1424 -570
rect 212 -573 332 -572
rect 527 -573 1277 -572
rect 212 -575 423 -574
rect 562 -575 773 -574
rect 793 -575 885 -574
rect 898 -575 1060 -574
rect 1255 -575 1277 -574
rect 240 -577 290 -576
rect 338 -577 423 -576
rect 635 -577 1095 -576
rect 1234 -577 1256 -576
rect 1503 -577 1508 -576
rect 289 -579 300 -578
rect 579 -579 636 -578
rect 639 -579 752 -578
rect 772 -579 850 -578
rect 856 -579 934 -578
rect 968 -579 976 -578
rect 1094 -579 1116 -578
rect 1206 -579 1235 -578
rect 639 -581 675 -580
rect 688 -581 808 -580
rect 849 -581 997 -580
rect 1101 -581 1116 -580
rect 1143 -581 1207 -580
rect 555 -583 675 -582
rect 698 -583 1004 -582
rect 1031 -583 1102 -582
rect 51 -585 699 -584
rect 702 -585 808 -584
rect 866 -585 1144 -584
rect 513 -587 556 -586
rect 660 -587 682 -586
rect 702 -587 846 -586
rect 877 -587 976 -586
rect 1024 -587 1032 -586
rect 86 -589 661 -588
rect 737 -589 745 -588
rect 870 -589 878 -588
rect 884 -589 895 -588
rect 926 -589 955 -588
rect 1010 -589 1025 -588
rect 86 -591 601 -590
rect 744 -591 822 -590
rect 912 -591 927 -590
rect 940 -591 1011 -590
rect 453 -593 941 -592
rect 821 -595 1487 -594
rect 912 -597 1375 -596
rect 1353 -599 1375 -598
rect 110 -601 1354 -600
rect 9 -612 454 -611
rect 492 -612 591 -611
rect 604 -612 633 -611
rect 653 -612 657 -611
rect 674 -612 710 -611
rect 761 -612 948 -611
rect 1017 -612 1053 -611
rect 1339 -612 1529 -611
rect 1535 -612 1788 -611
rect 9 -614 269 -613
rect 303 -614 318 -613
rect 320 -614 381 -613
rect 408 -614 713 -613
rect 786 -614 822 -613
rect 824 -614 962 -613
rect 1241 -614 1340 -613
rect 1346 -614 1620 -613
rect 1668 -614 1802 -613
rect 16 -616 94 -615
rect 114 -616 185 -615
rect 233 -616 262 -615
rect 303 -616 325 -615
rect 362 -616 650 -615
rect 653 -616 668 -615
rect 677 -616 1431 -615
rect 1437 -616 1592 -615
rect 1738 -616 1823 -615
rect 30 -618 59 -617
rect 72 -618 458 -617
rect 544 -618 612 -617
rect 660 -618 962 -617
rect 1087 -618 1347 -617
rect 1388 -618 1536 -617
rect 1556 -618 1658 -617
rect 1759 -618 1795 -617
rect 30 -620 118 -619
rect 145 -620 269 -619
rect 352 -620 458 -619
rect 569 -620 591 -619
rect 604 -620 717 -619
rect 786 -620 1000 -619
rect 1157 -620 1242 -619
rect 1325 -620 1438 -619
rect 1444 -620 1578 -619
rect 1766 -620 1858 -619
rect 37 -622 871 -621
rect 873 -622 1389 -621
rect 1409 -622 1543 -621
rect 44 -624 97 -623
rect 114 -624 1263 -623
rect 1290 -624 1410 -623
rect 1416 -624 1564 -623
rect 44 -626 500 -625
rect 667 -626 703 -625
rect 709 -626 1571 -625
rect 51 -628 73 -627
rect 79 -628 83 -627
rect 128 -628 353 -627
rect 373 -628 430 -627
rect 499 -628 507 -627
rect 681 -628 703 -627
rect 793 -628 913 -627
rect 933 -628 1193 -627
rect 1206 -628 1263 -627
rect 1269 -628 1417 -627
rect 1423 -628 1557 -627
rect 51 -630 104 -629
rect 128 -630 136 -629
rect 149 -630 325 -629
rect 373 -630 384 -629
rect 408 -630 423 -629
rect 429 -630 472 -629
rect 509 -630 1207 -629
rect 1227 -630 1326 -629
rect 1451 -630 1585 -629
rect 58 -632 66 -631
rect 79 -632 108 -631
rect 135 -632 1634 -631
rect 65 -634 143 -633
rect 149 -634 213 -633
rect 243 -634 444 -633
rect 681 -634 752 -633
rect 796 -634 1466 -633
rect 1472 -634 1550 -633
rect 142 -636 766 -635
rect 800 -636 822 -635
rect 842 -636 1102 -635
rect 1108 -636 1158 -635
rect 1178 -636 1270 -635
rect 1353 -636 1473 -635
rect 1479 -636 1613 -635
rect 100 -638 1109 -637
rect 1129 -638 1228 -637
rect 1360 -638 1466 -637
rect 1468 -638 1480 -637
rect 1486 -638 1627 -637
rect 100 -640 192 -639
rect 212 -640 468 -639
rect 562 -640 801 -639
rect 849 -640 1515 -639
rect 156 -642 892 -641
rect 894 -642 1403 -641
rect 1458 -642 1599 -641
rect 156 -644 402 -643
rect 415 -644 514 -643
rect 562 -644 731 -643
rect 737 -644 766 -643
rect 782 -644 1459 -643
rect 1493 -644 1641 -643
rect 163 -646 493 -645
rect 513 -646 549 -645
rect 569 -646 843 -645
rect 845 -646 1515 -645
rect 163 -648 647 -647
rect 660 -648 738 -647
rect 852 -648 1214 -647
rect 1255 -648 1361 -647
rect 1374 -648 1487 -647
rect 1500 -648 1662 -647
rect 170 -650 528 -649
rect 593 -650 850 -649
rect 863 -650 1431 -649
rect 1507 -650 1648 -649
rect 170 -652 1291 -651
rect 1297 -652 1508 -651
rect 173 -654 619 -653
rect 646 -654 720 -653
rect 723 -654 752 -653
rect 870 -654 923 -653
rect 989 -654 1088 -653
rect 1115 -654 1214 -653
rect 1248 -654 1256 -653
rect 1311 -654 1375 -653
rect 1381 -654 1494 -653
rect 187 -656 1445 -655
rect 191 -658 199 -657
rect 236 -658 416 -657
rect 422 -658 531 -657
rect 635 -658 990 -657
rect 996 -658 1102 -657
rect 1136 -658 1354 -657
rect 1367 -658 1501 -657
rect 198 -660 339 -659
rect 366 -660 472 -659
rect 520 -660 549 -659
rect 656 -660 724 -659
rect 730 -660 745 -659
rect 877 -660 948 -659
rect 1024 -660 1137 -659
rect 1164 -660 1249 -659
rect 1276 -660 1382 -659
rect 61 -662 1025 -661
rect 1031 -662 1179 -661
rect 1185 -662 1277 -661
rect 1283 -662 1368 -661
rect 236 -664 584 -663
rect 625 -664 745 -663
rect 828 -664 878 -663
rect 898 -664 934 -663
rect 1038 -664 1298 -663
rect 1318 -664 1403 -663
rect 240 -666 367 -665
rect 387 -666 619 -665
rect 625 -666 1021 -665
rect 1059 -666 1193 -665
rect 1199 -666 1452 -665
rect 240 -668 832 -667
rect 856 -668 1060 -667
rect 1066 -668 1116 -667
rect 1171 -668 1284 -667
rect 152 -670 857 -669
rect 908 -670 1606 -669
rect 254 -672 867 -671
rect 926 -672 1032 -671
rect 1045 -672 1200 -671
rect 1234 -672 1319 -671
rect 261 -674 346 -673
rect 387 -674 601 -673
rect 688 -674 864 -673
rect 884 -674 927 -673
rect 954 -674 1046 -673
rect 1073 -674 1186 -673
rect 331 -676 339 -675
rect 345 -676 482 -675
rect 520 -676 542 -675
rect 586 -676 899 -675
rect 940 -676 1074 -675
rect 1080 -676 1130 -675
rect 1143 -676 1172 -675
rect 275 -678 332 -677
rect 401 -678 640 -677
rect 691 -678 916 -677
rect 975 -678 1039 -677
rect 1150 -678 1235 -677
rect 275 -680 395 -679
rect 432 -680 1312 -679
rect 394 -682 780 -681
rect 793 -682 941 -681
rect 982 -682 1081 -681
rect 247 -684 780 -683
rect 814 -684 983 -683
rect 1003 -684 1151 -683
rect 247 -686 290 -685
rect 443 -686 577 -685
rect 597 -686 640 -685
rect 695 -686 1123 -685
rect 289 -688 297 -687
rect 464 -688 528 -687
rect 541 -688 612 -687
rect 695 -688 972 -687
rect 1010 -688 1067 -687
rect 1122 -688 1396 -687
rect 23 -690 465 -689
rect 555 -690 577 -689
rect 597 -690 1144 -689
rect 1304 -690 1396 -689
rect 23 -692 311 -691
rect 698 -692 1424 -691
rect 121 -694 311 -693
rect 740 -694 1165 -693
rect 1220 -694 1305 -693
rect 121 -696 451 -695
rect 772 -696 976 -695
rect 1094 -696 1221 -695
rect 219 -698 297 -697
rect 450 -698 479 -697
rect 758 -698 773 -697
rect 807 -698 815 -697
rect 828 -698 1522 -697
rect 86 -700 220 -699
rect 254 -700 479 -699
rect 506 -700 1522 -699
rect 86 -702 227 -701
rect 621 -702 808 -701
rect 835 -702 955 -701
rect 968 -702 1095 -701
rect 226 -704 759 -703
rect 884 -704 902 -703
rect 905 -704 1004 -703
rect 359 -706 836 -705
rect 919 -706 1011 -705
rect 359 -708 486 -707
rect 485 -710 1672 -709
rect 9 -721 94 -720
rect 114 -721 1784 -720
rect 1787 -721 1893 -720
rect 9 -723 423 -722
rect 439 -723 556 -722
rect 562 -723 650 -722
rect 709 -723 1298 -722
rect 1458 -723 1844 -722
rect 1857 -723 1886 -722
rect 16 -725 118 -724
rect 121 -725 125 -724
rect 128 -725 139 -724
rect 170 -725 181 -724
rect 254 -725 258 -724
rect 303 -725 307 -724
rect 422 -725 720 -724
rect 723 -725 738 -724
rect 740 -725 1592 -724
rect 1605 -725 1739 -724
rect 1801 -725 1858 -724
rect 37 -727 234 -726
rect 254 -727 528 -726
rect 548 -727 563 -726
rect 586 -727 997 -726
rect 999 -727 1564 -726
rect 1577 -727 1732 -726
rect 1822 -727 1851 -726
rect 37 -729 573 -728
rect 597 -729 1452 -728
rect 1486 -729 1676 -728
rect 1794 -729 1823 -728
rect 58 -731 545 -730
rect 555 -731 1592 -730
rect 1612 -731 1760 -730
rect 30 -733 59 -732
rect 79 -733 115 -732
rect 121 -733 234 -732
rect 268 -733 528 -732
rect 618 -733 1298 -732
rect 1360 -733 1452 -732
rect 1493 -733 1606 -732
rect 1626 -733 1788 -732
rect 30 -735 101 -734
rect 135 -735 146 -734
rect 170 -735 178 -734
rect 201 -735 1564 -734
rect 1570 -735 1578 -734
rect 1584 -735 1767 -734
rect 93 -737 185 -736
rect 268 -737 416 -736
rect 443 -737 507 -736
rect 520 -737 542 -736
rect 614 -737 619 -736
rect 621 -737 1487 -736
rect 1542 -737 1690 -736
rect 65 -739 521 -738
rect 628 -739 731 -738
rect 779 -739 1473 -738
rect 1479 -739 1585 -738
rect 1633 -739 1795 -738
rect 65 -741 517 -740
rect 632 -741 731 -740
rect 758 -741 1473 -740
rect 1549 -741 1746 -740
rect 100 -743 290 -742
rect 303 -743 388 -742
rect 443 -743 486 -742
rect 495 -743 829 -742
rect 831 -743 1669 -742
rect 1671 -743 1718 -742
rect 107 -745 185 -744
rect 275 -745 416 -744
rect 450 -745 486 -744
rect 590 -745 633 -744
rect 674 -745 710 -744
rect 712 -745 1802 -744
rect 107 -747 472 -746
rect 478 -747 976 -746
rect 1034 -747 1830 -746
rect 135 -749 500 -748
rect 653 -749 675 -748
rect 681 -749 738 -748
rect 779 -749 1711 -748
rect 173 -751 458 -750
rect 464 -751 1074 -750
rect 1143 -751 1697 -750
rect 96 -753 465 -752
rect 478 -753 668 -752
rect 716 -753 1200 -752
rect 1234 -753 1361 -752
rect 1367 -753 1459 -752
rect 1465 -753 1543 -752
rect 1549 -753 1599 -752
rect 1633 -753 1662 -752
rect 156 -755 458 -754
rect 467 -755 668 -754
rect 723 -755 941 -754
rect 1045 -755 1144 -754
rect 1178 -755 1200 -754
rect 1234 -755 1305 -754
rect 1339 -755 1480 -754
rect 1556 -755 1704 -754
rect 51 -757 157 -756
rect 275 -757 283 -756
rect 289 -757 601 -756
rect 639 -757 682 -756
rect 782 -757 906 -756
rect 919 -757 962 -756
rect 1073 -757 1221 -756
rect 1241 -757 1368 -756
rect 1381 -757 1494 -756
rect 1556 -757 1781 -756
rect 282 -759 318 -758
rect 324 -759 717 -758
rect 793 -759 1410 -758
rect 1444 -759 1613 -758
rect 1640 -759 1774 -758
rect 296 -761 829 -760
rect 835 -761 1046 -760
rect 1080 -761 1179 -760
rect 1195 -761 1683 -760
rect 324 -763 909 -762
rect 922 -763 1753 -762
rect 345 -765 622 -764
rect 772 -765 794 -764
rect 800 -765 804 -764
rect 807 -765 941 -764
rect 1052 -765 1081 -764
rect 1094 -765 1221 -764
rect 1262 -765 1340 -764
rect 1388 -765 1599 -764
rect 1647 -765 1809 -764
rect 345 -767 367 -766
rect 373 -767 962 -766
rect 1136 -767 1242 -766
rect 1269 -767 1382 -766
rect 1402 -767 1571 -766
rect 310 -769 367 -768
rect 373 -769 402 -768
rect 436 -769 472 -768
rect 492 -769 500 -768
rect 569 -769 640 -768
rect 695 -769 773 -768
rect 800 -769 871 -768
rect 884 -769 1627 -768
rect 54 -771 311 -770
rect 401 -771 409 -770
rect 450 -771 920 -770
rect 933 -771 1095 -770
rect 1157 -771 1263 -770
rect 1276 -771 1389 -770
rect 1430 -771 1648 -770
rect 142 -773 934 -772
rect 954 -773 1053 -772
rect 1101 -773 1158 -772
rect 1283 -773 1445 -772
rect 1465 -773 1529 -772
rect 142 -775 199 -774
rect 359 -775 409 -774
rect 492 -775 535 -774
rect 576 -775 654 -774
rect 803 -775 871 -774
rect 898 -775 1305 -774
rect 1318 -775 1403 -774
rect 1521 -775 1641 -774
rect 44 -777 577 -776
rect 604 -777 808 -776
rect 814 -777 836 -776
rect 842 -777 1354 -776
rect 1437 -777 1522 -776
rect 177 -779 899 -778
rect 901 -779 1620 -778
rect 198 -781 360 -780
rect 534 -781 689 -780
rect 824 -781 1515 -780
rect 548 -783 843 -782
rect 845 -783 1725 -782
rect 583 -785 605 -784
rect 611 -785 696 -784
rect 782 -785 1515 -784
rect 163 -787 612 -786
rect 625 -787 815 -786
rect 849 -787 1018 -786
rect 1020 -787 1438 -786
rect 1507 -787 1620 -786
rect 163 -789 1424 -788
rect 583 -791 591 -790
rect 625 -791 1662 -790
rect 646 -793 885 -792
rect 912 -793 955 -792
rect 1010 -793 1270 -792
rect 1290 -793 1837 -792
rect 212 -795 1011 -794
rect 1031 -795 1137 -794
rect 1185 -795 1284 -794
rect 1311 -795 1424 -794
rect 296 -797 1032 -796
rect 1038 -797 1102 -796
rect 1108 -797 1291 -796
rect 1325 -797 1410 -796
rect 1416 -797 1508 -796
rect 166 -799 1326 -798
rect 1332 -799 1354 -798
rect 1374 -799 1417 -798
rect 429 -801 647 -800
rect 744 -801 850 -800
rect 926 -801 1018 -800
rect 1087 -801 1186 -800
rect 1192 -801 1312 -800
rect 1346 -801 1431 -800
rect 79 -803 1088 -802
rect 1115 -803 1277 -802
rect 352 -805 430 -804
rect 509 -805 1039 -804
rect 1066 -805 1116 -804
rect 1213 -805 1319 -804
rect 338 -807 353 -806
rect 691 -807 927 -806
rect 947 -807 1067 -806
rect 1227 -807 1333 -806
rect 82 -809 339 -808
rect 744 -809 752 -808
rect 761 -809 1214 -808
rect 1248 -809 1375 -808
rect 702 -811 752 -810
rect 761 -811 1207 -810
rect 1255 -811 1529 -810
rect 789 -813 948 -812
rect 971 -813 1347 -812
rect 821 -815 913 -814
rect 982 -815 1207 -814
rect 821 -817 1501 -816
rect 863 -819 983 -818
rect 989 -819 1109 -818
rect 1129 -819 1249 -818
rect 1395 -819 1501 -818
rect 765 -821 864 -820
rect 989 -821 1655 -820
rect 226 -823 766 -822
rect 1003 -823 1130 -822
rect 1150 -823 1228 -822
rect 226 -825 262 -824
rect 1024 -825 1256 -824
rect 240 -827 1004 -826
rect 1150 -827 1165 -826
rect 1171 -827 1396 -826
rect 72 -829 1165 -828
rect 1192 -829 1655 -828
rect 72 -831 150 -830
rect 240 -831 248 -830
rect 261 -831 332 -830
rect 891 -831 1025 -830
rect 1059 -831 1172 -830
rect 44 -833 150 -832
rect 205 -833 248 -832
rect 331 -833 381 -832
rect 877 -833 892 -832
rect 968 -833 1060 -832
rect 191 -835 206 -834
rect 380 -835 514 -834
rect 660 -835 878 -834
rect 128 -837 192 -836
rect 212 -837 514 -836
rect 579 -837 661 -836
rect 856 -837 969 -836
rect 786 -839 857 -838
rect 786 -841 1536 -840
rect 1122 -843 1536 -842
rect 558 -845 1123 -844
rect 86 -847 559 -846
rect 86 -849 220 -848
rect 23 -851 220 -850
rect 23 -853 395 -852
rect 187 -855 395 -854
rect 2 -866 69 -865
rect 86 -866 90 -865
rect 110 -866 1235 -865
rect 1591 -866 1595 -865
rect 1724 -866 1865 -865
rect 1885 -866 1914 -865
rect 37 -868 80 -867
rect 86 -868 206 -867
rect 261 -868 265 -867
rect 310 -868 944 -867
rect 1006 -868 1767 -867
rect 1780 -868 1823 -867
rect 1829 -868 1942 -867
rect 30 -870 80 -869
rect 114 -870 122 -869
rect 135 -870 514 -869
rect 516 -870 1669 -869
rect 1703 -870 1767 -869
rect 1787 -870 1830 -869
rect 1836 -870 1949 -869
rect 30 -872 227 -871
rect 261 -872 276 -871
rect 310 -872 451 -871
rect 460 -872 1921 -871
rect 37 -874 73 -873
rect 121 -874 129 -873
rect 156 -874 822 -873
rect 828 -874 1613 -873
rect 1633 -874 1886 -873
rect 1892 -874 1956 -873
rect 51 -876 115 -875
rect 163 -876 248 -875
rect 275 -876 304 -875
rect 338 -876 437 -875
rect 450 -876 748 -875
rect 779 -876 1067 -875
rect 1083 -876 1732 -875
rect 1759 -876 1872 -875
rect 47 -878 1067 -877
rect 1108 -878 1112 -877
rect 1153 -878 1676 -877
rect 1717 -878 1788 -877
rect 1801 -878 1935 -877
rect 51 -880 94 -879
rect 177 -880 1025 -879
rect 1031 -880 1599 -879
rect 1619 -880 1676 -879
rect 1752 -880 1760 -879
rect 1843 -880 1907 -879
rect 65 -882 549 -881
rect 572 -882 1326 -881
rect 1353 -882 1599 -881
rect 1633 -882 1879 -881
rect 65 -884 1014 -883
rect 1031 -884 1529 -883
rect 1556 -884 1613 -883
rect 1654 -884 1725 -883
rect 1794 -884 1844 -883
rect 1850 -884 1882 -883
rect 72 -886 234 -885
rect 247 -886 430 -885
rect 492 -886 654 -885
rect 684 -886 829 -885
rect 915 -886 1326 -885
rect 1360 -886 1620 -885
rect 1661 -886 1718 -885
rect 1738 -886 1795 -885
rect 1857 -886 1893 -885
rect 93 -888 164 -887
rect 177 -888 682 -887
rect 688 -888 1480 -887
rect 1500 -888 1557 -887
rect 1577 -888 1837 -887
rect 128 -890 234 -889
rect 268 -890 437 -889
rect 492 -890 563 -889
rect 576 -890 878 -889
rect 919 -890 1074 -889
rect 1108 -890 1179 -889
rect 1297 -890 1354 -889
rect 1381 -890 1655 -889
rect 1668 -890 1746 -889
rect 1808 -890 1858 -889
rect 156 -892 1361 -891
rect 1430 -892 1480 -891
rect 1521 -892 1578 -891
rect 1591 -892 1711 -891
rect 180 -894 381 -893
rect 387 -894 692 -893
rect 705 -894 962 -893
rect 985 -894 1781 -893
rect 58 -896 381 -895
rect 429 -896 591 -895
rect 604 -896 654 -895
rect 688 -896 990 -895
rect 1003 -896 1025 -895
rect 1034 -896 1445 -895
rect 1451 -896 1501 -895
rect 1521 -896 1585 -895
rect 1605 -896 1662 -895
rect 1689 -896 1739 -895
rect 187 -898 598 -897
rect 604 -898 1564 -897
rect 1640 -898 1690 -897
rect 1696 -898 1753 -897
rect 191 -900 864 -899
rect 877 -900 1193 -899
rect 1374 -900 1431 -899
rect 1465 -900 1802 -899
rect 198 -902 556 -901
rect 583 -902 675 -901
rect 723 -902 1235 -901
rect 1402 -902 1445 -901
rect 1465 -902 1543 -901
rect 1549 -902 1851 -901
rect 170 -904 199 -903
rect 201 -904 283 -903
rect 338 -904 444 -903
rect 478 -904 598 -903
rect 618 -904 717 -903
rect 726 -904 1697 -903
rect 170 -906 325 -905
rect 394 -906 444 -905
rect 485 -906 563 -905
rect 586 -906 1046 -905
rect 1059 -906 1529 -905
rect 1535 -906 1606 -905
rect 1647 -906 1711 -905
rect 184 -908 395 -907
rect 408 -908 486 -907
rect 495 -908 780 -907
rect 782 -908 1704 -907
rect 184 -910 332 -909
rect 506 -910 549 -909
rect 590 -910 647 -909
rect 674 -910 1039 -909
rect 1041 -910 1571 -909
rect 205 -912 220 -911
rect 240 -912 325 -911
rect 422 -912 507 -911
rect 513 -912 850 -911
rect 856 -912 1382 -911
rect 1409 -912 1452 -911
rect 1472 -912 1746 -911
rect 212 -914 479 -913
rect 527 -914 559 -913
rect 618 -914 825 -913
rect 831 -914 1375 -913
rect 1395 -914 1410 -913
rect 1416 -914 1571 -913
rect 142 -916 213 -915
rect 240 -916 346 -915
rect 415 -916 423 -915
rect 499 -916 528 -915
rect 534 -916 584 -915
rect 621 -916 1823 -915
rect 226 -918 535 -917
rect 537 -918 1207 -917
rect 1255 -918 1417 -917
rect 1423 -918 1550 -917
rect 1563 -918 1900 -917
rect 268 -920 601 -919
rect 625 -920 752 -919
rect 758 -920 1046 -919
rect 1059 -920 1298 -919
rect 1318 -920 1424 -919
rect 1486 -920 1536 -919
rect 282 -922 360 -921
rect 415 -922 1095 -921
rect 1115 -922 1256 -921
rect 1276 -922 1319 -921
rect 1346 -922 1403 -921
rect 1486 -922 1917 -921
rect 289 -924 332 -923
rect 359 -924 1784 -923
rect 289 -926 353 -925
rect 499 -926 755 -925
rect 758 -926 773 -925
rect 775 -926 1585 -925
rect 254 -928 353 -927
rect 541 -928 577 -927
rect 625 -928 661 -927
rect 709 -928 850 -927
rect 856 -928 976 -927
rect 1017 -928 1074 -927
rect 1087 -928 1116 -927
rect 1129 -928 1179 -927
rect 1276 -928 1389 -927
rect 1493 -928 1543 -927
rect 58 -930 542 -929
rect 639 -930 1018 -929
rect 1052 -930 1088 -929
rect 1094 -930 1102 -929
rect 1122 -930 1130 -929
rect 1164 -930 1193 -929
rect 1283 -930 1347 -929
rect 1367 -930 1473 -929
rect 1493 -930 1683 -929
rect 254 -932 570 -931
rect 639 -932 801 -931
rect 814 -932 1102 -931
rect 1171 -932 1207 -931
rect 1241 -932 1284 -931
rect 1304 -932 1368 -931
rect 1507 -932 1641 -931
rect 1682 -932 1819 -931
rect 142 -934 815 -933
rect 821 -934 843 -933
rect 863 -934 913 -933
rect 922 -934 1732 -933
rect 296 -936 409 -935
rect 520 -936 710 -935
rect 716 -936 731 -935
rect 740 -936 1809 -935
rect 296 -938 472 -937
rect 544 -938 570 -937
rect 646 -938 906 -937
rect 922 -938 1928 -937
rect 166 -940 906 -939
rect 947 -940 990 -939
rect 1003 -940 1165 -939
rect 1311 -940 1389 -939
rect 1458 -940 1508 -939
rect 1594 -940 1648 -939
rect 317 -942 346 -941
rect 401 -942 472 -941
rect 660 -942 941 -941
rect 947 -942 983 -941
rect 1062 -942 1515 -941
rect 149 -944 318 -943
rect 401 -944 458 -943
rect 464 -944 521 -943
rect 702 -944 1242 -943
rect 1262 -944 1312 -943
rect 100 -946 150 -945
rect 373 -946 703 -945
rect 730 -946 1011 -945
rect 1143 -946 1172 -945
rect 1213 -946 1459 -945
rect 9 -948 101 -947
rect 107 -948 374 -947
rect 390 -948 465 -947
rect 744 -948 787 -947
rect 789 -948 843 -947
rect 891 -948 1053 -947
rect 1080 -948 1144 -947
rect 1157 -948 1305 -947
rect 9 -950 24 -949
rect 44 -950 108 -949
rect 135 -950 458 -949
rect 611 -950 787 -949
rect 800 -950 941 -949
rect 954 -950 976 -949
rect 1010 -950 1774 -949
rect 23 -952 195 -951
rect 611 -952 696 -951
rect 744 -952 1291 -951
rect 667 -954 696 -953
rect 761 -954 1515 -953
rect 667 -956 871 -955
rect 884 -956 955 -955
rect 961 -956 997 -955
rect 1034 -956 1774 -955
rect 765 -958 983 -957
rect 996 -958 1039 -957
rect 1080 -958 1816 -957
rect 737 -960 766 -959
rect 772 -960 1270 -959
rect 807 -962 892 -961
rect 1157 -962 1396 -961
rect 793 -964 808 -963
rect 835 -964 871 -963
rect 884 -964 899 -963
rect 1185 -964 1214 -963
rect 1227 -964 1270 -963
rect 54 -966 836 -965
rect 1150 -966 1186 -965
rect 1248 -966 1291 -965
rect 236 -968 1249 -967
rect 1262 -968 1627 -967
rect 439 -970 899 -969
rect 1437 -970 1627 -969
rect 793 -972 1161 -971
rect 1332 -972 1438 -971
rect 1199 -974 1333 -973
rect 628 -976 1200 -975
rect 47 -987 703 -986
rect 733 -987 773 -986
rect 775 -987 822 -986
rect 866 -987 1424 -986
rect 1745 -987 1900 -986
rect 1927 -987 1977 -986
rect 58 -989 454 -988
rect 457 -989 538 -988
rect 541 -989 626 -988
rect 656 -989 1417 -988
rect 1710 -989 1746 -988
rect 1867 -989 1893 -988
rect 1927 -989 1935 -988
rect 1941 -989 1963 -988
rect 58 -991 171 -990
rect 240 -991 685 -990
rect 709 -991 822 -990
rect 870 -991 916 -990
rect 919 -991 1431 -990
rect 1710 -991 1767 -990
rect 1878 -991 1907 -990
rect 1948 -991 1970 -990
rect 68 -993 395 -992
rect 443 -993 458 -992
rect 485 -993 605 -992
rect 625 -993 1438 -992
rect 1584 -993 1879 -992
rect 1948 -993 1956 -992
rect 30 -995 395 -994
rect 485 -995 619 -994
rect 674 -995 710 -994
rect 716 -995 773 -994
rect 779 -995 1417 -994
rect 1493 -995 1585 -994
rect 30 -997 52 -996
rect 72 -997 391 -996
rect 513 -997 605 -996
rect 667 -997 717 -996
rect 737 -997 759 -996
rect 761 -997 1725 -996
rect 51 -999 409 -998
rect 478 -999 668 -998
rect 674 -999 1193 -998
rect 1241 -999 1245 -998
rect 1276 -999 1424 -998
rect 1493 -999 1501 -998
rect 1724 -999 1886 -998
rect 72 -1001 636 -1000
rect 681 -1001 1179 -1000
rect 1241 -1001 1270 -1000
rect 1276 -1001 1291 -1000
rect 1409 -1001 1431 -1000
rect 1500 -1001 1508 -1000
rect 82 -1003 1018 -1002
rect 1020 -1003 1256 -1002
rect 1367 -1003 1410 -1002
rect 1507 -1003 1515 -1002
rect 86 -1005 146 -1004
rect 149 -1005 171 -1004
rect 240 -1005 402 -1004
rect 408 -1005 493 -1004
rect 513 -1005 612 -1004
rect 646 -1005 1179 -1004
rect 1244 -1005 1270 -1004
rect 1514 -1005 1571 -1004
rect 9 -1007 87 -1006
rect 93 -1007 220 -1006
rect 282 -1007 727 -1006
rect 737 -1007 1438 -1006
rect 1535 -1007 1571 -1006
rect 9 -1009 227 -1008
rect 282 -1009 437 -1008
rect 478 -1009 780 -1008
rect 786 -1009 958 -1008
rect 968 -1009 1291 -1008
rect 1535 -1009 1599 -1008
rect 79 -1011 150 -1010
rect 156 -1011 444 -1010
rect 492 -1011 731 -1010
rect 747 -1011 1459 -1010
rect 1598 -1011 1634 -1010
rect 79 -1013 1235 -1012
rect 1255 -1013 1298 -1012
rect 1451 -1013 1459 -1012
rect 68 -1015 1452 -1014
rect 96 -1017 759 -1016
rect 863 -1017 871 -1016
rect 891 -1017 1368 -1016
rect 107 -1019 129 -1018
rect 142 -1019 160 -1018
rect 226 -1019 661 -1018
rect 681 -1019 1529 -1018
rect 128 -1021 311 -1020
rect 345 -1021 437 -1020
rect 506 -1021 969 -1020
rect 982 -1021 1865 -1020
rect 142 -1023 192 -1022
rect 268 -1023 787 -1022
rect 842 -1023 892 -1022
rect 894 -1023 899 -1022
rect 912 -1023 1473 -1022
rect 37 -1025 269 -1024
rect 296 -1025 535 -1024
rect 565 -1025 612 -1024
rect 632 -1025 661 -1024
rect 702 -1025 731 -1024
rect 751 -1025 1774 -1024
rect 37 -1027 472 -1026
rect 499 -1027 535 -1026
rect 569 -1027 1084 -1026
rect 1108 -1027 1158 -1026
rect 1160 -1027 1851 -1026
rect 156 -1029 1063 -1028
rect 1108 -1029 1123 -1028
rect 1136 -1029 1529 -1028
rect 1773 -1029 1921 -1028
rect 191 -1031 237 -1030
rect 303 -1031 346 -1030
rect 387 -1031 563 -1030
rect 579 -1031 1634 -1030
rect 198 -1033 297 -1032
rect 380 -1033 388 -1032
rect 397 -1033 913 -1032
rect 919 -1033 927 -1032
rect 940 -1033 1872 -1032
rect 121 -1035 199 -1034
rect 205 -1035 472 -1034
rect 499 -1035 528 -1034
rect 618 -1035 1137 -1034
rect 1139 -1035 1809 -1034
rect 100 -1037 528 -1036
rect 646 -1037 850 -1036
rect 877 -1037 899 -1036
rect 905 -1037 1851 -1036
rect 44 -1039 101 -1038
rect 114 -1039 122 -1038
rect 219 -1039 927 -1038
rect 954 -1039 1007 -1038
rect 1010 -1039 1767 -1038
rect 1808 -1039 1830 -1038
rect 114 -1041 178 -1040
rect 205 -1041 955 -1040
rect 982 -1041 997 -1040
rect 1010 -1041 1053 -1040
rect 1059 -1041 1550 -1040
rect 1591 -1041 1830 -1040
rect 177 -1043 430 -1042
rect 450 -1043 507 -1042
rect 520 -1043 570 -1042
rect 688 -1043 941 -1042
rect 961 -1043 997 -1042
rect 1013 -1043 1193 -1042
rect 1220 -1043 1235 -1042
rect 1297 -1043 1305 -1042
rect 1360 -1043 1872 -1042
rect 233 -1045 451 -1044
rect 520 -1045 923 -1044
rect 985 -1045 1655 -1044
rect 254 -1047 304 -1046
rect 352 -1047 430 -1046
rect 688 -1047 1154 -1046
rect 1206 -1047 1221 -1046
rect 1262 -1047 1655 -1046
rect 254 -1049 325 -1048
rect 352 -1049 650 -1048
rect 695 -1049 1154 -1048
rect 1199 -1049 1207 -1048
rect 1213 -1049 1263 -1048
rect 1304 -1049 1312 -1048
rect 1353 -1049 1361 -1048
rect 1472 -1049 1480 -1048
rect 1549 -1049 1788 -1048
rect 366 -1051 381 -1050
rect 401 -1051 423 -1050
rect 607 -1051 696 -1050
rect 723 -1051 1200 -1050
rect 1213 -1051 1284 -1050
rect 1479 -1051 1557 -1050
rect 1591 -1051 1690 -1050
rect 1787 -1051 1816 -1050
rect 275 -1053 423 -1052
rect 653 -1053 724 -1052
rect 751 -1053 857 -1052
rect 877 -1053 885 -1052
rect 1003 -1053 1354 -1052
rect 1465 -1053 1557 -1052
rect 1563 -1053 1690 -1052
rect 1815 -1053 1844 -1052
rect 16 -1055 885 -1054
rect 1003 -1055 1046 -1054
rect 1048 -1055 1802 -1054
rect 16 -1057 216 -1056
rect 275 -1057 318 -1056
rect 324 -1057 1046 -1056
rect 1052 -1057 1074 -1056
rect 1122 -1057 1130 -1056
rect 1150 -1057 1683 -1056
rect 1696 -1057 1844 -1056
rect 317 -1059 745 -1058
rect 782 -1059 1284 -1058
rect 1563 -1059 1627 -1058
rect 1682 -1059 1739 -1058
rect 1759 -1059 1802 -1058
rect 338 -1061 1130 -1060
rect 1150 -1061 1466 -1060
rect 1626 -1061 1648 -1060
rect 1696 -1061 1753 -1060
rect 331 -1063 339 -1062
rect 366 -1063 633 -1062
rect 744 -1063 801 -1062
rect 807 -1063 857 -1062
rect 1017 -1063 1739 -1062
rect 135 -1065 332 -1064
rect 765 -1065 808 -1064
rect 835 -1065 906 -1064
rect 1031 -1065 1760 -1064
rect 135 -1067 416 -1066
rect 597 -1067 766 -1066
rect 793 -1067 962 -1066
rect 1038 -1067 1102 -1066
rect 1227 -1067 1312 -1066
rect 1612 -1067 1648 -1066
rect 359 -1069 598 -1068
rect 628 -1069 836 -1068
rect 842 -1069 1116 -1068
rect 1227 -1069 1837 -1068
rect 359 -1071 374 -1070
rect 415 -1071 465 -1070
rect 639 -1071 794 -1070
rect 800 -1071 1035 -1070
rect 1041 -1071 1641 -1070
rect 1836 -1071 1858 -1070
rect 247 -1073 465 -1072
rect 639 -1073 755 -1072
rect 828 -1073 1102 -1072
rect 1115 -1073 1165 -1072
rect 1521 -1073 1613 -1072
rect 1640 -1073 1662 -1072
rect 1822 -1073 1858 -1072
rect 184 -1075 248 -1074
rect 289 -1075 374 -1074
rect 653 -1075 1522 -1074
rect 1661 -1075 1704 -1074
rect 163 -1077 185 -1076
rect 212 -1077 290 -1076
rect 684 -1077 1823 -1076
rect 23 -1079 213 -1078
rect 849 -1079 1382 -1078
rect 1675 -1079 1704 -1078
rect 23 -1081 311 -1080
rect 947 -1081 1032 -1080
rect 1059 -1081 1095 -1080
rect 1143 -1081 1165 -1080
rect 1381 -1081 1389 -1080
rect 1675 -1081 1732 -1080
rect 163 -1083 591 -1082
rect 947 -1083 976 -1082
rect 1024 -1083 1039 -1082
rect 1066 -1083 1095 -1082
rect 1143 -1083 1186 -1082
rect 1388 -1083 1396 -1082
rect 1577 -1083 1732 -1082
rect 555 -1085 591 -1084
rect 863 -1085 1067 -1084
rect 1073 -1085 1088 -1084
rect 1185 -1085 1231 -1084
rect 1339 -1085 1396 -1084
rect 1542 -1085 1578 -1084
rect 555 -1087 577 -1086
rect 740 -1087 1088 -1086
rect 1332 -1087 1340 -1086
rect 1542 -1087 1606 -1086
rect 576 -1089 1249 -1088
rect 1325 -1089 1333 -1088
rect 1605 -1089 1718 -1088
rect 740 -1091 1620 -1090
rect 1717 -1091 1781 -1090
rect 65 -1093 1620 -1092
rect 1780 -1093 1795 -1092
rect 2 -1095 66 -1094
rect 828 -1095 1231 -1094
rect 1248 -1095 1403 -1094
rect 1668 -1095 1795 -1094
rect 110 -1097 1669 -1096
rect 933 -1099 976 -1098
rect 1024 -1099 1172 -1098
rect 1318 -1099 1326 -1098
rect 1402 -1099 1487 -1098
rect 572 -1101 934 -1100
rect 1080 -1101 1753 -1100
rect 789 -1103 1319 -1102
rect 1486 -1103 1882 -1102
rect 814 -1105 1172 -1104
rect 814 -1107 944 -1106
rect 1080 -1107 1903 -1106
rect 2 -1118 73 -1117
rect 128 -1118 675 -1117
rect 716 -1118 930 -1117
rect 933 -1118 1151 -1117
rect 1153 -1118 1830 -1117
rect 1843 -1118 1868 -1117
rect 1878 -1118 1921 -1117
rect 1948 -1118 1956 -1117
rect 1976 -1118 1991 -1117
rect 16 -1120 223 -1119
rect 233 -1120 654 -1119
rect 656 -1120 773 -1119
rect 775 -1120 871 -1119
rect 880 -1120 1368 -1119
rect 1549 -1120 1893 -1119
rect 1969 -1120 1977 -1119
rect 16 -1122 115 -1121
rect 135 -1122 773 -1121
rect 779 -1122 857 -1121
rect 866 -1122 1025 -1121
rect 1045 -1122 1200 -1121
rect 1318 -1122 1907 -1121
rect 1962 -1122 1970 -1121
rect 23 -1124 566 -1123
rect 572 -1124 661 -1123
rect 674 -1124 703 -1123
rect 716 -1124 1081 -1123
rect 1132 -1124 1571 -1123
rect 1584 -1124 1886 -1123
rect 30 -1126 41 -1125
rect 44 -1126 934 -1125
rect 957 -1126 1704 -1125
rect 1759 -1126 1879 -1125
rect 30 -1128 199 -1127
rect 219 -1128 535 -1127
rect 562 -1128 843 -1127
rect 870 -1128 1291 -1127
rect 1311 -1128 1319 -1127
rect 1367 -1128 1389 -1127
rect 1451 -1128 1571 -1127
rect 1591 -1128 1760 -1127
rect 1780 -1128 1900 -1127
rect 61 -1130 269 -1129
rect 282 -1130 755 -1129
rect 758 -1130 1004 -1129
rect 1010 -1130 1025 -1129
rect 1045 -1130 1732 -1129
rect 1780 -1130 1788 -1129
rect 1808 -1130 1830 -1129
rect 1836 -1130 1844 -1129
rect 1871 -1130 1963 -1129
rect 65 -1132 528 -1131
rect 562 -1132 1231 -1131
rect 1360 -1132 1389 -1131
rect 1500 -1132 1550 -1131
rect 1591 -1132 1599 -1131
rect 1689 -1132 1732 -1131
rect 1787 -1132 1802 -1131
rect 1822 -1132 1865 -1131
rect 65 -1134 416 -1133
rect 422 -1134 454 -1133
rect 464 -1134 682 -1133
rect 695 -1134 703 -1133
rect 730 -1134 748 -1133
rect 751 -1134 1452 -1133
rect 1458 -1134 1501 -1133
rect 1542 -1134 1872 -1133
rect 72 -1136 395 -1135
rect 415 -1136 587 -1135
rect 625 -1136 654 -1135
rect 660 -1136 976 -1135
rect 996 -1136 1011 -1135
rect 1017 -1136 1578 -1135
rect 1598 -1136 1613 -1135
rect 1682 -1136 1823 -1135
rect 100 -1138 129 -1137
rect 131 -1138 682 -1137
rect 695 -1138 724 -1137
rect 730 -1138 766 -1137
rect 782 -1138 1263 -1137
rect 1423 -1138 1683 -1137
rect 1696 -1138 1837 -1137
rect 9 -1140 101 -1139
rect 114 -1140 790 -1139
rect 810 -1140 1032 -1139
rect 1080 -1140 1102 -1139
rect 1139 -1140 1193 -1139
rect 1402 -1140 1424 -1139
rect 1458 -1140 1487 -1139
rect 1493 -1140 1543 -1139
rect 1563 -1140 1578 -1139
rect 1605 -1140 1690 -1139
rect 1724 -1140 1865 -1139
rect 9 -1142 426 -1141
rect 429 -1142 857 -1141
rect 859 -1142 1263 -1141
rect 1381 -1142 1403 -1141
rect 1444 -1142 1494 -1141
rect 1521 -1142 1697 -1141
rect 1794 -1142 1809 -1141
rect 79 -1144 1564 -1143
rect 1605 -1144 1627 -1143
rect 1668 -1144 1725 -1143
rect 1752 -1144 1795 -1143
rect 121 -1146 136 -1145
rect 159 -1146 311 -1145
rect 331 -1146 535 -1145
rect 555 -1146 626 -1145
rect 723 -1146 745 -1145
rect 761 -1146 1291 -1145
rect 1444 -1146 1480 -1145
rect 1486 -1146 1557 -1145
rect 1612 -1146 1634 -1145
rect 1668 -1146 1816 -1145
rect 121 -1148 783 -1147
rect 814 -1148 843 -1147
rect 863 -1148 1382 -1147
rect 1437 -1148 1480 -1147
rect 1507 -1148 1557 -1147
rect 1626 -1148 1641 -1147
rect 1745 -1148 1753 -1147
rect 180 -1150 853 -1149
rect 863 -1150 878 -1149
rect 894 -1150 1648 -1149
rect 1717 -1150 1746 -1149
rect 198 -1152 318 -1151
rect 359 -1152 629 -1151
rect 670 -1152 1508 -1151
rect 1514 -1152 1641 -1151
rect 1647 -1152 1676 -1151
rect 1717 -1152 1739 -1151
rect 82 -1154 318 -1153
rect 359 -1154 381 -1153
rect 422 -1154 1130 -1153
rect 1136 -1154 1676 -1153
rect 1710 -1154 1739 -1153
rect 233 -1156 248 -1155
rect 261 -1156 293 -1155
rect 303 -1156 332 -1155
rect 366 -1156 370 -1155
rect 373 -1156 395 -1155
rect 436 -1156 524 -1155
rect 555 -1156 668 -1155
rect 684 -1156 1816 -1155
rect 51 -1158 374 -1157
rect 380 -1158 801 -1157
rect 873 -1158 1585 -1157
rect 1633 -1158 1662 -1157
rect 51 -1160 741 -1159
rect 779 -1160 1438 -1159
rect 1465 -1160 1515 -1159
rect 1521 -1160 1655 -1159
rect 240 -1162 248 -1161
rect 268 -1162 276 -1161
rect 282 -1162 346 -1161
rect 366 -1162 388 -1161
rect 436 -1162 913 -1161
rect 926 -1162 1361 -1161
rect 1472 -1162 1655 -1161
rect 163 -1164 346 -1163
rect 352 -1164 927 -1163
rect 975 -1164 983 -1163
rect 989 -1164 997 -1163
rect 1003 -1164 1221 -1163
rect 1248 -1164 1473 -1163
rect 1535 -1164 1662 -1163
rect 58 -1166 353 -1165
rect 446 -1166 1704 -1165
rect 163 -1168 458 -1167
rect 464 -1168 542 -1167
rect 583 -1168 787 -1167
rect 912 -1168 1130 -1167
rect 1160 -1168 1914 -1167
rect 142 -1170 542 -1169
rect 583 -1170 1032 -1169
rect 1038 -1170 1221 -1169
rect 1241 -1170 1249 -1169
rect 142 -1172 230 -1171
rect 240 -1172 297 -1171
rect 303 -1172 909 -1171
rect 961 -1172 990 -1171
rect 1017 -1172 1466 -1171
rect 254 -1174 297 -1173
rect 313 -1174 1137 -1173
rect 1164 -1174 1193 -1173
rect 1234 -1174 1242 -1173
rect 212 -1176 255 -1175
rect 275 -1176 339 -1175
rect 450 -1176 1802 -1175
rect 37 -1178 451 -1177
rect 453 -1178 1200 -1177
rect 1213 -1178 1235 -1177
rect 289 -1180 577 -1179
rect 590 -1180 815 -1179
rect 849 -1180 1039 -1179
rect 1048 -1180 1711 -1179
rect 107 -1182 1049 -1181
rect 1087 -1182 1312 -1181
rect 107 -1184 892 -1183
rect 982 -1184 1053 -1183
rect 1059 -1184 1088 -1183
rect 1094 -1184 1102 -1183
rect 1115 -1184 1165 -1183
rect 156 -1186 591 -1185
rect 632 -1186 1536 -1185
rect 324 -1188 633 -1187
rect 667 -1188 1529 -1187
rect 324 -1190 486 -1189
rect 516 -1190 1228 -1189
rect 338 -1192 605 -1191
rect 709 -1192 801 -1191
rect 821 -1192 850 -1191
rect 877 -1192 1060 -1191
rect 1108 -1192 1116 -1191
rect 1157 -1192 1214 -1191
rect 37 -1194 605 -1193
rect 709 -1194 808 -1193
rect 891 -1194 899 -1193
rect 1052 -1194 1067 -1193
rect 1108 -1194 1284 -1193
rect 408 -1196 1284 -1195
rect 408 -1198 689 -1197
rect 733 -1198 1851 -1197
rect 443 -1200 1095 -1199
rect 1157 -1200 1410 -1199
rect 212 -1202 444 -1201
rect 457 -1202 507 -1201
rect 576 -1202 619 -1201
rect 737 -1202 1179 -1201
rect 1181 -1202 1851 -1201
rect 44 -1204 1179 -1203
rect 1185 -1204 1529 -1203
rect 289 -1206 619 -1205
rect 744 -1206 822 -1205
rect 898 -1206 906 -1205
rect 1066 -1206 1074 -1205
rect 1143 -1206 1186 -1205
rect 1395 -1206 1410 -1205
rect 471 -1208 528 -1207
rect 611 -1208 689 -1207
rect 747 -1208 766 -1207
rect 807 -1208 955 -1207
rect 1143 -1208 1256 -1207
rect 1374 -1208 1396 -1207
rect 429 -1210 472 -1209
rect 474 -1210 500 -1209
rect 506 -1210 640 -1209
rect 905 -1210 1858 -1209
rect 124 -1212 500 -1211
rect 513 -1212 738 -1211
rect 940 -1212 1074 -1211
rect 1255 -1212 1340 -1211
rect 1353 -1212 1375 -1211
rect 1619 -1212 1858 -1211
rect 82 -1214 1620 -1213
rect 478 -1216 752 -1215
rect 940 -1216 965 -1215
rect 1325 -1216 1340 -1215
rect 1346 -1216 1354 -1215
rect 177 -1218 479 -1217
rect 485 -1218 549 -1217
rect 579 -1218 612 -1217
rect 947 -1218 955 -1217
rect 1297 -1218 1326 -1217
rect 1332 -1218 1347 -1217
rect 177 -1220 1172 -1219
rect 1297 -1220 1305 -1219
rect 520 -1222 1172 -1221
rect 1304 -1222 1431 -1221
rect 93 -1224 521 -1223
rect 548 -1224 969 -1223
rect 1416 -1224 1431 -1223
rect 47 -1226 1417 -1225
rect 93 -1228 150 -1227
rect 569 -1228 1333 -1227
rect 149 -1230 206 -1229
rect 492 -1230 570 -1229
rect 597 -1230 640 -1229
rect 828 -1230 969 -1229
rect 58 -1232 598 -1231
rect 828 -1232 885 -1231
rect 919 -1232 948 -1231
rect 191 -1234 206 -1233
rect 492 -1234 1021 -1233
rect 170 -1236 192 -1235
rect 646 -1236 920 -1235
rect 170 -1238 647 -1237
rect 835 -1238 885 -1237
rect 793 -1240 836 -1239
rect 226 -1242 794 -1241
rect 23 -1253 94 -1252
rect 107 -1253 146 -1252
rect 163 -1253 227 -1252
rect 247 -1253 262 -1252
rect 282 -1253 454 -1252
rect 457 -1253 671 -1252
rect 688 -1253 780 -1252
rect 793 -1253 1077 -1252
rect 1111 -1253 1879 -1252
rect 1906 -1253 1949 -1252
rect 1962 -1253 1998 -1252
rect 30 -1255 447 -1254
rect 457 -1255 598 -1254
rect 628 -1255 787 -1254
rect 821 -1255 1067 -1254
rect 1129 -1255 1823 -1254
rect 1843 -1255 1907 -1254
rect 1913 -1255 1942 -1254
rect 1976 -1255 1984 -1254
rect 30 -1257 209 -1256
rect 226 -1257 514 -1256
rect 541 -1257 598 -1256
rect 604 -1257 822 -1256
rect 838 -1257 1473 -1256
rect 1675 -1257 1844 -1256
rect 1920 -1257 1935 -1256
rect 1955 -1257 1977 -1256
rect 37 -1259 45 -1258
rect 58 -1259 794 -1258
rect 856 -1259 1760 -1258
rect 40 -1261 1655 -1260
rect 1759 -1261 1914 -1260
rect 44 -1263 577 -1262
rect 586 -1263 850 -1262
rect 856 -1263 874 -1262
rect 908 -1263 1221 -1262
rect 1269 -1263 1273 -1262
rect 1290 -1263 1921 -1262
rect 58 -1265 1858 -1264
rect 61 -1267 1522 -1266
rect 1612 -1267 1655 -1266
rect 1787 -1267 1858 -1266
rect 65 -1269 283 -1268
rect 289 -1269 402 -1268
rect 415 -1269 514 -1268
rect 562 -1269 1074 -1268
rect 1129 -1269 1137 -1268
rect 1178 -1269 1886 -1268
rect 51 -1271 66 -1270
rect 79 -1271 339 -1270
rect 352 -1271 657 -1270
rect 688 -1271 724 -1270
rect 775 -1271 1851 -1270
rect 9 -1273 80 -1272
rect 82 -1273 605 -1272
rect 646 -1273 1133 -1272
rect 1171 -1273 1179 -1272
rect 1220 -1273 1235 -1272
rect 1269 -1273 1277 -1272
rect 1290 -1273 1298 -1272
rect 1388 -1273 1392 -1272
rect 1458 -1273 1473 -1272
rect 1542 -1273 1613 -1272
rect 1626 -1273 1676 -1272
rect 1787 -1273 1917 -1272
rect 9 -1275 801 -1274
rect 824 -1275 850 -1274
rect 870 -1275 913 -1274
rect 922 -1275 1893 -1274
rect 2 -1277 801 -1276
rect 912 -1277 1109 -1276
rect 1122 -1277 1137 -1276
rect 1171 -1277 1522 -1276
rect 1808 -1277 1851 -1276
rect 86 -1279 171 -1278
rect 177 -1279 612 -1278
rect 681 -1279 724 -1278
rect 779 -1279 1070 -1278
rect 1073 -1279 1662 -1278
rect 1829 -1279 1886 -1278
rect 54 -1281 87 -1280
rect 93 -1281 143 -1280
rect 149 -1281 178 -1280
rect 247 -1281 1095 -1280
rect 1234 -1281 1263 -1280
rect 1297 -1281 1333 -1280
rect 1388 -1281 1410 -1280
rect 1437 -1281 1459 -1280
rect 1486 -1281 1627 -1280
rect 1773 -1281 1830 -1280
rect 107 -1283 549 -1282
rect 611 -1283 619 -1282
rect 653 -1283 682 -1282
rect 877 -1283 1123 -1282
rect 1143 -1283 1263 -1282
rect 1416 -1283 1438 -1282
rect 1479 -1283 1487 -1282
rect 1493 -1283 1543 -1282
rect 1591 -1283 1662 -1282
rect 1745 -1283 1774 -1282
rect 110 -1285 1823 -1284
rect 121 -1287 230 -1286
rect 254 -1287 580 -1286
rect 618 -1287 892 -1286
rect 926 -1287 1879 -1286
rect 152 -1289 262 -1288
rect 296 -1289 300 -1288
rect 317 -1289 542 -1288
rect 548 -1289 941 -1288
rect 964 -1289 1683 -1288
rect 156 -1291 1893 -1290
rect 156 -1293 661 -1292
rect 712 -1293 1683 -1292
rect 128 -1295 661 -1294
rect 877 -1295 1025 -1294
rect 1038 -1295 1158 -1294
rect 1244 -1295 1494 -1294
rect 1563 -1295 1592 -1294
rect 1605 -1295 1746 -1294
rect 75 -1297 1025 -1296
rect 1045 -1297 1088 -1296
rect 1094 -1297 1116 -1296
rect 1143 -1297 1186 -1296
rect 1255 -1297 1333 -1296
rect 1416 -1297 1424 -1296
rect 1465 -1297 1480 -1296
rect 124 -1299 1088 -1298
rect 1185 -1299 1837 -1298
rect 128 -1301 843 -1300
rect 891 -1301 948 -1300
rect 961 -1301 1039 -1300
rect 1055 -1301 1809 -1300
rect 163 -1303 241 -1302
rect 254 -1303 671 -1302
rect 842 -1303 899 -1302
rect 929 -1303 1606 -1302
rect 1780 -1303 1837 -1302
rect 170 -1305 381 -1304
rect 394 -1305 426 -1304
rect 443 -1305 1312 -1304
rect 1423 -1305 1508 -1304
rect 1766 -1305 1781 -1304
rect 205 -1307 241 -1306
rect 268 -1307 395 -1306
rect 401 -1307 556 -1306
rect 807 -1307 899 -1306
rect 929 -1307 1564 -1306
rect 1752 -1307 1767 -1306
rect 184 -1309 206 -1308
rect 233 -1309 269 -1308
rect 296 -1309 332 -1308
rect 338 -1309 409 -1308
rect 422 -1309 1802 -1308
rect 184 -1311 304 -1310
rect 310 -1311 556 -1310
rect 807 -1311 1081 -1310
rect 1108 -1311 1508 -1310
rect 1696 -1311 1753 -1310
rect 100 -1313 311 -1312
rect 317 -1313 388 -1312
rect 408 -1313 521 -1312
rect 534 -1313 563 -1312
rect 810 -1313 1802 -1312
rect 72 -1315 388 -1314
rect 422 -1315 668 -1314
rect 947 -1315 955 -1314
rect 961 -1315 990 -1314
rect 1017 -1315 1872 -1314
rect 51 -1317 668 -1316
rect 954 -1317 976 -1316
rect 989 -1317 1032 -1316
rect 1066 -1317 1312 -1316
rect 1391 -1317 1410 -1316
rect 1451 -1317 1466 -1316
rect 1668 -1317 1872 -1316
rect 72 -1319 570 -1318
rect 968 -1319 1116 -1318
rect 1255 -1319 1375 -1318
rect 1598 -1319 1669 -1318
rect 1696 -1319 1704 -1318
rect 100 -1321 265 -1320
rect 352 -1321 360 -1320
rect 366 -1321 381 -1320
rect 443 -1321 773 -1320
rect 968 -1321 1021 -1320
rect 1031 -1321 1326 -1320
rect 1360 -1321 1452 -1320
rect 142 -1323 304 -1322
rect 324 -1323 360 -1322
rect 366 -1323 517 -1322
rect 534 -1323 766 -1322
rect 772 -1323 815 -1322
rect 975 -1323 983 -1322
rect 996 -1323 1018 -1322
rect 1080 -1323 1165 -1322
rect 1304 -1323 1361 -1322
rect 1374 -1323 1396 -1322
rect 1444 -1323 1599 -1322
rect 233 -1325 493 -1324
rect 530 -1325 1445 -1324
rect 275 -1327 325 -1326
rect 373 -1327 416 -1326
rect 450 -1327 815 -1326
rect 859 -1327 1305 -1326
rect 1325 -1327 1340 -1326
rect 212 -1329 276 -1328
rect 373 -1329 678 -1328
rect 765 -1329 836 -1328
rect 859 -1329 1704 -1328
rect 198 -1331 213 -1330
rect 436 -1331 451 -1330
rect 464 -1331 647 -1330
rect 905 -1331 983 -1330
rect 996 -1331 1900 -1330
rect 198 -1333 640 -1332
rect 884 -1333 906 -1332
rect 1164 -1333 1214 -1332
rect 1227 -1333 1396 -1332
rect 1864 -1333 1900 -1332
rect 436 -1335 759 -1334
rect 884 -1335 920 -1334
rect 1059 -1335 1214 -1334
rect 1227 -1335 1249 -1334
rect 1318 -1335 1340 -1334
rect 1815 -1335 1865 -1334
rect 464 -1337 717 -1336
rect 751 -1337 759 -1336
rect 1052 -1337 1060 -1336
rect 1248 -1337 1347 -1336
rect 1794 -1337 1816 -1336
rect 471 -1339 1004 -1338
rect 1318 -1339 1403 -1338
rect 1647 -1339 1795 -1338
rect 474 -1341 626 -1340
rect 639 -1341 675 -1340
rect 716 -1341 738 -1340
rect 744 -1341 752 -1340
rect 1003 -1341 1182 -1340
rect 1346 -1341 1354 -1340
rect 1647 -1341 1739 -1340
rect 114 -1343 675 -1342
rect 737 -1343 1011 -1342
rect 1052 -1343 1403 -1342
rect 1717 -1343 1739 -1342
rect 114 -1345 346 -1344
rect 478 -1345 521 -1344
rect 569 -1345 710 -1344
rect 943 -1345 1718 -1344
rect 159 -1347 346 -1346
rect 478 -1347 500 -1346
rect 590 -1347 836 -1346
rect 1353 -1347 1368 -1346
rect 173 -1349 1011 -1348
rect 1367 -1349 1382 -1348
rect 485 -1351 584 -1350
rect 625 -1351 696 -1350
rect 709 -1351 787 -1350
rect 1241 -1351 1382 -1350
rect 219 -1353 696 -1352
rect 1241 -1353 1641 -1352
rect 191 -1355 220 -1354
rect 432 -1355 584 -1354
rect 1556 -1355 1641 -1354
rect 191 -1357 566 -1356
rect 1535 -1357 1557 -1356
rect 485 -1359 703 -1358
rect 1528 -1359 1536 -1358
rect 429 -1361 703 -1360
rect 1514 -1361 1529 -1360
rect 429 -1363 1620 -1362
rect 492 -1365 507 -1364
rect 527 -1365 591 -1364
rect 1500 -1365 1515 -1364
rect 1570 -1365 1620 -1364
rect 499 -1367 934 -1366
rect 1500 -1367 1634 -1366
rect 506 -1369 633 -1368
rect 933 -1369 1000 -1368
rect 1549 -1369 1571 -1368
rect 1577 -1369 1634 -1368
rect 527 -1371 1284 -1370
rect 1549 -1371 1732 -1370
rect 632 -1373 829 -1372
rect 919 -1373 1578 -1372
rect 1724 -1373 1732 -1372
rect 744 -1375 1284 -1374
rect 1710 -1375 1725 -1374
rect 828 -1377 864 -1376
rect 1584 -1377 1711 -1376
rect 653 -1379 864 -1378
rect 1199 -1379 1585 -1378
rect 1192 -1381 1200 -1380
rect 1192 -1383 1207 -1382
rect 180 -1385 1207 -1384
rect 2 -1396 209 -1395
rect 485 -1396 920 -1395
rect 940 -1396 1648 -1395
rect 1899 -1396 1963 -1395
rect 1976 -1396 2026 -1395
rect 9 -1398 216 -1397
rect 485 -1398 493 -1397
rect 527 -1398 647 -1397
rect 674 -1398 682 -1397
rect 712 -1398 913 -1397
rect 947 -1398 1000 -1397
rect 1003 -1398 1014 -1397
rect 1038 -1398 1074 -1397
rect 1104 -1398 1543 -1397
rect 1647 -1398 1823 -1397
rect 1913 -1398 1928 -1397
rect 1941 -1398 2012 -1397
rect 9 -1400 262 -1399
rect 527 -1400 923 -1399
rect 926 -1400 1039 -1399
rect 1052 -1400 1809 -1399
rect 1822 -1400 1921 -1399
rect 1948 -1400 1956 -1399
rect 1983 -1400 1987 -1399
rect 1997 -1400 2019 -1399
rect 16 -1402 153 -1401
rect 184 -1402 1186 -1401
rect 1241 -1402 1795 -1401
rect 1843 -1402 1949 -1401
rect 1983 -1402 1991 -1401
rect 16 -1404 122 -1403
rect 142 -1404 1683 -1403
rect 1780 -1404 1844 -1403
rect 1864 -1404 1928 -1403
rect 30 -1406 958 -1405
rect 968 -1406 1445 -1405
rect 1577 -1406 1809 -1405
rect 1864 -1406 1879 -1405
rect 1916 -1406 1935 -1405
rect 30 -1408 619 -1407
rect 632 -1408 668 -1407
rect 677 -1408 962 -1407
rect 975 -1408 1053 -1407
rect 1055 -1408 1382 -1407
rect 1444 -1408 1592 -1407
rect 1605 -1408 1683 -1407
rect 1738 -1408 1781 -1407
rect 1787 -1408 1879 -1407
rect 1885 -1408 1935 -1407
rect 47 -1410 1543 -1409
rect 1556 -1410 1606 -1409
rect 1661 -1410 1739 -1409
rect 1794 -1410 1858 -1409
rect 51 -1412 1900 -1411
rect 51 -1414 101 -1413
rect 107 -1414 234 -1413
rect 450 -1414 633 -1413
rect 814 -1414 969 -1413
rect 975 -1414 1308 -1413
rect 1335 -1414 1907 -1413
rect 58 -1416 500 -1415
rect 548 -1416 682 -1415
rect 814 -1416 829 -1415
rect 849 -1416 941 -1415
rect 947 -1416 1361 -1415
rect 1437 -1416 1592 -1415
rect 1801 -1416 1907 -1415
rect 58 -1418 248 -1417
rect 408 -1418 549 -1417
rect 562 -1418 710 -1417
rect 744 -1418 829 -1417
rect 905 -1418 913 -1417
rect 922 -1418 1942 -1417
rect 65 -1420 73 -1419
rect 79 -1420 262 -1419
rect 408 -1420 507 -1419
rect 562 -1420 710 -1419
rect 744 -1420 836 -1419
rect 842 -1420 906 -1419
rect 926 -1420 934 -1419
rect 961 -1420 1179 -1419
rect 1185 -1420 1263 -1419
rect 1283 -1420 1837 -1419
rect 1850 -1420 1858 -1419
rect 79 -1422 836 -1421
rect 884 -1422 934 -1421
rect 985 -1422 1410 -1421
rect 1521 -1422 1557 -1421
rect 1577 -1422 1655 -1421
rect 1703 -1422 1802 -1421
rect 82 -1424 1137 -1423
rect 1164 -1424 1242 -1423
rect 1283 -1424 1326 -1423
rect 1346 -1424 1361 -1423
rect 1374 -1424 1410 -1423
rect 1507 -1424 1522 -1423
rect 1535 -1424 1662 -1423
rect 1703 -1424 1774 -1423
rect 86 -1426 185 -1425
rect 194 -1426 696 -1425
rect 751 -1426 843 -1425
rect 982 -1426 1137 -1425
rect 1150 -1426 1165 -1425
rect 1171 -1426 1452 -1425
rect 1479 -1426 1508 -1425
rect 1549 -1426 1851 -1425
rect 93 -1428 101 -1427
rect 114 -1428 433 -1427
rect 450 -1428 580 -1427
rect 583 -1428 696 -1427
rect 786 -1428 850 -1427
rect 982 -1428 1641 -1427
rect 1717 -1428 1774 -1427
rect 93 -1430 150 -1429
rect 198 -1430 244 -1429
rect 247 -1430 951 -1429
rect 996 -1430 1382 -1429
rect 1388 -1430 1452 -1429
rect 1549 -1430 1627 -1429
rect 1640 -1430 1998 -1429
rect 114 -1432 437 -1431
rect 492 -1432 668 -1431
rect 807 -1432 1172 -1431
rect 1178 -1432 1396 -1431
rect 1759 -1432 1837 -1431
rect 121 -1434 132 -1433
rect 145 -1434 1914 -1433
rect 145 -1436 1207 -1435
rect 1248 -1436 1326 -1435
rect 1346 -1436 1473 -1435
rect 1752 -1436 1760 -1435
rect 149 -1438 1109 -1437
rect 1111 -1438 1613 -1437
rect 198 -1440 283 -1439
rect 310 -1440 787 -1439
rect 793 -1440 808 -1439
rect 929 -1440 1473 -1439
rect 1493 -1440 1753 -1439
rect 37 -1442 283 -1441
rect 303 -1442 311 -1441
rect 373 -1442 437 -1441
rect 506 -1442 514 -1441
rect 569 -1442 944 -1441
rect 954 -1442 997 -1441
rect 1003 -1442 1046 -1441
rect 1066 -1442 1711 -1441
rect 37 -1444 76 -1443
rect 86 -1444 955 -1443
rect 1006 -1444 1200 -1443
rect 1248 -1444 1291 -1443
rect 1367 -1444 1396 -1443
rect 1493 -1444 1571 -1443
rect 1633 -1444 1711 -1443
rect 1986 -1444 1991 -1443
rect 110 -1446 304 -1445
rect 338 -1446 374 -1445
rect 387 -1446 1207 -1445
rect 1255 -1446 1389 -1445
rect 1528 -1446 1571 -1445
rect 128 -1448 1634 -1447
rect 128 -1450 136 -1449
rect 205 -1450 227 -1449
rect 233 -1450 1305 -1449
rect 1367 -1450 1424 -1449
rect 1486 -1450 1529 -1449
rect 1563 -1450 1613 -1449
rect 135 -1452 178 -1451
rect 226 -1452 332 -1451
rect 338 -1452 521 -1451
rect 555 -1452 570 -1451
rect 576 -1452 860 -1451
rect 1010 -1452 1718 -1451
rect 296 -1454 332 -1453
rect 387 -1454 395 -1453
rect 422 -1454 584 -1453
rect 590 -1454 647 -1453
rect 663 -1454 1438 -1453
rect 163 -1456 395 -1455
rect 415 -1456 423 -1455
rect 513 -1456 612 -1455
rect 618 -1456 629 -1455
rect 793 -1456 801 -1455
rect 898 -1456 1011 -1455
rect 1024 -1456 1886 -1455
rect 163 -1458 255 -1457
rect 415 -1458 458 -1457
rect 478 -1458 801 -1457
rect 821 -1458 899 -1457
rect 1031 -1458 1627 -1457
rect 212 -1460 458 -1459
rect 520 -1460 689 -1459
rect 702 -1460 822 -1459
rect 989 -1460 1032 -1459
rect 1034 -1460 1655 -1459
rect 177 -1462 213 -1461
rect 219 -1462 297 -1461
rect 443 -1462 479 -1461
rect 534 -1462 703 -1461
rect 751 -1462 1025 -1461
rect 1087 -1462 1536 -1461
rect 191 -1464 535 -1463
rect 555 -1464 2008 -1463
rect 191 -1466 773 -1465
rect 989 -1466 1018 -1465
rect 1087 -1466 1095 -1465
rect 1108 -1466 1480 -1465
rect 219 -1468 290 -1467
rect 359 -1468 444 -1467
rect 576 -1468 780 -1467
rect 863 -1468 1018 -1467
rect 1080 -1468 1095 -1467
rect 1111 -1468 1291 -1467
rect 1304 -1468 1830 -1467
rect 254 -1470 269 -1469
rect 275 -1470 290 -1469
rect 324 -1470 360 -1469
rect 590 -1470 857 -1469
rect 1080 -1470 1266 -1469
rect 1286 -1470 1340 -1469
rect 1402 -1470 1424 -1469
rect 1731 -1470 1830 -1469
rect 240 -1472 269 -1471
rect 275 -1472 353 -1471
rect 597 -1472 657 -1471
rect 670 -1472 1403 -1471
rect 1724 -1472 1732 -1471
rect 324 -1474 402 -1473
rect 464 -1474 598 -1473
rect 604 -1474 885 -1473
rect 1115 -1474 1263 -1473
rect 1339 -1474 1459 -1473
rect 1696 -1474 1725 -1473
rect 352 -1476 640 -1475
rect 653 -1476 864 -1475
rect 1118 -1476 1746 -1475
rect 401 -1478 503 -1477
rect 541 -1478 640 -1477
rect 653 -1478 1133 -1477
rect 1143 -1478 1151 -1477
rect 1160 -1478 1487 -1477
rect 1675 -1478 1746 -1477
rect 44 -1480 542 -1479
rect 604 -1480 713 -1479
rect 758 -1480 773 -1479
rect 779 -1480 892 -1479
rect 1059 -1480 1144 -1479
rect 1199 -1480 1214 -1479
rect 1220 -1480 1256 -1479
rect 1416 -1480 1459 -1479
rect 1584 -1480 1676 -1479
rect 44 -1482 1921 -1481
rect 170 -1484 759 -1483
rect 856 -1484 1116 -1483
rect 1122 -1484 1564 -1483
rect 61 -1486 171 -1485
rect 464 -1486 531 -1485
rect 611 -1486 1077 -1485
rect 1101 -1486 1123 -1485
rect 1157 -1486 1214 -1485
rect 1244 -1486 1697 -1485
rect 61 -1488 66 -1487
rect 628 -1488 717 -1487
rect 870 -1488 892 -1487
rect 1059 -1488 1130 -1487
rect 1157 -1488 1872 -1487
rect 471 -1490 871 -1489
rect 1101 -1490 1312 -1489
rect 1318 -1490 1417 -1489
rect 1815 -1490 1872 -1489
rect 366 -1492 472 -1491
rect 688 -1492 731 -1491
rect 1129 -1492 1375 -1491
rect 1668 -1492 1816 -1491
rect 366 -1494 381 -1493
rect 716 -1494 738 -1493
rect 1192 -1494 1221 -1493
rect 1297 -1494 1319 -1493
rect 1598 -1494 1669 -1493
rect 380 -1496 766 -1495
rect 1192 -1496 1788 -1495
rect 660 -1498 766 -1497
rect 1269 -1498 1298 -1497
rect 1311 -1498 1515 -1497
rect 1598 -1498 1690 -1497
rect 156 -1500 661 -1499
rect 723 -1500 738 -1499
rect 1269 -1500 1277 -1499
rect 1619 -1500 1690 -1499
rect 156 -1502 430 -1501
rect 730 -1502 755 -1501
rect 1069 -1502 1620 -1501
rect 240 -1504 724 -1503
rect 1069 -1504 1501 -1503
rect 317 -1506 430 -1505
rect 1234 -1506 1277 -1505
rect 1465 -1506 1501 -1505
rect 317 -1508 346 -1507
rect 1227 -1508 1235 -1507
rect 1430 -1508 1466 -1507
rect 166 -1510 346 -1509
rect 625 -1510 1228 -1509
rect 1353 -1510 1431 -1509
rect 625 -1512 1585 -1511
rect 1332 -1514 1354 -1513
rect 1332 -1516 1515 -1515
rect 2 -1527 48 -1526
rect 58 -1527 1725 -1526
rect 1808 -1527 1812 -1526
rect 1948 -1527 1970 -1526
rect 1979 -1527 1991 -1526
rect 2 -1529 178 -1528
rect 180 -1529 255 -1528
rect 338 -1529 752 -1528
rect 754 -1529 1662 -1528
rect 1689 -1529 1725 -1528
rect 1766 -1529 1949 -1528
rect 1955 -1529 1973 -1528
rect 1983 -1529 2001 -1528
rect 23 -1531 69 -1530
rect 82 -1531 1105 -1530
rect 1108 -1531 1830 -1530
rect 23 -1533 199 -1532
rect 233 -1533 325 -1532
rect 338 -1533 360 -1532
rect 485 -1533 661 -1532
rect 663 -1533 752 -1532
rect 768 -1533 815 -1532
rect 884 -1533 1161 -1532
rect 1192 -1533 1235 -1532
rect 1262 -1533 1347 -1532
rect 1356 -1533 1732 -1532
rect 1808 -1533 1879 -1532
rect 30 -1535 920 -1534
rect 954 -1535 1851 -1534
rect 30 -1537 248 -1536
rect 254 -1537 1056 -1536
rect 1101 -1537 1340 -1536
rect 1346 -1537 1361 -1536
rect 1503 -1537 1837 -1536
rect 37 -1539 500 -1538
rect 502 -1539 1039 -1538
rect 1108 -1539 1336 -1538
rect 1339 -1539 1354 -1538
rect 1360 -1539 1382 -1538
rect 1591 -1539 2005 -1538
rect 37 -1541 52 -1540
rect 58 -1541 108 -1540
rect 117 -1541 122 -1540
rect 142 -1541 304 -1540
rect 324 -1541 444 -1540
rect 499 -1541 556 -1540
rect 593 -1541 689 -1540
rect 709 -1541 878 -1540
rect 905 -1541 948 -1540
rect 957 -1541 1690 -1540
rect 1703 -1541 1767 -1540
rect 1811 -1541 1879 -1540
rect 9 -1543 52 -1542
rect 86 -1543 108 -1542
rect 121 -1543 185 -1542
rect 194 -1543 1207 -1542
rect 1234 -1543 1256 -1542
rect 1262 -1543 1287 -1542
rect 1353 -1543 1529 -1542
rect 1577 -1543 1704 -1542
rect 1717 -1543 1851 -1542
rect 9 -1545 157 -1544
rect 184 -1545 545 -1544
rect 555 -1545 703 -1544
rect 712 -1545 1543 -1544
rect 1577 -1545 1613 -1544
rect 1661 -1545 1977 -1544
rect 44 -1547 101 -1546
rect 142 -1547 629 -1546
rect 667 -1547 1172 -1546
rect 1199 -1547 1256 -1546
rect 1265 -1547 1963 -1546
rect 1976 -1547 2026 -1546
rect 16 -1549 45 -1548
rect 79 -1549 101 -1548
rect 114 -1549 668 -1548
rect 674 -1549 1039 -1548
rect 1111 -1549 1823 -1548
rect 1829 -1549 1886 -1548
rect 16 -1551 90 -1550
rect 145 -1551 199 -1550
rect 226 -1551 248 -1550
rect 289 -1551 486 -1550
rect 618 -1551 1102 -1550
rect 1118 -1551 1186 -1550
rect 1199 -1551 1214 -1550
rect 1374 -1551 1382 -1550
rect 1493 -1551 1592 -1550
rect 1612 -1551 1620 -1550
rect 1731 -1551 1753 -1550
rect 1794 -1551 1886 -1550
rect 86 -1553 699 -1552
rect 702 -1553 822 -1552
rect 835 -1553 878 -1552
rect 961 -1553 1333 -1552
rect 1374 -1553 1396 -1552
rect 1493 -1553 1669 -1552
rect 1822 -1553 1907 -1552
rect 128 -1555 146 -1554
rect 156 -1555 220 -1554
rect 226 -1555 1116 -1554
rect 1129 -1555 1882 -1554
rect 1906 -1555 1935 -1554
rect 93 -1557 129 -1556
rect 191 -1557 220 -1556
rect 233 -1557 311 -1556
rect 345 -1557 671 -1556
rect 681 -1557 1305 -1556
rect 1307 -1557 1753 -1556
rect 1871 -1557 1935 -1556
rect 65 -1559 94 -1558
rect 163 -1559 192 -1558
rect 205 -1559 346 -1558
rect 415 -1559 822 -1558
rect 849 -1559 906 -1558
rect 971 -1559 1284 -1558
rect 1307 -1559 1858 -1558
rect 1871 -1559 1921 -1558
rect 163 -1561 661 -1560
rect 663 -1561 1795 -1560
rect 205 -1563 521 -1562
rect 646 -1563 675 -1562
rect 681 -1563 829 -1562
rect 863 -1563 1718 -1562
rect 268 -1565 311 -1564
rect 397 -1565 647 -1564
rect 670 -1565 843 -1564
rect 1003 -1565 1802 -1564
rect 268 -1567 570 -1566
rect 583 -1567 843 -1566
rect 968 -1567 1004 -1566
rect 1073 -1567 1116 -1566
rect 1132 -1567 1312 -1566
rect 1332 -1567 1865 -1566
rect 282 -1569 521 -1568
rect 569 -1569 577 -1568
rect 583 -1569 731 -1568
rect 800 -1569 1130 -1568
rect 1132 -1569 1550 -1568
rect 1619 -1569 1634 -1568
rect 1647 -1569 1858 -1568
rect 1864 -1569 1914 -1568
rect 282 -1571 451 -1570
rect 457 -1571 713 -1570
rect 723 -1571 1210 -1570
rect 1213 -1571 1445 -1570
rect 1507 -1571 1634 -1570
rect 1647 -1571 1655 -1570
rect 1668 -1571 1697 -1570
rect 1787 -1571 1802 -1570
rect 1913 -1571 1942 -1570
rect 261 -1573 451 -1572
rect 464 -1573 689 -1572
rect 723 -1573 983 -1572
rect 1024 -1573 1074 -1572
rect 1150 -1573 1193 -1572
rect 1283 -1573 1627 -1572
rect 1654 -1573 1683 -1572
rect 1696 -1573 1844 -1572
rect 1941 -1573 2012 -1572
rect 261 -1575 1070 -1574
rect 1171 -1575 1242 -1574
rect 1311 -1575 1319 -1574
rect 1395 -1575 1403 -1574
rect 1444 -1575 1466 -1574
rect 1521 -1575 1529 -1574
rect 1542 -1575 1564 -1574
rect 1626 -1575 1711 -1574
rect 1787 -1575 1928 -1574
rect 65 -1577 1711 -1576
rect 1843 -1577 1921 -1576
rect 289 -1579 367 -1578
rect 418 -1579 850 -1578
rect 919 -1579 1508 -1578
rect 1521 -1579 1606 -1578
rect 296 -1581 360 -1580
rect 366 -1581 430 -1580
rect 443 -1581 654 -1580
rect 730 -1581 976 -1580
rect 1006 -1581 1683 -1580
rect 114 -1583 654 -1582
rect 772 -1583 801 -1582
rect 807 -1583 955 -1582
rect 968 -1583 990 -1582
rect 1024 -1583 1137 -1582
rect 1185 -1583 1249 -1582
rect 1290 -1583 1466 -1582
rect 1549 -1583 1557 -1582
rect 1563 -1583 1585 -1582
rect 1598 -1583 1928 -1582
rect 296 -1585 986 -1584
rect 989 -1585 1091 -1584
rect 1220 -1585 1249 -1584
rect 1290 -1585 1298 -1584
rect 1402 -1585 1417 -1584
rect 1535 -1585 1585 -1584
rect 1598 -1585 1641 -1584
rect 303 -1587 332 -1586
rect 422 -1587 458 -1586
rect 478 -1587 619 -1586
rect 765 -1587 773 -1586
rect 793 -1587 808 -1586
rect 817 -1587 1837 -1586
rect 212 -1589 423 -1588
rect 429 -1589 951 -1588
rect 1031 -1589 1151 -1588
rect 1164 -1589 1298 -1588
rect 1367 -1589 1536 -1588
rect 1570 -1589 1606 -1588
rect 170 -1591 213 -1590
rect 317 -1591 465 -1590
rect 478 -1591 514 -1590
rect 597 -1591 864 -1590
rect 922 -1591 1641 -1590
rect 317 -1593 612 -1592
rect 793 -1593 857 -1592
rect 884 -1593 923 -1592
rect 926 -1593 983 -1592
rect 1010 -1593 1032 -1592
rect 1059 -1593 1319 -1592
rect 1367 -1593 1389 -1592
rect 1416 -1593 1424 -1592
rect 79 -1595 1011 -1594
rect 1080 -1595 1165 -1594
rect 1195 -1595 1571 -1594
rect 331 -1597 388 -1596
rect 513 -1597 542 -1596
rect 611 -1597 741 -1596
rect 828 -1597 1137 -1596
rect 1220 -1597 1277 -1596
rect 1388 -1597 1452 -1596
rect 387 -1599 815 -1598
rect 856 -1599 892 -1598
rect 912 -1599 927 -1598
rect 933 -1599 976 -1598
rect 1080 -1599 1228 -1598
rect 1241 -1599 1816 -1598
rect 177 -1601 934 -1600
rect 940 -1601 1060 -1600
rect 1227 -1601 1410 -1600
rect 1423 -1601 1431 -1600
rect 1451 -1601 1473 -1600
rect 1815 -1601 1900 -1600
rect 352 -1603 1431 -1602
rect 1458 -1603 1473 -1602
rect 352 -1605 563 -1604
rect 870 -1605 1277 -1604
rect 1458 -1605 1480 -1604
rect 380 -1607 941 -1606
rect 1094 -1607 1410 -1606
rect 1479 -1607 1487 -1606
rect 380 -1609 493 -1608
rect 534 -1609 598 -1608
rect 786 -1609 871 -1608
rect 891 -1609 1179 -1608
rect 1206 -1609 1900 -1608
rect 394 -1611 493 -1610
rect 541 -1611 577 -1610
rect 744 -1611 787 -1610
rect 898 -1611 913 -1610
rect 1045 -1611 1095 -1610
rect 1244 -1611 1557 -1610
rect 173 -1613 745 -1612
rect 898 -1613 1067 -1612
rect 1087 -1613 1179 -1612
rect 1486 -1613 1501 -1612
rect 82 -1615 1088 -1614
rect 1500 -1615 1676 -1614
rect 394 -1617 836 -1616
rect 1017 -1617 1067 -1616
rect 1675 -1617 1739 -1616
rect 471 -1619 535 -1618
rect 562 -1619 1158 -1618
rect 1738 -1619 1746 -1618
rect 471 -1621 528 -1620
rect 779 -1621 1018 -1620
rect 1045 -1621 1336 -1620
rect 1745 -1621 1774 -1620
rect 408 -1623 528 -1622
rect 695 -1623 780 -1622
rect 1143 -1623 1158 -1622
rect 1759 -1623 1774 -1622
rect 408 -1625 591 -1624
rect 1052 -1625 1144 -1624
rect 1759 -1625 2008 -1624
rect 590 -1627 717 -1626
rect 1052 -1627 1893 -1626
rect 240 -1629 1893 -1628
rect 240 -1631 402 -1630
rect 716 -1631 759 -1630
rect 401 -1633 437 -1632
rect 737 -1633 759 -1632
rect 373 -1635 437 -1634
rect 625 -1635 738 -1634
rect 275 -1637 374 -1636
rect 604 -1637 626 -1636
rect 149 -1639 276 -1638
rect 604 -1639 640 -1638
rect 149 -1641 171 -1640
rect 632 -1641 640 -1640
rect 632 -1643 832 -1642
rect 9 -1654 664 -1653
rect 670 -1654 717 -1653
rect 737 -1654 1557 -1653
rect 1843 -1654 1935 -1653
rect 1937 -1654 1977 -1653
rect 9 -1656 129 -1655
rect 131 -1656 1102 -1655
rect 1206 -1656 1704 -1655
rect 1815 -1656 1844 -1655
rect 1850 -1656 1935 -1655
rect 1941 -1656 1970 -1655
rect 44 -1658 80 -1657
rect 86 -1658 276 -1657
rect 324 -1658 559 -1657
rect 590 -1658 832 -1657
rect 842 -1658 1105 -1657
rect 1206 -1658 1291 -1657
rect 1332 -1658 1816 -1657
rect 1850 -1658 1858 -1657
rect 1944 -1658 1963 -1657
rect 37 -1660 45 -1659
rect 65 -1660 178 -1659
rect 180 -1660 360 -1659
rect 422 -1660 426 -1659
rect 485 -1660 685 -1659
rect 709 -1660 1396 -1659
rect 1468 -1660 1697 -1659
rect 1857 -1660 1865 -1659
rect 1948 -1660 1956 -1659
rect 37 -1662 59 -1661
rect 68 -1662 535 -1661
rect 541 -1662 773 -1661
rect 793 -1662 1039 -1661
rect 1055 -1662 1298 -1661
rect 1332 -1662 1417 -1661
rect 1468 -1662 1711 -1661
rect 1822 -1662 1865 -1661
rect 1941 -1662 1949 -1661
rect 58 -1664 430 -1663
rect 478 -1664 486 -1663
rect 534 -1664 626 -1663
rect 688 -1664 710 -1663
rect 712 -1664 1039 -1663
rect 1076 -1664 1354 -1663
rect 1395 -1664 1403 -1663
rect 1416 -1664 1424 -1663
rect 1500 -1664 1781 -1663
rect 1794 -1664 1823 -1663
rect 72 -1666 83 -1665
rect 89 -1666 1690 -1665
rect 1696 -1666 1760 -1665
rect 1766 -1666 1795 -1665
rect 72 -1668 661 -1667
rect 688 -1668 990 -1667
rect 1083 -1668 1921 -1667
rect 117 -1670 1165 -1669
rect 1220 -1670 1291 -1669
rect 1297 -1670 1466 -1669
rect 1556 -1670 1564 -1669
rect 1640 -1670 1690 -1669
rect 1731 -1670 1760 -1669
rect 1906 -1670 1921 -1669
rect 128 -1672 969 -1671
rect 985 -1672 1214 -1671
rect 1286 -1672 1928 -1671
rect 156 -1674 395 -1673
rect 422 -1674 500 -1673
rect 523 -1674 1781 -1673
rect 1899 -1674 1907 -1673
rect 114 -1676 395 -1675
rect 429 -1676 437 -1675
rect 499 -1676 1284 -1675
rect 1335 -1676 1739 -1675
rect 1752 -1676 1767 -1675
rect 1892 -1676 1900 -1675
rect 114 -1678 444 -1677
rect 541 -1678 741 -1677
rect 751 -1678 1403 -1677
rect 1423 -1678 1438 -1677
rect 1521 -1678 1564 -1677
rect 1619 -1678 1641 -1677
rect 1654 -1678 1704 -1677
rect 1717 -1678 1732 -1677
rect 1752 -1678 1774 -1677
rect 1787 -1678 1893 -1677
rect 149 -1680 437 -1679
rect 443 -1680 647 -1679
rect 660 -1680 941 -1679
rect 943 -1680 1725 -1679
rect 121 -1682 150 -1681
rect 156 -1682 318 -1681
rect 324 -1682 409 -1681
rect 481 -1682 752 -1681
rect 765 -1682 864 -1681
rect 901 -1682 1025 -1681
rect 1087 -1682 1473 -1681
rect 1493 -1682 1620 -1681
rect 1626 -1682 1739 -1681
rect 121 -1684 815 -1683
rect 828 -1684 1112 -1683
rect 1185 -1684 1214 -1683
rect 1241 -1684 1655 -1683
rect 1675 -1684 1788 -1683
rect 184 -1686 668 -1685
rect 702 -1686 794 -1685
rect 831 -1686 1319 -1685
rect 1339 -1686 1438 -1685
rect 1472 -1686 1480 -1685
rect 1591 -1686 1627 -1685
rect 1682 -1686 1711 -1685
rect 187 -1688 1277 -1687
rect 1311 -1688 1494 -1687
rect 1542 -1688 1592 -1687
rect 1668 -1688 1683 -1687
rect 100 -1690 1543 -1689
rect 1661 -1690 1669 -1689
rect 2 -1692 101 -1691
rect 201 -1692 650 -1691
rect 716 -1692 1074 -1691
rect 1101 -1692 1676 -1691
rect 205 -1694 209 -1693
rect 254 -1694 398 -1693
rect 408 -1694 563 -1693
rect 583 -1694 626 -1693
rect 639 -1694 815 -1693
rect 842 -1694 878 -1693
rect 919 -1694 1585 -1693
rect 1661 -1694 1746 -1693
rect 191 -1696 255 -1695
rect 275 -1696 451 -1695
rect 520 -1696 703 -1695
rect 737 -1696 811 -1695
rect 863 -1696 913 -1695
rect 919 -1696 1210 -1695
rect 1241 -1696 1501 -1695
rect 1584 -1696 1599 -1695
rect 1745 -1696 1837 -1695
rect 191 -1698 419 -1697
rect 576 -1698 640 -1697
rect 740 -1698 1431 -1697
rect 1479 -1698 1487 -1697
rect 1598 -1698 1613 -1697
rect 1808 -1698 1837 -1697
rect 198 -1700 451 -1699
rect 527 -1700 577 -1699
rect 583 -1700 682 -1699
rect 768 -1700 990 -1699
rect 1024 -1700 1137 -1699
rect 1185 -1700 1200 -1699
rect 1244 -1700 1718 -1699
rect 198 -1702 850 -1701
rect 877 -1702 962 -1701
rect 968 -1702 1046 -1701
rect 1073 -1702 1830 -1701
rect 205 -1704 493 -1703
rect 527 -1704 633 -1703
rect 681 -1704 1774 -1703
rect 219 -1706 1046 -1705
rect 1129 -1706 1809 -1705
rect 219 -1708 262 -1707
rect 317 -1708 339 -1707
rect 359 -1708 458 -1707
rect 492 -1708 731 -1707
rect 772 -1708 1067 -1707
rect 1122 -1708 1130 -1707
rect 1132 -1708 1830 -1707
rect 261 -1710 507 -1709
rect 590 -1710 598 -1709
rect 604 -1710 668 -1709
rect 786 -1710 1284 -1709
rect 1311 -1710 1466 -1709
rect 1612 -1710 1648 -1709
rect 310 -1712 339 -1711
rect 373 -1712 419 -1711
rect 425 -1712 787 -1711
rect 849 -1712 899 -1711
rect 912 -1712 927 -1711
rect 933 -1712 1522 -1711
rect 282 -1714 311 -1713
rect 373 -1714 402 -1713
rect 457 -1714 465 -1713
rect 506 -1714 724 -1713
rect 922 -1714 948 -1713
rect 961 -1714 1004 -1713
rect 1041 -1714 1123 -1713
rect 1136 -1714 1158 -1713
rect 1199 -1714 1249 -1713
rect 1269 -1714 1277 -1713
rect 1318 -1714 1928 -1713
rect 142 -1716 402 -1715
rect 569 -1716 605 -1715
rect 632 -1716 699 -1715
rect 723 -1716 871 -1715
rect 943 -1716 1088 -1715
rect 1157 -1716 1193 -1715
rect 1244 -1716 1606 -1715
rect 93 -1718 143 -1717
rect 194 -1718 1606 -1717
rect 93 -1720 601 -1719
rect 653 -1720 927 -1719
rect 947 -1720 983 -1719
rect 996 -1720 1004 -1719
rect 1066 -1720 1151 -1719
rect 1192 -1720 1347 -1719
rect 1353 -1720 1634 -1719
rect 16 -1722 983 -1721
rect 1010 -1722 1634 -1721
rect 16 -1724 171 -1723
rect 184 -1724 1011 -1723
rect 1150 -1724 1179 -1723
rect 1248 -1724 1326 -1723
rect 1339 -1724 1515 -1723
rect 170 -1726 269 -1725
rect 397 -1726 822 -1725
rect 870 -1726 906 -1725
rect 971 -1726 1487 -1725
rect 1507 -1726 1515 -1725
rect 233 -1728 465 -1727
rect 569 -1728 612 -1727
rect 646 -1728 997 -1727
rect 1171 -1728 1179 -1727
rect 1227 -1728 1326 -1727
rect 1356 -1728 1725 -1727
rect 233 -1730 304 -1729
rect 597 -1730 1165 -1729
rect 1220 -1730 1357 -1729
rect 1388 -1730 1431 -1729
rect 1507 -1730 1578 -1729
rect 240 -1732 304 -1731
rect 611 -1732 619 -1731
rect 653 -1732 1305 -1731
rect 1388 -1732 1445 -1731
rect 226 -1734 619 -1733
rect 821 -1734 836 -1733
rect 891 -1734 1347 -1733
rect 1444 -1734 1536 -1733
rect 226 -1736 332 -1735
rect 807 -1736 836 -1735
rect 891 -1736 955 -1735
rect 1080 -1736 1172 -1735
rect 1227 -1736 1235 -1735
rect 1269 -1736 1361 -1735
rect 1528 -1736 1536 -1735
rect 240 -1738 416 -1737
rect 898 -1738 1578 -1737
rect 247 -1740 283 -1739
rect 331 -1740 353 -1739
rect 905 -1740 976 -1739
rect 1234 -1740 1368 -1739
rect 1528 -1740 1550 -1739
rect 247 -1742 346 -1741
rect 352 -1742 549 -1741
rect 933 -1742 1081 -1741
rect 1304 -1742 1648 -1741
rect 268 -1744 367 -1743
rect 513 -1744 549 -1743
rect 954 -1744 1879 -1743
rect 23 -1746 367 -1745
rect 513 -1746 675 -1745
rect 975 -1746 1018 -1745
rect 1307 -1746 1879 -1745
rect 23 -1748 545 -1747
rect 674 -1748 780 -1747
rect 1052 -1748 1308 -1747
rect 1360 -1748 1364 -1747
rect 1367 -1748 1459 -1747
rect 289 -1750 346 -1749
rect 744 -1750 1018 -1749
rect 1052 -1750 1109 -1749
rect 1374 -1750 1459 -1749
rect 289 -1752 381 -1751
rect 744 -1752 759 -1751
rect 779 -1752 1032 -1751
rect 1374 -1752 1382 -1751
rect 1409 -1752 1550 -1751
rect 107 -1754 381 -1753
rect 758 -1754 885 -1753
rect 1031 -1754 1095 -1753
rect 1115 -1754 1410 -1753
rect 107 -1756 136 -1755
rect 695 -1756 1095 -1755
rect 1115 -1756 1144 -1755
rect 1381 -1756 1847 -1755
rect 135 -1758 164 -1757
rect 565 -1758 1144 -1757
rect 163 -1760 213 -1759
rect 695 -1760 1060 -1759
rect 212 -1762 388 -1761
rect 1059 -1762 1256 -1761
rect 296 -1764 388 -1763
rect 516 -1764 1256 -1763
rect 296 -1766 472 -1765
rect 30 -1768 472 -1767
rect 30 -1770 556 -1769
rect 555 -1772 888 -1771
rect 65 -1783 76 -1782
rect 93 -1783 146 -1782
rect 170 -1783 524 -1782
rect 527 -1783 531 -1782
rect 555 -1783 794 -1782
rect 810 -1783 1928 -1782
rect 1955 -1783 1998 -1782
rect 2011 -1783 2019 -1782
rect 65 -1785 276 -1784
rect 282 -1785 482 -1784
rect 506 -1785 556 -1784
rect 597 -1785 871 -1784
rect 884 -1785 1690 -1784
rect 1878 -1785 1956 -1784
rect 1962 -1785 2019 -1784
rect 93 -1787 108 -1786
rect 114 -1787 192 -1786
rect 198 -1787 878 -1786
rect 884 -1787 2005 -1786
rect 107 -1789 500 -1788
rect 527 -1789 1074 -1788
rect 1080 -1789 1690 -1788
rect 1878 -1789 1942 -1788
rect 1969 -1789 2026 -1788
rect 114 -1791 213 -1790
rect 254 -1791 692 -1790
rect 695 -1791 927 -1790
rect 943 -1791 1494 -1790
rect 1566 -1791 1886 -1790
rect 1892 -1791 1963 -1790
rect 58 -1793 213 -1792
rect 254 -1793 290 -1792
rect 310 -1793 808 -1792
rect 870 -1793 934 -1792
rect 985 -1793 1571 -1792
rect 1829 -1793 1886 -1792
rect 1899 -1793 1970 -1792
rect 16 -1795 59 -1794
rect 128 -1795 136 -1794
rect 138 -1795 290 -1794
rect 352 -1795 489 -1794
rect 499 -1795 626 -1794
rect 649 -1795 815 -1794
rect 898 -1795 1039 -1794
rect 1059 -1795 1077 -1794
rect 1080 -1795 1088 -1794
rect 1090 -1795 1207 -1794
rect 1209 -1795 1627 -1794
rect 1731 -1795 1830 -1794
rect 1843 -1795 1893 -1794
rect 1906 -1795 1984 -1794
rect 9 -1797 136 -1796
rect 142 -1797 311 -1796
rect 352 -1797 360 -1796
rect 366 -1797 563 -1796
rect 583 -1797 598 -1796
rect 600 -1797 703 -1796
rect 719 -1797 731 -1796
rect 751 -1797 878 -1796
rect 908 -1797 1095 -1796
rect 1104 -1797 1445 -1796
rect 1468 -1797 1921 -1796
rect 16 -1799 52 -1798
rect 121 -1799 626 -1798
rect 639 -1799 703 -1798
rect 730 -1799 1382 -1798
rect 1409 -1799 1991 -1798
rect 37 -1801 52 -1800
rect 79 -1801 122 -1800
rect 131 -1801 367 -1800
rect 387 -1801 640 -1800
rect 681 -1801 794 -1800
rect 814 -1801 843 -1800
rect 954 -1801 1039 -1800
rect 1059 -1801 1291 -1800
rect 1304 -1801 1774 -1800
rect 1850 -1801 1907 -1800
rect 1913 -1801 1921 -1800
rect 37 -1803 143 -1802
rect 156 -1803 283 -1802
rect 387 -1803 510 -1802
rect 562 -1803 605 -1802
rect 632 -1803 682 -1802
rect 684 -1803 937 -1802
rect 1017 -1803 1095 -1802
rect 1104 -1803 1214 -1802
rect 1244 -1803 1641 -1802
rect 1717 -1803 1774 -1802
rect 1815 -1803 1851 -1802
rect 1871 -1803 1942 -1802
rect 79 -1805 654 -1804
rect 765 -1805 843 -1804
rect 1073 -1805 1172 -1804
rect 1248 -1805 1291 -1804
rect 1304 -1805 1438 -1804
rect 1535 -1805 1844 -1804
rect 156 -1807 409 -1806
rect 415 -1807 920 -1806
rect 1108 -1807 1977 -1806
rect 170 -1809 983 -1808
rect 1111 -1809 1193 -1808
rect 1269 -1809 1354 -1808
rect 1360 -1809 1739 -1808
rect 1745 -1809 1900 -1808
rect 177 -1811 276 -1810
rect 401 -1811 941 -1810
rect 1136 -1811 1172 -1810
rect 1185 -1811 1249 -1810
rect 1262 -1811 1270 -1810
rect 1283 -1811 1361 -1810
rect 1363 -1811 1928 -1810
rect 177 -1813 395 -1812
rect 404 -1813 416 -1812
rect 429 -1813 514 -1812
rect 583 -1813 1102 -1812
rect 1115 -1813 1137 -1812
rect 1150 -1813 1186 -1812
rect 1276 -1813 1284 -1812
rect 1307 -1813 1788 -1812
rect 1794 -1813 1872 -1812
rect 191 -1815 220 -1814
rect 240 -1815 395 -1814
rect 408 -1815 1126 -1814
rect 1150 -1815 1445 -1814
rect 1535 -1815 1781 -1814
rect 1822 -1815 1914 -1814
rect 201 -1817 297 -1816
rect 380 -1817 402 -1816
rect 429 -1817 549 -1816
rect 604 -1817 724 -1816
rect 751 -1817 1109 -1816
rect 1157 -1817 1193 -1816
rect 1311 -1817 1494 -1816
rect 1563 -1817 1571 -1816
rect 1577 -1817 1746 -1816
rect 1759 -1817 1781 -1816
rect 1801 -1817 1823 -1816
rect 187 -1819 1802 -1818
rect 219 -1821 444 -1820
rect 450 -1821 696 -1820
rect 723 -1821 829 -1820
rect 831 -1821 1438 -1820
rect 1598 -1821 1816 -1820
rect 23 -1823 829 -1822
rect 863 -1823 1312 -1822
rect 1318 -1823 1704 -1822
rect 1738 -1823 1753 -1822
rect 1766 -1823 1795 -1822
rect 23 -1825 615 -1824
rect 632 -1825 668 -1824
rect 765 -1825 864 -1824
rect 891 -1825 941 -1824
rect 975 -1825 1158 -1824
rect 1164 -1825 1214 -1824
rect 1321 -1825 1627 -1824
rect 1654 -1825 1718 -1824
rect 72 -1827 451 -1826
rect 464 -1827 521 -1826
rect 541 -1827 549 -1826
rect 576 -1827 668 -1826
rect 768 -1827 1459 -1826
rect 1486 -1827 1767 -1826
rect 44 -1829 73 -1828
rect 100 -1829 976 -1828
rect 1024 -1829 1165 -1828
rect 1178 -1829 1263 -1828
rect 1325 -1829 1382 -1828
rect 1409 -1829 1550 -1828
rect 1598 -1829 1662 -1828
rect 1696 -1829 1704 -1828
rect 30 -1831 1025 -1830
rect 1083 -1831 1753 -1830
rect 30 -1833 227 -1832
rect 240 -1833 339 -1832
rect 373 -1833 444 -1832
rect 464 -1833 612 -1832
rect 772 -1833 1018 -1832
rect 1143 -1833 1179 -1832
rect 1255 -1833 1326 -1832
rect 1339 -1833 1578 -1832
rect 1605 -1833 1641 -1832
rect 1661 -1833 1837 -1832
rect 44 -1835 398 -1834
rect 436 -1835 654 -1834
rect 772 -1835 997 -1834
rect 1122 -1835 1144 -1834
rect 1199 -1835 1256 -1834
rect 1430 -1835 1732 -1834
rect 1808 -1835 1837 -1834
rect 184 -1837 1319 -1836
rect 1451 -1837 1459 -1836
rect 1479 -1837 1487 -1836
rect 1633 -1837 1655 -1836
rect 1682 -1837 1697 -1836
rect 1710 -1837 1809 -1836
rect 163 -1839 185 -1838
rect 205 -1839 374 -1838
rect 380 -1839 423 -1838
rect 485 -1839 542 -1838
rect 558 -1839 1200 -1838
rect 1234 -1839 1340 -1838
rect 1367 -1839 1480 -1838
rect 1542 -1839 1711 -1838
rect 163 -1841 517 -1840
rect 520 -1841 689 -1840
rect 891 -1841 1242 -1840
rect 1367 -1841 1375 -1840
rect 1388 -1841 1452 -1840
rect 1556 -1841 1634 -1840
rect 1668 -1841 1683 -1840
rect 205 -1843 234 -1842
rect 261 -1843 360 -1842
rect 478 -1843 1543 -1842
rect 1556 -1843 1945 -1842
rect 149 -1845 262 -1844
rect 296 -1845 479 -1844
rect 485 -1845 1788 -1844
rect 149 -1847 888 -1846
rect 912 -1847 920 -1846
rect 933 -1847 1760 -1846
rect 226 -1849 346 -1848
rect 492 -1849 888 -1848
rect 912 -1849 962 -1848
rect 996 -1849 1004 -1848
rect 1045 -1849 1431 -1848
rect 1647 -1849 1669 -1848
rect 233 -1851 269 -1850
rect 331 -1851 437 -1850
rect 492 -1851 619 -1850
rect 779 -1851 1004 -1850
rect 1031 -1851 1046 -1850
rect 1122 -1851 1865 -1850
rect 86 -1853 269 -1852
rect 324 -1853 332 -1852
rect 513 -1853 1154 -1852
rect 1220 -1853 1235 -1852
rect 1241 -1853 1466 -1852
rect 1612 -1853 1648 -1852
rect 86 -1855 1224 -1854
rect 1374 -1855 1396 -1854
rect 1423 -1855 1613 -1854
rect 247 -1857 346 -1856
rect 530 -1857 1116 -1856
rect 1346 -1857 1396 -1856
rect 1416 -1857 1424 -1856
rect 1465 -1857 1529 -1856
rect 247 -1859 2015 -1858
rect 317 -1861 325 -1860
rect 579 -1861 1550 -1860
rect 317 -1863 458 -1862
rect 611 -1863 1606 -1862
rect 198 -1865 458 -1864
rect 618 -1865 787 -1864
rect 905 -1865 962 -1864
rect 1031 -1865 1067 -1864
rect 1111 -1865 1865 -1864
rect 422 -1867 906 -1866
rect 954 -1867 1221 -1866
rect 1297 -1867 1347 -1866
rect 1388 -1867 1403 -1866
rect 1416 -1867 1935 -1866
rect 779 -1869 857 -1868
rect 1052 -1869 1067 -1868
rect 1227 -1869 1298 -1868
rect 1332 -1869 1403 -1868
rect 1528 -1869 1592 -1868
rect 1857 -1869 1935 -1868
rect 61 -1871 1228 -1870
rect 1507 -1871 1592 -1870
rect 68 -1873 1858 -1872
rect 103 -1875 857 -1874
rect 989 -1875 1053 -1874
rect 1507 -1875 1515 -1874
rect 534 -1877 990 -1876
rect 1472 -1877 1515 -1876
rect 534 -1879 759 -1878
rect 786 -1879 850 -1878
rect 1472 -1879 1676 -1878
rect 674 -1881 850 -1880
rect 1675 -1881 1725 -1880
rect 418 -1883 1725 -1882
rect 674 -1885 710 -1884
rect 737 -1885 1333 -1884
rect 565 -1887 710 -1886
rect 758 -1887 822 -1886
rect 646 -1889 738 -1888
rect 821 -1889 836 -1888
rect 569 -1891 647 -1890
rect 800 -1891 836 -1890
rect 471 -1893 570 -1892
rect 716 -1893 801 -1892
rect 471 -1895 1949 -1894
rect 716 -1897 927 -1896
rect 1563 -1897 1949 -1896
rect 2 -1908 227 -1907
rect 313 -1908 451 -1907
rect 478 -1908 556 -1907
rect 562 -1908 577 -1907
rect 614 -1908 990 -1907
rect 1024 -1908 1382 -1907
rect 1454 -1908 1872 -1907
rect 5 -1910 69 -1909
rect 79 -1910 510 -1909
rect 537 -1910 1116 -1909
rect 1153 -1910 1809 -1909
rect 1871 -1910 1900 -1909
rect 9 -1912 38 -1911
rect 44 -1912 139 -1911
rect 142 -1912 1445 -1911
rect 1535 -1912 1809 -1911
rect 1899 -1912 1949 -1911
rect 37 -1914 542 -1913
rect 555 -1914 738 -1913
rect 744 -1914 1102 -1913
rect 1108 -1914 1298 -1913
rect 1367 -1914 1382 -1913
rect 1444 -1914 1452 -1913
rect 1535 -1914 2012 -1913
rect 44 -1916 290 -1915
rect 317 -1916 745 -1915
rect 828 -1916 934 -1915
rect 964 -1916 1312 -1915
rect 1451 -1916 1529 -1915
rect 1563 -1916 1571 -1915
rect 1948 -1916 1977 -1915
rect 58 -1918 696 -1917
rect 716 -1918 738 -1917
rect 772 -1918 1571 -1917
rect 1976 -1918 2019 -1917
rect 79 -1920 472 -1919
rect 481 -1920 1242 -1919
rect 1283 -1920 1312 -1919
rect 1528 -1920 1753 -1919
rect 23 -1922 472 -1921
rect 485 -1922 909 -1921
rect 919 -1922 934 -1921
rect 982 -1922 1634 -1921
rect 23 -1924 115 -1923
rect 135 -1924 727 -1923
rect 730 -1924 895 -1923
rect 905 -1924 1816 -1923
rect 86 -1926 290 -1925
rect 317 -1926 759 -1925
rect 779 -1926 906 -1925
rect 982 -1926 1137 -1925
rect 1143 -1926 1242 -1925
rect 1293 -1926 1844 -1925
rect 100 -1928 269 -1927
rect 338 -1928 829 -1927
rect 845 -1928 1158 -1927
rect 1199 -1928 1368 -1927
rect 1566 -1928 1585 -1927
rect 1633 -1928 1655 -1927
rect 1815 -1928 1823 -1927
rect 1843 -1928 1886 -1927
rect 100 -1930 528 -1929
rect 562 -1930 584 -1929
rect 632 -1930 769 -1929
rect 779 -1930 857 -1929
rect 880 -1930 1039 -1929
rect 1090 -1930 1991 -1929
rect 30 -1932 528 -1931
rect 583 -1932 598 -1931
rect 660 -1932 664 -1931
rect 688 -1932 1396 -1931
rect 1472 -1932 1655 -1931
rect 1822 -1932 1837 -1931
rect 1885 -1932 1928 -1931
rect 1990 -1932 2026 -1931
rect 30 -1934 514 -1933
rect 660 -1934 668 -1933
rect 681 -1934 689 -1933
rect 698 -1934 1284 -1933
rect 1297 -1934 1494 -1933
rect 1584 -1934 1606 -1933
rect 1836 -1934 1851 -1933
rect 1927 -1934 1956 -1933
rect 16 -1936 514 -1935
rect 674 -1936 682 -1935
rect 709 -1936 717 -1935
rect 719 -1936 815 -1935
rect 856 -1936 1081 -1935
rect 1094 -1936 1116 -1935
rect 1129 -1936 1144 -1935
rect 1157 -1936 1172 -1935
rect 1206 -1936 1217 -1935
rect 1220 -1936 1732 -1935
rect 1955 -1936 1984 -1935
rect 65 -1938 633 -1937
rect 674 -1938 703 -1937
rect 709 -1938 1060 -1937
rect 1066 -1938 1081 -1937
rect 1094 -1938 1319 -1937
rect 1395 -1938 1501 -1937
rect 1661 -1938 1851 -1937
rect 103 -1940 976 -1939
rect 989 -1940 1032 -1939
rect 1052 -1940 1060 -1939
rect 1108 -1940 1515 -1939
rect 16 -1942 1032 -1941
rect 1136 -1942 1179 -1941
rect 1206 -1942 1522 -1941
rect 107 -1944 115 -1943
rect 135 -1944 388 -1943
rect 401 -1944 1210 -1943
rect 1220 -1944 1417 -1943
rect 1472 -1944 1543 -1943
rect 93 -1946 388 -1945
rect 415 -1946 542 -1945
rect 639 -1946 703 -1945
rect 730 -1946 1879 -1945
rect 51 -1948 94 -1947
rect 107 -1948 986 -1947
rect 1003 -1948 1067 -1947
rect 1164 -1948 1200 -1947
rect 1223 -1948 1921 -1947
rect 51 -1950 692 -1949
rect 733 -1950 1753 -1949
rect 1878 -1950 1907 -1949
rect 1920 -1950 1998 -1949
rect 142 -1952 1830 -1951
rect 1906 -1952 1935 -1951
rect 145 -1954 241 -1953
rect 408 -1954 416 -1953
rect 464 -1954 640 -1953
rect 758 -1954 962 -1953
rect 1010 -1954 1025 -1953
rect 1027 -1954 1802 -1953
rect 1934 -1954 1963 -1953
rect 86 -1956 146 -1955
rect 198 -1956 262 -1955
rect 408 -1956 752 -1955
rect 800 -1956 1053 -1955
rect 1164 -1956 1249 -1955
rect 1262 -1956 1501 -1955
rect 1521 -1956 1550 -1955
rect 1787 -1956 1830 -1955
rect 170 -1958 262 -1957
rect 464 -1958 776 -1957
rect 807 -1958 1039 -1957
rect 1171 -1958 1256 -1957
rect 1265 -1958 1732 -1957
rect 1794 -1958 1802 -1957
rect 170 -1960 776 -1959
rect 807 -1960 836 -1959
rect 849 -1960 1130 -1959
rect 1178 -1960 1186 -1959
rect 1216 -1960 1550 -1959
rect 1598 -1960 1795 -1959
rect 198 -1962 1263 -1961
rect 1290 -1962 1319 -1961
rect 1416 -1962 1424 -1961
rect 1479 -1962 1515 -1961
rect 1542 -1962 1557 -1961
rect 212 -1964 244 -1963
rect 268 -1964 1291 -1963
rect 1409 -1964 1424 -1963
rect 1465 -1964 1557 -1963
rect 184 -1966 213 -1965
rect 226 -1966 304 -1965
rect 485 -1966 654 -1965
rect 814 -1966 1333 -1965
rect 1388 -1966 1410 -1965
rect 1486 -1966 1494 -1965
rect 1507 -1966 1599 -1965
rect 184 -1968 192 -1967
rect 205 -1968 304 -1967
rect 457 -1968 654 -1967
rect 821 -1968 836 -1967
rect 849 -1968 1074 -1967
rect 1087 -1968 1466 -1967
rect 1486 -1968 1648 -1967
rect 163 -1970 192 -1969
rect 205 -1970 580 -1969
rect 618 -1970 752 -1969
rect 793 -1970 1074 -1969
rect 1087 -1970 1354 -1969
rect 1360 -1970 1508 -1969
rect 1647 -1970 1690 -1969
rect 72 -1972 164 -1971
rect 341 -1972 619 -1971
rect 793 -1972 955 -1971
rect 961 -1972 1788 -1971
rect 61 -1974 73 -1973
rect 380 -1974 458 -1973
rect 499 -1974 598 -1973
rect 821 -1974 1193 -1973
rect 1237 -1974 1280 -1973
rect 1325 -1974 1333 -1973
rect 1374 -1974 1389 -1973
rect 1689 -1974 1760 -1973
rect 380 -1976 437 -1975
rect 443 -1976 500 -1975
rect 506 -1976 1249 -1975
rect 1269 -1976 1361 -1975
rect 247 -1978 437 -1977
rect 754 -1978 1270 -1977
rect 1276 -1978 1480 -1977
rect 177 -1980 1277 -1979
rect 1304 -1980 1326 -1979
rect 1339 -1980 1375 -1979
rect 177 -1982 367 -1981
rect 863 -1982 1004 -1981
rect 1150 -1982 1760 -1981
rect 247 -1984 325 -1983
rect 352 -1984 444 -1983
rect 611 -1984 1151 -1983
rect 1192 -1984 1914 -1983
rect 254 -1986 367 -1985
rect 611 -1986 818 -1985
rect 863 -1986 2005 -1985
rect 254 -1988 311 -1987
rect 324 -1988 423 -1987
rect 866 -1988 1963 -1987
rect 275 -1990 507 -1989
rect 877 -1990 976 -1989
rect 996 -1990 1011 -1989
rect 1255 -1990 1914 -1989
rect 275 -1992 871 -1991
rect 877 -1992 1578 -1991
rect 296 -1994 311 -1993
rect 345 -1994 423 -1993
rect 842 -1994 871 -1993
rect 884 -1994 1613 -1993
rect 121 -1996 297 -1995
rect 345 -1996 489 -1995
rect 604 -1996 885 -1995
rect 887 -1996 1984 -1995
rect 121 -1998 430 -1997
rect 604 -1998 1046 -1997
rect 1339 -1998 1347 -1997
rect 1577 -1998 1592 -1997
rect 1612 -1998 1676 -1997
rect 219 -2000 430 -1999
rect 842 -2000 1711 -1999
rect 219 -2002 535 -2001
rect 912 -2002 955 -2001
rect 968 -2002 997 -2001
rect 1017 -2002 1046 -2001
rect 1111 -2002 1711 -2001
rect 352 -2004 570 -2003
rect 800 -2004 969 -2003
rect 1017 -2004 1438 -2003
rect 1591 -2004 1669 -2003
rect 1675 -2004 1704 -2003
rect 492 -2006 570 -2005
rect 912 -2006 937 -2005
rect 1111 -2006 1354 -2005
rect 1402 -2006 1438 -2005
rect 1668 -2006 1697 -2005
rect 1703 -2006 1739 -2005
rect 359 -2008 493 -2007
rect 520 -2008 535 -2007
rect 723 -2008 1403 -2007
rect 1640 -2008 1697 -2007
rect 331 -2010 360 -2009
rect 394 -2010 521 -2009
rect 530 -2010 1739 -2009
rect 149 -2012 332 -2011
rect 723 -2012 1662 -2011
rect 149 -2014 223 -2013
rect 233 -2014 395 -2013
rect 919 -2014 1305 -2013
rect 1640 -2014 1683 -2013
rect 233 -2016 283 -2015
rect 922 -2016 1606 -2015
rect 1682 -2016 1725 -2015
rect 282 -2018 374 -2017
rect 926 -2018 1186 -2017
rect 1234 -2018 1347 -2017
rect 1724 -2018 1767 -2017
rect 373 -2020 1123 -2019
rect 1766 -2020 1774 -2019
rect 898 -2022 927 -2021
rect 940 -2022 1123 -2021
rect 1773 -2022 1781 -2021
rect 625 -2024 941 -2023
rect 1619 -2024 1781 -2023
rect 548 -2026 626 -2025
rect 786 -2026 899 -2025
rect 1619 -2026 1718 -2025
rect 548 -2028 647 -2027
rect 772 -2028 787 -2027
rect 1626 -2028 1718 -2027
rect 590 -2030 647 -2029
rect 1626 -2030 1865 -2029
rect 590 -2032 766 -2031
rect 1104 -2032 1865 -2031
rect 765 -2034 892 -2033
rect 891 -2036 1858 -2035
rect 1857 -2038 1893 -2037
rect 1892 -2040 1942 -2039
rect 1941 -2042 1970 -2041
rect 761 -2044 1970 -2043
rect 2 -2055 339 -2054
rect 352 -2055 727 -2054
rect 733 -2055 1102 -2054
rect 1108 -2055 1515 -2054
rect 1920 -2055 1977 -2054
rect 2 -2057 206 -2056
rect 219 -2057 538 -2056
rect 548 -2057 815 -2056
rect 817 -2057 983 -2056
rect 1087 -2057 1235 -2056
rect 1237 -2057 1494 -2056
rect 23 -2059 143 -2058
rect 149 -2059 220 -2058
rect 222 -2059 703 -2058
rect 723 -2059 927 -2058
rect 961 -2059 1501 -2058
rect 9 -2061 143 -2060
rect 177 -2061 241 -2060
rect 352 -2061 395 -2060
rect 401 -2061 703 -2060
rect 723 -2061 997 -2060
rect 1087 -2061 1186 -2060
rect 1241 -2061 1263 -2060
rect 1265 -2061 1851 -2060
rect 23 -2063 111 -2062
rect 117 -2063 1508 -2062
rect 1850 -2063 1928 -2062
rect 30 -2065 314 -2064
rect 394 -2065 710 -2064
rect 751 -2065 1130 -2064
rect 1139 -2065 1438 -2064
rect 1493 -2065 1606 -2064
rect 30 -2067 510 -2066
rect 520 -2067 650 -2066
rect 695 -2067 1039 -2066
rect 1101 -2067 1179 -2066
rect 1241 -2067 1305 -2066
rect 1360 -2067 1455 -2066
rect 1500 -2067 1760 -2066
rect 37 -2069 440 -2068
rect 450 -2069 500 -2068
rect 530 -2069 1403 -2068
rect 1437 -2069 1473 -2068
rect 1507 -2069 1711 -2068
rect 1759 -2069 1858 -2068
rect 51 -2071 699 -2070
rect 751 -2071 1109 -2070
rect 1129 -2071 1137 -2070
rect 1143 -2071 1263 -2070
rect 1290 -2071 1354 -2070
rect 1363 -2071 1830 -2070
rect 1857 -2071 1942 -2070
rect 51 -2073 262 -2072
rect 303 -2073 402 -2072
rect 408 -2073 839 -2072
rect 845 -2073 1515 -2072
rect 1605 -2073 1774 -2072
rect 1829 -2073 1900 -2072
rect 65 -2075 1403 -2074
rect 1710 -2075 1837 -2074
rect 1899 -2075 1991 -2074
rect 65 -2077 381 -2076
rect 415 -2077 731 -2076
rect 761 -2077 787 -2076
rect 807 -2077 815 -2076
rect 891 -2077 1032 -2076
rect 1038 -2077 1053 -2076
rect 1143 -2077 1214 -2076
rect 1255 -2077 1312 -2076
rect 1353 -2077 1571 -2076
rect 1773 -2077 1844 -2076
rect 44 -2079 381 -2078
rect 422 -2079 451 -2078
rect 492 -2079 500 -2078
rect 548 -2079 563 -2078
rect 583 -2079 808 -2078
rect 919 -2079 1599 -2078
rect 1843 -2079 1914 -2078
rect 44 -2081 87 -2080
rect 89 -2081 325 -2080
rect 422 -2081 976 -2080
rect 978 -2081 1375 -2080
rect 1475 -2081 1837 -2080
rect 68 -2083 472 -2082
rect 492 -2083 542 -2082
rect 562 -2083 1112 -2082
rect 1160 -2083 1305 -2082
rect 1311 -2083 1389 -2082
rect 1570 -2083 1662 -2082
rect 1717 -2083 1914 -2082
rect 79 -2085 83 -2084
rect 86 -2085 514 -2084
rect 583 -2085 647 -2084
rect 695 -2085 717 -2084
rect 730 -2085 965 -2084
rect 968 -2085 1480 -2084
rect 1661 -2085 1725 -2084
rect 79 -2087 136 -2086
rect 163 -2087 304 -2086
rect 436 -2087 514 -2086
rect 590 -2087 1399 -2086
rect 1479 -2087 1585 -2086
rect 1633 -2087 1725 -2086
rect 93 -2089 521 -2088
rect 593 -2089 745 -2088
rect 772 -2089 1067 -2088
rect 1171 -2089 1186 -2088
rect 1213 -2089 1340 -2088
rect 1374 -2089 1907 -2088
rect 33 -2091 745 -2090
rect 772 -2091 1112 -2090
rect 1171 -2091 1347 -2090
rect 1388 -2091 1459 -2090
rect 1584 -2091 1669 -2090
rect 1675 -2091 1907 -2090
rect 93 -2093 388 -2092
rect 467 -2093 969 -2092
rect 971 -2093 1424 -2092
rect 1458 -2093 1543 -2092
rect 1675 -2093 1732 -2092
rect 96 -2095 391 -2094
rect 597 -2095 850 -2094
rect 852 -2095 1634 -2094
rect 1703 -2095 1732 -2094
rect 16 -2097 850 -2096
rect 905 -2097 920 -2096
rect 922 -2097 1123 -2096
rect 1178 -2097 1417 -2096
rect 1542 -2097 1620 -2096
rect 1703 -2097 1795 -2096
rect 16 -2099 244 -2098
rect 247 -2099 262 -2098
rect 268 -2099 409 -2098
rect 506 -2099 598 -2098
rect 604 -2099 710 -2098
rect 779 -2099 892 -2098
rect 926 -2099 934 -2098
rect 954 -2099 962 -2098
rect 975 -2099 1011 -2098
rect 1031 -2099 1207 -2098
rect 1220 -2099 1340 -2098
rect 1346 -2099 1924 -2098
rect 128 -2101 150 -2100
rect 163 -2101 311 -2100
rect 324 -2101 591 -2100
rect 618 -2101 717 -2100
rect 786 -2101 1165 -2100
rect 1192 -2101 1207 -2100
rect 1220 -2101 1284 -2100
rect 1395 -2101 1424 -2100
rect 1619 -2101 1767 -2100
rect 1794 -2101 1816 -2100
rect 107 -2103 129 -2102
rect 135 -2103 157 -2102
rect 177 -2103 290 -2102
rect 341 -2103 619 -2102
rect 639 -2103 759 -2102
rect 884 -2103 906 -2102
rect 933 -2103 1018 -2102
rect 1052 -2103 1697 -2102
rect 1717 -2103 1746 -2102
rect 1766 -2103 1823 -2102
rect 156 -2105 185 -2104
rect 191 -2105 472 -2104
rect 506 -2105 780 -2104
rect 870 -2105 885 -2104
rect 954 -2105 1298 -2104
rect 1409 -2105 1669 -2104
rect 1696 -2105 1970 -2104
rect 184 -2107 843 -2106
rect 982 -2107 1004 -2106
rect 1010 -2107 1060 -2106
rect 1066 -2107 1746 -2106
rect 1815 -2107 1893 -2106
rect 191 -2109 360 -2108
rect 485 -2109 843 -2108
rect 989 -2109 1018 -2108
rect 1059 -2109 1158 -2108
rect 1192 -2109 1326 -2108
rect 1409 -2109 1466 -2108
rect 1822 -2109 1949 -2108
rect 198 -2111 311 -2110
rect 485 -2111 570 -2110
rect 576 -2111 605 -2110
rect 611 -2111 1165 -2110
rect 1248 -2111 1417 -2110
rect 1465 -2111 1578 -2110
rect 1892 -2111 1984 -2110
rect 198 -2113 227 -2112
rect 236 -2113 864 -2112
rect 989 -2113 1046 -2112
rect 1115 -2113 1123 -2112
rect 1157 -2113 1879 -2112
rect 205 -2115 972 -2114
rect 996 -2115 1025 -2114
rect 1045 -2115 1378 -2114
rect 1577 -2115 1809 -2114
rect 226 -2117 234 -2116
rect 247 -2117 346 -2116
rect 527 -2117 1284 -2116
rect 1325 -2117 1382 -2116
rect 1738 -2117 1879 -2116
rect 212 -2119 234 -2118
rect 268 -2119 374 -2118
rect 527 -2119 878 -2118
rect 1003 -2119 1074 -2118
rect 1115 -2119 1200 -2118
rect 1248 -2119 1368 -2118
rect 1381 -2119 1592 -2118
rect 1738 -2119 1802 -2118
rect 1808 -2119 1935 -2118
rect 145 -2121 1368 -2120
rect 1591 -2121 1683 -2120
rect 1801 -2121 1886 -2120
rect 170 -2123 374 -2122
rect 415 -2123 878 -2122
rect 1024 -2123 1522 -2122
rect 1682 -2123 1753 -2122
rect 1885 -2123 1963 -2122
rect 40 -2125 171 -2124
rect 212 -2125 367 -2124
rect 576 -2125 654 -2124
rect 737 -2125 759 -2124
rect 863 -2125 1070 -2124
rect 1073 -2125 1081 -2124
rect 1199 -2125 1277 -2124
rect 1486 -2125 1522 -2124
rect 1689 -2125 1753 -2124
rect 114 -2127 367 -2126
rect 611 -2127 626 -2126
rect 628 -2127 871 -2126
rect 894 -2127 1277 -2126
rect 1486 -2127 1550 -2126
rect 1689 -2127 1788 -2126
rect 282 -2129 360 -2128
rect 625 -2129 801 -2128
rect 1080 -2129 1781 -2128
rect 1787 -2129 1872 -2128
rect 100 -2131 283 -2130
rect 289 -2131 867 -2130
rect 1255 -2131 1361 -2130
rect 1549 -2131 1557 -2130
rect 1780 -2131 1865 -2130
rect 1871 -2131 1956 -2130
rect 100 -2133 1452 -2132
rect 1556 -2133 1648 -2132
rect 296 -2135 570 -2134
rect 639 -2135 857 -2134
rect 1269 -2135 1298 -2134
rect 1451 -2135 1599 -2134
rect 1612 -2135 1648 -2134
rect 254 -2137 297 -2136
rect 317 -2137 857 -2136
rect 1269 -2137 1333 -2136
rect 82 -2139 255 -2138
rect 317 -2139 332 -2138
rect 345 -2139 444 -2138
rect 646 -2139 1095 -2138
rect 1293 -2139 1613 -2138
rect 331 -2141 479 -2140
rect 653 -2141 675 -2140
rect 737 -2141 794 -2140
rect 800 -2141 822 -2140
rect 940 -2141 1095 -2140
rect 1332 -2141 1445 -2140
rect 443 -2143 766 -2142
rect 793 -2143 899 -2142
rect 1444 -2143 1536 -2142
rect 275 -2145 899 -2144
rect 1430 -2145 1536 -2144
rect 275 -2147 829 -2146
rect 1430 -2147 1529 -2146
rect 453 -2149 829 -2148
rect 1528 -2149 1641 -2148
rect 457 -2151 479 -2150
rect 667 -2151 941 -2150
rect 1626 -2151 1641 -2150
rect 457 -2153 661 -2152
rect 667 -2153 689 -2152
rect 754 -2153 1865 -2152
rect 555 -2155 689 -2154
rect 765 -2155 1396 -2154
rect 1563 -2155 1627 -2154
rect 555 -2157 633 -2156
rect 660 -2157 1091 -2156
rect 1563 -2157 1655 -2156
rect 404 -2159 1655 -2158
rect 429 -2161 633 -2160
rect 674 -2161 682 -2160
rect 821 -2161 836 -2160
rect 429 -2163 437 -2162
rect 534 -2163 836 -2162
rect 534 -2165 881 -2164
rect 681 -2167 1084 -2166
rect 880 -2169 1151 -2168
rect 1150 -2171 1228 -2170
rect 1227 -2173 1319 -2172
rect 912 -2175 1319 -2174
rect 121 -2177 913 -2176
rect 72 -2179 122 -2178
rect 72 -2181 465 -2180
rect 58 -2183 465 -2182
rect 58 -2185 388 -2184
rect 2 -2196 41 -2195
rect 58 -2196 216 -2195
rect 222 -2196 1140 -2195
rect 1178 -2196 1452 -2195
rect 1454 -2196 1809 -2195
rect 12 -2198 17 -2197
rect 33 -2198 521 -2197
rect 527 -2198 762 -2197
rect 817 -2198 1039 -2197
rect 1055 -2198 1319 -2197
rect 1360 -2198 1487 -2197
rect 1713 -2198 1725 -2197
rect 1727 -2198 1907 -2197
rect 16 -2200 304 -2199
rect 317 -2200 342 -2199
rect 352 -2200 626 -2199
rect 646 -2200 892 -2199
rect 950 -2200 1879 -2199
rect 37 -2202 850 -2201
rect 877 -2202 1298 -2201
rect 1318 -2202 1459 -2201
rect 1475 -2202 1760 -2201
rect 23 -2204 38 -2203
rect 44 -2204 59 -2203
rect 68 -2204 297 -2203
rect 303 -2204 563 -2203
rect 572 -2204 885 -2203
rect 891 -2204 1305 -2203
rect 1395 -2204 1788 -2203
rect 23 -2206 192 -2205
rect 254 -2206 1084 -2205
rect 1108 -2206 1263 -2205
rect 1276 -2206 1287 -2205
rect 1304 -2206 1823 -2205
rect 44 -2208 129 -2207
rect 163 -2208 1126 -2207
rect 1136 -2208 1221 -2207
rect 1255 -2208 1263 -2207
rect 1276 -2208 1326 -2207
rect 1395 -2208 1606 -2207
rect 1787 -2208 1795 -2207
rect 1822 -2208 1893 -2207
rect 107 -2210 276 -2209
rect 282 -2210 339 -2209
rect 352 -2210 598 -2209
rect 670 -2210 1886 -2209
rect 107 -2212 815 -2211
rect 877 -2212 920 -2211
rect 954 -2212 1298 -2211
rect 1325 -2212 1445 -2211
rect 1458 -2212 1480 -2211
rect 1605 -2212 1648 -2211
rect 1794 -2212 1900 -2211
rect 110 -2214 325 -2213
rect 387 -2214 479 -2213
rect 520 -2214 717 -2213
rect 786 -2214 1487 -2213
rect 1640 -2214 1648 -2213
rect 117 -2216 150 -2215
rect 163 -2216 248 -2215
rect 254 -2216 332 -2215
rect 408 -2216 479 -2215
rect 527 -2216 612 -2215
rect 737 -2216 787 -2215
rect 793 -2216 850 -2215
rect 880 -2216 1501 -2215
rect 1640 -2216 1746 -2215
rect 128 -2218 136 -2217
rect 170 -2218 388 -2217
rect 408 -2218 486 -2217
rect 544 -2218 913 -2217
rect 919 -2218 948 -2217
rect 968 -2218 1578 -2217
rect 1745 -2218 1914 -2217
rect 135 -2220 185 -2219
rect 191 -2220 976 -2219
rect 999 -2220 1536 -2219
rect 170 -2222 269 -2221
rect 289 -2222 325 -2221
rect 331 -2222 465 -2221
rect 471 -2222 1081 -2221
rect 1108 -2222 1284 -2221
rect 1353 -2222 1578 -2221
rect 79 -2224 290 -2223
rect 296 -2224 444 -2223
rect 457 -2224 510 -2223
rect 562 -2224 724 -2223
rect 737 -2224 864 -2223
rect 912 -2224 927 -2223
rect 968 -2224 1004 -2223
rect 1038 -2224 1102 -2223
rect 1111 -2224 1627 -2223
rect 51 -2226 458 -2225
rect 485 -2226 493 -2225
rect 569 -2226 717 -2225
rect 796 -2226 955 -2225
rect 971 -2226 1095 -2225
rect 1101 -2226 1151 -2225
rect 1178 -2226 1340 -2225
rect 1353 -2226 1417 -2225
rect 1444 -2226 1494 -2225
rect 1500 -2226 1592 -2225
rect 1626 -2226 1739 -2225
rect 30 -2228 52 -2227
rect 79 -2228 101 -2227
rect 142 -2228 269 -2227
rect 380 -2228 570 -2227
rect 590 -2228 1242 -2227
rect 1279 -2228 1550 -2227
rect 1591 -2228 1676 -2227
rect 1696 -2228 1739 -2227
rect 30 -2230 1025 -2229
rect 1031 -2230 1340 -2229
rect 1398 -2230 1872 -2229
rect 65 -2232 101 -2231
rect 177 -2232 472 -2231
rect 576 -2232 591 -2231
rect 597 -2232 633 -2231
rect 639 -2232 794 -2231
rect 926 -2232 962 -2231
rect 989 -2232 1004 -2231
rect 1010 -2232 1032 -2231
rect 1052 -2232 1361 -2231
rect 1402 -2232 1620 -2231
rect 1675 -2232 1830 -2231
rect 86 -2234 178 -2233
rect 184 -2234 220 -2233
rect 226 -2234 248 -2233
rect 261 -2234 318 -2233
rect 415 -2234 493 -2233
rect 506 -2234 962 -2233
rect 989 -2234 1018 -2233
rect 1024 -2234 1060 -2233
rect 1066 -2234 1186 -2233
rect 1188 -2234 1333 -2233
rect 1402 -2234 1431 -2233
rect 1479 -2234 1564 -2233
rect 1619 -2234 1704 -2233
rect 1829 -2234 1851 -2233
rect 86 -2236 395 -2235
rect 415 -2236 468 -2235
rect 506 -2236 773 -2235
rect 800 -2236 1060 -2235
rect 1087 -2236 1151 -2235
rect 1192 -2236 1242 -2235
rect 1283 -2236 1389 -2235
rect 1430 -2236 1515 -2235
rect 1535 -2236 1690 -2235
rect 1696 -2236 1816 -2235
rect 173 -2238 773 -2237
rect 1010 -2238 1165 -2237
rect 1192 -2238 1291 -2237
rect 1332 -2238 1424 -2237
rect 1493 -2238 1543 -2237
rect 1549 -2238 1774 -2237
rect 93 -2240 1424 -2239
rect 1514 -2240 1571 -2239
rect 1689 -2240 1844 -2239
rect 93 -2242 125 -2241
rect 198 -2242 283 -2241
rect 394 -2242 542 -2241
rect 576 -2242 948 -2241
rect 975 -2242 1291 -2241
rect 1542 -2242 1585 -2241
rect 1703 -2242 1858 -2241
rect 198 -2244 402 -2243
rect 429 -2244 633 -2243
rect 649 -2244 1417 -2243
rect 1563 -2244 1634 -2243
rect 1773 -2244 1802 -2243
rect 205 -2246 276 -2245
rect 345 -2246 402 -2245
rect 429 -2246 843 -2245
rect 1052 -2246 1347 -2245
rect 1570 -2246 1655 -2245
rect 72 -2248 346 -2247
rect 366 -2248 542 -2247
rect 611 -2248 654 -2247
rect 656 -2248 1095 -2247
rect 1122 -2248 1161 -2247
rect 1164 -2248 1235 -2247
rect 1346 -2248 1438 -2247
rect 1584 -2248 1662 -2247
rect 72 -2250 122 -2249
rect 156 -2250 206 -2249
rect 208 -2250 724 -2249
rect 744 -2250 1235 -2249
rect 1286 -2250 1662 -2249
rect 121 -2252 143 -2251
rect 156 -2252 1669 -2251
rect 212 -2254 381 -2253
rect 443 -2254 451 -2253
rect 618 -2254 801 -2253
rect 842 -2254 906 -2253
rect 1087 -2254 1116 -2253
rect 1122 -2254 1711 -2253
rect 212 -2256 759 -2255
rect 765 -2256 1018 -2255
rect 1115 -2256 1130 -2255
rect 1213 -2256 1256 -2255
rect 1293 -2256 1669 -2255
rect 1710 -2256 1760 -2255
rect 219 -2258 437 -2257
rect 450 -2258 500 -2257
rect 618 -2258 934 -2257
rect 1129 -2258 1207 -2257
rect 1220 -2258 1410 -2257
rect 1437 -2258 1522 -2257
rect 1633 -2258 1837 -2257
rect 226 -2260 241 -2259
rect 261 -2260 360 -2259
rect 366 -2260 556 -2259
rect 628 -2260 1207 -2259
rect 1409 -2260 1557 -2259
rect 236 -2262 1655 -2261
rect 240 -2264 1753 -2263
rect 310 -2266 360 -2265
rect 422 -2266 934 -2265
rect 1521 -2266 1683 -2265
rect 1752 -2266 1865 -2265
rect 159 -2268 311 -2267
rect 373 -2268 423 -2267
rect 436 -2268 871 -2267
rect 905 -2268 941 -2267
rect 1556 -2268 1613 -2267
rect 1682 -2268 1781 -2267
rect 373 -2270 549 -2269
rect 555 -2270 682 -2269
rect 709 -2270 864 -2269
rect 870 -2270 899 -2269
rect 940 -2270 983 -2269
rect 1612 -2270 1767 -2269
rect 390 -2272 1781 -2271
rect 499 -2274 535 -2273
rect 548 -2274 605 -2273
rect 639 -2274 759 -2273
rect 765 -2274 857 -2273
rect 898 -2274 1158 -2273
rect 1731 -2274 1767 -2273
rect 89 -2276 535 -2275
rect 604 -2276 675 -2275
rect 677 -2276 1389 -2275
rect 1472 -2276 1732 -2275
rect 653 -2278 1046 -2277
rect 1157 -2278 1228 -2277
rect 660 -2280 682 -2279
rect 702 -2280 710 -2279
rect 744 -2280 808 -2279
rect 821 -2280 857 -2279
rect 982 -2280 997 -2279
rect 1185 -2280 1473 -2279
rect 9 -2282 997 -2281
rect 1227 -2282 1312 -2281
rect 660 -2284 668 -2283
rect 674 -2284 1074 -2283
rect 1311 -2284 1382 -2283
rect 688 -2286 703 -2285
rect 751 -2286 1046 -2285
rect 1073 -2286 1144 -2285
rect 583 -2288 689 -2287
rect 751 -2288 825 -2287
rect 835 -2288 1382 -2287
rect 513 -2290 584 -2289
rect 807 -2290 829 -2289
rect 835 -2290 888 -2289
rect 978 -2290 1144 -2289
rect 65 -2292 514 -2291
rect 821 -2292 1214 -2291
rect 828 -2294 1200 -2293
rect 1199 -2296 1375 -2295
rect 1374 -2298 1466 -2297
rect 1465 -2300 1529 -2299
rect 1507 -2302 1529 -2301
rect 1507 -2304 1599 -2303
rect 1069 -2306 1599 -2305
rect 1069 -2308 1172 -2307
rect 1171 -2310 1270 -2309
rect 1269 -2312 1368 -2311
rect 149 -2314 1368 -2313
rect 9 -2325 171 -2324
rect 177 -2325 1728 -2324
rect 1731 -2325 1746 -2324
rect 1748 -2325 1823 -2324
rect 9 -2327 493 -2326
rect 499 -2327 818 -2326
rect 821 -2327 1207 -2326
rect 1216 -2327 1452 -2326
rect 1577 -2327 1732 -2326
rect 1755 -2327 1767 -2326
rect 1780 -2327 1802 -2326
rect 16 -2329 619 -2328
rect 625 -2329 1053 -2328
rect 1069 -2329 1256 -2328
rect 1276 -2329 1294 -2328
rect 1307 -2329 1459 -2328
rect 1738 -2329 1767 -2328
rect 1787 -2329 1809 -2328
rect 16 -2331 433 -2330
rect 439 -2331 458 -2330
rect 460 -2331 591 -2330
rect 625 -2331 906 -2330
rect 947 -2331 1039 -2330
rect 1052 -2331 1487 -2330
rect 1675 -2331 1739 -2330
rect 1759 -2331 1781 -2330
rect 1787 -2331 1795 -2330
rect 1797 -2331 1830 -2330
rect 30 -2333 115 -2332
rect 142 -2333 213 -2332
rect 233 -2333 388 -2332
rect 408 -2333 734 -2332
rect 793 -2333 808 -2332
rect 814 -2333 976 -2332
rect 996 -2333 1578 -2332
rect 1619 -2333 1676 -2332
rect 1759 -2333 1774 -2332
rect 30 -2335 150 -2334
rect 159 -2335 325 -2334
rect 352 -2335 668 -2334
rect 698 -2335 843 -2334
rect 863 -2335 976 -2334
rect 1020 -2335 1242 -2334
rect 1248 -2335 1277 -2334
rect 1290 -2335 1550 -2334
rect 1619 -2335 1690 -2334
rect 1717 -2335 1774 -2334
rect 44 -2337 237 -2336
rect 282 -2337 465 -2336
rect 471 -2337 619 -2336
rect 646 -2337 843 -2336
rect 884 -2337 1004 -2336
rect 1017 -2337 1242 -2336
rect 1321 -2337 1326 -2336
rect 1342 -2337 1711 -2336
rect 44 -2339 227 -2338
rect 303 -2339 531 -2338
rect 544 -2339 640 -2338
rect 646 -2339 888 -2338
rect 905 -2339 913 -2338
rect 947 -2339 962 -2338
rect 1038 -2339 1060 -2338
rect 1066 -2339 1291 -2338
rect 1370 -2339 1396 -2338
rect 1423 -2339 1452 -2338
rect 1486 -2339 1494 -2338
rect 1542 -2339 1550 -2338
rect 1633 -2339 1690 -2338
rect 51 -2341 1004 -2340
rect 1010 -2341 1060 -2340
rect 1066 -2341 1081 -2340
rect 1115 -2341 1515 -2340
rect 1521 -2341 1634 -2340
rect 37 -2343 1081 -2342
rect 1115 -2343 1179 -2342
rect 1188 -2343 1683 -2342
rect 37 -2345 241 -2344
rect 310 -2345 458 -2344
rect 467 -2345 1424 -2344
rect 1430 -2345 1459 -2344
rect 1465 -2345 1494 -2344
rect 1521 -2345 1557 -2344
rect 1640 -2345 1683 -2344
rect 51 -2347 244 -2346
rect 310 -2347 447 -2346
rect 450 -2347 465 -2346
rect 478 -2347 493 -2346
rect 534 -2347 962 -2346
rect 1010 -2347 1095 -2346
rect 1157 -2347 1161 -2346
rect 1171 -2347 1207 -2346
rect 1213 -2347 1256 -2346
rect 1283 -2347 1326 -2346
rect 1360 -2347 1396 -2346
rect 1437 -2347 1466 -2346
rect 1479 -2347 1515 -2346
rect 1640 -2347 1704 -2346
rect 58 -2349 83 -2348
rect 86 -2349 678 -2348
rect 723 -2349 997 -2348
rect 1017 -2349 1172 -2348
rect 1227 -2349 1249 -2348
rect 1339 -2349 1361 -2348
rect 1416 -2349 1438 -2348
rect 1444 -2349 1480 -2348
rect 1500 -2349 1557 -2348
rect 1661 -2349 1704 -2348
rect 58 -2351 220 -2350
rect 296 -2351 678 -2350
rect 772 -2351 1179 -2350
rect 1227 -2351 1795 -2350
rect 65 -2353 486 -2352
rect 513 -2353 535 -2352
rect 562 -2353 825 -2352
rect 831 -2353 1543 -2352
rect 1626 -2353 1662 -2352
rect 72 -2355 111 -2354
rect 114 -2355 199 -2354
rect 205 -2355 500 -2354
rect 541 -2355 563 -2354
rect 583 -2355 591 -2354
rect 604 -2355 640 -2354
rect 667 -2355 703 -2354
rect 772 -2355 787 -2354
rect 856 -2355 888 -2354
rect 912 -2355 927 -2354
rect 1055 -2355 1284 -2354
rect 1332 -2355 1445 -2354
rect 1591 -2355 1627 -2354
rect 72 -2357 101 -2356
rect 107 -2357 409 -2356
rect 415 -2357 472 -2356
rect 478 -2357 682 -2356
rect 786 -2357 808 -2356
rect 856 -2357 871 -2356
rect 926 -2357 1270 -2356
rect 1339 -2357 1648 -2356
rect 79 -2359 227 -2358
rect 289 -2359 297 -2358
rect 324 -2359 528 -2358
rect 541 -2359 689 -2358
rect 863 -2359 885 -2358
rect 1094 -2359 1165 -2358
rect 1199 -2359 1333 -2358
rect 1388 -2359 1417 -2358
rect 1528 -2359 1592 -2358
rect 1605 -2359 1648 -2358
rect 86 -2361 94 -2360
rect 96 -2361 1718 -2360
rect 93 -2363 125 -2362
rect 135 -2363 304 -2362
rect 352 -2363 1119 -2362
rect 1150 -2363 1200 -2362
rect 1269 -2363 1319 -2362
rect 1388 -2363 1697 -2362
rect 100 -2365 164 -2364
rect 170 -2365 423 -2364
rect 429 -2365 724 -2364
rect 870 -2365 878 -2364
rect 1150 -2365 1214 -2364
rect 1563 -2365 1606 -2364
rect 1654 -2365 1697 -2364
rect 121 -2367 514 -2366
rect 520 -2367 689 -2366
rect 877 -2367 941 -2366
rect 1157 -2367 1221 -2366
rect 1507 -2367 1564 -2366
rect 1598 -2367 1655 -2366
rect 107 -2369 941 -2368
rect 1083 -2369 1508 -2368
rect 1598 -2369 1669 -2368
rect 131 -2371 136 -2370
rect 142 -2371 1000 -2370
rect 1164 -2371 1613 -2370
rect 149 -2373 577 -2372
rect 583 -2373 969 -2372
rect 1192 -2373 1221 -2372
rect 1535 -2373 1669 -2372
rect 156 -2375 199 -2374
rect 212 -2375 216 -2374
rect 219 -2375 437 -2374
rect 450 -2375 738 -2374
rect 968 -2375 983 -2374
rect 1160 -2375 1193 -2374
rect 1535 -2375 1571 -2374
rect 1584 -2375 1613 -2374
rect 156 -2377 1186 -2376
rect 1402 -2377 1585 -2376
rect 163 -2379 731 -2378
rect 737 -2379 780 -2378
rect 891 -2379 1186 -2378
rect 1374 -2379 1403 -2378
rect 1570 -2379 1753 -2378
rect 177 -2381 276 -2380
rect 366 -2381 430 -2380
rect 436 -2381 654 -2380
rect 681 -2381 696 -2380
rect 730 -2381 1501 -2380
rect 184 -2383 283 -2382
rect 366 -2383 381 -2382
rect 387 -2383 822 -2382
rect 891 -2383 920 -2382
rect 982 -2383 1032 -2382
rect 1346 -2383 1375 -2382
rect 184 -2385 360 -2384
rect 390 -2385 703 -2384
rect 828 -2385 1347 -2384
rect 191 -2387 241 -2386
rect 261 -2387 423 -2386
rect 485 -2387 549 -2386
rect 572 -2387 780 -2386
rect 828 -2387 1725 -2386
rect 23 -2389 192 -2388
rect 205 -2389 1753 -2388
rect 261 -2391 444 -2390
rect 520 -2391 850 -2390
rect 919 -2391 934 -2390
rect 1031 -2391 1046 -2390
rect 275 -2393 318 -2392
rect 338 -2393 360 -2392
rect 394 -2393 416 -2392
rect 527 -2393 1431 -2392
rect 289 -2395 444 -2394
rect 548 -2395 710 -2394
rect 800 -2395 850 -2394
rect 933 -2395 955 -2394
rect 1045 -2395 1305 -2394
rect 317 -2397 507 -2396
rect 569 -2397 710 -2396
rect 765 -2397 801 -2396
rect 835 -2397 955 -2396
rect 1262 -2397 1305 -2396
rect 268 -2399 507 -2398
rect 555 -2399 766 -2398
rect 835 -2399 1168 -2398
rect 268 -2401 332 -2400
rect 338 -2401 899 -2400
rect 1143 -2401 1263 -2400
rect 331 -2403 675 -2402
rect 695 -2403 1392 -2402
rect 254 -2405 675 -2404
rect 898 -2405 1714 -2404
rect 117 -2407 255 -2406
rect 341 -2407 381 -2406
rect 404 -2407 1529 -2406
rect 345 -2409 395 -2408
rect 569 -2409 612 -2408
rect 656 -2409 1144 -2408
rect 373 -2411 556 -2410
rect 576 -2411 1123 -2410
rect 373 -2413 797 -2412
rect 1108 -2413 1123 -2412
rect 597 -2415 612 -2414
rect 1073 -2415 1109 -2414
rect 345 -2417 598 -2416
rect 604 -2417 661 -2416
rect 1073 -2417 1368 -2416
rect 660 -2419 951 -2418
rect 1367 -2419 1473 -2418
rect 1311 -2421 1473 -2420
rect 1311 -2423 1354 -2422
rect 1297 -2425 1354 -2424
rect 1297 -2427 1410 -2426
rect 1381 -2429 1410 -2428
rect 1234 -2431 1382 -2430
rect 758 -2433 1235 -2432
rect 744 -2435 759 -2434
rect 744 -2437 752 -2436
rect 716 -2439 752 -2438
rect 9 -2450 598 -2449
rect 723 -2450 1018 -2449
rect 1020 -2450 1487 -2449
rect 1741 -2450 1774 -2449
rect 1808 -2450 1816 -2449
rect 16 -2452 24 -2451
rect 44 -2452 388 -2451
rect 408 -2452 720 -2451
rect 726 -2452 1718 -2451
rect 1752 -2452 1760 -2451
rect 1773 -2452 1795 -2451
rect 1801 -2452 1809 -2451
rect 16 -2454 678 -2453
rect 807 -2454 811 -2453
rect 828 -2454 853 -2453
rect 884 -2454 913 -2453
rect 950 -2454 1382 -2453
rect 1619 -2454 1718 -2453
rect 1759 -2454 1767 -2453
rect 44 -2456 150 -2455
rect 159 -2456 433 -2455
rect 439 -2456 1095 -2455
rect 1132 -2456 1522 -2455
rect 1570 -2456 1767 -2455
rect 51 -2458 545 -2457
rect 583 -2458 787 -2457
rect 807 -2458 955 -2457
rect 982 -2458 1119 -2457
rect 1150 -2458 1487 -2457
rect 1521 -2458 1543 -2457
rect 1619 -2458 1669 -2457
rect 51 -2460 577 -2459
rect 597 -2460 822 -2459
rect 828 -2460 864 -2459
rect 884 -2460 927 -2459
rect 940 -2460 955 -2459
rect 968 -2460 983 -2459
rect 1055 -2460 1249 -2459
rect 1325 -2460 1340 -2459
rect 1381 -2460 1396 -2459
rect 1542 -2460 1557 -2459
rect 1668 -2460 1711 -2459
rect 58 -2462 402 -2461
rect 408 -2462 713 -2461
rect 786 -2462 843 -2461
rect 887 -2462 1732 -2461
rect 58 -2464 262 -2463
rect 324 -2464 724 -2463
rect 821 -2464 1046 -2463
rect 1076 -2464 1697 -2463
rect 30 -2466 262 -2465
rect 275 -2466 325 -2465
rect 352 -2466 1396 -2465
rect 1556 -2466 1676 -2465
rect 1689 -2466 1711 -2465
rect 30 -2468 213 -2467
rect 226 -2468 402 -2467
rect 429 -2468 612 -2467
rect 842 -2468 1067 -2467
rect 1087 -2468 1095 -2467
rect 1150 -2468 1179 -2467
rect 1195 -2468 1634 -2467
rect 1640 -2468 1732 -2467
rect 65 -2470 391 -2469
rect 450 -2470 517 -2469
rect 530 -2470 570 -2469
rect 600 -2470 1179 -2469
rect 1325 -2470 1375 -2469
rect 1640 -2470 1655 -2469
rect 1675 -2470 1725 -2469
rect 65 -2472 318 -2471
rect 352 -2472 1168 -2471
rect 1332 -2472 1802 -2471
rect 72 -2474 388 -2473
rect 457 -2474 584 -2473
rect 600 -2474 696 -2473
rect 905 -2474 913 -2473
rect 940 -2474 1060 -2473
rect 1066 -2474 1130 -2473
rect 1160 -2474 1662 -2473
rect 1689 -2474 1739 -2473
rect 72 -2476 195 -2475
rect 198 -2476 213 -2475
rect 226 -2476 948 -2475
rect 971 -2476 1375 -2475
rect 1598 -2476 1725 -2475
rect 1738 -2476 1781 -2475
rect 82 -2478 234 -2477
rect 243 -2478 1011 -2477
rect 1048 -2478 1662 -2477
rect 1696 -2478 1788 -2477
rect 93 -2480 381 -2479
rect 443 -2480 1599 -2479
rect 1654 -2480 1683 -2479
rect 93 -2482 269 -2481
rect 275 -2482 395 -2481
rect 443 -2482 507 -2481
rect 513 -2482 591 -2481
rect 681 -2482 696 -2481
rect 740 -2482 948 -2481
rect 996 -2482 1011 -2481
rect 1087 -2482 1389 -2481
rect 96 -2484 346 -2483
rect 366 -2484 395 -2483
rect 457 -2484 850 -2483
rect 877 -2484 906 -2483
rect 989 -2484 997 -2483
rect 1129 -2484 1249 -2483
rect 1255 -2484 1683 -2483
rect 37 -2486 346 -2485
rect 366 -2486 619 -2485
rect 653 -2486 682 -2485
rect 810 -2486 1060 -2485
rect 1115 -2486 1256 -2485
rect 1321 -2486 1781 -2485
rect 37 -2488 115 -2487
rect 128 -2488 290 -2487
rect 317 -2488 461 -2487
rect 471 -2488 528 -2487
rect 541 -2488 661 -2487
rect 849 -2488 927 -2487
rect 989 -2488 1319 -2487
rect 1332 -2488 1494 -2487
rect 100 -2490 115 -2489
rect 128 -2490 283 -2489
rect 289 -2490 304 -2489
rect 415 -2490 472 -2489
rect 478 -2490 591 -2489
rect 604 -2490 661 -2489
rect 1115 -2490 1298 -2489
rect 1318 -2490 1361 -2489
rect 1367 -2490 1494 -2489
rect 100 -2492 1347 -2491
rect 1367 -2492 1466 -2491
rect 107 -2494 339 -2493
rect 478 -2494 738 -2493
rect 1003 -2494 1347 -2493
rect 1388 -2494 1403 -2493
rect 1465 -2494 1480 -2493
rect 107 -2496 1186 -2495
rect 1241 -2496 1788 -2495
rect 110 -2498 1018 -2497
rect 1101 -2498 1186 -2497
rect 1241 -2498 1291 -2497
rect 1402 -2498 1410 -2497
rect 1479 -2498 1508 -2497
rect 103 -2500 1102 -2499
rect 1157 -2500 1298 -2499
rect 1409 -2500 1417 -2499
rect 131 -2502 864 -2501
rect 1164 -2502 1312 -2501
rect 1416 -2502 1438 -2501
rect 135 -2504 437 -2503
rect 485 -2504 577 -2503
rect 604 -2504 1021 -2503
rect 1164 -2504 1200 -2503
rect 1269 -2504 1361 -2503
rect 1437 -2504 1452 -2503
rect 135 -2506 1046 -2505
rect 1080 -2506 1270 -2505
rect 1290 -2506 1515 -2505
rect 142 -2508 416 -2507
rect 436 -2508 1032 -2507
rect 1080 -2508 1137 -2507
rect 1311 -2508 1700 -2507
rect 121 -2510 143 -2509
rect 149 -2510 1634 -2509
rect 121 -2512 157 -2511
rect 163 -2512 381 -2511
rect 485 -2512 836 -2511
rect 1024 -2512 1032 -2511
rect 1122 -2512 1200 -2511
rect 1514 -2512 1529 -2511
rect 152 -2514 612 -2513
rect 639 -2514 654 -2513
rect 674 -2514 1452 -2513
rect 1528 -2514 1704 -2513
rect 163 -2516 1053 -2515
rect 1073 -2516 1704 -2515
rect 170 -2518 339 -2517
rect 492 -2518 832 -2517
rect 1108 -2518 1123 -2517
rect 170 -2520 1144 -2519
rect 173 -2522 311 -2521
rect 492 -2522 500 -2521
rect 506 -2522 689 -2521
rect 702 -2522 1025 -2521
rect 1108 -2522 1193 -2521
rect 191 -2524 878 -2523
rect 1143 -2524 1207 -2523
rect 191 -2526 871 -2525
rect 1192 -2526 1445 -2525
rect 198 -2528 559 -2527
rect 569 -2528 962 -2527
rect 1206 -2528 1221 -2527
rect 1444 -2528 1459 -2527
rect 219 -2530 619 -2529
rect 667 -2530 703 -2529
rect 737 -2530 1571 -2529
rect 219 -2532 465 -2531
rect 499 -2532 535 -2531
rect 674 -2532 710 -2531
rect 789 -2532 836 -2531
rect 870 -2532 934 -2531
rect 961 -2532 976 -2531
rect 1220 -2532 1277 -2531
rect 233 -2534 241 -2533
rect 247 -2534 451 -2533
rect 464 -2534 549 -2533
rect 688 -2534 752 -2533
rect 975 -2534 1172 -2533
rect 1276 -2534 1473 -2533
rect 247 -2536 1158 -2535
rect 1171 -2536 1536 -2535
rect 254 -2538 304 -2537
rect 310 -2538 629 -2537
rect 709 -2538 1004 -2537
rect 1472 -2538 1501 -2537
rect 1535 -2538 1550 -2537
rect 254 -2540 374 -2539
rect 513 -2540 556 -2539
rect 730 -2540 934 -2539
rect 1500 -2540 1564 -2539
rect 268 -2542 717 -2541
rect 730 -2542 1175 -2541
rect 1549 -2542 1578 -2541
rect 282 -2544 332 -2543
rect 359 -2544 374 -2543
rect 520 -2544 556 -2543
rect 716 -2544 759 -2543
rect 1563 -2544 1585 -2543
rect 177 -2546 332 -2545
rect 520 -2546 801 -2545
rect 1577 -2546 1592 -2545
rect 177 -2548 206 -2547
rect 527 -2548 563 -2547
rect 625 -2548 801 -2547
rect 1584 -2548 1606 -2547
rect 184 -2550 360 -2549
rect 534 -2550 745 -2549
rect 751 -2550 1214 -2549
rect 1591 -2550 1648 -2549
rect 184 -2552 342 -2551
rect 548 -2552 993 -2551
rect 1213 -2552 1228 -2551
rect 1283 -2552 1648 -2551
rect 205 -2554 423 -2553
rect 562 -2554 640 -2553
rect 744 -2554 766 -2553
rect 968 -2554 1228 -2553
rect 1262 -2554 1284 -2553
rect 1605 -2554 1613 -2553
rect 156 -2556 423 -2555
rect 625 -2556 1459 -2555
rect 1612 -2556 1627 -2555
rect 79 -2558 1627 -2557
rect 79 -2560 297 -2559
rect 758 -2560 773 -2559
rect 1262 -2560 1431 -2559
rect 296 -2562 405 -2561
rect 765 -2562 780 -2561
rect 1234 -2562 1431 -2561
rect 772 -2564 794 -2563
rect 1234 -2564 1305 -2563
rect 110 -2566 1305 -2565
rect 670 -2568 794 -2567
rect 779 -2570 899 -2569
rect 891 -2572 899 -2571
rect 453 -2574 892 -2573
rect 9 -2585 444 -2584
rect 450 -2585 1060 -2584
rect 1062 -2585 1277 -2584
rect 1293 -2585 1340 -2584
rect 1510 -2585 1592 -2584
rect 1738 -2585 1781 -2584
rect 44 -2587 629 -2586
rect 639 -2587 808 -2586
rect 852 -2587 997 -2586
rect 1020 -2587 1109 -2586
rect 1115 -2587 1312 -2586
rect 1339 -2587 1375 -2586
rect 1769 -2587 1784 -2586
rect 44 -2589 780 -2588
rect 807 -2589 829 -2588
rect 866 -2589 1508 -2588
rect 107 -2591 367 -2590
rect 443 -2591 584 -2590
rect 660 -2591 713 -2590
rect 726 -2591 1648 -2590
rect 79 -2593 108 -2592
rect 121 -2593 241 -2592
rect 243 -2593 283 -2592
rect 292 -2593 598 -2592
rect 660 -2593 871 -2592
rect 915 -2593 1354 -2592
rect 1507 -2593 1536 -2592
rect 1647 -2593 1655 -2592
rect 79 -2595 843 -2594
rect 947 -2595 1245 -2594
rect 1276 -2595 1305 -2594
rect 1311 -2595 1389 -2594
rect 1654 -2595 1777 -2594
rect 121 -2597 129 -2596
rect 149 -2597 388 -2596
rect 457 -2597 671 -2596
rect 695 -2597 713 -2596
rect 737 -2597 1487 -2596
rect 68 -2599 150 -2598
rect 156 -2599 255 -2598
rect 275 -2599 559 -2598
rect 642 -2599 1536 -2598
rect 86 -2601 129 -2600
rect 142 -2601 276 -2600
rect 282 -2601 290 -2600
rect 296 -2601 587 -2600
rect 681 -2601 738 -2600
rect 765 -2601 780 -2600
rect 842 -2601 885 -2600
rect 968 -2601 1431 -2600
rect 1486 -2601 1543 -2600
rect 86 -2603 101 -2602
rect 103 -2603 290 -2602
rect 296 -2603 1018 -2602
rect 1048 -2603 1291 -2602
rect 1304 -2603 1361 -2602
rect 1430 -2603 1445 -2602
rect 1542 -2603 1571 -2602
rect 37 -2605 101 -2604
rect 142 -2605 437 -2604
rect 453 -2605 682 -2604
rect 695 -2605 878 -2604
rect 905 -2605 969 -2604
rect 971 -2605 1704 -2604
rect 37 -2607 846 -2606
rect 856 -2607 878 -2606
rect 905 -2607 951 -2606
rect 989 -2607 1039 -2606
rect 1073 -2607 1095 -2606
rect 1108 -2607 1144 -2606
rect 1157 -2607 1221 -2606
rect 1262 -2607 1389 -2606
rect 1444 -2607 1459 -2606
rect 1570 -2607 1599 -2606
rect 1675 -2607 1704 -2606
rect 156 -2609 199 -2608
rect 205 -2609 451 -2608
rect 492 -2609 766 -2608
rect 775 -2609 1375 -2608
rect 1458 -2609 1515 -2608
rect 1598 -2609 1620 -2608
rect 1675 -2609 1718 -2608
rect 159 -2611 927 -2610
rect 940 -2611 1144 -2610
rect 1174 -2611 1333 -2610
rect 1353 -2611 1410 -2610
rect 1514 -2611 1700 -2610
rect 1710 -2611 1718 -2610
rect 170 -2613 1249 -2612
rect 1409 -2613 1606 -2612
rect 1689 -2613 1711 -2612
rect 170 -2615 605 -2614
rect 702 -2615 741 -2614
rect 856 -2615 1053 -2614
rect 1066 -2615 1333 -2614
rect 1556 -2615 1606 -2614
rect 1689 -2615 1767 -2614
rect 173 -2617 1102 -2616
rect 1118 -2617 1592 -2616
rect 177 -2619 255 -2618
rect 303 -2619 458 -2618
rect 492 -2619 731 -2618
rect 828 -2619 1767 -2618
rect 23 -2621 178 -2620
rect 184 -2621 668 -2620
rect 702 -2621 787 -2620
rect 870 -2621 1053 -2620
rect 1076 -2621 1186 -2620
rect 1220 -2621 1319 -2620
rect 1556 -2621 1585 -2620
rect 184 -2623 199 -2622
rect 205 -2623 346 -2622
rect 387 -2623 689 -2622
rect 709 -2623 1207 -2622
rect 1241 -2623 1263 -2622
rect 1584 -2623 1613 -2622
rect 226 -2625 1021 -2624
rect 1024 -2625 1039 -2624
rect 1094 -2625 1151 -2624
rect 1241 -2625 1368 -2624
rect 1612 -2625 1627 -2624
rect 30 -2627 227 -2626
rect 303 -2627 486 -2626
rect 513 -2627 605 -2626
rect 646 -2627 668 -2626
rect 723 -2627 1361 -2626
rect 1367 -2627 1494 -2626
rect 1626 -2627 1634 -2626
rect 30 -2629 66 -2628
rect 310 -2629 426 -2628
rect 436 -2629 717 -2628
rect 730 -2629 745 -2628
rect 786 -2629 1172 -2628
rect 1248 -2629 1322 -2628
rect 1479 -2629 1494 -2628
rect 1633 -2629 1732 -2628
rect 58 -2631 514 -2630
rect 520 -2631 853 -2630
rect 912 -2631 927 -2630
rect 933 -2631 1207 -2630
rect 1731 -2631 1746 -2630
rect 58 -2633 801 -2632
rect 835 -2633 934 -2632
rect 940 -2633 1396 -2632
rect 1745 -2633 1753 -2632
rect 110 -2635 311 -2634
rect 338 -2635 367 -2634
rect 380 -2635 689 -2634
rect 716 -2635 1319 -2634
rect 1395 -2635 1417 -2634
rect 1752 -2635 1760 -2634
rect 135 -2637 836 -2636
rect 919 -2637 1186 -2636
rect 1416 -2637 1473 -2636
rect 1759 -2637 1774 -2636
rect 135 -2639 234 -2638
rect 338 -2639 402 -2638
rect 408 -2639 990 -2638
rect 996 -2639 1011 -2638
rect 1017 -2639 1683 -2638
rect 72 -2641 234 -2640
rect 345 -2641 353 -2640
rect 359 -2641 381 -2640
rect 394 -2641 402 -2640
rect 422 -2641 486 -2640
rect 520 -2641 1662 -2640
rect 72 -2643 465 -2642
rect 523 -2643 570 -2642
rect 646 -2643 654 -2642
rect 674 -2643 724 -2642
rect 800 -2643 979 -2642
rect 1003 -2643 1067 -2642
rect 1101 -2643 1165 -2642
rect 1171 -2643 1298 -2642
rect 1472 -2643 1522 -2642
rect 152 -2645 1662 -2644
rect 201 -2647 1480 -2646
rect 1521 -2647 1550 -2646
rect 268 -2649 675 -2648
rect 891 -2649 1011 -2648
rect 1024 -2649 1081 -2648
rect 1122 -2649 1137 -2648
rect 1139 -2649 1739 -2648
rect 268 -2651 1161 -2650
rect 1297 -2651 1326 -2650
rect 1549 -2651 1578 -2650
rect 324 -2653 353 -2652
rect 359 -2653 430 -2652
rect 464 -2653 794 -2652
rect 821 -2653 1137 -2652
rect 1325 -2653 1620 -2652
rect 324 -2655 549 -2654
rect 569 -2655 591 -2654
rect 625 -2655 892 -2654
rect 912 -2655 1081 -2654
rect 1122 -2655 1179 -2654
rect 1577 -2655 1742 -2654
rect 163 -2657 549 -2656
rect 590 -2657 619 -2656
rect 625 -2657 850 -2656
rect 954 -2657 1004 -2656
rect 1087 -2657 1179 -2656
rect 163 -2659 220 -2658
rect 373 -2659 409 -2658
rect 415 -2659 430 -2658
rect 506 -2659 619 -2658
rect 632 -2659 654 -2658
rect 772 -2659 794 -2658
rect 814 -2659 822 -2658
rect 849 -2659 1683 -2658
rect 219 -2661 248 -2660
rect 331 -2661 374 -2660
rect 394 -2661 752 -2660
rect 814 -2661 1200 -2660
rect 93 -2663 332 -2662
rect 415 -2663 1196 -2662
rect 1199 -2663 1214 -2662
rect 93 -2665 115 -2664
rect 191 -2665 248 -2664
rect 478 -2665 773 -2664
rect 863 -2665 955 -2664
rect 961 -2665 1165 -2664
rect 1195 -2665 1501 -2664
rect 114 -2667 209 -2666
rect 471 -2667 479 -2666
rect 506 -2667 563 -2666
rect 597 -2667 633 -2666
rect 635 -2667 752 -2666
rect 961 -2667 983 -2666
rect 1045 -2667 1088 -2666
rect 1132 -2667 1669 -2666
rect 191 -2669 213 -2668
rect 471 -2669 1151 -2668
rect 1213 -2669 1802 -2668
rect 51 -2671 213 -2670
rect 499 -2671 563 -2670
rect 975 -2671 983 -2670
rect 1045 -2671 1347 -2670
rect 1500 -2671 1788 -2670
rect 1801 -2671 1809 -2670
rect 51 -2673 423 -2672
rect 499 -2673 584 -2672
rect 975 -2673 1032 -2672
rect 1346 -2673 1382 -2672
rect 1528 -2673 1669 -2672
rect 1787 -2673 1795 -2672
rect 1808 -2673 1816 -2672
rect 527 -2675 531 -2674
rect 534 -2675 745 -2674
rect 1381 -2675 1403 -2674
rect 1696 -2675 1795 -2674
rect 527 -2677 542 -2676
rect 555 -2677 1697 -2676
rect 530 -2679 542 -2678
rect 555 -2679 577 -2678
rect 611 -2679 1032 -2678
rect 1192 -2679 1403 -2678
rect 534 -2681 1056 -2680
rect 576 -2683 1774 -2682
rect 611 -2685 1130 -2684
rect 709 -2687 1529 -2686
rect 1055 -2689 1641 -2688
rect 1059 -2691 1130 -2690
rect 1269 -2691 1641 -2690
rect 1234 -2693 1270 -2692
rect 1227 -2695 1235 -2694
rect 1227 -2697 1284 -2696
rect 1255 -2699 1284 -2698
rect 1255 -2701 1452 -2700
rect 1423 -2703 1452 -2702
rect 1423 -2705 1438 -2704
rect 1192 -2707 1438 -2706
rect 30 -2718 713 -2717
rect 737 -2718 773 -2717
rect 842 -2718 1494 -2717
rect 1769 -2718 1809 -2717
rect 44 -2720 69 -2719
rect 72 -2720 643 -2719
rect 712 -2720 1196 -2719
rect 1290 -2720 1361 -2719
rect 1433 -2720 1452 -2719
rect 1493 -2720 1508 -2719
rect 1780 -2720 1802 -2719
rect 58 -2722 73 -2721
rect 96 -2722 143 -2721
rect 198 -2722 1777 -2721
rect 1783 -2722 1788 -2721
rect 58 -2724 591 -2723
rect 621 -2724 738 -2723
rect 775 -2724 1508 -2723
rect 65 -2726 1126 -2725
rect 1129 -2726 1203 -2725
rect 1297 -2726 1361 -2725
rect 100 -2728 104 -2727
rect 107 -2728 524 -2727
rect 534 -2728 888 -2727
rect 891 -2728 979 -2727
rect 1003 -2728 1326 -2727
rect 1328 -2728 1676 -2727
rect 100 -2730 157 -2729
rect 198 -2730 209 -2729
rect 289 -2730 374 -2729
rect 401 -2730 423 -2729
rect 425 -2730 605 -2729
rect 660 -2730 892 -2729
rect 919 -2730 1235 -2729
rect 1297 -2730 1340 -2729
rect 1346 -2730 1452 -2729
rect 1675 -2730 1718 -2729
rect 107 -2732 444 -2731
rect 464 -2732 1182 -2731
rect 1318 -2732 1606 -2731
rect 142 -2734 668 -2733
rect 842 -2734 857 -2733
rect 863 -2734 1207 -2733
rect 1318 -2734 1438 -2733
rect 1605 -2734 1627 -2733
rect 149 -2736 157 -2735
rect 201 -2736 262 -2735
rect 292 -2736 514 -2735
rect 534 -2736 745 -2735
rect 849 -2736 1284 -2735
rect 1325 -2736 1424 -2735
rect 1437 -2736 1550 -2735
rect 1626 -2736 1648 -2735
rect 103 -2738 150 -2737
rect 205 -2738 220 -2737
rect 226 -2738 374 -2737
rect 436 -2738 633 -2737
rect 660 -2738 664 -2737
rect 667 -2738 955 -2737
rect 1003 -2738 1070 -2737
rect 1080 -2738 1242 -2737
rect 1332 -2738 1774 -2737
rect 128 -2740 220 -2739
rect 226 -2740 612 -2739
rect 632 -2740 654 -2739
rect 705 -2740 1333 -2739
rect 1346 -2740 1354 -2739
rect 1549 -2740 1585 -2739
rect 1647 -2740 1683 -2739
rect 1773 -2740 1795 -2739
rect 79 -2742 129 -2741
rect 170 -2742 654 -2741
rect 716 -2742 857 -2741
rect 863 -2742 1214 -2741
rect 1241 -2742 1389 -2741
rect 1584 -2742 1613 -2741
rect 1682 -2742 1725 -2741
rect 61 -2744 1214 -2743
rect 1237 -2744 1613 -2743
rect 79 -2746 94 -2745
rect 170 -2746 360 -2745
rect 436 -2746 640 -2745
rect 716 -2746 780 -2745
rect 852 -2746 878 -2745
rect 884 -2746 1165 -2745
rect 1283 -2746 1725 -2745
rect 37 -2748 360 -2747
rect 443 -2748 542 -2747
rect 562 -2748 640 -2747
rect 695 -2748 780 -2747
rect 877 -2748 1322 -2747
rect 1388 -2748 1431 -2747
rect 37 -2750 87 -2749
rect 261 -2750 1354 -2749
rect 9 -2752 87 -2751
rect 303 -2752 860 -2751
rect 884 -2752 1063 -2751
rect 1080 -2752 1095 -2751
rect 1118 -2752 1662 -2751
rect 44 -2754 94 -2753
rect 303 -2754 367 -2753
rect 464 -2754 787 -2753
rect 919 -2754 990 -2753
rect 1010 -2754 1053 -2753
rect 1087 -2754 1343 -2753
rect 1661 -2754 1753 -2753
rect 268 -2756 367 -2755
rect 478 -2756 482 -2755
rect 513 -2756 528 -2755
rect 541 -2756 598 -2755
rect 611 -2756 724 -2755
rect 744 -2756 794 -2755
rect 940 -2756 1207 -2755
rect 1720 -2756 1753 -2755
rect 135 -2758 269 -2757
rect 331 -2758 566 -2757
rect 569 -2758 916 -2757
rect 940 -2758 1154 -2757
rect 1164 -2758 1200 -2757
rect 135 -2760 234 -2759
rect 310 -2760 332 -2759
rect 338 -2760 402 -2759
rect 527 -2760 829 -2759
rect 954 -2760 962 -2759
rect 982 -2760 990 -2759
rect 1013 -2760 1424 -2759
rect 51 -2762 234 -2761
rect 310 -2762 1011 -2761
rect 1017 -2762 1760 -2761
rect 51 -2764 388 -2763
rect 562 -2764 703 -2763
rect 786 -2764 1046 -2763
rect 1052 -2764 1074 -2763
rect 1094 -2764 1571 -2763
rect 1745 -2764 1760 -2763
rect 324 -2766 703 -2765
rect 866 -2766 1571 -2765
rect 324 -2768 353 -2767
rect 355 -2768 836 -2767
rect 961 -2768 1144 -2767
rect 1150 -2768 1690 -2767
rect 338 -2770 458 -2769
rect 569 -2770 626 -2769
rect 695 -2770 731 -2769
rect 821 -2770 836 -2769
rect 982 -2770 1179 -2769
rect 1199 -2770 1515 -2769
rect 1633 -2770 1690 -2769
rect 345 -2772 423 -2771
rect 457 -2772 832 -2771
rect 1031 -2772 1046 -2771
rect 1073 -2772 1277 -2771
rect 1430 -2772 1746 -2771
rect 345 -2774 1060 -2773
rect 1143 -2774 1249 -2773
rect 1276 -2774 1312 -2773
rect 1514 -2774 1543 -2773
rect 1633 -2774 1655 -2773
rect 380 -2776 388 -2775
rect 499 -2776 626 -2775
rect 751 -2776 1249 -2775
rect 1311 -2776 1459 -2775
rect 1542 -2776 1557 -2775
rect 380 -2778 409 -2777
rect 478 -2778 500 -2777
rect 583 -2778 1375 -2777
rect 1458 -2778 1473 -2777
rect 1556 -2778 1697 -2777
rect 408 -2780 507 -2779
rect 583 -2780 724 -2779
rect 807 -2780 822 -2779
rect 996 -2780 1060 -2779
rect 1129 -2780 1655 -2779
rect 1696 -2780 1732 -2779
rect 415 -2782 507 -2781
rect 520 -2782 808 -2781
rect 1031 -2782 1480 -2781
rect 1500 -2782 1732 -2781
rect 415 -2784 430 -2783
rect 520 -2784 577 -2783
rect 590 -2784 1718 -2783
rect 247 -2786 577 -2785
rect 597 -2786 689 -2785
rect 1150 -2786 1172 -2785
rect 1178 -2786 1564 -2785
rect 247 -2788 472 -2787
rect 548 -2788 997 -2787
rect 1171 -2788 1228 -2787
rect 1374 -2788 1767 -2787
rect 177 -2790 549 -2789
rect 607 -2790 794 -2789
rect 947 -2790 1228 -2789
rect 1402 -2790 1767 -2789
rect 121 -2792 178 -2791
rect 296 -2792 689 -2791
rect 1402 -2792 1592 -2791
rect 121 -2794 241 -2793
rect 296 -2794 682 -2793
rect 1465 -2794 1564 -2793
rect 1591 -2794 1620 -2793
rect 212 -2796 241 -2795
rect 317 -2796 430 -2795
rect 471 -2796 486 -2795
rect 618 -2796 731 -2795
rect 1465 -2796 1487 -2795
rect 1619 -2796 1704 -2795
rect 212 -2798 283 -2797
rect 317 -2798 1186 -2797
rect 1472 -2798 1522 -2797
rect 1703 -2798 1739 -2797
rect 254 -2800 283 -2799
rect 485 -2800 556 -2799
rect 618 -2800 752 -2799
rect 912 -2800 1522 -2799
rect 163 -2802 556 -2801
rect 635 -2802 948 -2801
rect 975 -2802 1487 -2801
rect 163 -2804 192 -2803
rect 254 -2804 871 -2803
rect 912 -2804 927 -2803
rect 975 -2804 1039 -2803
rect 1185 -2804 1263 -2803
rect 1381 -2804 1739 -2803
rect 191 -2806 493 -2805
rect 681 -2806 766 -2805
rect 926 -2806 969 -2805
rect 1038 -2806 1116 -2805
rect 1255 -2806 1263 -2805
rect 1381 -2806 1445 -2805
rect 1479 -2806 1529 -2805
rect 450 -2808 493 -2807
rect 709 -2808 766 -2807
rect 968 -2808 1025 -2807
rect 1087 -2808 1116 -2807
rect 1255 -2808 1305 -2807
rect 1444 -2808 1641 -2807
rect 394 -2810 451 -2809
rect 709 -2810 846 -2809
rect 1024 -2810 1067 -2809
rect 1304 -2810 1368 -2809
rect 1528 -2810 1578 -2809
rect 1640 -2810 1669 -2809
rect 394 -2812 675 -2811
rect 1066 -2812 1221 -2811
rect 1367 -2812 1396 -2811
rect 1577 -2812 1599 -2811
rect 1668 -2812 1711 -2811
rect 674 -2814 759 -2813
rect 1020 -2814 1396 -2813
rect 1500 -2814 1711 -2813
rect 758 -2816 801 -2815
rect 1020 -2816 1193 -2815
rect 1220 -2816 1270 -2815
rect 1535 -2816 1599 -2815
rect 800 -2818 934 -2817
rect 1136 -2818 1270 -2817
rect 1409 -2818 1536 -2817
rect 814 -2820 934 -2819
rect 1136 -2820 1245 -2819
rect 1409 -2820 1417 -2819
rect 814 -2822 1714 -2821
rect 905 -2824 1417 -2823
rect 898 -2826 906 -2825
rect 1157 -2826 1193 -2825
rect 733 -2828 899 -2827
rect 1122 -2828 1158 -2827
rect 23 -2839 290 -2838
rect 331 -2839 584 -2838
rect 621 -2839 1032 -2838
rect 1097 -2839 1669 -2838
rect 1713 -2839 1760 -2838
rect 44 -2841 559 -2840
rect 656 -2841 1417 -2840
rect 1433 -2841 1690 -2840
rect 1717 -2841 1774 -2840
rect 79 -2843 584 -2842
rect 660 -2843 1249 -2842
rect 1283 -2843 1676 -2842
rect 1720 -2843 1767 -2842
rect 93 -2845 1249 -2844
rect 1339 -2845 1613 -2844
rect 1654 -2845 1676 -2844
rect 1727 -2845 1753 -2844
rect 93 -2847 122 -2846
rect 128 -2847 829 -2846
rect 859 -2847 1697 -2846
rect 96 -2849 706 -2848
rect 712 -2849 787 -2848
rect 824 -2849 1508 -2848
rect 1598 -2849 1697 -2848
rect 100 -2851 619 -2850
rect 681 -2851 997 -2850
rect 1013 -2851 1389 -2850
rect 1465 -2851 1508 -2850
rect 1591 -2851 1599 -2850
rect 1647 -2851 1655 -2850
rect 37 -2853 682 -2852
rect 730 -2853 878 -2852
rect 915 -2853 1333 -2852
rect 1342 -2853 1564 -2852
rect 1640 -2853 1648 -2852
rect 51 -2855 101 -2854
rect 107 -2855 857 -2854
rect 870 -2855 906 -2854
rect 947 -2855 1018 -2854
rect 1024 -2855 1130 -2854
rect 1150 -2855 1284 -2854
rect 1353 -2855 1683 -2854
rect 51 -2857 73 -2856
rect 107 -2857 1158 -2856
rect 1178 -2857 1704 -2856
rect 72 -2859 325 -2858
rect 359 -2859 710 -2858
rect 765 -2859 857 -2858
rect 877 -2859 1011 -2858
rect 1024 -2859 1515 -2858
rect 1661 -2859 1683 -2858
rect 1703 -2859 1725 -2858
rect 121 -2861 192 -2860
rect 226 -2861 353 -2860
rect 366 -2861 482 -2860
rect 520 -2861 1056 -2860
rect 1101 -2861 1151 -2860
rect 1199 -2861 1277 -2860
rect 1353 -2861 1375 -2860
rect 1381 -2861 1417 -2860
rect 1444 -2861 1592 -2860
rect 1640 -2861 1662 -2860
rect 65 -2863 521 -2862
rect 555 -2863 1046 -2862
rect 1066 -2863 1102 -2862
rect 1115 -2863 1165 -2862
rect 1202 -2863 1452 -2862
rect 1514 -2863 1529 -2862
rect 65 -2865 262 -2864
rect 275 -2865 356 -2864
rect 366 -2865 381 -2864
rect 429 -2865 433 -2864
rect 464 -2865 1179 -2864
rect 1227 -2865 1690 -2864
rect 128 -2867 230 -2866
rect 247 -2867 1000 -2866
rect 1066 -2867 1235 -2866
rect 1237 -2867 1501 -2866
rect 135 -2869 412 -2868
rect 429 -2869 542 -2868
rect 555 -2869 647 -2868
rect 674 -2869 1116 -2868
rect 1125 -2869 1543 -2868
rect 142 -2871 703 -2870
rect 737 -2871 766 -2870
rect 779 -2871 948 -2870
rect 968 -2871 1046 -2870
rect 1136 -2871 1277 -2870
rect 1311 -2871 1452 -2870
rect 1500 -2871 1522 -2870
rect 1535 -2871 1543 -2870
rect 86 -2873 143 -2872
rect 145 -2873 1613 -2872
rect 86 -2875 115 -2874
rect 170 -2875 587 -2874
rect 604 -2875 1130 -2874
rect 1164 -2875 1172 -2874
rect 1227 -2875 1732 -2874
rect 58 -2877 115 -2876
rect 156 -2877 171 -2876
rect 226 -2877 468 -2876
rect 562 -2877 1564 -2876
rect 58 -2879 783 -2878
rect 786 -2879 1028 -2878
rect 1171 -2879 1396 -2878
rect 1437 -2879 1529 -2878
rect 156 -2881 185 -2880
rect 240 -2881 248 -2880
rect 254 -2881 867 -2880
rect 971 -2881 1298 -2880
rect 1311 -2881 1711 -2880
rect 149 -2883 255 -2882
rect 261 -2883 374 -2882
rect 380 -2883 566 -2882
rect 576 -2883 619 -2882
rect 646 -2883 808 -2882
rect 821 -2883 871 -2882
rect 982 -2883 1137 -2882
rect 1234 -2883 1305 -2882
rect 1318 -2883 1396 -2882
rect 1423 -2883 1438 -2882
rect 1444 -2883 1578 -2882
rect 149 -2885 339 -2884
rect 373 -2885 388 -2884
rect 394 -2885 465 -2884
rect 562 -2885 570 -2884
rect 576 -2885 850 -2884
rect 898 -2885 983 -2884
rect 989 -2885 1011 -2884
rect 1255 -2885 1298 -2884
rect 1318 -2885 1739 -2884
rect 184 -2887 626 -2886
rect 667 -2887 899 -2886
rect 933 -2887 1424 -2886
rect 1479 -2887 1522 -2886
rect 1570 -2887 1578 -2886
rect 233 -2889 388 -2888
rect 394 -2889 423 -2888
rect 432 -2889 542 -2888
rect 590 -2889 605 -2888
rect 625 -2889 874 -2888
rect 1143 -2889 1256 -2888
rect 1262 -2889 1389 -2888
rect 1458 -2889 1480 -2888
rect 1486 -2889 1536 -2888
rect 1570 -2889 1585 -2888
rect 233 -2891 1123 -2890
rect 1185 -2891 1263 -2890
rect 1269 -2891 1305 -2890
rect 1325 -2891 1382 -2890
rect 1409 -2891 1585 -2890
rect 240 -2893 269 -2892
rect 275 -2893 815 -2892
rect 828 -2893 836 -2892
rect 849 -2893 1361 -2892
rect 1367 -2893 1375 -2892
rect 1472 -2893 1487 -2892
rect 268 -2895 640 -2894
rect 653 -2895 1144 -2894
rect 1185 -2895 1193 -2894
rect 1213 -2895 1361 -2894
rect 1472 -2895 1494 -2894
rect 282 -2897 360 -2896
rect 415 -2897 423 -2896
rect 439 -2897 1410 -2896
rect 198 -2899 416 -2898
rect 527 -2899 570 -2898
rect 590 -2899 717 -2898
rect 737 -2899 941 -2898
rect 1059 -2899 1193 -2898
rect 1220 -2899 1270 -2898
rect 1325 -2899 1347 -2898
rect 1356 -2899 1620 -2898
rect 110 -2901 717 -2900
rect 751 -2901 934 -2900
rect 1052 -2901 1060 -2900
rect 1069 -2901 1459 -2900
rect 198 -2903 206 -2902
rect 212 -2903 283 -2902
rect 289 -2903 311 -2902
rect 317 -2903 990 -2902
rect 1052 -2903 1557 -2902
rect 163 -2905 206 -2904
rect 212 -2905 1287 -2904
rect 1290 -2905 1347 -2904
rect 1402 -2905 1557 -2904
rect 163 -2907 1158 -2906
rect 1206 -2907 1620 -2906
rect 303 -2909 318 -2908
rect 324 -2909 402 -2908
rect 506 -2909 528 -2908
rect 653 -2909 1669 -2908
rect 208 -2911 304 -2910
rect 310 -2911 458 -2910
rect 506 -2911 598 -2910
rect 663 -2911 815 -2910
rect 835 -2911 1088 -2910
rect 1094 -2911 1494 -2910
rect 219 -2913 458 -2912
rect 667 -2913 1032 -2912
rect 1073 -2913 1291 -2912
rect 1402 -2913 1746 -2912
rect 219 -2915 969 -2914
rect 1038 -2915 1074 -2914
rect 1080 -2915 1123 -2914
rect 1241 -2915 1368 -2914
rect 338 -2917 409 -2916
rect 436 -2917 598 -2916
rect 674 -2917 853 -2916
rect 891 -2917 1214 -2916
rect 191 -2919 437 -2918
rect 688 -2919 752 -2918
rect 800 -2919 906 -2918
rect 961 -2919 1207 -2918
rect 331 -2921 853 -2920
rect 926 -2921 962 -2920
rect 975 -2921 1039 -2920
rect 1108 -2921 1221 -2920
rect 345 -2923 640 -2922
rect 688 -2923 1021 -2922
rect 1108 -2923 1431 -2922
rect 177 -2925 346 -2924
rect 401 -2925 451 -2924
rect 695 -2925 801 -2924
rect 807 -2925 885 -2924
rect 919 -2925 976 -2924
rect 1003 -2925 1081 -2924
rect 1430 -2925 1606 -2924
rect 177 -2927 486 -2926
rect 534 -2927 696 -2926
rect 723 -2927 1088 -2926
rect 1605 -2927 1627 -2926
rect 443 -2929 451 -2928
rect 485 -2929 538 -2928
rect 723 -2929 759 -2928
rect 793 -2929 920 -2928
rect 926 -2929 1203 -2928
rect 1626 -2929 1634 -2928
rect 443 -2931 514 -2930
rect 733 -2931 1634 -2930
rect 478 -2933 514 -2932
rect 744 -2933 794 -2932
rect 842 -2933 892 -2932
rect 478 -2935 944 -2934
rect 492 -2937 535 -2936
rect 611 -2937 745 -2936
rect 758 -2937 773 -2936
rect 863 -2937 1004 -2936
rect 492 -2939 661 -2938
rect 663 -2939 843 -2938
rect 863 -2939 1242 -2938
rect 548 -2941 773 -2940
rect 884 -2941 913 -2940
rect 82 -2943 549 -2942
rect 611 -2943 633 -2942
rect 912 -2943 1466 -2942
rect 296 -2945 633 -2944
rect 166 -2947 297 -2946
rect 30 -2958 94 -2957
rect 100 -2958 437 -2957
rect 439 -2958 815 -2957
rect 821 -2958 857 -2957
rect 863 -2958 1585 -2957
rect 1640 -2958 1697 -2957
rect 37 -2960 290 -2959
rect 303 -2960 307 -2959
rect 369 -2960 454 -2959
rect 541 -2960 654 -2959
rect 663 -2960 1214 -2959
rect 1332 -2960 1508 -2959
rect 1577 -2960 1704 -2959
rect 44 -2962 395 -2961
rect 450 -2962 542 -2961
rect 548 -2962 815 -2961
rect 842 -2962 1025 -2961
rect 1027 -2962 1690 -2961
rect 23 -2964 451 -2963
rect 499 -2964 549 -2963
rect 611 -2964 654 -2963
rect 674 -2964 979 -2963
rect 1020 -2964 1221 -2963
rect 1332 -2964 1382 -2963
rect 1458 -2964 1641 -2963
rect 72 -2966 412 -2965
rect 499 -2966 689 -2965
rect 740 -2966 1144 -2965
rect 1171 -2966 1382 -2965
rect 1458 -2966 1466 -2965
rect 1577 -2966 1606 -2965
rect 51 -2968 73 -2967
rect 79 -2968 458 -2967
rect 569 -2968 612 -2967
rect 618 -2968 843 -2967
rect 849 -2968 1116 -2967
rect 1150 -2968 1172 -2967
rect 1199 -2968 1529 -2967
rect 1605 -2968 1648 -2967
rect 51 -2970 213 -2969
rect 219 -2970 997 -2969
rect 1010 -2970 1144 -2969
rect 1199 -2970 1242 -2969
rect 1339 -2970 1585 -2969
rect 1647 -2970 1683 -2969
rect 65 -2972 220 -2971
rect 261 -2972 395 -2971
rect 408 -2972 458 -2971
rect 492 -2972 570 -2971
rect 604 -2972 619 -2971
rect 674 -2972 794 -2971
rect 835 -2972 1151 -2971
rect 1164 -2972 1242 -2971
rect 1339 -2972 1389 -2971
rect 1465 -2972 1487 -2971
rect 65 -2974 209 -2973
rect 261 -2974 514 -2973
rect 604 -2974 759 -2973
rect 782 -2974 1536 -2973
rect 82 -2976 1179 -2975
rect 1213 -2976 1256 -2975
rect 1297 -2976 1389 -2975
rect 1486 -2976 1494 -2975
rect 1535 -2976 1564 -2975
rect 93 -2978 563 -2977
rect 793 -2978 927 -2977
rect 943 -2978 1417 -2977
rect 1430 -2978 1564 -2977
rect 79 -2980 1417 -2979
rect 1430 -2980 1669 -2979
rect 100 -2982 661 -2981
rect 835 -2982 990 -2981
rect 996 -2982 1039 -2981
rect 1052 -2982 1060 -2981
rect 1094 -2982 1319 -2981
rect 1493 -2982 1515 -2981
rect 107 -2984 1025 -2983
rect 1031 -2984 1592 -2983
rect 107 -2986 444 -2985
rect 562 -2986 867 -2985
rect 901 -2986 1424 -2985
rect 1514 -2986 1550 -2985
rect 1591 -2986 1634 -2985
rect 110 -2988 255 -2987
rect 268 -2988 1098 -2987
rect 1115 -2988 1130 -2987
rect 1136 -2988 1179 -2987
rect 1202 -2988 1634 -2987
rect 121 -2990 622 -2989
rect 660 -2990 731 -2989
rect 849 -2990 885 -2989
rect 926 -2990 948 -2989
rect 982 -2990 1039 -2989
rect 1045 -2990 1130 -2989
rect 1136 -2990 1361 -2989
rect 1423 -2990 1676 -2989
rect 82 -2992 1046 -2991
rect 1055 -2992 1522 -2991
rect 1549 -2992 1571 -2991
rect 121 -2994 360 -2993
rect 408 -2994 416 -2993
rect 443 -2994 668 -2993
rect 852 -2994 920 -2993
rect 947 -2994 955 -2993
rect 989 -2994 1074 -2993
rect 1122 -2994 1165 -2993
rect 1220 -2994 1263 -2993
rect 1297 -2994 1354 -2993
rect 1521 -2994 1557 -2993
rect 1570 -2994 1599 -2993
rect 89 -2996 1123 -2995
rect 1255 -2996 1291 -2995
rect 1318 -2996 1368 -2995
rect 1598 -2996 1627 -2995
rect 142 -2998 983 -2997
rect 1010 -2998 1228 -2997
rect 1262 -2998 1312 -2997
rect 1367 -2998 1396 -2997
rect 1626 -2998 1662 -2997
rect 145 -3000 584 -2999
rect 632 -3000 731 -2999
rect 856 -3000 871 -2999
rect 877 -3000 920 -2999
rect 954 -3000 962 -2999
rect 968 -3000 1074 -2999
rect 1227 -3000 1347 -2999
rect 156 -3002 255 -3001
rect 268 -3002 381 -3001
rect 415 -3002 423 -3001
rect 506 -3002 1361 -3001
rect 156 -3004 787 -3003
rect 880 -3004 1354 -3003
rect 163 -3006 934 -3005
rect 961 -3006 1336 -3005
rect 1346 -3006 1707 -3005
rect 86 -3008 164 -3007
rect 170 -3008 227 -3007
rect 282 -3008 381 -3007
rect 401 -3008 507 -3007
rect 583 -3008 941 -3007
rect 968 -3008 976 -3007
rect 1017 -3008 1032 -3007
rect 1034 -3008 1613 -3007
rect 86 -3010 1620 -3009
rect 128 -3012 227 -3011
rect 275 -3012 283 -3011
rect 289 -3012 577 -3011
rect 632 -3012 864 -3011
rect 884 -3012 1109 -3011
rect 1234 -3012 1312 -3011
rect 1612 -3012 1655 -3011
rect 58 -3014 577 -3013
rect 639 -3014 668 -3013
rect 702 -3014 878 -3013
rect 898 -3014 934 -3013
rect 1059 -3014 1088 -3013
rect 1108 -3014 1207 -3013
rect 1234 -3014 1277 -3013
rect 58 -3016 136 -3015
rect 138 -3016 276 -3015
rect 303 -3016 479 -3015
rect 513 -3016 1018 -3015
rect 1192 -3016 1655 -3015
rect 128 -3018 696 -3017
rect 702 -3018 724 -3017
rect 789 -3018 941 -3017
rect 1185 -3018 1193 -3017
rect 1206 -3018 1249 -3017
rect 170 -3020 192 -3019
rect 205 -3020 297 -3019
rect 317 -3020 423 -3019
rect 478 -3020 556 -3019
rect 639 -3020 647 -3019
rect 656 -3020 1291 -3019
rect 61 -3022 297 -3021
rect 306 -3022 556 -3021
rect 646 -3022 1102 -3021
rect 1248 -3022 1284 -3021
rect 177 -3024 692 -3023
rect 709 -3024 871 -3023
rect 898 -3024 1067 -3023
rect 1283 -3024 1326 -3023
rect 177 -3026 374 -3025
rect 401 -3026 430 -3025
rect 681 -3026 1277 -3025
rect 1325 -3026 1375 -3025
rect 114 -3028 430 -3027
rect 464 -3028 682 -3027
rect 688 -3028 1102 -3027
rect 1374 -3028 1403 -3027
rect 149 -3030 465 -3029
rect 709 -3030 752 -3029
rect 912 -3030 1557 -3029
rect 149 -3032 1158 -3031
rect 1304 -3032 1403 -3031
rect 187 -3034 1529 -3033
rect 191 -3036 199 -3035
rect 205 -3036 388 -3035
rect 716 -3036 1158 -3035
rect 1269 -3036 1305 -3035
rect 310 -3038 318 -3037
rect 338 -3038 374 -3037
rect 387 -3038 528 -3037
rect 716 -3038 745 -3037
rect 751 -3038 773 -3037
rect 1003 -3038 1186 -3037
rect 1269 -3038 1438 -3037
rect 184 -3040 745 -3039
rect 1066 -3040 1081 -3039
rect 184 -3042 801 -3041
rect 1080 -3042 1410 -3041
rect 310 -3044 626 -3043
rect 723 -3044 759 -3043
rect 800 -3044 1620 -3043
rect 324 -3046 339 -3045
rect 345 -3046 626 -3045
rect 1409 -3046 1452 -3045
rect 324 -3048 332 -3047
rect 345 -3048 696 -3047
rect 786 -3048 1452 -3047
rect 331 -3050 367 -3049
rect 485 -3050 1438 -3049
rect 114 -3052 367 -3051
rect 485 -3052 591 -3051
rect 352 -3054 493 -3053
rect 520 -3054 773 -3053
rect 152 -3056 353 -3055
rect 359 -3056 538 -3055
rect 590 -3056 916 -3055
rect 471 -3058 521 -3057
rect 527 -3058 766 -3057
rect 915 -3058 1480 -3057
rect 471 -3060 738 -3059
rect 765 -3060 808 -3059
rect 1479 -3060 1501 -3059
rect 534 -3062 1004 -3061
rect 1500 -3062 1543 -3061
rect 233 -3064 535 -3063
rect 737 -3064 1396 -3063
rect 1444 -3064 1543 -3063
rect 233 -3066 241 -3065
rect 807 -3066 829 -3065
rect 1444 -3066 1473 -3065
rect 240 -3068 248 -3067
rect 828 -3068 1508 -3067
rect 247 -3070 780 -3069
rect 831 -3070 1473 -3069
rect 597 -3072 780 -3071
rect 597 -3074 636 -3073
rect 30 -3085 475 -3084
rect 478 -3085 636 -3084
rect 646 -3085 976 -3084
rect 999 -3085 1634 -3084
rect 37 -3087 87 -3086
rect 114 -3087 213 -3086
rect 215 -3087 255 -3086
rect 275 -3087 801 -3086
rect 814 -3087 1088 -3086
rect 1090 -3087 1389 -3086
rect 1475 -3087 1571 -3086
rect 61 -3089 626 -3088
rect 656 -3089 780 -3088
rect 789 -3089 843 -3088
rect 877 -3089 1172 -3088
rect 1388 -3089 1564 -3088
rect 65 -3091 80 -3090
rect 82 -3091 437 -3090
rect 471 -3091 804 -3090
rect 842 -3091 983 -3090
rect 1020 -3091 1459 -3090
rect 79 -3093 696 -3092
rect 716 -3093 916 -3092
rect 933 -3093 1091 -3092
rect 1171 -3093 1340 -3092
rect 1444 -3093 1459 -3092
rect 86 -3095 178 -3094
rect 184 -3095 951 -3094
rect 975 -3095 1032 -3094
rect 1062 -3095 1585 -3094
rect 117 -3097 1277 -3096
rect 1339 -3097 1529 -3096
rect 131 -3099 206 -3098
rect 219 -3099 223 -3098
rect 254 -3099 927 -3098
rect 933 -3099 1200 -3098
rect 1276 -3099 1431 -3098
rect 135 -3101 164 -3100
rect 177 -3101 241 -3100
rect 282 -3101 395 -3100
rect 404 -3101 437 -3100
rect 453 -3101 927 -3100
rect 940 -3101 1200 -3100
rect 1423 -3101 1445 -3100
rect 51 -3103 283 -3102
rect 303 -3103 503 -3102
rect 527 -3103 626 -3102
rect 674 -3103 762 -3102
rect 779 -3103 1039 -3102
rect 1083 -3103 1368 -3102
rect 1423 -3103 1606 -3102
rect 93 -3105 304 -3104
rect 345 -3105 353 -3104
rect 366 -3105 584 -3104
rect 593 -3105 661 -3104
rect 674 -3105 745 -3104
rect 758 -3105 920 -3104
rect 940 -3105 1060 -3104
rect 1367 -3105 1543 -3104
rect 1605 -3105 1648 -3104
rect 93 -3107 738 -3106
rect 744 -3107 892 -3106
rect 919 -3107 1053 -3106
rect 1430 -3107 1613 -3106
rect 135 -3109 682 -3108
rect 684 -3109 1361 -3108
rect 142 -3111 1487 -3110
rect 142 -3113 773 -3112
rect 793 -3113 797 -3112
rect 800 -3113 839 -3112
rect 877 -3113 1025 -3112
rect 1031 -3113 1088 -3112
rect 1360 -3113 1536 -3112
rect 145 -3115 171 -3114
rect 184 -3115 514 -3114
rect 534 -3115 829 -3114
rect 838 -3115 1067 -3114
rect 1486 -3115 1627 -3114
rect 121 -3117 535 -3116
rect 562 -3117 647 -3116
rect 660 -3117 783 -3116
rect 793 -3117 1641 -3116
rect 100 -3119 122 -3118
rect 149 -3119 1396 -3118
rect 89 -3121 101 -3120
rect 152 -3121 269 -3120
rect 348 -3121 381 -3120
rect 394 -3121 507 -3120
rect 562 -3121 822 -3120
rect 828 -3121 969 -3120
rect 982 -3121 1130 -3120
rect 44 -3123 269 -3122
rect 352 -3123 591 -3122
rect 618 -3123 703 -3122
rect 716 -3123 836 -3122
rect 947 -3123 1165 -3122
rect 152 -3125 787 -3124
rect 821 -3125 1102 -3124
rect 1129 -3125 1284 -3124
rect 156 -3127 507 -3126
rect 576 -3127 1060 -3126
rect 1066 -3127 1235 -3126
rect 1283 -3127 1466 -3126
rect 156 -3129 654 -3128
rect 688 -3129 724 -3128
rect 730 -3129 815 -3128
rect 835 -3129 1354 -3128
rect 163 -3131 741 -3130
rect 772 -3131 1074 -3130
rect 1164 -3131 1270 -3130
rect 170 -3133 402 -3132
rect 429 -3133 584 -3132
rect 653 -3133 689 -3132
rect 691 -3133 1599 -3132
rect 191 -3135 202 -3134
rect 219 -3135 444 -3134
rect 457 -3135 514 -3134
rect 579 -3135 1102 -3134
rect 1234 -3135 1410 -3134
rect 128 -3137 458 -3136
rect 478 -3137 752 -3136
rect 786 -3137 899 -3136
rect 947 -3137 1403 -3136
rect 1409 -3137 1515 -3136
rect 72 -3139 129 -3138
rect 191 -3139 248 -3138
rect 261 -3139 444 -3138
rect 492 -3139 528 -3138
rect 681 -3139 724 -3138
rect 730 -3139 850 -3138
rect 898 -3139 990 -3138
rect 1003 -3139 1074 -3138
rect 1269 -3139 1522 -3138
rect 72 -3141 227 -3140
rect 233 -3141 248 -3140
rect 261 -3141 290 -3140
rect 366 -3141 416 -3140
rect 432 -3141 465 -3140
rect 492 -3141 549 -3140
rect 695 -3141 825 -3140
rect 849 -3141 955 -3140
rect 968 -3141 1228 -3140
rect 1297 -3141 1515 -3140
rect 198 -3143 1081 -3142
rect 1178 -3143 1298 -3142
rect 1325 -3143 1522 -3142
rect 149 -3145 1081 -3144
rect 1178 -3145 1312 -3144
rect 1325 -3145 1501 -3144
rect 198 -3147 871 -3146
rect 954 -3147 1151 -3146
rect 1227 -3147 1417 -3146
rect 222 -3149 290 -3148
rect 369 -3149 409 -3148
rect 537 -3149 1417 -3148
rect 226 -3151 605 -3150
rect 702 -3151 857 -3150
rect 870 -3151 1413 -3150
rect 233 -3153 612 -3152
rect 737 -3153 766 -3152
rect 856 -3153 885 -3152
rect 989 -3153 1438 -3152
rect 373 -3155 416 -3154
rect 548 -3155 668 -3154
rect 751 -3155 906 -3154
rect 1003 -3155 1158 -3154
rect 1311 -3155 1480 -3154
rect 107 -3157 374 -3156
rect 380 -3157 542 -3156
rect 597 -3157 605 -3156
rect 611 -3157 710 -3156
rect 765 -3157 1014 -3156
rect 1024 -3157 1116 -3156
rect 1122 -3157 1501 -3156
rect 107 -3159 640 -3158
rect 667 -3159 864 -3158
rect 884 -3159 1011 -3158
rect 1038 -3159 1249 -3158
rect 1402 -3159 1592 -3158
rect 387 -3161 465 -3160
rect 471 -3161 864 -3160
rect 905 -3161 913 -3160
rect 1052 -3161 1221 -3160
rect 1248 -3161 1508 -3160
rect 387 -3163 1144 -3162
rect 1150 -3163 1214 -3162
rect 1220 -3163 1382 -3162
rect 1437 -3163 1620 -3162
rect 401 -3165 521 -3164
rect 590 -3165 598 -3164
rect 632 -3165 1214 -3164
rect 1304 -3165 1508 -3164
rect 114 -3167 521 -3166
rect 632 -3167 962 -3166
rect 978 -3167 1305 -3166
rect 1381 -3167 1557 -3166
rect 408 -3169 570 -3168
rect 639 -3169 1207 -3168
rect 429 -3171 570 -3170
rect 709 -3171 808 -3170
rect 912 -3171 1046 -3170
rect 1094 -3171 1116 -3170
rect 1122 -3171 1319 -3170
rect 576 -3173 808 -3172
rect 961 -3173 1109 -3172
rect 1136 -3173 1158 -3172
rect 1185 -3173 1480 -3172
rect 1045 -3175 1193 -3174
rect 1206 -3175 1375 -3174
rect 1094 -3177 1263 -3176
rect 1318 -3177 1494 -3176
rect 996 -3179 1494 -3178
rect 996 -3181 1396 -3180
rect 1017 -3183 1263 -3182
rect 1374 -3183 1550 -3182
rect 1017 -3185 1291 -3184
rect 1108 -3187 1655 -3186
rect 1136 -3189 1256 -3188
rect 1290 -3189 1473 -3188
rect 1143 -3191 1242 -3190
rect 1255 -3191 1452 -3190
rect 450 -3193 1452 -3192
rect 310 -3195 451 -3194
rect 1185 -3195 1333 -3194
rect 310 -3197 332 -3196
rect 621 -3197 1333 -3196
rect 331 -3199 423 -3198
rect 1192 -3199 1347 -3198
rect 422 -3201 486 -3200
rect 1241 -3201 1578 -3200
rect 296 -3203 486 -3202
rect 1346 -3203 1466 -3202
rect 296 -3205 339 -3204
rect 338 -3207 360 -3206
rect 359 -3209 556 -3208
rect 499 -3211 556 -3210
rect 275 -3213 500 -3212
rect 65 -3224 115 -3223
rect 121 -3224 500 -3223
rect 502 -3224 717 -3223
rect 779 -3224 871 -3223
rect 880 -3224 1032 -3223
rect 1059 -3224 1333 -3223
rect 1346 -3224 1480 -3223
rect 1584 -3224 1606 -3223
rect 72 -3226 472 -3225
rect 485 -3226 580 -3225
rect 593 -3226 675 -3225
rect 684 -3226 787 -3225
rect 800 -3226 1357 -3225
rect 1409 -3226 1522 -3225
rect 86 -3228 402 -3227
rect 404 -3228 528 -3227
rect 544 -3228 556 -3227
rect 576 -3228 612 -3227
rect 625 -3228 797 -3227
rect 800 -3228 850 -3227
rect 894 -3228 1158 -3227
rect 1185 -3228 1210 -3227
rect 1297 -3228 1494 -3227
rect 142 -3230 577 -3229
rect 611 -3230 738 -3229
rect 849 -3230 955 -3229
rect 999 -3230 1004 -3229
rect 1010 -3230 1270 -3229
rect 1300 -3230 1466 -3229
rect 149 -3232 192 -3231
rect 212 -3232 241 -3231
rect 243 -3232 318 -3231
rect 324 -3232 1014 -3231
rect 1020 -3232 1137 -3231
rect 1269 -3232 1382 -3231
rect 1458 -3232 1532 -3231
rect 107 -3234 213 -3233
rect 226 -3234 486 -3233
rect 492 -3234 773 -3233
rect 905 -3234 986 -3233
rect 1010 -3234 1207 -3233
rect 1325 -3234 1329 -3233
rect 1332 -3234 1389 -3233
rect 152 -3236 360 -3235
rect 387 -3236 391 -3235
rect 415 -3236 542 -3235
rect 544 -3236 836 -3235
rect 905 -3236 1249 -3235
rect 1325 -3236 1361 -3235
rect 1381 -3236 1508 -3235
rect 156 -3238 528 -3237
rect 541 -3238 948 -3237
rect 954 -3238 1200 -3237
rect 1346 -3238 1424 -3237
rect 170 -3240 493 -3239
rect 499 -3240 549 -3239
rect 555 -3240 605 -3239
rect 625 -3240 808 -3239
rect 940 -3240 997 -3239
rect 1031 -3240 1221 -3239
rect 1349 -3240 1515 -3239
rect 93 -3242 171 -3241
rect 177 -3242 349 -3241
rect 359 -3242 395 -3241
rect 429 -3242 451 -3241
rect 457 -3242 591 -3241
rect 604 -3242 668 -3241
rect 705 -3242 1018 -3241
rect 1087 -3242 1319 -3241
rect 1353 -3242 1487 -3241
rect 191 -3244 206 -3243
rect 226 -3244 839 -3243
rect 940 -3244 983 -3243
rect 996 -3244 1172 -3243
rect 1199 -3244 1242 -3243
rect 1283 -3244 1354 -3243
rect 1388 -3244 1396 -3243
rect 205 -3246 633 -3245
rect 653 -3246 703 -3245
rect 709 -3246 825 -3245
rect 919 -3246 1284 -3245
rect 247 -3248 496 -3247
rect 520 -3248 780 -3247
rect 919 -3248 1081 -3247
rect 1090 -3248 1179 -3247
rect 1220 -3248 1438 -3247
rect 135 -3250 248 -3249
rect 254 -3250 678 -3249
rect 709 -3250 902 -3249
rect 947 -3250 1116 -3249
rect 1129 -3250 1189 -3249
rect 1234 -3250 1242 -3249
rect 128 -3252 136 -3251
rect 254 -3252 703 -3251
rect 716 -3252 829 -3251
rect 891 -3252 1179 -3251
rect 1234 -3252 1305 -3251
rect 261 -3254 395 -3253
rect 429 -3254 790 -3253
rect 828 -3254 1501 -3253
rect 261 -3256 332 -3255
rect 338 -3256 440 -3255
rect 450 -3256 479 -3255
rect 520 -3256 570 -3255
rect 632 -3256 731 -3255
rect 737 -3256 1074 -3255
rect 1080 -3256 1263 -3255
rect 1304 -3256 1476 -3255
rect 198 -3258 731 -3257
rect 751 -3258 1137 -3257
rect 1171 -3258 1277 -3257
rect 79 -3260 199 -3259
rect 275 -3260 332 -3259
rect 352 -3260 479 -3259
rect 548 -3260 661 -3259
rect 667 -3260 745 -3259
rect 751 -3260 1228 -3259
rect 1276 -3260 1375 -3259
rect 184 -3262 276 -3261
rect 282 -3262 339 -3261
rect 352 -3262 409 -3261
rect 422 -3262 570 -3261
rect 660 -3262 682 -3261
rect 723 -3262 808 -3261
rect 891 -3262 1263 -3261
rect 163 -3264 409 -3263
rect 422 -3264 619 -3263
rect 681 -3264 696 -3263
rect 723 -3264 843 -3263
rect 968 -3264 1004 -3263
rect 1052 -3264 1319 -3263
rect 100 -3266 164 -3265
rect 184 -3266 535 -3265
rect 618 -3266 990 -3265
rect 1045 -3266 1053 -3265
rect 1073 -3266 1144 -3265
rect 1213 -3266 1228 -3265
rect 282 -3268 951 -3267
rect 968 -3268 1039 -3267
rect 1045 -3268 1256 -3267
rect 296 -3270 325 -3269
rect 373 -3270 416 -3269
rect 457 -3270 794 -3269
rect 814 -3270 1039 -3269
rect 1094 -3270 1259 -3269
rect 296 -3272 381 -3271
rect 387 -3272 444 -3271
rect 471 -3272 531 -3271
rect 534 -3272 983 -3271
rect 1094 -3272 1291 -3271
rect 303 -3274 374 -3273
rect 380 -3274 514 -3273
rect 695 -3274 878 -3273
rect 1101 -3274 1158 -3273
rect 1290 -3274 1445 -3273
rect 303 -3276 311 -3275
rect 317 -3276 346 -3275
rect 443 -3276 647 -3275
rect 744 -3276 822 -3275
rect 842 -3276 1340 -3275
rect 177 -3278 346 -3277
rect 513 -3278 584 -3277
rect 758 -3278 878 -3277
rect 1101 -3278 1417 -3277
rect 289 -3280 311 -3279
rect 464 -3280 584 -3279
rect 758 -3280 885 -3279
rect 1115 -3280 1431 -3279
rect 289 -3282 437 -3281
rect 464 -3282 689 -3281
rect 772 -3282 1266 -3281
rect 1311 -3282 1340 -3281
rect 366 -3284 437 -3283
rect 793 -3284 962 -3283
rect 1129 -3284 1165 -3283
rect 1311 -3284 1368 -3283
rect 219 -3286 367 -3285
rect 814 -3286 1025 -3285
rect 1143 -3286 1151 -3285
rect 1164 -3286 1193 -3285
rect 1328 -3286 1361 -3285
rect 219 -3288 563 -3287
rect 821 -3288 934 -3287
rect 1150 -3288 1256 -3287
rect 506 -3290 563 -3289
rect 856 -3290 885 -3289
rect 915 -3290 962 -3289
rect 1192 -3290 1403 -3289
rect 506 -3292 766 -3291
rect 856 -3292 899 -3291
rect 926 -3292 1025 -3291
rect 765 -3294 913 -3293
rect 926 -3294 1067 -3293
rect 863 -3296 990 -3295
rect 1066 -3296 1214 -3295
rect 639 -3298 864 -3297
rect 912 -3298 976 -3297
rect 639 -3300 657 -3299
rect 933 -3300 1109 -3299
rect 835 -3302 1109 -3301
rect 975 -3304 1123 -3303
rect 1122 -3306 1452 -3305
rect 131 -3317 136 -3316
rect 163 -3317 580 -3316
rect 590 -3317 689 -3316
rect 691 -3317 1158 -3316
rect 1178 -3317 1529 -3316
rect 1577 -3317 1585 -3316
rect 205 -3319 542 -3318
rect 590 -3319 843 -3318
rect 870 -3319 1193 -3318
rect 1209 -3319 1277 -3318
rect 1360 -3319 1375 -3318
rect 233 -3321 493 -3320
rect 506 -3321 804 -3320
rect 870 -3321 986 -3320
rect 1003 -3321 1109 -3320
rect 1111 -3321 1291 -3320
rect 212 -3323 507 -3322
rect 513 -3323 545 -3322
rect 614 -3323 1151 -3322
rect 1153 -3323 1235 -3322
rect 1248 -3323 1326 -3322
rect 247 -3325 444 -3324
rect 464 -3325 675 -3324
rect 705 -3325 878 -3324
rect 880 -3325 1137 -3324
rect 1192 -3325 1284 -3324
rect 198 -3327 248 -3326
rect 268 -3327 619 -3326
rect 621 -3327 909 -3326
rect 915 -3327 1144 -3326
rect 1199 -3327 1249 -3326
rect 1262 -3327 1312 -3326
rect 240 -3329 269 -3328
rect 310 -3329 402 -3328
rect 436 -3329 472 -3328
rect 485 -3329 951 -3328
rect 961 -3329 1158 -3328
rect 1171 -3329 1200 -3328
rect 1213 -3329 1242 -3328
rect 1311 -3329 1333 -3328
rect 177 -3331 241 -3330
rect 359 -3331 514 -3330
rect 523 -3331 689 -3330
rect 716 -3331 878 -3330
rect 894 -3331 1217 -3330
rect 1234 -3331 1319 -3330
rect 1332 -3331 1382 -3330
rect 359 -3333 367 -3332
rect 380 -3333 444 -3332
rect 471 -3333 500 -3332
rect 618 -3333 710 -3332
rect 716 -3333 780 -3332
rect 789 -3333 801 -3332
rect 901 -3333 941 -3332
rect 947 -3333 1137 -3332
rect 1171 -3333 1298 -3332
rect 1353 -3333 1382 -3332
rect 170 -3335 500 -3334
rect 632 -3335 899 -3334
rect 947 -3335 969 -3334
rect 982 -3335 1165 -3334
rect 1213 -3335 1319 -3334
rect 275 -3337 367 -3336
rect 380 -3337 447 -3336
rect 478 -3337 486 -3336
rect 632 -3337 724 -3336
rect 730 -3337 874 -3336
rect 898 -3337 927 -3336
rect 961 -3337 1102 -3336
rect 1164 -3337 1270 -3336
rect 394 -3339 465 -3338
rect 478 -3339 521 -3338
rect 639 -3339 780 -3338
rect 891 -3339 927 -3338
rect 982 -3339 1123 -3338
rect 1241 -3339 1340 -3338
rect 345 -3341 395 -3340
rect 401 -3341 416 -3340
rect 576 -3341 640 -3340
rect 667 -3341 843 -3340
rect 996 -3341 1102 -3340
rect 282 -3343 346 -3342
rect 548 -3343 577 -3342
rect 667 -3343 745 -3342
rect 758 -3343 969 -3342
rect 1003 -3343 1088 -3342
rect 1094 -3343 1123 -3342
rect 184 -3345 283 -3344
rect 317 -3345 416 -3344
rect 530 -3345 1088 -3344
rect 226 -3347 549 -3346
rect 583 -3347 759 -3346
rect 863 -3347 997 -3346
rect 1013 -3347 1221 -3346
rect 219 -3349 584 -3348
rect 674 -3349 829 -3348
rect 1024 -3349 1130 -3348
rect 317 -3351 332 -3350
rect 408 -3351 864 -3350
rect 1024 -3351 1228 -3350
rect 296 -3353 332 -3352
rect 373 -3353 409 -3352
rect 709 -3353 773 -3352
rect 828 -3353 885 -3352
rect 1031 -3353 1035 -3352
rect 1038 -3353 1186 -3352
rect 191 -3355 297 -3354
rect 660 -3355 773 -3354
rect 814 -3355 885 -3354
rect 989 -3355 1039 -3354
rect 1045 -3355 1144 -3354
rect 1185 -3355 1207 -3354
rect 261 -3357 374 -3356
rect 660 -3357 766 -3356
rect 849 -3357 990 -3356
rect 1031 -3357 1116 -3356
rect 1206 -3357 1252 -3356
rect 681 -3359 815 -3358
rect 1034 -3359 1116 -3358
rect 681 -3361 1063 -3360
rect 1066 -3361 1095 -3360
rect 702 -3363 766 -3362
rect 786 -3363 850 -3362
rect 1045 -3363 1074 -3362
rect 1080 -3363 1130 -3362
rect 646 -3365 703 -3364
rect 723 -3365 794 -3364
rect 856 -3365 1081 -3364
rect 611 -3367 794 -3366
rect 856 -3367 1168 -3366
rect 254 -3369 612 -3368
rect 646 -3369 752 -3368
rect 786 -3369 801 -3368
rect 933 -3369 1074 -3368
rect 737 -3371 941 -3370
rect 1052 -3371 1109 -3370
rect 737 -3373 808 -3372
rect 933 -3373 1021 -3372
rect 1066 -3373 1266 -3372
rect 387 -3375 1021 -3374
rect 1265 -3375 1347 -3374
rect 387 -3377 458 -3376
rect 597 -3377 808 -3376
rect 450 -3379 458 -3378
rect 597 -3379 696 -3378
rect 744 -3379 822 -3378
rect 450 -3381 528 -3380
rect 695 -3381 836 -3380
rect 527 -3383 535 -3382
rect 562 -3383 836 -3382
rect 534 -3385 556 -3384
rect 562 -3385 570 -3384
rect 751 -3385 913 -3384
rect 555 -3387 626 -3386
rect 821 -3387 920 -3386
rect 569 -3389 605 -3388
rect 625 -3389 654 -3388
rect 912 -3389 955 -3388
rect 422 -3391 654 -3390
rect 919 -3391 976 -3390
rect 338 -3393 423 -3392
rect 604 -3393 906 -3392
rect 954 -3393 1018 -3392
rect 338 -3395 353 -3394
rect 905 -3395 1011 -3394
rect 324 -3397 353 -3396
rect 975 -3397 1060 -3396
rect 303 -3399 325 -3398
rect 1059 -3399 1305 -3398
rect 289 -3401 304 -3400
rect 289 -3403 311 -3402
rect 240 -3414 262 -3413
rect 268 -3414 293 -3413
rect 338 -3414 356 -3413
rect 376 -3414 451 -3413
rect 457 -3414 475 -3413
rect 485 -3414 612 -3413
rect 663 -3414 1039 -3413
rect 1041 -3414 1046 -3413
rect 1052 -3414 1074 -3413
rect 1111 -3414 1193 -3413
rect 1199 -3414 1214 -3413
rect 1248 -3414 1270 -3413
rect 1304 -3414 1312 -3413
rect 1318 -3414 1347 -3413
rect 1374 -3414 1396 -3413
rect 247 -3416 290 -3415
rect 317 -3416 458 -3415
rect 499 -3416 605 -3415
rect 702 -3416 811 -3415
rect 824 -3416 983 -3415
rect 989 -3416 1056 -3415
rect 1073 -3416 1102 -3415
rect 1122 -3416 1126 -3415
rect 1129 -3416 1161 -3415
rect 1185 -3416 1193 -3415
rect 1318 -3416 1333 -3415
rect 1381 -3416 1385 -3415
rect 282 -3418 318 -3417
rect 324 -3418 339 -3417
rect 352 -3418 374 -3417
rect 394 -3418 500 -3417
rect 513 -3418 657 -3417
rect 702 -3418 738 -3417
rect 793 -3418 804 -3417
rect 863 -3418 1266 -3417
rect 1381 -3418 1389 -3417
rect 366 -3420 395 -3419
rect 415 -3420 514 -3419
rect 520 -3420 528 -3419
rect 562 -3420 731 -3419
rect 733 -3420 787 -3419
rect 800 -3420 815 -3419
rect 842 -3420 864 -3419
rect 884 -3420 892 -3419
rect 898 -3420 1000 -3419
rect 1017 -3420 1032 -3419
rect 1080 -3420 1200 -3419
rect 359 -3422 521 -3421
rect 562 -3422 591 -3421
rect 625 -3422 731 -3421
rect 751 -3422 885 -3421
rect 898 -3422 906 -3421
rect 919 -3422 990 -3421
rect 996 -3422 1011 -3421
rect 1024 -3422 1172 -3421
rect 359 -3424 510 -3423
rect 576 -3424 598 -3423
rect 625 -3424 647 -3423
rect 681 -3424 738 -3423
rect 758 -3424 787 -3423
rect 807 -3424 843 -3423
rect 849 -3424 892 -3423
rect 919 -3424 962 -3423
rect 968 -3424 1168 -3423
rect 366 -3426 388 -3425
rect 415 -3426 437 -3425
rect 443 -3426 587 -3425
rect 597 -3426 696 -3425
rect 751 -3426 850 -3425
rect 877 -3426 1011 -3425
rect 1031 -3426 1151 -3425
rect 1153 -3426 1207 -3425
rect 303 -3428 444 -3427
rect 450 -3428 479 -3427
rect 492 -3428 605 -3427
rect 618 -3428 696 -3427
rect 758 -3428 822 -3427
rect 877 -3428 895 -3427
rect 940 -3428 1018 -3427
rect 1087 -3428 1214 -3427
rect 380 -3430 388 -3429
rect 408 -3430 437 -3429
rect 464 -3430 528 -3429
rect 548 -3430 808 -3429
rect 814 -3430 829 -3429
rect 912 -3430 941 -3429
rect 954 -3430 983 -3429
rect 1003 -3430 1025 -3429
rect 1101 -3430 1116 -3429
rect 1122 -3430 1137 -3429
rect 1157 -3430 1235 -3429
rect 331 -3432 381 -3431
rect 401 -3432 465 -3431
rect 471 -3432 479 -3431
rect 492 -3432 535 -3431
rect 548 -3432 556 -3431
rect 579 -3432 1081 -3431
rect 1094 -3432 1116 -3431
rect 1129 -3432 1301 -3431
rect 299 -3434 402 -3433
rect 422 -3434 524 -3433
rect 534 -3434 542 -3433
rect 646 -3434 661 -3433
rect 681 -3434 710 -3433
rect 772 -3434 906 -3433
rect 912 -3434 927 -3433
rect 933 -3434 955 -3433
rect 961 -3434 976 -3433
rect 1003 -3434 1067 -3433
rect 1136 -3434 1144 -3433
rect 1206 -3434 1242 -3433
rect 345 -3436 423 -3435
rect 471 -3436 542 -3435
rect 709 -3436 745 -3435
rect 765 -3436 976 -3435
rect 1384 -3436 1389 -3435
rect 310 -3438 346 -3437
rect 485 -3438 661 -3437
rect 716 -3438 766 -3437
rect 779 -3438 794 -3437
rect 821 -3438 1217 -3437
rect 310 -3440 353 -3439
rect 506 -3440 556 -3439
rect 653 -3440 780 -3439
rect 828 -3440 836 -3439
rect 933 -3440 997 -3439
rect 506 -3442 622 -3441
rect 674 -3442 717 -3441
rect 723 -3442 773 -3441
rect 835 -3442 948 -3441
rect 667 -3444 675 -3443
rect 723 -3444 853 -3443
rect 870 -3444 948 -3443
rect 614 -3446 668 -3445
rect 744 -3446 857 -3445
rect 870 -3446 1021 -3445
rect 583 -3448 857 -3447
rect 583 -3450 927 -3449
rect 261 -3461 269 -3460
rect 296 -3461 311 -3460
rect 317 -3461 356 -3460
rect 359 -3461 412 -3460
rect 439 -3461 657 -3460
rect 660 -3461 734 -3460
rect 800 -3461 808 -3460
rect 821 -3461 829 -3460
rect 842 -3461 916 -3460
rect 940 -3461 944 -3460
rect 947 -3461 1007 -3460
rect 1010 -3461 1060 -3460
rect 1066 -3461 1074 -3460
rect 1087 -3461 1102 -3460
rect 1115 -3461 1119 -3460
rect 1143 -3461 1158 -3460
rect 1181 -3461 1417 -3460
rect 373 -3463 391 -3462
rect 401 -3463 584 -3462
rect 611 -3463 720 -3462
rect 786 -3463 801 -3462
rect 807 -3463 815 -3462
rect 828 -3463 871 -3462
rect 940 -3463 962 -3462
rect 968 -3463 983 -3462
rect 989 -3463 1011 -3462
rect 1017 -3463 1046 -3462
rect 1073 -3463 1130 -3462
rect 1185 -3463 1207 -3462
rect 1213 -3463 1249 -3462
rect 1269 -3463 1277 -3462
rect 1297 -3463 1319 -3462
rect 1374 -3463 1382 -3462
rect 345 -3465 374 -3464
rect 380 -3465 409 -3464
rect 520 -3465 591 -3464
rect 618 -3465 626 -3464
rect 632 -3465 664 -3464
rect 667 -3465 755 -3464
rect 765 -3465 787 -3464
rect 852 -3465 920 -3464
rect 954 -3465 962 -3464
rect 975 -3465 1039 -3464
rect 1080 -3465 1270 -3464
rect 1300 -3465 1305 -3464
rect 1346 -3465 1382 -3464
rect 366 -3467 381 -3466
rect 387 -3467 426 -3466
rect 506 -3467 591 -3466
rect 618 -3467 724 -3466
rect 758 -3467 766 -3466
rect 772 -3467 815 -3466
rect 856 -3467 948 -3466
rect 975 -3467 1004 -3466
rect 1115 -3467 1123 -3466
rect 1199 -3467 1235 -3466
rect 338 -3469 367 -3468
rect 450 -3469 507 -3468
rect 527 -3469 622 -3468
rect 653 -3469 682 -3468
rect 695 -3469 759 -3468
rect 891 -3469 920 -3468
rect 926 -3469 1081 -3468
rect 1118 -3469 1123 -3468
rect 429 -3471 451 -3470
rect 499 -3471 528 -3470
rect 534 -3471 633 -3470
rect 653 -3471 1091 -3470
rect 394 -3473 430 -3472
rect 457 -3473 500 -3472
rect 534 -3473 608 -3472
rect 695 -3473 745 -3472
rect 884 -3473 892 -3472
rect 905 -3473 927 -3472
rect 1003 -3473 1179 -3472
rect 436 -3475 458 -3474
rect 541 -3475 587 -3474
rect 702 -3475 717 -3474
rect 723 -3475 752 -3474
rect 863 -3475 885 -3474
rect 898 -3475 906 -3474
rect 478 -3477 542 -3476
rect 548 -3477 594 -3476
rect 688 -3477 703 -3476
rect 709 -3477 822 -3476
rect 898 -3477 913 -3476
rect 464 -3479 479 -3478
rect 548 -3479 577 -3478
rect 646 -3479 710 -3478
rect 730 -3479 773 -3478
rect 779 -3479 913 -3478
rect 555 -3481 584 -3480
rect 674 -3481 689 -3480
rect 730 -3481 836 -3480
rect 492 -3483 556 -3482
rect 562 -3483 577 -3482
rect 744 -3483 997 -3482
rect 443 -3485 493 -3484
rect 513 -3485 563 -3484
rect 569 -3485 647 -3484
rect 996 -3485 1032 -3484
rect 415 -3487 444 -3486
rect 569 -3487 598 -3486
rect 422 -3489 514 -3488
rect 422 -3491 472 -3490
rect 268 -3502 283 -3501
rect 285 -3502 297 -3501
rect 366 -3502 388 -3501
rect 390 -3502 395 -3501
rect 408 -3502 440 -3501
rect 450 -3502 482 -3501
rect 506 -3502 566 -3501
rect 583 -3502 598 -3501
rect 632 -3502 727 -3501
rect 733 -3502 1182 -3501
rect 1234 -3502 1280 -3501
rect 1374 -3502 1382 -3501
rect 1384 -3502 1389 -3501
rect 1416 -3502 1501 -3501
rect 373 -3504 402 -3503
rect 443 -3504 451 -3503
rect 457 -3504 465 -3503
rect 492 -3504 507 -3503
rect 520 -3504 549 -3503
rect 562 -3504 584 -3503
rect 590 -3504 657 -3503
rect 674 -3504 696 -3503
rect 737 -3504 755 -3503
rect 758 -3504 780 -3503
rect 786 -3504 790 -3503
rect 821 -3504 864 -3503
rect 905 -3504 913 -3503
rect 947 -3504 1035 -3503
rect 1045 -3504 1049 -3503
rect 1059 -3504 1091 -3503
rect 1122 -3504 1130 -3503
rect 1157 -3504 1165 -3503
rect 1178 -3504 1186 -3503
rect 1248 -3504 1263 -3503
rect 1269 -3504 1340 -3503
rect 429 -3506 444 -3505
rect 478 -3506 493 -3505
rect 527 -3506 559 -3505
rect 576 -3506 591 -3505
rect 646 -3506 731 -3505
rect 758 -3506 773 -3505
rect 786 -3506 794 -3505
rect 800 -3506 822 -3505
rect 842 -3506 1018 -3505
rect 1020 -3506 1074 -3505
rect 1080 -3506 1144 -3505
rect 429 -3508 479 -3507
rect 499 -3508 528 -3507
rect 541 -3508 549 -3507
rect 576 -3508 619 -3507
rect 639 -3508 647 -3507
rect 653 -3508 745 -3507
rect 765 -3508 773 -3507
rect 800 -3508 808 -3507
rect 884 -3508 906 -3507
rect 957 -3508 997 -3507
rect 1010 -3508 1042 -3507
rect 1045 -3508 1053 -3507
rect 1062 -3508 1067 -3507
rect 485 -3510 500 -3509
rect 513 -3510 542 -3509
rect 688 -3510 696 -3509
rect 709 -3510 731 -3509
rect 807 -3510 815 -3509
rect 877 -3510 885 -3509
rect 961 -3510 965 -3509
rect 968 -3510 976 -3509
rect 1024 -3510 1032 -3509
rect 1038 -3510 1074 -3509
rect 471 -3512 486 -3511
rect 513 -3512 535 -3511
rect 709 -3512 717 -3511
rect 765 -3512 1039 -3511
rect 1048 -3512 1053 -3511
rect 534 -3514 570 -3513
rect 814 -3514 829 -3513
rect 877 -3514 899 -3513
rect 954 -3514 962 -3513
rect 555 -3516 570 -3515
rect 891 -3516 899 -3515
rect 926 -3516 955 -3515
rect 926 -3518 934 -3517
rect 919 -3520 934 -3519
rect 919 -3522 948 -3521
rect 387 -3533 391 -3532
rect 408 -3533 430 -3532
rect 450 -3533 458 -3532
rect 464 -3533 475 -3532
rect 506 -3533 521 -3532
rect 558 -3533 1109 -3532
rect 1157 -3533 1165 -3532
rect 1262 -3533 1280 -3532
rect 1339 -3533 1361 -3532
rect 1381 -3533 1389 -3532
rect 1500 -3533 1581 -3532
rect 387 -3535 402 -3534
rect 443 -3535 451 -3534
rect 506 -3535 514 -3534
rect 565 -3535 654 -3534
rect 660 -3535 675 -3534
rect 695 -3535 706 -3534
rect 730 -3535 738 -3534
rect 796 -3535 801 -3534
rect 807 -3535 825 -3534
rect 884 -3535 892 -3534
rect 926 -3535 951 -3534
rect 957 -3535 969 -3534
rect 1038 -3535 1046 -3534
rect 1052 -3535 1060 -3534
rect 1073 -3535 1112 -3534
rect 1143 -3535 1165 -3534
rect 394 -3537 402 -3536
rect 499 -3537 514 -3536
rect 565 -3537 577 -3536
rect 604 -3537 608 -3536
rect 646 -3537 664 -3536
rect 667 -3537 766 -3536
rect 779 -3537 801 -3536
rect 877 -3537 885 -3536
rect 919 -3537 927 -3536
rect 933 -3537 937 -3536
rect 390 -3539 395 -3538
rect 492 -3539 500 -3538
rect 576 -3539 591 -3538
rect 702 -3539 710 -3538
rect 772 -3539 780 -3538
rect 793 -3539 808 -3538
rect 863 -3539 878 -3538
rect 485 -3541 493 -3540
rect 590 -3541 598 -3540
rect 772 -3541 843 -3540
rect 583 -3543 598 -3542
rect 555 -3545 584 -3544
rect 541 -3547 556 -3546
rect 534 -3549 542 -3548
rect 534 -3551 563 -3550
rect 401 -3562 405 -3561
rect 457 -3562 465 -3561
rect 474 -3562 479 -3561
rect 499 -3562 514 -3561
rect 527 -3562 542 -3561
rect 555 -3562 563 -3561
rect 569 -3562 577 -3561
rect 579 -3562 598 -3561
rect 632 -3562 668 -3561
rect 702 -3562 710 -3561
rect 737 -3562 748 -3561
rect 758 -3562 766 -3561
rect 768 -3562 780 -3561
rect 786 -3562 797 -3561
rect 877 -3562 895 -3561
rect 901 -3562 906 -3561
rect 926 -3562 951 -3561
rect 1111 -3562 1116 -3561
rect 1132 -3562 1137 -3561
rect 1164 -3562 1172 -3561
rect 1178 -3562 1186 -3561
rect 1192 -3562 1200 -3561
rect 1391 -3562 1396 -3561
rect 380 -3564 402 -3563
rect 450 -3564 458 -3563
rect 502 -3564 507 -3563
rect 530 -3564 535 -3563
rect 548 -3564 563 -3563
rect 576 -3564 584 -3563
rect 758 -3564 773 -3563
rect 793 -3564 808 -3563
rect 891 -3564 899 -3563
rect 933 -3564 941 -3563
rect 1129 -3564 1137 -3563
rect 1388 -3564 1396 -3563
rect 807 -3566 815 -3565
rect 1360 -3566 1389 -3565
rect 387 -3577 402 -3576
rect 457 -3577 465 -3576
rect 492 -3577 503 -3576
rect 562 -3577 580 -3576
rect 590 -3577 598 -3576
rect 600 -3577 633 -3576
rect 747 -3577 759 -3576
rect 800 -3577 811 -3576
rect 884 -3577 899 -3576
rect 1129 -3577 1137 -3576
rect 1171 -3577 1182 -3576
rect 1195 -3577 1200 -3576
rect 1388 -3577 1396 -3576
rect 397 -3579 409 -3578
rect 1178 -3579 1186 -3578
<< m2contact >>
rect 233 0 234 1
rect 436 0 437 1
rect 443 0 444 1
rect 457 0 458 1
rect 527 0 528 1
rect 548 0 549 1
rect 555 0 556 1
rect 754 0 755 1
rect 877 0 878 1
rect 954 0 955 1
rect 345 -2 346 -1
rect 352 -2 353 -1
rect 359 -2 360 -1
rect 467 -2 468 -1
rect 604 -2 605 -1
rect 614 -2 615 -1
rect 653 -2 654 -1
rect 677 -2 678 -1
rect 716 -2 717 -1
rect 800 -2 801 -1
rect 380 -4 381 -3
rect 534 -4 535 -3
rect 670 -4 671 -3
rect 688 -4 689 -3
rect 401 -6 402 -5
rect 460 -6 461 -5
rect 408 -8 409 -7
rect 432 -8 433 -7
rect 453 -8 454 -7
rect 471 -8 472 -7
rect 415 -10 416 -9
rect 506 -10 507 -9
rect 422 -12 423 -11
rect 450 -12 451 -11
rect 145 -23 146 -22
rect 149 -23 150 -22
rect 156 -23 157 -22
rect 233 -23 234 -22
rect 261 -23 262 -22
rect 306 -23 307 -22
rect 324 -23 325 -22
rect 359 -23 360 -22
rect 373 -23 374 -22
rect 408 -23 409 -22
rect 425 -23 426 -22
rect 443 -23 444 -22
rect 450 -23 451 -22
rect 555 -23 556 -22
rect 590 -23 591 -22
rect 821 -23 822 -22
rect 842 -23 843 -22
rect 884 -23 885 -22
rect 954 -23 955 -22
rect 989 -23 990 -22
rect 226 -25 227 -24
rect 236 -25 237 -24
rect 282 -25 283 -24
rect 390 -25 391 -24
rect 394 -25 395 -24
rect 415 -25 416 -24
rect 429 -25 430 -24
rect 443 -25 444 -24
rect 460 -25 461 -24
rect 555 -25 556 -24
rect 618 -25 619 -24
rect 632 -25 633 -24
rect 653 -25 654 -24
rect 667 -25 668 -24
rect 677 -25 678 -24
rect 681 -25 682 -24
rect 688 -25 689 -24
rect 702 -25 703 -24
rect 712 -25 713 -24
rect 772 -25 773 -24
rect 800 -25 801 -24
rect 828 -25 829 -24
rect 331 -27 332 -26
rect 380 -27 381 -26
rect 408 -27 409 -26
rect 562 -27 563 -26
rect 653 -27 654 -26
rect 670 -27 671 -26
rect 677 -27 678 -26
rect 730 -27 731 -26
rect 751 -27 752 -26
rect 996 -27 997 -26
rect 338 -29 339 -28
rect 345 -29 346 -28
rect 380 -29 381 -28
rect 401 -29 402 -28
rect 436 -29 437 -28
rect 660 -29 661 -28
rect 688 -29 689 -28
rect 719 -29 720 -28
rect 758 -29 759 -28
rect 898 -29 899 -28
rect 401 -31 402 -30
rect 422 -31 423 -30
rect 432 -31 433 -30
rect 436 -31 437 -30
rect 460 -31 461 -30
rect 744 -31 745 -30
rect 814 -31 815 -30
rect 880 -31 881 -30
rect 464 -33 465 -32
rect 597 -33 598 -32
rect 716 -33 717 -32
rect 754 -33 755 -32
rect 471 -35 472 -34
rect 478 -35 479 -34
rect 492 -35 493 -34
rect 506 -35 507 -34
rect 509 -35 510 -34
rect 611 -35 612 -34
rect 471 -37 472 -36
rect 516 -37 517 -36
rect 520 -37 521 -36
rect 639 -37 640 -36
rect 495 -39 496 -38
rect 499 -39 500 -38
rect 513 -39 514 -38
rect 625 -39 626 -38
rect 523 -41 524 -40
rect 541 -41 542 -40
rect 551 -41 552 -40
rect 576 -41 577 -40
rect 530 -43 531 -42
rect 548 -43 549 -42
rect 534 -45 535 -44
rect 646 -45 647 -44
rect 527 -47 528 -46
rect 534 -47 535 -46
rect 537 -47 538 -46
rect 583 -47 584 -46
rect 464 -49 465 -48
rect 527 -49 528 -48
rect 128 -60 129 -59
rect 156 -60 157 -59
rect 191 -60 192 -59
rect 198 -60 199 -59
rect 205 -60 206 -59
rect 226 -60 227 -59
rect 254 -60 255 -59
rect 432 -60 433 -59
rect 474 -60 475 -59
rect 737 -60 738 -59
rect 744 -60 745 -59
rect 870 -60 871 -59
rect 884 -60 885 -59
rect 940 -60 941 -59
rect 989 -60 990 -59
rect 1010 -60 1011 -59
rect 219 -62 220 -61
rect 282 -62 283 -61
rect 289 -62 290 -61
rect 324 -62 325 -61
rect 345 -62 346 -61
rect 422 -62 423 -61
rect 478 -62 479 -61
rect 488 -62 489 -61
rect 492 -62 493 -61
rect 709 -62 710 -61
rect 716 -62 717 -61
rect 744 -62 745 -61
rect 751 -62 752 -61
rect 887 -62 888 -61
rect 898 -62 899 -61
rect 954 -62 955 -61
rect 996 -62 997 -61
rect 1087 -62 1088 -61
rect 261 -64 262 -63
rect 268 -64 269 -63
rect 275 -64 276 -63
rect 457 -64 458 -63
rect 478 -64 479 -63
rect 590 -64 591 -63
rect 625 -64 626 -63
rect 695 -64 696 -63
rect 730 -64 731 -63
rect 786 -64 787 -63
rect 796 -64 797 -63
rect 863 -64 864 -63
rect 936 -64 937 -63
rect 947 -64 948 -63
rect 247 -66 248 -65
rect 261 -66 262 -65
rect 282 -66 283 -65
rect 460 -66 461 -65
rect 506 -66 507 -65
rect 520 -66 521 -65
rect 551 -66 552 -65
rect 677 -66 678 -65
rect 688 -66 689 -65
rect 716 -66 717 -65
rect 772 -66 773 -65
rect 835 -66 836 -65
rect 296 -68 297 -67
rect 408 -68 409 -67
rect 422 -68 423 -67
rect 436 -68 437 -67
rect 506 -68 507 -67
rect 593 -68 594 -67
rect 625 -68 626 -67
rect 810 -68 811 -67
rect 817 -68 818 -67
rect 856 -68 857 -67
rect 303 -70 304 -69
rect 338 -70 339 -69
rect 352 -70 353 -69
rect 415 -70 416 -69
rect 555 -70 556 -69
rect 674 -70 675 -69
rect 702 -70 703 -69
rect 730 -70 731 -69
rect 779 -70 780 -69
rect 884 -70 885 -69
rect 306 -72 307 -71
rect 359 -72 360 -71
rect 366 -72 367 -71
rect 401 -72 402 -71
rect 415 -72 416 -71
rect 516 -72 517 -71
rect 555 -72 556 -71
rect 576 -72 577 -71
rect 583 -72 584 -71
rect 688 -72 689 -71
rect 800 -72 801 -71
rect 828 -72 829 -71
rect 310 -74 311 -73
rect 450 -74 451 -73
rect 530 -74 531 -73
rect 583 -74 584 -73
rect 590 -74 591 -73
rect 618 -74 619 -73
rect 646 -74 647 -73
rect 709 -74 710 -73
rect 807 -74 808 -73
rect 842 -74 843 -73
rect 317 -76 318 -75
rect 331 -76 332 -75
rect 338 -76 339 -75
rect 464 -76 465 -75
rect 541 -76 542 -75
rect 576 -76 577 -75
rect 597 -76 598 -75
rect 702 -76 703 -75
rect 712 -76 713 -75
rect 842 -76 843 -75
rect 324 -78 325 -77
rect 373 -78 374 -77
rect 376 -78 377 -77
rect 380 -78 381 -77
rect 387 -78 388 -77
rect 436 -78 437 -77
rect 464 -78 465 -77
rect 471 -78 472 -77
rect 499 -78 500 -77
rect 541 -78 542 -77
rect 604 -78 605 -77
rect 618 -78 619 -77
rect 649 -78 650 -77
rect 793 -78 794 -77
rect 814 -78 815 -77
rect 828 -78 829 -77
rect 331 -80 332 -79
rect 443 -80 444 -79
rect 534 -80 535 -79
rect 597 -80 598 -79
rect 660 -80 661 -79
rect 723 -80 724 -79
rect 821 -80 822 -79
rect 891 -80 892 -79
rect 334 -82 335 -81
rect 499 -82 500 -81
rect 513 -82 514 -81
rect 534 -82 535 -81
rect 569 -82 570 -81
rect 604 -82 605 -81
rect 611 -82 612 -81
rect 660 -82 661 -81
rect 373 -84 374 -83
rect 380 -84 381 -83
rect 387 -84 388 -83
rect 523 -84 524 -83
rect 548 -84 549 -83
rect 569 -84 570 -83
rect 632 -84 633 -83
rect 821 -84 822 -83
rect 401 -86 402 -85
rect 429 -86 430 -85
rect 562 -86 563 -85
rect 611 -86 612 -85
rect 411 -88 412 -87
rect 450 -88 451 -87
rect 562 -88 563 -87
rect 653 -88 654 -87
rect 653 -90 654 -89
rect 667 -90 668 -89
rect 667 -92 668 -91
rect 681 -92 682 -91
rect 639 -94 640 -93
rect 681 -94 682 -93
rect 639 -96 640 -95
rect 758 -96 759 -95
rect 89 -107 90 -106
rect 93 -107 94 -106
rect 114 -107 115 -106
rect 128 -107 129 -106
rect 135 -107 136 -106
rect 219 -107 220 -106
rect 226 -107 227 -106
rect 292 -107 293 -106
rect 345 -107 346 -106
rect 362 -107 363 -106
rect 373 -107 374 -106
rect 394 -107 395 -106
rect 408 -107 409 -106
rect 467 -107 468 -106
rect 471 -107 472 -106
rect 488 -107 489 -106
rect 513 -107 514 -106
rect 548 -107 549 -106
rect 611 -107 612 -106
rect 646 -107 647 -106
rect 656 -107 657 -106
rect 744 -107 745 -106
rect 793 -107 794 -106
rect 821 -107 822 -106
rect 828 -107 829 -106
rect 912 -107 913 -106
rect 940 -107 941 -106
rect 996 -107 997 -106
rect 1010 -107 1011 -106
rect 1038 -107 1039 -106
rect 1087 -107 1088 -106
rect 1129 -107 1130 -106
rect 1195 -107 1196 -106
rect 1220 -107 1221 -106
rect 142 -109 143 -108
rect 254 -109 255 -108
rect 261 -109 262 -108
rect 471 -109 472 -108
rect 481 -109 482 -108
rect 551 -109 552 -108
rect 646 -109 647 -108
rect 716 -109 717 -108
rect 723 -109 724 -108
rect 849 -109 850 -108
rect 856 -109 857 -108
rect 898 -109 899 -108
rect 947 -109 948 -108
rect 968 -109 969 -108
rect 156 -111 157 -110
rect 331 -111 332 -110
rect 380 -111 381 -110
rect 383 -111 384 -110
rect 394 -111 395 -110
rect 639 -111 640 -110
rect 674 -111 675 -110
rect 758 -111 759 -110
rect 810 -111 811 -110
rect 940 -111 941 -110
rect 954 -111 955 -110
rect 982 -111 983 -110
rect 163 -113 164 -112
rect 205 -113 206 -112
rect 219 -113 220 -112
rect 303 -113 304 -112
rect 310 -113 311 -112
rect 373 -113 374 -112
rect 380 -113 381 -112
rect 443 -113 444 -112
rect 450 -113 451 -112
rect 457 -113 458 -112
rect 485 -113 486 -112
rect 509 -113 510 -112
rect 513 -113 514 -112
rect 933 -113 934 -112
rect 170 -115 171 -114
rect 355 -115 356 -114
rect 376 -115 377 -114
rect 485 -115 486 -114
rect 530 -115 531 -114
rect 548 -115 549 -114
rect 576 -115 577 -114
rect 639 -115 640 -114
rect 681 -115 682 -114
rect 723 -115 724 -114
rect 744 -115 745 -114
rect 800 -115 801 -114
rect 817 -115 818 -114
rect 828 -115 829 -114
rect 835 -115 836 -114
rect 919 -115 920 -114
rect 177 -117 178 -116
rect 338 -117 339 -116
rect 352 -117 353 -116
rect 457 -117 458 -116
rect 537 -117 538 -116
rect 625 -117 626 -116
rect 660 -117 661 -116
rect 800 -117 801 -116
rect 824 -117 825 -116
rect 1010 -117 1011 -116
rect 184 -119 185 -118
rect 191 -119 192 -118
rect 198 -119 199 -118
rect 247 -119 248 -118
rect 250 -119 251 -118
rect 310 -119 311 -118
rect 317 -119 318 -118
rect 331 -119 332 -118
rect 338 -119 339 -118
rect 632 -119 633 -118
rect 698 -119 699 -118
rect 905 -119 906 -118
rect 191 -121 192 -120
rect 275 -121 276 -120
rect 289 -121 290 -120
rect 429 -121 430 -120
rect 450 -121 451 -120
rect 502 -121 503 -120
rect 576 -121 577 -120
rect 653 -121 654 -120
rect 709 -121 710 -120
rect 807 -121 808 -120
rect 842 -121 843 -120
rect 961 -121 962 -120
rect 208 -123 209 -122
rect 317 -123 318 -122
rect 383 -123 384 -122
rect 443 -123 444 -122
rect 460 -123 461 -122
rect 632 -123 633 -122
rect 716 -123 717 -122
rect 768 -123 769 -122
rect 779 -123 780 -122
rect 835 -123 836 -122
rect 856 -123 857 -122
rect 877 -123 878 -122
rect 880 -123 881 -122
rect 926 -123 927 -122
rect 243 -125 244 -124
rect 345 -125 346 -124
rect 408 -125 409 -124
rect 422 -125 423 -124
rect 590 -125 591 -124
rect 674 -125 675 -124
rect 796 -125 797 -124
rect 842 -125 843 -124
rect 863 -125 864 -124
rect 954 -125 955 -124
rect 247 -127 248 -126
rect 520 -127 521 -126
rect 569 -127 570 -126
rect 590 -127 591 -126
rect 597 -127 598 -126
rect 681 -127 682 -126
rect 814 -127 815 -126
rect 863 -127 864 -126
rect 870 -127 871 -126
rect 975 -127 976 -126
rect 254 -129 255 -128
rect 282 -129 283 -128
rect 296 -129 297 -128
rect 422 -129 423 -128
rect 432 -129 433 -128
rect 597 -129 598 -128
rect 611 -129 612 -128
rect 660 -129 661 -128
rect 737 -129 738 -128
rect 814 -129 815 -128
rect 884 -129 885 -128
rect 1136 -129 1137 -128
rect 261 -131 262 -130
rect 474 -131 475 -130
rect 520 -131 521 -130
rect 947 -131 948 -130
rect 268 -133 269 -132
rect 303 -133 304 -132
rect 432 -133 433 -132
rect 464 -133 465 -132
rect 618 -133 619 -132
rect 709 -133 710 -132
rect 786 -133 787 -132
rect 870 -133 871 -132
rect 268 -135 269 -134
rect 366 -135 367 -134
rect 415 -135 416 -134
rect 464 -135 465 -134
rect 618 -135 619 -134
rect 751 -135 752 -134
rect 275 -137 276 -136
rect 562 -137 563 -136
rect 625 -137 626 -136
rect 667 -137 668 -136
rect 688 -137 689 -136
rect 751 -137 752 -136
rect 282 -139 283 -138
rect 387 -139 388 -138
rect 401 -139 402 -138
rect 415 -139 416 -138
rect 534 -139 535 -138
rect 562 -139 563 -138
rect 649 -139 650 -138
rect 779 -139 780 -138
rect 296 -141 297 -140
rect 478 -141 479 -140
rect 534 -141 535 -140
rect 555 -141 556 -140
rect 667 -141 668 -140
rect 793 -141 794 -140
rect 366 -143 367 -142
rect 653 -143 654 -142
rect 702 -143 703 -142
rect 737 -143 738 -142
rect 352 -145 353 -144
rect 702 -145 703 -144
rect 730 -145 731 -144
rect 786 -145 787 -144
rect 387 -147 388 -146
rect 436 -147 437 -146
rect 478 -147 479 -146
rect 569 -147 570 -146
rect 695 -147 696 -146
rect 730 -147 731 -146
rect 401 -149 402 -148
rect 527 -149 528 -148
rect 359 -151 360 -150
rect 527 -151 528 -150
rect 359 -153 360 -152
rect 772 -153 773 -152
rect 436 -155 437 -154
rect 541 -155 542 -154
rect 492 -157 493 -156
rect 555 -157 556 -156
rect 492 -159 493 -158
rect 506 -159 507 -158
rect 541 -159 542 -158
rect 604 -159 605 -158
rect 499 -161 500 -160
rect 604 -161 605 -160
rect 499 -163 500 -162
rect 887 -163 888 -162
rect 506 -165 507 -164
rect 688 -165 689 -164
rect 51 -176 52 -175
rect 163 -176 164 -175
rect 177 -176 178 -175
rect 506 -176 507 -175
rect 516 -176 517 -175
rect 1157 -176 1158 -175
rect 1220 -176 1221 -175
rect 1227 -176 1228 -175
rect 58 -178 59 -177
rect 261 -178 262 -177
rect 296 -178 297 -177
rect 499 -178 500 -177
rect 530 -178 531 -177
rect 828 -178 829 -177
rect 849 -178 850 -177
rect 884 -178 885 -177
rect 887 -178 888 -177
rect 1087 -178 1088 -177
rect 1097 -178 1098 -177
rect 1150 -178 1151 -177
rect 65 -180 66 -179
rect 450 -180 451 -179
rect 457 -180 458 -179
rect 481 -180 482 -179
rect 544 -180 545 -179
rect 723 -180 724 -179
rect 737 -180 738 -179
rect 1031 -180 1032 -179
rect 1038 -180 1039 -179
rect 1108 -180 1109 -179
rect 1118 -180 1119 -179
rect 1195 -180 1196 -179
rect 72 -182 73 -181
rect 156 -182 157 -181
rect 163 -182 164 -181
rect 432 -182 433 -181
rect 443 -182 444 -181
rect 499 -182 500 -181
rect 541 -182 542 -181
rect 737 -182 738 -181
rect 772 -182 773 -181
rect 1024 -182 1025 -181
rect 1129 -182 1130 -181
rect 1171 -182 1172 -181
rect 79 -184 80 -183
rect 464 -184 465 -183
rect 474 -184 475 -183
rect 1283 -184 1284 -183
rect 86 -186 87 -185
rect 240 -186 241 -185
rect 261 -186 262 -185
rect 352 -186 353 -185
rect 366 -186 367 -185
rect 495 -186 496 -185
rect 548 -186 549 -185
rect 723 -186 724 -185
rect 772 -186 773 -185
rect 821 -186 822 -185
rect 863 -186 864 -185
rect 1038 -186 1039 -185
rect 1125 -186 1126 -185
rect 1129 -186 1130 -185
rect 1136 -186 1137 -185
rect 1255 -186 1256 -185
rect 93 -188 94 -187
rect 100 -188 101 -187
rect 107 -188 108 -187
rect 114 -188 115 -187
rect 121 -188 122 -187
rect 513 -188 514 -187
rect 548 -188 549 -187
rect 614 -188 615 -187
rect 653 -188 654 -187
rect 835 -188 836 -187
rect 870 -188 871 -187
rect 1052 -188 1053 -187
rect 93 -190 94 -189
rect 170 -190 171 -189
rect 177 -190 178 -189
rect 191 -190 192 -189
rect 212 -190 213 -189
rect 303 -190 304 -189
rect 317 -190 318 -189
rect 352 -190 353 -189
rect 380 -190 381 -189
rect 509 -190 510 -189
rect 614 -190 615 -189
rect 758 -190 759 -189
rect 789 -190 790 -189
rect 842 -190 843 -189
rect 877 -190 878 -189
rect 891 -190 892 -189
rect 905 -190 906 -189
rect 1017 -190 1018 -189
rect 117 -192 118 -191
rect 170 -192 171 -191
rect 184 -192 185 -191
rect 201 -192 202 -191
rect 219 -192 220 -191
rect 359 -192 360 -191
rect 380 -192 381 -191
rect 527 -192 528 -191
rect 569 -192 570 -191
rect 842 -192 843 -191
rect 880 -192 881 -191
rect 898 -192 899 -191
rect 905 -192 906 -191
rect 968 -192 969 -191
rect 975 -192 976 -191
rect 1080 -192 1081 -191
rect 128 -194 129 -193
rect 268 -194 269 -193
rect 292 -194 293 -193
rect 366 -194 367 -193
rect 383 -194 384 -193
rect 513 -194 514 -193
rect 656 -194 657 -193
rect 975 -194 976 -193
rect 996 -194 997 -193
rect 1101 -194 1102 -193
rect 142 -196 143 -195
rect 215 -196 216 -195
rect 219 -196 220 -195
rect 282 -196 283 -195
rect 296 -196 297 -195
rect 583 -196 584 -195
rect 688 -196 689 -195
rect 835 -196 836 -195
rect 898 -196 899 -195
rect 940 -196 941 -195
rect 954 -196 955 -195
rect 1073 -196 1074 -195
rect 142 -198 143 -197
rect 149 -198 150 -197
rect 156 -198 157 -197
rect 593 -198 594 -197
rect 688 -198 689 -197
rect 856 -198 857 -197
rect 933 -198 934 -197
rect 1143 -198 1144 -197
rect 149 -200 150 -199
rect 408 -200 409 -199
rect 415 -200 416 -199
rect 446 -200 447 -199
rect 457 -200 458 -199
rect 632 -200 633 -199
rect 681 -200 682 -199
rect 856 -200 857 -199
rect 940 -200 941 -199
rect 961 -200 962 -199
rect 968 -200 969 -199
rect 982 -200 983 -199
rect 996 -200 997 -199
rect 1059 -200 1060 -199
rect 184 -202 185 -201
rect 198 -202 199 -201
rect 254 -202 255 -201
rect 282 -202 283 -201
rect 303 -202 304 -201
rect 520 -202 521 -201
rect 632 -202 633 -201
rect 674 -202 675 -201
rect 681 -202 682 -201
rect 919 -202 920 -201
rect 999 -202 1000 -201
rect 1066 -202 1067 -201
rect 191 -204 192 -203
rect 205 -204 206 -203
rect 254 -204 255 -203
rect 324 -204 325 -203
rect 345 -204 346 -203
rect 408 -204 409 -203
rect 429 -204 430 -203
rect 534 -204 535 -203
rect 562 -204 563 -203
rect 674 -204 675 -203
rect 698 -204 699 -203
rect 1003 -204 1004 -203
rect 1010 -204 1011 -203
rect 1136 -204 1137 -203
rect 268 -206 269 -205
rect 387 -206 388 -205
rect 394 -206 395 -205
rect 450 -206 451 -205
rect 492 -206 493 -205
rect 583 -206 584 -205
rect 709 -206 710 -205
rect 863 -206 864 -205
rect 947 -206 948 -205
rect 1010 -206 1011 -205
rect 275 -208 276 -207
rect 415 -208 416 -207
rect 509 -208 510 -207
rect 653 -208 654 -207
rect 716 -208 717 -207
rect 1045 -208 1046 -207
rect 208 -210 209 -209
rect 275 -210 276 -209
rect 289 -210 290 -209
rect 324 -210 325 -209
rect 345 -210 346 -209
rect 362 -210 363 -209
rect 387 -210 388 -209
rect 523 -210 524 -209
rect 534 -210 535 -209
rect 730 -210 731 -209
rect 744 -210 745 -209
rect 870 -210 871 -209
rect 243 -212 244 -211
rect 289 -212 290 -211
rect 310 -212 311 -211
rect 394 -212 395 -211
rect 422 -212 423 -211
rect 730 -212 731 -211
rect 751 -212 752 -211
rect 982 -212 983 -211
rect 135 -214 136 -213
rect 243 -214 244 -213
rect 310 -214 311 -213
rect 331 -214 332 -213
rect 359 -214 360 -213
rect 831 -214 832 -213
rect 135 -216 136 -215
rect 233 -216 234 -215
rect 317 -216 318 -215
rect 338 -216 339 -215
rect 422 -216 423 -215
rect 569 -216 570 -215
rect 604 -216 605 -215
rect 709 -216 710 -215
rect 765 -216 766 -215
rect 891 -216 892 -215
rect 233 -218 234 -217
rect 758 -218 759 -217
rect 765 -218 766 -217
rect 926 -218 927 -217
rect 247 -220 248 -219
rect 338 -220 339 -219
rect 471 -220 472 -219
rect 926 -220 927 -219
rect 247 -222 248 -221
rect 544 -222 545 -221
rect 562 -222 563 -221
rect 590 -222 591 -221
rect 604 -222 605 -221
rect 625 -222 626 -221
rect 660 -222 661 -221
rect 751 -222 752 -221
rect 768 -222 769 -221
rect 919 -222 920 -221
rect 331 -224 332 -223
rect 579 -224 580 -223
rect 702 -224 703 -223
rect 744 -224 745 -223
rect 779 -224 780 -223
rect 933 -224 934 -223
rect 436 -226 437 -225
rect 471 -226 472 -225
rect 478 -226 479 -225
rect 590 -226 591 -225
rect 611 -226 612 -225
rect 779 -226 780 -225
rect 793 -226 794 -225
rect 961 -226 962 -225
rect 236 -228 237 -227
rect 436 -228 437 -227
rect 520 -228 521 -227
rect 576 -228 577 -227
rect 611 -228 612 -227
rect 947 -228 948 -227
rect 226 -230 227 -229
rect 236 -230 237 -229
rect 541 -230 542 -229
rect 625 -230 626 -229
rect 793 -230 794 -229
rect 912 -230 913 -229
rect 226 -232 227 -231
rect 373 -232 374 -231
rect 555 -232 556 -231
rect 660 -232 661 -231
rect 719 -232 720 -231
rect 912 -232 913 -231
rect 373 -234 374 -233
rect 443 -234 444 -233
rect 555 -234 556 -233
rect 695 -234 696 -233
rect 796 -234 797 -233
rect 1164 -234 1165 -233
rect 572 -236 573 -235
rect 695 -236 696 -235
rect 800 -236 801 -235
rect 849 -236 850 -235
rect 502 -238 503 -237
rect 800 -238 801 -237
rect 807 -238 808 -237
rect 989 -238 990 -237
rect 618 -240 619 -239
rect 702 -240 703 -239
rect 786 -240 787 -239
rect 807 -240 808 -239
rect 814 -240 815 -239
rect 954 -240 955 -239
rect 460 -242 461 -241
rect 618 -242 619 -241
rect 597 -244 598 -243
rect 814 -244 815 -243
rect 597 -246 598 -245
rect 667 -246 668 -245
rect 485 -248 486 -247
rect 667 -248 668 -247
rect 401 -250 402 -249
rect 485 -250 486 -249
rect 401 -252 402 -251
rect 467 -252 468 -251
rect 44 -263 45 -262
rect 296 -263 297 -262
rect 383 -263 384 -262
rect 541 -263 542 -262
rect 548 -263 549 -262
rect 590 -263 591 -262
rect 593 -263 594 -262
rect 947 -263 948 -262
rect 989 -263 990 -262
rect 1381 -263 1382 -262
rect 51 -265 52 -264
rect 236 -265 237 -264
rect 285 -265 286 -264
rect 1150 -265 1151 -264
rect 1164 -265 1165 -264
rect 1346 -265 1347 -264
rect 51 -267 52 -266
rect 429 -267 430 -266
rect 460 -267 461 -266
rect 667 -267 668 -266
rect 681 -267 682 -266
rect 947 -267 948 -266
rect 996 -267 997 -266
rect 1157 -267 1158 -266
rect 1202 -267 1203 -266
rect 1353 -267 1354 -266
rect 58 -269 59 -268
rect 341 -269 342 -268
rect 415 -269 416 -268
rect 464 -269 465 -268
rect 471 -269 472 -268
rect 751 -269 752 -268
rect 772 -269 773 -268
rect 821 -269 822 -268
rect 828 -269 829 -268
rect 1213 -269 1214 -268
rect 1255 -269 1256 -268
rect 1374 -269 1375 -268
rect 61 -271 62 -270
rect 72 -271 73 -270
rect 86 -271 87 -270
rect 471 -271 472 -270
rect 474 -271 475 -270
rect 835 -271 836 -270
rect 842 -271 843 -270
rect 1290 -271 1291 -270
rect 72 -273 73 -272
rect 93 -273 94 -272
rect 96 -273 97 -272
rect 121 -273 122 -272
rect 142 -273 143 -272
rect 415 -273 416 -272
rect 474 -273 475 -272
rect 1325 -273 1326 -272
rect 65 -275 66 -274
rect 142 -275 143 -274
rect 156 -275 157 -274
rect 233 -275 234 -274
rect 338 -275 339 -274
rect 429 -275 430 -274
rect 506 -275 507 -274
rect 1234 -275 1235 -274
rect 1283 -275 1284 -274
rect 1591 -275 1592 -274
rect 65 -277 66 -276
rect 453 -277 454 -276
rect 509 -277 510 -276
rect 856 -277 857 -276
rect 863 -277 864 -276
rect 1339 -277 1340 -276
rect 86 -279 87 -278
rect 138 -279 139 -278
rect 163 -279 164 -278
rect 467 -279 468 -278
rect 513 -279 514 -278
rect 1388 -279 1389 -278
rect 107 -281 108 -280
rect 296 -281 297 -280
rect 387 -281 388 -280
rect 513 -281 514 -280
rect 527 -281 528 -280
rect 1360 -281 1361 -280
rect 107 -283 108 -282
rect 457 -283 458 -282
rect 527 -283 528 -282
rect 583 -283 584 -282
rect 614 -283 615 -282
rect 982 -283 983 -282
rect 1024 -283 1025 -282
rect 1206 -283 1207 -282
rect 93 -285 94 -284
rect 457 -285 458 -284
rect 499 -285 500 -284
rect 583 -285 584 -284
rect 632 -285 633 -284
rect 835 -285 836 -284
rect 863 -285 864 -284
rect 1094 -285 1095 -284
rect 1101 -285 1102 -284
rect 1367 -285 1368 -284
rect 121 -287 122 -286
rect 156 -287 157 -286
rect 163 -287 164 -286
rect 205 -287 206 -286
rect 215 -287 216 -286
rect 1262 -287 1263 -286
rect 170 -289 171 -288
rect 282 -289 283 -288
rect 352 -289 353 -288
rect 387 -289 388 -288
rect 450 -289 451 -288
rect 506 -289 507 -288
rect 509 -289 510 -288
rect 632 -289 633 -288
rect 667 -289 668 -288
rect 1276 -289 1277 -288
rect 198 -291 199 -290
rect 548 -291 549 -290
rect 576 -291 577 -290
rect 828 -291 829 -290
rect 891 -291 892 -290
rect 894 -291 895 -290
rect 905 -291 906 -290
rect 989 -291 990 -290
rect 1038 -291 1039 -290
rect 1283 -291 1284 -290
rect 135 -293 136 -292
rect 576 -293 577 -292
rect 579 -293 580 -292
rect 639 -293 640 -292
rect 681 -293 682 -292
rect 716 -293 717 -292
rect 723 -293 724 -292
rect 842 -293 843 -292
rect 891 -293 892 -292
rect 898 -293 899 -292
rect 912 -293 913 -292
rect 1241 -293 1242 -292
rect 201 -295 202 -294
rect 380 -295 381 -294
rect 408 -295 409 -294
rect 450 -295 451 -294
rect 478 -295 479 -294
rect 639 -295 640 -294
rect 688 -295 689 -294
rect 821 -295 822 -294
rect 894 -295 895 -294
rect 898 -295 899 -294
rect 933 -295 934 -294
rect 1094 -295 1095 -294
rect 1101 -295 1102 -294
rect 1143 -295 1144 -294
rect 1171 -295 1172 -294
rect 1255 -295 1256 -294
rect 114 -297 115 -296
rect 933 -297 934 -296
rect 1045 -297 1046 -296
rect 1297 -297 1298 -296
rect 205 -299 206 -298
rect 530 -299 531 -298
rect 544 -299 545 -298
rect 716 -299 717 -298
rect 744 -299 745 -298
rect 982 -299 983 -298
rect 1052 -299 1053 -298
rect 1304 -299 1305 -298
rect 282 -301 283 -300
rect 345 -301 346 -300
rect 359 -301 360 -300
rect 478 -301 479 -300
rect 499 -301 500 -300
rect 1395 -301 1396 -300
rect 275 -303 276 -302
rect 345 -303 346 -302
rect 359 -303 360 -302
rect 373 -303 374 -302
rect 443 -303 444 -302
rect 1171 -303 1172 -302
rect 198 -305 199 -304
rect 443 -305 444 -304
rect 611 -305 612 -304
rect 1038 -305 1039 -304
rect 1059 -305 1060 -304
rect 1150 -305 1151 -304
rect 317 -307 318 -306
rect 352 -307 353 -306
rect 373 -307 374 -306
rect 422 -307 423 -306
rect 611 -307 612 -306
rect 1031 -307 1032 -306
rect 1073 -307 1074 -306
rect 1332 -307 1333 -306
rect 58 -309 59 -308
rect 1031 -309 1032 -308
rect 1073 -309 1074 -308
rect 1097 -309 1098 -308
rect 1108 -309 1109 -308
rect 1318 -309 1319 -308
rect 324 -311 325 -310
rect 408 -311 409 -310
rect 422 -311 423 -310
rect 555 -311 556 -310
rect 614 -311 615 -310
rect 723 -311 724 -310
rect 747 -311 748 -310
rect 1003 -311 1004 -310
rect 1017 -311 1018 -310
rect 1108 -311 1109 -310
rect 1115 -311 1116 -310
rect 1129 -311 1130 -310
rect 1136 -311 1137 -310
rect 1311 -311 1312 -310
rect 173 -313 174 -312
rect 1115 -313 1116 -312
rect 1118 -313 1119 -312
rect 1248 -313 1249 -312
rect 324 -315 325 -314
rect 733 -315 734 -314
rect 751 -315 752 -314
rect 1185 -315 1186 -314
rect 492 -317 493 -316
rect 1129 -317 1130 -316
rect 226 -319 227 -318
rect 492 -319 493 -318
rect 555 -319 556 -318
rect 793 -319 794 -318
rect 800 -319 801 -318
rect 905 -319 906 -318
rect 968 -319 969 -318
rect 1059 -319 1060 -318
rect 1066 -319 1067 -318
rect 1136 -319 1137 -318
rect 149 -321 150 -320
rect 226 -321 227 -320
rect 495 -321 496 -320
rect 800 -321 801 -320
rect 814 -321 815 -320
rect 1024 -321 1025 -320
rect 1080 -321 1081 -320
rect 1164 -321 1165 -320
rect 149 -323 150 -322
rect 243 -323 244 -322
rect 618 -323 619 -322
rect 688 -323 689 -322
rect 695 -323 696 -322
rect 912 -323 913 -322
rect 919 -323 920 -322
rect 968 -323 969 -322
rect 975 -323 976 -322
rect 1045 -323 1046 -322
rect 1087 -323 1088 -322
rect 1220 -323 1221 -322
rect 607 -325 608 -324
rect 618 -325 619 -324
rect 625 -325 626 -324
rect 695 -325 696 -324
rect 705 -325 706 -324
rect 1178 -325 1179 -324
rect 520 -327 521 -326
rect 625 -327 626 -326
rect 670 -327 671 -326
rect 1052 -327 1053 -326
rect 1122 -327 1123 -326
rect 1192 -327 1193 -326
rect 520 -329 521 -328
rect 534 -329 535 -328
rect 674 -329 675 -328
rect 793 -329 794 -328
rect 870 -329 871 -328
rect 1003 -329 1004 -328
rect 366 -331 367 -330
rect 534 -331 535 -330
rect 562 -331 563 -330
rect 870 -331 871 -330
rect 926 -331 927 -330
rect 1087 -331 1088 -330
rect 191 -333 192 -332
rect 562 -333 563 -332
rect 653 -333 654 -332
rect 674 -333 675 -332
rect 709 -333 710 -332
rect 814 -333 815 -332
rect 884 -333 885 -332
rect 926 -333 927 -332
rect 961 -333 962 -332
rect 1122 -333 1123 -332
rect 79 -335 80 -334
rect 709 -335 710 -334
rect 712 -335 713 -334
rect 1269 -335 1270 -334
rect 79 -337 80 -336
rect 331 -337 332 -336
rect 439 -337 440 -336
rect 653 -337 654 -336
rect 730 -337 731 -336
rect 919 -337 920 -336
rect 975 -337 976 -336
rect 1010 -337 1011 -336
rect 177 -339 178 -338
rect 191 -339 192 -338
rect 254 -339 255 -338
rect 366 -339 367 -338
rect 730 -339 731 -338
rect 1017 -339 1018 -338
rect 177 -341 178 -340
rect 247 -341 248 -340
rect 331 -341 332 -340
rect 572 -341 573 -340
rect 754 -341 755 -340
rect 884 -341 885 -340
rect 999 -341 1000 -340
rect 1080 -341 1081 -340
rect 208 -343 209 -342
rect 254 -343 255 -342
rect 758 -343 759 -342
rect 1066 -343 1067 -342
rect 646 -345 647 -344
rect 758 -345 759 -344
rect 779 -345 780 -344
rect 856 -345 857 -344
rect 877 -345 878 -344
rect 961 -345 962 -344
rect 194 -347 195 -346
rect 646 -347 647 -346
rect 660 -347 661 -346
rect 779 -347 780 -346
rect 786 -347 787 -346
rect 1143 -347 1144 -346
rect 117 -349 118 -348
rect 786 -349 787 -348
rect 789 -349 790 -348
rect 954 -349 955 -348
rect 117 -351 118 -350
rect 240 -351 241 -350
rect 569 -351 570 -350
rect 877 -351 878 -350
rect 940 -351 941 -350
rect 954 -351 955 -350
rect 569 -353 570 -352
rect 1157 -353 1158 -352
rect 604 -355 605 -354
rect 660 -355 661 -354
rect 737 -355 738 -354
rect 940 -355 941 -354
rect 485 -357 486 -356
rect 737 -357 738 -356
rect 849 -357 850 -356
rect 1010 -357 1011 -356
rect 401 -359 402 -358
rect 485 -359 486 -358
rect 597 -359 598 -358
rect 604 -359 605 -358
rect 765 -359 766 -358
rect 849 -359 850 -358
rect 289 -361 290 -360
rect 597 -361 598 -360
rect 702 -361 703 -360
rect 765 -361 766 -360
rect 275 -363 276 -362
rect 702 -363 703 -362
rect 289 -365 290 -364
rect 303 -365 304 -364
rect 338 -365 339 -364
rect 401 -365 402 -364
rect 303 -367 304 -366
rect 394 -367 395 -366
rect 268 -369 269 -368
rect 394 -369 395 -368
rect 268 -371 269 -370
rect 310 -371 311 -370
rect 261 -373 262 -372
rect 310 -373 311 -372
rect 219 -375 220 -374
rect 261 -375 262 -374
rect 219 -377 220 -376
rect 436 -377 437 -376
rect 128 -379 129 -378
rect 436 -379 437 -378
rect 100 -381 101 -380
rect 128 -381 129 -380
rect 100 -383 101 -382
rect 411 -383 412 -382
rect 23 -394 24 -393
rect 233 -394 234 -393
rect 247 -394 248 -393
rect 453 -394 454 -393
rect 506 -394 507 -393
rect 1290 -394 1291 -393
rect 1297 -394 1298 -393
rect 1444 -394 1445 -393
rect 1591 -394 1592 -393
rect 1710 -394 1711 -393
rect 30 -396 31 -395
rect 443 -396 444 -395
rect 450 -396 451 -395
rect 1486 -396 1487 -395
rect 37 -398 38 -397
rect 100 -398 101 -397
rect 107 -398 108 -397
rect 362 -398 363 -397
rect 408 -398 409 -397
rect 583 -398 584 -397
rect 597 -398 598 -397
rect 730 -398 731 -397
rect 1143 -398 1144 -397
rect 1451 -398 1452 -397
rect 58 -400 59 -399
rect 275 -400 276 -399
rect 317 -400 318 -399
rect 387 -400 388 -399
rect 429 -400 430 -399
rect 523 -400 524 -399
rect 530 -400 531 -399
rect 744 -400 745 -399
rect 1031 -400 1032 -399
rect 1143 -400 1144 -399
rect 1164 -400 1165 -399
rect 1465 -400 1466 -399
rect 82 -402 83 -401
rect 576 -402 577 -401
rect 607 -402 608 -401
rect 1339 -402 1340 -401
rect 1346 -402 1347 -401
rect 1500 -402 1501 -401
rect 86 -404 87 -403
rect 408 -404 409 -403
rect 429 -404 430 -403
rect 758 -404 759 -403
rect 933 -404 934 -403
rect 1031 -404 1032 -403
rect 1052 -404 1053 -403
rect 1164 -404 1165 -403
rect 1171 -404 1172 -403
rect 1339 -404 1340 -403
rect 1353 -404 1354 -403
rect 1479 -404 1480 -403
rect 86 -406 87 -405
rect 583 -406 584 -405
rect 611 -406 612 -405
rect 793 -406 794 -405
rect 807 -406 808 -405
rect 1052 -406 1053 -405
rect 1066 -406 1067 -405
rect 1171 -406 1172 -405
rect 1178 -406 1179 -405
rect 1297 -406 1298 -405
rect 1304 -406 1305 -405
rect 1409 -406 1410 -405
rect 89 -408 90 -407
rect 128 -408 129 -407
rect 135 -408 136 -407
rect 933 -408 934 -407
rect 982 -408 983 -407
rect 1066 -408 1067 -407
rect 1073 -408 1074 -407
rect 1178 -408 1179 -407
rect 1220 -408 1221 -407
rect 1493 -408 1494 -407
rect 93 -410 94 -409
rect 103 -410 104 -409
rect 110 -410 111 -409
rect 919 -410 920 -409
rect 982 -410 983 -409
rect 1080 -410 1081 -409
rect 1094 -410 1095 -409
rect 1220 -410 1221 -409
rect 1227 -410 1228 -409
rect 1290 -410 1291 -409
rect 1311 -410 1312 -409
rect 1416 -410 1417 -409
rect 96 -412 97 -411
rect 681 -412 682 -411
rect 695 -412 696 -411
rect 793 -412 794 -411
rect 905 -412 906 -411
rect 1094 -412 1095 -411
rect 1115 -412 1116 -411
rect 1227 -412 1228 -411
rect 1269 -412 1270 -411
rect 1423 -412 1424 -411
rect 100 -414 101 -413
rect 1248 -414 1249 -413
rect 1269 -414 1270 -413
rect 1398 -414 1399 -413
rect 114 -416 115 -415
rect 261 -416 262 -415
rect 268 -416 269 -415
rect 285 -416 286 -415
rect 324 -416 325 -415
rect 474 -416 475 -415
rect 481 -416 482 -415
rect 1073 -416 1074 -415
rect 1136 -416 1137 -415
rect 1346 -416 1347 -415
rect 1353 -416 1354 -415
rect 1524 -416 1525 -415
rect 65 -418 66 -417
rect 268 -418 269 -417
rect 324 -418 325 -417
rect 569 -418 570 -417
rect 576 -418 577 -417
rect 688 -418 689 -417
rect 695 -418 696 -417
rect 737 -418 738 -417
rect 747 -418 748 -417
rect 1311 -418 1312 -417
rect 1318 -418 1319 -417
rect 1430 -418 1431 -417
rect 65 -420 66 -419
rect 359 -420 360 -419
rect 366 -420 367 -419
rect 387 -420 388 -419
rect 436 -420 437 -419
rect 527 -420 528 -419
rect 534 -420 535 -419
rect 593 -420 594 -419
rect 618 -420 619 -419
rect 730 -420 731 -419
rect 733 -420 734 -419
rect 1304 -420 1305 -419
rect 1325 -420 1326 -419
rect 1472 -420 1473 -419
rect 79 -422 80 -421
rect 366 -422 367 -421
rect 401 -422 402 -421
rect 436 -422 437 -421
rect 439 -422 440 -421
rect 744 -422 745 -421
rect 758 -422 759 -421
rect 842 -422 843 -421
rect 884 -422 885 -421
rect 1325 -422 1326 -421
rect 1332 -422 1333 -421
rect 1458 -422 1459 -421
rect 79 -424 80 -423
rect 359 -424 360 -423
rect 474 -424 475 -423
rect 1136 -424 1137 -423
rect 1192 -424 1193 -423
rect 1332 -424 1333 -423
rect 1374 -424 1375 -423
rect 1507 -424 1508 -423
rect 121 -426 122 -425
rect 299 -426 300 -425
rect 331 -426 332 -425
rect 401 -426 402 -425
rect 485 -426 486 -425
rect 506 -426 507 -425
rect 534 -426 535 -425
rect 1318 -426 1319 -425
rect 121 -428 122 -427
rect 499 -428 500 -427
rect 541 -428 542 -427
rect 569 -428 570 -427
rect 639 -428 640 -427
rect 751 -428 752 -427
rect 842 -428 843 -427
rect 1122 -428 1123 -427
rect 1206 -428 1207 -427
rect 1374 -428 1375 -427
rect 124 -430 125 -429
rect 1129 -430 1130 -429
rect 1276 -430 1277 -429
rect 1402 -430 1403 -429
rect 128 -432 129 -431
rect 135 -432 136 -431
rect 163 -432 164 -431
rect 166 -432 167 -431
rect 170 -432 171 -431
rect 418 -432 419 -431
rect 464 -432 465 -431
rect 485 -432 486 -431
rect 492 -432 493 -431
rect 541 -432 542 -431
rect 653 -432 654 -431
rect 751 -432 752 -431
rect 856 -432 857 -431
rect 884 -432 885 -431
rect 919 -432 920 -431
rect 926 -432 927 -431
rect 954 -432 955 -431
rect 1248 -432 1249 -431
rect 1283 -432 1284 -431
rect 1437 -432 1438 -431
rect 51 -434 52 -433
rect 653 -434 654 -433
rect 660 -434 661 -433
rect 667 -434 668 -433
rect 670 -434 671 -433
rect 1388 -434 1389 -433
rect 51 -436 52 -435
rect 303 -436 304 -435
rect 331 -436 332 -435
rect 471 -436 472 -435
rect 478 -436 479 -435
rect 499 -436 500 -435
rect 509 -436 510 -435
rect 856 -436 857 -435
rect 898 -436 899 -435
rect 954 -436 955 -435
rect 968 -436 969 -435
rect 1129 -436 1130 -435
rect 1255 -436 1256 -435
rect 1388 -436 1389 -435
rect 163 -438 164 -437
rect 289 -438 290 -437
rect 303 -438 304 -437
rect 394 -438 395 -437
rect 443 -438 444 -437
rect 492 -438 493 -437
rect 604 -438 605 -437
rect 926 -438 927 -437
rect 989 -438 990 -437
rect 1115 -438 1116 -437
rect 1150 -438 1151 -437
rect 1255 -438 1256 -437
rect 1283 -438 1284 -437
rect 1367 -438 1368 -437
rect 166 -440 167 -439
rect 289 -440 290 -439
rect 352 -440 353 -439
rect 527 -440 528 -439
rect 562 -440 563 -439
rect 604 -440 605 -439
rect 625 -440 626 -439
rect 660 -440 661 -439
rect 674 -440 675 -439
rect 681 -440 682 -439
rect 702 -440 703 -439
rect 1381 -440 1382 -439
rect 26 -442 27 -441
rect 562 -442 563 -441
rect 632 -442 633 -441
rect 674 -442 675 -441
rect 712 -442 713 -441
rect 1276 -442 1277 -441
rect 142 -444 143 -443
rect 625 -444 626 -443
rect 632 -444 633 -443
rect 1514 -444 1515 -443
rect 142 -446 143 -445
rect 296 -446 297 -445
rect 352 -446 353 -445
rect 555 -446 556 -445
rect 716 -446 717 -445
rect 807 -446 808 -445
rect 863 -446 864 -445
rect 968 -446 969 -445
rect 1010 -446 1011 -445
rect 1122 -446 1123 -445
rect 1213 -446 1214 -445
rect 1367 -446 1368 -445
rect 117 -448 118 -447
rect 716 -448 717 -447
rect 800 -448 801 -447
rect 863 -448 864 -447
rect 877 -448 878 -447
rect 989 -448 990 -447
rect 1017 -448 1018 -447
rect 1206 -448 1207 -447
rect 1241 -448 1242 -447
rect 1381 -448 1382 -447
rect 170 -450 171 -449
rect 422 -450 423 -449
rect 464 -450 465 -449
rect 590 -450 591 -449
rect 649 -450 650 -449
rect 877 -450 878 -449
rect 891 -450 892 -449
rect 1010 -450 1011 -449
rect 1017 -450 1018 -449
rect 1101 -450 1102 -449
rect 1108 -450 1109 -449
rect 1213 -450 1214 -449
rect 180 -452 181 -451
rect 702 -452 703 -451
rect 709 -452 710 -451
rect 1241 -452 1242 -451
rect 187 -454 188 -453
rect 422 -454 423 -453
rect 478 -454 479 -453
rect 1360 -454 1361 -453
rect 194 -456 195 -455
rect 611 -456 612 -455
rect 779 -456 780 -455
rect 891 -456 892 -455
rect 898 -456 899 -455
rect 1528 -456 1529 -455
rect 198 -458 199 -457
rect 905 -458 906 -457
rect 996 -458 997 -457
rect 1108 -458 1109 -457
rect 1199 -458 1200 -457
rect 1360 -458 1361 -457
rect 184 -460 185 -459
rect 198 -460 199 -459
rect 205 -460 206 -459
rect 261 -460 262 -459
rect 282 -460 283 -459
rect 737 -460 738 -459
rect 870 -460 871 -459
rect 996 -460 997 -459
rect 1003 -460 1004 -459
rect 1101 -460 1102 -459
rect 1185 -460 1186 -459
rect 1199 -460 1200 -459
rect 205 -462 206 -461
rect 513 -462 514 -461
rect 520 -462 521 -461
rect 555 -462 556 -461
rect 590 -462 591 -461
rect 821 -462 822 -461
rect 870 -462 871 -461
rect 947 -462 948 -461
rect 1003 -462 1004 -461
rect 1395 -462 1396 -461
rect 44 -464 45 -463
rect 821 -464 822 -463
rect 849 -464 850 -463
rect 947 -464 948 -463
rect 1038 -464 1039 -463
rect 1150 -464 1151 -463
rect 1262 -464 1263 -463
rect 1395 -464 1396 -463
rect 44 -466 45 -465
rect 226 -466 227 -465
rect 254 -466 255 -465
rect 275 -466 276 -465
rect 282 -466 283 -465
rect 495 -466 496 -465
rect 520 -466 521 -465
rect 1024 -466 1025 -465
rect 1045 -466 1046 -465
rect 1080 -466 1081 -465
rect 1087 -466 1088 -465
rect 1185 -466 1186 -465
rect 191 -468 192 -467
rect 226 -468 227 -467
rect 254 -468 255 -467
rect 614 -468 615 -467
rect 635 -468 636 -467
rect 1262 -468 1263 -467
rect 191 -470 192 -469
rect 513 -470 514 -469
rect 723 -470 724 -469
rect 779 -470 780 -469
rect 786 -470 787 -469
rect 849 -470 850 -469
rect 940 -470 941 -469
rect 1045 -470 1046 -469
rect 1087 -470 1088 -469
rect 1157 -470 1158 -469
rect 138 -472 139 -471
rect 786 -472 787 -471
rect 961 -472 962 -471
rect 1038 -472 1039 -471
rect 1059 -472 1060 -471
rect 1157 -472 1158 -471
rect 138 -474 139 -473
rect 618 -474 619 -473
rect 723 -474 724 -473
rect 814 -474 815 -473
rect 828 -474 829 -473
rect 1059 -474 1060 -473
rect 215 -476 216 -475
rect 688 -476 689 -475
rect 828 -476 829 -475
rect 1234 -476 1235 -475
rect 107 -478 108 -477
rect 1234 -478 1235 -477
rect 219 -480 220 -479
rect 639 -480 640 -479
rect 835 -480 836 -479
rect 961 -480 962 -479
rect 975 -480 976 -479
rect 1024 -480 1025 -479
rect 338 -482 339 -481
rect 814 -482 815 -481
rect 912 -482 913 -481
rect 975 -482 976 -481
rect 338 -484 339 -483
rect 345 -484 346 -483
rect 380 -484 381 -483
rect 394 -484 395 -483
rect 548 -484 549 -483
rect 912 -484 913 -483
rect 149 -486 150 -485
rect 380 -486 381 -485
rect 457 -486 458 -485
rect 548 -486 549 -485
rect 597 -486 598 -485
rect 940 -486 941 -485
rect 149 -488 150 -487
rect 177 -488 178 -487
rect 310 -488 311 -487
rect 345 -488 346 -487
rect 457 -488 458 -487
rect 646 -488 647 -487
rect 765 -488 766 -487
rect 835 -488 836 -487
rect 177 -490 178 -489
rect 212 -490 213 -489
rect 310 -490 311 -489
rect 415 -490 416 -489
rect 646 -490 647 -489
rect 800 -490 801 -489
rect 212 -492 213 -491
rect 240 -492 241 -491
rect 373 -492 374 -491
rect 765 -492 766 -491
rect 219 -494 220 -493
rect 240 -494 241 -493
rect 320 -494 321 -493
rect 373 -494 374 -493
rect 9 -505 10 -504
rect 282 -505 283 -504
rect 317 -505 318 -504
rect 415 -505 416 -504
rect 450 -505 451 -504
rect 863 -505 864 -504
rect 873 -505 874 -504
rect 982 -505 983 -504
rect 1136 -505 1137 -504
rect 1192 -505 1193 -504
rect 1269 -505 1270 -504
rect 1272 -505 1273 -504
rect 1468 -505 1469 -504
rect 1556 -505 1557 -504
rect 1710 -505 1711 -504
rect 1759 -505 1760 -504
rect 23 -507 24 -506
rect 51 -507 52 -506
rect 58 -507 59 -506
rect 100 -507 101 -506
rect 103 -507 104 -506
rect 324 -507 325 -506
rect 359 -507 360 -506
rect 408 -507 409 -506
rect 450 -507 451 -506
rect 569 -507 570 -506
rect 583 -507 584 -506
rect 607 -507 608 -506
rect 618 -507 619 -506
rect 982 -507 983 -506
rect 1129 -507 1130 -506
rect 1136 -507 1137 -506
rect 1269 -507 1270 -506
rect 1304 -507 1305 -506
rect 1486 -507 1487 -506
rect 1521 -507 1522 -506
rect 1528 -507 1529 -506
rect 1766 -507 1767 -506
rect 37 -509 38 -508
rect 184 -509 185 -508
rect 194 -509 195 -508
rect 1164 -509 1165 -508
rect 1500 -509 1501 -508
rect 1503 -509 1504 -508
rect 1514 -509 1515 -508
rect 1738 -509 1739 -508
rect 61 -511 62 -510
rect 1262 -511 1263 -510
rect 1458 -511 1459 -510
rect 1514 -511 1515 -510
rect 79 -513 80 -512
rect 324 -513 325 -512
rect 362 -513 363 -512
rect 751 -513 752 -512
rect 758 -513 759 -512
rect 1360 -513 1361 -512
rect 1451 -513 1452 -512
rect 1458 -513 1459 -512
rect 1500 -513 1501 -512
rect 1507 -513 1508 -512
rect 72 -515 73 -514
rect 79 -515 80 -514
rect 103 -515 104 -514
rect 408 -515 409 -514
rect 453 -515 454 -514
rect 597 -515 598 -514
rect 618 -515 619 -514
rect 1073 -515 1074 -514
rect 1122 -515 1123 -514
rect 1129 -515 1130 -514
rect 1150 -515 1151 -514
rect 1164 -515 1165 -514
rect 1325 -515 1326 -514
rect 1360 -515 1361 -514
rect 1430 -515 1431 -514
rect 1451 -515 1452 -514
rect 72 -517 73 -516
rect 114 -517 115 -516
rect 128 -517 129 -516
rect 219 -517 220 -516
rect 222 -517 223 -516
rect 688 -517 689 -516
rect 709 -517 710 -516
rect 1220 -517 1221 -516
rect 1402 -517 1403 -516
rect 1430 -517 1431 -516
rect 107 -519 108 -518
rect 121 -519 122 -518
rect 128 -519 129 -518
rect 394 -519 395 -518
rect 401 -519 402 -518
rect 474 -519 475 -518
rect 481 -519 482 -518
rect 800 -519 801 -518
rect 824 -519 825 -518
rect 1248 -519 1249 -518
rect 114 -521 115 -520
rect 537 -521 538 -520
rect 548 -521 549 -520
rect 569 -521 570 -520
rect 583 -521 584 -520
rect 961 -521 962 -520
rect 1052 -521 1053 -520
rect 1122 -521 1123 -520
rect 1185 -521 1186 -520
rect 1220 -521 1221 -520
rect 121 -523 122 -522
rect 338 -523 339 -522
rect 341 -523 342 -522
rect 548 -523 549 -522
rect 590 -523 591 -522
rect 828 -523 829 -522
rect 831 -523 832 -522
rect 1150 -523 1151 -522
rect 1199 -523 1200 -522
rect 1325 -523 1326 -522
rect 138 -525 139 -524
rect 1444 -525 1445 -524
rect 152 -527 153 -526
rect 586 -527 587 -526
rect 593 -527 594 -526
rect 1073 -527 1074 -526
rect 1080 -527 1081 -526
rect 1402 -527 1403 -526
rect 1416 -527 1417 -526
rect 1444 -527 1445 -526
rect 156 -529 157 -528
rect 187 -529 188 -528
rect 243 -529 244 -528
rect 359 -529 360 -528
rect 373 -529 374 -528
rect 534 -529 535 -528
rect 593 -529 594 -528
rect 1199 -529 1200 -528
rect 1213 -529 1214 -528
rect 1248 -529 1249 -528
rect 1395 -529 1396 -528
rect 1416 -529 1417 -528
rect 44 -531 45 -530
rect 534 -531 535 -530
rect 597 -531 598 -530
rect 814 -531 815 -530
rect 828 -531 829 -530
rect 835 -531 836 -530
rect 842 -531 843 -530
rect 1262 -531 1263 -530
rect 1367 -531 1368 -530
rect 1395 -531 1396 -530
rect 44 -533 45 -532
rect 901 -533 902 -532
rect 947 -533 948 -532
rect 950 -533 951 -532
rect 961 -533 962 -532
rect 1066 -533 1067 -532
rect 1178 -533 1179 -532
rect 1213 -533 1214 -532
rect 1332 -533 1333 -532
rect 1367 -533 1368 -532
rect 93 -535 94 -534
rect 156 -535 157 -534
rect 177 -535 178 -534
rect 198 -535 199 -534
rect 268 -535 269 -534
rect 296 -535 297 -534
rect 317 -535 318 -534
rect 765 -535 766 -534
rect 779 -535 780 -534
rect 800 -535 801 -534
rect 842 -535 843 -534
rect 1437 -535 1438 -534
rect 93 -537 94 -536
rect 142 -537 143 -536
rect 180 -537 181 -536
rect 205 -537 206 -536
rect 268 -537 269 -536
rect 520 -537 521 -536
rect 530 -537 531 -536
rect 730 -537 731 -536
rect 761 -537 762 -536
rect 1185 -537 1186 -536
rect 1318 -537 1319 -536
rect 1332 -537 1333 -536
rect 1409 -537 1410 -536
rect 1437 -537 1438 -536
rect 65 -539 66 -538
rect 520 -539 521 -538
rect 530 -539 531 -538
rect 646 -539 647 -538
rect 667 -539 668 -538
rect 712 -539 713 -538
rect 716 -539 717 -538
rect 758 -539 759 -538
rect 765 -539 766 -538
rect 1339 -539 1340 -538
rect 1388 -539 1389 -538
rect 1409 -539 1410 -538
rect 65 -541 66 -540
rect 135 -541 136 -540
rect 142 -541 143 -540
rect 457 -541 458 -540
rect 460 -541 461 -540
rect 1423 -541 1424 -540
rect 135 -543 136 -542
rect 149 -543 150 -542
rect 191 -543 192 -542
rect 457 -543 458 -542
rect 464 -543 465 -542
rect 649 -543 650 -542
rect 653 -543 654 -542
rect 667 -543 668 -542
rect 677 -543 678 -542
rect 716 -543 717 -542
rect 723 -543 724 -542
rect 814 -543 815 -542
rect 915 -543 916 -542
rect 1388 -543 1389 -542
rect 149 -545 150 -544
rect 310 -545 311 -544
rect 352 -545 353 -544
rect 653 -545 654 -544
rect 681 -545 682 -544
rect 723 -545 724 -544
rect 730 -545 731 -544
rect 793 -545 794 -544
rect 947 -545 948 -544
rect 989 -545 990 -544
rect 1017 -545 1018 -544
rect 1080 -545 1081 -544
rect 1157 -545 1158 -544
rect 1178 -545 1179 -544
rect 1297 -545 1298 -544
rect 1318 -545 1319 -544
rect 1339 -545 1340 -544
rect 1381 -545 1382 -544
rect 198 -547 199 -546
rect 254 -547 255 -546
rect 275 -547 276 -546
rect 282 -547 283 -546
rect 310 -547 311 -546
rect 506 -547 507 -546
rect 516 -547 517 -546
rect 709 -547 710 -546
rect 779 -547 780 -546
rect 1472 -547 1473 -546
rect 30 -549 31 -548
rect 506 -549 507 -548
rect 516 -549 517 -548
rect 1157 -549 1158 -548
rect 1297 -549 1298 -548
rect 1346 -549 1347 -548
rect 1472 -549 1473 -548
rect 1479 -549 1480 -548
rect 163 -551 164 -550
rect 275 -551 276 -550
rect 366 -551 367 -550
rect 373 -551 374 -550
rect 380 -551 381 -550
rect 401 -551 402 -550
rect 464 -551 465 -550
rect 695 -551 696 -550
rect 786 -551 787 -550
rect 835 -551 836 -550
rect 954 -551 955 -550
rect 1017 -551 1018 -550
rect 1038 -551 1039 -550
rect 1066 -551 1067 -550
rect 1283 -551 1284 -550
rect 1479 -551 1480 -550
rect 163 -553 164 -552
rect 261 -553 262 -552
rect 366 -553 367 -552
rect 485 -553 486 -552
rect 492 -553 493 -552
rect 891 -553 892 -552
rect 919 -553 920 -552
rect 1038 -553 1039 -552
rect 1052 -553 1053 -552
rect 1311 -553 1312 -552
rect 1346 -553 1347 -552
rect 1465 -553 1466 -552
rect 205 -555 206 -554
rect 247 -555 248 -554
rect 254 -555 255 -554
rect 576 -555 577 -554
rect 625 -555 626 -554
rect 852 -555 853 -554
rect 891 -555 892 -554
rect 1535 -555 1536 -554
rect 30 -557 31 -556
rect 247 -557 248 -556
rect 261 -557 262 -556
rect 478 -557 479 -556
rect 485 -557 486 -556
rect 611 -557 612 -556
rect 625 -557 626 -556
rect 737 -557 738 -556
rect 786 -557 787 -556
rect 1003 -557 1004 -556
rect 1241 -557 1242 -556
rect 1283 -557 1284 -556
rect 1290 -557 1291 -556
rect 1311 -557 1312 -556
rect 170 -559 171 -558
rect 611 -559 612 -558
rect 632 -559 633 -558
rect 996 -559 997 -558
rect 1087 -559 1088 -558
rect 1290 -559 1291 -558
rect 170 -561 171 -560
rect 429 -561 430 -560
rect 436 -561 437 -560
rect 478 -561 479 -560
rect 492 -561 493 -560
rect 856 -561 857 -560
rect 919 -561 920 -560
rect 1059 -561 1060 -560
rect 1087 -561 1088 -560
rect 1227 -561 1228 -560
rect 226 -563 227 -562
rect 352 -563 353 -562
rect 387 -563 388 -562
rect 394 -563 395 -562
rect 418 -563 419 -562
rect 1241 -563 1242 -562
rect 226 -565 227 -564
rect 443 -565 444 -564
rect 471 -565 472 -564
rect 562 -565 563 -564
rect 576 -565 577 -564
rect 1108 -565 1109 -564
rect 1195 -565 1196 -564
rect 1227 -565 1228 -564
rect 233 -567 234 -566
rect 443 -567 444 -566
rect 495 -567 496 -566
rect 968 -567 969 -566
rect 1055 -567 1056 -566
rect 1108 -567 1109 -566
rect 303 -569 304 -568
rect 387 -569 388 -568
rect 523 -569 524 -568
rect 1381 -569 1382 -568
rect 240 -571 241 -570
rect 303 -571 304 -570
rect 331 -571 332 -570
rect 436 -571 437 -570
rect 527 -571 528 -570
rect 1423 -571 1424 -570
rect 212 -573 213 -572
rect 331 -573 332 -572
rect 527 -573 528 -572
rect 1276 -573 1277 -572
rect 212 -575 213 -574
rect 422 -575 423 -574
rect 562 -575 563 -574
rect 772 -575 773 -574
rect 793 -575 794 -574
rect 884 -575 885 -574
rect 898 -575 899 -574
rect 1059 -575 1060 -574
rect 1255 -575 1256 -574
rect 1276 -575 1277 -574
rect 240 -577 241 -576
rect 289 -577 290 -576
rect 338 -577 339 -576
rect 422 -577 423 -576
rect 635 -577 636 -576
rect 1094 -577 1095 -576
rect 1234 -577 1235 -576
rect 1255 -577 1256 -576
rect 1503 -577 1504 -576
rect 1507 -577 1508 -576
rect 289 -579 290 -578
rect 299 -579 300 -578
rect 579 -579 580 -578
rect 635 -579 636 -578
rect 639 -579 640 -578
rect 751 -579 752 -578
rect 772 -579 773 -578
rect 849 -579 850 -578
rect 856 -579 857 -578
rect 933 -579 934 -578
rect 968 -579 969 -578
rect 975 -579 976 -578
rect 1094 -579 1095 -578
rect 1115 -579 1116 -578
rect 1206 -579 1207 -578
rect 1234 -579 1235 -578
rect 639 -581 640 -580
rect 674 -581 675 -580
rect 688 -581 689 -580
rect 807 -581 808 -580
rect 849 -581 850 -580
rect 996 -581 997 -580
rect 1101 -581 1102 -580
rect 1115 -581 1116 -580
rect 1143 -581 1144 -580
rect 1206 -581 1207 -580
rect 555 -583 556 -582
rect 674 -583 675 -582
rect 698 -583 699 -582
rect 1003 -583 1004 -582
rect 1031 -583 1032 -582
rect 1101 -583 1102 -582
rect 51 -585 52 -584
rect 698 -585 699 -584
rect 702 -585 703 -584
rect 807 -585 808 -584
rect 866 -585 867 -584
rect 1143 -585 1144 -584
rect 513 -587 514 -586
rect 555 -587 556 -586
rect 660 -587 661 -586
rect 681 -587 682 -586
rect 702 -587 703 -586
rect 845 -587 846 -586
rect 877 -587 878 -586
rect 975 -587 976 -586
rect 1024 -587 1025 -586
rect 1031 -587 1032 -586
rect 86 -589 87 -588
rect 660 -589 661 -588
rect 737 -589 738 -588
rect 744 -589 745 -588
rect 870 -589 871 -588
rect 877 -589 878 -588
rect 884 -589 885 -588
rect 894 -589 895 -588
rect 926 -589 927 -588
rect 954 -589 955 -588
rect 1010 -589 1011 -588
rect 1024 -589 1025 -588
rect 86 -591 87 -590
rect 600 -591 601 -590
rect 744 -591 745 -590
rect 821 -591 822 -590
rect 912 -591 913 -590
rect 926 -591 927 -590
rect 940 -591 941 -590
rect 1010 -591 1011 -590
rect 453 -593 454 -592
rect 940 -593 941 -592
rect 821 -595 822 -594
rect 1486 -595 1487 -594
rect 912 -597 913 -596
rect 1374 -597 1375 -596
rect 1353 -599 1354 -598
rect 1374 -599 1375 -598
rect 110 -601 111 -600
rect 1353 -601 1354 -600
rect 9 -612 10 -611
rect 453 -612 454 -611
rect 492 -612 493 -611
rect 590 -612 591 -611
rect 604 -612 605 -611
rect 632 -612 633 -611
rect 653 -612 654 -611
rect 656 -612 657 -611
rect 674 -612 675 -611
rect 709 -612 710 -611
rect 761 -612 762 -611
rect 947 -612 948 -611
rect 1017 -612 1018 -611
rect 1052 -612 1053 -611
rect 1339 -612 1340 -611
rect 1528 -612 1529 -611
rect 1535 -612 1536 -611
rect 1787 -612 1788 -611
rect 9 -614 10 -613
rect 268 -614 269 -613
rect 303 -614 304 -613
rect 317 -614 318 -613
rect 320 -614 321 -613
rect 380 -614 381 -613
rect 408 -614 409 -613
rect 712 -614 713 -613
rect 786 -614 787 -613
rect 821 -614 822 -613
rect 824 -614 825 -613
rect 961 -614 962 -613
rect 1241 -614 1242 -613
rect 1339 -614 1340 -613
rect 1346 -614 1347 -613
rect 1619 -614 1620 -613
rect 1668 -614 1669 -613
rect 1801 -614 1802 -613
rect 16 -616 17 -615
rect 93 -616 94 -615
rect 114 -616 115 -615
rect 184 -616 185 -615
rect 233 -616 234 -615
rect 261 -616 262 -615
rect 303 -616 304 -615
rect 324 -616 325 -615
rect 362 -616 363 -615
rect 649 -616 650 -615
rect 653 -616 654 -615
rect 667 -616 668 -615
rect 677 -616 678 -615
rect 1430 -616 1431 -615
rect 1437 -616 1438 -615
rect 1591 -616 1592 -615
rect 1738 -616 1739 -615
rect 1822 -616 1823 -615
rect 30 -618 31 -617
rect 58 -618 59 -617
rect 72 -618 73 -617
rect 457 -618 458 -617
rect 544 -618 545 -617
rect 611 -618 612 -617
rect 660 -618 661 -617
rect 961 -618 962 -617
rect 1087 -618 1088 -617
rect 1346 -618 1347 -617
rect 1388 -618 1389 -617
rect 1535 -618 1536 -617
rect 1556 -618 1557 -617
rect 1657 -618 1658 -617
rect 1759 -618 1760 -617
rect 1794 -618 1795 -617
rect 30 -620 31 -619
rect 117 -620 118 -619
rect 145 -620 146 -619
rect 268 -620 269 -619
rect 352 -620 353 -619
rect 457 -620 458 -619
rect 569 -620 570 -619
rect 590 -620 591 -619
rect 604 -620 605 -619
rect 716 -620 717 -619
rect 786 -620 787 -619
rect 999 -620 1000 -619
rect 1157 -620 1158 -619
rect 1241 -620 1242 -619
rect 1325 -620 1326 -619
rect 1437 -620 1438 -619
rect 1444 -620 1445 -619
rect 1577 -620 1578 -619
rect 1766 -620 1767 -619
rect 1857 -620 1858 -619
rect 37 -622 38 -621
rect 870 -622 871 -621
rect 873 -622 874 -621
rect 1388 -622 1389 -621
rect 1409 -622 1410 -621
rect 1542 -622 1543 -621
rect 44 -624 45 -623
rect 96 -624 97 -623
rect 114 -624 115 -623
rect 1262 -624 1263 -623
rect 1290 -624 1291 -623
rect 1409 -624 1410 -623
rect 1416 -624 1417 -623
rect 1563 -624 1564 -623
rect 44 -626 45 -625
rect 499 -626 500 -625
rect 667 -626 668 -625
rect 702 -626 703 -625
rect 709 -626 710 -625
rect 1570 -626 1571 -625
rect 51 -628 52 -627
rect 72 -628 73 -627
rect 79 -628 80 -627
rect 82 -628 83 -627
rect 128 -628 129 -627
rect 352 -628 353 -627
rect 373 -628 374 -627
rect 429 -628 430 -627
rect 499 -628 500 -627
rect 506 -628 507 -627
rect 681 -628 682 -627
rect 702 -628 703 -627
rect 793 -628 794 -627
rect 912 -628 913 -627
rect 933 -628 934 -627
rect 1192 -628 1193 -627
rect 1206 -628 1207 -627
rect 1262 -628 1263 -627
rect 1269 -628 1270 -627
rect 1416 -628 1417 -627
rect 1423 -628 1424 -627
rect 1556 -628 1557 -627
rect 51 -630 52 -629
rect 103 -630 104 -629
rect 128 -630 129 -629
rect 135 -630 136 -629
rect 149 -630 150 -629
rect 324 -630 325 -629
rect 373 -630 374 -629
rect 383 -630 384 -629
rect 408 -630 409 -629
rect 422 -630 423 -629
rect 429 -630 430 -629
rect 471 -630 472 -629
rect 509 -630 510 -629
rect 1206 -630 1207 -629
rect 1227 -630 1228 -629
rect 1325 -630 1326 -629
rect 1451 -630 1452 -629
rect 1584 -630 1585 -629
rect 58 -632 59 -631
rect 65 -632 66 -631
rect 79 -632 80 -631
rect 107 -632 108 -631
rect 135 -632 136 -631
rect 1633 -632 1634 -631
rect 65 -634 66 -633
rect 142 -634 143 -633
rect 149 -634 150 -633
rect 212 -634 213 -633
rect 243 -634 244 -633
rect 443 -634 444 -633
rect 681 -634 682 -633
rect 751 -634 752 -633
rect 796 -634 797 -633
rect 1465 -634 1466 -633
rect 1472 -634 1473 -633
rect 1549 -634 1550 -633
rect 142 -636 143 -635
rect 765 -636 766 -635
rect 800 -636 801 -635
rect 821 -636 822 -635
rect 842 -636 843 -635
rect 1101 -636 1102 -635
rect 1108 -636 1109 -635
rect 1157 -636 1158 -635
rect 1178 -636 1179 -635
rect 1269 -636 1270 -635
rect 1353 -636 1354 -635
rect 1472 -636 1473 -635
rect 1479 -636 1480 -635
rect 1612 -636 1613 -635
rect 100 -638 101 -637
rect 1108 -638 1109 -637
rect 1129 -638 1130 -637
rect 1227 -638 1228 -637
rect 1360 -638 1361 -637
rect 1465 -638 1466 -637
rect 1468 -638 1469 -637
rect 1479 -638 1480 -637
rect 1486 -638 1487 -637
rect 1626 -638 1627 -637
rect 100 -640 101 -639
rect 191 -640 192 -639
rect 212 -640 213 -639
rect 467 -640 468 -639
rect 562 -640 563 -639
rect 800 -640 801 -639
rect 849 -640 850 -639
rect 1514 -640 1515 -639
rect 156 -642 157 -641
rect 891 -642 892 -641
rect 894 -642 895 -641
rect 1402 -642 1403 -641
rect 1458 -642 1459 -641
rect 1598 -642 1599 -641
rect 156 -644 157 -643
rect 401 -644 402 -643
rect 415 -644 416 -643
rect 513 -644 514 -643
rect 562 -644 563 -643
rect 730 -644 731 -643
rect 737 -644 738 -643
rect 765 -644 766 -643
rect 782 -644 783 -643
rect 1458 -644 1459 -643
rect 1493 -644 1494 -643
rect 1640 -644 1641 -643
rect 163 -646 164 -645
rect 492 -646 493 -645
rect 513 -646 514 -645
rect 548 -646 549 -645
rect 569 -646 570 -645
rect 842 -646 843 -645
rect 845 -646 846 -645
rect 1514 -646 1515 -645
rect 163 -648 164 -647
rect 646 -648 647 -647
rect 660 -648 661 -647
rect 737 -648 738 -647
rect 852 -648 853 -647
rect 1213 -648 1214 -647
rect 1255 -648 1256 -647
rect 1360 -648 1361 -647
rect 1374 -648 1375 -647
rect 1486 -648 1487 -647
rect 1500 -648 1501 -647
rect 1661 -648 1662 -647
rect 170 -650 171 -649
rect 527 -650 528 -649
rect 593 -650 594 -649
rect 849 -650 850 -649
rect 863 -650 864 -649
rect 1430 -650 1431 -649
rect 1507 -650 1508 -649
rect 1647 -650 1648 -649
rect 170 -652 171 -651
rect 1290 -652 1291 -651
rect 1297 -652 1298 -651
rect 1507 -652 1508 -651
rect 173 -654 174 -653
rect 618 -654 619 -653
rect 646 -654 647 -653
rect 719 -654 720 -653
rect 723 -654 724 -653
rect 751 -654 752 -653
rect 870 -654 871 -653
rect 922 -654 923 -653
rect 989 -654 990 -653
rect 1087 -654 1088 -653
rect 1115 -654 1116 -653
rect 1213 -654 1214 -653
rect 1248 -654 1249 -653
rect 1255 -654 1256 -653
rect 1311 -654 1312 -653
rect 1374 -654 1375 -653
rect 1381 -654 1382 -653
rect 1493 -654 1494 -653
rect 187 -656 188 -655
rect 1444 -656 1445 -655
rect 191 -658 192 -657
rect 198 -658 199 -657
rect 236 -658 237 -657
rect 415 -658 416 -657
rect 422 -658 423 -657
rect 530 -658 531 -657
rect 635 -658 636 -657
rect 989 -658 990 -657
rect 996 -658 997 -657
rect 1101 -658 1102 -657
rect 1136 -658 1137 -657
rect 1353 -658 1354 -657
rect 1367 -658 1368 -657
rect 1500 -658 1501 -657
rect 198 -660 199 -659
rect 338 -660 339 -659
rect 366 -660 367 -659
rect 471 -660 472 -659
rect 520 -660 521 -659
rect 548 -660 549 -659
rect 656 -660 657 -659
rect 723 -660 724 -659
rect 730 -660 731 -659
rect 744 -660 745 -659
rect 877 -660 878 -659
rect 947 -660 948 -659
rect 1024 -660 1025 -659
rect 1136 -660 1137 -659
rect 1164 -660 1165 -659
rect 1248 -660 1249 -659
rect 1276 -660 1277 -659
rect 1381 -660 1382 -659
rect 61 -662 62 -661
rect 1024 -662 1025 -661
rect 1031 -662 1032 -661
rect 1178 -662 1179 -661
rect 1185 -662 1186 -661
rect 1276 -662 1277 -661
rect 1283 -662 1284 -661
rect 1367 -662 1368 -661
rect 236 -664 237 -663
rect 583 -664 584 -663
rect 625 -664 626 -663
rect 744 -664 745 -663
rect 828 -664 829 -663
rect 877 -664 878 -663
rect 898 -664 899 -663
rect 933 -664 934 -663
rect 1038 -664 1039 -663
rect 1297 -664 1298 -663
rect 1318 -664 1319 -663
rect 1402 -664 1403 -663
rect 240 -666 241 -665
rect 366 -666 367 -665
rect 387 -666 388 -665
rect 618 -666 619 -665
rect 625 -666 626 -665
rect 1020 -666 1021 -665
rect 1059 -666 1060 -665
rect 1192 -666 1193 -665
rect 1199 -666 1200 -665
rect 1451 -666 1452 -665
rect 240 -668 241 -667
rect 831 -668 832 -667
rect 856 -668 857 -667
rect 1059 -668 1060 -667
rect 1066 -668 1067 -667
rect 1115 -668 1116 -667
rect 1171 -668 1172 -667
rect 1283 -668 1284 -667
rect 152 -670 153 -669
rect 856 -670 857 -669
rect 908 -670 909 -669
rect 1605 -670 1606 -669
rect 254 -672 255 -671
rect 866 -672 867 -671
rect 926 -672 927 -671
rect 1031 -672 1032 -671
rect 1045 -672 1046 -671
rect 1199 -672 1200 -671
rect 1234 -672 1235 -671
rect 1318 -672 1319 -671
rect 261 -674 262 -673
rect 345 -674 346 -673
rect 387 -674 388 -673
rect 600 -674 601 -673
rect 688 -674 689 -673
rect 863 -674 864 -673
rect 884 -674 885 -673
rect 926 -674 927 -673
rect 954 -674 955 -673
rect 1045 -674 1046 -673
rect 1073 -674 1074 -673
rect 1185 -674 1186 -673
rect 331 -676 332 -675
rect 338 -676 339 -675
rect 345 -676 346 -675
rect 481 -676 482 -675
rect 520 -676 521 -675
rect 541 -676 542 -675
rect 586 -676 587 -675
rect 898 -676 899 -675
rect 940 -676 941 -675
rect 1073 -676 1074 -675
rect 1080 -676 1081 -675
rect 1129 -676 1130 -675
rect 1143 -676 1144 -675
rect 1171 -676 1172 -675
rect 275 -678 276 -677
rect 331 -678 332 -677
rect 401 -678 402 -677
rect 639 -678 640 -677
rect 691 -678 692 -677
rect 915 -678 916 -677
rect 975 -678 976 -677
rect 1038 -678 1039 -677
rect 1150 -678 1151 -677
rect 1234 -678 1235 -677
rect 275 -680 276 -679
rect 394 -680 395 -679
rect 432 -680 433 -679
rect 1311 -680 1312 -679
rect 394 -682 395 -681
rect 779 -682 780 -681
rect 793 -682 794 -681
rect 940 -682 941 -681
rect 982 -682 983 -681
rect 1080 -682 1081 -681
rect 247 -684 248 -683
rect 779 -684 780 -683
rect 814 -684 815 -683
rect 982 -684 983 -683
rect 1003 -684 1004 -683
rect 1150 -684 1151 -683
rect 247 -686 248 -685
rect 289 -686 290 -685
rect 443 -686 444 -685
rect 576 -686 577 -685
rect 597 -686 598 -685
rect 639 -686 640 -685
rect 695 -686 696 -685
rect 1122 -686 1123 -685
rect 289 -688 290 -687
rect 296 -688 297 -687
rect 464 -688 465 -687
rect 527 -688 528 -687
rect 541 -688 542 -687
rect 611 -688 612 -687
rect 695 -688 696 -687
rect 971 -688 972 -687
rect 1010 -688 1011 -687
rect 1066 -688 1067 -687
rect 1122 -688 1123 -687
rect 1395 -688 1396 -687
rect 23 -690 24 -689
rect 464 -690 465 -689
rect 555 -690 556 -689
rect 576 -690 577 -689
rect 597 -690 598 -689
rect 1143 -690 1144 -689
rect 1304 -690 1305 -689
rect 1395 -690 1396 -689
rect 23 -692 24 -691
rect 310 -692 311 -691
rect 698 -692 699 -691
rect 1423 -692 1424 -691
rect 121 -694 122 -693
rect 310 -694 311 -693
rect 740 -694 741 -693
rect 1164 -694 1165 -693
rect 1220 -694 1221 -693
rect 1304 -694 1305 -693
rect 121 -696 122 -695
rect 450 -696 451 -695
rect 772 -696 773 -695
rect 975 -696 976 -695
rect 1094 -696 1095 -695
rect 1220 -696 1221 -695
rect 219 -698 220 -697
rect 296 -698 297 -697
rect 450 -698 451 -697
rect 478 -698 479 -697
rect 758 -698 759 -697
rect 772 -698 773 -697
rect 807 -698 808 -697
rect 814 -698 815 -697
rect 828 -698 829 -697
rect 1521 -698 1522 -697
rect 86 -700 87 -699
rect 219 -700 220 -699
rect 254 -700 255 -699
rect 478 -700 479 -699
rect 506 -700 507 -699
rect 1521 -700 1522 -699
rect 86 -702 87 -701
rect 226 -702 227 -701
rect 621 -702 622 -701
rect 807 -702 808 -701
rect 835 -702 836 -701
rect 954 -702 955 -701
rect 968 -702 969 -701
rect 1094 -702 1095 -701
rect 226 -704 227 -703
rect 758 -704 759 -703
rect 884 -704 885 -703
rect 901 -704 902 -703
rect 905 -704 906 -703
rect 1003 -704 1004 -703
rect 359 -706 360 -705
rect 835 -706 836 -705
rect 919 -706 920 -705
rect 1010 -706 1011 -705
rect 359 -708 360 -707
rect 485 -708 486 -707
rect 485 -710 486 -709
rect 1671 -710 1672 -709
rect 9 -721 10 -720
rect 93 -721 94 -720
rect 114 -721 115 -720
rect 1783 -721 1784 -720
rect 1787 -721 1788 -720
rect 1892 -721 1893 -720
rect 9 -723 10 -722
rect 422 -723 423 -722
rect 439 -723 440 -722
rect 555 -723 556 -722
rect 562 -723 563 -722
rect 649 -723 650 -722
rect 709 -723 710 -722
rect 1297 -723 1298 -722
rect 1458 -723 1459 -722
rect 1843 -723 1844 -722
rect 1857 -723 1858 -722
rect 1885 -723 1886 -722
rect 16 -725 17 -724
rect 117 -725 118 -724
rect 121 -725 122 -724
rect 124 -725 125 -724
rect 128 -725 129 -724
rect 138 -725 139 -724
rect 170 -725 171 -724
rect 180 -725 181 -724
rect 254 -725 255 -724
rect 257 -725 258 -724
rect 303 -725 304 -724
rect 306 -725 307 -724
rect 422 -725 423 -724
rect 719 -725 720 -724
rect 723 -725 724 -724
rect 737 -725 738 -724
rect 740 -725 741 -724
rect 1591 -725 1592 -724
rect 1605 -725 1606 -724
rect 1738 -725 1739 -724
rect 1801 -725 1802 -724
rect 1857 -725 1858 -724
rect 37 -727 38 -726
rect 233 -727 234 -726
rect 254 -727 255 -726
rect 527 -727 528 -726
rect 548 -727 549 -726
rect 562 -727 563 -726
rect 586 -727 587 -726
rect 996 -727 997 -726
rect 999 -727 1000 -726
rect 1563 -727 1564 -726
rect 1577 -727 1578 -726
rect 1731 -727 1732 -726
rect 1822 -727 1823 -726
rect 1850 -727 1851 -726
rect 37 -729 38 -728
rect 572 -729 573 -728
rect 597 -729 598 -728
rect 1451 -729 1452 -728
rect 1486 -729 1487 -728
rect 1675 -729 1676 -728
rect 1794 -729 1795 -728
rect 1822 -729 1823 -728
rect 58 -731 59 -730
rect 544 -731 545 -730
rect 555 -731 556 -730
rect 1591 -731 1592 -730
rect 1612 -731 1613 -730
rect 1759 -731 1760 -730
rect 30 -733 31 -732
rect 58 -733 59 -732
rect 79 -733 80 -732
rect 114 -733 115 -732
rect 121 -733 122 -732
rect 233 -733 234 -732
rect 268 -733 269 -732
rect 527 -733 528 -732
rect 618 -733 619 -732
rect 1297 -733 1298 -732
rect 1360 -733 1361 -732
rect 1451 -733 1452 -732
rect 1493 -733 1494 -732
rect 1605 -733 1606 -732
rect 1626 -733 1627 -732
rect 1787 -733 1788 -732
rect 30 -735 31 -734
rect 100 -735 101 -734
rect 135 -735 136 -734
rect 145 -735 146 -734
rect 170 -735 171 -734
rect 177 -735 178 -734
rect 201 -735 202 -734
rect 1563 -735 1564 -734
rect 1570 -735 1571 -734
rect 1577 -735 1578 -734
rect 1584 -735 1585 -734
rect 1766 -735 1767 -734
rect 93 -737 94 -736
rect 184 -737 185 -736
rect 268 -737 269 -736
rect 415 -737 416 -736
rect 443 -737 444 -736
rect 506 -737 507 -736
rect 520 -737 521 -736
rect 541 -737 542 -736
rect 614 -737 615 -736
rect 618 -737 619 -736
rect 621 -737 622 -736
rect 1486 -737 1487 -736
rect 1542 -737 1543 -736
rect 1689 -737 1690 -736
rect 65 -739 66 -738
rect 520 -739 521 -738
rect 628 -739 629 -738
rect 730 -739 731 -738
rect 779 -739 780 -738
rect 1472 -739 1473 -738
rect 1479 -739 1480 -738
rect 1584 -739 1585 -738
rect 1633 -739 1634 -738
rect 1794 -739 1795 -738
rect 65 -741 66 -740
rect 516 -741 517 -740
rect 632 -741 633 -740
rect 730 -741 731 -740
rect 758 -741 759 -740
rect 1472 -741 1473 -740
rect 1549 -741 1550 -740
rect 1745 -741 1746 -740
rect 100 -743 101 -742
rect 289 -743 290 -742
rect 303 -743 304 -742
rect 387 -743 388 -742
rect 443 -743 444 -742
rect 485 -743 486 -742
rect 495 -743 496 -742
rect 828 -743 829 -742
rect 831 -743 832 -742
rect 1668 -743 1669 -742
rect 1671 -743 1672 -742
rect 1717 -743 1718 -742
rect 107 -745 108 -744
rect 184 -745 185 -744
rect 275 -745 276 -744
rect 415 -745 416 -744
rect 450 -745 451 -744
rect 485 -745 486 -744
rect 590 -745 591 -744
rect 632 -745 633 -744
rect 674 -745 675 -744
rect 709 -745 710 -744
rect 712 -745 713 -744
rect 1801 -745 1802 -744
rect 107 -747 108 -746
rect 471 -747 472 -746
rect 478 -747 479 -746
rect 975 -747 976 -746
rect 1034 -747 1035 -746
rect 1829 -747 1830 -746
rect 135 -749 136 -748
rect 499 -749 500 -748
rect 653 -749 654 -748
rect 674 -749 675 -748
rect 681 -749 682 -748
rect 737 -749 738 -748
rect 779 -749 780 -748
rect 1710 -749 1711 -748
rect 173 -751 174 -750
rect 457 -751 458 -750
rect 464 -751 465 -750
rect 1073 -751 1074 -750
rect 1143 -751 1144 -750
rect 1696 -751 1697 -750
rect 96 -753 97 -752
rect 464 -753 465 -752
rect 478 -753 479 -752
rect 667 -753 668 -752
rect 716 -753 717 -752
rect 1199 -753 1200 -752
rect 1234 -753 1235 -752
rect 1360 -753 1361 -752
rect 1367 -753 1368 -752
rect 1458 -753 1459 -752
rect 1465 -753 1466 -752
rect 1542 -753 1543 -752
rect 1549 -753 1550 -752
rect 1598 -753 1599 -752
rect 1633 -753 1634 -752
rect 1661 -753 1662 -752
rect 156 -755 157 -754
rect 457 -755 458 -754
rect 467 -755 468 -754
rect 667 -755 668 -754
rect 723 -755 724 -754
rect 940 -755 941 -754
rect 1045 -755 1046 -754
rect 1143 -755 1144 -754
rect 1178 -755 1179 -754
rect 1199 -755 1200 -754
rect 1234 -755 1235 -754
rect 1304 -755 1305 -754
rect 1339 -755 1340 -754
rect 1479 -755 1480 -754
rect 1556 -755 1557 -754
rect 1703 -755 1704 -754
rect 51 -757 52 -756
rect 156 -757 157 -756
rect 275 -757 276 -756
rect 282 -757 283 -756
rect 289 -757 290 -756
rect 600 -757 601 -756
rect 639 -757 640 -756
rect 681 -757 682 -756
rect 782 -757 783 -756
rect 905 -757 906 -756
rect 919 -757 920 -756
rect 961 -757 962 -756
rect 1073 -757 1074 -756
rect 1220 -757 1221 -756
rect 1241 -757 1242 -756
rect 1367 -757 1368 -756
rect 1381 -757 1382 -756
rect 1493 -757 1494 -756
rect 1556 -757 1557 -756
rect 1780 -757 1781 -756
rect 282 -759 283 -758
rect 317 -759 318 -758
rect 324 -759 325 -758
rect 716 -759 717 -758
rect 793 -759 794 -758
rect 1409 -759 1410 -758
rect 1444 -759 1445 -758
rect 1612 -759 1613 -758
rect 1640 -759 1641 -758
rect 1773 -759 1774 -758
rect 296 -761 297 -760
rect 828 -761 829 -760
rect 835 -761 836 -760
rect 1045 -761 1046 -760
rect 1080 -761 1081 -760
rect 1178 -761 1179 -760
rect 1195 -761 1196 -760
rect 1682 -761 1683 -760
rect 324 -763 325 -762
rect 908 -763 909 -762
rect 922 -763 923 -762
rect 1752 -763 1753 -762
rect 345 -765 346 -764
rect 621 -765 622 -764
rect 772 -765 773 -764
rect 793 -765 794 -764
rect 800 -765 801 -764
rect 803 -765 804 -764
rect 807 -765 808 -764
rect 940 -765 941 -764
rect 1052 -765 1053 -764
rect 1080 -765 1081 -764
rect 1094 -765 1095 -764
rect 1220 -765 1221 -764
rect 1262 -765 1263 -764
rect 1339 -765 1340 -764
rect 1388 -765 1389 -764
rect 1598 -765 1599 -764
rect 1647 -765 1648 -764
rect 1808 -765 1809 -764
rect 345 -767 346 -766
rect 366 -767 367 -766
rect 373 -767 374 -766
rect 961 -767 962 -766
rect 1136 -767 1137 -766
rect 1241 -767 1242 -766
rect 1269 -767 1270 -766
rect 1381 -767 1382 -766
rect 1402 -767 1403 -766
rect 1570 -767 1571 -766
rect 310 -769 311 -768
rect 366 -769 367 -768
rect 373 -769 374 -768
rect 401 -769 402 -768
rect 436 -769 437 -768
rect 471 -769 472 -768
rect 492 -769 493 -768
rect 499 -769 500 -768
rect 569 -769 570 -768
rect 639 -769 640 -768
rect 695 -769 696 -768
rect 772 -769 773 -768
rect 800 -769 801 -768
rect 870 -769 871 -768
rect 884 -769 885 -768
rect 1626 -769 1627 -768
rect 54 -771 55 -770
rect 310 -771 311 -770
rect 401 -771 402 -770
rect 408 -771 409 -770
rect 450 -771 451 -770
rect 919 -771 920 -770
rect 933 -771 934 -770
rect 1094 -771 1095 -770
rect 1157 -771 1158 -770
rect 1262 -771 1263 -770
rect 1276 -771 1277 -770
rect 1388 -771 1389 -770
rect 1430 -771 1431 -770
rect 1647 -771 1648 -770
rect 142 -773 143 -772
rect 933 -773 934 -772
rect 954 -773 955 -772
rect 1052 -773 1053 -772
rect 1101 -773 1102 -772
rect 1157 -773 1158 -772
rect 1283 -773 1284 -772
rect 1444 -773 1445 -772
rect 1465 -773 1466 -772
rect 1528 -773 1529 -772
rect 142 -775 143 -774
rect 198 -775 199 -774
rect 359 -775 360 -774
rect 408 -775 409 -774
rect 492 -775 493 -774
rect 534 -775 535 -774
rect 576 -775 577 -774
rect 653 -775 654 -774
rect 803 -775 804 -774
rect 870 -775 871 -774
rect 898 -775 899 -774
rect 1304 -775 1305 -774
rect 1318 -775 1319 -774
rect 1402 -775 1403 -774
rect 1521 -775 1522 -774
rect 1640 -775 1641 -774
rect 44 -777 45 -776
rect 576 -777 577 -776
rect 604 -777 605 -776
rect 807 -777 808 -776
rect 814 -777 815 -776
rect 835 -777 836 -776
rect 842 -777 843 -776
rect 1353 -777 1354 -776
rect 1437 -777 1438 -776
rect 1521 -777 1522 -776
rect 177 -779 178 -778
rect 898 -779 899 -778
rect 901 -779 902 -778
rect 1619 -779 1620 -778
rect 198 -781 199 -780
rect 359 -781 360 -780
rect 534 -781 535 -780
rect 688 -781 689 -780
rect 824 -781 825 -780
rect 1514 -781 1515 -780
rect 548 -783 549 -782
rect 842 -783 843 -782
rect 845 -783 846 -782
rect 1724 -783 1725 -782
rect 583 -785 584 -784
rect 604 -785 605 -784
rect 611 -785 612 -784
rect 695 -785 696 -784
rect 782 -785 783 -784
rect 1514 -785 1515 -784
rect 163 -787 164 -786
rect 611 -787 612 -786
rect 625 -787 626 -786
rect 814 -787 815 -786
rect 849 -787 850 -786
rect 1017 -787 1018 -786
rect 1020 -787 1021 -786
rect 1437 -787 1438 -786
rect 1507 -787 1508 -786
rect 1619 -787 1620 -786
rect 163 -789 164 -788
rect 1423 -789 1424 -788
rect 583 -791 584 -790
rect 590 -791 591 -790
rect 625 -791 626 -790
rect 1661 -791 1662 -790
rect 646 -793 647 -792
rect 884 -793 885 -792
rect 912 -793 913 -792
rect 954 -793 955 -792
rect 1010 -793 1011 -792
rect 1269 -793 1270 -792
rect 1290 -793 1291 -792
rect 1836 -793 1837 -792
rect 212 -795 213 -794
rect 1010 -795 1011 -794
rect 1031 -795 1032 -794
rect 1136 -795 1137 -794
rect 1185 -795 1186 -794
rect 1283 -795 1284 -794
rect 1311 -795 1312 -794
rect 1423 -795 1424 -794
rect 296 -797 297 -796
rect 1031 -797 1032 -796
rect 1038 -797 1039 -796
rect 1101 -797 1102 -796
rect 1108 -797 1109 -796
rect 1290 -797 1291 -796
rect 1325 -797 1326 -796
rect 1409 -797 1410 -796
rect 1416 -797 1417 -796
rect 1507 -797 1508 -796
rect 166 -799 167 -798
rect 1325 -799 1326 -798
rect 1332 -799 1333 -798
rect 1353 -799 1354 -798
rect 1374 -799 1375 -798
rect 1416 -799 1417 -798
rect 429 -801 430 -800
rect 646 -801 647 -800
rect 744 -801 745 -800
rect 849 -801 850 -800
rect 926 -801 927 -800
rect 1017 -801 1018 -800
rect 1087 -801 1088 -800
rect 1185 -801 1186 -800
rect 1192 -801 1193 -800
rect 1311 -801 1312 -800
rect 1346 -801 1347 -800
rect 1430 -801 1431 -800
rect 79 -803 80 -802
rect 1087 -803 1088 -802
rect 1115 -803 1116 -802
rect 1276 -803 1277 -802
rect 352 -805 353 -804
rect 429 -805 430 -804
rect 509 -805 510 -804
rect 1038 -805 1039 -804
rect 1066 -805 1067 -804
rect 1115 -805 1116 -804
rect 1213 -805 1214 -804
rect 1318 -805 1319 -804
rect 338 -807 339 -806
rect 352 -807 353 -806
rect 691 -807 692 -806
rect 926 -807 927 -806
rect 947 -807 948 -806
rect 1066 -807 1067 -806
rect 1227 -807 1228 -806
rect 1332 -807 1333 -806
rect 82 -809 83 -808
rect 338 -809 339 -808
rect 744 -809 745 -808
rect 751 -809 752 -808
rect 761 -809 762 -808
rect 1213 -809 1214 -808
rect 1248 -809 1249 -808
rect 1374 -809 1375 -808
rect 702 -811 703 -810
rect 751 -811 752 -810
rect 761 -811 762 -810
rect 1206 -811 1207 -810
rect 1255 -811 1256 -810
rect 1528 -811 1529 -810
rect 789 -813 790 -812
rect 947 -813 948 -812
rect 971 -813 972 -812
rect 1346 -813 1347 -812
rect 821 -815 822 -814
rect 912 -815 913 -814
rect 982 -815 983 -814
rect 1206 -815 1207 -814
rect 821 -817 822 -816
rect 1500 -817 1501 -816
rect 863 -819 864 -818
rect 982 -819 983 -818
rect 989 -819 990 -818
rect 1108 -819 1109 -818
rect 1129 -819 1130 -818
rect 1248 -819 1249 -818
rect 1395 -819 1396 -818
rect 1500 -819 1501 -818
rect 765 -821 766 -820
rect 863 -821 864 -820
rect 989 -821 990 -820
rect 1654 -821 1655 -820
rect 226 -823 227 -822
rect 765 -823 766 -822
rect 1003 -823 1004 -822
rect 1129 -823 1130 -822
rect 1150 -823 1151 -822
rect 1227 -823 1228 -822
rect 226 -825 227 -824
rect 261 -825 262 -824
rect 1024 -825 1025 -824
rect 1255 -825 1256 -824
rect 240 -827 241 -826
rect 1003 -827 1004 -826
rect 1150 -827 1151 -826
rect 1164 -827 1165 -826
rect 1171 -827 1172 -826
rect 1395 -827 1396 -826
rect 72 -829 73 -828
rect 1164 -829 1165 -828
rect 1192 -829 1193 -828
rect 1654 -829 1655 -828
rect 72 -831 73 -830
rect 149 -831 150 -830
rect 240 -831 241 -830
rect 247 -831 248 -830
rect 261 -831 262 -830
rect 331 -831 332 -830
rect 891 -831 892 -830
rect 1024 -831 1025 -830
rect 1059 -831 1060 -830
rect 1171 -831 1172 -830
rect 44 -833 45 -832
rect 149 -833 150 -832
rect 205 -833 206 -832
rect 247 -833 248 -832
rect 331 -833 332 -832
rect 380 -833 381 -832
rect 877 -833 878 -832
rect 891 -833 892 -832
rect 968 -833 969 -832
rect 1059 -833 1060 -832
rect 191 -835 192 -834
rect 205 -835 206 -834
rect 380 -835 381 -834
rect 513 -835 514 -834
rect 660 -835 661 -834
rect 877 -835 878 -834
rect 128 -837 129 -836
rect 191 -837 192 -836
rect 212 -837 213 -836
rect 513 -837 514 -836
rect 579 -837 580 -836
rect 660 -837 661 -836
rect 856 -837 857 -836
rect 968 -837 969 -836
rect 786 -839 787 -838
rect 856 -839 857 -838
rect 786 -841 787 -840
rect 1535 -841 1536 -840
rect 1122 -843 1123 -842
rect 1535 -843 1536 -842
rect 558 -845 559 -844
rect 1122 -845 1123 -844
rect 86 -847 87 -846
rect 558 -847 559 -846
rect 86 -849 87 -848
rect 219 -849 220 -848
rect 23 -851 24 -850
rect 219 -851 220 -850
rect 23 -853 24 -852
rect 394 -853 395 -852
rect 187 -855 188 -854
rect 394 -855 395 -854
rect 2 -866 3 -865
rect 68 -866 69 -865
rect 86 -866 87 -865
rect 89 -866 90 -865
rect 110 -866 111 -865
rect 1234 -866 1235 -865
rect 1591 -866 1592 -865
rect 1594 -866 1595 -865
rect 1724 -866 1725 -865
rect 1864 -866 1865 -865
rect 1885 -866 1886 -865
rect 1913 -866 1914 -865
rect 37 -868 38 -867
rect 79 -868 80 -867
rect 86 -868 87 -867
rect 205 -868 206 -867
rect 261 -868 262 -867
rect 264 -868 265 -867
rect 310 -868 311 -867
rect 943 -868 944 -867
rect 1006 -868 1007 -867
rect 1766 -868 1767 -867
rect 1780 -868 1781 -867
rect 1822 -868 1823 -867
rect 1829 -868 1830 -867
rect 1941 -868 1942 -867
rect 30 -870 31 -869
rect 79 -870 80 -869
rect 114 -870 115 -869
rect 121 -870 122 -869
rect 135 -870 136 -869
rect 513 -870 514 -869
rect 516 -870 517 -869
rect 1668 -870 1669 -869
rect 1703 -870 1704 -869
rect 1766 -870 1767 -869
rect 1787 -870 1788 -869
rect 1829 -870 1830 -869
rect 1836 -870 1837 -869
rect 1948 -870 1949 -869
rect 30 -872 31 -871
rect 226 -872 227 -871
rect 261 -872 262 -871
rect 275 -872 276 -871
rect 310 -872 311 -871
rect 450 -872 451 -871
rect 460 -872 461 -871
rect 1920 -872 1921 -871
rect 37 -874 38 -873
rect 72 -874 73 -873
rect 121 -874 122 -873
rect 128 -874 129 -873
rect 156 -874 157 -873
rect 821 -874 822 -873
rect 828 -874 829 -873
rect 1612 -874 1613 -873
rect 1633 -874 1634 -873
rect 1885 -874 1886 -873
rect 1892 -874 1893 -873
rect 1955 -874 1956 -873
rect 51 -876 52 -875
rect 114 -876 115 -875
rect 163 -876 164 -875
rect 247 -876 248 -875
rect 275 -876 276 -875
rect 303 -876 304 -875
rect 338 -876 339 -875
rect 436 -876 437 -875
rect 450 -876 451 -875
rect 747 -876 748 -875
rect 779 -876 780 -875
rect 1066 -876 1067 -875
rect 1083 -876 1084 -875
rect 1731 -876 1732 -875
rect 1759 -876 1760 -875
rect 1871 -876 1872 -875
rect 47 -878 48 -877
rect 1066 -878 1067 -877
rect 1108 -878 1109 -877
rect 1111 -878 1112 -877
rect 1153 -878 1154 -877
rect 1675 -878 1676 -877
rect 1717 -878 1718 -877
rect 1787 -878 1788 -877
rect 1801 -878 1802 -877
rect 1934 -878 1935 -877
rect 51 -880 52 -879
rect 93 -880 94 -879
rect 177 -880 178 -879
rect 1024 -880 1025 -879
rect 1031 -880 1032 -879
rect 1598 -880 1599 -879
rect 1619 -880 1620 -879
rect 1675 -880 1676 -879
rect 1752 -880 1753 -879
rect 1759 -880 1760 -879
rect 1843 -880 1844 -879
rect 1906 -880 1907 -879
rect 65 -882 66 -881
rect 548 -882 549 -881
rect 572 -882 573 -881
rect 1325 -882 1326 -881
rect 1353 -882 1354 -881
rect 1598 -882 1599 -881
rect 1633 -882 1634 -881
rect 1878 -882 1879 -881
rect 65 -884 66 -883
rect 1013 -884 1014 -883
rect 1031 -884 1032 -883
rect 1528 -884 1529 -883
rect 1556 -884 1557 -883
rect 1612 -884 1613 -883
rect 1654 -884 1655 -883
rect 1724 -884 1725 -883
rect 1794 -884 1795 -883
rect 1843 -884 1844 -883
rect 1850 -884 1851 -883
rect 1881 -884 1882 -883
rect 72 -886 73 -885
rect 233 -886 234 -885
rect 247 -886 248 -885
rect 429 -886 430 -885
rect 492 -886 493 -885
rect 653 -886 654 -885
rect 684 -886 685 -885
rect 828 -886 829 -885
rect 915 -886 916 -885
rect 1325 -886 1326 -885
rect 1360 -886 1361 -885
rect 1619 -886 1620 -885
rect 1661 -886 1662 -885
rect 1717 -886 1718 -885
rect 1738 -886 1739 -885
rect 1794 -886 1795 -885
rect 1857 -886 1858 -885
rect 1892 -886 1893 -885
rect 93 -888 94 -887
rect 163 -888 164 -887
rect 177 -888 178 -887
rect 681 -888 682 -887
rect 688 -888 689 -887
rect 1479 -888 1480 -887
rect 1500 -888 1501 -887
rect 1556 -888 1557 -887
rect 1577 -888 1578 -887
rect 1836 -888 1837 -887
rect 128 -890 129 -889
rect 233 -890 234 -889
rect 268 -890 269 -889
rect 436 -890 437 -889
rect 492 -890 493 -889
rect 562 -890 563 -889
rect 576 -890 577 -889
rect 877 -890 878 -889
rect 919 -890 920 -889
rect 1073 -890 1074 -889
rect 1108 -890 1109 -889
rect 1178 -890 1179 -889
rect 1297 -890 1298 -889
rect 1353 -890 1354 -889
rect 1381 -890 1382 -889
rect 1654 -890 1655 -889
rect 1668 -890 1669 -889
rect 1745 -890 1746 -889
rect 1808 -890 1809 -889
rect 1857 -890 1858 -889
rect 156 -892 157 -891
rect 1360 -892 1361 -891
rect 1430 -892 1431 -891
rect 1479 -892 1480 -891
rect 1521 -892 1522 -891
rect 1577 -892 1578 -891
rect 1591 -892 1592 -891
rect 1710 -892 1711 -891
rect 180 -894 181 -893
rect 380 -894 381 -893
rect 387 -894 388 -893
rect 691 -894 692 -893
rect 705 -894 706 -893
rect 961 -894 962 -893
rect 985 -894 986 -893
rect 1780 -894 1781 -893
rect 58 -896 59 -895
rect 380 -896 381 -895
rect 429 -896 430 -895
rect 590 -896 591 -895
rect 604 -896 605 -895
rect 653 -896 654 -895
rect 688 -896 689 -895
rect 989 -896 990 -895
rect 1003 -896 1004 -895
rect 1024 -896 1025 -895
rect 1034 -896 1035 -895
rect 1444 -896 1445 -895
rect 1451 -896 1452 -895
rect 1500 -896 1501 -895
rect 1521 -896 1522 -895
rect 1584 -896 1585 -895
rect 1605 -896 1606 -895
rect 1661 -896 1662 -895
rect 1689 -896 1690 -895
rect 1738 -896 1739 -895
rect 187 -898 188 -897
rect 597 -898 598 -897
rect 604 -898 605 -897
rect 1563 -898 1564 -897
rect 1640 -898 1641 -897
rect 1689 -898 1690 -897
rect 1696 -898 1697 -897
rect 1752 -898 1753 -897
rect 191 -900 192 -899
rect 863 -900 864 -899
rect 877 -900 878 -899
rect 1192 -900 1193 -899
rect 1374 -900 1375 -899
rect 1430 -900 1431 -899
rect 1465 -900 1466 -899
rect 1801 -900 1802 -899
rect 198 -902 199 -901
rect 555 -902 556 -901
rect 583 -902 584 -901
rect 674 -902 675 -901
rect 723 -902 724 -901
rect 1234 -902 1235 -901
rect 1402 -902 1403 -901
rect 1444 -902 1445 -901
rect 1465 -902 1466 -901
rect 1542 -902 1543 -901
rect 1549 -902 1550 -901
rect 1850 -902 1851 -901
rect 170 -904 171 -903
rect 198 -904 199 -903
rect 201 -904 202 -903
rect 282 -904 283 -903
rect 338 -904 339 -903
rect 443 -904 444 -903
rect 478 -904 479 -903
rect 597 -904 598 -903
rect 618 -904 619 -903
rect 716 -904 717 -903
rect 726 -904 727 -903
rect 1696 -904 1697 -903
rect 170 -906 171 -905
rect 324 -906 325 -905
rect 394 -906 395 -905
rect 443 -906 444 -905
rect 485 -906 486 -905
rect 562 -906 563 -905
rect 586 -906 587 -905
rect 1045 -906 1046 -905
rect 1059 -906 1060 -905
rect 1528 -906 1529 -905
rect 1535 -906 1536 -905
rect 1605 -906 1606 -905
rect 1647 -906 1648 -905
rect 1710 -906 1711 -905
rect 184 -908 185 -907
rect 394 -908 395 -907
rect 408 -908 409 -907
rect 485 -908 486 -907
rect 495 -908 496 -907
rect 779 -908 780 -907
rect 782 -908 783 -907
rect 1703 -908 1704 -907
rect 184 -910 185 -909
rect 331 -910 332 -909
rect 506 -910 507 -909
rect 548 -910 549 -909
rect 590 -910 591 -909
rect 646 -910 647 -909
rect 674 -910 675 -909
rect 1038 -910 1039 -909
rect 1041 -910 1042 -909
rect 1570 -910 1571 -909
rect 205 -912 206 -911
rect 219 -912 220 -911
rect 240 -912 241 -911
rect 324 -912 325 -911
rect 422 -912 423 -911
rect 506 -912 507 -911
rect 513 -912 514 -911
rect 849 -912 850 -911
rect 856 -912 857 -911
rect 1381 -912 1382 -911
rect 1409 -912 1410 -911
rect 1451 -912 1452 -911
rect 1472 -912 1473 -911
rect 1745 -912 1746 -911
rect 212 -914 213 -913
rect 478 -914 479 -913
rect 527 -914 528 -913
rect 558 -914 559 -913
rect 618 -914 619 -913
rect 824 -914 825 -913
rect 831 -914 832 -913
rect 1374 -914 1375 -913
rect 1395 -914 1396 -913
rect 1409 -914 1410 -913
rect 1416 -914 1417 -913
rect 1570 -914 1571 -913
rect 142 -916 143 -915
rect 212 -916 213 -915
rect 240 -916 241 -915
rect 345 -916 346 -915
rect 415 -916 416 -915
rect 422 -916 423 -915
rect 499 -916 500 -915
rect 527 -916 528 -915
rect 534 -916 535 -915
rect 583 -916 584 -915
rect 621 -916 622 -915
rect 1822 -916 1823 -915
rect 226 -918 227 -917
rect 534 -918 535 -917
rect 537 -918 538 -917
rect 1206 -918 1207 -917
rect 1255 -918 1256 -917
rect 1416 -918 1417 -917
rect 1423 -918 1424 -917
rect 1549 -918 1550 -917
rect 1563 -918 1564 -917
rect 1899 -918 1900 -917
rect 268 -920 269 -919
rect 600 -920 601 -919
rect 625 -920 626 -919
rect 751 -920 752 -919
rect 758 -920 759 -919
rect 1045 -920 1046 -919
rect 1059 -920 1060 -919
rect 1297 -920 1298 -919
rect 1318 -920 1319 -919
rect 1423 -920 1424 -919
rect 1486 -920 1487 -919
rect 1535 -920 1536 -919
rect 282 -922 283 -921
rect 359 -922 360 -921
rect 415 -922 416 -921
rect 1094 -922 1095 -921
rect 1115 -922 1116 -921
rect 1255 -922 1256 -921
rect 1276 -922 1277 -921
rect 1318 -922 1319 -921
rect 1346 -922 1347 -921
rect 1402 -922 1403 -921
rect 1486 -922 1487 -921
rect 1916 -922 1917 -921
rect 289 -924 290 -923
rect 331 -924 332 -923
rect 359 -924 360 -923
rect 1783 -924 1784 -923
rect 289 -926 290 -925
rect 352 -926 353 -925
rect 499 -926 500 -925
rect 754 -926 755 -925
rect 758 -926 759 -925
rect 772 -926 773 -925
rect 775 -926 776 -925
rect 1584 -926 1585 -925
rect 254 -928 255 -927
rect 352 -928 353 -927
rect 541 -928 542 -927
rect 576 -928 577 -927
rect 625 -928 626 -927
rect 660 -928 661 -927
rect 709 -928 710 -927
rect 849 -928 850 -927
rect 856 -928 857 -927
rect 975 -928 976 -927
rect 1017 -928 1018 -927
rect 1073 -928 1074 -927
rect 1087 -928 1088 -927
rect 1115 -928 1116 -927
rect 1129 -928 1130 -927
rect 1178 -928 1179 -927
rect 1276 -928 1277 -927
rect 1388 -928 1389 -927
rect 1493 -928 1494 -927
rect 1542 -928 1543 -927
rect 58 -930 59 -929
rect 541 -930 542 -929
rect 639 -930 640 -929
rect 1017 -930 1018 -929
rect 1052 -930 1053 -929
rect 1087 -930 1088 -929
rect 1094 -930 1095 -929
rect 1101 -930 1102 -929
rect 1122 -930 1123 -929
rect 1129 -930 1130 -929
rect 1164 -930 1165 -929
rect 1192 -930 1193 -929
rect 1283 -930 1284 -929
rect 1346 -930 1347 -929
rect 1367 -930 1368 -929
rect 1472 -930 1473 -929
rect 1493 -930 1494 -929
rect 1682 -930 1683 -929
rect 254 -932 255 -931
rect 569 -932 570 -931
rect 639 -932 640 -931
rect 800 -932 801 -931
rect 814 -932 815 -931
rect 1101 -932 1102 -931
rect 1171 -932 1172 -931
rect 1206 -932 1207 -931
rect 1241 -932 1242 -931
rect 1283 -932 1284 -931
rect 1304 -932 1305 -931
rect 1367 -932 1368 -931
rect 1507 -932 1508 -931
rect 1640 -932 1641 -931
rect 1682 -932 1683 -931
rect 1818 -932 1819 -931
rect 142 -934 143 -933
rect 814 -934 815 -933
rect 821 -934 822 -933
rect 842 -934 843 -933
rect 863 -934 864 -933
rect 912 -934 913 -933
rect 922 -934 923 -933
rect 1731 -934 1732 -933
rect 296 -936 297 -935
rect 408 -936 409 -935
rect 520 -936 521 -935
rect 709 -936 710 -935
rect 716 -936 717 -935
rect 730 -936 731 -935
rect 740 -936 741 -935
rect 1808 -936 1809 -935
rect 296 -938 297 -937
rect 471 -938 472 -937
rect 544 -938 545 -937
rect 569 -938 570 -937
rect 646 -938 647 -937
rect 905 -938 906 -937
rect 922 -938 923 -937
rect 1927 -938 1928 -937
rect 166 -940 167 -939
rect 905 -940 906 -939
rect 947 -940 948 -939
rect 989 -940 990 -939
rect 1003 -940 1004 -939
rect 1164 -940 1165 -939
rect 1311 -940 1312 -939
rect 1388 -940 1389 -939
rect 1458 -940 1459 -939
rect 1507 -940 1508 -939
rect 1594 -940 1595 -939
rect 1647 -940 1648 -939
rect 317 -942 318 -941
rect 345 -942 346 -941
rect 401 -942 402 -941
rect 471 -942 472 -941
rect 660 -942 661 -941
rect 940 -942 941 -941
rect 947 -942 948 -941
rect 982 -942 983 -941
rect 1062 -942 1063 -941
rect 1514 -942 1515 -941
rect 149 -944 150 -943
rect 317 -944 318 -943
rect 401 -944 402 -943
rect 457 -944 458 -943
rect 464 -944 465 -943
rect 520 -944 521 -943
rect 702 -944 703 -943
rect 1241 -944 1242 -943
rect 1262 -944 1263 -943
rect 1311 -944 1312 -943
rect 100 -946 101 -945
rect 149 -946 150 -945
rect 373 -946 374 -945
rect 702 -946 703 -945
rect 730 -946 731 -945
rect 1010 -946 1011 -945
rect 1143 -946 1144 -945
rect 1171 -946 1172 -945
rect 1213 -946 1214 -945
rect 1458 -946 1459 -945
rect 9 -948 10 -947
rect 100 -948 101 -947
rect 107 -948 108 -947
rect 373 -948 374 -947
rect 390 -948 391 -947
rect 464 -948 465 -947
rect 744 -948 745 -947
rect 786 -948 787 -947
rect 789 -948 790 -947
rect 842 -948 843 -947
rect 891 -948 892 -947
rect 1052 -948 1053 -947
rect 1080 -948 1081 -947
rect 1143 -948 1144 -947
rect 1157 -948 1158 -947
rect 1304 -948 1305 -947
rect 9 -950 10 -949
rect 23 -950 24 -949
rect 44 -950 45 -949
rect 107 -950 108 -949
rect 135 -950 136 -949
rect 457 -950 458 -949
rect 611 -950 612 -949
rect 786 -950 787 -949
rect 800 -950 801 -949
rect 940 -950 941 -949
rect 954 -950 955 -949
rect 975 -950 976 -949
rect 1010 -950 1011 -949
rect 1773 -950 1774 -949
rect 23 -952 24 -951
rect 194 -952 195 -951
rect 611 -952 612 -951
rect 695 -952 696 -951
rect 744 -952 745 -951
rect 1290 -952 1291 -951
rect 667 -954 668 -953
rect 695 -954 696 -953
rect 761 -954 762 -953
rect 1514 -954 1515 -953
rect 667 -956 668 -955
rect 870 -956 871 -955
rect 884 -956 885 -955
rect 954 -956 955 -955
rect 961 -956 962 -955
rect 996 -956 997 -955
rect 1034 -956 1035 -955
rect 1773 -956 1774 -955
rect 765 -958 766 -957
rect 982 -958 983 -957
rect 996 -958 997 -957
rect 1038 -958 1039 -957
rect 1080 -958 1081 -957
rect 1815 -958 1816 -957
rect 737 -960 738 -959
rect 765 -960 766 -959
rect 772 -960 773 -959
rect 1269 -960 1270 -959
rect 807 -962 808 -961
rect 891 -962 892 -961
rect 1157 -962 1158 -961
rect 1395 -962 1396 -961
rect 793 -964 794 -963
rect 807 -964 808 -963
rect 835 -964 836 -963
rect 870 -964 871 -963
rect 884 -964 885 -963
rect 898 -964 899 -963
rect 1185 -964 1186 -963
rect 1213 -964 1214 -963
rect 1227 -964 1228 -963
rect 1269 -964 1270 -963
rect 54 -966 55 -965
rect 835 -966 836 -965
rect 1150 -966 1151 -965
rect 1185 -966 1186 -965
rect 1248 -966 1249 -965
rect 1290 -966 1291 -965
rect 236 -968 237 -967
rect 1248 -968 1249 -967
rect 1262 -968 1263 -967
rect 1626 -968 1627 -967
rect 439 -970 440 -969
rect 898 -970 899 -969
rect 1437 -970 1438 -969
rect 1626 -970 1627 -969
rect 793 -972 794 -971
rect 1160 -972 1161 -971
rect 1332 -972 1333 -971
rect 1437 -972 1438 -971
rect 1199 -974 1200 -973
rect 1332 -974 1333 -973
rect 628 -976 629 -975
rect 1199 -976 1200 -975
rect 47 -987 48 -986
rect 702 -987 703 -986
rect 733 -987 734 -986
rect 772 -987 773 -986
rect 775 -987 776 -986
rect 821 -987 822 -986
rect 866 -987 867 -986
rect 1423 -987 1424 -986
rect 1745 -987 1746 -986
rect 1899 -987 1900 -986
rect 1927 -987 1928 -986
rect 1976 -987 1977 -986
rect 58 -989 59 -988
rect 453 -989 454 -988
rect 457 -989 458 -988
rect 537 -989 538 -988
rect 541 -989 542 -988
rect 625 -989 626 -988
rect 656 -989 657 -988
rect 1416 -989 1417 -988
rect 1710 -989 1711 -988
rect 1745 -989 1746 -988
rect 1867 -989 1868 -988
rect 1892 -989 1893 -988
rect 1927 -989 1928 -988
rect 1934 -989 1935 -988
rect 1941 -989 1942 -988
rect 1962 -989 1963 -988
rect 58 -991 59 -990
rect 170 -991 171 -990
rect 240 -991 241 -990
rect 684 -991 685 -990
rect 709 -991 710 -990
rect 821 -991 822 -990
rect 870 -991 871 -990
rect 915 -991 916 -990
rect 919 -991 920 -990
rect 1430 -991 1431 -990
rect 1710 -991 1711 -990
rect 1766 -991 1767 -990
rect 1878 -991 1879 -990
rect 1906 -991 1907 -990
rect 1948 -991 1949 -990
rect 1969 -991 1970 -990
rect 68 -993 69 -992
rect 394 -993 395 -992
rect 443 -993 444 -992
rect 457 -993 458 -992
rect 485 -993 486 -992
rect 604 -993 605 -992
rect 625 -993 626 -992
rect 1437 -993 1438 -992
rect 1584 -993 1585 -992
rect 1878 -993 1879 -992
rect 1948 -993 1949 -992
rect 1955 -993 1956 -992
rect 30 -995 31 -994
rect 394 -995 395 -994
rect 485 -995 486 -994
rect 618 -995 619 -994
rect 674 -995 675 -994
rect 709 -995 710 -994
rect 716 -995 717 -994
rect 772 -995 773 -994
rect 779 -995 780 -994
rect 1416 -995 1417 -994
rect 1493 -995 1494 -994
rect 1584 -995 1585 -994
rect 30 -997 31 -996
rect 51 -997 52 -996
rect 72 -997 73 -996
rect 390 -997 391 -996
rect 513 -997 514 -996
rect 604 -997 605 -996
rect 667 -997 668 -996
rect 716 -997 717 -996
rect 737 -997 738 -996
rect 758 -997 759 -996
rect 761 -997 762 -996
rect 1724 -997 1725 -996
rect 51 -999 52 -998
rect 408 -999 409 -998
rect 478 -999 479 -998
rect 667 -999 668 -998
rect 674 -999 675 -998
rect 1192 -999 1193 -998
rect 1241 -999 1242 -998
rect 1244 -999 1245 -998
rect 1276 -999 1277 -998
rect 1423 -999 1424 -998
rect 1493 -999 1494 -998
rect 1500 -999 1501 -998
rect 1724 -999 1725 -998
rect 1885 -999 1886 -998
rect 72 -1001 73 -1000
rect 635 -1001 636 -1000
rect 681 -1001 682 -1000
rect 1178 -1001 1179 -1000
rect 1241 -1001 1242 -1000
rect 1269 -1001 1270 -1000
rect 1276 -1001 1277 -1000
rect 1290 -1001 1291 -1000
rect 1409 -1001 1410 -1000
rect 1430 -1001 1431 -1000
rect 1500 -1001 1501 -1000
rect 1507 -1001 1508 -1000
rect 82 -1003 83 -1002
rect 1017 -1003 1018 -1002
rect 1020 -1003 1021 -1002
rect 1255 -1003 1256 -1002
rect 1367 -1003 1368 -1002
rect 1409 -1003 1410 -1002
rect 1507 -1003 1508 -1002
rect 1514 -1003 1515 -1002
rect 86 -1005 87 -1004
rect 145 -1005 146 -1004
rect 149 -1005 150 -1004
rect 170 -1005 171 -1004
rect 240 -1005 241 -1004
rect 401 -1005 402 -1004
rect 408 -1005 409 -1004
rect 492 -1005 493 -1004
rect 513 -1005 514 -1004
rect 611 -1005 612 -1004
rect 646 -1005 647 -1004
rect 1178 -1005 1179 -1004
rect 1244 -1005 1245 -1004
rect 1269 -1005 1270 -1004
rect 1514 -1005 1515 -1004
rect 1570 -1005 1571 -1004
rect 9 -1007 10 -1006
rect 86 -1007 87 -1006
rect 93 -1007 94 -1006
rect 219 -1007 220 -1006
rect 282 -1007 283 -1006
rect 726 -1007 727 -1006
rect 737 -1007 738 -1006
rect 1437 -1007 1438 -1006
rect 1535 -1007 1536 -1006
rect 1570 -1007 1571 -1006
rect 9 -1009 10 -1008
rect 226 -1009 227 -1008
rect 282 -1009 283 -1008
rect 436 -1009 437 -1008
rect 478 -1009 479 -1008
rect 779 -1009 780 -1008
rect 786 -1009 787 -1008
rect 957 -1009 958 -1008
rect 968 -1009 969 -1008
rect 1290 -1009 1291 -1008
rect 1535 -1009 1536 -1008
rect 1598 -1009 1599 -1008
rect 79 -1011 80 -1010
rect 149 -1011 150 -1010
rect 156 -1011 157 -1010
rect 443 -1011 444 -1010
rect 492 -1011 493 -1010
rect 730 -1011 731 -1010
rect 747 -1011 748 -1010
rect 1458 -1011 1459 -1010
rect 1598 -1011 1599 -1010
rect 1633 -1011 1634 -1010
rect 79 -1013 80 -1012
rect 1234 -1013 1235 -1012
rect 1255 -1013 1256 -1012
rect 1297 -1013 1298 -1012
rect 1451 -1013 1452 -1012
rect 1458 -1013 1459 -1012
rect 68 -1015 69 -1014
rect 1451 -1015 1452 -1014
rect 96 -1017 97 -1016
rect 758 -1017 759 -1016
rect 863 -1017 864 -1016
rect 870 -1017 871 -1016
rect 891 -1017 892 -1016
rect 1367 -1017 1368 -1016
rect 107 -1019 108 -1018
rect 128 -1019 129 -1018
rect 142 -1019 143 -1018
rect 159 -1019 160 -1018
rect 226 -1019 227 -1018
rect 660 -1019 661 -1018
rect 681 -1019 682 -1018
rect 1528 -1019 1529 -1018
rect 128 -1021 129 -1020
rect 310 -1021 311 -1020
rect 345 -1021 346 -1020
rect 436 -1021 437 -1020
rect 506 -1021 507 -1020
rect 968 -1021 969 -1020
rect 982 -1021 983 -1020
rect 1864 -1021 1865 -1020
rect 142 -1023 143 -1022
rect 191 -1023 192 -1022
rect 268 -1023 269 -1022
rect 786 -1023 787 -1022
rect 842 -1023 843 -1022
rect 891 -1023 892 -1022
rect 894 -1023 895 -1022
rect 898 -1023 899 -1022
rect 912 -1023 913 -1022
rect 1472 -1023 1473 -1022
rect 37 -1025 38 -1024
rect 268 -1025 269 -1024
rect 296 -1025 297 -1024
rect 534 -1025 535 -1024
rect 565 -1025 566 -1024
rect 611 -1025 612 -1024
rect 632 -1025 633 -1024
rect 660 -1025 661 -1024
rect 702 -1025 703 -1024
rect 730 -1025 731 -1024
rect 751 -1025 752 -1024
rect 1773 -1025 1774 -1024
rect 37 -1027 38 -1026
rect 471 -1027 472 -1026
rect 499 -1027 500 -1026
rect 534 -1027 535 -1026
rect 569 -1027 570 -1026
rect 1083 -1027 1084 -1026
rect 1108 -1027 1109 -1026
rect 1157 -1027 1158 -1026
rect 1160 -1027 1161 -1026
rect 1850 -1027 1851 -1026
rect 156 -1029 157 -1028
rect 1062 -1029 1063 -1028
rect 1108 -1029 1109 -1028
rect 1122 -1029 1123 -1028
rect 1136 -1029 1137 -1028
rect 1528 -1029 1529 -1028
rect 1773 -1029 1774 -1028
rect 1920 -1029 1921 -1028
rect 191 -1031 192 -1030
rect 236 -1031 237 -1030
rect 303 -1031 304 -1030
rect 345 -1031 346 -1030
rect 387 -1031 388 -1030
rect 562 -1031 563 -1030
rect 579 -1031 580 -1030
rect 1633 -1031 1634 -1030
rect 198 -1033 199 -1032
rect 296 -1033 297 -1032
rect 380 -1033 381 -1032
rect 387 -1033 388 -1032
rect 397 -1033 398 -1032
rect 912 -1033 913 -1032
rect 919 -1033 920 -1032
rect 926 -1033 927 -1032
rect 940 -1033 941 -1032
rect 1871 -1033 1872 -1032
rect 121 -1035 122 -1034
rect 198 -1035 199 -1034
rect 205 -1035 206 -1034
rect 471 -1035 472 -1034
rect 499 -1035 500 -1034
rect 527 -1035 528 -1034
rect 618 -1035 619 -1034
rect 1136 -1035 1137 -1034
rect 1139 -1035 1140 -1034
rect 1808 -1035 1809 -1034
rect 100 -1037 101 -1036
rect 527 -1037 528 -1036
rect 646 -1037 647 -1036
rect 849 -1037 850 -1036
rect 877 -1037 878 -1036
rect 898 -1037 899 -1036
rect 905 -1037 906 -1036
rect 1850 -1037 1851 -1036
rect 44 -1039 45 -1038
rect 100 -1039 101 -1038
rect 114 -1039 115 -1038
rect 121 -1039 122 -1038
rect 219 -1039 220 -1038
rect 926 -1039 927 -1038
rect 954 -1039 955 -1038
rect 1006 -1039 1007 -1038
rect 1010 -1039 1011 -1038
rect 1766 -1039 1767 -1038
rect 1808 -1039 1809 -1038
rect 1829 -1039 1830 -1038
rect 114 -1041 115 -1040
rect 177 -1041 178 -1040
rect 205 -1041 206 -1040
rect 954 -1041 955 -1040
rect 982 -1041 983 -1040
rect 996 -1041 997 -1040
rect 1010 -1041 1011 -1040
rect 1052 -1041 1053 -1040
rect 1059 -1041 1060 -1040
rect 1549 -1041 1550 -1040
rect 1591 -1041 1592 -1040
rect 1829 -1041 1830 -1040
rect 177 -1043 178 -1042
rect 429 -1043 430 -1042
rect 450 -1043 451 -1042
rect 506 -1043 507 -1042
rect 520 -1043 521 -1042
rect 569 -1043 570 -1042
rect 688 -1043 689 -1042
rect 940 -1043 941 -1042
rect 961 -1043 962 -1042
rect 996 -1043 997 -1042
rect 1013 -1043 1014 -1042
rect 1192 -1043 1193 -1042
rect 1220 -1043 1221 -1042
rect 1234 -1043 1235 -1042
rect 1297 -1043 1298 -1042
rect 1304 -1043 1305 -1042
rect 1360 -1043 1361 -1042
rect 1871 -1043 1872 -1042
rect 233 -1045 234 -1044
rect 450 -1045 451 -1044
rect 520 -1045 521 -1044
rect 922 -1045 923 -1044
rect 985 -1045 986 -1044
rect 1654 -1045 1655 -1044
rect 254 -1047 255 -1046
rect 303 -1047 304 -1046
rect 352 -1047 353 -1046
rect 429 -1047 430 -1046
rect 688 -1047 689 -1046
rect 1153 -1047 1154 -1046
rect 1206 -1047 1207 -1046
rect 1220 -1047 1221 -1046
rect 1262 -1047 1263 -1046
rect 1654 -1047 1655 -1046
rect 254 -1049 255 -1048
rect 324 -1049 325 -1048
rect 352 -1049 353 -1048
rect 649 -1049 650 -1048
rect 695 -1049 696 -1048
rect 1153 -1049 1154 -1048
rect 1199 -1049 1200 -1048
rect 1206 -1049 1207 -1048
rect 1213 -1049 1214 -1048
rect 1262 -1049 1263 -1048
rect 1304 -1049 1305 -1048
rect 1311 -1049 1312 -1048
rect 1353 -1049 1354 -1048
rect 1360 -1049 1361 -1048
rect 1472 -1049 1473 -1048
rect 1479 -1049 1480 -1048
rect 1549 -1049 1550 -1048
rect 1787 -1049 1788 -1048
rect 366 -1051 367 -1050
rect 380 -1051 381 -1050
rect 401 -1051 402 -1050
rect 422 -1051 423 -1050
rect 607 -1051 608 -1050
rect 695 -1051 696 -1050
rect 723 -1051 724 -1050
rect 1199 -1051 1200 -1050
rect 1213 -1051 1214 -1050
rect 1283 -1051 1284 -1050
rect 1479 -1051 1480 -1050
rect 1556 -1051 1557 -1050
rect 1591 -1051 1592 -1050
rect 1689 -1051 1690 -1050
rect 1787 -1051 1788 -1050
rect 1815 -1051 1816 -1050
rect 275 -1053 276 -1052
rect 422 -1053 423 -1052
rect 653 -1053 654 -1052
rect 723 -1053 724 -1052
rect 751 -1053 752 -1052
rect 856 -1053 857 -1052
rect 877 -1053 878 -1052
rect 884 -1053 885 -1052
rect 1003 -1053 1004 -1052
rect 1353 -1053 1354 -1052
rect 1465 -1053 1466 -1052
rect 1556 -1053 1557 -1052
rect 1563 -1053 1564 -1052
rect 1689 -1053 1690 -1052
rect 1815 -1053 1816 -1052
rect 1843 -1053 1844 -1052
rect 16 -1055 17 -1054
rect 884 -1055 885 -1054
rect 1003 -1055 1004 -1054
rect 1045 -1055 1046 -1054
rect 1048 -1055 1049 -1054
rect 1801 -1055 1802 -1054
rect 16 -1057 17 -1056
rect 215 -1057 216 -1056
rect 275 -1057 276 -1056
rect 317 -1057 318 -1056
rect 324 -1057 325 -1056
rect 1045 -1057 1046 -1056
rect 1052 -1057 1053 -1056
rect 1073 -1057 1074 -1056
rect 1122 -1057 1123 -1056
rect 1129 -1057 1130 -1056
rect 1150 -1057 1151 -1056
rect 1682 -1057 1683 -1056
rect 1696 -1057 1697 -1056
rect 1843 -1057 1844 -1056
rect 317 -1059 318 -1058
rect 744 -1059 745 -1058
rect 782 -1059 783 -1058
rect 1283 -1059 1284 -1058
rect 1563 -1059 1564 -1058
rect 1626 -1059 1627 -1058
rect 1682 -1059 1683 -1058
rect 1738 -1059 1739 -1058
rect 1759 -1059 1760 -1058
rect 1801 -1059 1802 -1058
rect 338 -1061 339 -1060
rect 1129 -1061 1130 -1060
rect 1150 -1061 1151 -1060
rect 1465 -1061 1466 -1060
rect 1626 -1061 1627 -1060
rect 1647 -1061 1648 -1060
rect 1696 -1061 1697 -1060
rect 1752 -1061 1753 -1060
rect 331 -1063 332 -1062
rect 338 -1063 339 -1062
rect 366 -1063 367 -1062
rect 632 -1063 633 -1062
rect 744 -1063 745 -1062
rect 800 -1063 801 -1062
rect 807 -1063 808 -1062
rect 856 -1063 857 -1062
rect 1017 -1063 1018 -1062
rect 1738 -1063 1739 -1062
rect 135 -1065 136 -1064
rect 331 -1065 332 -1064
rect 765 -1065 766 -1064
rect 807 -1065 808 -1064
rect 835 -1065 836 -1064
rect 905 -1065 906 -1064
rect 1031 -1065 1032 -1064
rect 1759 -1065 1760 -1064
rect 135 -1067 136 -1066
rect 415 -1067 416 -1066
rect 597 -1067 598 -1066
rect 765 -1067 766 -1066
rect 793 -1067 794 -1066
rect 961 -1067 962 -1066
rect 1038 -1067 1039 -1066
rect 1101 -1067 1102 -1066
rect 1227 -1067 1228 -1066
rect 1311 -1067 1312 -1066
rect 1612 -1067 1613 -1066
rect 1647 -1067 1648 -1066
rect 359 -1069 360 -1068
rect 597 -1069 598 -1068
rect 628 -1069 629 -1068
rect 835 -1069 836 -1068
rect 842 -1069 843 -1068
rect 1115 -1069 1116 -1068
rect 1227 -1069 1228 -1068
rect 1836 -1069 1837 -1068
rect 359 -1071 360 -1070
rect 373 -1071 374 -1070
rect 415 -1071 416 -1070
rect 464 -1071 465 -1070
rect 639 -1071 640 -1070
rect 793 -1071 794 -1070
rect 800 -1071 801 -1070
rect 1034 -1071 1035 -1070
rect 1041 -1071 1042 -1070
rect 1640 -1071 1641 -1070
rect 1836 -1071 1837 -1070
rect 1857 -1071 1858 -1070
rect 247 -1073 248 -1072
rect 464 -1073 465 -1072
rect 639 -1073 640 -1072
rect 754 -1073 755 -1072
rect 828 -1073 829 -1072
rect 1101 -1073 1102 -1072
rect 1115 -1073 1116 -1072
rect 1164 -1073 1165 -1072
rect 1521 -1073 1522 -1072
rect 1612 -1073 1613 -1072
rect 1640 -1073 1641 -1072
rect 1661 -1073 1662 -1072
rect 1822 -1073 1823 -1072
rect 1857 -1073 1858 -1072
rect 184 -1075 185 -1074
rect 247 -1075 248 -1074
rect 289 -1075 290 -1074
rect 373 -1075 374 -1074
rect 653 -1075 654 -1074
rect 1521 -1075 1522 -1074
rect 1661 -1075 1662 -1074
rect 1703 -1075 1704 -1074
rect 163 -1077 164 -1076
rect 184 -1077 185 -1076
rect 212 -1077 213 -1076
rect 289 -1077 290 -1076
rect 684 -1077 685 -1076
rect 1822 -1077 1823 -1076
rect 23 -1079 24 -1078
rect 212 -1079 213 -1078
rect 849 -1079 850 -1078
rect 1381 -1079 1382 -1078
rect 1675 -1079 1676 -1078
rect 1703 -1079 1704 -1078
rect 23 -1081 24 -1080
rect 310 -1081 311 -1080
rect 947 -1081 948 -1080
rect 1031 -1081 1032 -1080
rect 1059 -1081 1060 -1080
rect 1094 -1081 1095 -1080
rect 1143 -1081 1144 -1080
rect 1164 -1081 1165 -1080
rect 1381 -1081 1382 -1080
rect 1388 -1081 1389 -1080
rect 1675 -1081 1676 -1080
rect 1731 -1081 1732 -1080
rect 163 -1083 164 -1082
rect 590 -1083 591 -1082
rect 947 -1083 948 -1082
rect 975 -1083 976 -1082
rect 1024 -1083 1025 -1082
rect 1038 -1083 1039 -1082
rect 1066 -1083 1067 -1082
rect 1094 -1083 1095 -1082
rect 1143 -1083 1144 -1082
rect 1185 -1083 1186 -1082
rect 1388 -1083 1389 -1082
rect 1395 -1083 1396 -1082
rect 1577 -1083 1578 -1082
rect 1731 -1083 1732 -1082
rect 555 -1085 556 -1084
rect 590 -1085 591 -1084
rect 863 -1085 864 -1084
rect 1066 -1085 1067 -1084
rect 1073 -1085 1074 -1084
rect 1087 -1085 1088 -1084
rect 1185 -1085 1186 -1084
rect 1230 -1085 1231 -1084
rect 1339 -1085 1340 -1084
rect 1395 -1085 1396 -1084
rect 1542 -1085 1543 -1084
rect 1577 -1085 1578 -1084
rect 555 -1087 556 -1086
rect 576 -1087 577 -1086
rect 740 -1087 741 -1086
rect 1087 -1087 1088 -1086
rect 1332 -1087 1333 -1086
rect 1339 -1087 1340 -1086
rect 1542 -1087 1543 -1086
rect 1605 -1087 1606 -1086
rect 576 -1089 577 -1088
rect 1248 -1089 1249 -1088
rect 1325 -1089 1326 -1088
rect 1332 -1089 1333 -1088
rect 1605 -1089 1606 -1088
rect 1717 -1089 1718 -1088
rect 740 -1091 741 -1090
rect 1619 -1091 1620 -1090
rect 1717 -1091 1718 -1090
rect 1780 -1091 1781 -1090
rect 65 -1093 66 -1092
rect 1619 -1093 1620 -1092
rect 1780 -1093 1781 -1092
rect 1794 -1093 1795 -1092
rect 2 -1095 3 -1094
rect 65 -1095 66 -1094
rect 828 -1095 829 -1094
rect 1230 -1095 1231 -1094
rect 1248 -1095 1249 -1094
rect 1402 -1095 1403 -1094
rect 1668 -1095 1669 -1094
rect 1794 -1095 1795 -1094
rect 110 -1097 111 -1096
rect 1668 -1097 1669 -1096
rect 933 -1099 934 -1098
rect 975 -1099 976 -1098
rect 1024 -1099 1025 -1098
rect 1171 -1099 1172 -1098
rect 1318 -1099 1319 -1098
rect 1325 -1099 1326 -1098
rect 1402 -1099 1403 -1098
rect 1486 -1099 1487 -1098
rect 572 -1101 573 -1100
rect 933 -1101 934 -1100
rect 1080 -1101 1081 -1100
rect 1752 -1101 1753 -1100
rect 789 -1103 790 -1102
rect 1318 -1103 1319 -1102
rect 1486 -1103 1487 -1102
rect 1881 -1103 1882 -1102
rect 814 -1105 815 -1104
rect 1171 -1105 1172 -1104
rect 814 -1107 815 -1106
rect 943 -1107 944 -1106
rect 1080 -1107 1081 -1106
rect 1902 -1107 1903 -1106
rect 2 -1118 3 -1117
rect 72 -1118 73 -1117
rect 128 -1118 129 -1117
rect 674 -1118 675 -1117
rect 716 -1118 717 -1117
rect 929 -1118 930 -1117
rect 933 -1118 934 -1117
rect 1150 -1118 1151 -1117
rect 1153 -1118 1154 -1117
rect 1829 -1118 1830 -1117
rect 1843 -1118 1844 -1117
rect 1867 -1118 1868 -1117
rect 1878 -1118 1879 -1117
rect 1920 -1118 1921 -1117
rect 1948 -1118 1949 -1117
rect 1955 -1118 1956 -1117
rect 1976 -1118 1977 -1117
rect 1990 -1118 1991 -1117
rect 16 -1120 17 -1119
rect 222 -1120 223 -1119
rect 233 -1120 234 -1119
rect 653 -1120 654 -1119
rect 656 -1120 657 -1119
rect 772 -1120 773 -1119
rect 775 -1120 776 -1119
rect 870 -1120 871 -1119
rect 880 -1120 881 -1119
rect 1367 -1120 1368 -1119
rect 1549 -1120 1550 -1119
rect 1892 -1120 1893 -1119
rect 1969 -1120 1970 -1119
rect 1976 -1120 1977 -1119
rect 16 -1122 17 -1121
rect 114 -1122 115 -1121
rect 135 -1122 136 -1121
rect 772 -1122 773 -1121
rect 779 -1122 780 -1121
rect 856 -1122 857 -1121
rect 866 -1122 867 -1121
rect 1024 -1122 1025 -1121
rect 1045 -1122 1046 -1121
rect 1199 -1122 1200 -1121
rect 1318 -1122 1319 -1121
rect 1906 -1122 1907 -1121
rect 1962 -1122 1963 -1121
rect 1969 -1122 1970 -1121
rect 23 -1124 24 -1123
rect 565 -1124 566 -1123
rect 572 -1124 573 -1123
rect 660 -1124 661 -1123
rect 674 -1124 675 -1123
rect 702 -1124 703 -1123
rect 716 -1124 717 -1123
rect 1080 -1124 1081 -1123
rect 1132 -1124 1133 -1123
rect 1570 -1124 1571 -1123
rect 1584 -1124 1585 -1123
rect 1885 -1124 1886 -1123
rect 30 -1126 31 -1125
rect 40 -1126 41 -1125
rect 44 -1126 45 -1125
rect 933 -1126 934 -1125
rect 957 -1126 958 -1125
rect 1703 -1126 1704 -1125
rect 1759 -1126 1760 -1125
rect 1878 -1126 1879 -1125
rect 30 -1128 31 -1127
rect 198 -1128 199 -1127
rect 219 -1128 220 -1127
rect 534 -1128 535 -1127
rect 562 -1128 563 -1127
rect 842 -1128 843 -1127
rect 870 -1128 871 -1127
rect 1290 -1128 1291 -1127
rect 1311 -1128 1312 -1127
rect 1318 -1128 1319 -1127
rect 1367 -1128 1368 -1127
rect 1388 -1128 1389 -1127
rect 1451 -1128 1452 -1127
rect 1570 -1128 1571 -1127
rect 1591 -1128 1592 -1127
rect 1759 -1128 1760 -1127
rect 1780 -1128 1781 -1127
rect 1899 -1128 1900 -1127
rect 61 -1130 62 -1129
rect 268 -1130 269 -1129
rect 282 -1130 283 -1129
rect 754 -1130 755 -1129
rect 758 -1130 759 -1129
rect 1003 -1130 1004 -1129
rect 1010 -1130 1011 -1129
rect 1024 -1130 1025 -1129
rect 1045 -1130 1046 -1129
rect 1731 -1130 1732 -1129
rect 1780 -1130 1781 -1129
rect 1787 -1130 1788 -1129
rect 1808 -1130 1809 -1129
rect 1829 -1130 1830 -1129
rect 1836 -1130 1837 -1129
rect 1843 -1130 1844 -1129
rect 1871 -1130 1872 -1129
rect 1962 -1130 1963 -1129
rect 65 -1132 66 -1131
rect 527 -1132 528 -1131
rect 562 -1132 563 -1131
rect 1230 -1132 1231 -1131
rect 1360 -1132 1361 -1131
rect 1388 -1132 1389 -1131
rect 1500 -1132 1501 -1131
rect 1549 -1132 1550 -1131
rect 1591 -1132 1592 -1131
rect 1598 -1132 1599 -1131
rect 1689 -1132 1690 -1131
rect 1731 -1132 1732 -1131
rect 1787 -1132 1788 -1131
rect 1801 -1132 1802 -1131
rect 1822 -1132 1823 -1131
rect 1864 -1132 1865 -1131
rect 65 -1134 66 -1133
rect 415 -1134 416 -1133
rect 422 -1134 423 -1133
rect 453 -1134 454 -1133
rect 464 -1134 465 -1133
rect 681 -1134 682 -1133
rect 695 -1134 696 -1133
rect 702 -1134 703 -1133
rect 730 -1134 731 -1133
rect 747 -1134 748 -1133
rect 751 -1134 752 -1133
rect 1451 -1134 1452 -1133
rect 1458 -1134 1459 -1133
rect 1500 -1134 1501 -1133
rect 1542 -1134 1543 -1133
rect 1871 -1134 1872 -1133
rect 72 -1136 73 -1135
rect 394 -1136 395 -1135
rect 415 -1136 416 -1135
rect 586 -1136 587 -1135
rect 625 -1136 626 -1135
rect 653 -1136 654 -1135
rect 660 -1136 661 -1135
rect 975 -1136 976 -1135
rect 996 -1136 997 -1135
rect 1010 -1136 1011 -1135
rect 1017 -1136 1018 -1135
rect 1577 -1136 1578 -1135
rect 1598 -1136 1599 -1135
rect 1612 -1136 1613 -1135
rect 1682 -1136 1683 -1135
rect 1822 -1136 1823 -1135
rect 100 -1138 101 -1137
rect 128 -1138 129 -1137
rect 131 -1138 132 -1137
rect 681 -1138 682 -1137
rect 695 -1138 696 -1137
rect 723 -1138 724 -1137
rect 730 -1138 731 -1137
rect 765 -1138 766 -1137
rect 782 -1138 783 -1137
rect 1262 -1138 1263 -1137
rect 1423 -1138 1424 -1137
rect 1682 -1138 1683 -1137
rect 1696 -1138 1697 -1137
rect 1836 -1138 1837 -1137
rect 9 -1140 10 -1139
rect 100 -1140 101 -1139
rect 114 -1140 115 -1139
rect 789 -1140 790 -1139
rect 810 -1140 811 -1139
rect 1031 -1140 1032 -1139
rect 1080 -1140 1081 -1139
rect 1101 -1140 1102 -1139
rect 1139 -1140 1140 -1139
rect 1192 -1140 1193 -1139
rect 1402 -1140 1403 -1139
rect 1423 -1140 1424 -1139
rect 1458 -1140 1459 -1139
rect 1486 -1140 1487 -1139
rect 1493 -1140 1494 -1139
rect 1542 -1140 1543 -1139
rect 1563 -1140 1564 -1139
rect 1577 -1140 1578 -1139
rect 1605 -1140 1606 -1139
rect 1689 -1140 1690 -1139
rect 1724 -1140 1725 -1139
rect 1864 -1140 1865 -1139
rect 9 -1142 10 -1141
rect 425 -1142 426 -1141
rect 429 -1142 430 -1141
rect 856 -1142 857 -1141
rect 859 -1142 860 -1141
rect 1262 -1142 1263 -1141
rect 1381 -1142 1382 -1141
rect 1402 -1142 1403 -1141
rect 1444 -1142 1445 -1141
rect 1493 -1142 1494 -1141
rect 1521 -1142 1522 -1141
rect 1696 -1142 1697 -1141
rect 1794 -1142 1795 -1141
rect 1808 -1142 1809 -1141
rect 79 -1144 80 -1143
rect 1563 -1144 1564 -1143
rect 1605 -1144 1606 -1143
rect 1626 -1144 1627 -1143
rect 1668 -1144 1669 -1143
rect 1724 -1144 1725 -1143
rect 1752 -1144 1753 -1143
rect 1794 -1144 1795 -1143
rect 121 -1146 122 -1145
rect 135 -1146 136 -1145
rect 159 -1146 160 -1145
rect 310 -1146 311 -1145
rect 331 -1146 332 -1145
rect 534 -1146 535 -1145
rect 555 -1146 556 -1145
rect 625 -1146 626 -1145
rect 723 -1146 724 -1145
rect 744 -1146 745 -1145
rect 761 -1146 762 -1145
rect 1290 -1146 1291 -1145
rect 1444 -1146 1445 -1145
rect 1479 -1146 1480 -1145
rect 1486 -1146 1487 -1145
rect 1556 -1146 1557 -1145
rect 1612 -1146 1613 -1145
rect 1633 -1146 1634 -1145
rect 1668 -1146 1669 -1145
rect 1815 -1146 1816 -1145
rect 121 -1148 122 -1147
rect 782 -1148 783 -1147
rect 814 -1148 815 -1147
rect 842 -1148 843 -1147
rect 863 -1148 864 -1147
rect 1381 -1148 1382 -1147
rect 1437 -1148 1438 -1147
rect 1479 -1148 1480 -1147
rect 1507 -1148 1508 -1147
rect 1556 -1148 1557 -1147
rect 1626 -1148 1627 -1147
rect 1640 -1148 1641 -1147
rect 1745 -1148 1746 -1147
rect 1752 -1148 1753 -1147
rect 180 -1150 181 -1149
rect 852 -1150 853 -1149
rect 863 -1150 864 -1149
rect 877 -1150 878 -1149
rect 894 -1150 895 -1149
rect 1647 -1150 1648 -1149
rect 1717 -1150 1718 -1149
rect 1745 -1150 1746 -1149
rect 198 -1152 199 -1151
rect 317 -1152 318 -1151
rect 359 -1152 360 -1151
rect 628 -1152 629 -1151
rect 670 -1152 671 -1151
rect 1507 -1152 1508 -1151
rect 1514 -1152 1515 -1151
rect 1640 -1152 1641 -1151
rect 1647 -1152 1648 -1151
rect 1675 -1152 1676 -1151
rect 1717 -1152 1718 -1151
rect 1738 -1152 1739 -1151
rect 82 -1154 83 -1153
rect 317 -1154 318 -1153
rect 359 -1154 360 -1153
rect 380 -1154 381 -1153
rect 422 -1154 423 -1153
rect 1129 -1154 1130 -1153
rect 1136 -1154 1137 -1153
rect 1675 -1154 1676 -1153
rect 1710 -1154 1711 -1153
rect 1738 -1154 1739 -1153
rect 233 -1156 234 -1155
rect 247 -1156 248 -1155
rect 261 -1156 262 -1155
rect 292 -1156 293 -1155
rect 303 -1156 304 -1155
rect 331 -1156 332 -1155
rect 366 -1156 367 -1155
rect 369 -1156 370 -1155
rect 373 -1156 374 -1155
rect 394 -1156 395 -1155
rect 436 -1156 437 -1155
rect 523 -1156 524 -1155
rect 555 -1156 556 -1155
rect 667 -1156 668 -1155
rect 684 -1156 685 -1155
rect 1815 -1156 1816 -1155
rect 51 -1158 52 -1157
rect 373 -1158 374 -1157
rect 380 -1158 381 -1157
rect 800 -1158 801 -1157
rect 873 -1158 874 -1157
rect 1584 -1158 1585 -1157
rect 1633 -1158 1634 -1157
rect 1661 -1158 1662 -1157
rect 51 -1160 52 -1159
rect 740 -1160 741 -1159
rect 779 -1160 780 -1159
rect 1437 -1160 1438 -1159
rect 1465 -1160 1466 -1159
rect 1514 -1160 1515 -1159
rect 1521 -1160 1522 -1159
rect 1654 -1160 1655 -1159
rect 240 -1162 241 -1161
rect 247 -1162 248 -1161
rect 268 -1162 269 -1161
rect 275 -1162 276 -1161
rect 282 -1162 283 -1161
rect 345 -1162 346 -1161
rect 366 -1162 367 -1161
rect 387 -1162 388 -1161
rect 436 -1162 437 -1161
rect 912 -1162 913 -1161
rect 926 -1162 927 -1161
rect 1360 -1162 1361 -1161
rect 1472 -1162 1473 -1161
rect 1654 -1162 1655 -1161
rect 163 -1164 164 -1163
rect 345 -1164 346 -1163
rect 352 -1164 353 -1163
rect 926 -1164 927 -1163
rect 975 -1164 976 -1163
rect 982 -1164 983 -1163
rect 989 -1164 990 -1163
rect 996 -1164 997 -1163
rect 1003 -1164 1004 -1163
rect 1220 -1164 1221 -1163
rect 1248 -1164 1249 -1163
rect 1472 -1164 1473 -1163
rect 1535 -1164 1536 -1163
rect 1661 -1164 1662 -1163
rect 58 -1166 59 -1165
rect 352 -1166 353 -1165
rect 446 -1166 447 -1165
rect 1703 -1166 1704 -1165
rect 163 -1168 164 -1167
rect 457 -1168 458 -1167
rect 464 -1168 465 -1167
rect 541 -1168 542 -1167
rect 583 -1168 584 -1167
rect 786 -1168 787 -1167
rect 912 -1168 913 -1167
rect 1129 -1168 1130 -1167
rect 1160 -1168 1161 -1167
rect 1913 -1168 1914 -1167
rect 142 -1170 143 -1169
rect 541 -1170 542 -1169
rect 583 -1170 584 -1169
rect 1031 -1170 1032 -1169
rect 1038 -1170 1039 -1169
rect 1220 -1170 1221 -1169
rect 1241 -1170 1242 -1169
rect 1248 -1170 1249 -1169
rect 142 -1172 143 -1171
rect 229 -1172 230 -1171
rect 240 -1172 241 -1171
rect 296 -1172 297 -1171
rect 303 -1172 304 -1171
rect 908 -1172 909 -1171
rect 961 -1172 962 -1171
rect 989 -1172 990 -1171
rect 1017 -1172 1018 -1171
rect 1465 -1172 1466 -1171
rect 254 -1174 255 -1173
rect 296 -1174 297 -1173
rect 313 -1174 314 -1173
rect 1136 -1174 1137 -1173
rect 1164 -1174 1165 -1173
rect 1192 -1174 1193 -1173
rect 1234 -1174 1235 -1173
rect 1241 -1174 1242 -1173
rect 212 -1176 213 -1175
rect 254 -1176 255 -1175
rect 275 -1176 276 -1175
rect 338 -1176 339 -1175
rect 450 -1176 451 -1175
rect 1801 -1176 1802 -1175
rect 37 -1178 38 -1177
rect 450 -1178 451 -1177
rect 453 -1178 454 -1177
rect 1199 -1178 1200 -1177
rect 1213 -1178 1214 -1177
rect 1234 -1178 1235 -1177
rect 289 -1180 290 -1179
rect 576 -1180 577 -1179
rect 590 -1180 591 -1179
rect 814 -1180 815 -1179
rect 849 -1180 850 -1179
rect 1038 -1180 1039 -1179
rect 1048 -1180 1049 -1179
rect 1710 -1180 1711 -1179
rect 107 -1182 108 -1181
rect 1048 -1182 1049 -1181
rect 1087 -1182 1088 -1181
rect 1311 -1182 1312 -1181
rect 107 -1184 108 -1183
rect 891 -1184 892 -1183
rect 982 -1184 983 -1183
rect 1052 -1184 1053 -1183
rect 1059 -1184 1060 -1183
rect 1087 -1184 1088 -1183
rect 1094 -1184 1095 -1183
rect 1101 -1184 1102 -1183
rect 1115 -1184 1116 -1183
rect 1164 -1184 1165 -1183
rect 156 -1186 157 -1185
rect 590 -1186 591 -1185
rect 632 -1186 633 -1185
rect 1535 -1186 1536 -1185
rect 324 -1188 325 -1187
rect 632 -1188 633 -1187
rect 667 -1188 668 -1187
rect 1528 -1188 1529 -1187
rect 324 -1190 325 -1189
rect 485 -1190 486 -1189
rect 516 -1190 517 -1189
rect 1227 -1190 1228 -1189
rect 338 -1192 339 -1191
rect 604 -1192 605 -1191
rect 709 -1192 710 -1191
rect 800 -1192 801 -1191
rect 821 -1192 822 -1191
rect 849 -1192 850 -1191
rect 877 -1192 878 -1191
rect 1059 -1192 1060 -1191
rect 1108 -1192 1109 -1191
rect 1115 -1192 1116 -1191
rect 1157 -1192 1158 -1191
rect 1213 -1192 1214 -1191
rect 37 -1194 38 -1193
rect 604 -1194 605 -1193
rect 709 -1194 710 -1193
rect 807 -1194 808 -1193
rect 891 -1194 892 -1193
rect 898 -1194 899 -1193
rect 1052 -1194 1053 -1193
rect 1066 -1194 1067 -1193
rect 1108 -1194 1109 -1193
rect 1283 -1194 1284 -1193
rect 408 -1196 409 -1195
rect 1283 -1196 1284 -1195
rect 408 -1198 409 -1197
rect 688 -1198 689 -1197
rect 733 -1198 734 -1197
rect 1850 -1198 1851 -1197
rect 443 -1200 444 -1199
rect 1094 -1200 1095 -1199
rect 1157 -1200 1158 -1199
rect 1409 -1200 1410 -1199
rect 212 -1202 213 -1201
rect 443 -1202 444 -1201
rect 457 -1202 458 -1201
rect 506 -1202 507 -1201
rect 576 -1202 577 -1201
rect 618 -1202 619 -1201
rect 737 -1202 738 -1201
rect 1178 -1202 1179 -1201
rect 1181 -1202 1182 -1201
rect 1850 -1202 1851 -1201
rect 44 -1204 45 -1203
rect 1178 -1204 1179 -1203
rect 1185 -1204 1186 -1203
rect 1528 -1204 1529 -1203
rect 289 -1206 290 -1205
rect 618 -1206 619 -1205
rect 744 -1206 745 -1205
rect 821 -1206 822 -1205
rect 898 -1206 899 -1205
rect 905 -1206 906 -1205
rect 1066 -1206 1067 -1205
rect 1073 -1206 1074 -1205
rect 1143 -1206 1144 -1205
rect 1185 -1206 1186 -1205
rect 1395 -1206 1396 -1205
rect 1409 -1206 1410 -1205
rect 471 -1208 472 -1207
rect 527 -1208 528 -1207
rect 611 -1208 612 -1207
rect 688 -1208 689 -1207
rect 747 -1208 748 -1207
rect 765 -1208 766 -1207
rect 807 -1208 808 -1207
rect 954 -1208 955 -1207
rect 1143 -1208 1144 -1207
rect 1255 -1208 1256 -1207
rect 1374 -1208 1375 -1207
rect 1395 -1208 1396 -1207
rect 429 -1210 430 -1209
rect 471 -1210 472 -1209
rect 474 -1210 475 -1209
rect 499 -1210 500 -1209
rect 506 -1210 507 -1209
rect 639 -1210 640 -1209
rect 905 -1210 906 -1209
rect 1857 -1210 1858 -1209
rect 124 -1212 125 -1211
rect 499 -1212 500 -1211
rect 513 -1212 514 -1211
rect 737 -1212 738 -1211
rect 940 -1212 941 -1211
rect 1073 -1212 1074 -1211
rect 1255 -1212 1256 -1211
rect 1339 -1212 1340 -1211
rect 1353 -1212 1354 -1211
rect 1374 -1212 1375 -1211
rect 1619 -1212 1620 -1211
rect 1857 -1212 1858 -1211
rect 82 -1214 83 -1213
rect 1619 -1214 1620 -1213
rect 478 -1216 479 -1215
rect 751 -1216 752 -1215
rect 940 -1216 941 -1215
rect 964 -1216 965 -1215
rect 1325 -1216 1326 -1215
rect 1339 -1216 1340 -1215
rect 1346 -1216 1347 -1215
rect 1353 -1216 1354 -1215
rect 177 -1218 178 -1217
rect 478 -1218 479 -1217
rect 485 -1218 486 -1217
rect 548 -1218 549 -1217
rect 579 -1218 580 -1217
rect 611 -1218 612 -1217
rect 947 -1218 948 -1217
rect 954 -1218 955 -1217
rect 1297 -1218 1298 -1217
rect 1325 -1218 1326 -1217
rect 1332 -1218 1333 -1217
rect 1346 -1218 1347 -1217
rect 177 -1220 178 -1219
rect 1171 -1220 1172 -1219
rect 1297 -1220 1298 -1219
rect 1304 -1220 1305 -1219
rect 520 -1222 521 -1221
rect 1171 -1222 1172 -1221
rect 1304 -1222 1305 -1221
rect 1430 -1222 1431 -1221
rect 93 -1224 94 -1223
rect 520 -1224 521 -1223
rect 548 -1224 549 -1223
rect 968 -1224 969 -1223
rect 1416 -1224 1417 -1223
rect 1430 -1224 1431 -1223
rect 47 -1226 48 -1225
rect 1416 -1226 1417 -1225
rect 93 -1228 94 -1227
rect 149 -1228 150 -1227
rect 569 -1228 570 -1227
rect 1332 -1228 1333 -1227
rect 149 -1230 150 -1229
rect 205 -1230 206 -1229
rect 492 -1230 493 -1229
rect 569 -1230 570 -1229
rect 597 -1230 598 -1229
rect 639 -1230 640 -1229
rect 828 -1230 829 -1229
rect 968 -1230 969 -1229
rect 58 -1232 59 -1231
rect 597 -1232 598 -1231
rect 828 -1232 829 -1231
rect 884 -1232 885 -1231
rect 919 -1232 920 -1231
rect 947 -1232 948 -1231
rect 191 -1234 192 -1233
rect 205 -1234 206 -1233
rect 492 -1234 493 -1233
rect 1020 -1234 1021 -1233
rect 170 -1236 171 -1235
rect 191 -1236 192 -1235
rect 646 -1236 647 -1235
rect 919 -1236 920 -1235
rect 170 -1238 171 -1237
rect 646 -1238 647 -1237
rect 835 -1238 836 -1237
rect 884 -1238 885 -1237
rect 793 -1240 794 -1239
rect 835 -1240 836 -1239
rect 226 -1242 227 -1241
rect 793 -1242 794 -1241
rect 23 -1253 24 -1252
rect 93 -1253 94 -1252
rect 107 -1253 108 -1252
rect 145 -1253 146 -1252
rect 163 -1253 164 -1252
rect 226 -1253 227 -1252
rect 247 -1253 248 -1252
rect 261 -1253 262 -1252
rect 282 -1253 283 -1252
rect 453 -1253 454 -1252
rect 457 -1253 458 -1252
rect 670 -1253 671 -1252
rect 688 -1253 689 -1252
rect 779 -1253 780 -1252
rect 793 -1253 794 -1252
rect 1076 -1253 1077 -1252
rect 1111 -1253 1112 -1252
rect 1878 -1253 1879 -1252
rect 1906 -1253 1907 -1252
rect 1948 -1253 1949 -1252
rect 1962 -1253 1963 -1252
rect 1997 -1253 1998 -1252
rect 30 -1255 31 -1254
rect 446 -1255 447 -1254
rect 457 -1255 458 -1254
rect 597 -1255 598 -1254
rect 628 -1255 629 -1254
rect 786 -1255 787 -1254
rect 821 -1255 822 -1254
rect 1066 -1255 1067 -1254
rect 1129 -1255 1130 -1254
rect 1822 -1255 1823 -1254
rect 1843 -1255 1844 -1254
rect 1906 -1255 1907 -1254
rect 1913 -1255 1914 -1254
rect 1941 -1255 1942 -1254
rect 1976 -1255 1977 -1254
rect 1983 -1255 1984 -1254
rect 30 -1257 31 -1256
rect 208 -1257 209 -1256
rect 226 -1257 227 -1256
rect 513 -1257 514 -1256
rect 541 -1257 542 -1256
rect 597 -1257 598 -1256
rect 604 -1257 605 -1256
rect 821 -1257 822 -1256
rect 838 -1257 839 -1256
rect 1472 -1257 1473 -1256
rect 1675 -1257 1676 -1256
rect 1843 -1257 1844 -1256
rect 1920 -1257 1921 -1256
rect 1934 -1257 1935 -1256
rect 1955 -1257 1956 -1256
rect 1976 -1257 1977 -1256
rect 37 -1259 38 -1258
rect 44 -1259 45 -1258
rect 58 -1259 59 -1258
rect 793 -1259 794 -1258
rect 856 -1259 857 -1258
rect 1759 -1259 1760 -1258
rect 40 -1261 41 -1260
rect 1654 -1261 1655 -1260
rect 1759 -1261 1760 -1260
rect 1913 -1261 1914 -1260
rect 44 -1263 45 -1262
rect 576 -1263 577 -1262
rect 586 -1263 587 -1262
rect 849 -1263 850 -1262
rect 856 -1263 857 -1262
rect 873 -1263 874 -1262
rect 908 -1263 909 -1262
rect 1220 -1263 1221 -1262
rect 1269 -1263 1270 -1262
rect 1272 -1263 1273 -1262
rect 1290 -1263 1291 -1262
rect 1920 -1263 1921 -1262
rect 58 -1265 59 -1264
rect 1857 -1265 1858 -1264
rect 61 -1267 62 -1266
rect 1521 -1267 1522 -1266
rect 1612 -1267 1613 -1266
rect 1654 -1267 1655 -1266
rect 1787 -1267 1788 -1266
rect 1857 -1267 1858 -1266
rect 65 -1269 66 -1268
rect 282 -1269 283 -1268
rect 289 -1269 290 -1268
rect 401 -1269 402 -1268
rect 415 -1269 416 -1268
rect 513 -1269 514 -1268
rect 562 -1269 563 -1268
rect 1073 -1269 1074 -1268
rect 1129 -1269 1130 -1268
rect 1136 -1269 1137 -1268
rect 1178 -1269 1179 -1268
rect 1885 -1269 1886 -1268
rect 51 -1271 52 -1270
rect 65 -1271 66 -1270
rect 79 -1271 80 -1270
rect 338 -1271 339 -1270
rect 352 -1271 353 -1270
rect 656 -1271 657 -1270
rect 688 -1271 689 -1270
rect 723 -1271 724 -1270
rect 775 -1271 776 -1270
rect 1850 -1271 1851 -1270
rect 9 -1273 10 -1272
rect 79 -1273 80 -1272
rect 82 -1273 83 -1272
rect 604 -1273 605 -1272
rect 646 -1273 647 -1272
rect 1132 -1273 1133 -1272
rect 1171 -1273 1172 -1272
rect 1178 -1273 1179 -1272
rect 1220 -1273 1221 -1272
rect 1234 -1273 1235 -1272
rect 1269 -1273 1270 -1272
rect 1276 -1273 1277 -1272
rect 1290 -1273 1291 -1272
rect 1297 -1273 1298 -1272
rect 1388 -1273 1389 -1272
rect 1391 -1273 1392 -1272
rect 1458 -1273 1459 -1272
rect 1472 -1273 1473 -1272
rect 1542 -1273 1543 -1272
rect 1612 -1273 1613 -1272
rect 1626 -1273 1627 -1272
rect 1675 -1273 1676 -1272
rect 1787 -1273 1788 -1272
rect 1916 -1273 1917 -1272
rect 9 -1275 10 -1274
rect 800 -1275 801 -1274
rect 824 -1275 825 -1274
rect 849 -1275 850 -1274
rect 870 -1275 871 -1274
rect 912 -1275 913 -1274
rect 922 -1275 923 -1274
rect 1892 -1275 1893 -1274
rect 2 -1277 3 -1276
rect 800 -1277 801 -1276
rect 912 -1277 913 -1276
rect 1108 -1277 1109 -1276
rect 1122 -1277 1123 -1276
rect 1136 -1277 1137 -1276
rect 1171 -1277 1172 -1276
rect 1521 -1277 1522 -1276
rect 1808 -1277 1809 -1276
rect 1850 -1277 1851 -1276
rect 86 -1279 87 -1278
rect 170 -1279 171 -1278
rect 177 -1279 178 -1278
rect 611 -1279 612 -1278
rect 681 -1279 682 -1278
rect 723 -1279 724 -1278
rect 779 -1279 780 -1278
rect 1069 -1279 1070 -1278
rect 1073 -1279 1074 -1278
rect 1661 -1279 1662 -1278
rect 1829 -1279 1830 -1278
rect 1885 -1279 1886 -1278
rect 54 -1281 55 -1280
rect 86 -1281 87 -1280
rect 93 -1281 94 -1280
rect 142 -1281 143 -1280
rect 149 -1281 150 -1280
rect 177 -1281 178 -1280
rect 247 -1281 248 -1280
rect 1094 -1281 1095 -1280
rect 1234 -1281 1235 -1280
rect 1262 -1281 1263 -1280
rect 1297 -1281 1298 -1280
rect 1332 -1281 1333 -1280
rect 1388 -1281 1389 -1280
rect 1409 -1281 1410 -1280
rect 1437 -1281 1438 -1280
rect 1458 -1281 1459 -1280
rect 1486 -1281 1487 -1280
rect 1626 -1281 1627 -1280
rect 1773 -1281 1774 -1280
rect 1829 -1281 1830 -1280
rect 107 -1283 108 -1282
rect 548 -1283 549 -1282
rect 611 -1283 612 -1282
rect 618 -1283 619 -1282
rect 653 -1283 654 -1282
rect 681 -1283 682 -1282
rect 877 -1283 878 -1282
rect 1122 -1283 1123 -1282
rect 1143 -1283 1144 -1282
rect 1262 -1283 1263 -1282
rect 1416 -1283 1417 -1282
rect 1437 -1283 1438 -1282
rect 1479 -1283 1480 -1282
rect 1486 -1283 1487 -1282
rect 1493 -1283 1494 -1282
rect 1542 -1283 1543 -1282
rect 1591 -1283 1592 -1282
rect 1661 -1283 1662 -1282
rect 1745 -1283 1746 -1282
rect 1773 -1283 1774 -1282
rect 110 -1285 111 -1284
rect 1822 -1285 1823 -1284
rect 121 -1287 122 -1286
rect 229 -1287 230 -1286
rect 254 -1287 255 -1286
rect 579 -1287 580 -1286
rect 618 -1287 619 -1286
rect 891 -1287 892 -1286
rect 926 -1287 927 -1286
rect 1878 -1287 1879 -1286
rect 152 -1289 153 -1288
rect 261 -1289 262 -1288
rect 296 -1289 297 -1288
rect 299 -1289 300 -1288
rect 317 -1289 318 -1288
rect 541 -1289 542 -1288
rect 548 -1289 549 -1288
rect 940 -1289 941 -1288
rect 964 -1289 965 -1288
rect 1682 -1289 1683 -1288
rect 156 -1291 157 -1290
rect 1892 -1291 1893 -1290
rect 156 -1293 157 -1292
rect 660 -1293 661 -1292
rect 712 -1293 713 -1292
rect 1682 -1293 1683 -1292
rect 128 -1295 129 -1294
rect 660 -1295 661 -1294
rect 877 -1295 878 -1294
rect 1024 -1295 1025 -1294
rect 1038 -1295 1039 -1294
rect 1157 -1295 1158 -1294
rect 1244 -1295 1245 -1294
rect 1493 -1295 1494 -1294
rect 1563 -1295 1564 -1294
rect 1591 -1295 1592 -1294
rect 1605 -1295 1606 -1294
rect 1745 -1295 1746 -1294
rect 75 -1297 76 -1296
rect 1024 -1297 1025 -1296
rect 1045 -1297 1046 -1296
rect 1087 -1297 1088 -1296
rect 1094 -1297 1095 -1296
rect 1115 -1297 1116 -1296
rect 1143 -1297 1144 -1296
rect 1185 -1297 1186 -1296
rect 1255 -1297 1256 -1296
rect 1332 -1297 1333 -1296
rect 1416 -1297 1417 -1296
rect 1423 -1297 1424 -1296
rect 1465 -1297 1466 -1296
rect 1479 -1297 1480 -1296
rect 124 -1299 125 -1298
rect 1087 -1299 1088 -1298
rect 1185 -1299 1186 -1298
rect 1836 -1299 1837 -1298
rect 128 -1301 129 -1300
rect 842 -1301 843 -1300
rect 891 -1301 892 -1300
rect 947 -1301 948 -1300
rect 961 -1301 962 -1300
rect 1038 -1301 1039 -1300
rect 1055 -1301 1056 -1300
rect 1808 -1301 1809 -1300
rect 163 -1303 164 -1302
rect 240 -1303 241 -1302
rect 254 -1303 255 -1302
rect 670 -1303 671 -1302
rect 842 -1303 843 -1302
rect 898 -1303 899 -1302
rect 929 -1303 930 -1302
rect 1605 -1303 1606 -1302
rect 1780 -1303 1781 -1302
rect 1836 -1303 1837 -1302
rect 170 -1305 171 -1304
rect 380 -1305 381 -1304
rect 394 -1305 395 -1304
rect 425 -1305 426 -1304
rect 443 -1305 444 -1304
rect 1311 -1305 1312 -1304
rect 1423 -1305 1424 -1304
rect 1507 -1305 1508 -1304
rect 1766 -1305 1767 -1304
rect 1780 -1305 1781 -1304
rect 205 -1307 206 -1306
rect 240 -1307 241 -1306
rect 268 -1307 269 -1306
rect 394 -1307 395 -1306
rect 401 -1307 402 -1306
rect 555 -1307 556 -1306
rect 807 -1307 808 -1306
rect 898 -1307 899 -1306
rect 929 -1307 930 -1306
rect 1563 -1307 1564 -1306
rect 1752 -1307 1753 -1306
rect 1766 -1307 1767 -1306
rect 184 -1309 185 -1308
rect 205 -1309 206 -1308
rect 233 -1309 234 -1308
rect 268 -1309 269 -1308
rect 296 -1309 297 -1308
rect 331 -1309 332 -1308
rect 338 -1309 339 -1308
rect 408 -1309 409 -1308
rect 422 -1309 423 -1308
rect 1801 -1309 1802 -1308
rect 184 -1311 185 -1310
rect 303 -1311 304 -1310
rect 310 -1311 311 -1310
rect 555 -1311 556 -1310
rect 807 -1311 808 -1310
rect 1080 -1311 1081 -1310
rect 1108 -1311 1109 -1310
rect 1507 -1311 1508 -1310
rect 1696 -1311 1697 -1310
rect 1752 -1311 1753 -1310
rect 100 -1313 101 -1312
rect 310 -1313 311 -1312
rect 317 -1313 318 -1312
rect 387 -1313 388 -1312
rect 408 -1313 409 -1312
rect 520 -1313 521 -1312
rect 534 -1313 535 -1312
rect 562 -1313 563 -1312
rect 810 -1313 811 -1312
rect 1801 -1313 1802 -1312
rect 72 -1315 73 -1314
rect 387 -1315 388 -1314
rect 422 -1315 423 -1314
rect 667 -1315 668 -1314
rect 947 -1315 948 -1314
rect 954 -1315 955 -1314
rect 961 -1315 962 -1314
rect 989 -1315 990 -1314
rect 1017 -1315 1018 -1314
rect 1871 -1315 1872 -1314
rect 51 -1317 52 -1316
rect 667 -1317 668 -1316
rect 954 -1317 955 -1316
rect 975 -1317 976 -1316
rect 989 -1317 990 -1316
rect 1031 -1317 1032 -1316
rect 1066 -1317 1067 -1316
rect 1311 -1317 1312 -1316
rect 1391 -1317 1392 -1316
rect 1409 -1317 1410 -1316
rect 1451 -1317 1452 -1316
rect 1465 -1317 1466 -1316
rect 1668 -1317 1669 -1316
rect 1871 -1317 1872 -1316
rect 72 -1319 73 -1318
rect 569 -1319 570 -1318
rect 968 -1319 969 -1318
rect 1115 -1319 1116 -1318
rect 1255 -1319 1256 -1318
rect 1374 -1319 1375 -1318
rect 1598 -1319 1599 -1318
rect 1668 -1319 1669 -1318
rect 1696 -1319 1697 -1318
rect 1703 -1319 1704 -1318
rect 100 -1321 101 -1320
rect 264 -1321 265 -1320
rect 352 -1321 353 -1320
rect 359 -1321 360 -1320
rect 366 -1321 367 -1320
rect 380 -1321 381 -1320
rect 443 -1321 444 -1320
rect 772 -1321 773 -1320
rect 968 -1321 969 -1320
rect 1020 -1321 1021 -1320
rect 1031 -1321 1032 -1320
rect 1325 -1321 1326 -1320
rect 1360 -1321 1361 -1320
rect 1451 -1321 1452 -1320
rect 142 -1323 143 -1322
rect 303 -1323 304 -1322
rect 324 -1323 325 -1322
rect 359 -1323 360 -1322
rect 366 -1323 367 -1322
rect 516 -1323 517 -1322
rect 534 -1323 535 -1322
rect 765 -1323 766 -1322
rect 772 -1323 773 -1322
rect 814 -1323 815 -1322
rect 975 -1323 976 -1322
rect 982 -1323 983 -1322
rect 996 -1323 997 -1322
rect 1017 -1323 1018 -1322
rect 1080 -1323 1081 -1322
rect 1164 -1323 1165 -1322
rect 1304 -1323 1305 -1322
rect 1360 -1323 1361 -1322
rect 1374 -1323 1375 -1322
rect 1395 -1323 1396 -1322
rect 1444 -1323 1445 -1322
rect 1598 -1323 1599 -1322
rect 233 -1325 234 -1324
rect 492 -1325 493 -1324
rect 530 -1325 531 -1324
rect 1444 -1325 1445 -1324
rect 275 -1327 276 -1326
rect 324 -1327 325 -1326
rect 373 -1327 374 -1326
rect 415 -1327 416 -1326
rect 450 -1327 451 -1326
rect 814 -1327 815 -1326
rect 859 -1327 860 -1326
rect 1304 -1327 1305 -1326
rect 1325 -1327 1326 -1326
rect 1339 -1327 1340 -1326
rect 212 -1329 213 -1328
rect 275 -1329 276 -1328
rect 373 -1329 374 -1328
rect 677 -1329 678 -1328
rect 765 -1329 766 -1328
rect 835 -1329 836 -1328
rect 859 -1329 860 -1328
rect 1703 -1329 1704 -1328
rect 198 -1331 199 -1330
rect 212 -1331 213 -1330
rect 436 -1331 437 -1330
rect 450 -1331 451 -1330
rect 464 -1331 465 -1330
rect 646 -1331 647 -1330
rect 905 -1331 906 -1330
rect 982 -1331 983 -1330
rect 996 -1331 997 -1330
rect 1899 -1331 1900 -1330
rect 198 -1333 199 -1332
rect 639 -1333 640 -1332
rect 884 -1333 885 -1332
rect 905 -1333 906 -1332
rect 1164 -1333 1165 -1332
rect 1213 -1333 1214 -1332
rect 1227 -1333 1228 -1332
rect 1395 -1333 1396 -1332
rect 1864 -1333 1865 -1332
rect 1899 -1333 1900 -1332
rect 436 -1335 437 -1334
rect 758 -1335 759 -1334
rect 884 -1335 885 -1334
rect 919 -1335 920 -1334
rect 1059 -1335 1060 -1334
rect 1213 -1335 1214 -1334
rect 1227 -1335 1228 -1334
rect 1248 -1335 1249 -1334
rect 1318 -1335 1319 -1334
rect 1339 -1335 1340 -1334
rect 1815 -1335 1816 -1334
rect 1864 -1335 1865 -1334
rect 464 -1337 465 -1336
rect 716 -1337 717 -1336
rect 751 -1337 752 -1336
rect 758 -1337 759 -1336
rect 1052 -1337 1053 -1336
rect 1059 -1337 1060 -1336
rect 1248 -1337 1249 -1336
rect 1346 -1337 1347 -1336
rect 1794 -1337 1795 -1336
rect 1815 -1337 1816 -1336
rect 471 -1339 472 -1338
rect 1003 -1339 1004 -1338
rect 1318 -1339 1319 -1338
rect 1402 -1339 1403 -1338
rect 1647 -1339 1648 -1338
rect 1794 -1339 1795 -1338
rect 474 -1341 475 -1340
rect 625 -1341 626 -1340
rect 639 -1341 640 -1340
rect 674 -1341 675 -1340
rect 716 -1341 717 -1340
rect 737 -1341 738 -1340
rect 744 -1341 745 -1340
rect 751 -1341 752 -1340
rect 1003 -1341 1004 -1340
rect 1181 -1341 1182 -1340
rect 1346 -1341 1347 -1340
rect 1353 -1341 1354 -1340
rect 1647 -1341 1648 -1340
rect 1738 -1341 1739 -1340
rect 114 -1343 115 -1342
rect 674 -1343 675 -1342
rect 737 -1343 738 -1342
rect 1010 -1343 1011 -1342
rect 1052 -1343 1053 -1342
rect 1402 -1343 1403 -1342
rect 1717 -1343 1718 -1342
rect 1738 -1343 1739 -1342
rect 114 -1345 115 -1344
rect 345 -1345 346 -1344
rect 478 -1345 479 -1344
rect 520 -1345 521 -1344
rect 569 -1345 570 -1344
rect 709 -1345 710 -1344
rect 943 -1345 944 -1344
rect 1717 -1345 1718 -1344
rect 159 -1347 160 -1346
rect 345 -1347 346 -1346
rect 478 -1347 479 -1346
rect 499 -1347 500 -1346
rect 590 -1347 591 -1346
rect 835 -1347 836 -1346
rect 1353 -1347 1354 -1346
rect 1367 -1347 1368 -1346
rect 173 -1349 174 -1348
rect 1010 -1349 1011 -1348
rect 1367 -1349 1368 -1348
rect 1381 -1349 1382 -1348
rect 485 -1351 486 -1350
rect 583 -1351 584 -1350
rect 625 -1351 626 -1350
rect 695 -1351 696 -1350
rect 709 -1351 710 -1350
rect 786 -1351 787 -1350
rect 1241 -1351 1242 -1350
rect 1381 -1351 1382 -1350
rect 219 -1353 220 -1352
rect 695 -1353 696 -1352
rect 1241 -1353 1242 -1352
rect 1640 -1353 1641 -1352
rect 191 -1355 192 -1354
rect 219 -1355 220 -1354
rect 432 -1355 433 -1354
rect 583 -1355 584 -1354
rect 1556 -1355 1557 -1354
rect 1640 -1355 1641 -1354
rect 191 -1357 192 -1356
rect 565 -1357 566 -1356
rect 1535 -1357 1536 -1356
rect 1556 -1357 1557 -1356
rect 485 -1359 486 -1358
rect 702 -1359 703 -1358
rect 1528 -1359 1529 -1358
rect 1535 -1359 1536 -1358
rect 429 -1361 430 -1360
rect 702 -1361 703 -1360
rect 1514 -1361 1515 -1360
rect 1528 -1361 1529 -1360
rect 429 -1363 430 -1362
rect 1619 -1363 1620 -1362
rect 492 -1365 493 -1364
rect 506 -1365 507 -1364
rect 527 -1365 528 -1364
rect 590 -1365 591 -1364
rect 1500 -1365 1501 -1364
rect 1514 -1365 1515 -1364
rect 1570 -1365 1571 -1364
rect 1619 -1365 1620 -1364
rect 499 -1367 500 -1366
rect 933 -1367 934 -1366
rect 1500 -1367 1501 -1366
rect 1633 -1367 1634 -1366
rect 506 -1369 507 -1368
rect 632 -1369 633 -1368
rect 933 -1369 934 -1368
rect 999 -1369 1000 -1368
rect 1549 -1369 1550 -1368
rect 1570 -1369 1571 -1368
rect 1577 -1369 1578 -1368
rect 1633 -1369 1634 -1368
rect 527 -1371 528 -1370
rect 1283 -1371 1284 -1370
rect 1549 -1371 1550 -1370
rect 1731 -1371 1732 -1370
rect 632 -1373 633 -1372
rect 828 -1373 829 -1372
rect 919 -1373 920 -1372
rect 1577 -1373 1578 -1372
rect 1724 -1373 1725 -1372
rect 1731 -1373 1732 -1372
rect 744 -1375 745 -1374
rect 1283 -1375 1284 -1374
rect 1710 -1375 1711 -1374
rect 1724 -1375 1725 -1374
rect 828 -1377 829 -1376
rect 863 -1377 864 -1376
rect 1584 -1377 1585 -1376
rect 1710 -1377 1711 -1376
rect 653 -1379 654 -1378
rect 863 -1379 864 -1378
rect 1199 -1379 1200 -1378
rect 1584 -1379 1585 -1378
rect 1192 -1381 1193 -1380
rect 1199 -1381 1200 -1380
rect 1192 -1383 1193 -1382
rect 1206 -1383 1207 -1382
rect 180 -1385 181 -1384
rect 1206 -1385 1207 -1384
rect 2 -1396 3 -1395
rect 208 -1396 209 -1395
rect 485 -1396 486 -1395
rect 919 -1396 920 -1395
rect 940 -1396 941 -1395
rect 1647 -1396 1648 -1395
rect 1899 -1396 1900 -1395
rect 1962 -1396 1963 -1395
rect 1976 -1396 1977 -1395
rect 2025 -1396 2026 -1395
rect 9 -1398 10 -1397
rect 215 -1398 216 -1397
rect 485 -1398 486 -1397
rect 492 -1398 493 -1397
rect 527 -1398 528 -1397
rect 646 -1398 647 -1397
rect 674 -1398 675 -1397
rect 681 -1398 682 -1397
rect 712 -1398 713 -1397
rect 912 -1398 913 -1397
rect 947 -1398 948 -1397
rect 999 -1398 1000 -1397
rect 1003 -1398 1004 -1397
rect 1013 -1398 1014 -1397
rect 1038 -1398 1039 -1397
rect 1073 -1398 1074 -1397
rect 1104 -1398 1105 -1397
rect 1542 -1398 1543 -1397
rect 1647 -1398 1648 -1397
rect 1822 -1398 1823 -1397
rect 1913 -1398 1914 -1397
rect 1927 -1398 1928 -1397
rect 1941 -1398 1942 -1397
rect 2011 -1398 2012 -1397
rect 9 -1400 10 -1399
rect 261 -1400 262 -1399
rect 527 -1400 528 -1399
rect 922 -1400 923 -1399
rect 926 -1400 927 -1399
rect 1038 -1400 1039 -1399
rect 1052 -1400 1053 -1399
rect 1808 -1400 1809 -1399
rect 1822 -1400 1823 -1399
rect 1920 -1400 1921 -1399
rect 1948 -1400 1949 -1399
rect 1955 -1400 1956 -1399
rect 1983 -1400 1984 -1399
rect 1986 -1400 1987 -1399
rect 1997 -1400 1998 -1399
rect 2018 -1400 2019 -1399
rect 16 -1402 17 -1401
rect 152 -1402 153 -1401
rect 184 -1402 185 -1401
rect 1185 -1402 1186 -1401
rect 1241 -1402 1242 -1401
rect 1794 -1402 1795 -1401
rect 1843 -1402 1844 -1401
rect 1948 -1402 1949 -1401
rect 1983 -1402 1984 -1401
rect 1990 -1402 1991 -1401
rect 16 -1404 17 -1403
rect 121 -1404 122 -1403
rect 142 -1404 143 -1403
rect 1682 -1404 1683 -1403
rect 1780 -1404 1781 -1403
rect 1843 -1404 1844 -1403
rect 1864 -1404 1865 -1403
rect 1927 -1404 1928 -1403
rect 30 -1406 31 -1405
rect 957 -1406 958 -1405
rect 968 -1406 969 -1405
rect 1444 -1406 1445 -1405
rect 1577 -1406 1578 -1405
rect 1808 -1406 1809 -1405
rect 1864 -1406 1865 -1405
rect 1878 -1406 1879 -1405
rect 1916 -1406 1917 -1405
rect 1934 -1406 1935 -1405
rect 30 -1408 31 -1407
rect 618 -1408 619 -1407
rect 632 -1408 633 -1407
rect 667 -1408 668 -1407
rect 677 -1408 678 -1407
rect 961 -1408 962 -1407
rect 975 -1408 976 -1407
rect 1052 -1408 1053 -1407
rect 1055 -1408 1056 -1407
rect 1381 -1408 1382 -1407
rect 1444 -1408 1445 -1407
rect 1591 -1408 1592 -1407
rect 1605 -1408 1606 -1407
rect 1682 -1408 1683 -1407
rect 1738 -1408 1739 -1407
rect 1780 -1408 1781 -1407
rect 1787 -1408 1788 -1407
rect 1878 -1408 1879 -1407
rect 1885 -1408 1886 -1407
rect 1934 -1408 1935 -1407
rect 47 -1410 48 -1409
rect 1542 -1410 1543 -1409
rect 1556 -1410 1557 -1409
rect 1605 -1410 1606 -1409
rect 1661 -1410 1662 -1409
rect 1738 -1410 1739 -1409
rect 1794 -1410 1795 -1409
rect 1857 -1410 1858 -1409
rect 51 -1412 52 -1411
rect 1899 -1412 1900 -1411
rect 51 -1414 52 -1413
rect 100 -1414 101 -1413
rect 107 -1414 108 -1413
rect 233 -1414 234 -1413
rect 450 -1414 451 -1413
rect 632 -1414 633 -1413
rect 814 -1414 815 -1413
rect 968 -1414 969 -1413
rect 975 -1414 976 -1413
rect 1307 -1414 1308 -1413
rect 1335 -1414 1336 -1413
rect 1906 -1414 1907 -1413
rect 58 -1416 59 -1415
rect 499 -1416 500 -1415
rect 548 -1416 549 -1415
rect 681 -1416 682 -1415
rect 814 -1416 815 -1415
rect 828 -1416 829 -1415
rect 849 -1416 850 -1415
rect 940 -1416 941 -1415
rect 947 -1416 948 -1415
rect 1360 -1416 1361 -1415
rect 1437 -1416 1438 -1415
rect 1591 -1416 1592 -1415
rect 1801 -1416 1802 -1415
rect 1906 -1416 1907 -1415
rect 58 -1418 59 -1417
rect 247 -1418 248 -1417
rect 408 -1418 409 -1417
rect 548 -1418 549 -1417
rect 562 -1418 563 -1417
rect 709 -1418 710 -1417
rect 744 -1418 745 -1417
rect 828 -1418 829 -1417
rect 905 -1418 906 -1417
rect 912 -1418 913 -1417
rect 922 -1418 923 -1417
rect 1941 -1418 1942 -1417
rect 65 -1420 66 -1419
rect 72 -1420 73 -1419
rect 79 -1420 80 -1419
rect 261 -1420 262 -1419
rect 408 -1420 409 -1419
rect 506 -1420 507 -1419
rect 562 -1420 563 -1419
rect 709 -1420 710 -1419
rect 744 -1420 745 -1419
rect 835 -1420 836 -1419
rect 842 -1420 843 -1419
rect 905 -1420 906 -1419
rect 926 -1420 927 -1419
rect 933 -1420 934 -1419
rect 961 -1420 962 -1419
rect 1178 -1420 1179 -1419
rect 1185 -1420 1186 -1419
rect 1262 -1420 1263 -1419
rect 1283 -1420 1284 -1419
rect 1836 -1420 1837 -1419
rect 1850 -1420 1851 -1419
rect 1857 -1420 1858 -1419
rect 79 -1422 80 -1421
rect 835 -1422 836 -1421
rect 884 -1422 885 -1421
rect 933 -1422 934 -1421
rect 985 -1422 986 -1421
rect 1409 -1422 1410 -1421
rect 1521 -1422 1522 -1421
rect 1556 -1422 1557 -1421
rect 1577 -1422 1578 -1421
rect 1654 -1422 1655 -1421
rect 1703 -1422 1704 -1421
rect 1801 -1422 1802 -1421
rect 82 -1424 83 -1423
rect 1136 -1424 1137 -1423
rect 1164 -1424 1165 -1423
rect 1241 -1424 1242 -1423
rect 1283 -1424 1284 -1423
rect 1325 -1424 1326 -1423
rect 1346 -1424 1347 -1423
rect 1360 -1424 1361 -1423
rect 1374 -1424 1375 -1423
rect 1409 -1424 1410 -1423
rect 1507 -1424 1508 -1423
rect 1521 -1424 1522 -1423
rect 1535 -1424 1536 -1423
rect 1661 -1424 1662 -1423
rect 1703 -1424 1704 -1423
rect 1773 -1424 1774 -1423
rect 86 -1426 87 -1425
rect 184 -1426 185 -1425
rect 194 -1426 195 -1425
rect 695 -1426 696 -1425
rect 751 -1426 752 -1425
rect 842 -1426 843 -1425
rect 982 -1426 983 -1425
rect 1136 -1426 1137 -1425
rect 1150 -1426 1151 -1425
rect 1164 -1426 1165 -1425
rect 1171 -1426 1172 -1425
rect 1451 -1426 1452 -1425
rect 1479 -1426 1480 -1425
rect 1507 -1426 1508 -1425
rect 1549 -1426 1550 -1425
rect 1850 -1426 1851 -1425
rect 93 -1428 94 -1427
rect 100 -1428 101 -1427
rect 114 -1428 115 -1427
rect 432 -1428 433 -1427
rect 450 -1428 451 -1427
rect 579 -1428 580 -1427
rect 583 -1428 584 -1427
rect 695 -1428 696 -1427
rect 786 -1428 787 -1427
rect 849 -1428 850 -1427
rect 982 -1428 983 -1427
rect 1640 -1428 1641 -1427
rect 1717 -1428 1718 -1427
rect 1773 -1428 1774 -1427
rect 93 -1430 94 -1429
rect 149 -1430 150 -1429
rect 198 -1430 199 -1429
rect 243 -1430 244 -1429
rect 247 -1430 248 -1429
rect 950 -1430 951 -1429
rect 996 -1430 997 -1429
rect 1381 -1430 1382 -1429
rect 1388 -1430 1389 -1429
rect 1451 -1430 1452 -1429
rect 1549 -1430 1550 -1429
rect 1626 -1430 1627 -1429
rect 1640 -1430 1641 -1429
rect 1997 -1430 1998 -1429
rect 114 -1432 115 -1431
rect 436 -1432 437 -1431
rect 492 -1432 493 -1431
rect 667 -1432 668 -1431
rect 807 -1432 808 -1431
rect 1171 -1432 1172 -1431
rect 1178 -1432 1179 -1431
rect 1395 -1432 1396 -1431
rect 1759 -1432 1760 -1431
rect 1836 -1432 1837 -1431
rect 121 -1434 122 -1433
rect 131 -1434 132 -1433
rect 145 -1434 146 -1433
rect 1913 -1434 1914 -1433
rect 145 -1436 146 -1435
rect 1206 -1436 1207 -1435
rect 1248 -1436 1249 -1435
rect 1325 -1436 1326 -1435
rect 1346 -1436 1347 -1435
rect 1472 -1436 1473 -1435
rect 1752 -1436 1753 -1435
rect 1759 -1436 1760 -1435
rect 149 -1438 150 -1437
rect 1108 -1438 1109 -1437
rect 1111 -1438 1112 -1437
rect 1612 -1438 1613 -1437
rect 198 -1440 199 -1439
rect 282 -1440 283 -1439
rect 310 -1440 311 -1439
rect 786 -1440 787 -1439
rect 793 -1440 794 -1439
rect 807 -1440 808 -1439
rect 929 -1440 930 -1439
rect 1472 -1440 1473 -1439
rect 1493 -1440 1494 -1439
rect 1752 -1440 1753 -1439
rect 37 -1442 38 -1441
rect 282 -1442 283 -1441
rect 303 -1442 304 -1441
rect 310 -1442 311 -1441
rect 373 -1442 374 -1441
rect 436 -1442 437 -1441
rect 506 -1442 507 -1441
rect 513 -1442 514 -1441
rect 569 -1442 570 -1441
rect 943 -1442 944 -1441
rect 954 -1442 955 -1441
rect 996 -1442 997 -1441
rect 1003 -1442 1004 -1441
rect 1045 -1442 1046 -1441
rect 1066 -1442 1067 -1441
rect 1710 -1442 1711 -1441
rect 37 -1444 38 -1443
rect 75 -1444 76 -1443
rect 86 -1444 87 -1443
rect 954 -1444 955 -1443
rect 1006 -1444 1007 -1443
rect 1199 -1444 1200 -1443
rect 1248 -1444 1249 -1443
rect 1290 -1444 1291 -1443
rect 1367 -1444 1368 -1443
rect 1395 -1444 1396 -1443
rect 1493 -1444 1494 -1443
rect 1570 -1444 1571 -1443
rect 1633 -1444 1634 -1443
rect 1710 -1444 1711 -1443
rect 1986 -1444 1987 -1443
rect 1990 -1444 1991 -1443
rect 110 -1446 111 -1445
rect 303 -1446 304 -1445
rect 338 -1446 339 -1445
rect 373 -1446 374 -1445
rect 387 -1446 388 -1445
rect 1206 -1446 1207 -1445
rect 1255 -1446 1256 -1445
rect 1388 -1446 1389 -1445
rect 1528 -1446 1529 -1445
rect 1570 -1446 1571 -1445
rect 128 -1448 129 -1447
rect 1633 -1448 1634 -1447
rect 128 -1450 129 -1449
rect 135 -1450 136 -1449
rect 205 -1450 206 -1449
rect 226 -1450 227 -1449
rect 233 -1450 234 -1449
rect 1304 -1450 1305 -1449
rect 1367 -1450 1368 -1449
rect 1423 -1450 1424 -1449
rect 1486 -1450 1487 -1449
rect 1528 -1450 1529 -1449
rect 1563 -1450 1564 -1449
rect 1612 -1450 1613 -1449
rect 135 -1452 136 -1451
rect 177 -1452 178 -1451
rect 226 -1452 227 -1451
rect 331 -1452 332 -1451
rect 338 -1452 339 -1451
rect 520 -1452 521 -1451
rect 555 -1452 556 -1451
rect 569 -1452 570 -1451
rect 576 -1452 577 -1451
rect 859 -1452 860 -1451
rect 1010 -1452 1011 -1451
rect 1717 -1452 1718 -1451
rect 296 -1454 297 -1453
rect 331 -1454 332 -1453
rect 387 -1454 388 -1453
rect 394 -1454 395 -1453
rect 422 -1454 423 -1453
rect 583 -1454 584 -1453
rect 590 -1454 591 -1453
rect 646 -1454 647 -1453
rect 663 -1454 664 -1453
rect 1437 -1454 1438 -1453
rect 163 -1456 164 -1455
rect 394 -1456 395 -1455
rect 415 -1456 416 -1455
rect 422 -1456 423 -1455
rect 513 -1456 514 -1455
rect 611 -1456 612 -1455
rect 618 -1456 619 -1455
rect 628 -1456 629 -1455
rect 793 -1456 794 -1455
rect 800 -1456 801 -1455
rect 898 -1456 899 -1455
rect 1010 -1456 1011 -1455
rect 1024 -1456 1025 -1455
rect 1885 -1456 1886 -1455
rect 163 -1458 164 -1457
rect 254 -1458 255 -1457
rect 415 -1458 416 -1457
rect 457 -1458 458 -1457
rect 478 -1458 479 -1457
rect 800 -1458 801 -1457
rect 821 -1458 822 -1457
rect 898 -1458 899 -1457
rect 1031 -1458 1032 -1457
rect 1626 -1458 1627 -1457
rect 212 -1460 213 -1459
rect 457 -1460 458 -1459
rect 520 -1460 521 -1459
rect 688 -1460 689 -1459
rect 702 -1460 703 -1459
rect 821 -1460 822 -1459
rect 989 -1460 990 -1459
rect 1031 -1460 1032 -1459
rect 1034 -1460 1035 -1459
rect 1654 -1460 1655 -1459
rect 177 -1462 178 -1461
rect 212 -1462 213 -1461
rect 219 -1462 220 -1461
rect 296 -1462 297 -1461
rect 443 -1462 444 -1461
rect 478 -1462 479 -1461
rect 534 -1462 535 -1461
rect 702 -1462 703 -1461
rect 751 -1462 752 -1461
rect 1024 -1462 1025 -1461
rect 1087 -1462 1088 -1461
rect 1535 -1462 1536 -1461
rect 191 -1464 192 -1463
rect 534 -1464 535 -1463
rect 555 -1464 556 -1463
rect 2007 -1464 2008 -1463
rect 191 -1466 192 -1465
rect 772 -1466 773 -1465
rect 989 -1466 990 -1465
rect 1017 -1466 1018 -1465
rect 1087 -1466 1088 -1465
rect 1094 -1466 1095 -1465
rect 1108 -1466 1109 -1465
rect 1479 -1466 1480 -1465
rect 219 -1468 220 -1467
rect 289 -1468 290 -1467
rect 359 -1468 360 -1467
rect 443 -1468 444 -1467
rect 576 -1468 577 -1467
rect 779 -1468 780 -1467
rect 863 -1468 864 -1467
rect 1017 -1468 1018 -1467
rect 1080 -1468 1081 -1467
rect 1094 -1468 1095 -1467
rect 1111 -1468 1112 -1467
rect 1290 -1468 1291 -1467
rect 1304 -1468 1305 -1467
rect 1829 -1468 1830 -1467
rect 254 -1470 255 -1469
rect 268 -1470 269 -1469
rect 275 -1470 276 -1469
rect 289 -1470 290 -1469
rect 324 -1470 325 -1469
rect 359 -1470 360 -1469
rect 590 -1470 591 -1469
rect 856 -1470 857 -1469
rect 1080 -1470 1081 -1469
rect 1265 -1470 1266 -1469
rect 1286 -1470 1287 -1469
rect 1339 -1470 1340 -1469
rect 1402 -1470 1403 -1469
rect 1423 -1470 1424 -1469
rect 1731 -1470 1732 -1469
rect 1829 -1470 1830 -1469
rect 240 -1472 241 -1471
rect 268 -1472 269 -1471
rect 275 -1472 276 -1471
rect 352 -1472 353 -1471
rect 597 -1472 598 -1471
rect 656 -1472 657 -1471
rect 670 -1472 671 -1471
rect 1402 -1472 1403 -1471
rect 1724 -1472 1725 -1471
rect 1731 -1472 1732 -1471
rect 324 -1474 325 -1473
rect 401 -1474 402 -1473
rect 464 -1474 465 -1473
rect 597 -1474 598 -1473
rect 604 -1474 605 -1473
rect 884 -1474 885 -1473
rect 1115 -1474 1116 -1473
rect 1262 -1474 1263 -1473
rect 1339 -1474 1340 -1473
rect 1458 -1474 1459 -1473
rect 1696 -1474 1697 -1473
rect 1724 -1474 1725 -1473
rect 352 -1476 353 -1475
rect 639 -1476 640 -1475
rect 653 -1476 654 -1475
rect 863 -1476 864 -1475
rect 1118 -1476 1119 -1475
rect 1745 -1476 1746 -1475
rect 401 -1478 402 -1477
rect 502 -1478 503 -1477
rect 541 -1478 542 -1477
rect 639 -1478 640 -1477
rect 653 -1478 654 -1477
rect 1132 -1478 1133 -1477
rect 1143 -1478 1144 -1477
rect 1150 -1478 1151 -1477
rect 1160 -1478 1161 -1477
rect 1486 -1478 1487 -1477
rect 1675 -1478 1676 -1477
rect 1745 -1478 1746 -1477
rect 44 -1480 45 -1479
rect 541 -1480 542 -1479
rect 604 -1480 605 -1479
rect 712 -1480 713 -1479
rect 758 -1480 759 -1479
rect 772 -1480 773 -1479
rect 779 -1480 780 -1479
rect 891 -1480 892 -1479
rect 1059 -1480 1060 -1479
rect 1143 -1480 1144 -1479
rect 1199 -1480 1200 -1479
rect 1213 -1480 1214 -1479
rect 1220 -1480 1221 -1479
rect 1255 -1480 1256 -1479
rect 1416 -1480 1417 -1479
rect 1458 -1480 1459 -1479
rect 1584 -1480 1585 -1479
rect 1675 -1480 1676 -1479
rect 44 -1482 45 -1481
rect 1920 -1482 1921 -1481
rect 170 -1484 171 -1483
rect 758 -1484 759 -1483
rect 856 -1484 857 -1483
rect 1115 -1484 1116 -1483
rect 1122 -1484 1123 -1483
rect 1563 -1484 1564 -1483
rect 61 -1486 62 -1485
rect 170 -1486 171 -1485
rect 464 -1486 465 -1485
rect 530 -1486 531 -1485
rect 611 -1486 612 -1485
rect 1076 -1486 1077 -1485
rect 1101 -1486 1102 -1485
rect 1122 -1486 1123 -1485
rect 1157 -1486 1158 -1485
rect 1213 -1486 1214 -1485
rect 1244 -1486 1245 -1485
rect 1696 -1486 1697 -1485
rect 61 -1488 62 -1487
rect 65 -1488 66 -1487
rect 628 -1488 629 -1487
rect 716 -1488 717 -1487
rect 870 -1488 871 -1487
rect 891 -1488 892 -1487
rect 1059 -1488 1060 -1487
rect 1129 -1488 1130 -1487
rect 1157 -1488 1158 -1487
rect 1871 -1488 1872 -1487
rect 471 -1490 472 -1489
rect 870 -1490 871 -1489
rect 1101 -1490 1102 -1489
rect 1311 -1490 1312 -1489
rect 1318 -1490 1319 -1489
rect 1416 -1490 1417 -1489
rect 1815 -1490 1816 -1489
rect 1871 -1490 1872 -1489
rect 366 -1492 367 -1491
rect 471 -1492 472 -1491
rect 688 -1492 689 -1491
rect 730 -1492 731 -1491
rect 1129 -1492 1130 -1491
rect 1374 -1492 1375 -1491
rect 1668 -1492 1669 -1491
rect 1815 -1492 1816 -1491
rect 366 -1494 367 -1493
rect 380 -1494 381 -1493
rect 716 -1494 717 -1493
rect 737 -1494 738 -1493
rect 1192 -1494 1193 -1493
rect 1220 -1494 1221 -1493
rect 1297 -1494 1298 -1493
rect 1318 -1494 1319 -1493
rect 1598 -1494 1599 -1493
rect 1668 -1494 1669 -1493
rect 380 -1496 381 -1495
rect 765 -1496 766 -1495
rect 1192 -1496 1193 -1495
rect 1787 -1496 1788 -1495
rect 660 -1498 661 -1497
rect 765 -1498 766 -1497
rect 1269 -1498 1270 -1497
rect 1297 -1498 1298 -1497
rect 1311 -1498 1312 -1497
rect 1514 -1498 1515 -1497
rect 1598 -1498 1599 -1497
rect 1689 -1498 1690 -1497
rect 156 -1500 157 -1499
rect 660 -1500 661 -1499
rect 723 -1500 724 -1499
rect 737 -1500 738 -1499
rect 1269 -1500 1270 -1499
rect 1276 -1500 1277 -1499
rect 1619 -1500 1620 -1499
rect 1689 -1500 1690 -1499
rect 156 -1502 157 -1501
rect 429 -1502 430 -1501
rect 730 -1502 731 -1501
rect 754 -1502 755 -1501
rect 1069 -1502 1070 -1501
rect 1619 -1502 1620 -1501
rect 240 -1504 241 -1503
rect 723 -1504 724 -1503
rect 1069 -1504 1070 -1503
rect 1500 -1504 1501 -1503
rect 317 -1506 318 -1505
rect 429 -1506 430 -1505
rect 1234 -1506 1235 -1505
rect 1276 -1506 1277 -1505
rect 1465 -1506 1466 -1505
rect 1500 -1506 1501 -1505
rect 317 -1508 318 -1507
rect 345 -1508 346 -1507
rect 1227 -1508 1228 -1507
rect 1234 -1508 1235 -1507
rect 1430 -1508 1431 -1507
rect 1465 -1508 1466 -1507
rect 166 -1510 167 -1509
rect 345 -1510 346 -1509
rect 625 -1510 626 -1509
rect 1227 -1510 1228 -1509
rect 1353 -1510 1354 -1509
rect 1430 -1510 1431 -1509
rect 625 -1512 626 -1511
rect 1584 -1512 1585 -1511
rect 1332 -1514 1333 -1513
rect 1353 -1514 1354 -1513
rect 1332 -1516 1333 -1515
rect 1514 -1516 1515 -1515
rect 2 -1527 3 -1526
rect 47 -1527 48 -1526
rect 58 -1527 59 -1526
rect 1724 -1527 1725 -1526
rect 1808 -1527 1809 -1526
rect 1811 -1527 1812 -1526
rect 1948 -1527 1949 -1526
rect 1969 -1527 1970 -1526
rect 1979 -1527 1980 -1526
rect 1990 -1527 1991 -1526
rect 2 -1529 3 -1528
rect 177 -1529 178 -1528
rect 180 -1529 181 -1528
rect 254 -1529 255 -1528
rect 338 -1529 339 -1528
rect 751 -1529 752 -1528
rect 754 -1529 755 -1528
rect 1661 -1529 1662 -1528
rect 1689 -1529 1690 -1528
rect 1724 -1529 1725 -1528
rect 1766 -1529 1767 -1528
rect 1948 -1529 1949 -1528
rect 1955 -1529 1956 -1528
rect 1972 -1529 1973 -1528
rect 1983 -1529 1984 -1528
rect 2000 -1529 2001 -1528
rect 23 -1531 24 -1530
rect 68 -1531 69 -1530
rect 82 -1531 83 -1530
rect 1104 -1531 1105 -1530
rect 1108 -1531 1109 -1530
rect 1829 -1531 1830 -1530
rect 23 -1533 24 -1532
rect 198 -1533 199 -1532
rect 233 -1533 234 -1532
rect 324 -1533 325 -1532
rect 338 -1533 339 -1532
rect 359 -1533 360 -1532
rect 485 -1533 486 -1532
rect 660 -1533 661 -1532
rect 663 -1533 664 -1532
rect 751 -1533 752 -1532
rect 768 -1533 769 -1532
rect 814 -1533 815 -1532
rect 884 -1533 885 -1532
rect 1160 -1533 1161 -1532
rect 1192 -1533 1193 -1532
rect 1234 -1533 1235 -1532
rect 1262 -1533 1263 -1532
rect 1346 -1533 1347 -1532
rect 1356 -1533 1357 -1532
rect 1731 -1533 1732 -1532
rect 1808 -1533 1809 -1532
rect 1878 -1533 1879 -1532
rect 30 -1535 31 -1534
rect 919 -1535 920 -1534
rect 954 -1535 955 -1534
rect 1850 -1535 1851 -1534
rect 30 -1537 31 -1536
rect 247 -1537 248 -1536
rect 254 -1537 255 -1536
rect 1055 -1537 1056 -1536
rect 1101 -1537 1102 -1536
rect 1339 -1537 1340 -1536
rect 1346 -1537 1347 -1536
rect 1360 -1537 1361 -1536
rect 1503 -1537 1504 -1536
rect 1836 -1537 1837 -1536
rect 37 -1539 38 -1538
rect 499 -1539 500 -1538
rect 502 -1539 503 -1538
rect 1038 -1539 1039 -1538
rect 1108 -1539 1109 -1538
rect 1335 -1539 1336 -1538
rect 1339 -1539 1340 -1538
rect 1353 -1539 1354 -1538
rect 1360 -1539 1361 -1538
rect 1381 -1539 1382 -1538
rect 1591 -1539 1592 -1538
rect 2004 -1539 2005 -1538
rect 37 -1541 38 -1540
rect 51 -1541 52 -1540
rect 58 -1541 59 -1540
rect 107 -1541 108 -1540
rect 117 -1541 118 -1540
rect 121 -1541 122 -1540
rect 142 -1541 143 -1540
rect 303 -1541 304 -1540
rect 324 -1541 325 -1540
rect 443 -1541 444 -1540
rect 499 -1541 500 -1540
rect 555 -1541 556 -1540
rect 593 -1541 594 -1540
rect 688 -1541 689 -1540
rect 709 -1541 710 -1540
rect 877 -1541 878 -1540
rect 905 -1541 906 -1540
rect 947 -1541 948 -1540
rect 957 -1541 958 -1540
rect 1689 -1541 1690 -1540
rect 1703 -1541 1704 -1540
rect 1766 -1541 1767 -1540
rect 1811 -1541 1812 -1540
rect 1878 -1541 1879 -1540
rect 9 -1543 10 -1542
rect 51 -1543 52 -1542
rect 86 -1543 87 -1542
rect 107 -1543 108 -1542
rect 121 -1543 122 -1542
rect 184 -1543 185 -1542
rect 194 -1543 195 -1542
rect 1206 -1543 1207 -1542
rect 1234 -1543 1235 -1542
rect 1255 -1543 1256 -1542
rect 1262 -1543 1263 -1542
rect 1286 -1543 1287 -1542
rect 1353 -1543 1354 -1542
rect 1528 -1543 1529 -1542
rect 1577 -1543 1578 -1542
rect 1703 -1543 1704 -1542
rect 1717 -1543 1718 -1542
rect 1850 -1543 1851 -1542
rect 9 -1545 10 -1544
rect 156 -1545 157 -1544
rect 184 -1545 185 -1544
rect 544 -1545 545 -1544
rect 555 -1545 556 -1544
rect 702 -1545 703 -1544
rect 712 -1545 713 -1544
rect 1542 -1545 1543 -1544
rect 1577 -1545 1578 -1544
rect 1612 -1545 1613 -1544
rect 1661 -1545 1662 -1544
rect 1976 -1545 1977 -1544
rect 44 -1547 45 -1546
rect 100 -1547 101 -1546
rect 142 -1547 143 -1546
rect 628 -1547 629 -1546
rect 667 -1547 668 -1546
rect 1171 -1547 1172 -1546
rect 1199 -1547 1200 -1546
rect 1255 -1547 1256 -1546
rect 1265 -1547 1266 -1546
rect 1962 -1547 1963 -1546
rect 1976 -1547 1977 -1546
rect 2025 -1547 2026 -1546
rect 16 -1549 17 -1548
rect 44 -1549 45 -1548
rect 79 -1549 80 -1548
rect 100 -1549 101 -1548
rect 114 -1549 115 -1548
rect 667 -1549 668 -1548
rect 674 -1549 675 -1548
rect 1038 -1549 1039 -1548
rect 1111 -1549 1112 -1548
rect 1822 -1549 1823 -1548
rect 1829 -1549 1830 -1548
rect 1885 -1549 1886 -1548
rect 16 -1551 17 -1550
rect 89 -1551 90 -1550
rect 145 -1551 146 -1550
rect 198 -1551 199 -1550
rect 226 -1551 227 -1550
rect 247 -1551 248 -1550
rect 289 -1551 290 -1550
rect 485 -1551 486 -1550
rect 618 -1551 619 -1550
rect 1101 -1551 1102 -1550
rect 1118 -1551 1119 -1550
rect 1185 -1551 1186 -1550
rect 1199 -1551 1200 -1550
rect 1213 -1551 1214 -1550
rect 1374 -1551 1375 -1550
rect 1381 -1551 1382 -1550
rect 1493 -1551 1494 -1550
rect 1591 -1551 1592 -1550
rect 1612 -1551 1613 -1550
rect 1619 -1551 1620 -1550
rect 1731 -1551 1732 -1550
rect 1752 -1551 1753 -1550
rect 1794 -1551 1795 -1550
rect 1885 -1551 1886 -1550
rect 86 -1553 87 -1552
rect 698 -1553 699 -1552
rect 702 -1553 703 -1552
rect 821 -1553 822 -1552
rect 835 -1553 836 -1552
rect 877 -1553 878 -1552
rect 961 -1553 962 -1552
rect 1332 -1553 1333 -1552
rect 1374 -1553 1375 -1552
rect 1395 -1553 1396 -1552
rect 1493 -1553 1494 -1552
rect 1668 -1553 1669 -1552
rect 1822 -1553 1823 -1552
rect 1906 -1553 1907 -1552
rect 128 -1555 129 -1554
rect 145 -1555 146 -1554
rect 156 -1555 157 -1554
rect 219 -1555 220 -1554
rect 226 -1555 227 -1554
rect 1115 -1555 1116 -1554
rect 1129 -1555 1130 -1554
rect 1881 -1555 1882 -1554
rect 1906 -1555 1907 -1554
rect 1934 -1555 1935 -1554
rect 93 -1557 94 -1556
rect 128 -1557 129 -1556
rect 191 -1557 192 -1556
rect 219 -1557 220 -1556
rect 233 -1557 234 -1556
rect 310 -1557 311 -1556
rect 345 -1557 346 -1556
rect 670 -1557 671 -1556
rect 681 -1557 682 -1556
rect 1304 -1557 1305 -1556
rect 1307 -1557 1308 -1556
rect 1752 -1557 1753 -1556
rect 1871 -1557 1872 -1556
rect 1934 -1557 1935 -1556
rect 65 -1559 66 -1558
rect 93 -1559 94 -1558
rect 163 -1559 164 -1558
rect 191 -1559 192 -1558
rect 205 -1559 206 -1558
rect 345 -1559 346 -1558
rect 415 -1559 416 -1558
rect 821 -1559 822 -1558
rect 849 -1559 850 -1558
rect 905 -1559 906 -1558
rect 971 -1559 972 -1558
rect 1283 -1559 1284 -1558
rect 1307 -1559 1308 -1558
rect 1857 -1559 1858 -1558
rect 1871 -1559 1872 -1558
rect 1920 -1559 1921 -1558
rect 163 -1561 164 -1560
rect 660 -1561 661 -1560
rect 663 -1561 664 -1560
rect 1794 -1561 1795 -1560
rect 205 -1563 206 -1562
rect 520 -1563 521 -1562
rect 646 -1563 647 -1562
rect 674 -1563 675 -1562
rect 681 -1563 682 -1562
rect 828 -1563 829 -1562
rect 863 -1563 864 -1562
rect 1717 -1563 1718 -1562
rect 268 -1565 269 -1564
rect 310 -1565 311 -1564
rect 397 -1565 398 -1564
rect 646 -1565 647 -1564
rect 670 -1565 671 -1564
rect 842 -1565 843 -1564
rect 1003 -1565 1004 -1564
rect 1801 -1565 1802 -1564
rect 268 -1567 269 -1566
rect 569 -1567 570 -1566
rect 583 -1567 584 -1566
rect 842 -1567 843 -1566
rect 968 -1567 969 -1566
rect 1003 -1567 1004 -1566
rect 1073 -1567 1074 -1566
rect 1115 -1567 1116 -1566
rect 1132 -1567 1133 -1566
rect 1311 -1567 1312 -1566
rect 1332 -1567 1333 -1566
rect 1864 -1567 1865 -1566
rect 282 -1569 283 -1568
rect 520 -1569 521 -1568
rect 569 -1569 570 -1568
rect 576 -1569 577 -1568
rect 583 -1569 584 -1568
rect 730 -1569 731 -1568
rect 800 -1569 801 -1568
rect 1129 -1569 1130 -1568
rect 1132 -1569 1133 -1568
rect 1549 -1569 1550 -1568
rect 1619 -1569 1620 -1568
rect 1633 -1569 1634 -1568
rect 1647 -1569 1648 -1568
rect 1857 -1569 1858 -1568
rect 1864 -1569 1865 -1568
rect 1913 -1569 1914 -1568
rect 282 -1571 283 -1570
rect 450 -1571 451 -1570
rect 457 -1571 458 -1570
rect 712 -1571 713 -1570
rect 723 -1571 724 -1570
rect 1209 -1571 1210 -1570
rect 1213 -1571 1214 -1570
rect 1444 -1571 1445 -1570
rect 1507 -1571 1508 -1570
rect 1633 -1571 1634 -1570
rect 1647 -1571 1648 -1570
rect 1654 -1571 1655 -1570
rect 1668 -1571 1669 -1570
rect 1696 -1571 1697 -1570
rect 1787 -1571 1788 -1570
rect 1801 -1571 1802 -1570
rect 1913 -1571 1914 -1570
rect 1941 -1571 1942 -1570
rect 261 -1573 262 -1572
rect 450 -1573 451 -1572
rect 464 -1573 465 -1572
rect 688 -1573 689 -1572
rect 723 -1573 724 -1572
rect 982 -1573 983 -1572
rect 1024 -1573 1025 -1572
rect 1073 -1573 1074 -1572
rect 1150 -1573 1151 -1572
rect 1192 -1573 1193 -1572
rect 1283 -1573 1284 -1572
rect 1626 -1573 1627 -1572
rect 1654 -1573 1655 -1572
rect 1682 -1573 1683 -1572
rect 1696 -1573 1697 -1572
rect 1843 -1573 1844 -1572
rect 1941 -1573 1942 -1572
rect 2011 -1573 2012 -1572
rect 261 -1575 262 -1574
rect 1069 -1575 1070 -1574
rect 1171 -1575 1172 -1574
rect 1241 -1575 1242 -1574
rect 1311 -1575 1312 -1574
rect 1318 -1575 1319 -1574
rect 1395 -1575 1396 -1574
rect 1402 -1575 1403 -1574
rect 1444 -1575 1445 -1574
rect 1465 -1575 1466 -1574
rect 1521 -1575 1522 -1574
rect 1528 -1575 1529 -1574
rect 1542 -1575 1543 -1574
rect 1563 -1575 1564 -1574
rect 1626 -1575 1627 -1574
rect 1710 -1575 1711 -1574
rect 1787 -1575 1788 -1574
rect 1927 -1575 1928 -1574
rect 65 -1577 66 -1576
rect 1710 -1577 1711 -1576
rect 1843 -1577 1844 -1576
rect 1920 -1577 1921 -1576
rect 289 -1579 290 -1578
rect 366 -1579 367 -1578
rect 418 -1579 419 -1578
rect 849 -1579 850 -1578
rect 919 -1579 920 -1578
rect 1507 -1579 1508 -1578
rect 1521 -1579 1522 -1578
rect 1605 -1579 1606 -1578
rect 296 -1581 297 -1580
rect 359 -1581 360 -1580
rect 366 -1581 367 -1580
rect 429 -1581 430 -1580
rect 443 -1581 444 -1580
rect 653 -1581 654 -1580
rect 730 -1581 731 -1580
rect 975 -1581 976 -1580
rect 1006 -1581 1007 -1580
rect 1682 -1581 1683 -1580
rect 114 -1583 115 -1582
rect 653 -1583 654 -1582
rect 772 -1583 773 -1582
rect 800 -1583 801 -1582
rect 807 -1583 808 -1582
rect 954 -1583 955 -1582
rect 968 -1583 969 -1582
rect 989 -1583 990 -1582
rect 1024 -1583 1025 -1582
rect 1136 -1583 1137 -1582
rect 1185 -1583 1186 -1582
rect 1248 -1583 1249 -1582
rect 1290 -1583 1291 -1582
rect 1465 -1583 1466 -1582
rect 1549 -1583 1550 -1582
rect 1556 -1583 1557 -1582
rect 1563 -1583 1564 -1582
rect 1584 -1583 1585 -1582
rect 1598 -1583 1599 -1582
rect 1927 -1583 1928 -1582
rect 296 -1585 297 -1584
rect 985 -1585 986 -1584
rect 989 -1585 990 -1584
rect 1090 -1585 1091 -1584
rect 1220 -1585 1221 -1584
rect 1248 -1585 1249 -1584
rect 1290 -1585 1291 -1584
rect 1297 -1585 1298 -1584
rect 1402 -1585 1403 -1584
rect 1416 -1585 1417 -1584
rect 1535 -1585 1536 -1584
rect 1584 -1585 1585 -1584
rect 1598 -1585 1599 -1584
rect 1640 -1585 1641 -1584
rect 303 -1587 304 -1586
rect 331 -1587 332 -1586
rect 422 -1587 423 -1586
rect 457 -1587 458 -1586
rect 478 -1587 479 -1586
rect 618 -1587 619 -1586
rect 765 -1587 766 -1586
rect 772 -1587 773 -1586
rect 793 -1587 794 -1586
rect 807 -1587 808 -1586
rect 817 -1587 818 -1586
rect 1836 -1587 1837 -1586
rect 212 -1589 213 -1588
rect 422 -1589 423 -1588
rect 429 -1589 430 -1588
rect 950 -1589 951 -1588
rect 1031 -1589 1032 -1588
rect 1150 -1589 1151 -1588
rect 1164 -1589 1165 -1588
rect 1297 -1589 1298 -1588
rect 1367 -1589 1368 -1588
rect 1535 -1589 1536 -1588
rect 1570 -1589 1571 -1588
rect 1605 -1589 1606 -1588
rect 170 -1591 171 -1590
rect 212 -1591 213 -1590
rect 317 -1591 318 -1590
rect 464 -1591 465 -1590
rect 478 -1591 479 -1590
rect 513 -1591 514 -1590
rect 597 -1591 598 -1590
rect 863 -1591 864 -1590
rect 922 -1591 923 -1590
rect 1640 -1591 1641 -1590
rect 317 -1593 318 -1592
rect 611 -1593 612 -1592
rect 793 -1593 794 -1592
rect 856 -1593 857 -1592
rect 884 -1593 885 -1592
rect 922 -1593 923 -1592
rect 926 -1593 927 -1592
rect 982 -1593 983 -1592
rect 1010 -1593 1011 -1592
rect 1031 -1593 1032 -1592
rect 1059 -1593 1060 -1592
rect 1318 -1593 1319 -1592
rect 1367 -1593 1368 -1592
rect 1388 -1593 1389 -1592
rect 1416 -1593 1417 -1592
rect 1423 -1593 1424 -1592
rect 79 -1595 80 -1594
rect 1010 -1595 1011 -1594
rect 1080 -1595 1081 -1594
rect 1164 -1595 1165 -1594
rect 1195 -1595 1196 -1594
rect 1570 -1595 1571 -1594
rect 331 -1597 332 -1596
rect 387 -1597 388 -1596
rect 513 -1597 514 -1596
rect 541 -1597 542 -1596
rect 611 -1597 612 -1596
rect 740 -1597 741 -1596
rect 828 -1597 829 -1596
rect 1136 -1597 1137 -1596
rect 1220 -1597 1221 -1596
rect 1276 -1597 1277 -1596
rect 1388 -1597 1389 -1596
rect 1451 -1597 1452 -1596
rect 387 -1599 388 -1598
rect 814 -1599 815 -1598
rect 856 -1599 857 -1598
rect 891 -1599 892 -1598
rect 912 -1599 913 -1598
rect 926 -1599 927 -1598
rect 933 -1599 934 -1598
rect 975 -1599 976 -1598
rect 1080 -1599 1081 -1598
rect 1227 -1599 1228 -1598
rect 1241 -1599 1242 -1598
rect 1815 -1599 1816 -1598
rect 177 -1601 178 -1600
rect 933 -1601 934 -1600
rect 940 -1601 941 -1600
rect 1059 -1601 1060 -1600
rect 1227 -1601 1228 -1600
rect 1409 -1601 1410 -1600
rect 1423 -1601 1424 -1600
rect 1430 -1601 1431 -1600
rect 1451 -1601 1452 -1600
rect 1472 -1601 1473 -1600
rect 1815 -1601 1816 -1600
rect 1899 -1601 1900 -1600
rect 352 -1603 353 -1602
rect 1430 -1603 1431 -1602
rect 1458 -1603 1459 -1602
rect 1472 -1603 1473 -1602
rect 352 -1605 353 -1604
rect 562 -1605 563 -1604
rect 870 -1605 871 -1604
rect 1276 -1605 1277 -1604
rect 1458 -1605 1459 -1604
rect 1479 -1605 1480 -1604
rect 380 -1607 381 -1606
rect 940 -1607 941 -1606
rect 1094 -1607 1095 -1606
rect 1409 -1607 1410 -1606
rect 1479 -1607 1480 -1606
rect 1486 -1607 1487 -1606
rect 380 -1609 381 -1608
rect 492 -1609 493 -1608
rect 534 -1609 535 -1608
rect 597 -1609 598 -1608
rect 786 -1609 787 -1608
rect 870 -1609 871 -1608
rect 891 -1609 892 -1608
rect 1178 -1609 1179 -1608
rect 1206 -1609 1207 -1608
rect 1899 -1609 1900 -1608
rect 394 -1611 395 -1610
rect 492 -1611 493 -1610
rect 541 -1611 542 -1610
rect 576 -1611 577 -1610
rect 744 -1611 745 -1610
rect 786 -1611 787 -1610
rect 898 -1611 899 -1610
rect 912 -1611 913 -1610
rect 1045 -1611 1046 -1610
rect 1094 -1611 1095 -1610
rect 1244 -1611 1245 -1610
rect 1556 -1611 1557 -1610
rect 173 -1613 174 -1612
rect 744 -1613 745 -1612
rect 898 -1613 899 -1612
rect 1066 -1613 1067 -1612
rect 1087 -1613 1088 -1612
rect 1178 -1613 1179 -1612
rect 1486 -1613 1487 -1612
rect 1500 -1613 1501 -1612
rect 82 -1615 83 -1614
rect 1087 -1615 1088 -1614
rect 1500 -1615 1501 -1614
rect 1675 -1615 1676 -1614
rect 394 -1617 395 -1616
rect 835 -1617 836 -1616
rect 1017 -1617 1018 -1616
rect 1066 -1617 1067 -1616
rect 1675 -1617 1676 -1616
rect 1738 -1617 1739 -1616
rect 471 -1619 472 -1618
rect 534 -1619 535 -1618
rect 562 -1619 563 -1618
rect 1157 -1619 1158 -1618
rect 1738 -1619 1739 -1618
rect 1745 -1619 1746 -1618
rect 471 -1621 472 -1620
rect 527 -1621 528 -1620
rect 779 -1621 780 -1620
rect 1017 -1621 1018 -1620
rect 1045 -1621 1046 -1620
rect 1335 -1621 1336 -1620
rect 1745 -1621 1746 -1620
rect 1773 -1621 1774 -1620
rect 408 -1623 409 -1622
rect 527 -1623 528 -1622
rect 695 -1623 696 -1622
rect 779 -1623 780 -1622
rect 1143 -1623 1144 -1622
rect 1157 -1623 1158 -1622
rect 1759 -1623 1760 -1622
rect 1773 -1623 1774 -1622
rect 408 -1625 409 -1624
rect 590 -1625 591 -1624
rect 1052 -1625 1053 -1624
rect 1143 -1625 1144 -1624
rect 1759 -1625 1760 -1624
rect 2007 -1625 2008 -1624
rect 590 -1627 591 -1626
rect 716 -1627 717 -1626
rect 1052 -1627 1053 -1626
rect 1892 -1627 1893 -1626
rect 240 -1629 241 -1628
rect 1892 -1629 1893 -1628
rect 240 -1631 241 -1630
rect 401 -1631 402 -1630
rect 716 -1631 717 -1630
rect 758 -1631 759 -1630
rect 401 -1633 402 -1632
rect 436 -1633 437 -1632
rect 737 -1633 738 -1632
rect 758 -1633 759 -1632
rect 373 -1635 374 -1634
rect 436 -1635 437 -1634
rect 625 -1635 626 -1634
rect 737 -1635 738 -1634
rect 275 -1637 276 -1636
rect 373 -1637 374 -1636
rect 604 -1637 605 -1636
rect 625 -1637 626 -1636
rect 149 -1639 150 -1638
rect 275 -1639 276 -1638
rect 604 -1639 605 -1638
rect 639 -1639 640 -1638
rect 149 -1641 150 -1640
rect 170 -1641 171 -1640
rect 632 -1641 633 -1640
rect 639 -1641 640 -1640
rect 632 -1643 633 -1642
rect 831 -1643 832 -1642
rect 9 -1654 10 -1653
rect 663 -1654 664 -1653
rect 670 -1654 671 -1653
rect 716 -1654 717 -1653
rect 737 -1654 738 -1653
rect 1556 -1654 1557 -1653
rect 1843 -1654 1844 -1653
rect 1934 -1654 1935 -1653
rect 1937 -1654 1938 -1653
rect 1976 -1654 1977 -1653
rect 9 -1656 10 -1655
rect 128 -1656 129 -1655
rect 131 -1656 132 -1655
rect 1101 -1656 1102 -1655
rect 1206 -1656 1207 -1655
rect 1703 -1656 1704 -1655
rect 1815 -1656 1816 -1655
rect 1843 -1656 1844 -1655
rect 1850 -1656 1851 -1655
rect 1934 -1656 1935 -1655
rect 1941 -1656 1942 -1655
rect 1969 -1656 1970 -1655
rect 44 -1658 45 -1657
rect 79 -1658 80 -1657
rect 86 -1658 87 -1657
rect 275 -1658 276 -1657
rect 324 -1658 325 -1657
rect 558 -1658 559 -1657
rect 590 -1658 591 -1657
rect 831 -1658 832 -1657
rect 842 -1658 843 -1657
rect 1104 -1658 1105 -1657
rect 1206 -1658 1207 -1657
rect 1290 -1658 1291 -1657
rect 1332 -1658 1333 -1657
rect 1815 -1658 1816 -1657
rect 1850 -1658 1851 -1657
rect 1857 -1658 1858 -1657
rect 1944 -1658 1945 -1657
rect 1962 -1658 1963 -1657
rect 37 -1660 38 -1659
rect 44 -1660 45 -1659
rect 65 -1660 66 -1659
rect 177 -1660 178 -1659
rect 180 -1660 181 -1659
rect 359 -1660 360 -1659
rect 422 -1660 423 -1659
rect 425 -1660 426 -1659
rect 485 -1660 486 -1659
rect 684 -1660 685 -1659
rect 709 -1660 710 -1659
rect 1395 -1660 1396 -1659
rect 1468 -1660 1469 -1659
rect 1696 -1660 1697 -1659
rect 1857 -1660 1858 -1659
rect 1864 -1660 1865 -1659
rect 1948 -1660 1949 -1659
rect 1955 -1660 1956 -1659
rect 37 -1662 38 -1661
rect 58 -1662 59 -1661
rect 68 -1662 69 -1661
rect 534 -1662 535 -1661
rect 541 -1662 542 -1661
rect 772 -1662 773 -1661
rect 793 -1662 794 -1661
rect 1038 -1662 1039 -1661
rect 1055 -1662 1056 -1661
rect 1297 -1662 1298 -1661
rect 1332 -1662 1333 -1661
rect 1416 -1662 1417 -1661
rect 1468 -1662 1469 -1661
rect 1710 -1662 1711 -1661
rect 1822 -1662 1823 -1661
rect 1864 -1662 1865 -1661
rect 1941 -1662 1942 -1661
rect 1948 -1662 1949 -1661
rect 58 -1664 59 -1663
rect 429 -1664 430 -1663
rect 478 -1664 479 -1663
rect 485 -1664 486 -1663
rect 534 -1664 535 -1663
rect 625 -1664 626 -1663
rect 688 -1664 689 -1663
rect 709 -1664 710 -1663
rect 712 -1664 713 -1663
rect 1038 -1664 1039 -1663
rect 1076 -1664 1077 -1663
rect 1353 -1664 1354 -1663
rect 1395 -1664 1396 -1663
rect 1402 -1664 1403 -1663
rect 1416 -1664 1417 -1663
rect 1423 -1664 1424 -1663
rect 1500 -1664 1501 -1663
rect 1780 -1664 1781 -1663
rect 1794 -1664 1795 -1663
rect 1822 -1664 1823 -1663
rect 72 -1666 73 -1665
rect 82 -1666 83 -1665
rect 89 -1666 90 -1665
rect 1689 -1666 1690 -1665
rect 1696 -1666 1697 -1665
rect 1759 -1666 1760 -1665
rect 1766 -1666 1767 -1665
rect 1794 -1666 1795 -1665
rect 72 -1668 73 -1667
rect 660 -1668 661 -1667
rect 688 -1668 689 -1667
rect 989 -1668 990 -1667
rect 1083 -1668 1084 -1667
rect 1920 -1668 1921 -1667
rect 117 -1670 118 -1669
rect 1164 -1670 1165 -1669
rect 1220 -1670 1221 -1669
rect 1290 -1670 1291 -1669
rect 1297 -1670 1298 -1669
rect 1465 -1670 1466 -1669
rect 1556 -1670 1557 -1669
rect 1563 -1670 1564 -1669
rect 1640 -1670 1641 -1669
rect 1689 -1670 1690 -1669
rect 1731 -1670 1732 -1669
rect 1759 -1670 1760 -1669
rect 1906 -1670 1907 -1669
rect 1920 -1670 1921 -1669
rect 128 -1672 129 -1671
rect 968 -1672 969 -1671
rect 985 -1672 986 -1671
rect 1213 -1672 1214 -1671
rect 1286 -1672 1287 -1671
rect 1927 -1672 1928 -1671
rect 156 -1674 157 -1673
rect 394 -1674 395 -1673
rect 422 -1674 423 -1673
rect 499 -1674 500 -1673
rect 523 -1674 524 -1673
rect 1780 -1674 1781 -1673
rect 1899 -1674 1900 -1673
rect 1906 -1674 1907 -1673
rect 114 -1676 115 -1675
rect 394 -1676 395 -1675
rect 429 -1676 430 -1675
rect 436 -1676 437 -1675
rect 499 -1676 500 -1675
rect 1283 -1676 1284 -1675
rect 1335 -1676 1336 -1675
rect 1738 -1676 1739 -1675
rect 1752 -1676 1753 -1675
rect 1766 -1676 1767 -1675
rect 1892 -1676 1893 -1675
rect 1899 -1676 1900 -1675
rect 114 -1678 115 -1677
rect 443 -1678 444 -1677
rect 541 -1678 542 -1677
rect 740 -1678 741 -1677
rect 751 -1678 752 -1677
rect 1402 -1678 1403 -1677
rect 1423 -1678 1424 -1677
rect 1437 -1678 1438 -1677
rect 1521 -1678 1522 -1677
rect 1563 -1678 1564 -1677
rect 1619 -1678 1620 -1677
rect 1640 -1678 1641 -1677
rect 1654 -1678 1655 -1677
rect 1703 -1678 1704 -1677
rect 1717 -1678 1718 -1677
rect 1731 -1678 1732 -1677
rect 1752 -1678 1753 -1677
rect 1773 -1678 1774 -1677
rect 1787 -1678 1788 -1677
rect 1892 -1678 1893 -1677
rect 149 -1680 150 -1679
rect 436 -1680 437 -1679
rect 443 -1680 444 -1679
rect 646 -1680 647 -1679
rect 660 -1680 661 -1679
rect 940 -1680 941 -1679
rect 943 -1680 944 -1679
rect 1724 -1680 1725 -1679
rect 121 -1682 122 -1681
rect 149 -1682 150 -1681
rect 156 -1682 157 -1681
rect 317 -1682 318 -1681
rect 324 -1682 325 -1681
rect 408 -1682 409 -1681
rect 481 -1682 482 -1681
rect 751 -1682 752 -1681
rect 765 -1682 766 -1681
rect 863 -1682 864 -1681
rect 901 -1682 902 -1681
rect 1024 -1682 1025 -1681
rect 1087 -1682 1088 -1681
rect 1472 -1682 1473 -1681
rect 1493 -1682 1494 -1681
rect 1619 -1682 1620 -1681
rect 1626 -1682 1627 -1681
rect 1738 -1682 1739 -1681
rect 121 -1684 122 -1683
rect 814 -1684 815 -1683
rect 828 -1684 829 -1683
rect 1111 -1684 1112 -1683
rect 1185 -1684 1186 -1683
rect 1213 -1684 1214 -1683
rect 1241 -1684 1242 -1683
rect 1654 -1684 1655 -1683
rect 1675 -1684 1676 -1683
rect 1787 -1684 1788 -1683
rect 184 -1686 185 -1685
rect 667 -1686 668 -1685
rect 702 -1686 703 -1685
rect 793 -1686 794 -1685
rect 831 -1686 832 -1685
rect 1318 -1686 1319 -1685
rect 1339 -1686 1340 -1685
rect 1437 -1686 1438 -1685
rect 1472 -1686 1473 -1685
rect 1479 -1686 1480 -1685
rect 1591 -1686 1592 -1685
rect 1626 -1686 1627 -1685
rect 1682 -1686 1683 -1685
rect 1710 -1686 1711 -1685
rect 187 -1688 188 -1687
rect 1276 -1688 1277 -1687
rect 1311 -1688 1312 -1687
rect 1493 -1688 1494 -1687
rect 1542 -1688 1543 -1687
rect 1591 -1688 1592 -1687
rect 1668 -1688 1669 -1687
rect 1682 -1688 1683 -1687
rect 100 -1690 101 -1689
rect 1542 -1690 1543 -1689
rect 1661 -1690 1662 -1689
rect 1668 -1690 1669 -1689
rect 2 -1692 3 -1691
rect 100 -1692 101 -1691
rect 201 -1692 202 -1691
rect 649 -1692 650 -1691
rect 716 -1692 717 -1691
rect 1073 -1692 1074 -1691
rect 1101 -1692 1102 -1691
rect 1675 -1692 1676 -1691
rect 205 -1694 206 -1693
rect 208 -1694 209 -1693
rect 254 -1694 255 -1693
rect 397 -1694 398 -1693
rect 408 -1694 409 -1693
rect 562 -1694 563 -1693
rect 583 -1694 584 -1693
rect 625 -1694 626 -1693
rect 639 -1694 640 -1693
rect 814 -1694 815 -1693
rect 842 -1694 843 -1693
rect 877 -1694 878 -1693
rect 919 -1694 920 -1693
rect 1584 -1694 1585 -1693
rect 1661 -1694 1662 -1693
rect 1745 -1694 1746 -1693
rect 191 -1696 192 -1695
rect 254 -1696 255 -1695
rect 275 -1696 276 -1695
rect 450 -1696 451 -1695
rect 520 -1696 521 -1695
rect 702 -1696 703 -1695
rect 737 -1696 738 -1695
rect 810 -1696 811 -1695
rect 863 -1696 864 -1695
rect 912 -1696 913 -1695
rect 919 -1696 920 -1695
rect 1209 -1696 1210 -1695
rect 1241 -1696 1242 -1695
rect 1500 -1696 1501 -1695
rect 1584 -1696 1585 -1695
rect 1598 -1696 1599 -1695
rect 1745 -1696 1746 -1695
rect 1836 -1696 1837 -1695
rect 191 -1698 192 -1697
rect 418 -1698 419 -1697
rect 576 -1698 577 -1697
rect 639 -1698 640 -1697
rect 740 -1698 741 -1697
rect 1430 -1698 1431 -1697
rect 1479 -1698 1480 -1697
rect 1486 -1698 1487 -1697
rect 1598 -1698 1599 -1697
rect 1612 -1698 1613 -1697
rect 1808 -1698 1809 -1697
rect 1836 -1698 1837 -1697
rect 198 -1700 199 -1699
rect 450 -1700 451 -1699
rect 527 -1700 528 -1699
rect 576 -1700 577 -1699
rect 583 -1700 584 -1699
rect 681 -1700 682 -1699
rect 768 -1700 769 -1699
rect 989 -1700 990 -1699
rect 1024 -1700 1025 -1699
rect 1136 -1700 1137 -1699
rect 1185 -1700 1186 -1699
rect 1199 -1700 1200 -1699
rect 1244 -1700 1245 -1699
rect 1717 -1700 1718 -1699
rect 198 -1702 199 -1701
rect 849 -1702 850 -1701
rect 877 -1702 878 -1701
rect 961 -1702 962 -1701
rect 968 -1702 969 -1701
rect 1045 -1702 1046 -1701
rect 1073 -1702 1074 -1701
rect 1829 -1702 1830 -1701
rect 205 -1704 206 -1703
rect 492 -1704 493 -1703
rect 527 -1704 528 -1703
rect 632 -1704 633 -1703
rect 681 -1704 682 -1703
rect 1773 -1704 1774 -1703
rect 219 -1706 220 -1705
rect 1045 -1706 1046 -1705
rect 1129 -1706 1130 -1705
rect 1808 -1706 1809 -1705
rect 219 -1708 220 -1707
rect 261 -1708 262 -1707
rect 317 -1708 318 -1707
rect 338 -1708 339 -1707
rect 359 -1708 360 -1707
rect 457 -1708 458 -1707
rect 492 -1708 493 -1707
rect 730 -1708 731 -1707
rect 772 -1708 773 -1707
rect 1066 -1708 1067 -1707
rect 1122 -1708 1123 -1707
rect 1129 -1708 1130 -1707
rect 1132 -1708 1133 -1707
rect 1829 -1708 1830 -1707
rect 261 -1710 262 -1709
rect 506 -1710 507 -1709
rect 590 -1710 591 -1709
rect 597 -1710 598 -1709
rect 604 -1710 605 -1709
rect 667 -1710 668 -1709
rect 786 -1710 787 -1709
rect 1283 -1710 1284 -1709
rect 1311 -1710 1312 -1709
rect 1465 -1710 1466 -1709
rect 1612 -1710 1613 -1709
rect 1647 -1710 1648 -1709
rect 310 -1712 311 -1711
rect 338 -1712 339 -1711
rect 373 -1712 374 -1711
rect 418 -1712 419 -1711
rect 425 -1712 426 -1711
rect 786 -1712 787 -1711
rect 849 -1712 850 -1711
rect 898 -1712 899 -1711
rect 912 -1712 913 -1711
rect 926 -1712 927 -1711
rect 933 -1712 934 -1711
rect 1521 -1712 1522 -1711
rect 282 -1714 283 -1713
rect 310 -1714 311 -1713
rect 373 -1714 374 -1713
rect 401 -1714 402 -1713
rect 457 -1714 458 -1713
rect 464 -1714 465 -1713
rect 506 -1714 507 -1713
rect 723 -1714 724 -1713
rect 922 -1714 923 -1713
rect 947 -1714 948 -1713
rect 961 -1714 962 -1713
rect 1003 -1714 1004 -1713
rect 1041 -1714 1042 -1713
rect 1122 -1714 1123 -1713
rect 1136 -1714 1137 -1713
rect 1157 -1714 1158 -1713
rect 1199 -1714 1200 -1713
rect 1248 -1714 1249 -1713
rect 1269 -1714 1270 -1713
rect 1276 -1714 1277 -1713
rect 1318 -1714 1319 -1713
rect 1927 -1714 1928 -1713
rect 142 -1716 143 -1715
rect 401 -1716 402 -1715
rect 569 -1716 570 -1715
rect 604 -1716 605 -1715
rect 632 -1716 633 -1715
rect 698 -1716 699 -1715
rect 723 -1716 724 -1715
rect 870 -1716 871 -1715
rect 943 -1716 944 -1715
rect 1087 -1716 1088 -1715
rect 1157 -1716 1158 -1715
rect 1192 -1716 1193 -1715
rect 1244 -1716 1245 -1715
rect 1605 -1716 1606 -1715
rect 93 -1718 94 -1717
rect 142 -1718 143 -1717
rect 194 -1718 195 -1717
rect 1605 -1718 1606 -1717
rect 93 -1720 94 -1719
rect 600 -1720 601 -1719
rect 653 -1720 654 -1719
rect 926 -1720 927 -1719
rect 947 -1720 948 -1719
rect 982 -1720 983 -1719
rect 996 -1720 997 -1719
rect 1003 -1720 1004 -1719
rect 1066 -1720 1067 -1719
rect 1150 -1720 1151 -1719
rect 1192 -1720 1193 -1719
rect 1346 -1720 1347 -1719
rect 1353 -1720 1354 -1719
rect 1633 -1720 1634 -1719
rect 16 -1722 17 -1721
rect 982 -1722 983 -1721
rect 1010 -1722 1011 -1721
rect 1633 -1722 1634 -1721
rect 16 -1724 17 -1723
rect 170 -1724 171 -1723
rect 184 -1724 185 -1723
rect 1010 -1724 1011 -1723
rect 1150 -1724 1151 -1723
rect 1178 -1724 1179 -1723
rect 1248 -1724 1249 -1723
rect 1325 -1724 1326 -1723
rect 1339 -1724 1340 -1723
rect 1514 -1724 1515 -1723
rect 170 -1726 171 -1725
rect 268 -1726 269 -1725
rect 397 -1726 398 -1725
rect 821 -1726 822 -1725
rect 870 -1726 871 -1725
rect 905 -1726 906 -1725
rect 971 -1726 972 -1725
rect 1486 -1726 1487 -1725
rect 1507 -1726 1508 -1725
rect 1514 -1726 1515 -1725
rect 233 -1728 234 -1727
rect 464 -1728 465 -1727
rect 569 -1728 570 -1727
rect 611 -1728 612 -1727
rect 646 -1728 647 -1727
rect 996 -1728 997 -1727
rect 1171 -1728 1172 -1727
rect 1178 -1728 1179 -1727
rect 1227 -1728 1228 -1727
rect 1325 -1728 1326 -1727
rect 1356 -1728 1357 -1727
rect 1724 -1728 1725 -1727
rect 233 -1730 234 -1729
rect 303 -1730 304 -1729
rect 597 -1730 598 -1729
rect 1164 -1730 1165 -1729
rect 1220 -1730 1221 -1729
rect 1356 -1730 1357 -1729
rect 1388 -1730 1389 -1729
rect 1430 -1730 1431 -1729
rect 1507 -1730 1508 -1729
rect 1577 -1730 1578 -1729
rect 240 -1732 241 -1731
rect 303 -1732 304 -1731
rect 611 -1732 612 -1731
rect 618 -1732 619 -1731
rect 653 -1732 654 -1731
rect 1304 -1732 1305 -1731
rect 1388 -1732 1389 -1731
rect 1444 -1732 1445 -1731
rect 226 -1734 227 -1733
rect 618 -1734 619 -1733
rect 821 -1734 822 -1733
rect 835 -1734 836 -1733
rect 891 -1734 892 -1733
rect 1346 -1734 1347 -1733
rect 1444 -1734 1445 -1733
rect 1535 -1734 1536 -1733
rect 226 -1736 227 -1735
rect 331 -1736 332 -1735
rect 807 -1736 808 -1735
rect 835 -1736 836 -1735
rect 891 -1736 892 -1735
rect 954 -1736 955 -1735
rect 1080 -1736 1081 -1735
rect 1171 -1736 1172 -1735
rect 1227 -1736 1228 -1735
rect 1234 -1736 1235 -1735
rect 1269 -1736 1270 -1735
rect 1360 -1736 1361 -1735
rect 1528 -1736 1529 -1735
rect 1535 -1736 1536 -1735
rect 240 -1738 241 -1737
rect 415 -1738 416 -1737
rect 898 -1738 899 -1737
rect 1577 -1738 1578 -1737
rect 247 -1740 248 -1739
rect 282 -1740 283 -1739
rect 331 -1740 332 -1739
rect 352 -1740 353 -1739
rect 905 -1740 906 -1739
rect 975 -1740 976 -1739
rect 1234 -1740 1235 -1739
rect 1367 -1740 1368 -1739
rect 1528 -1740 1529 -1739
rect 1549 -1740 1550 -1739
rect 247 -1742 248 -1741
rect 345 -1742 346 -1741
rect 352 -1742 353 -1741
rect 548 -1742 549 -1741
rect 933 -1742 934 -1741
rect 1080 -1742 1081 -1741
rect 1304 -1742 1305 -1741
rect 1647 -1742 1648 -1741
rect 268 -1744 269 -1743
rect 366 -1744 367 -1743
rect 513 -1744 514 -1743
rect 548 -1744 549 -1743
rect 954 -1744 955 -1743
rect 1878 -1744 1879 -1743
rect 23 -1746 24 -1745
rect 366 -1746 367 -1745
rect 513 -1746 514 -1745
rect 674 -1746 675 -1745
rect 975 -1746 976 -1745
rect 1017 -1746 1018 -1745
rect 1307 -1746 1308 -1745
rect 1878 -1746 1879 -1745
rect 23 -1748 24 -1747
rect 544 -1748 545 -1747
rect 674 -1748 675 -1747
rect 779 -1748 780 -1747
rect 1052 -1748 1053 -1747
rect 1307 -1748 1308 -1747
rect 1360 -1748 1361 -1747
rect 1363 -1748 1364 -1747
rect 1367 -1748 1368 -1747
rect 1458 -1748 1459 -1747
rect 289 -1750 290 -1749
rect 345 -1750 346 -1749
rect 744 -1750 745 -1749
rect 1017 -1750 1018 -1749
rect 1052 -1750 1053 -1749
rect 1108 -1750 1109 -1749
rect 1374 -1750 1375 -1749
rect 1458 -1750 1459 -1749
rect 289 -1752 290 -1751
rect 380 -1752 381 -1751
rect 744 -1752 745 -1751
rect 758 -1752 759 -1751
rect 779 -1752 780 -1751
rect 1031 -1752 1032 -1751
rect 1374 -1752 1375 -1751
rect 1381 -1752 1382 -1751
rect 1409 -1752 1410 -1751
rect 1549 -1752 1550 -1751
rect 107 -1754 108 -1753
rect 380 -1754 381 -1753
rect 758 -1754 759 -1753
rect 884 -1754 885 -1753
rect 1031 -1754 1032 -1753
rect 1094 -1754 1095 -1753
rect 1115 -1754 1116 -1753
rect 1409 -1754 1410 -1753
rect 107 -1756 108 -1755
rect 135 -1756 136 -1755
rect 695 -1756 696 -1755
rect 1094 -1756 1095 -1755
rect 1115 -1756 1116 -1755
rect 1143 -1756 1144 -1755
rect 1381 -1756 1382 -1755
rect 1846 -1756 1847 -1755
rect 135 -1758 136 -1757
rect 163 -1758 164 -1757
rect 565 -1758 566 -1757
rect 1143 -1758 1144 -1757
rect 163 -1760 164 -1759
rect 212 -1760 213 -1759
rect 695 -1760 696 -1759
rect 1059 -1760 1060 -1759
rect 212 -1762 213 -1761
rect 387 -1762 388 -1761
rect 1059 -1762 1060 -1761
rect 1255 -1762 1256 -1761
rect 296 -1764 297 -1763
rect 387 -1764 388 -1763
rect 516 -1764 517 -1763
rect 1255 -1764 1256 -1763
rect 296 -1766 297 -1765
rect 471 -1766 472 -1765
rect 30 -1768 31 -1767
rect 471 -1768 472 -1767
rect 30 -1770 31 -1769
rect 555 -1770 556 -1769
rect 555 -1772 556 -1771
rect 887 -1772 888 -1771
rect 65 -1783 66 -1782
rect 75 -1783 76 -1782
rect 93 -1783 94 -1782
rect 145 -1783 146 -1782
rect 170 -1783 171 -1782
rect 523 -1783 524 -1782
rect 527 -1783 528 -1782
rect 530 -1783 531 -1782
rect 555 -1783 556 -1782
rect 793 -1783 794 -1782
rect 810 -1783 811 -1782
rect 1927 -1783 1928 -1782
rect 1955 -1783 1956 -1782
rect 1997 -1783 1998 -1782
rect 2011 -1783 2012 -1782
rect 2018 -1783 2019 -1782
rect 65 -1785 66 -1784
rect 275 -1785 276 -1784
rect 282 -1785 283 -1784
rect 481 -1785 482 -1784
rect 506 -1785 507 -1784
rect 555 -1785 556 -1784
rect 597 -1785 598 -1784
rect 870 -1785 871 -1784
rect 884 -1785 885 -1784
rect 1689 -1785 1690 -1784
rect 1878 -1785 1879 -1784
rect 1955 -1785 1956 -1784
rect 1962 -1785 1963 -1784
rect 2018 -1785 2019 -1784
rect 93 -1787 94 -1786
rect 107 -1787 108 -1786
rect 114 -1787 115 -1786
rect 191 -1787 192 -1786
rect 198 -1787 199 -1786
rect 877 -1787 878 -1786
rect 884 -1787 885 -1786
rect 2004 -1787 2005 -1786
rect 107 -1789 108 -1788
rect 499 -1789 500 -1788
rect 527 -1789 528 -1788
rect 1073 -1789 1074 -1788
rect 1080 -1789 1081 -1788
rect 1689 -1789 1690 -1788
rect 1878 -1789 1879 -1788
rect 1941 -1789 1942 -1788
rect 1969 -1789 1970 -1788
rect 2025 -1789 2026 -1788
rect 114 -1791 115 -1790
rect 212 -1791 213 -1790
rect 254 -1791 255 -1790
rect 691 -1791 692 -1790
rect 695 -1791 696 -1790
rect 926 -1791 927 -1790
rect 943 -1791 944 -1790
rect 1493 -1791 1494 -1790
rect 1566 -1791 1567 -1790
rect 1885 -1791 1886 -1790
rect 1892 -1791 1893 -1790
rect 1962 -1791 1963 -1790
rect 58 -1793 59 -1792
rect 212 -1793 213 -1792
rect 254 -1793 255 -1792
rect 289 -1793 290 -1792
rect 310 -1793 311 -1792
rect 807 -1793 808 -1792
rect 870 -1793 871 -1792
rect 933 -1793 934 -1792
rect 985 -1793 986 -1792
rect 1570 -1793 1571 -1792
rect 1829 -1793 1830 -1792
rect 1885 -1793 1886 -1792
rect 1899 -1793 1900 -1792
rect 1969 -1793 1970 -1792
rect 16 -1795 17 -1794
rect 58 -1795 59 -1794
rect 128 -1795 129 -1794
rect 135 -1795 136 -1794
rect 138 -1795 139 -1794
rect 289 -1795 290 -1794
rect 352 -1795 353 -1794
rect 488 -1795 489 -1794
rect 499 -1795 500 -1794
rect 625 -1795 626 -1794
rect 649 -1795 650 -1794
rect 814 -1795 815 -1794
rect 898 -1795 899 -1794
rect 1038 -1795 1039 -1794
rect 1059 -1795 1060 -1794
rect 1076 -1795 1077 -1794
rect 1080 -1795 1081 -1794
rect 1087 -1795 1088 -1794
rect 1090 -1795 1091 -1794
rect 1206 -1795 1207 -1794
rect 1209 -1795 1210 -1794
rect 1626 -1795 1627 -1794
rect 1731 -1795 1732 -1794
rect 1829 -1795 1830 -1794
rect 1843 -1795 1844 -1794
rect 1892 -1795 1893 -1794
rect 1906 -1795 1907 -1794
rect 1983 -1795 1984 -1794
rect 9 -1797 10 -1796
rect 135 -1797 136 -1796
rect 142 -1797 143 -1796
rect 310 -1797 311 -1796
rect 352 -1797 353 -1796
rect 359 -1797 360 -1796
rect 366 -1797 367 -1796
rect 562 -1797 563 -1796
rect 583 -1797 584 -1796
rect 597 -1797 598 -1796
rect 600 -1797 601 -1796
rect 702 -1797 703 -1796
rect 719 -1797 720 -1796
rect 730 -1797 731 -1796
rect 751 -1797 752 -1796
rect 877 -1797 878 -1796
rect 908 -1797 909 -1796
rect 1094 -1797 1095 -1796
rect 1104 -1797 1105 -1796
rect 1444 -1797 1445 -1796
rect 1468 -1797 1469 -1796
rect 1920 -1797 1921 -1796
rect 16 -1799 17 -1798
rect 51 -1799 52 -1798
rect 121 -1799 122 -1798
rect 625 -1799 626 -1798
rect 639 -1799 640 -1798
rect 702 -1799 703 -1798
rect 730 -1799 731 -1798
rect 1381 -1799 1382 -1798
rect 1409 -1799 1410 -1798
rect 1990 -1799 1991 -1798
rect 37 -1801 38 -1800
rect 51 -1801 52 -1800
rect 79 -1801 80 -1800
rect 121 -1801 122 -1800
rect 131 -1801 132 -1800
rect 366 -1801 367 -1800
rect 387 -1801 388 -1800
rect 639 -1801 640 -1800
rect 681 -1801 682 -1800
rect 793 -1801 794 -1800
rect 814 -1801 815 -1800
rect 842 -1801 843 -1800
rect 954 -1801 955 -1800
rect 1038 -1801 1039 -1800
rect 1059 -1801 1060 -1800
rect 1290 -1801 1291 -1800
rect 1304 -1801 1305 -1800
rect 1773 -1801 1774 -1800
rect 1850 -1801 1851 -1800
rect 1906 -1801 1907 -1800
rect 1913 -1801 1914 -1800
rect 1920 -1801 1921 -1800
rect 37 -1803 38 -1802
rect 142 -1803 143 -1802
rect 156 -1803 157 -1802
rect 282 -1803 283 -1802
rect 387 -1803 388 -1802
rect 509 -1803 510 -1802
rect 562 -1803 563 -1802
rect 604 -1803 605 -1802
rect 632 -1803 633 -1802
rect 681 -1803 682 -1802
rect 684 -1803 685 -1802
rect 936 -1803 937 -1802
rect 1017 -1803 1018 -1802
rect 1094 -1803 1095 -1802
rect 1104 -1803 1105 -1802
rect 1213 -1803 1214 -1802
rect 1244 -1803 1245 -1802
rect 1640 -1803 1641 -1802
rect 1717 -1803 1718 -1802
rect 1773 -1803 1774 -1802
rect 1815 -1803 1816 -1802
rect 1850 -1803 1851 -1802
rect 1871 -1803 1872 -1802
rect 1941 -1803 1942 -1802
rect 79 -1805 80 -1804
rect 653 -1805 654 -1804
rect 765 -1805 766 -1804
rect 842 -1805 843 -1804
rect 1073 -1805 1074 -1804
rect 1171 -1805 1172 -1804
rect 1248 -1805 1249 -1804
rect 1290 -1805 1291 -1804
rect 1304 -1805 1305 -1804
rect 1437 -1805 1438 -1804
rect 1535 -1805 1536 -1804
rect 1843 -1805 1844 -1804
rect 156 -1807 157 -1806
rect 408 -1807 409 -1806
rect 415 -1807 416 -1806
rect 919 -1807 920 -1806
rect 1108 -1807 1109 -1806
rect 1976 -1807 1977 -1806
rect 170 -1809 171 -1808
rect 982 -1809 983 -1808
rect 1111 -1809 1112 -1808
rect 1192 -1809 1193 -1808
rect 1269 -1809 1270 -1808
rect 1353 -1809 1354 -1808
rect 1360 -1809 1361 -1808
rect 1738 -1809 1739 -1808
rect 1745 -1809 1746 -1808
rect 1899 -1809 1900 -1808
rect 177 -1811 178 -1810
rect 275 -1811 276 -1810
rect 401 -1811 402 -1810
rect 940 -1811 941 -1810
rect 1136 -1811 1137 -1810
rect 1171 -1811 1172 -1810
rect 1185 -1811 1186 -1810
rect 1248 -1811 1249 -1810
rect 1262 -1811 1263 -1810
rect 1269 -1811 1270 -1810
rect 1283 -1811 1284 -1810
rect 1360 -1811 1361 -1810
rect 1363 -1811 1364 -1810
rect 1927 -1811 1928 -1810
rect 177 -1813 178 -1812
rect 394 -1813 395 -1812
rect 404 -1813 405 -1812
rect 415 -1813 416 -1812
rect 429 -1813 430 -1812
rect 513 -1813 514 -1812
rect 583 -1813 584 -1812
rect 1101 -1813 1102 -1812
rect 1115 -1813 1116 -1812
rect 1136 -1813 1137 -1812
rect 1150 -1813 1151 -1812
rect 1185 -1813 1186 -1812
rect 1276 -1813 1277 -1812
rect 1283 -1813 1284 -1812
rect 1307 -1813 1308 -1812
rect 1787 -1813 1788 -1812
rect 1794 -1813 1795 -1812
rect 1871 -1813 1872 -1812
rect 191 -1815 192 -1814
rect 219 -1815 220 -1814
rect 240 -1815 241 -1814
rect 394 -1815 395 -1814
rect 408 -1815 409 -1814
rect 1125 -1815 1126 -1814
rect 1150 -1815 1151 -1814
rect 1444 -1815 1445 -1814
rect 1535 -1815 1536 -1814
rect 1780 -1815 1781 -1814
rect 1822 -1815 1823 -1814
rect 1913 -1815 1914 -1814
rect 201 -1817 202 -1816
rect 296 -1817 297 -1816
rect 380 -1817 381 -1816
rect 401 -1817 402 -1816
rect 429 -1817 430 -1816
rect 548 -1817 549 -1816
rect 604 -1817 605 -1816
rect 723 -1817 724 -1816
rect 751 -1817 752 -1816
rect 1108 -1817 1109 -1816
rect 1157 -1817 1158 -1816
rect 1192 -1817 1193 -1816
rect 1311 -1817 1312 -1816
rect 1493 -1817 1494 -1816
rect 1563 -1817 1564 -1816
rect 1570 -1817 1571 -1816
rect 1577 -1817 1578 -1816
rect 1745 -1817 1746 -1816
rect 1759 -1817 1760 -1816
rect 1780 -1817 1781 -1816
rect 1801 -1817 1802 -1816
rect 1822 -1817 1823 -1816
rect 187 -1819 188 -1818
rect 1801 -1819 1802 -1818
rect 219 -1821 220 -1820
rect 443 -1821 444 -1820
rect 450 -1821 451 -1820
rect 695 -1821 696 -1820
rect 723 -1821 724 -1820
rect 828 -1821 829 -1820
rect 831 -1821 832 -1820
rect 1437 -1821 1438 -1820
rect 1598 -1821 1599 -1820
rect 1815 -1821 1816 -1820
rect 23 -1823 24 -1822
rect 828 -1823 829 -1822
rect 863 -1823 864 -1822
rect 1311 -1823 1312 -1822
rect 1318 -1823 1319 -1822
rect 1703 -1823 1704 -1822
rect 1738 -1823 1739 -1822
rect 1752 -1823 1753 -1822
rect 1766 -1823 1767 -1822
rect 1794 -1823 1795 -1822
rect 23 -1825 24 -1824
rect 614 -1825 615 -1824
rect 632 -1825 633 -1824
rect 667 -1825 668 -1824
rect 765 -1825 766 -1824
rect 863 -1825 864 -1824
rect 891 -1825 892 -1824
rect 940 -1825 941 -1824
rect 975 -1825 976 -1824
rect 1157 -1825 1158 -1824
rect 1164 -1825 1165 -1824
rect 1213 -1825 1214 -1824
rect 1321 -1825 1322 -1824
rect 1626 -1825 1627 -1824
rect 1654 -1825 1655 -1824
rect 1717 -1825 1718 -1824
rect 72 -1827 73 -1826
rect 450 -1827 451 -1826
rect 464 -1827 465 -1826
rect 520 -1827 521 -1826
rect 541 -1827 542 -1826
rect 548 -1827 549 -1826
rect 576 -1827 577 -1826
rect 667 -1827 668 -1826
rect 768 -1827 769 -1826
rect 1458 -1827 1459 -1826
rect 1486 -1827 1487 -1826
rect 1766 -1827 1767 -1826
rect 44 -1829 45 -1828
rect 72 -1829 73 -1828
rect 100 -1829 101 -1828
rect 975 -1829 976 -1828
rect 1024 -1829 1025 -1828
rect 1164 -1829 1165 -1828
rect 1178 -1829 1179 -1828
rect 1262 -1829 1263 -1828
rect 1325 -1829 1326 -1828
rect 1381 -1829 1382 -1828
rect 1409 -1829 1410 -1828
rect 1549 -1829 1550 -1828
rect 1598 -1829 1599 -1828
rect 1661 -1829 1662 -1828
rect 1696 -1829 1697 -1828
rect 1703 -1829 1704 -1828
rect 30 -1831 31 -1830
rect 1024 -1831 1025 -1830
rect 1083 -1831 1084 -1830
rect 1752 -1831 1753 -1830
rect 30 -1833 31 -1832
rect 226 -1833 227 -1832
rect 240 -1833 241 -1832
rect 338 -1833 339 -1832
rect 373 -1833 374 -1832
rect 443 -1833 444 -1832
rect 464 -1833 465 -1832
rect 611 -1833 612 -1832
rect 772 -1833 773 -1832
rect 1017 -1833 1018 -1832
rect 1143 -1833 1144 -1832
rect 1178 -1833 1179 -1832
rect 1255 -1833 1256 -1832
rect 1325 -1833 1326 -1832
rect 1339 -1833 1340 -1832
rect 1577 -1833 1578 -1832
rect 1605 -1833 1606 -1832
rect 1640 -1833 1641 -1832
rect 1661 -1833 1662 -1832
rect 1836 -1833 1837 -1832
rect 44 -1835 45 -1834
rect 397 -1835 398 -1834
rect 436 -1835 437 -1834
rect 653 -1835 654 -1834
rect 772 -1835 773 -1834
rect 996 -1835 997 -1834
rect 1122 -1835 1123 -1834
rect 1143 -1835 1144 -1834
rect 1199 -1835 1200 -1834
rect 1255 -1835 1256 -1834
rect 1430 -1835 1431 -1834
rect 1731 -1835 1732 -1834
rect 1808 -1835 1809 -1834
rect 1836 -1835 1837 -1834
rect 184 -1837 185 -1836
rect 1318 -1837 1319 -1836
rect 1451 -1837 1452 -1836
rect 1458 -1837 1459 -1836
rect 1479 -1837 1480 -1836
rect 1486 -1837 1487 -1836
rect 1633 -1837 1634 -1836
rect 1654 -1837 1655 -1836
rect 1682 -1837 1683 -1836
rect 1696 -1837 1697 -1836
rect 1710 -1837 1711 -1836
rect 1808 -1837 1809 -1836
rect 163 -1839 164 -1838
rect 184 -1839 185 -1838
rect 205 -1839 206 -1838
rect 373 -1839 374 -1838
rect 380 -1839 381 -1838
rect 422 -1839 423 -1838
rect 485 -1839 486 -1838
rect 541 -1839 542 -1838
rect 558 -1839 559 -1838
rect 1199 -1839 1200 -1838
rect 1234 -1839 1235 -1838
rect 1339 -1839 1340 -1838
rect 1367 -1839 1368 -1838
rect 1479 -1839 1480 -1838
rect 1542 -1839 1543 -1838
rect 1710 -1839 1711 -1838
rect 163 -1841 164 -1840
rect 516 -1841 517 -1840
rect 520 -1841 521 -1840
rect 688 -1841 689 -1840
rect 891 -1841 892 -1840
rect 1241 -1841 1242 -1840
rect 1367 -1841 1368 -1840
rect 1374 -1841 1375 -1840
rect 1388 -1841 1389 -1840
rect 1451 -1841 1452 -1840
rect 1556 -1841 1557 -1840
rect 1633 -1841 1634 -1840
rect 1668 -1841 1669 -1840
rect 1682 -1841 1683 -1840
rect 205 -1843 206 -1842
rect 233 -1843 234 -1842
rect 261 -1843 262 -1842
rect 359 -1843 360 -1842
rect 478 -1843 479 -1842
rect 1542 -1843 1543 -1842
rect 1556 -1843 1557 -1842
rect 1944 -1843 1945 -1842
rect 149 -1845 150 -1844
rect 261 -1845 262 -1844
rect 296 -1845 297 -1844
rect 478 -1845 479 -1844
rect 485 -1845 486 -1844
rect 1787 -1845 1788 -1844
rect 149 -1847 150 -1846
rect 887 -1847 888 -1846
rect 912 -1847 913 -1846
rect 919 -1847 920 -1846
rect 933 -1847 934 -1846
rect 1759 -1847 1760 -1846
rect 226 -1849 227 -1848
rect 345 -1849 346 -1848
rect 492 -1849 493 -1848
rect 887 -1849 888 -1848
rect 912 -1849 913 -1848
rect 961 -1849 962 -1848
rect 996 -1849 997 -1848
rect 1003 -1849 1004 -1848
rect 1045 -1849 1046 -1848
rect 1430 -1849 1431 -1848
rect 1647 -1849 1648 -1848
rect 1668 -1849 1669 -1848
rect 233 -1851 234 -1850
rect 268 -1851 269 -1850
rect 331 -1851 332 -1850
rect 436 -1851 437 -1850
rect 492 -1851 493 -1850
rect 618 -1851 619 -1850
rect 779 -1851 780 -1850
rect 1003 -1851 1004 -1850
rect 1031 -1851 1032 -1850
rect 1045 -1851 1046 -1850
rect 1122 -1851 1123 -1850
rect 1864 -1851 1865 -1850
rect 86 -1853 87 -1852
rect 268 -1853 269 -1852
rect 324 -1853 325 -1852
rect 331 -1853 332 -1852
rect 513 -1853 514 -1852
rect 1153 -1853 1154 -1852
rect 1220 -1853 1221 -1852
rect 1234 -1853 1235 -1852
rect 1241 -1853 1242 -1852
rect 1465 -1853 1466 -1852
rect 1612 -1853 1613 -1852
rect 1647 -1853 1648 -1852
rect 86 -1855 87 -1854
rect 1223 -1855 1224 -1854
rect 1374 -1855 1375 -1854
rect 1395 -1855 1396 -1854
rect 1423 -1855 1424 -1854
rect 1612 -1855 1613 -1854
rect 247 -1857 248 -1856
rect 345 -1857 346 -1856
rect 530 -1857 531 -1856
rect 1115 -1857 1116 -1856
rect 1346 -1857 1347 -1856
rect 1395 -1857 1396 -1856
rect 1416 -1857 1417 -1856
rect 1423 -1857 1424 -1856
rect 1465 -1857 1466 -1856
rect 1528 -1857 1529 -1856
rect 247 -1859 248 -1858
rect 2014 -1859 2015 -1858
rect 317 -1861 318 -1860
rect 324 -1861 325 -1860
rect 579 -1861 580 -1860
rect 1549 -1861 1550 -1860
rect 317 -1863 318 -1862
rect 457 -1863 458 -1862
rect 611 -1863 612 -1862
rect 1605 -1863 1606 -1862
rect 198 -1865 199 -1864
rect 457 -1865 458 -1864
rect 618 -1865 619 -1864
rect 786 -1865 787 -1864
rect 905 -1865 906 -1864
rect 961 -1865 962 -1864
rect 1031 -1865 1032 -1864
rect 1066 -1865 1067 -1864
rect 1111 -1865 1112 -1864
rect 1864 -1865 1865 -1864
rect 422 -1867 423 -1866
rect 905 -1867 906 -1866
rect 954 -1867 955 -1866
rect 1220 -1867 1221 -1866
rect 1297 -1867 1298 -1866
rect 1346 -1867 1347 -1866
rect 1388 -1867 1389 -1866
rect 1402 -1867 1403 -1866
rect 1416 -1867 1417 -1866
rect 1934 -1867 1935 -1866
rect 779 -1869 780 -1868
rect 856 -1869 857 -1868
rect 1052 -1869 1053 -1868
rect 1066 -1869 1067 -1868
rect 1227 -1869 1228 -1868
rect 1297 -1869 1298 -1868
rect 1332 -1869 1333 -1868
rect 1402 -1869 1403 -1868
rect 1528 -1869 1529 -1868
rect 1591 -1869 1592 -1868
rect 1857 -1869 1858 -1868
rect 1934 -1869 1935 -1868
rect 61 -1871 62 -1870
rect 1227 -1871 1228 -1870
rect 1507 -1871 1508 -1870
rect 1591 -1871 1592 -1870
rect 68 -1873 69 -1872
rect 1857 -1873 1858 -1872
rect 103 -1875 104 -1874
rect 856 -1875 857 -1874
rect 989 -1875 990 -1874
rect 1052 -1875 1053 -1874
rect 1507 -1875 1508 -1874
rect 1514 -1875 1515 -1874
rect 534 -1877 535 -1876
rect 989 -1877 990 -1876
rect 1472 -1877 1473 -1876
rect 1514 -1877 1515 -1876
rect 534 -1879 535 -1878
rect 758 -1879 759 -1878
rect 786 -1879 787 -1878
rect 849 -1879 850 -1878
rect 1472 -1879 1473 -1878
rect 1675 -1879 1676 -1878
rect 674 -1881 675 -1880
rect 849 -1881 850 -1880
rect 1675 -1881 1676 -1880
rect 1724 -1881 1725 -1880
rect 418 -1883 419 -1882
rect 1724 -1883 1725 -1882
rect 674 -1885 675 -1884
rect 709 -1885 710 -1884
rect 737 -1885 738 -1884
rect 1332 -1885 1333 -1884
rect 565 -1887 566 -1886
rect 709 -1887 710 -1886
rect 758 -1887 759 -1886
rect 821 -1887 822 -1886
rect 646 -1889 647 -1888
rect 737 -1889 738 -1888
rect 821 -1889 822 -1888
rect 835 -1889 836 -1888
rect 569 -1891 570 -1890
rect 646 -1891 647 -1890
rect 800 -1891 801 -1890
rect 835 -1891 836 -1890
rect 471 -1893 472 -1892
rect 569 -1893 570 -1892
rect 716 -1893 717 -1892
rect 800 -1893 801 -1892
rect 471 -1895 472 -1894
rect 1948 -1895 1949 -1894
rect 716 -1897 717 -1896
rect 926 -1897 927 -1896
rect 1563 -1897 1564 -1896
rect 1948 -1897 1949 -1896
rect 2 -1908 3 -1907
rect 226 -1908 227 -1907
rect 313 -1908 314 -1907
rect 450 -1908 451 -1907
rect 478 -1908 479 -1907
rect 555 -1908 556 -1907
rect 562 -1908 563 -1907
rect 576 -1908 577 -1907
rect 614 -1908 615 -1907
rect 989 -1908 990 -1907
rect 1024 -1908 1025 -1907
rect 1381 -1908 1382 -1907
rect 1454 -1908 1455 -1907
rect 1871 -1908 1872 -1907
rect 5 -1910 6 -1909
rect 68 -1910 69 -1909
rect 79 -1910 80 -1909
rect 509 -1910 510 -1909
rect 537 -1910 538 -1909
rect 1115 -1910 1116 -1909
rect 1153 -1910 1154 -1909
rect 1808 -1910 1809 -1909
rect 1871 -1910 1872 -1909
rect 1899 -1910 1900 -1909
rect 9 -1912 10 -1911
rect 37 -1912 38 -1911
rect 44 -1912 45 -1911
rect 138 -1912 139 -1911
rect 142 -1912 143 -1911
rect 1444 -1912 1445 -1911
rect 1535 -1912 1536 -1911
rect 1808 -1912 1809 -1911
rect 1899 -1912 1900 -1911
rect 1948 -1912 1949 -1911
rect 37 -1914 38 -1913
rect 541 -1914 542 -1913
rect 555 -1914 556 -1913
rect 737 -1914 738 -1913
rect 744 -1914 745 -1913
rect 1101 -1914 1102 -1913
rect 1108 -1914 1109 -1913
rect 1297 -1914 1298 -1913
rect 1367 -1914 1368 -1913
rect 1381 -1914 1382 -1913
rect 1444 -1914 1445 -1913
rect 1451 -1914 1452 -1913
rect 1535 -1914 1536 -1913
rect 2011 -1914 2012 -1913
rect 44 -1916 45 -1915
rect 289 -1916 290 -1915
rect 317 -1916 318 -1915
rect 744 -1916 745 -1915
rect 828 -1916 829 -1915
rect 933 -1916 934 -1915
rect 964 -1916 965 -1915
rect 1311 -1916 1312 -1915
rect 1451 -1916 1452 -1915
rect 1528 -1916 1529 -1915
rect 1563 -1916 1564 -1915
rect 1570 -1916 1571 -1915
rect 1948 -1916 1949 -1915
rect 1976 -1916 1977 -1915
rect 58 -1918 59 -1917
rect 695 -1918 696 -1917
rect 716 -1918 717 -1917
rect 737 -1918 738 -1917
rect 772 -1918 773 -1917
rect 1570 -1918 1571 -1917
rect 1976 -1918 1977 -1917
rect 2018 -1918 2019 -1917
rect 79 -1920 80 -1919
rect 471 -1920 472 -1919
rect 481 -1920 482 -1919
rect 1241 -1920 1242 -1919
rect 1283 -1920 1284 -1919
rect 1311 -1920 1312 -1919
rect 1528 -1920 1529 -1919
rect 1752 -1920 1753 -1919
rect 23 -1922 24 -1921
rect 471 -1922 472 -1921
rect 485 -1922 486 -1921
rect 908 -1922 909 -1921
rect 919 -1922 920 -1921
rect 933 -1922 934 -1921
rect 982 -1922 983 -1921
rect 1633 -1922 1634 -1921
rect 23 -1924 24 -1923
rect 114 -1924 115 -1923
rect 135 -1924 136 -1923
rect 726 -1924 727 -1923
rect 730 -1924 731 -1923
rect 894 -1924 895 -1923
rect 905 -1924 906 -1923
rect 1815 -1924 1816 -1923
rect 86 -1926 87 -1925
rect 289 -1926 290 -1925
rect 317 -1926 318 -1925
rect 758 -1926 759 -1925
rect 779 -1926 780 -1925
rect 905 -1926 906 -1925
rect 982 -1926 983 -1925
rect 1136 -1926 1137 -1925
rect 1143 -1926 1144 -1925
rect 1241 -1926 1242 -1925
rect 1293 -1926 1294 -1925
rect 1843 -1926 1844 -1925
rect 100 -1928 101 -1927
rect 268 -1928 269 -1927
rect 338 -1928 339 -1927
rect 828 -1928 829 -1927
rect 845 -1928 846 -1927
rect 1157 -1928 1158 -1927
rect 1199 -1928 1200 -1927
rect 1367 -1928 1368 -1927
rect 1566 -1928 1567 -1927
rect 1584 -1928 1585 -1927
rect 1633 -1928 1634 -1927
rect 1654 -1928 1655 -1927
rect 1815 -1928 1816 -1927
rect 1822 -1928 1823 -1927
rect 1843 -1928 1844 -1927
rect 1885 -1928 1886 -1927
rect 100 -1930 101 -1929
rect 527 -1930 528 -1929
rect 562 -1930 563 -1929
rect 583 -1930 584 -1929
rect 632 -1930 633 -1929
rect 768 -1930 769 -1929
rect 779 -1930 780 -1929
rect 856 -1930 857 -1929
rect 880 -1930 881 -1929
rect 1038 -1930 1039 -1929
rect 1090 -1930 1091 -1929
rect 1990 -1930 1991 -1929
rect 30 -1932 31 -1931
rect 527 -1932 528 -1931
rect 583 -1932 584 -1931
rect 597 -1932 598 -1931
rect 660 -1932 661 -1931
rect 663 -1932 664 -1931
rect 688 -1932 689 -1931
rect 1395 -1932 1396 -1931
rect 1472 -1932 1473 -1931
rect 1654 -1932 1655 -1931
rect 1822 -1932 1823 -1931
rect 1836 -1932 1837 -1931
rect 1885 -1932 1886 -1931
rect 1927 -1932 1928 -1931
rect 1990 -1932 1991 -1931
rect 2025 -1932 2026 -1931
rect 30 -1934 31 -1933
rect 513 -1934 514 -1933
rect 660 -1934 661 -1933
rect 667 -1934 668 -1933
rect 681 -1934 682 -1933
rect 688 -1934 689 -1933
rect 698 -1934 699 -1933
rect 1283 -1934 1284 -1933
rect 1297 -1934 1298 -1933
rect 1493 -1934 1494 -1933
rect 1584 -1934 1585 -1933
rect 1605 -1934 1606 -1933
rect 1836 -1934 1837 -1933
rect 1850 -1934 1851 -1933
rect 1927 -1934 1928 -1933
rect 1955 -1934 1956 -1933
rect 16 -1936 17 -1935
rect 513 -1936 514 -1935
rect 674 -1936 675 -1935
rect 681 -1936 682 -1935
rect 709 -1936 710 -1935
rect 716 -1936 717 -1935
rect 719 -1936 720 -1935
rect 814 -1936 815 -1935
rect 856 -1936 857 -1935
rect 1080 -1936 1081 -1935
rect 1094 -1936 1095 -1935
rect 1115 -1936 1116 -1935
rect 1129 -1936 1130 -1935
rect 1143 -1936 1144 -1935
rect 1157 -1936 1158 -1935
rect 1171 -1936 1172 -1935
rect 1206 -1936 1207 -1935
rect 1216 -1936 1217 -1935
rect 1220 -1936 1221 -1935
rect 1731 -1936 1732 -1935
rect 1955 -1936 1956 -1935
rect 1983 -1936 1984 -1935
rect 65 -1938 66 -1937
rect 632 -1938 633 -1937
rect 674 -1938 675 -1937
rect 702 -1938 703 -1937
rect 709 -1938 710 -1937
rect 1059 -1938 1060 -1937
rect 1066 -1938 1067 -1937
rect 1080 -1938 1081 -1937
rect 1094 -1938 1095 -1937
rect 1318 -1938 1319 -1937
rect 1395 -1938 1396 -1937
rect 1500 -1938 1501 -1937
rect 1661 -1938 1662 -1937
rect 1850 -1938 1851 -1937
rect 103 -1940 104 -1939
rect 975 -1940 976 -1939
rect 989 -1940 990 -1939
rect 1031 -1940 1032 -1939
rect 1052 -1940 1053 -1939
rect 1059 -1940 1060 -1939
rect 1108 -1940 1109 -1939
rect 1514 -1940 1515 -1939
rect 16 -1942 17 -1941
rect 1031 -1942 1032 -1941
rect 1136 -1942 1137 -1941
rect 1178 -1942 1179 -1941
rect 1206 -1942 1207 -1941
rect 1521 -1942 1522 -1941
rect 107 -1944 108 -1943
rect 114 -1944 115 -1943
rect 135 -1944 136 -1943
rect 387 -1944 388 -1943
rect 401 -1944 402 -1943
rect 1209 -1944 1210 -1943
rect 1220 -1944 1221 -1943
rect 1416 -1944 1417 -1943
rect 1472 -1944 1473 -1943
rect 1542 -1944 1543 -1943
rect 93 -1946 94 -1945
rect 387 -1946 388 -1945
rect 415 -1946 416 -1945
rect 541 -1946 542 -1945
rect 639 -1946 640 -1945
rect 702 -1946 703 -1945
rect 730 -1946 731 -1945
rect 1878 -1946 1879 -1945
rect 51 -1948 52 -1947
rect 93 -1948 94 -1947
rect 107 -1948 108 -1947
rect 985 -1948 986 -1947
rect 1003 -1948 1004 -1947
rect 1066 -1948 1067 -1947
rect 1164 -1948 1165 -1947
rect 1199 -1948 1200 -1947
rect 1223 -1948 1224 -1947
rect 1920 -1948 1921 -1947
rect 51 -1950 52 -1949
rect 691 -1950 692 -1949
rect 733 -1950 734 -1949
rect 1752 -1950 1753 -1949
rect 1878 -1950 1879 -1949
rect 1906 -1950 1907 -1949
rect 1920 -1950 1921 -1949
rect 1997 -1950 1998 -1949
rect 142 -1952 143 -1951
rect 1829 -1952 1830 -1951
rect 1906 -1952 1907 -1951
rect 1934 -1952 1935 -1951
rect 145 -1954 146 -1953
rect 240 -1954 241 -1953
rect 408 -1954 409 -1953
rect 415 -1954 416 -1953
rect 464 -1954 465 -1953
rect 639 -1954 640 -1953
rect 758 -1954 759 -1953
rect 961 -1954 962 -1953
rect 1010 -1954 1011 -1953
rect 1024 -1954 1025 -1953
rect 1027 -1954 1028 -1953
rect 1801 -1954 1802 -1953
rect 1934 -1954 1935 -1953
rect 1962 -1954 1963 -1953
rect 86 -1956 87 -1955
rect 145 -1956 146 -1955
rect 198 -1956 199 -1955
rect 261 -1956 262 -1955
rect 408 -1956 409 -1955
rect 751 -1956 752 -1955
rect 800 -1956 801 -1955
rect 1052 -1956 1053 -1955
rect 1164 -1956 1165 -1955
rect 1248 -1956 1249 -1955
rect 1262 -1956 1263 -1955
rect 1500 -1956 1501 -1955
rect 1521 -1956 1522 -1955
rect 1549 -1956 1550 -1955
rect 1787 -1956 1788 -1955
rect 1829 -1956 1830 -1955
rect 170 -1958 171 -1957
rect 261 -1958 262 -1957
rect 464 -1958 465 -1957
rect 775 -1958 776 -1957
rect 807 -1958 808 -1957
rect 1038 -1958 1039 -1957
rect 1171 -1958 1172 -1957
rect 1255 -1958 1256 -1957
rect 1265 -1958 1266 -1957
rect 1731 -1958 1732 -1957
rect 1794 -1958 1795 -1957
rect 1801 -1958 1802 -1957
rect 170 -1960 171 -1959
rect 775 -1960 776 -1959
rect 807 -1960 808 -1959
rect 835 -1960 836 -1959
rect 849 -1960 850 -1959
rect 1129 -1960 1130 -1959
rect 1178 -1960 1179 -1959
rect 1185 -1960 1186 -1959
rect 1216 -1960 1217 -1959
rect 1549 -1960 1550 -1959
rect 1598 -1960 1599 -1959
rect 1794 -1960 1795 -1959
rect 198 -1962 199 -1961
rect 1262 -1962 1263 -1961
rect 1290 -1962 1291 -1961
rect 1318 -1962 1319 -1961
rect 1416 -1962 1417 -1961
rect 1423 -1962 1424 -1961
rect 1479 -1962 1480 -1961
rect 1514 -1962 1515 -1961
rect 1542 -1962 1543 -1961
rect 1556 -1962 1557 -1961
rect 212 -1964 213 -1963
rect 243 -1964 244 -1963
rect 268 -1964 269 -1963
rect 1290 -1964 1291 -1963
rect 1409 -1964 1410 -1963
rect 1423 -1964 1424 -1963
rect 1465 -1964 1466 -1963
rect 1556 -1964 1557 -1963
rect 184 -1966 185 -1965
rect 212 -1966 213 -1965
rect 226 -1966 227 -1965
rect 303 -1966 304 -1965
rect 485 -1966 486 -1965
rect 653 -1966 654 -1965
rect 814 -1966 815 -1965
rect 1332 -1966 1333 -1965
rect 1388 -1966 1389 -1965
rect 1409 -1966 1410 -1965
rect 1486 -1966 1487 -1965
rect 1493 -1966 1494 -1965
rect 1507 -1966 1508 -1965
rect 1598 -1966 1599 -1965
rect 184 -1968 185 -1967
rect 191 -1968 192 -1967
rect 205 -1968 206 -1967
rect 303 -1968 304 -1967
rect 457 -1968 458 -1967
rect 653 -1968 654 -1967
rect 821 -1968 822 -1967
rect 835 -1968 836 -1967
rect 849 -1968 850 -1967
rect 1073 -1968 1074 -1967
rect 1087 -1968 1088 -1967
rect 1465 -1968 1466 -1967
rect 1486 -1968 1487 -1967
rect 1647 -1968 1648 -1967
rect 163 -1970 164 -1969
rect 191 -1970 192 -1969
rect 205 -1970 206 -1969
rect 579 -1970 580 -1969
rect 618 -1970 619 -1969
rect 751 -1970 752 -1969
rect 793 -1970 794 -1969
rect 1073 -1970 1074 -1969
rect 1087 -1970 1088 -1969
rect 1353 -1970 1354 -1969
rect 1360 -1970 1361 -1969
rect 1507 -1970 1508 -1969
rect 1647 -1970 1648 -1969
rect 1689 -1970 1690 -1969
rect 72 -1972 73 -1971
rect 163 -1972 164 -1971
rect 341 -1972 342 -1971
rect 618 -1972 619 -1971
rect 793 -1972 794 -1971
rect 954 -1972 955 -1971
rect 961 -1972 962 -1971
rect 1787 -1972 1788 -1971
rect 61 -1974 62 -1973
rect 72 -1974 73 -1973
rect 380 -1974 381 -1973
rect 457 -1974 458 -1973
rect 499 -1974 500 -1973
rect 597 -1974 598 -1973
rect 821 -1974 822 -1973
rect 1192 -1974 1193 -1973
rect 1237 -1974 1238 -1973
rect 1279 -1974 1280 -1973
rect 1325 -1974 1326 -1973
rect 1332 -1974 1333 -1973
rect 1374 -1974 1375 -1973
rect 1388 -1974 1389 -1973
rect 1689 -1974 1690 -1973
rect 1759 -1974 1760 -1973
rect 380 -1976 381 -1975
rect 436 -1976 437 -1975
rect 443 -1976 444 -1975
rect 499 -1976 500 -1975
rect 506 -1976 507 -1975
rect 1248 -1976 1249 -1975
rect 1269 -1976 1270 -1975
rect 1360 -1976 1361 -1975
rect 247 -1978 248 -1977
rect 436 -1978 437 -1977
rect 754 -1978 755 -1977
rect 1269 -1978 1270 -1977
rect 1276 -1978 1277 -1977
rect 1479 -1978 1480 -1977
rect 177 -1980 178 -1979
rect 1276 -1980 1277 -1979
rect 1304 -1980 1305 -1979
rect 1325 -1980 1326 -1979
rect 1339 -1980 1340 -1979
rect 1374 -1980 1375 -1979
rect 177 -1982 178 -1981
rect 366 -1982 367 -1981
rect 863 -1982 864 -1981
rect 1003 -1982 1004 -1981
rect 1150 -1982 1151 -1981
rect 1759 -1982 1760 -1981
rect 247 -1984 248 -1983
rect 324 -1984 325 -1983
rect 352 -1984 353 -1983
rect 443 -1984 444 -1983
rect 611 -1984 612 -1983
rect 1150 -1984 1151 -1983
rect 1192 -1984 1193 -1983
rect 1913 -1984 1914 -1983
rect 254 -1986 255 -1985
rect 366 -1986 367 -1985
rect 611 -1986 612 -1985
rect 817 -1986 818 -1985
rect 863 -1986 864 -1985
rect 2004 -1986 2005 -1985
rect 254 -1988 255 -1987
rect 310 -1988 311 -1987
rect 324 -1988 325 -1987
rect 422 -1988 423 -1987
rect 866 -1988 867 -1987
rect 1962 -1988 1963 -1987
rect 275 -1990 276 -1989
rect 506 -1990 507 -1989
rect 877 -1990 878 -1989
rect 975 -1990 976 -1989
rect 996 -1990 997 -1989
rect 1010 -1990 1011 -1989
rect 1255 -1990 1256 -1989
rect 1913 -1990 1914 -1989
rect 275 -1992 276 -1991
rect 870 -1992 871 -1991
rect 877 -1992 878 -1991
rect 1577 -1992 1578 -1991
rect 296 -1994 297 -1993
rect 310 -1994 311 -1993
rect 345 -1994 346 -1993
rect 422 -1994 423 -1993
rect 842 -1994 843 -1993
rect 870 -1994 871 -1993
rect 884 -1994 885 -1993
rect 1612 -1994 1613 -1993
rect 121 -1996 122 -1995
rect 296 -1996 297 -1995
rect 345 -1996 346 -1995
rect 488 -1996 489 -1995
rect 604 -1996 605 -1995
rect 884 -1996 885 -1995
rect 887 -1996 888 -1995
rect 1983 -1996 1984 -1995
rect 121 -1998 122 -1997
rect 429 -1998 430 -1997
rect 604 -1998 605 -1997
rect 1045 -1998 1046 -1997
rect 1339 -1998 1340 -1997
rect 1346 -1998 1347 -1997
rect 1577 -1998 1578 -1997
rect 1591 -1998 1592 -1997
rect 1612 -1998 1613 -1997
rect 1675 -1998 1676 -1997
rect 219 -2000 220 -1999
rect 429 -2000 430 -1999
rect 842 -2000 843 -1999
rect 1710 -2000 1711 -1999
rect 219 -2002 220 -2001
rect 534 -2002 535 -2001
rect 912 -2002 913 -2001
rect 954 -2002 955 -2001
rect 968 -2002 969 -2001
rect 996 -2002 997 -2001
rect 1017 -2002 1018 -2001
rect 1045 -2002 1046 -2001
rect 1111 -2002 1112 -2001
rect 1710 -2002 1711 -2001
rect 352 -2004 353 -2003
rect 569 -2004 570 -2003
rect 800 -2004 801 -2003
rect 968 -2004 969 -2003
rect 1017 -2004 1018 -2003
rect 1437 -2004 1438 -2003
rect 1591 -2004 1592 -2003
rect 1668 -2004 1669 -2003
rect 1675 -2004 1676 -2003
rect 1703 -2004 1704 -2003
rect 492 -2006 493 -2005
rect 569 -2006 570 -2005
rect 912 -2006 913 -2005
rect 936 -2006 937 -2005
rect 1111 -2006 1112 -2005
rect 1353 -2006 1354 -2005
rect 1402 -2006 1403 -2005
rect 1437 -2006 1438 -2005
rect 1668 -2006 1669 -2005
rect 1696 -2006 1697 -2005
rect 1703 -2006 1704 -2005
rect 1738 -2006 1739 -2005
rect 359 -2008 360 -2007
rect 492 -2008 493 -2007
rect 520 -2008 521 -2007
rect 534 -2008 535 -2007
rect 723 -2008 724 -2007
rect 1402 -2008 1403 -2007
rect 1640 -2008 1641 -2007
rect 1696 -2008 1697 -2007
rect 331 -2010 332 -2009
rect 359 -2010 360 -2009
rect 394 -2010 395 -2009
rect 520 -2010 521 -2009
rect 530 -2010 531 -2009
rect 1738 -2010 1739 -2009
rect 149 -2012 150 -2011
rect 331 -2012 332 -2011
rect 723 -2012 724 -2011
rect 1661 -2012 1662 -2011
rect 149 -2014 150 -2013
rect 222 -2014 223 -2013
rect 233 -2014 234 -2013
rect 394 -2014 395 -2013
rect 919 -2014 920 -2013
rect 1304 -2014 1305 -2013
rect 1640 -2014 1641 -2013
rect 1682 -2014 1683 -2013
rect 233 -2016 234 -2015
rect 282 -2016 283 -2015
rect 922 -2016 923 -2015
rect 1605 -2016 1606 -2015
rect 1682 -2016 1683 -2015
rect 1724 -2016 1725 -2015
rect 282 -2018 283 -2017
rect 373 -2018 374 -2017
rect 926 -2018 927 -2017
rect 1185 -2018 1186 -2017
rect 1234 -2018 1235 -2017
rect 1346 -2018 1347 -2017
rect 1724 -2018 1725 -2017
rect 1766 -2018 1767 -2017
rect 373 -2020 374 -2019
rect 1122 -2020 1123 -2019
rect 1766 -2020 1767 -2019
rect 1773 -2020 1774 -2019
rect 898 -2022 899 -2021
rect 926 -2022 927 -2021
rect 940 -2022 941 -2021
rect 1122 -2022 1123 -2021
rect 1773 -2022 1774 -2021
rect 1780 -2022 1781 -2021
rect 625 -2024 626 -2023
rect 940 -2024 941 -2023
rect 1619 -2024 1620 -2023
rect 1780 -2024 1781 -2023
rect 548 -2026 549 -2025
rect 625 -2026 626 -2025
rect 786 -2026 787 -2025
rect 898 -2026 899 -2025
rect 1619 -2026 1620 -2025
rect 1717 -2026 1718 -2025
rect 548 -2028 549 -2027
rect 646 -2028 647 -2027
rect 772 -2028 773 -2027
rect 786 -2028 787 -2027
rect 1626 -2028 1627 -2027
rect 1717 -2028 1718 -2027
rect 590 -2030 591 -2029
rect 646 -2030 647 -2029
rect 1626 -2030 1627 -2029
rect 1864 -2030 1865 -2029
rect 590 -2032 591 -2031
rect 765 -2032 766 -2031
rect 1104 -2032 1105 -2031
rect 1864 -2032 1865 -2031
rect 765 -2034 766 -2033
rect 891 -2034 892 -2033
rect 891 -2036 892 -2035
rect 1857 -2036 1858 -2035
rect 1857 -2038 1858 -2037
rect 1892 -2038 1893 -2037
rect 1892 -2040 1893 -2039
rect 1941 -2040 1942 -2039
rect 1941 -2042 1942 -2041
rect 1969 -2042 1970 -2041
rect 761 -2044 762 -2043
rect 1969 -2044 1970 -2043
rect 2 -2055 3 -2054
rect 338 -2055 339 -2054
rect 352 -2055 353 -2054
rect 726 -2055 727 -2054
rect 733 -2055 734 -2054
rect 1101 -2055 1102 -2054
rect 1108 -2055 1109 -2054
rect 1514 -2055 1515 -2054
rect 1920 -2055 1921 -2054
rect 1976 -2055 1977 -2054
rect 2 -2057 3 -2056
rect 205 -2057 206 -2056
rect 219 -2057 220 -2056
rect 537 -2057 538 -2056
rect 548 -2057 549 -2056
rect 814 -2057 815 -2056
rect 817 -2057 818 -2056
rect 982 -2057 983 -2056
rect 1087 -2057 1088 -2056
rect 1234 -2057 1235 -2056
rect 1237 -2057 1238 -2056
rect 1493 -2057 1494 -2056
rect 23 -2059 24 -2058
rect 142 -2059 143 -2058
rect 149 -2059 150 -2058
rect 219 -2059 220 -2058
rect 222 -2059 223 -2058
rect 702 -2059 703 -2058
rect 723 -2059 724 -2058
rect 926 -2059 927 -2058
rect 961 -2059 962 -2058
rect 1500 -2059 1501 -2058
rect 9 -2061 10 -2060
rect 142 -2061 143 -2060
rect 177 -2061 178 -2060
rect 240 -2061 241 -2060
rect 352 -2061 353 -2060
rect 394 -2061 395 -2060
rect 401 -2061 402 -2060
rect 702 -2061 703 -2060
rect 723 -2061 724 -2060
rect 996 -2061 997 -2060
rect 1087 -2061 1088 -2060
rect 1185 -2061 1186 -2060
rect 1241 -2061 1242 -2060
rect 1262 -2061 1263 -2060
rect 1265 -2061 1266 -2060
rect 1850 -2061 1851 -2060
rect 23 -2063 24 -2062
rect 110 -2063 111 -2062
rect 117 -2063 118 -2062
rect 1507 -2063 1508 -2062
rect 1850 -2063 1851 -2062
rect 1927 -2063 1928 -2062
rect 30 -2065 31 -2064
rect 313 -2065 314 -2064
rect 394 -2065 395 -2064
rect 709 -2065 710 -2064
rect 751 -2065 752 -2064
rect 1129 -2065 1130 -2064
rect 1139 -2065 1140 -2064
rect 1437 -2065 1438 -2064
rect 1493 -2065 1494 -2064
rect 1605 -2065 1606 -2064
rect 30 -2067 31 -2066
rect 509 -2067 510 -2066
rect 520 -2067 521 -2066
rect 649 -2067 650 -2066
rect 695 -2067 696 -2066
rect 1038 -2067 1039 -2066
rect 1101 -2067 1102 -2066
rect 1178 -2067 1179 -2066
rect 1241 -2067 1242 -2066
rect 1304 -2067 1305 -2066
rect 1360 -2067 1361 -2066
rect 1454 -2067 1455 -2066
rect 1500 -2067 1501 -2066
rect 1759 -2067 1760 -2066
rect 37 -2069 38 -2068
rect 439 -2069 440 -2068
rect 450 -2069 451 -2068
rect 499 -2069 500 -2068
rect 530 -2069 531 -2068
rect 1402 -2069 1403 -2068
rect 1437 -2069 1438 -2068
rect 1472 -2069 1473 -2068
rect 1507 -2069 1508 -2068
rect 1710 -2069 1711 -2068
rect 1759 -2069 1760 -2068
rect 1857 -2069 1858 -2068
rect 51 -2071 52 -2070
rect 698 -2071 699 -2070
rect 751 -2071 752 -2070
rect 1108 -2071 1109 -2070
rect 1129 -2071 1130 -2070
rect 1136 -2071 1137 -2070
rect 1143 -2071 1144 -2070
rect 1262 -2071 1263 -2070
rect 1290 -2071 1291 -2070
rect 1353 -2071 1354 -2070
rect 1363 -2071 1364 -2070
rect 1829 -2071 1830 -2070
rect 1857 -2071 1858 -2070
rect 1941 -2071 1942 -2070
rect 51 -2073 52 -2072
rect 261 -2073 262 -2072
rect 303 -2073 304 -2072
rect 401 -2073 402 -2072
rect 408 -2073 409 -2072
rect 838 -2073 839 -2072
rect 845 -2073 846 -2072
rect 1514 -2073 1515 -2072
rect 1605 -2073 1606 -2072
rect 1773 -2073 1774 -2072
rect 1829 -2073 1830 -2072
rect 1899 -2073 1900 -2072
rect 65 -2075 66 -2074
rect 1402 -2075 1403 -2074
rect 1710 -2075 1711 -2074
rect 1836 -2075 1837 -2074
rect 1899 -2075 1900 -2074
rect 1990 -2075 1991 -2074
rect 65 -2077 66 -2076
rect 380 -2077 381 -2076
rect 415 -2077 416 -2076
rect 730 -2077 731 -2076
rect 761 -2077 762 -2076
rect 786 -2077 787 -2076
rect 807 -2077 808 -2076
rect 814 -2077 815 -2076
rect 891 -2077 892 -2076
rect 1031 -2077 1032 -2076
rect 1038 -2077 1039 -2076
rect 1052 -2077 1053 -2076
rect 1143 -2077 1144 -2076
rect 1213 -2077 1214 -2076
rect 1255 -2077 1256 -2076
rect 1311 -2077 1312 -2076
rect 1353 -2077 1354 -2076
rect 1570 -2077 1571 -2076
rect 1773 -2077 1774 -2076
rect 1843 -2077 1844 -2076
rect 44 -2079 45 -2078
rect 380 -2079 381 -2078
rect 422 -2079 423 -2078
rect 450 -2079 451 -2078
rect 492 -2079 493 -2078
rect 499 -2079 500 -2078
rect 548 -2079 549 -2078
rect 562 -2079 563 -2078
rect 583 -2079 584 -2078
rect 807 -2079 808 -2078
rect 919 -2079 920 -2078
rect 1598 -2079 1599 -2078
rect 1843 -2079 1844 -2078
rect 1913 -2079 1914 -2078
rect 44 -2081 45 -2080
rect 86 -2081 87 -2080
rect 89 -2081 90 -2080
rect 324 -2081 325 -2080
rect 422 -2081 423 -2080
rect 975 -2081 976 -2080
rect 978 -2081 979 -2080
rect 1374 -2081 1375 -2080
rect 1475 -2081 1476 -2080
rect 1836 -2081 1837 -2080
rect 68 -2083 69 -2082
rect 471 -2083 472 -2082
rect 492 -2083 493 -2082
rect 541 -2083 542 -2082
rect 562 -2083 563 -2082
rect 1111 -2083 1112 -2082
rect 1160 -2083 1161 -2082
rect 1304 -2083 1305 -2082
rect 1311 -2083 1312 -2082
rect 1388 -2083 1389 -2082
rect 1570 -2083 1571 -2082
rect 1661 -2083 1662 -2082
rect 1717 -2083 1718 -2082
rect 1913 -2083 1914 -2082
rect 79 -2085 80 -2084
rect 82 -2085 83 -2084
rect 86 -2085 87 -2084
rect 513 -2085 514 -2084
rect 583 -2085 584 -2084
rect 646 -2085 647 -2084
rect 695 -2085 696 -2084
rect 716 -2085 717 -2084
rect 730 -2085 731 -2084
rect 964 -2085 965 -2084
rect 968 -2085 969 -2084
rect 1479 -2085 1480 -2084
rect 1661 -2085 1662 -2084
rect 1724 -2085 1725 -2084
rect 79 -2087 80 -2086
rect 135 -2087 136 -2086
rect 163 -2087 164 -2086
rect 303 -2087 304 -2086
rect 436 -2087 437 -2086
rect 513 -2087 514 -2086
rect 590 -2087 591 -2086
rect 1398 -2087 1399 -2086
rect 1479 -2087 1480 -2086
rect 1584 -2087 1585 -2086
rect 1633 -2087 1634 -2086
rect 1724 -2087 1725 -2086
rect 93 -2089 94 -2088
rect 520 -2089 521 -2088
rect 593 -2089 594 -2088
rect 744 -2089 745 -2088
rect 772 -2089 773 -2088
rect 1066 -2089 1067 -2088
rect 1171 -2089 1172 -2088
rect 1185 -2089 1186 -2088
rect 1213 -2089 1214 -2088
rect 1339 -2089 1340 -2088
rect 1374 -2089 1375 -2088
rect 1906 -2089 1907 -2088
rect 33 -2091 34 -2090
rect 744 -2091 745 -2090
rect 772 -2091 773 -2090
rect 1111 -2091 1112 -2090
rect 1171 -2091 1172 -2090
rect 1346 -2091 1347 -2090
rect 1388 -2091 1389 -2090
rect 1458 -2091 1459 -2090
rect 1584 -2091 1585 -2090
rect 1668 -2091 1669 -2090
rect 1675 -2091 1676 -2090
rect 1906 -2091 1907 -2090
rect 93 -2093 94 -2092
rect 387 -2093 388 -2092
rect 467 -2093 468 -2092
rect 968 -2093 969 -2092
rect 971 -2093 972 -2092
rect 1423 -2093 1424 -2092
rect 1458 -2093 1459 -2092
rect 1542 -2093 1543 -2092
rect 1675 -2093 1676 -2092
rect 1731 -2093 1732 -2092
rect 96 -2095 97 -2094
rect 390 -2095 391 -2094
rect 597 -2095 598 -2094
rect 849 -2095 850 -2094
rect 852 -2095 853 -2094
rect 1633 -2095 1634 -2094
rect 1703 -2095 1704 -2094
rect 1731 -2095 1732 -2094
rect 16 -2097 17 -2096
rect 849 -2097 850 -2096
rect 905 -2097 906 -2096
rect 919 -2097 920 -2096
rect 922 -2097 923 -2096
rect 1122 -2097 1123 -2096
rect 1178 -2097 1179 -2096
rect 1416 -2097 1417 -2096
rect 1542 -2097 1543 -2096
rect 1619 -2097 1620 -2096
rect 1703 -2097 1704 -2096
rect 1794 -2097 1795 -2096
rect 16 -2099 17 -2098
rect 243 -2099 244 -2098
rect 247 -2099 248 -2098
rect 261 -2099 262 -2098
rect 268 -2099 269 -2098
rect 408 -2099 409 -2098
rect 506 -2099 507 -2098
rect 597 -2099 598 -2098
rect 604 -2099 605 -2098
rect 709 -2099 710 -2098
rect 779 -2099 780 -2098
rect 891 -2099 892 -2098
rect 926 -2099 927 -2098
rect 933 -2099 934 -2098
rect 954 -2099 955 -2098
rect 961 -2099 962 -2098
rect 975 -2099 976 -2098
rect 1010 -2099 1011 -2098
rect 1031 -2099 1032 -2098
rect 1206 -2099 1207 -2098
rect 1220 -2099 1221 -2098
rect 1339 -2099 1340 -2098
rect 1346 -2099 1347 -2098
rect 1923 -2099 1924 -2098
rect 128 -2101 129 -2100
rect 149 -2101 150 -2100
rect 163 -2101 164 -2100
rect 310 -2101 311 -2100
rect 324 -2101 325 -2100
rect 590 -2101 591 -2100
rect 618 -2101 619 -2100
rect 716 -2101 717 -2100
rect 786 -2101 787 -2100
rect 1164 -2101 1165 -2100
rect 1192 -2101 1193 -2100
rect 1206 -2101 1207 -2100
rect 1220 -2101 1221 -2100
rect 1283 -2101 1284 -2100
rect 1395 -2101 1396 -2100
rect 1423 -2101 1424 -2100
rect 1619 -2101 1620 -2100
rect 1766 -2101 1767 -2100
rect 1794 -2101 1795 -2100
rect 1815 -2101 1816 -2100
rect 107 -2103 108 -2102
rect 128 -2103 129 -2102
rect 135 -2103 136 -2102
rect 156 -2103 157 -2102
rect 177 -2103 178 -2102
rect 289 -2103 290 -2102
rect 341 -2103 342 -2102
rect 618 -2103 619 -2102
rect 639 -2103 640 -2102
rect 758 -2103 759 -2102
rect 884 -2103 885 -2102
rect 905 -2103 906 -2102
rect 933 -2103 934 -2102
rect 1017 -2103 1018 -2102
rect 1052 -2103 1053 -2102
rect 1696 -2103 1697 -2102
rect 1717 -2103 1718 -2102
rect 1745 -2103 1746 -2102
rect 1766 -2103 1767 -2102
rect 1822 -2103 1823 -2102
rect 156 -2105 157 -2104
rect 184 -2105 185 -2104
rect 191 -2105 192 -2104
rect 471 -2105 472 -2104
rect 506 -2105 507 -2104
rect 779 -2105 780 -2104
rect 870 -2105 871 -2104
rect 884 -2105 885 -2104
rect 954 -2105 955 -2104
rect 1297 -2105 1298 -2104
rect 1409 -2105 1410 -2104
rect 1668 -2105 1669 -2104
rect 1696 -2105 1697 -2104
rect 1969 -2105 1970 -2104
rect 184 -2107 185 -2106
rect 842 -2107 843 -2106
rect 982 -2107 983 -2106
rect 1003 -2107 1004 -2106
rect 1010 -2107 1011 -2106
rect 1059 -2107 1060 -2106
rect 1066 -2107 1067 -2106
rect 1745 -2107 1746 -2106
rect 1815 -2107 1816 -2106
rect 1892 -2107 1893 -2106
rect 191 -2109 192 -2108
rect 359 -2109 360 -2108
rect 485 -2109 486 -2108
rect 842 -2109 843 -2108
rect 989 -2109 990 -2108
rect 1017 -2109 1018 -2108
rect 1059 -2109 1060 -2108
rect 1157 -2109 1158 -2108
rect 1192 -2109 1193 -2108
rect 1325 -2109 1326 -2108
rect 1409 -2109 1410 -2108
rect 1465 -2109 1466 -2108
rect 1822 -2109 1823 -2108
rect 1948 -2109 1949 -2108
rect 198 -2111 199 -2110
rect 310 -2111 311 -2110
rect 485 -2111 486 -2110
rect 569 -2111 570 -2110
rect 576 -2111 577 -2110
rect 604 -2111 605 -2110
rect 611 -2111 612 -2110
rect 1164 -2111 1165 -2110
rect 1248 -2111 1249 -2110
rect 1416 -2111 1417 -2110
rect 1465 -2111 1466 -2110
rect 1577 -2111 1578 -2110
rect 1892 -2111 1893 -2110
rect 1983 -2111 1984 -2110
rect 198 -2113 199 -2112
rect 226 -2113 227 -2112
rect 236 -2113 237 -2112
rect 863 -2113 864 -2112
rect 989 -2113 990 -2112
rect 1045 -2113 1046 -2112
rect 1115 -2113 1116 -2112
rect 1122 -2113 1123 -2112
rect 1157 -2113 1158 -2112
rect 1878 -2113 1879 -2112
rect 205 -2115 206 -2114
rect 971 -2115 972 -2114
rect 996 -2115 997 -2114
rect 1024 -2115 1025 -2114
rect 1045 -2115 1046 -2114
rect 1377 -2115 1378 -2114
rect 1577 -2115 1578 -2114
rect 1808 -2115 1809 -2114
rect 226 -2117 227 -2116
rect 233 -2117 234 -2116
rect 247 -2117 248 -2116
rect 345 -2117 346 -2116
rect 527 -2117 528 -2116
rect 1283 -2117 1284 -2116
rect 1325 -2117 1326 -2116
rect 1381 -2117 1382 -2116
rect 1738 -2117 1739 -2116
rect 1878 -2117 1879 -2116
rect 212 -2119 213 -2118
rect 233 -2119 234 -2118
rect 268 -2119 269 -2118
rect 373 -2119 374 -2118
rect 527 -2119 528 -2118
rect 877 -2119 878 -2118
rect 1003 -2119 1004 -2118
rect 1073 -2119 1074 -2118
rect 1115 -2119 1116 -2118
rect 1199 -2119 1200 -2118
rect 1248 -2119 1249 -2118
rect 1367 -2119 1368 -2118
rect 1381 -2119 1382 -2118
rect 1591 -2119 1592 -2118
rect 1738 -2119 1739 -2118
rect 1801 -2119 1802 -2118
rect 1808 -2119 1809 -2118
rect 1934 -2119 1935 -2118
rect 145 -2121 146 -2120
rect 1367 -2121 1368 -2120
rect 1591 -2121 1592 -2120
rect 1682 -2121 1683 -2120
rect 1801 -2121 1802 -2120
rect 1885 -2121 1886 -2120
rect 170 -2123 171 -2122
rect 373 -2123 374 -2122
rect 415 -2123 416 -2122
rect 877 -2123 878 -2122
rect 1024 -2123 1025 -2122
rect 1521 -2123 1522 -2122
rect 1682 -2123 1683 -2122
rect 1752 -2123 1753 -2122
rect 1885 -2123 1886 -2122
rect 1962 -2123 1963 -2122
rect 40 -2125 41 -2124
rect 170 -2125 171 -2124
rect 212 -2125 213 -2124
rect 366 -2125 367 -2124
rect 576 -2125 577 -2124
rect 653 -2125 654 -2124
rect 737 -2125 738 -2124
rect 758 -2125 759 -2124
rect 863 -2125 864 -2124
rect 1069 -2125 1070 -2124
rect 1073 -2125 1074 -2124
rect 1080 -2125 1081 -2124
rect 1199 -2125 1200 -2124
rect 1276 -2125 1277 -2124
rect 1486 -2125 1487 -2124
rect 1521 -2125 1522 -2124
rect 1689 -2125 1690 -2124
rect 1752 -2125 1753 -2124
rect 114 -2127 115 -2126
rect 366 -2127 367 -2126
rect 611 -2127 612 -2126
rect 625 -2127 626 -2126
rect 628 -2127 629 -2126
rect 870 -2127 871 -2126
rect 894 -2127 895 -2126
rect 1276 -2127 1277 -2126
rect 1486 -2127 1487 -2126
rect 1549 -2127 1550 -2126
rect 1689 -2127 1690 -2126
rect 1787 -2127 1788 -2126
rect 282 -2129 283 -2128
rect 359 -2129 360 -2128
rect 625 -2129 626 -2128
rect 800 -2129 801 -2128
rect 1080 -2129 1081 -2128
rect 1780 -2129 1781 -2128
rect 1787 -2129 1788 -2128
rect 1871 -2129 1872 -2128
rect 100 -2131 101 -2130
rect 282 -2131 283 -2130
rect 289 -2131 290 -2130
rect 866 -2131 867 -2130
rect 1255 -2131 1256 -2130
rect 1360 -2131 1361 -2130
rect 1549 -2131 1550 -2130
rect 1556 -2131 1557 -2130
rect 1780 -2131 1781 -2130
rect 1864 -2131 1865 -2130
rect 1871 -2131 1872 -2130
rect 1955 -2131 1956 -2130
rect 100 -2133 101 -2132
rect 1451 -2133 1452 -2132
rect 1556 -2133 1557 -2132
rect 1647 -2133 1648 -2132
rect 296 -2135 297 -2134
rect 569 -2135 570 -2134
rect 639 -2135 640 -2134
rect 856 -2135 857 -2134
rect 1269 -2135 1270 -2134
rect 1297 -2135 1298 -2134
rect 1451 -2135 1452 -2134
rect 1598 -2135 1599 -2134
rect 1612 -2135 1613 -2134
rect 1647 -2135 1648 -2134
rect 254 -2137 255 -2136
rect 296 -2137 297 -2136
rect 317 -2137 318 -2136
rect 856 -2137 857 -2136
rect 1269 -2137 1270 -2136
rect 1332 -2137 1333 -2136
rect 82 -2139 83 -2138
rect 254 -2139 255 -2138
rect 317 -2139 318 -2138
rect 331 -2139 332 -2138
rect 345 -2139 346 -2138
rect 443 -2139 444 -2138
rect 646 -2139 647 -2138
rect 1094 -2139 1095 -2138
rect 1293 -2139 1294 -2138
rect 1612 -2139 1613 -2138
rect 331 -2141 332 -2140
rect 478 -2141 479 -2140
rect 653 -2141 654 -2140
rect 674 -2141 675 -2140
rect 737 -2141 738 -2140
rect 793 -2141 794 -2140
rect 800 -2141 801 -2140
rect 821 -2141 822 -2140
rect 940 -2141 941 -2140
rect 1094 -2141 1095 -2140
rect 1332 -2141 1333 -2140
rect 1444 -2141 1445 -2140
rect 443 -2143 444 -2142
rect 765 -2143 766 -2142
rect 793 -2143 794 -2142
rect 898 -2143 899 -2142
rect 1444 -2143 1445 -2142
rect 1535 -2143 1536 -2142
rect 275 -2145 276 -2144
rect 898 -2145 899 -2144
rect 1430 -2145 1431 -2144
rect 1535 -2145 1536 -2144
rect 275 -2147 276 -2146
rect 828 -2147 829 -2146
rect 1430 -2147 1431 -2146
rect 1528 -2147 1529 -2146
rect 453 -2149 454 -2148
rect 828 -2149 829 -2148
rect 1528 -2149 1529 -2148
rect 1640 -2149 1641 -2148
rect 457 -2151 458 -2150
rect 478 -2151 479 -2150
rect 667 -2151 668 -2150
rect 940 -2151 941 -2150
rect 1626 -2151 1627 -2150
rect 1640 -2151 1641 -2150
rect 457 -2153 458 -2152
rect 660 -2153 661 -2152
rect 667 -2153 668 -2152
rect 688 -2153 689 -2152
rect 754 -2153 755 -2152
rect 1864 -2153 1865 -2152
rect 555 -2155 556 -2154
rect 688 -2155 689 -2154
rect 765 -2155 766 -2154
rect 1395 -2155 1396 -2154
rect 1563 -2155 1564 -2154
rect 1626 -2155 1627 -2154
rect 555 -2157 556 -2156
rect 632 -2157 633 -2156
rect 660 -2157 661 -2156
rect 1090 -2157 1091 -2156
rect 1563 -2157 1564 -2156
rect 1654 -2157 1655 -2156
rect 404 -2159 405 -2158
rect 1654 -2159 1655 -2158
rect 429 -2161 430 -2160
rect 632 -2161 633 -2160
rect 674 -2161 675 -2160
rect 681 -2161 682 -2160
rect 821 -2161 822 -2160
rect 835 -2161 836 -2160
rect 429 -2163 430 -2162
rect 436 -2163 437 -2162
rect 534 -2163 535 -2162
rect 835 -2163 836 -2162
rect 534 -2165 535 -2164
rect 880 -2165 881 -2164
rect 681 -2167 682 -2166
rect 1083 -2167 1084 -2166
rect 880 -2169 881 -2168
rect 1150 -2169 1151 -2168
rect 1150 -2171 1151 -2170
rect 1227 -2171 1228 -2170
rect 1227 -2173 1228 -2172
rect 1318 -2173 1319 -2172
rect 912 -2175 913 -2174
rect 1318 -2175 1319 -2174
rect 121 -2177 122 -2176
rect 912 -2177 913 -2176
rect 72 -2179 73 -2178
rect 121 -2179 122 -2178
rect 72 -2181 73 -2180
rect 464 -2181 465 -2180
rect 58 -2183 59 -2182
rect 464 -2183 465 -2182
rect 58 -2185 59 -2184
rect 387 -2185 388 -2184
rect 2 -2196 3 -2195
rect 40 -2196 41 -2195
rect 58 -2196 59 -2195
rect 215 -2196 216 -2195
rect 222 -2196 223 -2195
rect 1139 -2196 1140 -2195
rect 1178 -2196 1179 -2195
rect 1451 -2196 1452 -2195
rect 1454 -2196 1455 -2195
rect 1808 -2196 1809 -2195
rect 12 -2198 13 -2197
rect 16 -2198 17 -2197
rect 33 -2198 34 -2197
rect 520 -2198 521 -2197
rect 527 -2198 528 -2197
rect 761 -2198 762 -2197
rect 817 -2198 818 -2197
rect 1038 -2198 1039 -2197
rect 1055 -2198 1056 -2197
rect 1318 -2198 1319 -2197
rect 1360 -2198 1361 -2197
rect 1486 -2198 1487 -2197
rect 1713 -2198 1714 -2197
rect 1724 -2198 1725 -2197
rect 1727 -2198 1728 -2197
rect 1906 -2198 1907 -2197
rect 16 -2200 17 -2199
rect 303 -2200 304 -2199
rect 317 -2200 318 -2199
rect 341 -2200 342 -2199
rect 352 -2200 353 -2199
rect 625 -2200 626 -2199
rect 646 -2200 647 -2199
rect 891 -2200 892 -2199
rect 950 -2200 951 -2199
rect 1878 -2200 1879 -2199
rect 37 -2202 38 -2201
rect 849 -2202 850 -2201
rect 877 -2202 878 -2201
rect 1297 -2202 1298 -2201
rect 1318 -2202 1319 -2201
rect 1458 -2202 1459 -2201
rect 1475 -2202 1476 -2201
rect 1759 -2202 1760 -2201
rect 23 -2204 24 -2203
rect 37 -2204 38 -2203
rect 44 -2204 45 -2203
rect 58 -2204 59 -2203
rect 68 -2204 69 -2203
rect 296 -2204 297 -2203
rect 303 -2204 304 -2203
rect 562 -2204 563 -2203
rect 572 -2204 573 -2203
rect 884 -2204 885 -2203
rect 891 -2204 892 -2203
rect 1304 -2204 1305 -2203
rect 1395 -2204 1396 -2203
rect 1787 -2204 1788 -2203
rect 23 -2206 24 -2205
rect 191 -2206 192 -2205
rect 254 -2206 255 -2205
rect 1083 -2206 1084 -2205
rect 1108 -2206 1109 -2205
rect 1262 -2206 1263 -2205
rect 1276 -2206 1277 -2205
rect 1286 -2206 1287 -2205
rect 1304 -2206 1305 -2205
rect 1822 -2206 1823 -2205
rect 44 -2208 45 -2207
rect 128 -2208 129 -2207
rect 163 -2208 164 -2207
rect 1125 -2208 1126 -2207
rect 1136 -2208 1137 -2207
rect 1220 -2208 1221 -2207
rect 1255 -2208 1256 -2207
rect 1262 -2208 1263 -2207
rect 1276 -2208 1277 -2207
rect 1325 -2208 1326 -2207
rect 1395 -2208 1396 -2207
rect 1605 -2208 1606 -2207
rect 1787 -2208 1788 -2207
rect 1794 -2208 1795 -2207
rect 1822 -2208 1823 -2207
rect 1892 -2208 1893 -2207
rect 107 -2210 108 -2209
rect 275 -2210 276 -2209
rect 282 -2210 283 -2209
rect 338 -2210 339 -2209
rect 352 -2210 353 -2209
rect 597 -2210 598 -2209
rect 670 -2210 671 -2209
rect 1885 -2210 1886 -2209
rect 107 -2212 108 -2211
rect 814 -2212 815 -2211
rect 877 -2212 878 -2211
rect 919 -2212 920 -2211
rect 954 -2212 955 -2211
rect 1297 -2212 1298 -2211
rect 1325 -2212 1326 -2211
rect 1444 -2212 1445 -2211
rect 1458 -2212 1459 -2211
rect 1479 -2212 1480 -2211
rect 1605 -2212 1606 -2211
rect 1647 -2212 1648 -2211
rect 1794 -2212 1795 -2211
rect 1899 -2212 1900 -2211
rect 110 -2214 111 -2213
rect 324 -2214 325 -2213
rect 387 -2214 388 -2213
rect 478 -2214 479 -2213
rect 520 -2214 521 -2213
rect 716 -2214 717 -2213
rect 786 -2214 787 -2213
rect 1486 -2214 1487 -2213
rect 1640 -2214 1641 -2213
rect 1647 -2214 1648 -2213
rect 117 -2216 118 -2215
rect 149 -2216 150 -2215
rect 163 -2216 164 -2215
rect 247 -2216 248 -2215
rect 254 -2216 255 -2215
rect 331 -2216 332 -2215
rect 408 -2216 409 -2215
rect 478 -2216 479 -2215
rect 527 -2216 528 -2215
rect 611 -2216 612 -2215
rect 737 -2216 738 -2215
rect 786 -2216 787 -2215
rect 793 -2216 794 -2215
rect 849 -2216 850 -2215
rect 880 -2216 881 -2215
rect 1500 -2216 1501 -2215
rect 1640 -2216 1641 -2215
rect 1745 -2216 1746 -2215
rect 128 -2218 129 -2217
rect 135 -2218 136 -2217
rect 170 -2218 171 -2217
rect 387 -2218 388 -2217
rect 408 -2218 409 -2217
rect 485 -2218 486 -2217
rect 544 -2218 545 -2217
rect 912 -2218 913 -2217
rect 919 -2218 920 -2217
rect 947 -2218 948 -2217
rect 968 -2218 969 -2217
rect 1577 -2218 1578 -2217
rect 1745 -2218 1746 -2217
rect 1913 -2218 1914 -2217
rect 135 -2220 136 -2219
rect 184 -2220 185 -2219
rect 191 -2220 192 -2219
rect 975 -2220 976 -2219
rect 999 -2220 1000 -2219
rect 1535 -2220 1536 -2219
rect 170 -2222 171 -2221
rect 268 -2222 269 -2221
rect 289 -2222 290 -2221
rect 324 -2222 325 -2221
rect 331 -2222 332 -2221
rect 464 -2222 465 -2221
rect 471 -2222 472 -2221
rect 1080 -2222 1081 -2221
rect 1108 -2222 1109 -2221
rect 1283 -2222 1284 -2221
rect 1353 -2222 1354 -2221
rect 1577 -2222 1578 -2221
rect 79 -2224 80 -2223
rect 289 -2224 290 -2223
rect 296 -2224 297 -2223
rect 443 -2224 444 -2223
rect 457 -2224 458 -2223
rect 509 -2224 510 -2223
rect 562 -2224 563 -2223
rect 723 -2224 724 -2223
rect 737 -2224 738 -2223
rect 863 -2224 864 -2223
rect 912 -2224 913 -2223
rect 926 -2224 927 -2223
rect 968 -2224 969 -2223
rect 1003 -2224 1004 -2223
rect 1038 -2224 1039 -2223
rect 1101 -2224 1102 -2223
rect 1111 -2224 1112 -2223
rect 1626 -2224 1627 -2223
rect 51 -2226 52 -2225
rect 457 -2226 458 -2225
rect 485 -2226 486 -2225
rect 492 -2226 493 -2225
rect 569 -2226 570 -2225
rect 716 -2226 717 -2225
rect 796 -2226 797 -2225
rect 954 -2226 955 -2225
rect 971 -2226 972 -2225
rect 1094 -2226 1095 -2225
rect 1101 -2226 1102 -2225
rect 1150 -2226 1151 -2225
rect 1178 -2226 1179 -2225
rect 1339 -2226 1340 -2225
rect 1353 -2226 1354 -2225
rect 1416 -2226 1417 -2225
rect 1444 -2226 1445 -2225
rect 1493 -2226 1494 -2225
rect 1500 -2226 1501 -2225
rect 1591 -2226 1592 -2225
rect 1626 -2226 1627 -2225
rect 1738 -2226 1739 -2225
rect 30 -2228 31 -2227
rect 51 -2228 52 -2227
rect 79 -2228 80 -2227
rect 100 -2228 101 -2227
rect 142 -2228 143 -2227
rect 268 -2228 269 -2227
rect 380 -2228 381 -2227
rect 569 -2228 570 -2227
rect 590 -2228 591 -2227
rect 1241 -2228 1242 -2227
rect 1279 -2228 1280 -2227
rect 1549 -2228 1550 -2227
rect 1591 -2228 1592 -2227
rect 1675 -2228 1676 -2227
rect 1696 -2228 1697 -2227
rect 1738 -2228 1739 -2227
rect 30 -2230 31 -2229
rect 1024 -2230 1025 -2229
rect 1031 -2230 1032 -2229
rect 1339 -2230 1340 -2229
rect 1398 -2230 1399 -2229
rect 1871 -2230 1872 -2229
rect 65 -2232 66 -2231
rect 100 -2232 101 -2231
rect 177 -2232 178 -2231
rect 471 -2232 472 -2231
rect 576 -2232 577 -2231
rect 590 -2232 591 -2231
rect 597 -2232 598 -2231
rect 632 -2232 633 -2231
rect 639 -2232 640 -2231
rect 793 -2232 794 -2231
rect 926 -2232 927 -2231
rect 961 -2232 962 -2231
rect 989 -2232 990 -2231
rect 1003 -2232 1004 -2231
rect 1010 -2232 1011 -2231
rect 1031 -2232 1032 -2231
rect 1052 -2232 1053 -2231
rect 1360 -2232 1361 -2231
rect 1402 -2232 1403 -2231
rect 1619 -2232 1620 -2231
rect 1675 -2232 1676 -2231
rect 1829 -2232 1830 -2231
rect 86 -2234 87 -2233
rect 177 -2234 178 -2233
rect 184 -2234 185 -2233
rect 219 -2234 220 -2233
rect 226 -2234 227 -2233
rect 247 -2234 248 -2233
rect 261 -2234 262 -2233
rect 317 -2234 318 -2233
rect 415 -2234 416 -2233
rect 492 -2234 493 -2233
rect 506 -2234 507 -2233
rect 961 -2234 962 -2233
rect 989 -2234 990 -2233
rect 1017 -2234 1018 -2233
rect 1024 -2234 1025 -2233
rect 1059 -2234 1060 -2233
rect 1066 -2234 1067 -2233
rect 1185 -2234 1186 -2233
rect 1188 -2234 1189 -2233
rect 1332 -2234 1333 -2233
rect 1402 -2234 1403 -2233
rect 1430 -2234 1431 -2233
rect 1479 -2234 1480 -2233
rect 1563 -2234 1564 -2233
rect 1619 -2234 1620 -2233
rect 1703 -2234 1704 -2233
rect 1829 -2234 1830 -2233
rect 1850 -2234 1851 -2233
rect 86 -2236 87 -2235
rect 394 -2236 395 -2235
rect 415 -2236 416 -2235
rect 467 -2236 468 -2235
rect 506 -2236 507 -2235
rect 772 -2236 773 -2235
rect 800 -2236 801 -2235
rect 1059 -2236 1060 -2235
rect 1087 -2236 1088 -2235
rect 1150 -2236 1151 -2235
rect 1192 -2236 1193 -2235
rect 1241 -2236 1242 -2235
rect 1283 -2236 1284 -2235
rect 1388 -2236 1389 -2235
rect 1430 -2236 1431 -2235
rect 1514 -2236 1515 -2235
rect 1535 -2236 1536 -2235
rect 1689 -2236 1690 -2235
rect 1696 -2236 1697 -2235
rect 1815 -2236 1816 -2235
rect 173 -2238 174 -2237
rect 772 -2238 773 -2237
rect 1010 -2238 1011 -2237
rect 1164 -2238 1165 -2237
rect 1192 -2238 1193 -2237
rect 1290 -2238 1291 -2237
rect 1332 -2238 1333 -2237
rect 1423 -2238 1424 -2237
rect 1493 -2238 1494 -2237
rect 1542 -2238 1543 -2237
rect 1549 -2238 1550 -2237
rect 1773 -2238 1774 -2237
rect 93 -2240 94 -2239
rect 1423 -2240 1424 -2239
rect 1514 -2240 1515 -2239
rect 1570 -2240 1571 -2239
rect 1689 -2240 1690 -2239
rect 1843 -2240 1844 -2239
rect 93 -2242 94 -2241
rect 124 -2242 125 -2241
rect 198 -2242 199 -2241
rect 282 -2242 283 -2241
rect 394 -2242 395 -2241
rect 541 -2242 542 -2241
rect 576 -2242 577 -2241
rect 947 -2242 948 -2241
rect 975 -2242 976 -2241
rect 1290 -2242 1291 -2241
rect 1542 -2242 1543 -2241
rect 1584 -2242 1585 -2241
rect 1703 -2242 1704 -2241
rect 1857 -2242 1858 -2241
rect 198 -2244 199 -2243
rect 401 -2244 402 -2243
rect 429 -2244 430 -2243
rect 632 -2244 633 -2243
rect 649 -2244 650 -2243
rect 1416 -2244 1417 -2243
rect 1563 -2244 1564 -2243
rect 1633 -2244 1634 -2243
rect 1773 -2244 1774 -2243
rect 1801 -2244 1802 -2243
rect 205 -2246 206 -2245
rect 275 -2246 276 -2245
rect 345 -2246 346 -2245
rect 401 -2246 402 -2245
rect 429 -2246 430 -2245
rect 842 -2246 843 -2245
rect 1052 -2246 1053 -2245
rect 1346 -2246 1347 -2245
rect 1570 -2246 1571 -2245
rect 1654 -2246 1655 -2245
rect 72 -2248 73 -2247
rect 345 -2248 346 -2247
rect 366 -2248 367 -2247
rect 541 -2248 542 -2247
rect 611 -2248 612 -2247
rect 653 -2248 654 -2247
rect 656 -2248 657 -2247
rect 1094 -2248 1095 -2247
rect 1122 -2248 1123 -2247
rect 1160 -2248 1161 -2247
rect 1164 -2248 1165 -2247
rect 1234 -2248 1235 -2247
rect 1346 -2248 1347 -2247
rect 1437 -2248 1438 -2247
rect 1584 -2248 1585 -2247
rect 1661 -2248 1662 -2247
rect 72 -2250 73 -2249
rect 121 -2250 122 -2249
rect 156 -2250 157 -2249
rect 205 -2250 206 -2249
rect 208 -2250 209 -2249
rect 723 -2250 724 -2249
rect 744 -2250 745 -2249
rect 1234 -2250 1235 -2249
rect 1286 -2250 1287 -2249
rect 1661 -2250 1662 -2249
rect 121 -2252 122 -2251
rect 142 -2252 143 -2251
rect 156 -2252 157 -2251
rect 1668 -2252 1669 -2251
rect 212 -2254 213 -2253
rect 380 -2254 381 -2253
rect 443 -2254 444 -2253
rect 450 -2254 451 -2253
rect 618 -2254 619 -2253
rect 800 -2254 801 -2253
rect 842 -2254 843 -2253
rect 905 -2254 906 -2253
rect 1087 -2254 1088 -2253
rect 1115 -2254 1116 -2253
rect 1122 -2254 1123 -2253
rect 1710 -2254 1711 -2253
rect 212 -2256 213 -2255
rect 758 -2256 759 -2255
rect 765 -2256 766 -2255
rect 1017 -2256 1018 -2255
rect 1115 -2256 1116 -2255
rect 1129 -2256 1130 -2255
rect 1213 -2256 1214 -2255
rect 1255 -2256 1256 -2255
rect 1293 -2256 1294 -2255
rect 1668 -2256 1669 -2255
rect 1710 -2256 1711 -2255
rect 1759 -2256 1760 -2255
rect 219 -2258 220 -2257
rect 436 -2258 437 -2257
rect 450 -2258 451 -2257
rect 499 -2258 500 -2257
rect 618 -2258 619 -2257
rect 933 -2258 934 -2257
rect 1129 -2258 1130 -2257
rect 1206 -2258 1207 -2257
rect 1220 -2258 1221 -2257
rect 1409 -2258 1410 -2257
rect 1437 -2258 1438 -2257
rect 1521 -2258 1522 -2257
rect 1633 -2258 1634 -2257
rect 1836 -2258 1837 -2257
rect 226 -2260 227 -2259
rect 240 -2260 241 -2259
rect 261 -2260 262 -2259
rect 359 -2260 360 -2259
rect 366 -2260 367 -2259
rect 555 -2260 556 -2259
rect 628 -2260 629 -2259
rect 1206 -2260 1207 -2259
rect 1409 -2260 1410 -2259
rect 1556 -2260 1557 -2259
rect 236 -2262 237 -2261
rect 1654 -2262 1655 -2261
rect 240 -2264 241 -2263
rect 1752 -2264 1753 -2263
rect 310 -2266 311 -2265
rect 359 -2266 360 -2265
rect 422 -2266 423 -2265
rect 933 -2266 934 -2265
rect 1521 -2266 1522 -2265
rect 1682 -2266 1683 -2265
rect 1752 -2266 1753 -2265
rect 1864 -2266 1865 -2265
rect 159 -2268 160 -2267
rect 310 -2268 311 -2267
rect 373 -2268 374 -2267
rect 422 -2268 423 -2267
rect 436 -2268 437 -2267
rect 870 -2268 871 -2267
rect 905 -2268 906 -2267
rect 940 -2268 941 -2267
rect 1556 -2268 1557 -2267
rect 1612 -2268 1613 -2267
rect 1682 -2268 1683 -2267
rect 1780 -2268 1781 -2267
rect 373 -2270 374 -2269
rect 548 -2270 549 -2269
rect 555 -2270 556 -2269
rect 681 -2270 682 -2269
rect 709 -2270 710 -2269
rect 863 -2270 864 -2269
rect 870 -2270 871 -2269
rect 898 -2270 899 -2269
rect 940 -2270 941 -2269
rect 982 -2270 983 -2269
rect 1612 -2270 1613 -2269
rect 1766 -2270 1767 -2269
rect 390 -2272 391 -2271
rect 1780 -2272 1781 -2271
rect 499 -2274 500 -2273
rect 534 -2274 535 -2273
rect 548 -2274 549 -2273
rect 604 -2274 605 -2273
rect 639 -2274 640 -2273
rect 758 -2274 759 -2273
rect 765 -2274 766 -2273
rect 856 -2274 857 -2273
rect 898 -2274 899 -2273
rect 1157 -2274 1158 -2273
rect 1731 -2274 1732 -2273
rect 1766 -2274 1767 -2273
rect 89 -2276 90 -2275
rect 534 -2276 535 -2275
rect 604 -2276 605 -2275
rect 674 -2276 675 -2275
rect 677 -2276 678 -2275
rect 1388 -2276 1389 -2275
rect 1472 -2276 1473 -2275
rect 1731 -2276 1732 -2275
rect 653 -2278 654 -2277
rect 1045 -2278 1046 -2277
rect 1157 -2278 1158 -2277
rect 1227 -2278 1228 -2277
rect 660 -2280 661 -2279
rect 681 -2280 682 -2279
rect 702 -2280 703 -2279
rect 709 -2280 710 -2279
rect 744 -2280 745 -2279
rect 807 -2280 808 -2279
rect 821 -2280 822 -2279
rect 856 -2280 857 -2279
rect 982 -2280 983 -2279
rect 996 -2280 997 -2279
rect 1185 -2280 1186 -2279
rect 1472 -2280 1473 -2279
rect 9 -2282 10 -2281
rect 996 -2282 997 -2281
rect 1227 -2282 1228 -2281
rect 1311 -2282 1312 -2281
rect 660 -2284 661 -2283
rect 667 -2284 668 -2283
rect 674 -2284 675 -2283
rect 1073 -2284 1074 -2283
rect 1311 -2284 1312 -2283
rect 1381 -2284 1382 -2283
rect 688 -2286 689 -2285
rect 702 -2286 703 -2285
rect 751 -2286 752 -2285
rect 1045 -2286 1046 -2285
rect 1073 -2286 1074 -2285
rect 1143 -2286 1144 -2285
rect 583 -2288 584 -2287
rect 688 -2288 689 -2287
rect 751 -2288 752 -2287
rect 824 -2288 825 -2287
rect 835 -2288 836 -2287
rect 1381 -2288 1382 -2287
rect 513 -2290 514 -2289
rect 583 -2290 584 -2289
rect 807 -2290 808 -2289
rect 828 -2290 829 -2289
rect 835 -2290 836 -2289
rect 887 -2290 888 -2289
rect 978 -2290 979 -2289
rect 1143 -2290 1144 -2289
rect 65 -2292 66 -2291
rect 513 -2292 514 -2291
rect 821 -2292 822 -2291
rect 1213 -2292 1214 -2291
rect 828 -2294 829 -2293
rect 1199 -2294 1200 -2293
rect 1199 -2296 1200 -2295
rect 1374 -2296 1375 -2295
rect 1374 -2298 1375 -2297
rect 1465 -2298 1466 -2297
rect 1465 -2300 1466 -2299
rect 1528 -2300 1529 -2299
rect 1507 -2302 1508 -2301
rect 1528 -2302 1529 -2301
rect 1507 -2304 1508 -2303
rect 1598 -2304 1599 -2303
rect 1069 -2306 1070 -2305
rect 1598 -2306 1599 -2305
rect 1069 -2308 1070 -2307
rect 1171 -2308 1172 -2307
rect 1171 -2310 1172 -2309
rect 1269 -2310 1270 -2309
rect 1269 -2312 1270 -2311
rect 1367 -2312 1368 -2311
rect 149 -2314 150 -2313
rect 1367 -2314 1368 -2313
rect 9 -2325 10 -2324
rect 170 -2325 171 -2324
rect 177 -2325 178 -2324
rect 1727 -2325 1728 -2324
rect 1731 -2325 1732 -2324
rect 1745 -2325 1746 -2324
rect 1748 -2325 1749 -2324
rect 1822 -2325 1823 -2324
rect 9 -2327 10 -2326
rect 492 -2327 493 -2326
rect 499 -2327 500 -2326
rect 817 -2327 818 -2326
rect 821 -2327 822 -2326
rect 1206 -2327 1207 -2326
rect 1216 -2327 1217 -2326
rect 1451 -2327 1452 -2326
rect 1577 -2327 1578 -2326
rect 1731 -2327 1732 -2326
rect 1755 -2327 1756 -2326
rect 1766 -2327 1767 -2326
rect 1780 -2327 1781 -2326
rect 1801 -2327 1802 -2326
rect 16 -2329 17 -2328
rect 618 -2329 619 -2328
rect 625 -2329 626 -2328
rect 1052 -2329 1053 -2328
rect 1069 -2329 1070 -2328
rect 1255 -2329 1256 -2328
rect 1276 -2329 1277 -2328
rect 1293 -2329 1294 -2328
rect 1307 -2329 1308 -2328
rect 1458 -2329 1459 -2328
rect 1738 -2329 1739 -2328
rect 1766 -2329 1767 -2328
rect 1787 -2329 1788 -2328
rect 1808 -2329 1809 -2328
rect 16 -2331 17 -2330
rect 432 -2331 433 -2330
rect 439 -2331 440 -2330
rect 457 -2331 458 -2330
rect 460 -2331 461 -2330
rect 590 -2331 591 -2330
rect 625 -2331 626 -2330
rect 905 -2331 906 -2330
rect 947 -2331 948 -2330
rect 1038 -2331 1039 -2330
rect 1052 -2331 1053 -2330
rect 1486 -2331 1487 -2330
rect 1675 -2331 1676 -2330
rect 1738 -2331 1739 -2330
rect 1759 -2331 1760 -2330
rect 1780 -2331 1781 -2330
rect 1787 -2331 1788 -2330
rect 1794 -2331 1795 -2330
rect 1797 -2331 1798 -2330
rect 1829 -2331 1830 -2330
rect 30 -2333 31 -2332
rect 114 -2333 115 -2332
rect 142 -2333 143 -2332
rect 212 -2333 213 -2332
rect 233 -2333 234 -2332
rect 387 -2333 388 -2332
rect 408 -2333 409 -2332
rect 733 -2333 734 -2332
rect 793 -2333 794 -2332
rect 807 -2333 808 -2332
rect 814 -2333 815 -2332
rect 975 -2333 976 -2332
rect 996 -2333 997 -2332
rect 1577 -2333 1578 -2332
rect 1619 -2333 1620 -2332
rect 1675 -2333 1676 -2332
rect 1759 -2333 1760 -2332
rect 1773 -2333 1774 -2332
rect 30 -2335 31 -2334
rect 149 -2335 150 -2334
rect 159 -2335 160 -2334
rect 324 -2335 325 -2334
rect 352 -2335 353 -2334
rect 667 -2335 668 -2334
rect 698 -2335 699 -2334
rect 842 -2335 843 -2334
rect 863 -2335 864 -2334
rect 975 -2335 976 -2334
rect 1020 -2335 1021 -2334
rect 1241 -2335 1242 -2334
rect 1248 -2335 1249 -2334
rect 1276 -2335 1277 -2334
rect 1290 -2335 1291 -2334
rect 1549 -2335 1550 -2334
rect 1619 -2335 1620 -2334
rect 1689 -2335 1690 -2334
rect 1717 -2335 1718 -2334
rect 1773 -2335 1774 -2334
rect 44 -2337 45 -2336
rect 236 -2337 237 -2336
rect 282 -2337 283 -2336
rect 464 -2337 465 -2336
rect 471 -2337 472 -2336
rect 618 -2337 619 -2336
rect 646 -2337 647 -2336
rect 842 -2337 843 -2336
rect 884 -2337 885 -2336
rect 1003 -2337 1004 -2336
rect 1017 -2337 1018 -2336
rect 1241 -2337 1242 -2336
rect 1321 -2337 1322 -2336
rect 1325 -2337 1326 -2336
rect 1342 -2337 1343 -2336
rect 1710 -2337 1711 -2336
rect 44 -2339 45 -2338
rect 226 -2339 227 -2338
rect 303 -2339 304 -2338
rect 530 -2339 531 -2338
rect 544 -2339 545 -2338
rect 639 -2339 640 -2338
rect 646 -2339 647 -2338
rect 887 -2339 888 -2338
rect 905 -2339 906 -2338
rect 912 -2339 913 -2338
rect 947 -2339 948 -2338
rect 961 -2339 962 -2338
rect 1038 -2339 1039 -2338
rect 1059 -2339 1060 -2338
rect 1066 -2339 1067 -2338
rect 1290 -2339 1291 -2338
rect 1370 -2339 1371 -2338
rect 1395 -2339 1396 -2338
rect 1423 -2339 1424 -2338
rect 1451 -2339 1452 -2338
rect 1486 -2339 1487 -2338
rect 1493 -2339 1494 -2338
rect 1542 -2339 1543 -2338
rect 1549 -2339 1550 -2338
rect 1633 -2339 1634 -2338
rect 1689 -2339 1690 -2338
rect 51 -2341 52 -2340
rect 1003 -2341 1004 -2340
rect 1010 -2341 1011 -2340
rect 1059 -2341 1060 -2340
rect 1066 -2341 1067 -2340
rect 1080 -2341 1081 -2340
rect 1115 -2341 1116 -2340
rect 1514 -2341 1515 -2340
rect 1521 -2341 1522 -2340
rect 1633 -2341 1634 -2340
rect 37 -2343 38 -2342
rect 1080 -2343 1081 -2342
rect 1115 -2343 1116 -2342
rect 1178 -2343 1179 -2342
rect 1188 -2343 1189 -2342
rect 1682 -2343 1683 -2342
rect 37 -2345 38 -2344
rect 240 -2345 241 -2344
rect 310 -2345 311 -2344
rect 457 -2345 458 -2344
rect 467 -2345 468 -2344
rect 1423 -2345 1424 -2344
rect 1430 -2345 1431 -2344
rect 1458 -2345 1459 -2344
rect 1465 -2345 1466 -2344
rect 1493 -2345 1494 -2344
rect 1521 -2345 1522 -2344
rect 1556 -2345 1557 -2344
rect 1640 -2345 1641 -2344
rect 1682 -2345 1683 -2344
rect 51 -2347 52 -2346
rect 243 -2347 244 -2346
rect 310 -2347 311 -2346
rect 446 -2347 447 -2346
rect 450 -2347 451 -2346
rect 464 -2347 465 -2346
rect 478 -2347 479 -2346
rect 492 -2347 493 -2346
rect 534 -2347 535 -2346
rect 961 -2347 962 -2346
rect 1010 -2347 1011 -2346
rect 1094 -2347 1095 -2346
rect 1157 -2347 1158 -2346
rect 1160 -2347 1161 -2346
rect 1171 -2347 1172 -2346
rect 1206 -2347 1207 -2346
rect 1213 -2347 1214 -2346
rect 1255 -2347 1256 -2346
rect 1283 -2347 1284 -2346
rect 1325 -2347 1326 -2346
rect 1360 -2347 1361 -2346
rect 1395 -2347 1396 -2346
rect 1437 -2347 1438 -2346
rect 1465 -2347 1466 -2346
rect 1479 -2347 1480 -2346
rect 1514 -2347 1515 -2346
rect 1640 -2347 1641 -2346
rect 1703 -2347 1704 -2346
rect 58 -2349 59 -2348
rect 82 -2349 83 -2348
rect 86 -2349 87 -2348
rect 677 -2349 678 -2348
rect 723 -2349 724 -2348
rect 996 -2349 997 -2348
rect 1017 -2349 1018 -2348
rect 1171 -2349 1172 -2348
rect 1227 -2349 1228 -2348
rect 1248 -2349 1249 -2348
rect 1339 -2349 1340 -2348
rect 1360 -2349 1361 -2348
rect 1416 -2349 1417 -2348
rect 1437 -2349 1438 -2348
rect 1444 -2349 1445 -2348
rect 1479 -2349 1480 -2348
rect 1500 -2349 1501 -2348
rect 1556 -2349 1557 -2348
rect 1661 -2349 1662 -2348
rect 1703 -2349 1704 -2348
rect 58 -2351 59 -2350
rect 219 -2351 220 -2350
rect 296 -2351 297 -2350
rect 677 -2351 678 -2350
rect 772 -2351 773 -2350
rect 1178 -2351 1179 -2350
rect 1227 -2351 1228 -2350
rect 1794 -2351 1795 -2350
rect 65 -2353 66 -2352
rect 485 -2353 486 -2352
rect 513 -2353 514 -2352
rect 534 -2353 535 -2352
rect 562 -2353 563 -2352
rect 824 -2353 825 -2352
rect 831 -2353 832 -2352
rect 1542 -2353 1543 -2352
rect 1626 -2353 1627 -2352
rect 1661 -2353 1662 -2352
rect 72 -2355 73 -2354
rect 110 -2355 111 -2354
rect 114 -2355 115 -2354
rect 198 -2355 199 -2354
rect 205 -2355 206 -2354
rect 499 -2355 500 -2354
rect 541 -2355 542 -2354
rect 562 -2355 563 -2354
rect 583 -2355 584 -2354
rect 590 -2355 591 -2354
rect 604 -2355 605 -2354
rect 639 -2355 640 -2354
rect 667 -2355 668 -2354
rect 702 -2355 703 -2354
rect 772 -2355 773 -2354
rect 786 -2355 787 -2354
rect 856 -2355 857 -2354
rect 887 -2355 888 -2354
rect 912 -2355 913 -2354
rect 926 -2355 927 -2354
rect 1055 -2355 1056 -2354
rect 1283 -2355 1284 -2354
rect 1332 -2355 1333 -2354
rect 1444 -2355 1445 -2354
rect 1591 -2355 1592 -2354
rect 1626 -2355 1627 -2354
rect 72 -2357 73 -2356
rect 100 -2357 101 -2356
rect 107 -2357 108 -2356
rect 408 -2357 409 -2356
rect 415 -2357 416 -2356
rect 471 -2357 472 -2356
rect 478 -2357 479 -2356
rect 681 -2357 682 -2356
rect 786 -2357 787 -2356
rect 807 -2357 808 -2356
rect 856 -2357 857 -2356
rect 870 -2357 871 -2356
rect 926 -2357 927 -2356
rect 1269 -2357 1270 -2356
rect 1339 -2357 1340 -2356
rect 1647 -2357 1648 -2356
rect 79 -2359 80 -2358
rect 226 -2359 227 -2358
rect 289 -2359 290 -2358
rect 296 -2359 297 -2358
rect 324 -2359 325 -2358
rect 527 -2359 528 -2358
rect 541 -2359 542 -2358
rect 688 -2359 689 -2358
rect 863 -2359 864 -2358
rect 884 -2359 885 -2358
rect 1094 -2359 1095 -2358
rect 1164 -2359 1165 -2358
rect 1199 -2359 1200 -2358
rect 1332 -2359 1333 -2358
rect 1388 -2359 1389 -2358
rect 1416 -2359 1417 -2358
rect 1528 -2359 1529 -2358
rect 1591 -2359 1592 -2358
rect 1605 -2359 1606 -2358
rect 1647 -2359 1648 -2358
rect 86 -2361 87 -2360
rect 93 -2361 94 -2360
rect 96 -2361 97 -2360
rect 1717 -2361 1718 -2360
rect 93 -2363 94 -2362
rect 124 -2363 125 -2362
rect 135 -2363 136 -2362
rect 303 -2363 304 -2362
rect 352 -2363 353 -2362
rect 1118 -2363 1119 -2362
rect 1150 -2363 1151 -2362
rect 1199 -2363 1200 -2362
rect 1269 -2363 1270 -2362
rect 1318 -2363 1319 -2362
rect 1388 -2363 1389 -2362
rect 1696 -2363 1697 -2362
rect 100 -2365 101 -2364
rect 163 -2365 164 -2364
rect 170 -2365 171 -2364
rect 422 -2365 423 -2364
rect 429 -2365 430 -2364
rect 723 -2365 724 -2364
rect 870 -2365 871 -2364
rect 877 -2365 878 -2364
rect 1150 -2365 1151 -2364
rect 1213 -2365 1214 -2364
rect 1563 -2365 1564 -2364
rect 1605 -2365 1606 -2364
rect 1654 -2365 1655 -2364
rect 1696 -2365 1697 -2364
rect 121 -2367 122 -2366
rect 513 -2367 514 -2366
rect 520 -2367 521 -2366
rect 688 -2367 689 -2366
rect 877 -2367 878 -2366
rect 940 -2367 941 -2366
rect 1157 -2367 1158 -2366
rect 1220 -2367 1221 -2366
rect 1507 -2367 1508 -2366
rect 1563 -2367 1564 -2366
rect 1598 -2367 1599 -2366
rect 1654 -2367 1655 -2366
rect 107 -2369 108 -2368
rect 940 -2369 941 -2368
rect 1083 -2369 1084 -2368
rect 1507 -2369 1508 -2368
rect 1598 -2369 1599 -2368
rect 1668 -2369 1669 -2368
rect 131 -2371 132 -2370
rect 135 -2371 136 -2370
rect 142 -2371 143 -2370
rect 999 -2371 1000 -2370
rect 1164 -2371 1165 -2370
rect 1612 -2371 1613 -2370
rect 149 -2373 150 -2372
rect 576 -2373 577 -2372
rect 583 -2373 584 -2372
rect 968 -2373 969 -2372
rect 1192 -2373 1193 -2372
rect 1220 -2373 1221 -2372
rect 1535 -2373 1536 -2372
rect 1668 -2373 1669 -2372
rect 156 -2375 157 -2374
rect 198 -2375 199 -2374
rect 212 -2375 213 -2374
rect 215 -2375 216 -2374
rect 219 -2375 220 -2374
rect 436 -2375 437 -2374
rect 450 -2375 451 -2374
rect 737 -2375 738 -2374
rect 968 -2375 969 -2374
rect 982 -2375 983 -2374
rect 1160 -2375 1161 -2374
rect 1192 -2375 1193 -2374
rect 1535 -2375 1536 -2374
rect 1570 -2375 1571 -2374
rect 1584 -2375 1585 -2374
rect 1612 -2375 1613 -2374
rect 156 -2377 157 -2376
rect 1185 -2377 1186 -2376
rect 1402 -2377 1403 -2376
rect 1584 -2377 1585 -2376
rect 163 -2379 164 -2378
rect 730 -2379 731 -2378
rect 737 -2379 738 -2378
rect 779 -2379 780 -2378
rect 891 -2379 892 -2378
rect 1185 -2379 1186 -2378
rect 1374 -2379 1375 -2378
rect 1402 -2379 1403 -2378
rect 1570 -2379 1571 -2378
rect 1752 -2379 1753 -2378
rect 177 -2381 178 -2380
rect 275 -2381 276 -2380
rect 366 -2381 367 -2380
rect 429 -2381 430 -2380
rect 436 -2381 437 -2380
rect 653 -2381 654 -2380
rect 681 -2381 682 -2380
rect 695 -2381 696 -2380
rect 730 -2381 731 -2380
rect 1500 -2381 1501 -2380
rect 184 -2383 185 -2382
rect 282 -2383 283 -2382
rect 366 -2383 367 -2382
rect 380 -2383 381 -2382
rect 387 -2383 388 -2382
rect 821 -2383 822 -2382
rect 891 -2383 892 -2382
rect 919 -2383 920 -2382
rect 982 -2383 983 -2382
rect 1031 -2383 1032 -2382
rect 1346 -2383 1347 -2382
rect 1374 -2383 1375 -2382
rect 184 -2385 185 -2384
rect 359 -2385 360 -2384
rect 390 -2385 391 -2384
rect 702 -2385 703 -2384
rect 828 -2385 829 -2384
rect 1346 -2385 1347 -2384
rect 191 -2387 192 -2386
rect 240 -2387 241 -2386
rect 261 -2387 262 -2386
rect 422 -2387 423 -2386
rect 485 -2387 486 -2386
rect 548 -2387 549 -2386
rect 572 -2387 573 -2386
rect 779 -2387 780 -2386
rect 828 -2387 829 -2386
rect 1724 -2387 1725 -2386
rect 23 -2389 24 -2388
rect 191 -2389 192 -2388
rect 205 -2389 206 -2388
rect 1752 -2389 1753 -2388
rect 261 -2391 262 -2390
rect 443 -2391 444 -2390
rect 520 -2391 521 -2390
rect 849 -2391 850 -2390
rect 919 -2391 920 -2390
rect 933 -2391 934 -2390
rect 1031 -2391 1032 -2390
rect 1045 -2391 1046 -2390
rect 275 -2393 276 -2392
rect 317 -2393 318 -2392
rect 338 -2393 339 -2392
rect 359 -2393 360 -2392
rect 394 -2393 395 -2392
rect 415 -2393 416 -2392
rect 527 -2393 528 -2392
rect 1430 -2393 1431 -2392
rect 289 -2395 290 -2394
rect 443 -2395 444 -2394
rect 548 -2395 549 -2394
rect 709 -2395 710 -2394
rect 800 -2395 801 -2394
rect 849 -2395 850 -2394
rect 933 -2395 934 -2394
rect 954 -2395 955 -2394
rect 1045 -2395 1046 -2394
rect 1304 -2395 1305 -2394
rect 317 -2397 318 -2396
rect 506 -2397 507 -2396
rect 569 -2397 570 -2396
rect 709 -2397 710 -2396
rect 765 -2397 766 -2396
rect 800 -2397 801 -2396
rect 835 -2397 836 -2396
rect 954 -2397 955 -2396
rect 1262 -2397 1263 -2396
rect 1304 -2397 1305 -2396
rect 268 -2399 269 -2398
rect 506 -2399 507 -2398
rect 555 -2399 556 -2398
rect 765 -2399 766 -2398
rect 835 -2399 836 -2398
rect 1167 -2399 1168 -2398
rect 268 -2401 269 -2400
rect 331 -2401 332 -2400
rect 338 -2401 339 -2400
rect 898 -2401 899 -2400
rect 1143 -2401 1144 -2400
rect 1262 -2401 1263 -2400
rect 331 -2403 332 -2402
rect 674 -2403 675 -2402
rect 695 -2403 696 -2402
rect 1391 -2403 1392 -2402
rect 254 -2405 255 -2404
rect 674 -2405 675 -2404
rect 898 -2405 899 -2404
rect 1713 -2405 1714 -2404
rect 117 -2407 118 -2406
rect 254 -2407 255 -2406
rect 341 -2407 342 -2406
rect 380 -2407 381 -2406
rect 404 -2407 405 -2406
rect 1528 -2407 1529 -2406
rect 345 -2409 346 -2408
rect 394 -2409 395 -2408
rect 569 -2409 570 -2408
rect 611 -2409 612 -2408
rect 656 -2409 657 -2408
rect 1143 -2409 1144 -2408
rect 373 -2411 374 -2410
rect 555 -2411 556 -2410
rect 576 -2411 577 -2410
rect 1122 -2411 1123 -2410
rect 373 -2413 374 -2412
rect 796 -2413 797 -2412
rect 1108 -2413 1109 -2412
rect 1122 -2413 1123 -2412
rect 597 -2415 598 -2414
rect 611 -2415 612 -2414
rect 1073 -2415 1074 -2414
rect 1108 -2415 1109 -2414
rect 345 -2417 346 -2416
rect 597 -2417 598 -2416
rect 604 -2417 605 -2416
rect 660 -2417 661 -2416
rect 1073 -2417 1074 -2416
rect 1367 -2417 1368 -2416
rect 660 -2419 661 -2418
rect 950 -2419 951 -2418
rect 1367 -2419 1368 -2418
rect 1472 -2419 1473 -2418
rect 1311 -2421 1312 -2420
rect 1472 -2421 1473 -2420
rect 1311 -2423 1312 -2422
rect 1353 -2423 1354 -2422
rect 1297 -2425 1298 -2424
rect 1353 -2425 1354 -2424
rect 1297 -2427 1298 -2426
rect 1409 -2427 1410 -2426
rect 1381 -2429 1382 -2428
rect 1409 -2429 1410 -2428
rect 1234 -2431 1235 -2430
rect 1381 -2431 1382 -2430
rect 758 -2433 759 -2432
rect 1234 -2433 1235 -2432
rect 744 -2435 745 -2434
rect 758 -2435 759 -2434
rect 744 -2437 745 -2436
rect 751 -2437 752 -2436
rect 716 -2439 717 -2438
rect 751 -2439 752 -2438
rect 9 -2450 10 -2449
rect 597 -2450 598 -2449
rect 723 -2450 724 -2449
rect 1017 -2450 1018 -2449
rect 1020 -2450 1021 -2449
rect 1486 -2450 1487 -2449
rect 1741 -2450 1742 -2449
rect 1773 -2450 1774 -2449
rect 1808 -2450 1809 -2449
rect 1815 -2450 1816 -2449
rect 16 -2452 17 -2451
rect 23 -2452 24 -2451
rect 44 -2452 45 -2451
rect 387 -2452 388 -2451
rect 408 -2452 409 -2451
rect 719 -2452 720 -2451
rect 726 -2452 727 -2451
rect 1717 -2452 1718 -2451
rect 1752 -2452 1753 -2451
rect 1759 -2452 1760 -2451
rect 1773 -2452 1774 -2451
rect 1794 -2452 1795 -2451
rect 1801 -2452 1802 -2451
rect 1808 -2452 1809 -2451
rect 16 -2454 17 -2453
rect 677 -2454 678 -2453
rect 807 -2454 808 -2453
rect 810 -2454 811 -2453
rect 828 -2454 829 -2453
rect 852 -2454 853 -2453
rect 884 -2454 885 -2453
rect 912 -2454 913 -2453
rect 950 -2454 951 -2453
rect 1381 -2454 1382 -2453
rect 1619 -2454 1620 -2453
rect 1717 -2454 1718 -2453
rect 1759 -2454 1760 -2453
rect 1766 -2454 1767 -2453
rect 44 -2456 45 -2455
rect 149 -2456 150 -2455
rect 159 -2456 160 -2455
rect 432 -2456 433 -2455
rect 439 -2456 440 -2455
rect 1094 -2456 1095 -2455
rect 1132 -2456 1133 -2455
rect 1521 -2456 1522 -2455
rect 1570 -2456 1571 -2455
rect 1766 -2456 1767 -2455
rect 51 -2458 52 -2457
rect 544 -2458 545 -2457
rect 583 -2458 584 -2457
rect 786 -2458 787 -2457
rect 807 -2458 808 -2457
rect 954 -2458 955 -2457
rect 982 -2458 983 -2457
rect 1118 -2458 1119 -2457
rect 1150 -2458 1151 -2457
rect 1486 -2458 1487 -2457
rect 1521 -2458 1522 -2457
rect 1542 -2458 1543 -2457
rect 1619 -2458 1620 -2457
rect 1668 -2458 1669 -2457
rect 51 -2460 52 -2459
rect 576 -2460 577 -2459
rect 597 -2460 598 -2459
rect 821 -2460 822 -2459
rect 828 -2460 829 -2459
rect 863 -2460 864 -2459
rect 884 -2460 885 -2459
rect 926 -2460 927 -2459
rect 940 -2460 941 -2459
rect 954 -2460 955 -2459
rect 968 -2460 969 -2459
rect 982 -2460 983 -2459
rect 1055 -2460 1056 -2459
rect 1248 -2460 1249 -2459
rect 1325 -2460 1326 -2459
rect 1339 -2460 1340 -2459
rect 1381 -2460 1382 -2459
rect 1395 -2460 1396 -2459
rect 1542 -2460 1543 -2459
rect 1556 -2460 1557 -2459
rect 1668 -2460 1669 -2459
rect 1710 -2460 1711 -2459
rect 58 -2462 59 -2461
rect 401 -2462 402 -2461
rect 408 -2462 409 -2461
rect 712 -2462 713 -2461
rect 786 -2462 787 -2461
rect 842 -2462 843 -2461
rect 887 -2462 888 -2461
rect 1731 -2462 1732 -2461
rect 58 -2464 59 -2463
rect 261 -2464 262 -2463
rect 324 -2464 325 -2463
rect 723 -2464 724 -2463
rect 821 -2464 822 -2463
rect 1045 -2464 1046 -2463
rect 1076 -2464 1077 -2463
rect 1696 -2464 1697 -2463
rect 30 -2466 31 -2465
rect 261 -2466 262 -2465
rect 275 -2466 276 -2465
rect 324 -2466 325 -2465
rect 352 -2466 353 -2465
rect 1395 -2466 1396 -2465
rect 1556 -2466 1557 -2465
rect 1675 -2466 1676 -2465
rect 1689 -2466 1690 -2465
rect 1710 -2466 1711 -2465
rect 30 -2468 31 -2467
rect 212 -2468 213 -2467
rect 226 -2468 227 -2467
rect 401 -2468 402 -2467
rect 429 -2468 430 -2467
rect 611 -2468 612 -2467
rect 842 -2468 843 -2467
rect 1066 -2468 1067 -2467
rect 1087 -2468 1088 -2467
rect 1094 -2468 1095 -2467
rect 1150 -2468 1151 -2467
rect 1178 -2468 1179 -2467
rect 1195 -2468 1196 -2467
rect 1633 -2468 1634 -2467
rect 1640 -2468 1641 -2467
rect 1731 -2468 1732 -2467
rect 65 -2470 66 -2469
rect 390 -2470 391 -2469
rect 450 -2470 451 -2469
rect 516 -2470 517 -2469
rect 530 -2470 531 -2469
rect 569 -2470 570 -2469
rect 600 -2470 601 -2469
rect 1178 -2470 1179 -2469
rect 1325 -2470 1326 -2469
rect 1374 -2470 1375 -2469
rect 1640 -2470 1641 -2469
rect 1654 -2470 1655 -2469
rect 1675 -2470 1676 -2469
rect 1724 -2470 1725 -2469
rect 65 -2472 66 -2471
rect 317 -2472 318 -2471
rect 352 -2472 353 -2471
rect 1167 -2472 1168 -2471
rect 1332 -2472 1333 -2471
rect 1801 -2472 1802 -2471
rect 72 -2474 73 -2473
rect 387 -2474 388 -2473
rect 457 -2474 458 -2473
rect 583 -2474 584 -2473
rect 600 -2474 601 -2473
rect 695 -2474 696 -2473
rect 905 -2474 906 -2473
rect 912 -2474 913 -2473
rect 940 -2474 941 -2473
rect 1059 -2474 1060 -2473
rect 1066 -2474 1067 -2473
rect 1129 -2474 1130 -2473
rect 1160 -2474 1161 -2473
rect 1661 -2474 1662 -2473
rect 1689 -2474 1690 -2473
rect 1738 -2474 1739 -2473
rect 72 -2476 73 -2475
rect 194 -2476 195 -2475
rect 198 -2476 199 -2475
rect 212 -2476 213 -2475
rect 226 -2476 227 -2475
rect 947 -2476 948 -2475
rect 971 -2476 972 -2475
rect 1374 -2476 1375 -2475
rect 1598 -2476 1599 -2475
rect 1724 -2476 1725 -2475
rect 1738 -2476 1739 -2475
rect 1780 -2476 1781 -2475
rect 82 -2478 83 -2477
rect 233 -2478 234 -2477
rect 243 -2478 244 -2477
rect 1010 -2478 1011 -2477
rect 1048 -2478 1049 -2477
rect 1661 -2478 1662 -2477
rect 1696 -2478 1697 -2477
rect 1787 -2478 1788 -2477
rect 93 -2480 94 -2479
rect 380 -2480 381 -2479
rect 443 -2480 444 -2479
rect 1598 -2480 1599 -2479
rect 1654 -2480 1655 -2479
rect 1682 -2480 1683 -2479
rect 93 -2482 94 -2481
rect 268 -2482 269 -2481
rect 275 -2482 276 -2481
rect 394 -2482 395 -2481
rect 443 -2482 444 -2481
rect 506 -2482 507 -2481
rect 513 -2482 514 -2481
rect 590 -2482 591 -2481
rect 681 -2482 682 -2481
rect 695 -2482 696 -2481
rect 740 -2482 741 -2481
rect 947 -2482 948 -2481
rect 996 -2482 997 -2481
rect 1010 -2482 1011 -2481
rect 1087 -2482 1088 -2481
rect 1388 -2482 1389 -2481
rect 96 -2484 97 -2483
rect 345 -2484 346 -2483
rect 366 -2484 367 -2483
rect 394 -2484 395 -2483
rect 457 -2484 458 -2483
rect 849 -2484 850 -2483
rect 877 -2484 878 -2483
rect 905 -2484 906 -2483
rect 989 -2484 990 -2483
rect 996 -2484 997 -2483
rect 1129 -2484 1130 -2483
rect 1248 -2484 1249 -2483
rect 1255 -2484 1256 -2483
rect 1682 -2484 1683 -2483
rect 37 -2486 38 -2485
rect 345 -2486 346 -2485
rect 366 -2486 367 -2485
rect 618 -2486 619 -2485
rect 653 -2486 654 -2485
rect 681 -2486 682 -2485
rect 810 -2486 811 -2485
rect 1059 -2486 1060 -2485
rect 1115 -2486 1116 -2485
rect 1255 -2486 1256 -2485
rect 1321 -2486 1322 -2485
rect 1780 -2486 1781 -2485
rect 37 -2488 38 -2487
rect 114 -2488 115 -2487
rect 128 -2488 129 -2487
rect 289 -2488 290 -2487
rect 317 -2488 318 -2487
rect 460 -2488 461 -2487
rect 471 -2488 472 -2487
rect 527 -2488 528 -2487
rect 541 -2488 542 -2487
rect 660 -2488 661 -2487
rect 849 -2488 850 -2487
rect 926 -2488 927 -2487
rect 989 -2488 990 -2487
rect 1318 -2488 1319 -2487
rect 1332 -2488 1333 -2487
rect 1493 -2488 1494 -2487
rect 100 -2490 101 -2489
rect 114 -2490 115 -2489
rect 128 -2490 129 -2489
rect 282 -2490 283 -2489
rect 289 -2490 290 -2489
rect 303 -2490 304 -2489
rect 415 -2490 416 -2489
rect 471 -2490 472 -2489
rect 478 -2490 479 -2489
rect 590 -2490 591 -2489
rect 604 -2490 605 -2489
rect 660 -2490 661 -2489
rect 1115 -2490 1116 -2489
rect 1297 -2490 1298 -2489
rect 1318 -2490 1319 -2489
rect 1360 -2490 1361 -2489
rect 1367 -2490 1368 -2489
rect 1493 -2490 1494 -2489
rect 100 -2492 101 -2491
rect 1346 -2492 1347 -2491
rect 1367 -2492 1368 -2491
rect 1465 -2492 1466 -2491
rect 107 -2494 108 -2493
rect 338 -2494 339 -2493
rect 478 -2494 479 -2493
rect 737 -2494 738 -2493
rect 1003 -2494 1004 -2493
rect 1346 -2494 1347 -2493
rect 1388 -2494 1389 -2493
rect 1402 -2494 1403 -2493
rect 1465 -2494 1466 -2493
rect 1479 -2494 1480 -2493
rect 107 -2496 108 -2495
rect 1185 -2496 1186 -2495
rect 1241 -2496 1242 -2495
rect 1787 -2496 1788 -2495
rect 110 -2498 111 -2497
rect 1017 -2498 1018 -2497
rect 1101 -2498 1102 -2497
rect 1185 -2498 1186 -2497
rect 1241 -2498 1242 -2497
rect 1290 -2498 1291 -2497
rect 1402 -2498 1403 -2497
rect 1409 -2498 1410 -2497
rect 1479 -2498 1480 -2497
rect 1507 -2498 1508 -2497
rect 103 -2500 104 -2499
rect 1101 -2500 1102 -2499
rect 1157 -2500 1158 -2499
rect 1297 -2500 1298 -2499
rect 1409 -2500 1410 -2499
rect 1416 -2500 1417 -2499
rect 131 -2502 132 -2501
rect 863 -2502 864 -2501
rect 1164 -2502 1165 -2501
rect 1311 -2502 1312 -2501
rect 1416 -2502 1417 -2501
rect 1437 -2502 1438 -2501
rect 135 -2504 136 -2503
rect 436 -2504 437 -2503
rect 485 -2504 486 -2503
rect 576 -2504 577 -2503
rect 604 -2504 605 -2503
rect 1020 -2504 1021 -2503
rect 1164 -2504 1165 -2503
rect 1199 -2504 1200 -2503
rect 1269 -2504 1270 -2503
rect 1360 -2504 1361 -2503
rect 1437 -2504 1438 -2503
rect 1451 -2504 1452 -2503
rect 135 -2506 136 -2505
rect 1045 -2506 1046 -2505
rect 1080 -2506 1081 -2505
rect 1269 -2506 1270 -2505
rect 1290 -2506 1291 -2505
rect 1514 -2506 1515 -2505
rect 142 -2508 143 -2507
rect 415 -2508 416 -2507
rect 436 -2508 437 -2507
rect 1031 -2508 1032 -2507
rect 1080 -2508 1081 -2507
rect 1136 -2508 1137 -2507
rect 1311 -2508 1312 -2507
rect 1699 -2508 1700 -2507
rect 121 -2510 122 -2509
rect 142 -2510 143 -2509
rect 149 -2510 150 -2509
rect 1633 -2510 1634 -2509
rect 121 -2512 122 -2511
rect 156 -2512 157 -2511
rect 163 -2512 164 -2511
rect 380 -2512 381 -2511
rect 485 -2512 486 -2511
rect 835 -2512 836 -2511
rect 1024 -2512 1025 -2511
rect 1031 -2512 1032 -2511
rect 1122 -2512 1123 -2511
rect 1199 -2512 1200 -2511
rect 1514 -2512 1515 -2511
rect 1528 -2512 1529 -2511
rect 152 -2514 153 -2513
rect 611 -2514 612 -2513
rect 639 -2514 640 -2513
rect 653 -2514 654 -2513
rect 674 -2514 675 -2513
rect 1451 -2514 1452 -2513
rect 1528 -2514 1529 -2513
rect 1703 -2514 1704 -2513
rect 163 -2516 164 -2515
rect 1052 -2516 1053 -2515
rect 1073 -2516 1074 -2515
rect 1703 -2516 1704 -2515
rect 170 -2518 171 -2517
rect 338 -2518 339 -2517
rect 492 -2518 493 -2517
rect 831 -2518 832 -2517
rect 1108 -2518 1109 -2517
rect 1122 -2518 1123 -2517
rect 170 -2520 171 -2519
rect 1143 -2520 1144 -2519
rect 173 -2522 174 -2521
rect 310 -2522 311 -2521
rect 492 -2522 493 -2521
rect 499 -2522 500 -2521
rect 506 -2522 507 -2521
rect 688 -2522 689 -2521
rect 702 -2522 703 -2521
rect 1024 -2522 1025 -2521
rect 1108 -2522 1109 -2521
rect 1192 -2522 1193 -2521
rect 191 -2524 192 -2523
rect 877 -2524 878 -2523
rect 1143 -2524 1144 -2523
rect 1206 -2524 1207 -2523
rect 191 -2526 192 -2525
rect 870 -2526 871 -2525
rect 1192 -2526 1193 -2525
rect 1444 -2526 1445 -2525
rect 198 -2528 199 -2527
rect 558 -2528 559 -2527
rect 569 -2528 570 -2527
rect 961 -2528 962 -2527
rect 1206 -2528 1207 -2527
rect 1220 -2528 1221 -2527
rect 1444 -2528 1445 -2527
rect 1458 -2528 1459 -2527
rect 219 -2530 220 -2529
rect 618 -2530 619 -2529
rect 667 -2530 668 -2529
rect 702 -2530 703 -2529
rect 737 -2530 738 -2529
rect 1570 -2530 1571 -2529
rect 219 -2532 220 -2531
rect 464 -2532 465 -2531
rect 499 -2532 500 -2531
rect 534 -2532 535 -2531
rect 674 -2532 675 -2531
rect 709 -2532 710 -2531
rect 789 -2532 790 -2531
rect 835 -2532 836 -2531
rect 870 -2532 871 -2531
rect 933 -2532 934 -2531
rect 961 -2532 962 -2531
rect 975 -2532 976 -2531
rect 1220 -2532 1221 -2531
rect 1276 -2532 1277 -2531
rect 233 -2534 234 -2533
rect 240 -2534 241 -2533
rect 247 -2534 248 -2533
rect 450 -2534 451 -2533
rect 464 -2534 465 -2533
rect 548 -2534 549 -2533
rect 688 -2534 689 -2533
rect 751 -2534 752 -2533
rect 975 -2534 976 -2533
rect 1171 -2534 1172 -2533
rect 1276 -2534 1277 -2533
rect 1472 -2534 1473 -2533
rect 247 -2536 248 -2535
rect 1157 -2536 1158 -2535
rect 1171 -2536 1172 -2535
rect 1535 -2536 1536 -2535
rect 254 -2538 255 -2537
rect 303 -2538 304 -2537
rect 310 -2538 311 -2537
rect 628 -2538 629 -2537
rect 709 -2538 710 -2537
rect 1003 -2538 1004 -2537
rect 1472 -2538 1473 -2537
rect 1500 -2538 1501 -2537
rect 1535 -2538 1536 -2537
rect 1549 -2538 1550 -2537
rect 254 -2540 255 -2539
rect 373 -2540 374 -2539
rect 513 -2540 514 -2539
rect 555 -2540 556 -2539
rect 730 -2540 731 -2539
rect 933 -2540 934 -2539
rect 1500 -2540 1501 -2539
rect 1563 -2540 1564 -2539
rect 268 -2542 269 -2541
rect 716 -2542 717 -2541
rect 730 -2542 731 -2541
rect 1174 -2542 1175 -2541
rect 1549 -2542 1550 -2541
rect 1577 -2542 1578 -2541
rect 282 -2544 283 -2543
rect 331 -2544 332 -2543
rect 359 -2544 360 -2543
rect 373 -2544 374 -2543
rect 520 -2544 521 -2543
rect 555 -2544 556 -2543
rect 716 -2544 717 -2543
rect 758 -2544 759 -2543
rect 1563 -2544 1564 -2543
rect 1584 -2544 1585 -2543
rect 177 -2546 178 -2545
rect 331 -2546 332 -2545
rect 520 -2546 521 -2545
rect 800 -2546 801 -2545
rect 1577 -2546 1578 -2545
rect 1591 -2546 1592 -2545
rect 177 -2548 178 -2547
rect 205 -2548 206 -2547
rect 527 -2548 528 -2547
rect 562 -2548 563 -2547
rect 625 -2548 626 -2547
rect 800 -2548 801 -2547
rect 1584 -2548 1585 -2547
rect 1605 -2548 1606 -2547
rect 184 -2550 185 -2549
rect 359 -2550 360 -2549
rect 534 -2550 535 -2549
rect 744 -2550 745 -2549
rect 751 -2550 752 -2549
rect 1213 -2550 1214 -2549
rect 1591 -2550 1592 -2549
rect 1647 -2550 1648 -2549
rect 184 -2552 185 -2551
rect 341 -2552 342 -2551
rect 548 -2552 549 -2551
rect 992 -2552 993 -2551
rect 1213 -2552 1214 -2551
rect 1227 -2552 1228 -2551
rect 1283 -2552 1284 -2551
rect 1647 -2552 1648 -2551
rect 205 -2554 206 -2553
rect 422 -2554 423 -2553
rect 562 -2554 563 -2553
rect 639 -2554 640 -2553
rect 744 -2554 745 -2553
rect 765 -2554 766 -2553
rect 968 -2554 969 -2553
rect 1227 -2554 1228 -2553
rect 1262 -2554 1263 -2553
rect 1283 -2554 1284 -2553
rect 1605 -2554 1606 -2553
rect 1612 -2554 1613 -2553
rect 156 -2556 157 -2555
rect 422 -2556 423 -2555
rect 625 -2556 626 -2555
rect 1458 -2556 1459 -2555
rect 1612 -2556 1613 -2555
rect 1626 -2556 1627 -2555
rect 79 -2558 80 -2557
rect 1626 -2558 1627 -2557
rect 79 -2560 80 -2559
rect 296 -2560 297 -2559
rect 758 -2560 759 -2559
rect 772 -2560 773 -2559
rect 1262 -2560 1263 -2559
rect 1430 -2560 1431 -2559
rect 296 -2562 297 -2561
rect 404 -2562 405 -2561
rect 765 -2562 766 -2561
rect 779 -2562 780 -2561
rect 1234 -2562 1235 -2561
rect 1430 -2562 1431 -2561
rect 772 -2564 773 -2563
rect 793 -2564 794 -2563
rect 1234 -2564 1235 -2563
rect 1304 -2564 1305 -2563
rect 110 -2566 111 -2565
rect 1304 -2566 1305 -2565
rect 670 -2568 671 -2567
rect 793 -2568 794 -2567
rect 779 -2570 780 -2569
rect 898 -2570 899 -2569
rect 891 -2572 892 -2571
rect 898 -2572 899 -2571
rect 453 -2574 454 -2573
rect 891 -2574 892 -2573
rect 9 -2585 10 -2584
rect 443 -2585 444 -2584
rect 450 -2585 451 -2584
rect 1059 -2585 1060 -2584
rect 1062 -2585 1063 -2584
rect 1276 -2585 1277 -2584
rect 1293 -2585 1294 -2584
rect 1339 -2585 1340 -2584
rect 1510 -2585 1511 -2584
rect 1591 -2585 1592 -2584
rect 1738 -2585 1739 -2584
rect 1780 -2585 1781 -2584
rect 44 -2587 45 -2586
rect 628 -2587 629 -2586
rect 639 -2587 640 -2586
rect 807 -2587 808 -2586
rect 852 -2587 853 -2586
rect 996 -2587 997 -2586
rect 1020 -2587 1021 -2586
rect 1108 -2587 1109 -2586
rect 1115 -2587 1116 -2586
rect 1311 -2587 1312 -2586
rect 1339 -2587 1340 -2586
rect 1374 -2587 1375 -2586
rect 1769 -2587 1770 -2586
rect 1783 -2587 1784 -2586
rect 44 -2589 45 -2588
rect 779 -2589 780 -2588
rect 807 -2589 808 -2588
rect 828 -2589 829 -2588
rect 866 -2589 867 -2588
rect 1507 -2589 1508 -2588
rect 107 -2591 108 -2590
rect 366 -2591 367 -2590
rect 443 -2591 444 -2590
rect 583 -2591 584 -2590
rect 660 -2591 661 -2590
rect 712 -2591 713 -2590
rect 726 -2591 727 -2590
rect 1647 -2591 1648 -2590
rect 79 -2593 80 -2592
rect 107 -2593 108 -2592
rect 121 -2593 122 -2592
rect 240 -2593 241 -2592
rect 243 -2593 244 -2592
rect 282 -2593 283 -2592
rect 292 -2593 293 -2592
rect 597 -2593 598 -2592
rect 660 -2593 661 -2592
rect 870 -2593 871 -2592
rect 915 -2593 916 -2592
rect 1353 -2593 1354 -2592
rect 1507 -2593 1508 -2592
rect 1535 -2593 1536 -2592
rect 1647 -2593 1648 -2592
rect 1654 -2593 1655 -2592
rect 79 -2595 80 -2594
rect 842 -2595 843 -2594
rect 947 -2595 948 -2594
rect 1244 -2595 1245 -2594
rect 1276 -2595 1277 -2594
rect 1304 -2595 1305 -2594
rect 1311 -2595 1312 -2594
rect 1388 -2595 1389 -2594
rect 1654 -2595 1655 -2594
rect 1776 -2595 1777 -2594
rect 121 -2597 122 -2596
rect 128 -2597 129 -2596
rect 149 -2597 150 -2596
rect 387 -2597 388 -2596
rect 457 -2597 458 -2596
rect 670 -2597 671 -2596
rect 695 -2597 696 -2596
rect 712 -2597 713 -2596
rect 737 -2597 738 -2596
rect 1486 -2597 1487 -2596
rect 68 -2599 69 -2598
rect 149 -2599 150 -2598
rect 156 -2599 157 -2598
rect 254 -2599 255 -2598
rect 275 -2599 276 -2598
rect 558 -2599 559 -2598
rect 642 -2599 643 -2598
rect 1535 -2599 1536 -2598
rect 86 -2601 87 -2600
rect 128 -2601 129 -2600
rect 142 -2601 143 -2600
rect 275 -2601 276 -2600
rect 282 -2601 283 -2600
rect 289 -2601 290 -2600
rect 296 -2601 297 -2600
rect 586 -2601 587 -2600
rect 681 -2601 682 -2600
rect 737 -2601 738 -2600
rect 765 -2601 766 -2600
rect 779 -2601 780 -2600
rect 842 -2601 843 -2600
rect 884 -2601 885 -2600
rect 968 -2601 969 -2600
rect 1430 -2601 1431 -2600
rect 1486 -2601 1487 -2600
rect 1542 -2601 1543 -2600
rect 86 -2603 87 -2602
rect 100 -2603 101 -2602
rect 103 -2603 104 -2602
rect 289 -2603 290 -2602
rect 296 -2603 297 -2602
rect 1017 -2603 1018 -2602
rect 1048 -2603 1049 -2602
rect 1290 -2603 1291 -2602
rect 1304 -2603 1305 -2602
rect 1360 -2603 1361 -2602
rect 1430 -2603 1431 -2602
rect 1444 -2603 1445 -2602
rect 1542 -2603 1543 -2602
rect 1570 -2603 1571 -2602
rect 37 -2605 38 -2604
rect 100 -2605 101 -2604
rect 142 -2605 143 -2604
rect 436 -2605 437 -2604
rect 453 -2605 454 -2604
rect 681 -2605 682 -2604
rect 695 -2605 696 -2604
rect 877 -2605 878 -2604
rect 905 -2605 906 -2604
rect 968 -2605 969 -2604
rect 971 -2605 972 -2604
rect 1703 -2605 1704 -2604
rect 37 -2607 38 -2606
rect 845 -2607 846 -2606
rect 856 -2607 857 -2606
rect 877 -2607 878 -2606
rect 905 -2607 906 -2606
rect 950 -2607 951 -2606
rect 989 -2607 990 -2606
rect 1038 -2607 1039 -2606
rect 1073 -2607 1074 -2606
rect 1094 -2607 1095 -2606
rect 1108 -2607 1109 -2606
rect 1143 -2607 1144 -2606
rect 1157 -2607 1158 -2606
rect 1220 -2607 1221 -2606
rect 1262 -2607 1263 -2606
rect 1388 -2607 1389 -2606
rect 1444 -2607 1445 -2606
rect 1458 -2607 1459 -2606
rect 1570 -2607 1571 -2606
rect 1598 -2607 1599 -2606
rect 1675 -2607 1676 -2606
rect 1703 -2607 1704 -2606
rect 156 -2609 157 -2608
rect 198 -2609 199 -2608
rect 205 -2609 206 -2608
rect 450 -2609 451 -2608
rect 492 -2609 493 -2608
rect 765 -2609 766 -2608
rect 775 -2609 776 -2608
rect 1374 -2609 1375 -2608
rect 1458 -2609 1459 -2608
rect 1514 -2609 1515 -2608
rect 1598 -2609 1599 -2608
rect 1619 -2609 1620 -2608
rect 1675 -2609 1676 -2608
rect 1717 -2609 1718 -2608
rect 159 -2611 160 -2610
rect 926 -2611 927 -2610
rect 940 -2611 941 -2610
rect 1143 -2611 1144 -2610
rect 1174 -2611 1175 -2610
rect 1332 -2611 1333 -2610
rect 1353 -2611 1354 -2610
rect 1409 -2611 1410 -2610
rect 1514 -2611 1515 -2610
rect 1699 -2611 1700 -2610
rect 1710 -2611 1711 -2610
rect 1717 -2611 1718 -2610
rect 170 -2613 171 -2612
rect 1248 -2613 1249 -2612
rect 1409 -2613 1410 -2612
rect 1605 -2613 1606 -2612
rect 1689 -2613 1690 -2612
rect 1710 -2613 1711 -2612
rect 170 -2615 171 -2614
rect 604 -2615 605 -2614
rect 702 -2615 703 -2614
rect 740 -2615 741 -2614
rect 856 -2615 857 -2614
rect 1052 -2615 1053 -2614
rect 1066 -2615 1067 -2614
rect 1332 -2615 1333 -2614
rect 1556 -2615 1557 -2614
rect 1605 -2615 1606 -2614
rect 1689 -2615 1690 -2614
rect 1766 -2615 1767 -2614
rect 173 -2617 174 -2616
rect 1101 -2617 1102 -2616
rect 1118 -2617 1119 -2616
rect 1591 -2617 1592 -2616
rect 177 -2619 178 -2618
rect 254 -2619 255 -2618
rect 303 -2619 304 -2618
rect 457 -2619 458 -2618
rect 492 -2619 493 -2618
rect 730 -2619 731 -2618
rect 828 -2619 829 -2618
rect 1766 -2619 1767 -2618
rect 23 -2621 24 -2620
rect 177 -2621 178 -2620
rect 184 -2621 185 -2620
rect 667 -2621 668 -2620
rect 702 -2621 703 -2620
rect 786 -2621 787 -2620
rect 870 -2621 871 -2620
rect 1052 -2621 1053 -2620
rect 1076 -2621 1077 -2620
rect 1185 -2621 1186 -2620
rect 1220 -2621 1221 -2620
rect 1318 -2621 1319 -2620
rect 1556 -2621 1557 -2620
rect 1584 -2621 1585 -2620
rect 184 -2623 185 -2622
rect 198 -2623 199 -2622
rect 205 -2623 206 -2622
rect 345 -2623 346 -2622
rect 387 -2623 388 -2622
rect 688 -2623 689 -2622
rect 709 -2623 710 -2622
rect 1206 -2623 1207 -2622
rect 1241 -2623 1242 -2622
rect 1262 -2623 1263 -2622
rect 1584 -2623 1585 -2622
rect 1612 -2623 1613 -2622
rect 226 -2625 227 -2624
rect 1020 -2625 1021 -2624
rect 1024 -2625 1025 -2624
rect 1038 -2625 1039 -2624
rect 1094 -2625 1095 -2624
rect 1150 -2625 1151 -2624
rect 1241 -2625 1242 -2624
rect 1367 -2625 1368 -2624
rect 1612 -2625 1613 -2624
rect 1626 -2625 1627 -2624
rect 30 -2627 31 -2626
rect 226 -2627 227 -2626
rect 303 -2627 304 -2626
rect 485 -2627 486 -2626
rect 513 -2627 514 -2626
rect 604 -2627 605 -2626
rect 646 -2627 647 -2626
rect 667 -2627 668 -2626
rect 723 -2627 724 -2626
rect 1360 -2627 1361 -2626
rect 1367 -2627 1368 -2626
rect 1493 -2627 1494 -2626
rect 1626 -2627 1627 -2626
rect 1633 -2627 1634 -2626
rect 30 -2629 31 -2628
rect 65 -2629 66 -2628
rect 310 -2629 311 -2628
rect 425 -2629 426 -2628
rect 436 -2629 437 -2628
rect 716 -2629 717 -2628
rect 730 -2629 731 -2628
rect 744 -2629 745 -2628
rect 786 -2629 787 -2628
rect 1171 -2629 1172 -2628
rect 1248 -2629 1249 -2628
rect 1321 -2629 1322 -2628
rect 1479 -2629 1480 -2628
rect 1493 -2629 1494 -2628
rect 1633 -2629 1634 -2628
rect 1731 -2629 1732 -2628
rect 58 -2631 59 -2630
rect 513 -2631 514 -2630
rect 520 -2631 521 -2630
rect 852 -2631 853 -2630
rect 912 -2631 913 -2630
rect 926 -2631 927 -2630
rect 933 -2631 934 -2630
rect 1206 -2631 1207 -2630
rect 1731 -2631 1732 -2630
rect 1745 -2631 1746 -2630
rect 58 -2633 59 -2632
rect 800 -2633 801 -2632
rect 835 -2633 836 -2632
rect 933 -2633 934 -2632
rect 940 -2633 941 -2632
rect 1395 -2633 1396 -2632
rect 1745 -2633 1746 -2632
rect 1752 -2633 1753 -2632
rect 110 -2635 111 -2634
rect 310 -2635 311 -2634
rect 338 -2635 339 -2634
rect 366 -2635 367 -2634
rect 380 -2635 381 -2634
rect 688 -2635 689 -2634
rect 716 -2635 717 -2634
rect 1318 -2635 1319 -2634
rect 1395 -2635 1396 -2634
rect 1416 -2635 1417 -2634
rect 1752 -2635 1753 -2634
rect 1759 -2635 1760 -2634
rect 135 -2637 136 -2636
rect 835 -2637 836 -2636
rect 919 -2637 920 -2636
rect 1185 -2637 1186 -2636
rect 1416 -2637 1417 -2636
rect 1472 -2637 1473 -2636
rect 1759 -2637 1760 -2636
rect 1773 -2637 1774 -2636
rect 135 -2639 136 -2638
rect 233 -2639 234 -2638
rect 338 -2639 339 -2638
rect 401 -2639 402 -2638
rect 408 -2639 409 -2638
rect 989 -2639 990 -2638
rect 996 -2639 997 -2638
rect 1010 -2639 1011 -2638
rect 1017 -2639 1018 -2638
rect 1682 -2639 1683 -2638
rect 72 -2641 73 -2640
rect 233 -2641 234 -2640
rect 345 -2641 346 -2640
rect 352 -2641 353 -2640
rect 359 -2641 360 -2640
rect 380 -2641 381 -2640
rect 394 -2641 395 -2640
rect 401 -2641 402 -2640
rect 422 -2641 423 -2640
rect 485 -2641 486 -2640
rect 520 -2641 521 -2640
rect 1661 -2641 1662 -2640
rect 72 -2643 73 -2642
rect 464 -2643 465 -2642
rect 523 -2643 524 -2642
rect 569 -2643 570 -2642
rect 646 -2643 647 -2642
rect 653 -2643 654 -2642
rect 674 -2643 675 -2642
rect 723 -2643 724 -2642
rect 800 -2643 801 -2642
rect 978 -2643 979 -2642
rect 1003 -2643 1004 -2642
rect 1066 -2643 1067 -2642
rect 1101 -2643 1102 -2642
rect 1164 -2643 1165 -2642
rect 1171 -2643 1172 -2642
rect 1297 -2643 1298 -2642
rect 1472 -2643 1473 -2642
rect 1521 -2643 1522 -2642
rect 152 -2645 153 -2644
rect 1661 -2645 1662 -2644
rect 201 -2647 202 -2646
rect 1479 -2647 1480 -2646
rect 1521 -2647 1522 -2646
rect 1549 -2647 1550 -2646
rect 268 -2649 269 -2648
rect 674 -2649 675 -2648
rect 891 -2649 892 -2648
rect 1010 -2649 1011 -2648
rect 1024 -2649 1025 -2648
rect 1080 -2649 1081 -2648
rect 1122 -2649 1123 -2648
rect 1136 -2649 1137 -2648
rect 1139 -2649 1140 -2648
rect 1738 -2649 1739 -2648
rect 268 -2651 269 -2650
rect 1160 -2651 1161 -2650
rect 1297 -2651 1298 -2650
rect 1325 -2651 1326 -2650
rect 1549 -2651 1550 -2650
rect 1577 -2651 1578 -2650
rect 324 -2653 325 -2652
rect 352 -2653 353 -2652
rect 359 -2653 360 -2652
rect 429 -2653 430 -2652
rect 464 -2653 465 -2652
rect 793 -2653 794 -2652
rect 821 -2653 822 -2652
rect 1136 -2653 1137 -2652
rect 1325 -2653 1326 -2652
rect 1619 -2653 1620 -2652
rect 324 -2655 325 -2654
rect 548 -2655 549 -2654
rect 569 -2655 570 -2654
rect 590 -2655 591 -2654
rect 625 -2655 626 -2654
rect 891 -2655 892 -2654
rect 912 -2655 913 -2654
rect 1080 -2655 1081 -2654
rect 1122 -2655 1123 -2654
rect 1178 -2655 1179 -2654
rect 1577 -2655 1578 -2654
rect 1741 -2655 1742 -2654
rect 163 -2657 164 -2656
rect 548 -2657 549 -2656
rect 590 -2657 591 -2656
rect 618 -2657 619 -2656
rect 625 -2657 626 -2656
rect 849 -2657 850 -2656
rect 954 -2657 955 -2656
rect 1003 -2657 1004 -2656
rect 1087 -2657 1088 -2656
rect 1178 -2657 1179 -2656
rect 163 -2659 164 -2658
rect 219 -2659 220 -2658
rect 373 -2659 374 -2658
rect 408 -2659 409 -2658
rect 415 -2659 416 -2658
rect 429 -2659 430 -2658
rect 506 -2659 507 -2658
rect 618 -2659 619 -2658
rect 632 -2659 633 -2658
rect 653 -2659 654 -2658
rect 772 -2659 773 -2658
rect 793 -2659 794 -2658
rect 814 -2659 815 -2658
rect 821 -2659 822 -2658
rect 849 -2659 850 -2658
rect 1682 -2659 1683 -2658
rect 219 -2661 220 -2660
rect 247 -2661 248 -2660
rect 331 -2661 332 -2660
rect 373 -2661 374 -2660
rect 394 -2661 395 -2660
rect 751 -2661 752 -2660
rect 814 -2661 815 -2660
rect 1199 -2661 1200 -2660
rect 93 -2663 94 -2662
rect 331 -2663 332 -2662
rect 415 -2663 416 -2662
rect 1195 -2663 1196 -2662
rect 1199 -2663 1200 -2662
rect 1213 -2663 1214 -2662
rect 93 -2665 94 -2664
rect 114 -2665 115 -2664
rect 191 -2665 192 -2664
rect 247 -2665 248 -2664
rect 478 -2665 479 -2664
rect 772 -2665 773 -2664
rect 863 -2665 864 -2664
rect 954 -2665 955 -2664
rect 961 -2665 962 -2664
rect 1164 -2665 1165 -2664
rect 1195 -2665 1196 -2664
rect 1500 -2665 1501 -2664
rect 114 -2667 115 -2666
rect 208 -2667 209 -2666
rect 471 -2667 472 -2666
rect 478 -2667 479 -2666
rect 506 -2667 507 -2666
rect 562 -2667 563 -2666
rect 597 -2667 598 -2666
rect 632 -2667 633 -2666
rect 635 -2667 636 -2666
rect 751 -2667 752 -2666
rect 961 -2667 962 -2666
rect 982 -2667 983 -2666
rect 1045 -2667 1046 -2666
rect 1087 -2667 1088 -2666
rect 1132 -2667 1133 -2666
rect 1668 -2667 1669 -2666
rect 191 -2669 192 -2668
rect 212 -2669 213 -2668
rect 471 -2669 472 -2668
rect 1150 -2669 1151 -2668
rect 1213 -2669 1214 -2668
rect 1801 -2669 1802 -2668
rect 51 -2671 52 -2670
rect 212 -2671 213 -2670
rect 499 -2671 500 -2670
rect 562 -2671 563 -2670
rect 975 -2671 976 -2670
rect 982 -2671 983 -2670
rect 1045 -2671 1046 -2670
rect 1346 -2671 1347 -2670
rect 1500 -2671 1501 -2670
rect 1787 -2671 1788 -2670
rect 1801 -2671 1802 -2670
rect 1808 -2671 1809 -2670
rect 51 -2673 52 -2672
rect 422 -2673 423 -2672
rect 499 -2673 500 -2672
rect 583 -2673 584 -2672
rect 975 -2673 976 -2672
rect 1031 -2673 1032 -2672
rect 1346 -2673 1347 -2672
rect 1381 -2673 1382 -2672
rect 1528 -2673 1529 -2672
rect 1668 -2673 1669 -2672
rect 1787 -2673 1788 -2672
rect 1794 -2673 1795 -2672
rect 1808 -2673 1809 -2672
rect 1815 -2673 1816 -2672
rect 527 -2675 528 -2674
rect 530 -2675 531 -2674
rect 534 -2675 535 -2674
rect 744 -2675 745 -2674
rect 1381 -2675 1382 -2674
rect 1402 -2675 1403 -2674
rect 1696 -2675 1697 -2674
rect 1794 -2675 1795 -2674
rect 527 -2677 528 -2676
rect 541 -2677 542 -2676
rect 555 -2677 556 -2676
rect 1696 -2677 1697 -2676
rect 530 -2679 531 -2678
rect 541 -2679 542 -2678
rect 555 -2679 556 -2678
rect 576 -2679 577 -2678
rect 611 -2679 612 -2678
rect 1031 -2679 1032 -2678
rect 1192 -2679 1193 -2678
rect 1402 -2679 1403 -2678
rect 534 -2681 535 -2680
rect 1055 -2681 1056 -2680
rect 576 -2683 577 -2682
rect 1773 -2683 1774 -2682
rect 611 -2685 612 -2684
rect 1129 -2685 1130 -2684
rect 709 -2687 710 -2686
rect 1528 -2687 1529 -2686
rect 1055 -2689 1056 -2688
rect 1640 -2689 1641 -2688
rect 1059 -2691 1060 -2690
rect 1129 -2691 1130 -2690
rect 1269 -2691 1270 -2690
rect 1640 -2691 1641 -2690
rect 1234 -2693 1235 -2692
rect 1269 -2693 1270 -2692
rect 1227 -2695 1228 -2694
rect 1234 -2695 1235 -2694
rect 1227 -2697 1228 -2696
rect 1283 -2697 1284 -2696
rect 1255 -2699 1256 -2698
rect 1283 -2699 1284 -2698
rect 1255 -2701 1256 -2700
rect 1451 -2701 1452 -2700
rect 1423 -2703 1424 -2702
rect 1451 -2703 1452 -2702
rect 1423 -2705 1424 -2704
rect 1437 -2705 1438 -2704
rect 1192 -2707 1193 -2706
rect 1437 -2707 1438 -2706
rect 30 -2718 31 -2717
rect 712 -2718 713 -2717
rect 737 -2718 738 -2717
rect 772 -2718 773 -2717
rect 842 -2718 843 -2717
rect 1493 -2718 1494 -2717
rect 1769 -2718 1770 -2717
rect 1808 -2718 1809 -2717
rect 44 -2720 45 -2719
rect 68 -2720 69 -2719
rect 72 -2720 73 -2719
rect 642 -2720 643 -2719
rect 712 -2720 713 -2719
rect 1195 -2720 1196 -2719
rect 1290 -2720 1291 -2719
rect 1360 -2720 1361 -2719
rect 1433 -2720 1434 -2719
rect 1451 -2720 1452 -2719
rect 1493 -2720 1494 -2719
rect 1507 -2720 1508 -2719
rect 1780 -2720 1781 -2719
rect 1801 -2720 1802 -2719
rect 58 -2722 59 -2721
rect 72 -2722 73 -2721
rect 96 -2722 97 -2721
rect 142 -2722 143 -2721
rect 198 -2722 199 -2721
rect 1776 -2722 1777 -2721
rect 1783 -2722 1784 -2721
rect 1787 -2722 1788 -2721
rect 58 -2724 59 -2723
rect 590 -2724 591 -2723
rect 621 -2724 622 -2723
rect 737 -2724 738 -2723
rect 775 -2724 776 -2723
rect 1507 -2724 1508 -2723
rect 65 -2726 66 -2725
rect 1125 -2726 1126 -2725
rect 1129 -2726 1130 -2725
rect 1202 -2726 1203 -2725
rect 1297 -2726 1298 -2725
rect 1360 -2726 1361 -2725
rect 100 -2728 101 -2727
rect 103 -2728 104 -2727
rect 107 -2728 108 -2727
rect 523 -2728 524 -2727
rect 534 -2728 535 -2727
rect 887 -2728 888 -2727
rect 891 -2728 892 -2727
rect 978 -2728 979 -2727
rect 1003 -2728 1004 -2727
rect 1325 -2728 1326 -2727
rect 1328 -2728 1329 -2727
rect 1675 -2728 1676 -2727
rect 100 -2730 101 -2729
rect 156 -2730 157 -2729
rect 198 -2730 199 -2729
rect 208 -2730 209 -2729
rect 289 -2730 290 -2729
rect 373 -2730 374 -2729
rect 401 -2730 402 -2729
rect 422 -2730 423 -2729
rect 425 -2730 426 -2729
rect 604 -2730 605 -2729
rect 660 -2730 661 -2729
rect 891 -2730 892 -2729
rect 919 -2730 920 -2729
rect 1234 -2730 1235 -2729
rect 1297 -2730 1298 -2729
rect 1339 -2730 1340 -2729
rect 1346 -2730 1347 -2729
rect 1451 -2730 1452 -2729
rect 1675 -2730 1676 -2729
rect 1717 -2730 1718 -2729
rect 107 -2732 108 -2731
rect 443 -2732 444 -2731
rect 464 -2732 465 -2731
rect 1181 -2732 1182 -2731
rect 1318 -2732 1319 -2731
rect 1605 -2732 1606 -2731
rect 142 -2734 143 -2733
rect 667 -2734 668 -2733
rect 842 -2734 843 -2733
rect 856 -2734 857 -2733
rect 863 -2734 864 -2733
rect 1206 -2734 1207 -2733
rect 1318 -2734 1319 -2733
rect 1437 -2734 1438 -2733
rect 1605 -2734 1606 -2733
rect 1626 -2734 1627 -2733
rect 149 -2736 150 -2735
rect 156 -2736 157 -2735
rect 201 -2736 202 -2735
rect 261 -2736 262 -2735
rect 292 -2736 293 -2735
rect 513 -2736 514 -2735
rect 534 -2736 535 -2735
rect 744 -2736 745 -2735
rect 849 -2736 850 -2735
rect 1283 -2736 1284 -2735
rect 1325 -2736 1326 -2735
rect 1423 -2736 1424 -2735
rect 1437 -2736 1438 -2735
rect 1549 -2736 1550 -2735
rect 1626 -2736 1627 -2735
rect 1647 -2736 1648 -2735
rect 103 -2738 104 -2737
rect 149 -2738 150 -2737
rect 205 -2738 206 -2737
rect 219 -2738 220 -2737
rect 226 -2738 227 -2737
rect 373 -2738 374 -2737
rect 436 -2738 437 -2737
rect 632 -2738 633 -2737
rect 660 -2738 661 -2737
rect 663 -2738 664 -2737
rect 667 -2738 668 -2737
rect 954 -2738 955 -2737
rect 1003 -2738 1004 -2737
rect 1069 -2738 1070 -2737
rect 1080 -2738 1081 -2737
rect 1241 -2738 1242 -2737
rect 1332 -2738 1333 -2737
rect 1773 -2738 1774 -2737
rect 128 -2740 129 -2739
rect 219 -2740 220 -2739
rect 226 -2740 227 -2739
rect 611 -2740 612 -2739
rect 632 -2740 633 -2739
rect 653 -2740 654 -2739
rect 705 -2740 706 -2739
rect 1332 -2740 1333 -2739
rect 1346 -2740 1347 -2739
rect 1353 -2740 1354 -2739
rect 1549 -2740 1550 -2739
rect 1584 -2740 1585 -2739
rect 1647 -2740 1648 -2739
rect 1682 -2740 1683 -2739
rect 1773 -2740 1774 -2739
rect 1794 -2740 1795 -2739
rect 79 -2742 80 -2741
rect 128 -2742 129 -2741
rect 170 -2742 171 -2741
rect 653 -2742 654 -2741
rect 716 -2742 717 -2741
rect 856 -2742 857 -2741
rect 863 -2742 864 -2741
rect 1213 -2742 1214 -2741
rect 1241 -2742 1242 -2741
rect 1388 -2742 1389 -2741
rect 1584 -2742 1585 -2741
rect 1612 -2742 1613 -2741
rect 1682 -2742 1683 -2741
rect 1724 -2742 1725 -2741
rect 61 -2744 62 -2743
rect 1213 -2744 1214 -2743
rect 1237 -2744 1238 -2743
rect 1612 -2744 1613 -2743
rect 79 -2746 80 -2745
rect 93 -2746 94 -2745
rect 170 -2746 171 -2745
rect 359 -2746 360 -2745
rect 436 -2746 437 -2745
rect 639 -2746 640 -2745
rect 716 -2746 717 -2745
rect 779 -2746 780 -2745
rect 852 -2746 853 -2745
rect 877 -2746 878 -2745
rect 884 -2746 885 -2745
rect 1164 -2746 1165 -2745
rect 1283 -2746 1284 -2745
rect 1724 -2746 1725 -2745
rect 37 -2748 38 -2747
rect 359 -2748 360 -2747
rect 443 -2748 444 -2747
rect 541 -2748 542 -2747
rect 562 -2748 563 -2747
rect 639 -2748 640 -2747
rect 695 -2748 696 -2747
rect 779 -2748 780 -2747
rect 877 -2748 878 -2747
rect 1321 -2748 1322 -2747
rect 1388 -2748 1389 -2747
rect 1430 -2748 1431 -2747
rect 37 -2750 38 -2749
rect 86 -2750 87 -2749
rect 261 -2750 262 -2749
rect 1353 -2750 1354 -2749
rect 9 -2752 10 -2751
rect 86 -2752 87 -2751
rect 303 -2752 304 -2751
rect 859 -2752 860 -2751
rect 884 -2752 885 -2751
rect 1062 -2752 1063 -2751
rect 1080 -2752 1081 -2751
rect 1094 -2752 1095 -2751
rect 1118 -2752 1119 -2751
rect 1661 -2752 1662 -2751
rect 44 -2754 45 -2753
rect 93 -2754 94 -2753
rect 303 -2754 304 -2753
rect 366 -2754 367 -2753
rect 464 -2754 465 -2753
rect 786 -2754 787 -2753
rect 919 -2754 920 -2753
rect 989 -2754 990 -2753
rect 1010 -2754 1011 -2753
rect 1052 -2754 1053 -2753
rect 1087 -2754 1088 -2753
rect 1342 -2754 1343 -2753
rect 1661 -2754 1662 -2753
rect 1752 -2754 1753 -2753
rect 268 -2756 269 -2755
rect 366 -2756 367 -2755
rect 478 -2756 479 -2755
rect 481 -2756 482 -2755
rect 513 -2756 514 -2755
rect 527 -2756 528 -2755
rect 541 -2756 542 -2755
rect 597 -2756 598 -2755
rect 611 -2756 612 -2755
rect 723 -2756 724 -2755
rect 744 -2756 745 -2755
rect 793 -2756 794 -2755
rect 940 -2756 941 -2755
rect 1206 -2756 1207 -2755
rect 1720 -2756 1721 -2755
rect 1752 -2756 1753 -2755
rect 135 -2758 136 -2757
rect 268 -2758 269 -2757
rect 331 -2758 332 -2757
rect 565 -2758 566 -2757
rect 569 -2758 570 -2757
rect 915 -2758 916 -2757
rect 940 -2758 941 -2757
rect 1153 -2758 1154 -2757
rect 1164 -2758 1165 -2757
rect 1199 -2758 1200 -2757
rect 135 -2760 136 -2759
rect 233 -2760 234 -2759
rect 310 -2760 311 -2759
rect 331 -2760 332 -2759
rect 338 -2760 339 -2759
rect 401 -2760 402 -2759
rect 527 -2760 528 -2759
rect 828 -2760 829 -2759
rect 954 -2760 955 -2759
rect 961 -2760 962 -2759
rect 982 -2760 983 -2759
rect 989 -2760 990 -2759
rect 1013 -2760 1014 -2759
rect 1423 -2760 1424 -2759
rect 51 -2762 52 -2761
rect 233 -2762 234 -2761
rect 310 -2762 311 -2761
rect 1010 -2762 1011 -2761
rect 1017 -2762 1018 -2761
rect 1759 -2762 1760 -2761
rect 51 -2764 52 -2763
rect 387 -2764 388 -2763
rect 562 -2764 563 -2763
rect 702 -2764 703 -2763
rect 786 -2764 787 -2763
rect 1045 -2764 1046 -2763
rect 1052 -2764 1053 -2763
rect 1073 -2764 1074 -2763
rect 1094 -2764 1095 -2763
rect 1570 -2764 1571 -2763
rect 1745 -2764 1746 -2763
rect 1759 -2764 1760 -2763
rect 324 -2766 325 -2765
rect 702 -2766 703 -2765
rect 866 -2766 867 -2765
rect 1570 -2766 1571 -2765
rect 324 -2768 325 -2767
rect 352 -2768 353 -2767
rect 355 -2768 356 -2767
rect 835 -2768 836 -2767
rect 961 -2768 962 -2767
rect 1143 -2768 1144 -2767
rect 1150 -2768 1151 -2767
rect 1689 -2768 1690 -2767
rect 338 -2770 339 -2769
rect 457 -2770 458 -2769
rect 569 -2770 570 -2769
rect 625 -2770 626 -2769
rect 695 -2770 696 -2769
rect 730 -2770 731 -2769
rect 821 -2770 822 -2769
rect 835 -2770 836 -2769
rect 982 -2770 983 -2769
rect 1178 -2770 1179 -2769
rect 1199 -2770 1200 -2769
rect 1514 -2770 1515 -2769
rect 1633 -2770 1634 -2769
rect 1689 -2770 1690 -2769
rect 345 -2772 346 -2771
rect 422 -2772 423 -2771
rect 457 -2772 458 -2771
rect 831 -2772 832 -2771
rect 1031 -2772 1032 -2771
rect 1045 -2772 1046 -2771
rect 1073 -2772 1074 -2771
rect 1276 -2772 1277 -2771
rect 1430 -2772 1431 -2771
rect 1745 -2772 1746 -2771
rect 345 -2774 346 -2773
rect 1059 -2774 1060 -2773
rect 1143 -2774 1144 -2773
rect 1248 -2774 1249 -2773
rect 1276 -2774 1277 -2773
rect 1311 -2774 1312 -2773
rect 1514 -2774 1515 -2773
rect 1542 -2774 1543 -2773
rect 1633 -2774 1634 -2773
rect 1654 -2774 1655 -2773
rect 380 -2776 381 -2775
rect 387 -2776 388 -2775
rect 499 -2776 500 -2775
rect 625 -2776 626 -2775
rect 751 -2776 752 -2775
rect 1248 -2776 1249 -2775
rect 1311 -2776 1312 -2775
rect 1458 -2776 1459 -2775
rect 1542 -2776 1543 -2775
rect 1556 -2776 1557 -2775
rect 380 -2778 381 -2777
rect 408 -2778 409 -2777
rect 478 -2778 479 -2777
rect 499 -2778 500 -2777
rect 583 -2778 584 -2777
rect 1374 -2778 1375 -2777
rect 1458 -2778 1459 -2777
rect 1472 -2778 1473 -2777
rect 1556 -2778 1557 -2777
rect 1696 -2778 1697 -2777
rect 408 -2780 409 -2779
rect 506 -2780 507 -2779
rect 583 -2780 584 -2779
rect 723 -2780 724 -2779
rect 807 -2780 808 -2779
rect 821 -2780 822 -2779
rect 996 -2780 997 -2779
rect 1059 -2780 1060 -2779
rect 1129 -2780 1130 -2779
rect 1654 -2780 1655 -2779
rect 1696 -2780 1697 -2779
rect 1731 -2780 1732 -2779
rect 415 -2782 416 -2781
rect 506 -2782 507 -2781
rect 520 -2782 521 -2781
rect 807 -2782 808 -2781
rect 1031 -2782 1032 -2781
rect 1479 -2782 1480 -2781
rect 1500 -2782 1501 -2781
rect 1731 -2782 1732 -2781
rect 415 -2784 416 -2783
rect 429 -2784 430 -2783
rect 520 -2784 521 -2783
rect 576 -2784 577 -2783
rect 590 -2784 591 -2783
rect 1717 -2784 1718 -2783
rect 247 -2786 248 -2785
rect 576 -2786 577 -2785
rect 597 -2786 598 -2785
rect 688 -2786 689 -2785
rect 1150 -2786 1151 -2785
rect 1171 -2786 1172 -2785
rect 1178 -2786 1179 -2785
rect 1563 -2786 1564 -2785
rect 247 -2788 248 -2787
rect 471 -2788 472 -2787
rect 548 -2788 549 -2787
rect 996 -2788 997 -2787
rect 1171 -2788 1172 -2787
rect 1227 -2788 1228 -2787
rect 1374 -2788 1375 -2787
rect 1766 -2788 1767 -2787
rect 177 -2790 178 -2789
rect 548 -2790 549 -2789
rect 607 -2790 608 -2789
rect 793 -2790 794 -2789
rect 947 -2790 948 -2789
rect 1227 -2790 1228 -2789
rect 1402 -2790 1403 -2789
rect 1766 -2790 1767 -2789
rect 121 -2792 122 -2791
rect 177 -2792 178 -2791
rect 296 -2792 297 -2791
rect 688 -2792 689 -2791
rect 1402 -2792 1403 -2791
rect 1591 -2792 1592 -2791
rect 121 -2794 122 -2793
rect 240 -2794 241 -2793
rect 296 -2794 297 -2793
rect 681 -2794 682 -2793
rect 1465 -2794 1466 -2793
rect 1563 -2794 1564 -2793
rect 1591 -2794 1592 -2793
rect 1619 -2794 1620 -2793
rect 212 -2796 213 -2795
rect 240 -2796 241 -2795
rect 317 -2796 318 -2795
rect 429 -2796 430 -2795
rect 471 -2796 472 -2795
rect 485 -2796 486 -2795
rect 618 -2796 619 -2795
rect 730 -2796 731 -2795
rect 1465 -2796 1466 -2795
rect 1486 -2796 1487 -2795
rect 1619 -2796 1620 -2795
rect 1703 -2796 1704 -2795
rect 212 -2798 213 -2797
rect 282 -2798 283 -2797
rect 317 -2798 318 -2797
rect 1185 -2798 1186 -2797
rect 1472 -2798 1473 -2797
rect 1521 -2798 1522 -2797
rect 1703 -2798 1704 -2797
rect 1738 -2798 1739 -2797
rect 254 -2800 255 -2799
rect 282 -2800 283 -2799
rect 485 -2800 486 -2799
rect 555 -2800 556 -2799
rect 618 -2800 619 -2799
rect 751 -2800 752 -2799
rect 912 -2800 913 -2799
rect 1521 -2800 1522 -2799
rect 163 -2802 164 -2801
rect 555 -2802 556 -2801
rect 635 -2802 636 -2801
rect 947 -2802 948 -2801
rect 975 -2802 976 -2801
rect 1486 -2802 1487 -2801
rect 163 -2804 164 -2803
rect 191 -2804 192 -2803
rect 254 -2804 255 -2803
rect 870 -2804 871 -2803
rect 912 -2804 913 -2803
rect 926 -2804 927 -2803
rect 975 -2804 976 -2803
rect 1038 -2804 1039 -2803
rect 1185 -2804 1186 -2803
rect 1262 -2804 1263 -2803
rect 1381 -2804 1382 -2803
rect 1738 -2804 1739 -2803
rect 191 -2806 192 -2805
rect 492 -2806 493 -2805
rect 681 -2806 682 -2805
rect 765 -2806 766 -2805
rect 926 -2806 927 -2805
rect 968 -2806 969 -2805
rect 1038 -2806 1039 -2805
rect 1115 -2806 1116 -2805
rect 1255 -2806 1256 -2805
rect 1262 -2806 1263 -2805
rect 1381 -2806 1382 -2805
rect 1444 -2806 1445 -2805
rect 1479 -2806 1480 -2805
rect 1528 -2806 1529 -2805
rect 450 -2808 451 -2807
rect 492 -2808 493 -2807
rect 709 -2808 710 -2807
rect 765 -2808 766 -2807
rect 968 -2808 969 -2807
rect 1024 -2808 1025 -2807
rect 1087 -2808 1088 -2807
rect 1115 -2808 1116 -2807
rect 1255 -2808 1256 -2807
rect 1304 -2808 1305 -2807
rect 1444 -2808 1445 -2807
rect 1640 -2808 1641 -2807
rect 394 -2810 395 -2809
rect 450 -2810 451 -2809
rect 709 -2810 710 -2809
rect 845 -2810 846 -2809
rect 1024 -2810 1025 -2809
rect 1066 -2810 1067 -2809
rect 1304 -2810 1305 -2809
rect 1367 -2810 1368 -2809
rect 1528 -2810 1529 -2809
rect 1577 -2810 1578 -2809
rect 1640 -2810 1641 -2809
rect 1668 -2810 1669 -2809
rect 394 -2812 395 -2811
rect 674 -2812 675 -2811
rect 1066 -2812 1067 -2811
rect 1220 -2812 1221 -2811
rect 1367 -2812 1368 -2811
rect 1395 -2812 1396 -2811
rect 1577 -2812 1578 -2811
rect 1598 -2812 1599 -2811
rect 1668 -2812 1669 -2811
rect 1710 -2812 1711 -2811
rect 674 -2814 675 -2813
rect 758 -2814 759 -2813
rect 1020 -2814 1021 -2813
rect 1395 -2814 1396 -2813
rect 1500 -2814 1501 -2813
rect 1710 -2814 1711 -2813
rect 758 -2816 759 -2815
rect 800 -2816 801 -2815
rect 1020 -2816 1021 -2815
rect 1192 -2816 1193 -2815
rect 1220 -2816 1221 -2815
rect 1269 -2816 1270 -2815
rect 1535 -2816 1536 -2815
rect 1598 -2816 1599 -2815
rect 800 -2818 801 -2817
rect 933 -2818 934 -2817
rect 1136 -2818 1137 -2817
rect 1269 -2818 1270 -2817
rect 1409 -2818 1410 -2817
rect 1535 -2818 1536 -2817
rect 814 -2820 815 -2819
rect 933 -2820 934 -2819
rect 1136 -2820 1137 -2819
rect 1244 -2820 1245 -2819
rect 1409 -2820 1410 -2819
rect 1416 -2820 1417 -2819
rect 814 -2822 815 -2821
rect 1713 -2822 1714 -2821
rect 905 -2824 906 -2823
rect 1416 -2824 1417 -2823
rect 898 -2826 899 -2825
rect 905 -2826 906 -2825
rect 1157 -2826 1158 -2825
rect 1192 -2826 1193 -2825
rect 733 -2828 734 -2827
rect 898 -2828 899 -2827
rect 1122 -2828 1123 -2827
rect 1157 -2828 1158 -2827
rect 23 -2839 24 -2838
rect 289 -2839 290 -2838
rect 331 -2839 332 -2838
rect 583 -2839 584 -2838
rect 621 -2839 622 -2838
rect 1031 -2839 1032 -2838
rect 1097 -2839 1098 -2838
rect 1668 -2839 1669 -2838
rect 1713 -2839 1714 -2838
rect 1759 -2839 1760 -2838
rect 44 -2841 45 -2840
rect 558 -2841 559 -2840
rect 656 -2841 657 -2840
rect 1416 -2841 1417 -2840
rect 1433 -2841 1434 -2840
rect 1689 -2841 1690 -2840
rect 1717 -2841 1718 -2840
rect 1773 -2841 1774 -2840
rect 79 -2843 80 -2842
rect 583 -2843 584 -2842
rect 660 -2843 661 -2842
rect 1248 -2843 1249 -2842
rect 1283 -2843 1284 -2842
rect 1675 -2843 1676 -2842
rect 1720 -2843 1721 -2842
rect 1766 -2843 1767 -2842
rect 93 -2845 94 -2844
rect 1248 -2845 1249 -2844
rect 1339 -2845 1340 -2844
rect 1612 -2845 1613 -2844
rect 1654 -2845 1655 -2844
rect 1675 -2845 1676 -2844
rect 1727 -2845 1728 -2844
rect 1752 -2845 1753 -2844
rect 93 -2847 94 -2846
rect 121 -2847 122 -2846
rect 128 -2847 129 -2846
rect 828 -2847 829 -2846
rect 859 -2847 860 -2846
rect 1696 -2847 1697 -2846
rect 96 -2849 97 -2848
rect 705 -2849 706 -2848
rect 712 -2849 713 -2848
rect 786 -2849 787 -2848
rect 824 -2849 825 -2848
rect 1507 -2849 1508 -2848
rect 1598 -2849 1599 -2848
rect 1696 -2849 1697 -2848
rect 100 -2851 101 -2850
rect 618 -2851 619 -2850
rect 681 -2851 682 -2850
rect 996 -2851 997 -2850
rect 1013 -2851 1014 -2850
rect 1388 -2851 1389 -2850
rect 1465 -2851 1466 -2850
rect 1507 -2851 1508 -2850
rect 1591 -2851 1592 -2850
rect 1598 -2851 1599 -2850
rect 1647 -2851 1648 -2850
rect 1654 -2851 1655 -2850
rect 37 -2853 38 -2852
rect 681 -2853 682 -2852
rect 730 -2853 731 -2852
rect 877 -2853 878 -2852
rect 915 -2853 916 -2852
rect 1332 -2853 1333 -2852
rect 1342 -2853 1343 -2852
rect 1563 -2853 1564 -2852
rect 1640 -2853 1641 -2852
rect 1647 -2853 1648 -2852
rect 51 -2855 52 -2854
rect 100 -2855 101 -2854
rect 107 -2855 108 -2854
rect 856 -2855 857 -2854
rect 870 -2855 871 -2854
rect 905 -2855 906 -2854
rect 947 -2855 948 -2854
rect 1017 -2855 1018 -2854
rect 1024 -2855 1025 -2854
rect 1129 -2855 1130 -2854
rect 1150 -2855 1151 -2854
rect 1283 -2855 1284 -2854
rect 1353 -2855 1354 -2854
rect 1682 -2855 1683 -2854
rect 51 -2857 52 -2856
rect 72 -2857 73 -2856
rect 107 -2857 108 -2856
rect 1157 -2857 1158 -2856
rect 1178 -2857 1179 -2856
rect 1703 -2857 1704 -2856
rect 72 -2859 73 -2858
rect 324 -2859 325 -2858
rect 359 -2859 360 -2858
rect 709 -2859 710 -2858
rect 765 -2859 766 -2858
rect 856 -2859 857 -2858
rect 877 -2859 878 -2858
rect 1010 -2859 1011 -2858
rect 1024 -2859 1025 -2858
rect 1514 -2859 1515 -2858
rect 1661 -2859 1662 -2858
rect 1682 -2859 1683 -2858
rect 1703 -2859 1704 -2858
rect 1724 -2859 1725 -2858
rect 121 -2861 122 -2860
rect 191 -2861 192 -2860
rect 226 -2861 227 -2860
rect 352 -2861 353 -2860
rect 366 -2861 367 -2860
rect 481 -2861 482 -2860
rect 520 -2861 521 -2860
rect 1055 -2861 1056 -2860
rect 1101 -2861 1102 -2860
rect 1150 -2861 1151 -2860
rect 1199 -2861 1200 -2860
rect 1276 -2861 1277 -2860
rect 1353 -2861 1354 -2860
rect 1374 -2861 1375 -2860
rect 1381 -2861 1382 -2860
rect 1416 -2861 1417 -2860
rect 1444 -2861 1445 -2860
rect 1591 -2861 1592 -2860
rect 1640 -2861 1641 -2860
rect 1661 -2861 1662 -2860
rect 65 -2863 66 -2862
rect 520 -2863 521 -2862
rect 555 -2863 556 -2862
rect 1045 -2863 1046 -2862
rect 1066 -2863 1067 -2862
rect 1101 -2863 1102 -2862
rect 1115 -2863 1116 -2862
rect 1164 -2863 1165 -2862
rect 1202 -2863 1203 -2862
rect 1451 -2863 1452 -2862
rect 1514 -2863 1515 -2862
rect 1528 -2863 1529 -2862
rect 65 -2865 66 -2864
rect 261 -2865 262 -2864
rect 275 -2865 276 -2864
rect 355 -2865 356 -2864
rect 366 -2865 367 -2864
rect 380 -2865 381 -2864
rect 429 -2865 430 -2864
rect 432 -2865 433 -2864
rect 464 -2865 465 -2864
rect 1178 -2865 1179 -2864
rect 1227 -2865 1228 -2864
rect 1689 -2865 1690 -2864
rect 128 -2867 129 -2866
rect 229 -2867 230 -2866
rect 247 -2867 248 -2866
rect 999 -2867 1000 -2866
rect 1066 -2867 1067 -2866
rect 1234 -2867 1235 -2866
rect 1237 -2867 1238 -2866
rect 1500 -2867 1501 -2866
rect 135 -2869 136 -2868
rect 411 -2869 412 -2868
rect 429 -2869 430 -2868
rect 541 -2869 542 -2868
rect 555 -2869 556 -2868
rect 646 -2869 647 -2868
rect 674 -2869 675 -2868
rect 1115 -2869 1116 -2868
rect 1125 -2869 1126 -2868
rect 1542 -2869 1543 -2868
rect 142 -2871 143 -2870
rect 702 -2871 703 -2870
rect 737 -2871 738 -2870
rect 765 -2871 766 -2870
rect 779 -2871 780 -2870
rect 947 -2871 948 -2870
rect 968 -2871 969 -2870
rect 1045 -2871 1046 -2870
rect 1136 -2871 1137 -2870
rect 1276 -2871 1277 -2870
rect 1311 -2871 1312 -2870
rect 1451 -2871 1452 -2870
rect 1500 -2871 1501 -2870
rect 1521 -2871 1522 -2870
rect 1535 -2871 1536 -2870
rect 1542 -2871 1543 -2870
rect 86 -2873 87 -2872
rect 142 -2873 143 -2872
rect 145 -2873 146 -2872
rect 1612 -2873 1613 -2872
rect 86 -2875 87 -2874
rect 114 -2875 115 -2874
rect 170 -2875 171 -2874
rect 586 -2875 587 -2874
rect 604 -2875 605 -2874
rect 1129 -2875 1130 -2874
rect 1164 -2875 1165 -2874
rect 1171 -2875 1172 -2874
rect 1227 -2875 1228 -2874
rect 1731 -2875 1732 -2874
rect 58 -2877 59 -2876
rect 114 -2877 115 -2876
rect 156 -2877 157 -2876
rect 170 -2877 171 -2876
rect 226 -2877 227 -2876
rect 467 -2877 468 -2876
rect 562 -2877 563 -2876
rect 1563 -2877 1564 -2876
rect 58 -2879 59 -2878
rect 782 -2879 783 -2878
rect 786 -2879 787 -2878
rect 1027 -2879 1028 -2878
rect 1171 -2879 1172 -2878
rect 1395 -2879 1396 -2878
rect 1437 -2879 1438 -2878
rect 1528 -2879 1529 -2878
rect 156 -2881 157 -2880
rect 184 -2881 185 -2880
rect 240 -2881 241 -2880
rect 247 -2881 248 -2880
rect 254 -2881 255 -2880
rect 866 -2881 867 -2880
rect 971 -2881 972 -2880
rect 1297 -2881 1298 -2880
rect 1311 -2881 1312 -2880
rect 1710 -2881 1711 -2880
rect 149 -2883 150 -2882
rect 254 -2883 255 -2882
rect 261 -2883 262 -2882
rect 373 -2883 374 -2882
rect 380 -2883 381 -2882
rect 565 -2883 566 -2882
rect 576 -2883 577 -2882
rect 618 -2883 619 -2882
rect 646 -2883 647 -2882
rect 807 -2883 808 -2882
rect 821 -2883 822 -2882
rect 870 -2883 871 -2882
rect 982 -2883 983 -2882
rect 1136 -2883 1137 -2882
rect 1234 -2883 1235 -2882
rect 1304 -2883 1305 -2882
rect 1318 -2883 1319 -2882
rect 1395 -2883 1396 -2882
rect 1423 -2883 1424 -2882
rect 1437 -2883 1438 -2882
rect 1444 -2883 1445 -2882
rect 1577 -2883 1578 -2882
rect 149 -2885 150 -2884
rect 338 -2885 339 -2884
rect 373 -2885 374 -2884
rect 387 -2885 388 -2884
rect 394 -2885 395 -2884
rect 464 -2885 465 -2884
rect 562 -2885 563 -2884
rect 569 -2885 570 -2884
rect 576 -2885 577 -2884
rect 849 -2885 850 -2884
rect 898 -2885 899 -2884
rect 982 -2885 983 -2884
rect 989 -2885 990 -2884
rect 1010 -2885 1011 -2884
rect 1255 -2885 1256 -2884
rect 1297 -2885 1298 -2884
rect 1318 -2885 1319 -2884
rect 1738 -2885 1739 -2884
rect 184 -2887 185 -2886
rect 625 -2887 626 -2886
rect 667 -2887 668 -2886
rect 898 -2887 899 -2886
rect 933 -2887 934 -2886
rect 1423 -2887 1424 -2886
rect 1479 -2887 1480 -2886
rect 1521 -2887 1522 -2886
rect 1570 -2887 1571 -2886
rect 1577 -2887 1578 -2886
rect 233 -2889 234 -2888
rect 387 -2889 388 -2888
rect 394 -2889 395 -2888
rect 422 -2889 423 -2888
rect 432 -2889 433 -2888
rect 541 -2889 542 -2888
rect 590 -2889 591 -2888
rect 604 -2889 605 -2888
rect 625 -2889 626 -2888
rect 873 -2889 874 -2888
rect 1143 -2889 1144 -2888
rect 1255 -2889 1256 -2888
rect 1262 -2889 1263 -2888
rect 1388 -2889 1389 -2888
rect 1458 -2889 1459 -2888
rect 1479 -2889 1480 -2888
rect 1486 -2889 1487 -2888
rect 1535 -2889 1536 -2888
rect 1570 -2889 1571 -2888
rect 1584 -2889 1585 -2888
rect 233 -2891 234 -2890
rect 1122 -2891 1123 -2890
rect 1185 -2891 1186 -2890
rect 1262 -2891 1263 -2890
rect 1269 -2891 1270 -2890
rect 1304 -2891 1305 -2890
rect 1325 -2891 1326 -2890
rect 1381 -2891 1382 -2890
rect 1409 -2891 1410 -2890
rect 1584 -2891 1585 -2890
rect 240 -2893 241 -2892
rect 268 -2893 269 -2892
rect 275 -2893 276 -2892
rect 814 -2893 815 -2892
rect 828 -2893 829 -2892
rect 835 -2893 836 -2892
rect 849 -2893 850 -2892
rect 1360 -2893 1361 -2892
rect 1367 -2893 1368 -2892
rect 1374 -2893 1375 -2892
rect 1472 -2893 1473 -2892
rect 1486 -2893 1487 -2892
rect 268 -2895 269 -2894
rect 639 -2895 640 -2894
rect 653 -2895 654 -2894
rect 1143 -2895 1144 -2894
rect 1185 -2895 1186 -2894
rect 1192 -2895 1193 -2894
rect 1213 -2895 1214 -2894
rect 1360 -2895 1361 -2894
rect 1472 -2895 1473 -2894
rect 1493 -2895 1494 -2894
rect 282 -2897 283 -2896
rect 359 -2897 360 -2896
rect 415 -2897 416 -2896
rect 422 -2897 423 -2896
rect 439 -2897 440 -2896
rect 1409 -2897 1410 -2896
rect 198 -2899 199 -2898
rect 415 -2899 416 -2898
rect 527 -2899 528 -2898
rect 569 -2899 570 -2898
rect 590 -2899 591 -2898
rect 716 -2899 717 -2898
rect 737 -2899 738 -2898
rect 940 -2899 941 -2898
rect 1059 -2899 1060 -2898
rect 1192 -2899 1193 -2898
rect 1220 -2899 1221 -2898
rect 1269 -2899 1270 -2898
rect 1325 -2899 1326 -2898
rect 1346 -2899 1347 -2898
rect 1356 -2899 1357 -2898
rect 1619 -2899 1620 -2898
rect 110 -2901 111 -2900
rect 716 -2901 717 -2900
rect 751 -2901 752 -2900
rect 933 -2901 934 -2900
rect 1052 -2901 1053 -2900
rect 1059 -2901 1060 -2900
rect 1069 -2901 1070 -2900
rect 1458 -2901 1459 -2900
rect 198 -2903 199 -2902
rect 205 -2903 206 -2902
rect 212 -2903 213 -2902
rect 282 -2903 283 -2902
rect 289 -2903 290 -2902
rect 310 -2903 311 -2902
rect 317 -2903 318 -2902
rect 989 -2903 990 -2902
rect 1052 -2903 1053 -2902
rect 1556 -2903 1557 -2902
rect 163 -2905 164 -2904
rect 205 -2905 206 -2904
rect 212 -2905 213 -2904
rect 1286 -2905 1287 -2904
rect 1290 -2905 1291 -2904
rect 1346 -2905 1347 -2904
rect 1402 -2905 1403 -2904
rect 1556 -2905 1557 -2904
rect 163 -2907 164 -2906
rect 1157 -2907 1158 -2906
rect 1206 -2907 1207 -2906
rect 1619 -2907 1620 -2906
rect 303 -2909 304 -2908
rect 317 -2909 318 -2908
rect 324 -2909 325 -2908
rect 401 -2909 402 -2908
rect 506 -2909 507 -2908
rect 527 -2909 528 -2908
rect 653 -2909 654 -2908
rect 1668 -2909 1669 -2908
rect 208 -2911 209 -2910
rect 303 -2911 304 -2910
rect 310 -2911 311 -2910
rect 457 -2911 458 -2910
rect 506 -2911 507 -2910
rect 597 -2911 598 -2910
rect 663 -2911 664 -2910
rect 814 -2911 815 -2910
rect 835 -2911 836 -2910
rect 1087 -2911 1088 -2910
rect 1094 -2911 1095 -2910
rect 1493 -2911 1494 -2910
rect 219 -2913 220 -2912
rect 457 -2913 458 -2912
rect 667 -2913 668 -2912
rect 1031 -2913 1032 -2912
rect 1073 -2913 1074 -2912
rect 1290 -2913 1291 -2912
rect 1402 -2913 1403 -2912
rect 1745 -2913 1746 -2912
rect 219 -2915 220 -2914
rect 968 -2915 969 -2914
rect 1038 -2915 1039 -2914
rect 1073 -2915 1074 -2914
rect 1080 -2915 1081 -2914
rect 1122 -2915 1123 -2914
rect 1241 -2915 1242 -2914
rect 1367 -2915 1368 -2914
rect 338 -2917 339 -2916
rect 408 -2917 409 -2916
rect 436 -2917 437 -2916
rect 597 -2917 598 -2916
rect 674 -2917 675 -2916
rect 852 -2917 853 -2916
rect 891 -2917 892 -2916
rect 1213 -2917 1214 -2916
rect 191 -2919 192 -2918
rect 436 -2919 437 -2918
rect 688 -2919 689 -2918
rect 751 -2919 752 -2918
rect 800 -2919 801 -2918
rect 905 -2919 906 -2918
rect 961 -2919 962 -2918
rect 1206 -2919 1207 -2918
rect 331 -2921 332 -2920
rect 852 -2921 853 -2920
rect 926 -2921 927 -2920
rect 961 -2921 962 -2920
rect 975 -2921 976 -2920
rect 1038 -2921 1039 -2920
rect 1108 -2921 1109 -2920
rect 1220 -2921 1221 -2920
rect 345 -2923 346 -2922
rect 639 -2923 640 -2922
rect 688 -2923 689 -2922
rect 1020 -2923 1021 -2922
rect 1108 -2923 1109 -2922
rect 1430 -2923 1431 -2922
rect 177 -2925 178 -2924
rect 345 -2925 346 -2924
rect 401 -2925 402 -2924
rect 450 -2925 451 -2924
rect 695 -2925 696 -2924
rect 800 -2925 801 -2924
rect 807 -2925 808 -2924
rect 884 -2925 885 -2924
rect 919 -2925 920 -2924
rect 975 -2925 976 -2924
rect 1003 -2925 1004 -2924
rect 1080 -2925 1081 -2924
rect 1430 -2925 1431 -2924
rect 1605 -2925 1606 -2924
rect 177 -2927 178 -2926
rect 485 -2927 486 -2926
rect 534 -2927 535 -2926
rect 695 -2927 696 -2926
rect 723 -2927 724 -2926
rect 1087 -2927 1088 -2926
rect 1605 -2927 1606 -2926
rect 1626 -2927 1627 -2926
rect 443 -2929 444 -2928
rect 450 -2929 451 -2928
rect 485 -2929 486 -2928
rect 537 -2929 538 -2928
rect 723 -2929 724 -2928
rect 758 -2929 759 -2928
rect 793 -2929 794 -2928
rect 919 -2929 920 -2928
rect 926 -2929 927 -2928
rect 1202 -2929 1203 -2928
rect 1626 -2929 1627 -2928
rect 1633 -2929 1634 -2928
rect 443 -2931 444 -2930
rect 513 -2931 514 -2930
rect 733 -2931 734 -2930
rect 1633 -2931 1634 -2930
rect 478 -2933 479 -2932
rect 513 -2933 514 -2932
rect 744 -2933 745 -2932
rect 793 -2933 794 -2932
rect 842 -2933 843 -2932
rect 891 -2933 892 -2932
rect 478 -2935 479 -2934
rect 943 -2935 944 -2934
rect 492 -2937 493 -2936
rect 534 -2937 535 -2936
rect 611 -2937 612 -2936
rect 744 -2937 745 -2936
rect 758 -2937 759 -2936
rect 772 -2937 773 -2936
rect 863 -2937 864 -2936
rect 1003 -2937 1004 -2936
rect 492 -2939 493 -2938
rect 660 -2939 661 -2938
rect 663 -2939 664 -2938
rect 842 -2939 843 -2938
rect 863 -2939 864 -2938
rect 1241 -2939 1242 -2938
rect 548 -2941 549 -2940
rect 772 -2941 773 -2940
rect 884 -2941 885 -2940
rect 912 -2941 913 -2940
rect 82 -2943 83 -2942
rect 548 -2943 549 -2942
rect 611 -2943 612 -2942
rect 632 -2943 633 -2942
rect 912 -2943 913 -2942
rect 1465 -2943 1466 -2942
rect 296 -2945 297 -2944
rect 632 -2945 633 -2944
rect 166 -2947 167 -2946
rect 296 -2947 297 -2946
rect 30 -2958 31 -2957
rect 93 -2958 94 -2957
rect 100 -2958 101 -2957
rect 436 -2958 437 -2957
rect 439 -2958 440 -2957
rect 814 -2958 815 -2957
rect 821 -2958 822 -2957
rect 856 -2958 857 -2957
rect 863 -2958 864 -2957
rect 1584 -2958 1585 -2957
rect 1640 -2958 1641 -2957
rect 1696 -2958 1697 -2957
rect 37 -2960 38 -2959
rect 289 -2960 290 -2959
rect 303 -2960 304 -2959
rect 306 -2960 307 -2959
rect 369 -2960 370 -2959
rect 453 -2960 454 -2959
rect 541 -2960 542 -2959
rect 653 -2960 654 -2959
rect 663 -2960 664 -2959
rect 1213 -2960 1214 -2959
rect 1332 -2960 1333 -2959
rect 1507 -2960 1508 -2959
rect 1577 -2960 1578 -2959
rect 1703 -2960 1704 -2959
rect 44 -2962 45 -2961
rect 394 -2962 395 -2961
rect 450 -2962 451 -2961
rect 541 -2962 542 -2961
rect 548 -2962 549 -2961
rect 814 -2962 815 -2961
rect 842 -2962 843 -2961
rect 1024 -2962 1025 -2961
rect 1027 -2962 1028 -2961
rect 1689 -2962 1690 -2961
rect 23 -2964 24 -2963
rect 450 -2964 451 -2963
rect 499 -2964 500 -2963
rect 548 -2964 549 -2963
rect 611 -2964 612 -2963
rect 653 -2964 654 -2963
rect 674 -2964 675 -2963
rect 978 -2964 979 -2963
rect 1020 -2964 1021 -2963
rect 1220 -2964 1221 -2963
rect 1332 -2964 1333 -2963
rect 1381 -2964 1382 -2963
rect 1458 -2964 1459 -2963
rect 1640 -2964 1641 -2963
rect 72 -2966 73 -2965
rect 411 -2966 412 -2965
rect 499 -2966 500 -2965
rect 688 -2966 689 -2965
rect 740 -2966 741 -2965
rect 1143 -2966 1144 -2965
rect 1171 -2966 1172 -2965
rect 1381 -2966 1382 -2965
rect 1458 -2966 1459 -2965
rect 1465 -2966 1466 -2965
rect 1577 -2966 1578 -2965
rect 1605 -2966 1606 -2965
rect 51 -2968 52 -2967
rect 72 -2968 73 -2967
rect 79 -2968 80 -2967
rect 457 -2968 458 -2967
rect 569 -2968 570 -2967
rect 611 -2968 612 -2967
rect 618 -2968 619 -2967
rect 842 -2968 843 -2967
rect 849 -2968 850 -2967
rect 1115 -2968 1116 -2967
rect 1150 -2968 1151 -2967
rect 1171 -2968 1172 -2967
rect 1199 -2968 1200 -2967
rect 1528 -2968 1529 -2967
rect 1605 -2968 1606 -2967
rect 1647 -2968 1648 -2967
rect 51 -2970 52 -2969
rect 212 -2970 213 -2969
rect 219 -2970 220 -2969
rect 996 -2970 997 -2969
rect 1010 -2970 1011 -2969
rect 1143 -2970 1144 -2969
rect 1199 -2970 1200 -2969
rect 1241 -2970 1242 -2969
rect 1339 -2970 1340 -2969
rect 1584 -2970 1585 -2969
rect 1647 -2970 1648 -2969
rect 1682 -2970 1683 -2969
rect 65 -2972 66 -2971
rect 219 -2972 220 -2971
rect 261 -2972 262 -2971
rect 394 -2972 395 -2971
rect 408 -2972 409 -2971
rect 457 -2972 458 -2971
rect 492 -2972 493 -2971
rect 569 -2972 570 -2971
rect 604 -2972 605 -2971
rect 618 -2972 619 -2971
rect 674 -2972 675 -2971
rect 793 -2972 794 -2971
rect 835 -2972 836 -2971
rect 1150 -2972 1151 -2971
rect 1164 -2972 1165 -2971
rect 1241 -2972 1242 -2971
rect 1339 -2972 1340 -2971
rect 1388 -2972 1389 -2971
rect 1465 -2972 1466 -2971
rect 1486 -2972 1487 -2971
rect 65 -2974 66 -2973
rect 208 -2974 209 -2973
rect 261 -2974 262 -2973
rect 513 -2974 514 -2973
rect 604 -2974 605 -2973
rect 758 -2974 759 -2973
rect 782 -2974 783 -2973
rect 1535 -2974 1536 -2973
rect 82 -2976 83 -2975
rect 1178 -2976 1179 -2975
rect 1213 -2976 1214 -2975
rect 1255 -2976 1256 -2975
rect 1297 -2976 1298 -2975
rect 1388 -2976 1389 -2975
rect 1486 -2976 1487 -2975
rect 1493 -2976 1494 -2975
rect 1535 -2976 1536 -2975
rect 1563 -2976 1564 -2975
rect 93 -2978 94 -2977
rect 562 -2978 563 -2977
rect 793 -2978 794 -2977
rect 926 -2978 927 -2977
rect 943 -2978 944 -2977
rect 1416 -2978 1417 -2977
rect 1430 -2978 1431 -2977
rect 1563 -2978 1564 -2977
rect 79 -2980 80 -2979
rect 1416 -2980 1417 -2979
rect 1430 -2980 1431 -2979
rect 1668 -2980 1669 -2979
rect 100 -2982 101 -2981
rect 660 -2982 661 -2981
rect 835 -2982 836 -2981
rect 989 -2982 990 -2981
rect 996 -2982 997 -2981
rect 1038 -2982 1039 -2981
rect 1052 -2982 1053 -2981
rect 1059 -2982 1060 -2981
rect 1094 -2982 1095 -2981
rect 1318 -2982 1319 -2981
rect 1493 -2982 1494 -2981
rect 1514 -2982 1515 -2981
rect 107 -2984 108 -2983
rect 1024 -2984 1025 -2983
rect 1031 -2984 1032 -2983
rect 1591 -2984 1592 -2983
rect 107 -2986 108 -2985
rect 443 -2986 444 -2985
rect 562 -2986 563 -2985
rect 866 -2986 867 -2985
rect 901 -2986 902 -2985
rect 1423 -2986 1424 -2985
rect 1514 -2986 1515 -2985
rect 1549 -2986 1550 -2985
rect 1591 -2986 1592 -2985
rect 1633 -2986 1634 -2985
rect 110 -2988 111 -2987
rect 254 -2988 255 -2987
rect 268 -2988 269 -2987
rect 1097 -2988 1098 -2987
rect 1115 -2988 1116 -2987
rect 1129 -2988 1130 -2987
rect 1136 -2988 1137 -2987
rect 1178 -2988 1179 -2987
rect 1202 -2988 1203 -2987
rect 1633 -2988 1634 -2987
rect 121 -2990 122 -2989
rect 621 -2990 622 -2989
rect 660 -2990 661 -2989
rect 730 -2990 731 -2989
rect 849 -2990 850 -2989
rect 884 -2990 885 -2989
rect 926 -2990 927 -2989
rect 947 -2990 948 -2989
rect 982 -2990 983 -2989
rect 1038 -2990 1039 -2989
rect 1045 -2990 1046 -2989
rect 1129 -2990 1130 -2989
rect 1136 -2990 1137 -2989
rect 1360 -2990 1361 -2989
rect 1423 -2990 1424 -2989
rect 1675 -2990 1676 -2989
rect 82 -2992 83 -2991
rect 1045 -2992 1046 -2991
rect 1055 -2992 1056 -2991
rect 1521 -2992 1522 -2991
rect 1549 -2992 1550 -2991
rect 1570 -2992 1571 -2991
rect 121 -2994 122 -2993
rect 359 -2994 360 -2993
rect 408 -2994 409 -2993
rect 415 -2994 416 -2993
rect 443 -2994 444 -2993
rect 667 -2994 668 -2993
rect 852 -2994 853 -2993
rect 919 -2994 920 -2993
rect 947 -2994 948 -2993
rect 954 -2994 955 -2993
rect 989 -2994 990 -2993
rect 1073 -2994 1074 -2993
rect 1122 -2994 1123 -2993
rect 1164 -2994 1165 -2993
rect 1220 -2994 1221 -2993
rect 1262 -2994 1263 -2993
rect 1297 -2994 1298 -2993
rect 1353 -2994 1354 -2993
rect 1521 -2994 1522 -2993
rect 1556 -2994 1557 -2993
rect 1570 -2994 1571 -2993
rect 1598 -2994 1599 -2993
rect 89 -2996 90 -2995
rect 1122 -2996 1123 -2995
rect 1255 -2996 1256 -2995
rect 1290 -2996 1291 -2995
rect 1318 -2996 1319 -2995
rect 1367 -2996 1368 -2995
rect 1598 -2996 1599 -2995
rect 1626 -2996 1627 -2995
rect 142 -2998 143 -2997
rect 982 -2998 983 -2997
rect 1010 -2998 1011 -2997
rect 1227 -2998 1228 -2997
rect 1262 -2998 1263 -2997
rect 1311 -2998 1312 -2997
rect 1367 -2998 1368 -2997
rect 1395 -2998 1396 -2997
rect 1626 -2998 1627 -2997
rect 1661 -2998 1662 -2997
rect 145 -3000 146 -2999
rect 583 -3000 584 -2999
rect 632 -3000 633 -2999
rect 730 -3000 731 -2999
rect 856 -3000 857 -2999
rect 870 -3000 871 -2999
rect 877 -3000 878 -2999
rect 919 -3000 920 -2999
rect 954 -3000 955 -2999
rect 961 -3000 962 -2999
rect 968 -3000 969 -2999
rect 1073 -3000 1074 -2999
rect 1227 -3000 1228 -2999
rect 1346 -3000 1347 -2999
rect 156 -3002 157 -3001
rect 254 -3002 255 -3001
rect 268 -3002 269 -3001
rect 380 -3002 381 -3001
rect 415 -3002 416 -3001
rect 422 -3002 423 -3001
rect 506 -3002 507 -3001
rect 1360 -3002 1361 -3001
rect 156 -3004 157 -3003
rect 786 -3004 787 -3003
rect 880 -3004 881 -3003
rect 1353 -3004 1354 -3003
rect 163 -3006 164 -3005
rect 933 -3006 934 -3005
rect 961 -3006 962 -3005
rect 1335 -3006 1336 -3005
rect 1346 -3006 1347 -3005
rect 1706 -3006 1707 -3005
rect 86 -3008 87 -3007
rect 163 -3008 164 -3007
rect 170 -3008 171 -3007
rect 226 -3008 227 -3007
rect 282 -3008 283 -3007
rect 380 -3008 381 -3007
rect 401 -3008 402 -3007
rect 506 -3008 507 -3007
rect 583 -3008 584 -3007
rect 940 -3008 941 -3007
rect 968 -3008 969 -3007
rect 975 -3008 976 -3007
rect 1017 -3008 1018 -3007
rect 1031 -3008 1032 -3007
rect 1034 -3008 1035 -3007
rect 1612 -3008 1613 -3007
rect 86 -3010 87 -3009
rect 1619 -3010 1620 -3009
rect 128 -3012 129 -3011
rect 226 -3012 227 -3011
rect 275 -3012 276 -3011
rect 282 -3012 283 -3011
rect 289 -3012 290 -3011
rect 576 -3012 577 -3011
rect 632 -3012 633 -3011
rect 863 -3012 864 -3011
rect 884 -3012 885 -3011
rect 1108 -3012 1109 -3011
rect 1234 -3012 1235 -3011
rect 1311 -3012 1312 -3011
rect 1612 -3012 1613 -3011
rect 1654 -3012 1655 -3011
rect 58 -3014 59 -3013
rect 576 -3014 577 -3013
rect 639 -3014 640 -3013
rect 667 -3014 668 -3013
rect 702 -3014 703 -3013
rect 877 -3014 878 -3013
rect 898 -3014 899 -3013
rect 933 -3014 934 -3013
rect 1059 -3014 1060 -3013
rect 1087 -3014 1088 -3013
rect 1108 -3014 1109 -3013
rect 1206 -3014 1207 -3013
rect 1234 -3014 1235 -3013
rect 1276 -3014 1277 -3013
rect 58 -3016 59 -3015
rect 135 -3016 136 -3015
rect 138 -3016 139 -3015
rect 275 -3016 276 -3015
rect 303 -3016 304 -3015
rect 478 -3016 479 -3015
rect 513 -3016 514 -3015
rect 1017 -3016 1018 -3015
rect 1192 -3016 1193 -3015
rect 1654 -3016 1655 -3015
rect 128 -3018 129 -3017
rect 695 -3018 696 -3017
rect 702 -3018 703 -3017
rect 723 -3018 724 -3017
rect 789 -3018 790 -3017
rect 940 -3018 941 -3017
rect 1185 -3018 1186 -3017
rect 1192 -3018 1193 -3017
rect 1206 -3018 1207 -3017
rect 1248 -3018 1249 -3017
rect 170 -3020 171 -3019
rect 191 -3020 192 -3019
rect 205 -3020 206 -3019
rect 296 -3020 297 -3019
rect 317 -3020 318 -3019
rect 422 -3020 423 -3019
rect 478 -3020 479 -3019
rect 555 -3020 556 -3019
rect 639 -3020 640 -3019
rect 646 -3020 647 -3019
rect 656 -3020 657 -3019
rect 1290 -3020 1291 -3019
rect 61 -3022 62 -3021
rect 296 -3022 297 -3021
rect 306 -3022 307 -3021
rect 555 -3022 556 -3021
rect 646 -3022 647 -3021
rect 1101 -3022 1102 -3021
rect 1248 -3022 1249 -3021
rect 1283 -3022 1284 -3021
rect 177 -3024 178 -3023
rect 691 -3024 692 -3023
rect 709 -3024 710 -3023
rect 870 -3024 871 -3023
rect 898 -3024 899 -3023
rect 1066 -3024 1067 -3023
rect 1283 -3024 1284 -3023
rect 1325 -3024 1326 -3023
rect 177 -3026 178 -3025
rect 373 -3026 374 -3025
rect 401 -3026 402 -3025
rect 429 -3026 430 -3025
rect 681 -3026 682 -3025
rect 1276 -3026 1277 -3025
rect 1325 -3026 1326 -3025
rect 1374 -3026 1375 -3025
rect 114 -3028 115 -3027
rect 429 -3028 430 -3027
rect 464 -3028 465 -3027
rect 681 -3028 682 -3027
rect 688 -3028 689 -3027
rect 1101 -3028 1102 -3027
rect 1374 -3028 1375 -3027
rect 1402 -3028 1403 -3027
rect 149 -3030 150 -3029
rect 464 -3030 465 -3029
rect 709 -3030 710 -3029
rect 751 -3030 752 -3029
rect 912 -3030 913 -3029
rect 1556 -3030 1557 -3029
rect 149 -3032 150 -3031
rect 1157 -3032 1158 -3031
rect 1304 -3032 1305 -3031
rect 1402 -3032 1403 -3031
rect 187 -3034 188 -3033
rect 1528 -3034 1529 -3033
rect 191 -3036 192 -3035
rect 198 -3036 199 -3035
rect 205 -3036 206 -3035
rect 387 -3036 388 -3035
rect 716 -3036 717 -3035
rect 1157 -3036 1158 -3035
rect 1269 -3036 1270 -3035
rect 1304 -3036 1305 -3035
rect 310 -3038 311 -3037
rect 317 -3038 318 -3037
rect 338 -3038 339 -3037
rect 373 -3038 374 -3037
rect 387 -3038 388 -3037
rect 527 -3038 528 -3037
rect 716 -3038 717 -3037
rect 744 -3038 745 -3037
rect 751 -3038 752 -3037
rect 772 -3038 773 -3037
rect 1003 -3038 1004 -3037
rect 1185 -3038 1186 -3037
rect 1269 -3038 1270 -3037
rect 1437 -3038 1438 -3037
rect 184 -3040 185 -3039
rect 744 -3040 745 -3039
rect 1066 -3040 1067 -3039
rect 1080 -3040 1081 -3039
rect 184 -3042 185 -3041
rect 800 -3042 801 -3041
rect 1080 -3042 1081 -3041
rect 1409 -3042 1410 -3041
rect 310 -3044 311 -3043
rect 625 -3044 626 -3043
rect 723 -3044 724 -3043
rect 758 -3044 759 -3043
rect 800 -3044 801 -3043
rect 1619 -3044 1620 -3043
rect 324 -3046 325 -3045
rect 338 -3046 339 -3045
rect 345 -3046 346 -3045
rect 625 -3046 626 -3045
rect 1409 -3046 1410 -3045
rect 1451 -3046 1452 -3045
rect 324 -3048 325 -3047
rect 331 -3048 332 -3047
rect 345 -3048 346 -3047
rect 695 -3048 696 -3047
rect 786 -3048 787 -3047
rect 1451 -3048 1452 -3047
rect 331 -3050 332 -3049
rect 366 -3050 367 -3049
rect 485 -3050 486 -3049
rect 1437 -3050 1438 -3049
rect 114 -3052 115 -3051
rect 366 -3052 367 -3051
rect 485 -3052 486 -3051
rect 590 -3052 591 -3051
rect 352 -3054 353 -3053
rect 492 -3054 493 -3053
rect 520 -3054 521 -3053
rect 772 -3054 773 -3053
rect 152 -3056 153 -3055
rect 352 -3056 353 -3055
rect 359 -3056 360 -3055
rect 537 -3056 538 -3055
rect 590 -3056 591 -3055
rect 915 -3056 916 -3055
rect 471 -3058 472 -3057
rect 520 -3058 521 -3057
rect 527 -3058 528 -3057
rect 765 -3058 766 -3057
rect 915 -3058 916 -3057
rect 1479 -3058 1480 -3057
rect 471 -3060 472 -3059
rect 737 -3060 738 -3059
rect 765 -3060 766 -3059
rect 807 -3060 808 -3059
rect 1479 -3060 1480 -3059
rect 1500 -3060 1501 -3059
rect 534 -3062 535 -3061
rect 1003 -3062 1004 -3061
rect 1500 -3062 1501 -3061
rect 1542 -3062 1543 -3061
rect 233 -3064 234 -3063
rect 534 -3064 535 -3063
rect 737 -3064 738 -3063
rect 1395 -3064 1396 -3063
rect 1444 -3064 1445 -3063
rect 1542 -3064 1543 -3063
rect 233 -3066 234 -3065
rect 240 -3066 241 -3065
rect 807 -3066 808 -3065
rect 828 -3066 829 -3065
rect 1444 -3066 1445 -3065
rect 1472 -3066 1473 -3065
rect 240 -3068 241 -3067
rect 247 -3068 248 -3067
rect 828 -3068 829 -3067
rect 1507 -3068 1508 -3067
rect 247 -3070 248 -3069
rect 779 -3070 780 -3069
rect 831 -3070 832 -3069
rect 1472 -3070 1473 -3069
rect 597 -3072 598 -3071
rect 779 -3072 780 -3071
rect 597 -3074 598 -3073
rect 635 -3074 636 -3073
rect 30 -3085 31 -3084
rect 474 -3085 475 -3084
rect 478 -3085 479 -3084
rect 635 -3085 636 -3084
rect 646 -3085 647 -3084
rect 975 -3085 976 -3084
rect 999 -3085 1000 -3084
rect 1633 -3085 1634 -3084
rect 37 -3087 38 -3086
rect 86 -3087 87 -3086
rect 114 -3087 115 -3086
rect 212 -3087 213 -3086
rect 215 -3087 216 -3086
rect 254 -3087 255 -3086
rect 275 -3087 276 -3086
rect 800 -3087 801 -3086
rect 814 -3087 815 -3086
rect 1087 -3087 1088 -3086
rect 1090 -3087 1091 -3086
rect 1388 -3087 1389 -3086
rect 1475 -3087 1476 -3086
rect 1570 -3087 1571 -3086
rect 61 -3089 62 -3088
rect 625 -3089 626 -3088
rect 656 -3089 657 -3088
rect 779 -3089 780 -3088
rect 789 -3089 790 -3088
rect 842 -3089 843 -3088
rect 877 -3089 878 -3088
rect 1171 -3089 1172 -3088
rect 1388 -3089 1389 -3088
rect 1563 -3089 1564 -3088
rect 65 -3091 66 -3090
rect 79 -3091 80 -3090
rect 82 -3091 83 -3090
rect 436 -3091 437 -3090
rect 471 -3091 472 -3090
rect 803 -3091 804 -3090
rect 842 -3091 843 -3090
rect 982 -3091 983 -3090
rect 1020 -3091 1021 -3090
rect 1458 -3091 1459 -3090
rect 79 -3093 80 -3092
rect 695 -3093 696 -3092
rect 716 -3093 717 -3092
rect 915 -3093 916 -3092
rect 933 -3093 934 -3092
rect 1090 -3093 1091 -3092
rect 1171 -3093 1172 -3092
rect 1339 -3093 1340 -3092
rect 1444 -3093 1445 -3092
rect 1458 -3093 1459 -3092
rect 86 -3095 87 -3094
rect 177 -3095 178 -3094
rect 184 -3095 185 -3094
rect 950 -3095 951 -3094
rect 975 -3095 976 -3094
rect 1031 -3095 1032 -3094
rect 1062 -3095 1063 -3094
rect 1584 -3095 1585 -3094
rect 117 -3097 118 -3096
rect 1276 -3097 1277 -3096
rect 1339 -3097 1340 -3096
rect 1528 -3097 1529 -3096
rect 131 -3099 132 -3098
rect 205 -3099 206 -3098
rect 219 -3099 220 -3098
rect 222 -3099 223 -3098
rect 254 -3099 255 -3098
rect 926 -3099 927 -3098
rect 933 -3099 934 -3098
rect 1199 -3099 1200 -3098
rect 1276 -3099 1277 -3098
rect 1430 -3099 1431 -3098
rect 135 -3101 136 -3100
rect 163 -3101 164 -3100
rect 177 -3101 178 -3100
rect 240 -3101 241 -3100
rect 282 -3101 283 -3100
rect 394 -3101 395 -3100
rect 404 -3101 405 -3100
rect 436 -3101 437 -3100
rect 453 -3101 454 -3100
rect 926 -3101 927 -3100
rect 940 -3101 941 -3100
rect 1199 -3101 1200 -3100
rect 1423 -3101 1424 -3100
rect 1444 -3101 1445 -3100
rect 51 -3103 52 -3102
rect 282 -3103 283 -3102
rect 303 -3103 304 -3102
rect 502 -3103 503 -3102
rect 527 -3103 528 -3102
rect 625 -3103 626 -3102
rect 674 -3103 675 -3102
rect 761 -3103 762 -3102
rect 779 -3103 780 -3102
rect 1038 -3103 1039 -3102
rect 1083 -3103 1084 -3102
rect 1367 -3103 1368 -3102
rect 1423 -3103 1424 -3102
rect 1605 -3103 1606 -3102
rect 93 -3105 94 -3104
rect 303 -3105 304 -3104
rect 345 -3105 346 -3104
rect 352 -3105 353 -3104
rect 366 -3105 367 -3104
rect 583 -3105 584 -3104
rect 593 -3105 594 -3104
rect 660 -3105 661 -3104
rect 674 -3105 675 -3104
rect 744 -3105 745 -3104
rect 758 -3105 759 -3104
rect 919 -3105 920 -3104
rect 940 -3105 941 -3104
rect 1059 -3105 1060 -3104
rect 1367 -3105 1368 -3104
rect 1542 -3105 1543 -3104
rect 1605 -3105 1606 -3104
rect 1647 -3105 1648 -3104
rect 93 -3107 94 -3106
rect 737 -3107 738 -3106
rect 744 -3107 745 -3106
rect 891 -3107 892 -3106
rect 919 -3107 920 -3106
rect 1052 -3107 1053 -3106
rect 1430 -3107 1431 -3106
rect 1612 -3107 1613 -3106
rect 135 -3109 136 -3108
rect 681 -3109 682 -3108
rect 684 -3109 685 -3108
rect 1360 -3109 1361 -3108
rect 142 -3111 143 -3110
rect 1486 -3111 1487 -3110
rect 142 -3113 143 -3112
rect 772 -3113 773 -3112
rect 793 -3113 794 -3112
rect 796 -3113 797 -3112
rect 800 -3113 801 -3112
rect 838 -3113 839 -3112
rect 877 -3113 878 -3112
rect 1024 -3113 1025 -3112
rect 1031 -3113 1032 -3112
rect 1087 -3113 1088 -3112
rect 1360 -3113 1361 -3112
rect 1535 -3113 1536 -3112
rect 145 -3115 146 -3114
rect 170 -3115 171 -3114
rect 184 -3115 185 -3114
rect 513 -3115 514 -3114
rect 534 -3115 535 -3114
rect 828 -3115 829 -3114
rect 838 -3115 839 -3114
rect 1066 -3115 1067 -3114
rect 1486 -3115 1487 -3114
rect 1626 -3115 1627 -3114
rect 121 -3117 122 -3116
rect 534 -3117 535 -3116
rect 562 -3117 563 -3116
rect 646 -3117 647 -3116
rect 660 -3117 661 -3116
rect 782 -3117 783 -3116
rect 793 -3117 794 -3116
rect 1640 -3117 1641 -3116
rect 100 -3119 101 -3118
rect 121 -3119 122 -3118
rect 149 -3119 150 -3118
rect 1395 -3119 1396 -3118
rect 89 -3121 90 -3120
rect 100 -3121 101 -3120
rect 152 -3121 153 -3120
rect 268 -3121 269 -3120
rect 348 -3121 349 -3120
rect 380 -3121 381 -3120
rect 394 -3121 395 -3120
rect 506 -3121 507 -3120
rect 562 -3121 563 -3120
rect 821 -3121 822 -3120
rect 828 -3121 829 -3120
rect 968 -3121 969 -3120
rect 982 -3121 983 -3120
rect 1129 -3121 1130 -3120
rect 44 -3123 45 -3122
rect 268 -3123 269 -3122
rect 352 -3123 353 -3122
rect 590 -3123 591 -3122
rect 618 -3123 619 -3122
rect 702 -3123 703 -3122
rect 716 -3123 717 -3122
rect 835 -3123 836 -3122
rect 947 -3123 948 -3122
rect 1164 -3123 1165 -3122
rect 152 -3125 153 -3124
rect 786 -3125 787 -3124
rect 821 -3125 822 -3124
rect 1101 -3125 1102 -3124
rect 1129 -3125 1130 -3124
rect 1283 -3125 1284 -3124
rect 156 -3127 157 -3126
rect 506 -3127 507 -3126
rect 576 -3127 577 -3126
rect 1059 -3127 1060 -3126
rect 1066 -3127 1067 -3126
rect 1234 -3127 1235 -3126
rect 1283 -3127 1284 -3126
rect 1465 -3127 1466 -3126
rect 156 -3129 157 -3128
rect 653 -3129 654 -3128
rect 688 -3129 689 -3128
rect 723 -3129 724 -3128
rect 730 -3129 731 -3128
rect 814 -3129 815 -3128
rect 835 -3129 836 -3128
rect 1353 -3129 1354 -3128
rect 163 -3131 164 -3130
rect 740 -3131 741 -3130
rect 772 -3131 773 -3130
rect 1073 -3131 1074 -3130
rect 1164 -3131 1165 -3130
rect 1269 -3131 1270 -3130
rect 170 -3133 171 -3132
rect 401 -3133 402 -3132
rect 429 -3133 430 -3132
rect 583 -3133 584 -3132
rect 653 -3133 654 -3132
rect 688 -3133 689 -3132
rect 691 -3133 692 -3132
rect 1598 -3133 1599 -3132
rect 191 -3135 192 -3134
rect 201 -3135 202 -3134
rect 219 -3135 220 -3134
rect 443 -3135 444 -3134
rect 457 -3135 458 -3134
rect 513 -3135 514 -3134
rect 579 -3135 580 -3134
rect 1101 -3135 1102 -3134
rect 1234 -3135 1235 -3134
rect 1409 -3135 1410 -3134
rect 128 -3137 129 -3136
rect 457 -3137 458 -3136
rect 478 -3137 479 -3136
rect 751 -3137 752 -3136
rect 786 -3137 787 -3136
rect 898 -3137 899 -3136
rect 947 -3137 948 -3136
rect 1402 -3137 1403 -3136
rect 1409 -3137 1410 -3136
rect 1514 -3137 1515 -3136
rect 72 -3139 73 -3138
rect 128 -3139 129 -3138
rect 191 -3139 192 -3138
rect 247 -3139 248 -3138
rect 261 -3139 262 -3138
rect 443 -3139 444 -3138
rect 492 -3139 493 -3138
rect 527 -3139 528 -3138
rect 681 -3139 682 -3138
rect 723 -3139 724 -3138
rect 730 -3139 731 -3138
rect 849 -3139 850 -3138
rect 898 -3139 899 -3138
rect 989 -3139 990 -3138
rect 1003 -3139 1004 -3138
rect 1073 -3139 1074 -3138
rect 1269 -3139 1270 -3138
rect 1521 -3139 1522 -3138
rect 72 -3141 73 -3140
rect 226 -3141 227 -3140
rect 233 -3141 234 -3140
rect 247 -3141 248 -3140
rect 261 -3141 262 -3140
rect 289 -3141 290 -3140
rect 366 -3141 367 -3140
rect 415 -3141 416 -3140
rect 432 -3141 433 -3140
rect 464 -3141 465 -3140
rect 492 -3141 493 -3140
rect 548 -3141 549 -3140
rect 695 -3141 696 -3140
rect 824 -3141 825 -3140
rect 849 -3141 850 -3140
rect 954 -3141 955 -3140
rect 968 -3141 969 -3140
rect 1227 -3141 1228 -3140
rect 1297 -3141 1298 -3140
rect 1514 -3141 1515 -3140
rect 198 -3143 199 -3142
rect 1080 -3143 1081 -3142
rect 1178 -3143 1179 -3142
rect 1297 -3143 1298 -3142
rect 1325 -3143 1326 -3142
rect 1521 -3143 1522 -3142
rect 149 -3145 150 -3144
rect 1080 -3145 1081 -3144
rect 1178 -3145 1179 -3144
rect 1311 -3145 1312 -3144
rect 1325 -3145 1326 -3144
rect 1500 -3145 1501 -3144
rect 198 -3147 199 -3146
rect 870 -3147 871 -3146
rect 954 -3147 955 -3146
rect 1150 -3147 1151 -3146
rect 1227 -3147 1228 -3146
rect 1416 -3147 1417 -3146
rect 222 -3149 223 -3148
rect 289 -3149 290 -3148
rect 369 -3149 370 -3148
rect 408 -3149 409 -3148
rect 537 -3149 538 -3148
rect 1416 -3149 1417 -3148
rect 226 -3151 227 -3150
rect 604 -3151 605 -3150
rect 702 -3151 703 -3150
rect 856 -3151 857 -3150
rect 870 -3151 871 -3150
rect 1412 -3151 1413 -3150
rect 233 -3153 234 -3152
rect 611 -3153 612 -3152
rect 737 -3153 738 -3152
rect 765 -3153 766 -3152
rect 856 -3153 857 -3152
rect 884 -3153 885 -3152
rect 989 -3153 990 -3152
rect 1437 -3153 1438 -3152
rect 373 -3155 374 -3154
rect 415 -3155 416 -3154
rect 548 -3155 549 -3154
rect 667 -3155 668 -3154
rect 751 -3155 752 -3154
rect 905 -3155 906 -3154
rect 1003 -3155 1004 -3154
rect 1157 -3155 1158 -3154
rect 1311 -3155 1312 -3154
rect 1479 -3155 1480 -3154
rect 107 -3157 108 -3156
rect 373 -3157 374 -3156
rect 380 -3157 381 -3156
rect 541 -3157 542 -3156
rect 597 -3157 598 -3156
rect 604 -3157 605 -3156
rect 611 -3157 612 -3156
rect 709 -3157 710 -3156
rect 765 -3157 766 -3156
rect 1013 -3157 1014 -3156
rect 1024 -3157 1025 -3156
rect 1115 -3157 1116 -3156
rect 1122 -3157 1123 -3156
rect 1500 -3157 1501 -3156
rect 107 -3159 108 -3158
rect 639 -3159 640 -3158
rect 667 -3159 668 -3158
rect 863 -3159 864 -3158
rect 884 -3159 885 -3158
rect 1010 -3159 1011 -3158
rect 1038 -3159 1039 -3158
rect 1248 -3159 1249 -3158
rect 1402 -3159 1403 -3158
rect 1591 -3159 1592 -3158
rect 387 -3161 388 -3160
rect 464 -3161 465 -3160
rect 471 -3161 472 -3160
rect 863 -3161 864 -3160
rect 905 -3161 906 -3160
rect 912 -3161 913 -3160
rect 1052 -3161 1053 -3160
rect 1220 -3161 1221 -3160
rect 1248 -3161 1249 -3160
rect 1507 -3161 1508 -3160
rect 387 -3163 388 -3162
rect 1143 -3163 1144 -3162
rect 1150 -3163 1151 -3162
rect 1213 -3163 1214 -3162
rect 1220 -3163 1221 -3162
rect 1381 -3163 1382 -3162
rect 1437 -3163 1438 -3162
rect 1619 -3163 1620 -3162
rect 401 -3165 402 -3164
rect 520 -3165 521 -3164
rect 590 -3165 591 -3164
rect 597 -3165 598 -3164
rect 632 -3165 633 -3164
rect 1213 -3165 1214 -3164
rect 1304 -3165 1305 -3164
rect 1507 -3165 1508 -3164
rect 114 -3167 115 -3166
rect 520 -3167 521 -3166
rect 632 -3167 633 -3166
rect 961 -3167 962 -3166
rect 978 -3167 979 -3166
rect 1304 -3167 1305 -3166
rect 1381 -3167 1382 -3166
rect 1556 -3167 1557 -3166
rect 408 -3169 409 -3168
rect 569 -3169 570 -3168
rect 639 -3169 640 -3168
rect 1206 -3169 1207 -3168
rect 429 -3171 430 -3170
rect 569 -3171 570 -3170
rect 709 -3171 710 -3170
rect 807 -3171 808 -3170
rect 912 -3171 913 -3170
rect 1045 -3171 1046 -3170
rect 1094 -3171 1095 -3170
rect 1115 -3171 1116 -3170
rect 1122 -3171 1123 -3170
rect 1318 -3171 1319 -3170
rect 576 -3173 577 -3172
rect 807 -3173 808 -3172
rect 961 -3173 962 -3172
rect 1108 -3173 1109 -3172
rect 1136 -3173 1137 -3172
rect 1157 -3173 1158 -3172
rect 1185 -3173 1186 -3172
rect 1479 -3173 1480 -3172
rect 1045 -3175 1046 -3174
rect 1192 -3175 1193 -3174
rect 1206 -3175 1207 -3174
rect 1374 -3175 1375 -3174
rect 1094 -3177 1095 -3176
rect 1262 -3177 1263 -3176
rect 1318 -3177 1319 -3176
rect 1493 -3177 1494 -3176
rect 996 -3179 997 -3178
rect 1493 -3179 1494 -3178
rect 996 -3181 997 -3180
rect 1395 -3181 1396 -3180
rect 1017 -3183 1018 -3182
rect 1262 -3183 1263 -3182
rect 1374 -3183 1375 -3182
rect 1549 -3183 1550 -3182
rect 1017 -3185 1018 -3184
rect 1290 -3185 1291 -3184
rect 1108 -3187 1109 -3186
rect 1654 -3187 1655 -3186
rect 1136 -3189 1137 -3188
rect 1255 -3189 1256 -3188
rect 1290 -3189 1291 -3188
rect 1472 -3189 1473 -3188
rect 1143 -3191 1144 -3190
rect 1241 -3191 1242 -3190
rect 1255 -3191 1256 -3190
rect 1451 -3191 1452 -3190
rect 450 -3193 451 -3192
rect 1451 -3193 1452 -3192
rect 310 -3195 311 -3194
rect 450 -3195 451 -3194
rect 1185 -3195 1186 -3194
rect 1332 -3195 1333 -3194
rect 310 -3197 311 -3196
rect 331 -3197 332 -3196
rect 621 -3197 622 -3196
rect 1332 -3197 1333 -3196
rect 331 -3199 332 -3198
rect 422 -3199 423 -3198
rect 1192 -3199 1193 -3198
rect 1346 -3199 1347 -3198
rect 422 -3201 423 -3200
rect 485 -3201 486 -3200
rect 1241 -3201 1242 -3200
rect 1577 -3201 1578 -3200
rect 296 -3203 297 -3202
rect 485 -3203 486 -3202
rect 1346 -3203 1347 -3202
rect 1465 -3203 1466 -3202
rect 296 -3205 297 -3204
rect 338 -3205 339 -3204
rect 338 -3207 339 -3206
rect 359 -3207 360 -3206
rect 359 -3209 360 -3208
rect 555 -3209 556 -3208
rect 499 -3211 500 -3210
rect 555 -3211 556 -3210
rect 275 -3213 276 -3212
rect 499 -3213 500 -3212
rect 65 -3224 66 -3223
rect 114 -3224 115 -3223
rect 121 -3224 122 -3223
rect 499 -3224 500 -3223
rect 502 -3224 503 -3223
rect 716 -3224 717 -3223
rect 779 -3224 780 -3223
rect 870 -3224 871 -3223
rect 880 -3224 881 -3223
rect 1031 -3224 1032 -3223
rect 1059 -3224 1060 -3223
rect 1332 -3224 1333 -3223
rect 1346 -3224 1347 -3223
rect 1479 -3224 1480 -3223
rect 1584 -3224 1585 -3223
rect 1605 -3224 1606 -3223
rect 72 -3226 73 -3225
rect 471 -3226 472 -3225
rect 485 -3226 486 -3225
rect 579 -3226 580 -3225
rect 593 -3226 594 -3225
rect 674 -3226 675 -3225
rect 684 -3226 685 -3225
rect 786 -3226 787 -3225
rect 800 -3226 801 -3225
rect 1356 -3226 1357 -3225
rect 1409 -3226 1410 -3225
rect 1521 -3226 1522 -3225
rect 86 -3228 87 -3227
rect 401 -3228 402 -3227
rect 404 -3228 405 -3227
rect 527 -3228 528 -3227
rect 544 -3228 545 -3227
rect 555 -3228 556 -3227
rect 576 -3228 577 -3227
rect 611 -3228 612 -3227
rect 625 -3228 626 -3227
rect 796 -3228 797 -3227
rect 800 -3228 801 -3227
rect 849 -3228 850 -3227
rect 894 -3228 895 -3227
rect 1157 -3228 1158 -3227
rect 1185 -3228 1186 -3227
rect 1209 -3228 1210 -3227
rect 1297 -3228 1298 -3227
rect 1493 -3228 1494 -3227
rect 142 -3230 143 -3229
rect 576 -3230 577 -3229
rect 611 -3230 612 -3229
rect 737 -3230 738 -3229
rect 849 -3230 850 -3229
rect 954 -3230 955 -3229
rect 999 -3230 1000 -3229
rect 1003 -3230 1004 -3229
rect 1010 -3230 1011 -3229
rect 1269 -3230 1270 -3229
rect 1300 -3230 1301 -3229
rect 1465 -3230 1466 -3229
rect 149 -3232 150 -3231
rect 191 -3232 192 -3231
rect 212 -3232 213 -3231
rect 240 -3232 241 -3231
rect 243 -3232 244 -3231
rect 317 -3232 318 -3231
rect 324 -3232 325 -3231
rect 1013 -3232 1014 -3231
rect 1020 -3232 1021 -3231
rect 1136 -3232 1137 -3231
rect 1269 -3232 1270 -3231
rect 1381 -3232 1382 -3231
rect 1458 -3232 1459 -3231
rect 1531 -3232 1532 -3231
rect 107 -3234 108 -3233
rect 212 -3234 213 -3233
rect 226 -3234 227 -3233
rect 485 -3234 486 -3233
rect 492 -3234 493 -3233
rect 772 -3234 773 -3233
rect 905 -3234 906 -3233
rect 985 -3234 986 -3233
rect 1010 -3234 1011 -3233
rect 1206 -3234 1207 -3233
rect 1325 -3234 1326 -3233
rect 1328 -3234 1329 -3233
rect 1332 -3234 1333 -3233
rect 1388 -3234 1389 -3233
rect 152 -3236 153 -3235
rect 359 -3236 360 -3235
rect 387 -3236 388 -3235
rect 390 -3236 391 -3235
rect 415 -3236 416 -3235
rect 541 -3236 542 -3235
rect 544 -3236 545 -3235
rect 835 -3236 836 -3235
rect 905 -3236 906 -3235
rect 1248 -3236 1249 -3235
rect 1325 -3236 1326 -3235
rect 1360 -3236 1361 -3235
rect 1381 -3236 1382 -3235
rect 1507 -3236 1508 -3235
rect 156 -3238 157 -3237
rect 527 -3238 528 -3237
rect 541 -3238 542 -3237
rect 947 -3238 948 -3237
rect 954 -3238 955 -3237
rect 1199 -3238 1200 -3237
rect 1346 -3238 1347 -3237
rect 1423 -3238 1424 -3237
rect 170 -3240 171 -3239
rect 492 -3240 493 -3239
rect 499 -3240 500 -3239
rect 548 -3240 549 -3239
rect 555 -3240 556 -3239
rect 604 -3240 605 -3239
rect 625 -3240 626 -3239
rect 807 -3240 808 -3239
rect 940 -3240 941 -3239
rect 996 -3240 997 -3239
rect 1031 -3240 1032 -3239
rect 1220 -3240 1221 -3239
rect 1349 -3240 1350 -3239
rect 1514 -3240 1515 -3239
rect 93 -3242 94 -3241
rect 170 -3242 171 -3241
rect 177 -3242 178 -3241
rect 348 -3242 349 -3241
rect 359 -3242 360 -3241
rect 394 -3242 395 -3241
rect 429 -3242 430 -3241
rect 450 -3242 451 -3241
rect 457 -3242 458 -3241
rect 590 -3242 591 -3241
rect 604 -3242 605 -3241
rect 667 -3242 668 -3241
rect 705 -3242 706 -3241
rect 1017 -3242 1018 -3241
rect 1087 -3242 1088 -3241
rect 1318 -3242 1319 -3241
rect 1353 -3242 1354 -3241
rect 1486 -3242 1487 -3241
rect 191 -3244 192 -3243
rect 205 -3244 206 -3243
rect 226 -3244 227 -3243
rect 838 -3244 839 -3243
rect 940 -3244 941 -3243
rect 982 -3244 983 -3243
rect 996 -3244 997 -3243
rect 1171 -3244 1172 -3243
rect 1199 -3244 1200 -3243
rect 1241 -3244 1242 -3243
rect 1283 -3244 1284 -3243
rect 1353 -3244 1354 -3243
rect 1388 -3244 1389 -3243
rect 1395 -3244 1396 -3243
rect 205 -3246 206 -3245
rect 632 -3246 633 -3245
rect 653 -3246 654 -3245
rect 702 -3246 703 -3245
rect 709 -3246 710 -3245
rect 824 -3246 825 -3245
rect 919 -3246 920 -3245
rect 1283 -3246 1284 -3245
rect 247 -3248 248 -3247
rect 495 -3248 496 -3247
rect 520 -3248 521 -3247
rect 779 -3248 780 -3247
rect 919 -3248 920 -3247
rect 1080 -3248 1081 -3247
rect 1090 -3248 1091 -3247
rect 1178 -3248 1179 -3247
rect 1220 -3248 1221 -3247
rect 1437 -3248 1438 -3247
rect 135 -3250 136 -3249
rect 247 -3250 248 -3249
rect 254 -3250 255 -3249
rect 677 -3250 678 -3249
rect 709 -3250 710 -3249
rect 901 -3250 902 -3249
rect 947 -3250 948 -3249
rect 1115 -3250 1116 -3249
rect 1129 -3250 1130 -3249
rect 1188 -3250 1189 -3249
rect 1234 -3250 1235 -3249
rect 1241 -3250 1242 -3249
rect 128 -3252 129 -3251
rect 135 -3252 136 -3251
rect 254 -3252 255 -3251
rect 702 -3252 703 -3251
rect 716 -3252 717 -3251
rect 828 -3252 829 -3251
rect 891 -3252 892 -3251
rect 1178 -3252 1179 -3251
rect 1234 -3252 1235 -3251
rect 1304 -3252 1305 -3251
rect 261 -3254 262 -3253
rect 394 -3254 395 -3253
rect 429 -3254 430 -3253
rect 789 -3254 790 -3253
rect 828 -3254 829 -3253
rect 1500 -3254 1501 -3253
rect 261 -3256 262 -3255
rect 331 -3256 332 -3255
rect 338 -3256 339 -3255
rect 439 -3256 440 -3255
rect 450 -3256 451 -3255
rect 478 -3256 479 -3255
rect 520 -3256 521 -3255
rect 569 -3256 570 -3255
rect 632 -3256 633 -3255
rect 730 -3256 731 -3255
rect 737 -3256 738 -3255
rect 1073 -3256 1074 -3255
rect 1080 -3256 1081 -3255
rect 1262 -3256 1263 -3255
rect 1304 -3256 1305 -3255
rect 1475 -3256 1476 -3255
rect 198 -3258 199 -3257
rect 730 -3258 731 -3257
rect 751 -3258 752 -3257
rect 1136 -3258 1137 -3257
rect 1171 -3258 1172 -3257
rect 1276 -3258 1277 -3257
rect 79 -3260 80 -3259
rect 198 -3260 199 -3259
rect 275 -3260 276 -3259
rect 331 -3260 332 -3259
rect 352 -3260 353 -3259
rect 478 -3260 479 -3259
rect 548 -3260 549 -3259
rect 660 -3260 661 -3259
rect 667 -3260 668 -3259
rect 744 -3260 745 -3259
rect 751 -3260 752 -3259
rect 1227 -3260 1228 -3259
rect 1276 -3260 1277 -3259
rect 1374 -3260 1375 -3259
rect 184 -3262 185 -3261
rect 275 -3262 276 -3261
rect 282 -3262 283 -3261
rect 338 -3262 339 -3261
rect 352 -3262 353 -3261
rect 408 -3262 409 -3261
rect 422 -3262 423 -3261
rect 569 -3262 570 -3261
rect 660 -3262 661 -3261
rect 681 -3262 682 -3261
rect 723 -3262 724 -3261
rect 807 -3262 808 -3261
rect 891 -3262 892 -3261
rect 1262 -3262 1263 -3261
rect 163 -3264 164 -3263
rect 408 -3264 409 -3263
rect 422 -3264 423 -3263
rect 618 -3264 619 -3263
rect 681 -3264 682 -3263
rect 695 -3264 696 -3263
rect 723 -3264 724 -3263
rect 842 -3264 843 -3263
rect 968 -3264 969 -3263
rect 1003 -3264 1004 -3263
rect 1052 -3264 1053 -3263
rect 1318 -3264 1319 -3263
rect 100 -3266 101 -3265
rect 163 -3266 164 -3265
rect 184 -3266 185 -3265
rect 534 -3266 535 -3265
rect 618 -3266 619 -3265
rect 989 -3266 990 -3265
rect 1045 -3266 1046 -3265
rect 1052 -3266 1053 -3265
rect 1073 -3266 1074 -3265
rect 1143 -3266 1144 -3265
rect 1213 -3266 1214 -3265
rect 1227 -3266 1228 -3265
rect 282 -3268 283 -3267
rect 950 -3268 951 -3267
rect 968 -3268 969 -3267
rect 1038 -3268 1039 -3267
rect 1045 -3268 1046 -3267
rect 1255 -3268 1256 -3267
rect 296 -3270 297 -3269
rect 324 -3270 325 -3269
rect 373 -3270 374 -3269
rect 415 -3270 416 -3269
rect 457 -3270 458 -3269
rect 793 -3270 794 -3269
rect 814 -3270 815 -3269
rect 1038 -3270 1039 -3269
rect 1094 -3270 1095 -3269
rect 1258 -3270 1259 -3269
rect 296 -3272 297 -3271
rect 380 -3272 381 -3271
rect 387 -3272 388 -3271
rect 443 -3272 444 -3271
rect 471 -3272 472 -3271
rect 530 -3272 531 -3271
rect 534 -3272 535 -3271
rect 982 -3272 983 -3271
rect 1094 -3272 1095 -3271
rect 1290 -3272 1291 -3271
rect 303 -3274 304 -3273
rect 373 -3274 374 -3273
rect 380 -3274 381 -3273
rect 513 -3274 514 -3273
rect 695 -3274 696 -3273
rect 877 -3274 878 -3273
rect 1101 -3274 1102 -3273
rect 1157 -3274 1158 -3273
rect 1290 -3274 1291 -3273
rect 1444 -3274 1445 -3273
rect 303 -3276 304 -3275
rect 310 -3276 311 -3275
rect 317 -3276 318 -3275
rect 345 -3276 346 -3275
rect 443 -3276 444 -3275
rect 646 -3276 647 -3275
rect 744 -3276 745 -3275
rect 821 -3276 822 -3275
rect 842 -3276 843 -3275
rect 1339 -3276 1340 -3275
rect 177 -3278 178 -3277
rect 345 -3278 346 -3277
rect 513 -3278 514 -3277
rect 583 -3278 584 -3277
rect 758 -3278 759 -3277
rect 877 -3278 878 -3277
rect 1101 -3278 1102 -3277
rect 1416 -3278 1417 -3277
rect 289 -3280 290 -3279
rect 310 -3280 311 -3279
rect 464 -3280 465 -3279
rect 583 -3280 584 -3279
rect 758 -3280 759 -3279
rect 884 -3280 885 -3279
rect 1115 -3280 1116 -3279
rect 1430 -3280 1431 -3279
rect 289 -3282 290 -3281
rect 436 -3282 437 -3281
rect 464 -3282 465 -3281
rect 688 -3282 689 -3281
rect 772 -3282 773 -3281
rect 1265 -3282 1266 -3281
rect 1311 -3282 1312 -3281
rect 1339 -3282 1340 -3281
rect 366 -3284 367 -3283
rect 436 -3284 437 -3283
rect 793 -3284 794 -3283
rect 961 -3284 962 -3283
rect 1129 -3284 1130 -3283
rect 1164 -3284 1165 -3283
rect 1311 -3284 1312 -3283
rect 1367 -3284 1368 -3283
rect 219 -3286 220 -3285
rect 366 -3286 367 -3285
rect 814 -3286 815 -3285
rect 1024 -3286 1025 -3285
rect 1143 -3286 1144 -3285
rect 1150 -3286 1151 -3285
rect 1164 -3286 1165 -3285
rect 1192 -3286 1193 -3285
rect 1328 -3286 1329 -3285
rect 1360 -3286 1361 -3285
rect 219 -3288 220 -3287
rect 562 -3288 563 -3287
rect 821 -3288 822 -3287
rect 933 -3288 934 -3287
rect 1150 -3288 1151 -3287
rect 1255 -3288 1256 -3287
rect 506 -3290 507 -3289
rect 562 -3290 563 -3289
rect 856 -3290 857 -3289
rect 884 -3290 885 -3289
rect 915 -3290 916 -3289
rect 961 -3290 962 -3289
rect 1192 -3290 1193 -3289
rect 1402 -3290 1403 -3289
rect 506 -3292 507 -3291
rect 765 -3292 766 -3291
rect 856 -3292 857 -3291
rect 898 -3292 899 -3291
rect 926 -3292 927 -3291
rect 1024 -3292 1025 -3291
rect 765 -3294 766 -3293
rect 912 -3294 913 -3293
rect 926 -3294 927 -3293
rect 1066 -3294 1067 -3293
rect 863 -3296 864 -3295
rect 989 -3296 990 -3295
rect 1066 -3296 1067 -3295
rect 1213 -3296 1214 -3295
rect 639 -3298 640 -3297
rect 863 -3298 864 -3297
rect 912 -3298 913 -3297
rect 975 -3298 976 -3297
rect 639 -3300 640 -3299
rect 656 -3300 657 -3299
rect 933 -3300 934 -3299
rect 1108 -3300 1109 -3299
rect 835 -3302 836 -3301
rect 1108 -3302 1109 -3301
rect 975 -3304 976 -3303
rect 1122 -3304 1123 -3303
rect 1122 -3306 1123 -3305
rect 1451 -3306 1452 -3305
rect 131 -3317 132 -3316
rect 135 -3317 136 -3316
rect 163 -3317 164 -3316
rect 579 -3317 580 -3316
rect 590 -3317 591 -3316
rect 688 -3317 689 -3316
rect 691 -3317 692 -3316
rect 1157 -3317 1158 -3316
rect 1178 -3317 1179 -3316
rect 1528 -3317 1529 -3316
rect 1577 -3317 1578 -3316
rect 1584 -3317 1585 -3316
rect 205 -3319 206 -3318
rect 541 -3319 542 -3318
rect 590 -3319 591 -3318
rect 842 -3319 843 -3318
rect 870 -3319 871 -3318
rect 1192 -3319 1193 -3318
rect 1209 -3319 1210 -3318
rect 1276 -3319 1277 -3318
rect 1360 -3319 1361 -3318
rect 1374 -3319 1375 -3318
rect 233 -3321 234 -3320
rect 492 -3321 493 -3320
rect 506 -3321 507 -3320
rect 803 -3321 804 -3320
rect 870 -3321 871 -3320
rect 985 -3321 986 -3320
rect 1003 -3321 1004 -3320
rect 1108 -3321 1109 -3320
rect 1111 -3321 1112 -3320
rect 1290 -3321 1291 -3320
rect 212 -3323 213 -3322
rect 506 -3323 507 -3322
rect 513 -3323 514 -3322
rect 544 -3323 545 -3322
rect 614 -3323 615 -3322
rect 1150 -3323 1151 -3322
rect 1153 -3323 1154 -3322
rect 1234 -3323 1235 -3322
rect 1248 -3323 1249 -3322
rect 1325 -3323 1326 -3322
rect 247 -3325 248 -3324
rect 443 -3325 444 -3324
rect 464 -3325 465 -3324
rect 674 -3325 675 -3324
rect 705 -3325 706 -3324
rect 877 -3325 878 -3324
rect 880 -3325 881 -3324
rect 1136 -3325 1137 -3324
rect 1192 -3325 1193 -3324
rect 1283 -3325 1284 -3324
rect 198 -3327 199 -3326
rect 247 -3327 248 -3326
rect 268 -3327 269 -3326
rect 618 -3327 619 -3326
rect 621 -3327 622 -3326
rect 908 -3327 909 -3326
rect 915 -3327 916 -3326
rect 1143 -3327 1144 -3326
rect 1199 -3327 1200 -3326
rect 1248 -3327 1249 -3326
rect 1262 -3327 1263 -3326
rect 1311 -3327 1312 -3326
rect 240 -3329 241 -3328
rect 268 -3329 269 -3328
rect 310 -3329 311 -3328
rect 401 -3329 402 -3328
rect 436 -3329 437 -3328
rect 471 -3329 472 -3328
rect 485 -3329 486 -3328
rect 950 -3329 951 -3328
rect 961 -3329 962 -3328
rect 1157 -3329 1158 -3328
rect 1171 -3329 1172 -3328
rect 1199 -3329 1200 -3328
rect 1213 -3329 1214 -3328
rect 1241 -3329 1242 -3328
rect 1311 -3329 1312 -3328
rect 1332 -3329 1333 -3328
rect 177 -3331 178 -3330
rect 240 -3331 241 -3330
rect 359 -3331 360 -3330
rect 513 -3331 514 -3330
rect 523 -3331 524 -3330
rect 688 -3331 689 -3330
rect 716 -3331 717 -3330
rect 877 -3331 878 -3330
rect 894 -3331 895 -3330
rect 1216 -3331 1217 -3330
rect 1234 -3331 1235 -3330
rect 1318 -3331 1319 -3330
rect 1332 -3331 1333 -3330
rect 1381 -3331 1382 -3330
rect 359 -3333 360 -3332
rect 366 -3333 367 -3332
rect 380 -3333 381 -3332
rect 443 -3333 444 -3332
rect 471 -3333 472 -3332
rect 499 -3333 500 -3332
rect 618 -3333 619 -3332
rect 709 -3333 710 -3332
rect 716 -3333 717 -3332
rect 779 -3333 780 -3332
rect 789 -3333 790 -3332
rect 800 -3333 801 -3332
rect 901 -3333 902 -3332
rect 940 -3333 941 -3332
rect 947 -3333 948 -3332
rect 1136 -3333 1137 -3332
rect 1171 -3333 1172 -3332
rect 1297 -3333 1298 -3332
rect 1353 -3333 1354 -3332
rect 1381 -3333 1382 -3332
rect 170 -3335 171 -3334
rect 499 -3335 500 -3334
rect 632 -3335 633 -3334
rect 898 -3335 899 -3334
rect 947 -3335 948 -3334
rect 968 -3335 969 -3334
rect 982 -3335 983 -3334
rect 1164 -3335 1165 -3334
rect 1213 -3335 1214 -3334
rect 1318 -3335 1319 -3334
rect 275 -3337 276 -3336
rect 366 -3337 367 -3336
rect 380 -3337 381 -3336
rect 446 -3337 447 -3336
rect 478 -3337 479 -3336
rect 485 -3337 486 -3336
rect 632 -3337 633 -3336
rect 723 -3337 724 -3336
rect 730 -3337 731 -3336
rect 873 -3337 874 -3336
rect 898 -3337 899 -3336
rect 926 -3337 927 -3336
rect 961 -3337 962 -3336
rect 1101 -3337 1102 -3336
rect 1164 -3337 1165 -3336
rect 1269 -3337 1270 -3336
rect 394 -3339 395 -3338
rect 464 -3339 465 -3338
rect 478 -3339 479 -3338
rect 520 -3339 521 -3338
rect 639 -3339 640 -3338
rect 779 -3339 780 -3338
rect 891 -3339 892 -3338
rect 926 -3339 927 -3338
rect 982 -3339 983 -3338
rect 1122 -3339 1123 -3338
rect 1241 -3339 1242 -3338
rect 1339 -3339 1340 -3338
rect 345 -3341 346 -3340
rect 394 -3341 395 -3340
rect 401 -3341 402 -3340
rect 415 -3341 416 -3340
rect 576 -3341 577 -3340
rect 639 -3341 640 -3340
rect 667 -3341 668 -3340
rect 842 -3341 843 -3340
rect 996 -3341 997 -3340
rect 1101 -3341 1102 -3340
rect 282 -3343 283 -3342
rect 345 -3343 346 -3342
rect 548 -3343 549 -3342
rect 576 -3343 577 -3342
rect 667 -3343 668 -3342
rect 744 -3343 745 -3342
rect 758 -3343 759 -3342
rect 968 -3343 969 -3342
rect 1003 -3343 1004 -3342
rect 1087 -3343 1088 -3342
rect 1094 -3343 1095 -3342
rect 1122 -3343 1123 -3342
rect 184 -3345 185 -3344
rect 282 -3345 283 -3344
rect 317 -3345 318 -3344
rect 415 -3345 416 -3344
rect 530 -3345 531 -3344
rect 1087 -3345 1088 -3344
rect 226 -3347 227 -3346
rect 548 -3347 549 -3346
rect 583 -3347 584 -3346
rect 758 -3347 759 -3346
rect 863 -3347 864 -3346
rect 996 -3347 997 -3346
rect 1013 -3347 1014 -3346
rect 1220 -3347 1221 -3346
rect 219 -3349 220 -3348
rect 583 -3349 584 -3348
rect 674 -3349 675 -3348
rect 828 -3349 829 -3348
rect 1024 -3349 1025 -3348
rect 1129 -3349 1130 -3348
rect 317 -3351 318 -3350
rect 331 -3351 332 -3350
rect 408 -3351 409 -3350
rect 863 -3351 864 -3350
rect 1024 -3351 1025 -3350
rect 1227 -3351 1228 -3350
rect 296 -3353 297 -3352
rect 331 -3353 332 -3352
rect 373 -3353 374 -3352
rect 408 -3353 409 -3352
rect 709 -3353 710 -3352
rect 772 -3353 773 -3352
rect 828 -3353 829 -3352
rect 884 -3353 885 -3352
rect 1031 -3353 1032 -3352
rect 1034 -3353 1035 -3352
rect 1038 -3353 1039 -3352
rect 1185 -3353 1186 -3352
rect 191 -3355 192 -3354
rect 296 -3355 297 -3354
rect 660 -3355 661 -3354
rect 772 -3355 773 -3354
rect 814 -3355 815 -3354
rect 884 -3355 885 -3354
rect 989 -3355 990 -3354
rect 1038 -3355 1039 -3354
rect 1045 -3355 1046 -3354
rect 1143 -3355 1144 -3354
rect 1185 -3355 1186 -3354
rect 1206 -3355 1207 -3354
rect 261 -3357 262 -3356
rect 373 -3357 374 -3356
rect 660 -3357 661 -3356
rect 765 -3357 766 -3356
rect 849 -3357 850 -3356
rect 989 -3357 990 -3356
rect 1031 -3357 1032 -3356
rect 1115 -3357 1116 -3356
rect 1206 -3357 1207 -3356
rect 1251 -3357 1252 -3356
rect 681 -3359 682 -3358
rect 814 -3359 815 -3358
rect 1034 -3359 1035 -3358
rect 1115 -3359 1116 -3358
rect 681 -3361 682 -3360
rect 1062 -3361 1063 -3360
rect 1066 -3361 1067 -3360
rect 1094 -3361 1095 -3360
rect 702 -3363 703 -3362
rect 765 -3363 766 -3362
rect 786 -3363 787 -3362
rect 849 -3363 850 -3362
rect 1045 -3363 1046 -3362
rect 1073 -3363 1074 -3362
rect 1080 -3363 1081 -3362
rect 1129 -3363 1130 -3362
rect 646 -3365 647 -3364
rect 702 -3365 703 -3364
rect 723 -3365 724 -3364
rect 793 -3365 794 -3364
rect 856 -3365 857 -3364
rect 1080 -3365 1081 -3364
rect 611 -3367 612 -3366
rect 793 -3367 794 -3366
rect 856 -3367 857 -3366
rect 1167 -3367 1168 -3366
rect 254 -3369 255 -3368
rect 611 -3369 612 -3368
rect 646 -3369 647 -3368
rect 751 -3369 752 -3368
rect 786 -3369 787 -3368
rect 800 -3369 801 -3368
rect 933 -3369 934 -3368
rect 1073 -3369 1074 -3368
rect 737 -3371 738 -3370
rect 940 -3371 941 -3370
rect 1052 -3371 1053 -3370
rect 1108 -3371 1109 -3370
rect 737 -3373 738 -3372
rect 807 -3373 808 -3372
rect 933 -3373 934 -3372
rect 1020 -3373 1021 -3372
rect 1066 -3373 1067 -3372
rect 1265 -3373 1266 -3372
rect 387 -3375 388 -3374
rect 1020 -3375 1021 -3374
rect 1265 -3375 1266 -3374
rect 1346 -3375 1347 -3374
rect 387 -3377 388 -3376
rect 457 -3377 458 -3376
rect 597 -3377 598 -3376
rect 807 -3377 808 -3376
rect 450 -3379 451 -3378
rect 457 -3379 458 -3378
rect 597 -3379 598 -3378
rect 695 -3379 696 -3378
rect 744 -3379 745 -3378
rect 821 -3379 822 -3378
rect 450 -3381 451 -3380
rect 527 -3381 528 -3380
rect 695 -3381 696 -3380
rect 835 -3381 836 -3380
rect 527 -3383 528 -3382
rect 534 -3383 535 -3382
rect 562 -3383 563 -3382
rect 835 -3383 836 -3382
rect 534 -3385 535 -3384
rect 555 -3385 556 -3384
rect 562 -3385 563 -3384
rect 569 -3385 570 -3384
rect 751 -3385 752 -3384
rect 912 -3385 913 -3384
rect 555 -3387 556 -3386
rect 625 -3387 626 -3386
rect 821 -3387 822 -3386
rect 919 -3387 920 -3386
rect 569 -3389 570 -3388
rect 604 -3389 605 -3388
rect 625 -3389 626 -3388
rect 653 -3389 654 -3388
rect 912 -3389 913 -3388
rect 954 -3389 955 -3388
rect 422 -3391 423 -3390
rect 653 -3391 654 -3390
rect 919 -3391 920 -3390
rect 975 -3391 976 -3390
rect 338 -3393 339 -3392
rect 422 -3393 423 -3392
rect 604 -3393 605 -3392
rect 905 -3393 906 -3392
rect 954 -3393 955 -3392
rect 1017 -3393 1018 -3392
rect 338 -3395 339 -3394
rect 352 -3395 353 -3394
rect 905 -3395 906 -3394
rect 1010 -3395 1011 -3394
rect 324 -3397 325 -3396
rect 352 -3397 353 -3396
rect 975 -3397 976 -3396
rect 1059 -3397 1060 -3396
rect 303 -3399 304 -3398
rect 324 -3399 325 -3398
rect 1059 -3399 1060 -3398
rect 1304 -3399 1305 -3398
rect 289 -3401 290 -3400
rect 303 -3401 304 -3400
rect 289 -3403 290 -3402
rect 310 -3403 311 -3402
rect 240 -3414 241 -3413
rect 261 -3414 262 -3413
rect 268 -3414 269 -3413
rect 292 -3414 293 -3413
rect 338 -3414 339 -3413
rect 355 -3414 356 -3413
rect 376 -3414 377 -3413
rect 450 -3414 451 -3413
rect 457 -3414 458 -3413
rect 474 -3414 475 -3413
rect 485 -3414 486 -3413
rect 611 -3414 612 -3413
rect 663 -3414 664 -3413
rect 1038 -3414 1039 -3413
rect 1041 -3414 1042 -3413
rect 1045 -3414 1046 -3413
rect 1052 -3414 1053 -3413
rect 1073 -3414 1074 -3413
rect 1111 -3414 1112 -3413
rect 1192 -3414 1193 -3413
rect 1199 -3414 1200 -3413
rect 1213 -3414 1214 -3413
rect 1248 -3414 1249 -3413
rect 1269 -3414 1270 -3413
rect 1304 -3414 1305 -3413
rect 1311 -3414 1312 -3413
rect 1318 -3414 1319 -3413
rect 1346 -3414 1347 -3413
rect 1374 -3414 1375 -3413
rect 1395 -3414 1396 -3413
rect 247 -3416 248 -3415
rect 289 -3416 290 -3415
rect 317 -3416 318 -3415
rect 457 -3416 458 -3415
rect 499 -3416 500 -3415
rect 604 -3416 605 -3415
rect 702 -3416 703 -3415
rect 810 -3416 811 -3415
rect 824 -3416 825 -3415
rect 982 -3416 983 -3415
rect 989 -3416 990 -3415
rect 1055 -3416 1056 -3415
rect 1073 -3416 1074 -3415
rect 1101 -3416 1102 -3415
rect 1122 -3416 1123 -3415
rect 1125 -3416 1126 -3415
rect 1129 -3416 1130 -3415
rect 1160 -3416 1161 -3415
rect 1185 -3416 1186 -3415
rect 1192 -3416 1193 -3415
rect 1318 -3416 1319 -3415
rect 1332 -3416 1333 -3415
rect 1381 -3416 1382 -3415
rect 1384 -3416 1385 -3415
rect 282 -3418 283 -3417
rect 317 -3418 318 -3417
rect 324 -3418 325 -3417
rect 338 -3418 339 -3417
rect 352 -3418 353 -3417
rect 373 -3418 374 -3417
rect 394 -3418 395 -3417
rect 499 -3418 500 -3417
rect 513 -3418 514 -3417
rect 656 -3418 657 -3417
rect 702 -3418 703 -3417
rect 737 -3418 738 -3417
rect 793 -3418 794 -3417
rect 803 -3418 804 -3417
rect 863 -3418 864 -3417
rect 1265 -3418 1266 -3417
rect 1381 -3418 1382 -3417
rect 1388 -3418 1389 -3417
rect 366 -3420 367 -3419
rect 394 -3420 395 -3419
rect 415 -3420 416 -3419
rect 513 -3420 514 -3419
rect 520 -3420 521 -3419
rect 527 -3420 528 -3419
rect 562 -3420 563 -3419
rect 730 -3420 731 -3419
rect 733 -3420 734 -3419
rect 786 -3420 787 -3419
rect 800 -3420 801 -3419
rect 814 -3420 815 -3419
rect 842 -3420 843 -3419
rect 863 -3420 864 -3419
rect 884 -3420 885 -3419
rect 891 -3420 892 -3419
rect 898 -3420 899 -3419
rect 999 -3420 1000 -3419
rect 1017 -3420 1018 -3419
rect 1031 -3420 1032 -3419
rect 1080 -3420 1081 -3419
rect 1199 -3420 1200 -3419
rect 359 -3422 360 -3421
rect 520 -3422 521 -3421
rect 562 -3422 563 -3421
rect 590 -3422 591 -3421
rect 625 -3422 626 -3421
rect 730 -3422 731 -3421
rect 751 -3422 752 -3421
rect 884 -3422 885 -3421
rect 898 -3422 899 -3421
rect 905 -3422 906 -3421
rect 919 -3422 920 -3421
rect 989 -3422 990 -3421
rect 996 -3422 997 -3421
rect 1010 -3422 1011 -3421
rect 1024 -3422 1025 -3421
rect 1171 -3422 1172 -3421
rect 359 -3424 360 -3423
rect 509 -3424 510 -3423
rect 576 -3424 577 -3423
rect 597 -3424 598 -3423
rect 625 -3424 626 -3423
rect 646 -3424 647 -3423
rect 681 -3424 682 -3423
rect 737 -3424 738 -3423
rect 758 -3424 759 -3423
rect 786 -3424 787 -3423
rect 807 -3424 808 -3423
rect 842 -3424 843 -3423
rect 849 -3424 850 -3423
rect 891 -3424 892 -3423
rect 919 -3424 920 -3423
rect 961 -3424 962 -3423
rect 968 -3424 969 -3423
rect 1167 -3424 1168 -3423
rect 366 -3426 367 -3425
rect 387 -3426 388 -3425
rect 415 -3426 416 -3425
rect 436 -3426 437 -3425
rect 443 -3426 444 -3425
rect 586 -3426 587 -3425
rect 597 -3426 598 -3425
rect 695 -3426 696 -3425
rect 751 -3426 752 -3425
rect 849 -3426 850 -3425
rect 877 -3426 878 -3425
rect 1010 -3426 1011 -3425
rect 1031 -3426 1032 -3425
rect 1150 -3426 1151 -3425
rect 1153 -3426 1154 -3425
rect 1206 -3426 1207 -3425
rect 303 -3428 304 -3427
rect 443 -3428 444 -3427
rect 450 -3428 451 -3427
rect 478 -3428 479 -3427
rect 492 -3428 493 -3427
rect 604 -3428 605 -3427
rect 618 -3428 619 -3427
rect 695 -3428 696 -3427
rect 758 -3428 759 -3427
rect 821 -3428 822 -3427
rect 877 -3428 878 -3427
rect 894 -3428 895 -3427
rect 940 -3428 941 -3427
rect 1017 -3428 1018 -3427
rect 1087 -3428 1088 -3427
rect 1213 -3428 1214 -3427
rect 380 -3430 381 -3429
rect 387 -3430 388 -3429
rect 408 -3430 409 -3429
rect 436 -3430 437 -3429
rect 464 -3430 465 -3429
rect 527 -3430 528 -3429
rect 548 -3430 549 -3429
rect 807 -3430 808 -3429
rect 814 -3430 815 -3429
rect 828 -3430 829 -3429
rect 912 -3430 913 -3429
rect 940 -3430 941 -3429
rect 954 -3430 955 -3429
rect 982 -3430 983 -3429
rect 1003 -3430 1004 -3429
rect 1024 -3430 1025 -3429
rect 1101 -3430 1102 -3429
rect 1115 -3430 1116 -3429
rect 1122 -3430 1123 -3429
rect 1136 -3430 1137 -3429
rect 1157 -3430 1158 -3429
rect 1234 -3430 1235 -3429
rect 331 -3432 332 -3431
rect 380 -3432 381 -3431
rect 401 -3432 402 -3431
rect 464 -3432 465 -3431
rect 471 -3432 472 -3431
rect 478 -3432 479 -3431
rect 492 -3432 493 -3431
rect 534 -3432 535 -3431
rect 548 -3432 549 -3431
rect 555 -3432 556 -3431
rect 579 -3432 580 -3431
rect 1080 -3432 1081 -3431
rect 1094 -3432 1095 -3431
rect 1115 -3432 1116 -3431
rect 1129 -3432 1130 -3431
rect 1300 -3432 1301 -3431
rect 299 -3434 300 -3433
rect 401 -3434 402 -3433
rect 422 -3434 423 -3433
rect 523 -3434 524 -3433
rect 534 -3434 535 -3433
rect 541 -3434 542 -3433
rect 646 -3434 647 -3433
rect 660 -3434 661 -3433
rect 681 -3434 682 -3433
rect 709 -3434 710 -3433
rect 772 -3434 773 -3433
rect 905 -3434 906 -3433
rect 912 -3434 913 -3433
rect 926 -3434 927 -3433
rect 933 -3434 934 -3433
rect 954 -3434 955 -3433
rect 961 -3434 962 -3433
rect 975 -3434 976 -3433
rect 1003 -3434 1004 -3433
rect 1066 -3434 1067 -3433
rect 1136 -3434 1137 -3433
rect 1143 -3434 1144 -3433
rect 1206 -3434 1207 -3433
rect 1241 -3434 1242 -3433
rect 345 -3436 346 -3435
rect 422 -3436 423 -3435
rect 471 -3436 472 -3435
rect 541 -3436 542 -3435
rect 709 -3436 710 -3435
rect 744 -3436 745 -3435
rect 765 -3436 766 -3435
rect 975 -3436 976 -3435
rect 1384 -3436 1385 -3435
rect 1388 -3436 1389 -3435
rect 310 -3438 311 -3437
rect 345 -3438 346 -3437
rect 485 -3438 486 -3437
rect 660 -3438 661 -3437
rect 716 -3438 717 -3437
rect 765 -3438 766 -3437
rect 779 -3438 780 -3437
rect 793 -3438 794 -3437
rect 821 -3438 822 -3437
rect 1216 -3438 1217 -3437
rect 310 -3440 311 -3439
rect 352 -3440 353 -3439
rect 506 -3440 507 -3439
rect 555 -3440 556 -3439
rect 653 -3440 654 -3439
rect 779 -3440 780 -3439
rect 828 -3440 829 -3439
rect 835 -3440 836 -3439
rect 933 -3440 934 -3439
rect 996 -3440 997 -3439
rect 506 -3442 507 -3441
rect 621 -3442 622 -3441
rect 674 -3442 675 -3441
rect 716 -3442 717 -3441
rect 723 -3442 724 -3441
rect 772 -3442 773 -3441
rect 835 -3442 836 -3441
rect 947 -3442 948 -3441
rect 667 -3444 668 -3443
rect 674 -3444 675 -3443
rect 723 -3444 724 -3443
rect 852 -3444 853 -3443
rect 870 -3444 871 -3443
rect 947 -3444 948 -3443
rect 614 -3446 615 -3445
rect 667 -3446 668 -3445
rect 744 -3446 745 -3445
rect 856 -3446 857 -3445
rect 870 -3446 871 -3445
rect 1020 -3446 1021 -3445
rect 583 -3448 584 -3447
rect 856 -3448 857 -3447
rect 583 -3450 584 -3449
rect 926 -3450 927 -3449
rect 261 -3461 262 -3460
rect 268 -3461 269 -3460
rect 296 -3461 297 -3460
rect 310 -3461 311 -3460
rect 317 -3461 318 -3460
rect 355 -3461 356 -3460
rect 359 -3461 360 -3460
rect 411 -3461 412 -3460
rect 439 -3461 440 -3460
rect 656 -3461 657 -3460
rect 660 -3461 661 -3460
rect 733 -3461 734 -3460
rect 800 -3461 801 -3460
rect 807 -3461 808 -3460
rect 821 -3461 822 -3460
rect 828 -3461 829 -3460
rect 842 -3461 843 -3460
rect 915 -3461 916 -3460
rect 940 -3461 941 -3460
rect 943 -3461 944 -3460
rect 947 -3461 948 -3460
rect 1006 -3461 1007 -3460
rect 1010 -3461 1011 -3460
rect 1059 -3461 1060 -3460
rect 1066 -3461 1067 -3460
rect 1073 -3461 1074 -3460
rect 1087 -3461 1088 -3460
rect 1101 -3461 1102 -3460
rect 1115 -3461 1116 -3460
rect 1118 -3461 1119 -3460
rect 1143 -3461 1144 -3460
rect 1157 -3461 1158 -3460
rect 1181 -3461 1182 -3460
rect 1416 -3461 1417 -3460
rect 373 -3463 374 -3462
rect 390 -3463 391 -3462
rect 401 -3463 402 -3462
rect 583 -3463 584 -3462
rect 611 -3463 612 -3462
rect 719 -3463 720 -3462
rect 786 -3463 787 -3462
rect 800 -3463 801 -3462
rect 807 -3463 808 -3462
rect 814 -3463 815 -3462
rect 828 -3463 829 -3462
rect 870 -3463 871 -3462
rect 940 -3463 941 -3462
rect 961 -3463 962 -3462
rect 968 -3463 969 -3462
rect 982 -3463 983 -3462
rect 989 -3463 990 -3462
rect 1010 -3463 1011 -3462
rect 1017 -3463 1018 -3462
rect 1045 -3463 1046 -3462
rect 1073 -3463 1074 -3462
rect 1129 -3463 1130 -3462
rect 1185 -3463 1186 -3462
rect 1206 -3463 1207 -3462
rect 1213 -3463 1214 -3462
rect 1248 -3463 1249 -3462
rect 1269 -3463 1270 -3462
rect 1276 -3463 1277 -3462
rect 1297 -3463 1298 -3462
rect 1318 -3463 1319 -3462
rect 1374 -3463 1375 -3462
rect 1381 -3463 1382 -3462
rect 345 -3465 346 -3464
rect 373 -3465 374 -3464
rect 380 -3465 381 -3464
rect 408 -3465 409 -3464
rect 520 -3465 521 -3464
rect 590 -3465 591 -3464
rect 618 -3465 619 -3464
rect 625 -3465 626 -3464
rect 632 -3465 633 -3464
rect 663 -3465 664 -3464
rect 667 -3465 668 -3464
rect 754 -3465 755 -3464
rect 765 -3465 766 -3464
rect 786 -3465 787 -3464
rect 852 -3465 853 -3464
rect 919 -3465 920 -3464
rect 954 -3465 955 -3464
rect 961 -3465 962 -3464
rect 975 -3465 976 -3464
rect 1038 -3465 1039 -3464
rect 1080 -3465 1081 -3464
rect 1269 -3465 1270 -3464
rect 1300 -3465 1301 -3464
rect 1304 -3465 1305 -3464
rect 1346 -3465 1347 -3464
rect 1381 -3465 1382 -3464
rect 366 -3467 367 -3466
rect 380 -3467 381 -3466
rect 387 -3467 388 -3466
rect 425 -3467 426 -3466
rect 506 -3467 507 -3466
rect 590 -3467 591 -3466
rect 618 -3467 619 -3466
rect 723 -3467 724 -3466
rect 758 -3467 759 -3466
rect 765 -3467 766 -3466
rect 772 -3467 773 -3466
rect 814 -3467 815 -3466
rect 856 -3467 857 -3466
rect 947 -3467 948 -3466
rect 975 -3467 976 -3466
rect 1003 -3467 1004 -3466
rect 1115 -3467 1116 -3466
rect 1122 -3467 1123 -3466
rect 1199 -3467 1200 -3466
rect 1234 -3467 1235 -3466
rect 338 -3469 339 -3468
rect 366 -3469 367 -3468
rect 450 -3469 451 -3468
rect 506 -3469 507 -3468
rect 527 -3469 528 -3468
rect 621 -3469 622 -3468
rect 653 -3469 654 -3468
rect 681 -3469 682 -3468
rect 695 -3469 696 -3468
rect 758 -3469 759 -3468
rect 891 -3469 892 -3468
rect 919 -3469 920 -3468
rect 926 -3469 927 -3468
rect 1080 -3469 1081 -3468
rect 1118 -3469 1119 -3468
rect 1122 -3469 1123 -3468
rect 429 -3471 430 -3470
rect 450 -3471 451 -3470
rect 499 -3471 500 -3470
rect 527 -3471 528 -3470
rect 534 -3471 535 -3470
rect 632 -3471 633 -3470
rect 653 -3471 654 -3470
rect 1090 -3471 1091 -3470
rect 394 -3473 395 -3472
rect 429 -3473 430 -3472
rect 457 -3473 458 -3472
rect 499 -3473 500 -3472
rect 534 -3473 535 -3472
rect 607 -3473 608 -3472
rect 695 -3473 696 -3472
rect 744 -3473 745 -3472
rect 884 -3473 885 -3472
rect 891 -3473 892 -3472
rect 905 -3473 906 -3472
rect 926 -3473 927 -3472
rect 1003 -3473 1004 -3472
rect 1178 -3473 1179 -3472
rect 436 -3475 437 -3474
rect 457 -3475 458 -3474
rect 541 -3475 542 -3474
rect 586 -3475 587 -3474
rect 702 -3475 703 -3474
rect 716 -3475 717 -3474
rect 723 -3475 724 -3474
rect 751 -3475 752 -3474
rect 863 -3475 864 -3474
rect 884 -3475 885 -3474
rect 898 -3475 899 -3474
rect 905 -3475 906 -3474
rect 478 -3477 479 -3476
rect 541 -3477 542 -3476
rect 548 -3477 549 -3476
rect 593 -3477 594 -3476
rect 688 -3477 689 -3476
rect 702 -3477 703 -3476
rect 709 -3477 710 -3476
rect 821 -3477 822 -3476
rect 898 -3477 899 -3476
rect 912 -3477 913 -3476
rect 464 -3479 465 -3478
rect 478 -3479 479 -3478
rect 548 -3479 549 -3478
rect 576 -3479 577 -3478
rect 646 -3479 647 -3478
rect 709 -3479 710 -3478
rect 730 -3479 731 -3478
rect 772 -3479 773 -3478
rect 779 -3479 780 -3478
rect 912 -3479 913 -3478
rect 555 -3481 556 -3480
rect 583 -3481 584 -3480
rect 674 -3481 675 -3480
rect 688 -3481 689 -3480
rect 730 -3481 731 -3480
rect 835 -3481 836 -3480
rect 492 -3483 493 -3482
rect 555 -3483 556 -3482
rect 562 -3483 563 -3482
rect 576 -3483 577 -3482
rect 744 -3483 745 -3482
rect 996 -3483 997 -3482
rect 443 -3485 444 -3484
rect 492 -3485 493 -3484
rect 513 -3485 514 -3484
rect 562 -3485 563 -3484
rect 569 -3485 570 -3484
rect 646 -3485 647 -3484
rect 996 -3485 997 -3484
rect 1031 -3485 1032 -3484
rect 415 -3487 416 -3486
rect 443 -3487 444 -3486
rect 569 -3487 570 -3486
rect 597 -3487 598 -3486
rect 422 -3489 423 -3488
rect 513 -3489 514 -3488
rect 422 -3491 423 -3490
rect 471 -3491 472 -3490
rect 268 -3502 269 -3501
rect 282 -3502 283 -3501
rect 285 -3502 286 -3501
rect 296 -3502 297 -3501
rect 366 -3502 367 -3501
rect 387 -3502 388 -3501
rect 390 -3502 391 -3501
rect 394 -3502 395 -3501
rect 408 -3502 409 -3501
rect 439 -3502 440 -3501
rect 450 -3502 451 -3501
rect 481 -3502 482 -3501
rect 506 -3502 507 -3501
rect 565 -3502 566 -3501
rect 583 -3502 584 -3501
rect 597 -3502 598 -3501
rect 632 -3502 633 -3501
rect 726 -3502 727 -3501
rect 733 -3502 734 -3501
rect 1181 -3502 1182 -3501
rect 1234 -3502 1235 -3501
rect 1279 -3502 1280 -3501
rect 1374 -3502 1375 -3501
rect 1381 -3502 1382 -3501
rect 1384 -3502 1385 -3501
rect 1388 -3502 1389 -3501
rect 1416 -3502 1417 -3501
rect 1500 -3502 1501 -3501
rect 373 -3504 374 -3503
rect 401 -3504 402 -3503
rect 443 -3504 444 -3503
rect 450 -3504 451 -3503
rect 457 -3504 458 -3503
rect 464 -3504 465 -3503
rect 492 -3504 493 -3503
rect 506 -3504 507 -3503
rect 520 -3504 521 -3503
rect 548 -3504 549 -3503
rect 562 -3504 563 -3503
rect 583 -3504 584 -3503
rect 590 -3504 591 -3503
rect 656 -3504 657 -3503
rect 674 -3504 675 -3503
rect 695 -3504 696 -3503
rect 737 -3504 738 -3503
rect 754 -3504 755 -3503
rect 758 -3504 759 -3503
rect 779 -3504 780 -3503
rect 786 -3504 787 -3503
rect 789 -3504 790 -3503
rect 821 -3504 822 -3503
rect 863 -3504 864 -3503
rect 905 -3504 906 -3503
rect 912 -3504 913 -3503
rect 947 -3504 948 -3503
rect 1034 -3504 1035 -3503
rect 1045 -3504 1046 -3503
rect 1048 -3504 1049 -3503
rect 1059 -3504 1060 -3503
rect 1090 -3504 1091 -3503
rect 1122 -3504 1123 -3503
rect 1129 -3504 1130 -3503
rect 1157 -3504 1158 -3503
rect 1164 -3504 1165 -3503
rect 1178 -3504 1179 -3503
rect 1185 -3504 1186 -3503
rect 1248 -3504 1249 -3503
rect 1262 -3504 1263 -3503
rect 1269 -3504 1270 -3503
rect 1339 -3504 1340 -3503
rect 429 -3506 430 -3505
rect 443 -3506 444 -3505
rect 478 -3506 479 -3505
rect 492 -3506 493 -3505
rect 527 -3506 528 -3505
rect 558 -3506 559 -3505
rect 576 -3506 577 -3505
rect 590 -3506 591 -3505
rect 646 -3506 647 -3505
rect 730 -3506 731 -3505
rect 758 -3506 759 -3505
rect 772 -3506 773 -3505
rect 786 -3506 787 -3505
rect 793 -3506 794 -3505
rect 800 -3506 801 -3505
rect 821 -3506 822 -3505
rect 842 -3506 843 -3505
rect 1017 -3506 1018 -3505
rect 1020 -3506 1021 -3505
rect 1073 -3506 1074 -3505
rect 1080 -3506 1081 -3505
rect 1143 -3506 1144 -3505
rect 429 -3508 430 -3507
rect 478 -3508 479 -3507
rect 499 -3508 500 -3507
rect 527 -3508 528 -3507
rect 541 -3508 542 -3507
rect 548 -3508 549 -3507
rect 576 -3508 577 -3507
rect 618 -3508 619 -3507
rect 639 -3508 640 -3507
rect 646 -3508 647 -3507
rect 653 -3508 654 -3507
rect 744 -3508 745 -3507
rect 765 -3508 766 -3507
rect 772 -3508 773 -3507
rect 800 -3508 801 -3507
rect 807 -3508 808 -3507
rect 884 -3508 885 -3507
rect 905 -3508 906 -3507
rect 957 -3508 958 -3507
rect 996 -3508 997 -3507
rect 1010 -3508 1011 -3507
rect 1041 -3508 1042 -3507
rect 1045 -3508 1046 -3507
rect 1052 -3508 1053 -3507
rect 1062 -3508 1063 -3507
rect 1066 -3508 1067 -3507
rect 485 -3510 486 -3509
rect 499 -3510 500 -3509
rect 513 -3510 514 -3509
rect 541 -3510 542 -3509
rect 688 -3510 689 -3509
rect 695 -3510 696 -3509
rect 709 -3510 710 -3509
rect 730 -3510 731 -3509
rect 807 -3510 808 -3509
rect 814 -3510 815 -3509
rect 877 -3510 878 -3509
rect 884 -3510 885 -3509
rect 961 -3510 962 -3509
rect 964 -3510 965 -3509
rect 968 -3510 969 -3509
rect 975 -3510 976 -3509
rect 1024 -3510 1025 -3509
rect 1031 -3510 1032 -3509
rect 1038 -3510 1039 -3509
rect 1073 -3510 1074 -3509
rect 471 -3512 472 -3511
rect 485 -3512 486 -3511
rect 513 -3512 514 -3511
rect 534 -3512 535 -3511
rect 709 -3512 710 -3511
rect 716 -3512 717 -3511
rect 765 -3512 766 -3511
rect 1038 -3512 1039 -3511
rect 1048 -3512 1049 -3511
rect 1052 -3512 1053 -3511
rect 534 -3514 535 -3513
rect 569 -3514 570 -3513
rect 814 -3514 815 -3513
rect 828 -3514 829 -3513
rect 877 -3514 878 -3513
rect 898 -3514 899 -3513
rect 954 -3514 955 -3513
rect 961 -3514 962 -3513
rect 555 -3516 556 -3515
rect 569 -3516 570 -3515
rect 891 -3516 892 -3515
rect 898 -3516 899 -3515
rect 926 -3516 927 -3515
rect 954 -3516 955 -3515
rect 926 -3518 927 -3517
rect 933 -3518 934 -3517
rect 919 -3520 920 -3519
rect 933 -3520 934 -3519
rect 919 -3522 920 -3521
rect 947 -3522 948 -3521
rect 387 -3533 388 -3532
rect 390 -3533 391 -3532
rect 408 -3533 409 -3532
rect 429 -3533 430 -3532
rect 450 -3533 451 -3532
rect 457 -3533 458 -3532
rect 464 -3533 465 -3532
rect 474 -3533 475 -3532
rect 506 -3533 507 -3532
rect 520 -3533 521 -3532
rect 558 -3533 559 -3532
rect 1108 -3533 1109 -3532
rect 1157 -3533 1158 -3532
rect 1164 -3533 1165 -3532
rect 1262 -3533 1263 -3532
rect 1279 -3533 1280 -3532
rect 1339 -3533 1340 -3532
rect 1360 -3533 1361 -3532
rect 1381 -3533 1382 -3532
rect 1388 -3533 1389 -3532
rect 1500 -3533 1501 -3532
rect 1580 -3533 1581 -3532
rect 387 -3535 388 -3534
rect 401 -3535 402 -3534
rect 443 -3535 444 -3534
rect 450 -3535 451 -3534
rect 506 -3535 507 -3534
rect 513 -3535 514 -3534
rect 565 -3535 566 -3534
rect 653 -3535 654 -3534
rect 660 -3535 661 -3534
rect 674 -3535 675 -3534
rect 695 -3535 696 -3534
rect 705 -3535 706 -3534
rect 730 -3535 731 -3534
rect 737 -3535 738 -3534
rect 796 -3535 797 -3534
rect 800 -3535 801 -3534
rect 807 -3535 808 -3534
rect 824 -3535 825 -3534
rect 884 -3535 885 -3534
rect 891 -3535 892 -3534
rect 926 -3535 927 -3534
rect 950 -3535 951 -3534
rect 957 -3535 958 -3534
rect 968 -3535 969 -3534
rect 1038 -3535 1039 -3534
rect 1045 -3535 1046 -3534
rect 1052 -3535 1053 -3534
rect 1059 -3535 1060 -3534
rect 1073 -3535 1074 -3534
rect 1111 -3535 1112 -3534
rect 1143 -3535 1144 -3534
rect 1164 -3535 1165 -3534
rect 394 -3537 395 -3536
rect 401 -3537 402 -3536
rect 499 -3537 500 -3536
rect 513 -3537 514 -3536
rect 565 -3537 566 -3536
rect 576 -3537 577 -3536
rect 604 -3537 605 -3536
rect 607 -3537 608 -3536
rect 646 -3537 647 -3536
rect 663 -3537 664 -3536
rect 667 -3537 668 -3536
rect 765 -3537 766 -3536
rect 779 -3537 780 -3536
rect 800 -3537 801 -3536
rect 877 -3537 878 -3536
rect 884 -3537 885 -3536
rect 919 -3537 920 -3536
rect 926 -3537 927 -3536
rect 933 -3537 934 -3536
rect 936 -3537 937 -3536
rect 390 -3539 391 -3538
rect 394 -3539 395 -3538
rect 492 -3539 493 -3538
rect 499 -3539 500 -3538
rect 576 -3539 577 -3538
rect 590 -3539 591 -3538
rect 702 -3539 703 -3538
rect 709 -3539 710 -3538
rect 772 -3539 773 -3538
rect 779 -3539 780 -3538
rect 793 -3539 794 -3538
rect 807 -3539 808 -3538
rect 863 -3539 864 -3538
rect 877 -3539 878 -3538
rect 485 -3541 486 -3540
rect 492 -3541 493 -3540
rect 590 -3541 591 -3540
rect 597 -3541 598 -3540
rect 772 -3541 773 -3540
rect 842 -3541 843 -3540
rect 583 -3543 584 -3542
rect 597 -3543 598 -3542
rect 555 -3545 556 -3544
rect 583 -3545 584 -3544
rect 541 -3547 542 -3546
rect 555 -3547 556 -3546
rect 534 -3549 535 -3548
rect 541 -3549 542 -3548
rect 534 -3551 535 -3550
rect 562 -3551 563 -3550
rect 401 -3562 402 -3561
rect 404 -3562 405 -3561
rect 457 -3562 458 -3561
rect 464 -3562 465 -3561
rect 474 -3562 475 -3561
rect 478 -3562 479 -3561
rect 499 -3562 500 -3561
rect 513 -3562 514 -3561
rect 527 -3562 528 -3561
rect 541 -3562 542 -3561
rect 555 -3562 556 -3561
rect 562 -3562 563 -3561
rect 569 -3562 570 -3561
rect 576 -3562 577 -3561
rect 579 -3562 580 -3561
rect 597 -3562 598 -3561
rect 632 -3562 633 -3561
rect 667 -3562 668 -3561
rect 702 -3562 703 -3561
rect 709 -3562 710 -3561
rect 737 -3562 738 -3561
rect 747 -3562 748 -3561
rect 758 -3562 759 -3561
rect 765 -3562 766 -3561
rect 768 -3562 769 -3561
rect 779 -3562 780 -3561
rect 786 -3562 787 -3561
rect 796 -3562 797 -3561
rect 877 -3562 878 -3561
rect 894 -3562 895 -3561
rect 901 -3562 902 -3561
rect 905 -3562 906 -3561
rect 926 -3562 927 -3561
rect 950 -3562 951 -3561
rect 1111 -3562 1112 -3561
rect 1115 -3562 1116 -3561
rect 1132 -3562 1133 -3561
rect 1136 -3562 1137 -3561
rect 1164 -3562 1165 -3561
rect 1171 -3562 1172 -3561
rect 1178 -3562 1179 -3561
rect 1185 -3562 1186 -3561
rect 1192 -3562 1193 -3561
rect 1199 -3562 1200 -3561
rect 1391 -3562 1392 -3561
rect 1395 -3562 1396 -3561
rect 380 -3564 381 -3563
rect 401 -3564 402 -3563
rect 450 -3564 451 -3563
rect 457 -3564 458 -3563
rect 502 -3564 503 -3563
rect 506 -3564 507 -3563
rect 530 -3564 531 -3563
rect 534 -3564 535 -3563
rect 548 -3564 549 -3563
rect 562 -3564 563 -3563
rect 576 -3564 577 -3563
rect 583 -3564 584 -3563
rect 758 -3564 759 -3563
rect 772 -3564 773 -3563
rect 793 -3564 794 -3563
rect 807 -3564 808 -3563
rect 891 -3564 892 -3563
rect 898 -3564 899 -3563
rect 933 -3564 934 -3563
rect 940 -3564 941 -3563
rect 1129 -3564 1130 -3563
rect 1136 -3564 1137 -3563
rect 1388 -3564 1389 -3563
rect 1395 -3564 1396 -3563
rect 807 -3566 808 -3565
rect 814 -3566 815 -3565
rect 1360 -3566 1361 -3565
rect 1388 -3566 1389 -3565
rect 387 -3577 388 -3576
rect 401 -3577 402 -3576
rect 457 -3577 458 -3576
rect 464 -3577 465 -3576
rect 492 -3577 493 -3576
rect 502 -3577 503 -3576
rect 562 -3577 563 -3576
rect 579 -3577 580 -3576
rect 590 -3577 591 -3576
rect 597 -3577 598 -3576
rect 600 -3577 601 -3576
rect 632 -3577 633 -3576
rect 747 -3577 748 -3576
rect 758 -3577 759 -3576
rect 800 -3577 801 -3576
rect 810 -3577 811 -3576
rect 884 -3577 885 -3576
rect 898 -3577 899 -3576
rect 1129 -3577 1130 -3576
rect 1136 -3577 1137 -3576
rect 1171 -3577 1172 -3576
rect 1181 -3577 1182 -3576
rect 1195 -3577 1196 -3576
rect 1199 -3577 1200 -3576
rect 1388 -3577 1389 -3576
rect 1395 -3577 1396 -3576
rect 397 -3579 398 -3578
rect 408 -3579 409 -3578
rect 1178 -3579 1179 -3578
rect 1185 -3579 1186 -3578
<< metal2 >>
rect 233 -13 234 1
rect 436 -13 437 1
rect 443 -13 444 1
rect 457 -13 458 1
rect 527 -13 528 1
rect 548 -13 549 1
rect 555 -13 556 1
rect 754 -13 755 1
rect 877 -13 878 1
rect 954 -13 955 1
rect 345 -13 346 -1
rect 352 -13 353 -1
rect 359 -13 360 -1
rect 467 -13 468 -1
rect 604 -13 605 -1
rect 614 -13 615 -1
rect 653 -13 654 -1
rect 677 -13 678 -1
rect 716 -13 717 -1
rect 800 -13 801 -1
rect 380 -13 381 -3
rect 534 -13 535 -3
rect 670 -13 671 -3
rect 688 -13 689 -3
rect 401 -13 402 -5
rect 460 -13 461 -5
rect 408 -13 409 -7
rect 432 -13 433 -7
rect 453 -13 454 -7
rect 471 -13 472 -7
rect 415 -13 416 -9
rect 506 -13 507 -9
rect 422 -13 423 -11
rect 450 -13 451 -11
rect 145 -50 146 -22
rect 149 -50 150 -22
rect 156 -50 157 -22
rect 233 -23 234 -21
rect 261 -50 262 -22
rect 306 -50 307 -22
rect 324 -50 325 -22
rect 359 -23 360 -21
rect 373 -50 374 -22
rect 408 -23 409 -21
rect 425 -50 426 -22
rect 443 -23 444 -21
rect 450 -50 451 -22
rect 555 -23 556 -21
rect 590 -50 591 -22
rect 821 -50 822 -22
rect 842 -50 843 -22
rect 884 -50 885 -22
rect 954 -23 955 -21
rect 989 -50 990 -22
rect 226 -50 227 -24
rect 236 -50 237 -24
rect 282 -50 283 -24
rect 390 -50 391 -24
rect 394 -50 395 -24
rect 415 -25 416 -21
rect 429 -50 430 -24
rect 443 -50 444 -24
rect 460 -25 461 -21
rect 555 -50 556 -24
rect 604 -25 605 -21
rect 604 -50 605 -24
rect 604 -25 605 -21
rect 604 -50 605 -24
rect 618 -50 619 -24
rect 632 -50 633 -24
rect 653 -25 654 -21
rect 667 -50 668 -24
rect 677 -25 678 -21
rect 681 -50 682 -24
rect 688 -25 689 -21
rect 702 -50 703 -24
rect 712 -50 713 -24
rect 772 -50 773 -24
rect 800 -25 801 -21
rect 828 -50 829 -24
rect 331 -50 332 -26
rect 380 -27 381 -21
rect 408 -50 409 -26
rect 562 -50 563 -26
rect 653 -50 654 -26
rect 670 -27 671 -21
rect 677 -50 678 -26
rect 730 -50 731 -26
rect 751 -27 752 -21
rect 996 -50 997 -26
rect 338 -50 339 -28
rect 345 -29 346 -21
rect 380 -50 381 -28
rect 401 -29 402 -21
rect 436 -29 437 -21
rect 660 -50 661 -28
rect 688 -50 689 -28
rect 719 -29 720 -21
rect 758 -50 759 -28
rect 898 -50 899 -28
rect 401 -50 402 -30
rect 422 -31 423 -21
rect 432 -31 433 -21
rect 436 -50 437 -30
rect 460 -50 461 -30
rect 744 -50 745 -30
rect 814 -50 815 -30
rect 880 -31 881 -21
rect 464 -33 465 -21
rect 597 -50 598 -32
rect 716 -50 717 -32
rect 754 -33 755 -21
rect 471 -35 472 -21
rect 478 -50 479 -34
rect 492 -50 493 -34
rect 506 -50 507 -34
rect 509 -35 510 -21
rect 611 -50 612 -34
rect 471 -50 472 -36
rect 516 -50 517 -36
rect 520 -50 521 -36
rect 639 -50 640 -36
rect 495 -50 496 -38
rect 499 -50 500 -38
rect 513 -50 514 -38
rect 625 -50 626 -38
rect 523 -50 524 -40
rect 541 -50 542 -40
rect 551 -41 552 -21
rect 576 -50 577 -40
rect 530 -50 531 -42
rect 548 -50 549 -42
rect 534 -45 535 -21
rect 646 -50 647 -44
rect 527 -47 528 -21
rect 534 -50 535 -46
rect 537 -47 538 -21
rect 583 -50 584 -46
rect 464 -50 465 -48
rect 527 -50 528 -48
rect 128 -97 129 -59
rect 156 -60 157 -58
rect 191 -97 192 -59
rect 198 -97 199 -59
rect 205 -97 206 -59
rect 226 -60 227 -58
rect 254 -97 255 -59
rect 432 -97 433 -59
rect 474 -97 475 -59
rect 737 -97 738 -59
rect 744 -60 745 -58
rect 870 -97 871 -59
rect 884 -60 885 -58
rect 940 -97 941 -59
rect 989 -60 990 -58
rect 1010 -97 1011 -59
rect 149 -62 150 -58
rect 149 -97 150 -61
rect 149 -62 150 -58
rect 149 -97 150 -61
rect 219 -97 220 -61
rect 282 -62 283 -58
rect 289 -97 290 -61
rect 324 -62 325 -58
rect 345 -97 346 -61
rect 422 -62 423 -58
rect 478 -62 479 -58
rect 488 -97 489 -61
rect 492 -97 493 -61
rect 709 -62 710 -58
rect 716 -62 717 -58
rect 744 -97 745 -61
rect 751 -97 752 -61
rect 887 -97 888 -61
rect 898 -62 899 -58
rect 954 -97 955 -61
rect 996 -62 997 -58
rect 1087 -97 1088 -61
rect 261 -64 262 -58
rect 268 -97 269 -63
rect 275 -97 276 -63
rect 457 -64 458 -58
rect 478 -97 479 -63
rect 590 -64 591 -58
rect 625 -64 626 -58
rect 695 -97 696 -63
rect 730 -64 731 -58
rect 786 -97 787 -63
rect 796 -97 797 -63
rect 863 -97 864 -63
rect 936 -64 937 -58
rect 947 -97 948 -63
rect 247 -97 248 -65
rect 261 -97 262 -65
rect 282 -97 283 -65
rect 460 -66 461 -58
rect 506 -66 507 -58
rect 520 -97 521 -65
rect 551 -97 552 -65
rect 677 -66 678 -58
rect 688 -66 689 -58
rect 716 -97 717 -65
rect 772 -66 773 -58
rect 835 -97 836 -65
rect 296 -97 297 -67
rect 408 -68 409 -58
rect 422 -97 423 -67
rect 436 -68 437 -58
rect 506 -97 507 -67
rect 593 -68 594 -58
rect 625 -97 626 -67
rect 810 -97 811 -67
rect 817 -97 818 -67
rect 856 -97 857 -67
rect 303 -97 304 -69
rect 338 -70 339 -58
rect 352 -97 353 -69
rect 415 -70 416 -58
rect 555 -70 556 -58
rect 674 -97 675 -69
rect 702 -70 703 -58
rect 730 -97 731 -69
rect 779 -97 780 -69
rect 884 -97 885 -69
rect 306 -72 307 -58
rect 359 -97 360 -71
rect 366 -97 367 -71
rect 401 -72 402 -58
rect 415 -97 416 -71
rect 516 -72 517 -58
rect 555 -97 556 -71
rect 576 -72 577 -58
rect 583 -72 584 -58
rect 688 -97 689 -71
rect 800 -97 801 -71
rect 828 -72 829 -58
rect 310 -97 311 -73
rect 450 -74 451 -58
rect 530 -97 531 -73
rect 583 -97 584 -73
rect 590 -97 591 -73
rect 618 -74 619 -58
rect 646 -74 647 -58
rect 709 -97 710 -73
rect 807 -97 808 -73
rect 842 -74 843 -58
rect 317 -97 318 -75
rect 331 -76 332 -58
rect 338 -97 339 -75
rect 464 -76 465 -58
rect 541 -76 542 -58
rect 576 -97 577 -75
rect 597 -76 598 -58
rect 702 -97 703 -75
rect 712 -76 713 -58
rect 842 -97 843 -75
rect 324 -97 325 -77
rect 373 -78 374 -58
rect 376 -97 377 -77
rect 380 -78 381 -58
rect 387 -78 388 -58
rect 436 -97 437 -77
rect 464 -97 465 -77
rect 471 -78 472 -58
rect 499 -78 500 -58
rect 541 -97 542 -77
rect 604 -78 605 -58
rect 618 -97 619 -77
rect 649 -97 650 -77
rect 793 -97 794 -77
rect 814 -78 815 -58
rect 828 -97 829 -77
rect 331 -97 332 -79
rect 443 -97 444 -79
rect 534 -80 535 -58
rect 597 -97 598 -79
rect 660 -80 661 -58
rect 723 -97 724 -79
rect 821 -80 822 -58
rect 891 -97 892 -79
rect 334 -97 335 -81
rect 499 -97 500 -81
rect 513 -97 514 -81
rect 534 -97 535 -81
rect 569 -82 570 -58
rect 604 -97 605 -81
rect 611 -82 612 -58
rect 660 -97 661 -81
rect 373 -97 374 -83
rect 380 -97 381 -83
rect 387 -97 388 -83
rect 523 -84 524 -58
rect 548 -84 549 -58
rect 569 -97 570 -83
rect 632 -97 633 -83
rect 821 -97 822 -83
rect 394 -86 395 -58
rect 394 -97 395 -85
rect 394 -86 395 -58
rect 394 -97 395 -85
rect 401 -97 402 -85
rect 429 -86 430 -58
rect 562 -86 563 -58
rect 611 -97 612 -85
rect 411 -97 412 -87
rect 450 -97 451 -87
rect 562 -97 563 -87
rect 653 -88 654 -58
rect 653 -97 654 -89
rect 667 -90 668 -58
rect 667 -97 668 -91
rect 681 -92 682 -58
rect 639 -94 640 -58
rect 681 -97 682 -93
rect 639 -97 640 -95
rect 758 -96 759 -58
rect 89 -107 90 -105
rect 93 -166 94 -106
rect 114 -166 115 -106
rect 128 -107 129 -105
rect 135 -166 136 -106
rect 219 -107 220 -105
rect 226 -166 227 -106
rect 292 -107 293 -105
rect 324 -107 325 -105
rect 324 -166 325 -106
rect 324 -107 325 -105
rect 324 -166 325 -106
rect 345 -107 346 -105
rect 362 -166 363 -106
rect 373 -107 374 -105
rect 394 -107 395 -105
rect 408 -107 409 -105
rect 467 -166 468 -106
rect 471 -107 472 -105
rect 488 -107 489 -105
rect 513 -107 514 -105
rect 548 -107 549 -105
rect 583 -107 584 -105
rect 583 -166 584 -106
rect 583 -107 584 -105
rect 583 -166 584 -106
rect 611 -107 612 -105
rect 646 -107 647 -105
rect 656 -166 657 -106
rect 744 -107 745 -105
rect 793 -107 794 -105
rect 821 -166 822 -106
rect 828 -107 829 -105
rect 912 -166 913 -106
rect 940 -107 941 -105
rect 996 -166 997 -106
rect 1010 -107 1011 -105
rect 1038 -166 1039 -106
rect 1087 -107 1088 -105
rect 1129 -166 1130 -106
rect 1195 -166 1196 -106
rect 1220 -166 1221 -106
rect 142 -166 143 -108
rect 254 -109 255 -105
rect 261 -109 262 -105
rect 471 -166 472 -108
rect 481 -166 482 -108
rect 551 -109 552 -105
rect 646 -166 647 -108
rect 716 -109 717 -105
rect 723 -109 724 -105
rect 849 -166 850 -108
rect 856 -109 857 -105
rect 898 -166 899 -108
rect 947 -109 948 -105
rect 968 -166 969 -108
rect 149 -111 150 -105
rect 149 -166 150 -110
rect 149 -111 150 -105
rect 149 -166 150 -110
rect 156 -166 157 -110
rect 331 -111 332 -105
rect 380 -111 381 -105
rect 383 -123 384 -110
rect 394 -166 395 -110
rect 639 -111 640 -105
rect 674 -111 675 -105
rect 758 -166 759 -110
rect 810 -111 811 -105
rect 940 -166 941 -110
rect 954 -111 955 -105
rect 982 -166 983 -110
rect 163 -166 164 -112
rect 205 -113 206 -105
rect 219 -166 220 -112
rect 303 -113 304 -105
rect 310 -113 311 -105
rect 373 -166 374 -112
rect 380 -166 381 -112
rect 443 -113 444 -105
rect 450 -113 451 -105
rect 457 -113 458 -105
rect 485 -113 486 -105
rect 509 -166 510 -112
rect 513 -166 514 -112
rect 933 -166 934 -112
rect 170 -166 171 -114
rect 355 -166 356 -114
rect 376 -115 377 -105
rect 485 -166 486 -114
rect 530 -115 531 -105
rect 548 -166 549 -114
rect 576 -115 577 -105
rect 639 -166 640 -114
rect 681 -115 682 -105
rect 723 -166 724 -114
rect 744 -166 745 -114
rect 800 -115 801 -105
rect 817 -115 818 -105
rect 828 -166 829 -114
rect 835 -115 836 -105
rect 919 -166 920 -114
rect 177 -166 178 -116
rect 338 -117 339 -105
rect 352 -117 353 -105
rect 457 -166 458 -116
rect 537 -117 538 -105
rect 625 -117 626 -105
rect 660 -117 661 -105
rect 800 -166 801 -116
rect 824 -117 825 -105
rect 1010 -166 1011 -116
rect 184 -166 185 -118
rect 191 -119 192 -105
rect 198 -166 199 -118
rect 247 -119 248 -105
rect 250 -119 251 -105
rect 310 -166 311 -118
rect 317 -119 318 -105
rect 331 -166 332 -118
rect 338 -166 339 -118
rect 632 -119 633 -105
rect 698 -166 699 -118
rect 905 -166 906 -118
rect 191 -166 192 -120
rect 275 -121 276 -105
rect 289 -166 290 -120
rect 429 -166 430 -120
rect 450 -166 451 -120
rect 502 -166 503 -120
rect 576 -166 577 -120
rect 653 -121 654 -105
rect 709 -121 710 -105
rect 807 -166 808 -120
rect 842 -121 843 -105
rect 961 -166 962 -120
rect 208 -166 209 -122
rect 317 -166 318 -122
rect 443 -166 444 -122
rect 460 -123 461 -105
rect 632 -166 633 -122
rect 716 -166 717 -122
rect 768 -166 769 -122
rect 779 -123 780 -105
rect 835 -166 836 -122
rect 856 -166 857 -122
rect 877 -166 878 -122
rect 880 -166 881 -122
rect 926 -166 927 -122
rect 243 -166 244 -124
rect 345 -166 346 -124
rect 408 -166 409 -124
rect 422 -125 423 -105
rect 590 -125 591 -105
rect 674 -166 675 -124
rect 796 -125 797 -105
rect 842 -166 843 -124
rect 863 -125 864 -105
rect 954 -166 955 -124
rect 247 -166 248 -126
rect 520 -127 521 -105
rect 569 -127 570 -105
rect 590 -166 591 -126
rect 597 -127 598 -105
rect 681 -166 682 -126
rect 814 -127 815 -105
rect 863 -166 864 -126
rect 870 -127 871 -105
rect 975 -166 976 -126
rect 254 -166 255 -128
rect 282 -129 283 -105
rect 296 -129 297 -105
rect 422 -166 423 -128
rect 432 -129 433 -105
rect 597 -166 598 -128
rect 611 -166 612 -128
rect 660 -166 661 -128
rect 737 -129 738 -105
rect 814 -166 815 -128
rect 884 -129 885 -105
rect 1136 -166 1137 -128
rect 261 -166 262 -130
rect 474 -131 475 -105
rect 520 -166 521 -130
rect 947 -166 948 -130
rect 268 -133 269 -105
rect 303 -166 304 -132
rect 432 -166 433 -132
rect 464 -133 465 -105
rect 618 -133 619 -105
rect 709 -166 710 -132
rect 786 -133 787 -105
rect 870 -166 871 -132
rect 891 -133 892 -105
rect 891 -166 892 -132
rect 891 -133 892 -105
rect 891 -166 892 -132
rect 268 -166 269 -134
rect 366 -135 367 -105
rect 415 -135 416 -105
rect 464 -166 465 -134
rect 618 -166 619 -134
rect 751 -135 752 -105
rect 275 -166 276 -136
rect 562 -137 563 -105
rect 625 -166 626 -136
rect 667 -137 668 -105
rect 688 -137 689 -105
rect 751 -166 752 -136
rect 282 -166 283 -138
rect 387 -139 388 -105
rect 401 -139 402 -105
rect 415 -166 416 -138
rect 534 -139 535 -105
rect 562 -166 563 -138
rect 649 -139 650 -105
rect 779 -166 780 -138
rect 296 -166 297 -140
rect 478 -141 479 -105
rect 534 -166 535 -140
rect 555 -141 556 -105
rect 667 -166 668 -140
rect 793 -166 794 -140
rect 366 -166 367 -142
rect 653 -166 654 -142
rect 702 -143 703 -105
rect 737 -166 738 -142
rect 352 -166 353 -144
rect 702 -166 703 -144
rect 730 -145 731 -105
rect 786 -166 787 -144
rect 387 -166 388 -146
rect 436 -147 437 -105
rect 478 -166 479 -146
rect 569 -166 570 -146
rect 695 -147 696 -105
rect 730 -166 731 -146
rect 401 -166 402 -148
rect 527 -149 528 -105
rect 359 -151 360 -105
rect 527 -166 528 -150
rect 359 -166 360 -152
rect 772 -166 773 -152
rect 436 -166 437 -154
rect 541 -155 542 -105
rect 492 -157 493 -105
rect 555 -166 556 -156
rect 492 -166 493 -158
rect 506 -159 507 -105
rect 541 -166 542 -158
rect 604 -159 605 -105
rect 499 -161 500 -105
rect 604 -166 605 -160
rect 499 -166 500 -162
rect 887 -166 888 -162
rect 506 -166 507 -164
rect 688 -166 689 -164
rect 51 -253 52 -175
rect 163 -176 164 -174
rect 177 -176 178 -174
rect 506 -253 507 -175
rect 516 -176 517 -174
rect 1157 -253 1158 -175
rect 1220 -176 1221 -174
rect 1227 -253 1228 -175
rect 58 -253 59 -177
rect 261 -178 262 -174
rect 296 -178 297 -174
rect 499 -178 500 -174
rect 530 -253 531 -177
rect 828 -178 829 -174
rect 849 -178 850 -174
rect 884 -253 885 -177
rect 887 -178 888 -174
rect 1087 -253 1088 -177
rect 1097 -253 1098 -177
rect 1150 -253 1151 -177
rect 65 -253 66 -179
rect 450 -180 451 -174
rect 457 -180 458 -174
rect 481 -180 482 -174
rect 544 -180 545 -174
rect 723 -180 724 -174
rect 737 -180 738 -174
rect 1031 -253 1032 -179
rect 1038 -180 1039 -174
rect 1108 -253 1109 -179
rect 1118 -253 1119 -179
rect 1195 -180 1196 -174
rect 72 -253 73 -181
rect 156 -182 157 -174
rect 163 -253 164 -181
rect 432 -182 433 -174
rect 443 -182 444 -174
rect 499 -253 500 -181
rect 541 -182 542 -174
rect 737 -253 738 -181
rect 772 -182 773 -174
rect 1024 -253 1025 -181
rect 1129 -182 1130 -174
rect 1171 -253 1172 -181
rect 79 -253 80 -183
rect 464 -184 465 -174
rect 474 -253 475 -183
rect 1283 -253 1284 -183
rect 86 -253 87 -185
rect 240 -186 241 -174
rect 261 -253 262 -185
rect 352 -186 353 -174
rect 366 -186 367 -174
rect 495 -253 496 -185
rect 548 -186 549 -174
rect 723 -253 724 -185
rect 772 -253 773 -185
rect 821 -253 822 -185
rect 863 -186 864 -174
rect 1038 -253 1039 -185
rect 1125 -253 1126 -185
rect 1129 -253 1130 -185
rect 1136 -186 1137 -174
rect 1255 -253 1256 -185
rect 93 -188 94 -174
rect 100 -253 101 -187
rect 107 -253 108 -187
rect 114 -188 115 -174
rect 121 -253 122 -187
rect 513 -188 514 -174
rect 548 -253 549 -187
rect 614 -188 615 -174
rect 639 -188 640 -174
rect 639 -253 640 -187
rect 639 -188 640 -174
rect 639 -253 640 -187
rect 646 -188 647 -174
rect 646 -253 647 -187
rect 646 -188 647 -174
rect 646 -253 647 -187
rect 653 -188 654 -174
rect 835 -188 836 -174
rect 870 -188 871 -174
rect 1052 -253 1053 -187
rect 93 -253 94 -189
rect 170 -190 171 -174
rect 177 -253 178 -189
rect 191 -190 192 -174
rect 212 -253 213 -189
rect 303 -190 304 -174
rect 317 -190 318 -174
rect 352 -253 353 -189
rect 380 -190 381 -174
rect 509 -190 510 -174
rect 614 -253 615 -189
rect 758 -190 759 -174
rect 789 -253 790 -189
rect 842 -190 843 -174
rect 877 -253 878 -189
rect 891 -190 892 -174
rect 905 -190 906 -174
rect 1017 -253 1018 -189
rect 117 -253 118 -191
rect 170 -253 171 -191
rect 184 -192 185 -174
rect 201 -253 202 -191
rect 219 -192 220 -174
rect 359 -192 360 -174
rect 380 -253 381 -191
rect 527 -192 528 -174
rect 569 -192 570 -174
rect 842 -253 843 -191
rect 880 -192 881 -174
rect 898 -192 899 -174
rect 905 -253 906 -191
rect 968 -192 969 -174
rect 975 -192 976 -174
rect 1080 -253 1081 -191
rect 128 -253 129 -193
rect 268 -194 269 -174
rect 292 -253 293 -193
rect 366 -253 367 -193
rect 383 -253 384 -193
rect 513 -253 514 -193
rect 656 -194 657 -174
rect 975 -253 976 -193
rect 996 -194 997 -174
rect 1101 -253 1102 -193
rect 142 -196 143 -174
rect 215 -196 216 -174
rect 219 -253 220 -195
rect 282 -196 283 -174
rect 296 -253 297 -195
rect 583 -196 584 -174
rect 688 -196 689 -174
rect 835 -253 836 -195
rect 898 -253 899 -195
rect 940 -196 941 -174
rect 954 -196 955 -174
rect 1073 -253 1074 -195
rect 142 -253 143 -197
rect 149 -198 150 -174
rect 156 -253 157 -197
rect 593 -253 594 -197
rect 688 -253 689 -197
rect 856 -198 857 -174
rect 933 -198 934 -174
rect 1143 -253 1144 -197
rect 149 -253 150 -199
rect 408 -200 409 -174
rect 415 -200 416 -174
rect 446 -253 447 -199
rect 457 -253 458 -199
rect 632 -200 633 -174
rect 681 -200 682 -174
rect 856 -253 857 -199
rect 940 -253 941 -199
rect 961 -200 962 -174
rect 968 -253 969 -199
rect 982 -200 983 -174
rect 996 -253 997 -199
rect 1059 -253 1060 -199
rect 184 -253 185 -201
rect 198 -202 199 -174
rect 254 -202 255 -174
rect 282 -253 283 -201
rect 303 -253 304 -201
rect 520 -202 521 -174
rect 632 -253 633 -201
rect 674 -202 675 -174
rect 681 -253 682 -201
rect 919 -202 920 -174
rect 999 -253 1000 -201
rect 1066 -253 1067 -201
rect 191 -253 192 -203
rect 205 -253 206 -203
rect 254 -253 255 -203
rect 324 -204 325 -174
rect 345 -204 346 -174
rect 408 -253 409 -203
rect 429 -253 430 -203
rect 534 -204 535 -174
rect 562 -204 563 -174
rect 674 -253 675 -203
rect 698 -204 699 -174
rect 1003 -253 1004 -203
rect 1010 -204 1011 -174
rect 1136 -253 1137 -203
rect 268 -253 269 -205
rect 387 -206 388 -174
rect 394 -206 395 -174
rect 450 -253 451 -205
rect 492 -206 493 -174
rect 583 -253 584 -205
rect 709 -206 710 -174
rect 863 -253 864 -205
rect 947 -206 948 -174
rect 1010 -253 1011 -205
rect 275 -208 276 -174
rect 415 -253 416 -207
rect 509 -253 510 -207
rect 653 -253 654 -207
rect 716 -208 717 -174
rect 1045 -253 1046 -207
rect 208 -210 209 -174
rect 275 -253 276 -209
rect 289 -210 290 -174
rect 324 -253 325 -209
rect 345 -253 346 -209
rect 362 -210 363 -174
rect 387 -253 388 -209
rect 523 -210 524 -174
rect 534 -253 535 -209
rect 730 -210 731 -174
rect 744 -210 745 -174
rect 870 -253 871 -209
rect 243 -212 244 -174
rect 289 -253 290 -211
rect 310 -212 311 -174
rect 394 -253 395 -211
rect 422 -212 423 -174
rect 730 -253 731 -211
rect 751 -212 752 -174
rect 982 -253 983 -211
rect 135 -214 136 -174
rect 243 -253 244 -213
rect 310 -253 311 -213
rect 331 -214 332 -174
rect 359 -253 360 -213
rect 831 -253 832 -213
rect 135 -253 136 -215
rect 233 -216 234 -174
rect 317 -253 318 -215
rect 338 -216 339 -174
rect 422 -253 423 -215
rect 569 -253 570 -215
rect 604 -216 605 -174
rect 709 -253 710 -215
rect 765 -216 766 -174
rect 891 -253 892 -215
rect 233 -253 234 -217
rect 758 -253 759 -217
rect 765 -253 766 -217
rect 926 -218 927 -174
rect 247 -220 248 -174
rect 338 -253 339 -219
rect 471 -220 472 -174
rect 926 -253 927 -219
rect 247 -253 248 -221
rect 544 -253 545 -221
rect 562 -253 563 -221
rect 590 -222 591 -174
rect 604 -253 605 -221
rect 625 -222 626 -174
rect 660 -222 661 -174
rect 751 -253 752 -221
rect 768 -222 769 -174
rect 919 -253 920 -221
rect 331 -253 332 -223
rect 579 -253 580 -223
rect 702 -224 703 -174
rect 744 -253 745 -223
rect 779 -224 780 -174
rect 933 -253 934 -223
rect 436 -226 437 -174
rect 471 -253 472 -225
rect 478 -253 479 -225
rect 590 -253 591 -225
rect 611 -226 612 -174
rect 779 -253 780 -225
rect 793 -226 794 -174
rect 961 -253 962 -225
rect 236 -228 237 -174
rect 436 -253 437 -227
rect 520 -253 521 -227
rect 576 -228 577 -174
rect 611 -253 612 -227
rect 947 -253 948 -227
rect 226 -230 227 -174
rect 236 -253 237 -229
rect 541 -253 542 -229
rect 625 -253 626 -229
rect 793 -253 794 -229
rect 912 -230 913 -174
rect 226 -253 227 -231
rect 373 -232 374 -174
rect 555 -232 556 -174
rect 660 -253 661 -231
rect 719 -253 720 -231
rect 912 -253 913 -231
rect 373 -253 374 -233
rect 443 -253 444 -233
rect 555 -253 556 -233
rect 695 -234 696 -174
rect 796 -234 797 -174
rect 1164 -253 1165 -233
rect 572 -253 573 -235
rect 695 -253 696 -235
rect 800 -236 801 -174
rect 849 -253 850 -235
rect 502 -238 503 -174
rect 800 -253 801 -237
rect 807 -238 808 -174
rect 989 -253 990 -237
rect 618 -240 619 -174
rect 702 -253 703 -239
rect 786 -240 787 -174
rect 807 -253 808 -239
rect 814 -240 815 -174
rect 954 -253 955 -239
rect 460 -253 461 -241
rect 618 -253 619 -241
rect 597 -244 598 -174
rect 814 -253 815 -243
rect 597 -253 598 -245
rect 667 -246 668 -174
rect 485 -248 486 -174
rect 667 -253 668 -247
rect 401 -250 402 -174
rect 485 -253 486 -249
rect 401 -253 402 -251
rect 467 -253 468 -251
rect 44 -384 45 -262
rect 296 -263 297 -261
rect 383 -263 384 -261
rect 541 -384 542 -262
rect 548 -263 549 -261
rect 590 -384 591 -262
rect 593 -263 594 -261
rect 947 -263 948 -261
rect 989 -263 990 -261
rect 1381 -384 1382 -262
rect 51 -265 52 -261
rect 236 -265 237 -261
rect 285 -384 286 -264
rect 1150 -265 1151 -261
rect 1164 -265 1165 -261
rect 1346 -384 1347 -264
rect 51 -384 52 -266
rect 429 -267 430 -261
rect 460 -267 461 -261
rect 667 -267 668 -261
rect 681 -267 682 -261
rect 947 -384 948 -266
rect 996 -384 997 -266
rect 1157 -267 1158 -261
rect 1202 -384 1203 -266
rect 1353 -384 1354 -266
rect 58 -269 59 -261
rect 341 -384 342 -268
rect 415 -269 416 -261
rect 464 -384 465 -268
rect 471 -269 472 -261
rect 751 -269 752 -261
rect 772 -384 773 -268
rect 821 -269 822 -261
rect 828 -269 829 -261
rect 1213 -384 1214 -268
rect 1227 -269 1228 -261
rect 1227 -384 1228 -268
rect 1227 -269 1228 -261
rect 1227 -384 1228 -268
rect 1255 -269 1256 -261
rect 1374 -384 1375 -268
rect 61 -384 62 -270
rect 72 -271 73 -261
rect 86 -271 87 -261
rect 471 -384 472 -270
rect 474 -271 475 -261
rect 835 -271 836 -261
rect 842 -271 843 -261
rect 1290 -384 1291 -270
rect 72 -384 73 -272
rect 93 -273 94 -261
rect 96 -384 97 -272
rect 121 -273 122 -261
rect 142 -273 143 -261
rect 415 -384 416 -272
rect 474 -384 475 -272
rect 1325 -384 1326 -272
rect 65 -275 66 -261
rect 142 -384 143 -274
rect 156 -275 157 -261
rect 233 -275 234 -261
rect 338 -275 339 -261
rect 429 -384 430 -274
rect 506 -275 507 -261
rect 1234 -384 1235 -274
rect 1283 -275 1284 -261
rect 1591 -384 1592 -274
rect 65 -384 66 -276
rect 453 -384 454 -276
rect 509 -277 510 -261
rect 856 -277 857 -261
rect 863 -277 864 -261
rect 1339 -384 1340 -276
rect 86 -384 87 -278
rect 138 -384 139 -278
rect 163 -279 164 -261
rect 467 -279 468 -261
rect 513 -279 514 -261
rect 1388 -384 1389 -278
rect 107 -281 108 -261
rect 296 -384 297 -280
rect 387 -281 388 -261
rect 513 -384 514 -280
rect 527 -281 528 -261
rect 1360 -384 1361 -280
rect 107 -384 108 -282
rect 457 -283 458 -261
rect 527 -384 528 -282
rect 583 -283 584 -261
rect 614 -283 615 -261
rect 982 -283 983 -261
rect 1024 -283 1025 -261
rect 1206 -384 1207 -282
rect 93 -384 94 -284
rect 457 -384 458 -284
rect 499 -285 500 -261
rect 583 -384 584 -284
rect 632 -285 633 -261
rect 835 -384 836 -284
rect 863 -384 864 -284
rect 1094 -285 1095 -261
rect 1101 -285 1102 -261
rect 1367 -384 1368 -284
rect 121 -384 122 -286
rect 156 -384 157 -286
rect 163 -384 164 -286
rect 205 -287 206 -261
rect 215 -287 216 -261
rect 1262 -384 1263 -286
rect 170 -384 171 -288
rect 282 -289 283 -261
rect 352 -289 353 -261
rect 387 -384 388 -288
rect 450 -289 451 -261
rect 506 -384 507 -288
rect 509 -384 510 -288
rect 632 -384 633 -288
rect 667 -384 668 -288
rect 1276 -384 1277 -288
rect 184 -291 185 -261
rect 184 -384 185 -290
rect 184 -291 185 -261
rect 184 -384 185 -290
rect 198 -291 199 -261
rect 548 -384 549 -290
rect 576 -291 577 -261
rect 828 -384 829 -290
rect 891 -291 892 -261
rect 894 -295 895 -290
rect 905 -291 906 -261
rect 989 -384 990 -290
rect 1038 -291 1039 -261
rect 1283 -384 1284 -290
rect 135 -293 136 -261
rect 576 -384 577 -292
rect 579 -293 580 -261
rect 639 -293 640 -261
rect 681 -384 682 -292
rect 716 -293 717 -261
rect 723 -293 724 -261
rect 842 -384 843 -292
rect 891 -384 892 -292
rect 898 -293 899 -261
rect 912 -293 913 -261
rect 1241 -384 1242 -292
rect 201 -384 202 -294
rect 380 -384 381 -294
rect 408 -295 409 -261
rect 450 -384 451 -294
rect 478 -295 479 -261
rect 639 -384 640 -294
rect 688 -295 689 -261
rect 821 -384 822 -294
rect 898 -384 899 -294
rect 933 -295 934 -261
rect 1094 -384 1095 -294
rect 1101 -384 1102 -294
rect 1143 -295 1144 -261
rect 1171 -295 1172 -261
rect 1255 -384 1256 -294
rect 114 -384 115 -296
rect 933 -384 934 -296
rect 1045 -297 1046 -261
rect 1297 -384 1298 -296
rect 205 -384 206 -298
rect 530 -299 531 -261
rect 544 -299 545 -261
rect 716 -384 717 -298
rect 744 -299 745 -261
rect 982 -384 983 -298
rect 1052 -299 1053 -261
rect 1304 -384 1305 -298
rect 282 -384 283 -300
rect 345 -301 346 -261
rect 359 -301 360 -261
rect 478 -384 479 -300
rect 499 -384 500 -300
rect 1395 -384 1396 -300
rect 275 -303 276 -261
rect 345 -384 346 -302
rect 359 -384 360 -302
rect 373 -303 374 -261
rect 443 -303 444 -261
rect 1171 -384 1172 -302
rect 198 -384 199 -304
rect 443 -384 444 -304
rect 611 -305 612 -261
rect 1038 -384 1039 -304
rect 1059 -305 1060 -261
rect 1150 -384 1151 -304
rect 317 -307 318 -261
rect 352 -384 353 -306
rect 373 -384 374 -306
rect 422 -307 423 -261
rect 611 -384 612 -306
rect 1031 -307 1032 -261
rect 1073 -307 1074 -261
rect 1332 -384 1333 -306
rect 58 -384 59 -308
rect 1031 -384 1032 -308
rect 1073 -384 1074 -308
rect 1097 -309 1098 -261
rect 1108 -309 1109 -261
rect 1318 -384 1319 -308
rect 324 -311 325 -261
rect 408 -384 409 -310
rect 422 -384 423 -310
rect 555 -311 556 -261
rect 614 -384 615 -310
rect 723 -384 724 -310
rect 747 -384 748 -310
rect 1003 -311 1004 -261
rect 1017 -311 1018 -261
rect 1108 -384 1109 -310
rect 1115 -311 1116 -261
rect 1129 -311 1130 -261
rect 1136 -311 1137 -261
rect 1311 -384 1312 -310
rect 173 -313 174 -261
rect 1115 -384 1116 -312
rect 1118 -313 1119 -261
rect 1248 -384 1249 -312
rect 324 -384 325 -314
rect 733 -384 734 -314
rect 751 -384 752 -314
rect 1185 -384 1186 -314
rect 492 -317 493 -261
rect 1129 -384 1130 -316
rect 226 -319 227 -261
rect 492 -384 493 -318
rect 555 -384 556 -318
rect 793 -319 794 -261
rect 800 -319 801 -261
rect 905 -384 906 -318
rect 968 -319 969 -261
rect 1059 -384 1060 -318
rect 1066 -319 1067 -261
rect 1136 -384 1137 -318
rect 149 -321 150 -261
rect 226 -384 227 -320
rect 495 -321 496 -261
rect 800 -384 801 -320
rect 807 -321 808 -261
rect 807 -384 808 -320
rect 807 -321 808 -261
rect 807 -384 808 -320
rect 814 -321 815 -261
rect 1024 -384 1025 -320
rect 1080 -321 1081 -261
rect 1164 -384 1165 -320
rect 149 -384 150 -322
rect 243 -323 244 -261
rect 618 -323 619 -261
rect 688 -384 689 -322
rect 695 -323 696 -261
rect 912 -384 913 -322
rect 919 -323 920 -261
rect 968 -384 969 -322
rect 975 -323 976 -261
rect 1045 -384 1046 -322
rect 1087 -323 1088 -261
rect 1220 -384 1221 -322
rect 607 -384 608 -324
rect 618 -384 619 -324
rect 625 -325 626 -261
rect 695 -384 696 -324
rect 705 -384 706 -324
rect 1178 -384 1179 -324
rect 520 -327 521 -261
rect 625 -384 626 -326
rect 670 -384 671 -326
rect 1052 -384 1053 -326
rect 1122 -327 1123 -261
rect 1192 -384 1193 -326
rect 520 -384 521 -328
rect 534 -329 535 -261
rect 674 -329 675 -261
rect 793 -384 794 -328
rect 870 -329 871 -261
rect 1003 -384 1004 -328
rect 366 -331 367 -261
rect 534 -384 535 -330
rect 562 -331 563 -261
rect 870 -384 871 -330
rect 926 -331 927 -261
rect 1087 -384 1088 -330
rect 191 -333 192 -261
rect 562 -384 563 -332
rect 653 -333 654 -261
rect 674 -384 675 -332
rect 709 -333 710 -261
rect 814 -384 815 -332
rect 884 -333 885 -261
rect 926 -384 927 -332
rect 961 -333 962 -261
rect 1122 -384 1123 -332
rect 79 -335 80 -261
rect 709 -384 710 -334
rect 712 -384 713 -334
rect 1269 -384 1270 -334
rect 79 -384 80 -336
rect 331 -337 332 -261
rect 439 -384 440 -336
rect 653 -384 654 -336
rect 730 -337 731 -261
rect 919 -384 920 -336
rect 975 -384 976 -336
rect 1010 -337 1011 -261
rect 177 -339 178 -261
rect 191 -384 192 -338
rect 254 -339 255 -261
rect 366 -384 367 -338
rect 730 -384 731 -338
rect 1017 -384 1018 -338
rect 177 -384 178 -340
rect 247 -341 248 -261
rect 331 -384 332 -340
rect 572 -341 573 -261
rect 754 -384 755 -340
rect 884 -384 885 -340
rect 999 -341 1000 -261
rect 1080 -384 1081 -340
rect 208 -384 209 -342
rect 254 -384 255 -342
rect 758 -343 759 -261
rect 1066 -384 1067 -342
rect 646 -345 647 -261
rect 758 -384 759 -344
rect 779 -345 780 -261
rect 856 -384 857 -344
rect 877 -345 878 -261
rect 961 -384 962 -344
rect 194 -347 195 -261
rect 646 -384 647 -346
rect 660 -347 661 -261
rect 779 -384 780 -346
rect 786 -347 787 -261
rect 1143 -384 1144 -346
rect 117 -349 118 -261
rect 786 -384 787 -348
rect 789 -349 790 -261
rect 954 -349 955 -261
rect 117 -384 118 -350
rect 240 -384 241 -350
rect 569 -351 570 -261
rect 877 -384 878 -350
rect 940 -351 941 -261
rect 954 -384 955 -350
rect 569 -384 570 -352
rect 1157 -384 1158 -352
rect 604 -355 605 -261
rect 660 -384 661 -354
rect 737 -355 738 -261
rect 940 -384 941 -354
rect 485 -357 486 -261
rect 737 -384 738 -356
rect 849 -357 850 -261
rect 1010 -384 1011 -356
rect 401 -359 402 -261
rect 485 -384 486 -358
rect 597 -359 598 -261
rect 604 -384 605 -358
rect 765 -359 766 -261
rect 849 -384 850 -358
rect 289 -361 290 -261
rect 597 -384 598 -360
rect 702 -361 703 -261
rect 765 -384 766 -360
rect 275 -384 276 -362
rect 702 -384 703 -362
rect 289 -384 290 -364
rect 303 -365 304 -261
rect 338 -384 339 -364
rect 401 -384 402 -364
rect 303 -384 304 -366
rect 394 -367 395 -261
rect 268 -369 269 -261
rect 394 -384 395 -368
rect 268 -384 269 -370
rect 310 -371 311 -261
rect 261 -373 262 -261
rect 310 -384 311 -372
rect 219 -375 220 -261
rect 261 -384 262 -374
rect 219 -384 220 -376
rect 436 -377 437 -261
rect 128 -379 129 -261
rect 436 -384 437 -378
rect 100 -381 101 -261
rect 128 -384 129 -380
rect 100 -384 101 -382
rect 411 -384 412 -382
rect 23 -495 24 -393
rect 233 -495 234 -393
rect 247 -495 248 -393
rect 453 -495 454 -393
rect 506 -394 507 -392
rect 1290 -394 1291 -392
rect 1297 -394 1298 -392
rect 1444 -495 1445 -393
rect 1591 -394 1592 -392
rect 1710 -495 1711 -393
rect 30 -495 31 -395
rect 443 -396 444 -392
rect 450 -396 451 -392
rect 1486 -495 1487 -395
rect 37 -495 38 -397
rect 100 -398 101 -392
rect 107 -398 108 -392
rect 362 -495 363 -397
rect 408 -398 409 -392
rect 583 -398 584 -392
rect 597 -398 598 -392
rect 730 -398 731 -392
rect 772 -398 773 -392
rect 772 -495 773 -397
rect 772 -398 773 -392
rect 772 -495 773 -397
rect 1143 -398 1144 -392
rect 1451 -495 1452 -397
rect 58 -495 59 -399
rect 275 -400 276 -392
rect 317 -495 318 -399
rect 387 -400 388 -392
rect 429 -400 430 -392
rect 523 -495 524 -399
rect 530 -495 531 -399
rect 744 -400 745 -392
rect 1031 -400 1032 -392
rect 1143 -495 1144 -399
rect 1164 -400 1165 -392
rect 1465 -495 1466 -399
rect 72 -402 73 -392
rect 72 -495 73 -401
rect 72 -402 73 -392
rect 72 -495 73 -401
rect 82 -495 83 -401
rect 576 -402 577 -392
rect 607 -402 608 -392
rect 1339 -402 1340 -392
rect 1346 -402 1347 -392
rect 1500 -495 1501 -401
rect 86 -404 87 -392
rect 408 -495 409 -403
rect 429 -495 430 -403
rect 758 -404 759 -392
rect 933 -404 934 -392
rect 1031 -495 1032 -403
rect 1052 -404 1053 -392
rect 1164 -495 1165 -403
rect 1171 -404 1172 -392
rect 1339 -495 1340 -403
rect 1353 -404 1354 -392
rect 1479 -495 1480 -403
rect 86 -495 87 -405
rect 583 -495 584 -405
rect 611 -406 612 -392
rect 793 -406 794 -392
rect 807 -406 808 -392
rect 1052 -495 1053 -405
rect 1066 -406 1067 -392
rect 1171 -495 1172 -405
rect 1178 -406 1179 -392
rect 1297 -495 1298 -405
rect 1304 -406 1305 -392
rect 1409 -495 1410 -405
rect 89 -495 90 -407
rect 128 -408 129 -392
rect 135 -408 136 -392
rect 933 -495 934 -407
rect 982 -408 983 -392
rect 1066 -495 1067 -407
rect 1073 -408 1074 -392
rect 1178 -495 1179 -407
rect 1220 -408 1221 -392
rect 1493 -495 1494 -407
rect 93 -495 94 -409
rect 103 -495 104 -409
rect 110 -495 111 -409
rect 919 -410 920 -392
rect 982 -495 983 -409
rect 1080 -410 1081 -392
rect 1094 -410 1095 -392
rect 1220 -495 1221 -409
rect 1227 -410 1228 -392
rect 1290 -495 1291 -409
rect 1311 -410 1312 -392
rect 1416 -495 1417 -409
rect 96 -412 97 -392
rect 681 -412 682 -392
rect 695 -412 696 -392
rect 793 -495 794 -411
rect 905 -412 906 -392
rect 1094 -495 1095 -411
rect 1115 -412 1116 -392
rect 1227 -495 1228 -411
rect 1269 -412 1270 -392
rect 1423 -495 1424 -411
rect 100 -495 101 -413
rect 1248 -414 1249 -392
rect 1269 -495 1270 -413
rect 1398 -414 1399 -392
rect 114 -495 115 -415
rect 261 -416 262 -392
rect 268 -416 269 -392
rect 285 -416 286 -392
rect 324 -416 325 -392
rect 474 -416 475 -392
rect 481 -495 482 -415
rect 1073 -495 1074 -415
rect 1136 -416 1137 -392
rect 1346 -495 1347 -415
rect 1353 -495 1354 -415
rect 1524 -495 1525 -415
rect 65 -418 66 -392
rect 268 -495 269 -417
rect 324 -495 325 -417
rect 569 -418 570 -392
rect 576 -495 577 -417
rect 688 -418 689 -392
rect 695 -495 696 -417
rect 737 -418 738 -392
rect 747 -418 748 -392
rect 1311 -495 1312 -417
rect 1318 -418 1319 -392
rect 1430 -495 1431 -417
rect 65 -495 66 -419
rect 359 -420 360 -392
rect 366 -420 367 -392
rect 387 -495 388 -419
rect 436 -420 437 -392
rect 527 -420 528 -392
rect 534 -420 535 -392
rect 593 -495 594 -419
rect 618 -420 619 -392
rect 730 -495 731 -419
rect 733 -420 734 -392
rect 1304 -495 1305 -419
rect 1325 -420 1326 -392
rect 1472 -495 1473 -419
rect 79 -422 80 -392
rect 366 -495 367 -421
rect 401 -422 402 -392
rect 436 -495 437 -421
rect 439 -422 440 -392
rect 744 -495 745 -421
rect 758 -495 759 -421
rect 842 -422 843 -392
rect 884 -422 885 -392
rect 1325 -495 1326 -421
rect 1332 -422 1333 -392
rect 1458 -495 1459 -421
rect 79 -495 80 -423
rect 359 -495 360 -423
rect 474 -495 475 -423
rect 1136 -495 1137 -423
rect 1192 -424 1193 -392
rect 1332 -495 1333 -423
rect 1374 -424 1375 -392
rect 1507 -495 1508 -423
rect 121 -426 122 -392
rect 299 -495 300 -425
rect 331 -426 332 -392
rect 401 -495 402 -425
rect 485 -426 486 -392
rect 506 -495 507 -425
rect 534 -495 535 -425
rect 1318 -495 1319 -425
rect 121 -495 122 -427
rect 499 -428 500 -392
rect 541 -428 542 -392
rect 569 -495 570 -427
rect 639 -428 640 -392
rect 751 -428 752 -392
rect 842 -495 843 -427
rect 1122 -428 1123 -392
rect 1206 -428 1207 -392
rect 1374 -495 1375 -427
rect 124 -430 125 -392
rect 1129 -430 1130 -392
rect 1276 -430 1277 -392
rect 1402 -495 1403 -429
rect 128 -495 129 -431
rect 135 -495 136 -431
rect 156 -432 157 -392
rect 156 -495 157 -431
rect 156 -432 157 -392
rect 156 -495 157 -431
rect 163 -432 164 -392
rect 166 -440 167 -431
rect 170 -432 171 -392
rect 418 -495 419 -431
rect 464 -432 465 -392
rect 485 -495 486 -431
rect 492 -432 493 -392
rect 541 -495 542 -431
rect 653 -432 654 -392
rect 751 -495 752 -431
rect 856 -432 857 -392
rect 884 -495 885 -431
rect 919 -495 920 -431
rect 926 -432 927 -392
rect 954 -432 955 -392
rect 1248 -495 1249 -431
rect 1283 -432 1284 -392
rect 1437 -495 1438 -431
rect 51 -434 52 -392
rect 653 -495 654 -433
rect 660 -434 661 -392
rect 667 -495 668 -433
rect 670 -434 671 -392
rect 1388 -434 1389 -392
rect 51 -495 52 -435
rect 303 -436 304 -392
rect 331 -495 332 -435
rect 471 -495 472 -435
rect 478 -436 479 -392
rect 499 -495 500 -435
rect 509 -436 510 -392
rect 856 -495 857 -435
rect 898 -436 899 -392
rect 954 -495 955 -435
rect 968 -436 969 -392
rect 1129 -495 1130 -435
rect 1255 -436 1256 -392
rect 1388 -495 1389 -435
rect 163 -495 164 -437
rect 289 -438 290 -392
rect 303 -495 304 -437
rect 394 -438 395 -392
rect 443 -495 444 -437
rect 492 -495 493 -437
rect 604 -438 605 -392
rect 926 -495 927 -437
rect 989 -438 990 -392
rect 1115 -495 1116 -437
rect 1150 -438 1151 -392
rect 1255 -495 1256 -437
rect 1283 -495 1284 -437
rect 1367 -438 1368 -392
rect 289 -495 290 -439
rect 352 -440 353 -392
rect 527 -495 528 -439
rect 562 -440 563 -392
rect 604 -495 605 -439
rect 625 -440 626 -392
rect 660 -495 661 -439
rect 674 -440 675 -392
rect 681 -495 682 -439
rect 702 -440 703 -392
rect 1381 -440 1382 -392
rect 26 -495 27 -441
rect 562 -495 563 -441
rect 632 -442 633 -392
rect 674 -495 675 -441
rect 712 -442 713 -392
rect 1276 -495 1277 -441
rect 142 -444 143 -392
rect 625 -495 626 -443
rect 632 -495 633 -443
rect 1514 -495 1515 -443
rect 142 -495 143 -445
rect 296 -446 297 -392
rect 352 -495 353 -445
rect 555 -446 556 -392
rect 716 -446 717 -392
rect 807 -495 808 -445
rect 863 -446 864 -392
rect 968 -495 969 -445
rect 1010 -446 1011 -392
rect 1122 -495 1123 -445
rect 1213 -446 1214 -392
rect 1367 -495 1368 -445
rect 117 -448 118 -392
rect 716 -495 717 -447
rect 800 -448 801 -392
rect 863 -495 864 -447
rect 877 -448 878 -392
rect 989 -495 990 -447
rect 1017 -448 1018 -392
rect 1206 -495 1207 -447
rect 1241 -448 1242 -392
rect 1381 -495 1382 -447
rect 170 -495 171 -449
rect 422 -450 423 -392
rect 464 -495 465 -449
rect 590 -450 591 -392
rect 649 -495 650 -449
rect 877 -495 878 -449
rect 891 -450 892 -392
rect 1010 -495 1011 -449
rect 1017 -495 1018 -449
rect 1101 -450 1102 -392
rect 1108 -450 1109 -392
rect 1213 -495 1214 -449
rect 180 -495 181 -451
rect 702 -495 703 -451
rect 709 -495 710 -451
rect 1241 -495 1242 -451
rect 187 -495 188 -453
rect 422 -495 423 -453
rect 478 -495 479 -453
rect 1360 -454 1361 -392
rect 194 -495 195 -455
rect 611 -495 612 -455
rect 779 -456 780 -392
rect 891 -495 892 -455
rect 898 -495 899 -455
rect 1528 -495 1529 -455
rect 198 -458 199 -392
rect 905 -495 906 -457
rect 996 -458 997 -392
rect 1108 -495 1109 -457
rect 1199 -458 1200 -392
rect 1360 -495 1361 -457
rect 184 -460 185 -392
rect 198 -495 199 -459
rect 205 -460 206 -392
rect 261 -495 262 -459
rect 282 -460 283 -392
rect 737 -495 738 -459
rect 870 -460 871 -392
rect 996 -495 997 -459
rect 1003 -460 1004 -392
rect 1101 -495 1102 -459
rect 1185 -460 1186 -392
rect 1199 -495 1200 -459
rect 205 -495 206 -461
rect 513 -462 514 -392
rect 520 -462 521 -392
rect 555 -495 556 -461
rect 590 -495 591 -461
rect 821 -462 822 -392
rect 870 -495 871 -461
rect 947 -462 948 -392
rect 1003 -495 1004 -461
rect 1395 -462 1396 -392
rect 44 -464 45 -392
rect 821 -495 822 -463
rect 849 -464 850 -392
rect 947 -495 948 -463
rect 1038 -464 1039 -392
rect 1150 -495 1151 -463
rect 1262 -464 1263 -392
rect 1395 -495 1396 -463
rect 44 -495 45 -465
rect 226 -466 227 -392
rect 254 -466 255 -392
rect 275 -495 276 -465
rect 282 -495 283 -465
rect 495 -495 496 -465
rect 520 -495 521 -465
rect 1024 -466 1025 -392
rect 1045 -466 1046 -392
rect 1080 -495 1081 -465
rect 1087 -466 1088 -392
rect 1185 -495 1186 -465
rect 191 -468 192 -392
rect 226 -495 227 -467
rect 254 -495 255 -467
rect 614 -468 615 -392
rect 635 -495 636 -467
rect 1262 -495 1263 -467
rect 191 -495 192 -469
rect 513 -495 514 -469
rect 723 -470 724 -392
rect 779 -495 780 -469
rect 786 -470 787 -392
rect 849 -495 850 -469
rect 940 -470 941 -392
rect 1045 -495 1046 -469
rect 1087 -495 1088 -469
rect 1157 -470 1158 -392
rect 138 -472 139 -392
rect 786 -495 787 -471
rect 961 -472 962 -392
rect 1038 -495 1039 -471
rect 1059 -472 1060 -392
rect 1157 -495 1158 -471
rect 138 -495 139 -473
rect 618 -495 619 -473
rect 723 -495 724 -473
rect 814 -474 815 -392
rect 828 -474 829 -392
rect 1059 -495 1060 -473
rect 215 -476 216 -392
rect 688 -495 689 -475
rect 828 -495 829 -475
rect 1234 -476 1235 -392
rect 107 -495 108 -477
rect 1234 -495 1235 -477
rect 219 -480 220 -392
rect 639 -495 640 -479
rect 835 -480 836 -392
rect 961 -495 962 -479
rect 975 -480 976 -392
rect 1024 -495 1025 -479
rect 338 -482 339 -392
rect 814 -495 815 -481
rect 912 -482 913 -392
rect 975 -495 976 -481
rect 338 -495 339 -483
rect 345 -484 346 -392
rect 380 -484 381 -392
rect 394 -495 395 -483
rect 548 -484 549 -392
rect 912 -495 913 -483
rect 149 -486 150 -392
rect 380 -495 381 -485
rect 457 -486 458 -392
rect 548 -495 549 -485
rect 597 -495 598 -485
rect 940 -495 941 -485
rect 149 -495 150 -487
rect 177 -488 178 -392
rect 310 -488 311 -392
rect 345 -495 346 -487
rect 457 -495 458 -487
rect 646 -488 647 -392
rect 765 -488 766 -392
rect 835 -495 836 -487
rect 177 -495 178 -489
rect 212 -490 213 -392
rect 310 -495 311 -489
rect 415 -490 416 -392
rect 646 -495 647 -489
rect 800 -495 801 -489
rect 212 -495 213 -491
rect 240 -492 241 -392
rect 373 -492 374 -392
rect 765 -495 766 -491
rect 219 -495 220 -493
rect 240 -495 241 -493
rect 320 -494 321 -392
rect 373 -495 374 -493
rect 9 -602 10 -504
rect 282 -505 283 -503
rect 317 -505 318 -503
rect 415 -602 416 -504
rect 450 -505 451 -503
rect 863 -505 864 -503
rect 873 -602 874 -504
rect 982 -505 983 -503
rect 1045 -505 1046 -503
rect 1045 -602 1046 -504
rect 1045 -505 1046 -503
rect 1045 -602 1046 -504
rect 1136 -505 1137 -503
rect 1192 -602 1193 -504
rect 1269 -505 1270 -503
rect 1272 -505 1273 -503
rect 1468 -602 1469 -504
rect 1556 -602 1557 -504
rect 1710 -505 1711 -503
rect 1759 -602 1760 -504
rect 23 -602 24 -506
rect 51 -507 52 -503
rect 58 -507 59 -503
rect 100 -507 101 -503
rect 103 -507 104 -503
rect 324 -507 325 -503
rect 345 -507 346 -503
rect 345 -602 346 -506
rect 345 -507 346 -503
rect 345 -602 346 -506
rect 359 -507 360 -503
rect 408 -507 409 -503
rect 450 -602 451 -506
rect 569 -507 570 -503
rect 583 -507 584 -503
rect 607 -577 608 -506
rect 618 -507 619 -503
rect 982 -602 983 -506
rect 1129 -507 1130 -503
rect 1136 -602 1137 -506
rect 1171 -507 1172 -503
rect 1171 -602 1172 -506
rect 1171 -507 1172 -503
rect 1171 -602 1172 -506
rect 1269 -602 1270 -506
rect 1304 -507 1305 -503
rect 1486 -507 1487 -503
rect 1521 -602 1522 -506
rect 1528 -507 1529 -503
rect 1766 -602 1767 -506
rect 37 -509 38 -503
rect 184 -602 185 -508
rect 194 -509 195 -503
rect 1164 -509 1165 -503
rect 1493 -509 1494 -503
rect 1493 -602 1494 -508
rect 1493 -509 1494 -503
rect 1493 -602 1494 -508
rect 1500 -509 1501 -503
rect 1503 -509 1504 -503
rect 1514 -509 1515 -503
rect 1738 -602 1739 -508
rect 61 -602 62 -510
rect 1262 -511 1263 -503
rect 1458 -511 1459 -503
rect 1514 -602 1515 -510
rect 79 -513 80 -503
rect 324 -602 325 -512
rect 362 -513 363 -503
rect 751 -513 752 -503
rect 758 -513 759 -503
rect 1360 -513 1361 -503
rect 1451 -513 1452 -503
rect 1458 -602 1459 -512
rect 1500 -602 1501 -512
rect 1507 -513 1508 -503
rect 72 -515 73 -503
rect 79 -602 80 -514
rect 103 -602 104 -514
rect 408 -602 409 -514
rect 453 -515 454 -503
rect 597 -515 598 -503
rect 604 -515 605 -503
rect 604 -602 605 -514
rect 604 -515 605 -503
rect 604 -602 605 -514
rect 618 -602 619 -514
rect 1073 -515 1074 -503
rect 1122 -515 1123 -503
rect 1129 -602 1130 -514
rect 1150 -515 1151 -503
rect 1164 -602 1165 -514
rect 1325 -515 1326 -503
rect 1360 -602 1361 -514
rect 1430 -515 1431 -503
rect 1451 -602 1452 -514
rect 72 -602 73 -516
rect 114 -517 115 -503
rect 128 -517 129 -503
rect 219 -602 220 -516
rect 222 -517 223 -503
rect 688 -517 689 -503
rect 709 -517 710 -503
rect 1220 -517 1221 -503
rect 1402 -517 1403 -503
rect 1430 -602 1431 -516
rect 107 -602 108 -518
rect 121 -519 122 -503
rect 128 -602 129 -518
rect 394 -519 395 -503
rect 401 -519 402 -503
rect 474 -519 475 -503
rect 481 -519 482 -503
rect 800 -519 801 -503
rect 824 -602 825 -518
rect 1248 -519 1249 -503
rect 114 -602 115 -520
rect 537 -521 538 -503
rect 541 -521 542 -503
rect 541 -602 542 -520
rect 541 -521 542 -503
rect 541 -602 542 -520
rect 548 -521 549 -503
rect 569 -602 570 -520
rect 583 -602 584 -520
rect 961 -521 962 -503
rect 1052 -521 1053 -503
rect 1122 -602 1123 -520
rect 1185 -521 1186 -503
rect 1220 -602 1221 -520
rect 121 -602 122 -522
rect 338 -523 339 -503
rect 341 -602 342 -522
rect 548 -602 549 -522
rect 590 -602 591 -522
rect 828 -523 829 -503
rect 831 -523 832 -503
rect 1150 -602 1151 -522
rect 1199 -523 1200 -503
rect 1325 -602 1326 -522
rect 138 -525 139 -503
rect 1444 -525 1445 -503
rect 152 -602 153 -526
rect 586 -602 587 -526
rect 593 -527 594 -503
rect 1073 -602 1074 -526
rect 1080 -527 1081 -503
rect 1402 -602 1403 -526
rect 1416 -527 1417 -503
rect 1444 -602 1445 -526
rect 156 -529 157 -503
rect 187 -529 188 -503
rect 243 -602 244 -528
rect 359 -602 360 -528
rect 373 -529 374 -503
rect 534 -529 535 -503
rect 593 -602 594 -528
rect 1199 -602 1200 -528
rect 1213 -529 1214 -503
rect 1248 -602 1249 -528
rect 1395 -529 1396 -503
rect 1416 -602 1417 -528
rect 44 -531 45 -503
rect 534 -602 535 -530
rect 597 -602 598 -530
rect 814 -531 815 -503
rect 828 -602 829 -530
rect 835 -531 836 -503
rect 842 -531 843 -503
rect 1262 -602 1263 -530
rect 1367 -531 1368 -503
rect 1395 -602 1396 -530
rect 44 -602 45 -532
rect 901 -533 902 -503
rect 905 -533 906 -503
rect 905 -602 906 -532
rect 905 -533 906 -503
rect 905 -602 906 -532
rect 947 -533 948 -503
rect 950 -577 951 -532
rect 961 -602 962 -532
rect 1066 -533 1067 -503
rect 1178 -533 1179 -503
rect 1213 -602 1214 -532
rect 1332 -533 1333 -503
rect 1367 -602 1368 -532
rect 93 -535 94 -503
rect 156 -602 157 -534
rect 177 -602 178 -534
rect 198 -535 199 -503
rect 268 -535 269 -503
rect 296 -602 297 -534
rect 317 -602 318 -534
rect 765 -535 766 -503
rect 779 -535 780 -503
rect 800 -602 801 -534
rect 842 -602 843 -534
rect 1437 -535 1438 -503
rect 93 -602 94 -536
rect 142 -537 143 -503
rect 180 -537 181 -503
rect 205 -537 206 -503
rect 268 -602 269 -536
rect 520 -537 521 -503
rect 530 -537 531 -503
rect 730 -537 731 -503
rect 761 -537 762 -503
rect 1185 -602 1186 -536
rect 1318 -537 1319 -503
rect 1332 -602 1333 -536
rect 1409 -537 1410 -503
rect 1437 -602 1438 -536
rect 65 -539 66 -503
rect 520 -602 521 -538
rect 530 -602 531 -538
rect 646 -602 647 -538
rect 667 -539 668 -503
rect 712 -539 713 -503
rect 716 -539 717 -503
rect 758 -602 759 -538
rect 765 -602 766 -538
rect 1339 -539 1340 -503
rect 1388 -539 1389 -503
rect 1409 -602 1410 -538
rect 65 -602 66 -540
rect 135 -541 136 -503
rect 142 -602 143 -540
rect 457 -541 458 -503
rect 460 -602 461 -540
rect 1423 -541 1424 -503
rect 135 -602 136 -542
rect 149 -543 150 -503
rect 191 -602 192 -542
rect 457 -602 458 -542
rect 464 -543 465 -503
rect 649 -543 650 -503
rect 653 -543 654 -503
rect 667 -602 668 -542
rect 677 -602 678 -542
rect 716 -602 717 -542
rect 723 -543 724 -503
rect 814 -602 815 -542
rect 915 -602 916 -542
rect 1388 -602 1389 -542
rect 149 -602 150 -544
rect 310 -545 311 -503
rect 352 -545 353 -503
rect 653 -602 654 -544
rect 681 -545 682 -503
rect 723 -602 724 -544
rect 730 -602 731 -544
rect 793 -545 794 -503
rect 947 -602 948 -544
rect 1017 -545 1018 -503
rect 1080 -602 1081 -544
rect 1157 -545 1158 -503
rect 1178 -602 1179 -544
rect 1297 -545 1298 -503
rect 1318 -602 1319 -544
rect 1339 -602 1340 -544
rect 1381 -545 1382 -503
rect 198 -602 199 -546
rect 254 -547 255 -503
rect 275 -547 276 -503
rect 282 -602 283 -546
rect 310 -602 311 -546
rect 506 -547 507 -503
rect 516 -547 517 -503
rect 709 -602 710 -546
rect 779 -602 780 -546
rect 1472 -547 1473 -503
rect 30 -549 31 -503
rect 506 -602 507 -548
rect 516 -602 517 -548
rect 1157 -602 1158 -548
rect 1297 -602 1298 -548
rect 1346 -549 1347 -503
rect 1472 -602 1473 -548
rect 1479 -549 1480 -503
rect 163 -551 164 -503
rect 275 -602 276 -550
rect 366 -551 367 -503
rect 373 -602 374 -550
rect 380 -551 381 -503
rect 401 -602 402 -550
rect 464 -602 465 -550
rect 695 -551 696 -503
rect 786 -551 787 -503
rect 835 -602 836 -550
rect 954 -551 955 -503
rect 1017 -602 1018 -550
rect 1038 -551 1039 -503
rect 1066 -602 1067 -550
rect 1283 -551 1284 -503
rect 1479 -602 1480 -550
rect 163 -602 164 -552
rect 261 -553 262 -503
rect 366 -602 367 -552
rect 485 -553 486 -503
rect 492 -553 493 -503
rect 891 -553 892 -503
rect 919 -553 920 -503
rect 1038 -602 1039 -552
rect 1052 -602 1053 -552
rect 1311 -553 1312 -503
rect 1346 -602 1347 -552
rect 1465 -553 1466 -503
rect 205 -602 206 -554
rect 247 -555 248 -503
rect 254 -602 255 -554
rect 576 -555 577 -503
rect 625 -555 626 -503
rect 852 -602 853 -554
rect 891 -602 892 -554
rect 1535 -602 1536 -554
rect 30 -602 31 -556
rect 247 -602 248 -556
rect 261 -602 262 -556
rect 478 -557 479 -503
rect 485 -602 486 -556
rect 611 -557 612 -503
rect 625 -602 626 -556
rect 737 -557 738 -503
rect 786 -602 787 -556
rect 1003 -557 1004 -503
rect 1241 -557 1242 -503
rect 1283 -602 1284 -556
rect 1290 -557 1291 -503
rect 1311 -602 1312 -556
rect 170 -559 171 -503
rect 611 -602 612 -558
rect 632 -602 633 -558
rect 996 -559 997 -503
rect 1087 -559 1088 -503
rect 1290 -602 1291 -558
rect 170 -602 171 -560
rect 429 -561 430 -503
rect 436 -561 437 -503
rect 478 -602 479 -560
rect 492 -602 493 -560
rect 856 -561 857 -503
rect 919 -602 920 -560
rect 1059 -561 1060 -503
rect 1087 -602 1088 -560
rect 1227 -561 1228 -503
rect 226 -563 227 -503
rect 352 -602 353 -562
rect 387 -563 388 -503
rect 394 -602 395 -562
rect 418 -563 419 -503
rect 1241 -602 1242 -562
rect 226 -602 227 -564
rect 443 -565 444 -503
rect 471 -602 472 -564
rect 562 -565 563 -503
rect 576 -602 577 -564
rect 1108 -565 1109 -503
rect 1195 -565 1196 -503
rect 1227 -602 1228 -564
rect 233 -567 234 -503
rect 443 -602 444 -566
rect 495 -567 496 -503
rect 968 -567 969 -503
rect 1055 -602 1056 -566
rect 1108 -602 1109 -566
rect 303 -569 304 -503
rect 387 -602 388 -568
rect 499 -569 500 -503
rect 499 -602 500 -568
rect 499 -569 500 -503
rect 499 -602 500 -568
rect 523 -569 524 -503
rect 1381 -602 1382 -568
rect 240 -571 241 -503
rect 303 -602 304 -570
rect 331 -571 332 -503
rect 436 -602 437 -570
rect 527 -571 528 -503
rect 1423 -602 1424 -570
rect 212 -573 213 -503
rect 331 -602 332 -572
rect 527 -602 528 -572
rect 1276 -573 1277 -503
rect 212 -602 213 -574
rect 422 -575 423 -503
rect 562 -602 563 -574
rect 772 -575 773 -503
rect 793 -602 794 -574
rect 884 -575 885 -503
rect 1059 -602 1060 -574
rect 1255 -575 1256 -503
rect 1276 -602 1277 -574
rect 240 -602 241 -576
rect 289 -577 290 -503
rect 338 -602 339 -576
rect 422 -602 423 -576
rect 635 -577 636 -503
rect 1094 -577 1095 -503
rect 1234 -577 1235 -503
rect 1255 -602 1256 -576
rect 1503 -602 1504 -576
rect 1507 -602 1508 -576
rect 289 -602 290 -578
rect 299 -579 300 -503
rect 579 -602 580 -578
rect 635 -602 636 -578
rect 639 -579 640 -503
rect 751 -602 752 -578
rect 772 -602 773 -578
rect 849 -579 850 -503
rect 856 -602 857 -578
rect 933 -579 934 -503
rect 968 -602 969 -578
rect 975 -579 976 -503
rect 1094 -602 1095 -578
rect 1115 -579 1116 -503
rect 1206 -579 1207 -503
rect 1234 -602 1235 -578
rect 639 -602 640 -580
rect 674 -581 675 -503
rect 688 -602 689 -580
rect 807 -581 808 -503
rect 849 -602 850 -580
rect 996 -602 997 -580
rect 1101 -581 1102 -503
rect 1115 -602 1116 -580
rect 1143 -581 1144 -503
rect 1206 -602 1207 -580
rect 555 -583 556 -503
rect 674 -602 675 -582
rect 698 -583 699 -503
rect 1003 -602 1004 -582
rect 1031 -583 1032 -503
rect 1101 -602 1102 -582
rect 51 -602 52 -584
rect 698 -602 699 -584
rect 702 -585 703 -503
rect 807 -602 808 -584
rect 866 -602 867 -584
rect 1143 -602 1144 -584
rect 513 -602 514 -586
rect 555 -602 556 -586
rect 660 -587 661 -503
rect 681 -602 682 -586
rect 702 -602 703 -586
rect 845 -602 846 -586
rect 877 -587 878 -503
rect 975 -602 976 -586
rect 1024 -587 1025 -503
rect 1031 -602 1032 -586
rect 86 -589 87 -503
rect 660 -602 661 -588
rect 737 -602 738 -588
rect 744 -589 745 -503
rect 870 -589 871 -503
rect 877 -602 878 -588
rect 884 -602 885 -588
rect 894 -602 895 -588
rect 926 -589 927 -503
rect 954 -602 955 -588
rect 1010 -589 1011 -503
rect 1024 -602 1025 -588
rect 86 -602 87 -590
rect 600 -591 601 -503
rect 744 -602 745 -590
rect 821 -591 822 -503
rect 912 -591 913 -503
rect 926 -602 927 -590
rect 940 -591 941 -503
rect 1010 -602 1011 -590
rect 453 -602 454 -592
rect 940 -602 941 -592
rect 821 -602 822 -594
rect 1486 -602 1487 -594
rect 912 -602 913 -596
rect 1374 -597 1375 -503
rect 1353 -599 1354 -503
rect 1374 -602 1375 -598
rect 110 -601 111 -503
rect 1353 -602 1354 -600
rect 9 -612 10 -610
rect 453 -612 454 -610
rect 492 -612 493 -610
rect 590 -612 591 -610
rect 604 -612 605 -610
rect 632 -711 633 -611
rect 653 -612 654 -610
rect 656 -612 657 -610
rect 674 -711 675 -611
rect 709 -612 710 -610
rect 761 -711 762 -611
rect 947 -612 948 -610
rect 1017 -612 1018 -610
rect 1052 -711 1053 -611
rect 1332 -612 1333 -610
rect 1332 -711 1333 -611
rect 1332 -612 1333 -610
rect 1332 -711 1333 -611
rect 1339 -612 1340 -610
rect 1528 -711 1529 -611
rect 1535 -612 1536 -610
rect 1787 -711 1788 -611
rect 9 -711 10 -613
rect 268 -614 269 -610
rect 282 -614 283 -610
rect 282 -711 283 -613
rect 282 -614 283 -610
rect 282 -711 283 -613
rect 303 -614 304 -610
rect 317 -711 318 -613
rect 320 -614 321 -610
rect 380 -711 381 -613
rect 408 -614 409 -610
rect 712 -711 713 -613
rect 786 -614 787 -610
rect 821 -614 822 -610
rect 824 -614 825 -610
rect 961 -614 962 -610
rect 1241 -614 1242 -610
rect 1339 -711 1340 -613
rect 1346 -614 1347 -610
rect 1619 -711 1620 -613
rect 1668 -711 1669 -613
rect 1801 -711 1802 -613
rect 16 -711 17 -615
rect 93 -616 94 -610
rect 114 -616 115 -610
rect 184 -616 185 -610
rect 205 -616 206 -610
rect 205 -711 206 -615
rect 205 -616 206 -610
rect 205 -711 206 -615
rect 233 -616 234 -610
rect 261 -616 262 -610
rect 303 -711 304 -615
rect 324 -616 325 -610
rect 362 -711 363 -615
rect 649 -711 650 -615
rect 653 -711 654 -615
rect 667 -616 668 -610
rect 677 -616 678 -610
rect 1430 -616 1431 -610
rect 1437 -616 1438 -610
rect 1591 -711 1592 -615
rect 1738 -616 1739 -610
rect 1822 -711 1823 -615
rect 30 -618 31 -610
rect 58 -618 59 -610
rect 72 -618 73 -610
rect 457 -618 458 -610
rect 534 -618 535 -610
rect 534 -711 535 -617
rect 534 -618 535 -610
rect 534 -711 535 -617
rect 544 -711 545 -617
rect 611 -618 612 -610
rect 660 -618 661 -610
rect 961 -711 962 -617
rect 1087 -618 1088 -610
rect 1346 -711 1347 -617
rect 1388 -618 1389 -610
rect 1535 -711 1536 -617
rect 1556 -618 1557 -610
rect 1657 -711 1658 -617
rect 1759 -618 1760 -610
rect 1794 -711 1795 -617
rect 30 -711 31 -619
rect 117 -711 118 -619
rect 145 -711 146 -619
rect 268 -711 269 -619
rect 352 -620 353 -610
rect 457 -711 458 -619
rect 569 -620 570 -610
rect 590 -711 591 -619
rect 604 -711 605 -619
rect 716 -620 717 -610
rect 786 -711 787 -619
rect 999 -711 1000 -619
rect 1157 -620 1158 -610
rect 1241 -711 1242 -619
rect 1325 -620 1326 -610
rect 1437 -711 1438 -619
rect 1444 -620 1445 -610
rect 1577 -711 1578 -619
rect 1766 -620 1767 -610
rect 1857 -711 1858 -619
rect 37 -711 38 -621
rect 870 -622 871 -610
rect 873 -622 874 -610
rect 1388 -711 1389 -621
rect 1409 -622 1410 -610
rect 1542 -711 1543 -621
rect 44 -624 45 -610
rect 96 -711 97 -623
rect 114 -711 115 -623
rect 1262 -624 1263 -610
rect 1290 -624 1291 -610
rect 1409 -711 1410 -623
rect 1416 -624 1417 -610
rect 1563 -711 1564 -623
rect 44 -711 45 -625
rect 499 -626 500 -610
rect 667 -711 668 -625
rect 702 -626 703 -610
rect 709 -711 710 -625
rect 1570 -711 1571 -625
rect 51 -628 52 -610
rect 72 -711 73 -627
rect 79 -628 80 -610
rect 82 -660 83 -627
rect 128 -628 129 -610
rect 352 -711 353 -627
rect 373 -628 374 -610
rect 429 -628 430 -610
rect 436 -628 437 -610
rect 436 -711 437 -627
rect 436 -628 437 -610
rect 436 -711 437 -627
rect 499 -711 500 -627
rect 506 -628 507 -610
rect 681 -628 682 -610
rect 702 -711 703 -627
rect 793 -628 794 -610
rect 912 -711 913 -627
rect 933 -628 934 -610
rect 1192 -628 1193 -610
rect 1206 -628 1207 -610
rect 1262 -711 1263 -627
rect 1269 -628 1270 -610
rect 1416 -711 1417 -627
rect 1423 -628 1424 -610
rect 1556 -711 1557 -627
rect 51 -711 52 -629
rect 103 -630 104 -610
rect 128 -711 129 -629
rect 135 -630 136 -610
rect 149 -630 150 -610
rect 324 -711 325 -629
rect 373 -711 374 -629
rect 383 -630 384 -610
rect 408 -711 409 -629
rect 422 -630 423 -610
rect 429 -711 430 -629
rect 471 -630 472 -610
rect 509 -711 510 -629
rect 1206 -711 1207 -629
rect 1227 -630 1228 -610
rect 1325 -711 1326 -629
rect 1451 -630 1452 -610
rect 1584 -711 1585 -629
rect 58 -711 59 -631
rect 65 -632 66 -610
rect 79 -711 80 -631
rect 135 -711 136 -631
rect 1633 -711 1634 -631
rect 65 -711 66 -633
rect 142 -634 143 -610
rect 149 -711 150 -633
rect 212 -634 213 -610
rect 243 -634 244 -610
rect 443 -634 444 -610
rect 681 -711 682 -633
rect 751 -634 752 -610
rect 796 -711 797 -633
rect 1465 -634 1466 -610
rect 1472 -634 1473 -610
rect 1549 -711 1550 -633
rect 142 -711 143 -635
rect 765 -636 766 -610
rect 800 -636 801 -610
rect 821 -711 822 -635
rect 842 -636 843 -610
rect 1101 -636 1102 -610
rect 1108 -636 1109 -610
rect 1157 -711 1158 -635
rect 1178 -636 1179 -610
rect 1269 -711 1270 -635
rect 1353 -636 1354 -610
rect 1472 -711 1473 -635
rect 1479 -636 1480 -610
rect 1612 -711 1613 -635
rect 100 -638 101 -610
rect 1108 -711 1109 -637
rect 1129 -638 1130 -610
rect 1227 -711 1228 -637
rect 1360 -638 1361 -610
rect 1465 -711 1466 -637
rect 1468 -638 1469 -610
rect 1479 -711 1480 -637
rect 1486 -638 1487 -610
rect 1626 -711 1627 -637
rect 100 -711 101 -639
rect 191 -640 192 -610
rect 212 -711 213 -639
rect 467 -711 468 -639
rect 562 -640 563 -610
rect 800 -711 801 -639
rect 849 -640 850 -610
rect 1514 -640 1515 -610
rect 156 -642 157 -610
rect 891 -711 892 -641
rect 894 -642 895 -610
rect 1402 -642 1403 -610
rect 1458 -642 1459 -610
rect 1598 -711 1599 -641
rect 156 -711 157 -643
rect 401 -644 402 -610
rect 415 -644 416 -610
rect 513 -644 514 -610
rect 562 -711 563 -643
rect 730 -644 731 -610
rect 737 -644 738 -610
rect 765 -711 766 -643
rect 782 -711 783 -643
rect 1458 -711 1459 -643
rect 1493 -644 1494 -610
rect 1640 -711 1641 -643
rect 163 -646 164 -610
rect 492 -711 493 -645
rect 513 -711 514 -645
rect 548 -646 549 -610
rect 569 -711 570 -645
rect 842 -711 843 -645
rect 845 -711 846 -645
rect 1514 -711 1515 -645
rect 163 -711 164 -647
rect 646 -648 647 -610
rect 660 -711 661 -647
rect 737 -711 738 -647
rect 852 -648 853 -610
rect 1213 -648 1214 -610
rect 1255 -648 1256 -610
rect 1360 -711 1361 -647
rect 1374 -648 1375 -610
rect 1486 -711 1487 -647
rect 1500 -648 1501 -610
rect 1661 -711 1662 -647
rect 170 -650 171 -610
rect 527 -650 528 -610
rect 593 -650 594 -610
rect 849 -711 850 -649
rect 863 -650 864 -610
rect 1430 -711 1431 -649
rect 1507 -650 1508 -610
rect 1647 -711 1648 -649
rect 170 -711 171 -651
rect 1290 -711 1291 -651
rect 1297 -652 1298 -610
rect 1507 -711 1508 -651
rect 173 -711 174 -653
rect 618 -654 619 -610
rect 646 -711 647 -653
rect 719 -711 720 -653
rect 723 -654 724 -610
rect 751 -711 752 -653
rect 870 -711 871 -653
rect 922 -711 923 -653
rect 989 -654 990 -610
rect 1087 -711 1088 -653
rect 1115 -654 1116 -610
rect 1213 -711 1214 -653
rect 1248 -654 1249 -610
rect 1255 -711 1256 -653
rect 1311 -654 1312 -610
rect 1374 -711 1375 -653
rect 1381 -654 1382 -610
rect 1493 -711 1494 -653
rect 177 -656 178 -610
rect 177 -711 178 -655
rect 177 -656 178 -610
rect 177 -711 178 -655
rect 187 -656 188 -610
rect 1444 -711 1445 -655
rect 191 -711 192 -657
rect 198 -658 199 -610
rect 236 -658 237 -610
rect 415 -711 416 -657
rect 422 -711 423 -657
rect 530 -658 531 -610
rect 635 -658 636 -610
rect 989 -711 990 -657
rect 996 -658 997 -610
rect 1101 -711 1102 -657
rect 1136 -658 1137 -610
rect 1353 -711 1354 -657
rect 1367 -658 1368 -610
rect 1500 -711 1501 -657
rect 198 -711 199 -659
rect 338 -660 339 -610
rect 366 -660 367 -610
rect 471 -711 472 -659
rect 520 -660 521 -610
rect 548 -711 549 -659
rect 656 -711 657 -659
rect 723 -711 724 -659
rect 730 -711 731 -659
rect 744 -660 745 -610
rect 877 -660 878 -610
rect 947 -711 948 -659
rect 1024 -660 1025 -610
rect 1136 -711 1137 -659
rect 1164 -660 1165 -610
rect 1248 -711 1249 -659
rect 1276 -660 1277 -610
rect 1381 -711 1382 -659
rect 61 -662 62 -610
rect 1024 -711 1025 -661
rect 1031 -662 1032 -610
rect 1178 -711 1179 -661
rect 1185 -662 1186 -610
rect 1276 -711 1277 -661
rect 1283 -662 1284 -610
rect 1367 -711 1368 -661
rect 236 -711 237 -663
rect 583 -711 584 -663
rect 625 -664 626 -610
rect 744 -711 745 -663
rect 828 -664 829 -610
rect 877 -711 878 -663
rect 898 -664 899 -610
rect 933 -711 934 -663
rect 1038 -664 1039 -610
rect 1297 -711 1298 -663
rect 1318 -664 1319 -610
rect 1402 -711 1403 -663
rect 240 -666 241 -610
rect 366 -711 367 -665
rect 387 -666 388 -610
rect 618 -711 619 -665
rect 625 -711 626 -665
rect 1020 -711 1021 -665
rect 1059 -666 1060 -610
rect 1192 -711 1193 -665
rect 1199 -666 1200 -610
rect 1451 -711 1452 -665
rect 240 -711 241 -667
rect 831 -711 832 -667
rect 856 -668 857 -610
rect 1059 -711 1060 -667
rect 1066 -668 1067 -610
rect 1115 -711 1116 -667
rect 1171 -668 1172 -610
rect 1283 -711 1284 -667
rect 152 -670 153 -610
rect 856 -711 857 -669
rect 908 -711 909 -669
rect 1605 -711 1606 -669
rect 254 -672 255 -610
rect 866 -672 867 -610
rect 926 -672 927 -610
rect 1031 -711 1032 -671
rect 1045 -672 1046 -610
rect 1199 -711 1200 -671
rect 1234 -672 1235 -610
rect 1318 -711 1319 -671
rect 261 -711 262 -673
rect 345 -674 346 -610
rect 387 -711 388 -673
rect 600 -711 601 -673
rect 688 -674 689 -610
rect 863 -711 864 -673
rect 884 -674 885 -610
rect 926 -711 927 -673
rect 954 -674 955 -610
rect 1045 -711 1046 -673
rect 1073 -674 1074 -610
rect 1185 -711 1186 -673
rect 331 -676 332 -610
rect 338 -711 339 -675
rect 345 -711 346 -675
rect 481 -711 482 -675
rect 520 -711 521 -675
rect 541 -676 542 -610
rect 586 -676 587 -610
rect 898 -711 899 -675
rect 940 -676 941 -610
rect 1073 -711 1074 -675
rect 1080 -676 1081 -610
rect 1129 -711 1130 -675
rect 1143 -676 1144 -610
rect 1171 -711 1172 -675
rect 275 -678 276 -610
rect 331 -711 332 -677
rect 401 -711 402 -677
rect 639 -678 640 -610
rect 691 -711 692 -677
rect 915 -678 916 -610
rect 975 -678 976 -610
rect 1038 -711 1039 -677
rect 1150 -678 1151 -610
rect 1234 -711 1235 -677
rect 275 -711 276 -679
rect 394 -680 395 -610
rect 432 -680 433 -610
rect 1311 -711 1312 -679
rect 394 -711 395 -681
rect 779 -682 780 -610
rect 793 -711 794 -681
rect 940 -711 941 -681
rect 982 -682 983 -610
rect 1080 -711 1081 -681
rect 247 -684 248 -610
rect 779 -711 780 -683
rect 814 -684 815 -610
rect 982 -711 983 -683
rect 1003 -684 1004 -610
rect 1150 -711 1151 -683
rect 247 -711 248 -685
rect 289 -686 290 -610
rect 443 -711 444 -685
rect 576 -686 577 -610
rect 597 -686 598 -610
rect 639 -711 640 -685
rect 695 -686 696 -610
rect 1122 -686 1123 -610
rect 289 -711 290 -687
rect 296 -688 297 -610
rect 464 -688 465 -610
rect 527 -711 528 -687
rect 541 -711 542 -687
rect 611 -711 612 -687
rect 695 -711 696 -687
rect 971 -711 972 -687
rect 1010 -688 1011 -610
rect 1066 -711 1067 -687
rect 1122 -711 1123 -687
rect 1395 -688 1396 -610
rect 23 -690 24 -610
rect 464 -711 465 -689
rect 555 -690 556 -610
rect 576 -711 577 -689
rect 597 -711 598 -689
rect 1143 -711 1144 -689
rect 1304 -690 1305 -610
rect 1395 -711 1396 -689
rect 23 -711 24 -691
rect 310 -692 311 -610
rect 698 -692 699 -610
rect 1423 -711 1424 -691
rect 121 -694 122 -610
rect 310 -711 311 -693
rect 740 -711 741 -693
rect 1164 -711 1165 -693
rect 1220 -694 1221 -610
rect 1304 -711 1305 -693
rect 121 -711 122 -695
rect 450 -696 451 -610
rect 772 -696 773 -610
rect 975 -711 976 -695
rect 1094 -696 1095 -610
rect 1220 -711 1221 -695
rect 219 -698 220 -610
rect 296 -711 297 -697
rect 450 -711 451 -697
rect 478 -698 479 -610
rect 758 -698 759 -610
rect 772 -711 773 -697
rect 807 -698 808 -610
rect 814 -711 815 -697
rect 828 -711 829 -697
rect 1521 -698 1522 -610
rect 86 -700 87 -610
rect 219 -711 220 -699
rect 254 -711 255 -699
rect 478 -711 479 -699
rect 506 -711 507 -699
rect 1521 -711 1522 -699
rect 86 -711 87 -701
rect 226 -702 227 -610
rect 621 -711 622 -701
rect 807 -711 808 -701
rect 835 -702 836 -610
rect 954 -711 955 -701
rect 968 -702 969 -610
rect 1094 -711 1095 -701
rect 226 -711 227 -703
rect 758 -711 759 -703
rect 884 -711 885 -703
rect 901 -711 902 -703
rect 905 -704 906 -610
rect 1003 -711 1004 -703
rect 359 -706 360 -610
rect 835 -711 836 -705
rect 919 -706 920 -610
rect 1010 -711 1011 -705
rect 359 -711 360 -707
rect 485 -708 486 -610
rect 485 -711 486 -709
rect 1671 -711 1672 -709
rect 9 -721 10 -719
rect 93 -721 94 -719
rect 114 -721 115 -719
rect 1783 -856 1784 -720
rect 1787 -721 1788 -719
rect 1892 -856 1893 -720
rect 9 -856 10 -722
rect 422 -723 423 -719
rect 439 -856 440 -722
rect 555 -723 556 -719
rect 562 -723 563 -719
rect 649 -723 650 -719
rect 709 -723 710 -719
rect 1297 -723 1298 -719
rect 1458 -723 1459 -719
rect 1843 -856 1844 -722
rect 1857 -723 1858 -719
rect 1885 -856 1886 -722
rect 16 -725 17 -719
rect 117 -725 118 -719
rect 121 -725 122 -719
rect 124 -856 125 -724
rect 128 -725 129 -719
rect 138 -725 139 -719
rect 170 -725 171 -719
rect 180 -856 181 -724
rect 254 -725 255 -719
rect 257 -775 258 -724
rect 303 -725 304 -719
rect 306 -775 307 -724
rect 422 -856 423 -724
rect 719 -725 720 -719
rect 723 -725 724 -719
rect 737 -725 738 -719
rect 740 -725 741 -719
rect 1591 -725 1592 -719
rect 1605 -725 1606 -719
rect 1738 -856 1739 -724
rect 1801 -725 1802 -719
rect 1857 -856 1858 -724
rect 37 -727 38 -719
rect 233 -727 234 -719
rect 254 -856 255 -726
rect 527 -727 528 -719
rect 548 -727 549 -719
rect 562 -856 563 -726
rect 586 -856 587 -726
rect 996 -856 997 -726
rect 999 -727 1000 -719
rect 1563 -727 1564 -719
rect 1577 -727 1578 -719
rect 1731 -856 1732 -726
rect 1822 -727 1823 -719
rect 1850 -856 1851 -726
rect 37 -856 38 -728
rect 572 -856 573 -728
rect 597 -856 598 -728
rect 1451 -729 1452 -719
rect 1486 -729 1487 -719
rect 1675 -856 1676 -728
rect 1794 -729 1795 -719
rect 1822 -856 1823 -728
rect 58 -731 59 -719
rect 544 -731 545 -719
rect 555 -856 556 -730
rect 1591 -856 1592 -730
rect 1612 -731 1613 -719
rect 1759 -856 1760 -730
rect 30 -733 31 -719
rect 58 -856 59 -732
rect 79 -733 80 -719
rect 114 -856 115 -732
rect 121 -856 122 -732
rect 233 -856 234 -732
rect 268 -733 269 -719
rect 527 -856 528 -732
rect 618 -733 619 -719
rect 1297 -856 1298 -732
rect 1360 -733 1361 -719
rect 1451 -856 1452 -732
rect 1493 -733 1494 -719
rect 1605 -856 1606 -732
rect 1626 -733 1627 -719
rect 1787 -856 1788 -732
rect 30 -856 31 -734
rect 100 -735 101 -719
rect 135 -735 136 -719
rect 145 -735 146 -719
rect 170 -856 171 -734
rect 177 -735 178 -719
rect 201 -856 202 -734
rect 1563 -856 1564 -734
rect 1570 -735 1571 -719
rect 1577 -856 1578 -734
rect 1584 -735 1585 -719
rect 1766 -856 1767 -734
rect 93 -856 94 -736
rect 184 -737 185 -719
rect 268 -856 269 -736
rect 415 -737 416 -719
rect 443 -737 444 -719
rect 506 -856 507 -736
rect 520 -737 521 -719
rect 541 -856 542 -736
rect 614 -856 615 -736
rect 618 -856 619 -736
rect 621 -737 622 -719
rect 1486 -856 1487 -736
rect 1542 -737 1543 -719
rect 1689 -856 1690 -736
rect 65 -739 66 -719
rect 520 -856 521 -738
rect 628 -856 629 -738
rect 730 -739 731 -719
rect 779 -739 780 -719
rect 1472 -739 1473 -719
rect 1479 -739 1480 -719
rect 1584 -856 1585 -738
rect 1633 -739 1634 -719
rect 1794 -856 1795 -738
rect 65 -856 66 -740
rect 516 -856 517 -740
rect 632 -741 633 -719
rect 730 -856 731 -740
rect 758 -741 759 -719
rect 1472 -856 1473 -740
rect 1549 -741 1550 -719
rect 1745 -856 1746 -740
rect 100 -856 101 -742
rect 289 -743 290 -719
rect 303 -856 304 -742
rect 387 -743 388 -719
rect 443 -856 444 -742
rect 485 -743 486 -719
rect 495 -856 496 -742
rect 828 -743 829 -719
rect 831 -856 832 -742
rect 1668 -856 1669 -742
rect 1671 -743 1672 -719
rect 1717 -856 1718 -742
rect 107 -745 108 -719
rect 184 -856 185 -744
rect 275 -745 276 -719
rect 415 -856 416 -744
rect 450 -745 451 -719
rect 485 -856 486 -744
rect 590 -745 591 -719
rect 632 -856 633 -744
rect 674 -745 675 -719
rect 709 -856 710 -744
rect 712 -745 713 -719
rect 1801 -856 1802 -744
rect 107 -856 108 -746
rect 471 -747 472 -719
rect 478 -747 479 -719
rect 975 -747 976 -719
rect 1034 -856 1035 -746
rect 1829 -856 1830 -746
rect 135 -856 136 -748
rect 499 -749 500 -719
rect 653 -749 654 -719
rect 674 -856 675 -748
rect 681 -749 682 -719
rect 737 -856 738 -748
rect 779 -856 780 -748
rect 1710 -856 1711 -748
rect 173 -751 174 -719
rect 457 -751 458 -719
rect 464 -751 465 -719
rect 1073 -751 1074 -719
rect 1143 -751 1144 -719
rect 1696 -856 1697 -750
rect 96 -753 97 -719
rect 464 -856 465 -752
rect 478 -856 479 -752
rect 667 -753 668 -719
rect 716 -753 717 -719
rect 1199 -753 1200 -719
rect 1234 -753 1235 -719
rect 1360 -856 1361 -752
rect 1367 -753 1368 -719
rect 1458 -856 1459 -752
rect 1465 -753 1466 -719
rect 1542 -856 1543 -752
rect 1549 -856 1550 -752
rect 1598 -753 1599 -719
rect 1633 -856 1634 -752
rect 1661 -753 1662 -719
rect 156 -755 157 -719
rect 457 -856 458 -754
rect 467 -755 468 -719
rect 667 -856 668 -754
rect 723 -856 724 -754
rect 940 -755 941 -719
rect 1045 -755 1046 -719
rect 1143 -856 1144 -754
rect 1178 -755 1179 -719
rect 1199 -856 1200 -754
rect 1234 -856 1235 -754
rect 1304 -755 1305 -719
rect 1339 -755 1340 -719
rect 1479 -856 1480 -754
rect 1556 -755 1557 -719
rect 1703 -856 1704 -754
rect 51 -757 52 -719
rect 156 -856 157 -756
rect 275 -856 276 -756
rect 282 -757 283 -719
rect 289 -856 290 -756
rect 600 -757 601 -719
rect 639 -757 640 -719
rect 681 -856 682 -756
rect 782 -757 783 -719
rect 905 -856 906 -756
rect 919 -757 920 -719
rect 961 -757 962 -719
rect 1073 -856 1074 -756
rect 1220 -757 1221 -719
rect 1241 -757 1242 -719
rect 1367 -856 1368 -756
rect 1381 -757 1382 -719
rect 1493 -856 1494 -756
rect 1556 -856 1557 -756
rect 1780 -856 1781 -756
rect 282 -856 283 -758
rect 324 -759 325 -719
rect 716 -856 717 -758
rect 793 -759 794 -719
rect 1409 -759 1410 -719
rect 1444 -759 1445 -719
rect 1612 -856 1613 -758
rect 1640 -759 1641 -719
rect 1773 -856 1774 -758
rect 296 -761 297 -719
rect 828 -856 829 -760
rect 835 -761 836 -719
rect 1045 -856 1046 -760
rect 1080 -761 1081 -719
rect 1178 -856 1179 -760
rect 1195 -856 1196 -760
rect 1682 -856 1683 -760
rect 324 -856 325 -762
rect 908 -763 909 -719
rect 922 -763 923 -719
rect 1752 -856 1753 -762
rect 345 -765 346 -719
rect 621 -856 622 -764
rect 772 -765 773 -719
rect 793 -856 794 -764
rect 800 -765 801 -719
rect 803 -765 804 -719
rect 807 -765 808 -719
rect 940 -856 941 -764
rect 1052 -765 1053 -719
rect 1080 -856 1081 -764
rect 1094 -765 1095 -719
rect 1220 -856 1221 -764
rect 1262 -765 1263 -719
rect 1339 -856 1340 -764
rect 1388 -765 1389 -719
rect 1598 -856 1599 -764
rect 1647 -765 1648 -719
rect 1808 -856 1809 -764
rect 345 -856 346 -766
rect 366 -767 367 -719
rect 373 -767 374 -719
rect 961 -856 962 -766
rect 1136 -767 1137 -719
rect 1241 -856 1242 -766
rect 1269 -767 1270 -719
rect 1381 -856 1382 -766
rect 1402 -767 1403 -719
rect 1570 -856 1571 -766
rect 310 -769 311 -719
rect 366 -856 367 -768
rect 373 -856 374 -768
rect 401 -769 402 -719
rect 436 -769 437 -719
rect 471 -856 472 -768
rect 492 -769 493 -719
rect 499 -856 500 -768
rect 569 -769 570 -719
rect 639 -856 640 -768
rect 695 -769 696 -719
rect 772 -856 773 -768
rect 800 -856 801 -768
rect 870 -769 871 -719
rect 884 -769 885 -719
rect 1626 -856 1627 -768
rect 54 -856 55 -770
rect 310 -856 311 -770
rect 401 -856 402 -770
rect 408 -771 409 -719
rect 450 -856 451 -770
rect 919 -856 920 -770
rect 933 -771 934 -719
rect 1094 -856 1095 -770
rect 1157 -771 1158 -719
rect 1262 -856 1263 -770
rect 1276 -771 1277 -719
rect 1388 -856 1389 -770
rect 1430 -771 1431 -719
rect 1647 -856 1648 -770
rect 142 -773 143 -719
rect 933 -856 934 -772
rect 954 -773 955 -719
rect 1052 -856 1053 -772
rect 1101 -773 1102 -719
rect 1157 -856 1158 -772
rect 1283 -773 1284 -719
rect 1444 -856 1445 -772
rect 1465 -856 1466 -772
rect 1528 -773 1529 -719
rect 142 -856 143 -774
rect 198 -775 199 -719
rect 359 -775 360 -719
rect 408 -856 409 -774
rect 492 -856 493 -774
rect 534 -775 535 -719
rect 576 -775 577 -719
rect 653 -856 654 -774
rect 803 -856 804 -774
rect 870 -856 871 -774
rect 898 -775 899 -719
rect 1304 -856 1305 -774
rect 1318 -775 1319 -719
rect 1402 -856 1403 -774
rect 1521 -775 1522 -719
rect 1640 -856 1641 -774
rect 44 -777 45 -719
rect 576 -856 577 -776
rect 604 -777 605 -719
rect 807 -856 808 -776
rect 814 -777 815 -719
rect 835 -856 836 -776
rect 842 -777 843 -719
rect 1353 -777 1354 -719
rect 1437 -777 1438 -719
rect 1521 -856 1522 -776
rect 177 -856 178 -778
rect 898 -856 899 -778
rect 901 -779 902 -719
rect 1619 -779 1620 -719
rect 198 -856 199 -780
rect 359 -856 360 -780
rect 534 -856 535 -780
rect 688 -781 689 -719
rect 824 -856 825 -780
rect 1514 -781 1515 -719
rect 548 -856 549 -782
rect 842 -856 843 -782
rect 845 -783 846 -719
rect 1724 -856 1725 -782
rect 583 -785 584 -719
rect 604 -856 605 -784
rect 611 -785 612 -719
rect 695 -856 696 -784
rect 782 -856 783 -784
rect 1514 -856 1515 -784
rect 163 -787 164 -719
rect 611 -856 612 -786
rect 625 -787 626 -719
rect 814 -856 815 -786
rect 849 -787 850 -719
rect 1017 -787 1018 -719
rect 1020 -787 1021 -719
rect 1437 -856 1438 -786
rect 1507 -787 1508 -719
rect 1619 -856 1620 -786
rect 163 -856 164 -788
rect 1423 -789 1424 -719
rect 583 -856 584 -790
rect 590 -856 591 -790
rect 625 -856 626 -790
rect 1661 -856 1662 -790
rect 646 -793 647 -719
rect 884 -856 885 -792
rect 912 -793 913 -719
rect 954 -856 955 -792
rect 1010 -793 1011 -719
rect 1269 -856 1270 -792
rect 1290 -793 1291 -719
rect 1836 -856 1837 -792
rect 212 -795 213 -719
rect 1010 -856 1011 -794
rect 1031 -795 1032 -719
rect 1136 -856 1137 -794
rect 1185 -795 1186 -719
rect 1283 -856 1284 -794
rect 1311 -795 1312 -719
rect 1423 -856 1424 -794
rect 296 -856 297 -796
rect 1031 -856 1032 -796
rect 1038 -797 1039 -719
rect 1101 -856 1102 -796
rect 1108 -797 1109 -719
rect 1290 -856 1291 -796
rect 1325 -797 1326 -719
rect 1409 -856 1410 -796
rect 1416 -797 1417 -719
rect 1507 -856 1508 -796
rect 166 -856 167 -798
rect 1325 -856 1326 -798
rect 1332 -799 1333 -719
rect 1353 -856 1354 -798
rect 1374 -799 1375 -719
rect 1416 -856 1417 -798
rect 429 -801 430 -719
rect 646 -856 647 -800
rect 744 -801 745 -719
rect 849 -856 850 -800
rect 926 -801 927 -719
rect 1017 -856 1018 -800
rect 1087 -801 1088 -719
rect 1185 -856 1186 -800
rect 1192 -801 1193 -719
rect 1311 -856 1312 -800
rect 1346 -801 1347 -719
rect 1430 -856 1431 -800
rect 79 -856 80 -802
rect 1087 -856 1088 -802
rect 1115 -803 1116 -719
rect 1276 -856 1277 -802
rect 352 -805 353 -719
rect 429 -856 430 -804
rect 509 -805 510 -719
rect 1038 -856 1039 -804
rect 1066 -805 1067 -719
rect 1115 -856 1116 -804
rect 1213 -805 1214 -719
rect 1318 -856 1319 -804
rect 338 -807 339 -719
rect 352 -856 353 -806
rect 691 -856 692 -806
rect 926 -856 927 -806
rect 947 -807 948 -719
rect 1066 -856 1067 -806
rect 1227 -807 1228 -719
rect 1332 -856 1333 -806
rect 82 -856 83 -808
rect 338 -856 339 -808
rect 744 -856 745 -808
rect 751 -809 752 -719
rect 761 -809 762 -719
rect 1213 -856 1214 -808
rect 1248 -809 1249 -719
rect 1374 -856 1375 -808
rect 702 -811 703 -719
rect 751 -856 752 -810
rect 761 -856 762 -810
rect 1206 -811 1207 -719
rect 1255 -811 1256 -719
rect 1528 -856 1529 -810
rect 789 -856 790 -812
rect 947 -856 948 -812
rect 971 -813 972 -719
rect 1346 -856 1347 -812
rect 821 -815 822 -719
rect 912 -856 913 -814
rect 982 -815 983 -719
rect 1206 -856 1207 -814
rect 821 -856 822 -816
rect 1500 -817 1501 -719
rect 863 -819 864 -719
rect 982 -856 983 -818
rect 989 -819 990 -719
rect 1108 -856 1109 -818
rect 1129 -819 1130 -719
rect 1248 -856 1249 -818
rect 1395 -819 1396 -719
rect 1500 -856 1501 -818
rect 765 -821 766 -719
rect 863 -856 864 -820
rect 989 -856 990 -820
rect 1654 -821 1655 -719
rect 226 -823 227 -719
rect 765 -856 766 -822
rect 1003 -823 1004 -719
rect 1129 -856 1130 -822
rect 1150 -823 1151 -719
rect 1227 -856 1228 -822
rect 226 -856 227 -824
rect 261 -825 262 -719
rect 1024 -825 1025 -719
rect 1255 -856 1256 -824
rect 240 -827 241 -719
rect 1003 -856 1004 -826
rect 1150 -856 1151 -826
rect 1164 -827 1165 -719
rect 1171 -827 1172 -719
rect 1395 -856 1396 -826
rect 72 -829 73 -719
rect 1164 -856 1165 -828
rect 1192 -856 1193 -828
rect 1654 -856 1655 -828
rect 72 -856 73 -830
rect 149 -831 150 -719
rect 240 -856 241 -830
rect 247 -831 248 -719
rect 261 -856 262 -830
rect 331 -831 332 -719
rect 891 -831 892 -719
rect 1024 -856 1025 -830
rect 1059 -831 1060 -719
rect 1171 -856 1172 -830
rect 44 -856 45 -832
rect 149 -856 150 -832
rect 205 -833 206 -719
rect 247 -856 248 -832
rect 331 -856 332 -832
rect 380 -833 381 -719
rect 877 -833 878 -719
rect 891 -856 892 -832
rect 968 -833 969 -719
rect 1059 -856 1060 -832
rect 191 -835 192 -719
rect 205 -856 206 -834
rect 380 -856 381 -834
rect 513 -835 514 -719
rect 660 -835 661 -719
rect 877 -856 878 -834
rect 128 -856 129 -836
rect 191 -856 192 -836
rect 212 -856 213 -836
rect 513 -856 514 -836
rect 579 -856 580 -836
rect 660 -856 661 -836
rect 856 -837 857 -719
rect 968 -856 969 -836
rect 786 -839 787 -719
rect 856 -856 857 -838
rect 786 -856 787 -840
rect 1535 -841 1536 -719
rect 1122 -843 1123 -719
rect 1535 -856 1536 -842
rect 558 -845 559 -719
rect 1122 -856 1123 -844
rect 86 -847 87 -719
rect 558 -856 559 -846
rect 86 -856 87 -848
rect 219 -849 220 -719
rect 23 -851 24 -719
rect 219 -856 220 -850
rect 23 -856 24 -852
rect 394 -853 395 -719
rect 187 -855 188 -719
rect 394 -856 395 -854
rect 2 -977 3 -865
rect 68 -977 69 -865
rect 86 -866 87 -864
rect 89 -940 90 -865
rect 110 -977 111 -865
rect 1234 -866 1235 -864
rect 1339 -866 1340 -864
rect 1339 -977 1340 -865
rect 1339 -866 1340 -864
rect 1339 -977 1340 -865
rect 1591 -866 1592 -864
rect 1594 -866 1595 -864
rect 1724 -866 1725 -864
rect 1864 -977 1865 -865
rect 1885 -866 1886 -864
rect 1913 -977 1914 -865
rect 16 -868 17 -864
rect 16 -977 17 -867
rect 16 -868 17 -864
rect 16 -977 17 -867
rect 37 -868 38 -864
rect 79 -868 80 -864
rect 86 -977 87 -867
rect 205 -868 206 -864
rect 261 -868 262 -864
rect 264 -940 265 -867
rect 310 -868 311 -864
rect 943 -977 944 -867
rect 968 -868 969 -864
rect 968 -977 969 -867
rect 968 -868 969 -864
rect 968 -977 969 -867
rect 1006 -977 1007 -867
rect 1766 -868 1767 -864
rect 1780 -868 1781 -864
rect 1822 -868 1823 -864
rect 1829 -868 1830 -864
rect 1941 -977 1942 -867
rect 30 -870 31 -864
rect 79 -977 80 -869
rect 114 -870 115 -864
rect 121 -870 122 -864
rect 135 -870 136 -864
rect 513 -870 514 -864
rect 516 -870 517 -864
rect 1668 -870 1669 -864
rect 1703 -870 1704 -864
rect 1766 -977 1767 -869
rect 1787 -870 1788 -864
rect 1829 -977 1830 -869
rect 1836 -870 1837 -864
rect 1948 -977 1949 -869
rect 30 -977 31 -871
rect 226 -872 227 -864
rect 261 -977 262 -871
rect 275 -872 276 -864
rect 310 -977 311 -871
rect 450 -872 451 -864
rect 460 -977 461 -871
rect 1920 -977 1921 -871
rect 37 -977 38 -873
rect 72 -874 73 -864
rect 121 -977 122 -873
rect 128 -874 129 -864
rect 156 -874 157 -864
rect 821 -874 822 -864
rect 828 -874 829 -864
rect 1612 -874 1613 -864
rect 1633 -874 1634 -864
rect 1885 -977 1886 -873
rect 1892 -874 1893 -864
rect 1955 -977 1956 -873
rect 51 -876 52 -864
rect 114 -977 115 -875
rect 163 -876 164 -864
rect 247 -876 248 -864
rect 275 -977 276 -875
rect 338 -876 339 -864
rect 436 -876 437 -864
rect 450 -977 451 -875
rect 747 -977 748 -875
rect 779 -876 780 -864
rect 1066 -876 1067 -864
rect 1083 -977 1084 -875
rect 1731 -876 1732 -864
rect 1759 -876 1760 -864
rect 1871 -977 1872 -875
rect 47 -878 48 -864
rect 1066 -977 1067 -877
rect 1108 -878 1109 -864
rect 1111 -878 1112 -864
rect 1136 -878 1137 -864
rect 1136 -977 1137 -877
rect 1136 -878 1137 -864
rect 1136 -977 1137 -877
rect 1153 -977 1154 -877
rect 1675 -878 1676 -864
rect 1717 -878 1718 -864
rect 1787 -977 1788 -877
rect 1801 -878 1802 -864
rect 1934 -977 1935 -877
rect 51 -977 52 -879
rect 93 -880 94 -864
rect 177 -880 178 -864
rect 1024 -880 1025 -864
rect 1031 -880 1032 -864
rect 1598 -880 1599 -864
rect 1619 -880 1620 -864
rect 1675 -977 1676 -879
rect 1752 -880 1753 -864
rect 1759 -977 1760 -879
rect 1843 -880 1844 -864
rect 1906 -977 1907 -879
rect 65 -882 66 -864
rect 548 -882 549 -864
rect 572 -882 573 -864
rect 1325 -882 1326 -864
rect 1353 -882 1354 -864
rect 1598 -977 1599 -881
rect 1633 -977 1634 -881
rect 1878 -977 1879 -881
rect 65 -977 66 -883
rect 1013 -977 1014 -883
rect 1031 -977 1032 -883
rect 1528 -884 1529 -864
rect 1556 -884 1557 -864
rect 1612 -977 1613 -883
rect 1654 -884 1655 -864
rect 1724 -977 1725 -883
rect 1794 -884 1795 -864
rect 1843 -977 1844 -883
rect 1850 -884 1851 -864
rect 1881 -977 1882 -883
rect 72 -977 73 -885
rect 233 -886 234 -864
rect 247 -977 248 -885
rect 429 -886 430 -864
rect 492 -886 493 -864
rect 653 -886 654 -864
rect 684 -977 685 -885
rect 828 -977 829 -885
rect 915 -977 916 -885
rect 1325 -977 1326 -885
rect 1360 -886 1361 -864
rect 1619 -977 1620 -885
rect 1661 -886 1662 -864
rect 1717 -977 1718 -885
rect 1738 -886 1739 -864
rect 1794 -977 1795 -885
rect 1857 -886 1858 -864
rect 1892 -977 1893 -885
rect 93 -977 94 -887
rect 163 -977 164 -887
rect 177 -977 178 -887
rect 681 -888 682 -864
rect 688 -888 689 -864
rect 1479 -888 1480 -864
rect 1500 -888 1501 -864
rect 1556 -977 1557 -887
rect 1577 -888 1578 -864
rect 1836 -977 1837 -887
rect 128 -977 129 -889
rect 233 -977 234 -889
rect 268 -890 269 -864
rect 436 -977 437 -889
rect 492 -977 493 -889
rect 562 -890 563 -864
rect 576 -890 577 -864
rect 877 -890 878 -864
rect 919 -890 920 -864
rect 1073 -890 1074 -864
rect 1108 -977 1109 -889
rect 1178 -890 1179 -864
rect 1220 -890 1221 -864
rect 1220 -977 1221 -889
rect 1220 -890 1221 -864
rect 1220 -977 1221 -889
rect 1297 -890 1298 -864
rect 1353 -977 1354 -889
rect 1381 -890 1382 -864
rect 1654 -977 1655 -889
rect 1668 -977 1669 -889
rect 1745 -890 1746 -864
rect 1808 -890 1809 -864
rect 1857 -977 1858 -889
rect 156 -977 157 -891
rect 1360 -977 1361 -891
rect 1430 -892 1431 -864
rect 1479 -977 1480 -891
rect 1521 -892 1522 -864
rect 1577 -977 1578 -891
rect 1591 -977 1592 -891
rect 1710 -892 1711 -864
rect 180 -894 181 -864
rect 380 -894 381 -864
rect 387 -894 388 -864
rect 691 -894 692 -864
rect 705 -894 706 -864
rect 961 -894 962 -864
rect 985 -977 986 -893
rect 1780 -977 1781 -893
rect 58 -896 59 -864
rect 380 -977 381 -895
rect 429 -977 430 -895
rect 590 -896 591 -864
rect 604 -896 605 -864
rect 653 -977 654 -895
rect 688 -977 689 -895
rect 989 -896 990 -864
rect 1003 -896 1004 -864
rect 1024 -977 1025 -895
rect 1034 -896 1035 -864
rect 1444 -896 1445 -864
rect 1451 -896 1452 -864
rect 1500 -977 1501 -895
rect 1521 -977 1522 -895
rect 1584 -896 1585 -864
rect 1605 -896 1606 -864
rect 1661 -977 1662 -895
rect 1689 -896 1690 -864
rect 1738 -977 1739 -895
rect 187 -977 188 -897
rect 597 -898 598 -864
rect 604 -977 605 -897
rect 1563 -898 1564 -864
rect 1640 -898 1641 -864
rect 1689 -977 1690 -897
rect 1696 -898 1697 -864
rect 1752 -977 1753 -897
rect 191 -977 192 -899
rect 863 -900 864 -864
rect 877 -977 878 -899
rect 1192 -900 1193 -864
rect 1374 -900 1375 -864
rect 1430 -977 1431 -899
rect 1465 -900 1466 -864
rect 1801 -977 1802 -899
rect 198 -902 199 -864
rect 555 -977 556 -901
rect 583 -902 584 -864
rect 674 -902 675 -864
rect 723 -902 724 -864
rect 1234 -977 1235 -901
rect 1402 -902 1403 -864
rect 1444 -977 1445 -901
rect 1465 -977 1466 -901
rect 1542 -902 1543 -864
rect 1549 -902 1550 -864
rect 1850 -977 1851 -901
rect 170 -904 171 -864
rect 198 -977 199 -903
rect 201 -904 202 -864
rect 282 -904 283 -864
rect 338 -977 339 -903
rect 443 -904 444 -864
rect 478 -904 479 -864
rect 597 -977 598 -903
rect 618 -904 619 -864
rect 716 -904 717 -864
rect 726 -977 727 -903
rect 1696 -977 1697 -903
rect 170 -977 171 -905
rect 324 -906 325 -864
rect 366 -906 367 -864
rect 366 -977 367 -905
rect 366 -906 367 -864
rect 366 -977 367 -905
rect 394 -906 395 -864
rect 443 -977 444 -905
rect 485 -906 486 -864
rect 562 -977 563 -905
rect 586 -906 587 -864
rect 1045 -906 1046 -864
rect 1059 -906 1060 -864
rect 1528 -977 1529 -905
rect 1535 -906 1536 -864
rect 1605 -977 1606 -905
rect 1647 -906 1648 -864
rect 1710 -977 1711 -905
rect 184 -908 185 -864
rect 394 -977 395 -907
rect 408 -908 409 -864
rect 485 -977 486 -907
rect 495 -908 496 -864
rect 779 -977 780 -907
rect 782 -908 783 -864
rect 1703 -977 1704 -907
rect 184 -977 185 -909
rect 331 -910 332 -864
rect 506 -910 507 -864
rect 548 -977 549 -909
rect 590 -977 591 -909
rect 646 -910 647 -864
rect 674 -977 675 -909
rect 1038 -910 1039 -864
rect 1041 -977 1042 -909
rect 1570 -910 1571 -864
rect 205 -977 206 -911
rect 240 -912 241 -864
rect 324 -977 325 -911
rect 422 -912 423 -864
rect 506 -977 507 -911
rect 513 -977 514 -911
rect 849 -912 850 -864
rect 856 -912 857 -864
rect 1381 -977 1382 -911
rect 1409 -912 1410 -864
rect 1451 -977 1452 -911
rect 1472 -912 1473 -864
rect 1745 -977 1746 -911
rect 212 -914 213 -864
rect 478 -977 479 -913
rect 527 -914 528 -864
rect 558 -914 559 -864
rect 618 -977 619 -913
rect 824 -914 825 -864
rect 831 -914 832 -864
rect 1374 -977 1375 -913
rect 1395 -914 1396 -864
rect 1409 -977 1410 -913
rect 1416 -914 1417 -864
rect 1570 -977 1571 -913
rect 142 -916 143 -864
rect 212 -977 213 -915
rect 240 -977 241 -915
rect 345 -916 346 -864
rect 415 -916 416 -864
rect 422 -977 423 -915
rect 499 -916 500 -864
rect 527 -977 528 -915
rect 534 -916 535 -864
rect 583 -977 584 -915
rect 621 -916 622 -864
rect 1822 -977 1823 -915
rect 226 -977 227 -917
rect 534 -977 535 -917
rect 537 -977 538 -917
rect 1206 -918 1207 -864
rect 1255 -918 1256 -864
rect 1416 -977 1417 -917
rect 1423 -918 1424 -864
rect 1549 -977 1550 -917
rect 1563 -977 1564 -917
rect 1899 -977 1900 -917
rect 268 -977 269 -919
rect 600 -920 601 -864
rect 625 -920 626 -864
rect 751 -920 752 -864
rect 758 -920 759 -864
rect 1045 -977 1046 -919
rect 1059 -977 1060 -919
rect 1297 -977 1298 -919
rect 1318 -920 1319 -864
rect 1423 -977 1424 -919
rect 1486 -920 1487 -864
rect 1535 -977 1536 -919
rect 282 -977 283 -921
rect 359 -922 360 -864
rect 415 -977 416 -921
rect 1094 -922 1095 -864
rect 1115 -922 1116 -864
rect 1255 -977 1256 -921
rect 1276 -922 1277 -864
rect 1318 -977 1319 -921
rect 1346 -922 1347 -864
rect 1402 -977 1403 -921
rect 1486 -977 1487 -921
rect 1916 -977 1917 -921
rect 289 -924 290 -864
rect 331 -977 332 -923
rect 359 -977 360 -923
rect 1783 -924 1784 -864
rect 289 -977 290 -925
rect 352 -926 353 -864
rect 499 -977 500 -925
rect 754 -977 755 -925
rect 758 -977 759 -925
rect 772 -926 773 -864
rect 775 -977 776 -925
rect 1584 -977 1585 -925
rect 254 -928 255 -864
rect 352 -977 353 -927
rect 541 -928 542 -864
rect 576 -977 577 -927
rect 625 -977 626 -927
rect 660 -928 661 -864
rect 709 -928 710 -864
rect 849 -977 850 -927
rect 856 -977 857 -927
rect 975 -928 976 -864
rect 1017 -928 1018 -864
rect 1073 -977 1074 -927
rect 1087 -928 1088 -864
rect 1115 -977 1116 -927
rect 1129 -928 1130 -864
rect 1178 -977 1179 -927
rect 1276 -977 1277 -927
rect 1388 -928 1389 -864
rect 1493 -928 1494 -864
rect 1542 -977 1543 -927
rect 58 -977 59 -929
rect 541 -977 542 -929
rect 632 -930 633 -864
rect 632 -977 633 -929
rect 632 -930 633 -864
rect 632 -977 633 -929
rect 639 -930 640 -864
rect 1017 -977 1018 -929
rect 1052 -930 1053 -864
rect 1087 -977 1088 -929
rect 1094 -977 1095 -929
rect 1101 -930 1102 -864
rect 1122 -930 1123 -864
rect 1129 -977 1130 -929
rect 1164 -930 1165 -864
rect 1192 -977 1193 -929
rect 1283 -930 1284 -864
rect 1346 -977 1347 -929
rect 1367 -930 1368 -864
rect 1472 -977 1473 -929
rect 1493 -977 1494 -929
rect 1682 -930 1683 -864
rect 254 -977 255 -931
rect 569 -932 570 -864
rect 639 -977 640 -931
rect 800 -932 801 -864
rect 814 -932 815 -864
rect 1101 -977 1102 -931
rect 1171 -932 1172 -864
rect 1206 -977 1207 -931
rect 1241 -932 1242 -864
rect 1283 -977 1284 -931
rect 1304 -932 1305 -864
rect 1367 -977 1368 -931
rect 1507 -932 1508 -864
rect 1640 -977 1641 -931
rect 1682 -977 1683 -931
rect 1818 -932 1819 -864
rect 142 -977 143 -933
rect 814 -977 815 -933
rect 821 -977 822 -933
rect 842 -934 843 -864
rect 863 -977 864 -933
rect 912 -934 913 -864
rect 922 -934 923 -864
rect 1731 -977 1732 -933
rect 296 -936 297 -864
rect 408 -977 409 -935
rect 520 -936 521 -864
rect 709 -977 710 -935
rect 716 -977 717 -935
rect 730 -936 731 -864
rect 740 -977 741 -935
rect 1808 -977 1809 -935
rect 296 -977 297 -937
rect 471 -938 472 -864
rect 544 -977 545 -937
rect 569 -977 570 -937
rect 646 -977 647 -937
rect 905 -938 906 -864
rect 922 -977 923 -937
rect 1927 -977 1928 -937
rect 166 -940 167 -864
rect 905 -977 906 -939
rect 926 -940 927 -864
rect 926 -977 927 -939
rect 926 -940 927 -864
rect 926 -977 927 -939
rect 933 -940 934 -864
rect 933 -977 934 -939
rect 933 -940 934 -864
rect 933 -977 934 -939
rect 947 -940 948 -864
rect 989 -977 990 -939
rect 1003 -977 1004 -939
rect 1164 -977 1165 -939
rect 1311 -940 1312 -864
rect 1388 -977 1389 -939
rect 1458 -940 1459 -864
rect 1507 -977 1508 -939
rect 1594 -977 1595 -939
rect 1647 -977 1648 -939
rect 317 -942 318 -864
rect 345 -977 346 -941
rect 401 -942 402 -864
rect 471 -977 472 -941
rect 660 -977 661 -941
rect 940 -942 941 -864
rect 947 -977 948 -941
rect 982 -942 983 -864
rect 1062 -977 1063 -941
rect 1514 -942 1515 -864
rect 149 -944 150 -864
rect 317 -977 318 -943
rect 401 -977 402 -943
rect 457 -944 458 -864
rect 464 -944 465 -864
rect 520 -977 521 -943
rect 702 -944 703 -864
rect 1241 -977 1242 -943
rect 1262 -944 1263 -864
rect 1311 -977 1312 -943
rect 100 -946 101 -864
rect 149 -977 150 -945
rect 373 -946 374 -864
rect 702 -977 703 -945
rect 730 -977 731 -945
rect 1010 -946 1011 -864
rect 1143 -946 1144 -864
rect 1171 -977 1172 -945
rect 1213 -946 1214 -864
rect 1458 -977 1459 -945
rect 9 -948 10 -864
rect 100 -977 101 -947
rect 107 -948 108 -864
rect 373 -977 374 -947
rect 390 -977 391 -947
rect 464 -977 465 -947
rect 744 -948 745 -864
rect 786 -948 787 -864
rect 789 -948 790 -864
rect 842 -977 843 -947
rect 891 -948 892 -864
rect 1052 -977 1053 -947
rect 1080 -948 1081 -864
rect 1143 -977 1144 -947
rect 1157 -948 1158 -864
rect 1304 -977 1305 -947
rect 9 -977 10 -949
rect 23 -950 24 -864
rect 44 -977 45 -949
rect 107 -977 108 -949
rect 135 -977 136 -949
rect 457 -977 458 -949
rect 611 -950 612 -864
rect 786 -977 787 -949
rect 800 -977 801 -949
rect 940 -977 941 -949
rect 954 -950 955 -864
rect 975 -977 976 -949
rect 1010 -977 1011 -949
rect 1773 -950 1774 -864
rect 23 -977 24 -951
rect 194 -952 195 -864
rect 611 -977 612 -951
rect 695 -952 696 -864
rect 744 -977 745 -951
rect 1290 -952 1291 -864
rect 667 -954 668 -864
rect 695 -977 696 -953
rect 761 -954 762 -864
rect 1514 -977 1515 -953
rect 667 -977 668 -955
rect 870 -956 871 -864
rect 884 -956 885 -864
rect 954 -977 955 -955
rect 961 -977 962 -955
rect 996 -956 997 -864
rect 1034 -977 1035 -955
rect 1773 -977 1774 -955
rect 765 -958 766 -864
rect 982 -977 983 -957
rect 996 -977 997 -957
rect 1038 -977 1039 -957
rect 1080 -977 1081 -957
rect 1815 -977 1816 -957
rect 737 -960 738 -864
rect 765 -977 766 -959
rect 772 -977 773 -959
rect 1269 -960 1270 -864
rect 807 -962 808 -864
rect 891 -977 892 -961
rect 1157 -977 1158 -961
rect 1395 -977 1396 -961
rect 793 -964 794 -864
rect 807 -977 808 -963
rect 835 -964 836 -864
rect 870 -977 871 -963
rect 884 -977 885 -963
rect 898 -964 899 -864
rect 1185 -964 1186 -864
rect 1213 -977 1214 -963
rect 1227 -964 1228 -864
rect 1269 -977 1270 -963
rect 54 -966 55 -864
rect 835 -977 836 -965
rect 1150 -966 1151 -864
rect 1185 -977 1186 -965
rect 1248 -966 1249 -864
rect 1290 -977 1291 -965
rect 236 -977 237 -967
rect 1248 -977 1249 -967
rect 1262 -977 1263 -967
rect 1626 -968 1627 -864
rect 439 -970 440 -864
rect 898 -977 899 -969
rect 1437 -970 1438 -864
rect 1626 -977 1627 -969
rect 793 -977 794 -971
rect 1160 -977 1161 -971
rect 1332 -972 1333 -864
rect 1437 -977 1438 -971
rect 1199 -974 1200 -864
rect 1332 -977 1333 -973
rect 628 -976 629 -864
rect 1199 -977 1200 -975
rect 47 -1108 48 -986
rect 702 -987 703 -985
rect 733 -1108 734 -986
rect 772 -987 773 -985
rect 775 -987 776 -985
rect 821 -987 822 -985
rect 866 -1108 867 -986
rect 1423 -987 1424 -985
rect 1444 -987 1445 -985
rect 1444 -1108 1445 -986
rect 1444 -987 1445 -985
rect 1444 -1108 1445 -986
rect 1745 -987 1746 -985
rect 1899 -987 1900 -985
rect 1927 -987 1928 -985
rect 1976 -1108 1977 -986
rect 58 -989 59 -985
rect 453 -1108 454 -988
rect 457 -989 458 -985
rect 537 -989 538 -985
rect 541 -1108 542 -988
rect 625 -989 626 -985
rect 656 -1108 657 -988
rect 1416 -989 1417 -985
rect 1710 -989 1711 -985
rect 1745 -1108 1746 -988
rect 1867 -1108 1868 -988
rect 1892 -989 1893 -985
rect 1927 -1108 1928 -988
rect 1934 -989 1935 -985
rect 1941 -989 1942 -985
rect 1962 -1108 1963 -988
rect 58 -1108 59 -990
rect 170 -991 171 -985
rect 240 -991 241 -985
rect 684 -991 685 -985
rect 709 -991 710 -985
rect 821 -1108 822 -990
rect 870 -991 871 -985
rect 915 -991 916 -985
rect 919 -991 920 -985
rect 1430 -991 1431 -985
rect 1710 -1108 1711 -990
rect 1766 -991 1767 -985
rect 1878 -991 1879 -985
rect 1906 -991 1907 -985
rect 1948 -991 1949 -985
rect 1969 -1108 1970 -990
rect 68 -993 69 -985
rect 394 -993 395 -985
rect 443 -993 444 -985
rect 457 -1108 458 -992
rect 485 -993 486 -985
rect 604 -993 605 -985
rect 625 -1108 626 -992
rect 1437 -993 1438 -985
rect 1584 -993 1585 -985
rect 1878 -1108 1879 -992
rect 1948 -1108 1949 -992
rect 1955 -993 1956 -985
rect 30 -995 31 -985
rect 394 -1108 395 -994
rect 485 -1108 486 -994
rect 618 -995 619 -985
rect 674 -995 675 -985
rect 709 -1108 710 -994
rect 716 -995 717 -985
rect 772 -1108 773 -994
rect 779 -995 780 -985
rect 1416 -1108 1417 -994
rect 1493 -995 1494 -985
rect 1584 -1108 1585 -994
rect 30 -1108 31 -996
rect 51 -997 52 -985
rect 72 -997 73 -985
rect 390 -997 391 -985
rect 513 -997 514 -985
rect 604 -1108 605 -996
rect 667 -997 668 -985
rect 716 -1108 717 -996
rect 737 -997 738 -985
rect 758 -997 759 -985
rect 761 -1108 762 -996
rect 1724 -997 1725 -985
rect 51 -1108 52 -998
rect 408 -999 409 -985
rect 478 -999 479 -985
rect 667 -1108 668 -998
rect 674 -1108 675 -998
rect 1192 -999 1193 -985
rect 1241 -999 1242 -985
rect 1244 -1005 1245 -998
rect 1276 -999 1277 -985
rect 1423 -1108 1424 -998
rect 1493 -1108 1494 -998
rect 1500 -999 1501 -985
rect 1724 -1108 1725 -998
rect 1885 -999 1886 -985
rect 72 -1108 73 -1000
rect 635 -1108 636 -1000
rect 681 -1001 682 -985
rect 1178 -1001 1179 -985
rect 1241 -1108 1242 -1000
rect 1269 -1001 1270 -985
rect 1276 -1108 1277 -1000
rect 1290 -1001 1291 -985
rect 1346 -1001 1347 -985
rect 1346 -1108 1347 -1000
rect 1346 -1001 1347 -985
rect 1346 -1108 1347 -1000
rect 1374 -1001 1375 -985
rect 1374 -1108 1375 -1000
rect 1374 -1001 1375 -985
rect 1374 -1108 1375 -1000
rect 1409 -1001 1410 -985
rect 1430 -1108 1431 -1000
rect 1500 -1108 1501 -1000
rect 1507 -1001 1508 -985
rect 82 -1108 83 -1002
rect 1017 -1003 1018 -985
rect 1020 -1108 1021 -1002
rect 1255 -1003 1256 -985
rect 1367 -1003 1368 -985
rect 1409 -1108 1410 -1002
rect 1507 -1108 1508 -1002
rect 1514 -1003 1515 -985
rect 86 -1005 87 -985
rect 145 -1005 146 -985
rect 149 -1005 150 -985
rect 170 -1108 171 -1004
rect 240 -1108 241 -1004
rect 401 -1005 402 -985
rect 408 -1108 409 -1004
rect 492 -1005 493 -985
rect 513 -1108 514 -1004
rect 611 -1005 612 -985
rect 646 -1005 647 -985
rect 1178 -1108 1179 -1004
rect 1269 -1108 1270 -1004
rect 1514 -1108 1515 -1004
rect 1570 -1005 1571 -985
rect 9 -1007 10 -985
rect 86 -1108 87 -1006
rect 93 -1108 94 -1006
rect 219 -1007 220 -985
rect 261 -1007 262 -985
rect 261 -1108 262 -1006
rect 261 -1007 262 -985
rect 261 -1108 262 -1006
rect 282 -1007 283 -985
rect 726 -1007 727 -985
rect 737 -1108 738 -1006
rect 1437 -1108 1438 -1006
rect 1535 -1007 1536 -985
rect 1570 -1108 1571 -1006
rect 9 -1108 10 -1008
rect 226 -1009 227 -985
rect 282 -1108 283 -1008
rect 436 -1009 437 -985
rect 478 -1108 479 -1008
rect 779 -1108 780 -1008
rect 786 -1009 787 -985
rect 957 -1108 958 -1008
rect 968 -1009 969 -985
rect 1290 -1108 1291 -1008
rect 1535 -1108 1536 -1008
rect 1598 -1009 1599 -985
rect 79 -1011 80 -985
rect 149 -1108 150 -1010
rect 156 -1011 157 -985
rect 443 -1108 444 -1010
rect 492 -1108 493 -1010
rect 730 -1011 731 -985
rect 747 -1011 748 -985
rect 1458 -1011 1459 -985
rect 1598 -1108 1599 -1010
rect 1633 -1011 1634 -985
rect 79 -1108 80 -1012
rect 1234 -1013 1235 -985
rect 1255 -1108 1256 -1012
rect 1297 -1013 1298 -985
rect 1451 -1013 1452 -985
rect 1458 -1108 1459 -1012
rect 68 -1108 69 -1014
rect 1451 -1108 1452 -1014
rect 96 -1017 97 -985
rect 758 -1108 759 -1016
rect 863 -1017 864 -985
rect 870 -1108 871 -1016
rect 891 -1017 892 -985
rect 1367 -1108 1368 -1016
rect 107 -1108 108 -1018
rect 128 -1019 129 -985
rect 142 -1019 143 -985
rect 159 -1019 160 -985
rect 226 -1108 227 -1018
rect 660 -1019 661 -985
rect 681 -1108 682 -1018
rect 1528 -1019 1529 -985
rect 128 -1108 129 -1020
rect 310 -1021 311 -985
rect 345 -1021 346 -985
rect 436 -1108 437 -1020
rect 506 -1021 507 -985
rect 968 -1108 969 -1020
rect 982 -1021 983 -985
rect 1864 -1021 1865 -985
rect 142 -1108 143 -1022
rect 191 -1023 192 -985
rect 268 -1023 269 -985
rect 786 -1108 787 -1022
rect 842 -1023 843 -985
rect 891 -1108 892 -1022
rect 894 -1108 895 -1022
rect 898 -1023 899 -985
rect 912 -1023 913 -985
rect 1472 -1023 1473 -985
rect 37 -1025 38 -985
rect 268 -1108 269 -1024
rect 296 -1025 297 -985
rect 534 -1025 535 -985
rect 548 -1025 549 -985
rect 548 -1108 549 -1024
rect 548 -1025 549 -985
rect 548 -1108 549 -1024
rect 565 -1108 566 -1024
rect 611 -1108 612 -1024
rect 632 -1025 633 -985
rect 660 -1108 661 -1024
rect 702 -1108 703 -1024
rect 730 -1108 731 -1024
rect 751 -1025 752 -985
rect 1773 -1025 1774 -985
rect 37 -1108 38 -1026
rect 471 -1027 472 -985
rect 499 -1027 500 -985
rect 534 -1108 535 -1026
rect 569 -1027 570 -985
rect 1083 -1027 1084 -985
rect 1108 -1027 1109 -985
rect 1157 -1108 1158 -1026
rect 1160 -1027 1161 -985
rect 1850 -1027 1851 -985
rect 156 -1108 157 -1028
rect 1062 -1029 1063 -985
rect 1108 -1108 1109 -1028
rect 1122 -1029 1123 -985
rect 1136 -1029 1137 -985
rect 1528 -1108 1529 -1028
rect 1773 -1108 1774 -1028
rect 1920 -1029 1921 -985
rect 191 -1108 192 -1030
rect 236 -1031 237 -985
rect 303 -1031 304 -985
rect 345 -1108 346 -1030
rect 387 -1031 388 -985
rect 562 -1031 563 -985
rect 579 -1108 580 -1030
rect 1633 -1108 1634 -1030
rect 198 -1033 199 -985
rect 296 -1108 297 -1032
rect 380 -1033 381 -985
rect 387 -1108 388 -1032
rect 397 -1108 398 -1032
rect 912 -1108 913 -1032
rect 919 -1108 920 -1032
rect 926 -1033 927 -985
rect 940 -1033 941 -985
rect 1871 -1033 1872 -985
rect 121 -1035 122 -985
rect 198 -1108 199 -1034
rect 205 -1035 206 -985
rect 471 -1108 472 -1034
rect 499 -1108 500 -1034
rect 527 -1035 528 -985
rect 583 -1035 584 -985
rect 583 -1108 584 -1034
rect 583 -1035 584 -985
rect 583 -1108 584 -1034
rect 618 -1108 619 -1034
rect 1136 -1108 1137 -1034
rect 1139 -1108 1140 -1034
rect 1808 -1035 1809 -985
rect 100 -1037 101 -985
rect 527 -1108 528 -1036
rect 646 -1108 647 -1036
rect 849 -1037 850 -985
rect 877 -1037 878 -985
rect 898 -1108 899 -1036
rect 905 -1037 906 -985
rect 1850 -1108 1851 -1036
rect 44 -1039 45 -985
rect 100 -1108 101 -1038
rect 114 -1039 115 -985
rect 121 -1108 122 -1038
rect 219 -1108 220 -1038
rect 926 -1108 927 -1038
rect 954 -1039 955 -985
rect 1006 -1039 1007 -985
rect 1010 -1039 1011 -985
rect 1766 -1108 1767 -1038
rect 1808 -1108 1809 -1038
rect 1829 -1039 1830 -985
rect 114 -1108 115 -1040
rect 177 -1041 178 -985
rect 205 -1108 206 -1040
rect 954 -1108 955 -1040
rect 982 -1108 983 -1040
rect 996 -1041 997 -985
rect 1010 -1108 1011 -1040
rect 1052 -1041 1053 -985
rect 1059 -1041 1060 -985
rect 1549 -1041 1550 -985
rect 1591 -1041 1592 -985
rect 1829 -1108 1830 -1040
rect 177 -1108 178 -1042
rect 429 -1043 430 -985
rect 450 -1043 451 -985
rect 506 -1108 507 -1042
rect 520 -1043 521 -985
rect 569 -1108 570 -1042
rect 688 -1043 689 -985
rect 940 -1108 941 -1042
rect 961 -1043 962 -985
rect 996 -1108 997 -1042
rect 1013 -1043 1014 -985
rect 1192 -1108 1193 -1042
rect 1220 -1043 1221 -985
rect 1234 -1108 1235 -1042
rect 1297 -1108 1298 -1042
rect 1304 -1043 1305 -985
rect 1360 -1043 1361 -985
rect 1871 -1108 1872 -1042
rect 233 -1108 234 -1044
rect 450 -1108 451 -1044
rect 520 -1108 521 -1044
rect 922 -1045 923 -985
rect 985 -1045 986 -985
rect 1654 -1045 1655 -985
rect 254 -1047 255 -985
rect 303 -1108 304 -1046
rect 352 -1047 353 -985
rect 429 -1108 430 -1046
rect 688 -1108 689 -1046
rect 1153 -1047 1154 -985
rect 1206 -1047 1207 -985
rect 1220 -1108 1221 -1046
rect 1262 -1047 1263 -985
rect 1654 -1108 1655 -1046
rect 254 -1108 255 -1048
rect 324 -1049 325 -985
rect 352 -1108 353 -1048
rect 649 -1108 650 -1048
rect 695 -1049 696 -985
rect 1153 -1108 1154 -1048
rect 1199 -1049 1200 -985
rect 1206 -1108 1207 -1048
rect 1213 -1049 1214 -985
rect 1262 -1108 1263 -1048
rect 1304 -1108 1305 -1048
rect 1311 -1049 1312 -985
rect 1353 -1049 1354 -985
rect 1360 -1108 1361 -1048
rect 1472 -1108 1473 -1048
rect 1479 -1049 1480 -985
rect 1549 -1108 1550 -1048
rect 1787 -1049 1788 -985
rect 366 -1051 367 -985
rect 380 -1108 381 -1050
rect 401 -1108 402 -1050
rect 422 -1051 423 -985
rect 607 -1051 608 -985
rect 695 -1108 696 -1050
rect 723 -1051 724 -985
rect 1199 -1108 1200 -1050
rect 1213 -1108 1214 -1050
rect 1283 -1051 1284 -985
rect 1479 -1108 1480 -1050
rect 1556 -1051 1557 -985
rect 1591 -1108 1592 -1050
rect 1689 -1051 1690 -985
rect 1787 -1108 1788 -1050
rect 1815 -1051 1816 -985
rect 275 -1053 276 -985
rect 422 -1108 423 -1052
rect 653 -1053 654 -985
rect 723 -1108 724 -1052
rect 751 -1108 752 -1052
rect 856 -1053 857 -985
rect 877 -1108 878 -1052
rect 884 -1053 885 -985
rect 989 -1053 990 -985
rect 989 -1108 990 -1052
rect 989 -1053 990 -985
rect 989 -1108 990 -1052
rect 1003 -1053 1004 -985
rect 1353 -1108 1354 -1052
rect 1465 -1053 1466 -985
rect 1556 -1108 1557 -1052
rect 1563 -1053 1564 -985
rect 1689 -1108 1690 -1052
rect 1815 -1108 1816 -1052
rect 1843 -1053 1844 -985
rect 16 -1055 17 -985
rect 884 -1108 885 -1054
rect 1003 -1108 1004 -1054
rect 1045 -1055 1046 -985
rect 1048 -1108 1049 -1054
rect 1801 -1055 1802 -985
rect 16 -1108 17 -1056
rect 215 -1108 216 -1056
rect 275 -1108 276 -1056
rect 317 -1057 318 -985
rect 324 -1108 325 -1056
rect 1045 -1108 1046 -1056
rect 1052 -1108 1053 -1056
rect 1073 -1057 1074 -985
rect 1122 -1108 1123 -1056
rect 1129 -1057 1130 -985
rect 1150 -1057 1151 -985
rect 1682 -1057 1683 -985
rect 1696 -1057 1697 -985
rect 1843 -1108 1844 -1056
rect 317 -1108 318 -1058
rect 744 -1059 745 -985
rect 782 -1108 783 -1058
rect 1283 -1108 1284 -1058
rect 1563 -1108 1564 -1058
rect 1626 -1059 1627 -985
rect 1682 -1108 1683 -1058
rect 1738 -1059 1739 -985
rect 1759 -1059 1760 -985
rect 1801 -1108 1802 -1058
rect 338 -1061 339 -985
rect 1129 -1108 1130 -1060
rect 1150 -1108 1151 -1060
rect 1465 -1108 1466 -1060
rect 1626 -1108 1627 -1060
rect 1647 -1061 1648 -985
rect 1696 -1108 1697 -1060
rect 1752 -1061 1753 -985
rect 331 -1063 332 -985
rect 338 -1108 339 -1062
rect 366 -1108 367 -1062
rect 632 -1108 633 -1062
rect 744 -1108 745 -1062
rect 800 -1063 801 -985
rect 807 -1063 808 -985
rect 856 -1108 857 -1062
rect 1017 -1108 1018 -1062
rect 1738 -1108 1739 -1062
rect 135 -1065 136 -985
rect 331 -1108 332 -1064
rect 765 -1065 766 -985
rect 807 -1108 808 -1064
rect 835 -1065 836 -985
rect 905 -1108 906 -1064
rect 1031 -1065 1032 -985
rect 1759 -1108 1760 -1064
rect 135 -1108 136 -1066
rect 415 -1067 416 -985
rect 597 -1067 598 -985
rect 765 -1108 766 -1066
rect 793 -1067 794 -985
rect 961 -1108 962 -1066
rect 1038 -1067 1039 -985
rect 1101 -1067 1102 -985
rect 1227 -1067 1228 -985
rect 1311 -1108 1312 -1066
rect 1612 -1067 1613 -985
rect 1647 -1108 1648 -1066
rect 359 -1069 360 -985
rect 597 -1108 598 -1068
rect 628 -1108 629 -1068
rect 835 -1108 836 -1068
rect 842 -1108 843 -1068
rect 1115 -1069 1116 -985
rect 1227 -1108 1228 -1068
rect 1836 -1069 1837 -985
rect 359 -1108 360 -1070
rect 373 -1071 374 -985
rect 415 -1108 416 -1070
rect 464 -1071 465 -985
rect 639 -1071 640 -985
rect 793 -1108 794 -1070
rect 800 -1108 801 -1070
rect 1034 -1071 1035 -985
rect 1041 -1071 1042 -985
rect 1640 -1071 1641 -985
rect 1836 -1108 1837 -1070
rect 1857 -1071 1858 -985
rect 247 -1073 248 -985
rect 464 -1108 465 -1072
rect 639 -1108 640 -1072
rect 754 -1073 755 -985
rect 828 -1073 829 -985
rect 1101 -1108 1102 -1072
rect 1115 -1108 1116 -1072
rect 1164 -1073 1165 -985
rect 1521 -1073 1522 -985
rect 1612 -1108 1613 -1072
rect 1640 -1108 1641 -1072
rect 1661 -1073 1662 -985
rect 1822 -1073 1823 -985
rect 1857 -1108 1858 -1072
rect 184 -1075 185 -985
rect 247 -1108 248 -1074
rect 289 -1075 290 -985
rect 373 -1108 374 -1074
rect 653 -1108 654 -1074
rect 1521 -1108 1522 -1074
rect 1661 -1108 1662 -1074
rect 1703 -1075 1704 -985
rect 163 -1077 164 -985
rect 184 -1108 185 -1076
rect 212 -1077 213 -985
rect 289 -1108 290 -1076
rect 684 -1108 685 -1076
rect 1822 -1108 1823 -1076
rect 23 -1079 24 -985
rect 212 -1108 213 -1078
rect 849 -1108 850 -1078
rect 1381 -1079 1382 -985
rect 1675 -1079 1676 -985
rect 1703 -1108 1704 -1078
rect 23 -1108 24 -1080
rect 310 -1108 311 -1080
rect 947 -1081 948 -985
rect 1031 -1108 1032 -1080
rect 1059 -1108 1060 -1080
rect 1094 -1081 1095 -985
rect 1143 -1081 1144 -985
rect 1164 -1108 1165 -1080
rect 1381 -1108 1382 -1080
rect 1388 -1081 1389 -985
rect 1675 -1108 1676 -1080
rect 1731 -1081 1732 -985
rect 163 -1108 164 -1082
rect 590 -1083 591 -985
rect 947 -1108 948 -1082
rect 975 -1083 976 -985
rect 1024 -1083 1025 -985
rect 1038 -1108 1039 -1082
rect 1066 -1083 1067 -985
rect 1094 -1108 1095 -1082
rect 1143 -1108 1144 -1082
rect 1185 -1083 1186 -985
rect 1388 -1108 1389 -1082
rect 1395 -1083 1396 -985
rect 1577 -1083 1578 -985
rect 1731 -1108 1732 -1082
rect 555 -1085 556 -985
rect 590 -1108 591 -1084
rect 863 -1108 864 -1084
rect 1066 -1108 1067 -1084
rect 1073 -1108 1074 -1084
rect 1087 -1085 1088 -985
rect 1185 -1108 1186 -1084
rect 1230 -1085 1231 -985
rect 1339 -1085 1340 -985
rect 1395 -1108 1396 -1084
rect 1542 -1085 1543 -985
rect 1577 -1108 1578 -1084
rect 555 -1108 556 -1086
rect 576 -1087 577 -985
rect 740 -1087 741 -985
rect 1087 -1108 1088 -1086
rect 1332 -1087 1333 -985
rect 1339 -1108 1340 -1086
rect 1542 -1108 1543 -1086
rect 1605 -1087 1606 -985
rect 576 -1108 577 -1088
rect 1248 -1089 1249 -985
rect 1325 -1089 1326 -985
rect 1332 -1108 1333 -1088
rect 1605 -1108 1606 -1088
rect 1717 -1089 1718 -985
rect 740 -1108 741 -1090
rect 1619 -1091 1620 -985
rect 1717 -1108 1718 -1090
rect 1780 -1091 1781 -985
rect 65 -1093 66 -985
rect 1619 -1108 1620 -1092
rect 1780 -1108 1781 -1092
rect 1794 -1093 1795 -985
rect 2 -1095 3 -985
rect 65 -1108 66 -1094
rect 828 -1108 829 -1094
rect 1230 -1108 1231 -1094
rect 1248 -1108 1249 -1094
rect 1402 -1095 1403 -985
rect 1668 -1095 1669 -985
rect 1794 -1108 1795 -1094
rect 110 -1097 111 -985
rect 1668 -1108 1669 -1096
rect 933 -1099 934 -985
rect 975 -1108 976 -1098
rect 1024 -1108 1025 -1098
rect 1171 -1099 1172 -985
rect 1318 -1099 1319 -985
rect 1325 -1108 1326 -1098
rect 1402 -1108 1403 -1098
rect 1486 -1099 1487 -985
rect 572 -1108 573 -1100
rect 933 -1108 934 -1100
rect 1080 -1101 1081 -985
rect 1752 -1108 1753 -1100
rect 789 -1108 790 -1102
rect 1318 -1108 1319 -1102
rect 1486 -1108 1487 -1102
rect 1881 -1103 1882 -985
rect 814 -1105 815 -985
rect 1171 -1108 1172 -1104
rect 814 -1108 815 -1106
rect 943 -1107 944 -985
rect 1080 -1108 1081 -1106
rect 1902 -1107 1903 -985
rect 2 -1243 3 -1117
rect 72 -1118 73 -1116
rect 86 -1118 87 -1116
rect 86 -1243 87 -1117
rect 86 -1118 87 -1116
rect 86 -1243 87 -1117
rect 128 -1118 129 -1116
rect 674 -1118 675 -1116
rect 716 -1118 717 -1116
rect 929 -1243 930 -1117
rect 933 -1118 934 -1116
rect 1150 -1243 1151 -1117
rect 1153 -1118 1154 -1116
rect 1829 -1118 1830 -1116
rect 1843 -1118 1844 -1116
rect 1867 -1118 1868 -1116
rect 1878 -1118 1879 -1116
rect 1920 -1243 1921 -1117
rect 1927 -1118 1928 -1116
rect 1927 -1243 1928 -1117
rect 1927 -1118 1928 -1116
rect 1927 -1243 1928 -1117
rect 1948 -1118 1949 -1116
rect 1955 -1243 1956 -1117
rect 1976 -1118 1977 -1116
rect 1990 -1243 1991 -1117
rect 16 -1120 17 -1116
rect 222 -1120 223 -1116
rect 233 -1120 234 -1116
rect 653 -1120 654 -1116
rect 656 -1120 657 -1116
rect 772 -1120 773 -1116
rect 775 -1243 776 -1119
rect 870 -1120 871 -1116
rect 880 -1243 881 -1119
rect 1367 -1120 1368 -1116
rect 1549 -1120 1550 -1116
rect 1892 -1243 1893 -1119
rect 1969 -1120 1970 -1116
rect 1976 -1243 1977 -1119
rect 16 -1243 17 -1121
rect 114 -1122 115 -1116
rect 135 -1122 136 -1116
rect 772 -1243 773 -1121
rect 779 -1122 780 -1116
rect 856 -1122 857 -1116
rect 866 -1122 867 -1116
rect 1024 -1122 1025 -1116
rect 1045 -1122 1046 -1116
rect 1199 -1122 1200 -1116
rect 1206 -1122 1207 -1116
rect 1206 -1243 1207 -1121
rect 1206 -1122 1207 -1116
rect 1206 -1243 1207 -1121
rect 1269 -1122 1270 -1116
rect 1269 -1243 1270 -1121
rect 1269 -1122 1270 -1116
rect 1269 -1243 1270 -1121
rect 1276 -1122 1277 -1116
rect 1276 -1243 1277 -1121
rect 1276 -1122 1277 -1116
rect 1276 -1243 1277 -1121
rect 1318 -1122 1319 -1116
rect 1906 -1243 1907 -1121
rect 1962 -1122 1963 -1116
rect 1969 -1243 1970 -1121
rect 23 -1124 24 -1116
rect 565 -1124 566 -1116
rect 572 -1124 573 -1116
rect 660 -1124 661 -1116
rect 674 -1243 675 -1123
rect 702 -1124 703 -1116
rect 716 -1243 717 -1123
rect 1080 -1124 1081 -1116
rect 1122 -1124 1123 -1116
rect 1122 -1243 1123 -1123
rect 1122 -1124 1123 -1116
rect 1122 -1243 1123 -1123
rect 1132 -1243 1133 -1123
rect 1570 -1124 1571 -1116
rect 1584 -1124 1585 -1116
rect 1885 -1243 1886 -1123
rect 30 -1126 31 -1116
rect 40 -1243 41 -1125
rect 44 -1126 45 -1116
rect 933 -1243 934 -1125
rect 957 -1126 958 -1116
rect 1703 -1126 1704 -1116
rect 1759 -1126 1760 -1116
rect 1878 -1243 1879 -1125
rect 30 -1243 31 -1127
rect 198 -1128 199 -1116
rect 219 -1243 220 -1127
rect 534 -1128 535 -1116
rect 562 -1128 563 -1116
rect 842 -1128 843 -1116
rect 870 -1243 871 -1127
rect 1290 -1128 1291 -1116
rect 1311 -1128 1312 -1116
rect 1318 -1243 1319 -1127
rect 1367 -1243 1368 -1127
rect 1388 -1128 1389 -1116
rect 1451 -1128 1452 -1116
rect 1570 -1243 1571 -1127
rect 1591 -1128 1592 -1116
rect 1759 -1243 1760 -1127
rect 1766 -1128 1767 -1116
rect 1766 -1243 1767 -1127
rect 1766 -1128 1767 -1116
rect 1766 -1243 1767 -1127
rect 1773 -1128 1774 -1116
rect 1773 -1243 1774 -1127
rect 1773 -1128 1774 -1116
rect 1773 -1243 1774 -1127
rect 1780 -1128 1781 -1116
rect 1899 -1243 1900 -1127
rect 61 -1243 62 -1129
rect 268 -1130 269 -1116
rect 282 -1130 283 -1116
rect 754 -1130 755 -1116
rect 758 -1243 759 -1129
rect 1003 -1130 1004 -1116
rect 1010 -1130 1011 -1116
rect 1024 -1243 1025 -1129
rect 1045 -1243 1046 -1129
rect 1731 -1130 1732 -1116
rect 1780 -1243 1781 -1129
rect 1787 -1130 1788 -1116
rect 1808 -1130 1809 -1116
rect 1829 -1243 1830 -1129
rect 1836 -1130 1837 -1116
rect 1843 -1243 1844 -1129
rect 1871 -1130 1872 -1116
rect 1962 -1243 1963 -1129
rect 65 -1132 66 -1116
rect 527 -1132 528 -1116
rect 562 -1243 563 -1131
rect 1230 -1132 1231 -1116
rect 1360 -1132 1361 -1116
rect 1388 -1243 1389 -1131
rect 1500 -1132 1501 -1116
rect 1549 -1243 1550 -1131
rect 1591 -1243 1592 -1131
rect 1598 -1132 1599 -1116
rect 1689 -1132 1690 -1116
rect 1731 -1243 1732 -1131
rect 1787 -1243 1788 -1131
rect 1801 -1132 1802 -1116
rect 1822 -1132 1823 -1116
rect 1864 -1132 1865 -1116
rect 65 -1243 66 -1133
rect 415 -1134 416 -1116
rect 422 -1134 423 -1116
rect 453 -1134 454 -1116
rect 464 -1134 465 -1116
rect 681 -1134 682 -1116
rect 695 -1134 696 -1116
rect 702 -1243 703 -1133
rect 730 -1134 731 -1116
rect 747 -1134 748 -1116
rect 751 -1134 752 -1116
rect 1451 -1243 1452 -1133
rect 1458 -1134 1459 -1116
rect 1500 -1243 1501 -1133
rect 1542 -1134 1543 -1116
rect 1871 -1243 1872 -1133
rect 72 -1243 73 -1135
rect 394 -1136 395 -1116
rect 401 -1136 402 -1116
rect 401 -1243 402 -1135
rect 401 -1136 402 -1116
rect 401 -1243 402 -1135
rect 415 -1243 416 -1135
rect 586 -1243 587 -1135
rect 625 -1136 626 -1116
rect 653 -1243 654 -1135
rect 660 -1243 661 -1135
rect 975 -1136 976 -1116
rect 996 -1136 997 -1116
rect 1010 -1243 1011 -1135
rect 1017 -1136 1018 -1116
rect 1577 -1136 1578 -1116
rect 1598 -1243 1599 -1135
rect 1612 -1136 1613 -1116
rect 1682 -1136 1683 -1116
rect 1822 -1243 1823 -1135
rect 100 -1138 101 -1116
rect 128 -1243 129 -1137
rect 131 -1138 132 -1116
rect 681 -1243 682 -1137
rect 695 -1243 696 -1137
rect 723 -1138 724 -1116
rect 730 -1243 731 -1137
rect 765 -1138 766 -1116
rect 782 -1138 783 -1116
rect 1262 -1138 1263 -1116
rect 1423 -1138 1424 -1116
rect 1682 -1243 1683 -1137
rect 1696 -1138 1697 -1116
rect 1836 -1243 1837 -1137
rect 9 -1140 10 -1116
rect 100 -1243 101 -1139
rect 114 -1243 115 -1139
rect 789 -1140 790 -1116
rect 810 -1243 811 -1139
rect 1031 -1140 1032 -1116
rect 1080 -1243 1081 -1139
rect 1101 -1140 1102 -1116
rect 1139 -1140 1140 -1116
rect 1192 -1140 1193 -1116
rect 1402 -1140 1403 -1116
rect 1423 -1243 1424 -1139
rect 1458 -1243 1459 -1139
rect 1486 -1140 1487 -1116
rect 1493 -1140 1494 -1116
rect 1542 -1243 1543 -1139
rect 1563 -1140 1564 -1116
rect 1577 -1243 1578 -1139
rect 1605 -1140 1606 -1116
rect 1689 -1243 1690 -1139
rect 1724 -1140 1725 -1116
rect 1864 -1243 1865 -1139
rect 9 -1243 10 -1141
rect 425 -1243 426 -1141
rect 429 -1142 430 -1116
rect 856 -1243 857 -1141
rect 859 -1243 860 -1141
rect 1262 -1243 1263 -1141
rect 1381 -1142 1382 -1116
rect 1402 -1243 1403 -1141
rect 1444 -1142 1445 -1116
rect 1493 -1243 1494 -1141
rect 1521 -1142 1522 -1116
rect 1696 -1243 1697 -1141
rect 1794 -1142 1795 -1116
rect 1808 -1243 1809 -1141
rect 79 -1243 80 -1143
rect 1563 -1243 1564 -1143
rect 1605 -1243 1606 -1143
rect 1626 -1144 1627 -1116
rect 1668 -1144 1669 -1116
rect 1724 -1243 1725 -1143
rect 1752 -1144 1753 -1116
rect 1794 -1243 1795 -1143
rect 121 -1146 122 -1116
rect 135 -1243 136 -1145
rect 159 -1243 160 -1145
rect 310 -1243 311 -1145
rect 331 -1146 332 -1116
rect 534 -1243 535 -1145
rect 555 -1146 556 -1116
rect 625 -1243 626 -1145
rect 723 -1243 724 -1145
rect 744 -1146 745 -1116
rect 761 -1146 762 -1116
rect 1290 -1243 1291 -1145
rect 1444 -1243 1445 -1145
rect 1479 -1146 1480 -1116
rect 1486 -1243 1487 -1145
rect 1556 -1146 1557 -1116
rect 1612 -1243 1613 -1145
rect 1633 -1146 1634 -1116
rect 1668 -1243 1669 -1145
rect 1815 -1146 1816 -1116
rect 121 -1243 122 -1147
rect 782 -1243 783 -1147
rect 814 -1148 815 -1116
rect 842 -1243 843 -1147
rect 863 -1148 864 -1116
rect 1381 -1243 1382 -1147
rect 1437 -1148 1438 -1116
rect 1479 -1243 1480 -1147
rect 1507 -1148 1508 -1116
rect 1556 -1243 1557 -1147
rect 1626 -1243 1627 -1147
rect 1640 -1148 1641 -1116
rect 1745 -1148 1746 -1116
rect 1752 -1243 1753 -1147
rect 180 -1243 181 -1149
rect 852 -1150 853 -1116
rect 863 -1243 864 -1149
rect 877 -1150 878 -1116
rect 894 -1150 895 -1116
rect 1647 -1150 1648 -1116
rect 1717 -1150 1718 -1116
rect 1745 -1243 1746 -1149
rect 184 -1152 185 -1116
rect 184 -1243 185 -1151
rect 184 -1152 185 -1116
rect 184 -1243 185 -1151
rect 198 -1243 199 -1151
rect 317 -1152 318 -1116
rect 359 -1152 360 -1116
rect 628 -1152 629 -1116
rect 670 -1243 671 -1151
rect 1507 -1243 1508 -1151
rect 1514 -1152 1515 -1116
rect 1640 -1243 1641 -1151
rect 1647 -1243 1648 -1151
rect 1675 -1152 1676 -1116
rect 1717 -1243 1718 -1151
rect 1738 -1152 1739 -1116
rect 82 -1154 83 -1116
rect 317 -1243 318 -1153
rect 359 -1243 360 -1153
rect 380 -1154 381 -1116
rect 422 -1243 423 -1153
rect 1129 -1154 1130 -1116
rect 1136 -1154 1137 -1116
rect 1675 -1243 1676 -1153
rect 1710 -1154 1711 -1116
rect 1738 -1243 1739 -1153
rect 233 -1243 234 -1155
rect 247 -1156 248 -1116
rect 261 -1156 262 -1116
rect 292 -1243 293 -1155
rect 303 -1156 304 -1116
rect 331 -1243 332 -1155
rect 366 -1156 367 -1116
rect 369 -1208 370 -1155
rect 373 -1156 374 -1116
rect 394 -1243 395 -1155
rect 436 -1156 437 -1116
rect 523 -1156 524 -1116
rect 555 -1243 556 -1155
rect 667 -1156 668 -1116
rect 684 -1156 685 -1116
rect 1815 -1243 1816 -1155
rect 51 -1158 52 -1116
rect 373 -1243 374 -1157
rect 380 -1243 381 -1157
rect 800 -1158 801 -1116
rect 873 -1243 874 -1157
rect 1584 -1243 1585 -1157
rect 1633 -1243 1634 -1157
rect 1661 -1158 1662 -1116
rect 51 -1243 52 -1159
rect 740 -1160 741 -1116
rect 779 -1243 780 -1159
rect 1437 -1243 1438 -1159
rect 1465 -1160 1466 -1116
rect 1514 -1243 1515 -1159
rect 1521 -1243 1522 -1159
rect 1654 -1160 1655 -1116
rect 240 -1162 241 -1116
rect 247 -1243 248 -1161
rect 268 -1243 269 -1161
rect 275 -1162 276 -1116
rect 282 -1243 283 -1161
rect 345 -1162 346 -1116
rect 366 -1243 367 -1161
rect 436 -1243 437 -1161
rect 912 -1162 913 -1116
rect 926 -1162 927 -1116
rect 1360 -1243 1361 -1161
rect 1472 -1162 1473 -1116
rect 1654 -1243 1655 -1161
rect 163 -1164 164 -1116
rect 345 -1243 346 -1163
rect 352 -1164 353 -1116
rect 926 -1243 927 -1163
rect 975 -1243 976 -1163
rect 982 -1164 983 -1116
rect 989 -1164 990 -1116
rect 996 -1243 997 -1163
rect 1003 -1243 1004 -1163
rect 1220 -1164 1221 -1116
rect 1248 -1164 1249 -1116
rect 1472 -1243 1473 -1163
rect 1535 -1164 1536 -1116
rect 1661 -1243 1662 -1163
rect 58 -1166 59 -1116
rect 352 -1243 353 -1165
rect 446 -1243 447 -1165
rect 1703 -1243 1704 -1165
rect 163 -1243 164 -1167
rect 457 -1168 458 -1116
rect 464 -1243 465 -1167
rect 541 -1168 542 -1116
rect 583 -1168 584 -1116
rect 786 -1243 787 -1167
rect 912 -1243 913 -1167
rect 1129 -1243 1130 -1167
rect 1160 -1243 1161 -1167
rect 1913 -1243 1914 -1167
rect 142 -1170 143 -1116
rect 541 -1243 542 -1169
rect 583 -1243 584 -1169
rect 1031 -1243 1032 -1169
rect 1038 -1170 1039 -1116
rect 1220 -1243 1221 -1169
rect 1241 -1170 1242 -1116
rect 1248 -1243 1249 -1169
rect 142 -1243 143 -1171
rect 229 -1243 230 -1171
rect 240 -1243 241 -1171
rect 296 -1172 297 -1116
rect 303 -1243 304 -1171
rect 908 -1243 909 -1171
rect 961 -1172 962 -1116
rect 989 -1243 990 -1171
rect 1017 -1243 1018 -1171
rect 1465 -1243 1466 -1171
rect 254 -1174 255 -1116
rect 296 -1243 297 -1173
rect 313 -1174 314 -1116
rect 1136 -1243 1137 -1173
rect 1164 -1174 1165 -1116
rect 1192 -1243 1193 -1173
rect 1234 -1174 1235 -1116
rect 1241 -1243 1242 -1173
rect 212 -1176 213 -1116
rect 254 -1243 255 -1175
rect 275 -1243 276 -1175
rect 338 -1176 339 -1116
rect 450 -1176 451 -1116
rect 1801 -1243 1802 -1175
rect 37 -1178 38 -1116
rect 450 -1243 451 -1177
rect 453 -1243 454 -1177
rect 1199 -1243 1200 -1177
rect 1213 -1178 1214 -1116
rect 1234 -1243 1235 -1177
rect 289 -1180 290 -1116
rect 576 -1180 577 -1116
rect 590 -1180 591 -1116
rect 814 -1243 815 -1179
rect 849 -1180 850 -1116
rect 1038 -1243 1039 -1179
rect 1048 -1180 1049 -1116
rect 1710 -1243 1711 -1179
rect 107 -1182 108 -1116
rect 1048 -1243 1049 -1181
rect 1087 -1182 1088 -1116
rect 1311 -1243 1312 -1181
rect 107 -1243 108 -1183
rect 891 -1184 892 -1116
rect 982 -1243 983 -1183
rect 1052 -1184 1053 -1116
rect 1059 -1184 1060 -1116
rect 1087 -1243 1088 -1183
rect 1094 -1184 1095 -1116
rect 1101 -1243 1102 -1183
rect 1115 -1184 1116 -1116
rect 1164 -1243 1165 -1183
rect 156 -1186 157 -1116
rect 590 -1243 591 -1185
rect 632 -1186 633 -1116
rect 1535 -1243 1536 -1185
rect 324 -1188 325 -1116
rect 632 -1243 633 -1187
rect 667 -1243 668 -1187
rect 1528 -1188 1529 -1116
rect 324 -1243 325 -1189
rect 485 -1190 486 -1116
rect 516 -1243 517 -1189
rect 1227 -1243 1228 -1189
rect 338 -1243 339 -1191
rect 604 -1192 605 -1116
rect 709 -1192 710 -1116
rect 800 -1243 801 -1191
rect 821 -1192 822 -1116
rect 849 -1243 850 -1191
rect 877 -1243 878 -1191
rect 1059 -1243 1060 -1191
rect 1108 -1192 1109 -1116
rect 1115 -1243 1116 -1191
rect 1157 -1192 1158 -1116
rect 1213 -1243 1214 -1191
rect 37 -1243 38 -1193
rect 604 -1243 605 -1193
rect 709 -1243 710 -1193
rect 807 -1194 808 -1116
rect 891 -1243 892 -1193
rect 898 -1194 899 -1116
rect 1052 -1243 1053 -1193
rect 1066 -1194 1067 -1116
rect 1108 -1243 1109 -1193
rect 1283 -1194 1284 -1116
rect 408 -1196 409 -1116
rect 1283 -1243 1284 -1195
rect 408 -1243 409 -1197
rect 688 -1198 689 -1116
rect 733 -1198 734 -1116
rect 1850 -1198 1851 -1116
rect 443 -1200 444 -1116
rect 1094 -1243 1095 -1199
rect 1157 -1243 1158 -1199
rect 1409 -1200 1410 -1116
rect 212 -1243 213 -1201
rect 443 -1243 444 -1201
rect 457 -1243 458 -1201
rect 506 -1202 507 -1116
rect 576 -1243 577 -1201
rect 618 -1202 619 -1116
rect 737 -1202 738 -1116
rect 1178 -1202 1179 -1116
rect 1181 -1243 1182 -1201
rect 1850 -1243 1851 -1201
rect 44 -1243 45 -1203
rect 1178 -1243 1179 -1203
rect 1185 -1204 1186 -1116
rect 1528 -1243 1529 -1203
rect 289 -1243 290 -1205
rect 618 -1243 619 -1205
rect 744 -1243 745 -1205
rect 821 -1243 822 -1205
rect 898 -1243 899 -1205
rect 905 -1206 906 -1116
rect 1066 -1243 1067 -1205
rect 1073 -1206 1074 -1116
rect 1143 -1206 1144 -1116
rect 1185 -1243 1186 -1205
rect 1395 -1206 1396 -1116
rect 1409 -1243 1410 -1205
rect 471 -1208 472 -1116
rect 527 -1243 528 -1207
rect 611 -1208 612 -1116
rect 688 -1243 689 -1207
rect 747 -1243 748 -1207
rect 765 -1243 766 -1207
rect 807 -1243 808 -1207
rect 954 -1208 955 -1116
rect 1143 -1243 1144 -1207
rect 1255 -1208 1256 -1116
rect 1374 -1208 1375 -1116
rect 1395 -1243 1396 -1207
rect 429 -1243 430 -1209
rect 471 -1243 472 -1209
rect 474 -1243 475 -1209
rect 499 -1210 500 -1116
rect 506 -1243 507 -1209
rect 639 -1210 640 -1116
rect 905 -1243 906 -1209
rect 1857 -1210 1858 -1116
rect 124 -1243 125 -1211
rect 499 -1243 500 -1211
rect 513 -1212 514 -1116
rect 737 -1243 738 -1211
rect 940 -1212 941 -1116
rect 1073 -1243 1074 -1211
rect 1255 -1243 1256 -1211
rect 1339 -1212 1340 -1116
rect 1353 -1212 1354 -1116
rect 1374 -1243 1375 -1211
rect 1619 -1212 1620 -1116
rect 1857 -1243 1858 -1211
rect 82 -1243 83 -1213
rect 1619 -1243 1620 -1213
rect 478 -1216 479 -1116
rect 751 -1243 752 -1215
rect 940 -1243 941 -1215
rect 964 -1243 965 -1215
rect 1325 -1216 1326 -1116
rect 1339 -1243 1340 -1215
rect 1346 -1216 1347 -1116
rect 1353 -1243 1354 -1215
rect 177 -1218 178 -1116
rect 478 -1243 479 -1217
rect 485 -1243 486 -1217
rect 548 -1218 549 -1116
rect 579 -1218 580 -1116
rect 611 -1243 612 -1217
rect 947 -1218 948 -1116
rect 954 -1243 955 -1217
rect 1297 -1218 1298 -1116
rect 1325 -1243 1326 -1217
rect 1332 -1218 1333 -1116
rect 1346 -1243 1347 -1217
rect 177 -1243 178 -1219
rect 1171 -1220 1172 -1116
rect 1297 -1243 1298 -1219
rect 1304 -1220 1305 -1116
rect 520 -1222 521 -1116
rect 1171 -1243 1172 -1221
rect 1304 -1243 1305 -1221
rect 1430 -1222 1431 -1116
rect 93 -1224 94 -1116
rect 520 -1243 521 -1223
rect 548 -1243 549 -1223
rect 968 -1224 969 -1116
rect 1416 -1224 1417 -1116
rect 1430 -1243 1431 -1223
rect 47 -1226 48 -1116
rect 1416 -1243 1417 -1225
rect 93 -1243 94 -1227
rect 149 -1228 150 -1116
rect 569 -1228 570 -1116
rect 1332 -1243 1333 -1227
rect 149 -1243 150 -1229
rect 205 -1230 206 -1116
rect 492 -1230 493 -1116
rect 569 -1243 570 -1229
rect 597 -1230 598 -1116
rect 639 -1243 640 -1229
rect 828 -1230 829 -1116
rect 968 -1243 969 -1229
rect 58 -1243 59 -1231
rect 597 -1243 598 -1231
rect 828 -1243 829 -1231
rect 884 -1232 885 -1116
rect 919 -1232 920 -1116
rect 947 -1243 948 -1231
rect 191 -1234 192 -1116
rect 205 -1243 206 -1233
rect 492 -1243 493 -1233
rect 1020 -1234 1021 -1116
rect 170 -1236 171 -1116
rect 191 -1243 192 -1235
rect 646 -1236 647 -1116
rect 919 -1243 920 -1235
rect 170 -1243 171 -1237
rect 646 -1243 647 -1237
rect 835 -1238 836 -1116
rect 884 -1243 885 -1237
rect 793 -1240 794 -1116
rect 835 -1243 836 -1239
rect 226 -1242 227 -1116
rect 793 -1243 794 -1241
rect 16 -1253 17 -1251
rect 16 -1386 17 -1252
rect 16 -1253 17 -1251
rect 16 -1386 17 -1252
rect 23 -1386 24 -1252
rect 93 -1253 94 -1251
rect 107 -1253 108 -1251
rect 145 -1386 146 -1252
rect 163 -1253 164 -1251
rect 226 -1253 227 -1251
rect 247 -1253 248 -1251
rect 261 -1253 262 -1251
rect 282 -1253 283 -1251
rect 453 -1253 454 -1251
rect 457 -1253 458 -1251
rect 670 -1253 671 -1251
rect 688 -1253 689 -1251
rect 779 -1253 780 -1251
rect 793 -1253 794 -1251
rect 1076 -1386 1077 -1252
rect 1101 -1253 1102 -1251
rect 1101 -1386 1102 -1252
rect 1101 -1253 1102 -1251
rect 1101 -1386 1102 -1252
rect 1111 -1386 1112 -1252
rect 1878 -1253 1879 -1251
rect 1906 -1253 1907 -1251
rect 1948 -1386 1949 -1252
rect 1962 -1253 1963 -1251
rect 1997 -1386 1998 -1252
rect 30 -1255 31 -1251
rect 446 -1255 447 -1251
rect 457 -1386 458 -1254
rect 597 -1255 598 -1251
rect 628 -1386 629 -1254
rect 786 -1255 787 -1251
rect 821 -1255 822 -1251
rect 1066 -1255 1067 -1251
rect 1129 -1255 1130 -1251
rect 1822 -1255 1823 -1251
rect 1843 -1255 1844 -1251
rect 1906 -1386 1907 -1254
rect 1913 -1255 1914 -1251
rect 1941 -1386 1942 -1254
rect 1969 -1255 1970 -1251
rect 1969 -1386 1970 -1254
rect 1969 -1255 1970 -1251
rect 1969 -1386 1970 -1254
rect 1976 -1255 1977 -1251
rect 1983 -1386 1984 -1254
rect 1990 -1255 1991 -1251
rect 1990 -1386 1991 -1254
rect 1990 -1255 1991 -1251
rect 1990 -1386 1991 -1254
rect 30 -1386 31 -1256
rect 208 -1386 209 -1256
rect 226 -1386 227 -1256
rect 513 -1257 514 -1251
rect 541 -1257 542 -1251
rect 597 -1386 598 -1256
rect 604 -1257 605 -1251
rect 821 -1386 822 -1256
rect 838 -1386 839 -1256
rect 1472 -1257 1473 -1251
rect 1675 -1257 1676 -1251
rect 1843 -1386 1844 -1256
rect 1920 -1257 1921 -1251
rect 1934 -1386 1935 -1256
rect 1955 -1257 1956 -1251
rect 1976 -1386 1977 -1256
rect 37 -1386 38 -1258
rect 44 -1259 45 -1251
rect 58 -1259 59 -1251
rect 793 -1386 794 -1258
rect 856 -1259 857 -1251
rect 1759 -1259 1760 -1251
rect 1927 -1259 1928 -1251
rect 1927 -1386 1928 -1258
rect 1927 -1259 1928 -1251
rect 1927 -1386 1928 -1258
rect 40 -1261 41 -1251
rect 1654 -1261 1655 -1251
rect 1689 -1261 1690 -1251
rect 1689 -1386 1690 -1260
rect 1689 -1261 1690 -1251
rect 1689 -1386 1690 -1260
rect 1759 -1386 1760 -1260
rect 1913 -1386 1914 -1260
rect 44 -1386 45 -1262
rect 576 -1263 577 -1251
rect 586 -1263 587 -1251
rect 849 -1263 850 -1251
rect 856 -1386 857 -1262
rect 873 -1263 874 -1251
rect 908 -1263 909 -1251
rect 1220 -1263 1221 -1251
rect 1269 -1263 1270 -1251
rect 1272 -1317 1273 -1262
rect 1290 -1263 1291 -1251
rect 1920 -1386 1921 -1262
rect 58 -1386 59 -1264
rect 1857 -1265 1858 -1251
rect 61 -1267 62 -1251
rect 1521 -1267 1522 -1251
rect 1612 -1267 1613 -1251
rect 1654 -1386 1655 -1266
rect 1787 -1267 1788 -1251
rect 1857 -1386 1858 -1266
rect 65 -1269 66 -1251
rect 282 -1386 283 -1268
rect 289 -1386 290 -1268
rect 401 -1269 402 -1251
rect 415 -1269 416 -1251
rect 513 -1386 514 -1268
rect 562 -1269 563 -1251
rect 1073 -1269 1074 -1251
rect 1129 -1386 1130 -1268
rect 1136 -1269 1137 -1251
rect 1150 -1269 1151 -1251
rect 1150 -1386 1151 -1268
rect 1150 -1269 1151 -1251
rect 1150 -1386 1151 -1268
rect 1178 -1269 1179 -1251
rect 1885 -1269 1886 -1251
rect 51 -1271 52 -1251
rect 65 -1386 66 -1270
rect 79 -1271 80 -1251
rect 338 -1271 339 -1251
rect 352 -1271 353 -1251
rect 656 -1386 657 -1270
rect 688 -1386 689 -1270
rect 723 -1271 724 -1251
rect 730 -1271 731 -1251
rect 730 -1386 731 -1270
rect 730 -1271 731 -1251
rect 730 -1386 731 -1270
rect 775 -1271 776 -1251
rect 1850 -1271 1851 -1251
rect 9 -1273 10 -1251
rect 79 -1386 80 -1272
rect 82 -1273 83 -1251
rect 604 -1386 605 -1272
rect 646 -1273 647 -1251
rect 1132 -1273 1133 -1251
rect 1171 -1273 1172 -1251
rect 1178 -1386 1179 -1272
rect 1220 -1386 1221 -1272
rect 1234 -1273 1235 -1251
rect 1269 -1386 1270 -1272
rect 1276 -1273 1277 -1251
rect 1290 -1386 1291 -1272
rect 1297 -1273 1298 -1251
rect 1388 -1273 1389 -1251
rect 1391 -1273 1392 -1251
rect 1430 -1273 1431 -1251
rect 1430 -1386 1431 -1272
rect 1430 -1273 1431 -1251
rect 1430 -1386 1431 -1272
rect 1458 -1273 1459 -1251
rect 1472 -1386 1473 -1272
rect 1542 -1273 1543 -1251
rect 1612 -1386 1613 -1272
rect 1626 -1273 1627 -1251
rect 1675 -1386 1676 -1272
rect 1787 -1386 1788 -1272
rect 1916 -1386 1917 -1272
rect 9 -1386 10 -1274
rect 800 -1275 801 -1251
rect 824 -1275 825 -1251
rect 849 -1386 850 -1274
rect 870 -1386 871 -1274
rect 912 -1275 913 -1251
rect 922 -1386 923 -1274
rect 1892 -1275 1893 -1251
rect 2 -1277 3 -1251
rect 800 -1386 801 -1276
rect 912 -1386 913 -1276
rect 1108 -1277 1109 -1251
rect 1122 -1277 1123 -1251
rect 1136 -1386 1137 -1276
rect 1171 -1386 1172 -1276
rect 1521 -1386 1522 -1276
rect 1808 -1277 1809 -1251
rect 1850 -1386 1851 -1276
rect 86 -1279 87 -1251
rect 170 -1279 171 -1251
rect 177 -1279 178 -1251
rect 611 -1279 612 -1251
rect 681 -1279 682 -1251
rect 723 -1386 724 -1278
rect 779 -1386 780 -1278
rect 1069 -1386 1070 -1278
rect 1073 -1386 1074 -1278
rect 1661 -1279 1662 -1251
rect 1829 -1279 1830 -1251
rect 1885 -1386 1886 -1278
rect 54 -1386 55 -1280
rect 86 -1386 87 -1280
rect 93 -1386 94 -1280
rect 142 -1281 143 -1251
rect 149 -1281 150 -1251
rect 177 -1386 178 -1280
rect 247 -1386 248 -1280
rect 1094 -1281 1095 -1251
rect 1234 -1386 1235 -1280
rect 1262 -1281 1263 -1251
rect 1297 -1386 1298 -1280
rect 1332 -1281 1333 -1251
rect 1388 -1386 1389 -1280
rect 1409 -1281 1410 -1251
rect 1437 -1281 1438 -1251
rect 1458 -1386 1459 -1280
rect 1486 -1281 1487 -1251
rect 1626 -1386 1627 -1280
rect 1773 -1281 1774 -1251
rect 1829 -1386 1830 -1280
rect 107 -1386 108 -1282
rect 548 -1283 549 -1251
rect 611 -1386 612 -1282
rect 618 -1283 619 -1251
rect 653 -1283 654 -1251
rect 681 -1386 682 -1282
rect 877 -1283 878 -1251
rect 1122 -1386 1123 -1282
rect 1143 -1283 1144 -1251
rect 1262 -1386 1263 -1282
rect 1416 -1283 1417 -1251
rect 1437 -1386 1438 -1282
rect 1479 -1283 1480 -1251
rect 1486 -1386 1487 -1282
rect 1493 -1283 1494 -1251
rect 1542 -1386 1543 -1282
rect 1591 -1283 1592 -1251
rect 1661 -1386 1662 -1282
rect 1745 -1283 1746 -1251
rect 1773 -1386 1774 -1282
rect 110 -1386 111 -1284
rect 1822 -1386 1823 -1284
rect 121 -1386 122 -1286
rect 229 -1287 230 -1251
rect 254 -1287 255 -1251
rect 579 -1386 580 -1286
rect 618 -1386 619 -1286
rect 891 -1287 892 -1251
rect 926 -1287 927 -1251
rect 1878 -1386 1879 -1286
rect 135 -1289 136 -1251
rect 135 -1386 136 -1288
rect 135 -1289 136 -1251
rect 135 -1386 136 -1288
rect 152 -1386 153 -1288
rect 261 -1386 262 -1288
rect 296 -1289 297 -1251
rect 299 -1317 300 -1288
rect 317 -1289 318 -1251
rect 541 -1386 542 -1288
rect 548 -1386 549 -1288
rect 940 -1289 941 -1251
rect 964 -1289 965 -1251
rect 1682 -1289 1683 -1251
rect 156 -1291 157 -1251
rect 1892 -1386 1893 -1290
rect 156 -1386 157 -1292
rect 660 -1293 661 -1251
rect 712 -1386 713 -1292
rect 1682 -1386 1683 -1292
rect 128 -1295 129 -1251
rect 660 -1386 661 -1294
rect 877 -1386 878 -1294
rect 1024 -1295 1025 -1251
rect 1038 -1295 1039 -1251
rect 1157 -1386 1158 -1294
rect 1244 -1386 1245 -1294
rect 1493 -1386 1494 -1294
rect 1563 -1295 1564 -1251
rect 1591 -1386 1592 -1294
rect 1605 -1295 1606 -1251
rect 1745 -1386 1746 -1294
rect 75 -1386 76 -1296
rect 1024 -1386 1025 -1296
rect 1045 -1386 1046 -1296
rect 1087 -1297 1088 -1251
rect 1094 -1386 1095 -1296
rect 1115 -1297 1116 -1251
rect 1143 -1386 1144 -1296
rect 1185 -1297 1186 -1251
rect 1255 -1297 1256 -1251
rect 1332 -1386 1333 -1296
rect 1416 -1386 1417 -1296
rect 1423 -1297 1424 -1251
rect 1465 -1297 1466 -1251
rect 1479 -1386 1480 -1296
rect 124 -1299 125 -1251
rect 1087 -1386 1088 -1298
rect 1185 -1386 1186 -1298
rect 1836 -1299 1837 -1251
rect 128 -1386 129 -1300
rect 842 -1301 843 -1251
rect 891 -1386 892 -1300
rect 947 -1301 948 -1251
rect 961 -1301 962 -1251
rect 1038 -1386 1039 -1300
rect 1055 -1386 1056 -1300
rect 1808 -1386 1809 -1300
rect 163 -1386 164 -1302
rect 240 -1303 241 -1251
rect 254 -1386 255 -1302
rect 670 -1386 671 -1302
rect 842 -1386 843 -1302
rect 898 -1303 899 -1251
rect 929 -1303 930 -1251
rect 1605 -1386 1606 -1302
rect 1780 -1303 1781 -1251
rect 1836 -1386 1837 -1302
rect 170 -1386 171 -1304
rect 380 -1305 381 -1251
rect 394 -1305 395 -1251
rect 425 -1305 426 -1251
rect 443 -1305 444 -1251
rect 1311 -1305 1312 -1251
rect 1423 -1386 1424 -1304
rect 1507 -1305 1508 -1251
rect 1766 -1305 1767 -1251
rect 1780 -1386 1781 -1304
rect 205 -1307 206 -1251
rect 240 -1386 241 -1306
rect 268 -1307 269 -1251
rect 394 -1386 395 -1306
rect 401 -1386 402 -1306
rect 555 -1307 556 -1251
rect 807 -1307 808 -1251
rect 898 -1386 899 -1306
rect 929 -1386 930 -1306
rect 1563 -1386 1564 -1306
rect 1752 -1307 1753 -1251
rect 1766 -1386 1767 -1306
rect 184 -1309 185 -1251
rect 205 -1386 206 -1308
rect 233 -1309 234 -1251
rect 268 -1386 269 -1308
rect 296 -1386 297 -1308
rect 338 -1386 339 -1308
rect 408 -1309 409 -1251
rect 422 -1309 423 -1251
rect 1801 -1309 1802 -1251
rect 184 -1386 185 -1310
rect 303 -1311 304 -1251
rect 310 -1311 311 -1251
rect 555 -1386 556 -1310
rect 807 -1386 808 -1310
rect 1080 -1311 1081 -1251
rect 1108 -1386 1109 -1310
rect 1507 -1386 1508 -1310
rect 1696 -1311 1697 -1251
rect 1752 -1386 1753 -1310
rect 100 -1313 101 -1251
rect 310 -1386 311 -1312
rect 317 -1386 318 -1312
rect 387 -1313 388 -1251
rect 408 -1386 409 -1312
rect 520 -1313 521 -1251
rect 534 -1313 535 -1251
rect 562 -1386 563 -1312
rect 810 -1313 811 -1251
rect 1801 -1386 1802 -1312
rect 72 -1315 73 -1251
rect 387 -1386 388 -1314
rect 422 -1386 423 -1314
rect 667 -1315 668 -1251
rect 947 -1386 948 -1314
rect 954 -1315 955 -1251
rect 961 -1386 962 -1314
rect 989 -1315 990 -1251
rect 1017 -1315 1018 -1251
rect 1871 -1315 1872 -1251
rect 51 -1386 52 -1316
rect 667 -1386 668 -1316
rect 954 -1386 955 -1316
rect 975 -1317 976 -1251
rect 989 -1386 990 -1316
rect 1031 -1317 1032 -1251
rect 1066 -1386 1067 -1316
rect 1311 -1386 1312 -1316
rect 1391 -1386 1392 -1316
rect 1409 -1386 1410 -1316
rect 1451 -1317 1452 -1251
rect 1465 -1386 1466 -1316
rect 1668 -1317 1669 -1251
rect 1871 -1386 1872 -1316
rect 72 -1386 73 -1318
rect 569 -1319 570 -1251
rect 968 -1319 969 -1251
rect 1115 -1386 1116 -1318
rect 1255 -1386 1256 -1318
rect 1374 -1319 1375 -1251
rect 1598 -1319 1599 -1251
rect 1668 -1386 1669 -1318
rect 1696 -1386 1697 -1318
rect 1703 -1319 1704 -1251
rect 100 -1386 101 -1320
rect 264 -1321 265 -1251
rect 352 -1386 353 -1320
rect 359 -1321 360 -1251
rect 366 -1321 367 -1251
rect 380 -1386 381 -1320
rect 443 -1386 444 -1320
rect 772 -1321 773 -1251
rect 968 -1386 969 -1320
rect 1020 -1321 1021 -1251
rect 1031 -1386 1032 -1320
rect 1325 -1321 1326 -1251
rect 1360 -1321 1361 -1251
rect 1451 -1386 1452 -1320
rect 142 -1386 143 -1322
rect 303 -1386 304 -1322
rect 324 -1323 325 -1251
rect 359 -1386 360 -1322
rect 366 -1386 367 -1322
rect 516 -1323 517 -1251
rect 534 -1386 535 -1322
rect 765 -1323 766 -1251
rect 772 -1386 773 -1322
rect 814 -1323 815 -1251
rect 975 -1386 976 -1322
rect 982 -1323 983 -1251
rect 996 -1323 997 -1251
rect 1017 -1386 1018 -1322
rect 1080 -1386 1081 -1322
rect 1164 -1323 1165 -1251
rect 1304 -1323 1305 -1251
rect 1360 -1386 1361 -1322
rect 1374 -1386 1375 -1322
rect 1395 -1323 1396 -1251
rect 1444 -1323 1445 -1251
rect 1598 -1386 1599 -1322
rect 233 -1386 234 -1324
rect 492 -1325 493 -1251
rect 530 -1386 531 -1324
rect 1444 -1386 1445 -1324
rect 275 -1327 276 -1251
rect 324 -1386 325 -1326
rect 373 -1327 374 -1251
rect 415 -1386 416 -1326
rect 450 -1327 451 -1251
rect 814 -1386 815 -1326
rect 859 -1327 860 -1251
rect 1304 -1386 1305 -1326
rect 1325 -1386 1326 -1326
rect 1339 -1327 1340 -1251
rect 212 -1329 213 -1251
rect 275 -1386 276 -1328
rect 373 -1386 374 -1328
rect 677 -1386 678 -1328
rect 765 -1386 766 -1328
rect 835 -1329 836 -1251
rect 859 -1386 860 -1328
rect 1703 -1386 1704 -1328
rect 198 -1331 199 -1251
rect 212 -1386 213 -1330
rect 436 -1331 437 -1251
rect 450 -1386 451 -1330
rect 464 -1331 465 -1251
rect 646 -1386 647 -1330
rect 905 -1331 906 -1251
rect 982 -1386 983 -1330
rect 996 -1386 997 -1330
rect 1899 -1331 1900 -1251
rect 198 -1386 199 -1332
rect 639 -1333 640 -1251
rect 884 -1333 885 -1251
rect 905 -1386 906 -1332
rect 1164 -1386 1165 -1332
rect 1213 -1333 1214 -1251
rect 1227 -1333 1228 -1251
rect 1395 -1386 1396 -1332
rect 1864 -1333 1865 -1251
rect 1899 -1386 1900 -1332
rect 436 -1386 437 -1334
rect 758 -1335 759 -1251
rect 884 -1386 885 -1334
rect 919 -1335 920 -1251
rect 1059 -1335 1060 -1251
rect 1213 -1386 1214 -1334
rect 1227 -1386 1228 -1334
rect 1248 -1335 1249 -1251
rect 1318 -1335 1319 -1251
rect 1339 -1386 1340 -1334
rect 1815 -1335 1816 -1251
rect 1864 -1386 1865 -1334
rect 464 -1386 465 -1336
rect 716 -1337 717 -1251
rect 751 -1337 752 -1251
rect 758 -1386 759 -1336
rect 1052 -1337 1053 -1251
rect 1059 -1386 1060 -1336
rect 1248 -1386 1249 -1336
rect 1346 -1337 1347 -1251
rect 1794 -1337 1795 -1251
rect 1815 -1386 1816 -1336
rect 471 -1386 472 -1338
rect 1003 -1339 1004 -1251
rect 1318 -1386 1319 -1338
rect 1402 -1339 1403 -1251
rect 1647 -1339 1648 -1251
rect 1794 -1386 1795 -1338
rect 474 -1341 475 -1251
rect 625 -1341 626 -1251
rect 639 -1386 640 -1340
rect 674 -1341 675 -1251
rect 716 -1386 717 -1340
rect 737 -1341 738 -1251
rect 744 -1341 745 -1251
rect 751 -1386 752 -1340
rect 1003 -1386 1004 -1340
rect 1181 -1341 1182 -1251
rect 1346 -1386 1347 -1340
rect 1353 -1341 1354 -1251
rect 1647 -1386 1648 -1340
rect 1738 -1341 1739 -1251
rect 114 -1343 115 -1251
rect 674 -1386 675 -1342
rect 737 -1386 738 -1342
rect 1010 -1343 1011 -1251
rect 1052 -1386 1053 -1342
rect 1402 -1386 1403 -1342
rect 1717 -1343 1718 -1251
rect 1738 -1386 1739 -1342
rect 114 -1386 115 -1344
rect 345 -1345 346 -1251
rect 478 -1345 479 -1251
rect 520 -1386 521 -1344
rect 569 -1386 570 -1344
rect 709 -1345 710 -1251
rect 943 -1386 944 -1344
rect 1717 -1386 1718 -1344
rect 159 -1347 160 -1251
rect 345 -1386 346 -1346
rect 478 -1386 479 -1346
rect 499 -1347 500 -1251
rect 590 -1347 591 -1251
rect 835 -1386 836 -1346
rect 1353 -1386 1354 -1346
rect 1367 -1347 1368 -1251
rect 173 -1349 174 -1251
rect 1010 -1386 1011 -1348
rect 1367 -1386 1368 -1348
rect 1381 -1349 1382 -1251
rect 485 -1351 486 -1251
rect 583 -1351 584 -1251
rect 625 -1386 626 -1350
rect 695 -1351 696 -1251
rect 709 -1386 710 -1350
rect 786 -1386 787 -1350
rect 1241 -1351 1242 -1251
rect 1381 -1386 1382 -1350
rect 219 -1353 220 -1251
rect 695 -1386 696 -1352
rect 1241 -1386 1242 -1352
rect 1640 -1353 1641 -1251
rect 191 -1355 192 -1251
rect 219 -1386 220 -1354
rect 432 -1386 433 -1354
rect 583 -1386 584 -1354
rect 1556 -1355 1557 -1251
rect 1640 -1386 1641 -1354
rect 191 -1386 192 -1356
rect 565 -1357 566 -1251
rect 1535 -1357 1536 -1251
rect 1556 -1386 1557 -1356
rect 485 -1386 486 -1358
rect 702 -1359 703 -1251
rect 1528 -1359 1529 -1251
rect 1535 -1386 1536 -1358
rect 429 -1361 430 -1251
rect 702 -1386 703 -1360
rect 1514 -1361 1515 -1251
rect 1528 -1386 1529 -1360
rect 429 -1386 430 -1362
rect 1619 -1363 1620 -1251
rect 492 -1386 493 -1364
rect 506 -1365 507 -1251
rect 527 -1365 528 -1251
rect 590 -1386 591 -1364
rect 1500 -1365 1501 -1251
rect 1514 -1386 1515 -1364
rect 1570 -1365 1571 -1251
rect 1619 -1386 1620 -1364
rect 499 -1386 500 -1366
rect 933 -1367 934 -1251
rect 1500 -1386 1501 -1366
rect 1633 -1367 1634 -1251
rect 506 -1386 507 -1368
rect 632 -1369 633 -1251
rect 933 -1386 934 -1368
rect 999 -1386 1000 -1368
rect 1549 -1369 1550 -1251
rect 1570 -1386 1571 -1368
rect 1577 -1369 1578 -1251
rect 1633 -1386 1634 -1368
rect 527 -1386 528 -1370
rect 1283 -1371 1284 -1251
rect 1549 -1386 1550 -1370
rect 1731 -1371 1732 -1251
rect 632 -1386 633 -1372
rect 828 -1373 829 -1251
rect 919 -1386 920 -1372
rect 1577 -1386 1578 -1372
rect 1724 -1373 1725 -1251
rect 1731 -1386 1732 -1372
rect 744 -1386 745 -1374
rect 1283 -1386 1284 -1374
rect 1710 -1375 1711 -1251
rect 1724 -1386 1725 -1374
rect 828 -1386 829 -1376
rect 863 -1377 864 -1251
rect 1584 -1377 1585 -1251
rect 1710 -1386 1711 -1376
rect 653 -1386 654 -1378
rect 863 -1386 864 -1378
rect 1199 -1379 1200 -1251
rect 1584 -1386 1585 -1378
rect 1192 -1381 1193 -1251
rect 1199 -1386 1200 -1380
rect 1192 -1386 1193 -1382
rect 1206 -1383 1207 -1251
rect 180 -1385 181 -1251
rect 1206 -1386 1207 -1384
rect 2 -1517 3 -1395
rect 208 -1396 209 -1394
rect 485 -1396 486 -1394
rect 919 -1396 920 -1394
rect 940 -1396 941 -1394
rect 1647 -1396 1648 -1394
rect 1766 -1396 1767 -1394
rect 1766 -1517 1767 -1395
rect 1766 -1396 1767 -1394
rect 1766 -1517 1767 -1395
rect 1892 -1396 1893 -1394
rect 1892 -1517 1893 -1395
rect 1892 -1396 1893 -1394
rect 1892 -1517 1893 -1395
rect 1899 -1396 1900 -1394
rect 1962 -1517 1963 -1395
rect 1969 -1396 1970 -1394
rect 1969 -1517 1970 -1395
rect 1969 -1396 1970 -1394
rect 1969 -1517 1970 -1395
rect 1976 -1396 1977 -1394
rect 2025 -1517 2026 -1395
rect 9 -1398 10 -1394
rect 215 -1517 216 -1397
rect 485 -1517 486 -1397
rect 492 -1398 493 -1394
rect 527 -1398 528 -1394
rect 646 -1398 647 -1394
rect 674 -1517 675 -1397
rect 681 -1398 682 -1394
rect 712 -1398 713 -1394
rect 912 -1398 913 -1394
rect 947 -1398 948 -1394
rect 999 -1398 1000 -1394
rect 1003 -1398 1004 -1394
rect 1013 -1444 1014 -1397
rect 1038 -1398 1039 -1394
rect 1073 -1517 1074 -1397
rect 1104 -1517 1105 -1397
rect 1542 -1398 1543 -1394
rect 1647 -1517 1648 -1397
rect 1822 -1398 1823 -1394
rect 1913 -1398 1914 -1394
rect 1927 -1398 1928 -1394
rect 1941 -1398 1942 -1394
rect 2011 -1517 2012 -1397
rect 9 -1517 10 -1399
rect 261 -1400 262 -1394
rect 527 -1517 528 -1399
rect 922 -1400 923 -1394
rect 926 -1400 927 -1394
rect 1038 -1517 1039 -1399
rect 1052 -1400 1053 -1394
rect 1808 -1400 1809 -1394
rect 1822 -1517 1823 -1399
rect 1920 -1400 1921 -1394
rect 1948 -1400 1949 -1394
rect 1955 -1517 1956 -1399
rect 1983 -1400 1984 -1394
rect 1986 -1400 1987 -1394
rect 1997 -1400 1998 -1394
rect 2018 -1517 2019 -1399
rect 16 -1402 17 -1394
rect 152 -1402 153 -1394
rect 184 -1402 185 -1394
rect 1185 -1402 1186 -1394
rect 1241 -1402 1242 -1394
rect 1794 -1402 1795 -1394
rect 1843 -1402 1844 -1394
rect 1948 -1517 1949 -1401
rect 1983 -1517 1984 -1401
rect 1990 -1402 1991 -1394
rect 16 -1517 17 -1403
rect 121 -1404 122 -1394
rect 142 -1517 143 -1403
rect 1682 -1404 1683 -1394
rect 1780 -1404 1781 -1394
rect 1843 -1517 1844 -1403
rect 1864 -1404 1865 -1394
rect 1927 -1517 1928 -1403
rect 23 -1406 24 -1394
rect 23 -1517 24 -1405
rect 23 -1406 24 -1394
rect 23 -1517 24 -1405
rect 30 -1406 31 -1394
rect 957 -1517 958 -1405
rect 968 -1406 969 -1394
rect 1444 -1406 1445 -1394
rect 1577 -1406 1578 -1394
rect 1808 -1517 1809 -1405
rect 1864 -1517 1865 -1405
rect 1878 -1406 1879 -1394
rect 1916 -1406 1917 -1394
rect 1934 -1406 1935 -1394
rect 30 -1517 31 -1407
rect 618 -1408 619 -1394
rect 632 -1408 633 -1394
rect 667 -1408 668 -1394
rect 677 -1408 678 -1394
rect 961 -1408 962 -1394
rect 975 -1408 976 -1394
rect 1052 -1517 1053 -1407
rect 1055 -1408 1056 -1394
rect 1381 -1408 1382 -1394
rect 1444 -1517 1445 -1407
rect 1591 -1408 1592 -1394
rect 1605 -1408 1606 -1394
rect 1682 -1517 1683 -1407
rect 1738 -1408 1739 -1394
rect 1780 -1517 1781 -1407
rect 1787 -1408 1788 -1394
rect 1878 -1517 1879 -1407
rect 1885 -1408 1886 -1394
rect 1934 -1517 1935 -1407
rect 47 -1517 48 -1409
rect 1542 -1517 1543 -1409
rect 1556 -1410 1557 -1394
rect 1605 -1517 1606 -1409
rect 1661 -1410 1662 -1394
rect 1738 -1517 1739 -1409
rect 1794 -1517 1795 -1409
rect 1857 -1410 1858 -1394
rect 51 -1412 52 -1394
rect 1899 -1517 1900 -1411
rect 51 -1517 52 -1413
rect 100 -1414 101 -1394
rect 107 -1517 108 -1413
rect 233 -1414 234 -1394
rect 450 -1414 451 -1394
rect 632 -1517 633 -1413
rect 814 -1414 815 -1394
rect 968 -1517 969 -1413
rect 975 -1517 976 -1413
rect 1307 -1517 1308 -1413
rect 1335 -1517 1336 -1413
rect 1906 -1414 1907 -1394
rect 58 -1416 59 -1394
rect 499 -1416 500 -1394
rect 548 -1416 549 -1394
rect 681 -1517 682 -1415
rect 814 -1517 815 -1415
rect 828 -1416 829 -1394
rect 849 -1416 850 -1394
rect 940 -1517 941 -1415
rect 947 -1517 948 -1415
rect 1360 -1416 1361 -1394
rect 1437 -1416 1438 -1394
rect 1591 -1517 1592 -1415
rect 1801 -1416 1802 -1394
rect 1906 -1517 1907 -1415
rect 58 -1517 59 -1417
rect 247 -1418 248 -1394
rect 408 -1418 409 -1394
rect 548 -1517 549 -1417
rect 562 -1418 563 -1394
rect 709 -1418 710 -1394
rect 744 -1418 745 -1394
rect 828 -1517 829 -1417
rect 877 -1418 878 -1394
rect 877 -1517 878 -1417
rect 877 -1418 878 -1394
rect 877 -1517 878 -1417
rect 905 -1418 906 -1394
rect 912 -1517 913 -1417
rect 922 -1517 923 -1417
rect 1941 -1517 1942 -1417
rect 65 -1420 66 -1394
rect 72 -1517 73 -1419
rect 79 -1420 80 -1394
rect 261 -1517 262 -1419
rect 408 -1517 409 -1419
rect 506 -1420 507 -1394
rect 562 -1517 563 -1419
rect 709 -1517 710 -1419
rect 744 -1517 745 -1419
rect 835 -1420 836 -1394
rect 842 -1420 843 -1394
rect 905 -1517 906 -1419
rect 926 -1517 927 -1419
rect 933 -1420 934 -1394
rect 961 -1517 962 -1419
rect 1178 -1420 1179 -1394
rect 1185 -1517 1186 -1419
rect 1262 -1420 1263 -1394
rect 1283 -1420 1284 -1394
rect 1836 -1420 1837 -1394
rect 1850 -1420 1851 -1394
rect 1857 -1517 1858 -1419
rect 79 -1517 80 -1421
rect 835 -1517 836 -1421
rect 884 -1422 885 -1394
rect 933 -1517 934 -1421
rect 985 -1517 986 -1421
rect 1409 -1422 1410 -1394
rect 1521 -1422 1522 -1394
rect 1556 -1517 1557 -1421
rect 1577 -1517 1578 -1421
rect 1654 -1422 1655 -1394
rect 1703 -1422 1704 -1394
rect 1801 -1517 1802 -1421
rect 82 -1517 83 -1423
rect 1136 -1424 1137 -1394
rect 1164 -1424 1165 -1394
rect 1241 -1517 1242 -1423
rect 1283 -1517 1284 -1423
rect 1325 -1424 1326 -1394
rect 1346 -1424 1347 -1394
rect 1360 -1517 1361 -1423
rect 1374 -1424 1375 -1394
rect 1409 -1517 1410 -1423
rect 1507 -1424 1508 -1394
rect 1521 -1517 1522 -1423
rect 1535 -1424 1536 -1394
rect 1661 -1517 1662 -1423
rect 1703 -1517 1704 -1423
rect 1773 -1424 1774 -1394
rect 86 -1426 87 -1394
rect 184 -1517 185 -1425
rect 194 -1517 195 -1425
rect 695 -1426 696 -1394
rect 751 -1426 752 -1394
rect 842 -1517 843 -1425
rect 982 -1426 983 -1394
rect 1136 -1517 1137 -1425
rect 1150 -1426 1151 -1394
rect 1164 -1517 1165 -1425
rect 1171 -1426 1172 -1394
rect 1451 -1426 1452 -1394
rect 1479 -1426 1480 -1394
rect 1507 -1517 1508 -1425
rect 1549 -1426 1550 -1394
rect 1850 -1517 1851 -1425
rect 93 -1428 94 -1394
rect 100 -1517 101 -1427
rect 114 -1428 115 -1394
rect 432 -1428 433 -1394
rect 450 -1517 451 -1427
rect 579 -1428 580 -1394
rect 583 -1428 584 -1394
rect 695 -1517 696 -1427
rect 786 -1428 787 -1394
rect 849 -1517 850 -1427
rect 982 -1517 983 -1427
rect 1640 -1428 1641 -1394
rect 1717 -1428 1718 -1394
rect 1773 -1517 1774 -1427
rect 93 -1517 94 -1429
rect 149 -1430 150 -1394
rect 198 -1430 199 -1394
rect 243 -1517 244 -1429
rect 247 -1517 248 -1429
rect 950 -1517 951 -1429
rect 996 -1430 997 -1394
rect 1381 -1517 1382 -1429
rect 1388 -1430 1389 -1394
rect 1451 -1517 1452 -1429
rect 1549 -1517 1550 -1429
rect 1626 -1430 1627 -1394
rect 1640 -1517 1641 -1429
rect 1997 -1517 1998 -1429
rect 114 -1517 115 -1431
rect 436 -1432 437 -1394
rect 492 -1517 493 -1431
rect 667 -1517 668 -1431
rect 807 -1432 808 -1394
rect 1171 -1517 1172 -1431
rect 1178 -1517 1179 -1431
rect 1395 -1432 1396 -1394
rect 1759 -1432 1760 -1394
rect 1836 -1517 1837 -1431
rect 121 -1517 122 -1433
rect 131 -1434 132 -1394
rect 145 -1434 146 -1394
rect 1913 -1517 1914 -1433
rect 145 -1517 146 -1435
rect 1206 -1436 1207 -1394
rect 1248 -1436 1249 -1394
rect 1325 -1517 1326 -1435
rect 1346 -1517 1347 -1435
rect 1472 -1436 1473 -1394
rect 1752 -1436 1753 -1394
rect 1759 -1517 1760 -1435
rect 149 -1517 150 -1437
rect 1108 -1438 1109 -1394
rect 1111 -1438 1112 -1394
rect 1612 -1438 1613 -1394
rect 198 -1517 199 -1439
rect 282 -1440 283 -1394
rect 310 -1440 311 -1394
rect 786 -1517 787 -1439
rect 793 -1440 794 -1394
rect 807 -1517 808 -1439
rect 929 -1440 930 -1394
rect 1472 -1517 1473 -1439
rect 1493 -1440 1494 -1394
rect 1752 -1517 1753 -1439
rect 37 -1442 38 -1394
rect 282 -1517 283 -1441
rect 303 -1442 304 -1394
rect 310 -1517 311 -1441
rect 373 -1442 374 -1394
rect 436 -1517 437 -1441
rect 506 -1517 507 -1441
rect 513 -1442 514 -1394
rect 569 -1442 570 -1394
rect 943 -1442 944 -1394
rect 954 -1442 955 -1394
rect 996 -1517 997 -1441
rect 1003 -1517 1004 -1441
rect 1066 -1442 1067 -1394
rect 1710 -1442 1711 -1394
rect 37 -1517 38 -1443
rect 75 -1444 76 -1394
rect 86 -1517 87 -1443
rect 954 -1517 955 -1443
rect 1006 -1517 1007 -1443
rect 1199 -1444 1200 -1394
rect 1248 -1517 1249 -1443
rect 1290 -1444 1291 -1394
rect 1367 -1444 1368 -1394
rect 1395 -1517 1396 -1443
rect 1493 -1517 1494 -1443
rect 1570 -1444 1571 -1394
rect 1633 -1444 1634 -1394
rect 1710 -1517 1711 -1443
rect 1986 -1517 1987 -1443
rect 1990 -1517 1991 -1443
rect 110 -1446 111 -1394
rect 303 -1517 304 -1445
rect 338 -1446 339 -1394
rect 373 -1517 374 -1445
rect 387 -1446 388 -1394
rect 1206 -1517 1207 -1445
rect 1255 -1446 1256 -1394
rect 1388 -1517 1389 -1445
rect 1528 -1446 1529 -1394
rect 1570 -1517 1571 -1445
rect 128 -1448 129 -1394
rect 1633 -1517 1634 -1447
rect 128 -1517 129 -1449
rect 135 -1450 136 -1394
rect 205 -1517 206 -1449
rect 226 -1450 227 -1394
rect 233 -1517 234 -1449
rect 1304 -1450 1305 -1394
rect 1367 -1517 1368 -1449
rect 1423 -1450 1424 -1394
rect 1486 -1450 1487 -1394
rect 1528 -1517 1529 -1449
rect 1563 -1450 1564 -1394
rect 1612 -1517 1613 -1449
rect 135 -1517 136 -1451
rect 177 -1452 178 -1394
rect 226 -1517 227 -1451
rect 331 -1452 332 -1394
rect 338 -1517 339 -1451
rect 520 -1452 521 -1394
rect 555 -1452 556 -1394
rect 569 -1517 570 -1451
rect 576 -1452 577 -1394
rect 859 -1452 860 -1394
rect 1010 -1452 1011 -1394
rect 1717 -1517 1718 -1451
rect 296 -1454 297 -1394
rect 331 -1517 332 -1453
rect 387 -1517 388 -1453
rect 394 -1454 395 -1394
rect 422 -1454 423 -1394
rect 583 -1517 584 -1453
rect 590 -1454 591 -1394
rect 646 -1517 647 -1453
rect 663 -1517 664 -1453
rect 1437 -1517 1438 -1453
rect 163 -1456 164 -1394
rect 394 -1517 395 -1455
rect 415 -1456 416 -1394
rect 422 -1517 423 -1455
rect 513 -1517 514 -1455
rect 611 -1456 612 -1394
rect 618 -1517 619 -1455
rect 628 -1456 629 -1394
rect 793 -1517 794 -1455
rect 800 -1456 801 -1394
rect 898 -1456 899 -1394
rect 1010 -1517 1011 -1455
rect 1024 -1456 1025 -1394
rect 1885 -1517 1886 -1455
rect 163 -1517 164 -1457
rect 254 -1458 255 -1394
rect 415 -1517 416 -1457
rect 457 -1458 458 -1394
rect 478 -1458 479 -1394
rect 800 -1517 801 -1457
rect 821 -1458 822 -1394
rect 898 -1517 899 -1457
rect 1031 -1458 1032 -1394
rect 1626 -1517 1627 -1457
rect 212 -1460 213 -1394
rect 457 -1517 458 -1459
rect 520 -1517 521 -1459
rect 688 -1460 689 -1394
rect 702 -1460 703 -1394
rect 821 -1517 822 -1459
rect 989 -1460 990 -1394
rect 1031 -1517 1032 -1459
rect 1034 -1460 1035 -1394
rect 1654 -1517 1655 -1459
rect 177 -1517 178 -1461
rect 212 -1517 213 -1461
rect 219 -1462 220 -1394
rect 296 -1517 297 -1461
rect 443 -1462 444 -1394
rect 478 -1517 479 -1461
rect 534 -1462 535 -1394
rect 702 -1517 703 -1461
rect 751 -1517 752 -1461
rect 1024 -1517 1025 -1461
rect 1087 -1462 1088 -1394
rect 1535 -1517 1536 -1461
rect 191 -1464 192 -1394
rect 534 -1517 535 -1463
rect 555 -1517 556 -1463
rect 2007 -1517 2008 -1463
rect 191 -1517 192 -1465
rect 772 -1466 773 -1394
rect 989 -1517 990 -1465
rect 1017 -1466 1018 -1394
rect 1087 -1517 1088 -1465
rect 1094 -1466 1095 -1394
rect 1108 -1517 1109 -1465
rect 1479 -1517 1480 -1465
rect 219 -1517 220 -1467
rect 289 -1468 290 -1394
rect 359 -1468 360 -1394
rect 443 -1517 444 -1467
rect 576 -1517 577 -1467
rect 779 -1468 780 -1394
rect 863 -1468 864 -1394
rect 1017 -1517 1018 -1467
rect 1080 -1468 1081 -1394
rect 1094 -1517 1095 -1467
rect 1111 -1517 1112 -1467
rect 1290 -1517 1291 -1467
rect 1304 -1517 1305 -1467
rect 1829 -1468 1830 -1394
rect 254 -1517 255 -1469
rect 268 -1470 269 -1394
rect 275 -1470 276 -1394
rect 289 -1517 290 -1469
rect 324 -1470 325 -1394
rect 359 -1517 360 -1469
rect 590 -1517 591 -1469
rect 856 -1470 857 -1394
rect 1080 -1517 1081 -1469
rect 1265 -1517 1266 -1469
rect 1286 -1470 1287 -1394
rect 1339 -1470 1340 -1394
rect 1402 -1470 1403 -1394
rect 1423 -1517 1424 -1469
rect 1731 -1470 1732 -1394
rect 1829 -1517 1830 -1469
rect 240 -1472 241 -1394
rect 268 -1517 269 -1471
rect 275 -1517 276 -1471
rect 352 -1472 353 -1394
rect 597 -1472 598 -1394
rect 656 -1472 657 -1394
rect 670 -1517 671 -1471
rect 1402 -1517 1403 -1471
rect 1724 -1472 1725 -1394
rect 1731 -1517 1732 -1471
rect 324 -1517 325 -1473
rect 401 -1474 402 -1394
rect 464 -1474 465 -1394
rect 597 -1517 598 -1473
rect 604 -1474 605 -1394
rect 884 -1517 885 -1473
rect 1115 -1474 1116 -1394
rect 1262 -1517 1263 -1473
rect 1339 -1517 1340 -1473
rect 1458 -1474 1459 -1394
rect 1696 -1474 1697 -1394
rect 1724 -1517 1725 -1473
rect 352 -1517 353 -1475
rect 639 -1476 640 -1394
rect 653 -1476 654 -1394
rect 863 -1517 864 -1475
rect 1118 -1517 1119 -1475
rect 1745 -1476 1746 -1394
rect 401 -1517 402 -1477
rect 502 -1517 503 -1477
rect 541 -1478 542 -1394
rect 639 -1517 640 -1477
rect 653 -1517 654 -1477
rect 1132 -1517 1133 -1477
rect 1143 -1478 1144 -1394
rect 1150 -1517 1151 -1477
rect 1160 -1517 1161 -1477
rect 1486 -1517 1487 -1477
rect 1675 -1478 1676 -1394
rect 1745 -1517 1746 -1477
rect 44 -1480 45 -1394
rect 541 -1517 542 -1479
rect 604 -1517 605 -1479
rect 712 -1517 713 -1479
rect 758 -1480 759 -1394
rect 772 -1517 773 -1479
rect 779 -1517 780 -1479
rect 891 -1480 892 -1394
rect 1059 -1480 1060 -1394
rect 1143 -1517 1144 -1479
rect 1199 -1517 1200 -1479
rect 1213 -1480 1214 -1394
rect 1220 -1480 1221 -1394
rect 1255 -1517 1256 -1479
rect 1416 -1480 1417 -1394
rect 1458 -1517 1459 -1479
rect 1584 -1480 1585 -1394
rect 1675 -1517 1676 -1479
rect 44 -1517 45 -1481
rect 1920 -1517 1921 -1481
rect 170 -1484 171 -1394
rect 758 -1517 759 -1483
rect 856 -1517 857 -1483
rect 1115 -1517 1116 -1483
rect 1122 -1484 1123 -1394
rect 1563 -1517 1564 -1483
rect 61 -1486 62 -1394
rect 170 -1517 171 -1485
rect 464 -1517 465 -1485
rect 530 -1486 531 -1394
rect 611 -1517 612 -1485
rect 1076 -1486 1077 -1394
rect 1101 -1486 1102 -1394
rect 1122 -1517 1123 -1485
rect 1157 -1486 1158 -1394
rect 1213 -1517 1214 -1485
rect 1244 -1486 1245 -1394
rect 1696 -1517 1697 -1485
rect 61 -1517 62 -1487
rect 65 -1517 66 -1487
rect 628 -1517 629 -1487
rect 716 -1488 717 -1394
rect 870 -1488 871 -1394
rect 891 -1517 892 -1487
rect 1059 -1517 1060 -1487
rect 1129 -1488 1130 -1394
rect 1157 -1517 1158 -1487
rect 1871 -1488 1872 -1394
rect 471 -1490 472 -1394
rect 870 -1517 871 -1489
rect 1101 -1517 1102 -1489
rect 1311 -1490 1312 -1394
rect 1318 -1490 1319 -1394
rect 1416 -1517 1417 -1489
rect 1815 -1490 1816 -1394
rect 1871 -1517 1872 -1489
rect 366 -1492 367 -1394
rect 471 -1517 472 -1491
rect 688 -1517 689 -1491
rect 730 -1492 731 -1394
rect 1129 -1517 1130 -1491
rect 1374 -1517 1375 -1491
rect 1668 -1492 1669 -1394
rect 1815 -1517 1816 -1491
rect 366 -1517 367 -1493
rect 380 -1494 381 -1394
rect 716 -1517 717 -1493
rect 737 -1494 738 -1394
rect 1192 -1494 1193 -1394
rect 1220 -1517 1221 -1493
rect 1297 -1494 1298 -1394
rect 1318 -1517 1319 -1493
rect 1598 -1494 1599 -1394
rect 1668 -1517 1669 -1493
rect 380 -1517 381 -1495
rect 765 -1496 766 -1394
rect 1192 -1517 1193 -1495
rect 1787 -1517 1788 -1495
rect 660 -1498 661 -1394
rect 765 -1517 766 -1497
rect 1269 -1498 1270 -1394
rect 1297 -1517 1298 -1497
rect 1311 -1517 1312 -1497
rect 1514 -1498 1515 -1394
rect 1598 -1517 1599 -1497
rect 1689 -1498 1690 -1394
rect 156 -1500 157 -1394
rect 660 -1517 661 -1499
rect 723 -1500 724 -1394
rect 737 -1517 738 -1499
rect 1269 -1517 1270 -1499
rect 1276 -1500 1277 -1394
rect 1619 -1500 1620 -1394
rect 1689 -1517 1690 -1499
rect 156 -1517 157 -1501
rect 429 -1502 430 -1394
rect 730 -1517 731 -1501
rect 754 -1517 755 -1501
rect 1069 -1502 1070 -1394
rect 1619 -1517 1620 -1501
rect 240 -1517 241 -1503
rect 723 -1517 724 -1503
rect 1069 -1517 1070 -1503
rect 1500 -1504 1501 -1394
rect 317 -1506 318 -1394
rect 429 -1517 430 -1505
rect 1234 -1506 1235 -1394
rect 1276 -1517 1277 -1505
rect 1465 -1506 1466 -1394
rect 1500 -1517 1501 -1505
rect 317 -1517 318 -1507
rect 345 -1508 346 -1394
rect 1227 -1508 1228 -1394
rect 1234 -1517 1235 -1507
rect 1430 -1508 1431 -1394
rect 1465 -1517 1466 -1507
rect 166 -1510 167 -1394
rect 345 -1517 346 -1509
rect 625 -1510 626 -1394
rect 1227 -1517 1228 -1509
rect 1353 -1510 1354 -1394
rect 1430 -1517 1431 -1509
rect 625 -1517 626 -1511
rect 1584 -1517 1585 -1511
rect 1332 -1514 1333 -1394
rect 1353 -1517 1354 -1513
rect 1332 -1517 1333 -1515
rect 1514 -1517 1515 -1515
rect 2 -1527 3 -1525
rect 47 -1527 48 -1525
rect 58 -1527 59 -1525
rect 1724 -1527 1725 -1525
rect 1780 -1527 1781 -1525
rect 1780 -1644 1781 -1526
rect 1780 -1527 1781 -1525
rect 1780 -1644 1781 -1526
rect 1808 -1527 1809 -1525
rect 1811 -1541 1812 -1526
rect 1948 -1527 1949 -1525
rect 1969 -1527 1970 -1525
rect 1979 -1527 1980 -1525
rect 1990 -1527 1991 -1525
rect 2018 -1527 2019 -1525
rect 2018 -1644 2019 -1526
rect 2018 -1527 2019 -1525
rect 2018 -1644 2019 -1526
rect 2 -1644 3 -1528
rect 177 -1529 178 -1525
rect 180 -1644 181 -1528
rect 254 -1529 255 -1525
rect 338 -1529 339 -1525
rect 751 -1529 752 -1525
rect 754 -1529 755 -1525
rect 1661 -1529 1662 -1525
rect 1689 -1529 1690 -1525
rect 1724 -1644 1725 -1528
rect 1766 -1529 1767 -1525
rect 1948 -1644 1949 -1528
rect 1955 -1529 1956 -1525
rect 1972 -1529 1973 -1525
rect 1983 -1529 1984 -1525
rect 2000 -1529 2001 -1525
rect 23 -1531 24 -1525
rect 68 -1644 69 -1530
rect 72 -1531 73 -1525
rect 72 -1644 73 -1530
rect 72 -1531 73 -1525
rect 72 -1644 73 -1530
rect 82 -1531 83 -1525
rect 1104 -1531 1105 -1525
rect 1108 -1531 1109 -1525
rect 1829 -1531 1830 -1525
rect 23 -1644 24 -1532
rect 198 -1533 199 -1525
rect 233 -1533 234 -1525
rect 324 -1533 325 -1525
rect 338 -1644 339 -1532
rect 359 -1533 360 -1525
rect 485 -1533 486 -1525
rect 660 -1533 661 -1525
rect 663 -1533 664 -1525
rect 751 -1644 752 -1532
rect 768 -1644 769 -1532
rect 814 -1533 815 -1525
rect 884 -1533 885 -1525
rect 1160 -1533 1161 -1525
rect 1192 -1533 1193 -1525
rect 1234 -1533 1235 -1525
rect 1262 -1533 1263 -1525
rect 1346 -1533 1347 -1525
rect 1356 -1644 1357 -1532
rect 1731 -1533 1732 -1525
rect 1808 -1644 1809 -1532
rect 1878 -1533 1879 -1525
rect 30 -1535 31 -1525
rect 919 -1535 920 -1525
rect 954 -1535 955 -1525
rect 1850 -1535 1851 -1525
rect 30 -1644 31 -1536
rect 247 -1537 248 -1525
rect 254 -1644 255 -1536
rect 1055 -1644 1056 -1536
rect 1101 -1537 1102 -1525
rect 1339 -1537 1340 -1525
rect 1346 -1644 1347 -1536
rect 1360 -1537 1361 -1525
rect 1437 -1537 1438 -1525
rect 1437 -1644 1438 -1536
rect 1437 -1537 1438 -1525
rect 1437 -1644 1438 -1536
rect 1503 -1644 1504 -1536
rect 1836 -1537 1837 -1525
rect 37 -1539 38 -1525
rect 499 -1539 500 -1525
rect 502 -1539 503 -1525
rect 1038 -1539 1039 -1525
rect 1108 -1644 1109 -1538
rect 1335 -1539 1336 -1525
rect 1339 -1644 1340 -1538
rect 1353 -1539 1354 -1525
rect 1360 -1644 1361 -1538
rect 1381 -1539 1382 -1525
rect 1514 -1539 1515 -1525
rect 1514 -1644 1515 -1538
rect 1514 -1539 1515 -1525
rect 1514 -1644 1515 -1538
rect 1591 -1539 1592 -1525
rect 2004 -1539 2005 -1525
rect 37 -1644 38 -1540
rect 51 -1541 52 -1525
rect 58 -1644 59 -1540
rect 107 -1541 108 -1525
rect 117 -1644 118 -1540
rect 121 -1541 122 -1525
rect 135 -1541 136 -1525
rect 135 -1644 136 -1540
rect 135 -1541 136 -1525
rect 135 -1644 136 -1540
rect 142 -1541 143 -1525
rect 303 -1541 304 -1525
rect 324 -1644 325 -1540
rect 443 -1541 444 -1525
rect 499 -1644 500 -1540
rect 555 -1541 556 -1525
rect 593 -1541 594 -1525
rect 688 -1541 689 -1525
rect 709 -1541 710 -1525
rect 877 -1541 878 -1525
rect 905 -1541 906 -1525
rect 947 -1644 948 -1540
rect 957 -1541 958 -1525
rect 1689 -1644 1690 -1540
rect 1703 -1541 1704 -1525
rect 1766 -1644 1767 -1540
rect 1878 -1644 1879 -1540
rect 9 -1543 10 -1525
rect 51 -1644 52 -1542
rect 86 -1543 87 -1525
rect 107 -1644 108 -1542
rect 121 -1644 122 -1542
rect 184 -1543 185 -1525
rect 194 -1543 195 -1525
rect 1206 -1543 1207 -1525
rect 1234 -1644 1235 -1542
rect 1255 -1543 1256 -1525
rect 1262 -1644 1263 -1542
rect 1286 -1644 1287 -1542
rect 1325 -1543 1326 -1525
rect 1325 -1644 1326 -1542
rect 1325 -1543 1326 -1525
rect 1325 -1644 1326 -1542
rect 1353 -1644 1354 -1542
rect 1528 -1543 1529 -1525
rect 1577 -1543 1578 -1525
rect 1703 -1644 1704 -1542
rect 1717 -1543 1718 -1525
rect 1850 -1644 1851 -1542
rect 9 -1644 10 -1544
rect 156 -1545 157 -1525
rect 184 -1644 185 -1544
rect 544 -1644 545 -1544
rect 548 -1545 549 -1525
rect 548 -1644 549 -1544
rect 548 -1545 549 -1525
rect 548 -1644 549 -1544
rect 555 -1644 556 -1544
rect 702 -1545 703 -1525
rect 712 -1545 713 -1525
rect 1542 -1545 1543 -1525
rect 1577 -1644 1578 -1544
rect 1612 -1545 1613 -1525
rect 1661 -1644 1662 -1544
rect 1976 -1545 1977 -1525
rect 44 -1547 45 -1525
rect 100 -1547 101 -1525
rect 142 -1644 143 -1546
rect 628 -1547 629 -1525
rect 667 -1547 668 -1525
rect 1171 -1547 1172 -1525
rect 1199 -1547 1200 -1525
rect 1255 -1644 1256 -1546
rect 1265 -1547 1266 -1525
rect 1962 -1547 1963 -1525
rect 1976 -1644 1977 -1546
rect 2025 -1547 2026 -1525
rect 16 -1549 17 -1525
rect 44 -1644 45 -1548
rect 79 -1549 80 -1525
rect 100 -1644 101 -1548
rect 114 -1549 115 -1525
rect 667 -1644 668 -1548
rect 674 -1549 675 -1525
rect 1038 -1644 1039 -1548
rect 1111 -1549 1112 -1525
rect 1822 -1549 1823 -1525
rect 1829 -1644 1830 -1548
rect 1885 -1549 1886 -1525
rect 16 -1644 17 -1550
rect 89 -1644 90 -1550
rect 145 -1551 146 -1525
rect 198 -1644 199 -1550
rect 226 -1551 227 -1525
rect 247 -1644 248 -1550
rect 289 -1551 290 -1525
rect 485 -1644 486 -1550
rect 506 -1551 507 -1525
rect 506 -1644 507 -1550
rect 506 -1551 507 -1525
rect 506 -1644 507 -1550
rect 618 -1551 619 -1525
rect 1101 -1644 1102 -1550
rect 1118 -1551 1119 -1525
rect 1185 -1551 1186 -1525
rect 1199 -1644 1200 -1550
rect 1213 -1551 1214 -1525
rect 1269 -1551 1270 -1525
rect 1269 -1644 1270 -1550
rect 1269 -1551 1270 -1525
rect 1269 -1644 1270 -1550
rect 1374 -1551 1375 -1525
rect 1381 -1644 1382 -1550
rect 1493 -1551 1494 -1525
rect 1591 -1644 1592 -1550
rect 1612 -1644 1613 -1550
rect 1619 -1551 1620 -1525
rect 1731 -1644 1732 -1550
rect 1752 -1551 1753 -1525
rect 1794 -1551 1795 -1525
rect 1885 -1644 1886 -1550
rect 86 -1644 87 -1552
rect 698 -1644 699 -1552
rect 702 -1644 703 -1552
rect 821 -1553 822 -1525
rect 835 -1553 836 -1525
rect 877 -1644 878 -1552
rect 961 -1644 962 -1552
rect 1332 -1553 1333 -1525
rect 1374 -1644 1375 -1552
rect 1395 -1553 1396 -1525
rect 1493 -1644 1494 -1552
rect 1668 -1553 1669 -1525
rect 1822 -1644 1823 -1552
rect 1906 -1553 1907 -1525
rect 128 -1555 129 -1525
rect 145 -1644 146 -1554
rect 156 -1644 157 -1554
rect 219 -1555 220 -1525
rect 226 -1644 227 -1554
rect 1115 -1555 1116 -1525
rect 1122 -1555 1123 -1525
rect 1122 -1644 1123 -1554
rect 1122 -1555 1123 -1525
rect 1122 -1644 1123 -1554
rect 1129 -1555 1130 -1525
rect 1881 -1644 1882 -1554
rect 1906 -1644 1907 -1554
rect 1934 -1555 1935 -1525
rect 93 -1557 94 -1525
rect 128 -1644 129 -1556
rect 191 -1557 192 -1525
rect 219 -1644 220 -1556
rect 233 -1644 234 -1556
rect 310 -1557 311 -1525
rect 345 -1557 346 -1525
rect 670 -1557 671 -1525
rect 681 -1557 682 -1525
rect 1304 -1644 1305 -1556
rect 1307 -1557 1308 -1525
rect 1752 -1644 1753 -1556
rect 1871 -1557 1872 -1525
rect 1934 -1644 1935 -1556
rect 65 -1559 66 -1525
rect 93 -1644 94 -1558
rect 163 -1559 164 -1525
rect 191 -1644 192 -1558
rect 205 -1559 206 -1525
rect 345 -1644 346 -1558
rect 415 -1559 416 -1525
rect 821 -1644 822 -1558
rect 849 -1559 850 -1525
rect 905 -1644 906 -1558
rect 971 -1644 972 -1558
rect 1283 -1559 1284 -1525
rect 1307 -1644 1308 -1558
rect 1857 -1559 1858 -1525
rect 1871 -1644 1872 -1558
rect 1920 -1559 1921 -1525
rect 163 -1644 164 -1560
rect 660 -1644 661 -1560
rect 663 -1644 664 -1560
rect 1794 -1644 1795 -1560
rect 205 -1644 206 -1562
rect 520 -1563 521 -1525
rect 646 -1563 647 -1525
rect 674 -1644 675 -1562
rect 681 -1644 682 -1562
rect 828 -1563 829 -1525
rect 863 -1563 864 -1525
rect 1717 -1644 1718 -1562
rect 268 -1565 269 -1525
rect 310 -1644 311 -1564
rect 397 -1644 398 -1564
rect 646 -1644 647 -1564
rect 670 -1644 671 -1564
rect 842 -1565 843 -1525
rect 996 -1565 997 -1525
rect 996 -1644 997 -1564
rect 996 -1565 997 -1525
rect 996 -1644 997 -1564
rect 1003 -1565 1004 -1525
rect 1801 -1565 1802 -1525
rect 268 -1644 269 -1566
rect 569 -1567 570 -1525
rect 583 -1567 584 -1525
rect 842 -1644 843 -1566
rect 968 -1567 969 -1525
rect 1003 -1644 1004 -1566
rect 1073 -1567 1074 -1525
rect 1115 -1644 1116 -1566
rect 1132 -1567 1133 -1525
rect 1311 -1567 1312 -1525
rect 1332 -1644 1333 -1566
rect 1864 -1567 1865 -1525
rect 282 -1569 283 -1525
rect 520 -1644 521 -1568
rect 569 -1644 570 -1568
rect 576 -1569 577 -1525
rect 583 -1644 584 -1568
rect 730 -1569 731 -1525
rect 800 -1569 801 -1525
rect 1129 -1644 1130 -1568
rect 1132 -1644 1133 -1568
rect 1549 -1569 1550 -1525
rect 1619 -1644 1620 -1568
rect 1633 -1569 1634 -1525
rect 1647 -1569 1648 -1525
rect 1857 -1644 1858 -1568
rect 1864 -1644 1865 -1568
rect 1913 -1569 1914 -1525
rect 282 -1644 283 -1570
rect 450 -1571 451 -1525
rect 457 -1571 458 -1525
rect 712 -1644 713 -1570
rect 723 -1571 724 -1525
rect 1209 -1644 1210 -1570
rect 1213 -1644 1214 -1570
rect 1444 -1571 1445 -1525
rect 1507 -1571 1508 -1525
rect 1633 -1644 1634 -1570
rect 1647 -1644 1648 -1570
rect 1654 -1571 1655 -1525
rect 1668 -1644 1669 -1570
rect 1696 -1571 1697 -1525
rect 1787 -1571 1788 -1525
rect 1801 -1644 1802 -1570
rect 1913 -1644 1914 -1570
rect 1941 -1571 1942 -1525
rect 261 -1573 262 -1525
rect 450 -1644 451 -1572
rect 464 -1573 465 -1525
rect 688 -1644 689 -1572
rect 723 -1644 724 -1572
rect 982 -1573 983 -1525
rect 1024 -1573 1025 -1525
rect 1073 -1644 1074 -1572
rect 1150 -1573 1151 -1525
rect 1192 -1644 1193 -1572
rect 1283 -1644 1284 -1572
rect 1626 -1573 1627 -1525
rect 1654 -1644 1655 -1572
rect 1682 -1573 1683 -1525
rect 1696 -1644 1697 -1572
rect 1843 -1573 1844 -1525
rect 1941 -1644 1942 -1572
rect 2011 -1573 2012 -1525
rect 261 -1644 262 -1574
rect 1069 -1575 1070 -1525
rect 1171 -1644 1172 -1574
rect 1241 -1575 1242 -1525
rect 1311 -1644 1312 -1574
rect 1318 -1575 1319 -1525
rect 1395 -1644 1396 -1574
rect 1402 -1575 1403 -1525
rect 1444 -1644 1445 -1574
rect 1465 -1575 1466 -1525
rect 1521 -1575 1522 -1525
rect 1528 -1644 1529 -1574
rect 1542 -1644 1543 -1574
rect 1563 -1575 1564 -1525
rect 1626 -1644 1627 -1574
rect 1710 -1575 1711 -1525
rect 1787 -1644 1788 -1574
rect 1927 -1575 1928 -1525
rect 65 -1644 66 -1576
rect 1710 -1644 1711 -1576
rect 1843 -1644 1844 -1576
rect 1920 -1644 1921 -1576
rect 289 -1644 290 -1578
rect 366 -1579 367 -1525
rect 418 -1644 419 -1578
rect 849 -1644 850 -1578
rect 919 -1644 920 -1578
rect 1507 -1644 1508 -1578
rect 1521 -1644 1522 -1578
rect 1605 -1579 1606 -1525
rect 296 -1581 297 -1525
rect 359 -1644 360 -1580
rect 366 -1644 367 -1580
rect 429 -1581 430 -1525
rect 443 -1644 444 -1580
rect 653 -1581 654 -1525
rect 730 -1644 731 -1580
rect 975 -1581 976 -1525
rect 1006 -1581 1007 -1525
rect 1682 -1644 1683 -1580
rect 114 -1644 115 -1582
rect 653 -1644 654 -1582
rect 772 -1583 773 -1525
rect 800 -1644 801 -1582
rect 807 -1583 808 -1525
rect 954 -1644 955 -1582
rect 968 -1644 969 -1582
rect 989 -1583 990 -1525
rect 1024 -1644 1025 -1582
rect 1136 -1583 1137 -1525
rect 1185 -1644 1186 -1582
rect 1248 -1583 1249 -1525
rect 1290 -1583 1291 -1525
rect 1465 -1644 1466 -1582
rect 1549 -1644 1550 -1582
rect 1556 -1583 1557 -1525
rect 1563 -1644 1564 -1582
rect 1584 -1583 1585 -1525
rect 1598 -1583 1599 -1525
rect 1927 -1644 1928 -1582
rect 296 -1644 297 -1584
rect 985 -1585 986 -1525
rect 989 -1644 990 -1584
rect 1090 -1644 1091 -1584
rect 1220 -1585 1221 -1525
rect 1248 -1644 1249 -1584
rect 1290 -1644 1291 -1584
rect 1297 -1585 1298 -1525
rect 1402 -1644 1403 -1584
rect 1416 -1585 1417 -1525
rect 1535 -1585 1536 -1525
rect 1584 -1644 1585 -1584
rect 1598 -1644 1599 -1584
rect 1640 -1585 1641 -1525
rect 303 -1644 304 -1586
rect 331 -1587 332 -1525
rect 422 -1587 423 -1525
rect 457 -1644 458 -1586
rect 478 -1587 479 -1525
rect 618 -1644 619 -1586
rect 765 -1587 766 -1525
rect 772 -1644 773 -1586
rect 793 -1587 794 -1525
rect 807 -1644 808 -1586
rect 817 -1644 818 -1586
rect 1836 -1644 1837 -1586
rect 212 -1589 213 -1525
rect 422 -1644 423 -1588
rect 429 -1644 430 -1588
rect 950 -1589 951 -1525
rect 1031 -1589 1032 -1525
rect 1150 -1644 1151 -1588
rect 1164 -1589 1165 -1525
rect 1297 -1644 1298 -1588
rect 1367 -1589 1368 -1525
rect 1535 -1644 1536 -1588
rect 1570 -1589 1571 -1525
rect 1605 -1644 1606 -1588
rect 170 -1591 171 -1525
rect 212 -1644 213 -1590
rect 317 -1591 318 -1525
rect 464 -1644 465 -1590
rect 478 -1644 479 -1590
rect 513 -1591 514 -1525
rect 597 -1591 598 -1525
rect 863 -1644 864 -1590
rect 922 -1591 923 -1525
rect 1640 -1644 1641 -1590
rect 317 -1644 318 -1592
rect 611 -1593 612 -1525
rect 793 -1644 794 -1592
rect 856 -1593 857 -1525
rect 884 -1644 885 -1592
rect 922 -1644 923 -1592
rect 926 -1593 927 -1525
rect 982 -1644 983 -1592
rect 1010 -1593 1011 -1525
rect 1031 -1644 1032 -1592
rect 1059 -1593 1060 -1525
rect 1318 -1644 1319 -1592
rect 1367 -1644 1368 -1592
rect 1388 -1593 1389 -1525
rect 1416 -1644 1417 -1592
rect 1423 -1593 1424 -1525
rect 79 -1644 80 -1594
rect 1010 -1644 1011 -1594
rect 1080 -1595 1081 -1525
rect 1164 -1644 1165 -1594
rect 1195 -1595 1196 -1525
rect 1570 -1644 1571 -1594
rect 331 -1644 332 -1596
rect 387 -1597 388 -1525
rect 513 -1644 514 -1596
rect 541 -1597 542 -1525
rect 611 -1644 612 -1596
rect 740 -1644 741 -1596
rect 828 -1644 829 -1596
rect 1136 -1644 1137 -1596
rect 1220 -1644 1221 -1596
rect 1276 -1597 1277 -1525
rect 1388 -1644 1389 -1596
rect 1451 -1597 1452 -1525
rect 387 -1644 388 -1598
rect 814 -1644 815 -1598
rect 856 -1644 857 -1598
rect 891 -1599 892 -1525
rect 912 -1599 913 -1525
rect 926 -1644 927 -1598
rect 933 -1599 934 -1525
rect 975 -1644 976 -1598
rect 1080 -1644 1081 -1598
rect 1227 -1599 1228 -1525
rect 1241 -1644 1242 -1598
rect 1815 -1599 1816 -1525
rect 177 -1644 178 -1600
rect 933 -1644 934 -1600
rect 940 -1601 941 -1525
rect 1059 -1644 1060 -1600
rect 1227 -1644 1228 -1600
rect 1409 -1601 1410 -1525
rect 1423 -1644 1424 -1600
rect 1430 -1601 1431 -1525
rect 1451 -1644 1452 -1600
rect 1472 -1601 1473 -1525
rect 1815 -1644 1816 -1600
rect 1899 -1601 1900 -1525
rect 352 -1603 353 -1525
rect 1430 -1644 1431 -1602
rect 1458 -1603 1459 -1525
rect 1472 -1644 1473 -1602
rect 352 -1644 353 -1604
rect 562 -1605 563 -1525
rect 870 -1605 871 -1525
rect 1276 -1644 1277 -1604
rect 1458 -1644 1459 -1604
rect 1479 -1605 1480 -1525
rect 380 -1607 381 -1525
rect 940 -1644 941 -1606
rect 1094 -1607 1095 -1525
rect 1409 -1644 1410 -1606
rect 1479 -1644 1480 -1606
rect 1486 -1607 1487 -1525
rect 380 -1644 381 -1608
rect 492 -1609 493 -1525
rect 534 -1609 535 -1525
rect 597 -1644 598 -1608
rect 786 -1609 787 -1525
rect 870 -1644 871 -1608
rect 891 -1644 892 -1608
rect 1178 -1609 1179 -1525
rect 1206 -1644 1207 -1608
rect 1899 -1644 1900 -1608
rect 394 -1611 395 -1525
rect 492 -1644 493 -1610
rect 541 -1644 542 -1610
rect 576 -1644 577 -1610
rect 744 -1611 745 -1525
rect 786 -1644 787 -1610
rect 898 -1611 899 -1525
rect 912 -1644 913 -1610
rect 1045 -1611 1046 -1525
rect 1094 -1644 1095 -1610
rect 1244 -1644 1245 -1610
rect 1556 -1644 1557 -1610
rect 173 -1644 174 -1612
rect 744 -1644 745 -1612
rect 898 -1644 899 -1612
rect 1066 -1613 1067 -1525
rect 1087 -1613 1088 -1525
rect 1178 -1644 1179 -1612
rect 1486 -1644 1487 -1612
rect 1500 -1613 1501 -1525
rect 82 -1644 83 -1614
rect 1087 -1644 1088 -1614
rect 1500 -1644 1501 -1614
rect 1675 -1615 1676 -1525
rect 394 -1644 395 -1616
rect 835 -1644 836 -1616
rect 1017 -1617 1018 -1525
rect 1066 -1644 1067 -1616
rect 1675 -1644 1676 -1616
rect 1738 -1617 1739 -1525
rect 471 -1619 472 -1525
rect 534 -1644 535 -1618
rect 562 -1644 563 -1618
rect 1157 -1619 1158 -1525
rect 1738 -1644 1739 -1618
rect 1745 -1619 1746 -1525
rect 471 -1644 472 -1620
rect 527 -1621 528 -1525
rect 779 -1621 780 -1525
rect 1017 -1644 1018 -1620
rect 1045 -1644 1046 -1620
rect 1335 -1644 1336 -1620
rect 1745 -1644 1746 -1620
rect 1773 -1621 1774 -1525
rect 408 -1623 409 -1525
rect 527 -1644 528 -1622
rect 695 -1623 696 -1525
rect 779 -1644 780 -1622
rect 1143 -1623 1144 -1525
rect 1157 -1644 1158 -1622
rect 1759 -1623 1760 -1525
rect 1773 -1644 1774 -1622
rect 408 -1644 409 -1624
rect 590 -1625 591 -1525
rect 1052 -1625 1053 -1525
rect 1143 -1644 1144 -1624
rect 1759 -1644 1760 -1624
rect 2007 -1625 2008 -1525
rect 590 -1644 591 -1626
rect 716 -1627 717 -1525
rect 1052 -1644 1053 -1626
rect 1892 -1627 1893 -1525
rect 240 -1629 241 -1525
rect 1892 -1644 1893 -1628
rect 240 -1644 241 -1630
rect 401 -1631 402 -1525
rect 716 -1644 717 -1630
rect 758 -1631 759 -1525
rect 401 -1644 402 -1632
rect 436 -1633 437 -1525
rect 737 -1633 738 -1525
rect 758 -1644 759 -1632
rect 373 -1635 374 -1525
rect 436 -1644 437 -1634
rect 625 -1635 626 -1525
rect 737 -1644 738 -1634
rect 275 -1637 276 -1525
rect 373 -1644 374 -1636
rect 604 -1637 605 -1525
rect 625 -1644 626 -1636
rect 149 -1639 150 -1525
rect 275 -1644 276 -1638
rect 604 -1644 605 -1638
rect 639 -1639 640 -1525
rect 149 -1644 150 -1640
rect 170 -1644 171 -1640
rect 632 -1641 633 -1525
rect 639 -1644 640 -1640
rect 632 -1644 633 -1642
rect 831 -1644 832 -1642
rect 9 -1654 10 -1652
rect 663 -1654 664 -1652
rect 670 -1654 671 -1652
rect 716 -1654 717 -1652
rect 737 -1654 738 -1652
rect 1556 -1654 1557 -1652
rect 1570 -1654 1571 -1652
rect 1570 -1773 1571 -1653
rect 1570 -1654 1571 -1652
rect 1570 -1773 1571 -1653
rect 1801 -1654 1802 -1652
rect 1801 -1773 1802 -1653
rect 1801 -1654 1802 -1652
rect 1801 -1773 1802 -1653
rect 1843 -1654 1844 -1652
rect 1934 -1654 1935 -1652
rect 1937 -1773 1938 -1653
rect 1976 -1654 1977 -1652
rect 2018 -1654 2019 -1652
rect 2018 -1773 2019 -1653
rect 2018 -1654 2019 -1652
rect 2018 -1773 2019 -1653
rect 9 -1773 10 -1655
rect 128 -1656 129 -1652
rect 131 -1773 132 -1655
rect 1101 -1656 1102 -1652
rect 1206 -1656 1207 -1652
rect 1703 -1656 1704 -1652
rect 1815 -1656 1816 -1652
rect 1843 -1773 1844 -1655
rect 1850 -1656 1851 -1652
rect 1934 -1773 1935 -1655
rect 1941 -1656 1942 -1652
rect 1969 -1773 1970 -1655
rect 44 -1658 45 -1652
rect 79 -1773 80 -1657
rect 86 -1773 87 -1657
rect 275 -1658 276 -1652
rect 324 -1658 325 -1652
rect 558 -1773 559 -1657
rect 590 -1658 591 -1652
rect 831 -1658 832 -1652
rect 842 -1658 843 -1652
rect 1104 -1773 1105 -1657
rect 1206 -1773 1207 -1657
rect 1290 -1658 1291 -1652
rect 1332 -1658 1333 -1652
rect 1815 -1773 1816 -1657
rect 1850 -1773 1851 -1657
rect 1857 -1658 1858 -1652
rect 1871 -1658 1872 -1652
rect 1871 -1773 1872 -1657
rect 1871 -1658 1872 -1652
rect 1871 -1773 1872 -1657
rect 1885 -1658 1886 -1652
rect 1885 -1773 1886 -1657
rect 1885 -1658 1886 -1652
rect 1885 -1773 1886 -1657
rect 1913 -1658 1914 -1652
rect 1913 -1773 1914 -1657
rect 1913 -1658 1914 -1652
rect 1913 -1773 1914 -1657
rect 1944 -1773 1945 -1657
rect 1962 -1773 1963 -1657
rect 37 -1660 38 -1652
rect 44 -1773 45 -1659
rect 51 -1660 52 -1652
rect 51 -1773 52 -1659
rect 51 -1660 52 -1652
rect 51 -1773 52 -1659
rect 65 -1660 66 -1652
rect 177 -1773 178 -1659
rect 180 -1660 181 -1652
rect 359 -1660 360 -1652
rect 422 -1660 423 -1652
rect 425 -1712 426 -1659
rect 485 -1660 486 -1652
rect 684 -1773 685 -1659
rect 709 -1660 710 -1652
rect 1395 -1660 1396 -1652
rect 1451 -1660 1452 -1652
rect 1451 -1773 1452 -1659
rect 1451 -1660 1452 -1652
rect 1451 -1773 1452 -1659
rect 1468 -1660 1469 -1652
rect 1696 -1660 1697 -1652
rect 1857 -1773 1858 -1659
rect 1864 -1660 1865 -1652
rect 1948 -1660 1949 -1652
rect 1955 -1773 1956 -1659
rect 37 -1773 38 -1661
rect 58 -1662 59 -1652
rect 68 -1773 69 -1661
rect 534 -1662 535 -1652
rect 541 -1662 542 -1652
rect 772 -1662 773 -1652
rect 793 -1662 794 -1652
rect 1038 -1662 1039 -1652
rect 1055 -1662 1056 -1652
rect 1297 -1662 1298 -1652
rect 1332 -1773 1333 -1661
rect 1416 -1662 1417 -1652
rect 1468 -1773 1469 -1661
rect 1710 -1662 1711 -1652
rect 1822 -1662 1823 -1652
rect 1864 -1773 1865 -1661
rect 1941 -1773 1942 -1661
rect 1948 -1773 1949 -1661
rect 58 -1773 59 -1663
rect 429 -1664 430 -1652
rect 478 -1664 479 -1652
rect 485 -1773 486 -1663
rect 534 -1773 535 -1663
rect 625 -1664 626 -1652
rect 688 -1664 689 -1652
rect 709 -1773 710 -1663
rect 712 -1664 713 -1652
rect 1038 -1773 1039 -1663
rect 1076 -1773 1077 -1663
rect 1353 -1664 1354 -1652
rect 1395 -1773 1396 -1663
rect 1402 -1664 1403 -1652
rect 1416 -1773 1417 -1663
rect 1423 -1664 1424 -1652
rect 1500 -1664 1501 -1652
rect 1780 -1664 1781 -1652
rect 1794 -1664 1795 -1652
rect 1822 -1773 1823 -1663
rect 72 -1666 73 -1652
rect 82 -1666 83 -1652
rect 89 -1666 90 -1652
rect 1689 -1666 1690 -1652
rect 1696 -1773 1697 -1665
rect 1759 -1666 1760 -1652
rect 1766 -1666 1767 -1652
rect 1794 -1773 1795 -1665
rect 72 -1773 73 -1667
rect 660 -1668 661 -1652
rect 688 -1773 689 -1667
rect 989 -1668 990 -1652
rect 1083 -1773 1084 -1667
rect 1920 -1668 1921 -1652
rect 117 -1670 118 -1652
rect 1164 -1670 1165 -1652
rect 1220 -1670 1221 -1652
rect 1290 -1773 1291 -1669
rect 1297 -1773 1298 -1669
rect 1465 -1670 1466 -1652
rect 1556 -1773 1557 -1669
rect 1563 -1670 1564 -1652
rect 1640 -1670 1641 -1652
rect 1689 -1773 1690 -1669
rect 1731 -1670 1732 -1652
rect 1759 -1773 1760 -1669
rect 1906 -1670 1907 -1652
rect 1920 -1773 1921 -1669
rect 128 -1773 129 -1671
rect 968 -1672 969 -1652
rect 985 -1773 986 -1671
rect 1213 -1672 1214 -1652
rect 1262 -1672 1263 -1652
rect 1262 -1773 1263 -1671
rect 1262 -1672 1263 -1652
rect 1262 -1773 1263 -1671
rect 1286 -1672 1287 -1652
rect 1927 -1672 1928 -1652
rect 156 -1674 157 -1652
rect 394 -1674 395 -1652
rect 422 -1773 423 -1673
rect 499 -1674 500 -1652
rect 523 -1773 524 -1673
rect 1780 -1773 1781 -1673
rect 1899 -1674 1900 -1652
rect 1906 -1773 1907 -1673
rect 114 -1676 115 -1652
rect 394 -1773 395 -1675
rect 429 -1773 430 -1675
rect 436 -1676 437 -1652
rect 499 -1773 500 -1675
rect 1283 -1676 1284 -1652
rect 1335 -1676 1336 -1652
rect 1738 -1676 1739 -1652
rect 1752 -1676 1753 -1652
rect 1766 -1773 1767 -1675
rect 1892 -1676 1893 -1652
rect 1899 -1773 1900 -1675
rect 114 -1773 115 -1677
rect 443 -1678 444 -1652
rect 541 -1773 542 -1677
rect 740 -1678 741 -1652
rect 751 -1678 752 -1652
rect 1402 -1773 1403 -1677
rect 1423 -1773 1424 -1677
rect 1437 -1678 1438 -1652
rect 1521 -1678 1522 -1652
rect 1563 -1773 1564 -1677
rect 1619 -1678 1620 -1652
rect 1640 -1773 1641 -1677
rect 1654 -1678 1655 -1652
rect 1703 -1773 1704 -1677
rect 1717 -1678 1718 -1652
rect 1731 -1773 1732 -1677
rect 1752 -1773 1753 -1677
rect 1773 -1678 1774 -1652
rect 1787 -1678 1788 -1652
rect 1892 -1773 1893 -1677
rect 149 -1680 150 -1652
rect 436 -1773 437 -1679
rect 443 -1773 444 -1679
rect 646 -1680 647 -1652
rect 660 -1773 661 -1679
rect 940 -1680 941 -1652
rect 943 -1680 944 -1652
rect 1724 -1680 1725 -1652
rect 121 -1682 122 -1652
rect 149 -1773 150 -1681
rect 156 -1773 157 -1681
rect 317 -1682 318 -1652
rect 324 -1773 325 -1681
rect 408 -1682 409 -1652
rect 481 -1773 482 -1681
rect 751 -1773 752 -1681
rect 765 -1773 766 -1681
rect 863 -1682 864 -1652
rect 901 -1773 902 -1681
rect 1024 -1682 1025 -1652
rect 1087 -1682 1088 -1652
rect 1472 -1682 1473 -1652
rect 1493 -1682 1494 -1652
rect 1619 -1773 1620 -1681
rect 1626 -1682 1627 -1652
rect 1738 -1773 1739 -1681
rect 121 -1773 122 -1683
rect 814 -1684 815 -1652
rect 828 -1684 829 -1652
rect 1111 -1773 1112 -1683
rect 1185 -1684 1186 -1652
rect 1213 -1773 1214 -1683
rect 1241 -1684 1242 -1652
rect 1654 -1773 1655 -1683
rect 1675 -1684 1676 -1652
rect 1787 -1773 1788 -1683
rect 184 -1686 185 -1652
rect 667 -1686 668 -1652
rect 702 -1686 703 -1652
rect 793 -1773 794 -1685
rect 800 -1686 801 -1652
rect 800 -1773 801 -1685
rect 800 -1686 801 -1652
rect 800 -1773 801 -1685
rect 831 -1773 832 -1685
rect 1318 -1686 1319 -1652
rect 1339 -1686 1340 -1652
rect 1437 -1773 1438 -1685
rect 1472 -1773 1473 -1685
rect 1479 -1686 1480 -1652
rect 1591 -1686 1592 -1652
rect 1626 -1773 1627 -1685
rect 1682 -1686 1683 -1652
rect 1710 -1773 1711 -1685
rect 187 -1773 188 -1687
rect 1276 -1688 1277 -1652
rect 1311 -1688 1312 -1652
rect 1493 -1773 1494 -1687
rect 1542 -1688 1543 -1652
rect 1591 -1773 1592 -1687
rect 1668 -1688 1669 -1652
rect 1682 -1773 1683 -1687
rect 100 -1690 101 -1652
rect 1542 -1773 1543 -1689
rect 1661 -1690 1662 -1652
rect 1668 -1773 1669 -1689
rect 2 -1692 3 -1652
rect 100 -1773 101 -1691
rect 201 -1773 202 -1691
rect 649 -1773 650 -1691
rect 716 -1773 717 -1691
rect 1073 -1692 1074 -1652
rect 1101 -1773 1102 -1691
rect 1675 -1773 1676 -1691
rect 205 -1694 206 -1652
rect 208 -1712 209 -1693
rect 254 -1694 255 -1652
rect 397 -1694 398 -1652
rect 408 -1773 409 -1693
rect 562 -1694 563 -1652
rect 583 -1694 584 -1652
rect 625 -1773 626 -1693
rect 639 -1694 640 -1652
rect 814 -1773 815 -1693
rect 842 -1773 843 -1693
rect 877 -1694 878 -1652
rect 919 -1694 920 -1652
rect 1584 -1694 1585 -1652
rect 1661 -1773 1662 -1693
rect 1745 -1694 1746 -1652
rect 191 -1696 192 -1652
rect 254 -1773 255 -1695
rect 275 -1773 276 -1695
rect 450 -1696 451 -1652
rect 520 -1696 521 -1652
rect 702 -1773 703 -1695
rect 737 -1773 738 -1695
rect 810 -1773 811 -1695
rect 856 -1696 857 -1652
rect 856 -1773 857 -1695
rect 856 -1696 857 -1652
rect 856 -1773 857 -1695
rect 863 -1773 864 -1695
rect 912 -1696 913 -1652
rect 919 -1773 920 -1695
rect 1209 -1696 1210 -1652
rect 1241 -1773 1242 -1695
rect 1500 -1773 1501 -1695
rect 1584 -1773 1585 -1695
rect 1598 -1696 1599 -1652
rect 1745 -1773 1746 -1695
rect 1836 -1696 1837 -1652
rect 191 -1773 192 -1697
rect 418 -1698 419 -1652
rect 576 -1698 577 -1652
rect 639 -1773 640 -1697
rect 740 -1773 741 -1697
rect 1430 -1698 1431 -1652
rect 1479 -1773 1480 -1697
rect 1486 -1698 1487 -1652
rect 1598 -1773 1599 -1697
rect 1612 -1698 1613 -1652
rect 1808 -1698 1809 -1652
rect 1836 -1773 1837 -1697
rect 198 -1700 199 -1652
rect 450 -1773 451 -1699
rect 527 -1700 528 -1652
rect 576 -1773 577 -1699
rect 583 -1773 584 -1699
rect 681 -1700 682 -1652
rect 768 -1700 769 -1652
rect 989 -1773 990 -1699
rect 1024 -1773 1025 -1699
rect 1136 -1700 1137 -1652
rect 1185 -1773 1186 -1699
rect 1199 -1700 1200 -1652
rect 1244 -1700 1245 -1652
rect 1717 -1773 1718 -1699
rect 198 -1773 199 -1701
rect 849 -1702 850 -1652
rect 877 -1773 878 -1701
rect 961 -1702 962 -1652
rect 968 -1773 969 -1701
rect 1045 -1702 1046 -1652
rect 1073 -1773 1074 -1701
rect 1829 -1702 1830 -1652
rect 205 -1773 206 -1703
rect 492 -1704 493 -1652
rect 527 -1773 528 -1703
rect 632 -1704 633 -1652
rect 681 -1773 682 -1703
rect 1773 -1773 1774 -1703
rect 219 -1706 220 -1652
rect 1045 -1773 1046 -1705
rect 1129 -1706 1130 -1652
rect 1808 -1773 1809 -1705
rect 219 -1773 220 -1707
rect 261 -1708 262 -1652
rect 317 -1773 318 -1707
rect 338 -1708 339 -1652
rect 359 -1773 360 -1707
rect 457 -1708 458 -1652
rect 492 -1773 493 -1707
rect 730 -1708 731 -1652
rect 772 -1773 773 -1707
rect 1066 -1708 1067 -1652
rect 1122 -1708 1123 -1652
rect 1129 -1773 1130 -1707
rect 1132 -1708 1133 -1652
rect 1829 -1773 1830 -1707
rect 261 -1773 262 -1709
rect 506 -1710 507 -1652
rect 590 -1773 591 -1709
rect 597 -1710 598 -1652
rect 604 -1710 605 -1652
rect 667 -1773 668 -1709
rect 786 -1710 787 -1652
rect 1283 -1773 1284 -1709
rect 1311 -1773 1312 -1709
rect 1465 -1773 1466 -1709
rect 1612 -1773 1613 -1709
rect 1647 -1710 1648 -1652
rect 310 -1712 311 -1652
rect 338 -1773 339 -1711
rect 373 -1712 374 -1652
rect 418 -1773 419 -1711
rect 786 -1773 787 -1711
rect 849 -1773 850 -1711
rect 898 -1712 899 -1652
rect 912 -1773 913 -1711
rect 926 -1712 927 -1652
rect 933 -1712 934 -1652
rect 1521 -1773 1522 -1711
rect 282 -1714 283 -1652
rect 310 -1773 311 -1713
rect 373 -1773 374 -1713
rect 401 -1714 402 -1652
rect 457 -1773 458 -1713
rect 464 -1714 465 -1652
rect 506 -1773 507 -1713
rect 723 -1714 724 -1652
rect 922 -1714 923 -1652
rect 947 -1714 948 -1652
rect 961 -1773 962 -1713
rect 1003 -1714 1004 -1652
rect 1041 -1714 1042 -1652
rect 1122 -1773 1123 -1713
rect 1136 -1773 1137 -1713
rect 1157 -1714 1158 -1652
rect 1199 -1773 1200 -1713
rect 1248 -1714 1249 -1652
rect 1269 -1714 1270 -1652
rect 1276 -1773 1277 -1713
rect 1318 -1773 1319 -1713
rect 1927 -1773 1928 -1713
rect 142 -1716 143 -1652
rect 401 -1773 402 -1715
rect 569 -1716 570 -1652
rect 604 -1773 605 -1715
rect 632 -1773 633 -1715
rect 698 -1773 699 -1715
rect 723 -1773 724 -1715
rect 870 -1716 871 -1652
rect 943 -1773 944 -1715
rect 1087 -1773 1088 -1715
rect 1157 -1773 1158 -1715
rect 1192 -1716 1193 -1652
rect 1244 -1773 1245 -1715
rect 1605 -1716 1606 -1652
rect 93 -1718 94 -1652
rect 142 -1773 143 -1717
rect 194 -1773 195 -1717
rect 1605 -1773 1606 -1717
rect 93 -1773 94 -1719
rect 600 -1773 601 -1719
rect 653 -1720 654 -1652
rect 926 -1773 927 -1719
rect 947 -1773 948 -1719
rect 982 -1720 983 -1652
rect 996 -1720 997 -1652
rect 1003 -1773 1004 -1719
rect 1066 -1773 1067 -1719
rect 1150 -1720 1151 -1652
rect 1192 -1773 1193 -1719
rect 1346 -1720 1347 -1652
rect 1353 -1773 1354 -1719
rect 1633 -1720 1634 -1652
rect 16 -1722 17 -1652
rect 982 -1773 983 -1721
rect 1010 -1722 1011 -1652
rect 1633 -1773 1634 -1721
rect 16 -1773 17 -1723
rect 170 -1724 171 -1652
rect 184 -1773 185 -1723
rect 1010 -1773 1011 -1723
rect 1150 -1773 1151 -1723
rect 1178 -1724 1179 -1652
rect 1248 -1773 1249 -1723
rect 1325 -1724 1326 -1652
rect 1339 -1773 1340 -1723
rect 1514 -1724 1515 -1652
rect 170 -1773 171 -1725
rect 268 -1726 269 -1652
rect 397 -1773 398 -1725
rect 821 -1726 822 -1652
rect 870 -1773 871 -1725
rect 905 -1726 906 -1652
rect 971 -1726 972 -1652
rect 1486 -1773 1487 -1725
rect 1507 -1726 1508 -1652
rect 1514 -1773 1515 -1725
rect 233 -1728 234 -1652
rect 464 -1773 465 -1727
rect 569 -1773 570 -1727
rect 611 -1728 612 -1652
rect 646 -1773 647 -1727
rect 996 -1773 997 -1727
rect 1171 -1728 1172 -1652
rect 1178 -1773 1179 -1727
rect 1227 -1728 1228 -1652
rect 1325 -1773 1326 -1727
rect 1356 -1728 1357 -1652
rect 1724 -1773 1725 -1727
rect 233 -1773 234 -1729
rect 303 -1730 304 -1652
rect 597 -1773 598 -1729
rect 1164 -1773 1165 -1729
rect 1220 -1773 1221 -1729
rect 1356 -1773 1357 -1729
rect 1388 -1730 1389 -1652
rect 1430 -1773 1431 -1729
rect 1507 -1773 1508 -1729
rect 1577 -1730 1578 -1652
rect 240 -1732 241 -1652
rect 303 -1773 304 -1731
rect 611 -1773 612 -1731
rect 618 -1732 619 -1652
rect 653 -1773 654 -1731
rect 1304 -1732 1305 -1652
rect 1388 -1773 1389 -1731
rect 1444 -1732 1445 -1652
rect 226 -1734 227 -1652
rect 618 -1773 619 -1733
rect 821 -1773 822 -1733
rect 835 -1734 836 -1652
rect 891 -1734 892 -1652
rect 1346 -1773 1347 -1733
rect 1444 -1773 1445 -1733
rect 1535 -1734 1536 -1652
rect 226 -1773 227 -1735
rect 331 -1736 332 -1652
rect 807 -1736 808 -1652
rect 835 -1773 836 -1735
rect 891 -1773 892 -1735
rect 954 -1736 955 -1652
rect 1080 -1736 1081 -1652
rect 1171 -1773 1172 -1735
rect 1227 -1773 1228 -1735
rect 1234 -1736 1235 -1652
rect 1269 -1773 1270 -1735
rect 1360 -1736 1361 -1652
rect 1528 -1736 1529 -1652
rect 1535 -1773 1536 -1735
rect 240 -1773 241 -1737
rect 415 -1773 416 -1737
rect 898 -1773 899 -1737
rect 1577 -1773 1578 -1737
rect 247 -1740 248 -1652
rect 282 -1773 283 -1739
rect 331 -1773 332 -1739
rect 352 -1740 353 -1652
rect 905 -1773 906 -1739
rect 975 -1740 976 -1652
rect 1234 -1773 1235 -1739
rect 1367 -1740 1368 -1652
rect 1528 -1773 1529 -1739
rect 1549 -1740 1550 -1652
rect 247 -1773 248 -1741
rect 345 -1742 346 -1652
rect 352 -1773 353 -1741
rect 548 -1742 549 -1652
rect 933 -1773 934 -1741
rect 1080 -1773 1081 -1741
rect 1304 -1773 1305 -1741
rect 1647 -1773 1648 -1741
rect 268 -1773 269 -1743
rect 366 -1744 367 -1652
rect 513 -1744 514 -1652
rect 548 -1773 549 -1743
rect 954 -1773 955 -1743
rect 1878 -1744 1879 -1652
rect 23 -1746 24 -1652
rect 366 -1773 367 -1745
rect 513 -1773 514 -1745
rect 674 -1746 675 -1652
rect 975 -1773 976 -1745
rect 1017 -1746 1018 -1652
rect 1307 -1746 1308 -1652
rect 1878 -1773 1879 -1745
rect 23 -1773 24 -1747
rect 544 -1748 545 -1652
rect 674 -1773 675 -1747
rect 779 -1748 780 -1652
rect 1052 -1748 1053 -1652
rect 1307 -1773 1308 -1747
rect 1360 -1773 1361 -1747
rect 1363 -1773 1364 -1747
rect 1367 -1773 1368 -1747
rect 1458 -1748 1459 -1652
rect 289 -1750 290 -1652
rect 345 -1773 346 -1749
rect 744 -1750 745 -1652
rect 1017 -1773 1018 -1749
rect 1052 -1773 1053 -1749
rect 1108 -1750 1109 -1652
rect 1374 -1750 1375 -1652
rect 1458 -1773 1459 -1749
rect 289 -1773 290 -1751
rect 380 -1752 381 -1652
rect 744 -1773 745 -1751
rect 758 -1752 759 -1652
rect 779 -1773 780 -1751
rect 1031 -1752 1032 -1652
rect 1374 -1773 1375 -1751
rect 1381 -1752 1382 -1652
rect 1409 -1752 1410 -1652
rect 1549 -1773 1550 -1751
rect 107 -1754 108 -1652
rect 380 -1773 381 -1753
rect 758 -1773 759 -1753
rect 884 -1754 885 -1652
rect 1031 -1773 1032 -1753
rect 1094 -1754 1095 -1652
rect 1115 -1754 1116 -1652
rect 1409 -1773 1410 -1753
rect 107 -1773 108 -1755
rect 135 -1756 136 -1652
rect 695 -1756 696 -1652
rect 1094 -1773 1095 -1755
rect 1115 -1773 1116 -1755
rect 1143 -1756 1144 -1652
rect 1381 -1773 1382 -1755
rect 1846 -1756 1847 -1652
rect 135 -1773 136 -1757
rect 163 -1758 164 -1652
rect 565 -1773 566 -1757
rect 1143 -1773 1144 -1757
rect 163 -1773 164 -1759
rect 212 -1760 213 -1652
rect 695 -1773 696 -1759
rect 1059 -1760 1060 -1652
rect 212 -1773 213 -1761
rect 387 -1762 388 -1652
rect 1059 -1773 1060 -1761
rect 1255 -1762 1256 -1652
rect 296 -1764 297 -1652
rect 387 -1773 388 -1763
rect 516 -1773 517 -1763
rect 1255 -1773 1256 -1763
rect 296 -1773 297 -1765
rect 471 -1766 472 -1652
rect 30 -1768 31 -1652
rect 471 -1773 472 -1767
rect 30 -1773 31 -1769
rect 555 -1770 556 -1652
rect 555 -1773 556 -1771
rect 887 -1773 888 -1771
rect 65 -1783 66 -1781
rect 75 -1857 76 -1782
rect 93 -1783 94 -1781
rect 145 -1898 146 -1782
rect 170 -1783 171 -1781
rect 523 -1783 524 -1781
rect 527 -1783 528 -1781
rect 530 -1783 531 -1781
rect 555 -1783 556 -1781
rect 793 -1783 794 -1781
rect 810 -1783 811 -1781
rect 1927 -1783 1928 -1781
rect 1955 -1783 1956 -1781
rect 1997 -1898 1998 -1782
rect 2011 -1898 2012 -1782
rect 2018 -1783 2019 -1781
rect 65 -1898 66 -1784
rect 275 -1785 276 -1781
rect 282 -1785 283 -1781
rect 481 -1785 482 -1781
rect 506 -1785 507 -1781
rect 555 -1898 556 -1784
rect 590 -1785 591 -1781
rect 590 -1898 591 -1784
rect 590 -1785 591 -1781
rect 590 -1898 591 -1784
rect 597 -1785 598 -1781
rect 870 -1785 871 -1781
rect 884 -1785 885 -1781
rect 1689 -1785 1690 -1781
rect 1878 -1785 1879 -1781
rect 1955 -1898 1956 -1784
rect 1962 -1785 1963 -1781
rect 2018 -1898 2019 -1784
rect 93 -1898 94 -1786
rect 107 -1787 108 -1781
rect 114 -1787 115 -1781
rect 191 -1787 192 -1781
rect 198 -1787 199 -1781
rect 877 -1787 878 -1781
rect 884 -1898 885 -1786
rect 2004 -1898 2005 -1786
rect 107 -1898 108 -1788
rect 499 -1789 500 -1781
rect 527 -1898 528 -1788
rect 1073 -1789 1074 -1781
rect 1080 -1789 1081 -1781
rect 1689 -1898 1690 -1788
rect 1878 -1898 1879 -1788
rect 1941 -1789 1942 -1781
rect 1969 -1789 1970 -1781
rect 2025 -1898 2026 -1788
rect 114 -1898 115 -1790
rect 212 -1791 213 -1781
rect 254 -1791 255 -1781
rect 691 -1898 692 -1790
rect 695 -1791 696 -1781
rect 926 -1791 927 -1781
rect 943 -1791 944 -1781
rect 1493 -1791 1494 -1781
rect 1500 -1791 1501 -1781
rect 1500 -1898 1501 -1790
rect 1500 -1791 1501 -1781
rect 1500 -1898 1501 -1790
rect 1521 -1791 1522 -1781
rect 1521 -1898 1522 -1790
rect 1521 -1791 1522 -1781
rect 1521 -1898 1522 -1790
rect 1566 -1898 1567 -1790
rect 1885 -1791 1886 -1781
rect 1892 -1791 1893 -1781
rect 1962 -1898 1963 -1790
rect 58 -1793 59 -1781
rect 212 -1898 213 -1792
rect 254 -1898 255 -1792
rect 289 -1793 290 -1781
rect 303 -1793 304 -1781
rect 303 -1898 304 -1792
rect 303 -1793 304 -1781
rect 303 -1898 304 -1792
rect 310 -1793 311 -1781
rect 807 -1898 808 -1792
rect 870 -1898 871 -1792
rect 933 -1793 934 -1781
rect 947 -1793 948 -1781
rect 947 -1898 948 -1792
rect 947 -1793 948 -1781
rect 947 -1898 948 -1792
rect 968 -1793 969 -1781
rect 968 -1898 969 -1792
rect 968 -1793 969 -1781
rect 968 -1898 969 -1792
rect 985 -1898 986 -1792
rect 1570 -1793 1571 -1781
rect 1584 -1793 1585 -1781
rect 1584 -1898 1585 -1792
rect 1584 -1793 1585 -1781
rect 1584 -1898 1585 -1792
rect 1619 -1793 1620 -1781
rect 1619 -1898 1620 -1792
rect 1619 -1793 1620 -1781
rect 1619 -1898 1620 -1792
rect 1829 -1793 1830 -1781
rect 1885 -1898 1886 -1792
rect 1899 -1793 1900 -1781
rect 1969 -1898 1970 -1792
rect 16 -1795 17 -1781
rect 58 -1898 59 -1794
rect 128 -1898 129 -1794
rect 135 -1795 136 -1781
rect 138 -1898 139 -1794
rect 289 -1898 290 -1794
rect 352 -1795 353 -1781
rect 488 -1898 489 -1794
rect 499 -1898 500 -1794
rect 625 -1795 626 -1781
rect 649 -1795 650 -1781
rect 814 -1795 815 -1781
rect 898 -1898 899 -1794
rect 1038 -1795 1039 -1781
rect 1059 -1795 1060 -1781
rect 1076 -1795 1077 -1781
rect 1080 -1898 1081 -1794
rect 1087 -1795 1088 -1781
rect 1090 -1898 1091 -1794
rect 1206 -1795 1207 -1781
rect 1209 -1898 1210 -1794
rect 1626 -1795 1627 -1781
rect 1731 -1795 1732 -1781
rect 1829 -1898 1830 -1794
rect 1843 -1795 1844 -1781
rect 1892 -1898 1893 -1794
rect 1906 -1795 1907 -1781
rect 1983 -1898 1984 -1794
rect 9 -1797 10 -1781
rect 135 -1898 136 -1796
rect 142 -1797 143 -1781
rect 310 -1898 311 -1796
rect 352 -1898 353 -1796
rect 359 -1797 360 -1781
rect 366 -1797 367 -1781
rect 562 -1797 563 -1781
rect 583 -1797 584 -1781
rect 597 -1898 598 -1796
rect 600 -1797 601 -1781
rect 702 -1797 703 -1781
rect 719 -1898 720 -1796
rect 730 -1797 731 -1781
rect 744 -1797 745 -1781
rect 744 -1898 745 -1796
rect 744 -1797 745 -1781
rect 744 -1898 745 -1796
rect 751 -1797 752 -1781
rect 877 -1898 878 -1796
rect 908 -1898 909 -1796
rect 1094 -1797 1095 -1781
rect 1104 -1797 1105 -1781
rect 1444 -1797 1445 -1781
rect 1468 -1797 1469 -1781
rect 1920 -1797 1921 -1781
rect 16 -1898 17 -1798
rect 51 -1799 52 -1781
rect 121 -1799 122 -1781
rect 625 -1898 626 -1798
rect 639 -1799 640 -1781
rect 702 -1898 703 -1798
rect 730 -1898 731 -1798
rect 1381 -1799 1382 -1781
rect 1409 -1799 1410 -1781
rect 1990 -1898 1991 -1798
rect 37 -1801 38 -1781
rect 51 -1898 52 -1800
rect 79 -1801 80 -1781
rect 121 -1898 122 -1800
rect 131 -1801 132 -1781
rect 366 -1898 367 -1800
rect 387 -1801 388 -1781
rect 639 -1898 640 -1800
rect 660 -1801 661 -1781
rect 660 -1898 661 -1800
rect 660 -1801 661 -1781
rect 660 -1898 661 -1800
rect 681 -1801 682 -1781
rect 793 -1898 794 -1800
rect 814 -1898 815 -1800
rect 842 -1801 843 -1781
rect 954 -1801 955 -1781
rect 1038 -1898 1039 -1800
rect 1059 -1898 1060 -1800
rect 1290 -1801 1291 -1781
rect 1304 -1801 1305 -1781
rect 1773 -1801 1774 -1781
rect 1850 -1801 1851 -1781
rect 1906 -1898 1907 -1800
rect 1913 -1801 1914 -1781
rect 1920 -1898 1921 -1800
rect 37 -1898 38 -1802
rect 142 -1898 143 -1802
rect 156 -1803 157 -1781
rect 282 -1898 283 -1802
rect 387 -1898 388 -1802
rect 509 -1898 510 -1802
rect 562 -1898 563 -1802
rect 604 -1803 605 -1781
rect 632 -1803 633 -1781
rect 681 -1898 682 -1802
rect 684 -1803 685 -1781
rect 936 -1898 937 -1802
rect 1010 -1803 1011 -1781
rect 1010 -1898 1011 -1802
rect 1010 -1803 1011 -1781
rect 1010 -1898 1011 -1802
rect 1017 -1803 1018 -1781
rect 1094 -1898 1095 -1802
rect 1104 -1898 1105 -1802
rect 1213 -1803 1214 -1781
rect 1244 -1803 1245 -1781
rect 1640 -1803 1641 -1781
rect 1717 -1803 1718 -1781
rect 1773 -1898 1774 -1802
rect 1815 -1803 1816 -1781
rect 1850 -1898 1851 -1802
rect 1871 -1803 1872 -1781
rect 1941 -1898 1942 -1802
rect 79 -1898 80 -1804
rect 653 -1805 654 -1781
rect 765 -1805 766 -1781
rect 842 -1898 843 -1804
rect 1073 -1898 1074 -1804
rect 1171 -1805 1172 -1781
rect 1248 -1805 1249 -1781
rect 1290 -1898 1291 -1804
rect 1304 -1898 1305 -1804
rect 1437 -1805 1438 -1781
rect 1535 -1805 1536 -1781
rect 1843 -1898 1844 -1804
rect 156 -1898 157 -1806
rect 408 -1807 409 -1781
rect 415 -1807 416 -1781
rect 919 -1807 920 -1781
rect 1108 -1807 1109 -1781
rect 1976 -1898 1977 -1806
rect 170 -1898 171 -1808
rect 982 -1898 983 -1808
rect 1111 -1809 1112 -1781
rect 1192 -1809 1193 -1781
rect 1269 -1809 1270 -1781
rect 1353 -1898 1354 -1808
rect 1360 -1809 1361 -1781
rect 1738 -1809 1739 -1781
rect 1745 -1809 1746 -1781
rect 1899 -1898 1900 -1808
rect 177 -1811 178 -1781
rect 275 -1898 276 -1810
rect 401 -1811 402 -1781
rect 940 -1811 941 -1781
rect 1129 -1811 1130 -1781
rect 1129 -1898 1130 -1810
rect 1129 -1811 1130 -1781
rect 1129 -1898 1130 -1810
rect 1136 -1811 1137 -1781
rect 1171 -1898 1172 -1810
rect 1185 -1811 1186 -1781
rect 1248 -1898 1249 -1810
rect 1262 -1811 1263 -1781
rect 1269 -1898 1270 -1810
rect 1283 -1811 1284 -1781
rect 1360 -1898 1361 -1810
rect 1363 -1811 1364 -1781
rect 1927 -1898 1928 -1810
rect 177 -1898 178 -1812
rect 394 -1813 395 -1781
rect 404 -1898 405 -1812
rect 415 -1898 416 -1812
rect 429 -1813 430 -1781
rect 513 -1813 514 -1781
rect 583 -1898 584 -1812
rect 1101 -1898 1102 -1812
rect 1115 -1813 1116 -1781
rect 1136 -1898 1137 -1812
rect 1150 -1813 1151 -1781
rect 1185 -1898 1186 -1812
rect 1276 -1813 1277 -1781
rect 1283 -1898 1284 -1812
rect 1307 -1813 1308 -1781
rect 1787 -1813 1788 -1781
rect 1794 -1813 1795 -1781
rect 1871 -1898 1872 -1812
rect 191 -1898 192 -1814
rect 219 -1815 220 -1781
rect 240 -1815 241 -1781
rect 394 -1898 395 -1814
rect 408 -1898 409 -1814
rect 1125 -1898 1126 -1814
rect 1150 -1898 1151 -1814
rect 1444 -1898 1445 -1814
rect 1535 -1898 1536 -1814
rect 1780 -1815 1781 -1781
rect 1822 -1815 1823 -1781
rect 1913 -1898 1914 -1814
rect 201 -1898 202 -1816
rect 296 -1817 297 -1781
rect 380 -1817 381 -1781
rect 401 -1898 402 -1816
rect 429 -1898 430 -1816
rect 548 -1817 549 -1781
rect 604 -1898 605 -1816
rect 723 -1817 724 -1781
rect 751 -1898 752 -1816
rect 1108 -1898 1109 -1816
rect 1157 -1817 1158 -1781
rect 1192 -1898 1193 -1816
rect 1311 -1817 1312 -1781
rect 1493 -1898 1494 -1816
rect 1563 -1817 1564 -1781
rect 1570 -1898 1571 -1816
rect 1577 -1817 1578 -1781
rect 1745 -1898 1746 -1816
rect 1759 -1817 1760 -1781
rect 1780 -1898 1781 -1816
rect 1801 -1817 1802 -1781
rect 1822 -1898 1823 -1816
rect 187 -1819 188 -1781
rect 1801 -1898 1802 -1818
rect 219 -1898 220 -1820
rect 443 -1821 444 -1781
rect 450 -1821 451 -1781
rect 695 -1898 696 -1820
rect 723 -1898 724 -1820
rect 828 -1821 829 -1781
rect 831 -1821 832 -1781
rect 1437 -1898 1438 -1820
rect 1598 -1821 1599 -1781
rect 1815 -1898 1816 -1820
rect 23 -1823 24 -1781
rect 828 -1898 829 -1822
rect 863 -1823 864 -1781
rect 1311 -1898 1312 -1822
rect 1318 -1823 1319 -1781
rect 1703 -1823 1704 -1781
rect 1738 -1898 1739 -1822
rect 1752 -1823 1753 -1781
rect 1766 -1823 1767 -1781
rect 1794 -1898 1795 -1822
rect 23 -1898 24 -1824
rect 614 -1898 615 -1824
rect 632 -1898 633 -1824
rect 667 -1825 668 -1781
rect 765 -1898 766 -1824
rect 863 -1898 864 -1824
rect 891 -1825 892 -1781
rect 940 -1898 941 -1824
rect 975 -1825 976 -1781
rect 1157 -1898 1158 -1824
rect 1164 -1825 1165 -1781
rect 1213 -1898 1214 -1824
rect 1321 -1825 1322 -1781
rect 1626 -1898 1627 -1824
rect 1654 -1825 1655 -1781
rect 1717 -1898 1718 -1824
rect 72 -1827 73 -1781
rect 450 -1898 451 -1826
rect 464 -1827 465 -1781
rect 520 -1827 521 -1781
rect 541 -1827 542 -1781
rect 548 -1898 549 -1826
rect 576 -1827 577 -1781
rect 667 -1898 668 -1826
rect 768 -1898 769 -1826
rect 1458 -1827 1459 -1781
rect 1486 -1827 1487 -1781
rect 1766 -1898 1767 -1826
rect 44 -1829 45 -1781
rect 72 -1898 73 -1828
rect 100 -1829 101 -1781
rect 975 -1898 976 -1828
rect 1024 -1829 1025 -1781
rect 1164 -1898 1165 -1828
rect 1178 -1829 1179 -1781
rect 1262 -1898 1263 -1828
rect 1325 -1829 1326 -1781
rect 1381 -1898 1382 -1828
rect 1409 -1898 1410 -1828
rect 1549 -1829 1550 -1781
rect 1598 -1898 1599 -1828
rect 1661 -1829 1662 -1781
rect 1696 -1829 1697 -1781
rect 1703 -1898 1704 -1828
rect 30 -1831 31 -1781
rect 1024 -1898 1025 -1830
rect 1083 -1831 1084 -1781
rect 1752 -1898 1753 -1830
rect 30 -1898 31 -1832
rect 226 -1833 227 -1781
rect 240 -1898 241 -1832
rect 373 -1833 374 -1781
rect 443 -1898 444 -1832
rect 464 -1898 465 -1832
rect 611 -1833 612 -1781
rect 772 -1833 773 -1781
rect 1017 -1898 1018 -1832
rect 1143 -1833 1144 -1781
rect 1178 -1898 1179 -1832
rect 1255 -1833 1256 -1781
rect 1325 -1898 1326 -1832
rect 1339 -1833 1340 -1781
rect 1577 -1898 1578 -1832
rect 1605 -1833 1606 -1781
rect 1640 -1898 1641 -1832
rect 1661 -1898 1662 -1832
rect 1836 -1833 1837 -1781
rect 44 -1898 45 -1834
rect 397 -1835 398 -1781
rect 436 -1835 437 -1781
rect 653 -1898 654 -1834
rect 772 -1898 773 -1834
rect 996 -1835 997 -1781
rect 1122 -1835 1123 -1781
rect 1143 -1898 1144 -1834
rect 1199 -1835 1200 -1781
rect 1255 -1898 1256 -1834
rect 1430 -1835 1431 -1781
rect 1731 -1898 1732 -1834
rect 1808 -1835 1809 -1781
rect 1836 -1898 1837 -1834
rect 184 -1837 185 -1781
rect 1318 -1898 1319 -1836
rect 1451 -1837 1452 -1781
rect 1458 -1898 1459 -1836
rect 1479 -1837 1480 -1781
rect 1486 -1898 1487 -1836
rect 1633 -1837 1634 -1781
rect 1654 -1898 1655 -1836
rect 1682 -1837 1683 -1781
rect 1696 -1898 1697 -1836
rect 1710 -1837 1711 -1781
rect 1808 -1898 1809 -1836
rect 163 -1839 164 -1781
rect 184 -1898 185 -1838
rect 205 -1839 206 -1781
rect 373 -1898 374 -1838
rect 380 -1898 381 -1838
rect 422 -1839 423 -1781
rect 485 -1839 486 -1781
rect 541 -1898 542 -1838
rect 558 -1839 559 -1781
rect 1199 -1898 1200 -1838
rect 1234 -1839 1235 -1781
rect 1339 -1898 1340 -1838
rect 1367 -1839 1368 -1781
rect 1479 -1898 1480 -1838
rect 1542 -1839 1543 -1781
rect 1710 -1898 1711 -1838
rect 163 -1898 164 -1840
rect 516 -1841 517 -1781
rect 520 -1898 521 -1840
rect 688 -1841 689 -1781
rect 891 -1898 892 -1840
rect 1241 -1841 1242 -1781
rect 1367 -1898 1368 -1840
rect 1374 -1841 1375 -1781
rect 1388 -1841 1389 -1781
rect 1451 -1898 1452 -1840
rect 1556 -1841 1557 -1781
rect 1633 -1898 1634 -1840
rect 1668 -1841 1669 -1781
rect 1682 -1898 1683 -1840
rect 205 -1898 206 -1842
rect 233 -1843 234 -1781
rect 261 -1843 262 -1781
rect 359 -1898 360 -1842
rect 478 -1843 479 -1781
rect 1542 -1898 1543 -1842
rect 1556 -1898 1557 -1842
rect 1944 -1843 1945 -1781
rect 149 -1845 150 -1781
rect 261 -1898 262 -1844
rect 296 -1898 297 -1844
rect 478 -1898 479 -1844
rect 485 -1898 486 -1844
rect 1787 -1898 1788 -1844
rect 149 -1898 150 -1846
rect 887 -1847 888 -1781
rect 912 -1847 913 -1781
rect 919 -1898 920 -1846
rect 933 -1898 934 -1846
rect 1759 -1898 1760 -1846
rect 226 -1898 227 -1848
rect 345 -1849 346 -1781
rect 492 -1849 493 -1781
rect 887 -1898 888 -1848
rect 912 -1898 913 -1848
rect 961 -1849 962 -1781
rect 996 -1898 997 -1848
rect 1003 -1849 1004 -1781
rect 1045 -1849 1046 -1781
rect 1430 -1898 1431 -1848
rect 1647 -1849 1648 -1781
rect 1668 -1898 1669 -1848
rect 233 -1898 234 -1850
rect 268 -1851 269 -1781
rect 331 -1851 332 -1781
rect 436 -1898 437 -1850
rect 492 -1898 493 -1850
rect 618 -1851 619 -1781
rect 779 -1851 780 -1781
rect 1003 -1898 1004 -1850
rect 1031 -1851 1032 -1781
rect 1045 -1898 1046 -1850
rect 1122 -1898 1123 -1850
rect 1864 -1851 1865 -1781
rect 86 -1853 87 -1781
rect 268 -1898 269 -1852
rect 324 -1853 325 -1781
rect 331 -1898 332 -1852
rect 513 -1898 514 -1852
rect 1153 -1898 1154 -1852
rect 1220 -1853 1221 -1781
rect 1234 -1898 1235 -1852
rect 1241 -1898 1242 -1852
rect 1465 -1853 1466 -1781
rect 1612 -1853 1613 -1781
rect 1647 -1898 1648 -1852
rect 86 -1898 87 -1854
rect 1223 -1898 1224 -1854
rect 1374 -1898 1375 -1854
rect 1395 -1855 1396 -1781
rect 1423 -1855 1424 -1781
rect 1612 -1898 1613 -1854
rect 247 -1857 248 -1781
rect 345 -1898 346 -1856
rect 530 -1898 531 -1856
rect 1115 -1898 1116 -1856
rect 1346 -1857 1347 -1781
rect 1395 -1898 1396 -1856
rect 1416 -1857 1417 -1781
rect 1423 -1898 1424 -1856
rect 1465 -1898 1466 -1856
rect 1528 -1857 1529 -1781
rect 247 -1898 248 -1858
rect 2014 -1898 2015 -1858
rect 317 -1861 318 -1781
rect 324 -1898 325 -1860
rect 579 -1898 580 -1860
rect 1549 -1898 1550 -1860
rect 317 -1898 318 -1862
rect 457 -1863 458 -1781
rect 611 -1898 612 -1862
rect 1605 -1898 1606 -1862
rect 198 -1898 199 -1864
rect 457 -1898 458 -1864
rect 618 -1898 619 -1864
rect 786 -1865 787 -1781
rect 905 -1865 906 -1781
rect 961 -1898 962 -1864
rect 1031 -1898 1032 -1864
rect 1066 -1865 1067 -1781
rect 1111 -1898 1112 -1864
rect 1864 -1898 1865 -1864
rect 422 -1898 423 -1866
rect 905 -1898 906 -1866
rect 954 -1898 955 -1866
rect 1220 -1898 1221 -1866
rect 1297 -1867 1298 -1781
rect 1346 -1898 1347 -1866
rect 1388 -1898 1389 -1866
rect 1402 -1867 1403 -1781
rect 1416 -1898 1417 -1866
rect 1934 -1867 1935 -1781
rect 779 -1898 780 -1868
rect 856 -1869 857 -1781
rect 1052 -1869 1053 -1781
rect 1066 -1898 1067 -1868
rect 1227 -1869 1228 -1781
rect 1297 -1898 1298 -1868
rect 1332 -1869 1333 -1781
rect 1402 -1898 1403 -1868
rect 1528 -1898 1529 -1868
rect 1591 -1869 1592 -1781
rect 1857 -1869 1858 -1781
rect 1934 -1898 1935 -1868
rect 61 -1898 62 -1870
rect 1227 -1898 1228 -1870
rect 1507 -1871 1508 -1781
rect 1591 -1898 1592 -1870
rect 68 -1873 69 -1781
rect 1857 -1898 1858 -1872
rect 103 -1898 104 -1874
rect 856 -1898 857 -1874
rect 989 -1875 990 -1781
rect 1052 -1898 1053 -1874
rect 1507 -1898 1508 -1874
rect 1514 -1875 1515 -1781
rect 534 -1877 535 -1781
rect 989 -1898 990 -1876
rect 1472 -1877 1473 -1781
rect 1514 -1898 1515 -1876
rect 534 -1898 535 -1878
rect 758 -1879 759 -1781
rect 786 -1898 787 -1878
rect 849 -1879 850 -1781
rect 1472 -1898 1473 -1878
rect 1675 -1879 1676 -1781
rect 674 -1881 675 -1781
rect 849 -1898 850 -1880
rect 1675 -1898 1676 -1880
rect 1724 -1881 1725 -1781
rect 418 -1883 419 -1781
rect 1724 -1898 1725 -1882
rect 674 -1898 675 -1884
rect 709 -1885 710 -1781
rect 737 -1885 738 -1781
rect 1332 -1898 1333 -1884
rect 565 -1887 566 -1781
rect 709 -1898 710 -1886
rect 758 -1898 759 -1886
rect 821 -1887 822 -1781
rect 646 -1889 647 -1781
rect 737 -1898 738 -1888
rect 821 -1898 822 -1888
rect 835 -1889 836 -1781
rect 569 -1891 570 -1781
rect 646 -1898 647 -1890
rect 800 -1891 801 -1781
rect 835 -1898 836 -1890
rect 471 -1893 472 -1781
rect 569 -1898 570 -1892
rect 716 -1893 717 -1781
rect 800 -1898 801 -1892
rect 471 -1898 472 -1894
rect 1948 -1895 1949 -1781
rect 716 -1898 717 -1896
rect 926 -1898 927 -1896
rect 1563 -1898 1564 -1896
rect 1948 -1898 1949 -1896
rect 2 -2045 3 -1907
rect 226 -1908 227 -1906
rect 313 -2045 314 -1907
rect 450 -1908 451 -1906
rect 478 -2045 479 -1907
rect 555 -1908 556 -1906
rect 562 -1908 563 -1906
rect 576 -2045 577 -1907
rect 614 -1908 615 -1906
rect 989 -1908 990 -1906
rect 1024 -1908 1025 -1906
rect 1381 -1908 1382 -1906
rect 1430 -1908 1431 -1906
rect 1430 -2045 1431 -1907
rect 1430 -1908 1431 -1906
rect 1430 -2045 1431 -1907
rect 1454 -2045 1455 -1907
rect 1871 -1908 1872 -1906
rect 5 -1910 6 -1906
rect 68 -2045 69 -1909
rect 79 -1910 80 -1906
rect 509 -1910 510 -1906
rect 537 -2045 538 -1909
rect 1115 -1910 1116 -1906
rect 1153 -1910 1154 -1906
rect 1808 -1910 1809 -1906
rect 1871 -2045 1872 -1909
rect 1899 -1910 1900 -1906
rect 9 -2045 10 -1911
rect 37 -1912 38 -1906
rect 44 -1912 45 -1906
rect 138 -1912 139 -1906
rect 142 -1912 143 -1906
rect 1444 -1912 1445 -1906
rect 1458 -1912 1459 -1906
rect 1458 -2045 1459 -1911
rect 1458 -1912 1459 -1906
rect 1458 -2045 1459 -1911
rect 1535 -1912 1536 -1906
rect 1808 -2045 1809 -1911
rect 1899 -2045 1900 -1911
rect 1948 -1912 1949 -1906
rect 37 -2045 38 -1913
rect 541 -1914 542 -1906
rect 555 -2045 556 -1913
rect 737 -1914 738 -1906
rect 744 -1914 745 -1906
rect 1101 -2045 1102 -1913
rect 1108 -1914 1109 -1906
rect 1297 -1914 1298 -1906
rect 1367 -1914 1368 -1906
rect 1381 -2045 1382 -1913
rect 1444 -2045 1445 -1913
rect 1451 -1914 1452 -1906
rect 1535 -2045 1536 -1913
rect 2011 -1914 2012 -1906
rect 44 -2045 45 -1915
rect 289 -1916 290 -1906
rect 317 -1916 318 -1906
rect 744 -2045 745 -1915
rect 828 -1916 829 -1906
rect 933 -1916 934 -1906
rect 947 -1916 948 -1906
rect 947 -2045 948 -1915
rect 947 -1916 948 -1906
rect 947 -2045 948 -1915
rect 964 -2045 965 -1915
rect 1311 -1916 1312 -1906
rect 1451 -2045 1452 -1915
rect 1528 -1916 1529 -1906
rect 1563 -2045 1564 -1915
rect 1570 -1916 1571 -1906
rect 1745 -1916 1746 -1906
rect 1745 -2045 1746 -1915
rect 1745 -1916 1746 -1906
rect 1745 -2045 1746 -1915
rect 1948 -2045 1949 -1915
rect 1976 -1916 1977 -1906
rect 58 -2045 59 -1917
rect 695 -1918 696 -1906
rect 716 -1918 717 -1906
rect 737 -2045 738 -1917
rect 772 -1918 773 -1906
rect 1570 -2045 1571 -1917
rect 1976 -2045 1977 -1917
rect 2018 -1918 2019 -1906
rect 79 -2045 80 -1919
rect 471 -1920 472 -1906
rect 481 -1920 482 -1906
rect 1241 -1920 1242 -1906
rect 1283 -1920 1284 -1906
rect 1311 -2045 1312 -1919
rect 1528 -2045 1529 -1919
rect 1752 -1920 1753 -1906
rect 23 -1922 24 -1906
rect 471 -2045 472 -1921
rect 485 -1922 486 -1906
rect 908 -1922 909 -1906
rect 919 -1922 920 -1906
rect 933 -2045 934 -1921
rect 982 -1922 983 -1906
rect 1633 -1922 1634 -1906
rect 23 -2045 24 -1923
rect 114 -1924 115 -1906
rect 128 -1924 129 -1906
rect 128 -2045 129 -1923
rect 128 -1924 129 -1906
rect 128 -2045 129 -1923
rect 135 -1924 136 -1906
rect 726 -1924 727 -1906
rect 730 -1924 731 -1906
rect 894 -2045 895 -1923
rect 905 -1924 906 -1906
rect 1815 -1924 1816 -1906
rect 86 -1926 87 -1906
rect 289 -2045 290 -1925
rect 317 -2045 318 -1925
rect 758 -1926 759 -1906
rect 779 -1926 780 -1906
rect 905 -2045 906 -1925
rect 982 -2045 983 -1925
rect 1136 -1926 1137 -1906
rect 1143 -1926 1144 -1906
rect 1241 -2045 1242 -1925
rect 1293 -2045 1294 -1925
rect 1843 -1926 1844 -1906
rect 100 -1928 101 -1906
rect 268 -1928 269 -1906
rect 338 -1928 339 -1906
rect 828 -2045 829 -1927
rect 845 -2045 846 -1927
rect 1157 -1928 1158 -1906
rect 1199 -1928 1200 -1906
rect 1367 -2045 1368 -1927
rect 1566 -1928 1567 -1906
rect 1584 -1928 1585 -1906
rect 1633 -2045 1634 -1927
rect 1654 -1928 1655 -1906
rect 1815 -2045 1816 -1927
rect 1822 -1928 1823 -1906
rect 1843 -2045 1844 -1927
rect 1885 -1928 1886 -1906
rect 100 -2045 101 -1929
rect 527 -1930 528 -1906
rect 562 -2045 563 -1929
rect 583 -1930 584 -1906
rect 632 -1930 633 -1906
rect 768 -1930 769 -1906
rect 779 -2045 780 -1929
rect 856 -1930 857 -1906
rect 880 -2045 881 -1929
rect 1038 -1930 1039 -1906
rect 1090 -1930 1091 -1906
rect 1990 -1930 1991 -1906
rect 30 -1932 31 -1906
rect 527 -2045 528 -1931
rect 583 -2045 584 -1931
rect 597 -1932 598 -1906
rect 660 -1932 661 -1906
rect 663 -1960 664 -1931
rect 688 -1932 689 -1906
rect 1395 -1932 1396 -1906
rect 1472 -1932 1473 -1906
rect 1654 -2045 1655 -1931
rect 1822 -2045 1823 -1931
rect 1836 -1932 1837 -1906
rect 1885 -2045 1886 -1931
rect 1927 -1932 1928 -1906
rect 1990 -2045 1991 -1931
rect 2025 -1932 2026 -1906
rect 30 -2045 31 -1933
rect 513 -1934 514 -1906
rect 660 -2045 661 -1933
rect 681 -1934 682 -1906
rect 688 -2045 689 -1933
rect 698 -2045 699 -1933
rect 1283 -2045 1284 -1933
rect 1297 -2045 1298 -1933
rect 1493 -1934 1494 -1906
rect 1584 -2045 1585 -1933
rect 1605 -1934 1606 -1906
rect 1836 -2045 1837 -1933
rect 1850 -1934 1851 -1906
rect 1927 -2045 1928 -1933
rect 1955 -1934 1956 -1906
rect 16 -1936 17 -1906
rect 513 -2045 514 -1935
rect 674 -1936 675 -1906
rect 681 -2045 682 -1935
rect 709 -1936 710 -1906
rect 716 -2045 717 -1935
rect 719 -1936 720 -1906
rect 814 -1936 815 -1906
rect 856 -2045 857 -1935
rect 1080 -1936 1081 -1906
rect 1094 -1936 1095 -1906
rect 1115 -2045 1116 -1935
rect 1129 -1936 1130 -1906
rect 1143 -2045 1144 -1935
rect 1157 -2045 1158 -1935
rect 1171 -1936 1172 -1906
rect 1206 -1936 1207 -1906
rect 1216 -1936 1217 -1906
rect 1220 -1936 1221 -1906
rect 1731 -1936 1732 -1906
rect 1955 -2045 1956 -1935
rect 1983 -1936 1984 -1906
rect 65 -1938 66 -1906
rect 632 -2045 633 -1937
rect 674 -2045 675 -1937
rect 702 -1938 703 -1906
rect 709 -2045 710 -1937
rect 1059 -1938 1060 -1906
rect 1066 -1938 1067 -1906
rect 1080 -2045 1081 -1937
rect 1094 -2045 1095 -1937
rect 1318 -1938 1319 -1906
rect 1395 -2045 1396 -1937
rect 1500 -1938 1501 -1906
rect 1661 -1938 1662 -1906
rect 1850 -2045 1851 -1937
rect 103 -1940 104 -1906
rect 975 -1940 976 -1906
rect 989 -2045 990 -1939
rect 1031 -1940 1032 -1906
rect 1052 -1940 1053 -1906
rect 1059 -2045 1060 -1939
rect 1108 -2045 1109 -1939
rect 1514 -1940 1515 -1906
rect 16 -2045 17 -1941
rect 1031 -2045 1032 -1941
rect 1136 -2045 1137 -1941
rect 1178 -1942 1179 -1906
rect 1206 -2045 1207 -1941
rect 1521 -1942 1522 -1906
rect 107 -1944 108 -1906
rect 114 -2045 115 -1943
rect 135 -2045 136 -1943
rect 387 -1944 388 -1906
rect 401 -2045 402 -1943
rect 1209 -1944 1210 -1906
rect 1213 -1944 1214 -1906
rect 1213 -2045 1214 -1943
rect 1213 -1944 1214 -1906
rect 1213 -2045 1214 -1943
rect 1220 -2045 1221 -1943
rect 1416 -1944 1417 -1906
rect 1472 -2045 1473 -1943
rect 1542 -1944 1543 -1906
rect 93 -1946 94 -1906
rect 387 -2045 388 -1945
rect 415 -1946 416 -1906
rect 541 -2045 542 -1945
rect 639 -1946 640 -1906
rect 702 -2045 703 -1945
rect 730 -2045 731 -1945
rect 1878 -1946 1879 -1906
rect 51 -1948 52 -1906
rect 93 -2045 94 -1947
rect 107 -2045 108 -1947
rect 985 -1948 986 -1906
rect 1003 -1948 1004 -1906
rect 1066 -2045 1067 -1947
rect 1164 -1948 1165 -1906
rect 1199 -2045 1200 -1947
rect 1223 -1948 1224 -1906
rect 1920 -1948 1921 -1906
rect 51 -2045 52 -1949
rect 691 -1950 692 -1906
rect 733 -2045 734 -1949
rect 1752 -2045 1753 -1949
rect 1878 -2045 1879 -1949
rect 1906 -1950 1907 -1906
rect 1920 -2045 1921 -1949
rect 1997 -1950 1998 -1906
rect 142 -2045 143 -1951
rect 1829 -1952 1830 -1906
rect 1906 -2045 1907 -1951
rect 1934 -1952 1935 -1906
rect 145 -1954 146 -1906
rect 240 -1954 241 -1906
rect 408 -1954 409 -1906
rect 415 -2045 416 -1953
rect 464 -1954 465 -1906
rect 639 -2045 640 -1953
rect 758 -2045 759 -1953
rect 961 -1954 962 -1906
rect 1010 -1954 1011 -1906
rect 1024 -2045 1025 -1953
rect 1027 -1954 1028 -1906
rect 1801 -1954 1802 -1906
rect 1934 -2045 1935 -1953
rect 1962 -1954 1963 -1906
rect 86 -2045 87 -1955
rect 145 -2045 146 -1955
rect 156 -1956 157 -1906
rect 156 -2045 157 -1955
rect 156 -1956 157 -1906
rect 156 -2045 157 -1955
rect 198 -1956 199 -1906
rect 261 -1956 262 -1906
rect 408 -2045 409 -1955
rect 751 -1956 752 -1906
rect 800 -1956 801 -1906
rect 1052 -2045 1053 -1955
rect 1164 -2045 1165 -1955
rect 1248 -1956 1249 -1906
rect 1262 -1956 1263 -1906
rect 1500 -2045 1501 -1955
rect 1521 -2045 1522 -1955
rect 1549 -1956 1550 -1906
rect 1787 -1956 1788 -1906
rect 1829 -2045 1830 -1955
rect 170 -1958 171 -1906
rect 261 -2045 262 -1957
rect 464 -2045 465 -1957
rect 775 -1958 776 -1906
rect 807 -1958 808 -1906
rect 1038 -2045 1039 -1957
rect 1171 -2045 1172 -1957
rect 1255 -1958 1256 -1906
rect 1265 -2045 1266 -1957
rect 1731 -2045 1732 -1957
rect 1794 -1958 1795 -1906
rect 1801 -2045 1802 -1957
rect 170 -2045 171 -1959
rect 775 -2045 776 -1959
rect 807 -2045 808 -1959
rect 835 -1960 836 -1906
rect 849 -1960 850 -1906
rect 1129 -2045 1130 -1959
rect 1178 -2045 1179 -1959
rect 1185 -1960 1186 -1906
rect 1216 -2045 1217 -1959
rect 1549 -2045 1550 -1959
rect 1598 -1960 1599 -1906
rect 1794 -2045 1795 -1959
rect 198 -2045 199 -1961
rect 1262 -2045 1263 -1961
rect 1290 -1962 1291 -1906
rect 1318 -2045 1319 -1961
rect 1416 -2045 1417 -1961
rect 1423 -1962 1424 -1906
rect 1479 -1962 1480 -1906
rect 1514 -2045 1515 -1961
rect 1542 -2045 1543 -1961
rect 1556 -1962 1557 -1906
rect 212 -1964 213 -1906
rect 243 -2045 244 -1963
rect 268 -2045 269 -1963
rect 1290 -2045 1291 -1963
rect 1409 -1964 1410 -1906
rect 1423 -2045 1424 -1963
rect 1465 -1964 1466 -1906
rect 1556 -2045 1557 -1963
rect 184 -1966 185 -1906
rect 212 -2045 213 -1965
rect 226 -2045 227 -1965
rect 303 -1966 304 -1906
rect 485 -2045 486 -1965
rect 653 -1966 654 -1906
rect 814 -2045 815 -1965
rect 1332 -1966 1333 -1906
rect 1388 -1966 1389 -1906
rect 1409 -2045 1410 -1965
rect 1486 -1966 1487 -1906
rect 1493 -2045 1494 -1965
rect 1507 -1966 1508 -1906
rect 1598 -2045 1599 -1965
rect 184 -2045 185 -1967
rect 191 -1968 192 -1906
rect 205 -1968 206 -1906
rect 303 -2045 304 -1967
rect 457 -1968 458 -1906
rect 653 -2045 654 -1967
rect 821 -1968 822 -1906
rect 835 -2045 836 -1967
rect 849 -2045 850 -1967
rect 1073 -1968 1074 -1906
rect 1087 -1968 1088 -1906
rect 1465 -2045 1466 -1967
rect 1486 -2045 1487 -1967
rect 1647 -1968 1648 -1906
rect 163 -1970 164 -1906
rect 191 -2045 192 -1969
rect 205 -2045 206 -1969
rect 579 -1970 580 -1906
rect 618 -1970 619 -1906
rect 751 -2045 752 -1969
rect 793 -1970 794 -1906
rect 1073 -2045 1074 -1969
rect 1087 -2045 1088 -1969
rect 1353 -1970 1354 -1906
rect 1360 -1970 1361 -1906
rect 1507 -2045 1508 -1969
rect 1647 -2045 1648 -1969
rect 1689 -1970 1690 -1906
rect 72 -1972 73 -1906
rect 163 -2045 164 -1971
rect 341 -2045 342 -1971
rect 618 -2045 619 -1971
rect 793 -2045 794 -1971
rect 954 -1972 955 -1906
rect 961 -2045 962 -1971
rect 1787 -2045 1788 -1971
rect 61 -1974 62 -1906
rect 72 -2045 73 -1973
rect 380 -1974 381 -1906
rect 457 -2045 458 -1973
rect 499 -1974 500 -1906
rect 597 -2045 598 -1973
rect 821 -2045 822 -1973
rect 1192 -1974 1193 -1906
rect 1227 -1974 1228 -1906
rect 1227 -2045 1228 -1973
rect 1227 -1974 1228 -1906
rect 1227 -2045 1228 -1973
rect 1237 -2045 1238 -1973
rect 1279 -1974 1280 -1906
rect 1325 -1974 1326 -1906
rect 1332 -2045 1333 -1973
rect 1374 -1974 1375 -1906
rect 1388 -2045 1389 -1973
rect 1689 -2045 1690 -1973
rect 1759 -1974 1760 -1906
rect 380 -2045 381 -1975
rect 436 -1976 437 -1906
rect 443 -1976 444 -1906
rect 499 -2045 500 -1975
rect 506 -1976 507 -1906
rect 1248 -2045 1249 -1975
rect 1269 -1976 1270 -1906
rect 1360 -2045 1361 -1975
rect 247 -1978 248 -1906
rect 436 -2045 437 -1977
rect 754 -2045 755 -1977
rect 1269 -2045 1270 -1977
rect 1276 -1978 1277 -1906
rect 1479 -2045 1480 -1977
rect 177 -1980 178 -1906
rect 1276 -2045 1277 -1979
rect 1304 -1980 1305 -1906
rect 1325 -2045 1326 -1979
rect 1339 -1980 1340 -1906
rect 1374 -2045 1375 -1979
rect 177 -2045 178 -1981
rect 366 -1982 367 -1906
rect 863 -1982 864 -1906
rect 1003 -2045 1004 -1981
rect 1150 -1982 1151 -1906
rect 1759 -2045 1760 -1981
rect 247 -2045 248 -1983
rect 324 -1984 325 -1906
rect 352 -1984 353 -1906
rect 443 -2045 444 -1983
rect 611 -1984 612 -1906
rect 1150 -2045 1151 -1983
rect 1192 -2045 1193 -1983
rect 1913 -1984 1914 -1906
rect 254 -1986 255 -1906
rect 366 -2045 367 -1985
rect 611 -2045 612 -1985
rect 817 -2045 818 -1985
rect 863 -2045 864 -1985
rect 2004 -1986 2005 -1906
rect 254 -2045 255 -1987
rect 310 -1988 311 -1906
rect 324 -2045 325 -1987
rect 422 -1988 423 -1906
rect 866 -2045 867 -1987
rect 1962 -2045 1963 -1987
rect 275 -1990 276 -1906
rect 506 -2045 507 -1989
rect 877 -1990 878 -1906
rect 975 -2045 976 -1989
rect 996 -1990 997 -1906
rect 1010 -2045 1011 -1989
rect 1255 -2045 1256 -1989
rect 1913 -2045 1914 -1989
rect 275 -2045 276 -1991
rect 870 -1992 871 -1906
rect 877 -2045 878 -1991
rect 1577 -1992 1578 -1906
rect 296 -1994 297 -1906
rect 310 -2045 311 -1993
rect 345 -1994 346 -1906
rect 422 -2045 423 -1993
rect 842 -1994 843 -1906
rect 870 -2045 871 -1993
rect 884 -1994 885 -1906
rect 1612 -1994 1613 -1906
rect 121 -1996 122 -1906
rect 296 -2045 297 -1995
rect 345 -2045 346 -1995
rect 488 -1996 489 -1906
rect 604 -1996 605 -1906
rect 884 -2045 885 -1995
rect 887 -1996 888 -1906
rect 1983 -2045 1984 -1995
rect 121 -2045 122 -1997
rect 429 -1998 430 -1906
rect 604 -2045 605 -1997
rect 1045 -1998 1046 -1906
rect 1339 -2045 1340 -1997
rect 1346 -1998 1347 -1906
rect 1577 -2045 1578 -1997
rect 1591 -1998 1592 -1906
rect 1612 -2045 1613 -1997
rect 1675 -1998 1676 -1906
rect 219 -2000 220 -1906
rect 429 -2045 430 -1999
rect 842 -2045 843 -1999
rect 1710 -2000 1711 -1906
rect 219 -2045 220 -2001
rect 534 -2002 535 -1906
rect 912 -2002 913 -1906
rect 954 -2045 955 -2001
rect 968 -2002 969 -1906
rect 996 -2045 997 -2001
rect 1017 -2002 1018 -1906
rect 1045 -2045 1046 -2001
rect 1111 -2002 1112 -1906
rect 1710 -2045 1711 -2001
rect 352 -2045 353 -2003
rect 569 -2004 570 -1906
rect 800 -2045 801 -2003
rect 968 -2045 969 -2003
rect 1017 -2045 1018 -2003
rect 1437 -2004 1438 -1906
rect 1591 -2045 1592 -2003
rect 1668 -2004 1669 -1906
rect 1675 -2045 1676 -2003
rect 1703 -2004 1704 -1906
rect 492 -2006 493 -1906
rect 569 -2045 570 -2005
rect 912 -2045 913 -2005
rect 936 -2006 937 -1906
rect 1111 -2045 1112 -2005
rect 1353 -2045 1354 -2005
rect 1402 -2006 1403 -1906
rect 1437 -2045 1438 -2005
rect 1668 -2045 1669 -2005
rect 1696 -2006 1697 -1906
rect 1703 -2045 1704 -2005
rect 1738 -2006 1739 -1906
rect 359 -2008 360 -1906
rect 492 -2045 493 -2007
rect 520 -2008 521 -1906
rect 534 -2045 535 -2007
rect 723 -2008 724 -1906
rect 1402 -2045 1403 -2007
rect 1640 -2008 1641 -1906
rect 1696 -2045 1697 -2007
rect 331 -2010 332 -1906
rect 359 -2045 360 -2009
rect 394 -2010 395 -1906
rect 520 -2045 521 -2009
rect 530 -2045 531 -2009
rect 1738 -2045 1739 -2009
rect 149 -2012 150 -1906
rect 331 -2045 332 -2011
rect 723 -2045 724 -2011
rect 1661 -2045 1662 -2011
rect 149 -2045 150 -2013
rect 222 -2045 223 -2013
rect 233 -2014 234 -1906
rect 394 -2045 395 -2013
rect 919 -2045 920 -2013
rect 1304 -2045 1305 -2013
rect 1640 -2045 1641 -2013
rect 1682 -2014 1683 -1906
rect 233 -2045 234 -2015
rect 282 -2016 283 -1906
rect 922 -2045 923 -2015
rect 1605 -2045 1606 -2015
rect 1682 -2045 1683 -2015
rect 1724 -2016 1725 -1906
rect 282 -2045 283 -2017
rect 373 -2018 374 -1906
rect 926 -2018 927 -1906
rect 1185 -2045 1186 -2017
rect 1234 -2018 1235 -1906
rect 1346 -2045 1347 -2017
rect 1724 -2045 1725 -2017
rect 1766 -2018 1767 -1906
rect 373 -2045 374 -2019
rect 1122 -2020 1123 -1906
rect 1766 -2045 1767 -2019
rect 1773 -2020 1774 -1906
rect 898 -2022 899 -1906
rect 926 -2045 927 -2021
rect 940 -2022 941 -1906
rect 1122 -2045 1123 -2021
rect 1773 -2045 1774 -2021
rect 1780 -2022 1781 -1906
rect 625 -2024 626 -1906
rect 940 -2045 941 -2023
rect 1619 -2024 1620 -1906
rect 1780 -2045 1781 -2023
rect 548 -2026 549 -1906
rect 625 -2045 626 -2025
rect 786 -2026 787 -1906
rect 898 -2045 899 -2025
rect 1619 -2045 1620 -2025
rect 1717 -2026 1718 -1906
rect 548 -2045 549 -2027
rect 646 -2028 647 -1906
rect 772 -2045 773 -2027
rect 786 -2045 787 -2027
rect 1626 -2028 1627 -1906
rect 1717 -2045 1718 -2027
rect 590 -2030 591 -1906
rect 646 -2045 647 -2029
rect 1626 -2045 1627 -2029
rect 1864 -2030 1865 -1906
rect 590 -2045 591 -2031
rect 765 -2032 766 -1906
rect 1104 -2032 1105 -1906
rect 1864 -2045 1865 -2031
rect 765 -2045 766 -2033
rect 891 -2034 892 -1906
rect 891 -2045 892 -2035
rect 1857 -2036 1858 -1906
rect 1857 -2045 1858 -2037
rect 1892 -2038 1893 -1906
rect 1892 -2045 1893 -2039
rect 1941 -2040 1942 -1906
rect 1941 -2045 1942 -2041
rect 1969 -2042 1970 -1906
rect 761 -2045 762 -2043
rect 1969 -2045 1970 -2043
rect 2 -2055 3 -2053
rect 338 -2055 339 -2053
rect 352 -2055 353 -2053
rect 726 -2055 727 -2053
rect 733 -2055 734 -2053
rect 1101 -2055 1102 -2053
rect 1108 -2055 1109 -2053
rect 1514 -2055 1515 -2053
rect 1920 -2055 1921 -2053
rect 1976 -2055 1977 -2053
rect 2 -2186 3 -2056
rect 205 -2057 206 -2053
rect 219 -2057 220 -2053
rect 537 -2057 538 -2053
rect 548 -2057 549 -2053
rect 814 -2057 815 -2053
rect 817 -2057 818 -2053
rect 982 -2057 983 -2053
rect 1087 -2057 1088 -2053
rect 1234 -2186 1235 -2056
rect 1237 -2057 1238 -2053
rect 1493 -2057 1494 -2053
rect 23 -2059 24 -2053
rect 142 -2059 143 -2053
rect 149 -2059 150 -2053
rect 219 -2186 220 -2058
rect 222 -2059 223 -2053
rect 702 -2059 703 -2053
rect 723 -2059 724 -2053
rect 926 -2059 927 -2053
rect 947 -2059 948 -2053
rect 947 -2186 948 -2058
rect 947 -2059 948 -2053
rect 947 -2186 948 -2058
rect 961 -2059 962 -2053
rect 1500 -2059 1501 -2053
rect 9 -2061 10 -2053
rect 142 -2186 143 -2060
rect 177 -2061 178 -2053
rect 240 -2186 241 -2060
rect 352 -2186 353 -2060
rect 394 -2061 395 -2053
rect 401 -2061 402 -2053
rect 702 -2186 703 -2060
rect 723 -2186 724 -2060
rect 996 -2061 997 -2053
rect 1087 -2186 1088 -2060
rect 1185 -2061 1186 -2053
rect 1241 -2061 1242 -2053
rect 1262 -2061 1263 -2053
rect 1265 -2061 1266 -2053
rect 1850 -2061 1851 -2053
rect 23 -2186 24 -2062
rect 110 -2186 111 -2062
rect 117 -2063 118 -2053
rect 1507 -2063 1508 -2053
rect 1850 -2186 1851 -2062
rect 1927 -2063 1928 -2053
rect 30 -2065 31 -2053
rect 313 -2065 314 -2053
rect 394 -2186 395 -2064
rect 709 -2065 710 -2053
rect 751 -2065 752 -2053
rect 1129 -2065 1130 -2053
rect 1139 -2186 1140 -2064
rect 1437 -2065 1438 -2053
rect 1493 -2186 1494 -2064
rect 1605 -2065 1606 -2053
rect 30 -2186 31 -2066
rect 509 -2186 510 -2066
rect 520 -2067 521 -2053
rect 649 -2186 650 -2066
rect 695 -2067 696 -2053
rect 1038 -2067 1039 -2053
rect 1101 -2186 1102 -2066
rect 1178 -2067 1179 -2053
rect 1241 -2186 1242 -2066
rect 1304 -2067 1305 -2053
rect 1360 -2067 1361 -2053
rect 1454 -2186 1455 -2066
rect 1500 -2186 1501 -2066
rect 1759 -2067 1760 -2053
rect 37 -2069 38 -2053
rect 439 -2186 440 -2068
rect 450 -2069 451 -2053
rect 499 -2069 500 -2053
rect 530 -2069 531 -2053
rect 1402 -2069 1403 -2053
rect 1437 -2186 1438 -2068
rect 1472 -2069 1473 -2053
rect 1507 -2186 1508 -2068
rect 1710 -2069 1711 -2053
rect 1759 -2186 1760 -2068
rect 1857 -2069 1858 -2053
rect 51 -2071 52 -2053
rect 698 -2071 699 -2053
rect 751 -2186 752 -2070
rect 1108 -2186 1109 -2070
rect 1129 -2186 1130 -2070
rect 1136 -2071 1137 -2053
rect 1143 -2071 1144 -2053
rect 1262 -2186 1263 -2070
rect 1290 -2186 1291 -2070
rect 1353 -2071 1354 -2053
rect 1363 -2186 1364 -2070
rect 1829 -2071 1830 -2053
rect 1857 -2186 1858 -2070
rect 1941 -2071 1942 -2053
rect 51 -2186 52 -2072
rect 261 -2073 262 -2053
rect 303 -2073 304 -2053
rect 401 -2186 402 -2072
rect 408 -2073 409 -2053
rect 838 -2186 839 -2072
rect 845 -2073 846 -2053
rect 1514 -2186 1515 -2072
rect 1605 -2186 1606 -2072
rect 1773 -2073 1774 -2053
rect 1829 -2186 1830 -2072
rect 1899 -2073 1900 -2053
rect 65 -2075 66 -2053
rect 1402 -2186 1403 -2074
rect 1710 -2186 1711 -2074
rect 1836 -2075 1837 -2053
rect 1899 -2186 1900 -2074
rect 1990 -2075 1991 -2053
rect 65 -2186 66 -2076
rect 380 -2077 381 -2053
rect 415 -2077 416 -2053
rect 730 -2077 731 -2053
rect 761 -2077 762 -2053
rect 786 -2077 787 -2053
rect 807 -2077 808 -2053
rect 814 -2186 815 -2076
rect 891 -2077 892 -2053
rect 1031 -2077 1032 -2053
rect 1038 -2186 1039 -2076
rect 1052 -2077 1053 -2053
rect 1143 -2186 1144 -2076
rect 1213 -2077 1214 -2053
rect 1255 -2077 1256 -2053
rect 1311 -2077 1312 -2053
rect 1353 -2186 1354 -2076
rect 1570 -2077 1571 -2053
rect 1773 -2186 1774 -2076
rect 1843 -2077 1844 -2053
rect 44 -2079 45 -2053
rect 380 -2186 381 -2078
rect 422 -2079 423 -2053
rect 450 -2186 451 -2078
rect 492 -2079 493 -2053
rect 499 -2186 500 -2078
rect 548 -2186 549 -2078
rect 562 -2079 563 -2053
rect 583 -2079 584 -2053
rect 807 -2186 808 -2078
rect 919 -2079 920 -2053
rect 1598 -2079 1599 -2053
rect 1843 -2186 1844 -2078
rect 1913 -2079 1914 -2053
rect 44 -2186 45 -2080
rect 86 -2081 87 -2053
rect 89 -2186 90 -2080
rect 324 -2081 325 -2053
rect 422 -2186 423 -2080
rect 975 -2081 976 -2053
rect 978 -2186 979 -2080
rect 1374 -2081 1375 -2053
rect 1475 -2186 1476 -2080
rect 1836 -2186 1837 -2080
rect 68 -2083 69 -2053
rect 471 -2083 472 -2053
rect 492 -2186 493 -2082
rect 541 -2083 542 -2053
rect 562 -2186 563 -2082
rect 1111 -2083 1112 -2053
rect 1160 -2186 1161 -2082
rect 1304 -2186 1305 -2082
rect 1311 -2186 1312 -2082
rect 1388 -2083 1389 -2053
rect 1570 -2186 1571 -2082
rect 1661 -2083 1662 -2053
rect 1717 -2083 1718 -2053
rect 1913 -2186 1914 -2082
rect 79 -2085 80 -2053
rect 82 -2139 83 -2084
rect 86 -2186 87 -2084
rect 513 -2085 514 -2053
rect 583 -2186 584 -2084
rect 646 -2085 647 -2053
rect 695 -2186 696 -2084
rect 716 -2085 717 -2053
rect 730 -2186 731 -2084
rect 964 -2085 965 -2053
rect 968 -2085 969 -2053
rect 1479 -2085 1480 -2053
rect 1661 -2186 1662 -2084
rect 1724 -2085 1725 -2053
rect 79 -2186 80 -2086
rect 135 -2087 136 -2053
rect 163 -2087 164 -2053
rect 303 -2186 304 -2086
rect 436 -2087 437 -2053
rect 513 -2186 514 -2086
rect 590 -2087 591 -2053
rect 1398 -2186 1399 -2086
rect 1479 -2186 1480 -2086
rect 1584 -2087 1585 -2053
rect 1633 -2087 1634 -2053
rect 1724 -2186 1725 -2086
rect 93 -2089 94 -2053
rect 520 -2186 521 -2088
rect 593 -2186 594 -2088
rect 744 -2089 745 -2053
rect 772 -2089 773 -2053
rect 1066 -2089 1067 -2053
rect 1171 -2089 1172 -2053
rect 1185 -2186 1186 -2088
rect 1213 -2186 1214 -2088
rect 1339 -2089 1340 -2053
rect 1374 -2186 1375 -2088
rect 1906 -2089 1907 -2053
rect 33 -2186 34 -2090
rect 744 -2186 745 -2090
rect 772 -2186 773 -2090
rect 1111 -2186 1112 -2090
rect 1171 -2186 1172 -2090
rect 1346 -2091 1347 -2053
rect 1388 -2186 1389 -2090
rect 1458 -2091 1459 -2053
rect 1584 -2186 1585 -2090
rect 1668 -2091 1669 -2053
rect 1675 -2091 1676 -2053
rect 1906 -2186 1907 -2090
rect 93 -2186 94 -2092
rect 387 -2093 388 -2053
rect 467 -2186 468 -2092
rect 968 -2186 969 -2092
rect 971 -2093 972 -2053
rect 1423 -2093 1424 -2053
rect 1458 -2186 1459 -2092
rect 1542 -2093 1543 -2053
rect 1675 -2186 1676 -2092
rect 1731 -2093 1732 -2053
rect 96 -2186 97 -2094
rect 390 -2186 391 -2094
rect 597 -2095 598 -2053
rect 849 -2095 850 -2053
rect 852 -2095 853 -2053
rect 1633 -2186 1634 -2094
rect 1703 -2095 1704 -2053
rect 1731 -2186 1732 -2094
rect 16 -2097 17 -2053
rect 849 -2186 850 -2096
rect 905 -2097 906 -2053
rect 919 -2186 920 -2096
rect 922 -2097 923 -2053
rect 1122 -2097 1123 -2053
rect 1178 -2186 1179 -2096
rect 1416 -2097 1417 -2053
rect 1542 -2186 1543 -2096
rect 1619 -2097 1620 -2053
rect 1703 -2186 1704 -2096
rect 1794 -2097 1795 -2053
rect 16 -2186 17 -2098
rect 243 -2099 244 -2053
rect 247 -2099 248 -2053
rect 261 -2186 262 -2098
rect 268 -2099 269 -2053
rect 408 -2186 409 -2098
rect 506 -2099 507 -2053
rect 597 -2186 598 -2098
rect 604 -2099 605 -2053
rect 709 -2186 710 -2098
rect 779 -2099 780 -2053
rect 891 -2186 892 -2098
rect 926 -2186 927 -2098
rect 933 -2099 934 -2053
rect 954 -2099 955 -2053
rect 961 -2186 962 -2098
rect 975 -2186 976 -2098
rect 1010 -2099 1011 -2053
rect 1031 -2186 1032 -2098
rect 1206 -2099 1207 -2053
rect 1220 -2099 1221 -2053
rect 1339 -2186 1340 -2098
rect 1346 -2186 1347 -2098
rect 1923 -2099 1924 -2053
rect 128 -2101 129 -2053
rect 149 -2186 150 -2100
rect 163 -2186 164 -2100
rect 310 -2101 311 -2053
rect 324 -2186 325 -2100
rect 590 -2186 591 -2100
rect 618 -2101 619 -2053
rect 716 -2186 717 -2100
rect 786 -2186 787 -2100
rect 1164 -2101 1165 -2053
rect 1192 -2101 1193 -2053
rect 1206 -2186 1207 -2100
rect 1220 -2186 1221 -2100
rect 1283 -2101 1284 -2053
rect 1395 -2101 1396 -2053
rect 1423 -2186 1424 -2100
rect 1619 -2186 1620 -2100
rect 1766 -2101 1767 -2053
rect 1794 -2186 1795 -2100
rect 1815 -2101 1816 -2053
rect 107 -2103 108 -2053
rect 128 -2186 129 -2102
rect 135 -2186 136 -2102
rect 156 -2103 157 -2053
rect 177 -2186 178 -2102
rect 289 -2103 290 -2053
rect 341 -2186 342 -2102
rect 618 -2186 619 -2102
rect 639 -2103 640 -2053
rect 758 -2103 759 -2053
rect 884 -2103 885 -2053
rect 905 -2186 906 -2102
rect 933 -2186 934 -2102
rect 1017 -2103 1018 -2053
rect 1052 -2186 1053 -2102
rect 1696 -2103 1697 -2053
rect 1717 -2186 1718 -2102
rect 1745 -2103 1746 -2053
rect 1766 -2186 1767 -2102
rect 1822 -2103 1823 -2053
rect 156 -2186 157 -2104
rect 184 -2105 185 -2053
rect 191 -2105 192 -2053
rect 471 -2186 472 -2104
rect 506 -2186 507 -2104
rect 779 -2186 780 -2104
rect 870 -2105 871 -2053
rect 884 -2186 885 -2104
rect 954 -2186 955 -2104
rect 1297 -2105 1298 -2053
rect 1409 -2105 1410 -2053
rect 1668 -2186 1669 -2104
rect 1696 -2186 1697 -2104
rect 1969 -2105 1970 -2053
rect 184 -2186 185 -2106
rect 842 -2107 843 -2053
rect 982 -2186 983 -2106
rect 1003 -2107 1004 -2053
rect 1010 -2186 1011 -2106
rect 1059 -2107 1060 -2053
rect 1066 -2186 1067 -2106
rect 1745 -2186 1746 -2106
rect 1815 -2186 1816 -2106
rect 1892 -2107 1893 -2053
rect 191 -2186 192 -2108
rect 359 -2109 360 -2053
rect 485 -2109 486 -2053
rect 842 -2186 843 -2108
rect 989 -2109 990 -2053
rect 1017 -2186 1018 -2108
rect 1059 -2186 1060 -2108
rect 1157 -2109 1158 -2053
rect 1192 -2186 1193 -2108
rect 1325 -2109 1326 -2053
rect 1409 -2186 1410 -2108
rect 1465 -2109 1466 -2053
rect 1822 -2186 1823 -2108
rect 1948 -2109 1949 -2053
rect 198 -2111 199 -2053
rect 310 -2186 311 -2110
rect 485 -2186 486 -2110
rect 569 -2111 570 -2053
rect 576 -2111 577 -2053
rect 604 -2186 605 -2110
rect 611 -2111 612 -2053
rect 1164 -2186 1165 -2110
rect 1248 -2111 1249 -2053
rect 1416 -2186 1417 -2110
rect 1465 -2186 1466 -2110
rect 1577 -2111 1578 -2053
rect 1892 -2186 1893 -2110
rect 1983 -2111 1984 -2053
rect 198 -2186 199 -2112
rect 226 -2113 227 -2053
rect 236 -2186 237 -2112
rect 863 -2113 864 -2053
rect 989 -2186 990 -2112
rect 1045 -2113 1046 -2053
rect 1115 -2113 1116 -2053
rect 1122 -2186 1123 -2112
rect 1157 -2186 1158 -2112
rect 1878 -2113 1879 -2053
rect 205 -2186 206 -2114
rect 971 -2186 972 -2114
rect 996 -2186 997 -2114
rect 1024 -2115 1025 -2053
rect 1045 -2186 1046 -2114
rect 1377 -2186 1378 -2114
rect 1577 -2186 1578 -2114
rect 1808 -2115 1809 -2053
rect 226 -2186 227 -2116
rect 233 -2117 234 -2053
rect 247 -2186 248 -2116
rect 345 -2117 346 -2053
rect 527 -2117 528 -2053
rect 1283 -2186 1284 -2116
rect 1325 -2186 1326 -2116
rect 1381 -2117 1382 -2053
rect 1738 -2117 1739 -2053
rect 1878 -2186 1879 -2116
rect 212 -2119 213 -2053
rect 233 -2186 234 -2118
rect 268 -2186 269 -2118
rect 373 -2119 374 -2053
rect 527 -2186 528 -2118
rect 877 -2119 878 -2053
rect 1003 -2186 1004 -2118
rect 1073 -2119 1074 -2053
rect 1115 -2186 1116 -2118
rect 1199 -2119 1200 -2053
rect 1248 -2186 1249 -2118
rect 1367 -2119 1368 -2053
rect 1381 -2186 1382 -2118
rect 1591 -2119 1592 -2053
rect 1738 -2186 1739 -2118
rect 1801 -2119 1802 -2053
rect 1808 -2186 1809 -2118
rect 1934 -2119 1935 -2053
rect 145 -2121 146 -2053
rect 1367 -2186 1368 -2120
rect 1591 -2186 1592 -2120
rect 1682 -2121 1683 -2053
rect 1801 -2186 1802 -2120
rect 1885 -2121 1886 -2053
rect 170 -2123 171 -2053
rect 373 -2186 374 -2122
rect 415 -2186 416 -2122
rect 877 -2186 878 -2122
rect 1024 -2186 1025 -2122
rect 1521 -2123 1522 -2053
rect 1682 -2186 1683 -2122
rect 1752 -2123 1753 -2053
rect 1885 -2186 1886 -2122
rect 1962 -2123 1963 -2053
rect 40 -2186 41 -2124
rect 170 -2186 171 -2124
rect 212 -2186 213 -2124
rect 366 -2125 367 -2053
rect 576 -2186 577 -2124
rect 653 -2125 654 -2053
rect 737 -2125 738 -2053
rect 758 -2186 759 -2124
rect 863 -2186 864 -2124
rect 1069 -2186 1070 -2124
rect 1073 -2186 1074 -2124
rect 1080 -2125 1081 -2053
rect 1199 -2186 1200 -2124
rect 1276 -2125 1277 -2053
rect 1486 -2125 1487 -2053
rect 1521 -2186 1522 -2124
rect 1689 -2125 1690 -2053
rect 1752 -2186 1753 -2124
rect 114 -2127 115 -2053
rect 366 -2186 367 -2126
rect 611 -2186 612 -2126
rect 625 -2127 626 -2053
rect 628 -2186 629 -2126
rect 870 -2186 871 -2126
rect 894 -2127 895 -2053
rect 1276 -2186 1277 -2126
rect 1486 -2186 1487 -2126
rect 1549 -2127 1550 -2053
rect 1689 -2186 1690 -2126
rect 1787 -2127 1788 -2053
rect 282 -2129 283 -2053
rect 359 -2186 360 -2128
rect 625 -2186 626 -2128
rect 800 -2129 801 -2053
rect 1080 -2186 1081 -2128
rect 1780 -2129 1781 -2053
rect 1787 -2186 1788 -2128
rect 1871 -2129 1872 -2053
rect 100 -2131 101 -2053
rect 282 -2186 283 -2130
rect 289 -2186 290 -2130
rect 866 -2131 867 -2053
rect 1255 -2186 1256 -2130
rect 1360 -2186 1361 -2130
rect 1549 -2186 1550 -2130
rect 1556 -2131 1557 -2053
rect 1780 -2186 1781 -2130
rect 1864 -2131 1865 -2053
rect 1871 -2186 1872 -2130
rect 1955 -2131 1956 -2053
rect 100 -2186 101 -2132
rect 1451 -2133 1452 -2053
rect 1556 -2186 1557 -2132
rect 1647 -2133 1648 -2053
rect 296 -2135 297 -2053
rect 569 -2186 570 -2134
rect 639 -2186 640 -2134
rect 856 -2135 857 -2053
rect 1269 -2135 1270 -2053
rect 1297 -2186 1298 -2134
rect 1451 -2186 1452 -2134
rect 1598 -2186 1599 -2134
rect 1612 -2135 1613 -2053
rect 1647 -2186 1648 -2134
rect 254 -2137 255 -2053
rect 296 -2186 297 -2136
rect 317 -2137 318 -2053
rect 856 -2186 857 -2136
rect 1269 -2186 1270 -2136
rect 1332 -2137 1333 -2053
rect 254 -2186 255 -2138
rect 317 -2186 318 -2138
rect 331 -2139 332 -2053
rect 345 -2186 346 -2138
rect 443 -2139 444 -2053
rect 646 -2186 647 -2138
rect 1094 -2139 1095 -2053
rect 1293 -2139 1294 -2053
rect 1612 -2186 1613 -2138
rect 331 -2186 332 -2140
rect 478 -2141 479 -2053
rect 653 -2186 654 -2140
rect 674 -2141 675 -2053
rect 737 -2186 738 -2140
rect 793 -2141 794 -2053
rect 800 -2186 801 -2140
rect 821 -2141 822 -2053
rect 940 -2141 941 -2053
rect 1094 -2186 1095 -2140
rect 1332 -2186 1333 -2140
rect 1444 -2141 1445 -2053
rect 443 -2186 444 -2142
rect 765 -2143 766 -2053
rect 793 -2186 794 -2142
rect 898 -2143 899 -2053
rect 1444 -2186 1445 -2142
rect 1535 -2143 1536 -2053
rect 275 -2145 276 -2053
rect 898 -2186 899 -2144
rect 1430 -2145 1431 -2053
rect 1535 -2186 1536 -2144
rect 275 -2186 276 -2146
rect 828 -2147 829 -2053
rect 1430 -2186 1431 -2146
rect 1528 -2147 1529 -2053
rect 453 -2149 454 -2053
rect 828 -2186 829 -2148
rect 1528 -2186 1529 -2148
rect 1640 -2149 1641 -2053
rect 457 -2151 458 -2053
rect 478 -2186 479 -2150
rect 667 -2151 668 -2053
rect 940 -2186 941 -2150
rect 1626 -2151 1627 -2053
rect 1640 -2186 1641 -2150
rect 457 -2186 458 -2152
rect 660 -2153 661 -2053
rect 667 -2186 668 -2152
rect 688 -2153 689 -2053
rect 754 -2153 755 -2053
rect 1864 -2186 1865 -2152
rect 555 -2155 556 -2053
rect 688 -2186 689 -2154
rect 765 -2186 766 -2154
rect 1395 -2186 1396 -2154
rect 1563 -2155 1564 -2053
rect 1626 -2186 1627 -2154
rect 555 -2186 556 -2156
rect 632 -2157 633 -2053
rect 660 -2186 661 -2156
rect 1090 -2157 1091 -2053
rect 1563 -2186 1564 -2156
rect 1654 -2157 1655 -2053
rect 404 -2186 405 -2158
rect 1654 -2186 1655 -2158
rect 429 -2161 430 -2053
rect 632 -2186 633 -2160
rect 674 -2186 675 -2160
rect 681 -2161 682 -2053
rect 821 -2186 822 -2160
rect 835 -2161 836 -2053
rect 429 -2186 430 -2162
rect 436 -2186 437 -2162
rect 534 -2163 535 -2053
rect 835 -2186 836 -2162
rect 534 -2186 535 -2164
rect 880 -2165 881 -2053
rect 681 -2186 682 -2166
rect 1083 -2186 1084 -2166
rect 880 -2186 881 -2168
rect 1150 -2169 1151 -2053
rect 1150 -2186 1151 -2170
rect 1227 -2171 1228 -2053
rect 1227 -2186 1228 -2172
rect 1318 -2173 1319 -2053
rect 912 -2175 913 -2053
rect 1318 -2186 1319 -2174
rect 121 -2177 122 -2053
rect 912 -2186 913 -2176
rect 72 -2179 73 -2053
rect 121 -2186 122 -2178
rect 72 -2186 73 -2180
rect 464 -2181 465 -2053
rect 58 -2183 59 -2053
rect 464 -2186 465 -2182
rect 58 -2186 59 -2184
rect 387 -2186 388 -2184
rect 2 -2196 3 -2194
rect 40 -2196 41 -2194
rect 58 -2196 59 -2194
rect 215 -2315 216 -2195
rect 222 -2315 223 -2195
rect 1139 -2196 1140 -2194
rect 1178 -2196 1179 -2194
rect 1451 -2315 1452 -2195
rect 1454 -2196 1455 -2194
rect 1808 -2196 1809 -2194
rect 12 -2198 13 -2194
rect 16 -2198 17 -2194
rect 33 -2198 34 -2194
rect 520 -2198 521 -2194
rect 527 -2198 528 -2194
rect 761 -2315 762 -2197
rect 779 -2198 780 -2194
rect 779 -2315 780 -2197
rect 779 -2198 780 -2194
rect 779 -2315 780 -2197
rect 817 -2315 818 -2197
rect 1038 -2198 1039 -2194
rect 1055 -2198 1056 -2194
rect 1318 -2198 1319 -2194
rect 1360 -2198 1361 -2194
rect 1486 -2198 1487 -2194
rect 1713 -2315 1714 -2197
rect 1724 -2198 1725 -2194
rect 1727 -2315 1728 -2197
rect 1906 -2198 1907 -2194
rect 16 -2315 17 -2199
rect 303 -2200 304 -2194
rect 317 -2200 318 -2194
rect 341 -2200 342 -2194
rect 352 -2200 353 -2194
rect 625 -2315 626 -2199
rect 646 -2315 647 -2199
rect 891 -2200 892 -2194
rect 950 -2315 951 -2199
rect 1878 -2200 1879 -2194
rect 37 -2202 38 -2194
rect 849 -2202 850 -2194
rect 877 -2202 878 -2194
rect 1297 -2202 1298 -2194
rect 1318 -2315 1319 -2201
rect 1458 -2202 1459 -2194
rect 1475 -2202 1476 -2194
rect 1759 -2202 1760 -2194
rect 23 -2204 24 -2194
rect 37 -2315 38 -2203
rect 44 -2204 45 -2194
rect 58 -2315 59 -2203
rect 68 -2315 69 -2203
rect 296 -2204 297 -2194
rect 303 -2315 304 -2203
rect 562 -2204 563 -2194
rect 572 -2315 573 -2203
rect 884 -2204 885 -2194
rect 891 -2315 892 -2203
rect 1304 -2204 1305 -2194
rect 1395 -2204 1396 -2194
rect 1787 -2204 1788 -2194
rect 23 -2315 24 -2205
rect 191 -2206 192 -2194
rect 254 -2206 255 -2194
rect 1083 -2206 1084 -2194
rect 1108 -2206 1109 -2194
rect 1262 -2206 1263 -2194
rect 1276 -2206 1277 -2194
rect 1286 -2250 1287 -2205
rect 1304 -2315 1305 -2205
rect 1822 -2206 1823 -2194
rect 44 -2315 45 -2207
rect 128 -2208 129 -2194
rect 163 -2208 164 -2194
rect 1125 -2315 1126 -2207
rect 1136 -2315 1137 -2207
rect 1220 -2208 1221 -2194
rect 1248 -2208 1249 -2194
rect 1248 -2315 1249 -2207
rect 1248 -2208 1249 -2194
rect 1248 -2315 1249 -2207
rect 1255 -2208 1256 -2194
rect 1262 -2315 1263 -2207
rect 1276 -2315 1277 -2207
rect 1325 -2208 1326 -2194
rect 1395 -2315 1396 -2207
rect 1605 -2208 1606 -2194
rect 1717 -2208 1718 -2194
rect 1717 -2315 1718 -2207
rect 1717 -2208 1718 -2194
rect 1717 -2315 1718 -2207
rect 1787 -2315 1788 -2207
rect 1794 -2208 1795 -2194
rect 1822 -2315 1823 -2207
rect 1892 -2208 1893 -2194
rect 107 -2210 108 -2194
rect 275 -2210 276 -2194
rect 282 -2210 283 -2194
rect 338 -2315 339 -2209
rect 352 -2315 353 -2209
rect 597 -2210 598 -2194
rect 670 -2315 671 -2209
rect 1885 -2210 1886 -2194
rect 107 -2315 108 -2211
rect 814 -2212 815 -2194
rect 877 -2315 878 -2211
rect 919 -2212 920 -2194
rect 954 -2212 955 -2194
rect 1297 -2315 1298 -2211
rect 1325 -2315 1326 -2211
rect 1444 -2212 1445 -2194
rect 1458 -2315 1459 -2211
rect 1479 -2212 1480 -2194
rect 1605 -2315 1606 -2211
rect 1647 -2212 1648 -2194
rect 1794 -2315 1795 -2211
rect 1899 -2212 1900 -2194
rect 110 -2214 111 -2194
rect 324 -2214 325 -2194
rect 387 -2214 388 -2194
rect 478 -2214 479 -2194
rect 520 -2315 521 -2213
rect 716 -2214 717 -2194
rect 730 -2214 731 -2194
rect 730 -2315 731 -2213
rect 730 -2214 731 -2194
rect 730 -2315 731 -2213
rect 786 -2214 787 -2194
rect 1486 -2315 1487 -2213
rect 1640 -2214 1641 -2194
rect 1647 -2315 1648 -2213
rect 117 -2315 118 -2215
rect 149 -2216 150 -2194
rect 163 -2315 164 -2215
rect 247 -2216 248 -2194
rect 254 -2315 255 -2215
rect 331 -2216 332 -2194
rect 408 -2216 409 -2194
rect 478 -2315 479 -2215
rect 527 -2315 528 -2215
rect 611 -2216 612 -2194
rect 695 -2216 696 -2194
rect 695 -2315 696 -2215
rect 695 -2216 696 -2194
rect 695 -2315 696 -2215
rect 737 -2216 738 -2194
rect 786 -2315 787 -2215
rect 793 -2216 794 -2194
rect 849 -2315 850 -2215
rect 880 -2216 881 -2194
rect 1500 -2216 1501 -2194
rect 1640 -2315 1641 -2215
rect 1745 -2216 1746 -2194
rect 128 -2315 129 -2217
rect 135 -2218 136 -2194
rect 170 -2218 171 -2194
rect 387 -2315 388 -2217
rect 408 -2315 409 -2217
rect 485 -2218 486 -2194
rect 544 -2218 545 -2194
rect 912 -2218 913 -2194
rect 919 -2315 920 -2217
rect 947 -2218 948 -2194
rect 968 -2218 969 -2194
rect 1577 -2218 1578 -2194
rect 1745 -2315 1746 -2217
rect 1913 -2218 1914 -2194
rect 135 -2315 136 -2219
rect 184 -2220 185 -2194
rect 191 -2315 192 -2219
rect 975 -2220 976 -2194
rect 999 -2315 1000 -2219
rect 1535 -2220 1536 -2194
rect 170 -2315 171 -2221
rect 268 -2222 269 -2194
rect 289 -2222 290 -2194
rect 324 -2315 325 -2221
rect 331 -2315 332 -2221
rect 464 -2222 465 -2194
rect 471 -2222 472 -2194
rect 1080 -2315 1081 -2221
rect 1108 -2315 1109 -2221
rect 1283 -2222 1284 -2194
rect 1353 -2222 1354 -2194
rect 1577 -2315 1578 -2221
rect 79 -2224 80 -2194
rect 289 -2315 290 -2223
rect 296 -2315 297 -2223
rect 443 -2224 444 -2194
rect 457 -2224 458 -2194
rect 509 -2224 510 -2194
rect 562 -2315 563 -2223
rect 723 -2224 724 -2194
rect 737 -2315 738 -2223
rect 863 -2224 864 -2194
rect 912 -2315 913 -2223
rect 926 -2224 927 -2194
rect 968 -2315 969 -2223
rect 1003 -2224 1004 -2194
rect 1038 -2315 1039 -2223
rect 1101 -2224 1102 -2194
rect 1111 -2224 1112 -2194
rect 1626 -2224 1627 -2194
rect 51 -2226 52 -2194
rect 457 -2315 458 -2225
rect 485 -2315 486 -2225
rect 492 -2226 493 -2194
rect 569 -2226 570 -2194
rect 716 -2315 717 -2225
rect 796 -2315 797 -2225
rect 954 -2315 955 -2225
rect 971 -2226 972 -2194
rect 1094 -2226 1095 -2194
rect 1101 -2315 1102 -2225
rect 1150 -2226 1151 -2194
rect 1178 -2315 1179 -2225
rect 1339 -2226 1340 -2194
rect 1353 -2315 1354 -2225
rect 1416 -2226 1417 -2194
rect 1444 -2315 1445 -2225
rect 1493 -2226 1494 -2194
rect 1500 -2315 1501 -2225
rect 1591 -2226 1592 -2194
rect 1626 -2315 1627 -2225
rect 1738 -2226 1739 -2194
rect 30 -2228 31 -2194
rect 51 -2315 52 -2227
rect 79 -2315 80 -2227
rect 100 -2228 101 -2194
rect 142 -2228 143 -2194
rect 268 -2315 269 -2227
rect 380 -2228 381 -2194
rect 569 -2315 570 -2227
rect 590 -2228 591 -2194
rect 1241 -2228 1242 -2194
rect 1279 -2228 1280 -2194
rect 1549 -2228 1550 -2194
rect 1591 -2315 1592 -2227
rect 1675 -2228 1676 -2194
rect 1696 -2228 1697 -2194
rect 1738 -2315 1739 -2227
rect 30 -2315 31 -2229
rect 1024 -2230 1025 -2194
rect 1031 -2230 1032 -2194
rect 1339 -2315 1340 -2229
rect 1398 -2230 1399 -2194
rect 1871 -2230 1872 -2194
rect 65 -2232 66 -2194
rect 100 -2315 101 -2231
rect 177 -2232 178 -2194
rect 471 -2315 472 -2231
rect 576 -2232 577 -2194
rect 590 -2315 591 -2231
rect 597 -2315 598 -2231
rect 632 -2232 633 -2194
rect 639 -2232 640 -2194
rect 793 -2315 794 -2231
rect 926 -2315 927 -2231
rect 961 -2232 962 -2194
rect 989 -2232 990 -2194
rect 1003 -2315 1004 -2231
rect 1010 -2232 1011 -2194
rect 1031 -2315 1032 -2231
rect 1052 -2232 1053 -2194
rect 1360 -2315 1361 -2231
rect 1402 -2232 1403 -2194
rect 1619 -2232 1620 -2194
rect 1675 -2315 1676 -2231
rect 1829 -2232 1830 -2194
rect 86 -2234 87 -2194
rect 177 -2315 178 -2233
rect 184 -2315 185 -2233
rect 219 -2234 220 -2194
rect 226 -2234 227 -2194
rect 247 -2315 248 -2233
rect 261 -2234 262 -2194
rect 317 -2315 318 -2233
rect 415 -2234 416 -2194
rect 492 -2315 493 -2233
rect 506 -2234 507 -2194
rect 961 -2315 962 -2233
rect 989 -2315 990 -2233
rect 1017 -2234 1018 -2194
rect 1024 -2315 1025 -2233
rect 1059 -2234 1060 -2194
rect 1066 -2234 1067 -2194
rect 1185 -2234 1186 -2194
rect 1188 -2315 1189 -2233
rect 1332 -2234 1333 -2194
rect 1402 -2315 1403 -2233
rect 1430 -2234 1431 -2194
rect 1479 -2315 1480 -2233
rect 1563 -2234 1564 -2194
rect 1619 -2315 1620 -2233
rect 1703 -2234 1704 -2194
rect 1829 -2315 1830 -2233
rect 1850 -2234 1851 -2194
rect 86 -2315 87 -2235
rect 394 -2236 395 -2194
rect 415 -2315 416 -2235
rect 467 -2315 468 -2235
rect 506 -2315 507 -2235
rect 772 -2236 773 -2194
rect 800 -2236 801 -2194
rect 1059 -2315 1060 -2235
rect 1087 -2236 1088 -2194
rect 1150 -2315 1151 -2235
rect 1192 -2236 1193 -2194
rect 1241 -2315 1242 -2235
rect 1283 -2315 1284 -2235
rect 1388 -2236 1389 -2194
rect 1430 -2315 1431 -2235
rect 1514 -2236 1515 -2194
rect 1535 -2315 1536 -2235
rect 1689 -2236 1690 -2194
rect 1696 -2315 1697 -2235
rect 1815 -2236 1816 -2194
rect 173 -2315 174 -2237
rect 772 -2315 773 -2237
rect 1010 -2315 1011 -2237
rect 1164 -2238 1165 -2194
rect 1192 -2315 1193 -2237
rect 1290 -2238 1291 -2194
rect 1332 -2315 1333 -2237
rect 1423 -2238 1424 -2194
rect 1493 -2315 1494 -2237
rect 1542 -2238 1543 -2194
rect 1549 -2315 1550 -2237
rect 1773 -2238 1774 -2194
rect 93 -2240 94 -2194
rect 1423 -2315 1424 -2239
rect 1514 -2315 1515 -2239
rect 1570 -2240 1571 -2194
rect 1689 -2315 1690 -2239
rect 1843 -2240 1844 -2194
rect 93 -2315 94 -2241
rect 124 -2315 125 -2241
rect 198 -2242 199 -2194
rect 282 -2315 283 -2241
rect 394 -2315 395 -2241
rect 541 -2242 542 -2194
rect 576 -2315 577 -2241
rect 947 -2315 948 -2241
rect 975 -2315 976 -2241
rect 1290 -2315 1291 -2241
rect 1542 -2315 1543 -2241
rect 1584 -2242 1585 -2194
rect 1703 -2315 1704 -2241
rect 1857 -2242 1858 -2194
rect 198 -2315 199 -2243
rect 401 -2244 402 -2194
rect 429 -2244 430 -2194
rect 632 -2315 633 -2243
rect 649 -2244 650 -2194
rect 1416 -2315 1417 -2243
rect 1563 -2315 1564 -2243
rect 1633 -2244 1634 -2194
rect 1773 -2315 1774 -2243
rect 1801 -2244 1802 -2194
rect 205 -2246 206 -2194
rect 275 -2315 276 -2245
rect 345 -2246 346 -2194
rect 401 -2315 402 -2245
rect 429 -2315 430 -2245
rect 842 -2246 843 -2194
rect 1052 -2315 1053 -2245
rect 1346 -2246 1347 -2194
rect 1570 -2315 1571 -2245
rect 1654 -2246 1655 -2194
rect 72 -2248 73 -2194
rect 345 -2315 346 -2247
rect 366 -2248 367 -2194
rect 541 -2315 542 -2247
rect 611 -2315 612 -2247
rect 653 -2248 654 -2194
rect 656 -2315 657 -2247
rect 1094 -2315 1095 -2247
rect 1122 -2248 1123 -2194
rect 1160 -2248 1161 -2194
rect 1164 -2315 1165 -2247
rect 1234 -2248 1235 -2194
rect 1346 -2315 1347 -2247
rect 1437 -2248 1438 -2194
rect 1584 -2315 1585 -2247
rect 1661 -2248 1662 -2194
rect 72 -2315 73 -2249
rect 121 -2250 122 -2194
rect 156 -2250 157 -2194
rect 205 -2315 206 -2249
rect 208 -2315 209 -2249
rect 723 -2315 724 -2249
rect 744 -2250 745 -2194
rect 1234 -2315 1235 -2249
rect 1661 -2315 1662 -2249
rect 121 -2315 122 -2251
rect 142 -2315 143 -2251
rect 156 -2315 157 -2251
rect 1668 -2252 1669 -2194
rect 212 -2254 213 -2194
rect 380 -2315 381 -2253
rect 443 -2315 444 -2253
rect 450 -2254 451 -2194
rect 618 -2254 619 -2194
rect 800 -2315 801 -2253
rect 842 -2315 843 -2253
rect 905 -2254 906 -2194
rect 1087 -2315 1088 -2253
rect 1115 -2254 1116 -2194
rect 1122 -2315 1123 -2253
rect 1710 -2254 1711 -2194
rect 212 -2315 213 -2255
rect 758 -2256 759 -2194
rect 765 -2256 766 -2194
rect 1017 -2315 1018 -2255
rect 1115 -2315 1116 -2255
rect 1129 -2256 1130 -2194
rect 1213 -2256 1214 -2194
rect 1255 -2315 1256 -2255
rect 1293 -2315 1294 -2255
rect 1668 -2315 1669 -2255
rect 1710 -2315 1711 -2255
rect 1759 -2315 1760 -2255
rect 219 -2315 220 -2257
rect 436 -2258 437 -2194
rect 450 -2315 451 -2257
rect 499 -2258 500 -2194
rect 618 -2315 619 -2257
rect 933 -2258 934 -2194
rect 1129 -2315 1130 -2257
rect 1206 -2258 1207 -2194
rect 1220 -2315 1221 -2257
rect 1409 -2258 1410 -2194
rect 1437 -2315 1438 -2257
rect 1521 -2258 1522 -2194
rect 1633 -2315 1634 -2257
rect 1836 -2258 1837 -2194
rect 226 -2315 227 -2259
rect 240 -2260 241 -2194
rect 261 -2315 262 -2259
rect 359 -2260 360 -2194
rect 366 -2315 367 -2259
rect 555 -2260 556 -2194
rect 628 -2315 629 -2259
rect 1206 -2315 1207 -2259
rect 1409 -2315 1410 -2259
rect 1556 -2260 1557 -2194
rect 236 -2315 237 -2261
rect 1654 -2315 1655 -2261
rect 240 -2315 241 -2263
rect 1752 -2264 1753 -2194
rect 310 -2266 311 -2194
rect 359 -2315 360 -2265
rect 422 -2266 423 -2194
rect 933 -2315 934 -2265
rect 1521 -2315 1522 -2265
rect 1682 -2266 1683 -2194
rect 1752 -2315 1753 -2265
rect 1864 -2266 1865 -2194
rect 159 -2315 160 -2267
rect 310 -2315 311 -2267
rect 373 -2268 374 -2194
rect 422 -2315 423 -2267
rect 436 -2315 437 -2267
rect 870 -2268 871 -2194
rect 905 -2315 906 -2267
rect 940 -2268 941 -2194
rect 1556 -2315 1557 -2267
rect 1612 -2268 1613 -2194
rect 1682 -2315 1683 -2267
rect 1780 -2268 1781 -2194
rect 373 -2315 374 -2269
rect 548 -2270 549 -2194
rect 555 -2315 556 -2269
rect 681 -2270 682 -2194
rect 709 -2270 710 -2194
rect 863 -2315 864 -2269
rect 870 -2315 871 -2269
rect 898 -2270 899 -2194
rect 940 -2315 941 -2269
rect 982 -2270 983 -2194
rect 1612 -2315 1613 -2269
rect 1766 -2270 1767 -2194
rect 390 -2272 391 -2194
rect 1780 -2315 1781 -2271
rect 499 -2315 500 -2273
rect 534 -2274 535 -2194
rect 548 -2315 549 -2273
rect 604 -2274 605 -2194
rect 639 -2315 640 -2273
rect 758 -2315 759 -2273
rect 765 -2315 766 -2273
rect 856 -2274 857 -2194
rect 898 -2315 899 -2273
rect 1157 -2274 1158 -2194
rect 1731 -2274 1732 -2194
rect 1766 -2315 1767 -2273
rect 89 -2276 90 -2194
rect 534 -2315 535 -2275
rect 604 -2315 605 -2275
rect 674 -2276 675 -2194
rect 677 -2315 678 -2275
rect 1388 -2315 1389 -2275
rect 1472 -2276 1473 -2194
rect 1731 -2315 1732 -2275
rect 653 -2315 654 -2277
rect 1045 -2278 1046 -2194
rect 1157 -2315 1158 -2277
rect 1227 -2278 1228 -2194
rect 660 -2280 661 -2194
rect 681 -2315 682 -2279
rect 702 -2280 703 -2194
rect 709 -2315 710 -2279
rect 744 -2315 745 -2279
rect 807 -2280 808 -2194
rect 821 -2280 822 -2194
rect 856 -2315 857 -2279
rect 982 -2315 983 -2279
rect 996 -2280 997 -2194
rect 1185 -2315 1186 -2279
rect 1472 -2315 1473 -2279
rect 9 -2315 10 -2281
rect 996 -2315 997 -2281
rect 1227 -2315 1228 -2281
rect 1311 -2282 1312 -2194
rect 660 -2315 661 -2283
rect 667 -2284 668 -2194
rect 674 -2315 675 -2283
rect 1073 -2284 1074 -2194
rect 1311 -2315 1312 -2283
rect 1381 -2284 1382 -2194
rect 688 -2286 689 -2194
rect 702 -2315 703 -2285
rect 751 -2286 752 -2194
rect 1045 -2315 1046 -2285
rect 1073 -2315 1074 -2285
rect 1143 -2286 1144 -2194
rect 583 -2288 584 -2194
rect 688 -2315 689 -2287
rect 751 -2315 752 -2287
rect 824 -2315 825 -2287
rect 835 -2288 836 -2194
rect 1381 -2315 1382 -2287
rect 513 -2290 514 -2194
rect 583 -2315 584 -2289
rect 807 -2315 808 -2289
rect 828 -2290 829 -2194
rect 835 -2315 836 -2289
rect 887 -2315 888 -2289
rect 978 -2290 979 -2194
rect 1143 -2315 1144 -2289
rect 65 -2315 66 -2291
rect 513 -2315 514 -2291
rect 821 -2315 822 -2291
rect 1213 -2315 1214 -2291
rect 828 -2315 829 -2293
rect 1199 -2294 1200 -2194
rect 1199 -2315 1200 -2295
rect 1374 -2296 1375 -2194
rect 1374 -2315 1375 -2297
rect 1465 -2298 1466 -2194
rect 1465 -2315 1466 -2299
rect 1528 -2300 1529 -2194
rect 1507 -2302 1508 -2194
rect 1528 -2315 1529 -2301
rect 1507 -2315 1508 -2303
rect 1598 -2304 1599 -2194
rect 1069 -2306 1070 -2194
rect 1598 -2315 1599 -2305
rect 1069 -2315 1070 -2307
rect 1171 -2308 1172 -2194
rect 1171 -2315 1172 -2309
rect 1269 -2310 1270 -2194
rect 1269 -2315 1270 -2311
rect 1367 -2312 1368 -2194
rect 149 -2315 150 -2313
rect 1367 -2315 1368 -2313
rect 9 -2325 10 -2323
rect 170 -2325 171 -2323
rect 177 -2325 178 -2323
rect 1727 -2325 1728 -2323
rect 1731 -2325 1732 -2323
rect 1745 -2440 1746 -2324
rect 1748 -2325 1749 -2323
rect 1822 -2325 1823 -2323
rect 9 -2440 10 -2326
rect 492 -2327 493 -2323
rect 499 -2327 500 -2323
rect 817 -2327 818 -2323
rect 821 -2327 822 -2323
rect 1206 -2327 1207 -2323
rect 1216 -2440 1217 -2326
rect 1451 -2327 1452 -2323
rect 1577 -2327 1578 -2323
rect 1731 -2440 1732 -2326
rect 1755 -2440 1756 -2326
rect 1766 -2327 1767 -2323
rect 1780 -2327 1781 -2323
rect 1801 -2440 1802 -2326
rect 16 -2329 17 -2323
rect 618 -2329 619 -2323
rect 625 -2329 626 -2323
rect 1052 -2329 1053 -2323
rect 1069 -2329 1070 -2323
rect 1255 -2329 1256 -2323
rect 1276 -2329 1277 -2323
rect 1293 -2329 1294 -2323
rect 1307 -2329 1308 -2323
rect 1458 -2329 1459 -2323
rect 1738 -2329 1739 -2323
rect 1766 -2440 1767 -2328
rect 1787 -2329 1788 -2323
rect 1808 -2440 1809 -2328
rect 16 -2440 17 -2330
rect 432 -2440 433 -2330
rect 439 -2440 440 -2330
rect 457 -2331 458 -2323
rect 460 -2440 461 -2330
rect 590 -2331 591 -2323
rect 625 -2440 626 -2330
rect 905 -2331 906 -2323
rect 947 -2331 948 -2323
rect 1038 -2331 1039 -2323
rect 1052 -2440 1053 -2330
rect 1486 -2331 1487 -2323
rect 1675 -2331 1676 -2323
rect 1738 -2440 1739 -2330
rect 1759 -2331 1760 -2323
rect 1780 -2440 1781 -2330
rect 1787 -2440 1788 -2330
rect 1794 -2331 1795 -2323
rect 1797 -2440 1798 -2330
rect 1829 -2331 1830 -2323
rect 30 -2333 31 -2323
rect 114 -2333 115 -2323
rect 128 -2333 129 -2323
rect 128 -2440 129 -2332
rect 128 -2333 129 -2323
rect 128 -2440 129 -2332
rect 142 -2333 143 -2323
rect 212 -2333 213 -2323
rect 233 -2440 234 -2332
rect 387 -2333 388 -2323
rect 401 -2333 402 -2323
rect 401 -2440 402 -2332
rect 401 -2333 402 -2323
rect 401 -2440 402 -2332
rect 408 -2333 409 -2323
rect 733 -2440 734 -2332
rect 793 -2440 794 -2332
rect 807 -2333 808 -2323
rect 814 -2440 815 -2332
rect 975 -2333 976 -2323
rect 989 -2333 990 -2323
rect 989 -2440 990 -2332
rect 989 -2333 990 -2323
rect 989 -2440 990 -2332
rect 996 -2333 997 -2323
rect 1577 -2440 1578 -2332
rect 1619 -2333 1620 -2323
rect 1675 -2440 1676 -2332
rect 1759 -2440 1760 -2332
rect 1773 -2333 1774 -2323
rect 30 -2440 31 -2334
rect 149 -2335 150 -2323
rect 159 -2335 160 -2323
rect 324 -2335 325 -2323
rect 352 -2335 353 -2323
rect 667 -2335 668 -2323
rect 698 -2440 699 -2334
rect 842 -2335 843 -2323
rect 863 -2335 864 -2323
rect 975 -2440 976 -2334
rect 1020 -2440 1021 -2334
rect 1241 -2335 1242 -2323
rect 1248 -2335 1249 -2323
rect 1276 -2440 1277 -2334
rect 1290 -2335 1291 -2323
rect 1549 -2335 1550 -2323
rect 1619 -2440 1620 -2334
rect 1689 -2335 1690 -2323
rect 1717 -2335 1718 -2323
rect 1773 -2440 1774 -2334
rect 44 -2337 45 -2323
rect 236 -2337 237 -2323
rect 247 -2337 248 -2323
rect 247 -2440 248 -2336
rect 247 -2337 248 -2323
rect 247 -2440 248 -2336
rect 282 -2337 283 -2323
rect 464 -2337 465 -2323
rect 471 -2337 472 -2323
rect 618 -2440 619 -2336
rect 632 -2337 633 -2323
rect 632 -2440 633 -2336
rect 632 -2337 633 -2323
rect 632 -2440 633 -2336
rect 646 -2337 647 -2323
rect 842 -2440 843 -2336
rect 884 -2337 885 -2323
rect 1003 -2337 1004 -2323
rect 1017 -2337 1018 -2323
rect 1241 -2440 1242 -2336
rect 1321 -2440 1322 -2336
rect 1325 -2337 1326 -2323
rect 1342 -2440 1343 -2336
rect 1710 -2440 1711 -2336
rect 44 -2440 45 -2338
rect 226 -2339 227 -2323
rect 303 -2339 304 -2323
rect 530 -2440 531 -2338
rect 544 -2440 545 -2338
rect 639 -2339 640 -2323
rect 646 -2440 647 -2338
rect 887 -2339 888 -2323
rect 905 -2440 906 -2338
rect 912 -2339 913 -2323
rect 947 -2440 948 -2338
rect 961 -2339 962 -2323
rect 1024 -2339 1025 -2323
rect 1024 -2440 1025 -2338
rect 1024 -2339 1025 -2323
rect 1024 -2440 1025 -2338
rect 1038 -2440 1039 -2338
rect 1059 -2339 1060 -2323
rect 1066 -2339 1067 -2323
rect 1290 -2440 1291 -2338
rect 1370 -2339 1371 -2323
rect 1395 -2339 1396 -2323
rect 1423 -2339 1424 -2323
rect 1451 -2440 1452 -2338
rect 1486 -2440 1487 -2338
rect 1493 -2339 1494 -2323
rect 1542 -2339 1543 -2323
rect 1549 -2440 1550 -2338
rect 1633 -2339 1634 -2323
rect 1689 -2440 1690 -2338
rect 51 -2341 52 -2323
rect 1003 -2440 1004 -2340
rect 1010 -2341 1011 -2323
rect 1059 -2440 1060 -2340
rect 1066 -2440 1067 -2340
rect 1080 -2341 1081 -2323
rect 1087 -2341 1088 -2323
rect 1087 -2440 1088 -2340
rect 1087 -2341 1088 -2323
rect 1087 -2440 1088 -2340
rect 1101 -2341 1102 -2323
rect 1101 -2440 1102 -2340
rect 1101 -2341 1102 -2323
rect 1101 -2440 1102 -2340
rect 1115 -2341 1116 -2323
rect 1514 -2341 1515 -2323
rect 1521 -2341 1522 -2323
rect 1633 -2440 1634 -2340
rect 37 -2343 38 -2323
rect 1080 -2440 1081 -2342
rect 1115 -2440 1116 -2342
rect 1178 -2343 1179 -2323
rect 1188 -2343 1189 -2323
rect 1682 -2343 1683 -2323
rect 37 -2440 38 -2344
rect 240 -2345 241 -2323
rect 310 -2345 311 -2323
rect 457 -2440 458 -2344
rect 467 -2345 468 -2323
rect 1423 -2440 1424 -2344
rect 1430 -2345 1431 -2323
rect 1458 -2440 1459 -2344
rect 1465 -2345 1466 -2323
rect 1493 -2440 1494 -2344
rect 1521 -2440 1522 -2344
rect 1556 -2345 1557 -2323
rect 1640 -2345 1641 -2323
rect 1682 -2440 1683 -2344
rect 51 -2440 52 -2346
rect 243 -2347 244 -2323
rect 310 -2440 311 -2346
rect 446 -2440 447 -2346
rect 450 -2347 451 -2323
rect 464 -2440 465 -2346
rect 478 -2347 479 -2323
rect 492 -2440 493 -2346
rect 534 -2347 535 -2323
rect 961 -2440 962 -2346
rect 1010 -2440 1011 -2346
rect 1094 -2347 1095 -2323
rect 1129 -2347 1130 -2323
rect 1129 -2440 1130 -2346
rect 1129 -2347 1130 -2323
rect 1129 -2440 1130 -2346
rect 1136 -2347 1137 -2323
rect 1136 -2440 1137 -2346
rect 1136 -2347 1137 -2323
rect 1136 -2440 1137 -2346
rect 1157 -2347 1158 -2323
rect 1160 -2375 1161 -2346
rect 1171 -2347 1172 -2323
rect 1206 -2440 1207 -2346
rect 1213 -2347 1214 -2323
rect 1255 -2440 1256 -2346
rect 1283 -2347 1284 -2323
rect 1325 -2440 1326 -2346
rect 1360 -2347 1361 -2323
rect 1395 -2440 1396 -2346
rect 1437 -2347 1438 -2323
rect 1465 -2440 1466 -2346
rect 1479 -2347 1480 -2323
rect 1514 -2440 1515 -2346
rect 1640 -2440 1641 -2346
rect 1703 -2347 1704 -2323
rect 58 -2349 59 -2323
rect 82 -2440 83 -2348
rect 86 -2349 87 -2323
rect 677 -2349 678 -2323
rect 723 -2349 724 -2323
rect 996 -2440 997 -2348
rect 1017 -2440 1018 -2348
rect 1171 -2440 1172 -2348
rect 1227 -2349 1228 -2323
rect 1248 -2440 1249 -2348
rect 1339 -2349 1340 -2323
rect 1360 -2440 1361 -2348
rect 1416 -2349 1417 -2323
rect 1437 -2440 1438 -2348
rect 1444 -2349 1445 -2323
rect 1479 -2440 1480 -2348
rect 1500 -2349 1501 -2323
rect 1556 -2440 1557 -2348
rect 1661 -2349 1662 -2323
rect 1703 -2440 1704 -2348
rect 58 -2440 59 -2350
rect 219 -2351 220 -2323
rect 296 -2351 297 -2323
rect 677 -2440 678 -2350
rect 772 -2351 773 -2323
rect 1178 -2440 1179 -2350
rect 1227 -2440 1228 -2350
rect 1794 -2440 1795 -2350
rect 65 -2440 66 -2352
rect 485 -2353 486 -2323
rect 513 -2353 514 -2323
rect 534 -2440 535 -2352
rect 562 -2353 563 -2323
rect 824 -2353 825 -2323
rect 831 -2440 832 -2352
rect 1542 -2440 1543 -2352
rect 1626 -2353 1627 -2323
rect 1661 -2440 1662 -2352
rect 72 -2355 73 -2323
rect 110 -2440 111 -2354
rect 114 -2440 115 -2354
rect 198 -2355 199 -2323
rect 205 -2355 206 -2323
rect 499 -2440 500 -2354
rect 541 -2355 542 -2323
rect 562 -2440 563 -2354
rect 583 -2355 584 -2323
rect 590 -2440 591 -2354
rect 604 -2355 605 -2323
rect 639 -2440 640 -2354
rect 667 -2440 668 -2354
rect 702 -2355 703 -2323
rect 772 -2440 773 -2354
rect 786 -2355 787 -2323
rect 856 -2355 857 -2323
rect 887 -2440 888 -2354
rect 912 -2440 913 -2354
rect 926 -2355 927 -2323
rect 1055 -2440 1056 -2354
rect 1283 -2440 1284 -2354
rect 1332 -2355 1333 -2323
rect 1444 -2440 1445 -2354
rect 1591 -2355 1592 -2323
rect 1626 -2440 1627 -2354
rect 72 -2440 73 -2356
rect 100 -2357 101 -2323
rect 107 -2357 108 -2323
rect 408 -2440 409 -2356
rect 415 -2357 416 -2323
rect 471 -2440 472 -2356
rect 478 -2440 479 -2356
rect 681 -2357 682 -2323
rect 786 -2440 787 -2356
rect 807 -2440 808 -2356
rect 856 -2440 857 -2356
rect 870 -2357 871 -2323
rect 926 -2440 927 -2356
rect 1269 -2357 1270 -2323
rect 1339 -2440 1340 -2356
rect 1647 -2357 1648 -2323
rect 79 -2359 80 -2323
rect 226 -2440 227 -2358
rect 289 -2359 290 -2323
rect 296 -2440 297 -2358
rect 324 -2440 325 -2358
rect 527 -2359 528 -2323
rect 541 -2440 542 -2358
rect 688 -2359 689 -2323
rect 863 -2440 864 -2358
rect 884 -2440 885 -2358
rect 1094 -2440 1095 -2358
rect 1164 -2359 1165 -2323
rect 1199 -2359 1200 -2323
rect 1332 -2440 1333 -2358
rect 1388 -2359 1389 -2323
rect 1416 -2440 1417 -2358
rect 1528 -2359 1529 -2323
rect 1591 -2440 1592 -2358
rect 1605 -2359 1606 -2323
rect 1647 -2440 1648 -2358
rect 86 -2440 87 -2360
rect 93 -2361 94 -2323
rect 96 -2440 97 -2360
rect 1717 -2440 1718 -2360
rect 93 -2440 94 -2362
rect 124 -2363 125 -2323
rect 135 -2363 136 -2323
rect 303 -2440 304 -2362
rect 352 -2440 353 -2362
rect 1118 -2363 1119 -2323
rect 1150 -2363 1151 -2323
rect 1199 -2440 1200 -2362
rect 1269 -2440 1270 -2362
rect 1318 -2363 1319 -2323
rect 1388 -2440 1389 -2362
rect 1696 -2363 1697 -2323
rect 100 -2440 101 -2364
rect 163 -2365 164 -2323
rect 170 -2440 171 -2364
rect 422 -2365 423 -2323
rect 429 -2365 430 -2323
rect 723 -2440 724 -2364
rect 870 -2440 871 -2364
rect 877 -2365 878 -2323
rect 1150 -2440 1151 -2364
rect 1213 -2440 1214 -2364
rect 1563 -2365 1564 -2323
rect 1605 -2440 1606 -2364
rect 1654 -2365 1655 -2323
rect 1696 -2440 1697 -2364
rect 121 -2440 122 -2366
rect 513 -2440 514 -2366
rect 520 -2367 521 -2323
rect 688 -2440 689 -2366
rect 877 -2440 878 -2366
rect 940 -2367 941 -2323
rect 1157 -2440 1158 -2366
rect 1220 -2367 1221 -2323
rect 1507 -2367 1508 -2323
rect 1563 -2440 1564 -2366
rect 1598 -2367 1599 -2323
rect 1654 -2440 1655 -2366
rect 107 -2440 108 -2368
rect 940 -2440 941 -2368
rect 1083 -2440 1084 -2368
rect 1507 -2440 1508 -2368
rect 1598 -2440 1599 -2368
rect 1668 -2369 1669 -2323
rect 131 -2440 132 -2370
rect 135 -2440 136 -2370
rect 142 -2440 143 -2370
rect 999 -2371 1000 -2323
rect 1164 -2440 1165 -2370
rect 1612 -2371 1613 -2323
rect 149 -2440 150 -2372
rect 576 -2373 577 -2323
rect 583 -2440 584 -2372
rect 968 -2373 969 -2323
rect 1192 -2373 1193 -2323
rect 1220 -2440 1221 -2372
rect 1535 -2373 1536 -2323
rect 1668 -2440 1669 -2372
rect 156 -2375 157 -2323
rect 198 -2440 199 -2374
rect 212 -2440 213 -2374
rect 215 -2375 216 -2323
rect 219 -2440 220 -2374
rect 436 -2375 437 -2323
rect 450 -2440 451 -2374
rect 737 -2375 738 -2323
rect 968 -2440 969 -2374
rect 982 -2375 983 -2323
rect 1192 -2440 1193 -2374
rect 1535 -2440 1536 -2374
rect 1570 -2375 1571 -2323
rect 1584 -2375 1585 -2323
rect 1612 -2440 1613 -2374
rect 156 -2440 157 -2376
rect 1185 -2377 1186 -2323
rect 1402 -2377 1403 -2323
rect 1584 -2440 1585 -2376
rect 163 -2440 164 -2378
rect 730 -2379 731 -2323
rect 737 -2440 738 -2378
rect 779 -2379 780 -2323
rect 891 -2379 892 -2323
rect 1185 -2440 1186 -2378
rect 1374 -2379 1375 -2323
rect 1402 -2440 1403 -2378
rect 1570 -2440 1571 -2378
rect 1752 -2379 1753 -2323
rect 177 -2440 178 -2380
rect 275 -2381 276 -2323
rect 366 -2381 367 -2323
rect 429 -2440 430 -2380
rect 436 -2440 437 -2380
rect 653 -2440 654 -2380
rect 681 -2440 682 -2380
rect 695 -2381 696 -2323
rect 730 -2440 731 -2380
rect 1500 -2440 1501 -2380
rect 184 -2383 185 -2323
rect 282 -2440 283 -2382
rect 366 -2440 367 -2382
rect 380 -2383 381 -2323
rect 387 -2440 388 -2382
rect 821 -2440 822 -2382
rect 891 -2440 892 -2382
rect 919 -2383 920 -2323
rect 982 -2440 983 -2382
rect 1031 -2383 1032 -2323
rect 1346 -2383 1347 -2323
rect 1374 -2440 1375 -2382
rect 184 -2440 185 -2384
rect 359 -2385 360 -2323
rect 390 -2440 391 -2384
rect 702 -2440 703 -2384
rect 828 -2385 829 -2323
rect 1346 -2440 1347 -2384
rect 191 -2387 192 -2323
rect 240 -2440 241 -2386
rect 261 -2387 262 -2323
rect 422 -2440 423 -2386
rect 485 -2440 486 -2386
rect 548 -2387 549 -2323
rect 572 -2387 573 -2323
rect 779 -2440 780 -2386
rect 828 -2440 829 -2386
rect 1724 -2440 1725 -2386
rect 23 -2389 24 -2323
rect 191 -2440 192 -2388
rect 205 -2440 206 -2388
rect 1752 -2440 1753 -2388
rect 261 -2440 262 -2390
rect 443 -2391 444 -2323
rect 520 -2440 521 -2390
rect 849 -2391 850 -2323
rect 919 -2440 920 -2390
rect 933 -2391 934 -2323
rect 1031 -2440 1032 -2390
rect 1045 -2391 1046 -2323
rect 275 -2440 276 -2392
rect 317 -2393 318 -2323
rect 338 -2393 339 -2323
rect 359 -2440 360 -2392
rect 394 -2393 395 -2323
rect 415 -2440 416 -2392
rect 527 -2440 528 -2392
rect 1430 -2440 1431 -2392
rect 289 -2440 290 -2394
rect 443 -2440 444 -2394
rect 548 -2440 549 -2394
rect 709 -2395 710 -2323
rect 800 -2395 801 -2323
rect 849 -2440 850 -2394
rect 933 -2440 934 -2394
rect 954 -2395 955 -2323
rect 1045 -2440 1046 -2394
rect 1304 -2395 1305 -2323
rect 317 -2440 318 -2396
rect 506 -2397 507 -2323
rect 569 -2397 570 -2323
rect 709 -2440 710 -2396
rect 765 -2397 766 -2323
rect 800 -2440 801 -2396
rect 835 -2397 836 -2323
rect 954 -2440 955 -2396
rect 1262 -2397 1263 -2323
rect 1304 -2440 1305 -2396
rect 268 -2399 269 -2323
rect 506 -2440 507 -2398
rect 555 -2399 556 -2323
rect 765 -2440 766 -2398
rect 835 -2440 836 -2398
rect 1167 -2440 1168 -2398
rect 268 -2440 269 -2400
rect 331 -2401 332 -2323
rect 338 -2440 339 -2400
rect 898 -2401 899 -2323
rect 1143 -2401 1144 -2323
rect 1262 -2440 1263 -2400
rect 331 -2440 332 -2402
rect 674 -2403 675 -2323
rect 695 -2440 696 -2402
rect 1391 -2440 1392 -2402
rect 254 -2405 255 -2323
rect 674 -2440 675 -2404
rect 898 -2440 899 -2404
rect 1713 -2405 1714 -2323
rect 117 -2407 118 -2323
rect 254 -2440 255 -2406
rect 341 -2440 342 -2406
rect 380 -2440 381 -2406
rect 404 -2440 405 -2406
rect 1528 -2440 1529 -2406
rect 345 -2409 346 -2323
rect 394 -2440 395 -2408
rect 569 -2440 570 -2408
rect 611 -2409 612 -2323
rect 656 -2409 657 -2323
rect 1143 -2440 1144 -2408
rect 373 -2411 374 -2323
rect 555 -2440 556 -2410
rect 576 -2440 577 -2410
rect 1122 -2411 1123 -2323
rect 373 -2440 374 -2412
rect 796 -2413 797 -2323
rect 1108 -2413 1109 -2323
rect 1122 -2440 1123 -2412
rect 597 -2415 598 -2323
rect 611 -2440 612 -2414
rect 1073 -2415 1074 -2323
rect 1108 -2440 1109 -2414
rect 345 -2440 346 -2416
rect 597 -2440 598 -2416
rect 604 -2440 605 -2416
rect 660 -2417 661 -2323
rect 1073 -2440 1074 -2416
rect 1367 -2417 1368 -2323
rect 660 -2440 661 -2418
rect 950 -2419 951 -2323
rect 1367 -2440 1368 -2418
rect 1472 -2419 1473 -2323
rect 1311 -2421 1312 -2323
rect 1472 -2440 1473 -2420
rect 1311 -2440 1312 -2422
rect 1353 -2423 1354 -2323
rect 1297 -2425 1298 -2323
rect 1353 -2440 1354 -2424
rect 1297 -2440 1298 -2426
rect 1409 -2427 1410 -2323
rect 1381 -2429 1382 -2323
rect 1409 -2440 1410 -2428
rect 1234 -2431 1235 -2323
rect 1381 -2440 1382 -2430
rect 758 -2433 759 -2323
rect 1234 -2440 1235 -2432
rect 744 -2435 745 -2323
rect 758 -2440 759 -2434
rect 744 -2440 745 -2436
rect 751 -2437 752 -2323
rect 716 -2439 717 -2323
rect 751 -2440 752 -2438
rect 9 -2450 10 -2448
rect 597 -2450 598 -2448
rect 632 -2450 633 -2448
rect 632 -2575 633 -2449
rect 632 -2450 633 -2448
rect 632 -2575 633 -2449
rect 646 -2450 647 -2448
rect 646 -2575 647 -2449
rect 646 -2450 647 -2448
rect 646 -2575 647 -2449
rect 723 -2450 724 -2448
rect 1017 -2450 1018 -2448
rect 1020 -2450 1021 -2448
rect 1486 -2450 1487 -2448
rect 1741 -2575 1742 -2449
rect 1773 -2450 1774 -2448
rect 1808 -2450 1809 -2448
rect 1815 -2575 1816 -2449
rect 16 -2452 17 -2448
rect 23 -2575 24 -2451
rect 44 -2452 45 -2448
rect 387 -2452 388 -2448
rect 408 -2452 409 -2448
rect 719 -2452 720 -2448
rect 726 -2575 727 -2451
rect 1717 -2452 1718 -2448
rect 1745 -2452 1746 -2448
rect 1745 -2575 1746 -2451
rect 1745 -2452 1746 -2448
rect 1745 -2575 1746 -2451
rect 1752 -2575 1753 -2451
rect 1759 -2452 1760 -2448
rect 1773 -2575 1774 -2451
rect 1794 -2452 1795 -2448
rect 1801 -2452 1802 -2448
rect 1808 -2575 1809 -2451
rect 16 -2575 17 -2453
rect 677 -2454 678 -2448
rect 807 -2454 808 -2448
rect 810 -2486 811 -2453
rect 814 -2454 815 -2448
rect 814 -2575 815 -2453
rect 814 -2454 815 -2448
rect 814 -2575 815 -2453
rect 828 -2454 829 -2448
rect 852 -2575 853 -2453
rect 856 -2454 857 -2448
rect 856 -2575 857 -2453
rect 856 -2454 857 -2448
rect 856 -2575 857 -2453
rect 884 -2454 885 -2448
rect 912 -2454 913 -2448
rect 919 -2454 920 -2448
rect 919 -2575 920 -2453
rect 919 -2454 920 -2448
rect 919 -2575 920 -2453
rect 950 -2575 951 -2453
rect 1381 -2454 1382 -2448
rect 1423 -2454 1424 -2448
rect 1423 -2575 1424 -2453
rect 1423 -2454 1424 -2448
rect 1423 -2575 1424 -2453
rect 1619 -2454 1620 -2448
rect 1717 -2575 1718 -2453
rect 1759 -2575 1760 -2453
rect 1766 -2454 1767 -2448
rect 44 -2575 45 -2455
rect 149 -2456 150 -2448
rect 159 -2575 160 -2455
rect 432 -2456 433 -2448
rect 439 -2456 440 -2448
rect 1094 -2456 1095 -2448
rect 1132 -2575 1133 -2455
rect 1521 -2456 1522 -2448
rect 1570 -2456 1571 -2448
rect 1766 -2575 1767 -2455
rect 51 -2458 52 -2448
rect 544 -2458 545 -2448
rect 583 -2458 584 -2448
rect 786 -2458 787 -2448
rect 807 -2575 808 -2457
rect 954 -2458 955 -2448
rect 982 -2458 983 -2448
rect 1118 -2575 1119 -2457
rect 1150 -2458 1151 -2448
rect 1486 -2575 1487 -2457
rect 1521 -2575 1522 -2457
rect 1542 -2458 1543 -2448
rect 1619 -2575 1620 -2457
rect 1668 -2458 1669 -2448
rect 51 -2575 52 -2459
rect 576 -2460 577 -2448
rect 597 -2575 598 -2459
rect 821 -2460 822 -2448
rect 828 -2575 829 -2459
rect 863 -2460 864 -2448
rect 884 -2575 885 -2459
rect 926 -2460 927 -2448
rect 940 -2460 941 -2448
rect 954 -2575 955 -2459
rect 968 -2460 969 -2448
rect 982 -2575 983 -2459
rect 1038 -2460 1039 -2448
rect 1038 -2575 1039 -2459
rect 1038 -2460 1039 -2448
rect 1038 -2575 1039 -2459
rect 1055 -2575 1056 -2459
rect 1248 -2460 1249 -2448
rect 1325 -2460 1326 -2448
rect 1339 -2575 1340 -2459
rect 1353 -2460 1354 -2448
rect 1353 -2575 1354 -2459
rect 1353 -2460 1354 -2448
rect 1353 -2575 1354 -2459
rect 1381 -2575 1382 -2459
rect 1395 -2460 1396 -2448
rect 1542 -2575 1543 -2459
rect 1556 -2460 1557 -2448
rect 1668 -2575 1669 -2459
rect 1710 -2460 1711 -2448
rect 58 -2462 59 -2448
rect 401 -2462 402 -2448
rect 408 -2575 409 -2461
rect 712 -2575 713 -2461
rect 786 -2575 787 -2461
rect 842 -2462 843 -2448
rect 887 -2462 888 -2448
rect 1731 -2462 1732 -2448
rect 58 -2575 59 -2463
rect 261 -2464 262 -2448
rect 324 -2464 325 -2448
rect 723 -2575 724 -2463
rect 821 -2575 822 -2463
rect 1045 -2464 1046 -2448
rect 1076 -2575 1077 -2463
rect 1696 -2464 1697 -2448
rect 30 -2466 31 -2448
rect 261 -2575 262 -2465
rect 275 -2466 276 -2448
rect 324 -2575 325 -2465
rect 352 -2466 353 -2448
rect 1395 -2575 1396 -2465
rect 1556 -2575 1557 -2465
rect 1675 -2466 1676 -2448
rect 1689 -2466 1690 -2448
rect 1710 -2575 1711 -2465
rect 30 -2575 31 -2467
rect 212 -2468 213 -2448
rect 226 -2468 227 -2448
rect 401 -2575 402 -2467
rect 429 -2575 430 -2467
rect 611 -2468 612 -2448
rect 842 -2575 843 -2467
rect 1066 -2468 1067 -2448
rect 1087 -2468 1088 -2448
rect 1094 -2575 1095 -2467
rect 1150 -2575 1151 -2467
rect 1178 -2468 1179 -2448
rect 1195 -2575 1196 -2467
rect 1633 -2468 1634 -2448
rect 1640 -2468 1641 -2448
rect 1731 -2575 1732 -2467
rect 65 -2470 66 -2448
rect 390 -2470 391 -2448
rect 450 -2470 451 -2448
rect 516 -2470 517 -2448
rect 530 -2470 531 -2448
rect 569 -2470 570 -2448
rect 600 -2470 601 -2448
rect 1178 -2575 1179 -2469
rect 1325 -2575 1326 -2469
rect 1374 -2470 1375 -2448
rect 1640 -2575 1641 -2469
rect 1654 -2470 1655 -2448
rect 1675 -2575 1676 -2469
rect 1724 -2470 1725 -2448
rect 65 -2575 66 -2471
rect 317 -2472 318 -2448
rect 352 -2575 353 -2471
rect 1167 -2472 1168 -2448
rect 1332 -2472 1333 -2448
rect 1801 -2575 1802 -2471
rect 72 -2474 73 -2448
rect 387 -2575 388 -2473
rect 457 -2474 458 -2448
rect 583 -2575 584 -2473
rect 600 -2575 601 -2473
rect 695 -2474 696 -2448
rect 905 -2474 906 -2448
rect 912 -2575 913 -2473
rect 940 -2575 941 -2473
rect 1059 -2474 1060 -2448
rect 1066 -2575 1067 -2473
rect 1129 -2474 1130 -2448
rect 1160 -2575 1161 -2473
rect 1661 -2474 1662 -2448
rect 1689 -2575 1690 -2473
rect 1738 -2474 1739 -2448
rect 72 -2575 73 -2475
rect 194 -2476 195 -2448
rect 198 -2476 199 -2448
rect 212 -2575 213 -2475
rect 226 -2575 227 -2475
rect 947 -2476 948 -2448
rect 971 -2575 972 -2475
rect 1374 -2575 1375 -2475
rect 1598 -2476 1599 -2448
rect 1724 -2575 1725 -2475
rect 1738 -2575 1739 -2475
rect 1780 -2476 1781 -2448
rect 82 -2478 83 -2448
rect 233 -2478 234 -2448
rect 243 -2575 244 -2477
rect 1010 -2478 1011 -2448
rect 1048 -2575 1049 -2477
rect 1661 -2575 1662 -2477
rect 1696 -2575 1697 -2477
rect 1787 -2478 1788 -2448
rect 86 -2480 87 -2448
rect 86 -2575 87 -2479
rect 86 -2480 87 -2448
rect 86 -2575 87 -2479
rect 93 -2480 94 -2448
rect 380 -2480 381 -2448
rect 443 -2480 444 -2448
rect 1598 -2575 1599 -2479
rect 1654 -2575 1655 -2479
rect 1682 -2480 1683 -2448
rect 93 -2575 94 -2481
rect 268 -2482 269 -2448
rect 275 -2575 276 -2481
rect 394 -2482 395 -2448
rect 443 -2575 444 -2481
rect 506 -2482 507 -2448
rect 513 -2482 514 -2448
rect 590 -2482 591 -2448
rect 681 -2482 682 -2448
rect 695 -2575 696 -2481
rect 740 -2575 741 -2481
rect 947 -2575 948 -2481
rect 996 -2482 997 -2448
rect 1010 -2575 1011 -2481
rect 1087 -2575 1088 -2481
rect 1388 -2482 1389 -2448
rect 96 -2484 97 -2448
rect 345 -2484 346 -2448
rect 366 -2484 367 -2448
rect 394 -2575 395 -2483
rect 457 -2575 458 -2483
rect 849 -2484 850 -2448
rect 877 -2484 878 -2448
rect 905 -2575 906 -2483
rect 989 -2484 990 -2448
rect 996 -2575 997 -2483
rect 1129 -2575 1130 -2483
rect 1248 -2575 1249 -2483
rect 1255 -2484 1256 -2448
rect 1682 -2575 1683 -2483
rect 37 -2486 38 -2448
rect 345 -2575 346 -2485
rect 366 -2575 367 -2485
rect 618 -2486 619 -2448
rect 653 -2486 654 -2448
rect 681 -2575 682 -2485
rect 1059 -2575 1060 -2485
rect 1115 -2486 1116 -2448
rect 1255 -2575 1256 -2485
rect 1321 -2486 1322 -2448
rect 1780 -2575 1781 -2485
rect 37 -2575 38 -2487
rect 114 -2488 115 -2448
rect 128 -2488 129 -2448
rect 289 -2488 290 -2448
rect 317 -2575 318 -2487
rect 460 -2488 461 -2448
rect 471 -2488 472 -2448
rect 527 -2488 528 -2448
rect 541 -2575 542 -2487
rect 660 -2488 661 -2448
rect 849 -2575 850 -2487
rect 926 -2575 927 -2487
rect 989 -2575 990 -2487
rect 1318 -2488 1319 -2448
rect 1332 -2575 1333 -2487
rect 1493 -2488 1494 -2448
rect 100 -2490 101 -2448
rect 114 -2575 115 -2489
rect 128 -2575 129 -2489
rect 282 -2490 283 -2448
rect 289 -2575 290 -2489
rect 303 -2490 304 -2448
rect 415 -2490 416 -2448
rect 471 -2575 472 -2489
rect 478 -2490 479 -2448
rect 590 -2575 591 -2489
rect 604 -2490 605 -2448
rect 660 -2575 661 -2489
rect 1115 -2575 1116 -2489
rect 1297 -2490 1298 -2448
rect 1318 -2575 1319 -2489
rect 1360 -2490 1361 -2448
rect 1367 -2490 1368 -2448
rect 1493 -2575 1494 -2489
rect 100 -2575 101 -2491
rect 1346 -2492 1347 -2448
rect 1367 -2575 1368 -2491
rect 1465 -2492 1466 -2448
rect 107 -2494 108 -2448
rect 338 -2494 339 -2448
rect 478 -2575 479 -2493
rect 737 -2494 738 -2448
rect 1003 -2494 1004 -2448
rect 1346 -2575 1347 -2493
rect 1388 -2575 1389 -2493
rect 1402 -2494 1403 -2448
rect 1465 -2575 1466 -2493
rect 1479 -2494 1480 -2448
rect 107 -2575 108 -2495
rect 1185 -2496 1186 -2448
rect 1241 -2496 1242 -2448
rect 1787 -2575 1788 -2495
rect 110 -2498 111 -2448
rect 1017 -2575 1018 -2497
rect 1101 -2498 1102 -2448
rect 1185 -2575 1186 -2497
rect 1241 -2575 1242 -2497
rect 1290 -2498 1291 -2448
rect 1402 -2575 1403 -2497
rect 1409 -2498 1410 -2448
rect 1479 -2575 1480 -2497
rect 1507 -2498 1508 -2448
rect 103 -2575 104 -2499
rect 1101 -2575 1102 -2499
rect 1157 -2500 1158 -2448
rect 1297 -2575 1298 -2499
rect 1409 -2575 1410 -2499
rect 1416 -2500 1417 -2448
rect 131 -2502 132 -2448
rect 863 -2575 864 -2501
rect 1164 -2502 1165 -2448
rect 1311 -2502 1312 -2448
rect 1416 -2575 1417 -2501
rect 1437 -2502 1438 -2448
rect 135 -2504 136 -2448
rect 436 -2504 437 -2448
rect 485 -2504 486 -2448
rect 576 -2575 577 -2503
rect 604 -2575 605 -2503
rect 1020 -2575 1021 -2503
rect 1164 -2575 1165 -2503
rect 1199 -2504 1200 -2448
rect 1269 -2504 1270 -2448
rect 1360 -2575 1361 -2503
rect 1437 -2575 1438 -2503
rect 1451 -2504 1452 -2448
rect 135 -2575 136 -2505
rect 1045 -2575 1046 -2505
rect 1080 -2506 1081 -2448
rect 1269 -2575 1270 -2505
rect 1290 -2575 1291 -2505
rect 1514 -2506 1515 -2448
rect 142 -2508 143 -2448
rect 415 -2575 416 -2507
rect 436 -2575 437 -2507
rect 1031 -2508 1032 -2448
rect 1080 -2575 1081 -2507
rect 1136 -2508 1137 -2448
rect 1311 -2575 1312 -2507
rect 1699 -2575 1700 -2507
rect 121 -2510 122 -2448
rect 142 -2575 143 -2509
rect 149 -2575 150 -2509
rect 1633 -2575 1634 -2509
rect 121 -2575 122 -2511
rect 156 -2512 157 -2448
rect 163 -2512 164 -2448
rect 380 -2575 381 -2511
rect 485 -2575 486 -2511
rect 835 -2512 836 -2448
rect 1024 -2512 1025 -2448
rect 1031 -2575 1032 -2511
rect 1122 -2512 1123 -2448
rect 1199 -2575 1200 -2511
rect 1514 -2575 1515 -2511
rect 1528 -2512 1529 -2448
rect 152 -2575 153 -2513
rect 611 -2575 612 -2513
rect 639 -2514 640 -2448
rect 653 -2575 654 -2513
rect 674 -2514 675 -2448
rect 1451 -2575 1452 -2513
rect 1528 -2575 1529 -2513
rect 1703 -2514 1704 -2448
rect 163 -2575 164 -2515
rect 1052 -2575 1053 -2515
rect 1073 -2516 1074 -2448
rect 1703 -2575 1704 -2515
rect 170 -2518 171 -2448
rect 338 -2575 339 -2517
rect 492 -2518 493 -2448
rect 831 -2518 832 -2448
rect 1108 -2518 1109 -2448
rect 1122 -2575 1123 -2517
rect 170 -2575 171 -2519
rect 1143 -2520 1144 -2448
rect 173 -2575 174 -2521
rect 310 -2522 311 -2448
rect 492 -2575 493 -2521
rect 499 -2522 500 -2448
rect 506 -2575 507 -2521
rect 688 -2522 689 -2448
rect 702 -2522 703 -2448
rect 1024 -2575 1025 -2521
rect 1108 -2575 1109 -2521
rect 1192 -2522 1193 -2448
rect 191 -2524 192 -2448
rect 877 -2575 878 -2523
rect 1143 -2575 1144 -2523
rect 1206 -2524 1207 -2448
rect 191 -2575 192 -2525
rect 870 -2526 871 -2448
rect 1192 -2575 1193 -2525
rect 1444 -2526 1445 -2448
rect 198 -2575 199 -2527
rect 558 -2575 559 -2527
rect 569 -2575 570 -2527
rect 961 -2528 962 -2448
rect 1206 -2575 1207 -2527
rect 1220 -2528 1221 -2448
rect 1444 -2575 1445 -2527
rect 1458 -2528 1459 -2448
rect 219 -2530 220 -2448
rect 618 -2575 619 -2529
rect 667 -2530 668 -2448
rect 702 -2575 703 -2529
rect 737 -2575 738 -2529
rect 1570 -2575 1571 -2529
rect 219 -2575 220 -2531
rect 464 -2532 465 -2448
rect 499 -2575 500 -2531
rect 534 -2532 535 -2448
rect 674 -2575 675 -2531
rect 709 -2532 710 -2448
rect 789 -2532 790 -2448
rect 835 -2575 836 -2531
rect 870 -2575 871 -2531
rect 933 -2532 934 -2448
rect 961 -2575 962 -2531
rect 975 -2532 976 -2448
rect 1220 -2575 1221 -2531
rect 1276 -2532 1277 -2448
rect 233 -2575 234 -2533
rect 240 -2534 241 -2448
rect 247 -2534 248 -2448
rect 450 -2575 451 -2533
rect 464 -2575 465 -2533
rect 548 -2534 549 -2448
rect 688 -2575 689 -2533
rect 751 -2534 752 -2448
rect 975 -2575 976 -2533
rect 1171 -2534 1172 -2448
rect 1276 -2575 1277 -2533
rect 1472 -2534 1473 -2448
rect 247 -2575 248 -2535
rect 1157 -2575 1158 -2535
rect 1171 -2575 1172 -2535
rect 1535 -2536 1536 -2448
rect 254 -2538 255 -2448
rect 303 -2575 304 -2537
rect 310 -2575 311 -2537
rect 628 -2575 629 -2537
rect 709 -2575 710 -2537
rect 1003 -2575 1004 -2537
rect 1472 -2575 1473 -2537
rect 1500 -2538 1501 -2448
rect 1535 -2575 1536 -2537
rect 1549 -2538 1550 -2448
rect 254 -2575 255 -2539
rect 373 -2540 374 -2448
rect 513 -2575 514 -2539
rect 555 -2540 556 -2448
rect 730 -2540 731 -2448
rect 933 -2575 934 -2539
rect 1500 -2575 1501 -2539
rect 1563 -2540 1564 -2448
rect 268 -2575 269 -2541
rect 716 -2542 717 -2448
rect 730 -2575 731 -2541
rect 1174 -2575 1175 -2541
rect 1549 -2575 1550 -2541
rect 1577 -2542 1578 -2448
rect 282 -2575 283 -2543
rect 331 -2544 332 -2448
rect 359 -2544 360 -2448
rect 373 -2575 374 -2543
rect 520 -2544 521 -2448
rect 555 -2575 556 -2543
rect 716 -2575 717 -2543
rect 758 -2544 759 -2448
rect 1563 -2575 1564 -2543
rect 1584 -2544 1585 -2448
rect 177 -2546 178 -2448
rect 331 -2575 332 -2545
rect 520 -2575 521 -2545
rect 800 -2546 801 -2448
rect 1577 -2575 1578 -2545
rect 1591 -2546 1592 -2448
rect 177 -2575 178 -2547
rect 205 -2548 206 -2448
rect 527 -2575 528 -2547
rect 562 -2548 563 -2448
rect 625 -2548 626 -2448
rect 800 -2575 801 -2547
rect 1584 -2575 1585 -2547
rect 1605 -2548 1606 -2448
rect 184 -2550 185 -2448
rect 359 -2575 360 -2549
rect 534 -2575 535 -2549
rect 744 -2550 745 -2448
rect 751 -2575 752 -2549
rect 1213 -2550 1214 -2448
rect 1591 -2575 1592 -2549
rect 1647 -2550 1648 -2448
rect 184 -2575 185 -2551
rect 341 -2552 342 -2448
rect 548 -2575 549 -2551
rect 992 -2575 993 -2551
rect 1213 -2575 1214 -2551
rect 1227 -2552 1228 -2448
rect 1283 -2552 1284 -2448
rect 1647 -2575 1648 -2551
rect 205 -2575 206 -2553
rect 422 -2554 423 -2448
rect 562 -2575 563 -2553
rect 639 -2575 640 -2553
rect 744 -2575 745 -2553
rect 765 -2554 766 -2448
rect 968 -2575 969 -2553
rect 1227 -2575 1228 -2553
rect 1262 -2554 1263 -2448
rect 1283 -2575 1284 -2553
rect 1605 -2575 1606 -2553
rect 1612 -2554 1613 -2448
rect 156 -2575 157 -2555
rect 422 -2575 423 -2555
rect 625 -2575 626 -2555
rect 1458 -2575 1459 -2555
rect 1612 -2575 1613 -2555
rect 1626 -2556 1627 -2448
rect 79 -2558 80 -2448
rect 1626 -2575 1627 -2557
rect 79 -2575 80 -2559
rect 296 -2560 297 -2448
rect 758 -2575 759 -2559
rect 772 -2560 773 -2448
rect 1262 -2575 1263 -2559
rect 1430 -2560 1431 -2448
rect 296 -2575 297 -2561
rect 404 -2562 405 -2448
rect 765 -2575 766 -2561
rect 779 -2562 780 -2448
rect 1234 -2562 1235 -2448
rect 1430 -2575 1431 -2561
rect 772 -2575 773 -2563
rect 793 -2564 794 -2448
rect 1234 -2575 1235 -2563
rect 1304 -2564 1305 -2448
rect 110 -2575 111 -2565
rect 1304 -2575 1305 -2565
rect 670 -2575 671 -2567
rect 793 -2575 794 -2567
rect 779 -2575 780 -2569
rect 898 -2570 899 -2448
rect 891 -2572 892 -2448
rect 898 -2575 899 -2571
rect 453 -2575 454 -2573
rect 891 -2575 892 -2573
rect 9 -2708 10 -2584
rect 443 -2585 444 -2583
rect 450 -2585 451 -2583
rect 1059 -2585 1060 -2583
rect 1062 -2708 1063 -2584
rect 1276 -2585 1277 -2583
rect 1293 -2708 1294 -2584
rect 1339 -2585 1340 -2583
rect 1465 -2585 1466 -2583
rect 1465 -2708 1466 -2584
rect 1465 -2585 1466 -2583
rect 1465 -2708 1466 -2584
rect 1510 -2585 1511 -2583
rect 1591 -2585 1592 -2583
rect 1724 -2585 1725 -2583
rect 1724 -2708 1725 -2584
rect 1724 -2585 1725 -2583
rect 1724 -2708 1725 -2584
rect 1738 -2585 1739 -2583
rect 1780 -2585 1781 -2583
rect 16 -2587 17 -2583
rect 16 -2708 17 -2586
rect 16 -2587 17 -2583
rect 16 -2708 17 -2586
rect 44 -2587 45 -2583
rect 628 -2587 629 -2583
rect 639 -2587 640 -2583
rect 807 -2587 808 -2583
rect 852 -2587 853 -2583
rect 996 -2587 997 -2583
rect 1020 -2587 1021 -2583
rect 1108 -2587 1109 -2583
rect 1115 -2708 1116 -2586
rect 1311 -2587 1312 -2583
rect 1339 -2708 1340 -2586
rect 1374 -2587 1375 -2583
rect 1563 -2587 1564 -2583
rect 1563 -2708 1564 -2586
rect 1563 -2587 1564 -2583
rect 1563 -2708 1564 -2586
rect 1769 -2708 1770 -2586
rect 1783 -2708 1784 -2586
rect 44 -2708 45 -2588
rect 779 -2589 780 -2583
rect 807 -2708 808 -2588
rect 828 -2589 829 -2583
rect 866 -2708 867 -2588
rect 1507 -2589 1508 -2583
rect 107 -2591 108 -2583
rect 366 -2591 367 -2583
rect 443 -2708 444 -2590
rect 583 -2591 584 -2583
rect 660 -2591 661 -2583
rect 712 -2591 713 -2583
rect 726 -2591 727 -2583
rect 1647 -2591 1648 -2583
rect 79 -2593 80 -2583
rect 107 -2708 108 -2592
rect 121 -2593 122 -2583
rect 240 -2708 241 -2592
rect 243 -2593 244 -2583
rect 282 -2593 283 -2583
rect 292 -2708 293 -2592
rect 597 -2593 598 -2583
rect 660 -2708 661 -2592
rect 870 -2593 871 -2583
rect 898 -2593 899 -2583
rect 898 -2708 899 -2592
rect 898 -2593 899 -2583
rect 898 -2708 899 -2592
rect 915 -2708 916 -2592
rect 1353 -2593 1354 -2583
rect 1507 -2708 1508 -2592
rect 1535 -2593 1536 -2583
rect 1647 -2708 1648 -2592
rect 1654 -2593 1655 -2583
rect 79 -2708 80 -2594
rect 842 -2595 843 -2583
rect 947 -2708 948 -2594
rect 1244 -2708 1245 -2594
rect 1276 -2708 1277 -2594
rect 1304 -2595 1305 -2583
rect 1311 -2708 1312 -2594
rect 1388 -2595 1389 -2583
rect 1654 -2708 1655 -2594
rect 1776 -2708 1777 -2594
rect 121 -2708 122 -2596
rect 128 -2597 129 -2583
rect 149 -2597 150 -2583
rect 387 -2597 388 -2583
rect 457 -2597 458 -2583
rect 670 -2597 671 -2583
rect 695 -2597 696 -2583
rect 712 -2708 713 -2596
rect 737 -2597 738 -2583
rect 1486 -2597 1487 -2583
rect 68 -2708 69 -2598
rect 149 -2708 150 -2598
rect 156 -2599 157 -2583
rect 254 -2599 255 -2583
rect 261 -2599 262 -2583
rect 261 -2708 262 -2598
rect 261 -2599 262 -2583
rect 261 -2708 262 -2598
rect 275 -2599 276 -2583
rect 558 -2599 559 -2583
rect 642 -2708 643 -2598
rect 1535 -2708 1536 -2598
rect 86 -2601 87 -2583
rect 128 -2708 129 -2600
rect 142 -2601 143 -2583
rect 275 -2708 276 -2600
rect 282 -2708 283 -2600
rect 289 -2601 290 -2583
rect 296 -2601 297 -2583
rect 586 -2708 587 -2600
rect 681 -2601 682 -2583
rect 737 -2708 738 -2600
rect 758 -2601 759 -2583
rect 758 -2708 759 -2600
rect 758 -2601 759 -2583
rect 758 -2708 759 -2600
rect 765 -2601 766 -2583
rect 779 -2708 780 -2600
rect 842 -2708 843 -2600
rect 884 -2601 885 -2583
rect 968 -2601 969 -2583
rect 1430 -2601 1431 -2583
rect 1486 -2708 1487 -2600
rect 1542 -2601 1543 -2583
rect 86 -2708 87 -2602
rect 100 -2603 101 -2583
rect 103 -2603 104 -2583
rect 289 -2708 290 -2602
rect 296 -2708 297 -2602
rect 1017 -2603 1018 -2583
rect 1048 -2603 1049 -2583
rect 1290 -2603 1291 -2583
rect 1304 -2708 1305 -2602
rect 1360 -2603 1361 -2583
rect 1430 -2708 1431 -2602
rect 1444 -2603 1445 -2583
rect 1542 -2708 1543 -2602
rect 1570 -2603 1571 -2583
rect 37 -2605 38 -2583
rect 100 -2708 101 -2604
rect 142 -2708 143 -2604
rect 436 -2605 437 -2583
rect 453 -2605 454 -2583
rect 681 -2708 682 -2604
rect 695 -2708 696 -2604
rect 877 -2605 878 -2583
rect 905 -2605 906 -2583
rect 968 -2708 969 -2604
rect 971 -2605 972 -2583
rect 1703 -2605 1704 -2583
rect 37 -2708 38 -2606
rect 845 -2708 846 -2606
rect 856 -2607 857 -2583
rect 877 -2708 878 -2606
rect 905 -2708 906 -2606
rect 950 -2607 951 -2583
rect 989 -2607 990 -2583
rect 1038 -2607 1039 -2583
rect 1073 -2708 1074 -2606
rect 1094 -2607 1095 -2583
rect 1108 -2708 1109 -2606
rect 1143 -2607 1144 -2583
rect 1157 -2708 1158 -2606
rect 1220 -2607 1221 -2583
rect 1262 -2607 1263 -2583
rect 1388 -2708 1389 -2606
rect 1444 -2708 1445 -2606
rect 1458 -2607 1459 -2583
rect 1570 -2708 1571 -2606
rect 1598 -2607 1599 -2583
rect 1675 -2607 1676 -2583
rect 1703 -2708 1704 -2606
rect 156 -2708 157 -2608
rect 198 -2609 199 -2583
rect 205 -2609 206 -2583
rect 450 -2708 451 -2608
rect 492 -2609 493 -2583
rect 765 -2708 766 -2608
rect 775 -2708 776 -2608
rect 1374 -2708 1375 -2608
rect 1458 -2708 1459 -2608
rect 1514 -2609 1515 -2583
rect 1598 -2708 1599 -2608
rect 1619 -2609 1620 -2583
rect 1675 -2708 1676 -2608
rect 1717 -2609 1718 -2583
rect 159 -2611 160 -2583
rect 926 -2611 927 -2583
rect 940 -2611 941 -2583
rect 1143 -2708 1144 -2610
rect 1174 -2611 1175 -2583
rect 1332 -2611 1333 -2583
rect 1353 -2708 1354 -2610
rect 1409 -2611 1410 -2583
rect 1514 -2708 1515 -2610
rect 1699 -2611 1700 -2583
rect 1710 -2611 1711 -2583
rect 1717 -2708 1718 -2610
rect 170 -2613 171 -2583
rect 1248 -2613 1249 -2583
rect 1409 -2708 1410 -2612
rect 1605 -2613 1606 -2583
rect 1689 -2613 1690 -2583
rect 1710 -2708 1711 -2612
rect 170 -2708 171 -2614
rect 604 -2615 605 -2583
rect 702 -2615 703 -2583
rect 740 -2615 741 -2583
rect 856 -2708 857 -2614
rect 1052 -2615 1053 -2583
rect 1066 -2615 1067 -2583
rect 1332 -2708 1333 -2614
rect 1556 -2615 1557 -2583
rect 1605 -2708 1606 -2614
rect 1689 -2708 1690 -2614
rect 1766 -2615 1767 -2583
rect 173 -2617 174 -2583
rect 1101 -2617 1102 -2583
rect 1118 -2617 1119 -2583
rect 1591 -2708 1592 -2616
rect 177 -2619 178 -2583
rect 254 -2708 255 -2618
rect 303 -2619 304 -2583
rect 457 -2708 458 -2618
rect 492 -2708 493 -2618
rect 730 -2619 731 -2583
rect 828 -2708 829 -2618
rect 1766 -2708 1767 -2618
rect 23 -2621 24 -2583
rect 177 -2708 178 -2620
rect 184 -2621 185 -2583
rect 667 -2621 668 -2583
rect 702 -2708 703 -2620
rect 786 -2621 787 -2583
rect 870 -2708 871 -2620
rect 1052 -2708 1053 -2620
rect 1076 -2621 1077 -2583
rect 1185 -2621 1186 -2583
rect 1220 -2708 1221 -2620
rect 1318 -2621 1319 -2583
rect 1556 -2708 1557 -2620
rect 1584 -2621 1585 -2583
rect 184 -2708 185 -2622
rect 198 -2708 199 -2622
rect 205 -2708 206 -2622
rect 345 -2623 346 -2583
rect 387 -2708 388 -2622
rect 688 -2623 689 -2583
rect 709 -2623 710 -2583
rect 1206 -2623 1207 -2583
rect 1241 -2623 1242 -2583
rect 1262 -2708 1263 -2622
rect 1584 -2708 1585 -2622
rect 1612 -2623 1613 -2583
rect 226 -2625 227 -2583
rect 1020 -2708 1021 -2624
rect 1024 -2625 1025 -2583
rect 1038 -2708 1039 -2624
rect 1094 -2708 1095 -2624
rect 1150 -2625 1151 -2583
rect 1241 -2708 1242 -2624
rect 1367 -2625 1368 -2583
rect 1612 -2708 1613 -2624
rect 1626 -2625 1627 -2583
rect 30 -2627 31 -2583
rect 226 -2708 227 -2626
rect 303 -2708 304 -2626
rect 485 -2627 486 -2583
rect 513 -2627 514 -2583
rect 604 -2708 605 -2626
rect 646 -2627 647 -2583
rect 667 -2708 668 -2626
rect 723 -2627 724 -2583
rect 1360 -2708 1361 -2626
rect 1367 -2708 1368 -2626
rect 1493 -2627 1494 -2583
rect 1626 -2708 1627 -2626
rect 1633 -2627 1634 -2583
rect 30 -2708 31 -2628
rect 65 -2629 66 -2583
rect 310 -2629 311 -2583
rect 425 -2708 426 -2628
rect 436 -2708 437 -2628
rect 716 -2629 717 -2583
rect 730 -2708 731 -2628
rect 744 -2629 745 -2583
rect 786 -2708 787 -2628
rect 1171 -2629 1172 -2583
rect 1248 -2708 1249 -2628
rect 1321 -2708 1322 -2628
rect 1479 -2629 1480 -2583
rect 1493 -2708 1494 -2628
rect 1633 -2708 1634 -2628
rect 1731 -2629 1732 -2583
rect 58 -2631 59 -2583
rect 513 -2708 514 -2630
rect 520 -2631 521 -2583
rect 852 -2708 853 -2630
rect 912 -2631 913 -2583
rect 926 -2708 927 -2630
rect 933 -2631 934 -2583
rect 1206 -2708 1207 -2630
rect 1731 -2708 1732 -2630
rect 1745 -2631 1746 -2583
rect 58 -2708 59 -2632
rect 800 -2633 801 -2583
rect 835 -2633 836 -2583
rect 933 -2708 934 -2632
rect 940 -2708 941 -2632
rect 1395 -2633 1396 -2583
rect 1745 -2708 1746 -2632
rect 1752 -2633 1753 -2583
rect 110 -2635 111 -2583
rect 310 -2708 311 -2634
rect 317 -2635 318 -2583
rect 317 -2708 318 -2634
rect 317 -2635 318 -2583
rect 317 -2708 318 -2634
rect 338 -2635 339 -2583
rect 366 -2708 367 -2634
rect 380 -2635 381 -2583
rect 688 -2708 689 -2634
rect 716 -2708 717 -2634
rect 1318 -2708 1319 -2634
rect 1395 -2708 1396 -2634
rect 1416 -2635 1417 -2583
rect 1752 -2708 1753 -2634
rect 1759 -2635 1760 -2583
rect 135 -2637 136 -2583
rect 835 -2708 836 -2636
rect 919 -2637 920 -2583
rect 1185 -2708 1186 -2636
rect 1416 -2708 1417 -2636
rect 1472 -2637 1473 -2583
rect 1759 -2708 1760 -2636
rect 1773 -2637 1774 -2583
rect 135 -2708 136 -2638
rect 233 -2639 234 -2583
rect 338 -2708 339 -2638
rect 401 -2639 402 -2583
rect 408 -2639 409 -2583
rect 989 -2708 990 -2638
rect 996 -2708 997 -2638
rect 1010 -2639 1011 -2583
rect 1017 -2708 1018 -2638
rect 1682 -2639 1683 -2583
rect 72 -2641 73 -2583
rect 233 -2708 234 -2640
rect 345 -2708 346 -2640
rect 352 -2641 353 -2583
rect 359 -2641 360 -2583
rect 380 -2708 381 -2640
rect 394 -2641 395 -2583
rect 401 -2708 402 -2640
rect 422 -2641 423 -2583
rect 485 -2708 486 -2640
rect 520 -2708 521 -2640
rect 1661 -2641 1662 -2583
rect 72 -2708 73 -2642
rect 464 -2643 465 -2583
rect 523 -2708 524 -2642
rect 569 -2643 570 -2583
rect 646 -2708 647 -2642
rect 653 -2643 654 -2583
rect 674 -2643 675 -2583
rect 723 -2708 724 -2642
rect 800 -2708 801 -2642
rect 978 -2708 979 -2642
rect 1003 -2643 1004 -2583
rect 1066 -2708 1067 -2642
rect 1101 -2708 1102 -2642
rect 1164 -2643 1165 -2583
rect 1171 -2708 1172 -2642
rect 1297 -2643 1298 -2583
rect 1472 -2708 1473 -2642
rect 1521 -2643 1522 -2583
rect 152 -2645 153 -2583
rect 1661 -2708 1662 -2644
rect 201 -2708 202 -2646
rect 1479 -2708 1480 -2646
rect 1521 -2708 1522 -2646
rect 1549 -2647 1550 -2583
rect 268 -2649 269 -2583
rect 674 -2708 675 -2648
rect 891 -2649 892 -2583
rect 1010 -2708 1011 -2648
rect 1024 -2708 1025 -2648
rect 1080 -2649 1081 -2583
rect 1122 -2649 1123 -2583
rect 1136 -2649 1137 -2583
rect 1139 -2649 1140 -2583
rect 1738 -2708 1739 -2648
rect 268 -2708 269 -2650
rect 1160 -2651 1161 -2583
rect 1297 -2708 1298 -2650
rect 1325 -2651 1326 -2583
rect 1549 -2708 1550 -2650
rect 1577 -2651 1578 -2583
rect 324 -2653 325 -2583
rect 352 -2708 353 -2652
rect 359 -2708 360 -2652
rect 429 -2653 430 -2583
rect 464 -2708 465 -2652
rect 793 -2653 794 -2583
rect 821 -2653 822 -2583
rect 1136 -2708 1137 -2652
rect 1325 -2708 1326 -2652
rect 1619 -2708 1620 -2652
rect 324 -2708 325 -2654
rect 548 -2655 549 -2583
rect 569 -2708 570 -2654
rect 590 -2655 591 -2583
rect 625 -2655 626 -2583
rect 891 -2708 892 -2654
rect 912 -2708 913 -2654
rect 1080 -2708 1081 -2654
rect 1122 -2708 1123 -2654
rect 1178 -2655 1179 -2583
rect 1577 -2708 1578 -2654
rect 1741 -2655 1742 -2583
rect 163 -2657 164 -2583
rect 548 -2708 549 -2656
rect 590 -2708 591 -2656
rect 618 -2657 619 -2583
rect 625 -2708 626 -2656
rect 849 -2657 850 -2583
rect 954 -2657 955 -2583
rect 1003 -2708 1004 -2656
rect 1087 -2657 1088 -2583
rect 1178 -2708 1179 -2656
rect 163 -2708 164 -2658
rect 219 -2659 220 -2583
rect 373 -2659 374 -2583
rect 408 -2708 409 -2658
rect 415 -2659 416 -2583
rect 429 -2708 430 -2658
rect 506 -2659 507 -2583
rect 618 -2708 619 -2658
rect 632 -2659 633 -2583
rect 653 -2708 654 -2658
rect 772 -2659 773 -2583
rect 793 -2708 794 -2658
rect 814 -2659 815 -2583
rect 821 -2708 822 -2658
rect 849 -2708 850 -2658
rect 1682 -2708 1683 -2658
rect 219 -2708 220 -2660
rect 247 -2661 248 -2583
rect 331 -2661 332 -2583
rect 373 -2708 374 -2660
rect 394 -2708 395 -2660
rect 751 -2661 752 -2583
rect 814 -2708 815 -2660
rect 1199 -2661 1200 -2583
rect 93 -2663 94 -2583
rect 331 -2708 332 -2662
rect 415 -2708 416 -2662
rect 1195 -2663 1196 -2583
rect 1199 -2708 1200 -2662
rect 1213 -2663 1214 -2583
rect 93 -2708 94 -2664
rect 114 -2665 115 -2583
rect 191 -2665 192 -2583
rect 247 -2708 248 -2664
rect 478 -2665 479 -2583
rect 772 -2708 773 -2664
rect 863 -2665 864 -2583
rect 954 -2708 955 -2664
rect 961 -2665 962 -2583
rect 1164 -2708 1165 -2664
rect 1195 -2708 1196 -2664
rect 1500 -2665 1501 -2583
rect 114 -2708 115 -2666
rect 208 -2708 209 -2666
rect 471 -2667 472 -2583
rect 478 -2708 479 -2666
rect 506 -2708 507 -2666
rect 562 -2667 563 -2583
rect 597 -2708 598 -2666
rect 632 -2708 633 -2666
rect 635 -2708 636 -2666
rect 751 -2708 752 -2666
rect 961 -2708 962 -2666
rect 982 -2667 983 -2583
rect 1045 -2667 1046 -2583
rect 1087 -2708 1088 -2666
rect 1132 -2667 1133 -2583
rect 1668 -2667 1669 -2583
rect 191 -2708 192 -2668
rect 212 -2669 213 -2583
rect 471 -2708 472 -2668
rect 1150 -2708 1151 -2668
rect 1213 -2708 1214 -2668
rect 1801 -2669 1802 -2583
rect 51 -2671 52 -2583
rect 212 -2708 213 -2670
rect 499 -2671 500 -2583
rect 562 -2708 563 -2670
rect 975 -2671 976 -2583
rect 982 -2708 983 -2670
rect 1045 -2708 1046 -2670
rect 1346 -2671 1347 -2583
rect 1500 -2708 1501 -2670
rect 1787 -2671 1788 -2583
rect 1801 -2708 1802 -2670
rect 1808 -2671 1809 -2583
rect 51 -2708 52 -2672
rect 422 -2708 423 -2672
rect 499 -2708 500 -2672
rect 583 -2708 584 -2672
rect 975 -2708 976 -2672
rect 1031 -2673 1032 -2583
rect 1346 -2708 1347 -2672
rect 1381 -2673 1382 -2583
rect 1528 -2673 1529 -2583
rect 1668 -2708 1669 -2672
rect 1787 -2708 1788 -2672
rect 1794 -2673 1795 -2583
rect 1808 -2708 1809 -2672
rect 1815 -2673 1816 -2583
rect 527 -2675 528 -2583
rect 530 -2679 531 -2674
rect 534 -2675 535 -2583
rect 744 -2708 745 -2674
rect 1381 -2708 1382 -2674
rect 1402 -2675 1403 -2583
rect 1696 -2675 1697 -2583
rect 1794 -2708 1795 -2674
rect 527 -2708 528 -2676
rect 541 -2677 542 -2583
rect 555 -2677 556 -2583
rect 1696 -2708 1697 -2676
rect 541 -2708 542 -2678
rect 555 -2708 556 -2678
rect 576 -2679 577 -2583
rect 611 -2679 612 -2583
rect 1031 -2708 1032 -2678
rect 1192 -2679 1193 -2583
rect 1402 -2708 1403 -2678
rect 534 -2708 535 -2680
rect 1055 -2681 1056 -2583
rect 576 -2708 577 -2682
rect 1773 -2708 1774 -2682
rect 611 -2708 612 -2684
rect 1129 -2685 1130 -2583
rect 709 -2708 710 -2686
rect 1528 -2708 1529 -2686
rect 1055 -2708 1056 -2688
rect 1640 -2689 1641 -2583
rect 1059 -2708 1060 -2690
rect 1129 -2708 1130 -2690
rect 1269 -2691 1270 -2583
rect 1640 -2708 1641 -2690
rect 1234 -2693 1235 -2583
rect 1269 -2708 1270 -2692
rect 1227 -2695 1228 -2583
rect 1234 -2708 1235 -2694
rect 1227 -2708 1228 -2696
rect 1283 -2697 1284 -2583
rect 1255 -2699 1256 -2583
rect 1283 -2708 1284 -2698
rect 1255 -2708 1256 -2700
rect 1451 -2701 1452 -2583
rect 1423 -2703 1424 -2583
rect 1451 -2708 1452 -2702
rect 1423 -2708 1424 -2704
rect 1437 -2705 1438 -2583
rect 1192 -2708 1193 -2706
rect 1437 -2708 1438 -2706
rect 30 -2718 31 -2716
rect 712 -2718 713 -2716
rect 737 -2718 738 -2716
rect 772 -2829 773 -2717
rect 842 -2718 843 -2716
rect 1493 -2718 1494 -2716
rect 1769 -2718 1770 -2716
rect 1808 -2718 1809 -2716
rect 44 -2720 45 -2716
rect 68 -2720 69 -2716
rect 72 -2720 73 -2716
rect 642 -2720 643 -2716
rect 646 -2720 647 -2716
rect 646 -2829 647 -2719
rect 646 -2720 647 -2716
rect 646 -2829 647 -2719
rect 712 -2829 713 -2719
rect 1195 -2720 1196 -2716
rect 1290 -2829 1291 -2719
rect 1360 -2720 1361 -2716
rect 1433 -2829 1434 -2719
rect 1451 -2720 1452 -2716
rect 1493 -2829 1494 -2719
rect 1507 -2720 1508 -2716
rect 1780 -2720 1781 -2716
rect 1801 -2720 1802 -2716
rect 58 -2722 59 -2716
rect 72 -2829 73 -2721
rect 96 -2829 97 -2721
rect 142 -2722 143 -2716
rect 184 -2722 185 -2716
rect 184 -2829 185 -2721
rect 184 -2722 185 -2716
rect 184 -2829 185 -2721
rect 198 -2722 199 -2716
rect 1776 -2722 1777 -2716
rect 1783 -2722 1784 -2716
rect 1787 -2722 1788 -2716
rect 58 -2829 59 -2723
rect 590 -2724 591 -2716
rect 621 -2829 622 -2723
rect 737 -2829 738 -2723
rect 775 -2724 776 -2716
rect 1507 -2829 1508 -2723
rect 65 -2829 66 -2725
rect 1125 -2829 1126 -2725
rect 1129 -2726 1130 -2716
rect 1202 -2829 1203 -2725
rect 1297 -2726 1298 -2716
rect 1360 -2829 1361 -2725
rect 100 -2728 101 -2716
rect 103 -2738 104 -2727
rect 107 -2728 108 -2716
rect 523 -2728 524 -2716
rect 534 -2728 535 -2716
rect 887 -2728 888 -2716
rect 891 -2728 892 -2716
rect 978 -2728 979 -2716
rect 1003 -2728 1004 -2716
rect 1325 -2728 1326 -2716
rect 1328 -2728 1329 -2716
rect 1675 -2728 1676 -2716
rect 100 -2829 101 -2729
rect 156 -2730 157 -2716
rect 198 -2829 199 -2729
rect 208 -2730 209 -2716
rect 275 -2730 276 -2716
rect 275 -2829 276 -2729
rect 275 -2730 276 -2716
rect 275 -2829 276 -2729
rect 289 -2829 290 -2729
rect 373 -2730 374 -2716
rect 401 -2730 402 -2716
rect 422 -2730 423 -2716
rect 425 -2730 426 -2716
rect 604 -2829 605 -2729
rect 660 -2730 661 -2716
rect 891 -2829 892 -2729
rect 919 -2730 920 -2716
rect 1234 -2730 1235 -2716
rect 1297 -2829 1298 -2729
rect 1339 -2730 1340 -2716
rect 1346 -2730 1347 -2716
rect 1451 -2829 1452 -2729
rect 1675 -2829 1676 -2729
rect 1717 -2730 1718 -2716
rect 107 -2829 108 -2731
rect 443 -2732 444 -2716
rect 464 -2732 465 -2716
rect 1181 -2829 1182 -2731
rect 1318 -2732 1319 -2716
rect 1605 -2732 1606 -2716
rect 114 -2734 115 -2716
rect 114 -2829 115 -2733
rect 114 -2734 115 -2716
rect 114 -2829 115 -2733
rect 142 -2829 143 -2733
rect 667 -2734 668 -2716
rect 842 -2829 843 -2733
rect 856 -2734 857 -2716
rect 863 -2734 864 -2716
rect 1206 -2734 1207 -2716
rect 1318 -2829 1319 -2733
rect 1437 -2734 1438 -2716
rect 1605 -2829 1606 -2733
rect 1626 -2734 1627 -2716
rect 149 -2736 150 -2716
rect 156 -2829 157 -2735
rect 201 -2736 202 -2716
rect 261 -2736 262 -2716
rect 292 -2736 293 -2716
rect 513 -2736 514 -2716
rect 534 -2829 535 -2735
rect 744 -2736 745 -2716
rect 849 -2829 850 -2735
rect 1283 -2736 1284 -2716
rect 1325 -2829 1326 -2735
rect 1423 -2736 1424 -2716
rect 1437 -2829 1438 -2735
rect 1549 -2736 1550 -2716
rect 1626 -2829 1627 -2735
rect 1647 -2736 1648 -2716
rect 149 -2829 150 -2737
rect 205 -2829 206 -2737
rect 219 -2738 220 -2716
rect 226 -2738 227 -2716
rect 373 -2829 374 -2737
rect 436 -2738 437 -2716
rect 632 -2738 633 -2716
rect 660 -2829 661 -2737
rect 663 -2829 664 -2737
rect 667 -2829 668 -2737
rect 954 -2738 955 -2716
rect 1003 -2829 1004 -2737
rect 1069 -2829 1070 -2737
rect 1080 -2738 1081 -2716
rect 1241 -2738 1242 -2716
rect 1332 -2738 1333 -2716
rect 1773 -2738 1774 -2716
rect 128 -2740 129 -2716
rect 219 -2829 220 -2739
rect 226 -2829 227 -2739
rect 611 -2740 612 -2716
rect 632 -2829 633 -2739
rect 653 -2740 654 -2716
rect 705 -2829 706 -2739
rect 1332 -2829 1333 -2739
rect 1346 -2829 1347 -2739
rect 1353 -2740 1354 -2716
rect 1549 -2829 1550 -2739
rect 1584 -2740 1585 -2716
rect 1647 -2829 1648 -2739
rect 1682 -2740 1683 -2716
rect 1773 -2829 1774 -2739
rect 1794 -2740 1795 -2716
rect 79 -2742 80 -2716
rect 128 -2829 129 -2741
rect 170 -2742 171 -2716
rect 653 -2829 654 -2741
rect 716 -2742 717 -2716
rect 856 -2829 857 -2741
rect 863 -2829 864 -2741
rect 1213 -2742 1214 -2716
rect 1241 -2829 1242 -2741
rect 1388 -2742 1389 -2716
rect 1584 -2829 1585 -2741
rect 1612 -2742 1613 -2716
rect 1682 -2829 1683 -2741
rect 1724 -2742 1725 -2716
rect 61 -2744 62 -2716
rect 1213 -2829 1214 -2743
rect 1237 -2829 1238 -2743
rect 1612 -2829 1613 -2743
rect 79 -2829 80 -2745
rect 93 -2746 94 -2716
rect 170 -2829 171 -2745
rect 359 -2746 360 -2716
rect 436 -2829 437 -2745
rect 639 -2746 640 -2716
rect 716 -2829 717 -2745
rect 779 -2746 780 -2716
rect 852 -2829 853 -2745
rect 877 -2746 878 -2716
rect 884 -2746 885 -2716
rect 1164 -2746 1165 -2716
rect 1283 -2829 1284 -2745
rect 1724 -2829 1725 -2745
rect 37 -2748 38 -2716
rect 359 -2829 360 -2747
rect 443 -2829 444 -2747
rect 541 -2748 542 -2716
rect 562 -2748 563 -2716
rect 639 -2829 640 -2747
rect 695 -2748 696 -2716
rect 779 -2829 780 -2747
rect 877 -2829 878 -2747
rect 1321 -2748 1322 -2716
rect 1388 -2829 1389 -2747
rect 1430 -2748 1431 -2716
rect 37 -2829 38 -2749
rect 86 -2750 87 -2716
rect 261 -2829 262 -2749
rect 1353 -2829 1354 -2749
rect 9 -2752 10 -2716
rect 86 -2829 87 -2751
rect 303 -2752 304 -2716
rect 859 -2829 860 -2751
rect 884 -2829 885 -2751
rect 1062 -2752 1063 -2716
rect 1080 -2829 1081 -2751
rect 1094 -2752 1095 -2716
rect 1101 -2752 1102 -2716
rect 1101 -2829 1102 -2751
rect 1101 -2752 1102 -2716
rect 1101 -2829 1102 -2751
rect 1108 -2752 1109 -2716
rect 1108 -2829 1109 -2751
rect 1108 -2752 1109 -2716
rect 1108 -2829 1109 -2751
rect 1118 -2829 1119 -2751
rect 1661 -2752 1662 -2716
rect 44 -2829 45 -2753
rect 93 -2829 94 -2753
rect 303 -2829 304 -2753
rect 366 -2754 367 -2716
rect 464 -2829 465 -2753
rect 786 -2754 787 -2716
rect 919 -2829 920 -2753
rect 989 -2754 990 -2716
rect 1010 -2754 1011 -2716
rect 1052 -2754 1053 -2716
rect 1087 -2754 1088 -2716
rect 1342 -2829 1343 -2753
rect 1661 -2829 1662 -2753
rect 1752 -2754 1753 -2716
rect 268 -2756 269 -2716
rect 366 -2829 367 -2755
rect 478 -2756 479 -2716
rect 481 -2829 482 -2755
rect 513 -2829 514 -2755
rect 527 -2756 528 -2716
rect 541 -2829 542 -2755
rect 597 -2756 598 -2716
rect 611 -2829 612 -2755
rect 723 -2756 724 -2716
rect 744 -2829 745 -2755
rect 793 -2756 794 -2716
rect 940 -2756 941 -2716
rect 1206 -2829 1207 -2755
rect 1720 -2829 1721 -2755
rect 1752 -2829 1753 -2755
rect 135 -2758 136 -2716
rect 268 -2829 269 -2757
rect 331 -2758 332 -2716
rect 565 -2829 566 -2757
rect 569 -2758 570 -2716
rect 915 -2758 916 -2716
rect 940 -2829 941 -2757
rect 1153 -2758 1154 -2716
rect 1164 -2829 1165 -2757
rect 1199 -2758 1200 -2716
rect 135 -2829 136 -2759
rect 233 -2760 234 -2716
rect 310 -2760 311 -2716
rect 331 -2829 332 -2759
rect 338 -2760 339 -2716
rect 401 -2829 402 -2759
rect 527 -2829 528 -2759
rect 828 -2760 829 -2716
rect 954 -2829 955 -2759
rect 961 -2760 962 -2716
rect 982 -2760 983 -2716
rect 989 -2829 990 -2759
rect 1013 -2829 1014 -2759
rect 1423 -2829 1424 -2759
rect 51 -2762 52 -2716
rect 233 -2829 234 -2761
rect 310 -2829 311 -2761
rect 1010 -2829 1011 -2761
rect 1017 -2829 1018 -2761
rect 1759 -2762 1760 -2716
rect 51 -2829 52 -2763
rect 387 -2764 388 -2716
rect 562 -2829 563 -2763
rect 702 -2764 703 -2716
rect 786 -2829 787 -2763
rect 1045 -2764 1046 -2716
rect 1052 -2829 1053 -2763
rect 1073 -2764 1074 -2716
rect 1094 -2829 1095 -2763
rect 1570 -2764 1571 -2716
rect 1745 -2764 1746 -2716
rect 1759 -2829 1760 -2763
rect 324 -2766 325 -2716
rect 702 -2829 703 -2765
rect 866 -2766 867 -2716
rect 1570 -2829 1571 -2765
rect 324 -2829 325 -2767
rect 352 -2768 353 -2716
rect 355 -2829 356 -2767
rect 835 -2768 836 -2716
rect 961 -2829 962 -2767
rect 1143 -2768 1144 -2716
rect 1150 -2768 1151 -2716
rect 1689 -2768 1690 -2716
rect 338 -2829 339 -2769
rect 457 -2770 458 -2716
rect 569 -2829 570 -2769
rect 625 -2770 626 -2716
rect 695 -2829 696 -2769
rect 730 -2770 731 -2716
rect 821 -2770 822 -2716
rect 835 -2829 836 -2769
rect 982 -2829 983 -2769
rect 1178 -2770 1179 -2716
rect 1199 -2829 1200 -2769
rect 1514 -2770 1515 -2716
rect 1633 -2770 1634 -2716
rect 1689 -2829 1690 -2769
rect 345 -2772 346 -2716
rect 422 -2829 423 -2771
rect 457 -2829 458 -2771
rect 831 -2829 832 -2771
rect 1031 -2772 1032 -2716
rect 1045 -2829 1046 -2771
rect 1073 -2829 1074 -2771
rect 1276 -2772 1277 -2716
rect 1430 -2829 1431 -2771
rect 1745 -2829 1746 -2771
rect 345 -2829 346 -2773
rect 1059 -2774 1060 -2716
rect 1143 -2829 1144 -2773
rect 1248 -2774 1249 -2716
rect 1276 -2829 1277 -2773
rect 1311 -2774 1312 -2716
rect 1514 -2829 1515 -2773
rect 1542 -2774 1543 -2716
rect 1633 -2829 1634 -2773
rect 1654 -2774 1655 -2716
rect 380 -2776 381 -2716
rect 387 -2829 388 -2775
rect 499 -2776 500 -2716
rect 625 -2829 626 -2775
rect 751 -2776 752 -2716
rect 1248 -2829 1249 -2775
rect 1311 -2829 1312 -2775
rect 1458 -2776 1459 -2716
rect 1542 -2829 1543 -2775
rect 1556 -2776 1557 -2716
rect 380 -2829 381 -2777
rect 408 -2778 409 -2716
rect 478 -2829 479 -2777
rect 499 -2829 500 -2777
rect 583 -2778 584 -2716
rect 1374 -2778 1375 -2716
rect 1458 -2829 1459 -2777
rect 1472 -2778 1473 -2716
rect 1556 -2829 1557 -2777
rect 1696 -2778 1697 -2716
rect 408 -2829 409 -2779
rect 506 -2780 507 -2716
rect 583 -2829 584 -2779
rect 723 -2829 724 -2779
rect 807 -2780 808 -2716
rect 821 -2829 822 -2779
rect 996 -2780 997 -2716
rect 1059 -2829 1060 -2779
rect 1129 -2829 1130 -2779
rect 1654 -2829 1655 -2779
rect 1696 -2829 1697 -2779
rect 1731 -2780 1732 -2716
rect 415 -2782 416 -2716
rect 506 -2829 507 -2781
rect 520 -2782 521 -2716
rect 807 -2829 808 -2781
rect 1031 -2829 1032 -2781
rect 1479 -2782 1480 -2716
rect 1500 -2782 1501 -2716
rect 1731 -2829 1732 -2781
rect 415 -2829 416 -2783
rect 429 -2784 430 -2716
rect 520 -2829 521 -2783
rect 576 -2784 577 -2716
rect 590 -2829 591 -2783
rect 1717 -2829 1718 -2783
rect 247 -2786 248 -2716
rect 576 -2829 577 -2785
rect 597 -2829 598 -2785
rect 688 -2786 689 -2716
rect 1150 -2829 1151 -2785
rect 1171 -2786 1172 -2716
rect 1178 -2829 1179 -2785
rect 1563 -2786 1564 -2716
rect 247 -2829 248 -2787
rect 471 -2788 472 -2716
rect 548 -2788 549 -2716
rect 996 -2829 997 -2787
rect 1171 -2829 1172 -2787
rect 1227 -2788 1228 -2716
rect 1374 -2829 1375 -2787
rect 1766 -2788 1767 -2716
rect 177 -2790 178 -2716
rect 548 -2829 549 -2789
rect 607 -2790 608 -2716
rect 793 -2829 794 -2789
rect 947 -2790 948 -2716
rect 1227 -2829 1228 -2789
rect 1402 -2790 1403 -2716
rect 1766 -2829 1767 -2789
rect 121 -2792 122 -2716
rect 177 -2829 178 -2791
rect 296 -2792 297 -2716
rect 688 -2829 689 -2791
rect 1402 -2829 1403 -2791
rect 1591 -2792 1592 -2716
rect 121 -2829 122 -2793
rect 240 -2794 241 -2716
rect 296 -2829 297 -2793
rect 681 -2794 682 -2716
rect 1465 -2794 1466 -2716
rect 1563 -2829 1564 -2793
rect 1591 -2829 1592 -2793
rect 1619 -2794 1620 -2716
rect 212 -2796 213 -2716
rect 240 -2829 241 -2795
rect 317 -2796 318 -2716
rect 429 -2829 430 -2795
rect 471 -2829 472 -2795
rect 485 -2796 486 -2716
rect 618 -2796 619 -2716
rect 730 -2829 731 -2795
rect 1465 -2829 1466 -2795
rect 1486 -2796 1487 -2716
rect 1619 -2829 1620 -2795
rect 1703 -2796 1704 -2716
rect 212 -2829 213 -2797
rect 282 -2798 283 -2716
rect 317 -2829 318 -2797
rect 1185 -2798 1186 -2716
rect 1472 -2829 1473 -2797
rect 1521 -2798 1522 -2716
rect 1703 -2829 1704 -2797
rect 1738 -2798 1739 -2716
rect 254 -2800 255 -2716
rect 282 -2829 283 -2799
rect 485 -2829 486 -2799
rect 555 -2800 556 -2716
rect 618 -2829 619 -2799
rect 751 -2829 752 -2799
rect 912 -2800 913 -2716
rect 1521 -2829 1522 -2799
rect 163 -2802 164 -2716
rect 555 -2829 556 -2801
rect 635 -2802 636 -2716
rect 947 -2829 948 -2801
rect 975 -2802 976 -2716
rect 1486 -2829 1487 -2801
rect 163 -2829 164 -2803
rect 191 -2804 192 -2716
rect 254 -2829 255 -2803
rect 870 -2804 871 -2716
rect 912 -2829 913 -2803
rect 926 -2804 927 -2716
rect 975 -2829 976 -2803
rect 1038 -2804 1039 -2716
rect 1185 -2829 1186 -2803
rect 1262 -2804 1263 -2716
rect 1381 -2804 1382 -2716
rect 1738 -2829 1739 -2803
rect 191 -2829 192 -2805
rect 492 -2806 493 -2716
rect 681 -2829 682 -2805
rect 765 -2806 766 -2716
rect 926 -2829 927 -2805
rect 968 -2806 969 -2716
rect 1038 -2829 1039 -2805
rect 1115 -2806 1116 -2716
rect 1255 -2806 1256 -2716
rect 1262 -2829 1263 -2805
rect 1381 -2829 1382 -2805
rect 1444 -2806 1445 -2716
rect 1479 -2829 1480 -2805
rect 1528 -2806 1529 -2716
rect 450 -2808 451 -2716
rect 492 -2829 493 -2807
rect 709 -2808 710 -2716
rect 765 -2829 766 -2807
rect 968 -2829 969 -2807
rect 1024 -2808 1025 -2716
rect 1087 -2829 1088 -2807
rect 1115 -2829 1116 -2807
rect 1255 -2829 1256 -2807
rect 1304 -2808 1305 -2716
rect 1444 -2829 1445 -2807
rect 1640 -2808 1641 -2716
rect 394 -2810 395 -2716
rect 450 -2829 451 -2809
rect 709 -2829 710 -2809
rect 845 -2810 846 -2716
rect 1024 -2829 1025 -2809
rect 1066 -2810 1067 -2716
rect 1304 -2829 1305 -2809
rect 1367 -2810 1368 -2716
rect 1528 -2829 1529 -2809
rect 1577 -2810 1578 -2716
rect 1640 -2829 1641 -2809
rect 1668 -2810 1669 -2716
rect 394 -2829 395 -2811
rect 674 -2812 675 -2716
rect 1066 -2829 1067 -2811
rect 1220 -2812 1221 -2716
rect 1367 -2829 1368 -2811
rect 1395 -2812 1396 -2716
rect 1577 -2829 1578 -2811
rect 1598 -2812 1599 -2716
rect 1668 -2829 1669 -2811
rect 1710 -2812 1711 -2716
rect 674 -2829 675 -2813
rect 758 -2814 759 -2716
rect 1020 -2814 1021 -2716
rect 1395 -2829 1396 -2813
rect 1500 -2829 1501 -2813
rect 1710 -2829 1711 -2813
rect 758 -2829 759 -2815
rect 800 -2816 801 -2716
rect 1020 -2829 1021 -2815
rect 1192 -2816 1193 -2716
rect 1220 -2829 1221 -2815
rect 1269 -2816 1270 -2716
rect 1535 -2816 1536 -2716
rect 1598 -2829 1599 -2815
rect 800 -2829 801 -2817
rect 933 -2818 934 -2716
rect 1136 -2818 1137 -2716
rect 1269 -2829 1270 -2817
rect 1409 -2818 1410 -2716
rect 1535 -2829 1536 -2817
rect 814 -2820 815 -2716
rect 933 -2829 934 -2819
rect 1136 -2829 1137 -2819
rect 1244 -2820 1245 -2716
rect 1409 -2829 1410 -2819
rect 1416 -2820 1417 -2716
rect 814 -2829 815 -2821
rect 1713 -2829 1714 -2821
rect 905 -2824 906 -2716
rect 1416 -2829 1417 -2823
rect 898 -2826 899 -2716
rect 905 -2829 906 -2825
rect 1157 -2826 1158 -2716
rect 1192 -2829 1193 -2825
rect 733 -2829 734 -2827
rect 898 -2829 899 -2827
rect 1122 -2828 1123 -2716
rect 1157 -2829 1158 -2827
rect 23 -2948 24 -2838
rect 289 -2839 290 -2837
rect 331 -2839 332 -2837
rect 583 -2839 584 -2837
rect 621 -2839 622 -2837
rect 1031 -2839 1032 -2837
rect 1097 -2948 1098 -2838
rect 1668 -2839 1669 -2837
rect 1713 -2839 1714 -2837
rect 1759 -2839 1760 -2837
rect 44 -2841 45 -2837
rect 558 -2841 559 -2837
rect 656 -2948 657 -2840
rect 1416 -2841 1417 -2837
rect 1433 -2841 1434 -2837
rect 1689 -2841 1690 -2837
rect 1717 -2841 1718 -2837
rect 1773 -2841 1774 -2837
rect 79 -2843 80 -2837
rect 583 -2948 584 -2842
rect 660 -2843 661 -2837
rect 1248 -2843 1249 -2837
rect 1283 -2843 1284 -2837
rect 1675 -2843 1676 -2837
rect 1720 -2843 1721 -2837
rect 1766 -2843 1767 -2837
rect 93 -2845 94 -2837
rect 1248 -2948 1249 -2844
rect 1339 -2948 1340 -2844
rect 1612 -2845 1613 -2837
rect 1654 -2845 1655 -2837
rect 1675 -2948 1676 -2844
rect 1727 -2845 1728 -2837
rect 1752 -2845 1753 -2837
rect 93 -2948 94 -2846
rect 121 -2847 122 -2837
rect 128 -2847 129 -2837
rect 828 -2847 829 -2837
rect 859 -2847 860 -2837
rect 1696 -2847 1697 -2837
rect 96 -2849 97 -2837
rect 705 -2849 706 -2837
rect 712 -2849 713 -2837
rect 786 -2849 787 -2837
rect 824 -2948 825 -2848
rect 1507 -2849 1508 -2837
rect 1549 -2849 1550 -2837
rect 1549 -2948 1550 -2848
rect 1549 -2849 1550 -2837
rect 1549 -2948 1550 -2848
rect 1598 -2849 1599 -2837
rect 1696 -2948 1697 -2848
rect 100 -2851 101 -2837
rect 618 -2851 619 -2837
rect 681 -2851 682 -2837
rect 996 -2948 997 -2850
rect 1013 -2851 1014 -2837
rect 1388 -2851 1389 -2837
rect 1465 -2851 1466 -2837
rect 1507 -2948 1508 -2850
rect 1591 -2851 1592 -2837
rect 1598 -2948 1599 -2850
rect 1647 -2851 1648 -2837
rect 1654 -2948 1655 -2850
rect 37 -2853 38 -2837
rect 681 -2948 682 -2852
rect 730 -2948 731 -2852
rect 877 -2853 878 -2837
rect 915 -2948 916 -2852
rect 1332 -2853 1333 -2837
rect 1342 -2853 1343 -2837
rect 1563 -2853 1564 -2837
rect 1640 -2853 1641 -2837
rect 1647 -2948 1648 -2852
rect 51 -2855 52 -2837
rect 100 -2948 101 -2854
rect 107 -2855 108 -2837
rect 856 -2855 857 -2837
rect 870 -2855 871 -2837
rect 905 -2855 906 -2837
rect 947 -2855 948 -2837
rect 1017 -2948 1018 -2854
rect 1024 -2855 1025 -2837
rect 1129 -2855 1130 -2837
rect 1150 -2855 1151 -2837
rect 1283 -2948 1284 -2854
rect 1353 -2855 1354 -2837
rect 1682 -2855 1683 -2837
rect 51 -2948 52 -2856
rect 72 -2857 73 -2837
rect 107 -2948 108 -2856
rect 1157 -2857 1158 -2837
rect 1178 -2857 1179 -2837
rect 1703 -2857 1704 -2837
rect 72 -2948 73 -2858
rect 324 -2859 325 -2837
rect 359 -2859 360 -2837
rect 709 -2948 710 -2858
rect 765 -2859 766 -2837
rect 856 -2948 857 -2858
rect 877 -2948 878 -2858
rect 1010 -2859 1011 -2837
rect 1024 -2948 1025 -2858
rect 1514 -2859 1515 -2837
rect 1661 -2859 1662 -2837
rect 1682 -2948 1683 -2858
rect 1703 -2948 1704 -2858
rect 1724 -2859 1725 -2837
rect 121 -2948 122 -2860
rect 191 -2861 192 -2837
rect 226 -2861 227 -2837
rect 352 -2948 353 -2860
rect 366 -2861 367 -2837
rect 481 -2861 482 -2837
rect 499 -2861 500 -2837
rect 499 -2948 500 -2860
rect 499 -2861 500 -2837
rect 499 -2948 500 -2860
rect 520 -2861 521 -2837
rect 1055 -2948 1056 -2860
rect 1101 -2861 1102 -2837
rect 1150 -2948 1151 -2860
rect 1199 -2861 1200 -2837
rect 1276 -2861 1277 -2837
rect 1353 -2948 1354 -2860
rect 1374 -2861 1375 -2837
rect 1381 -2861 1382 -2837
rect 1416 -2948 1417 -2860
rect 1444 -2861 1445 -2837
rect 1591 -2948 1592 -2860
rect 1640 -2948 1641 -2860
rect 1661 -2948 1662 -2860
rect 65 -2863 66 -2837
rect 520 -2948 521 -2862
rect 555 -2863 556 -2837
rect 1045 -2863 1046 -2837
rect 1066 -2863 1067 -2837
rect 1101 -2948 1102 -2862
rect 1115 -2863 1116 -2837
rect 1164 -2863 1165 -2837
rect 1202 -2863 1203 -2837
rect 1451 -2863 1452 -2837
rect 1514 -2948 1515 -2862
rect 1528 -2863 1529 -2837
rect 65 -2948 66 -2864
rect 261 -2865 262 -2837
rect 275 -2865 276 -2837
rect 355 -2865 356 -2837
rect 366 -2948 367 -2864
rect 380 -2865 381 -2837
rect 429 -2865 430 -2837
rect 432 -2889 433 -2864
rect 464 -2865 465 -2837
rect 1178 -2948 1179 -2864
rect 1227 -2865 1228 -2837
rect 1689 -2948 1690 -2864
rect 128 -2948 129 -2866
rect 229 -2948 230 -2866
rect 247 -2867 248 -2837
rect 999 -2867 1000 -2837
rect 1066 -2948 1067 -2866
rect 1234 -2867 1235 -2837
rect 1237 -2867 1238 -2837
rect 1500 -2867 1501 -2837
rect 135 -2869 136 -2837
rect 411 -2948 412 -2868
rect 429 -2948 430 -2868
rect 541 -2869 542 -2837
rect 555 -2948 556 -2868
rect 646 -2869 647 -2837
rect 674 -2869 675 -2837
rect 1115 -2948 1116 -2868
rect 1125 -2869 1126 -2837
rect 1542 -2869 1543 -2837
rect 142 -2871 143 -2837
rect 702 -2948 703 -2870
rect 737 -2871 738 -2837
rect 765 -2948 766 -2870
rect 779 -2871 780 -2837
rect 947 -2948 948 -2870
rect 954 -2871 955 -2837
rect 954 -2948 955 -2870
rect 954 -2871 955 -2837
rect 954 -2948 955 -2870
rect 968 -2871 969 -2837
rect 1045 -2948 1046 -2870
rect 1136 -2871 1137 -2837
rect 1276 -2948 1277 -2870
rect 1311 -2871 1312 -2837
rect 1451 -2948 1452 -2870
rect 1500 -2948 1501 -2870
rect 1521 -2871 1522 -2837
rect 1535 -2871 1536 -2837
rect 1542 -2948 1543 -2870
rect 86 -2873 87 -2837
rect 142 -2948 143 -2872
rect 145 -2948 146 -2872
rect 1612 -2948 1613 -2872
rect 86 -2948 87 -2874
rect 114 -2875 115 -2837
rect 170 -2875 171 -2837
rect 586 -2875 587 -2837
rect 604 -2875 605 -2837
rect 1129 -2948 1130 -2874
rect 1164 -2948 1165 -2874
rect 1171 -2875 1172 -2837
rect 1227 -2948 1228 -2874
rect 1731 -2875 1732 -2837
rect 58 -2877 59 -2837
rect 114 -2948 115 -2876
rect 156 -2877 157 -2837
rect 170 -2948 171 -2876
rect 226 -2948 227 -2876
rect 467 -2948 468 -2876
rect 471 -2877 472 -2837
rect 471 -2948 472 -2876
rect 471 -2877 472 -2837
rect 471 -2948 472 -2876
rect 562 -2877 563 -2837
rect 1563 -2948 1564 -2876
rect 58 -2948 59 -2878
rect 782 -2948 783 -2878
rect 786 -2948 787 -2878
rect 1027 -2948 1028 -2878
rect 1171 -2948 1172 -2878
rect 1395 -2879 1396 -2837
rect 1437 -2879 1438 -2837
rect 1528 -2948 1529 -2878
rect 156 -2948 157 -2880
rect 184 -2881 185 -2837
rect 240 -2881 241 -2837
rect 247 -2948 248 -2880
rect 254 -2881 255 -2837
rect 866 -2948 867 -2880
rect 971 -2948 972 -2880
rect 1297 -2881 1298 -2837
rect 1311 -2948 1312 -2880
rect 1710 -2881 1711 -2837
rect 149 -2883 150 -2837
rect 254 -2948 255 -2882
rect 261 -2948 262 -2882
rect 373 -2883 374 -2837
rect 380 -2948 381 -2882
rect 565 -2883 566 -2837
rect 576 -2883 577 -2837
rect 618 -2948 619 -2882
rect 646 -2948 647 -2882
rect 807 -2883 808 -2837
rect 821 -2883 822 -2837
rect 870 -2948 871 -2882
rect 982 -2883 983 -2837
rect 1136 -2948 1137 -2882
rect 1234 -2948 1235 -2882
rect 1304 -2883 1305 -2837
rect 1318 -2883 1319 -2837
rect 1395 -2948 1396 -2882
rect 1423 -2883 1424 -2837
rect 1437 -2948 1438 -2882
rect 1444 -2948 1445 -2882
rect 1577 -2883 1578 -2837
rect 149 -2948 150 -2884
rect 338 -2885 339 -2837
rect 373 -2948 374 -2884
rect 387 -2885 388 -2837
rect 394 -2885 395 -2837
rect 464 -2948 465 -2884
rect 562 -2948 563 -2884
rect 569 -2885 570 -2837
rect 576 -2948 577 -2884
rect 849 -2885 850 -2837
rect 898 -2885 899 -2837
rect 982 -2948 983 -2884
rect 989 -2885 990 -2837
rect 1010 -2948 1011 -2884
rect 1255 -2885 1256 -2837
rect 1297 -2948 1298 -2884
rect 1318 -2948 1319 -2884
rect 1738 -2885 1739 -2837
rect 184 -2948 185 -2886
rect 625 -2887 626 -2837
rect 667 -2887 668 -2837
rect 898 -2948 899 -2886
rect 933 -2887 934 -2837
rect 1423 -2948 1424 -2886
rect 1479 -2887 1480 -2837
rect 1521 -2948 1522 -2886
rect 1570 -2887 1571 -2837
rect 1577 -2948 1578 -2886
rect 233 -2889 234 -2837
rect 387 -2948 388 -2888
rect 394 -2948 395 -2888
rect 422 -2889 423 -2837
rect 541 -2948 542 -2888
rect 590 -2889 591 -2837
rect 604 -2948 605 -2888
rect 625 -2948 626 -2888
rect 873 -2889 874 -2837
rect 1143 -2889 1144 -2837
rect 1255 -2948 1256 -2888
rect 1262 -2889 1263 -2837
rect 1388 -2948 1389 -2888
rect 1458 -2889 1459 -2837
rect 1479 -2948 1480 -2888
rect 1486 -2889 1487 -2837
rect 1535 -2948 1536 -2888
rect 1570 -2948 1571 -2888
rect 1584 -2889 1585 -2837
rect 233 -2948 234 -2890
rect 1122 -2891 1123 -2837
rect 1185 -2891 1186 -2837
rect 1262 -2948 1263 -2890
rect 1269 -2891 1270 -2837
rect 1304 -2948 1305 -2890
rect 1325 -2891 1326 -2837
rect 1381 -2948 1382 -2890
rect 1409 -2891 1410 -2837
rect 1584 -2948 1585 -2890
rect 240 -2948 241 -2892
rect 268 -2893 269 -2837
rect 275 -2948 276 -2892
rect 814 -2893 815 -2837
rect 828 -2948 829 -2892
rect 835 -2893 836 -2837
rect 849 -2948 850 -2892
rect 1360 -2893 1361 -2837
rect 1367 -2893 1368 -2837
rect 1374 -2948 1375 -2892
rect 1472 -2893 1473 -2837
rect 1486 -2948 1487 -2892
rect 268 -2948 269 -2894
rect 639 -2895 640 -2837
rect 653 -2895 654 -2837
rect 1143 -2948 1144 -2894
rect 1185 -2948 1186 -2894
rect 1192 -2895 1193 -2837
rect 1213 -2895 1214 -2837
rect 1360 -2948 1361 -2894
rect 1472 -2948 1473 -2894
rect 1493 -2895 1494 -2837
rect 282 -2897 283 -2837
rect 359 -2948 360 -2896
rect 415 -2897 416 -2837
rect 422 -2948 423 -2896
rect 439 -2948 440 -2896
rect 1409 -2948 1410 -2896
rect 198 -2899 199 -2837
rect 415 -2948 416 -2898
rect 527 -2899 528 -2837
rect 569 -2948 570 -2898
rect 590 -2948 591 -2898
rect 716 -2899 717 -2837
rect 737 -2948 738 -2898
rect 940 -2899 941 -2837
rect 1059 -2899 1060 -2837
rect 1192 -2948 1193 -2898
rect 1220 -2899 1221 -2837
rect 1269 -2948 1270 -2898
rect 1325 -2948 1326 -2898
rect 1346 -2899 1347 -2837
rect 1356 -2899 1357 -2837
rect 1619 -2899 1620 -2837
rect 110 -2948 111 -2900
rect 716 -2948 717 -2900
rect 751 -2901 752 -2837
rect 933 -2948 934 -2900
rect 1052 -2901 1053 -2837
rect 1059 -2948 1060 -2900
rect 1069 -2901 1070 -2837
rect 1458 -2948 1459 -2900
rect 198 -2948 199 -2902
rect 205 -2903 206 -2837
rect 212 -2903 213 -2837
rect 282 -2948 283 -2902
rect 289 -2948 290 -2902
rect 310 -2903 311 -2837
rect 317 -2903 318 -2837
rect 989 -2948 990 -2902
rect 1052 -2948 1053 -2902
rect 1556 -2903 1557 -2837
rect 163 -2905 164 -2837
rect 205 -2948 206 -2904
rect 212 -2948 213 -2904
rect 1286 -2905 1287 -2837
rect 1290 -2905 1291 -2837
rect 1346 -2948 1347 -2904
rect 1402 -2905 1403 -2837
rect 1556 -2948 1557 -2904
rect 163 -2948 164 -2906
rect 1157 -2948 1158 -2906
rect 1206 -2907 1207 -2837
rect 1619 -2948 1620 -2906
rect 303 -2909 304 -2837
rect 317 -2948 318 -2908
rect 324 -2948 325 -2908
rect 401 -2909 402 -2837
rect 506 -2909 507 -2837
rect 527 -2948 528 -2908
rect 653 -2948 654 -2908
rect 1668 -2948 1669 -2908
rect 208 -2948 209 -2910
rect 303 -2948 304 -2910
rect 310 -2948 311 -2910
rect 457 -2911 458 -2837
rect 506 -2948 507 -2910
rect 597 -2911 598 -2837
rect 663 -2911 664 -2837
rect 814 -2948 815 -2910
rect 835 -2948 836 -2910
rect 1087 -2911 1088 -2837
rect 1094 -2911 1095 -2837
rect 1493 -2948 1494 -2910
rect 219 -2913 220 -2837
rect 457 -2948 458 -2912
rect 667 -2948 668 -2912
rect 1031 -2948 1032 -2912
rect 1073 -2913 1074 -2837
rect 1290 -2948 1291 -2912
rect 1402 -2948 1403 -2912
rect 1745 -2913 1746 -2837
rect 219 -2948 220 -2914
rect 968 -2948 969 -2914
rect 1038 -2915 1039 -2837
rect 1073 -2948 1074 -2914
rect 1080 -2915 1081 -2837
rect 1122 -2948 1123 -2914
rect 1241 -2915 1242 -2837
rect 1367 -2948 1368 -2914
rect 338 -2948 339 -2916
rect 408 -2917 409 -2837
rect 436 -2917 437 -2837
rect 597 -2948 598 -2916
rect 674 -2948 675 -2916
rect 852 -2917 853 -2837
rect 891 -2917 892 -2837
rect 1213 -2948 1214 -2916
rect 191 -2948 192 -2918
rect 436 -2948 437 -2918
rect 688 -2919 689 -2837
rect 751 -2948 752 -2918
rect 800 -2919 801 -2837
rect 905 -2948 906 -2918
rect 961 -2919 962 -2837
rect 1206 -2948 1207 -2918
rect 331 -2948 332 -2920
rect 852 -2948 853 -2920
rect 926 -2921 927 -2837
rect 961 -2948 962 -2920
rect 975 -2921 976 -2837
rect 1038 -2948 1039 -2920
rect 1108 -2921 1109 -2837
rect 1220 -2948 1221 -2920
rect 345 -2923 346 -2837
rect 639 -2948 640 -2922
rect 688 -2948 689 -2922
rect 1020 -2923 1021 -2837
rect 1108 -2948 1109 -2922
rect 1430 -2923 1431 -2837
rect 177 -2925 178 -2837
rect 345 -2948 346 -2924
rect 401 -2948 402 -2924
rect 450 -2925 451 -2837
rect 695 -2925 696 -2837
rect 800 -2948 801 -2924
rect 807 -2948 808 -2924
rect 884 -2925 885 -2837
rect 919 -2925 920 -2837
rect 975 -2948 976 -2924
rect 1003 -2925 1004 -2837
rect 1080 -2948 1081 -2924
rect 1430 -2948 1431 -2924
rect 1605 -2925 1606 -2837
rect 177 -2948 178 -2926
rect 485 -2927 486 -2837
rect 534 -2927 535 -2837
rect 695 -2948 696 -2926
rect 723 -2927 724 -2837
rect 1087 -2948 1088 -2926
rect 1605 -2948 1606 -2926
rect 1626 -2927 1627 -2837
rect 443 -2929 444 -2837
rect 450 -2948 451 -2928
rect 485 -2948 486 -2928
rect 537 -2948 538 -2928
rect 723 -2948 724 -2928
rect 758 -2929 759 -2837
rect 793 -2929 794 -2837
rect 919 -2948 920 -2928
rect 926 -2948 927 -2928
rect 1202 -2948 1203 -2928
rect 1626 -2948 1627 -2928
rect 1633 -2929 1634 -2837
rect 443 -2948 444 -2930
rect 513 -2931 514 -2837
rect 733 -2931 734 -2837
rect 1633 -2948 1634 -2930
rect 478 -2933 479 -2837
rect 513 -2948 514 -2932
rect 744 -2933 745 -2837
rect 793 -2948 794 -2932
rect 842 -2933 843 -2837
rect 891 -2948 892 -2932
rect 478 -2948 479 -2934
rect 943 -2948 944 -2934
rect 492 -2937 493 -2837
rect 534 -2948 535 -2936
rect 611 -2937 612 -2837
rect 744 -2948 745 -2936
rect 758 -2948 759 -2936
rect 772 -2937 773 -2837
rect 863 -2937 864 -2837
rect 1003 -2948 1004 -2936
rect 492 -2948 493 -2938
rect 660 -2948 661 -2938
rect 663 -2948 664 -2938
rect 842 -2948 843 -2938
rect 863 -2948 864 -2938
rect 1241 -2948 1242 -2938
rect 548 -2941 549 -2837
rect 772 -2948 773 -2940
rect 884 -2948 885 -2940
rect 912 -2941 913 -2837
rect 82 -2948 83 -2942
rect 548 -2948 549 -2942
rect 611 -2948 612 -2942
rect 632 -2943 633 -2837
rect 912 -2948 913 -2942
rect 1465 -2948 1466 -2942
rect 296 -2945 297 -2837
rect 632 -2948 633 -2944
rect 166 -2948 167 -2946
rect 296 -2948 297 -2946
rect 30 -3075 31 -2957
rect 93 -2958 94 -2956
rect 100 -2958 101 -2956
rect 436 -3075 437 -2957
rect 439 -2958 440 -2956
rect 814 -2958 815 -2956
rect 821 -3075 822 -2957
rect 856 -2958 857 -2956
rect 863 -2958 864 -2956
rect 1584 -2958 1585 -2956
rect 1640 -2958 1641 -2956
rect 1696 -2958 1697 -2956
rect 37 -3075 38 -2959
rect 289 -2960 290 -2956
rect 303 -2960 304 -2956
rect 306 -3022 307 -2959
rect 369 -3075 370 -2959
rect 453 -3075 454 -2959
rect 541 -2960 542 -2956
rect 653 -2960 654 -2956
rect 663 -2960 664 -2956
rect 1213 -2960 1214 -2956
rect 1332 -2960 1333 -2956
rect 1507 -2960 1508 -2956
rect 1577 -2960 1578 -2956
rect 1703 -2960 1704 -2956
rect 44 -3075 45 -2961
rect 394 -2962 395 -2956
rect 450 -2962 451 -2956
rect 541 -3075 542 -2961
rect 548 -2962 549 -2956
rect 814 -3075 815 -2961
rect 842 -2962 843 -2956
rect 1024 -2962 1025 -2956
rect 1027 -2962 1028 -2956
rect 1689 -2962 1690 -2956
rect 23 -2964 24 -2956
rect 450 -3075 451 -2963
rect 499 -2964 500 -2956
rect 548 -3075 549 -2963
rect 611 -2964 612 -2956
rect 653 -3075 654 -2963
rect 674 -2964 675 -2956
rect 978 -3075 979 -2963
rect 1020 -3075 1021 -2963
rect 1220 -2964 1221 -2956
rect 1332 -3075 1333 -2963
rect 1381 -2964 1382 -2956
rect 1458 -2964 1459 -2956
rect 1640 -3075 1641 -2963
rect 72 -2966 73 -2956
rect 411 -2966 412 -2956
rect 499 -3075 500 -2965
rect 688 -2966 689 -2956
rect 740 -3075 741 -2965
rect 1143 -2966 1144 -2956
rect 1171 -2966 1172 -2956
rect 1381 -3075 1382 -2965
rect 1458 -3075 1459 -2965
rect 1465 -2966 1466 -2956
rect 1577 -3075 1578 -2965
rect 1605 -2966 1606 -2956
rect 51 -2968 52 -2956
rect 72 -3075 73 -2967
rect 79 -2968 80 -2956
rect 457 -2968 458 -2956
rect 569 -2968 570 -2956
rect 611 -3075 612 -2967
rect 618 -2968 619 -2956
rect 842 -3075 843 -2967
rect 849 -2968 850 -2956
rect 1115 -2968 1116 -2956
rect 1150 -2968 1151 -2956
rect 1171 -3075 1172 -2967
rect 1199 -2968 1200 -2956
rect 1528 -2968 1529 -2956
rect 1605 -3075 1606 -2967
rect 1647 -2968 1648 -2956
rect 51 -3075 52 -2969
rect 212 -2970 213 -2956
rect 219 -2970 220 -2956
rect 996 -2970 997 -2956
rect 1010 -2970 1011 -2956
rect 1143 -3075 1144 -2969
rect 1199 -3075 1200 -2969
rect 1241 -2970 1242 -2956
rect 1339 -2970 1340 -2956
rect 1584 -3075 1585 -2969
rect 1647 -3075 1648 -2969
rect 1682 -2970 1683 -2956
rect 65 -2972 66 -2956
rect 219 -3075 220 -2971
rect 261 -2972 262 -2956
rect 394 -3075 395 -2971
rect 408 -2972 409 -2956
rect 457 -3075 458 -2971
rect 492 -2972 493 -2956
rect 569 -3075 570 -2971
rect 604 -2972 605 -2956
rect 618 -3075 619 -2971
rect 674 -3075 675 -2971
rect 793 -2972 794 -2956
rect 835 -2972 836 -2956
rect 1150 -3075 1151 -2971
rect 1164 -2972 1165 -2956
rect 1241 -3075 1242 -2971
rect 1339 -3075 1340 -2971
rect 1388 -2972 1389 -2956
rect 1465 -3075 1466 -2971
rect 1486 -2972 1487 -2956
rect 65 -3075 66 -2973
rect 208 -3075 209 -2973
rect 261 -3075 262 -2973
rect 513 -2974 514 -2956
rect 604 -3075 605 -2973
rect 758 -2974 759 -2956
rect 782 -2974 783 -2956
rect 1535 -2974 1536 -2956
rect 82 -2976 83 -2956
rect 1178 -2976 1179 -2956
rect 1213 -3075 1214 -2975
rect 1255 -2976 1256 -2956
rect 1297 -2976 1298 -2956
rect 1388 -3075 1389 -2975
rect 1486 -3075 1487 -2975
rect 1493 -2976 1494 -2956
rect 1535 -3075 1536 -2975
rect 1563 -2976 1564 -2956
rect 93 -3075 94 -2977
rect 562 -2978 563 -2956
rect 793 -3075 794 -2977
rect 926 -2978 927 -2956
rect 943 -2978 944 -2956
rect 1416 -2978 1417 -2956
rect 1430 -2978 1431 -2956
rect 1563 -3075 1564 -2977
rect 79 -3075 80 -2979
rect 1416 -3075 1417 -2979
rect 1430 -3075 1431 -2979
rect 1668 -2980 1669 -2956
rect 100 -3075 101 -2981
rect 660 -2982 661 -2956
rect 835 -3075 836 -2981
rect 989 -2982 990 -2956
rect 996 -3075 997 -2981
rect 1038 -2982 1039 -2956
rect 1052 -3075 1053 -2981
rect 1059 -2982 1060 -2956
rect 1094 -3075 1095 -2981
rect 1318 -2982 1319 -2956
rect 1493 -3075 1494 -2981
rect 1514 -2982 1515 -2956
rect 107 -2984 108 -2956
rect 1024 -3075 1025 -2983
rect 1031 -2984 1032 -2956
rect 1591 -2984 1592 -2956
rect 107 -3075 108 -2985
rect 443 -2986 444 -2956
rect 562 -3075 563 -2985
rect 866 -2986 867 -2956
rect 891 -2986 892 -2956
rect 891 -3075 892 -2985
rect 891 -2986 892 -2956
rect 891 -3075 892 -2985
rect 901 -3075 902 -2985
rect 1423 -2986 1424 -2956
rect 1514 -3075 1515 -2985
rect 1549 -2986 1550 -2956
rect 1591 -3075 1592 -2985
rect 1633 -2986 1634 -2956
rect 110 -2988 111 -2956
rect 254 -2988 255 -2956
rect 268 -2988 269 -2956
rect 1097 -2988 1098 -2956
rect 1115 -3075 1116 -2987
rect 1129 -2988 1130 -2956
rect 1136 -2988 1137 -2956
rect 1178 -3075 1179 -2987
rect 1202 -2988 1203 -2956
rect 1633 -3075 1634 -2987
rect 121 -2990 122 -2956
rect 621 -3075 622 -2989
rect 660 -3075 661 -2989
rect 730 -2990 731 -2956
rect 849 -3075 850 -2989
rect 884 -2990 885 -2956
rect 905 -2990 906 -2956
rect 905 -3075 906 -2989
rect 905 -2990 906 -2956
rect 905 -3075 906 -2989
rect 926 -3075 927 -2989
rect 947 -2990 948 -2956
rect 982 -2990 983 -2956
rect 1038 -3075 1039 -2989
rect 1045 -2990 1046 -2956
rect 1129 -3075 1130 -2989
rect 1136 -3075 1137 -2989
rect 1360 -2990 1361 -2956
rect 1423 -3075 1424 -2989
rect 1675 -2990 1676 -2956
rect 82 -3075 83 -2991
rect 1045 -3075 1046 -2991
rect 1055 -2992 1056 -2956
rect 1521 -2992 1522 -2956
rect 1549 -3075 1550 -2991
rect 1570 -2992 1571 -2956
rect 121 -3075 122 -2993
rect 359 -2994 360 -2956
rect 408 -3075 409 -2993
rect 415 -2994 416 -2956
rect 443 -3075 444 -2993
rect 667 -2994 668 -2956
rect 852 -2994 853 -2956
rect 919 -2994 920 -2956
rect 947 -3075 948 -2993
rect 954 -2994 955 -2956
rect 989 -3075 990 -2993
rect 1073 -2994 1074 -2956
rect 1122 -2994 1123 -2956
rect 1164 -3075 1165 -2993
rect 1220 -3075 1221 -2993
rect 1262 -2994 1263 -2956
rect 1297 -3075 1298 -2993
rect 1353 -2994 1354 -2956
rect 1521 -3075 1522 -2993
rect 1556 -2994 1557 -2956
rect 1570 -3075 1571 -2993
rect 1598 -2994 1599 -2956
rect 89 -3075 90 -2995
rect 1122 -3075 1123 -2995
rect 1255 -3075 1256 -2995
rect 1290 -2996 1291 -2956
rect 1318 -3075 1319 -2995
rect 1367 -2996 1368 -2956
rect 1598 -3075 1599 -2995
rect 1626 -2996 1627 -2956
rect 142 -2998 143 -2956
rect 982 -3075 983 -2997
rect 1010 -3075 1011 -2997
rect 1227 -2998 1228 -2956
rect 1262 -3075 1263 -2997
rect 1311 -2998 1312 -2956
rect 1367 -3075 1368 -2997
rect 1395 -2998 1396 -2956
rect 1626 -3075 1627 -2997
rect 1661 -2998 1662 -2956
rect 145 -3075 146 -2999
rect 583 -3000 584 -2956
rect 632 -3000 633 -2956
rect 730 -3075 731 -2999
rect 856 -3075 857 -2999
rect 870 -3000 871 -2956
rect 877 -3000 878 -2956
rect 919 -3075 920 -2999
rect 954 -3075 955 -2999
rect 961 -3000 962 -2956
rect 968 -3000 969 -2956
rect 1073 -3075 1074 -2999
rect 1227 -3075 1228 -2999
rect 1346 -3000 1347 -2956
rect 156 -3002 157 -2956
rect 254 -3075 255 -3001
rect 268 -3075 269 -3001
rect 380 -3002 381 -2956
rect 415 -3075 416 -3001
rect 422 -3002 423 -2956
rect 506 -3002 507 -2956
rect 1360 -3075 1361 -3001
rect 156 -3075 157 -3003
rect 786 -3004 787 -2956
rect 880 -3075 881 -3003
rect 1353 -3075 1354 -3003
rect 163 -3006 164 -2956
rect 933 -3006 934 -2956
rect 961 -3075 962 -3005
rect 1335 -3006 1336 -2956
rect 1346 -3075 1347 -3005
rect 1706 -3006 1707 -2956
rect 86 -3008 87 -2956
rect 163 -3075 164 -3007
rect 170 -3008 171 -2956
rect 226 -3008 227 -2956
rect 282 -3008 283 -2956
rect 380 -3075 381 -3007
rect 401 -3008 402 -2956
rect 506 -3075 507 -3007
rect 583 -3075 584 -3007
rect 940 -3008 941 -2956
rect 968 -3075 969 -3007
rect 975 -3008 976 -2956
rect 1017 -3008 1018 -2956
rect 1031 -3075 1032 -3007
rect 1034 -3008 1035 -2956
rect 1612 -3008 1613 -2956
rect 86 -3075 87 -3009
rect 1619 -3010 1620 -2956
rect 128 -3012 129 -2956
rect 226 -3075 227 -3011
rect 275 -3012 276 -2956
rect 282 -3075 283 -3011
rect 289 -3075 290 -3011
rect 576 -3012 577 -2956
rect 632 -3075 633 -3011
rect 863 -3075 864 -3011
rect 884 -3075 885 -3011
rect 1108 -3012 1109 -2956
rect 1234 -3012 1235 -2956
rect 1311 -3075 1312 -3011
rect 1612 -3075 1613 -3011
rect 1654 -3012 1655 -2956
rect 58 -3014 59 -2956
rect 576 -3075 577 -3013
rect 639 -3014 640 -2956
rect 667 -3075 668 -3013
rect 702 -3014 703 -2956
rect 877 -3075 878 -3013
rect 898 -3014 899 -2956
rect 933 -3075 934 -3013
rect 1059 -3075 1060 -3013
rect 1087 -3014 1088 -2956
rect 1108 -3075 1109 -3013
rect 1206 -3014 1207 -2956
rect 1234 -3075 1235 -3013
rect 1276 -3014 1277 -2956
rect 58 -3075 59 -3015
rect 135 -3016 136 -2956
rect 138 -3016 139 -2956
rect 275 -3075 276 -3015
rect 303 -3075 304 -3015
rect 478 -3016 479 -2956
rect 513 -3075 514 -3015
rect 1017 -3075 1018 -3015
rect 1192 -3016 1193 -2956
rect 1654 -3075 1655 -3015
rect 128 -3075 129 -3017
rect 695 -3018 696 -2956
rect 702 -3075 703 -3017
rect 723 -3018 724 -2956
rect 789 -3075 790 -3017
rect 940 -3075 941 -3017
rect 1185 -3018 1186 -2956
rect 1192 -3075 1193 -3017
rect 1206 -3075 1207 -3017
rect 1248 -3018 1249 -2956
rect 170 -3075 171 -3019
rect 191 -3020 192 -2956
rect 205 -3020 206 -2956
rect 296 -3020 297 -2956
rect 317 -3020 318 -2956
rect 422 -3075 423 -3019
rect 478 -3075 479 -3019
rect 555 -3020 556 -2956
rect 639 -3075 640 -3019
rect 646 -3020 647 -2956
rect 656 -3020 657 -2956
rect 1290 -3075 1291 -3019
rect 61 -3075 62 -3021
rect 296 -3075 297 -3021
rect 555 -3075 556 -3021
rect 646 -3075 647 -3021
rect 1101 -3022 1102 -2956
rect 1248 -3075 1249 -3021
rect 1283 -3022 1284 -2956
rect 177 -3024 178 -2956
rect 691 -3075 692 -3023
rect 709 -3024 710 -2956
rect 870 -3075 871 -3023
rect 898 -3075 899 -3023
rect 1066 -3024 1067 -2956
rect 1283 -3075 1284 -3023
rect 1325 -3024 1326 -2956
rect 177 -3075 178 -3025
rect 373 -3026 374 -2956
rect 401 -3075 402 -3025
rect 429 -3026 430 -2956
rect 681 -3026 682 -2956
rect 1276 -3075 1277 -3025
rect 1325 -3075 1326 -3025
rect 1374 -3026 1375 -2956
rect 114 -3028 115 -2956
rect 429 -3075 430 -3027
rect 464 -3028 465 -2956
rect 681 -3075 682 -3027
rect 688 -3075 689 -3027
rect 1101 -3075 1102 -3027
rect 1374 -3075 1375 -3027
rect 1402 -3028 1403 -2956
rect 149 -3030 150 -2956
rect 464 -3075 465 -3029
rect 709 -3075 710 -3029
rect 751 -3030 752 -2956
rect 912 -3030 913 -2956
rect 1556 -3075 1557 -3029
rect 149 -3075 150 -3031
rect 1157 -3032 1158 -2956
rect 1304 -3032 1305 -2956
rect 1402 -3075 1403 -3031
rect 187 -3075 188 -3033
rect 1528 -3075 1529 -3033
rect 191 -3075 192 -3035
rect 198 -3036 199 -2956
rect 205 -3075 206 -3035
rect 387 -3036 388 -2956
rect 716 -3036 717 -2956
rect 1157 -3075 1158 -3035
rect 1269 -3036 1270 -2956
rect 1304 -3075 1305 -3035
rect 310 -3038 311 -2956
rect 317 -3075 318 -3037
rect 338 -3038 339 -2956
rect 373 -3075 374 -3037
rect 387 -3075 388 -3037
rect 527 -3038 528 -2956
rect 716 -3075 717 -3037
rect 744 -3038 745 -2956
rect 751 -3075 752 -3037
rect 772 -3038 773 -2956
rect 1003 -3038 1004 -2956
rect 1185 -3075 1186 -3037
rect 1269 -3075 1270 -3037
rect 1437 -3038 1438 -2956
rect 184 -3040 185 -2956
rect 744 -3075 745 -3039
rect 1066 -3075 1067 -3039
rect 1080 -3040 1081 -2956
rect 184 -3075 185 -3041
rect 800 -3042 801 -2956
rect 1080 -3075 1081 -3041
rect 1409 -3042 1410 -2956
rect 310 -3075 311 -3043
rect 625 -3044 626 -2956
rect 723 -3075 724 -3043
rect 758 -3075 759 -3043
rect 800 -3075 801 -3043
rect 1619 -3075 1620 -3043
rect 324 -3046 325 -2956
rect 338 -3075 339 -3045
rect 345 -3046 346 -2956
rect 625 -3075 626 -3045
rect 1409 -3075 1410 -3045
rect 1451 -3046 1452 -2956
rect 324 -3075 325 -3047
rect 331 -3048 332 -2956
rect 345 -3075 346 -3047
rect 695 -3075 696 -3047
rect 786 -3075 787 -3047
rect 1451 -3075 1452 -3047
rect 331 -3075 332 -3049
rect 366 -3050 367 -2956
rect 485 -3050 486 -2956
rect 1437 -3075 1438 -3049
rect 114 -3075 115 -3051
rect 366 -3075 367 -3051
rect 485 -3075 486 -3051
rect 590 -3052 591 -2956
rect 352 -3054 353 -2956
rect 492 -3075 493 -3053
rect 520 -3054 521 -2956
rect 772 -3075 773 -3053
rect 152 -3075 153 -3055
rect 352 -3075 353 -3055
rect 359 -3075 360 -3055
rect 537 -3056 538 -2956
rect 590 -3075 591 -3055
rect 915 -3056 916 -2956
rect 471 -3058 472 -2956
rect 520 -3075 521 -3057
rect 527 -3075 528 -3057
rect 765 -3058 766 -2956
rect 915 -3075 916 -3057
rect 1479 -3058 1480 -2956
rect 471 -3075 472 -3059
rect 737 -3060 738 -2956
rect 765 -3075 766 -3059
rect 807 -3060 808 -2956
rect 1479 -3075 1480 -3059
rect 1500 -3060 1501 -2956
rect 534 -3062 535 -2956
rect 1003 -3075 1004 -3061
rect 1500 -3075 1501 -3061
rect 1542 -3062 1543 -2956
rect 233 -3064 234 -2956
rect 534 -3075 535 -3063
rect 737 -3075 738 -3063
rect 1395 -3075 1396 -3063
rect 1444 -3064 1445 -2956
rect 1542 -3075 1543 -3063
rect 233 -3075 234 -3065
rect 240 -3066 241 -2956
rect 807 -3075 808 -3065
rect 828 -3066 829 -2956
rect 1444 -3075 1445 -3065
rect 1472 -3066 1473 -2956
rect 240 -3075 241 -3067
rect 247 -3068 248 -2956
rect 828 -3075 829 -3067
rect 1507 -3075 1508 -3067
rect 247 -3075 248 -3069
rect 779 -3070 780 -2956
rect 831 -3075 832 -3069
rect 1472 -3075 1473 -3069
rect 597 -3072 598 -2956
rect 779 -3075 780 -3071
rect 597 -3075 598 -3073
rect 635 -3075 636 -3073
rect 30 -3085 31 -3083
rect 474 -3214 475 -3084
rect 478 -3085 479 -3083
rect 635 -3085 636 -3083
rect 646 -3085 647 -3083
rect 975 -3085 976 -3083
rect 999 -3214 1000 -3084
rect 1633 -3085 1634 -3083
rect 37 -3087 38 -3083
rect 86 -3087 87 -3083
rect 114 -3087 115 -3083
rect 212 -3214 213 -3086
rect 215 -3087 216 -3083
rect 254 -3087 255 -3083
rect 275 -3087 276 -3083
rect 800 -3087 801 -3083
rect 814 -3087 815 -3083
rect 1087 -3087 1088 -3083
rect 1090 -3087 1091 -3083
rect 1388 -3087 1389 -3083
rect 1475 -3214 1476 -3086
rect 1570 -3087 1571 -3083
rect 61 -3089 62 -3083
rect 625 -3089 626 -3083
rect 656 -3214 657 -3088
rect 779 -3089 780 -3083
rect 789 -3089 790 -3083
rect 842 -3089 843 -3083
rect 877 -3089 878 -3083
rect 1171 -3089 1172 -3083
rect 1388 -3214 1389 -3088
rect 1563 -3089 1564 -3083
rect 65 -3091 66 -3083
rect 79 -3091 80 -3083
rect 82 -3091 83 -3083
rect 436 -3091 437 -3083
rect 471 -3091 472 -3083
rect 803 -3091 804 -3083
rect 842 -3214 843 -3090
rect 982 -3091 983 -3083
rect 1020 -3091 1021 -3083
rect 1458 -3091 1459 -3083
rect 79 -3214 80 -3092
rect 695 -3093 696 -3083
rect 716 -3093 717 -3083
rect 915 -3093 916 -3083
rect 933 -3093 934 -3083
rect 1090 -3214 1091 -3092
rect 1171 -3214 1172 -3092
rect 1339 -3093 1340 -3083
rect 1444 -3093 1445 -3083
rect 1458 -3214 1459 -3092
rect 86 -3214 87 -3094
rect 177 -3095 178 -3083
rect 184 -3095 185 -3083
rect 950 -3095 951 -3083
rect 975 -3214 976 -3094
rect 1031 -3095 1032 -3083
rect 1062 -3214 1063 -3094
rect 1584 -3095 1585 -3083
rect 117 -3214 118 -3096
rect 1276 -3097 1277 -3083
rect 1339 -3214 1340 -3096
rect 1528 -3097 1529 -3083
rect 131 -3214 132 -3098
rect 205 -3214 206 -3098
rect 219 -3099 220 -3083
rect 222 -3149 223 -3098
rect 254 -3214 255 -3098
rect 926 -3099 927 -3083
rect 933 -3214 934 -3098
rect 1199 -3099 1200 -3083
rect 1276 -3214 1277 -3098
rect 1430 -3099 1431 -3083
rect 135 -3101 136 -3083
rect 163 -3101 164 -3083
rect 177 -3214 178 -3100
rect 240 -3101 241 -3083
rect 282 -3101 283 -3083
rect 394 -3101 395 -3083
rect 404 -3214 405 -3100
rect 436 -3214 437 -3100
rect 453 -3101 454 -3083
rect 926 -3214 927 -3100
rect 940 -3101 941 -3083
rect 1199 -3214 1200 -3100
rect 1423 -3101 1424 -3083
rect 1444 -3214 1445 -3100
rect 51 -3103 52 -3083
rect 282 -3214 283 -3102
rect 303 -3103 304 -3083
rect 502 -3214 503 -3102
rect 527 -3103 528 -3083
rect 625 -3214 626 -3102
rect 674 -3103 675 -3083
rect 761 -3103 762 -3083
rect 779 -3214 780 -3102
rect 1038 -3103 1039 -3083
rect 1083 -3103 1084 -3083
rect 1367 -3103 1368 -3083
rect 1423 -3214 1424 -3102
rect 1605 -3103 1606 -3083
rect 93 -3105 94 -3083
rect 303 -3214 304 -3104
rect 317 -3105 318 -3083
rect 317 -3214 318 -3104
rect 317 -3105 318 -3083
rect 317 -3214 318 -3104
rect 324 -3105 325 -3083
rect 324 -3214 325 -3104
rect 324 -3105 325 -3083
rect 324 -3214 325 -3104
rect 345 -3214 346 -3104
rect 352 -3105 353 -3083
rect 366 -3105 367 -3083
rect 583 -3105 584 -3083
rect 593 -3214 594 -3104
rect 660 -3105 661 -3083
rect 674 -3214 675 -3104
rect 744 -3105 745 -3083
rect 758 -3214 759 -3104
rect 919 -3105 920 -3083
rect 940 -3214 941 -3104
rect 1059 -3105 1060 -3083
rect 1367 -3214 1368 -3104
rect 1542 -3105 1543 -3083
rect 1605 -3214 1606 -3104
rect 1647 -3105 1648 -3083
rect 93 -3214 94 -3106
rect 737 -3107 738 -3083
rect 744 -3214 745 -3106
rect 891 -3107 892 -3083
rect 919 -3214 920 -3106
rect 1052 -3107 1053 -3083
rect 1430 -3214 1431 -3106
rect 1612 -3107 1613 -3083
rect 135 -3214 136 -3108
rect 681 -3109 682 -3083
rect 684 -3214 685 -3108
rect 1360 -3109 1361 -3083
rect 142 -3111 143 -3083
rect 1486 -3111 1487 -3083
rect 142 -3214 143 -3112
rect 772 -3113 773 -3083
rect 793 -3113 794 -3083
rect 796 -3214 797 -3112
rect 800 -3214 801 -3112
rect 838 -3113 839 -3083
rect 877 -3214 878 -3112
rect 1024 -3113 1025 -3083
rect 1031 -3214 1032 -3112
rect 1087 -3214 1088 -3112
rect 1360 -3214 1361 -3112
rect 1535 -3113 1536 -3083
rect 145 -3115 146 -3083
rect 170 -3115 171 -3083
rect 184 -3214 185 -3114
rect 513 -3115 514 -3083
rect 534 -3115 535 -3083
rect 828 -3115 829 -3083
rect 838 -3214 839 -3114
rect 1066 -3115 1067 -3083
rect 1486 -3214 1487 -3114
rect 1626 -3115 1627 -3083
rect 121 -3117 122 -3083
rect 534 -3214 535 -3116
rect 562 -3117 563 -3083
rect 646 -3214 647 -3116
rect 660 -3214 661 -3116
rect 782 -3214 783 -3116
rect 793 -3214 794 -3116
rect 1640 -3117 1641 -3083
rect 100 -3119 101 -3083
rect 121 -3214 122 -3118
rect 149 -3119 150 -3083
rect 1395 -3119 1396 -3083
rect 89 -3121 90 -3083
rect 100 -3214 101 -3120
rect 152 -3121 153 -3083
rect 268 -3121 269 -3083
rect 348 -3121 349 -3083
rect 380 -3121 381 -3083
rect 394 -3214 395 -3120
rect 506 -3121 507 -3083
rect 562 -3214 563 -3120
rect 821 -3121 822 -3083
rect 828 -3214 829 -3120
rect 968 -3121 969 -3083
rect 982 -3214 983 -3120
rect 1129 -3121 1130 -3083
rect 44 -3123 45 -3083
rect 268 -3214 269 -3122
rect 352 -3214 353 -3122
rect 590 -3123 591 -3083
rect 618 -3214 619 -3122
rect 702 -3123 703 -3083
rect 716 -3214 717 -3122
rect 835 -3123 836 -3083
rect 947 -3123 948 -3083
rect 1164 -3123 1165 -3083
rect 152 -3214 153 -3124
rect 786 -3125 787 -3083
rect 821 -3214 822 -3124
rect 1101 -3125 1102 -3083
rect 1129 -3214 1130 -3124
rect 1283 -3125 1284 -3083
rect 156 -3127 157 -3083
rect 506 -3214 507 -3126
rect 576 -3127 577 -3083
rect 1059 -3214 1060 -3126
rect 1066 -3214 1067 -3126
rect 1234 -3127 1235 -3083
rect 1283 -3214 1284 -3126
rect 1465 -3127 1466 -3083
rect 156 -3214 157 -3128
rect 653 -3129 654 -3083
rect 688 -3129 689 -3083
rect 723 -3129 724 -3083
rect 730 -3129 731 -3083
rect 814 -3214 815 -3128
rect 835 -3214 836 -3128
rect 1353 -3129 1354 -3083
rect 163 -3214 164 -3130
rect 740 -3131 741 -3083
rect 772 -3214 773 -3130
rect 1073 -3131 1074 -3083
rect 1164 -3214 1165 -3130
rect 1269 -3131 1270 -3083
rect 170 -3214 171 -3132
rect 401 -3133 402 -3083
rect 429 -3133 430 -3083
rect 583 -3214 584 -3132
rect 653 -3214 654 -3132
rect 688 -3214 689 -3132
rect 691 -3133 692 -3083
rect 1598 -3133 1599 -3083
rect 191 -3135 192 -3083
rect 201 -3135 202 -3083
rect 219 -3214 220 -3134
rect 443 -3135 444 -3083
rect 457 -3135 458 -3083
rect 513 -3214 514 -3134
rect 579 -3214 580 -3134
rect 1101 -3214 1102 -3134
rect 1234 -3214 1235 -3134
rect 1409 -3135 1410 -3083
rect 128 -3137 129 -3083
rect 457 -3214 458 -3136
rect 478 -3214 479 -3136
rect 751 -3137 752 -3083
rect 786 -3214 787 -3136
rect 898 -3137 899 -3083
rect 947 -3214 948 -3136
rect 1402 -3137 1403 -3083
rect 1409 -3214 1410 -3136
rect 1514 -3137 1515 -3083
rect 72 -3139 73 -3083
rect 128 -3214 129 -3138
rect 191 -3214 192 -3138
rect 247 -3139 248 -3083
rect 261 -3139 262 -3083
rect 443 -3214 444 -3138
rect 492 -3139 493 -3083
rect 527 -3214 528 -3138
rect 681 -3214 682 -3138
rect 723 -3214 724 -3138
rect 730 -3214 731 -3138
rect 849 -3139 850 -3083
rect 898 -3214 899 -3138
rect 989 -3139 990 -3083
rect 1003 -3139 1004 -3083
rect 1073 -3214 1074 -3138
rect 1269 -3214 1270 -3138
rect 1521 -3139 1522 -3083
rect 72 -3214 73 -3140
rect 226 -3141 227 -3083
rect 233 -3141 234 -3083
rect 247 -3214 248 -3140
rect 261 -3214 262 -3140
rect 289 -3141 290 -3083
rect 366 -3214 367 -3140
rect 415 -3141 416 -3083
rect 432 -3214 433 -3140
rect 464 -3141 465 -3083
rect 492 -3214 493 -3140
rect 548 -3141 549 -3083
rect 695 -3214 696 -3140
rect 824 -3214 825 -3140
rect 849 -3214 850 -3140
rect 954 -3141 955 -3083
rect 968 -3214 969 -3140
rect 1227 -3141 1228 -3083
rect 1297 -3141 1298 -3083
rect 1514 -3214 1515 -3140
rect 198 -3143 199 -3083
rect 1080 -3143 1081 -3083
rect 1178 -3143 1179 -3083
rect 1297 -3214 1298 -3142
rect 1325 -3143 1326 -3083
rect 1521 -3214 1522 -3142
rect 149 -3214 150 -3144
rect 1080 -3214 1081 -3144
rect 1178 -3214 1179 -3144
rect 1311 -3145 1312 -3083
rect 1325 -3214 1326 -3144
rect 1500 -3145 1501 -3083
rect 198 -3214 199 -3146
rect 870 -3147 871 -3083
rect 954 -3214 955 -3146
rect 1150 -3147 1151 -3083
rect 1227 -3214 1228 -3146
rect 1416 -3147 1417 -3083
rect 289 -3214 290 -3148
rect 369 -3149 370 -3083
rect 408 -3149 409 -3083
rect 537 -3214 538 -3148
rect 1416 -3214 1417 -3148
rect 226 -3214 227 -3150
rect 604 -3151 605 -3083
rect 702 -3214 703 -3150
rect 856 -3151 857 -3083
rect 870 -3214 871 -3150
rect 1412 -3214 1413 -3150
rect 233 -3214 234 -3152
rect 611 -3153 612 -3083
rect 737 -3214 738 -3152
rect 765 -3153 766 -3083
rect 856 -3214 857 -3152
rect 884 -3153 885 -3083
rect 989 -3214 990 -3152
rect 1437 -3153 1438 -3083
rect 373 -3155 374 -3083
rect 415 -3214 416 -3154
rect 548 -3214 549 -3154
rect 667 -3155 668 -3083
rect 751 -3214 752 -3154
rect 905 -3155 906 -3083
rect 1003 -3214 1004 -3154
rect 1157 -3155 1158 -3083
rect 1311 -3214 1312 -3154
rect 1479 -3155 1480 -3083
rect 107 -3157 108 -3083
rect 373 -3214 374 -3156
rect 380 -3214 381 -3156
rect 541 -3157 542 -3083
rect 597 -3157 598 -3083
rect 604 -3214 605 -3156
rect 611 -3214 612 -3156
rect 709 -3157 710 -3083
rect 765 -3214 766 -3156
rect 1013 -3214 1014 -3156
rect 1024 -3214 1025 -3156
rect 1115 -3157 1116 -3083
rect 1122 -3157 1123 -3083
rect 1500 -3214 1501 -3156
rect 107 -3214 108 -3158
rect 639 -3159 640 -3083
rect 667 -3214 668 -3158
rect 863 -3159 864 -3083
rect 884 -3214 885 -3158
rect 1010 -3159 1011 -3083
rect 1038 -3214 1039 -3158
rect 1248 -3159 1249 -3083
rect 1402 -3214 1403 -3158
rect 1591 -3159 1592 -3083
rect 387 -3161 388 -3083
rect 464 -3214 465 -3160
rect 471 -3214 472 -3160
rect 863 -3214 864 -3160
rect 905 -3214 906 -3160
rect 912 -3161 913 -3083
rect 1052 -3214 1053 -3160
rect 1220 -3161 1221 -3083
rect 1248 -3214 1249 -3160
rect 1507 -3161 1508 -3083
rect 387 -3214 388 -3162
rect 1143 -3163 1144 -3083
rect 1150 -3214 1151 -3162
rect 1213 -3163 1214 -3083
rect 1220 -3214 1221 -3162
rect 1381 -3163 1382 -3083
rect 1437 -3214 1438 -3162
rect 1619 -3163 1620 -3083
rect 401 -3214 402 -3164
rect 520 -3165 521 -3083
rect 590 -3214 591 -3164
rect 597 -3214 598 -3164
rect 632 -3165 633 -3083
rect 1213 -3214 1214 -3164
rect 1304 -3165 1305 -3083
rect 1507 -3214 1508 -3164
rect 114 -3214 115 -3166
rect 520 -3214 521 -3166
rect 632 -3214 633 -3166
rect 961 -3167 962 -3083
rect 978 -3167 979 -3083
rect 1304 -3214 1305 -3166
rect 1381 -3214 1382 -3166
rect 1556 -3167 1557 -3083
rect 408 -3214 409 -3168
rect 569 -3169 570 -3083
rect 639 -3214 640 -3168
rect 1206 -3169 1207 -3083
rect 429 -3214 430 -3170
rect 569 -3214 570 -3170
rect 709 -3214 710 -3170
rect 807 -3171 808 -3083
rect 912 -3214 913 -3170
rect 1045 -3171 1046 -3083
rect 1094 -3171 1095 -3083
rect 1115 -3214 1116 -3170
rect 1122 -3214 1123 -3170
rect 1318 -3171 1319 -3083
rect 576 -3214 577 -3172
rect 807 -3214 808 -3172
rect 961 -3214 962 -3172
rect 1108 -3173 1109 -3083
rect 1136 -3173 1137 -3083
rect 1157 -3214 1158 -3172
rect 1185 -3173 1186 -3083
rect 1479 -3214 1480 -3172
rect 1045 -3214 1046 -3174
rect 1192 -3175 1193 -3083
rect 1206 -3214 1207 -3174
rect 1374 -3175 1375 -3083
rect 1094 -3214 1095 -3176
rect 1262 -3177 1263 -3083
rect 1318 -3214 1319 -3176
rect 1493 -3177 1494 -3083
rect 996 -3179 997 -3083
rect 1493 -3214 1494 -3178
rect 996 -3214 997 -3180
rect 1395 -3214 1396 -3180
rect 1017 -3183 1018 -3083
rect 1262 -3214 1263 -3182
rect 1374 -3214 1375 -3182
rect 1549 -3183 1550 -3083
rect 1017 -3214 1018 -3184
rect 1290 -3185 1291 -3083
rect 1108 -3214 1109 -3186
rect 1654 -3187 1655 -3083
rect 1136 -3214 1137 -3188
rect 1255 -3189 1256 -3083
rect 1290 -3214 1291 -3188
rect 1472 -3189 1473 -3083
rect 1143 -3214 1144 -3190
rect 1241 -3191 1242 -3083
rect 1255 -3214 1256 -3190
rect 1451 -3191 1452 -3083
rect 450 -3193 451 -3083
rect 1451 -3214 1452 -3192
rect 310 -3195 311 -3083
rect 450 -3214 451 -3194
rect 1185 -3214 1186 -3194
rect 1332 -3195 1333 -3083
rect 310 -3214 311 -3196
rect 331 -3197 332 -3083
rect 621 -3197 622 -3083
rect 1332 -3214 1333 -3196
rect 331 -3214 332 -3198
rect 422 -3199 423 -3083
rect 1192 -3214 1193 -3198
rect 1346 -3199 1347 -3083
rect 422 -3214 423 -3200
rect 485 -3201 486 -3083
rect 1241 -3214 1242 -3200
rect 1577 -3201 1578 -3083
rect 296 -3203 297 -3083
rect 485 -3214 486 -3202
rect 1346 -3214 1347 -3202
rect 1465 -3214 1466 -3202
rect 296 -3214 297 -3204
rect 338 -3205 339 -3083
rect 338 -3214 339 -3206
rect 359 -3207 360 -3083
rect 359 -3214 360 -3208
rect 555 -3209 556 -3083
rect 499 -3211 500 -3083
rect 555 -3214 556 -3210
rect 275 -3214 276 -3212
rect 499 -3214 500 -3212
rect 65 -3224 66 -3222
rect 114 -3224 115 -3222
rect 121 -3224 122 -3222
rect 499 -3224 500 -3222
rect 502 -3224 503 -3222
rect 716 -3224 717 -3222
rect 779 -3224 780 -3222
rect 870 -3224 871 -3222
rect 880 -3307 881 -3223
rect 1031 -3224 1032 -3222
rect 1059 -3307 1060 -3223
rect 1332 -3224 1333 -3222
rect 1346 -3224 1347 -3222
rect 1479 -3224 1480 -3222
rect 1584 -3307 1585 -3223
rect 1605 -3224 1606 -3222
rect 72 -3226 73 -3222
rect 471 -3226 472 -3222
rect 485 -3226 486 -3222
rect 579 -3226 580 -3222
rect 593 -3226 594 -3222
rect 674 -3226 675 -3222
rect 684 -3226 685 -3222
rect 786 -3226 787 -3222
rect 800 -3226 801 -3222
rect 1356 -3226 1357 -3222
rect 1409 -3226 1410 -3222
rect 1521 -3226 1522 -3222
rect 86 -3228 87 -3222
rect 401 -3228 402 -3222
rect 404 -3228 405 -3222
rect 527 -3228 528 -3222
rect 544 -3228 545 -3222
rect 555 -3228 556 -3222
rect 576 -3228 577 -3222
rect 611 -3228 612 -3222
rect 625 -3228 626 -3222
rect 796 -3228 797 -3222
rect 800 -3307 801 -3227
rect 849 -3228 850 -3222
rect 894 -3228 895 -3222
rect 1157 -3228 1158 -3222
rect 1185 -3228 1186 -3222
rect 1209 -3307 1210 -3227
rect 1297 -3307 1298 -3227
rect 1493 -3228 1494 -3222
rect 142 -3230 143 -3222
rect 576 -3307 577 -3229
rect 597 -3230 598 -3222
rect 597 -3307 598 -3229
rect 597 -3230 598 -3222
rect 597 -3307 598 -3229
rect 611 -3307 612 -3229
rect 737 -3230 738 -3222
rect 849 -3307 850 -3229
rect 954 -3230 955 -3222
rect 999 -3230 1000 -3222
rect 1003 -3230 1004 -3222
rect 1010 -3230 1011 -3222
rect 1269 -3230 1270 -3222
rect 1300 -3230 1301 -3222
rect 1465 -3230 1466 -3222
rect 149 -3232 150 -3222
rect 191 -3232 192 -3222
rect 212 -3232 213 -3222
rect 240 -3307 241 -3231
rect 243 -3232 244 -3222
rect 317 -3232 318 -3222
rect 324 -3232 325 -3222
rect 1013 -3232 1014 -3222
rect 1020 -3307 1021 -3231
rect 1136 -3232 1137 -3222
rect 1269 -3307 1270 -3231
rect 1381 -3232 1382 -3222
rect 1458 -3232 1459 -3222
rect 1531 -3307 1532 -3231
rect 107 -3234 108 -3222
rect 212 -3307 213 -3233
rect 226 -3234 227 -3222
rect 485 -3307 486 -3233
rect 492 -3234 493 -3222
rect 772 -3234 773 -3222
rect 905 -3234 906 -3222
rect 985 -3307 986 -3233
rect 1010 -3307 1011 -3233
rect 1206 -3234 1207 -3222
rect 1325 -3234 1326 -3222
rect 1328 -3234 1329 -3222
rect 1332 -3307 1333 -3233
rect 1388 -3234 1389 -3222
rect 152 -3236 153 -3222
rect 359 -3236 360 -3222
rect 387 -3236 388 -3222
rect 390 -3286 391 -3235
rect 415 -3236 416 -3222
rect 541 -3236 542 -3222
rect 544 -3307 545 -3235
rect 835 -3236 836 -3222
rect 905 -3307 906 -3235
rect 1248 -3236 1249 -3222
rect 1325 -3307 1326 -3235
rect 1360 -3236 1361 -3222
rect 1381 -3307 1382 -3235
rect 1507 -3236 1508 -3222
rect 156 -3238 157 -3222
rect 527 -3307 528 -3237
rect 541 -3307 542 -3237
rect 947 -3238 948 -3222
rect 954 -3307 955 -3237
rect 1199 -3238 1200 -3222
rect 1346 -3307 1347 -3237
rect 1423 -3238 1424 -3222
rect 170 -3240 171 -3222
rect 492 -3307 493 -3239
rect 499 -3307 500 -3239
rect 548 -3240 549 -3222
rect 555 -3307 556 -3239
rect 604 -3240 605 -3222
rect 625 -3307 626 -3239
rect 807 -3240 808 -3222
rect 940 -3240 941 -3222
rect 996 -3240 997 -3222
rect 1031 -3307 1032 -3239
rect 1220 -3240 1221 -3222
rect 1349 -3240 1350 -3222
rect 1514 -3240 1515 -3222
rect 93 -3242 94 -3222
rect 170 -3307 171 -3241
rect 177 -3242 178 -3222
rect 348 -3307 349 -3241
rect 359 -3307 360 -3241
rect 394 -3242 395 -3222
rect 429 -3242 430 -3222
rect 450 -3242 451 -3222
rect 457 -3242 458 -3222
rect 590 -3307 591 -3241
rect 604 -3307 605 -3241
rect 667 -3242 668 -3222
rect 705 -3307 706 -3241
rect 1017 -3242 1018 -3222
rect 1087 -3307 1088 -3241
rect 1318 -3242 1319 -3222
rect 1353 -3242 1354 -3222
rect 1486 -3242 1487 -3222
rect 191 -3307 192 -3243
rect 205 -3244 206 -3222
rect 226 -3307 227 -3243
rect 838 -3244 839 -3222
rect 940 -3307 941 -3243
rect 982 -3244 983 -3222
rect 996 -3307 997 -3243
rect 1171 -3244 1172 -3222
rect 1199 -3307 1200 -3243
rect 1241 -3244 1242 -3222
rect 1283 -3244 1284 -3222
rect 1353 -3307 1354 -3243
rect 1388 -3307 1389 -3243
rect 1395 -3244 1396 -3222
rect 205 -3307 206 -3245
rect 632 -3246 633 -3222
rect 653 -3307 654 -3245
rect 702 -3246 703 -3222
rect 709 -3246 710 -3222
rect 824 -3246 825 -3222
rect 919 -3246 920 -3222
rect 1283 -3307 1284 -3245
rect 233 -3248 234 -3222
rect 233 -3307 234 -3247
rect 233 -3248 234 -3222
rect 233 -3307 234 -3247
rect 247 -3248 248 -3222
rect 495 -3248 496 -3222
rect 520 -3248 521 -3222
rect 779 -3307 780 -3247
rect 919 -3307 920 -3247
rect 1080 -3248 1081 -3222
rect 1090 -3248 1091 -3222
rect 1178 -3248 1179 -3222
rect 1220 -3307 1221 -3247
rect 1437 -3248 1438 -3222
rect 135 -3250 136 -3222
rect 247 -3307 248 -3249
rect 254 -3250 255 -3222
rect 677 -3307 678 -3249
rect 709 -3307 710 -3249
rect 901 -3307 902 -3249
rect 947 -3307 948 -3249
rect 1115 -3250 1116 -3222
rect 1129 -3250 1130 -3222
rect 1188 -3307 1189 -3249
rect 1234 -3250 1235 -3222
rect 1241 -3307 1242 -3249
rect 128 -3252 129 -3222
rect 135 -3307 136 -3251
rect 254 -3307 255 -3251
rect 702 -3307 703 -3251
rect 716 -3307 717 -3251
rect 828 -3252 829 -3222
rect 891 -3252 892 -3222
rect 1178 -3307 1179 -3251
rect 1234 -3307 1235 -3251
rect 1304 -3252 1305 -3222
rect 261 -3254 262 -3222
rect 394 -3307 395 -3253
rect 429 -3307 430 -3253
rect 789 -3307 790 -3253
rect 828 -3307 829 -3253
rect 1500 -3254 1501 -3222
rect 261 -3307 262 -3255
rect 331 -3256 332 -3222
rect 338 -3256 339 -3222
rect 439 -3307 440 -3255
rect 450 -3307 451 -3255
rect 478 -3256 479 -3222
rect 520 -3307 521 -3255
rect 569 -3256 570 -3222
rect 632 -3307 633 -3255
rect 730 -3256 731 -3222
rect 737 -3307 738 -3255
rect 1073 -3256 1074 -3222
rect 1080 -3307 1081 -3255
rect 1262 -3256 1263 -3222
rect 1304 -3307 1305 -3255
rect 1475 -3256 1476 -3222
rect 198 -3258 199 -3222
rect 730 -3307 731 -3257
rect 751 -3258 752 -3222
rect 1136 -3307 1137 -3257
rect 1171 -3307 1172 -3257
rect 1276 -3258 1277 -3222
rect 79 -3260 80 -3222
rect 198 -3307 199 -3259
rect 268 -3260 269 -3222
rect 268 -3307 269 -3259
rect 268 -3260 269 -3222
rect 268 -3307 269 -3259
rect 275 -3260 276 -3222
rect 331 -3307 332 -3259
rect 352 -3260 353 -3222
rect 478 -3307 479 -3259
rect 548 -3307 549 -3259
rect 660 -3260 661 -3222
rect 667 -3307 668 -3259
rect 744 -3260 745 -3222
rect 751 -3307 752 -3259
rect 1227 -3260 1228 -3222
rect 1276 -3307 1277 -3259
rect 1374 -3260 1375 -3222
rect 184 -3262 185 -3222
rect 275 -3307 276 -3261
rect 282 -3262 283 -3222
rect 338 -3307 339 -3261
rect 352 -3307 353 -3261
rect 408 -3262 409 -3222
rect 422 -3262 423 -3222
rect 569 -3307 570 -3261
rect 660 -3307 661 -3261
rect 681 -3262 682 -3222
rect 723 -3262 724 -3222
rect 807 -3307 808 -3261
rect 891 -3307 892 -3261
rect 1262 -3307 1263 -3261
rect 163 -3264 164 -3222
rect 408 -3307 409 -3263
rect 422 -3307 423 -3263
rect 618 -3264 619 -3222
rect 681 -3307 682 -3263
rect 695 -3264 696 -3222
rect 723 -3307 724 -3263
rect 842 -3264 843 -3222
rect 968 -3264 969 -3222
rect 1003 -3307 1004 -3263
rect 1052 -3264 1053 -3222
rect 1318 -3307 1319 -3263
rect 100 -3266 101 -3222
rect 163 -3307 164 -3265
rect 184 -3307 185 -3265
rect 534 -3266 535 -3222
rect 618 -3307 619 -3265
rect 989 -3266 990 -3222
rect 1045 -3266 1046 -3222
rect 1052 -3307 1053 -3265
rect 1073 -3307 1074 -3265
rect 1143 -3266 1144 -3222
rect 1213 -3266 1214 -3222
rect 1227 -3307 1228 -3265
rect 282 -3307 283 -3267
rect 950 -3268 951 -3222
rect 968 -3307 969 -3267
rect 1038 -3268 1039 -3222
rect 1045 -3307 1046 -3267
rect 1255 -3268 1256 -3222
rect 296 -3270 297 -3222
rect 324 -3307 325 -3269
rect 373 -3270 374 -3222
rect 415 -3307 416 -3269
rect 457 -3307 458 -3269
rect 793 -3270 794 -3222
rect 814 -3270 815 -3222
rect 1038 -3307 1039 -3269
rect 1094 -3270 1095 -3222
rect 1258 -3307 1259 -3269
rect 296 -3307 297 -3271
rect 380 -3272 381 -3222
rect 387 -3307 388 -3271
rect 443 -3272 444 -3222
rect 471 -3307 472 -3271
rect 530 -3307 531 -3271
rect 534 -3307 535 -3271
rect 982 -3307 983 -3271
rect 1094 -3307 1095 -3271
rect 1290 -3272 1291 -3222
rect 303 -3274 304 -3222
rect 373 -3307 374 -3273
rect 380 -3307 381 -3273
rect 513 -3274 514 -3222
rect 695 -3307 696 -3273
rect 877 -3274 878 -3222
rect 1101 -3274 1102 -3222
rect 1157 -3307 1158 -3273
rect 1290 -3307 1291 -3273
rect 1444 -3274 1445 -3222
rect 303 -3307 304 -3275
rect 310 -3276 311 -3222
rect 317 -3307 318 -3275
rect 345 -3276 346 -3222
rect 443 -3307 444 -3275
rect 744 -3307 745 -3275
rect 821 -3276 822 -3222
rect 842 -3307 843 -3275
rect 1339 -3276 1340 -3222
rect 177 -3307 178 -3277
rect 345 -3307 346 -3277
rect 513 -3307 514 -3277
rect 583 -3278 584 -3222
rect 758 -3278 759 -3222
rect 877 -3307 878 -3277
rect 1101 -3307 1102 -3277
rect 1416 -3278 1417 -3222
rect 289 -3280 290 -3222
rect 310 -3307 311 -3279
rect 464 -3280 465 -3222
rect 583 -3307 584 -3279
rect 758 -3307 759 -3279
rect 884 -3280 885 -3222
rect 1115 -3307 1116 -3279
rect 1430 -3280 1431 -3222
rect 289 -3307 290 -3281
rect 436 -3282 437 -3222
rect 464 -3307 465 -3281
rect 688 -3282 689 -3222
rect 772 -3307 773 -3281
rect 1265 -3307 1266 -3281
rect 1311 -3282 1312 -3222
rect 1339 -3307 1340 -3281
rect 366 -3284 367 -3222
rect 436 -3307 437 -3283
rect 793 -3307 794 -3283
rect 961 -3284 962 -3222
rect 1129 -3307 1130 -3283
rect 1164 -3284 1165 -3222
rect 1311 -3307 1312 -3283
rect 1367 -3284 1368 -3222
rect 219 -3286 220 -3222
rect 366 -3307 367 -3285
rect 814 -3307 815 -3285
rect 1024 -3286 1025 -3222
rect 1143 -3307 1144 -3285
rect 1150 -3286 1151 -3222
rect 1164 -3307 1165 -3285
rect 1192 -3286 1193 -3222
rect 1328 -3307 1329 -3285
rect 1360 -3307 1361 -3285
rect 219 -3307 220 -3287
rect 562 -3288 563 -3222
rect 821 -3307 822 -3287
rect 933 -3288 934 -3222
rect 1150 -3307 1151 -3287
rect 1255 -3307 1256 -3287
rect 506 -3290 507 -3222
rect 562 -3307 563 -3289
rect 856 -3290 857 -3222
rect 884 -3307 885 -3289
rect 915 -3307 916 -3289
rect 961 -3307 962 -3289
rect 1192 -3307 1193 -3289
rect 1402 -3290 1403 -3222
rect 506 -3307 507 -3291
rect 765 -3292 766 -3222
rect 856 -3307 857 -3291
rect 898 -3292 899 -3222
rect 926 -3292 927 -3222
rect 1024 -3307 1025 -3291
rect 765 -3307 766 -3293
rect 912 -3294 913 -3222
rect 926 -3307 927 -3293
rect 1066 -3294 1067 -3222
rect 863 -3296 864 -3222
rect 989 -3307 990 -3295
rect 1066 -3307 1067 -3295
rect 1213 -3307 1214 -3295
rect 639 -3298 640 -3222
rect 863 -3307 864 -3297
rect 912 -3307 913 -3297
rect 975 -3298 976 -3222
rect 639 -3307 640 -3299
rect 656 -3300 657 -3222
rect 933 -3307 934 -3299
rect 1108 -3300 1109 -3222
rect 835 -3307 836 -3301
rect 1108 -3307 1109 -3301
rect 975 -3307 976 -3303
rect 1122 -3304 1123 -3222
rect 1122 -3307 1123 -3305
rect 1451 -3306 1452 -3222
rect 131 -3317 132 -3315
rect 135 -3317 136 -3315
rect 163 -3317 164 -3315
rect 579 -3404 580 -3316
rect 590 -3317 591 -3315
rect 688 -3317 689 -3315
rect 691 -3317 692 -3315
rect 1157 -3317 1158 -3315
rect 1178 -3317 1179 -3315
rect 1528 -3317 1529 -3315
rect 1577 -3404 1578 -3316
rect 1584 -3317 1585 -3315
rect 205 -3319 206 -3315
rect 541 -3404 542 -3318
rect 590 -3404 591 -3318
rect 842 -3319 843 -3315
rect 870 -3319 871 -3315
rect 1192 -3319 1193 -3315
rect 1209 -3319 1210 -3315
rect 1276 -3319 1277 -3315
rect 1360 -3319 1361 -3315
rect 1374 -3404 1375 -3318
rect 1388 -3319 1389 -3315
rect 1388 -3404 1389 -3318
rect 1388 -3319 1389 -3315
rect 1388 -3404 1389 -3318
rect 233 -3321 234 -3315
rect 492 -3404 493 -3320
rect 506 -3321 507 -3315
rect 803 -3404 804 -3320
rect 870 -3404 871 -3320
rect 985 -3321 986 -3315
rect 1003 -3321 1004 -3315
rect 1108 -3321 1109 -3315
rect 1111 -3321 1112 -3315
rect 1290 -3321 1291 -3315
rect 212 -3323 213 -3315
rect 506 -3404 507 -3322
rect 513 -3323 514 -3315
rect 544 -3323 545 -3315
rect 614 -3404 615 -3322
rect 1150 -3323 1151 -3315
rect 1153 -3404 1154 -3322
rect 1234 -3323 1235 -3315
rect 1248 -3323 1249 -3315
rect 1325 -3323 1326 -3315
rect 247 -3325 248 -3315
rect 443 -3325 444 -3315
rect 464 -3325 465 -3315
rect 674 -3325 675 -3315
rect 705 -3325 706 -3315
rect 877 -3325 878 -3315
rect 880 -3325 881 -3315
rect 1136 -3325 1137 -3315
rect 1192 -3404 1193 -3324
rect 1283 -3325 1284 -3315
rect 198 -3327 199 -3315
rect 247 -3404 248 -3326
rect 268 -3327 269 -3315
rect 618 -3327 619 -3315
rect 621 -3327 622 -3315
rect 908 -3327 909 -3315
rect 915 -3327 916 -3315
rect 1143 -3327 1144 -3315
rect 1199 -3327 1200 -3315
rect 1248 -3404 1249 -3326
rect 1262 -3327 1263 -3315
rect 1311 -3327 1312 -3315
rect 240 -3329 241 -3315
rect 268 -3404 269 -3328
rect 310 -3329 311 -3315
rect 401 -3329 402 -3315
rect 429 -3329 430 -3315
rect 429 -3404 430 -3328
rect 429 -3329 430 -3315
rect 429 -3404 430 -3328
rect 436 -3404 437 -3328
rect 471 -3329 472 -3315
rect 485 -3329 486 -3315
rect 950 -3404 951 -3328
rect 961 -3329 962 -3315
rect 1157 -3404 1158 -3328
rect 1171 -3329 1172 -3315
rect 1199 -3404 1200 -3328
rect 1213 -3329 1214 -3315
rect 1241 -3329 1242 -3315
rect 1311 -3404 1312 -3328
rect 1332 -3329 1333 -3315
rect 177 -3331 178 -3315
rect 240 -3404 241 -3330
rect 359 -3331 360 -3315
rect 513 -3404 514 -3330
rect 523 -3404 524 -3330
rect 688 -3404 689 -3330
rect 716 -3331 717 -3315
rect 877 -3404 878 -3330
rect 894 -3404 895 -3330
rect 1216 -3331 1217 -3315
rect 1234 -3404 1235 -3330
rect 1318 -3331 1319 -3315
rect 1332 -3404 1333 -3330
rect 1381 -3331 1382 -3315
rect 359 -3404 360 -3332
rect 366 -3333 367 -3315
rect 380 -3333 381 -3315
rect 443 -3404 444 -3332
rect 471 -3404 472 -3332
rect 499 -3333 500 -3315
rect 618 -3404 619 -3332
rect 709 -3333 710 -3315
rect 716 -3404 717 -3332
rect 779 -3333 780 -3315
rect 789 -3333 790 -3315
rect 800 -3333 801 -3315
rect 901 -3333 902 -3315
rect 940 -3333 941 -3315
rect 947 -3333 948 -3315
rect 1136 -3404 1137 -3332
rect 1171 -3404 1172 -3332
rect 1297 -3333 1298 -3315
rect 1353 -3333 1354 -3315
rect 1381 -3404 1382 -3332
rect 170 -3335 171 -3315
rect 499 -3404 500 -3334
rect 632 -3335 633 -3315
rect 898 -3335 899 -3315
rect 947 -3404 948 -3334
rect 968 -3335 969 -3315
rect 982 -3335 983 -3315
rect 1164 -3335 1165 -3315
rect 1213 -3404 1214 -3334
rect 1318 -3404 1319 -3334
rect 275 -3337 276 -3315
rect 366 -3404 367 -3336
rect 380 -3404 381 -3336
rect 446 -3337 447 -3315
rect 478 -3337 479 -3315
rect 485 -3404 486 -3336
rect 632 -3404 633 -3336
rect 723 -3337 724 -3315
rect 730 -3337 731 -3315
rect 873 -3337 874 -3315
rect 898 -3404 899 -3336
rect 926 -3337 927 -3315
rect 961 -3404 962 -3336
rect 1101 -3337 1102 -3315
rect 1164 -3404 1165 -3336
rect 1269 -3337 1270 -3315
rect 394 -3339 395 -3315
rect 464 -3404 465 -3338
rect 478 -3404 479 -3338
rect 520 -3339 521 -3315
rect 639 -3339 640 -3315
rect 779 -3404 780 -3338
rect 891 -3339 892 -3315
rect 926 -3404 927 -3338
rect 982 -3404 983 -3338
rect 1122 -3339 1123 -3315
rect 1241 -3404 1242 -3338
rect 1339 -3339 1340 -3315
rect 345 -3341 346 -3315
rect 394 -3404 395 -3340
rect 401 -3404 402 -3340
rect 415 -3341 416 -3315
rect 576 -3341 577 -3315
rect 639 -3404 640 -3340
rect 667 -3341 668 -3315
rect 842 -3404 843 -3340
rect 996 -3341 997 -3315
rect 1101 -3404 1102 -3340
rect 282 -3343 283 -3315
rect 345 -3404 346 -3342
rect 548 -3343 549 -3315
rect 576 -3404 577 -3342
rect 667 -3404 668 -3342
rect 744 -3343 745 -3315
rect 758 -3343 759 -3315
rect 968 -3404 969 -3342
rect 1003 -3404 1004 -3342
rect 1087 -3343 1088 -3315
rect 1094 -3343 1095 -3315
rect 1122 -3404 1123 -3342
rect 184 -3345 185 -3315
rect 282 -3404 283 -3344
rect 317 -3345 318 -3315
rect 415 -3404 416 -3344
rect 530 -3345 531 -3315
rect 1087 -3404 1088 -3344
rect 226 -3347 227 -3315
rect 548 -3404 549 -3346
rect 583 -3347 584 -3315
rect 758 -3404 759 -3346
rect 863 -3347 864 -3315
rect 996 -3404 997 -3346
rect 1013 -3404 1014 -3346
rect 1220 -3347 1221 -3315
rect 219 -3349 220 -3315
rect 583 -3404 584 -3348
rect 674 -3404 675 -3348
rect 828 -3349 829 -3315
rect 1024 -3349 1025 -3315
rect 1129 -3349 1130 -3315
rect 317 -3404 318 -3350
rect 331 -3351 332 -3315
rect 408 -3351 409 -3315
rect 863 -3404 864 -3350
rect 1024 -3404 1025 -3350
rect 1227 -3351 1228 -3315
rect 296 -3353 297 -3315
rect 331 -3404 332 -3352
rect 373 -3353 374 -3315
rect 408 -3404 409 -3352
rect 709 -3404 710 -3352
rect 772 -3353 773 -3315
rect 828 -3404 829 -3352
rect 884 -3353 885 -3315
rect 1031 -3353 1032 -3315
rect 1034 -3359 1035 -3352
rect 1038 -3353 1039 -3315
rect 1185 -3353 1186 -3315
rect 191 -3355 192 -3315
rect 296 -3404 297 -3354
rect 660 -3355 661 -3315
rect 772 -3404 773 -3354
rect 814 -3355 815 -3315
rect 884 -3404 885 -3354
rect 989 -3355 990 -3315
rect 1038 -3404 1039 -3354
rect 1045 -3355 1046 -3315
rect 1143 -3404 1144 -3354
rect 1185 -3404 1186 -3354
rect 1206 -3355 1207 -3315
rect 261 -3357 262 -3315
rect 373 -3404 374 -3356
rect 660 -3404 661 -3356
rect 765 -3357 766 -3315
rect 849 -3357 850 -3315
rect 989 -3404 990 -3356
rect 1031 -3404 1032 -3356
rect 1115 -3357 1116 -3315
rect 1206 -3404 1207 -3356
rect 1251 -3357 1252 -3315
rect 681 -3359 682 -3315
rect 814 -3404 815 -3358
rect 1115 -3404 1116 -3358
rect 681 -3404 682 -3360
rect 1062 -3404 1063 -3360
rect 1066 -3361 1067 -3315
rect 1094 -3404 1095 -3360
rect 702 -3363 703 -3315
rect 765 -3404 766 -3362
rect 786 -3363 787 -3315
rect 849 -3404 850 -3362
rect 1045 -3404 1046 -3362
rect 1073 -3363 1074 -3315
rect 1080 -3363 1081 -3315
rect 1129 -3404 1130 -3362
rect 646 -3365 647 -3315
rect 702 -3404 703 -3364
rect 723 -3404 724 -3364
rect 793 -3365 794 -3315
rect 856 -3365 857 -3315
rect 1080 -3404 1081 -3364
rect 611 -3367 612 -3315
rect 793 -3404 794 -3366
rect 856 -3404 857 -3366
rect 1167 -3404 1168 -3366
rect 254 -3369 255 -3315
rect 611 -3404 612 -3368
rect 646 -3404 647 -3368
rect 751 -3369 752 -3315
rect 786 -3404 787 -3368
rect 800 -3404 801 -3368
rect 933 -3369 934 -3315
rect 1073 -3404 1074 -3368
rect 737 -3371 738 -3315
rect 940 -3404 941 -3370
rect 1052 -3371 1053 -3315
rect 1108 -3404 1109 -3370
rect 737 -3404 738 -3372
rect 807 -3373 808 -3315
rect 933 -3404 934 -3372
rect 1020 -3373 1021 -3315
rect 1066 -3404 1067 -3372
rect 1265 -3373 1266 -3315
rect 387 -3375 388 -3315
rect 1020 -3404 1021 -3374
rect 1265 -3404 1266 -3374
rect 1346 -3375 1347 -3315
rect 387 -3404 388 -3376
rect 457 -3377 458 -3315
rect 597 -3377 598 -3315
rect 807 -3404 808 -3376
rect 450 -3379 451 -3315
rect 457 -3404 458 -3378
rect 597 -3404 598 -3378
rect 695 -3379 696 -3315
rect 744 -3404 745 -3378
rect 821 -3379 822 -3315
rect 450 -3404 451 -3380
rect 527 -3381 528 -3315
rect 695 -3404 696 -3380
rect 835 -3381 836 -3315
rect 527 -3404 528 -3382
rect 534 -3383 535 -3315
rect 562 -3383 563 -3315
rect 835 -3404 836 -3382
rect 534 -3404 535 -3384
rect 555 -3385 556 -3315
rect 562 -3404 563 -3384
rect 569 -3385 570 -3315
rect 751 -3404 752 -3384
rect 912 -3385 913 -3315
rect 555 -3404 556 -3386
rect 625 -3387 626 -3315
rect 821 -3404 822 -3386
rect 919 -3387 920 -3315
rect 569 -3404 570 -3388
rect 604 -3389 605 -3315
rect 625 -3404 626 -3388
rect 653 -3389 654 -3315
rect 912 -3404 913 -3388
rect 954 -3389 955 -3315
rect 422 -3391 423 -3315
rect 653 -3404 654 -3390
rect 919 -3404 920 -3390
rect 975 -3391 976 -3315
rect 338 -3393 339 -3315
rect 422 -3404 423 -3392
rect 604 -3404 605 -3392
rect 905 -3393 906 -3315
rect 954 -3404 955 -3392
rect 1017 -3404 1018 -3392
rect 338 -3404 339 -3394
rect 352 -3395 353 -3315
rect 905 -3404 906 -3394
rect 1010 -3395 1011 -3315
rect 324 -3397 325 -3315
rect 352 -3404 353 -3396
rect 975 -3404 976 -3396
rect 1059 -3397 1060 -3315
rect 303 -3399 304 -3315
rect 324 -3404 325 -3398
rect 1059 -3404 1060 -3398
rect 1304 -3399 1305 -3315
rect 289 -3401 290 -3315
rect 303 -3404 304 -3400
rect 289 -3404 290 -3402
rect 310 -3404 311 -3402
rect 240 -3414 241 -3412
rect 261 -3451 262 -3413
rect 268 -3414 269 -3412
rect 292 -3414 293 -3412
rect 338 -3414 339 -3412
rect 355 -3451 356 -3413
rect 376 -3414 377 -3412
rect 450 -3414 451 -3412
rect 457 -3414 458 -3412
rect 474 -3451 475 -3413
rect 485 -3414 486 -3412
rect 611 -3451 612 -3413
rect 632 -3414 633 -3412
rect 632 -3451 633 -3413
rect 632 -3414 633 -3412
rect 632 -3451 633 -3413
rect 639 -3414 640 -3412
rect 639 -3451 640 -3413
rect 639 -3414 640 -3412
rect 639 -3451 640 -3413
rect 663 -3451 664 -3413
rect 1038 -3414 1039 -3412
rect 1041 -3414 1042 -3412
rect 1045 -3414 1046 -3412
rect 1052 -3451 1053 -3413
rect 1073 -3414 1074 -3412
rect 1111 -3414 1112 -3412
rect 1192 -3414 1193 -3412
rect 1199 -3414 1200 -3412
rect 1213 -3414 1214 -3412
rect 1248 -3414 1249 -3412
rect 1269 -3451 1270 -3413
rect 1304 -3451 1305 -3413
rect 1311 -3414 1312 -3412
rect 1318 -3414 1319 -3412
rect 1346 -3451 1347 -3413
rect 1374 -3414 1375 -3412
rect 1395 -3451 1396 -3413
rect 1577 -3414 1578 -3412
rect 1577 -3451 1578 -3413
rect 1577 -3414 1578 -3412
rect 1577 -3451 1578 -3413
rect 247 -3416 248 -3412
rect 289 -3416 290 -3412
rect 317 -3416 318 -3412
rect 457 -3451 458 -3415
rect 499 -3416 500 -3412
rect 604 -3416 605 -3412
rect 688 -3416 689 -3412
rect 688 -3451 689 -3415
rect 688 -3416 689 -3412
rect 688 -3451 689 -3415
rect 702 -3416 703 -3412
rect 810 -3451 811 -3415
rect 824 -3451 825 -3415
rect 982 -3416 983 -3412
rect 989 -3416 990 -3412
rect 1055 -3416 1056 -3412
rect 1073 -3451 1074 -3415
rect 1101 -3416 1102 -3412
rect 1122 -3416 1123 -3412
rect 1125 -3436 1126 -3415
rect 1129 -3416 1130 -3412
rect 1160 -3416 1161 -3412
rect 1185 -3416 1186 -3412
rect 1192 -3451 1193 -3415
rect 1318 -3451 1319 -3415
rect 1332 -3416 1333 -3412
rect 1381 -3416 1382 -3412
rect 1384 -3416 1385 -3412
rect 282 -3418 283 -3412
rect 317 -3451 318 -3417
rect 324 -3418 325 -3412
rect 338 -3451 339 -3417
rect 352 -3418 353 -3412
rect 373 -3451 374 -3417
rect 394 -3418 395 -3412
rect 499 -3451 500 -3417
rect 513 -3418 514 -3412
rect 656 -3451 657 -3417
rect 702 -3451 703 -3417
rect 737 -3418 738 -3412
rect 793 -3418 794 -3412
rect 803 -3418 804 -3412
rect 863 -3418 864 -3412
rect 1265 -3418 1266 -3412
rect 1381 -3451 1382 -3417
rect 1388 -3418 1389 -3412
rect 366 -3420 367 -3412
rect 394 -3451 395 -3419
rect 415 -3420 416 -3412
rect 513 -3451 514 -3419
rect 520 -3420 521 -3412
rect 527 -3420 528 -3412
rect 562 -3420 563 -3412
rect 730 -3420 731 -3412
rect 733 -3420 734 -3412
rect 786 -3420 787 -3412
rect 800 -3451 801 -3419
rect 814 -3420 815 -3412
rect 842 -3420 843 -3412
rect 863 -3451 864 -3419
rect 884 -3420 885 -3412
rect 891 -3420 892 -3412
rect 898 -3420 899 -3412
rect 999 -3451 1000 -3419
rect 1017 -3420 1018 -3412
rect 1031 -3420 1032 -3412
rect 1080 -3420 1081 -3412
rect 1199 -3451 1200 -3419
rect 359 -3422 360 -3412
rect 520 -3451 521 -3421
rect 562 -3451 563 -3421
rect 590 -3422 591 -3412
rect 625 -3422 626 -3412
rect 730 -3451 731 -3421
rect 751 -3422 752 -3412
rect 884 -3451 885 -3421
rect 898 -3451 899 -3421
rect 905 -3422 906 -3412
rect 919 -3422 920 -3412
rect 989 -3451 990 -3421
rect 996 -3422 997 -3412
rect 1010 -3422 1011 -3412
rect 1024 -3422 1025 -3412
rect 1171 -3422 1172 -3412
rect 359 -3451 360 -3423
rect 509 -3451 510 -3423
rect 569 -3424 570 -3412
rect 569 -3451 570 -3423
rect 569 -3424 570 -3412
rect 569 -3451 570 -3423
rect 576 -3451 577 -3423
rect 597 -3424 598 -3412
rect 625 -3451 626 -3423
rect 646 -3424 647 -3412
rect 681 -3424 682 -3412
rect 737 -3451 738 -3423
rect 758 -3424 759 -3412
rect 786 -3451 787 -3423
rect 807 -3424 808 -3412
rect 842 -3451 843 -3423
rect 849 -3424 850 -3412
rect 891 -3451 892 -3423
rect 919 -3451 920 -3423
rect 961 -3424 962 -3412
rect 968 -3424 969 -3412
rect 1167 -3424 1168 -3412
rect 366 -3451 367 -3425
rect 387 -3426 388 -3412
rect 415 -3451 416 -3425
rect 436 -3426 437 -3412
rect 443 -3426 444 -3412
rect 586 -3451 587 -3425
rect 597 -3451 598 -3425
rect 695 -3426 696 -3412
rect 751 -3451 752 -3425
rect 849 -3451 850 -3425
rect 877 -3426 878 -3412
rect 1010 -3451 1011 -3425
rect 1031 -3451 1032 -3425
rect 1150 -3426 1151 -3412
rect 1153 -3426 1154 -3412
rect 1206 -3426 1207 -3412
rect 303 -3428 304 -3412
rect 443 -3451 444 -3427
rect 450 -3451 451 -3427
rect 478 -3428 479 -3412
rect 492 -3428 493 -3412
rect 604 -3451 605 -3427
rect 618 -3428 619 -3412
rect 695 -3451 696 -3427
rect 758 -3451 759 -3427
rect 821 -3428 822 -3412
rect 877 -3451 878 -3427
rect 894 -3428 895 -3412
rect 940 -3428 941 -3412
rect 1017 -3451 1018 -3427
rect 1087 -3428 1088 -3412
rect 1213 -3451 1214 -3427
rect 380 -3430 381 -3412
rect 387 -3451 388 -3429
rect 408 -3430 409 -3412
rect 436 -3451 437 -3429
rect 464 -3430 465 -3412
rect 527 -3451 528 -3429
rect 548 -3430 549 -3412
rect 807 -3451 808 -3429
rect 814 -3451 815 -3429
rect 828 -3430 829 -3412
rect 912 -3430 913 -3412
rect 940 -3451 941 -3429
rect 954 -3430 955 -3412
rect 982 -3451 983 -3429
rect 1003 -3430 1004 -3412
rect 1024 -3451 1025 -3429
rect 1101 -3451 1102 -3429
rect 1115 -3430 1116 -3412
rect 1122 -3451 1123 -3429
rect 1136 -3430 1137 -3412
rect 1157 -3430 1158 -3412
rect 1234 -3430 1235 -3412
rect 331 -3432 332 -3412
rect 380 -3451 381 -3431
rect 401 -3432 402 -3412
rect 464 -3451 465 -3431
rect 471 -3432 472 -3412
rect 478 -3451 479 -3431
rect 492 -3451 493 -3431
rect 534 -3432 535 -3412
rect 548 -3451 549 -3431
rect 555 -3432 556 -3412
rect 579 -3432 580 -3412
rect 1080 -3451 1081 -3431
rect 1094 -3432 1095 -3412
rect 1115 -3451 1116 -3431
rect 1129 -3451 1130 -3431
rect 1300 -3451 1301 -3431
rect 299 -3434 300 -3412
rect 401 -3451 402 -3433
rect 422 -3434 423 -3412
rect 523 -3434 524 -3412
rect 534 -3451 535 -3433
rect 541 -3434 542 -3412
rect 646 -3451 647 -3433
rect 660 -3434 661 -3412
rect 681 -3451 682 -3433
rect 709 -3434 710 -3412
rect 772 -3434 773 -3412
rect 905 -3451 906 -3433
rect 912 -3451 913 -3433
rect 926 -3434 927 -3412
rect 933 -3434 934 -3412
rect 954 -3451 955 -3433
rect 961 -3451 962 -3433
rect 975 -3434 976 -3412
rect 1003 -3451 1004 -3433
rect 1066 -3434 1067 -3412
rect 1136 -3451 1137 -3433
rect 1206 -3451 1207 -3433
rect 1241 -3434 1242 -3412
rect 345 -3436 346 -3412
rect 422 -3451 423 -3435
rect 429 -3436 430 -3412
rect 429 -3451 430 -3435
rect 429 -3436 430 -3412
rect 429 -3451 430 -3435
rect 471 -3451 472 -3435
rect 541 -3451 542 -3435
rect 709 -3451 710 -3435
rect 744 -3436 745 -3412
rect 765 -3436 766 -3412
rect 975 -3451 976 -3435
rect 1384 -3451 1385 -3435
rect 1388 -3451 1389 -3435
rect 310 -3438 311 -3412
rect 345 -3451 346 -3437
rect 485 -3451 486 -3437
rect 660 -3451 661 -3437
rect 716 -3438 717 -3412
rect 765 -3451 766 -3437
rect 779 -3438 780 -3412
rect 793 -3451 794 -3437
rect 821 -3451 822 -3437
rect 1216 -3438 1217 -3412
rect 310 -3451 311 -3439
rect 352 -3451 353 -3439
rect 506 -3440 507 -3412
rect 555 -3451 556 -3439
rect 653 -3440 654 -3412
rect 779 -3451 780 -3439
rect 828 -3451 829 -3439
rect 835 -3440 836 -3412
rect 933 -3451 934 -3439
rect 996 -3451 997 -3439
rect 506 -3451 507 -3441
rect 621 -3451 622 -3441
rect 674 -3442 675 -3412
rect 716 -3451 717 -3441
rect 723 -3442 724 -3412
rect 772 -3451 773 -3441
rect 835 -3451 836 -3441
rect 947 -3442 948 -3412
rect 667 -3444 668 -3412
rect 674 -3451 675 -3443
rect 723 -3451 724 -3443
rect 852 -3451 853 -3443
rect 870 -3444 871 -3412
rect 947 -3451 948 -3443
rect 614 -3446 615 -3412
rect 667 -3451 668 -3445
rect 744 -3451 745 -3445
rect 856 -3446 857 -3412
rect 870 -3451 871 -3445
rect 1020 -3446 1021 -3412
rect 583 -3448 584 -3412
rect 856 -3451 857 -3447
rect 583 -3451 584 -3449
rect 926 -3451 927 -3449
rect 261 -3461 262 -3459
rect 268 -3492 269 -3460
rect 296 -3492 297 -3460
rect 310 -3461 311 -3459
rect 317 -3461 318 -3459
rect 355 -3461 356 -3459
rect 359 -3461 360 -3459
rect 411 -3461 412 -3459
rect 439 -3492 440 -3460
rect 656 -3492 657 -3460
rect 660 -3461 661 -3459
rect 733 -3492 734 -3460
rect 737 -3461 738 -3459
rect 737 -3492 738 -3460
rect 737 -3461 738 -3459
rect 737 -3492 738 -3460
rect 793 -3461 794 -3459
rect 793 -3492 794 -3460
rect 793 -3461 794 -3459
rect 793 -3492 794 -3460
rect 800 -3461 801 -3459
rect 807 -3461 808 -3459
rect 821 -3461 822 -3459
rect 828 -3461 829 -3459
rect 842 -3461 843 -3459
rect 915 -3492 916 -3460
rect 933 -3461 934 -3459
rect 933 -3492 934 -3460
rect 933 -3461 934 -3459
rect 933 -3492 934 -3460
rect 940 -3461 941 -3459
rect 943 -3469 944 -3460
rect 947 -3461 948 -3459
rect 1006 -3492 1007 -3460
rect 1010 -3461 1011 -3459
rect 1059 -3492 1060 -3460
rect 1066 -3492 1067 -3460
rect 1073 -3461 1074 -3459
rect 1087 -3492 1088 -3460
rect 1101 -3461 1102 -3459
rect 1115 -3461 1116 -3459
rect 1118 -3461 1119 -3459
rect 1136 -3461 1137 -3459
rect 1136 -3492 1137 -3460
rect 1136 -3461 1137 -3459
rect 1136 -3492 1137 -3460
rect 1143 -3461 1144 -3459
rect 1157 -3492 1158 -3460
rect 1181 -3492 1182 -3460
rect 1416 -3492 1417 -3460
rect 1577 -3461 1578 -3459
rect 1577 -3492 1578 -3460
rect 1577 -3461 1578 -3459
rect 1577 -3492 1578 -3460
rect 373 -3463 374 -3459
rect 390 -3492 391 -3462
rect 401 -3463 402 -3459
rect 583 -3463 584 -3459
rect 604 -3463 605 -3459
rect 604 -3492 605 -3462
rect 604 -3463 605 -3459
rect 604 -3492 605 -3462
rect 611 -3463 612 -3459
rect 719 -3463 720 -3459
rect 786 -3463 787 -3459
rect 800 -3492 801 -3462
rect 807 -3492 808 -3462
rect 814 -3463 815 -3459
rect 828 -3492 829 -3462
rect 870 -3463 871 -3459
rect 877 -3463 878 -3459
rect 877 -3492 878 -3462
rect 877 -3463 878 -3459
rect 877 -3492 878 -3462
rect 940 -3492 941 -3462
rect 961 -3463 962 -3459
rect 968 -3463 969 -3459
rect 982 -3463 983 -3459
rect 989 -3463 990 -3459
rect 1010 -3492 1011 -3462
rect 1017 -3463 1018 -3459
rect 1045 -3492 1046 -3462
rect 1052 -3463 1053 -3459
rect 1052 -3492 1053 -3462
rect 1052 -3463 1053 -3459
rect 1052 -3492 1053 -3462
rect 1073 -3492 1074 -3462
rect 1129 -3463 1130 -3459
rect 1185 -3492 1186 -3462
rect 1206 -3463 1207 -3459
rect 1213 -3463 1214 -3459
rect 1248 -3492 1249 -3462
rect 1269 -3463 1270 -3459
rect 1276 -3492 1277 -3462
rect 1297 -3463 1298 -3459
rect 1318 -3463 1319 -3459
rect 1374 -3492 1375 -3462
rect 1381 -3463 1382 -3459
rect 1388 -3463 1389 -3459
rect 1388 -3492 1389 -3462
rect 1388 -3463 1389 -3459
rect 1388 -3492 1389 -3462
rect 1395 -3463 1396 -3459
rect 1395 -3492 1396 -3462
rect 1395 -3463 1396 -3459
rect 1395 -3492 1396 -3462
rect 345 -3465 346 -3459
rect 373 -3492 374 -3464
rect 380 -3465 381 -3459
rect 408 -3492 409 -3464
rect 485 -3465 486 -3459
rect 485 -3492 486 -3464
rect 485 -3465 486 -3459
rect 485 -3492 486 -3464
rect 520 -3465 521 -3459
rect 590 -3465 591 -3459
rect 618 -3465 619 -3459
rect 625 -3465 626 -3459
rect 632 -3465 633 -3459
rect 663 -3465 664 -3459
rect 667 -3465 668 -3459
rect 754 -3492 755 -3464
rect 765 -3465 766 -3459
rect 786 -3492 787 -3464
rect 852 -3465 853 -3459
rect 919 -3465 920 -3459
rect 961 -3492 962 -3464
rect 975 -3465 976 -3459
rect 1038 -3492 1039 -3464
rect 1080 -3465 1081 -3459
rect 1269 -3492 1270 -3464
rect 1300 -3465 1301 -3459
rect 1304 -3465 1305 -3459
rect 1346 -3465 1347 -3459
rect 1381 -3492 1382 -3464
rect 366 -3467 367 -3459
rect 380 -3492 381 -3466
rect 387 -3467 388 -3459
rect 425 -3492 426 -3466
rect 506 -3467 507 -3459
rect 590 -3492 591 -3466
rect 618 -3492 619 -3466
rect 723 -3467 724 -3459
rect 758 -3467 759 -3459
rect 765 -3492 766 -3466
rect 772 -3467 773 -3459
rect 814 -3492 815 -3466
rect 856 -3467 857 -3459
rect 947 -3492 948 -3466
rect 975 -3492 976 -3466
rect 1003 -3467 1004 -3459
rect 1024 -3467 1025 -3459
rect 1024 -3492 1025 -3466
rect 1024 -3467 1025 -3459
rect 1024 -3492 1025 -3466
rect 1115 -3492 1116 -3466
rect 1122 -3467 1123 -3459
rect 1192 -3467 1193 -3459
rect 1192 -3492 1193 -3466
rect 1192 -3467 1193 -3459
rect 1192 -3492 1193 -3466
rect 1199 -3467 1200 -3459
rect 1234 -3492 1235 -3466
rect 338 -3469 339 -3459
rect 366 -3492 367 -3468
rect 450 -3469 451 -3459
rect 506 -3492 507 -3468
rect 527 -3469 528 -3459
rect 621 -3469 622 -3459
rect 639 -3469 640 -3459
rect 639 -3492 640 -3468
rect 639 -3469 640 -3459
rect 639 -3492 640 -3468
rect 653 -3469 654 -3459
rect 681 -3469 682 -3459
rect 695 -3469 696 -3459
rect 758 -3492 759 -3468
rect 891 -3469 892 -3459
rect 919 -3492 920 -3468
rect 926 -3469 927 -3459
rect 1080 -3492 1081 -3468
rect 1118 -3492 1119 -3468
rect 1122 -3492 1123 -3468
rect 429 -3471 430 -3459
rect 450 -3492 451 -3470
rect 499 -3471 500 -3459
rect 527 -3492 528 -3470
rect 534 -3471 535 -3459
rect 632 -3492 633 -3470
rect 653 -3492 654 -3470
rect 1090 -3492 1091 -3470
rect 394 -3473 395 -3459
rect 429 -3492 430 -3472
rect 457 -3473 458 -3459
rect 499 -3492 500 -3472
rect 534 -3492 535 -3472
rect 607 -3473 608 -3459
rect 695 -3492 696 -3472
rect 744 -3473 745 -3459
rect 884 -3473 885 -3459
rect 891 -3492 892 -3472
rect 905 -3473 906 -3459
rect 926 -3492 927 -3472
rect 1003 -3492 1004 -3472
rect 1178 -3492 1179 -3472
rect 436 -3475 437 -3459
rect 457 -3492 458 -3474
rect 541 -3475 542 -3459
rect 586 -3475 587 -3459
rect 702 -3475 703 -3459
rect 716 -3492 717 -3474
rect 723 -3492 724 -3474
rect 751 -3475 752 -3459
rect 863 -3475 864 -3459
rect 884 -3492 885 -3474
rect 898 -3475 899 -3459
rect 905 -3492 906 -3474
rect 478 -3477 479 -3459
rect 541 -3492 542 -3476
rect 548 -3477 549 -3459
rect 593 -3477 594 -3459
rect 688 -3477 689 -3459
rect 702 -3492 703 -3476
rect 709 -3477 710 -3459
rect 821 -3492 822 -3476
rect 898 -3492 899 -3476
rect 912 -3477 913 -3459
rect 464 -3479 465 -3459
rect 478 -3492 479 -3478
rect 548 -3492 549 -3478
rect 576 -3479 577 -3459
rect 646 -3479 647 -3459
rect 709 -3492 710 -3478
rect 730 -3479 731 -3459
rect 772 -3492 773 -3478
rect 779 -3479 780 -3459
rect 912 -3492 913 -3478
rect 555 -3481 556 -3459
rect 583 -3492 584 -3480
rect 674 -3481 675 -3459
rect 688 -3492 689 -3480
rect 730 -3492 731 -3480
rect 835 -3481 836 -3459
rect 492 -3483 493 -3459
rect 555 -3492 556 -3482
rect 562 -3483 563 -3459
rect 576 -3492 577 -3482
rect 744 -3492 745 -3482
rect 996 -3483 997 -3459
rect 443 -3485 444 -3459
rect 492 -3492 493 -3484
rect 513 -3485 514 -3459
rect 562 -3492 563 -3484
rect 569 -3485 570 -3459
rect 646 -3492 647 -3484
rect 996 -3492 997 -3484
rect 1031 -3485 1032 -3459
rect 415 -3487 416 -3459
rect 443 -3492 444 -3486
rect 569 -3492 570 -3486
rect 597 -3487 598 -3459
rect 422 -3489 423 -3459
rect 513 -3492 514 -3488
rect 422 -3492 423 -3490
rect 471 -3492 472 -3490
rect 268 -3502 269 -3500
rect 282 -3502 283 -3500
rect 285 -3502 286 -3500
rect 296 -3502 297 -3500
rect 366 -3502 367 -3500
rect 387 -3523 388 -3501
rect 390 -3502 391 -3500
rect 394 -3523 395 -3501
rect 408 -3502 409 -3500
rect 439 -3502 440 -3500
rect 450 -3502 451 -3500
rect 481 -3523 482 -3501
rect 506 -3502 507 -3500
rect 565 -3523 566 -3501
rect 583 -3502 584 -3500
rect 597 -3523 598 -3501
rect 604 -3502 605 -3500
rect 604 -3523 605 -3501
rect 604 -3502 605 -3500
rect 604 -3523 605 -3501
rect 632 -3502 633 -3500
rect 726 -3502 727 -3500
rect 733 -3502 734 -3500
rect 1181 -3502 1182 -3500
rect 1192 -3502 1193 -3500
rect 1192 -3523 1193 -3501
rect 1192 -3502 1193 -3500
rect 1192 -3523 1193 -3501
rect 1234 -3502 1235 -3500
rect 1279 -3523 1280 -3501
rect 1374 -3502 1375 -3500
rect 1381 -3523 1382 -3501
rect 1384 -3502 1385 -3500
rect 1388 -3502 1389 -3500
rect 1395 -3502 1396 -3500
rect 1395 -3523 1396 -3501
rect 1395 -3502 1396 -3500
rect 1395 -3523 1396 -3501
rect 1416 -3502 1417 -3500
rect 1500 -3523 1501 -3501
rect 1577 -3502 1578 -3500
rect 1577 -3523 1578 -3501
rect 1577 -3502 1578 -3500
rect 1577 -3523 1578 -3501
rect 373 -3504 374 -3500
rect 401 -3523 402 -3503
rect 443 -3504 444 -3500
rect 450 -3523 451 -3503
rect 457 -3504 458 -3500
rect 464 -3523 465 -3503
rect 492 -3504 493 -3500
rect 506 -3523 507 -3503
rect 520 -3523 521 -3503
rect 548 -3504 549 -3500
rect 562 -3504 563 -3500
rect 583 -3523 584 -3503
rect 590 -3504 591 -3500
rect 656 -3504 657 -3500
rect 674 -3523 675 -3503
rect 695 -3504 696 -3500
rect 702 -3504 703 -3500
rect 702 -3523 703 -3503
rect 702 -3504 703 -3500
rect 702 -3523 703 -3503
rect 737 -3504 738 -3500
rect 754 -3504 755 -3500
rect 758 -3504 759 -3500
rect 779 -3523 780 -3503
rect 786 -3504 787 -3500
rect 789 -3512 790 -3503
rect 821 -3504 822 -3500
rect 863 -3523 864 -3503
rect 905 -3504 906 -3500
rect 912 -3504 913 -3500
rect 940 -3504 941 -3500
rect 940 -3523 941 -3503
rect 940 -3504 941 -3500
rect 940 -3523 941 -3503
rect 947 -3504 948 -3500
rect 1034 -3523 1035 -3503
rect 1045 -3504 1046 -3500
rect 1048 -3504 1049 -3500
rect 1059 -3504 1060 -3500
rect 1090 -3504 1091 -3500
rect 1115 -3504 1116 -3500
rect 1115 -3523 1116 -3503
rect 1115 -3504 1116 -3500
rect 1115 -3523 1116 -3503
rect 1122 -3504 1123 -3500
rect 1129 -3523 1130 -3503
rect 1136 -3504 1137 -3500
rect 1136 -3523 1137 -3503
rect 1136 -3504 1137 -3500
rect 1136 -3523 1137 -3503
rect 1157 -3504 1158 -3500
rect 1164 -3523 1165 -3503
rect 1178 -3523 1179 -3503
rect 1185 -3504 1186 -3500
rect 1248 -3504 1249 -3500
rect 1262 -3523 1263 -3503
rect 1269 -3504 1270 -3500
rect 1339 -3523 1340 -3503
rect 380 -3506 381 -3500
rect 380 -3523 381 -3505
rect 380 -3506 381 -3500
rect 380 -3523 381 -3505
rect 429 -3506 430 -3500
rect 443 -3523 444 -3505
rect 478 -3506 479 -3500
rect 492 -3523 493 -3505
rect 527 -3506 528 -3500
rect 558 -3523 559 -3505
rect 576 -3506 577 -3500
rect 590 -3523 591 -3505
rect 646 -3506 647 -3500
rect 730 -3506 731 -3500
rect 758 -3523 759 -3505
rect 772 -3506 773 -3500
rect 786 -3523 787 -3505
rect 800 -3506 801 -3500
rect 821 -3523 822 -3505
rect 842 -3523 843 -3505
rect 1017 -3523 1018 -3505
rect 1020 -3523 1021 -3505
rect 1073 -3506 1074 -3500
rect 1080 -3506 1081 -3500
rect 1143 -3523 1144 -3505
rect 1276 -3506 1277 -3500
rect 1276 -3523 1277 -3505
rect 1276 -3506 1277 -3500
rect 1276 -3523 1277 -3505
rect 429 -3523 430 -3507
rect 478 -3523 479 -3507
rect 499 -3508 500 -3500
rect 527 -3523 528 -3507
rect 541 -3508 542 -3500
rect 548 -3523 549 -3507
rect 576 -3523 577 -3507
rect 618 -3508 619 -3500
rect 639 -3508 640 -3500
rect 646 -3523 647 -3507
rect 653 -3523 654 -3507
rect 744 -3508 745 -3500
rect 765 -3508 766 -3500
rect 772 -3523 773 -3507
rect 800 -3523 801 -3507
rect 807 -3508 808 -3500
rect 884 -3508 885 -3500
rect 905 -3523 906 -3507
rect 957 -3523 958 -3507
rect 996 -3508 997 -3500
rect 1003 -3508 1004 -3500
rect 1003 -3523 1004 -3507
rect 1003 -3508 1004 -3500
rect 1003 -3523 1004 -3507
rect 1010 -3508 1011 -3500
rect 1041 -3523 1042 -3507
rect 1045 -3523 1046 -3507
rect 1052 -3508 1053 -3500
rect 1062 -3523 1063 -3507
rect 1066 -3508 1067 -3500
rect 485 -3510 486 -3500
rect 499 -3523 500 -3509
rect 513 -3510 514 -3500
rect 541 -3523 542 -3509
rect 688 -3510 689 -3500
rect 695 -3523 696 -3509
rect 709 -3510 710 -3500
rect 730 -3523 731 -3509
rect 807 -3523 808 -3509
rect 814 -3510 815 -3500
rect 877 -3510 878 -3500
rect 884 -3523 885 -3509
rect 961 -3510 962 -3500
rect 964 -3523 965 -3509
rect 968 -3523 969 -3509
rect 975 -3510 976 -3500
rect 1024 -3510 1025 -3500
rect 1031 -3523 1032 -3509
rect 1038 -3510 1039 -3500
rect 1073 -3523 1074 -3509
rect 471 -3512 472 -3500
rect 485 -3523 486 -3511
rect 513 -3523 514 -3511
rect 534 -3512 535 -3500
rect 709 -3523 710 -3511
rect 716 -3512 717 -3500
rect 765 -3523 766 -3511
rect 1038 -3523 1039 -3511
rect 1048 -3523 1049 -3511
rect 1052 -3523 1053 -3511
rect 534 -3523 535 -3513
rect 569 -3514 570 -3500
rect 814 -3523 815 -3513
rect 828 -3514 829 -3500
rect 877 -3523 878 -3513
rect 898 -3514 899 -3500
rect 954 -3514 955 -3500
rect 961 -3523 962 -3513
rect 555 -3516 556 -3500
rect 569 -3523 570 -3515
rect 891 -3516 892 -3500
rect 898 -3523 899 -3515
rect 926 -3516 927 -3500
rect 954 -3523 955 -3515
rect 926 -3523 927 -3517
rect 933 -3518 934 -3500
rect 919 -3520 920 -3500
rect 933 -3523 934 -3519
rect 919 -3523 920 -3521
rect 947 -3523 948 -3521
rect 380 -3533 381 -3531
rect 380 -3552 381 -3532
rect 380 -3533 381 -3531
rect 380 -3552 381 -3532
rect 387 -3533 388 -3531
rect 390 -3539 391 -3532
rect 408 -3552 409 -3532
rect 429 -3533 430 -3531
rect 450 -3533 451 -3531
rect 457 -3552 458 -3532
rect 464 -3533 465 -3531
rect 474 -3552 475 -3532
rect 478 -3533 479 -3531
rect 478 -3552 479 -3532
rect 478 -3533 479 -3531
rect 478 -3552 479 -3532
rect 506 -3533 507 -3531
rect 520 -3533 521 -3531
rect 527 -3533 528 -3531
rect 527 -3552 528 -3532
rect 527 -3533 528 -3531
rect 527 -3552 528 -3532
rect 548 -3533 549 -3531
rect 548 -3552 549 -3532
rect 548 -3533 549 -3531
rect 548 -3552 549 -3532
rect 558 -3533 559 -3531
rect 1108 -3552 1109 -3532
rect 1115 -3533 1116 -3531
rect 1115 -3552 1116 -3532
rect 1115 -3533 1116 -3531
rect 1115 -3552 1116 -3532
rect 1129 -3533 1130 -3531
rect 1129 -3552 1130 -3532
rect 1129 -3533 1130 -3531
rect 1129 -3552 1130 -3532
rect 1136 -3533 1137 -3531
rect 1136 -3552 1137 -3532
rect 1136 -3533 1137 -3531
rect 1136 -3552 1137 -3532
rect 1157 -3533 1158 -3531
rect 1164 -3533 1165 -3531
rect 1178 -3533 1179 -3531
rect 1178 -3552 1179 -3532
rect 1178 -3533 1179 -3531
rect 1178 -3552 1179 -3532
rect 1192 -3533 1193 -3531
rect 1192 -3552 1193 -3532
rect 1192 -3533 1193 -3531
rect 1192 -3552 1193 -3532
rect 1262 -3533 1263 -3531
rect 1279 -3533 1280 -3531
rect 1339 -3533 1340 -3531
rect 1360 -3552 1361 -3532
rect 1381 -3533 1382 -3531
rect 1388 -3552 1389 -3532
rect 1395 -3533 1396 -3531
rect 1395 -3552 1396 -3532
rect 1395 -3533 1396 -3531
rect 1395 -3552 1396 -3532
rect 1500 -3533 1501 -3531
rect 1580 -3533 1581 -3531
rect 387 -3552 388 -3534
rect 401 -3535 402 -3531
rect 443 -3535 444 -3531
rect 450 -3552 451 -3534
rect 506 -3552 507 -3534
rect 513 -3535 514 -3531
rect 565 -3535 566 -3531
rect 653 -3535 654 -3531
rect 660 -3552 661 -3534
rect 674 -3535 675 -3531
rect 695 -3535 696 -3531
rect 705 -3552 706 -3534
rect 730 -3535 731 -3531
rect 737 -3552 738 -3534
rect 758 -3535 759 -3531
rect 758 -3552 759 -3534
rect 758 -3535 759 -3531
rect 758 -3552 759 -3534
rect 786 -3535 787 -3531
rect 786 -3552 787 -3534
rect 786 -3535 787 -3531
rect 786 -3552 787 -3534
rect 796 -3552 797 -3534
rect 800 -3535 801 -3531
rect 807 -3535 808 -3531
rect 824 -3535 825 -3531
rect 884 -3535 885 -3531
rect 891 -3535 892 -3531
rect 898 -3535 899 -3531
rect 898 -3552 899 -3534
rect 898 -3535 899 -3531
rect 898 -3552 899 -3534
rect 905 -3535 906 -3531
rect 905 -3552 906 -3534
rect 905 -3535 906 -3531
rect 905 -3552 906 -3534
rect 926 -3535 927 -3531
rect 950 -3535 951 -3531
rect 957 -3535 958 -3531
rect 968 -3535 969 -3531
rect 1038 -3535 1039 -3531
rect 1045 -3535 1046 -3531
rect 1052 -3535 1053 -3531
rect 1059 -3535 1060 -3531
rect 1073 -3535 1074 -3531
rect 1111 -3552 1112 -3534
rect 1143 -3535 1144 -3531
rect 1164 -3552 1165 -3534
rect 394 -3537 395 -3531
rect 401 -3552 402 -3536
rect 499 -3537 500 -3531
rect 513 -3552 514 -3536
rect 565 -3552 566 -3536
rect 576 -3537 577 -3531
rect 604 -3537 605 -3531
rect 607 -3552 608 -3536
rect 646 -3537 647 -3531
rect 663 -3552 664 -3536
rect 667 -3552 668 -3536
rect 765 -3537 766 -3531
rect 779 -3537 780 -3531
rect 800 -3552 801 -3536
rect 814 -3537 815 -3531
rect 814 -3552 815 -3536
rect 814 -3537 815 -3531
rect 814 -3552 815 -3536
rect 877 -3537 878 -3531
rect 884 -3552 885 -3536
rect 919 -3537 920 -3531
rect 926 -3552 927 -3536
rect 933 -3537 934 -3531
rect 936 -3552 937 -3536
rect 940 -3537 941 -3531
rect 940 -3552 941 -3536
rect 940 -3537 941 -3531
rect 940 -3552 941 -3536
rect 394 -3552 395 -3538
rect 492 -3539 493 -3531
rect 499 -3552 500 -3538
rect 569 -3539 570 -3531
rect 569 -3552 570 -3538
rect 569 -3539 570 -3531
rect 569 -3552 570 -3538
rect 576 -3552 577 -3538
rect 590 -3539 591 -3531
rect 702 -3552 703 -3538
rect 709 -3539 710 -3531
rect 772 -3539 773 -3531
rect 779 -3552 780 -3538
rect 793 -3539 794 -3531
rect 807 -3552 808 -3538
rect 863 -3539 864 -3531
rect 877 -3552 878 -3538
rect 485 -3541 486 -3531
rect 492 -3552 493 -3540
rect 590 -3552 591 -3540
rect 597 -3541 598 -3531
rect 772 -3552 773 -3540
rect 842 -3541 843 -3531
rect 583 -3543 584 -3531
rect 597 -3552 598 -3542
rect 555 -3545 556 -3531
rect 583 -3552 584 -3544
rect 541 -3547 542 -3531
rect 555 -3552 556 -3546
rect 534 -3549 535 -3531
rect 541 -3552 542 -3548
rect 534 -3552 535 -3550
rect 562 -3551 563 -3531
rect 387 -3562 388 -3560
rect 387 -3567 388 -3561
rect 387 -3562 388 -3560
rect 387 -3567 388 -3561
rect 394 -3562 395 -3560
rect 394 -3567 395 -3561
rect 394 -3562 395 -3560
rect 394 -3567 395 -3561
rect 401 -3562 402 -3560
rect 404 -3567 405 -3561
rect 408 -3562 409 -3560
rect 408 -3567 409 -3561
rect 408 -3562 409 -3560
rect 408 -3567 409 -3561
rect 457 -3562 458 -3560
rect 464 -3567 465 -3561
rect 474 -3562 475 -3560
rect 478 -3562 479 -3560
rect 492 -3562 493 -3560
rect 492 -3567 493 -3561
rect 492 -3562 493 -3560
rect 492 -3567 493 -3561
rect 499 -3567 500 -3561
rect 513 -3562 514 -3560
rect 527 -3562 528 -3560
rect 541 -3562 542 -3560
rect 555 -3562 556 -3560
rect 562 -3562 563 -3560
rect 569 -3562 570 -3560
rect 576 -3562 577 -3560
rect 579 -3562 580 -3560
rect 597 -3562 598 -3560
rect 632 -3567 633 -3561
rect 667 -3562 668 -3560
rect 702 -3562 703 -3560
rect 709 -3562 710 -3560
rect 737 -3562 738 -3560
rect 747 -3567 748 -3561
rect 758 -3562 759 -3560
rect 765 -3562 766 -3560
rect 768 -3562 769 -3560
rect 779 -3562 780 -3560
rect 786 -3562 787 -3560
rect 796 -3562 797 -3560
rect 800 -3562 801 -3560
rect 800 -3567 801 -3561
rect 800 -3562 801 -3560
rect 800 -3567 801 -3561
rect 877 -3562 878 -3560
rect 894 -3567 895 -3561
rect 901 -3567 902 -3561
rect 905 -3562 906 -3560
rect 926 -3562 927 -3560
rect 950 -3562 951 -3560
rect 1111 -3562 1112 -3560
rect 1115 -3562 1116 -3560
rect 1132 -3567 1133 -3561
rect 1136 -3562 1137 -3560
rect 1164 -3562 1165 -3560
rect 1171 -3567 1172 -3561
rect 1178 -3562 1179 -3560
rect 1185 -3567 1186 -3561
rect 1192 -3562 1193 -3560
rect 1199 -3567 1200 -3561
rect 1391 -3567 1392 -3561
rect 1395 -3562 1396 -3560
rect 380 -3564 381 -3560
rect 401 -3567 402 -3563
rect 450 -3564 451 -3560
rect 457 -3567 458 -3563
rect 502 -3564 503 -3560
rect 506 -3564 507 -3560
rect 530 -3564 531 -3560
rect 534 -3564 535 -3560
rect 548 -3564 549 -3560
rect 562 -3567 563 -3563
rect 576 -3567 577 -3563
rect 583 -3564 584 -3560
rect 590 -3564 591 -3560
rect 590 -3567 591 -3563
rect 590 -3564 591 -3560
rect 590 -3567 591 -3563
rect 758 -3567 759 -3563
rect 772 -3564 773 -3560
rect 793 -3564 794 -3560
rect 807 -3564 808 -3560
rect 884 -3564 885 -3560
rect 884 -3567 885 -3563
rect 884 -3564 885 -3560
rect 884 -3567 885 -3563
rect 891 -3567 892 -3563
rect 898 -3564 899 -3560
rect 933 -3564 934 -3560
rect 940 -3564 941 -3560
rect 1129 -3564 1130 -3560
rect 1136 -3567 1137 -3563
rect 1388 -3564 1389 -3560
rect 1395 -3567 1396 -3563
rect 807 -3567 808 -3565
rect 814 -3566 815 -3560
rect 1360 -3566 1361 -3560
rect 1388 -3567 1389 -3565
rect 387 -3577 388 -3575
rect 401 -3577 402 -3575
rect 457 -3577 458 -3575
rect 464 -3577 465 -3575
rect 492 -3577 493 -3575
rect 502 -3577 503 -3575
rect 562 -3577 563 -3575
rect 579 -3577 580 -3575
rect 590 -3577 591 -3575
rect 597 -3577 598 -3575
rect 600 -3577 601 -3575
rect 632 -3577 633 -3575
rect 747 -3577 748 -3575
rect 758 -3577 759 -3575
rect 800 -3577 801 -3575
rect 810 -3577 811 -3575
rect 884 -3577 885 -3575
rect 898 -3577 899 -3575
rect 1129 -3577 1130 -3575
rect 1136 -3577 1137 -3575
rect 1171 -3577 1172 -3575
rect 1181 -3577 1182 -3575
rect 1195 -3577 1196 -3575
rect 1199 -3577 1200 -3575
rect 1388 -3577 1389 -3575
rect 1395 -3577 1396 -3575
rect 397 -3579 398 -3575
rect 408 -3579 409 -3575
rect 1178 -3579 1179 -3575
rect 1185 -3579 1186 -3575
<< labels >>
rlabel pdiffusion 3 -18 3 -18 0 cellNo=156
rlabel pdiffusion 10 -18 10 -18 0 cellNo=520
rlabel pdiffusion 17 -18 17 -18 0 cellNo=1001
rlabel pdiffusion 24 -18 24 -18 0 cellNo=1003
rlabel pdiffusion 31 -18 31 -18 0 cellNo=1182
rlabel pdiffusion 38 -18 38 -18 0 cellNo=1011
rlabel pdiffusion 45 -18 45 -18 0 cellNo=1016
rlabel pdiffusion 52 -18 52 -18 0 cellNo=1155
rlabel pdiffusion 59 -18 59 -18 0 cellNo=1025
rlabel pdiffusion 66 -18 66 -18 0 cellNo=1026
rlabel pdiffusion 73 -18 73 -18 0 cellNo=1132
rlabel pdiffusion 80 -18 80 -18 0 cellNo=1050
rlabel pdiffusion 87 -18 87 -18 0 cellNo=1072
rlabel pdiffusion 94 -18 94 -18 0 cellNo=1046
rlabel pdiffusion 101 -18 101 -18 0 cellNo=1058
rlabel pdiffusion 108 -18 108 -18 0 cellNo=1064
rlabel pdiffusion 115 -18 115 -18 0 cellNo=1080
rlabel pdiffusion 122 -18 122 -18 0 cellNo=1082
rlabel pdiffusion 129 -18 129 -18 0 cellNo=1120
rlabel pdiffusion 136 -18 136 -18 0 cellNo=1145
rlabel pdiffusion 234 -18 234 -18 0 feedthrough
rlabel pdiffusion 346 -18 346 -18 0 feedthrough
rlabel pdiffusion 353 -18 353 -18 0 cellNo=140
rlabel pdiffusion 360 -18 360 -18 0 feedthrough
rlabel pdiffusion 381 -18 381 -18 0 feedthrough
rlabel pdiffusion 402 -18 402 -18 0 feedthrough
rlabel pdiffusion 409 -18 409 -18 0 feedthrough
rlabel pdiffusion 416 -18 416 -18 0 feedthrough
rlabel pdiffusion 423 -18 423 -18 0 feedthrough
rlabel pdiffusion 430 -18 430 -18 0 cellNo=765
rlabel pdiffusion 437 -18 437 -18 0 cellNo=266
rlabel pdiffusion 444 -18 444 -18 0 feedthrough
rlabel pdiffusion 451 -18 451 -18 0 cellNo=189
rlabel pdiffusion 458 -18 458 -18 0 cellNo=739
rlabel pdiffusion 465 -18 465 -18 0 cellNo=62
rlabel pdiffusion 472 -18 472 -18 0 feedthrough
rlabel pdiffusion 507 -18 507 -18 0 cellNo=928
rlabel pdiffusion 528 -18 528 -18 0 feedthrough
rlabel pdiffusion 535 -18 535 -18 0 cellNo=965
rlabel pdiffusion 549 -18 549 -18 0 cellNo=789
rlabel pdiffusion 556 -18 556 -18 0 feedthrough
rlabel pdiffusion 605 -18 605 -18 0 feedthrough
rlabel pdiffusion 612 -18 612 -18 0 cellNo=118
rlabel pdiffusion 654 -18 654 -18 0 feedthrough
rlabel pdiffusion 668 -18 668 -18 0 cellNo=106
rlabel pdiffusion 675 -18 675 -18 0 cellNo=407
rlabel pdiffusion 689 -18 689 -18 0 feedthrough
rlabel pdiffusion 717 -18 717 -18 0 cellNo=766
rlabel pdiffusion 752 -18 752 -18 0 cellNo=497
rlabel pdiffusion 801 -18 801 -18 0 feedthrough
rlabel pdiffusion 878 -18 878 -18 0 cellNo=545
rlabel pdiffusion 955 -18 955 -18 0 feedthrough
rlabel pdiffusion 3 -55 3 -55 0 cellNo=1004
rlabel pdiffusion 10 -55 10 -55 0 cellNo=1008
rlabel pdiffusion 17 -55 17 -55 0 cellNo=1100
rlabel pdiffusion 24 -55 24 -55 0 cellNo=1075
rlabel pdiffusion 31 -55 31 -55 0 cellNo=1010
rlabel pdiffusion 38 -55 38 -55 0 cellNo=1015
rlabel pdiffusion 45 -55 45 -55 0 cellNo=1039
rlabel pdiffusion 52 -55 52 -55 0 cellNo=1062
rlabel pdiffusion 59 -55 59 -55 0 cellNo=1083
rlabel pdiffusion 66 -55 66 -55 0 cellNo=1092
rlabel pdiffusion 73 -55 73 -55 0 cellNo=1104
rlabel pdiffusion 80 -55 80 -55 0 cellNo=1114
rlabel pdiffusion 87 -55 87 -55 0 cellNo=1115
rlabel pdiffusion 94 -55 94 -55 0 cellNo=1137
rlabel pdiffusion 143 -55 143 -55 0 cellNo=486
rlabel pdiffusion 150 -55 150 -55 0 feedthrough
rlabel pdiffusion 157 -55 157 -55 0 feedthrough
rlabel pdiffusion 227 -55 227 -55 0 feedthrough
rlabel pdiffusion 234 -55 234 -55 0 cellNo=895
rlabel pdiffusion 262 -55 262 -55 0 feedthrough
rlabel pdiffusion 283 -55 283 -55 0 feedthrough
rlabel pdiffusion 304 -55 304 -55 0 cellNo=334
rlabel pdiffusion 325 -55 325 -55 0 feedthrough
rlabel pdiffusion 332 -55 332 -55 0 feedthrough
rlabel pdiffusion 339 -55 339 -55 0 feedthrough
rlabel pdiffusion 374 -55 374 -55 0 feedthrough
rlabel pdiffusion 381 -55 381 -55 0 feedthrough
rlabel pdiffusion 388 -55 388 -55 0 cellNo=214
rlabel pdiffusion 395 -55 395 -55 0 feedthrough
rlabel pdiffusion 402 -55 402 -55 0 feedthrough
rlabel pdiffusion 409 -55 409 -55 0 cellNo=400
rlabel pdiffusion 416 -55 416 -55 0 cellNo=97
rlabel pdiffusion 423 -55 423 -55 0 cellNo=22
rlabel pdiffusion 430 -55 430 -55 0 feedthrough
rlabel pdiffusion 437 -55 437 -55 0 feedthrough
rlabel pdiffusion 444 -55 444 -55 0 cellNo=332
rlabel pdiffusion 451 -55 451 -55 0 feedthrough
rlabel pdiffusion 458 -55 458 -55 0 cellNo=788
rlabel pdiffusion 465 -55 465 -55 0 feedthrough
rlabel pdiffusion 472 -55 472 -55 0 feedthrough
rlabel pdiffusion 479 -55 479 -55 0 feedthrough
rlabel pdiffusion 493 -55 493 -55 0 cellNo=271
rlabel pdiffusion 500 -55 500 -55 0 feedthrough
rlabel pdiffusion 507 -55 507 -55 0 feedthrough
rlabel pdiffusion 514 -55 514 -55 0 cellNo=591
rlabel pdiffusion 521 -55 521 -55 0 cellNo=992
rlabel pdiffusion 528 -55 528 -55 0 cellNo=76
rlabel pdiffusion 535 -55 535 -55 0 feedthrough
rlabel pdiffusion 542 -55 542 -55 0 feedthrough
rlabel pdiffusion 549 -55 549 -55 0 feedthrough
rlabel pdiffusion 556 -55 556 -55 0 feedthrough
rlabel pdiffusion 563 -55 563 -55 0 feedthrough
rlabel pdiffusion 570 -55 570 -55 0 cellNo=164
rlabel pdiffusion 577 -55 577 -55 0 feedthrough
rlabel pdiffusion 584 -55 584 -55 0 feedthrough
rlabel pdiffusion 591 -55 591 -55 0 cellNo=762
rlabel pdiffusion 598 -55 598 -55 0 feedthrough
rlabel pdiffusion 605 -55 605 -55 0 feedthrough
rlabel pdiffusion 612 -55 612 -55 0 feedthrough
rlabel pdiffusion 619 -55 619 -55 0 feedthrough
rlabel pdiffusion 626 -55 626 -55 0 feedthrough
rlabel pdiffusion 633 -55 633 -55 0 cellNo=430
rlabel pdiffusion 640 -55 640 -55 0 feedthrough
rlabel pdiffusion 647 -55 647 -55 0 feedthrough
rlabel pdiffusion 654 -55 654 -55 0 feedthrough
rlabel pdiffusion 661 -55 661 -55 0 feedthrough
rlabel pdiffusion 668 -55 668 -55 0 feedthrough
rlabel pdiffusion 675 -55 675 -55 0 cellNo=616
rlabel pdiffusion 682 -55 682 -55 0 feedthrough
rlabel pdiffusion 689 -55 689 -55 0 feedthrough
rlabel pdiffusion 703 -55 703 -55 0 feedthrough
rlabel pdiffusion 710 -55 710 -55 0 cellNo=818
rlabel pdiffusion 717 -55 717 -55 0 feedthrough
rlabel pdiffusion 731 -55 731 -55 0 feedthrough
rlabel pdiffusion 745 -55 745 -55 0 feedthrough
rlabel pdiffusion 759 -55 759 -55 0 cellNo=255
rlabel pdiffusion 773 -55 773 -55 0 feedthrough
rlabel pdiffusion 815 -55 815 -55 0 feedthrough
rlabel pdiffusion 822 -55 822 -55 0 feedthrough
rlabel pdiffusion 829 -55 829 -55 0 feedthrough
rlabel pdiffusion 843 -55 843 -55 0 feedthrough
rlabel pdiffusion 885 -55 885 -55 0 cellNo=729
rlabel pdiffusion 899 -55 899 -55 0 feedthrough
rlabel pdiffusion 934 -55 934 -55 0 cellNo=339
rlabel pdiffusion 990 -55 990 -55 0 feedthrough
rlabel pdiffusion 997 -55 997 -55 0 feedthrough
rlabel pdiffusion 3 -102 3 -102 0 cellNo=443
rlabel pdiffusion 10 -102 10 -102 0 cellNo=1097
rlabel pdiffusion 17 -102 17 -102 0 cellNo=1107
rlabel pdiffusion 24 -102 24 -102 0 cellNo=1009
rlabel pdiffusion 31 -102 31 -102 0 cellNo=1068
rlabel pdiffusion 38 -102 38 -102 0 cellNo=1033
rlabel pdiffusion 45 -102 45 -102 0 cellNo=1074
rlabel pdiffusion 52 -102 52 -102 0 cellNo=1110
rlabel pdiffusion 59 -102 59 -102 0 cellNo=1049
rlabel pdiffusion 66 -102 66 -102 0 cellNo=1055
rlabel pdiffusion 73 -102 73 -102 0 cellNo=1061
rlabel pdiffusion 80 -102 80 -102 0 cellNo=1071
rlabel pdiffusion 87 -102 87 -102 0 cellNo=906
rlabel pdiffusion 94 -102 94 -102 0 cellNo=1069
rlabel pdiffusion 101 -102 101 -102 0 cellNo=590
rlabel pdiffusion 108 -102 108 -102 0 cellNo=1091
rlabel pdiffusion 129 -102 129 -102 0 feedthrough
rlabel pdiffusion 150 -102 150 -102 0 feedthrough
rlabel pdiffusion 192 -102 192 -102 0 feedthrough
rlabel pdiffusion 199 -102 199 -102 0 cellNo=751
rlabel pdiffusion 206 -102 206 -102 0 feedthrough
rlabel pdiffusion 220 -102 220 -102 0 feedthrough
rlabel pdiffusion 248 -102 248 -102 0 cellNo=637
rlabel pdiffusion 255 -102 255 -102 0 feedthrough
rlabel pdiffusion 262 -102 262 -102 0 feedthrough
rlabel pdiffusion 269 -102 269 -102 0 feedthrough
rlabel pdiffusion 276 -102 276 -102 0 feedthrough
rlabel pdiffusion 283 -102 283 -102 0 feedthrough
rlabel pdiffusion 290 -102 290 -102 0 cellNo=102
rlabel pdiffusion 297 -102 297 -102 0 feedthrough
rlabel pdiffusion 304 -102 304 -102 0 feedthrough
rlabel pdiffusion 311 -102 311 -102 0 feedthrough
rlabel pdiffusion 318 -102 318 -102 0 feedthrough
rlabel pdiffusion 325 -102 325 -102 0 feedthrough
rlabel pdiffusion 332 -102 332 -102 0 cellNo=795
rlabel pdiffusion 339 -102 339 -102 0 feedthrough
rlabel pdiffusion 346 -102 346 -102 0 feedthrough
rlabel pdiffusion 353 -102 353 -102 0 feedthrough
rlabel pdiffusion 360 -102 360 -102 0 feedthrough
rlabel pdiffusion 367 -102 367 -102 0 feedthrough
rlabel pdiffusion 374 -102 374 -102 0 cellNo=71
rlabel pdiffusion 381 -102 381 -102 0 feedthrough
rlabel pdiffusion 388 -102 388 -102 0 feedthrough
rlabel pdiffusion 395 -102 395 -102 0 feedthrough
rlabel pdiffusion 402 -102 402 -102 0 feedthrough
rlabel pdiffusion 409 -102 409 -102 0 cellNo=816
rlabel pdiffusion 416 -102 416 -102 0 feedthrough
rlabel pdiffusion 423 -102 423 -102 0 feedthrough
rlabel pdiffusion 430 -102 430 -102 0 cellNo=539
rlabel pdiffusion 437 -102 437 -102 0 feedthrough
rlabel pdiffusion 444 -102 444 -102 0 feedthrough
rlabel pdiffusion 451 -102 451 -102 0 feedthrough
rlabel pdiffusion 458 -102 458 -102 0 cellNo=634
rlabel pdiffusion 465 -102 465 -102 0 feedthrough
rlabel pdiffusion 472 -102 472 -102 0 cellNo=798
rlabel pdiffusion 479 -102 479 -102 0 feedthrough
rlabel pdiffusion 486 -102 486 -102 0 cellNo=428
rlabel pdiffusion 493 -102 493 -102 0 feedthrough
rlabel pdiffusion 500 -102 500 -102 0 feedthrough
rlabel pdiffusion 507 -102 507 -102 0 feedthrough
rlabel pdiffusion 514 -102 514 -102 0 feedthrough
rlabel pdiffusion 521 -102 521 -102 0 feedthrough
rlabel pdiffusion 528 -102 528 -102 0 cellNo=916
rlabel pdiffusion 535 -102 535 -102 0 cellNo=719
rlabel pdiffusion 542 -102 542 -102 0 feedthrough
rlabel pdiffusion 549 -102 549 -102 0 cellNo=537
rlabel pdiffusion 556 -102 556 -102 0 feedthrough
rlabel pdiffusion 563 -102 563 -102 0 feedthrough
rlabel pdiffusion 570 -102 570 -102 0 feedthrough
rlabel pdiffusion 577 -102 577 -102 0 feedthrough
rlabel pdiffusion 584 -102 584 -102 0 feedthrough
rlabel pdiffusion 591 -102 591 -102 0 feedthrough
rlabel pdiffusion 598 -102 598 -102 0 feedthrough
rlabel pdiffusion 605 -102 605 -102 0 feedthrough
rlabel pdiffusion 612 -102 612 -102 0 feedthrough
rlabel pdiffusion 619 -102 619 -102 0 feedthrough
rlabel pdiffusion 626 -102 626 -102 0 feedthrough
rlabel pdiffusion 633 -102 633 -102 0 feedthrough
rlabel pdiffusion 640 -102 640 -102 0 feedthrough
rlabel pdiffusion 647 -102 647 -102 0 cellNo=814
rlabel pdiffusion 654 -102 654 -102 0 feedthrough
rlabel pdiffusion 661 -102 661 -102 0 feedthrough
rlabel pdiffusion 668 -102 668 -102 0 feedthrough
rlabel pdiffusion 675 -102 675 -102 0 feedthrough
rlabel pdiffusion 682 -102 682 -102 0 feedthrough
rlabel pdiffusion 689 -102 689 -102 0 feedthrough
rlabel pdiffusion 696 -102 696 -102 0 feedthrough
rlabel pdiffusion 703 -102 703 -102 0 feedthrough
rlabel pdiffusion 710 -102 710 -102 0 feedthrough
rlabel pdiffusion 717 -102 717 -102 0 feedthrough
rlabel pdiffusion 724 -102 724 -102 0 feedthrough
rlabel pdiffusion 731 -102 731 -102 0 feedthrough
rlabel pdiffusion 738 -102 738 -102 0 feedthrough
rlabel pdiffusion 745 -102 745 -102 0 feedthrough
rlabel pdiffusion 752 -102 752 -102 0 feedthrough
rlabel pdiffusion 780 -102 780 -102 0 feedthrough
rlabel pdiffusion 787 -102 787 -102 0 feedthrough
rlabel pdiffusion 794 -102 794 -102 0 cellNo=778
rlabel pdiffusion 801 -102 801 -102 0 feedthrough
rlabel pdiffusion 808 -102 808 -102 0 cellNo=584
rlabel pdiffusion 815 -102 815 -102 0 cellNo=792
rlabel pdiffusion 822 -102 822 -102 0 cellNo=380
rlabel pdiffusion 829 -102 829 -102 0 feedthrough
rlabel pdiffusion 836 -102 836 -102 0 feedthrough
rlabel pdiffusion 843 -102 843 -102 0 feedthrough
rlabel pdiffusion 857 -102 857 -102 0 feedthrough
rlabel pdiffusion 864 -102 864 -102 0 feedthrough
rlabel pdiffusion 871 -102 871 -102 0 feedthrough
rlabel pdiffusion 885 -102 885 -102 0 cellNo=859
rlabel pdiffusion 892 -102 892 -102 0 feedthrough
rlabel pdiffusion 941 -102 941 -102 0 feedthrough
rlabel pdiffusion 948 -102 948 -102 0 feedthrough
rlabel pdiffusion 955 -102 955 -102 0 feedthrough
rlabel pdiffusion 1011 -102 1011 -102 0 feedthrough
rlabel pdiffusion 1088 -102 1088 -102 0 feedthrough
rlabel pdiffusion 3 -171 3 -171 0 cellNo=1002
rlabel pdiffusion 10 -171 10 -171 0 cellNo=1027
rlabel pdiffusion 17 -171 17 -171 0 cellNo=1007
rlabel pdiffusion 24 -171 24 -171 0 cellNo=1014
rlabel pdiffusion 31 -171 31 -171 0 cellNo=1084
rlabel pdiffusion 38 -171 38 -171 0 cellNo=1096
rlabel pdiffusion 45 -171 45 -171 0 cellNo=1190
rlabel pdiffusion 52 -171 52 -171 0 cellNo=1111
rlabel pdiffusion 59 -171 59 -171 0 cellNo=1081
rlabel pdiffusion 66 -171 66 -171 0 cellNo=1103
rlabel pdiffusion 73 -171 73 -171 0 cellNo=1186
rlabel pdiffusion 80 -171 80 -171 0 cellNo=1189
rlabel pdiffusion 94 -171 94 -171 0 feedthrough
rlabel pdiffusion 115 -171 115 -171 0 feedthrough
rlabel pdiffusion 136 -171 136 -171 0 feedthrough
rlabel pdiffusion 143 -171 143 -171 0 feedthrough
rlabel pdiffusion 150 -171 150 -171 0 feedthrough
rlabel pdiffusion 157 -171 157 -171 0 feedthrough
rlabel pdiffusion 164 -171 164 -171 0 feedthrough
rlabel pdiffusion 171 -171 171 -171 0 feedthrough
rlabel pdiffusion 178 -171 178 -171 0 feedthrough
rlabel pdiffusion 185 -171 185 -171 0 feedthrough
rlabel pdiffusion 192 -171 192 -171 0 feedthrough
rlabel pdiffusion 199 -171 199 -171 0 feedthrough
rlabel pdiffusion 206 -171 206 -171 0 cellNo=834
rlabel pdiffusion 213 -171 213 -171 0 cellNo=862
rlabel pdiffusion 220 -171 220 -171 0 feedthrough
rlabel pdiffusion 227 -171 227 -171 0 feedthrough
rlabel pdiffusion 234 -171 234 -171 0 cellNo=728
rlabel pdiffusion 241 -171 241 -171 0 cellNo=636
rlabel pdiffusion 248 -171 248 -171 0 feedthrough
rlabel pdiffusion 255 -171 255 -171 0 feedthrough
rlabel pdiffusion 262 -171 262 -171 0 feedthrough
rlabel pdiffusion 269 -171 269 -171 0 feedthrough
rlabel pdiffusion 276 -171 276 -171 0 feedthrough
rlabel pdiffusion 283 -171 283 -171 0 feedthrough
rlabel pdiffusion 290 -171 290 -171 0 feedthrough
rlabel pdiffusion 297 -171 297 -171 0 feedthrough
rlabel pdiffusion 304 -171 304 -171 0 feedthrough
rlabel pdiffusion 311 -171 311 -171 0 feedthrough
rlabel pdiffusion 318 -171 318 -171 0 feedthrough
rlabel pdiffusion 325 -171 325 -171 0 feedthrough
rlabel pdiffusion 332 -171 332 -171 0 feedthrough
rlabel pdiffusion 339 -171 339 -171 0 feedthrough
rlabel pdiffusion 346 -171 346 -171 0 feedthrough
rlabel pdiffusion 353 -171 353 -171 0 cellNo=870
rlabel pdiffusion 360 -171 360 -171 0 cellNo=882
rlabel pdiffusion 367 -171 367 -171 0 feedthrough
rlabel pdiffusion 374 -171 374 -171 0 feedthrough
rlabel pdiffusion 381 -171 381 -171 0 feedthrough
rlabel pdiffusion 388 -171 388 -171 0 feedthrough
rlabel pdiffusion 395 -171 395 -171 0 feedthrough
rlabel pdiffusion 402 -171 402 -171 0 feedthrough
rlabel pdiffusion 409 -171 409 -171 0 feedthrough
rlabel pdiffusion 416 -171 416 -171 0 feedthrough
rlabel pdiffusion 423 -171 423 -171 0 feedthrough
rlabel pdiffusion 430 -171 430 -171 0 cellNo=493
rlabel pdiffusion 437 -171 437 -171 0 feedthrough
rlabel pdiffusion 444 -171 444 -171 0 feedthrough
rlabel pdiffusion 451 -171 451 -171 0 feedthrough
rlabel pdiffusion 458 -171 458 -171 0 feedthrough
rlabel pdiffusion 465 -171 465 -171 0 cellNo=296
rlabel pdiffusion 472 -171 472 -171 0 feedthrough
rlabel pdiffusion 479 -171 479 -171 0 cellNo=447
rlabel pdiffusion 486 -171 486 -171 0 feedthrough
rlabel pdiffusion 493 -171 493 -171 0 feedthrough
rlabel pdiffusion 500 -171 500 -171 0 cellNo=586
rlabel pdiffusion 507 -171 507 -171 0 cellNo=448
rlabel pdiffusion 514 -171 514 -171 0 cellNo=487
rlabel pdiffusion 521 -171 521 -171 0 cellNo=472
rlabel pdiffusion 528 -171 528 -171 0 feedthrough
rlabel pdiffusion 535 -171 535 -171 0 feedthrough
rlabel pdiffusion 542 -171 542 -171 0 cellNo=694
rlabel pdiffusion 549 -171 549 -171 0 feedthrough
rlabel pdiffusion 556 -171 556 -171 0 feedthrough
rlabel pdiffusion 563 -171 563 -171 0 feedthrough
rlabel pdiffusion 570 -171 570 -171 0 feedthrough
rlabel pdiffusion 577 -171 577 -171 0 feedthrough
rlabel pdiffusion 584 -171 584 -171 0 feedthrough
rlabel pdiffusion 591 -171 591 -171 0 feedthrough
rlabel pdiffusion 598 -171 598 -171 0 feedthrough
rlabel pdiffusion 605 -171 605 -171 0 feedthrough
rlabel pdiffusion 612 -171 612 -171 0 cellNo=677
rlabel pdiffusion 619 -171 619 -171 0 feedthrough
rlabel pdiffusion 626 -171 626 -171 0 feedthrough
rlabel pdiffusion 633 -171 633 -171 0 feedthrough
rlabel pdiffusion 640 -171 640 -171 0 feedthrough
rlabel pdiffusion 647 -171 647 -171 0 feedthrough
rlabel pdiffusion 654 -171 654 -171 0 cellNo=283
rlabel pdiffusion 661 -171 661 -171 0 feedthrough
rlabel pdiffusion 668 -171 668 -171 0 feedthrough
rlabel pdiffusion 675 -171 675 -171 0 feedthrough
rlabel pdiffusion 682 -171 682 -171 0 feedthrough
rlabel pdiffusion 689 -171 689 -171 0 feedthrough
rlabel pdiffusion 696 -171 696 -171 0 cellNo=712
rlabel pdiffusion 703 -171 703 -171 0 feedthrough
rlabel pdiffusion 710 -171 710 -171 0 feedthrough
rlabel pdiffusion 717 -171 717 -171 0 feedthrough
rlabel pdiffusion 724 -171 724 -171 0 feedthrough
rlabel pdiffusion 731 -171 731 -171 0 feedthrough
rlabel pdiffusion 738 -171 738 -171 0 feedthrough
rlabel pdiffusion 745 -171 745 -171 0 feedthrough
rlabel pdiffusion 752 -171 752 -171 0 feedthrough
rlabel pdiffusion 759 -171 759 -171 0 feedthrough
rlabel pdiffusion 766 -171 766 -171 0 cellNo=721
rlabel pdiffusion 773 -171 773 -171 0 feedthrough
rlabel pdiffusion 780 -171 780 -171 0 feedthrough
rlabel pdiffusion 787 -171 787 -171 0 feedthrough
rlabel pdiffusion 794 -171 794 -171 0 cellNo=458
rlabel pdiffusion 801 -171 801 -171 0 feedthrough
rlabel pdiffusion 808 -171 808 -171 0 feedthrough
rlabel pdiffusion 815 -171 815 -171 0 feedthrough
rlabel pdiffusion 822 -171 822 -171 0 cellNo=833
rlabel pdiffusion 829 -171 829 -171 0 feedthrough
rlabel pdiffusion 836 -171 836 -171 0 feedthrough
rlabel pdiffusion 843 -171 843 -171 0 feedthrough
rlabel pdiffusion 850 -171 850 -171 0 feedthrough
rlabel pdiffusion 857 -171 857 -171 0 feedthrough
rlabel pdiffusion 864 -171 864 -171 0 feedthrough
rlabel pdiffusion 871 -171 871 -171 0 feedthrough
rlabel pdiffusion 878 -171 878 -171 0 cellNo=774
rlabel pdiffusion 885 -171 885 -171 0 cellNo=3
rlabel pdiffusion 892 -171 892 -171 0 feedthrough
rlabel pdiffusion 899 -171 899 -171 0 feedthrough
rlabel pdiffusion 906 -171 906 -171 0 feedthrough
rlabel pdiffusion 913 -171 913 -171 0 feedthrough
rlabel pdiffusion 920 -171 920 -171 0 feedthrough
rlabel pdiffusion 927 -171 927 -171 0 feedthrough
rlabel pdiffusion 934 -171 934 -171 0 feedthrough
rlabel pdiffusion 941 -171 941 -171 0 feedthrough
rlabel pdiffusion 948 -171 948 -171 0 feedthrough
rlabel pdiffusion 955 -171 955 -171 0 feedthrough
rlabel pdiffusion 962 -171 962 -171 0 feedthrough
rlabel pdiffusion 969 -171 969 -171 0 feedthrough
rlabel pdiffusion 976 -171 976 -171 0 feedthrough
rlabel pdiffusion 983 -171 983 -171 0 feedthrough
rlabel pdiffusion 997 -171 997 -171 0 feedthrough
rlabel pdiffusion 1011 -171 1011 -171 0 feedthrough
rlabel pdiffusion 1039 -171 1039 -171 0 feedthrough
rlabel pdiffusion 1130 -171 1130 -171 0 feedthrough
rlabel pdiffusion 1137 -171 1137 -171 0 feedthrough
rlabel pdiffusion 1193 -171 1193 -171 0 cellNo=360
rlabel pdiffusion 1221 -171 1221 -171 0 feedthrough
rlabel pdiffusion 3 -258 3 -258 0 cellNo=1006
rlabel pdiffusion 10 -258 10 -258 0 cellNo=1113
rlabel pdiffusion 17 -258 17 -258 0 cellNo=1147
rlabel pdiffusion 24 -258 24 -258 0 cellNo=1070
rlabel pdiffusion 31 -258 31 -258 0 cellNo=1102
rlabel pdiffusion 38 -258 38 -258 0 cellNo=1143
rlabel pdiffusion 52 -258 52 -258 0 feedthrough
rlabel pdiffusion 59 -258 59 -258 0 feedthrough
rlabel pdiffusion 66 -258 66 -258 0 feedthrough
rlabel pdiffusion 73 -258 73 -258 0 feedthrough
rlabel pdiffusion 80 -258 80 -258 0 feedthrough
rlabel pdiffusion 87 -258 87 -258 0 feedthrough
rlabel pdiffusion 94 -258 94 -258 0 feedthrough
rlabel pdiffusion 101 -258 101 -258 0 feedthrough
rlabel pdiffusion 108 -258 108 -258 0 feedthrough
rlabel pdiffusion 115 -258 115 -258 0 cellNo=611
rlabel pdiffusion 122 -258 122 -258 0 feedthrough
rlabel pdiffusion 129 -258 129 -258 0 feedthrough
rlabel pdiffusion 136 -258 136 -258 0 feedthrough
rlabel pdiffusion 143 -258 143 -258 0 feedthrough
rlabel pdiffusion 150 -258 150 -258 0 feedthrough
rlabel pdiffusion 157 -258 157 -258 0 feedthrough
rlabel pdiffusion 164 -258 164 -258 0 feedthrough
rlabel pdiffusion 171 -258 171 -258 0 cellNo=294
rlabel pdiffusion 178 -258 178 -258 0 feedthrough
rlabel pdiffusion 185 -258 185 -258 0 feedthrough
rlabel pdiffusion 192 -258 192 -258 0 cellNo=864
rlabel pdiffusion 199 -258 199 -258 0 cellNo=295
rlabel pdiffusion 206 -258 206 -258 0 feedthrough
rlabel pdiffusion 213 -258 213 -258 0 cellNo=381
rlabel pdiffusion 220 -258 220 -258 0 feedthrough
rlabel pdiffusion 227 -258 227 -258 0 feedthrough
rlabel pdiffusion 234 -258 234 -258 0 cellNo=503
rlabel pdiffusion 241 -258 241 -258 0 cellNo=995
rlabel pdiffusion 248 -258 248 -258 0 feedthrough
rlabel pdiffusion 255 -258 255 -258 0 feedthrough
rlabel pdiffusion 262 -258 262 -258 0 feedthrough
rlabel pdiffusion 269 -258 269 -258 0 feedthrough
rlabel pdiffusion 276 -258 276 -258 0 feedthrough
rlabel pdiffusion 283 -258 283 -258 0 feedthrough
rlabel pdiffusion 290 -258 290 -258 0 cellNo=142
rlabel pdiffusion 297 -258 297 -258 0 feedthrough
rlabel pdiffusion 304 -258 304 -258 0 feedthrough
rlabel pdiffusion 311 -258 311 -258 0 feedthrough
rlabel pdiffusion 318 -258 318 -258 0 feedthrough
rlabel pdiffusion 325 -258 325 -258 0 feedthrough
rlabel pdiffusion 332 -258 332 -258 0 feedthrough
rlabel pdiffusion 339 -258 339 -258 0 feedthrough
rlabel pdiffusion 346 -258 346 -258 0 feedthrough
rlabel pdiffusion 353 -258 353 -258 0 feedthrough
rlabel pdiffusion 360 -258 360 -258 0 feedthrough
rlabel pdiffusion 367 -258 367 -258 0 feedthrough
rlabel pdiffusion 374 -258 374 -258 0 feedthrough
rlabel pdiffusion 381 -258 381 -258 0 cellNo=348
rlabel pdiffusion 388 -258 388 -258 0 feedthrough
rlabel pdiffusion 395 -258 395 -258 0 feedthrough
rlabel pdiffusion 402 -258 402 -258 0 feedthrough
rlabel pdiffusion 409 -258 409 -258 0 feedthrough
rlabel pdiffusion 416 -258 416 -258 0 feedthrough
rlabel pdiffusion 423 -258 423 -258 0 feedthrough
rlabel pdiffusion 430 -258 430 -258 0 feedthrough
rlabel pdiffusion 437 -258 437 -258 0 feedthrough
rlabel pdiffusion 444 -258 444 -258 0 cellNo=515
rlabel pdiffusion 451 -258 451 -258 0 feedthrough
rlabel pdiffusion 458 -258 458 -258 0 cellNo=874
rlabel pdiffusion 465 -258 465 -258 0 cellNo=274
rlabel pdiffusion 472 -258 472 -258 0 cellNo=297
rlabel pdiffusion 479 -258 479 -258 0 feedthrough
rlabel pdiffusion 486 -258 486 -258 0 feedthrough
rlabel pdiffusion 493 -258 493 -258 0 cellNo=77
rlabel pdiffusion 500 -258 500 -258 0 feedthrough
rlabel pdiffusion 507 -258 507 -258 0 cellNo=642
rlabel pdiffusion 514 -258 514 -258 0 feedthrough
rlabel pdiffusion 521 -258 521 -258 0 feedthrough
rlabel pdiffusion 528 -258 528 -258 0 cellNo=413
rlabel pdiffusion 535 -258 535 -258 0 feedthrough
rlabel pdiffusion 542 -258 542 -258 0 cellNo=9
rlabel pdiffusion 549 -258 549 -258 0 feedthrough
rlabel pdiffusion 556 -258 556 -258 0 feedthrough
rlabel pdiffusion 563 -258 563 -258 0 feedthrough
rlabel pdiffusion 570 -258 570 -258 0 cellNo=596
rlabel pdiffusion 577 -258 577 -258 0 cellNo=849
rlabel pdiffusion 584 -258 584 -258 0 feedthrough
rlabel pdiffusion 591 -258 591 -258 0 cellNo=11
rlabel pdiffusion 598 -258 598 -258 0 feedthrough
rlabel pdiffusion 605 -258 605 -258 0 feedthrough
rlabel pdiffusion 612 -258 612 -258 0 cellNo=390
rlabel pdiffusion 619 -258 619 -258 0 feedthrough
rlabel pdiffusion 626 -258 626 -258 0 feedthrough
rlabel pdiffusion 633 -258 633 -258 0 feedthrough
rlabel pdiffusion 640 -258 640 -258 0 feedthrough
rlabel pdiffusion 647 -258 647 -258 0 feedthrough
rlabel pdiffusion 654 -258 654 -258 0 feedthrough
rlabel pdiffusion 661 -258 661 -258 0 feedthrough
rlabel pdiffusion 668 -258 668 -258 0 feedthrough
rlabel pdiffusion 675 -258 675 -258 0 feedthrough
rlabel pdiffusion 682 -258 682 -258 0 feedthrough
rlabel pdiffusion 689 -258 689 -258 0 feedthrough
rlabel pdiffusion 696 -258 696 -258 0 feedthrough
rlabel pdiffusion 703 -258 703 -258 0 feedthrough
rlabel pdiffusion 710 -258 710 -258 0 feedthrough
rlabel pdiffusion 717 -258 717 -258 0 cellNo=956
rlabel pdiffusion 724 -258 724 -258 0 feedthrough
rlabel pdiffusion 731 -258 731 -258 0 feedthrough
rlabel pdiffusion 738 -258 738 -258 0 feedthrough
rlabel pdiffusion 745 -258 745 -258 0 feedthrough
rlabel pdiffusion 752 -258 752 -258 0 feedthrough
rlabel pdiffusion 759 -258 759 -258 0 feedthrough
rlabel pdiffusion 766 -258 766 -258 0 feedthrough
rlabel pdiffusion 773 -258 773 -258 0 cellNo=475
rlabel pdiffusion 780 -258 780 -258 0 feedthrough
rlabel pdiffusion 787 -258 787 -258 0 cellNo=764
rlabel pdiffusion 794 -258 794 -258 0 feedthrough
rlabel pdiffusion 801 -258 801 -258 0 feedthrough
rlabel pdiffusion 808 -258 808 -258 0 feedthrough
rlabel pdiffusion 815 -258 815 -258 0 feedthrough
rlabel pdiffusion 822 -258 822 -258 0 feedthrough
rlabel pdiffusion 829 -258 829 -258 0 cellNo=953
rlabel pdiffusion 836 -258 836 -258 0 feedthrough
rlabel pdiffusion 843 -258 843 -258 0 feedthrough
rlabel pdiffusion 850 -258 850 -258 0 feedthrough
rlabel pdiffusion 857 -258 857 -258 0 feedthrough
rlabel pdiffusion 864 -258 864 -258 0 feedthrough
rlabel pdiffusion 871 -258 871 -258 0 feedthrough
rlabel pdiffusion 878 -258 878 -258 0 feedthrough
rlabel pdiffusion 885 -258 885 -258 0 feedthrough
rlabel pdiffusion 892 -258 892 -258 0 feedthrough
rlabel pdiffusion 899 -258 899 -258 0 feedthrough
rlabel pdiffusion 906 -258 906 -258 0 feedthrough
rlabel pdiffusion 913 -258 913 -258 0 feedthrough
rlabel pdiffusion 920 -258 920 -258 0 feedthrough
rlabel pdiffusion 927 -258 927 -258 0 feedthrough
rlabel pdiffusion 934 -258 934 -258 0 feedthrough
rlabel pdiffusion 941 -258 941 -258 0 feedthrough
rlabel pdiffusion 948 -258 948 -258 0 feedthrough
rlabel pdiffusion 955 -258 955 -258 0 feedthrough
rlabel pdiffusion 962 -258 962 -258 0 feedthrough
rlabel pdiffusion 969 -258 969 -258 0 feedthrough
rlabel pdiffusion 976 -258 976 -258 0 feedthrough
rlabel pdiffusion 983 -258 983 -258 0 feedthrough
rlabel pdiffusion 990 -258 990 -258 0 feedthrough
rlabel pdiffusion 997 -258 997 -258 0 cellNo=710
rlabel pdiffusion 1004 -258 1004 -258 0 feedthrough
rlabel pdiffusion 1011 -258 1011 -258 0 feedthrough
rlabel pdiffusion 1018 -258 1018 -258 0 feedthrough
rlabel pdiffusion 1025 -258 1025 -258 0 feedthrough
rlabel pdiffusion 1032 -258 1032 -258 0 feedthrough
rlabel pdiffusion 1039 -258 1039 -258 0 feedthrough
rlabel pdiffusion 1046 -258 1046 -258 0 feedthrough
rlabel pdiffusion 1053 -258 1053 -258 0 feedthrough
rlabel pdiffusion 1060 -258 1060 -258 0 feedthrough
rlabel pdiffusion 1067 -258 1067 -258 0 feedthrough
rlabel pdiffusion 1074 -258 1074 -258 0 feedthrough
rlabel pdiffusion 1081 -258 1081 -258 0 feedthrough
rlabel pdiffusion 1088 -258 1088 -258 0 feedthrough
rlabel pdiffusion 1095 -258 1095 -258 0 cellNo=341
rlabel pdiffusion 1102 -258 1102 -258 0 feedthrough
rlabel pdiffusion 1109 -258 1109 -258 0 feedthrough
rlabel pdiffusion 1116 -258 1116 -258 0 cellNo=280
rlabel pdiffusion 1123 -258 1123 -258 0 cellNo=439
rlabel pdiffusion 1130 -258 1130 -258 0 feedthrough
rlabel pdiffusion 1137 -258 1137 -258 0 feedthrough
rlabel pdiffusion 1144 -258 1144 -258 0 feedthrough
rlabel pdiffusion 1151 -258 1151 -258 0 feedthrough
rlabel pdiffusion 1158 -258 1158 -258 0 feedthrough
rlabel pdiffusion 1165 -258 1165 -258 0 feedthrough
rlabel pdiffusion 1172 -258 1172 -258 0 feedthrough
rlabel pdiffusion 1228 -258 1228 -258 0 feedthrough
rlabel pdiffusion 1256 -258 1256 -258 0 feedthrough
rlabel pdiffusion 1284 -258 1284 -258 0 feedthrough
rlabel pdiffusion 3 -389 3 -389 0 cellNo=1005
rlabel pdiffusion 10 -389 10 -389 0 cellNo=1013
rlabel pdiffusion 17 -389 17 -389 0 cellNo=1022
rlabel pdiffusion 24 -389 24 -389 0 cellNo=1065
rlabel pdiffusion 31 -389 31 -389 0 cellNo=1020
rlabel pdiffusion 38 -389 38 -389 0 cellNo=1021
rlabel pdiffusion 45 -389 45 -389 0 feedthrough
rlabel pdiffusion 52 -389 52 -389 0 feedthrough
rlabel pdiffusion 59 -389 59 -389 0 cellNo=317
rlabel pdiffusion 66 -389 66 -389 0 feedthrough
rlabel pdiffusion 73 -389 73 -389 0 feedthrough
rlabel pdiffusion 80 -389 80 -389 0 feedthrough
rlabel pdiffusion 87 -389 87 -389 0 feedthrough
rlabel pdiffusion 94 -389 94 -389 0 cellNo=374
rlabel pdiffusion 101 -389 101 -389 0 feedthrough
rlabel pdiffusion 108 -389 108 -389 0 feedthrough
rlabel pdiffusion 115 -389 115 -389 0 cellNo=27
rlabel pdiffusion 122 -389 122 -389 0 cellNo=33
rlabel pdiffusion 129 -389 129 -389 0 feedthrough
rlabel pdiffusion 136 -389 136 -389 0 cellNo=362
rlabel pdiffusion 143 -389 143 -389 0 feedthrough
rlabel pdiffusion 150 -389 150 -389 0 feedthrough
rlabel pdiffusion 157 -389 157 -389 0 feedthrough
rlabel pdiffusion 164 -389 164 -389 0 feedthrough
rlabel pdiffusion 171 -389 171 -389 0 feedthrough
rlabel pdiffusion 178 -389 178 -389 0 feedthrough
rlabel pdiffusion 185 -389 185 -389 0 feedthrough
rlabel pdiffusion 192 -389 192 -389 0 feedthrough
rlabel pdiffusion 199 -389 199 -389 0 cellNo=505
rlabel pdiffusion 206 -389 206 -389 0 cellNo=826
rlabel pdiffusion 213 -389 213 -389 0 cellNo=499
rlabel pdiffusion 220 -389 220 -389 0 feedthrough
rlabel pdiffusion 227 -389 227 -389 0 feedthrough
rlabel pdiffusion 234 -389 234 -389 0 cellNo=1136
rlabel pdiffusion 241 -389 241 -389 0 feedthrough
rlabel pdiffusion 248 -389 248 -389 0 cellNo=1117
rlabel pdiffusion 255 -389 255 -389 0 feedthrough
rlabel pdiffusion 262 -389 262 -389 0 feedthrough
rlabel pdiffusion 269 -389 269 -389 0 feedthrough
rlabel pdiffusion 276 -389 276 -389 0 feedthrough
rlabel pdiffusion 283 -389 283 -389 0 cellNo=410
rlabel pdiffusion 290 -389 290 -389 0 feedthrough
rlabel pdiffusion 297 -389 297 -389 0 feedthrough
rlabel pdiffusion 304 -389 304 -389 0 feedthrough
rlabel pdiffusion 311 -389 311 -389 0 feedthrough
rlabel pdiffusion 318 -389 318 -389 0 cellNo=151
rlabel pdiffusion 325 -389 325 -389 0 feedthrough
rlabel pdiffusion 332 -389 332 -389 0 feedthrough
rlabel pdiffusion 339 -389 339 -389 0 cellNo=516
rlabel pdiffusion 346 -389 346 -389 0 feedthrough
rlabel pdiffusion 353 -389 353 -389 0 feedthrough
rlabel pdiffusion 360 -389 360 -389 0 feedthrough
rlabel pdiffusion 367 -389 367 -389 0 feedthrough
rlabel pdiffusion 374 -389 374 -389 0 feedthrough
rlabel pdiffusion 381 -389 381 -389 0 feedthrough
rlabel pdiffusion 388 -389 388 -389 0 feedthrough
rlabel pdiffusion 395 -389 395 -389 0 feedthrough
rlabel pdiffusion 402 -389 402 -389 0 feedthrough
rlabel pdiffusion 409 -389 409 -389 0 cellNo=158
rlabel pdiffusion 416 -389 416 -389 0 feedthrough
rlabel pdiffusion 423 -389 423 -389 0 feedthrough
rlabel pdiffusion 430 -389 430 -389 0 feedthrough
rlabel pdiffusion 437 -389 437 -389 0 cellNo=583
rlabel pdiffusion 444 -389 444 -389 0 feedthrough
rlabel pdiffusion 451 -389 451 -389 0 cellNo=686
rlabel pdiffusion 458 -389 458 -389 0 feedthrough
rlabel pdiffusion 465 -389 465 -389 0 feedthrough
rlabel pdiffusion 472 -389 472 -389 0 cellNo=455
rlabel pdiffusion 479 -389 479 -389 0 feedthrough
rlabel pdiffusion 486 -389 486 -389 0 feedthrough
rlabel pdiffusion 493 -389 493 -389 0 feedthrough
rlabel pdiffusion 500 -389 500 -389 0 feedthrough
rlabel pdiffusion 507 -389 507 -389 0 cellNo=848
rlabel pdiffusion 514 -389 514 -389 0 feedthrough
rlabel pdiffusion 521 -389 521 -389 0 feedthrough
rlabel pdiffusion 528 -389 528 -389 0 feedthrough
rlabel pdiffusion 535 -389 535 -389 0 feedthrough
rlabel pdiffusion 542 -389 542 -389 0 feedthrough
rlabel pdiffusion 549 -389 549 -389 0 feedthrough
rlabel pdiffusion 556 -389 556 -389 0 feedthrough
rlabel pdiffusion 563 -389 563 -389 0 feedthrough
rlabel pdiffusion 570 -389 570 -389 0 cellNo=7
rlabel pdiffusion 577 -389 577 -389 0 feedthrough
rlabel pdiffusion 584 -389 584 -389 0 feedthrough
rlabel pdiffusion 591 -389 591 -389 0 feedthrough
rlabel pdiffusion 598 -389 598 -389 0 feedthrough
rlabel pdiffusion 605 -389 605 -389 0 cellNo=408
rlabel pdiffusion 612 -389 612 -389 0 cellNo=577
rlabel pdiffusion 619 -389 619 -389 0 feedthrough
rlabel pdiffusion 626 -389 626 -389 0 feedthrough
rlabel pdiffusion 633 -389 633 -389 0 feedthrough
rlabel pdiffusion 640 -389 640 -389 0 feedthrough
rlabel pdiffusion 647 -389 647 -389 0 feedthrough
rlabel pdiffusion 654 -389 654 -389 0 feedthrough
rlabel pdiffusion 661 -389 661 -389 0 feedthrough
rlabel pdiffusion 668 -389 668 -389 0 cellNo=359
rlabel pdiffusion 675 -389 675 -389 0 feedthrough
rlabel pdiffusion 682 -389 682 -389 0 feedthrough
rlabel pdiffusion 689 -389 689 -389 0 feedthrough
rlabel pdiffusion 696 -389 696 -389 0 feedthrough
rlabel pdiffusion 703 -389 703 -389 0 cellNo=43
rlabel pdiffusion 710 -389 710 -389 0 cellNo=330
rlabel pdiffusion 717 -389 717 -389 0 feedthrough
rlabel pdiffusion 724 -389 724 -389 0 feedthrough
rlabel pdiffusion 731 -389 731 -389 0 cellNo=681
rlabel pdiffusion 738 -389 738 -389 0 feedthrough
rlabel pdiffusion 745 -389 745 -389 0 cellNo=215
rlabel pdiffusion 752 -389 752 -389 0 cellNo=624
rlabel pdiffusion 759 -389 759 -389 0 feedthrough
rlabel pdiffusion 766 -389 766 -389 0 feedthrough
rlabel pdiffusion 773 -389 773 -389 0 feedthrough
rlabel pdiffusion 780 -389 780 -389 0 feedthrough
rlabel pdiffusion 787 -389 787 -389 0 feedthrough
rlabel pdiffusion 794 -389 794 -389 0 feedthrough
rlabel pdiffusion 801 -389 801 -389 0 feedthrough
rlabel pdiffusion 808 -389 808 -389 0 feedthrough
rlabel pdiffusion 815 -389 815 -389 0 feedthrough
rlabel pdiffusion 822 -389 822 -389 0 feedthrough
rlabel pdiffusion 829 -389 829 -389 0 feedthrough
rlabel pdiffusion 836 -389 836 -389 0 feedthrough
rlabel pdiffusion 843 -389 843 -389 0 feedthrough
rlabel pdiffusion 850 -389 850 -389 0 feedthrough
rlabel pdiffusion 857 -389 857 -389 0 feedthrough
rlabel pdiffusion 864 -389 864 -389 0 feedthrough
rlabel pdiffusion 871 -389 871 -389 0 feedthrough
rlabel pdiffusion 878 -389 878 -389 0 feedthrough
rlabel pdiffusion 885 -389 885 -389 0 feedthrough
rlabel pdiffusion 892 -389 892 -389 0 feedthrough
rlabel pdiffusion 899 -389 899 -389 0 feedthrough
rlabel pdiffusion 906 -389 906 -389 0 feedthrough
rlabel pdiffusion 913 -389 913 -389 0 feedthrough
rlabel pdiffusion 920 -389 920 -389 0 feedthrough
rlabel pdiffusion 927 -389 927 -389 0 feedthrough
rlabel pdiffusion 934 -389 934 -389 0 feedthrough
rlabel pdiffusion 941 -389 941 -389 0 feedthrough
rlabel pdiffusion 948 -389 948 -389 0 feedthrough
rlabel pdiffusion 955 -389 955 -389 0 feedthrough
rlabel pdiffusion 962 -389 962 -389 0 feedthrough
rlabel pdiffusion 969 -389 969 -389 0 feedthrough
rlabel pdiffusion 976 -389 976 -389 0 feedthrough
rlabel pdiffusion 983 -389 983 -389 0 feedthrough
rlabel pdiffusion 990 -389 990 -389 0 feedthrough
rlabel pdiffusion 997 -389 997 -389 0 feedthrough
rlabel pdiffusion 1004 -389 1004 -389 0 feedthrough
rlabel pdiffusion 1011 -389 1011 -389 0 feedthrough
rlabel pdiffusion 1018 -389 1018 -389 0 feedthrough
rlabel pdiffusion 1025 -389 1025 -389 0 feedthrough
rlabel pdiffusion 1032 -389 1032 -389 0 feedthrough
rlabel pdiffusion 1039 -389 1039 -389 0 feedthrough
rlabel pdiffusion 1046 -389 1046 -389 0 feedthrough
rlabel pdiffusion 1053 -389 1053 -389 0 feedthrough
rlabel pdiffusion 1060 -389 1060 -389 0 feedthrough
rlabel pdiffusion 1067 -389 1067 -389 0 feedthrough
rlabel pdiffusion 1074 -389 1074 -389 0 feedthrough
rlabel pdiffusion 1081 -389 1081 -389 0 feedthrough
rlabel pdiffusion 1088 -389 1088 -389 0 feedthrough
rlabel pdiffusion 1095 -389 1095 -389 0 feedthrough
rlabel pdiffusion 1102 -389 1102 -389 0 feedthrough
rlabel pdiffusion 1109 -389 1109 -389 0 feedthrough
rlabel pdiffusion 1116 -389 1116 -389 0 feedthrough
rlabel pdiffusion 1123 -389 1123 -389 0 feedthrough
rlabel pdiffusion 1130 -389 1130 -389 0 feedthrough
rlabel pdiffusion 1137 -389 1137 -389 0 feedthrough
rlabel pdiffusion 1144 -389 1144 -389 0 feedthrough
rlabel pdiffusion 1151 -389 1151 -389 0 feedthrough
rlabel pdiffusion 1158 -389 1158 -389 0 feedthrough
rlabel pdiffusion 1165 -389 1165 -389 0 feedthrough
rlabel pdiffusion 1172 -389 1172 -389 0 feedthrough
rlabel pdiffusion 1179 -389 1179 -389 0 feedthrough
rlabel pdiffusion 1186 -389 1186 -389 0 feedthrough
rlabel pdiffusion 1193 -389 1193 -389 0 feedthrough
rlabel pdiffusion 1200 -389 1200 -389 0 cellNo=771
rlabel pdiffusion 1207 -389 1207 -389 0 feedthrough
rlabel pdiffusion 1214 -389 1214 -389 0 feedthrough
rlabel pdiffusion 1221 -389 1221 -389 0 feedthrough
rlabel pdiffusion 1228 -389 1228 -389 0 feedthrough
rlabel pdiffusion 1235 -389 1235 -389 0 feedthrough
rlabel pdiffusion 1242 -389 1242 -389 0 feedthrough
rlabel pdiffusion 1249 -389 1249 -389 0 feedthrough
rlabel pdiffusion 1256 -389 1256 -389 0 feedthrough
rlabel pdiffusion 1263 -389 1263 -389 0 feedthrough
rlabel pdiffusion 1270 -389 1270 -389 0 feedthrough
rlabel pdiffusion 1277 -389 1277 -389 0 feedthrough
rlabel pdiffusion 1284 -389 1284 -389 0 feedthrough
rlabel pdiffusion 1291 -389 1291 -389 0 feedthrough
rlabel pdiffusion 1298 -389 1298 -389 0 feedthrough
rlabel pdiffusion 1305 -389 1305 -389 0 feedthrough
rlabel pdiffusion 1312 -389 1312 -389 0 feedthrough
rlabel pdiffusion 1319 -389 1319 -389 0 feedthrough
rlabel pdiffusion 1326 -389 1326 -389 0 feedthrough
rlabel pdiffusion 1333 -389 1333 -389 0 feedthrough
rlabel pdiffusion 1340 -389 1340 -389 0 feedthrough
rlabel pdiffusion 1347 -389 1347 -389 0 feedthrough
rlabel pdiffusion 1354 -389 1354 -389 0 feedthrough
rlabel pdiffusion 1361 -389 1361 -389 0 feedthrough
rlabel pdiffusion 1368 -389 1368 -389 0 feedthrough
rlabel pdiffusion 1375 -389 1375 -389 0 feedthrough
rlabel pdiffusion 1382 -389 1382 -389 0 feedthrough
rlabel pdiffusion 1389 -389 1389 -389 0 feedthrough
rlabel pdiffusion 1396 -389 1396 -389 0 cellNo=357
rlabel pdiffusion 1592 -389 1592 -389 0 feedthrough
rlabel pdiffusion 3 -500 3 -500 0 cellNo=1012
rlabel pdiffusion 10 -500 10 -500 0 cellNo=1018
rlabel pdiffusion 17 -500 17 -500 0 cellNo=1142
rlabel pdiffusion 24 -500 24 -500 0 cellNo=846
rlabel pdiffusion 31 -500 31 -500 0 feedthrough
rlabel pdiffusion 38 -500 38 -500 0 feedthrough
rlabel pdiffusion 45 -500 45 -500 0 feedthrough
rlabel pdiffusion 52 -500 52 -500 0 feedthrough
rlabel pdiffusion 59 -500 59 -500 0 feedthrough
rlabel pdiffusion 66 -500 66 -500 0 feedthrough
rlabel pdiffusion 73 -500 73 -500 0 feedthrough
rlabel pdiffusion 80 -500 80 -500 0 cellNo=90
rlabel pdiffusion 87 -500 87 -500 0 cellNo=168
rlabel pdiffusion 94 -500 94 -500 0 feedthrough
rlabel pdiffusion 101 -500 101 -500 0 cellNo=172
rlabel pdiffusion 108 -500 108 -500 0 cellNo=141
rlabel pdiffusion 115 -500 115 -500 0 feedthrough
rlabel pdiffusion 122 -500 122 -500 0 feedthrough
rlabel pdiffusion 129 -500 129 -500 0 feedthrough
rlabel pdiffusion 136 -500 136 -500 0 cellNo=800
rlabel pdiffusion 143 -500 143 -500 0 feedthrough
rlabel pdiffusion 150 -500 150 -500 0 feedthrough
rlabel pdiffusion 157 -500 157 -500 0 feedthrough
rlabel pdiffusion 164 -500 164 -500 0 feedthrough
rlabel pdiffusion 171 -500 171 -500 0 feedthrough
rlabel pdiffusion 178 -500 178 -500 0 cellNo=512
rlabel pdiffusion 185 -500 185 -500 0 cellNo=411
rlabel pdiffusion 192 -500 192 -500 0 cellNo=602
rlabel pdiffusion 199 -500 199 -500 0 feedthrough
rlabel pdiffusion 206 -500 206 -500 0 feedthrough
rlabel pdiffusion 213 -500 213 -500 0 feedthrough
rlabel pdiffusion 220 -500 220 -500 0 cellNo=632
rlabel pdiffusion 227 -500 227 -500 0 feedthrough
rlabel pdiffusion 234 -500 234 -500 0 feedthrough
rlabel pdiffusion 241 -500 241 -500 0 feedthrough
rlabel pdiffusion 248 -500 248 -500 0 feedthrough
rlabel pdiffusion 255 -500 255 -500 0 feedthrough
rlabel pdiffusion 262 -500 262 -500 0 feedthrough
rlabel pdiffusion 269 -500 269 -500 0 feedthrough
rlabel pdiffusion 276 -500 276 -500 0 feedthrough
rlabel pdiffusion 283 -500 283 -500 0 feedthrough
rlabel pdiffusion 290 -500 290 -500 0 feedthrough
rlabel pdiffusion 297 -500 297 -500 0 cellNo=618
rlabel pdiffusion 304 -500 304 -500 0 feedthrough
rlabel pdiffusion 311 -500 311 -500 0 feedthrough
rlabel pdiffusion 318 -500 318 -500 0 feedthrough
rlabel pdiffusion 325 -500 325 -500 0 feedthrough
rlabel pdiffusion 332 -500 332 -500 0 feedthrough
rlabel pdiffusion 339 -500 339 -500 0 feedthrough
rlabel pdiffusion 346 -500 346 -500 0 feedthrough
rlabel pdiffusion 353 -500 353 -500 0 feedthrough
rlabel pdiffusion 360 -500 360 -500 0 cellNo=112
rlabel pdiffusion 367 -500 367 -500 0 feedthrough
rlabel pdiffusion 374 -500 374 -500 0 feedthrough
rlabel pdiffusion 381 -500 381 -500 0 feedthrough
rlabel pdiffusion 388 -500 388 -500 0 feedthrough
rlabel pdiffusion 395 -500 395 -500 0 feedthrough
rlabel pdiffusion 402 -500 402 -500 0 feedthrough
rlabel pdiffusion 409 -500 409 -500 0 feedthrough
rlabel pdiffusion 416 -500 416 -500 0 cellNo=24
rlabel pdiffusion 423 -500 423 -500 0 feedthrough
rlabel pdiffusion 430 -500 430 -500 0 feedthrough
rlabel pdiffusion 437 -500 437 -500 0 feedthrough
rlabel pdiffusion 444 -500 444 -500 0 feedthrough
rlabel pdiffusion 451 -500 451 -500 0 cellNo=405
rlabel pdiffusion 458 -500 458 -500 0 feedthrough
rlabel pdiffusion 465 -500 465 -500 0 feedthrough
rlabel pdiffusion 472 -500 472 -500 0 cellNo=894
rlabel pdiffusion 479 -500 479 -500 0 cellNo=37
rlabel pdiffusion 486 -500 486 -500 0 feedthrough
rlabel pdiffusion 493 -500 493 -500 0 cellNo=191
rlabel pdiffusion 500 -500 500 -500 0 feedthrough
rlabel pdiffusion 507 -500 507 -500 0 feedthrough
rlabel pdiffusion 514 -500 514 -500 0 cellNo=883
rlabel pdiffusion 521 -500 521 -500 0 cellNo=179
rlabel pdiffusion 528 -500 528 -500 0 cellNo=639
rlabel pdiffusion 535 -500 535 -500 0 cellNo=840
rlabel pdiffusion 542 -500 542 -500 0 feedthrough
rlabel pdiffusion 549 -500 549 -500 0 feedthrough
rlabel pdiffusion 556 -500 556 -500 0 feedthrough
rlabel pdiffusion 563 -500 563 -500 0 feedthrough
rlabel pdiffusion 570 -500 570 -500 0 feedthrough
rlabel pdiffusion 577 -500 577 -500 0 feedthrough
rlabel pdiffusion 584 -500 584 -500 0 feedthrough
rlabel pdiffusion 591 -500 591 -500 0 cellNo=672
rlabel pdiffusion 598 -500 598 -500 0 cellNo=206
rlabel pdiffusion 605 -500 605 -500 0 feedthrough
rlabel pdiffusion 612 -500 612 -500 0 feedthrough
rlabel pdiffusion 619 -500 619 -500 0 feedthrough
rlabel pdiffusion 626 -500 626 -500 0 feedthrough
rlabel pdiffusion 633 -500 633 -500 0 cellNo=452
rlabel pdiffusion 640 -500 640 -500 0 feedthrough
rlabel pdiffusion 647 -500 647 -500 0 cellNo=133
rlabel pdiffusion 654 -500 654 -500 0 feedthrough
rlabel pdiffusion 661 -500 661 -500 0 feedthrough
rlabel pdiffusion 668 -500 668 -500 0 feedthrough
rlabel pdiffusion 675 -500 675 -500 0 feedthrough
rlabel pdiffusion 682 -500 682 -500 0 feedthrough
rlabel pdiffusion 689 -500 689 -500 0 feedthrough
rlabel pdiffusion 696 -500 696 -500 0 cellNo=370
rlabel pdiffusion 703 -500 703 -500 0 feedthrough
rlabel pdiffusion 710 -500 710 -500 0 cellNo=291
rlabel pdiffusion 717 -500 717 -500 0 feedthrough
rlabel pdiffusion 724 -500 724 -500 0 feedthrough
rlabel pdiffusion 731 -500 731 -500 0 feedthrough
rlabel pdiffusion 738 -500 738 -500 0 feedthrough
rlabel pdiffusion 745 -500 745 -500 0 feedthrough
rlabel pdiffusion 752 -500 752 -500 0 feedthrough
rlabel pdiffusion 759 -500 759 -500 0 cellNo=527
rlabel pdiffusion 766 -500 766 -500 0 feedthrough
rlabel pdiffusion 773 -500 773 -500 0 feedthrough
rlabel pdiffusion 780 -500 780 -500 0 feedthrough
rlabel pdiffusion 787 -500 787 -500 0 feedthrough
rlabel pdiffusion 794 -500 794 -500 0 feedthrough
rlabel pdiffusion 801 -500 801 -500 0 feedthrough
rlabel pdiffusion 808 -500 808 -500 0 feedthrough
rlabel pdiffusion 815 -500 815 -500 0 feedthrough
rlabel pdiffusion 822 -500 822 -500 0 feedthrough
rlabel pdiffusion 829 -500 829 -500 0 cellNo=533
rlabel pdiffusion 836 -500 836 -500 0 feedthrough
rlabel pdiffusion 843 -500 843 -500 0 feedthrough
rlabel pdiffusion 850 -500 850 -500 0 feedthrough
rlabel pdiffusion 857 -500 857 -500 0 feedthrough
rlabel pdiffusion 864 -500 864 -500 0 feedthrough
rlabel pdiffusion 871 -500 871 -500 0 feedthrough
rlabel pdiffusion 878 -500 878 -500 0 feedthrough
rlabel pdiffusion 885 -500 885 -500 0 feedthrough
rlabel pdiffusion 892 -500 892 -500 0 feedthrough
rlabel pdiffusion 899 -500 899 -500 0 cellNo=892
rlabel pdiffusion 906 -500 906 -500 0 feedthrough
rlabel pdiffusion 913 -500 913 -500 0 feedthrough
rlabel pdiffusion 920 -500 920 -500 0 feedthrough
rlabel pdiffusion 927 -500 927 -500 0 feedthrough
rlabel pdiffusion 934 -500 934 -500 0 feedthrough
rlabel pdiffusion 941 -500 941 -500 0 feedthrough
rlabel pdiffusion 948 -500 948 -500 0 feedthrough
rlabel pdiffusion 955 -500 955 -500 0 feedthrough
rlabel pdiffusion 962 -500 962 -500 0 feedthrough
rlabel pdiffusion 969 -500 969 -500 0 feedthrough
rlabel pdiffusion 976 -500 976 -500 0 feedthrough
rlabel pdiffusion 983 -500 983 -500 0 feedthrough
rlabel pdiffusion 990 -500 990 -500 0 feedthrough
rlabel pdiffusion 997 -500 997 -500 0 feedthrough
rlabel pdiffusion 1004 -500 1004 -500 0 feedthrough
rlabel pdiffusion 1011 -500 1011 -500 0 feedthrough
rlabel pdiffusion 1018 -500 1018 -500 0 feedthrough
rlabel pdiffusion 1025 -500 1025 -500 0 feedthrough
rlabel pdiffusion 1032 -500 1032 -500 0 feedthrough
rlabel pdiffusion 1039 -500 1039 -500 0 feedthrough
rlabel pdiffusion 1046 -500 1046 -500 0 feedthrough
rlabel pdiffusion 1053 -500 1053 -500 0 feedthrough
rlabel pdiffusion 1060 -500 1060 -500 0 feedthrough
rlabel pdiffusion 1067 -500 1067 -500 0 feedthrough
rlabel pdiffusion 1074 -500 1074 -500 0 feedthrough
rlabel pdiffusion 1081 -500 1081 -500 0 feedthrough
rlabel pdiffusion 1088 -500 1088 -500 0 feedthrough
rlabel pdiffusion 1095 -500 1095 -500 0 feedthrough
rlabel pdiffusion 1102 -500 1102 -500 0 feedthrough
rlabel pdiffusion 1109 -500 1109 -500 0 feedthrough
rlabel pdiffusion 1116 -500 1116 -500 0 feedthrough
rlabel pdiffusion 1123 -500 1123 -500 0 feedthrough
rlabel pdiffusion 1130 -500 1130 -500 0 feedthrough
rlabel pdiffusion 1137 -500 1137 -500 0 feedthrough
rlabel pdiffusion 1144 -500 1144 -500 0 feedthrough
rlabel pdiffusion 1151 -500 1151 -500 0 feedthrough
rlabel pdiffusion 1158 -500 1158 -500 0 feedthrough
rlabel pdiffusion 1165 -500 1165 -500 0 feedthrough
rlabel pdiffusion 1172 -500 1172 -500 0 feedthrough
rlabel pdiffusion 1179 -500 1179 -500 0 feedthrough
rlabel pdiffusion 1186 -500 1186 -500 0 feedthrough
rlabel pdiffusion 1193 -500 1193 -500 0 cellNo=153
rlabel pdiffusion 1200 -500 1200 -500 0 feedthrough
rlabel pdiffusion 1207 -500 1207 -500 0 feedthrough
rlabel pdiffusion 1214 -500 1214 -500 0 feedthrough
rlabel pdiffusion 1221 -500 1221 -500 0 feedthrough
rlabel pdiffusion 1228 -500 1228 -500 0 feedthrough
rlabel pdiffusion 1235 -500 1235 -500 0 feedthrough
rlabel pdiffusion 1242 -500 1242 -500 0 feedthrough
rlabel pdiffusion 1249 -500 1249 -500 0 feedthrough
rlabel pdiffusion 1256 -500 1256 -500 0 feedthrough
rlabel pdiffusion 1263 -500 1263 -500 0 feedthrough
rlabel pdiffusion 1270 -500 1270 -500 0 feedthrough
rlabel pdiffusion 1277 -500 1277 -500 0 feedthrough
rlabel pdiffusion 1284 -500 1284 -500 0 feedthrough
rlabel pdiffusion 1291 -500 1291 -500 0 feedthrough
rlabel pdiffusion 1298 -500 1298 -500 0 feedthrough
rlabel pdiffusion 1305 -500 1305 -500 0 feedthrough
rlabel pdiffusion 1312 -500 1312 -500 0 feedthrough
rlabel pdiffusion 1319 -500 1319 -500 0 feedthrough
rlabel pdiffusion 1326 -500 1326 -500 0 feedthrough
rlabel pdiffusion 1333 -500 1333 -500 0 feedthrough
rlabel pdiffusion 1340 -500 1340 -500 0 feedthrough
rlabel pdiffusion 1347 -500 1347 -500 0 feedthrough
rlabel pdiffusion 1354 -500 1354 -500 0 feedthrough
rlabel pdiffusion 1361 -500 1361 -500 0 feedthrough
rlabel pdiffusion 1368 -500 1368 -500 0 feedthrough
rlabel pdiffusion 1375 -500 1375 -500 0 feedthrough
rlabel pdiffusion 1382 -500 1382 -500 0 feedthrough
rlabel pdiffusion 1389 -500 1389 -500 0 feedthrough
rlabel pdiffusion 1396 -500 1396 -500 0 feedthrough
rlabel pdiffusion 1403 -500 1403 -500 0 feedthrough
rlabel pdiffusion 1410 -500 1410 -500 0 feedthrough
rlabel pdiffusion 1417 -500 1417 -500 0 feedthrough
rlabel pdiffusion 1424 -500 1424 -500 0 feedthrough
rlabel pdiffusion 1431 -500 1431 -500 0 feedthrough
rlabel pdiffusion 1438 -500 1438 -500 0 feedthrough
rlabel pdiffusion 1445 -500 1445 -500 0 feedthrough
rlabel pdiffusion 1452 -500 1452 -500 0 feedthrough
rlabel pdiffusion 1459 -500 1459 -500 0 feedthrough
rlabel pdiffusion 1466 -500 1466 -500 0 feedthrough
rlabel pdiffusion 1473 -500 1473 -500 0 feedthrough
rlabel pdiffusion 1480 -500 1480 -500 0 feedthrough
rlabel pdiffusion 1487 -500 1487 -500 0 feedthrough
rlabel pdiffusion 1494 -500 1494 -500 0 feedthrough
rlabel pdiffusion 1501 -500 1501 -500 0 feedthrough
rlabel pdiffusion 1508 -500 1508 -500 0 feedthrough
rlabel pdiffusion 1515 -500 1515 -500 0 feedthrough
rlabel pdiffusion 1522 -500 1522 -500 0 cellNo=769
rlabel pdiffusion 1529 -500 1529 -500 0 feedthrough
rlabel pdiffusion 1711 -500 1711 -500 0 feedthrough
rlabel pdiffusion 3 -607 3 -607 0 cellNo=1017
rlabel pdiffusion 10 -607 10 -607 0 feedthrough
rlabel pdiffusion 17 -607 17 -607 0 cellNo=1079
rlabel pdiffusion 24 -607 24 -607 0 feedthrough
rlabel pdiffusion 31 -607 31 -607 0 cellNo=116
rlabel pdiffusion 38 -607 38 -607 0 cellNo=1077
rlabel pdiffusion 45 -607 45 -607 0 feedthrough
rlabel pdiffusion 52 -607 52 -607 0 feedthrough
rlabel pdiffusion 59 -607 59 -607 0 cellNo=257
rlabel pdiffusion 66 -607 66 -607 0 feedthrough
rlabel pdiffusion 73 -607 73 -607 0 feedthrough
rlabel pdiffusion 80 -607 80 -607 0 feedthrough
rlabel pdiffusion 87 -607 87 -607 0 feedthrough
rlabel pdiffusion 94 -607 94 -607 0 feedthrough
rlabel pdiffusion 101 -607 101 -607 0 cellNo=108
rlabel pdiffusion 108 -607 108 -607 0 feedthrough
rlabel pdiffusion 115 -607 115 -607 0 feedthrough
rlabel pdiffusion 122 -607 122 -607 0 feedthrough
rlabel pdiffusion 129 -607 129 -607 0 feedthrough
rlabel pdiffusion 136 -607 136 -607 0 feedthrough
rlabel pdiffusion 143 -607 143 -607 0 feedthrough
rlabel pdiffusion 150 -607 150 -607 0 cellNo=96
rlabel pdiffusion 157 -607 157 -607 0 feedthrough
rlabel pdiffusion 164 -607 164 -607 0 feedthrough
rlabel pdiffusion 171 -607 171 -607 0 feedthrough
rlabel pdiffusion 178 -607 178 -607 0 feedthrough
rlabel pdiffusion 185 -607 185 -607 0 cellNo=228
rlabel pdiffusion 192 -607 192 -607 0 feedthrough
rlabel pdiffusion 199 -607 199 -607 0 feedthrough
rlabel pdiffusion 206 -607 206 -607 0 feedthrough
rlabel pdiffusion 213 -607 213 -607 0 feedthrough
rlabel pdiffusion 220 -607 220 -607 0 feedthrough
rlabel pdiffusion 227 -607 227 -607 0 feedthrough
rlabel pdiffusion 234 -607 234 -607 0 cellNo=904
rlabel pdiffusion 241 -607 241 -607 0 cellNo=277
rlabel pdiffusion 248 -607 248 -607 0 feedthrough
rlabel pdiffusion 255 -607 255 -607 0 feedthrough
rlabel pdiffusion 262 -607 262 -607 0 feedthrough
rlabel pdiffusion 269 -607 269 -607 0 feedthrough
rlabel pdiffusion 276 -607 276 -607 0 feedthrough
rlabel pdiffusion 283 -607 283 -607 0 feedthrough
rlabel pdiffusion 290 -607 290 -607 0 feedthrough
rlabel pdiffusion 297 -607 297 -607 0 feedthrough
rlabel pdiffusion 304 -607 304 -607 0 feedthrough
rlabel pdiffusion 311 -607 311 -607 0 feedthrough
rlabel pdiffusion 318 -607 318 -607 0 cellNo=186
rlabel pdiffusion 325 -607 325 -607 0 feedthrough
rlabel pdiffusion 332 -607 332 -607 0 feedthrough
rlabel pdiffusion 339 -607 339 -607 0 cellNo=466
rlabel pdiffusion 346 -607 346 -607 0 feedthrough
rlabel pdiffusion 353 -607 353 -607 0 feedthrough
rlabel pdiffusion 360 -607 360 -607 0 feedthrough
rlabel pdiffusion 367 -607 367 -607 0 feedthrough
rlabel pdiffusion 374 -607 374 -607 0 feedthrough
rlabel pdiffusion 381 -607 381 -607 0 cellNo=397
rlabel pdiffusion 388 -607 388 -607 0 feedthrough
rlabel pdiffusion 395 -607 395 -607 0 feedthrough
rlabel pdiffusion 402 -607 402 -607 0 feedthrough
rlabel pdiffusion 409 -607 409 -607 0 feedthrough
rlabel pdiffusion 416 -607 416 -607 0 feedthrough
rlabel pdiffusion 423 -607 423 -607 0 feedthrough
rlabel pdiffusion 430 -607 430 -607 0 cellNo=23
rlabel pdiffusion 437 -607 437 -607 0 feedthrough
rlabel pdiffusion 444 -607 444 -607 0 feedthrough
rlabel pdiffusion 451 -607 451 -607 0 cellNo=449
rlabel pdiffusion 458 -607 458 -607 0 cellNo=613
rlabel pdiffusion 465 -607 465 -607 0 feedthrough
rlabel pdiffusion 472 -607 472 -607 0 feedthrough
rlabel pdiffusion 479 -607 479 -607 0 feedthrough
rlabel pdiffusion 486 -607 486 -607 0 feedthrough
rlabel pdiffusion 493 -607 493 -607 0 feedthrough
rlabel pdiffusion 500 -607 500 -607 0 feedthrough
rlabel pdiffusion 507 -607 507 -607 0 feedthrough
rlabel pdiffusion 514 -607 514 -607 0 cellNo=551
rlabel pdiffusion 521 -607 521 -607 0 feedthrough
rlabel pdiffusion 528 -607 528 -607 0 cellNo=160
rlabel pdiffusion 535 -607 535 -607 0 feedthrough
rlabel pdiffusion 542 -607 542 -607 0 feedthrough
rlabel pdiffusion 549 -607 549 -607 0 feedthrough
rlabel pdiffusion 556 -607 556 -607 0 feedthrough
rlabel pdiffusion 563 -607 563 -607 0 feedthrough
rlabel pdiffusion 570 -607 570 -607 0 feedthrough
rlabel pdiffusion 577 -607 577 -607 0 cellNo=832
rlabel pdiffusion 584 -607 584 -607 0 cellNo=318
rlabel pdiffusion 591 -607 591 -607 0 cellNo=885
rlabel pdiffusion 598 -607 598 -607 0 feedthrough
rlabel pdiffusion 605 -607 605 -607 0 feedthrough
rlabel pdiffusion 612 -607 612 -607 0 feedthrough
rlabel pdiffusion 619 -607 619 -607 0 feedthrough
rlabel pdiffusion 626 -607 626 -607 0 feedthrough
rlabel pdiffusion 633 -607 633 -607 0 cellNo=540
rlabel pdiffusion 640 -607 640 -607 0 feedthrough
rlabel pdiffusion 647 -607 647 -607 0 feedthrough
rlabel pdiffusion 654 -607 654 -607 0 feedthrough
rlabel pdiffusion 661 -607 661 -607 0 feedthrough
rlabel pdiffusion 668 -607 668 -607 0 feedthrough
rlabel pdiffusion 675 -607 675 -607 0 cellNo=306
rlabel pdiffusion 682 -607 682 -607 0 feedthrough
rlabel pdiffusion 689 -607 689 -607 0 feedthrough
rlabel pdiffusion 696 -607 696 -607 0 cellNo=281
rlabel pdiffusion 703 -607 703 -607 0 feedthrough
rlabel pdiffusion 710 -607 710 -607 0 feedthrough
rlabel pdiffusion 717 -607 717 -607 0 feedthrough
rlabel pdiffusion 724 -607 724 -607 0 feedthrough
rlabel pdiffusion 731 -607 731 -607 0 feedthrough
rlabel pdiffusion 738 -607 738 -607 0 feedthrough
rlabel pdiffusion 745 -607 745 -607 0 feedthrough
rlabel pdiffusion 752 -607 752 -607 0 feedthrough
rlabel pdiffusion 759 -607 759 -607 0 feedthrough
rlabel pdiffusion 766 -607 766 -607 0 feedthrough
rlabel pdiffusion 773 -607 773 -607 0 feedthrough
rlabel pdiffusion 780 -607 780 -607 0 cellNo=468
rlabel pdiffusion 787 -607 787 -607 0 feedthrough
rlabel pdiffusion 794 -607 794 -607 0 feedthrough
rlabel pdiffusion 801 -607 801 -607 0 feedthrough
rlabel pdiffusion 808 -607 808 -607 0 feedthrough
rlabel pdiffusion 815 -607 815 -607 0 feedthrough
rlabel pdiffusion 822 -607 822 -607 0 cellNo=741
rlabel pdiffusion 829 -607 829 -607 0 feedthrough
rlabel pdiffusion 836 -607 836 -607 0 feedthrough
rlabel pdiffusion 843 -607 843 -607 0 cellNo=149
rlabel pdiffusion 850 -607 850 -607 0 cellNo=463
rlabel pdiffusion 857 -607 857 -607 0 feedthrough
rlabel pdiffusion 864 -607 864 -607 0 cellNo=358
rlabel pdiffusion 871 -607 871 -607 0 cellNo=61
rlabel pdiffusion 878 -607 878 -607 0 feedthrough
rlabel pdiffusion 885 -607 885 -607 0 feedthrough
rlabel pdiffusion 892 -607 892 -607 0 cellNo=300
rlabel pdiffusion 899 -607 899 -607 0 feedthrough
rlabel pdiffusion 906 -607 906 -607 0 feedthrough
rlabel pdiffusion 913 -607 913 -607 0 cellNo=286
rlabel pdiffusion 920 -607 920 -607 0 feedthrough
rlabel pdiffusion 927 -607 927 -607 0 feedthrough
rlabel pdiffusion 934 -607 934 -607 0 cellNo=528
rlabel pdiffusion 941 -607 941 -607 0 feedthrough
rlabel pdiffusion 948 -607 948 -607 0 feedthrough
rlabel pdiffusion 955 -607 955 -607 0 feedthrough
rlabel pdiffusion 962 -607 962 -607 0 feedthrough
rlabel pdiffusion 969 -607 969 -607 0 feedthrough
rlabel pdiffusion 976 -607 976 -607 0 feedthrough
rlabel pdiffusion 983 -607 983 -607 0 feedthrough
rlabel pdiffusion 990 -607 990 -607 0 feedthrough
rlabel pdiffusion 997 -607 997 -607 0 feedthrough
rlabel pdiffusion 1004 -607 1004 -607 0 feedthrough
rlabel pdiffusion 1011 -607 1011 -607 0 feedthrough
rlabel pdiffusion 1018 -607 1018 -607 0 feedthrough
rlabel pdiffusion 1025 -607 1025 -607 0 feedthrough
rlabel pdiffusion 1032 -607 1032 -607 0 feedthrough
rlabel pdiffusion 1039 -607 1039 -607 0 feedthrough
rlabel pdiffusion 1046 -607 1046 -607 0 feedthrough
rlabel pdiffusion 1053 -607 1053 -607 0 cellNo=651
rlabel pdiffusion 1060 -607 1060 -607 0 feedthrough
rlabel pdiffusion 1067 -607 1067 -607 0 feedthrough
rlabel pdiffusion 1074 -607 1074 -607 0 feedthrough
rlabel pdiffusion 1081 -607 1081 -607 0 feedthrough
rlabel pdiffusion 1088 -607 1088 -607 0 feedthrough
rlabel pdiffusion 1095 -607 1095 -607 0 feedthrough
rlabel pdiffusion 1102 -607 1102 -607 0 feedthrough
rlabel pdiffusion 1109 -607 1109 -607 0 feedthrough
rlabel pdiffusion 1116 -607 1116 -607 0 feedthrough
rlabel pdiffusion 1123 -607 1123 -607 0 feedthrough
rlabel pdiffusion 1130 -607 1130 -607 0 feedthrough
rlabel pdiffusion 1137 -607 1137 -607 0 feedthrough
rlabel pdiffusion 1144 -607 1144 -607 0 feedthrough
rlabel pdiffusion 1151 -607 1151 -607 0 feedthrough
rlabel pdiffusion 1158 -607 1158 -607 0 feedthrough
rlabel pdiffusion 1165 -607 1165 -607 0 feedthrough
rlabel pdiffusion 1172 -607 1172 -607 0 feedthrough
rlabel pdiffusion 1179 -607 1179 -607 0 feedthrough
rlabel pdiffusion 1186 -607 1186 -607 0 feedthrough
rlabel pdiffusion 1193 -607 1193 -607 0 feedthrough
rlabel pdiffusion 1200 -607 1200 -607 0 feedthrough
rlabel pdiffusion 1207 -607 1207 -607 0 feedthrough
rlabel pdiffusion 1214 -607 1214 -607 0 feedthrough
rlabel pdiffusion 1221 -607 1221 -607 0 feedthrough
rlabel pdiffusion 1228 -607 1228 -607 0 feedthrough
rlabel pdiffusion 1235 -607 1235 -607 0 feedthrough
rlabel pdiffusion 1242 -607 1242 -607 0 feedthrough
rlabel pdiffusion 1249 -607 1249 -607 0 feedthrough
rlabel pdiffusion 1256 -607 1256 -607 0 feedthrough
rlabel pdiffusion 1263 -607 1263 -607 0 feedthrough
rlabel pdiffusion 1270 -607 1270 -607 0 feedthrough
rlabel pdiffusion 1277 -607 1277 -607 0 feedthrough
rlabel pdiffusion 1284 -607 1284 -607 0 feedthrough
rlabel pdiffusion 1291 -607 1291 -607 0 feedthrough
rlabel pdiffusion 1298 -607 1298 -607 0 feedthrough
rlabel pdiffusion 1305 -607 1305 -607 0 feedthrough
rlabel pdiffusion 1312 -607 1312 -607 0 feedthrough
rlabel pdiffusion 1319 -607 1319 -607 0 feedthrough
rlabel pdiffusion 1326 -607 1326 -607 0 feedthrough
rlabel pdiffusion 1333 -607 1333 -607 0 feedthrough
rlabel pdiffusion 1340 -607 1340 -607 0 feedthrough
rlabel pdiffusion 1347 -607 1347 -607 0 feedthrough
rlabel pdiffusion 1354 -607 1354 -607 0 feedthrough
rlabel pdiffusion 1361 -607 1361 -607 0 feedthrough
rlabel pdiffusion 1368 -607 1368 -607 0 feedthrough
rlabel pdiffusion 1375 -607 1375 -607 0 feedthrough
rlabel pdiffusion 1382 -607 1382 -607 0 feedthrough
rlabel pdiffusion 1389 -607 1389 -607 0 feedthrough
rlabel pdiffusion 1396 -607 1396 -607 0 feedthrough
rlabel pdiffusion 1403 -607 1403 -607 0 feedthrough
rlabel pdiffusion 1410 -607 1410 -607 0 feedthrough
rlabel pdiffusion 1417 -607 1417 -607 0 feedthrough
rlabel pdiffusion 1424 -607 1424 -607 0 feedthrough
rlabel pdiffusion 1431 -607 1431 -607 0 feedthrough
rlabel pdiffusion 1438 -607 1438 -607 0 feedthrough
rlabel pdiffusion 1445 -607 1445 -607 0 feedthrough
rlabel pdiffusion 1452 -607 1452 -607 0 feedthrough
rlabel pdiffusion 1459 -607 1459 -607 0 feedthrough
rlabel pdiffusion 1466 -607 1466 -607 0 cellNo=921
rlabel pdiffusion 1473 -607 1473 -607 0 feedthrough
rlabel pdiffusion 1480 -607 1480 -607 0 feedthrough
rlabel pdiffusion 1487 -607 1487 -607 0 feedthrough
rlabel pdiffusion 1494 -607 1494 -607 0 feedthrough
rlabel pdiffusion 1501 -607 1501 -607 0 feedthrough
rlabel pdiffusion 1508 -607 1508 -607 0 feedthrough
rlabel pdiffusion 1515 -607 1515 -607 0 feedthrough
rlabel pdiffusion 1522 -607 1522 -607 0 feedthrough
rlabel pdiffusion 1536 -607 1536 -607 0 feedthrough
rlabel pdiffusion 1557 -607 1557 -607 0 feedthrough
rlabel pdiffusion 1739 -607 1739 -607 0 feedthrough
rlabel pdiffusion 1760 -607 1760 -607 0 feedthrough
rlabel pdiffusion 1767 -607 1767 -607 0 feedthrough
rlabel pdiffusion 3 -716 3 -716 0 cellNo=1085
rlabel pdiffusion 10 -716 10 -716 0 feedthrough
rlabel pdiffusion 17 -716 17 -716 0 feedthrough
rlabel pdiffusion 24 -716 24 -716 0 feedthrough
rlabel pdiffusion 31 -716 31 -716 0 feedthrough
rlabel pdiffusion 38 -716 38 -716 0 feedthrough
rlabel pdiffusion 45 -716 45 -716 0 feedthrough
rlabel pdiffusion 52 -716 52 -716 0 feedthrough
rlabel pdiffusion 59 -716 59 -716 0 feedthrough
rlabel pdiffusion 66 -716 66 -716 0 feedthrough
rlabel pdiffusion 73 -716 73 -716 0 feedthrough
rlabel pdiffusion 80 -716 80 -716 0 feedthrough
rlabel pdiffusion 87 -716 87 -716 0 feedthrough
rlabel pdiffusion 94 -716 94 -716 0 cellNo=26
rlabel pdiffusion 101 -716 101 -716 0 feedthrough
rlabel pdiffusion 108 -716 108 -716 0 feedthrough
rlabel pdiffusion 115 -716 115 -716 0 cellNo=372
rlabel pdiffusion 122 -716 122 -716 0 feedthrough
rlabel pdiffusion 129 -716 129 -716 0 feedthrough
rlabel pdiffusion 136 -716 136 -716 0 cellNo=302
rlabel pdiffusion 143 -716 143 -716 0 cellNo=589
rlabel pdiffusion 150 -716 150 -716 0 feedthrough
rlabel pdiffusion 157 -716 157 -716 0 feedthrough
rlabel pdiffusion 164 -716 164 -716 0 feedthrough
rlabel pdiffusion 171 -716 171 -716 0 cellNo=453
rlabel pdiffusion 178 -716 178 -716 0 feedthrough
rlabel pdiffusion 185 -716 185 -716 0 cellNo=563
rlabel pdiffusion 192 -716 192 -716 0 feedthrough
rlabel pdiffusion 199 -716 199 -716 0 feedthrough
rlabel pdiffusion 206 -716 206 -716 0 feedthrough
rlabel pdiffusion 213 -716 213 -716 0 feedthrough
rlabel pdiffusion 220 -716 220 -716 0 feedthrough
rlabel pdiffusion 227 -716 227 -716 0 feedthrough
rlabel pdiffusion 234 -716 234 -716 0 cellNo=571
rlabel pdiffusion 241 -716 241 -716 0 feedthrough
rlabel pdiffusion 248 -716 248 -716 0 feedthrough
rlabel pdiffusion 255 -716 255 -716 0 feedthrough
rlabel pdiffusion 262 -716 262 -716 0 feedthrough
rlabel pdiffusion 269 -716 269 -716 0 feedthrough
rlabel pdiffusion 276 -716 276 -716 0 feedthrough
rlabel pdiffusion 283 -716 283 -716 0 feedthrough
rlabel pdiffusion 290 -716 290 -716 0 feedthrough
rlabel pdiffusion 297 -716 297 -716 0 feedthrough
rlabel pdiffusion 304 -716 304 -716 0 feedthrough
rlabel pdiffusion 311 -716 311 -716 0 feedthrough
rlabel pdiffusion 318 -716 318 -716 0 feedthrough
rlabel pdiffusion 325 -716 325 -716 0 feedthrough
rlabel pdiffusion 332 -716 332 -716 0 feedthrough
rlabel pdiffusion 339 -716 339 -716 0 feedthrough
rlabel pdiffusion 346 -716 346 -716 0 feedthrough
rlabel pdiffusion 353 -716 353 -716 0 feedthrough
rlabel pdiffusion 360 -716 360 -716 0 cellNo=513
rlabel pdiffusion 367 -716 367 -716 0 feedthrough
rlabel pdiffusion 374 -716 374 -716 0 feedthrough
rlabel pdiffusion 381 -716 381 -716 0 feedthrough
rlabel pdiffusion 388 -716 388 -716 0 feedthrough
rlabel pdiffusion 395 -716 395 -716 0 feedthrough
rlabel pdiffusion 402 -716 402 -716 0 feedthrough
rlabel pdiffusion 409 -716 409 -716 0 feedthrough
rlabel pdiffusion 416 -716 416 -716 0 feedthrough
rlabel pdiffusion 423 -716 423 -716 0 feedthrough
rlabel pdiffusion 430 -716 430 -716 0 feedthrough
rlabel pdiffusion 437 -716 437 -716 0 feedthrough
rlabel pdiffusion 444 -716 444 -716 0 feedthrough
rlabel pdiffusion 451 -716 451 -716 0 feedthrough
rlabel pdiffusion 458 -716 458 -716 0 feedthrough
rlabel pdiffusion 465 -716 465 -716 0 cellNo=750
rlabel pdiffusion 472 -716 472 -716 0 feedthrough
rlabel pdiffusion 479 -716 479 -716 0 cellNo=124
rlabel pdiffusion 486 -716 486 -716 0 feedthrough
rlabel pdiffusion 493 -716 493 -716 0 feedthrough
rlabel pdiffusion 500 -716 500 -716 0 feedthrough
rlabel pdiffusion 507 -716 507 -716 0 cellNo=289
rlabel pdiffusion 514 -716 514 -716 0 feedthrough
rlabel pdiffusion 521 -716 521 -716 0 feedthrough
rlabel pdiffusion 528 -716 528 -716 0 feedthrough
rlabel pdiffusion 535 -716 535 -716 0 feedthrough
rlabel pdiffusion 542 -716 542 -716 0 cellNo=958
rlabel pdiffusion 549 -716 549 -716 0 feedthrough
rlabel pdiffusion 556 -716 556 -716 0 cellNo=441
rlabel pdiffusion 563 -716 563 -716 0 feedthrough
rlabel pdiffusion 570 -716 570 -716 0 feedthrough
rlabel pdiffusion 577 -716 577 -716 0 feedthrough
rlabel pdiffusion 584 -716 584 -716 0 feedthrough
rlabel pdiffusion 591 -716 591 -716 0 feedthrough
rlabel pdiffusion 598 -716 598 -716 0 cellNo=200
rlabel pdiffusion 605 -716 605 -716 0 feedthrough
rlabel pdiffusion 612 -716 612 -716 0 feedthrough
rlabel pdiffusion 619 -716 619 -716 0 cellNo=595
rlabel pdiffusion 626 -716 626 -716 0 feedthrough
rlabel pdiffusion 633 -716 633 -716 0 feedthrough
rlabel pdiffusion 640 -716 640 -716 0 feedthrough
rlabel pdiffusion 647 -716 647 -716 0 cellNo=243
rlabel pdiffusion 654 -716 654 -716 0 feedthrough
rlabel pdiffusion 661 -716 661 -716 0 feedthrough
rlabel pdiffusion 668 -716 668 -716 0 feedthrough
rlabel pdiffusion 675 -716 675 -716 0 feedthrough
rlabel pdiffusion 682 -716 682 -716 0 feedthrough
rlabel pdiffusion 689 -716 689 -716 0 cellNo=312
rlabel pdiffusion 696 -716 696 -716 0 feedthrough
rlabel pdiffusion 703 -716 703 -716 0 feedthrough
rlabel pdiffusion 710 -716 710 -716 0 cellNo=6
rlabel pdiffusion 717 -716 717 -716 0 cellNo=234
rlabel pdiffusion 724 -716 724 -716 0 feedthrough
rlabel pdiffusion 731 -716 731 -716 0 feedthrough
rlabel pdiffusion 738 -716 738 -716 0 cellNo=313
rlabel pdiffusion 745 -716 745 -716 0 feedthrough
rlabel pdiffusion 752 -716 752 -716 0 feedthrough
rlabel pdiffusion 759 -716 759 -716 0 cellNo=101
rlabel pdiffusion 766 -716 766 -716 0 feedthrough
rlabel pdiffusion 773 -716 773 -716 0 feedthrough
rlabel pdiffusion 780 -716 780 -716 0 cellNo=572
rlabel pdiffusion 787 -716 787 -716 0 feedthrough
rlabel pdiffusion 794 -716 794 -716 0 cellNo=951
rlabel pdiffusion 801 -716 801 -716 0 feedthrough
rlabel pdiffusion 808 -716 808 -716 0 feedthrough
rlabel pdiffusion 815 -716 815 -716 0 feedthrough
rlabel pdiffusion 822 -716 822 -716 0 feedthrough
rlabel pdiffusion 829 -716 829 -716 0 cellNo=262
rlabel pdiffusion 836 -716 836 -716 0 feedthrough
rlabel pdiffusion 843 -716 843 -716 0 cellNo=604
rlabel pdiffusion 850 -716 850 -716 0 feedthrough
rlabel pdiffusion 857 -716 857 -716 0 feedthrough
rlabel pdiffusion 864 -716 864 -716 0 feedthrough
rlabel pdiffusion 871 -716 871 -716 0 feedthrough
rlabel pdiffusion 878 -716 878 -716 0 feedthrough
rlabel pdiffusion 885 -716 885 -716 0 feedthrough
rlabel pdiffusion 892 -716 892 -716 0 feedthrough
rlabel pdiffusion 899 -716 899 -716 0 cellNo=114
rlabel pdiffusion 906 -716 906 -716 0 cellNo=923
rlabel pdiffusion 913 -716 913 -716 0 feedthrough
rlabel pdiffusion 920 -716 920 -716 0 cellNo=808
rlabel pdiffusion 927 -716 927 -716 0 feedthrough
rlabel pdiffusion 934 -716 934 -716 0 feedthrough
rlabel pdiffusion 941 -716 941 -716 0 feedthrough
rlabel pdiffusion 948 -716 948 -716 0 feedthrough
rlabel pdiffusion 955 -716 955 -716 0 feedthrough
rlabel pdiffusion 962 -716 962 -716 0 feedthrough
rlabel pdiffusion 969 -716 969 -716 0 cellNo=492
rlabel pdiffusion 976 -716 976 -716 0 feedthrough
rlabel pdiffusion 983 -716 983 -716 0 feedthrough
rlabel pdiffusion 990 -716 990 -716 0 feedthrough
rlabel pdiffusion 997 -716 997 -716 0 cellNo=196
rlabel pdiffusion 1004 -716 1004 -716 0 feedthrough
rlabel pdiffusion 1011 -716 1011 -716 0 feedthrough
rlabel pdiffusion 1018 -716 1018 -716 0 cellNo=104
rlabel pdiffusion 1025 -716 1025 -716 0 feedthrough
rlabel pdiffusion 1032 -716 1032 -716 0 feedthrough
rlabel pdiffusion 1039 -716 1039 -716 0 feedthrough
rlabel pdiffusion 1046 -716 1046 -716 0 feedthrough
rlabel pdiffusion 1053 -716 1053 -716 0 feedthrough
rlabel pdiffusion 1060 -716 1060 -716 0 feedthrough
rlabel pdiffusion 1067 -716 1067 -716 0 feedthrough
rlabel pdiffusion 1074 -716 1074 -716 0 feedthrough
rlabel pdiffusion 1081 -716 1081 -716 0 feedthrough
rlabel pdiffusion 1088 -716 1088 -716 0 feedthrough
rlabel pdiffusion 1095 -716 1095 -716 0 feedthrough
rlabel pdiffusion 1102 -716 1102 -716 0 feedthrough
rlabel pdiffusion 1109 -716 1109 -716 0 feedthrough
rlabel pdiffusion 1116 -716 1116 -716 0 feedthrough
rlabel pdiffusion 1123 -716 1123 -716 0 cellNo=695
rlabel pdiffusion 1130 -716 1130 -716 0 feedthrough
rlabel pdiffusion 1137 -716 1137 -716 0 feedthrough
rlabel pdiffusion 1144 -716 1144 -716 0 feedthrough
rlabel pdiffusion 1151 -716 1151 -716 0 feedthrough
rlabel pdiffusion 1158 -716 1158 -716 0 feedthrough
rlabel pdiffusion 1165 -716 1165 -716 0 feedthrough
rlabel pdiffusion 1172 -716 1172 -716 0 feedthrough
rlabel pdiffusion 1179 -716 1179 -716 0 feedthrough
rlabel pdiffusion 1186 -716 1186 -716 0 feedthrough
rlabel pdiffusion 1193 -716 1193 -716 0 feedthrough
rlabel pdiffusion 1200 -716 1200 -716 0 feedthrough
rlabel pdiffusion 1207 -716 1207 -716 0 feedthrough
rlabel pdiffusion 1214 -716 1214 -716 0 feedthrough
rlabel pdiffusion 1221 -716 1221 -716 0 feedthrough
rlabel pdiffusion 1228 -716 1228 -716 0 feedthrough
rlabel pdiffusion 1235 -716 1235 -716 0 feedthrough
rlabel pdiffusion 1242 -716 1242 -716 0 feedthrough
rlabel pdiffusion 1249 -716 1249 -716 0 feedthrough
rlabel pdiffusion 1256 -716 1256 -716 0 feedthrough
rlabel pdiffusion 1263 -716 1263 -716 0 feedthrough
rlabel pdiffusion 1270 -716 1270 -716 0 feedthrough
rlabel pdiffusion 1277 -716 1277 -716 0 feedthrough
rlabel pdiffusion 1284 -716 1284 -716 0 feedthrough
rlabel pdiffusion 1291 -716 1291 -716 0 feedthrough
rlabel pdiffusion 1298 -716 1298 -716 0 feedthrough
rlabel pdiffusion 1305 -716 1305 -716 0 feedthrough
rlabel pdiffusion 1312 -716 1312 -716 0 feedthrough
rlabel pdiffusion 1319 -716 1319 -716 0 feedthrough
rlabel pdiffusion 1326 -716 1326 -716 0 feedthrough
rlabel pdiffusion 1333 -716 1333 -716 0 feedthrough
rlabel pdiffusion 1340 -716 1340 -716 0 feedthrough
rlabel pdiffusion 1347 -716 1347 -716 0 feedthrough
rlabel pdiffusion 1354 -716 1354 -716 0 feedthrough
rlabel pdiffusion 1361 -716 1361 -716 0 feedthrough
rlabel pdiffusion 1368 -716 1368 -716 0 feedthrough
rlabel pdiffusion 1375 -716 1375 -716 0 feedthrough
rlabel pdiffusion 1382 -716 1382 -716 0 feedthrough
rlabel pdiffusion 1389 -716 1389 -716 0 feedthrough
rlabel pdiffusion 1396 -716 1396 -716 0 feedthrough
rlabel pdiffusion 1403 -716 1403 -716 0 feedthrough
rlabel pdiffusion 1410 -716 1410 -716 0 feedthrough
rlabel pdiffusion 1417 -716 1417 -716 0 feedthrough
rlabel pdiffusion 1424 -716 1424 -716 0 feedthrough
rlabel pdiffusion 1431 -716 1431 -716 0 feedthrough
rlabel pdiffusion 1438 -716 1438 -716 0 feedthrough
rlabel pdiffusion 1445 -716 1445 -716 0 feedthrough
rlabel pdiffusion 1452 -716 1452 -716 0 feedthrough
rlabel pdiffusion 1459 -716 1459 -716 0 feedthrough
rlabel pdiffusion 1466 -716 1466 -716 0 feedthrough
rlabel pdiffusion 1473 -716 1473 -716 0 feedthrough
rlabel pdiffusion 1480 -716 1480 -716 0 feedthrough
rlabel pdiffusion 1487 -716 1487 -716 0 feedthrough
rlabel pdiffusion 1494 -716 1494 -716 0 feedthrough
rlabel pdiffusion 1501 -716 1501 -716 0 feedthrough
rlabel pdiffusion 1508 -716 1508 -716 0 feedthrough
rlabel pdiffusion 1515 -716 1515 -716 0 feedthrough
rlabel pdiffusion 1522 -716 1522 -716 0 feedthrough
rlabel pdiffusion 1529 -716 1529 -716 0 feedthrough
rlabel pdiffusion 1536 -716 1536 -716 0 feedthrough
rlabel pdiffusion 1543 -716 1543 -716 0 feedthrough
rlabel pdiffusion 1550 -716 1550 -716 0 feedthrough
rlabel pdiffusion 1557 -716 1557 -716 0 feedthrough
rlabel pdiffusion 1564 -716 1564 -716 0 feedthrough
rlabel pdiffusion 1571 -716 1571 -716 0 feedthrough
rlabel pdiffusion 1578 -716 1578 -716 0 feedthrough
rlabel pdiffusion 1585 -716 1585 -716 0 feedthrough
rlabel pdiffusion 1592 -716 1592 -716 0 feedthrough
rlabel pdiffusion 1599 -716 1599 -716 0 feedthrough
rlabel pdiffusion 1606 -716 1606 -716 0 feedthrough
rlabel pdiffusion 1613 -716 1613 -716 0 feedthrough
rlabel pdiffusion 1620 -716 1620 -716 0 feedthrough
rlabel pdiffusion 1627 -716 1627 -716 0 feedthrough
rlabel pdiffusion 1634 -716 1634 -716 0 feedthrough
rlabel pdiffusion 1641 -716 1641 -716 0 feedthrough
rlabel pdiffusion 1648 -716 1648 -716 0 feedthrough
rlabel pdiffusion 1655 -716 1655 -716 0 cellNo=320
rlabel pdiffusion 1662 -716 1662 -716 0 feedthrough
rlabel pdiffusion 1669 -716 1669 -716 0 cellNo=143
rlabel pdiffusion 1788 -716 1788 -716 0 feedthrough
rlabel pdiffusion 1795 -716 1795 -716 0 feedthrough
rlabel pdiffusion 1802 -716 1802 -716 0 feedthrough
rlabel pdiffusion 1823 -716 1823 -716 0 feedthrough
rlabel pdiffusion 1858 -716 1858 -716 0 feedthrough
rlabel pdiffusion 3 -861 3 -861 0 cellNo=1019
rlabel pdiffusion 10 -861 10 -861 0 feedthrough
rlabel pdiffusion 17 -861 17 -861 0 cellNo=431
rlabel pdiffusion 24 -861 24 -861 0 feedthrough
rlabel pdiffusion 31 -861 31 -861 0 feedthrough
rlabel pdiffusion 38 -861 38 -861 0 feedthrough
rlabel pdiffusion 45 -861 45 -861 0 cellNo=498
rlabel pdiffusion 52 -861 52 -861 0 cellNo=555
rlabel pdiffusion 59 -861 59 -861 0 feedthrough
rlabel pdiffusion 66 -861 66 -861 0 feedthrough
rlabel pdiffusion 73 -861 73 -861 0 feedthrough
rlabel pdiffusion 80 -861 80 -861 0 cellNo=190
rlabel pdiffusion 87 -861 87 -861 0 feedthrough
rlabel pdiffusion 94 -861 94 -861 0 feedthrough
rlabel pdiffusion 101 -861 101 -861 0 feedthrough
rlabel pdiffusion 108 -861 108 -861 0 feedthrough
rlabel pdiffusion 115 -861 115 -861 0 feedthrough
rlabel pdiffusion 122 -861 122 -861 0 cellNo=401
rlabel pdiffusion 129 -861 129 -861 0 feedthrough
rlabel pdiffusion 136 -861 136 -861 0 feedthrough
rlabel pdiffusion 143 -861 143 -861 0 feedthrough
rlabel pdiffusion 150 -861 150 -861 0 feedthrough
rlabel pdiffusion 157 -861 157 -861 0 feedthrough
rlabel pdiffusion 164 -861 164 -861 0 cellNo=830
rlabel pdiffusion 171 -861 171 -861 0 feedthrough
rlabel pdiffusion 178 -861 178 -861 0 cellNo=993
rlabel pdiffusion 185 -861 185 -861 0 feedthrough
rlabel pdiffusion 192 -861 192 -861 0 cellNo=52
rlabel pdiffusion 199 -861 199 -861 0 cellNo=980
rlabel pdiffusion 206 -861 206 -861 0 feedthrough
rlabel pdiffusion 213 -861 213 -861 0 feedthrough
rlabel pdiffusion 220 -861 220 -861 0 feedthrough
rlabel pdiffusion 227 -861 227 -861 0 feedthrough
rlabel pdiffusion 234 -861 234 -861 0 feedthrough
rlabel pdiffusion 241 -861 241 -861 0 feedthrough
rlabel pdiffusion 248 -861 248 -861 0 feedthrough
rlabel pdiffusion 255 -861 255 -861 0 feedthrough
rlabel pdiffusion 262 -861 262 -861 0 feedthrough
rlabel pdiffusion 269 -861 269 -861 0 feedthrough
rlabel pdiffusion 276 -861 276 -861 0 feedthrough
rlabel pdiffusion 283 -861 283 -861 0 feedthrough
rlabel pdiffusion 290 -861 290 -861 0 feedthrough
rlabel pdiffusion 297 -861 297 -861 0 feedthrough
rlabel pdiffusion 304 -861 304 -861 0 feedthrough
rlabel pdiffusion 311 -861 311 -861 0 feedthrough
rlabel pdiffusion 318 -861 318 -861 0 feedthrough
rlabel pdiffusion 325 -861 325 -861 0 feedthrough
rlabel pdiffusion 332 -861 332 -861 0 feedthrough
rlabel pdiffusion 339 -861 339 -861 0 feedthrough
rlabel pdiffusion 346 -861 346 -861 0 feedthrough
rlabel pdiffusion 353 -861 353 -861 0 feedthrough
rlabel pdiffusion 360 -861 360 -861 0 feedthrough
rlabel pdiffusion 367 -861 367 -861 0 feedthrough
rlabel pdiffusion 374 -861 374 -861 0 feedthrough
rlabel pdiffusion 381 -861 381 -861 0 feedthrough
rlabel pdiffusion 388 -861 388 -861 0 feedthrough
rlabel pdiffusion 395 -861 395 -861 0 feedthrough
rlabel pdiffusion 402 -861 402 -861 0 feedthrough
rlabel pdiffusion 409 -861 409 -861 0 feedthrough
rlabel pdiffusion 416 -861 416 -861 0 feedthrough
rlabel pdiffusion 423 -861 423 -861 0 feedthrough
rlabel pdiffusion 430 -861 430 -861 0 feedthrough
rlabel pdiffusion 437 -861 437 -861 0 cellNo=459
rlabel pdiffusion 444 -861 444 -861 0 feedthrough
rlabel pdiffusion 451 -861 451 -861 0 feedthrough
rlabel pdiffusion 458 -861 458 -861 0 feedthrough
rlabel pdiffusion 465 -861 465 -861 0 feedthrough
rlabel pdiffusion 472 -861 472 -861 0 feedthrough
rlabel pdiffusion 479 -861 479 -861 0 feedthrough
rlabel pdiffusion 486 -861 486 -861 0 feedthrough
rlabel pdiffusion 493 -861 493 -861 0 cellNo=227
rlabel pdiffusion 500 -861 500 -861 0 feedthrough
rlabel pdiffusion 507 -861 507 -861 0 feedthrough
rlabel pdiffusion 514 -861 514 -861 0 cellNo=747
rlabel pdiffusion 521 -861 521 -861 0 feedthrough
rlabel pdiffusion 528 -861 528 -861 0 feedthrough
rlabel pdiffusion 535 -861 535 -861 0 feedthrough
rlabel pdiffusion 542 -861 542 -861 0 feedthrough
rlabel pdiffusion 549 -861 549 -861 0 cellNo=342
rlabel pdiffusion 556 -861 556 -861 0 cellNo=50
rlabel pdiffusion 563 -861 563 -861 0 feedthrough
rlabel pdiffusion 570 -861 570 -861 0 cellNo=707
rlabel pdiffusion 577 -861 577 -861 0 cellNo=353
rlabel pdiffusion 584 -861 584 -861 0 cellNo=161
rlabel pdiffusion 591 -861 591 -861 0 feedthrough
rlabel pdiffusion 598 -861 598 -861 0 cellNo=259
rlabel pdiffusion 605 -861 605 -861 0 feedthrough
rlabel pdiffusion 612 -861 612 -861 0 cellNo=204
rlabel pdiffusion 619 -861 619 -861 0 cellNo=554
rlabel pdiffusion 626 -861 626 -861 0 cellNo=529
rlabel pdiffusion 633 -861 633 -861 0 feedthrough
rlabel pdiffusion 640 -861 640 -861 0 feedthrough
rlabel pdiffusion 647 -861 647 -861 0 feedthrough
rlabel pdiffusion 654 -861 654 -861 0 feedthrough
rlabel pdiffusion 661 -861 661 -861 0 feedthrough
rlabel pdiffusion 668 -861 668 -861 0 feedthrough
rlabel pdiffusion 675 -861 675 -861 0 feedthrough
rlabel pdiffusion 682 -861 682 -861 0 feedthrough
rlabel pdiffusion 689 -861 689 -861 0 cellNo=99
rlabel pdiffusion 696 -861 696 -861 0 feedthrough
rlabel pdiffusion 703 -861 703 -861 0 cellNo=620
rlabel pdiffusion 710 -861 710 -861 0 feedthrough
rlabel pdiffusion 717 -861 717 -861 0 feedthrough
rlabel pdiffusion 724 -861 724 -861 0 feedthrough
rlabel pdiffusion 731 -861 731 -861 0 feedthrough
rlabel pdiffusion 738 -861 738 -861 0 feedthrough
rlabel pdiffusion 745 -861 745 -861 0 feedthrough
rlabel pdiffusion 752 -861 752 -861 0 feedthrough
rlabel pdiffusion 759 -861 759 -861 0 cellNo=782
rlabel pdiffusion 766 -861 766 -861 0 feedthrough
rlabel pdiffusion 773 -861 773 -861 0 feedthrough
rlabel pdiffusion 780 -861 780 -861 0 cellNo=718
rlabel pdiffusion 787 -861 787 -861 0 cellNo=391
rlabel pdiffusion 794 -861 794 -861 0 feedthrough
rlabel pdiffusion 801 -861 801 -861 0 feedthrough
rlabel pdiffusion 808 -861 808 -861 0 feedthrough
rlabel pdiffusion 815 -861 815 -861 0 feedthrough
rlabel pdiffusion 822 -861 822 -861 0 cellNo=831
rlabel pdiffusion 829 -861 829 -861 0 cellNo=173
rlabel pdiffusion 836 -861 836 -861 0 feedthrough
rlabel pdiffusion 843 -861 843 -861 0 feedthrough
rlabel pdiffusion 850 -861 850 -861 0 feedthrough
rlabel pdiffusion 857 -861 857 -861 0 feedthrough
rlabel pdiffusion 864 -861 864 -861 0 feedthrough
rlabel pdiffusion 871 -861 871 -861 0 feedthrough
rlabel pdiffusion 878 -861 878 -861 0 feedthrough
rlabel pdiffusion 885 -861 885 -861 0 feedthrough
rlabel pdiffusion 892 -861 892 -861 0 feedthrough
rlabel pdiffusion 899 -861 899 -861 0 feedthrough
rlabel pdiffusion 906 -861 906 -861 0 feedthrough
rlabel pdiffusion 913 -861 913 -861 0 feedthrough
rlabel pdiffusion 920 -861 920 -861 0 cellNo=48
rlabel pdiffusion 927 -861 927 -861 0 feedthrough
rlabel pdiffusion 934 -861 934 -861 0 feedthrough
rlabel pdiffusion 941 -861 941 -861 0 feedthrough
rlabel pdiffusion 948 -861 948 -861 0 feedthrough
rlabel pdiffusion 955 -861 955 -861 0 feedthrough
rlabel pdiffusion 962 -861 962 -861 0 feedthrough
rlabel pdiffusion 969 -861 969 -861 0 feedthrough
rlabel pdiffusion 976 -861 976 -861 0 cellNo=474
rlabel pdiffusion 983 -861 983 -861 0 feedthrough
rlabel pdiffusion 990 -861 990 -861 0 feedthrough
rlabel pdiffusion 997 -861 997 -861 0 feedthrough
rlabel pdiffusion 1004 -861 1004 -861 0 feedthrough
rlabel pdiffusion 1011 -861 1011 -861 0 feedthrough
rlabel pdiffusion 1018 -861 1018 -861 0 feedthrough
rlabel pdiffusion 1025 -861 1025 -861 0 feedthrough
rlabel pdiffusion 1032 -861 1032 -861 0 cellNo=592
rlabel pdiffusion 1039 -861 1039 -861 0 feedthrough
rlabel pdiffusion 1046 -861 1046 -861 0 feedthrough
rlabel pdiffusion 1053 -861 1053 -861 0 feedthrough
rlabel pdiffusion 1060 -861 1060 -861 0 feedthrough
rlabel pdiffusion 1067 -861 1067 -861 0 feedthrough
rlabel pdiffusion 1074 -861 1074 -861 0 feedthrough
rlabel pdiffusion 1081 -861 1081 -861 0 feedthrough
rlabel pdiffusion 1088 -861 1088 -861 0 feedthrough
rlabel pdiffusion 1095 -861 1095 -861 0 feedthrough
rlabel pdiffusion 1102 -861 1102 -861 0 feedthrough
rlabel pdiffusion 1109 -861 1109 -861 0 feedthrough
rlabel pdiffusion 1116 -861 1116 -861 0 feedthrough
rlabel pdiffusion 1123 -861 1123 -861 0 feedthrough
rlabel pdiffusion 1130 -861 1130 -861 0 feedthrough
rlabel pdiffusion 1137 -861 1137 -861 0 feedthrough
rlabel pdiffusion 1144 -861 1144 -861 0 feedthrough
rlabel pdiffusion 1151 -861 1151 -861 0 feedthrough
rlabel pdiffusion 1158 -861 1158 -861 0 feedthrough
rlabel pdiffusion 1165 -861 1165 -861 0 feedthrough
rlabel pdiffusion 1172 -861 1172 -861 0 feedthrough
rlabel pdiffusion 1179 -861 1179 -861 0 feedthrough
rlabel pdiffusion 1186 -861 1186 -861 0 feedthrough
rlabel pdiffusion 1193 -861 1193 -861 0 cellNo=876
rlabel pdiffusion 1200 -861 1200 -861 0 feedthrough
rlabel pdiffusion 1207 -861 1207 -861 0 feedthrough
rlabel pdiffusion 1214 -861 1214 -861 0 feedthrough
rlabel pdiffusion 1221 -861 1221 -861 0 feedthrough
rlabel pdiffusion 1228 -861 1228 -861 0 feedthrough
rlabel pdiffusion 1235 -861 1235 -861 0 feedthrough
rlabel pdiffusion 1242 -861 1242 -861 0 feedthrough
rlabel pdiffusion 1249 -861 1249 -861 0 feedthrough
rlabel pdiffusion 1256 -861 1256 -861 0 feedthrough
rlabel pdiffusion 1263 -861 1263 -861 0 feedthrough
rlabel pdiffusion 1270 -861 1270 -861 0 feedthrough
rlabel pdiffusion 1277 -861 1277 -861 0 feedthrough
rlabel pdiffusion 1284 -861 1284 -861 0 feedthrough
rlabel pdiffusion 1291 -861 1291 -861 0 feedthrough
rlabel pdiffusion 1298 -861 1298 -861 0 feedthrough
rlabel pdiffusion 1305 -861 1305 -861 0 feedthrough
rlabel pdiffusion 1312 -861 1312 -861 0 feedthrough
rlabel pdiffusion 1319 -861 1319 -861 0 feedthrough
rlabel pdiffusion 1326 -861 1326 -861 0 feedthrough
rlabel pdiffusion 1333 -861 1333 -861 0 feedthrough
rlabel pdiffusion 1340 -861 1340 -861 0 feedthrough
rlabel pdiffusion 1347 -861 1347 -861 0 feedthrough
rlabel pdiffusion 1354 -861 1354 -861 0 feedthrough
rlabel pdiffusion 1361 -861 1361 -861 0 feedthrough
rlabel pdiffusion 1368 -861 1368 -861 0 feedthrough
rlabel pdiffusion 1375 -861 1375 -861 0 feedthrough
rlabel pdiffusion 1382 -861 1382 -861 0 feedthrough
rlabel pdiffusion 1389 -861 1389 -861 0 feedthrough
rlabel pdiffusion 1396 -861 1396 -861 0 feedthrough
rlabel pdiffusion 1403 -861 1403 -861 0 feedthrough
rlabel pdiffusion 1410 -861 1410 -861 0 feedthrough
rlabel pdiffusion 1417 -861 1417 -861 0 feedthrough
rlabel pdiffusion 1424 -861 1424 -861 0 feedthrough
rlabel pdiffusion 1431 -861 1431 -861 0 feedthrough
rlabel pdiffusion 1438 -861 1438 -861 0 feedthrough
rlabel pdiffusion 1445 -861 1445 -861 0 feedthrough
rlabel pdiffusion 1452 -861 1452 -861 0 feedthrough
rlabel pdiffusion 1459 -861 1459 -861 0 feedthrough
rlabel pdiffusion 1466 -861 1466 -861 0 feedthrough
rlabel pdiffusion 1473 -861 1473 -861 0 feedthrough
rlabel pdiffusion 1480 -861 1480 -861 0 feedthrough
rlabel pdiffusion 1487 -861 1487 -861 0 feedthrough
rlabel pdiffusion 1494 -861 1494 -861 0 feedthrough
rlabel pdiffusion 1501 -861 1501 -861 0 feedthrough
rlabel pdiffusion 1508 -861 1508 -861 0 feedthrough
rlabel pdiffusion 1515 -861 1515 -861 0 feedthrough
rlabel pdiffusion 1522 -861 1522 -861 0 feedthrough
rlabel pdiffusion 1529 -861 1529 -861 0 feedthrough
rlabel pdiffusion 1536 -861 1536 -861 0 feedthrough
rlabel pdiffusion 1543 -861 1543 -861 0 feedthrough
rlabel pdiffusion 1550 -861 1550 -861 0 feedthrough
rlabel pdiffusion 1557 -861 1557 -861 0 feedthrough
rlabel pdiffusion 1564 -861 1564 -861 0 feedthrough
rlabel pdiffusion 1571 -861 1571 -861 0 feedthrough
rlabel pdiffusion 1578 -861 1578 -861 0 feedthrough
rlabel pdiffusion 1585 -861 1585 -861 0 feedthrough
rlabel pdiffusion 1592 -861 1592 -861 0 feedthrough
rlabel pdiffusion 1599 -861 1599 -861 0 feedthrough
rlabel pdiffusion 1606 -861 1606 -861 0 feedthrough
rlabel pdiffusion 1613 -861 1613 -861 0 feedthrough
rlabel pdiffusion 1620 -861 1620 -861 0 feedthrough
rlabel pdiffusion 1627 -861 1627 -861 0 feedthrough
rlabel pdiffusion 1634 -861 1634 -861 0 feedthrough
rlabel pdiffusion 1641 -861 1641 -861 0 feedthrough
rlabel pdiffusion 1648 -861 1648 -861 0 feedthrough
rlabel pdiffusion 1655 -861 1655 -861 0 feedthrough
rlabel pdiffusion 1662 -861 1662 -861 0 feedthrough
rlabel pdiffusion 1669 -861 1669 -861 0 feedthrough
rlabel pdiffusion 1676 -861 1676 -861 0 feedthrough
rlabel pdiffusion 1683 -861 1683 -861 0 feedthrough
rlabel pdiffusion 1690 -861 1690 -861 0 feedthrough
rlabel pdiffusion 1697 -861 1697 -861 0 feedthrough
rlabel pdiffusion 1704 -861 1704 -861 0 feedthrough
rlabel pdiffusion 1711 -861 1711 -861 0 feedthrough
rlabel pdiffusion 1718 -861 1718 -861 0 feedthrough
rlabel pdiffusion 1725 -861 1725 -861 0 feedthrough
rlabel pdiffusion 1732 -861 1732 -861 0 feedthrough
rlabel pdiffusion 1739 -861 1739 -861 0 feedthrough
rlabel pdiffusion 1746 -861 1746 -861 0 feedthrough
rlabel pdiffusion 1753 -861 1753 -861 0 feedthrough
rlabel pdiffusion 1760 -861 1760 -861 0 feedthrough
rlabel pdiffusion 1767 -861 1767 -861 0 feedthrough
rlabel pdiffusion 1774 -861 1774 -861 0 feedthrough
rlabel pdiffusion 1781 -861 1781 -861 0 cellNo=824
rlabel pdiffusion 1788 -861 1788 -861 0 feedthrough
rlabel pdiffusion 1795 -861 1795 -861 0 feedthrough
rlabel pdiffusion 1802 -861 1802 -861 0 feedthrough
rlabel pdiffusion 1809 -861 1809 -861 0 feedthrough
rlabel pdiffusion 1816 -861 1816 -861 0 cellNo=340
rlabel pdiffusion 1823 -861 1823 -861 0 feedthrough
rlabel pdiffusion 1830 -861 1830 -861 0 feedthrough
rlabel pdiffusion 1837 -861 1837 -861 0 feedthrough
rlabel pdiffusion 1844 -861 1844 -861 0 feedthrough
rlabel pdiffusion 1851 -861 1851 -861 0 feedthrough
rlabel pdiffusion 1858 -861 1858 -861 0 feedthrough
rlabel pdiffusion 1886 -861 1886 -861 0 feedthrough
rlabel pdiffusion 1893 -861 1893 -861 0 feedthrough
rlabel pdiffusion 3 -982 3 -982 0 feedthrough
rlabel pdiffusion 10 -982 10 -982 0 feedthrough
rlabel pdiffusion 17 -982 17 -982 0 feedthrough
rlabel pdiffusion 24 -982 24 -982 0 feedthrough
rlabel pdiffusion 31 -982 31 -982 0 feedthrough
rlabel pdiffusion 38 -982 38 -982 0 feedthrough
rlabel pdiffusion 45 -982 45 -982 0 feedthrough
rlabel pdiffusion 52 -982 52 -982 0 feedthrough
rlabel pdiffusion 59 -982 59 -982 0 feedthrough
rlabel pdiffusion 66 -982 66 -982 0 cellNo=860
rlabel pdiffusion 73 -982 73 -982 0 feedthrough
rlabel pdiffusion 80 -982 80 -982 0 feedthrough
rlabel pdiffusion 87 -982 87 -982 0 feedthrough
rlabel pdiffusion 94 -982 94 -982 0 cellNo=514
rlabel pdiffusion 101 -982 101 -982 0 feedthrough
rlabel pdiffusion 108 -982 108 -982 0 cellNo=763
rlabel pdiffusion 115 -982 115 -982 0 feedthrough
rlabel pdiffusion 122 -982 122 -982 0 feedthrough
rlabel pdiffusion 129 -982 129 -982 0 feedthrough
rlabel pdiffusion 136 -982 136 -982 0 feedthrough
rlabel pdiffusion 143 -982 143 -982 0 cellNo=406
rlabel pdiffusion 150 -982 150 -982 0 feedthrough
rlabel pdiffusion 157 -982 157 -982 0 cellNo=287
rlabel pdiffusion 164 -982 164 -982 0 feedthrough
rlabel pdiffusion 171 -982 171 -982 0 feedthrough
rlabel pdiffusion 178 -982 178 -982 0 feedthrough
rlabel pdiffusion 185 -982 185 -982 0 cellNo=122
rlabel pdiffusion 192 -982 192 -982 0 feedthrough
rlabel pdiffusion 199 -982 199 -982 0 feedthrough
rlabel pdiffusion 206 -982 206 -982 0 feedthrough
rlabel pdiffusion 213 -982 213 -982 0 feedthrough
rlabel pdiffusion 220 -982 220 -982 0 feedthrough
rlabel pdiffusion 227 -982 227 -982 0 feedthrough
rlabel pdiffusion 234 -982 234 -982 0 cellNo=607
rlabel pdiffusion 241 -982 241 -982 0 feedthrough
rlabel pdiffusion 248 -982 248 -982 0 feedthrough
rlabel pdiffusion 255 -982 255 -982 0 feedthrough
rlabel pdiffusion 262 -982 262 -982 0 feedthrough
rlabel pdiffusion 269 -982 269 -982 0 feedthrough
rlabel pdiffusion 276 -982 276 -982 0 feedthrough
rlabel pdiffusion 283 -982 283 -982 0 feedthrough
rlabel pdiffusion 290 -982 290 -982 0 feedthrough
rlabel pdiffusion 297 -982 297 -982 0 feedthrough
rlabel pdiffusion 304 -982 304 -982 0 feedthrough
rlabel pdiffusion 311 -982 311 -982 0 feedthrough
rlabel pdiffusion 318 -982 318 -982 0 feedthrough
rlabel pdiffusion 325 -982 325 -982 0 feedthrough
rlabel pdiffusion 332 -982 332 -982 0 feedthrough
rlabel pdiffusion 339 -982 339 -982 0 feedthrough
rlabel pdiffusion 346 -982 346 -982 0 feedthrough
rlabel pdiffusion 353 -982 353 -982 0 feedthrough
rlabel pdiffusion 360 -982 360 -982 0 feedthrough
rlabel pdiffusion 367 -982 367 -982 0 feedthrough
rlabel pdiffusion 374 -982 374 -982 0 feedthrough
rlabel pdiffusion 381 -982 381 -982 0 feedthrough
rlabel pdiffusion 388 -982 388 -982 0 cellNo=451
rlabel pdiffusion 395 -982 395 -982 0 feedthrough
rlabel pdiffusion 402 -982 402 -982 0 feedthrough
rlabel pdiffusion 409 -982 409 -982 0 feedthrough
rlabel pdiffusion 416 -982 416 -982 0 feedthrough
rlabel pdiffusion 423 -982 423 -982 0 feedthrough
rlabel pdiffusion 430 -982 430 -982 0 feedthrough
rlabel pdiffusion 437 -982 437 -982 0 feedthrough
rlabel pdiffusion 444 -982 444 -982 0 feedthrough
rlabel pdiffusion 451 -982 451 -982 0 feedthrough
rlabel pdiffusion 458 -982 458 -982 0 cellNo=715
rlabel pdiffusion 465 -982 465 -982 0 feedthrough
rlabel pdiffusion 472 -982 472 -982 0 feedthrough
rlabel pdiffusion 479 -982 479 -982 0 feedthrough
rlabel pdiffusion 486 -982 486 -982 0 feedthrough
rlabel pdiffusion 493 -982 493 -982 0 feedthrough
rlabel pdiffusion 500 -982 500 -982 0 feedthrough
rlabel pdiffusion 507 -982 507 -982 0 feedthrough
rlabel pdiffusion 514 -982 514 -982 0 feedthrough
rlabel pdiffusion 521 -982 521 -982 0 feedthrough
rlabel pdiffusion 528 -982 528 -982 0 feedthrough
rlabel pdiffusion 535 -982 535 -982 0 cellNo=246
rlabel pdiffusion 542 -982 542 -982 0 cellNo=412
rlabel pdiffusion 549 -982 549 -982 0 feedthrough
rlabel pdiffusion 556 -982 556 -982 0 feedthrough
rlabel pdiffusion 563 -982 563 -982 0 feedthrough
rlabel pdiffusion 570 -982 570 -982 0 feedthrough
rlabel pdiffusion 577 -982 577 -982 0 feedthrough
rlabel pdiffusion 584 -982 584 -982 0 feedthrough
rlabel pdiffusion 591 -982 591 -982 0 feedthrough
rlabel pdiffusion 598 -982 598 -982 0 feedthrough
rlabel pdiffusion 605 -982 605 -982 0 cellNo=157
rlabel pdiffusion 612 -982 612 -982 0 feedthrough
rlabel pdiffusion 619 -982 619 -982 0 feedthrough
rlabel pdiffusion 626 -982 626 -982 0 feedthrough
rlabel pdiffusion 633 -982 633 -982 0 feedthrough
rlabel pdiffusion 640 -982 640 -982 0 feedthrough
rlabel pdiffusion 647 -982 647 -982 0 feedthrough
rlabel pdiffusion 654 -982 654 -982 0 feedthrough
rlabel pdiffusion 661 -982 661 -982 0 feedthrough
rlabel pdiffusion 668 -982 668 -982 0 feedthrough
rlabel pdiffusion 675 -982 675 -982 0 feedthrough
rlabel pdiffusion 682 -982 682 -982 0 cellNo=167
rlabel pdiffusion 689 -982 689 -982 0 feedthrough
rlabel pdiffusion 696 -982 696 -982 0 feedthrough
rlabel pdiffusion 703 -982 703 -982 0 feedthrough
rlabel pdiffusion 710 -982 710 -982 0 feedthrough
rlabel pdiffusion 717 -982 717 -982 0 feedthrough
rlabel pdiffusion 724 -982 724 -982 0 cellNo=659
rlabel pdiffusion 731 -982 731 -982 0 feedthrough
rlabel pdiffusion 738 -982 738 -982 0 cellNo=258
rlabel pdiffusion 745 -982 745 -982 0 cellNo=299
rlabel pdiffusion 752 -982 752 -982 0 cellNo=383
rlabel pdiffusion 759 -982 759 -982 0 feedthrough
rlabel pdiffusion 766 -982 766 -982 0 feedthrough
rlabel pdiffusion 773 -982 773 -982 0 cellNo=170
rlabel pdiffusion 780 -982 780 -982 0 feedthrough
rlabel pdiffusion 787 -982 787 -982 0 feedthrough
rlabel pdiffusion 794 -982 794 -982 0 feedthrough
rlabel pdiffusion 801 -982 801 -982 0 feedthrough
rlabel pdiffusion 808 -982 808 -982 0 feedthrough
rlabel pdiffusion 815 -982 815 -982 0 feedthrough
rlabel pdiffusion 822 -982 822 -982 0 feedthrough
rlabel pdiffusion 829 -982 829 -982 0 feedthrough
rlabel pdiffusion 836 -982 836 -982 0 feedthrough
rlabel pdiffusion 843 -982 843 -982 0 feedthrough
rlabel pdiffusion 850 -982 850 -982 0 feedthrough
rlabel pdiffusion 857 -982 857 -982 0 feedthrough
rlabel pdiffusion 864 -982 864 -982 0 feedthrough
rlabel pdiffusion 871 -982 871 -982 0 feedthrough
rlabel pdiffusion 878 -982 878 -982 0 feedthrough
rlabel pdiffusion 885 -982 885 -982 0 feedthrough
rlabel pdiffusion 892 -982 892 -982 0 feedthrough
rlabel pdiffusion 899 -982 899 -982 0 feedthrough
rlabel pdiffusion 906 -982 906 -982 0 feedthrough
rlabel pdiffusion 913 -982 913 -982 0 cellNo=538
rlabel pdiffusion 920 -982 920 -982 0 cellNo=815
rlabel pdiffusion 927 -982 927 -982 0 feedthrough
rlabel pdiffusion 934 -982 934 -982 0 feedthrough
rlabel pdiffusion 941 -982 941 -982 0 cellNo=89
rlabel pdiffusion 948 -982 948 -982 0 feedthrough
rlabel pdiffusion 955 -982 955 -982 0 feedthrough
rlabel pdiffusion 962 -982 962 -982 0 feedthrough
rlabel pdiffusion 969 -982 969 -982 0 feedthrough
rlabel pdiffusion 976 -982 976 -982 0 feedthrough
rlabel pdiffusion 983 -982 983 -982 0 cellNo=382
rlabel pdiffusion 990 -982 990 -982 0 feedthrough
rlabel pdiffusion 997 -982 997 -982 0 feedthrough
rlabel pdiffusion 1004 -982 1004 -982 0 cellNo=565
rlabel pdiffusion 1011 -982 1011 -982 0 cellNo=148
rlabel pdiffusion 1018 -982 1018 -982 0 feedthrough
rlabel pdiffusion 1025 -982 1025 -982 0 feedthrough
rlabel pdiffusion 1032 -982 1032 -982 0 cellNo=329
rlabel pdiffusion 1039 -982 1039 -982 0 cellNo=175
rlabel pdiffusion 1046 -982 1046 -982 0 feedthrough
rlabel pdiffusion 1053 -982 1053 -982 0 feedthrough
rlabel pdiffusion 1060 -982 1060 -982 0 cellNo=783
rlabel pdiffusion 1067 -982 1067 -982 0 feedthrough
rlabel pdiffusion 1074 -982 1074 -982 0 feedthrough
rlabel pdiffusion 1081 -982 1081 -982 0 cellNo=845
rlabel pdiffusion 1088 -982 1088 -982 0 feedthrough
rlabel pdiffusion 1095 -982 1095 -982 0 feedthrough
rlabel pdiffusion 1102 -982 1102 -982 0 feedthrough
rlabel pdiffusion 1109 -982 1109 -982 0 feedthrough
rlabel pdiffusion 1116 -982 1116 -982 0 feedthrough
rlabel pdiffusion 1123 -982 1123 -982 0 feedthrough
rlabel pdiffusion 1130 -982 1130 -982 0 feedthrough
rlabel pdiffusion 1137 -982 1137 -982 0 feedthrough
rlabel pdiffusion 1144 -982 1144 -982 0 feedthrough
rlabel pdiffusion 1151 -982 1151 -982 0 cellNo=685
rlabel pdiffusion 1158 -982 1158 -982 0 cellNo=755
rlabel pdiffusion 1165 -982 1165 -982 0 feedthrough
rlabel pdiffusion 1172 -982 1172 -982 0 feedthrough
rlabel pdiffusion 1179 -982 1179 -982 0 feedthrough
rlabel pdiffusion 1186 -982 1186 -982 0 feedthrough
rlabel pdiffusion 1193 -982 1193 -982 0 feedthrough
rlabel pdiffusion 1200 -982 1200 -982 0 feedthrough
rlabel pdiffusion 1207 -982 1207 -982 0 feedthrough
rlabel pdiffusion 1214 -982 1214 -982 0 feedthrough
rlabel pdiffusion 1221 -982 1221 -982 0 feedthrough
rlabel pdiffusion 1228 -982 1228 -982 0 cellNo=109
rlabel pdiffusion 1235 -982 1235 -982 0 feedthrough
rlabel pdiffusion 1242 -982 1242 -982 0 feedthrough
rlabel pdiffusion 1249 -982 1249 -982 0 feedthrough
rlabel pdiffusion 1256 -982 1256 -982 0 feedthrough
rlabel pdiffusion 1263 -982 1263 -982 0 feedthrough
rlabel pdiffusion 1270 -982 1270 -982 0 feedthrough
rlabel pdiffusion 1277 -982 1277 -982 0 feedthrough
rlabel pdiffusion 1284 -982 1284 -982 0 feedthrough
rlabel pdiffusion 1291 -982 1291 -982 0 feedthrough
rlabel pdiffusion 1298 -982 1298 -982 0 feedthrough
rlabel pdiffusion 1305 -982 1305 -982 0 feedthrough
rlabel pdiffusion 1312 -982 1312 -982 0 feedthrough
rlabel pdiffusion 1319 -982 1319 -982 0 feedthrough
rlabel pdiffusion 1326 -982 1326 -982 0 feedthrough
rlabel pdiffusion 1333 -982 1333 -982 0 feedthrough
rlabel pdiffusion 1340 -982 1340 -982 0 feedthrough
rlabel pdiffusion 1347 -982 1347 -982 0 feedthrough
rlabel pdiffusion 1354 -982 1354 -982 0 feedthrough
rlabel pdiffusion 1361 -982 1361 -982 0 feedthrough
rlabel pdiffusion 1368 -982 1368 -982 0 feedthrough
rlabel pdiffusion 1375 -982 1375 -982 0 feedthrough
rlabel pdiffusion 1382 -982 1382 -982 0 feedthrough
rlabel pdiffusion 1389 -982 1389 -982 0 feedthrough
rlabel pdiffusion 1396 -982 1396 -982 0 feedthrough
rlabel pdiffusion 1403 -982 1403 -982 0 feedthrough
rlabel pdiffusion 1410 -982 1410 -982 0 feedthrough
rlabel pdiffusion 1417 -982 1417 -982 0 feedthrough
rlabel pdiffusion 1424 -982 1424 -982 0 feedthrough
rlabel pdiffusion 1431 -982 1431 -982 0 feedthrough
rlabel pdiffusion 1438 -982 1438 -982 0 feedthrough
rlabel pdiffusion 1445 -982 1445 -982 0 feedthrough
rlabel pdiffusion 1452 -982 1452 -982 0 feedthrough
rlabel pdiffusion 1459 -982 1459 -982 0 feedthrough
rlabel pdiffusion 1466 -982 1466 -982 0 feedthrough
rlabel pdiffusion 1473 -982 1473 -982 0 feedthrough
rlabel pdiffusion 1480 -982 1480 -982 0 feedthrough
rlabel pdiffusion 1487 -982 1487 -982 0 feedthrough
rlabel pdiffusion 1494 -982 1494 -982 0 feedthrough
rlabel pdiffusion 1501 -982 1501 -982 0 feedthrough
rlabel pdiffusion 1508 -982 1508 -982 0 feedthrough
rlabel pdiffusion 1515 -982 1515 -982 0 feedthrough
rlabel pdiffusion 1522 -982 1522 -982 0 feedthrough
rlabel pdiffusion 1529 -982 1529 -982 0 feedthrough
rlabel pdiffusion 1536 -982 1536 -982 0 feedthrough
rlabel pdiffusion 1543 -982 1543 -982 0 feedthrough
rlabel pdiffusion 1550 -982 1550 -982 0 feedthrough
rlabel pdiffusion 1557 -982 1557 -982 0 feedthrough
rlabel pdiffusion 1564 -982 1564 -982 0 feedthrough
rlabel pdiffusion 1571 -982 1571 -982 0 feedthrough
rlabel pdiffusion 1578 -982 1578 -982 0 feedthrough
rlabel pdiffusion 1585 -982 1585 -982 0 feedthrough
rlabel pdiffusion 1592 -982 1592 -982 0 feedthrough
rlabel pdiffusion 1599 -982 1599 -982 0 feedthrough
rlabel pdiffusion 1606 -982 1606 -982 0 feedthrough
rlabel pdiffusion 1613 -982 1613 -982 0 feedthrough
rlabel pdiffusion 1620 -982 1620 -982 0 feedthrough
rlabel pdiffusion 1627 -982 1627 -982 0 feedthrough
rlabel pdiffusion 1634 -982 1634 -982 0 feedthrough
rlabel pdiffusion 1641 -982 1641 -982 0 feedthrough
rlabel pdiffusion 1648 -982 1648 -982 0 feedthrough
rlabel pdiffusion 1655 -982 1655 -982 0 feedthrough
rlabel pdiffusion 1662 -982 1662 -982 0 feedthrough
rlabel pdiffusion 1669 -982 1669 -982 0 feedthrough
rlabel pdiffusion 1676 -982 1676 -982 0 feedthrough
rlabel pdiffusion 1683 -982 1683 -982 0 feedthrough
rlabel pdiffusion 1690 -982 1690 -982 0 feedthrough
rlabel pdiffusion 1697 -982 1697 -982 0 feedthrough
rlabel pdiffusion 1704 -982 1704 -982 0 feedthrough
rlabel pdiffusion 1711 -982 1711 -982 0 feedthrough
rlabel pdiffusion 1718 -982 1718 -982 0 feedthrough
rlabel pdiffusion 1725 -982 1725 -982 0 feedthrough
rlabel pdiffusion 1732 -982 1732 -982 0 feedthrough
rlabel pdiffusion 1739 -982 1739 -982 0 feedthrough
rlabel pdiffusion 1746 -982 1746 -982 0 feedthrough
rlabel pdiffusion 1753 -982 1753 -982 0 feedthrough
rlabel pdiffusion 1760 -982 1760 -982 0 feedthrough
rlabel pdiffusion 1767 -982 1767 -982 0 feedthrough
rlabel pdiffusion 1774 -982 1774 -982 0 feedthrough
rlabel pdiffusion 1781 -982 1781 -982 0 feedthrough
rlabel pdiffusion 1788 -982 1788 -982 0 feedthrough
rlabel pdiffusion 1795 -982 1795 -982 0 feedthrough
rlabel pdiffusion 1802 -982 1802 -982 0 feedthrough
rlabel pdiffusion 1809 -982 1809 -982 0 feedthrough
rlabel pdiffusion 1816 -982 1816 -982 0 feedthrough
rlabel pdiffusion 1823 -982 1823 -982 0 feedthrough
rlabel pdiffusion 1830 -982 1830 -982 0 feedthrough
rlabel pdiffusion 1837 -982 1837 -982 0 feedthrough
rlabel pdiffusion 1844 -982 1844 -982 0 feedthrough
rlabel pdiffusion 1851 -982 1851 -982 0 feedthrough
rlabel pdiffusion 1858 -982 1858 -982 0 feedthrough
rlabel pdiffusion 1865 -982 1865 -982 0 feedthrough
rlabel pdiffusion 1872 -982 1872 -982 0 feedthrough
rlabel pdiffusion 1879 -982 1879 -982 0 cellNo=279
rlabel pdiffusion 1886 -982 1886 -982 0 feedthrough
rlabel pdiffusion 1893 -982 1893 -982 0 feedthrough
rlabel pdiffusion 1900 -982 1900 -982 0 cellNo=377
rlabel pdiffusion 1907 -982 1907 -982 0 feedthrough
rlabel pdiffusion 1914 -982 1914 -982 0 cellNo=679
rlabel pdiffusion 1921 -982 1921 -982 0 cellNo=568
rlabel pdiffusion 1928 -982 1928 -982 0 feedthrough
rlabel pdiffusion 1935 -982 1935 -982 0 feedthrough
rlabel pdiffusion 1942 -982 1942 -982 0 feedthrough
rlabel pdiffusion 1949 -982 1949 -982 0 feedthrough
rlabel pdiffusion 1956 -982 1956 -982 0 feedthrough
rlabel pdiffusion 3 -1113 3 -1113 0 cellNo=1023
rlabel pdiffusion 10 -1113 10 -1113 0 feedthrough
rlabel pdiffusion 17 -1113 17 -1113 0 feedthrough
rlabel pdiffusion 24 -1113 24 -1113 0 feedthrough
rlabel pdiffusion 31 -1113 31 -1113 0 feedthrough
rlabel pdiffusion 38 -1113 38 -1113 0 feedthrough
rlabel pdiffusion 45 -1113 45 -1113 0 cellNo=120
rlabel pdiffusion 52 -1113 52 -1113 0 feedthrough
rlabel pdiffusion 59 -1113 59 -1113 0 feedthrough
rlabel pdiffusion 66 -1113 66 -1113 0 cellNo=252
rlabel pdiffusion 73 -1113 73 -1113 0 feedthrough
rlabel pdiffusion 80 -1113 80 -1113 0 cellNo=319
rlabel pdiffusion 87 -1113 87 -1113 0 feedthrough
rlabel pdiffusion 94 -1113 94 -1113 0 feedthrough
rlabel pdiffusion 101 -1113 101 -1113 0 feedthrough
rlabel pdiffusion 108 -1113 108 -1113 0 feedthrough
rlabel pdiffusion 115 -1113 115 -1113 0 feedthrough
rlabel pdiffusion 122 -1113 122 -1113 0 feedthrough
rlabel pdiffusion 129 -1113 129 -1113 0 cellNo=21
rlabel pdiffusion 136 -1113 136 -1113 0 feedthrough
rlabel pdiffusion 143 -1113 143 -1113 0 feedthrough
rlabel pdiffusion 150 -1113 150 -1113 0 feedthrough
rlabel pdiffusion 157 -1113 157 -1113 0 feedthrough
rlabel pdiffusion 164 -1113 164 -1113 0 feedthrough
rlabel pdiffusion 171 -1113 171 -1113 0 feedthrough
rlabel pdiffusion 178 -1113 178 -1113 0 feedthrough
rlabel pdiffusion 185 -1113 185 -1113 0 feedthrough
rlabel pdiffusion 192 -1113 192 -1113 0 feedthrough
rlabel pdiffusion 199 -1113 199 -1113 0 feedthrough
rlabel pdiffusion 206 -1113 206 -1113 0 feedthrough
rlabel pdiffusion 213 -1113 213 -1113 0 cellNo=683
rlabel pdiffusion 220 -1113 220 -1113 0 cellNo=438
rlabel pdiffusion 227 -1113 227 -1113 0 feedthrough
rlabel pdiffusion 234 -1113 234 -1113 0 feedthrough
rlabel pdiffusion 241 -1113 241 -1113 0 feedthrough
rlabel pdiffusion 248 -1113 248 -1113 0 feedthrough
rlabel pdiffusion 255 -1113 255 -1113 0 feedthrough
rlabel pdiffusion 262 -1113 262 -1113 0 feedthrough
rlabel pdiffusion 269 -1113 269 -1113 0 feedthrough
rlabel pdiffusion 276 -1113 276 -1113 0 feedthrough
rlabel pdiffusion 283 -1113 283 -1113 0 feedthrough
rlabel pdiffusion 290 -1113 290 -1113 0 feedthrough
rlabel pdiffusion 297 -1113 297 -1113 0 feedthrough
rlabel pdiffusion 304 -1113 304 -1113 0 feedthrough
rlabel pdiffusion 311 -1113 311 -1113 0 cellNo=708
rlabel pdiffusion 318 -1113 318 -1113 0 feedthrough
rlabel pdiffusion 325 -1113 325 -1113 0 feedthrough
rlabel pdiffusion 332 -1113 332 -1113 0 feedthrough
rlabel pdiffusion 339 -1113 339 -1113 0 feedthrough
rlabel pdiffusion 346 -1113 346 -1113 0 feedthrough
rlabel pdiffusion 353 -1113 353 -1113 0 feedthrough
rlabel pdiffusion 360 -1113 360 -1113 0 feedthrough
rlabel pdiffusion 367 -1113 367 -1113 0 feedthrough
rlabel pdiffusion 374 -1113 374 -1113 0 feedthrough
rlabel pdiffusion 381 -1113 381 -1113 0 feedthrough
rlabel pdiffusion 388 -1113 388 -1113 0 feedthrough
rlabel pdiffusion 395 -1113 395 -1113 0 cellNo=293
rlabel pdiffusion 402 -1113 402 -1113 0 feedthrough
rlabel pdiffusion 409 -1113 409 -1113 0 feedthrough
rlabel pdiffusion 416 -1113 416 -1113 0 feedthrough
rlabel pdiffusion 423 -1113 423 -1113 0 feedthrough
rlabel pdiffusion 430 -1113 430 -1113 0 feedthrough
rlabel pdiffusion 437 -1113 437 -1113 0 feedthrough
rlabel pdiffusion 444 -1113 444 -1113 0 feedthrough
rlabel pdiffusion 451 -1113 451 -1113 0 cellNo=225
rlabel pdiffusion 458 -1113 458 -1113 0 feedthrough
rlabel pdiffusion 465 -1113 465 -1113 0 feedthrough
rlabel pdiffusion 472 -1113 472 -1113 0 feedthrough
rlabel pdiffusion 479 -1113 479 -1113 0 feedthrough
rlabel pdiffusion 486 -1113 486 -1113 0 feedthrough
rlabel pdiffusion 493 -1113 493 -1113 0 feedthrough
rlabel pdiffusion 500 -1113 500 -1113 0 feedthrough
rlabel pdiffusion 507 -1113 507 -1113 0 feedthrough
rlabel pdiffusion 514 -1113 514 -1113 0 feedthrough
rlabel pdiffusion 521 -1113 521 -1113 0 cellNo=791
rlabel pdiffusion 528 -1113 528 -1113 0 feedthrough
rlabel pdiffusion 535 -1113 535 -1113 0 feedthrough
rlabel pdiffusion 542 -1113 542 -1113 0 feedthrough
rlabel pdiffusion 549 -1113 549 -1113 0 feedthrough
rlabel pdiffusion 556 -1113 556 -1113 0 feedthrough
rlabel pdiffusion 563 -1113 563 -1113 0 cellNo=525
rlabel pdiffusion 570 -1113 570 -1113 0 cellNo=735
rlabel pdiffusion 577 -1113 577 -1113 0 cellNo=239
rlabel pdiffusion 584 -1113 584 -1113 0 feedthrough
rlabel pdiffusion 591 -1113 591 -1113 0 feedthrough
rlabel pdiffusion 598 -1113 598 -1113 0 feedthrough
rlabel pdiffusion 605 -1113 605 -1113 0 feedthrough
rlabel pdiffusion 612 -1113 612 -1113 0 feedthrough
rlabel pdiffusion 619 -1113 619 -1113 0 feedthrough
rlabel pdiffusion 626 -1113 626 -1113 0 cellNo=240
rlabel pdiffusion 633 -1113 633 -1113 0 cellNo=88
rlabel pdiffusion 640 -1113 640 -1113 0 feedthrough
rlabel pdiffusion 647 -1113 647 -1113 0 cellNo=197
rlabel pdiffusion 654 -1113 654 -1113 0 cellNo=666
rlabel pdiffusion 661 -1113 661 -1113 0 feedthrough
rlabel pdiffusion 668 -1113 668 -1113 0 feedthrough
rlabel pdiffusion 675 -1113 675 -1113 0 feedthrough
rlabel pdiffusion 682 -1113 682 -1113 0 cellNo=216
rlabel pdiffusion 689 -1113 689 -1113 0 feedthrough
rlabel pdiffusion 696 -1113 696 -1113 0 feedthrough
rlabel pdiffusion 703 -1113 703 -1113 0 feedthrough
rlabel pdiffusion 710 -1113 710 -1113 0 feedthrough
rlabel pdiffusion 717 -1113 717 -1113 0 feedthrough
rlabel pdiffusion 724 -1113 724 -1113 0 feedthrough
rlabel pdiffusion 731 -1113 731 -1113 0 cellNo=786
rlabel pdiffusion 738 -1113 738 -1113 0 cellNo=494
rlabel pdiffusion 745 -1113 745 -1113 0 feedthrough
rlabel pdiffusion 752 -1113 752 -1113 0 cellNo=39
rlabel pdiffusion 759 -1113 759 -1113 0 cellNo=250
rlabel pdiffusion 766 -1113 766 -1113 0 feedthrough
rlabel pdiffusion 773 -1113 773 -1113 0 feedthrough
rlabel pdiffusion 780 -1113 780 -1113 0 cellNo=433
rlabel pdiffusion 787 -1113 787 -1113 0 cellNo=905
rlabel pdiffusion 794 -1113 794 -1113 0 feedthrough
rlabel pdiffusion 801 -1113 801 -1113 0 feedthrough
rlabel pdiffusion 808 -1113 808 -1113 0 feedthrough
rlabel pdiffusion 815 -1113 815 -1113 0 feedthrough
rlabel pdiffusion 822 -1113 822 -1113 0 feedthrough
rlabel pdiffusion 829 -1113 829 -1113 0 feedthrough
rlabel pdiffusion 836 -1113 836 -1113 0 feedthrough
rlabel pdiffusion 843 -1113 843 -1113 0 feedthrough
rlabel pdiffusion 850 -1113 850 -1113 0 cellNo=902
rlabel pdiffusion 857 -1113 857 -1113 0 feedthrough
rlabel pdiffusion 864 -1113 864 -1113 0 cellNo=183
rlabel pdiffusion 871 -1113 871 -1113 0 feedthrough
rlabel pdiffusion 878 -1113 878 -1113 0 feedthrough
rlabel pdiffusion 885 -1113 885 -1113 0 feedthrough
rlabel pdiffusion 892 -1113 892 -1113 0 cellNo=479
rlabel pdiffusion 899 -1113 899 -1113 0 feedthrough
rlabel pdiffusion 906 -1113 906 -1113 0 feedthrough
rlabel pdiffusion 913 -1113 913 -1113 0 feedthrough
rlabel pdiffusion 920 -1113 920 -1113 0 feedthrough
rlabel pdiffusion 927 -1113 927 -1113 0 feedthrough
rlabel pdiffusion 934 -1113 934 -1113 0 feedthrough
rlabel pdiffusion 941 -1113 941 -1113 0 feedthrough
rlabel pdiffusion 948 -1113 948 -1113 0 feedthrough
rlabel pdiffusion 955 -1113 955 -1113 0 cellNo=454
rlabel pdiffusion 962 -1113 962 -1113 0 feedthrough
rlabel pdiffusion 969 -1113 969 -1113 0 feedthrough
rlabel pdiffusion 976 -1113 976 -1113 0 feedthrough
rlabel pdiffusion 983 -1113 983 -1113 0 feedthrough
rlabel pdiffusion 990 -1113 990 -1113 0 feedthrough
rlabel pdiffusion 997 -1113 997 -1113 0 feedthrough
rlabel pdiffusion 1004 -1113 1004 -1113 0 feedthrough
rlabel pdiffusion 1011 -1113 1011 -1113 0 feedthrough
rlabel pdiffusion 1018 -1113 1018 -1113 0 cellNo=367
rlabel pdiffusion 1025 -1113 1025 -1113 0 feedthrough
rlabel pdiffusion 1032 -1113 1032 -1113 0 feedthrough
rlabel pdiffusion 1039 -1113 1039 -1113 0 feedthrough
rlabel pdiffusion 1046 -1113 1046 -1113 0 cellNo=346
rlabel pdiffusion 1053 -1113 1053 -1113 0 feedthrough
rlabel pdiffusion 1060 -1113 1060 -1113 0 feedthrough
rlabel pdiffusion 1067 -1113 1067 -1113 0 feedthrough
rlabel pdiffusion 1074 -1113 1074 -1113 0 feedthrough
rlabel pdiffusion 1081 -1113 1081 -1113 0 feedthrough
rlabel pdiffusion 1088 -1113 1088 -1113 0 feedthrough
rlabel pdiffusion 1095 -1113 1095 -1113 0 feedthrough
rlabel pdiffusion 1102 -1113 1102 -1113 0 feedthrough
rlabel pdiffusion 1109 -1113 1109 -1113 0 feedthrough
rlabel pdiffusion 1116 -1113 1116 -1113 0 feedthrough
rlabel pdiffusion 1123 -1113 1123 -1113 0 feedthrough
rlabel pdiffusion 1130 -1113 1130 -1113 0 feedthrough
rlabel pdiffusion 1137 -1113 1137 -1113 0 cellNo=865
rlabel pdiffusion 1144 -1113 1144 -1113 0 feedthrough
rlabel pdiffusion 1151 -1113 1151 -1113 0 cellNo=219
rlabel pdiffusion 1158 -1113 1158 -1113 0 feedthrough
rlabel pdiffusion 1165 -1113 1165 -1113 0 feedthrough
rlabel pdiffusion 1172 -1113 1172 -1113 0 feedthrough
rlabel pdiffusion 1179 -1113 1179 -1113 0 feedthrough
rlabel pdiffusion 1186 -1113 1186 -1113 0 feedthrough
rlabel pdiffusion 1193 -1113 1193 -1113 0 feedthrough
rlabel pdiffusion 1200 -1113 1200 -1113 0 feedthrough
rlabel pdiffusion 1207 -1113 1207 -1113 0 feedthrough
rlabel pdiffusion 1214 -1113 1214 -1113 0 feedthrough
rlabel pdiffusion 1221 -1113 1221 -1113 0 feedthrough
rlabel pdiffusion 1228 -1113 1228 -1113 0 cellNo=244
rlabel pdiffusion 1235 -1113 1235 -1113 0 feedthrough
rlabel pdiffusion 1242 -1113 1242 -1113 0 feedthrough
rlabel pdiffusion 1249 -1113 1249 -1113 0 feedthrough
rlabel pdiffusion 1256 -1113 1256 -1113 0 feedthrough
rlabel pdiffusion 1263 -1113 1263 -1113 0 feedthrough
rlabel pdiffusion 1270 -1113 1270 -1113 0 feedthrough
rlabel pdiffusion 1277 -1113 1277 -1113 0 feedthrough
rlabel pdiffusion 1284 -1113 1284 -1113 0 feedthrough
rlabel pdiffusion 1291 -1113 1291 -1113 0 feedthrough
rlabel pdiffusion 1298 -1113 1298 -1113 0 feedthrough
rlabel pdiffusion 1305 -1113 1305 -1113 0 feedthrough
rlabel pdiffusion 1312 -1113 1312 -1113 0 feedthrough
rlabel pdiffusion 1319 -1113 1319 -1113 0 feedthrough
rlabel pdiffusion 1326 -1113 1326 -1113 0 feedthrough
rlabel pdiffusion 1333 -1113 1333 -1113 0 feedthrough
rlabel pdiffusion 1340 -1113 1340 -1113 0 feedthrough
rlabel pdiffusion 1347 -1113 1347 -1113 0 feedthrough
rlabel pdiffusion 1354 -1113 1354 -1113 0 feedthrough
rlabel pdiffusion 1361 -1113 1361 -1113 0 feedthrough
rlabel pdiffusion 1368 -1113 1368 -1113 0 feedthrough
rlabel pdiffusion 1375 -1113 1375 -1113 0 feedthrough
rlabel pdiffusion 1382 -1113 1382 -1113 0 feedthrough
rlabel pdiffusion 1389 -1113 1389 -1113 0 feedthrough
rlabel pdiffusion 1396 -1113 1396 -1113 0 feedthrough
rlabel pdiffusion 1403 -1113 1403 -1113 0 feedthrough
rlabel pdiffusion 1410 -1113 1410 -1113 0 feedthrough
rlabel pdiffusion 1417 -1113 1417 -1113 0 feedthrough
rlabel pdiffusion 1424 -1113 1424 -1113 0 feedthrough
rlabel pdiffusion 1431 -1113 1431 -1113 0 feedthrough
rlabel pdiffusion 1438 -1113 1438 -1113 0 feedthrough
rlabel pdiffusion 1445 -1113 1445 -1113 0 feedthrough
rlabel pdiffusion 1452 -1113 1452 -1113 0 feedthrough
rlabel pdiffusion 1459 -1113 1459 -1113 0 feedthrough
rlabel pdiffusion 1466 -1113 1466 -1113 0 feedthrough
rlabel pdiffusion 1473 -1113 1473 -1113 0 feedthrough
rlabel pdiffusion 1480 -1113 1480 -1113 0 feedthrough
rlabel pdiffusion 1487 -1113 1487 -1113 0 feedthrough
rlabel pdiffusion 1494 -1113 1494 -1113 0 feedthrough
rlabel pdiffusion 1501 -1113 1501 -1113 0 feedthrough
rlabel pdiffusion 1508 -1113 1508 -1113 0 feedthrough
rlabel pdiffusion 1515 -1113 1515 -1113 0 feedthrough
rlabel pdiffusion 1522 -1113 1522 -1113 0 feedthrough
rlabel pdiffusion 1529 -1113 1529 -1113 0 feedthrough
rlabel pdiffusion 1536 -1113 1536 -1113 0 feedthrough
rlabel pdiffusion 1543 -1113 1543 -1113 0 feedthrough
rlabel pdiffusion 1550 -1113 1550 -1113 0 feedthrough
rlabel pdiffusion 1557 -1113 1557 -1113 0 feedthrough
rlabel pdiffusion 1564 -1113 1564 -1113 0 feedthrough
rlabel pdiffusion 1571 -1113 1571 -1113 0 feedthrough
rlabel pdiffusion 1578 -1113 1578 -1113 0 feedthrough
rlabel pdiffusion 1585 -1113 1585 -1113 0 feedthrough
rlabel pdiffusion 1592 -1113 1592 -1113 0 feedthrough
rlabel pdiffusion 1599 -1113 1599 -1113 0 feedthrough
rlabel pdiffusion 1606 -1113 1606 -1113 0 feedthrough
rlabel pdiffusion 1613 -1113 1613 -1113 0 feedthrough
rlabel pdiffusion 1620 -1113 1620 -1113 0 feedthrough
rlabel pdiffusion 1627 -1113 1627 -1113 0 feedthrough
rlabel pdiffusion 1634 -1113 1634 -1113 0 feedthrough
rlabel pdiffusion 1641 -1113 1641 -1113 0 feedthrough
rlabel pdiffusion 1648 -1113 1648 -1113 0 feedthrough
rlabel pdiffusion 1655 -1113 1655 -1113 0 feedthrough
rlabel pdiffusion 1662 -1113 1662 -1113 0 feedthrough
rlabel pdiffusion 1669 -1113 1669 -1113 0 feedthrough
rlabel pdiffusion 1676 -1113 1676 -1113 0 feedthrough
rlabel pdiffusion 1683 -1113 1683 -1113 0 feedthrough
rlabel pdiffusion 1690 -1113 1690 -1113 0 feedthrough
rlabel pdiffusion 1697 -1113 1697 -1113 0 feedthrough
rlabel pdiffusion 1704 -1113 1704 -1113 0 feedthrough
rlabel pdiffusion 1711 -1113 1711 -1113 0 feedthrough
rlabel pdiffusion 1718 -1113 1718 -1113 0 feedthrough
rlabel pdiffusion 1725 -1113 1725 -1113 0 feedthrough
rlabel pdiffusion 1732 -1113 1732 -1113 0 feedthrough
rlabel pdiffusion 1739 -1113 1739 -1113 0 feedthrough
rlabel pdiffusion 1746 -1113 1746 -1113 0 feedthrough
rlabel pdiffusion 1753 -1113 1753 -1113 0 feedthrough
rlabel pdiffusion 1760 -1113 1760 -1113 0 feedthrough
rlabel pdiffusion 1767 -1113 1767 -1113 0 feedthrough
rlabel pdiffusion 1774 -1113 1774 -1113 0 feedthrough
rlabel pdiffusion 1781 -1113 1781 -1113 0 feedthrough
rlabel pdiffusion 1788 -1113 1788 -1113 0 feedthrough
rlabel pdiffusion 1795 -1113 1795 -1113 0 feedthrough
rlabel pdiffusion 1802 -1113 1802 -1113 0 feedthrough
rlabel pdiffusion 1809 -1113 1809 -1113 0 feedthrough
rlabel pdiffusion 1816 -1113 1816 -1113 0 feedthrough
rlabel pdiffusion 1823 -1113 1823 -1113 0 feedthrough
rlabel pdiffusion 1830 -1113 1830 -1113 0 feedthrough
rlabel pdiffusion 1837 -1113 1837 -1113 0 feedthrough
rlabel pdiffusion 1844 -1113 1844 -1113 0 feedthrough
rlabel pdiffusion 1851 -1113 1851 -1113 0 feedthrough
rlabel pdiffusion 1858 -1113 1858 -1113 0 feedthrough
rlabel pdiffusion 1865 -1113 1865 -1113 0 cellNo=779
rlabel pdiffusion 1872 -1113 1872 -1113 0 feedthrough
rlabel pdiffusion 1879 -1113 1879 -1113 0 feedthrough
rlabel pdiffusion 1928 -1113 1928 -1113 0 feedthrough
rlabel pdiffusion 1949 -1113 1949 -1113 0 feedthrough
rlabel pdiffusion 1963 -1113 1963 -1113 0 feedthrough
rlabel pdiffusion 1970 -1113 1970 -1113 0 feedthrough
rlabel pdiffusion 1977 -1113 1977 -1113 0 feedthrough
rlabel pdiffusion 3 -1248 3 -1248 0 feedthrough
rlabel pdiffusion 10 -1248 10 -1248 0 feedthrough
rlabel pdiffusion 17 -1248 17 -1248 0 feedthrough
rlabel pdiffusion 24 -1248 24 -1248 0 cellNo=1024
rlabel pdiffusion 31 -1248 31 -1248 0 feedthrough
rlabel pdiffusion 38 -1248 38 -1248 0 cellNo=725
rlabel pdiffusion 45 -1248 45 -1248 0 feedthrough
rlabel pdiffusion 52 -1248 52 -1248 0 feedthrough
rlabel pdiffusion 59 -1248 59 -1248 0 cellNo=773
rlabel pdiffusion 66 -1248 66 -1248 0 feedthrough
rlabel pdiffusion 73 -1248 73 -1248 0 feedthrough
rlabel pdiffusion 80 -1248 80 -1248 0 cellNo=222
rlabel pdiffusion 87 -1248 87 -1248 0 feedthrough
rlabel pdiffusion 94 -1248 94 -1248 0 feedthrough
rlabel pdiffusion 101 -1248 101 -1248 0 feedthrough
rlabel pdiffusion 108 -1248 108 -1248 0 feedthrough
rlabel pdiffusion 115 -1248 115 -1248 0 feedthrough
rlabel pdiffusion 122 -1248 122 -1248 0 cellNo=18
rlabel pdiffusion 129 -1248 129 -1248 0 feedthrough
rlabel pdiffusion 136 -1248 136 -1248 0 feedthrough
rlabel pdiffusion 143 -1248 143 -1248 0 feedthrough
rlabel pdiffusion 150 -1248 150 -1248 0 feedthrough
rlabel pdiffusion 157 -1248 157 -1248 0 cellNo=484
rlabel pdiffusion 164 -1248 164 -1248 0 feedthrough
rlabel pdiffusion 171 -1248 171 -1248 0 cellNo=314
rlabel pdiffusion 178 -1248 178 -1248 0 cellNo=195
rlabel pdiffusion 185 -1248 185 -1248 0 feedthrough
rlabel pdiffusion 192 -1248 192 -1248 0 feedthrough
rlabel pdiffusion 199 -1248 199 -1248 0 feedthrough
rlabel pdiffusion 206 -1248 206 -1248 0 feedthrough
rlabel pdiffusion 213 -1248 213 -1248 0 feedthrough
rlabel pdiffusion 220 -1248 220 -1248 0 feedthrough
rlabel pdiffusion 227 -1248 227 -1248 0 cellNo=858
rlabel pdiffusion 234 -1248 234 -1248 0 feedthrough
rlabel pdiffusion 241 -1248 241 -1248 0 feedthrough
rlabel pdiffusion 248 -1248 248 -1248 0 feedthrough
rlabel pdiffusion 255 -1248 255 -1248 0 feedthrough
rlabel pdiffusion 262 -1248 262 -1248 0 cellNo=387
rlabel pdiffusion 269 -1248 269 -1248 0 feedthrough
rlabel pdiffusion 276 -1248 276 -1248 0 feedthrough
rlabel pdiffusion 283 -1248 283 -1248 0 feedthrough
rlabel pdiffusion 290 -1248 290 -1248 0 cellNo=316
rlabel pdiffusion 297 -1248 297 -1248 0 feedthrough
rlabel pdiffusion 304 -1248 304 -1248 0 feedthrough
rlabel pdiffusion 311 -1248 311 -1248 0 feedthrough
rlabel pdiffusion 318 -1248 318 -1248 0 feedthrough
rlabel pdiffusion 325 -1248 325 -1248 0 feedthrough
rlabel pdiffusion 332 -1248 332 -1248 0 feedthrough
rlabel pdiffusion 339 -1248 339 -1248 0 feedthrough
rlabel pdiffusion 346 -1248 346 -1248 0 feedthrough
rlabel pdiffusion 353 -1248 353 -1248 0 feedthrough
rlabel pdiffusion 360 -1248 360 -1248 0 feedthrough
rlabel pdiffusion 367 -1248 367 -1248 0 feedthrough
rlabel pdiffusion 374 -1248 374 -1248 0 feedthrough
rlabel pdiffusion 381 -1248 381 -1248 0 feedthrough
rlabel pdiffusion 388 -1248 388 -1248 0 feedthrough
rlabel pdiffusion 395 -1248 395 -1248 0 feedthrough
rlabel pdiffusion 402 -1248 402 -1248 0 feedthrough
rlabel pdiffusion 409 -1248 409 -1248 0 feedthrough
rlabel pdiffusion 416 -1248 416 -1248 0 feedthrough
rlabel pdiffusion 423 -1248 423 -1248 0 cellNo=560
rlabel pdiffusion 430 -1248 430 -1248 0 feedthrough
rlabel pdiffusion 437 -1248 437 -1248 0 feedthrough
rlabel pdiffusion 444 -1248 444 -1248 0 cellNo=1
rlabel pdiffusion 451 -1248 451 -1248 0 cellNo=53
rlabel pdiffusion 458 -1248 458 -1248 0 feedthrough
rlabel pdiffusion 465 -1248 465 -1248 0 feedthrough
rlabel pdiffusion 472 -1248 472 -1248 0 cellNo=490
rlabel pdiffusion 479 -1248 479 -1248 0 feedthrough
rlabel pdiffusion 486 -1248 486 -1248 0 feedthrough
rlabel pdiffusion 493 -1248 493 -1248 0 feedthrough
rlabel pdiffusion 500 -1248 500 -1248 0 feedthrough
rlabel pdiffusion 507 -1248 507 -1248 0 feedthrough
rlabel pdiffusion 514 -1248 514 -1248 0 cellNo=178
rlabel pdiffusion 521 -1248 521 -1248 0 feedthrough
rlabel pdiffusion 528 -1248 528 -1248 0 feedthrough
rlabel pdiffusion 535 -1248 535 -1248 0 feedthrough
rlabel pdiffusion 542 -1248 542 -1248 0 feedthrough
rlabel pdiffusion 549 -1248 549 -1248 0 feedthrough
rlabel pdiffusion 556 -1248 556 -1248 0 feedthrough
rlabel pdiffusion 563 -1248 563 -1248 0 cellNo=119
rlabel pdiffusion 570 -1248 570 -1248 0 feedthrough
rlabel pdiffusion 577 -1248 577 -1248 0 feedthrough
rlabel pdiffusion 584 -1248 584 -1248 0 cellNo=549
rlabel pdiffusion 591 -1248 591 -1248 0 feedthrough
rlabel pdiffusion 598 -1248 598 -1248 0 feedthrough
rlabel pdiffusion 605 -1248 605 -1248 0 feedthrough
rlabel pdiffusion 612 -1248 612 -1248 0 feedthrough
rlabel pdiffusion 619 -1248 619 -1248 0 feedthrough
rlabel pdiffusion 626 -1248 626 -1248 0 feedthrough
rlabel pdiffusion 633 -1248 633 -1248 0 feedthrough
rlabel pdiffusion 640 -1248 640 -1248 0 feedthrough
rlabel pdiffusion 647 -1248 647 -1248 0 feedthrough
rlabel pdiffusion 654 -1248 654 -1248 0 feedthrough
rlabel pdiffusion 661 -1248 661 -1248 0 feedthrough
rlabel pdiffusion 668 -1248 668 -1248 0 cellNo=469
rlabel pdiffusion 675 -1248 675 -1248 0 feedthrough
rlabel pdiffusion 682 -1248 682 -1248 0 feedthrough
rlabel pdiffusion 689 -1248 689 -1248 0 feedthrough
rlabel pdiffusion 696 -1248 696 -1248 0 feedthrough
rlabel pdiffusion 703 -1248 703 -1248 0 feedthrough
rlabel pdiffusion 710 -1248 710 -1248 0 feedthrough
rlabel pdiffusion 717 -1248 717 -1248 0 feedthrough
rlabel pdiffusion 724 -1248 724 -1248 0 feedthrough
rlabel pdiffusion 731 -1248 731 -1248 0 feedthrough
rlabel pdiffusion 738 -1248 738 -1248 0 feedthrough
rlabel pdiffusion 745 -1248 745 -1248 0 feedthrough
rlabel pdiffusion 752 -1248 752 -1248 0 feedthrough
rlabel pdiffusion 759 -1248 759 -1248 0 feedthrough
rlabel pdiffusion 766 -1248 766 -1248 0 feedthrough
rlabel pdiffusion 773 -1248 773 -1248 0 cellNo=464
rlabel pdiffusion 780 -1248 780 -1248 0 cellNo=631
rlabel pdiffusion 787 -1248 787 -1248 0 feedthrough
rlabel pdiffusion 794 -1248 794 -1248 0 cellNo=63
rlabel pdiffusion 801 -1248 801 -1248 0 feedthrough
rlabel pdiffusion 808 -1248 808 -1248 0 cellNo=460
rlabel pdiffusion 815 -1248 815 -1248 0 feedthrough
rlabel pdiffusion 822 -1248 822 -1248 0 cellNo=948
rlabel pdiffusion 829 -1248 829 -1248 0 feedthrough
rlabel pdiffusion 836 -1248 836 -1248 0 feedthrough
rlabel pdiffusion 843 -1248 843 -1248 0 feedthrough
rlabel pdiffusion 850 -1248 850 -1248 0 feedthrough
rlabel pdiffusion 857 -1248 857 -1248 0 cellNo=509
rlabel pdiffusion 864 -1248 864 -1248 0 feedthrough
rlabel pdiffusion 871 -1248 871 -1248 0 cellNo=303
rlabel pdiffusion 878 -1248 878 -1248 0 cellNo=478
rlabel pdiffusion 885 -1248 885 -1248 0 feedthrough
rlabel pdiffusion 892 -1248 892 -1248 0 feedthrough
rlabel pdiffusion 899 -1248 899 -1248 0 feedthrough
rlabel pdiffusion 906 -1248 906 -1248 0 cellNo=210
rlabel pdiffusion 913 -1248 913 -1248 0 feedthrough
rlabel pdiffusion 920 -1248 920 -1248 0 feedthrough
rlabel pdiffusion 927 -1248 927 -1248 0 cellNo=205
rlabel pdiffusion 934 -1248 934 -1248 0 feedthrough
rlabel pdiffusion 941 -1248 941 -1248 0 feedthrough
rlabel pdiffusion 948 -1248 948 -1248 0 feedthrough
rlabel pdiffusion 955 -1248 955 -1248 0 feedthrough
rlabel pdiffusion 962 -1248 962 -1248 0 cellNo=429
rlabel pdiffusion 969 -1248 969 -1248 0 feedthrough
rlabel pdiffusion 976 -1248 976 -1248 0 feedthrough
rlabel pdiffusion 983 -1248 983 -1248 0 feedthrough
rlabel pdiffusion 990 -1248 990 -1248 0 feedthrough
rlabel pdiffusion 997 -1248 997 -1248 0 feedthrough
rlabel pdiffusion 1004 -1248 1004 -1248 0 feedthrough
rlabel pdiffusion 1011 -1248 1011 -1248 0 feedthrough
rlabel pdiffusion 1018 -1248 1018 -1248 0 cellNo=991
rlabel pdiffusion 1025 -1248 1025 -1248 0 feedthrough
rlabel pdiffusion 1032 -1248 1032 -1248 0 feedthrough
rlabel pdiffusion 1039 -1248 1039 -1248 0 feedthrough
rlabel pdiffusion 1046 -1248 1046 -1248 0 cellNo=56
rlabel pdiffusion 1053 -1248 1053 -1248 0 feedthrough
rlabel pdiffusion 1060 -1248 1060 -1248 0 feedthrough
rlabel pdiffusion 1067 -1248 1067 -1248 0 feedthrough
rlabel pdiffusion 1074 -1248 1074 -1248 0 feedthrough
rlabel pdiffusion 1081 -1248 1081 -1248 0 feedthrough
rlabel pdiffusion 1088 -1248 1088 -1248 0 feedthrough
rlabel pdiffusion 1095 -1248 1095 -1248 0 feedthrough
rlabel pdiffusion 1102 -1248 1102 -1248 0 feedthrough
rlabel pdiffusion 1109 -1248 1109 -1248 0 feedthrough
rlabel pdiffusion 1116 -1248 1116 -1248 0 feedthrough
rlabel pdiffusion 1123 -1248 1123 -1248 0 feedthrough
rlabel pdiffusion 1130 -1248 1130 -1248 0 cellNo=806
rlabel pdiffusion 1137 -1248 1137 -1248 0 feedthrough
rlabel pdiffusion 1144 -1248 1144 -1248 0 feedthrough
rlabel pdiffusion 1151 -1248 1151 -1248 0 feedthrough
rlabel pdiffusion 1158 -1248 1158 -1248 0 cellNo=369
rlabel pdiffusion 1165 -1248 1165 -1248 0 feedthrough
rlabel pdiffusion 1172 -1248 1172 -1248 0 feedthrough
rlabel pdiffusion 1179 -1248 1179 -1248 0 cellNo=957
rlabel pdiffusion 1186 -1248 1186 -1248 0 feedthrough
rlabel pdiffusion 1193 -1248 1193 -1248 0 feedthrough
rlabel pdiffusion 1200 -1248 1200 -1248 0 feedthrough
rlabel pdiffusion 1207 -1248 1207 -1248 0 feedthrough
rlabel pdiffusion 1214 -1248 1214 -1248 0 feedthrough
rlabel pdiffusion 1221 -1248 1221 -1248 0 feedthrough
rlabel pdiffusion 1228 -1248 1228 -1248 0 feedthrough
rlabel pdiffusion 1235 -1248 1235 -1248 0 feedthrough
rlabel pdiffusion 1242 -1248 1242 -1248 0 feedthrough
rlabel pdiffusion 1249 -1248 1249 -1248 0 feedthrough
rlabel pdiffusion 1256 -1248 1256 -1248 0 feedthrough
rlabel pdiffusion 1263 -1248 1263 -1248 0 feedthrough
rlabel pdiffusion 1270 -1248 1270 -1248 0 feedthrough
rlabel pdiffusion 1277 -1248 1277 -1248 0 feedthrough
rlabel pdiffusion 1284 -1248 1284 -1248 0 feedthrough
rlabel pdiffusion 1291 -1248 1291 -1248 0 feedthrough
rlabel pdiffusion 1298 -1248 1298 -1248 0 feedthrough
rlabel pdiffusion 1305 -1248 1305 -1248 0 feedthrough
rlabel pdiffusion 1312 -1248 1312 -1248 0 feedthrough
rlabel pdiffusion 1319 -1248 1319 -1248 0 feedthrough
rlabel pdiffusion 1326 -1248 1326 -1248 0 feedthrough
rlabel pdiffusion 1333 -1248 1333 -1248 0 feedthrough
rlabel pdiffusion 1340 -1248 1340 -1248 0 feedthrough
rlabel pdiffusion 1347 -1248 1347 -1248 0 feedthrough
rlabel pdiffusion 1354 -1248 1354 -1248 0 feedthrough
rlabel pdiffusion 1361 -1248 1361 -1248 0 feedthrough
rlabel pdiffusion 1368 -1248 1368 -1248 0 feedthrough
rlabel pdiffusion 1375 -1248 1375 -1248 0 feedthrough
rlabel pdiffusion 1382 -1248 1382 -1248 0 feedthrough
rlabel pdiffusion 1389 -1248 1389 -1248 0 feedthrough
rlabel pdiffusion 1396 -1248 1396 -1248 0 feedthrough
rlabel pdiffusion 1403 -1248 1403 -1248 0 feedthrough
rlabel pdiffusion 1410 -1248 1410 -1248 0 feedthrough
rlabel pdiffusion 1417 -1248 1417 -1248 0 feedthrough
rlabel pdiffusion 1424 -1248 1424 -1248 0 feedthrough
rlabel pdiffusion 1431 -1248 1431 -1248 0 feedthrough
rlabel pdiffusion 1438 -1248 1438 -1248 0 feedthrough
rlabel pdiffusion 1445 -1248 1445 -1248 0 feedthrough
rlabel pdiffusion 1452 -1248 1452 -1248 0 feedthrough
rlabel pdiffusion 1459 -1248 1459 -1248 0 feedthrough
rlabel pdiffusion 1466 -1248 1466 -1248 0 feedthrough
rlabel pdiffusion 1473 -1248 1473 -1248 0 feedthrough
rlabel pdiffusion 1480 -1248 1480 -1248 0 feedthrough
rlabel pdiffusion 1487 -1248 1487 -1248 0 feedthrough
rlabel pdiffusion 1494 -1248 1494 -1248 0 feedthrough
rlabel pdiffusion 1501 -1248 1501 -1248 0 feedthrough
rlabel pdiffusion 1508 -1248 1508 -1248 0 feedthrough
rlabel pdiffusion 1515 -1248 1515 -1248 0 feedthrough
rlabel pdiffusion 1522 -1248 1522 -1248 0 feedthrough
rlabel pdiffusion 1529 -1248 1529 -1248 0 feedthrough
rlabel pdiffusion 1536 -1248 1536 -1248 0 feedthrough
rlabel pdiffusion 1543 -1248 1543 -1248 0 feedthrough
rlabel pdiffusion 1550 -1248 1550 -1248 0 feedthrough
rlabel pdiffusion 1557 -1248 1557 -1248 0 feedthrough
rlabel pdiffusion 1564 -1248 1564 -1248 0 feedthrough
rlabel pdiffusion 1571 -1248 1571 -1248 0 feedthrough
rlabel pdiffusion 1578 -1248 1578 -1248 0 feedthrough
rlabel pdiffusion 1585 -1248 1585 -1248 0 feedthrough
rlabel pdiffusion 1592 -1248 1592 -1248 0 feedthrough
rlabel pdiffusion 1599 -1248 1599 -1248 0 feedthrough
rlabel pdiffusion 1606 -1248 1606 -1248 0 feedthrough
rlabel pdiffusion 1613 -1248 1613 -1248 0 feedthrough
rlabel pdiffusion 1620 -1248 1620 -1248 0 feedthrough
rlabel pdiffusion 1627 -1248 1627 -1248 0 feedthrough
rlabel pdiffusion 1634 -1248 1634 -1248 0 feedthrough
rlabel pdiffusion 1641 -1248 1641 -1248 0 feedthrough
rlabel pdiffusion 1648 -1248 1648 -1248 0 feedthrough
rlabel pdiffusion 1655 -1248 1655 -1248 0 feedthrough
rlabel pdiffusion 1662 -1248 1662 -1248 0 feedthrough
rlabel pdiffusion 1669 -1248 1669 -1248 0 feedthrough
rlabel pdiffusion 1676 -1248 1676 -1248 0 feedthrough
rlabel pdiffusion 1683 -1248 1683 -1248 0 feedthrough
rlabel pdiffusion 1690 -1248 1690 -1248 0 feedthrough
rlabel pdiffusion 1697 -1248 1697 -1248 0 feedthrough
rlabel pdiffusion 1704 -1248 1704 -1248 0 feedthrough
rlabel pdiffusion 1711 -1248 1711 -1248 0 feedthrough
rlabel pdiffusion 1718 -1248 1718 -1248 0 feedthrough
rlabel pdiffusion 1725 -1248 1725 -1248 0 feedthrough
rlabel pdiffusion 1732 -1248 1732 -1248 0 feedthrough
rlabel pdiffusion 1739 -1248 1739 -1248 0 feedthrough
rlabel pdiffusion 1746 -1248 1746 -1248 0 feedthrough
rlabel pdiffusion 1753 -1248 1753 -1248 0 feedthrough
rlabel pdiffusion 1760 -1248 1760 -1248 0 feedthrough
rlabel pdiffusion 1767 -1248 1767 -1248 0 feedthrough
rlabel pdiffusion 1774 -1248 1774 -1248 0 feedthrough
rlabel pdiffusion 1781 -1248 1781 -1248 0 feedthrough
rlabel pdiffusion 1788 -1248 1788 -1248 0 feedthrough
rlabel pdiffusion 1795 -1248 1795 -1248 0 feedthrough
rlabel pdiffusion 1802 -1248 1802 -1248 0 feedthrough
rlabel pdiffusion 1809 -1248 1809 -1248 0 feedthrough
rlabel pdiffusion 1816 -1248 1816 -1248 0 feedthrough
rlabel pdiffusion 1823 -1248 1823 -1248 0 feedthrough
rlabel pdiffusion 1830 -1248 1830 -1248 0 feedthrough
rlabel pdiffusion 1837 -1248 1837 -1248 0 feedthrough
rlabel pdiffusion 1844 -1248 1844 -1248 0 feedthrough
rlabel pdiffusion 1851 -1248 1851 -1248 0 feedthrough
rlabel pdiffusion 1858 -1248 1858 -1248 0 feedthrough
rlabel pdiffusion 1865 -1248 1865 -1248 0 feedthrough
rlabel pdiffusion 1872 -1248 1872 -1248 0 feedthrough
rlabel pdiffusion 1879 -1248 1879 -1248 0 feedthrough
rlabel pdiffusion 1886 -1248 1886 -1248 0 feedthrough
rlabel pdiffusion 1893 -1248 1893 -1248 0 feedthrough
rlabel pdiffusion 1900 -1248 1900 -1248 0 feedthrough
rlabel pdiffusion 1907 -1248 1907 -1248 0 feedthrough
rlabel pdiffusion 1914 -1248 1914 -1248 0 feedthrough
rlabel pdiffusion 1921 -1248 1921 -1248 0 feedthrough
rlabel pdiffusion 1928 -1248 1928 -1248 0 feedthrough
rlabel pdiffusion 1956 -1248 1956 -1248 0 feedthrough
rlabel pdiffusion 1963 -1248 1963 -1248 0 feedthrough
rlabel pdiffusion 1970 -1248 1970 -1248 0 feedthrough
rlabel pdiffusion 1977 -1248 1977 -1248 0 feedthrough
rlabel pdiffusion 1991 -1248 1991 -1248 0 feedthrough
rlabel pdiffusion 3 -1391 3 -1391 0 cellNo=1029
rlabel pdiffusion 10 -1391 10 -1391 0 feedthrough
rlabel pdiffusion 17 -1391 17 -1391 0 feedthrough
rlabel pdiffusion 24 -1391 24 -1391 0 feedthrough
rlabel pdiffusion 31 -1391 31 -1391 0 feedthrough
rlabel pdiffusion 38 -1391 38 -1391 0 feedthrough
rlabel pdiffusion 45 -1391 45 -1391 0 feedthrough
rlabel pdiffusion 52 -1391 52 -1391 0 cellNo=952
rlabel pdiffusion 59 -1391 59 -1391 0 cellNo=30
rlabel pdiffusion 66 -1391 66 -1391 0 feedthrough
rlabel pdiffusion 73 -1391 73 -1391 0 cellNo=998
rlabel pdiffusion 80 -1391 80 -1391 0 feedthrough
rlabel pdiffusion 87 -1391 87 -1391 0 feedthrough
rlabel pdiffusion 94 -1391 94 -1391 0 feedthrough
rlabel pdiffusion 101 -1391 101 -1391 0 feedthrough
rlabel pdiffusion 108 -1391 108 -1391 0 cellNo=194
rlabel pdiffusion 115 -1391 115 -1391 0 feedthrough
rlabel pdiffusion 122 -1391 122 -1391 0 feedthrough
rlabel pdiffusion 129 -1391 129 -1391 0 cellNo=32
rlabel pdiffusion 136 -1391 136 -1391 0 feedthrough
rlabel pdiffusion 143 -1391 143 -1391 0 cellNo=435
rlabel pdiffusion 150 -1391 150 -1391 0 cellNo=386
rlabel pdiffusion 157 -1391 157 -1391 0 feedthrough
rlabel pdiffusion 164 -1391 164 -1391 0 cellNo=507
rlabel pdiffusion 171 -1391 171 -1391 0 feedthrough
rlabel pdiffusion 178 -1391 178 -1391 0 feedthrough
rlabel pdiffusion 185 -1391 185 -1391 0 feedthrough
rlabel pdiffusion 192 -1391 192 -1391 0 feedthrough
rlabel pdiffusion 199 -1391 199 -1391 0 feedthrough
rlabel pdiffusion 206 -1391 206 -1391 0 cellNo=884
rlabel pdiffusion 213 -1391 213 -1391 0 feedthrough
rlabel pdiffusion 220 -1391 220 -1391 0 feedthrough
rlabel pdiffusion 227 -1391 227 -1391 0 feedthrough
rlabel pdiffusion 234 -1391 234 -1391 0 feedthrough
rlabel pdiffusion 241 -1391 241 -1391 0 feedthrough
rlabel pdiffusion 248 -1391 248 -1391 0 feedthrough
rlabel pdiffusion 255 -1391 255 -1391 0 feedthrough
rlabel pdiffusion 262 -1391 262 -1391 0 feedthrough
rlabel pdiffusion 269 -1391 269 -1391 0 feedthrough
rlabel pdiffusion 276 -1391 276 -1391 0 feedthrough
rlabel pdiffusion 283 -1391 283 -1391 0 feedthrough
rlabel pdiffusion 290 -1391 290 -1391 0 feedthrough
rlabel pdiffusion 297 -1391 297 -1391 0 feedthrough
rlabel pdiffusion 304 -1391 304 -1391 0 feedthrough
rlabel pdiffusion 311 -1391 311 -1391 0 feedthrough
rlabel pdiffusion 318 -1391 318 -1391 0 feedthrough
rlabel pdiffusion 325 -1391 325 -1391 0 feedthrough
rlabel pdiffusion 332 -1391 332 -1391 0 feedthrough
rlabel pdiffusion 339 -1391 339 -1391 0 feedthrough
rlabel pdiffusion 346 -1391 346 -1391 0 feedthrough
rlabel pdiffusion 353 -1391 353 -1391 0 feedthrough
rlabel pdiffusion 360 -1391 360 -1391 0 feedthrough
rlabel pdiffusion 367 -1391 367 -1391 0 feedthrough
rlabel pdiffusion 374 -1391 374 -1391 0 feedthrough
rlabel pdiffusion 381 -1391 381 -1391 0 feedthrough
rlabel pdiffusion 388 -1391 388 -1391 0 feedthrough
rlabel pdiffusion 395 -1391 395 -1391 0 feedthrough
rlabel pdiffusion 402 -1391 402 -1391 0 feedthrough
rlabel pdiffusion 409 -1391 409 -1391 0 feedthrough
rlabel pdiffusion 416 -1391 416 -1391 0 feedthrough
rlabel pdiffusion 423 -1391 423 -1391 0 feedthrough
rlabel pdiffusion 430 -1391 430 -1391 0 cellNo=181
rlabel pdiffusion 437 -1391 437 -1391 0 feedthrough
rlabel pdiffusion 444 -1391 444 -1391 0 feedthrough
rlabel pdiffusion 451 -1391 451 -1391 0 feedthrough
rlabel pdiffusion 458 -1391 458 -1391 0 feedthrough
rlabel pdiffusion 465 -1391 465 -1391 0 feedthrough
rlabel pdiffusion 472 -1391 472 -1391 0 feedthrough
rlabel pdiffusion 479 -1391 479 -1391 0 feedthrough
rlabel pdiffusion 486 -1391 486 -1391 0 feedthrough
rlabel pdiffusion 493 -1391 493 -1391 0 feedthrough
rlabel pdiffusion 500 -1391 500 -1391 0 feedthrough
rlabel pdiffusion 507 -1391 507 -1391 0 feedthrough
rlabel pdiffusion 514 -1391 514 -1391 0 feedthrough
rlabel pdiffusion 521 -1391 521 -1391 0 feedthrough
rlabel pdiffusion 528 -1391 528 -1391 0 cellNo=643
rlabel pdiffusion 535 -1391 535 -1391 0 feedthrough
rlabel pdiffusion 542 -1391 542 -1391 0 feedthrough
rlabel pdiffusion 549 -1391 549 -1391 0 feedthrough
rlabel pdiffusion 556 -1391 556 -1391 0 feedthrough
rlabel pdiffusion 563 -1391 563 -1391 0 feedthrough
rlabel pdiffusion 570 -1391 570 -1391 0 feedthrough
rlabel pdiffusion 577 -1391 577 -1391 0 cellNo=641
rlabel pdiffusion 584 -1391 584 -1391 0 feedthrough
rlabel pdiffusion 591 -1391 591 -1391 0 feedthrough
rlabel pdiffusion 598 -1391 598 -1391 0 feedthrough
rlabel pdiffusion 605 -1391 605 -1391 0 feedthrough
rlabel pdiffusion 612 -1391 612 -1391 0 feedthrough
rlabel pdiffusion 619 -1391 619 -1391 0 feedthrough
rlabel pdiffusion 626 -1391 626 -1391 0 cellNo=987
rlabel pdiffusion 633 -1391 633 -1391 0 feedthrough
rlabel pdiffusion 640 -1391 640 -1391 0 feedthrough
rlabel pdiffusion 647 -1391 647 -1391 0 feedthrough
rlabel pdiffusion 654 -1391 654 -1391 0 cellNo=558
rlabel pdiffusion 661 -1391 661 -1391 0 feedthrough
rlabel pdiffusion 668 -1391 668 -1391 0 cellNo=31
rlabel pdiffusion 675 -1391 675 -1391 0 cellNo=541
rlabel pdiffusion 682 -1391 682 -1391 0 feedthrough
rlabel pdiffusion 689 -1391 689 -1391 0 feedthrough
rlabel pdiffusion 696 -1391 696 -1391 0 feedthrough
rlabel pdiffusion 703 -1391 703 -1391 0 feedthrough
rlabel pdiffusion 710 -1391 710 -1391 0 cellNo=20
rlabel pdiffusion 717 -1391 717 -1391 0 feedthrough
rlabel pdiffusion 724 -1391 724 -1391 0 feedthrough
rlabel pdiffusion 731 -1391 731 -1391 0 feedthrough
rlabel pdiffusion 738 -1391 738 -1391 0 feedthrough
rlabel pdiffusion 745 -1391 745 -1391 0 feedthrough
rlabel pdiffusion 752 -1391 752 -1391 0 feedthrough
rlabel pdiffusion 759 -1391 759 -1391 0 feedthrough
rlabel pdiffusion 766 -1391 766 -1391 0 feedthrough
rlabel pdiffusion 773 -1391 773 -1391 0 feedthrough
rlabel pdiffusion 780 -1391 780 -1391 0 feedthrough
rlabel pdiffusion 787 -1391 787 -1391 0 feedthrough
rlabel pdiffusion 794 -1391 794 -1391 0 feedthrough
rlabel pdiffusion 801 -1391 801 -1391 0 feedthrough
rlabel pdiffusion 808 -1391 808 -1391 0 feedthrough
rlabel pdiffusion 815 -1391 815 -1391 0 feedthrough
rlabel pdiffusion 822 -1391 822 -1391 0 feedthrough
rlabel pdiffusion 829 -1391 829 -1391 0 feedthrough
rlabel pdiffusion 836 -1391 836 -1391 0 cellNo=732
rlabel pdiffusion 843 -1391 843 -1391 0 feedthrough
rlabel pdiffusion 850 -1391 850 -1391 0 feedthrough
rlabel pdiffusion 857 -1391 857 -1391 0 cellNo=163
rlabel pdiffusion 864 -1391 864 -1391 0 feedthrough
rlabel pdiffusion 871 -1391 871 -1391 0 feedthrough
rlabel pdiffusion 878 -1391 878 -1391 0 feedthrough
rlabel pdiffusion 885 -1391 885 -1391 0 feedthrough
rlabel pdiffusion 892 -1391 892 -1391 0 feedthrough
rlabel pdiffusion 899 -1391 899 -1391 0 feedthrough
rlabel pdiffusion 906 -1391 906 -1391 0 feedthrough
rlabel pdiffusion 913 -1391 913 -1391 0 feedthrough
rlabel pdiffusion 920 -1391 920 -1391 0 cellNo=496
rlabel pdiffusion 927 -1391 927 -1391 0 cellNo=680
rlabel pdiffusion 934 -1391 934 -1391 0 feedthrough
rlabel pdiffusion 941 -1391 941 -1391 0 cellNo=107
rlabel pdiffusion 948 -1391 948 -1391 0 feedthrough
rlabel pdiffusion 955 -1391 955 -1391 0 feedthrough
rlabel pdiffusion 962 -1391 962 -1391 0 feedthrough
rlabel pdiffusion 969 -1391 969 -1391 0 cellNo=93
rlabel pdiffusion 976 -1391 976 -1391 0 feedthrough
rlabel pdiffusion 983 -1391 983 -1391 0 feedthrough
rlabel pdiffusion 990 -1391 990 -1391 0 feedthrough
rlabel pdiffusion 997 -1391 997 -1391 0 cellNo=736
rlabel pdiffusion 1004 -1391 1004 -1391 0 feedthrough
rlabel pdiffusion 1011 -1391 1011 -1391 0 feedthrough
rlabel pdiffusion 1018 -1391 1018 -1391 0 feedthrough
rlabel pdiffusion 1025 -1391 1025 -1391 0 feedthrough
rlabel pdiffusion 1032 -1391 1032 -1391 0 cellNo=47
rlabel pdiffusion 1039 -1391 1039 -1391 0 feedthrough
rlabel pdiffusion 1046 -1391 1046 -1391 0 feedthrough
rlabel pdiffusion 1053 -1391 1053 -1391 0 cellNo=73
rlabel pdiffusion 1060 -1391 1060 -1391 0 feedthrough
rlabel pdiffusion 1067 -1391 1067 -1391 0 cellNo=981
rlabel pdiffusion 1074 -1391 1074 -1391 0 cellNo=345
rlabel pdiffusion 1081 -1391 1081 -1391 0 feedthrough
rlabel pdiffusion 1088 -1391 1088 -1391 0 feedthrough
rlabel pdiffusion 1095 -1391 1095 -1391 0 feedthrough
rlabel pdiffusion 1102 -1391 1102 -1391 0 feedthrough
rlabel pdiffusion 1109 -1391 1109 -1391 0 cellNo=349
rlabel pdiffusion 1116 -1391 1116 -1391 0 feedthrough
rlabel pdiffusion 1123 -1391 1123 -1391 0 feedthrough
rlabel pdiffusion 1130 -1391 1130 -1391 0 feedthrough
rlabel pdiffusion 1137 -1391 1137 -1391 0 feedthrough
rlabel pdiffusion 1144 -1391 1144 -1391 0 feedthrough
rlabel pdiffusion 1151 -1391 1151 -1391 0 feedthrough
rlabel pdiffusion 1158 -1391 1158 -1391 0 feedthrough
rlabel pdiffusion 1165 -1391 1165 -1391 0 feedthrough
rlabel pdiffusion 1172 -1391 1172 -1391 0 cellNo=878
rlabel pdiffusion 1179 -1391 1179 -1391 0 feedthrough
rlabel pdiffusion 1186 -1391 1186 -1391 0 cellNo=886
rlabel pdiffusion 1193 -1391 1193 -1391 0 feedthrough
rlabel pdiffusion 1200 -1391 1200 -1391 0 feedthrough
rlabel pdiffusion 1207 -1391 1207 -1391 0 feedthrough
rlabel pdiffusion 1214 -1391 1214 -1391 0 feedthrough
rlabel pdiffusion 1221 -1391 1221 -1391 0 feedthrough
rlabel pdiffusion 1228 -1391 1228 -1391 0 feedthrough
rlabel pdiffusion 1235 -1391 1235 -1391 0 feedthrough
rlabel pdiffusion 1242 -1391 1242 -1391 0 cellNo=852
rlabel pdiffusion 1249 -1391 1249 -1391 0 feedthrough
rlabel pdiffusion 1256 -1391 1256 -1391 0 feedthrough
rlabel pdiffusion 1263 -1391 1263 -1391 0 feedthrough
rlabel pdiffusion 1270 -1391 1270 -1391 0 feedthrough
rlabel pdiffusion 1277 -1391 1277 -1391 0 feedthrough
rlabel pdiffusion 1284 -1391 1284 -1391 0 cellNo=784
rlabel pdiffusion 1291 -1391 1291 -1391 0 feedthrough
rlabel pdiffusion 1298 -1391 1298 -1391 0 feedthrough
rlabel pdiffusion 1305 -1391 1305 -1391 0 feedthrough
rlabel pdiffusion 1312 -1391 1312 -1391 0 feedthrough
rlabel pdiffusion 1319 -1391 1319 -1391 0 feedthrough
rlabel pdiffusion 1326 -1391 1326 -1391 0 feedthrough
rlabel pdiffusion 1333 -1391 1333 -1391 0 feedthrough
rlabel pdiffusion 1340 -1391 1340 -1391 0 feedthrough
rlabel pdiffusion 1347 -1391 1347 -1391 0 feedthrough
rlabel pdiffusion 1354 -1391 1354 -1391 0 feedthrough
rlabel pdiffusion 1361 -1391 1361 -1391 0 feedthrough
rlabel pdiffusion 1368 -1391 1368 -1391 0 feedthrough
rlabel pdiffusion 1375 -1391 1375 -1391 0 feedthrough
rlabel pdiffusion 1382 -1391 1382 -1391 0 feedthrough
rlabel pdiffusion 1389 -1391 1389 -1391 0 feedthrough
rlabel pdiffusion 1396 -1391 1396 -1391 0 feedthrough
rlabel pdiffusion 1403 -1391 1403 -1391 0 feedthrough
rlabel pdiffusion 1410 -1391 1410 -1391 0 feedthrough
rlabel pdiffusion 1417 -1391 1417 -1391 0 feedthrough
rlabel pdiffusion 1424 -1391 1424 -1391 0 feedthrough
rlabel pdiffusion 1431 -1391 1431 -1391 0 feedthrough
rlabel pdiffusion 1438 -1391 1438 -1391 0 feedthrough
rlabel pdiffusion 1445 -1391 1445 -1391 0 feedthrough
rlabel pdiffusion 1452 -1391 1452 -1391 0 feedthrough
rlabel pdiffusion 1459 -1391 1459 -1391 0 feedthrough
rlabel pdiffusion 1466 -1391 1466 -1391 0 feedthrough
rlabel pdiffusion 1473 -1391 1473 -1391 0 feedthrough
rlabel pdiffusion 1480 -1391 1480 -1391 0 feedthrough
rlabel pdiffusion 1487 -1391 1487 -1391 0 feedthrough
rlabel pdiffusion 1494 -1391 1494 -1391 0 feedthrough
rlabel pdiffusion 1501 -1391 1501 -1391 0 feedthrough
rlabel pdiffusion 1508 -1391 1508 -1391 0 feedthrough
rlabel pdiffusion 1515 -1391 1515 -1391 0 feedthrough
rlabel pdiffusion 1522 -1391 1522 -1391 0 feedthrough
rlabel pdiffusion 1529 -1391 1529 -1391 0 feedthrough
rlabel pdiffusion 1536 -1391 1536 -1391 0 feedthrough
rlabel pdiffusion 1543 -1391 1543 -1391 0 feedthrough
rlabel pdiffusion 1550 -1391 1550 -1391 0 feedthrough
rlabel pdiffusion 1557 -1391 1557 -1391 0 feedthrough
rlabel pdiffusion 1564 -1391 1564 -1391 0 feedthrough
rlabel pdiffusion 1571 -1391 1571 -1391 0 feedthrough
rlabel pdiffusion 1578 -1391 1578 -1391 0 feedthrough
rlabel pdiffusion 1585 -1391 1585 -1391 0 feedthrough
rlabel pdiffusion 1592 -1391 1592 -1391 0 feedthrough
rlabel pdiffusion 1599 -1391 1599 -1391 0 feedthrough
rlabel pdiffusion 1606 -1391 1606 -1391 0 feedthrough
rlabel pdiffusion 1613 -1391 1613 -1391 0 feedthrough
rlabel pdiffusion 1620 -1391 1620 -1391 0 feedthrough
rlabel pdiffusion 1627 -1391 1627 -1391 0 feedthrough
rlabel pdiffusion 1634 -1391 1634 -1391 0 feedthrough
rlabel pdiffusion 1641 -1391 1641 -1391 0 feedthrough
rlabel pdiffusion 1648 -1391 1648 -1391 0 feedthrough
rlabel pdiffusion 1655 -1391 1655 -1391 0 feedthrough
rlabel pdiffusion 1662 -1391 1662 -1391 0 feedthrough
rlabel pdiffusion 1669 -1391 1669 -1391 0 feedthrough
rlabel pdiffusion 1676 -1391 1676 -1391 0 feedthrough
rlabel pdiffusion 1683 -1391 1683 -1391 0 feedthrough
rlabel pdiffusion 1690 -1391 1690 -1391 0 feedthrough
rlabel pdiffusion 1697 -1391 1697 -1391 0 feedthrough
rlabel pdiffusion 1704 -1391 1704 -1391 0 feedthrough
rlabel pdiffusion 1711 -1391 1711 -1391 0 feedthrough
rlabel pdiffusion 1718 -1391 1718 -1391 0 feedthrough
rlabel pdiffusion 1725 -1391 1725 -1391 0 feedthrough
rlabel pdiffusion 1732 -1391 1732 -1391 0 feedthrough
rlabel pdiffusion 1739 -1391 1739 -1391 0 feedthrough
rlabel pdiffusion 1746 -1391 1746 -1391 0 feedthrough
rlabel pdiffusion 1753 -1391 1753 -1391 0 feedthrough
rlabel pdiffusion 1760 -1391 1760 -1391 0 feedthrough
rlabel pdiffusion 1767 -1391 1767 -1391 0 feedthrough
rlabel pdiffusion 1774 -1391 1774 -1391 0 feedthrough
rlabel pdiffusion 1781 -1391 1781 -1391 0 feedthrough
rlabel pdiffusion 1788 -1391 1788 -1391 0 feedthrough
rlabel pdiffusion 1795 -1391 1795 -1391 0 feedthrough
rlabel pdiffusion 1802 -1391 1802 -1391 0 feedthrough
rlabel pdiffusion 1809 -1391 1809 -1391 0 feedthrough
rlabel pdiffusion 1816 -1391 1816 -1391 0 feedthrough
rlabel pdiffusion 1823 -1391 1823 -1391 0 feedthrough
rlabel pdiffusion 1830 -1391 1830 -1391 0 feedthrough
rlabel pdiffusion 1837 -1391 1837 -1391 0 feedthrough
rlabel pdiffusion 1844 -1391 1844 -1391 0 feedthrough
rlabel pdiffusion 1851 -1391 1851 -1391 0 feedthrough
rlabel pdiffusion 1858 -1391 1858 -1391 0 feedthrough
rlabel pdiffusion 1865 -1391 1865 -1391 0 feedthrough
rlabel pdiffusion 1872 -1391 1872 -1391 0 feedthrough
rlabel pdiffusion 1879 -1391 1879 -1391 0 feedthrough
rlabel pdiffusion 1886 -1391 1886 -1391 0 feedthrough
rlabel pdiffusion 1893 -1391 1893 -1391 0 feedthrough
rlabel pdiffusion 1900 -1391 1900 -1391 0 feedthrough
rlabel pdiffusion 1907 -1391 1907 -1391 0 feedthrough
rlabel pdiffusion 1914 -1391 1914 -1391 0 cellNo=245
rlabel pdiffusion 1921 -1391 1921 -1391 0 feedthrough
rlabel pdiffusion 1928 -1391 1928 -1391 0 feedthrough
rlabel pdiffusion 1935 -1391 1935 -1391 0 feedthrough
rlabel pdiffusion 1942 -1391 1942 -1391 0 feedthrough
rlabel pdiffusion 1949 -1391 1949 -1391 0 feedthrough
rlabel pdiffusion 1970 -1391 1970 -1391 0 feedthrough
rlabel pdiffusion 1977 -1391 1977 -1391 0 feedthrough
rlabel pdiffusion 1984 -1391 1984 -1391 0 feedthrough
rlabel pdiffusion 1991 -1391 1991 -1391 0 feedthrough
rlabel pdiffusion 1998 -1391 1998 -1391 0 feedthrough
rlabel pdiffusion 3 -1522 3 -1522 0 feedthrough
rlabel pdiffusion 10 -1522 10 -1522 0 feedthrough
rlabel pdiffusion 17 -1522 17 -1522 0 feedthrough
rlabel pdiffusion 24 -1522 24 -1522 0 feedthrough
rlabel pdiffusion 31 -1522 31 -1522 0 feedthrough
rlabel pdiffusion 38 -1522 38 -1522 0 feedthrough
rlabel pdiffusion 45 -1522 45 -1522 0 cellNo=152
rlabel pdiffusion 52 -1522 52 -1522 0 feedthrough
rlabel pdiffusion 59 -1522 59 -1522 0 cellNo=417
rlabel pdiffusion 66 -1522 66 -1522 0 feedthrough
rlabel pdiffusion 73 -1522 73 -1522 0 feedthrough
rlabel pdiffusion 80 -1522 80 -1522 0 cellNo=59
rlabel pdiffusion 87 -1522 87 -1522 0 feedthrough
rlabel pdiffusion 94 -1522 94 -1522 0 feedthrough
rlabel pdiffusion 101 -1522 101 -1522 0 feedthrough
rlabel pdiffusion 108 -1522 108 -1522 0 feedthrough
rlabel pdiffusion 115 -1522 115 -1522 0 feedthrough
rlabel pdiffusion 122 -1522 122 -1522 0 feedthrough
rlabel pdiffusion 129 -1522 129 -1522 0 feedthrough
rlabel pdiffusion 136 -1522 136 -1522 0 feedthrough
rlabel pdiffusion 143 -1522 143 -1522 0 cellNo=41
rlabel pdiffusion 150 -1522 150 -1522 0 feedthrough
rlabel pdiffusion 157 -1522 157 -1522 0 feedthrough
rlabel pdiffusion 164 -1522 164 -1522 0 feedthrough
rlabel pdiffusion 171 -1522 171 -1522 0 feedthrough
rlabel pdiffusion 178 -1522 178 -1522 0 feedthrough
rlabel pdiffusion 185 -1522 185 -1522 0 feedthrough
rlabel pdiffusion 192 -1522 192 -1522 0 cellNo=331
rlabel pdiffusion 199 -1522 199 -1522 0 feedthrough
rlabel pdiffusion 206 -1522 206 -1522 0 feedthrough
rlabel pdiffusion 213 -1522 213 -1522 0 cellNo=16
rlabel pdiffusion 220 -1522 220 -1522 0 feedthrough
rlabel pdiffusion 227 -1522 227 -1522 0 feedthrough
rlabel pdiffusion 234 -1522 234 -1522 0 cellNo=612
rlabel pdiffusion 241 -1522 241 -1522 0 cellNo=837
rlabel pdiffusion 248 -1522 248 -1522 0 feedthrough
rlabel pdiffusion 255 -1522 255 -1522 0 feedthrough
rlabel pdiffusion 262 -1522 262 -1522 0 feedthrough
rlabel pdiffusion 269 -1522 269 -1522 0 feedthrough
rlabel pdiffusion 276 -1522 276 -1522 0 feedthrough
rlabel pdiffusion 283 -1522 283 -1522 0 feedthrough
rlabel pdiffusion 290 -1522 290 -1522 0 feedthrough
rlabel pdiffusion 297 -1522 297 -1522 0 feedthrough
rlabel pdiffusion 304 -1522 304 -1522 0 feedthrough
rlabel pdiffusion 311 -1522 311 -1522 0 feedthrough
rlabel pdiffusion 318 -1522 318 -1522 0 feedthrough
rlabel pdiffusion 325 -1522 325 -1522 0 feedthrough
rlabel pdiffusion 332 -1522 332 -1522 0 feedthrough
rlabel pdiffusion 339 -1522 339 -1522 0 feedthrough
rlabel pdiffusion 346 -1522 346 -1522 0 feedthrough
rlabel pdiffusion 353 -1522 353 -1522 0 feedthrough
rlabel pdiffusion 360 -1522 360 -1522 0 feedthrough
rlabel pdiffusion 367 -1522 367 -1522 0 feedthrough
rlabel pdiffusion 374 -1522 374 -1522 0 feedthrough
rlabel pdiffusion 381 -1522 381 -1522 0 feedthrough
rlabel pdiffusion 388 -1522 388 -1522 0 feedthrough
rlabel pdiffusion 395 -1522 395 -1522 0 feedthrough
rlabel pdiffusion 402 -1522 402 -1522 0 feedthrough
rlabel pdiffusion 409 -1522 409 -1522 0 feedthrough
rlabel pdiffusion 416 -1522 416 -1522 0 feedthrough
rlabel pdiffusion 423 -1522 423 -1522 0 feedthrough
rlabel pdiffusion 430 -1522 430 -1522 0 feedthrough
rlabel pdiffusion 437 -1522 437 -1522 0 feedthrough
rlabel pdiffusion 444 -1522 444 -1522 0 feedthrough
rlabel pdiffusion 451 -1522 451 -1522 0 feedthrough
rlabel pdiffusion 458 -1522 458 -1522 0 feedthrough
rlabel pdiffusion 465 -1522 465 -1522 0 feedthrough
rlabel pdiffusion 472 -1522 472 -1522 0 feedthrough
rlabel pdiffusion 479 -1522 479 -1522 0 feedthrough
rlabel pdiffusion 486 -1522 486 -1522 0 feedthrough
rlabel pdiffusion 493 -1522 493 -1522 0 feedthrough
rlabel pdiffusion 500 -1522 500 -1522 0 cellNo=966
rlabel pdiffusion 507 -1522 507 -1522 0 feedthrough
rlabel pdiffusion 514 -1522 514 -1522 0 feedthrough
rlabel pdiffusion 521 -1522 521 -1522 0 feedthrough
rlabel pdiffusion 528 -1522 528 -1522 0 feedthrough
rlabel pdiffusion 535 -1522 535 -1522 0 feedthrough
rlabel pdiffusion 542 -1522 542 -1522 0 feedthrough
rlabel pdiffusion 549 -1522 549 -1522 0 feedthrough
rlabel pdiffusion 556 -1522 556 -1522 0 feedthrough
rlabel pdiffusion 563 -1522 563 -1522 0 feedthrough
rlabel pdiffusion 570 -1522 570 -1522 0 feedthrough
rlabel pdiffusion 577 -1522 577 -1522 0 feedthrough
rlabel pdiffusion 584 -1522 584 -1522 0 feedthrough
rlabel pdiffusion 591 -1522 591 -1522 0 cellNo=307
rlabel pdiffusion 598 -1522 598 -1522 0 feedthrough
rlabel pdiffusion 605 -1522 605 -1522 0 feedthrough
rlabel pdiffusion 612 -1522 612 -1522 0 feedthrough
rlabel pdiffusion 619 -1522 619 -1522 0 feedthrough
rlabel pdiffusion 626 -1522 626 -1522 0 cellNo=392
rlabel pdiffusion 633 -1522 633 -1522 0 feedthrough
rlabel pdiffusion 640 -1522 640 -1522 0 feedthrough
rlabel pdiffusion 647 -1522 647 -1522 0 feedthrough
rlabel pdiffusion 654 -1522 654 -1522 0 feedthrough
rlabel pdiffusion 661 -1522 661 -1522 0 cellNo=103
rlabel pdiffusion 668 -1522 668 -1522 0 cellNo=988
rlabel pdiffusion 675 -1522 675 -1522 0 feedthrough
rlabel pdiffusion 682 -1522 682 -1522 0 feedthrough
rlabel pdiffusion 689 -1522 689 -1522 0 feedthrough
rlabel pdiffusion 696 -1522 696 -1522 0 feedthrough
rlabel pdiffusion 703 -1522 703 -1522 0 feedthrough
rlabel pdiffusion 710 -1522 710 -1522 0 cellNo=552
rlabel pdiffusion 717 -1522 717 -1522 0 feedthrough
rlabel pdiffusion 724 -1522 724 -1522 0 feedthrough
rlabel pdiffusion 731 -1522 731 -1522 0 feedthrough
rlabel pdiffusion 738 -1522 738 -1522 0 feedthrough
rlabel pdiffusion 745 -1522 745 -1522 0 feedthrough
rlabel pdiffusion 752 -1522 752 -1522 0 cellNo=657
rlabel pdiffusion 759 -1522 759 -1522 0 feedthrough
rlabel pdiffusion 766 -1522 766 -1522 0 feedthrough
rlabel pdiffusion 773 -1522 773 -1522 0 feedthrough
rlabel pdiffusion 780 -1522 780 -1522 0 feedthrough
rlabel pdiffusion 787 -1522 787 -1522 0 feedthrough
rlabel pdiffusion 794 -1522 794 -1522 0 feedthrough
rlabel pdiffusion 801 -1522 801 -1522 0 feedthrough
rlabel pdiffusion 808 -1522 808 -1522 0 feedthrough
rlabel pdiffusion 815 -1522 815 -1522 0 feedthrough
rlabel pdiffusion 822 -1522 822 -1522 0 feedthrough
rlabel pdiffusion 829 -1522 829 -1522 0 feedthrough
rlabel pdiffusion 836 -1522 836 -1522 0 feedthrough
rlabel pdiffusion 843 -1522 843 -1522 0 feedthrough
rlabel pdiffusion 850 -1522 850 -1522 0 feedthrough
rlabel pdiffusion 857 -1522 857 -1522 0 feedthrough
rlabel pdiffusion 864 -1522 864 -1522 0 feedthrough
rlabel pdiffusion 871 -1522 871 -1522 0 feedthrough
rlabel pdiffusion 878 -1522 878 -1522 0 feedthrough
rlabel pdiffusion 885 -1522 885 -1522 0 feedthrough
rlabel pdiffusion 892 -1522 892 -1522 0 feedthrough
rlabel pdiffusion 899 -1522 899 -1522 0 feedthrough
rlabel pdiffusion 906 -1522 906 -1522 0 feedthrough
rlabel pdiffusion 913 -1522 913 -1522 0 feedthrough
rlabel pdiffusion 920 -1522 920 -1522 0 cellNo=363
rlabel pdiffusion 927 -1522 927 -1522 0 feedthrough
rlabel pdiffusion 934 -1522 934 -1522 0 feedthrough
rlabel pdiffusion 941 -1522 941 -1522 0 feedthrough
rlabel pdiffusion 948 -1522 948 -1522 0 cellNo=598
rlabel pdiffusion 955 -1522 955 -1522 0 cellNo=85
rlabel pdiffusion 962 -1522 962 -1522 0 cellNo=842
rlabel pdiffusion 969 -1522 969 -1522 0 feedthrough
rlabel pdiffusion 976 -1522 976 -1522 0 feedthrough
rlabel pdiffusion 983 -1522 983 -1522 0 cellNo=54
rlabel pdiffusion 990 -1522 990 -1522 0 feedthrough
rlabel pdiffusion 997 -1522 997 -1522 0 feedthrough
rlabel pdiffusion 1004 -1522 1004 -1522 0 cellNo=559
rlabel pdiffusion 1011 -1522 1011 -1522 0 feedthrough
rlabel pdiffusion 1018 -1522 1018 -1522 0 feedthrough
rlabel pdiffusion 1025 -1522 1025 -1522 0 feedthrough
rlabel pdiffusion 1032 -1522 1032 -1522 0 feedthrough
rlabel pdiffusion 1039 -1522 1039 -1522 0 feedthrough
rlabel pdiffusion 1046 -1522 1046 -1522 0 feedthrough
rlabel pdiffusion 1053 -1522 1053 -1522 0 feedthrough
rlabel pdiffusion 1060 -1522 1060 -1522 0 feedthrough
rlabel pdiffusion 1067 -1522 1067 -1522 0 cellNo=567
rlabel pdiffusion 1074 -1522 1074 -1522 0 feedthrough
rlabel pdiffusion 1081 -1522 1081 -1522 0 feedthrough
rlabel pdiffusion 1088 -1522 1088 -1522 0 feedthrough
rlabel pdiffusion 1095 -1522 1095 -1522 0 feedthrough
rlabel pdiffusion 1102 -1522 1102 -1522 0 cellNo=809
rlabel pdiffusion 1109 -1522 1109 -1522 0 cellNo=254
rlabel pdiffusion 1116 -1522 1116 -1522 0 cellNo=706
rlabel pdiffusion 1123 -1522 1123 -1522 0 feedthrough
rlabel pdiffusion 1130 -1522 1130 -1522 0 cellNo=261
rlabel pdiffusion 1137 -1522 1137 -1522 0 feedthrough
rlabel pdiffusion 1144 -1522 1144 -1522 0 feedthrough
rlabel pdiffusion 1151 -1522 1151 -1522 0 feedthrough
rlabel pdiffusion 1158 -1522 1158 -1522 0 cellNo=823
rlabel pdiffusion 1165 -1522 1165 -1522 0 feedthrough
rlabel pdiffusion 1172 -1522 1172 -1522 0 feedthrough
rlabel pdiffusion 1179 -1522 1179 -1522 0 feedthrough
rlabel pdiffusion 1186 -1522 1186 -1522 0 feedthrough
rlabel pdiffusion 1193 -1522 1193 -1522 0 cellNo=532
rlabel pdiffusion 1200 -1522 1200 -1522 0 feedthrough
rlabel pdiffusion 1207 -1522 1207 -1522 0 feedthrough
rlabel pdiffusion 1214 -1522 1214 -1522 0 feedthrough
rlabel pdiffusion 1221 -1522 1221 -1522 0 feedthrough
rlabel pdiffusion 1228 -1522 1228 -1522 0 feedthrough
rlabel pdiffusion 1235 -1522 1235 -1522 0 feedthrough
rlabel pdiffusion 1242 -1522 1242 -1522 0 feedthrough
rlabel pdiffusion 1249 -1522 1249 -1522 0 feedthrough
rlabel pdiffusion 1256 -1522 1256 -1522 0 feedthrough
rlabel pdiffusion 1263 -1522 1263 -1522 0 cellNo=364
rlabel pdiffusion 1270 -1522 1270 -1522 0 feedthrough
rlabel pdiffusion 1277 -1522 1277 -1522 0 feedthrough
rlabel pdiffusion 1284 -1522 1284 -1522 0 feedthrough
rlabel pdiffusion 1291 -1522 1291 -1522 0 feedthrough
rlabel pdiffusion 1298 -1522 1298 -1522 0 feedthrough
rlabel pdiffusion 1305 -1522 1305 -1522 0 cellNo=934
rlabel pdiffusion 1312 -1522 1312 -1522 0 feedthrough
rlabel pdiffusion 1319 -1522 1319 -1522 0 feedthrough
rlabel pdiffusion 1326 -1522 1326 -1522 0 feedthrough
rlabel pdiffusion 1333 -1522 1333 -1522 0 cellNo=201
rlabel pdiffusion 1340 -1522 1340 -1522 0 feedthrough
rlabel pdiffusion 1347 -1522 1347 -1522 0 feedthrough
rlabel pdiffusion 1354 -1522 1354 -1522 0 feedthrough
rlabel pdiffusion 1361 -1522 1361 -1522 0 feedthrough
rlabel pdiffusion 1368 -1522 1368 -1522 0 feedthrough
rlabel pdiffusion 1375 -1522 1375 -1522 0 feedthrough
rlabel pdiffusion 1382 -1522 1382 -1522 0 feedthrough
rlabel pdiffusion 1389 -1522 1389 -1522 0 feedthrough
rlabel pdiffusion 1396 -1522 1396 -1522 0 feedthrough
rlabel pdiffusion 1403 -1522 1403 -1522 0 feedthrough
rlabel pdiffusion 1410 -1522 1410 -1522 0 feedthrough
rlabel pdiffusion 1417 -1522 1417 -1522 0 feedthrough
rlabel pdiffusion 1424 -1522 1424 -1522 0 feedthrough
rlabel pdiffusion 1431 -1522 1431 -1522 0 feedthrough
rlabel pdiffusion 1438 -1522 1438 -1522 0 feedthrough
rlabel pdiffusion 1445 -1522 1445 -1522 0 feedthrough
rlabel pdiffusion 1452 -1522 1452 -1522 0 feedthrough
rlabel pdiffusion 1459 -1522 1459 -1522 0 feedthrough
rlabel pdiffusion 1466 -1522 1466 -1522 0 feedthrough
rlabel pdiffusion 1473 -1522 1473 -1522 0 feedthrough
rlabel pdiffusion 1480 -1522 1480 -1522 0 feedthrough
rlabel pdiffusion 1487 -1522 1487 -1522 0 feedthrough
rlabel pdiffusion 1494 -1522 1494 -1522 0 feedthrough
rlabel pdiffusion 1501 -1522 1501 -1522 0 feedthrough
rlabel pdiffusion 1508 -1522 1508 -1522 0 feedthrough
rlabel pdiffusion 1515 -1522 1515 -1522 0 feedthrough
rlabel pdiffusion 1522 -1522 1522 -1522 0 feedthrough
rlabel pdiffusion 1529 -1522 1529 -1522 0 feedthrough
rlabel pdiffusion 1536 -1522 1536 -1522 0 feedthrough
rlabel pdiffusion 1543 -1522 1543 -1522 0 feedthrough
rlabel pdiffusion 1550 -1522 1550 -1522 0 feedthrough
rlabel pdiffusion 1557 -1522 1557 -1522 0 feedthrough
rlabel pdiffusion 1564 -1522 1564 -1522 0 feedthrough
rlabel pdiffusion 1571 -1522 1571 -1522 0 feedthrough
rlabel pdiffusion 1578 -1522 1578 -1522 0 feedthrough
rlabel pdiffusion 1585 -1522 1585 -1522 0 feedthrough
rlabel pdiffusion 1592 -1522 1592 -1522 0 feedthrough
rlabel pdiffusion 1599 -1522 1599 -1522 0 feedthrough
rlabel pdiffusion 1606 -1522 1606 -1522 0 feedthrough
rlabel pdiffusion 1613 -1522 1613 -1522 0 feedthrough
rlabel pdiffusion 1620 -1522 1620 -1522 0 feedthrough
rlabel pdiffusion 1627 -1522 1627 -1522 0 feedthrough
rlabel pdiffusion 1634 -1522 1634 -1522 0 feedthrough
rlabel pdiffusion 1641 -1522 1641 -1522 0 feedthrough
rlabel pdiffusion 1648 -1522 1648 -1522 0 feedthrough
rlabel pdiffusion 1655 -1522 1655 -1522 0 feedthrough
rlabel pdiffusion 1662 -1522 1662 -1522 0 feedthrough
rlabel pdiffusion 1669 -1522 1669 -1522 0 feedthrough
rlabel pdiffusion 1676 -1522 1676 -1522 0 feedthrough
rlabel pdiffusion 1683 -1522 1683 -1522 0 feedthrough
rlabel pdiffusion 1690 -1522 1690 -1522 0 feedthrough
rlabel pdiffusion 1697 -1522 1697 -1522 0 feedthrough
rlabel pdiffusion 1704 -1522 1704 -1522 0 feedthrough
rlabel pdiffusion 1711 -1522 1711 -1522 0 feedthrough
rlabel pdiffusion 1718 -1522 1718 -1522 0 feedthrough
rlabel pdiffusion 1725 -1522 1725 -1522 0 feedthrough
rlabel pdiffusion 1732 -1522 1732 -1522 0 feedthrough
rlabel pdiffusion 1739 -1522 1739 -1522 0 feedthrough
rlabel pdiffusion 1746 -1522 1746 -1522 0 feedthrough
rlabel pdiffusion 1753 -1522 1753 -1522 0 feedthrough
rlabel pdiffusion 1760 -1522 1760 -1522 0 feedthrough
rlabel pdiffusion 1767 -1522 1767 -1522 0 feedthrough
rlabel pdiffusion 1774 -1522 1774 -1522 0 feedthrough
rlabel pdiffusion 1781 -1522 1781 -1522 0 feedthrough
rlabel pdiffusion 1788 -1522 1788 -1522 0 feedthrough
rlabel pdiffusion 1795 -1522 1795 -1522 0 feedthrough
rlabel pdiffusion 1802 -1522 1802 -1522 0 feedthrough
rlabel pdiffusion 1809 -1522 1809 -1522 0 feedthrough
rlabel pdiffusion 1816 -1522 1816 -1522 0 feedthrough
rlabel pdiffusion 1823 -1522 1823 -1522 0 feedthrough
rlabel pdiffusion 1830 -1522 1830 -1522 0 feedthrough
rlabel pdiffusion 1837 -1522 1837 -1522 0 feedthrough
rlabel pdiffusion 1844 -1522 1844 -1522 0 feedthrough
rlabel pdiffusion 1851 -1522 1851 -1522 0 feedthrough
rlabel pdiffusion 1858 -1522 1858 -1522 0 feedthrough
rlabel pdiffusion 1865 -1522 1865 -1522 0 feedthrough
rlabel pdiffusion 1872 -1522 1872 -1522 0 feedthrough
rlabel pdiffusion 1879 -1522 1879 -1522 0 feedthrough
rlabel pdiffusion 1886 -1522 1886 -1522 0 feedthrough
rlabel pdiffusion 1893 -1522 1893 -1522 0 feedthrough
rlabel pdiffusion 1900 -1522 1900 -1522 0 feedthrough
rlabel pdiffusion 1907 -1522 1907 -1522 0 feedthrough
rlabel pdiffusion 1914 -1522 1914 -1522 0 feedthrough
rlabel pdiffusion 1921 -1522 1921 -1522 0 feedthrough
rlabel pdiffusion 1928 -1522 1928 -1522 0 feedthrough
rlabel pdiffusion 1935 -1522 1935 -1522 0 feedthrough
rlabel pdiffusion 1942 -1522 1942 -1522 0 feedthrough
rlabel pdiffusion 1949 -1522 1949 -1522 0 feedthrough
rlabel pdiffusion 1956 -1522 1956 -1522 0 feedthrough
rlabel pdiffusion 1963 -1522 1963 -1522 0 feedthrough
rlabel pdiffusion 1970 -1522 1970 -1522 0 cellNo=521
rlabel pdiffusion 1977 -1522 1977 -1522 0 cellNo=488
rlabel pdiffusion 1984 -1522 1984 -1522 0 feedthrough
rlabel pdiffusion 1991 -1522 1991 -1522 0 feedthrough
rlabel pdiffusion 1998 -1522 1998 -1522 0 cellNo=232
rlabel pdiffusion 2005 -1522 2005 -1522 0 cellNo=999
rlabel pdiffusion 2012 -1522 2012 -1522 0 feedthrough
rlabel pdiffusion 2019 -1522 2019 -1522 0 feedthrough
rlabel pdiffusion 2026 -1522 2026 -1522 0 feedthrough
rlabel pdiffusion 3 -1649 3 -1649 0 feedthrough
rlabel pdiffusion 10 -1649 10 -1649 0 feedthrough
rlabel pdiffusion 17 -1649 17 -1649 0 feedthrough
rlabel pdiffusion 24 -1649 24 -1649 0 feedthrough
rlabel pdiffusion 31 -1649 31 -1649 0 feedthrough
rlabel pdiffusion 38 -1649 38 -1649 0 feedthrough
rlabel pdiffusion 45 -1649 45 -1649 0 feedthrough
rlabel pdiffusion 52 -1649 52 -1649 0 feedthrough
rlabel pdiffusion 59 -1649 59 -1649 0 feedthrough
rlabel pdiffusion 66 -1649 66 -1649 0 cellNo=84
rlabel pdiffusion 73 -1649 73 -1649 0 feedthrough
rlabel pdiffusion 80 -1649 80 -1649 0 cellNo=890
rlabel pdiffusion 87 -1649 87 -1649 0 cellNo=807
rlabel pdiffusion 94 -1649 94 -1649 0 feedthrough
rlabel pdiffusion 101 -1649 101 -1649 0 feedthrough
rlabel pdiffusion 108 -1649 108 -1649 0 feedthrough
rlabel pdiffusion 115 -1649 115 -1649 0 cellNo=692
rlabel pdiffusion 122 -1649 122 -1649 0 feedthrough
rlabel pdiffusion 129 -1649 129 -1649 0 feedthrough
rlabel pdiffusion 136 -1649 136 -1649 0 feedthrough
rlabel pdiffusion 143 -1649 143 -1649 0 cellNo=268
rlabel pdiffusion 150 -1649 150 -1649 0 feedthrough
rlabel pdiffusion 157 -1649 157 -1649 0 feedthrough
rlabel pdiffusion 164 -1649 164 -1649 0 feedthrough
rlabel pdiffusion 171 -1649 171 -1649 0 cellNo=856
rlabel pdiffusion 178 -1649 178 -1649 0 cellNo=309
rlabel pdiffusion 185 -1649 185 -1649 0 feedthrough
rlabel pdiffusion 192 -1649 192 -1649 0 feedthrough
rlabel pdiffusion 199 -1649 199 -1649 0 feedthrough
rlabel pdiffusion 206 -1649 206 -1649 0 feedthrough
rlabel pdiffusion 213 -1649 213 -1649 0 feedthrough
rlabel pdiffusion 220 -1649 220 -1649 0 feedthrough
rlabel pdiffusion 227 -1649 227 -1649 0 feedthrough
rlabel pdiffusion 234 -1649 234 -1649 0 feedthrough
rlabel pdiffusion 241 -1649 241 -1649 0 feedthrough
rlabel pdiffusion 248 -1649 248 -1649 0 feedthrough
rlabel pdiffusion 255 -1649 255 -1649 0 feedthrough
rlabel pdiffusion 262 -1649 262 -1649 0 feedthrough
rlabel pdiffusion 269 -1649 269 -1649 0 feedthrough
rlabel pdiffusion 276 -1649 276 -1649 0 feedthrough
rlabel pdiffusion 283 -1649 283 -1649 0 feedthrough
rlabel pdiffusion 290 -1649 290 -1649 0 feedthrough
rlabel pdiffusion 297 -1649 297 -1649 0 feedthrough
rlabel pdiffusion 304 -1649 304 -1649 0 feedthrough
rlabel pdiffusion 311 -1649 311 -1649 0 feedthrough
rlabel pdiffusion 318 -1649 318 -1649 0 feedthrough
rlabel pdiffusion 325 -1649 325 -1649 0 feedthrough
rlabel pdiffusion 332 -1649 332 -1649 0 feedthrough
rlabel pdiffusion 339 -1649 339 -1649 0 feedthrough
rlabel pdiffusion 346 -1649 346 -1649 0 feedthrough
rlabel pdiffusion 353 -1649 353 -1649 0 feedthrough
rlabel pdiffusion 360 -1649 360 -1649 0 feedthrough
rlabel pdiffusion 367 -1649 367 -1649 0 feedthrough
rlabel pdiffusion 374 -1649 374 -1649 0 feedthrough
rlabel pdiffusion 381 -1649 381 -1649 0 feedthrough
rlabel pdiffusion 388 -1649 388 -1649 0 feedthrough
rlabel pdiffusion 395 -1649 395 -1649 0 cellNo=40
rlabel pdiffusion 402 -1649 402 -1649 0 feedthrough
rlabel pdiffusion 409 -1649 409 -1649 0 feedthrough
rlabel pdiffusion 416 -1649 416 -1649 0 cellNo=25
rlabel pdiffusion 423 -1649 423 -1649 0 feedthrough
rlabel pdiffusion 430 -1649 430 -1649 0 feedthrough
rlabel pdiffusion 437 -1649 437 -1649 0 feedthrough
rlabel pdiffusion 444 -1649 444 -1649 0 feedthrough
rlabel pdiffusion 451 -1649 451 -1649 0 feedthrough
rlabel pdiffusion 458 -1649 458 -1649 0 feedthrough
rlabel pdiffusion 465 -1649 465 -1649 0 feedthrough
rlabel pdiffusion 472 -1649 472 -1649 0 feedthrough
rlabel pdiffusion 479 -1649 479 -1649 0 feedthrough
rlabel pdiffusion 486 -1649 486 -1649 0 feedthrough
rlabel pdiffusion 493 -1649 493 -1649 0 feedthrough
rlabel pdiffusion 500 -1649 500 -1649 0 feedthrough
rlabel pdiffusion 507 -1649 507 -1649 0 feedthrough
rlabel pdiffusion 514 -1649 514 -1649 0 feedthrough
rlabel pdiffusion 521 -1649 521 -1649 0 feedthrough
rlabel pdiffusion 528 -1649 528 -1649 0 feedthrough
rlabel pdiffusion 535 -1649 535 -1649 0 feedthrough
rlabel pdiffusion 542 -1649 542 -1649 0 cellNo=767
rlabel pdiffusion 549 -1649 549 -1649 0 feedthrough
rlabel pdiffusion 556 -1649 556 -1649 0 feedthrough
rlabel pdiffusion 563 -1649 563 -1649 0 feedthrough
rlabel pdiffusion 570 -1649 570 -1649 0 feedthrough
rlabel pdiffusion 577 -1649 577 -1649 0 feedthrough
rlabel pdiffusion 584 -1649 584 -1649 0 feedthrough
rlabel pdiffusion 591 -1649 591 -1649 0 feedthrough
rlabel pdiffusion 598 -1649 598 -1649 0 feedthrough
rlabel pdiffusion 605 -1649 605 -1649 0 feedthrough
rlabel pdiffusion 612 -1649 612 -1649 0 feedthrough
rlabel pdiffusion 619 -1649 619 -1649 0 feedthrough
rlabel pdiffusion 626 -1649 626 -1649 0 feedthrough
rlabel pdiffusion 633 -1649 633 -1649 0 feedthrough
rlabel pdiffusion 640 -1649 640 -1649 0 feedthrough
rlabel pdiffusion 647 -1649 647 -1649 0 feedthrough
rlabel pdiffusion 654 -1649 654 -1649 0 feedthrough
rlabel pdiffusion 661 -1649 661 -1649 0 cellNo=265
rlabel pdiffusion 668 -1649 668 -1649 0 cellNo=236
rlabel pdiffusion 675 -1649 675 -1649 0 feedthrough
rlabel pdiffusion 682 -1649 682 -1649 0 feedthrough
rlabel pdiffusion 689 -1649 689 -1649 0 feedthrough
rlabel pdiffusion 696 -1649 696 -1649 0 cellNo=614
rlabel pdiffusion 703 -1649 703 -1649 0 feedthrough
rlabel pdiffusion 710 -1649 710 -1649 0 cellNo=705
rlabel pdiffusion 717 -1649 717 -1649 0 feedthrough
rlabel pdiffusion 724 -1649 724 -1649 0 feedthrough
rlabel pdiffusion 731 -1649 731 -1649 0 feedthrough
rlabel pdiffusion 738 -1649 738 -1649 0 cellNo=889
rlabel pdiffusion 745 -1649 745 -1649 0 feedthrough
rlabel pdiffusion 752 -1649 752 -1649 0 feedthrough
rlabel pdiffusion 759 -1649 759 -1649 0 feedthrough
rlabel pdiffusion 766 -1649 766 -1649 0 cellNo=276
rlabel pdiffusion 773 -1649 773 -1649 0 feedthrough
rlabel pdiffusion 780 -1649 780 -1649 0 feedthrough
rlabel pdiffusion 787 -1649 787 -1649 0 feedthrough
rlabel pdiffusion 794 -1649 794 -1649 0 feedthrough
rlabel pdiffusion 801 -1649 801 -1649 0 feedthrough
rlabel pdiffusion 808 -1649 808 -1649 0 feedthrough
rlabel pdiffusion 815 -1649 815 -1649 0 cellNo=144
rlabel pdiffusion 822 -1649 822 -1649 0 feedthrough
rlabel pdiffusion 829 -1649 829 -1649 0 cellNo=820
rlabel pdiffusion 836 -1649 836 -1649 0 feedthrough
rlabel pdiffusion 843 -1649 843 -1649 0 feedthrough
rlabel pdiffusion 850 -1649 850 -1649 0 feedthrough
rlabel pdiffusion 857 -1649 857 -1649 0 feedthrough
rlabel pdiffusion 864 -1649 864 -1649 0 feedthrough
rlabel pdiffusion 871 -1649 871 -1649 0 feedthrough
rlabel pdiffusion 878 -1649 878 -1649 0 feedthrough
rlabel pdiffusion 885 -1649 885 -1649 0 feedthrough
rlabel pdiffusion 892 -1649 892 -1649 0 feedthrough
rlabel pdiffusion 899 -1649 899 -1649 0 feedthrough
rlabel pdiffusion 906 -1649 906 -1649 0 feedthrough
rlabel pdiffusion 913 -1649 913 -1649 0 feedthrough
rlabel pdiffusion 920 -1649 920 -1649 0 cellNo=446
rlabel pdiffusion 927 -1649 927 -1649 0 feedthrough
rlabel pdiffusion 934 -1649 934 -1649 0 feedthrough
rlabel pdiffusion 941 -1649 941 -1649 0 cellNo=235
rlabel pdiffusion 948 -1649 948 -1649 0 feedthrough
rlabel pdiffusion 955 -1649 955 -1649 0 feedthrough
rlabel pdiffusion 962 -1649 962 -1649 0 feedthrough
rlabel pdiffusion 969 -1649 969 -1649 0 cellNo=658
rlabel pdiffusion 976 -1649 976 -1649 0 feedthrough
rlabel pdiffusion 983 -1649 983 -1649 0 feedthrough
rlabel pdiffusion 990 -1649 990 -1649 0 feedthrough
rlabel pdiffusion 997 -1649 997 -1649 0 feedthrough
rlabel pdiffusion 1004 -1649 1004 -1649 0 feedthrough
rlabel pdiffusion 1011 -1649 1011 -1649 0 feedthrough
rlabel pdiffusion 1018 -1649 1018 -1649 0 feedthrough
rlabel pdiffusion 1025 -1649 1025 -1649 0 feedthrough
rlabel pdiffusion 1032 -1649 1032 -1649 0 feedthrough
rlabel pdiffusion 1039 -1649 1039 -1649 0 cellNo=45
rlabel pdiffusion 1046 -1649 1046 -1649 0 feedthrough
rlabel pdiffusion 1053 -1649 1053 -1649 0 cellNo=819
rlabel pdiffusion 1060 -1649 1060 -1649 0 feedthrough
rlabel pdiffusion 1067 -1649 1067 -1649 0 feedthrough
rlabel pdiffusion 1074 -1649 1074 -1649 0 feedthrough
rlabel pdiffusion 1081 -1649 1081 -1649 0 feedthrough
rlabel pdiffusion 1088 -1649 1088 -1649 0 cellNo=743
rlabel pdiffusion 1095 -1649 1095 -1649 0 feedthrough
rlabel pdiffusion 1102 -1649 1102 -1649 0 feedthrough
rlabel pdiffusion 1109 -1649 1109 -1649 0 feedthrough
rlabel pdiffusion 1116 -1649 1116 -1649 0 feedthrough
rlabel pdiffusion 1123 -1649 1123 -1649 0 feedthrough
rlabel pdiffusion 1130 -1649 1130 -1649 0 cellNo=990
rlabel pdiffusion 1137 -1649 1137 -1649 0 feedthrough
rlabel pdiffusion 1144 -1649 1144 -1649 0 feedthrough
rlabel pdiffusion 1151 -1649 1151 -1649 0 feedthrough
rlabel pdiffusion 1158 -1649 1158 -1649 0 feedthrough
rlabel pdiffusion 1165 -1649 1165 -1649 0 feedthrough
rlabel pdiffusion 1172 -1649 1172 -1649 0 feedthrough
rlabel pdiffusion 1179 -1649 1179 -1649 0 feedthrough
rlabel pdiffusion 1186 -1649 1186 -1649 0 feedthrough
rlabel pdiffusion 1193 -1649 1193 -1649 0 feedthrough
rlabel pdiffusion 1200 -1649 1200 -1649 0 feedthrough
rlabel pdiffusion 1207 -1649 1207 -1649 0 cellNo=110
rlabel pdiffusion 1214 -1649 1214 -1649 0 feedthrough
rlabel pdiffusion 1221 -1649 1221 -1649 0 feedthrough
rlabel pdiffusion 1228 -1649 1228 -1649 0 feedthrough
rlabel pdiffusion 1235 -1649 1235 -1649 0 feedthrough
rlabel pdiffusion 1242 -1649 1242 -1649 0 cellNo=335
rlabel pdiffusion 1249 -1649 1249 -1649 0 feedthrough
rlabel pdiffusion 1256 -1649 1256 -1649 0 feedthrough
rlabel pdiffusion 1263 -1649 1263 -1649 0 feedthrough
rlabel pdiffusion 1270 -1649 1270 -1649 0 feedthrough
rlabel pdiffusion 1277 -1649 1277 -1649 0 feedthrough
rlabel pdiffusion 1284 -1649 1284 -1649 0 cellNo=416
rlabel pdiffusion 1291 -1649 1291 -1649 0 feedthrough
rlabel pdiffusion 1298 -1649 1298 -1649 0 feedthrough
rlabel pdiffusion 1305 -1649 1305 -1649 0 cellNo=450
rlabel pdiffusion 1312 -1649 1312 -1649 0 feedthrough
rlabel pdiffusion 1319 -1649 1319 -1649 0 feedthrough
rlabel pdiffusion 1326 -1649 1326 -1649 0 feedthrough
rlabel pdiffusion 1333 -1649 1333 -1649 0 cellNo=480
rlabel pdiffusion 1340 -1649 1340 -1649 0 feedthrough
rlabel pdiffusion 1347 -1649 1347 -1649 0 feedthrough
rlabel pdiffusion 1354 -1649 1354 -1649 0 cellNo=12
rlabel pdiffusion 1361 -1649 1361 -1649 0 feedthrough
rlabel pdiffusion 1368 -1649 1368 -1649 0 feedthrough
rlabel pdiffusion 1375 -1649 1375 -1649 0 feedthrough
rlabel pdiffusion 1382 -1649 1382 -1649 0 feedthrough
rlabel pdiffusion 1389 -1649 1389 -1649 0 feedthrough
rlabel pdiffusion 1396 -1649 1396 -1649 0 feedthrough
rlabel pdiffusion 1403 -1649 1403 -1649 0 feedthrough
rlabel pdiffusion 1410 -1649 1410 -1649 0 feedthrough
rlabel pdiffusion 1417 -1649 1417 -1649 0 feedthrough
rlabel pdiffusion 1424 -1649 1424 -1649 0 feedthrough
rlabel pdiffusion 1431 -1649 1431 -1649 0 feedthrough
rlabel pdiffusion 1438 -1649 1438 -1649 0 feedthrough
rlabel pdiffusion 1445 -1649 1445 -1649 0 feedthrough
rlabel pdiffusion 1452 -1649 1452 -1649 0 feedthrough
rlabel pdiffusion 1459 -1649 1459 -1649 0 feedthrough
rlabel pdiffusion 1466 -1649 1466 -1649 0 cellNo=473
rlabel pdiffusion 1473 -1649 1473 -1649 0 feedthrough
rlabel pdiffusion 1480 -1649 1480 -1649 0 feedthrough
rlabel pdiffusion 1487 -1649 1487 -1649 0 feedthrough
rlabel pdiffusion 1494 -1649 1494 -1649 0 feedthrough
rlabel pdiffusion 1501 -1649 1501 -1649 0 cellNo=829
rlabel pdiffusion 1508 -1649 1508 -1649 0 feedthrough
rlabel pdiffusion 1515 -1649 1515 -1649 0 feedthrough
rlabel pdiffusion 1522 -1649 1522 -1649 0 feedthrough
rlabel pdiffusion 1529 -1649 1529 -1649 0 feedthrough
rlabel pdiffusion 1536 -1649 1536 -1649 0 feedthrough
rlabel pdiffusion 1543 -1649 1543 -1649 0 feedthrough
rlabel pdiffusion 1550 -1649 1550 -1649 0 feedthrough
rlabel pdiffusion 1557 -1649 1557 -1649 0 feedthrough
rlabel pdiffusion 1564 -1649 1564 -1649 0 feedthrough
rlabel pdiffusion 1571 -1649 1571 -1649 0 feedthrough
rlabel pdiffusion 1578 -1649 1578 -1649 0 feedthrough
rlabel pdiffusion 1585 -1649 1585 -1649 0 feedthrough
rlabel pdiffusion 1592 -1649 1592 -1649 0 feedthrough
rlabel pdiffusion 1599 -1649 1599 -1649 0 feedthrough
rlabel pdiffusion 1606 -1649 1606 -1649 0 feedthrough
rlabel pdiffusion 1613 -1649 1613 -1649 0 feedthrough
rlabel pdiffusion 1620 -1649 1620 -1649 0 feedthrough
rlabel pdiffusion 1627 -1649 1627 -1649 0 feedthrough
rlabel pdiffusion 1634 -1649 1634 -1649 0 feedthrough
rlabel pdiffusion 1641 -1649 1641 -1649 0 feedthrough
rlabel pdiffusion 1648 -1649 1648 -1649 0 feedthrough
rlabel pdiffusion 1655 -1649 1655 -1649 0 feedthrough
rlabel pdiffusion 1662 -1649 1662 -1649 0 feedthrough
rlabel pdiffusion 1669 -1649 1669 -1649 0 feedthrough
rlabel pdiffusion 1676 -1649 1676 -1649 0 feedthrough
rlabel pdiffusion 1683 -1649 1683 -1649 0 feedthrough
rlabel pdiffusion 1690 -1649 1690 -1649 0 feedthrough
rlabel pdiffusion 1697 -1649 1697 -1649 0 feedthrough
rlabel pdiffusion 1704 -1649 1704 -1649 0 feedthrough
rlabel pdiffusion 1711 -1649 1711 -1649 0 feedthrough
rlabel pdiffusion 1718 -1649 1718 -1649 0 feedthrough
rlabel pdiffusion 1725 -1649 1725 -1649 0 feedthrough
rlabel pdiffusion 1732 -1649 1732 -1649 0 feedthrough
rlabel pdiffusion 1739 -1649 1739 -1649 0 feedthrough
rlabel pdiffusion 1746 -1649 1746 -1649 0 feedthrough
rlabel pdiffusion 1753 -1649 1753 -1649 0 feedthrough
rlabel pdiffusion 1760 -1649 1760 -1649 0 feedthrough
rlabel pdiffusion 1767 -1649 1767 -1649 0 feedthrough
rlabel pdiffusion 1774 -1649 1774 -1649 0 feedthrough
rlabel pdiffusion 1781 -1649 1781 -1649 0 feedthrough
rlabel pdiffusion 1788 -1649 1788 -1649 0 feedthrough
rlabel pdiffusion 1795 -1649 1795 -1649 0 feedthrough
rlabel pdiffusion 1802 -1649 1802 -1649 0 feedthrough
rlabel pdiffusion 1809 -1649 1809 -1649 0 feedthrough
rlabel pdiffusion 1816 -1649 1816 -1649 0 feedthrough
rlabel pdiffusion 1823 -1649 1823 -1649 0 feedthrough
rlabel pdiffusion 1830 -1649 1830 -1649 0 feedthrough
rlabel pdiffusion 1837 -1649 1837 -1649 0 feedthrough
rlabel pdiffusion 1844 -1649 1844 -1649 0 cellNo=130
rlabel pdiffusion 1851 -1649 1851 -1649 0 feedthrough
rlabel pdiffusion 1858 -1649 1858 -1649 0 feedthrough
rlabel pdiffusion 1865 -1649 1865 -1649 0 feedthrough
rlabel pdiffusion 1872 -1649 1872 -1649 0 feedthrough
rlabel pdiffusion 1879 -1649 1879 -1649 0 cellNo=64
rlabel pdiffusion 1886 -1649 1886 -1649 0 feedthrough
rlabel pdiffusion 1893 -1649 1893 -1649 0 feedthrough
rlabel pdiffusion 1900 -1649 1900 -1649 0 feedthrough
rlabel pdiffusion 1907 -1649 1907 -1649 0 feedthrough
rlabel pdiffusion 1914 -1649 1914 -1649 0 feedthrough
rlabel pdiffusion 1921 -1649 1921 -1649 0 feedthrough
rlabel pdiffusion 1928 -1649 1928 -1649 0 feedthrough
rlabel pdiffusion 1935 -1649 1935 -1649 0 feedthrough
rlabel pdiffusion 1942 -1649 1942 -1649 0 feedthrough
rlabel pdiffusion 1949 -1649 1949 -1649 0 feedthrough
rlabel pdiffusion 1977 -1649 1977 -1649 0 feedthrough
rlabel pdiffusion 2019 -1649 2019 -1649 0 feedthrough
rlabel pdiffusion 10 -1778 10 -1778 0 feedthrough
rlabel pdiffusion 17 -1778 17 -1778 0 feedthrough
rlabel pdiffusion 24 -1778 24 -1778 0 feedthrough
rlabel pdiffusion 31 -1778 31 -1778 0 feedthrough
rlabel pdiffusion 38 -1778 38 -1778 0 feedthrough
rlabel pdiffusion 45 -1778 45 -1778 0 feedthrough
rlabel pdiffusion 52 -1778 52 -1778 0 feedthrough
rlabel pdiffusion 59 -1778 59 -1778 0 feedthrough
rlabel pdiffusion 66 -1778 66 -1778 0 cellNo=379
rlabel pdiffusion 73 -1778 73 -1778 0 feedthrough
rlabel pdiffusion 80 -1778 80 -1778 0 feedthrough
rlabel pdiffusion 87 -1778 87 -1778 0 feedthrough
rlabel pdiffusion 94 -1778 94 -1778 0 feedthrough
rlabel pdiffusion 101 -1778 101 -1778 0 feedthrough
rlabel pdiffusion 108 -1778 108 -1778 0 feedthrough
rlabel pdiffusion 115 -1778 115 -1778 0 feedthrough
rlabel pdiffusion 122 -1778 122 -1778 0 feedthrough
rlabel pdiffusion 129 -1778 129 -1778 0 cellNo=343
rlabel pdiffusion 136 -1778 136 -1778 0 feedthrough
rlabel pdiffusion 143 -1778 143 -1778 0 feedthrough
rlabel pdiffusion 150 -1778 150 -1778 0 feedthrough
rlabel pdiffusion 157 -1778 157 -1778 0 feedthrough
rlabel pdiffusion 164 -1778 164 -1778 0 feedthrough
rlabel pdiffusion 171 -1778 171 -1778 0 feedthrough
rlabel pdiffusion 178 -1778 178 -1778 0 feedthrough
rlabel pdiffusion 185 -1778 185 -1778 0 cellNo=208
rlabel pdiffusion 192 -1778 192 -1778 0 cellNo=169
rlabel pdiffusion 199 -1778 199 -1778 0 cellNo=70
rlabel pdiffusion 206 -1778 206 -1778 0 feedthrough
rlabel pdiffusion 213 -1778 213 -1778 0 feedthrough
rlabel pdiffusion 220 -1778 220 -1778 0 feedthrough
rlabel pdiffusion 227 -1778 227 -1778 0 feedthrough
rlabel pdiffusion 234 -1778 234 -1778 0 feedthrough
rlabel pdiffusion 241 -1778 241 -1778 0 feedthrough
rlabel pdiffusion 248 -1778 248 -1778 0 feedthrough
rlabel pdiffusion 255 -1778 255 -1778 0 feedthrough
rlabel pdiffusion 262 -1778 262 -1778 0 feedthrough
rlabel pdiffusion 269 -1778 269 -1778 0 feedthrough
rlabel pdiffusion 276 -1778 276 -1778 0 feedthrough
rlabel pdiffusion 283 -1778 283 -1778 0 feedthrough
rlabel pdiffusion 290 -1778 290 -1778 0 feedthrough
rlabel pdiffusion 297 -1778 297 -1778 0 feedthrough
rlabel pdiffusion 304 -1778 304 -1778 0 feedthrough
rlabel pdiffusion 311 -1778 311 -1778 0 feedthrough
rlabel pdiffusion 318 -1778 318 -1778 0 feedthrough
rlabel pdiffusion 325 -1778 325 -1778 0 feedthrough
rlabel pdiffusion 332 -1778 332 -1778 0 feedthrough
rlabel pdiffusion 339 -1778 339 -1778 0 feedthrough
rlabel pdiffusion 346 -1778 346 -1778 0 feedthrough
rlabel pdiffusion 353 -1778 353 -1778 0 feedthrough
rlabel pdiffusion 360 -1778 360 -1778 0 feedthrough
rlabel pdiffusion 367 -1778 367 -1778 0 feedthrough
rlabel pdiffusion 374 -1778 374 -1778 0 feedthrough
rlabel pdiffusion 381 -1778 381 -1778 0 feedthrough
rlabel pdiffusion 388 -1778 388 -1778 0 feedthrough
rlabel pdiffusion 395 -1778 395 -1778 0 cellNo=482
rlabel pdiffusion 402 -1778 402 -1778 0 feedthrough
rlabel pdiffusion 409 -1778 409 -1778 0 feedthrough
rlabel pdiffusion 416 -1778 416 -1778 0 cellNo=132
rlabel pdiffusion 423 -1778 423 -1778 0 feedthrough
rlabel pdiffusion 430 -1778 430 -1778 0 feedthrough
rlabel pdiffusion 437 -1778 437 -1778 0 feedthrough
rlabel pdiffusion 444 -1778 444 -1778 0 feedthrough
rlabel pdiffusion 451 -1778 451 -1778 0 feedthrough
rlabel pdiffusion 458 -1778 458 -1778 0 feedthrough
rlabel pdiffusion 465 -1778 465 -1778 0 feedthrough
rlabel pdiffusion 472 -1778 472 -1778 0 feedthrough
rlabel pdiffusion 479 -1778 479 -1778 0 cellNo=605
rlabel pdiffusion 486 -1778 486 -1778 0 feedthrough
rlabel pdiffusion 493 -1778 493 -1778 0 feedthrough
rlabel pdiffusion 500 -1778 500 -1778 0 feedthrough
rlabel pdiffusion 507 -1778 507 -1778 0 feedthrough
rlabel pdiffusion 514 -1778 514 -1778 0 cellNo=426
rlabel pdiffusion 521 -1778 521 -1778 0 cellNo=95
rlabel pdiffusion 528 -1778 528 -1778 0 feedthrough
rlabel pdiffusion 535 -1778 535 -1778 0 feedthrough
rlabel pdiffusion 542 -1778 542 -1778 0 feedthrough
rlabel pdiffusion 549 -1778 549 -1778 0 feedthrough
rlabel pdiffusion 556 -1778 556 -1778 0 cellNo=646
rlabel pdiffusion 563 -1778 563 -1778 0 cellNo=941
rlabel pdiffusion 570 -1778 570 -1778 0 feedthrough
rlabel pdiffusion 577 -1778 577 -1778 0 feedthrough
rlabel pdiffusion 584 -1778 584 -1778 0 feedthrough
rlabel pdiffusion 591 -1778 591 -1778 0 feedthrough
rlabel pdiffusion 598 -1778 598 -1778 0 cellNo=323
rlabel pdiffusion 605 -1778 605 -1778 0 feedthrough
rlabel pdiffusion 612 -1778 612 -1778 0 feedthrough
rlabel pdiffusion 619 -1778 619 -1778 0 feedthrough
rlabel pdiffusion 626 -1778 626 -1778 0 feedthrough
rlabel pdiffusion 633 -1778 633 -1778 0 feedthrough
rlabel pdiffusion 640 -1778 640 -1778 0 feedthrough
rlabel pdiffusion 647 -1778 647 -1778 0 cellNo=546
rlabel pdiffusion 654 -1778 654 -1778 0 feedthrough
rlabel pdiffusion 661 -1778 661 -1778 0 feedthrough
rlabel pdiffusion 668 -1778 668 -1778 0 feedthrough
rlabel pdiffusion 675 -1778 675 -1778 0 feedthrough
rlabel pdiffusion 682 -1778 682 -1778 0 cellNo=654
rlabel pdiffusion 689 -1778 689 -1778 0 feedthrough
rlabel pdiffusion 696 -1778 696 -1778 0 cellNo=649
rlabel pdiffusion 703 -1778 703 -1778 0 feedthrough
rlabel pdiffusion 710 -1778 710 -1778 0 feedthrough
rlabel pdiffusion 717 -1778 717 -1778 0 feedthrough
rlabel pdiffusion 724 -1778 724 -1778 0 feedthrough
rlabel pdiffusion 731 -1778 731 -1778 0 feedthrough
rlabel pdiffusion 738 -1778 738 -1778 0 cellNo=647
rlabel pdiffusion 745 -1778 745 -1778 0 feedthrough
rlabel pdiffusion 752 -1778 752 -1778 0 feedthrough
rlabel pdiffusion 759 -1778 759 -1778 0 feedthrough
rlabel pdiffusion 766 -1778 766 -1778 0 feedthrough
rlabel pdiffusion 773 -1778 773 -1778 0 feedthrough
rlabel pdiffusion 780 -1778 780 -1778 0 feedthrough
rlabel pdiffusion 787 -1778 787 -1778 0 feedthrough
rlabel pdiffusion 794 -1778 794 -1778 0 feedthrough
rlabel pdiffusion 801 -1778 801 -1778 0 feedthrough
rlabel pdiffusion 808 -1778 808 -1778 0 cellNo=336
rlabel pdiffusion 815 -1778 815 -1778 0 feedthrough
rlabel pdiffusion 822 -1778 822 -1778 0 feedthrough
rlabel pdiffusion 829 -1778 829 -1778 0 cellNo=432
rlabel pdiffusion 836 -1778 836 -1778 0 feedthrough
rlabel pdiffusion 843 -1778 843 -1778 0 feedthrough
rlabel pdiffusion 850 -1778 850 -1778 0 feedthrough
rlabel pdiffusion 857 -1778 857 -1778 0 feedthrough
rlabel pdiffusion 864 -1778 864 -1778 0 feedthrough
rlabel pdiffusion 871 -1778 871 -1778 0 feedthrough
rlabel pdiffusion 878 -1778 878 -1778 0 feedthrough
rlabel pdiffusion 885 -1778 885 -1778 0 cellNo=376
rlabel pdiffusion 892 -1778 892 -1778 0 feedthrough
rlabel pdiffusion 899 -1778 899 -1778 0 cellNo=311
rlabel pdiffusion 906 -1778 906 -1778 0 feedthrough
rlabel pdiffusion 913 -1778 913 -1778 0 feedthrough
rlabel pdiffusion 920 -1778 920 -1778 0 feedthrough
rlabel pdiffusion 927 -1778 927 -1778 0 feedthrough
rlabel pdiffusion 934 -1778 934 -1778 0 feedthrough
rlabel pdiffusion 941 -1778 941 -1778 0 cellNo=744
rlabel pdiffusion 948 -1778 948 -1778 0 feedthrough
rlabel pdiffusion 955 -1778 955 -1778 0 feedthrough
rlabel pdiffusion 962 -1778 962 -1778 0 feedthrough
rlabel pdiffusion 969 -1778 969 -1778 0 feedthrough
rlabel pdiffusion 976 -1778 976 -1778 0 feedthrough
rlabel pdiffusion 983 -1778 983 -1778 0 cellNo=919
rlabel pdiffusion 990 -1778 990 -1778 0 feedthrough
rlabel pdiffusion 997 -1778 997 -1778 0 feedthrough
rlabel pdiffusion 1004 -1778 1004 -1778 0 feedthrough
rlabel pdiffusion 1011 -1778 1011 -1778 0 feedthrough
rlabel pdiffusion 1018 -1778 1018 -1778 0 feedthrough
rlabel pdiffusion 1025 -1778 1025 -1778 0 feedthrough
rlabel pdiffusion 1032 -1778 1032 -1778 0 feedthrough
rlabel pdiffusion 1039 -1778 1039 -1778 0 feedthrough
rlabel pdiffusion 1046 -1778 1046 -1778 0 feedthrough
rlabel pdiffusion 1053 -1778 1053 -1778 0 feedthrough
rlabel pdiffusion 1060 -1778 1060 -1778 0 feedthrough
rlabel pdiffusion 1067 -1778 1067 -1778 0 feedthrough
rlabel pdiffusion 1074 -1778 1074 -1778 0 cellNo=697
rlabel pdiffusion 1081 -1778 1081 -1778 0 cellNo=298
rlabel pdiffusion 1088 -1778 1088 -1778 0 feedthrough
rlabel pdiffusion 1095 -1778 1095 -1778 0 feedthrough
rlabel pdiffusion 1102 -1778 1102 -1778 0 cellNo=393
rlabel pdiffusion 1109 -1778 1109 -1778 0 cellNo=14
rlabel pdiffusion 1116 -1778 1116 -1778 0 feedthrough
rlabel pdiffusion 1123 -1778 1123 -1778 0 feedthrough
rlabel pdiffusion 1130 -1778 1130 -1778 0 feedthrough
rlabel pdiffusion 1137 -1778 1137 -1778 0 feedthrough
rlabel pdiffusion 1144 -1778 1144 -1778 0 feedthrough
rlabel pdiffusion 1151 -1778 1151 -1778 0 feedthrough
rlabel pdiffusion 1158 -1778 1158 -1778 0 feedthrough
rlabel pdiffusion 1165 -1778 1165 -1778 0 feedthrough
rlabel pdiffusion 1172 -1778 1172 -1778 0 feedthrough
rlabel pdiffusion 1179 -1778 1179 -1778 0 feedthrough
rlabel pdiffusion 1186 -1778 1186 -1778 0 feedthrough
rlabel pdiffusion 1193 -1778 1193 -1778 0 feedthrough
rlabel pdiffusion 1200 -1778 1200 -1778 0 feedthrough
rlabel pdiffusion 1207 -1778 1207 -1778 0 feedthrough
rlabel pdiffusion 1214 -1778 1214 -1778 0 feedthrough
rlabel pdiffusion 1221 -1778 1221 -1778 0 feedthrough
rlabel pdiffusion 1228 -1778 1228 -1778 0 feedthrough
rlabel pdiffusion 1235 -1778 1235 -1778 0 feedthrough
rlabel pdiffusion 1242 -1778 1242 -1778 0 cellNo=72
rlabel pdiffusion 1249 -1778 1249 -1778 0 feedthrough
rlabel pdiffusion 1256 -1778 1256 -1778 0 feedthrough
rlabel pdiffusion 1263 -1778 1263 -1778 0 feedthrough
rlabel pdiffusion 1270 -1778 1270 -1778 0 feedthrough
rlabel pdiffusion 1277 -1778 1277 -1778 0 feedthrough
rlabel pdiffusion 1284 -1778 1284 -1778 0 feedthrough
rlabel pdiffusion 1291 -1778 1291 -1778 0 feedthrough
rlabel pdiffusion 1298 -1778 1298 -1778 0 feedthrough
rlabel pdiffusion 1305 -1778 1305 -1778 0 cellNo=354
rlabel pdiffusion 1312 -1778 1312 -1778 0 feedthrough
rlabel pdiffusion 1319 -1778 1319 -1778 0 cellNo=242
rlabel pdiffusion 1326 -1778 1326 -1778 0 feedthrough
rlabel pdiffusion 1333 -1778 1333 -1778 0 feedthrough
rlabel pdiffusion 1340 -1778 1340 -1778 0 feedthrough
rlabel pdiffusion 1347 -1778 1347 -1778 0 feedthrough
rlabel pdiffusion 1354 -1778 1354 -1778 0 cellNo=502
rlabel pdiffusion 1361 -1778 1361 -1778 0 cellNo=758
rlabel pdiffusion 1368 -1778 1368 -1778 0 feedthrough
rlabel pdiffusion 1375 -1778 1375 -1778 0 feedthrough
rlabel pdiffusion 1382 -1778 1382 -1778 0 feedthrough
rlabel pdiffusion 1389 -1778 1389 -1778 0 feedthrough
rlabel pdiffusion 1396 -1778 1396 -1778 0 feedthrough
rlabel pdiffusion 1403 -1778 1403 -1778 0 feedthrough
rlabel pdiffusion 1410 -1778 1410 -1778 0 feedthrough
rlabel pdiffusion 1417 -1778 1417 -1778 0 feedthrough
rlabel pdiffusion 1424 -1778 1424 -1778 0 feedthrough
rlabel pdiffusion 1431 -1778 1431 -1778 0 feedthrough
rlabel pdiffusion 1438 -1778 1438 -1778 0 feedthrough
rlabel pdiffusion 1445 -1778 1445 -1778 0 feedthrough
rlabel pdiffusion 1452 -1778 1452 -1778 0 feedthrough
rlabel pdiffusion 1459 -1778 1459 -1778 0 feedthrough
rlabel pdiffusion 1466 -1778 1466 -1778 0 cellNo=46
rlabel pdiffusion 1473 -1778 1473 -1778 0 feedthrough
rlabel pdiffusion 1480 -1778 1480 -1778 0 feedthrough
rlabel pdiffusion 1487 -1778 1487 -1778 0 feedthrough
rlabel pdiffusion 1494 -1778 1494 -1778 0 feedthrough
rlabel pdiffusion 1501 -1778 1501 -1778 0 feedthrough
rlabel pdiffusion 1508 -1778 1508 -1778 0 feedthrough
rlabel pdiffusion 1515 -1778 1515 -1778 0 feedthrough
rlabel pdiffusion 1522 -1778 1522 -1778 0 feedthrough
rlabel pdiffusion 1529 -1778 1529 -1778 0 feedthrough
rlabel pdiffusion 1536 -1778 1536 -1778 0 feedthrough
rlabel pdiffusion 1543 -1778 1543 -1778 0 feedthrough
rlabel pdiffusion 1550 -1778 1550 -1778 0 feedthrough
rlabel pdiffusion 1557 -1778 1557 -1778 0 feedthrough
rlabel pdiffusion 1564 -1778 1564 -1778 0 feedthrough
rlabel pdiffusion 1571 -1778 1571 -1778 0 feedthrough
rlabel pdiffusion 1578 -1778 1578 -1778 0 feedthrough
rlabel pdiffusion 1585 -1778 1585 -1778 0 feedthrough
rlabel pdiffusion 1592 -1778 1592 -1778 0 feedthrough
rlabel pdiffusion 1599 -1778 1599 -1778 0 feedthrough
rlabel pdiffusion 1606 -1778 1606 -1778 0 feedthrough
rlabel pdiffusion 1613 -1778 1613 -1778 0 feedthrough
rlabel pdiffusion 1620 -1778 1620 -1778 0 feedthrough
rlabel pdiffusion 1627 -1778 1627 -1778 0 feedthrough
rlabel pdiffusion 1634 -1778 1634 -1778 0 feedthrough
rlabel pdiffusion 1641 -1778 1641 -1778 0 feedthrough
rlabel pdiffusion 1648 -1778 1648 -1778 0 feedthrough
rlabel pdiffusion 1655 -1778 1655 -1778 0 feedthrough
rlabel pdiffusion 1662 -1778 1662 -1778 0 feedthrough
rlabel pdiffusion 1669 -1778 1669 -1778 0 feedthrough
rlabel pdiffusion 1676 -1778 1676 -1778 0 feedthrough
rlabel pdiffusion 1683 -1778 1683 -1778 0 feedthrough
rlabel pdiffusion 1690 -1778 1690 -1778 0 feedthrough
rlabel pdiffusion 1697 -1778 1697 -1778 0 feedthrough
rlabel pdiffusion 1704 -1778 1704 -1778 0 feedthrough
rlabel pdiffusion 1711 -1778 1711 -1778 0 feedthrough
rlabel pdiffusion 1718 -1778 1718 -1778 0 feedthrough
rlabel pdiffusion 1725 -1778 1725 -1778 0 feedthrough
rlabel pdiffusion 1732 -1778 1732 -1778 0 feedthrough
rlabel pdiffusion 1739 -1778 1739 -1778 0 feedthrough
rlabel pdiffusion 1746 -1778 1746 -1778 0 feedthrough
rlabel pdiffusion 1753 -1778 1753 -1778 0 feedthrough
rlabel pdiffusion 1760 -1778 1760 -1778 0 feedthrough
rlabel pdiffusion 1767 -1778 1767 -1778 0 feedthrough
rlabel pdiffusion 1774 -1778 1774 -1778 0 feedthrough
rlabel pdiffusion 1781 -1778 1781 -1778 0 feedthrough
rlabel pdiffusion 1788 -1778 1788 -1778 0 feedthrough
rlabel pdiffusion 1795 -1778 1795 -1778 0 feedthrough
rlabel pdiffusion 1802 -1778 1802 -1778 0 feedthrough
rlabel pdiffusion 1809 -1778 1809 -1778 0 feedthrough
rlabel pdiffusion 1816 -1778 1816 -1778 0 feedthrough
rlabel pdiffusion 1823 -1778 1823 -1778 0 feedthrough
rlabel pdiffusion 1830 -1778 1830 -1778 0 feedthrough
rlabel pdiffusion 1837 -1778 1837 -1778 0 feedthrough
rlabel pdiffusion 1844 -1778 1844 -1778 0 feedthrough
rlabel pdiffusion 1851 -1778 1851 -1778 0 feedthrough
rlabel pdiffusion 1858 -1778 1858 -1778 0 feedthrough
rlabel pdiffusion 1865 -1778 1865 -1778 0 feedthrough
rlabel pdiffusion 1872 -1778 1872 -1778 0 feedthrough
rlabel pdiffusion 1879 -1778 1879 -1778 0 feedthrough
rlabel pdiffusion 1886 -1778 1886 -1778 0 feedthrough
rlabel pdiffusion 1893 -1778 1893 -1778 0 feedthrough
rlabel pdiffusion 1900 -1778 1900 -1778 0 feedthrough
rlabel pdiffusion 1907 -1778 1907 -1778 0 feedthrough
rlabel pdiffusion 1914 -1778 1914 -1778 0 feedthrough
rlabel pdiffusion 1921 -1778 1921 -1778 0 feedthrough
rlabel pdiffusion 1928 -1778 1928 -1778 0 feedthrough
rlabel pdiffusion 1935 -1778 1935 -1778 0 cellNo=436
rlabel pdiffusion 1942 -1778 1942 -1778 0 cellNo=437
rlabel pdiffusion 1949 -1778 1949 -1778 0 feedthrough
rlabel pdiffusion 1956 -1778 1956 -1778 0 feedthrough
rlabel pdiffusion 1963 -1778 1963 -1778 0 feedthrough
rlabel pdiffusion 1970 -1778 1970 -1778 0 feedthrough
rlabel pdiffusion 2019 -1778 2019 -1778 0 feedthrough
rlabel pdiffusion 3 -1903 3 -1903 0 cellNo=920
rlabel pdiffusion 10 -1903 10 -1903 0 cellNo=1116
rlabel pdiffusion 17 -1903 17 -1903 0 feedthrough
rlabel pdiffusion 24 -1903 24 -1903 0 feedthrough
rlabel pdiffusion 31 -1903 31 -1903 0 feedthrough
rlabel pdiffusion 38 -1903 38 -1903 0 feedthrough
rlabel pdiffusion 45 -1903 45 -1903 0 feedthrough
rlabel pdiffusion 52 -1903 52 -1903 0 feedthrough
rlabel pdiffusion 59 -1903 59 -1903 0 cellNo=633
rlabel pdiffusion 66 -1903 66 -1903 0 feedthrough
rlabel pdiffusion 73 -1903 73 -1903 0 feedthrough
rlabel pdiffusion 80 -1903 80 -1903 0 feedthrough
rlabel pdiffusion 87 -1903 87 -1903 0 feedthrough
rlabel pdiffusion 94 -1903 94 -1903 0 feedthrough
rlabel pdiffusion 101 -1903 101 -1903 0 cellNo=574
rlabel pdiffusion 108 -1903 108 -1903 0 feedthrough
rlabel pdiffusion 115 -1903 115 -1903 0 feedthrough
rlabel pdiffusion 122 -1903 122 -1903 0 feedthrough
rlabel pdiffusion 129 -1903 129 -1903 0 feedthrough
rlabel pdiffusion 136 -1903 136 -1903 0 cellNo=740
rlabel pdiffusion 143 -1903 143 -1903 0 cellNo=398
rlabel pdiffusion 150 -1903 150 -1903 0 feedthrough
rlabel pdiffusion 157 -1903 157 -1903 0 feedthrough
rlabel pdiffusion 164 -1903 164 -1903 0 feedthrough
rlabel pdiffusion 171 -1903 171 -1903 0 feedthrough
rlabel pdiffusion 178 -1903 178 -1903 0 feedthrough
rlabel pdiffusion 185 -1903 185 -1903 0 feedthrough
rlabel pdiffusion 192 -1903 192 -1903 0 feedthrough
rlabel pdiffusion 199 -1903 199 -1903 0 cellNo=193
rlabel pdiffusion 206 -1903 206 -1903 0 feedthrough
rlabel pdiffusion 213 -1903 213 -1903 0 feedthrough
rlabel pdiffusion 220 -1903 220 -1903 0 feedthrough
rlabel pdiffusion 227 -1903 227 -1903 0 feedthrough
rlabel pdiffusion 234 -1903 234 -1903 0 feedthrough
rlabel pdiffusion 241 -1903 241 -1903 0 feedthrough
rlabel pdiffusion 248 -1903 248 -1903 0 feedthrough
rlabel pdiffusion 255 -1903 255 -1903 0 feedthrough
rlabel pdiffusion 262 -1903 262 -1903 0 feedthrough
rlabel pdiffusion 269 -1903 269 -1903 0 feedthrough
rlabel pdiffusion 276 -1903 276 -1903 0 feedthrough
rlabel pdiffusion 283 -1903 283 -1903 0 feedthrough
rlabel pdiffusion 290 -1903 290 -1903 0 feedthrough
rlabel pdiffusion 297 -1903 297 -1903 0 feedthrough
rlabel pdiffusion 304 -1903 304 -1903 0 feedthrough
rlabel pdiffusion 311 -1903 311 -1903 0 feedthrough
rlabel pdiffusion 318 -1903 318 -1903 0 feedthrough
rlabel pdiffusion 325 -1903 325 -1903 0 feedthrough
rlabel pdiffusion 332 -1903 332 -1903 0 feedthrough
rlabel pdiffusion 339 -1903 339 -1903 0 feedthrough
rlabel pdiffusion 346 -1903 346 -1903 0 feedthrough
rlabel pdiffusion 353 -1903 353 -1903 0 feedthrough
rlabel pdiffusion 360 -1903 360 -1903 0 feedthrough
rlabel pdiffusion 367 -1903 367 -1903 0 feedthrough
rlabel pdiffusion 374 -1903 374 -1903 0 feedthrough
rlabel pdiffusion 381 -1903 381 -1903 0 feedthrough
rlabel pdiffusion 388 -1903 388 -1903 0 feedthrough
rlabel pdiffusion 395 -1903 395 -1903 0 feedthrough
rlabel pdiffusion 402 -1903 402 -1903 0 cellNo=301
rlabel pdiffusion 409 -1903 409 -1903 0 feedthrough
rlabel pdiffusion 416 -1903 416 -1903 0 feedthrough
rlabel pdiffusion 423 -1903 423 -1903 0 feedthrough
rlabel pdiffusion 430 -1903 430 -1903 0 feedthrough
rlabel pdiffusion 437 -1903 437 -1903 0 feedthrough
rlabel pdiffusion 444 -1903 444 -1903 0 feedthrough
rlabel pdiffusion 451 -1903 451 -1903 0 feedthrough
rlabel pdiffusion 458 -1903 458 -1903 0 feedthrough
rlabel pdiffusion 465 -1903 465 -1903 0 feedthrough
rlabel pdiffusion 472 -1903 472 -1903 0 feedthrough
rlabel pdiffusion 479 -1903 479 -1903 0 cellNo=155
rlabel pdiffusion 486 -1903 486 -1903 0 cellNo=338
rlabel pdiffusion 493 -1903 493 -1903 0 feedthrough
rlabel pdiffusion 500 -1903 500 -1903 0 feedthrough
rlabel pdiffusion 507 -1903 507 -1903 0 cellNo=579
rlabel pdiffusion 514 -1903 514 -1903 0 feedthrough
rlabel pdiffusion 521 -1903 521 -1903 0 feedthrough
rlabel pdiffusion 528 -1903 528 -1903 0 feedthrough
rlabel pdiffusion 535 -1903 535 -1903 0 feedthrough
rlabel pdiffusion 542 -1903 542 -1903 0 feedthrough
rlabel pdiffusion 549 -1903 549 -1903 0 feedthrough
rlabel pdiffusion 556 -1903 556 -1903 0 feedthrough
rlabel pdiffusion 563 -1903 563 -1903 0 feedthrough
rlabel pdiffusion 570 -1903 570 -1903 0 feedthrough
rlabel pdiffusion 577 -1903 577 -1903 0 cellNo=674
rlabel pdiffusion 584 -1903 584 -1903 0 feedthrough
rlabel pdiffusion 591 -1903 591 -1903 0 feedthrough
rlabel pdiffusion 598 -1903 598 -1903 0 feedthrough
rlabel pdiffusion 605 -1903 605 -1903 0 feedthrough
rlabel pdiffusion 612 -1903 612 -1903 0 cellNo=444
rlabel pdiffusion 619 -1903 619 -1903 0 cellNo=978
rlabel pdiffusion 626 -1903 626 -1903 0 feedthrough
rlabel pdiffusion 633 -1903 633 -1903 0 feedthrough
rlabel pdiffusion 640 -1903 640 -1903 0 feedthrough
rlabel pdiffusion 647 -1903 647 -1903 0 feedthrough
rlabel pdiffusion 654 -1903 654 -1903 0 feedthrough
rlabel pdiffusion 661 -1903 661 -1903 0 feedthrough
rlabel pdiffusion 668 -1903 668 -1903 0 feedthrough
rlabel pdiffusion 675 -1903 675 -1903 0 feedthrough
rlabel pdiffusion 682 -1903 682 -1903 0 feedthrough
rlabel pdiffusion 689 -1903 689 -1903 0 cellNo=147
rlabel pdiffusion 696 -1903 696 -1903 0 feedthrough
rlabel pdiffusion 703 -1903 703 -1903 0 feedthrough
rlabel pdiffusion 710 -1903 710 -1903 0 feedthrough
rlabel pdiffusion 717 -1903 717 -1903 0 cellNo=927
rlabel pdiffusion 724 -1903 724 -1903 0 cellNo=881
rlabel pdiffusion 731 -1903 731 -1903 0 feedthrough
rlabel pdiffusion 738 -1903 738 -1903 0 feedthrough
rlabel pdiffusion 745 -1903 745 -1903 0 feedthrough
rlabel pdiffusion 752 -1903 752 -1903 0 feedthrough
rlabel pdiffusion 759 -1903 759 -1903 0 feedthrough
rlabel pdiffusion 766 -1903 766 -1903 0 cellNo=423
rlabel pdiffusion 773 -1903 773 -1903 0 cellNo=857
rlabel pdiffusion 780 -1903 780 -1903 0 feedthrough
rlabel pdiffusion 787 -1903 787 -1903 0 feedthrough
rlabel pdiffusion 794 -1903 794 -1903 0 feedthrough
rlabel pdiffusion 801 -1903 801 -1903 0 feedthrough
rlabel pdiffusion 808 -1903 808 -1903 0 feedthrough
rlabel pdiffusion 815 -1903 815 -1903 0 feedthrough
rlabel pdiffusion 822 -1903 822 -1903 0 feedthrough
rlabel pdiffusion 829 -1903 829 -1903 0 feedthrough
rlabel pdiffusion 836 -1903 836 -1903 0 feedthrough
rlabel pdiffusion 843 -1903 843 -1903 0 feedthrough
rlabel pdiffusion 850 -1903 850 -1903 0 feedthrough
rlabel pdiffusion 857 -1903 857 -1903 0 feedthrough
rlabel pdiffusion 864 -1903 864 -1903 0 feedthrough
rlabel pdiffusion 871 -1903 871 -1903 0 feedthrough
rlabel pdiffusion 878 -1903 878 -1903 0 feedthrough
rlabel pdiffusion 885 -1903 885 -1903 0 cellNo=913
rlabel pdiffusion 892 -1903 892 -1903 0 feedthrough
rlabel pdiffusion 899 -1903 899 -1903 0 feedthrough
rlabel pdiffusion 906 -1903 906 -1903 0 cellNo=553
rlabel pdiffusion 913 -1903 913 -1903 0 feedthrough
rlabel pdiffusion 920 -1903 920 -1903 0 feedthrough
rlabel pdiffusion 927 -1903 927 -1903 0 feedthrough
rlabel pdiffusion 934 -1903 934 -1903 0 cellNo=968
rlabel pdiffusion 941 -1903 941 -1903 0 feedthrough
rlabel pdiffusion 948 -1903 948 -1903 0 feedthrough
rlabel pdiffusion 955 -1903 955 -1903 0 feedthrough
rlabel pdiffusion 962 -1903 962 -1903 0 feedthrough
rlabel pdiffusion 969 -1903 969 -1903 0 feedthrough
rlabel pdiffusion 976 -1903 976 -1903 0 feedthrough
rlabel pdiffusion 983 -1903 983 -1903 0 cellNo=126
rlabel pdiffusion 990 -1903 990 -1903 0 feedthrough
rlabel pdiffusion 997 -1903 997 -1903 0 feedthrough
rlabel pdiffusion 1004 -1903 1004 -1903 0 feedthrough
rlabel pdiffusion 1011 -1903 1011 -1903 0 feedthrough
rlabel pdiffusion 1018 -1903 1018 -1903 0 feedthrough
rlabel pdiffusion 1025 -1903 1025 -1903 0 cellNo=738
rlabel pdiffusion 1032 -1903 1032 -1903 0 feedthrough
rlabel pdiffusion 1039 -1903 1039 -1903 0 feedthrough
rlabel pdiffusion 1046 -1903 1046 -1903 0 feedthrough
rlabel pdiffusion 1053 -1903 1053 -1903 0 feedthrough
rlabel pdiffusion 1060 -1903 1060 -1903 0 cellNo=518
rlabel pdiffusion 1067 -1903 1067 -1903 0 feedthrough
rlabel pdiffusion 1074 -1903 1074 -1903 0 feedthrough
rlabel pdiffusion 1081 -1903 1081 -1903 0 feedthrough
rlabel pdiffusion 1088 -1903 1088 -1903 0 cellNo=861
rlabel pdiffusion 1095 -1903 1095 -1903 0 feedthrough
rlabel pdiffusion 1102 -1903 1102 -1903 0 cellNo=716
rlabel pdiffusion 1109 -1903 1109 -1903 0 cellNo=963
rlabel pdiffusion 1116 -1903 1116 -1903 0 feedthrough
rlabel pdiffusion 1123 -1903 1123 -1903 0 cellNo=230
rlabel pdiffusion 1130 -1903 1130 -1903 0 feedthrough
rlabel pdiffusion 1137 -1903 1137 -1903 0 feedthrough
rlabel pdiffusion 1144 -1903 1144 -1903 0 feedthrough
rlabel pdiffusion 1151 -1903 1151 -1903 0 cellNo=278
rlabel pdiffusion 1158 -1903 1158 -1903 0 feedthrough
rlabel pdiffusion 1165 -1903 1165 -1903 0 feedthrough
rlabel pdiffusion 1172 -1903 1172 -1903 0 feedthrough
rlabel pdiffusion 1179 -1903 1179 -1903 0 feedthrough
rlabel pdiffusion 1186 -1903 1186 -1903 0 feedthrough
rlabel pdiffusion 1193 -1903 1193 -1903 0 feedthrough
rlabel pdiffusion 1200 -1903 1200 -1903 0 feedthrough
rlabel pdiffusion 1207 -1903 1207 -1903 0 cellNo=802
rlabel pdiffusion 1214 -1903 1214 -1903 0 feedthrough
rlabel pdiffusion 1221 -1903 1221 -1903 0 cellNo=229
rlabel pdiffusion 1228 -1903 1228 -1903 0 feedthrough
rlabel pdiffusion 1235 -1903 1235 -1903 0 feedthrough
rlabel pdiffusion 1242 -1903 1242 -1903 0 feedthrough
rlabel pdiffusion 1249 -1903 1249 -1903 0 feedthrough
rlabel pdiffusion 1256 -1903 1256 -1903 0 feedthrough
rlabel pdiffusion 1263 -1903 1263 -1903 0 feedthrough
rlabel pdiffusion 1270 -1903 1270 -1903 0 feedthrough
rlabel pdiffusion 1277 -1903 1277 -1903 0 cellNo=822
rlabel pdiffusion 1284 -1903 1284 -1903 0 feedthrough
rlabel pdiffusion 1291 -1903 1291 -1903 0 feedthrough
rlabel pdiffusion 1298 -1903 1298 -1903 0 feedthrough
rlabel pdiffusion 1305 -1903 1305 -1903 0 feedthrough
rlabel pdiffusion 1312 -1903 1312 -1903 0 feedthrough
rlabel pdiffusion 1319 -1903 1319 -1903 0 feedthrough
rlabel pdiffusion 1326 -1903 1326 -1903 0 feedthrough
rlabel pdiffusion 1333 -1903 1333 -1903 0 feedthrough
rlabel pdiffusion 1340 -1903 1340 -1903 0 feedthrough
rlabel pdiffusion 1347 -1903 1347 -1903 0 feedthrough
rlabel pdiffusion 1354 -1903 1354 -1903 0 feedthrough
rlabel pdiffusion 1361 -1903 1361 -1903 0 feedthrough
rlabel pdiffusion 1368 -1903 1368 -1903 0 feedthrough
rlabel pdiffusion 1375 -1903 1375 -1903 0 feedthrough
rlabel pdiffusion 1382 -1903 1382 -1903 0 feedthrough
rlabel pdiffusion 1389 -1903 1389 -1903 0 feedthrough
rlabel pdiffusion 1396 -1903 1396 -1903 0 feedthrough
rlabel pdiffusion 1403 -1903 1403 -1903 0 feedthrough
rlabel pdiffusion 1410 -1903 1410 -1903 0 feedthrough
rlabel pdiffusion 1417 -1903 1417 -1903 0 feedthrough
rlabel pdiffusion 1424 -1903 1424 -1903 0 feedthrough
rlabel pdiffusion 1431 -1903 1431 -1903 0 feedthrough
rlabel pdiffusion 1438 -1903 1438 -1903 0 feedthrough
rlabel pdiffusion 1445 -1903 1445 -1903 0 feedthrough
rlabel pdiffusion 1452 -1903 1452 -1903 0 feedthrough
rlabel pdiffusion 1459 -1903 1459 -1903 0 feedthrough
rlabel pdiffusion 1466 -1903 1466 -1903 0 feedthrough
rlabel pdiffusion 1473 -1903 1473 -1903 0 feedthrough
rlabel pdiffusion 1480 -1903 1480 -1903 0 feedthrough
rlabel pdiffusion 1487 -1903 1487 -1903 0 feedthrough
rlabel pdiffusion 1494 -1903 1494 -1903 0 feedthrough
rlabel pdiffusion 1501 -1903 1501 -1903 0 feedthrough
rlabel pdiffusion 1508 -1903 1508 -1903 0 feedthrough
rlabel pdiffusion 1515 -1903 1515 -1903 0 feedthrough
rlabel pdiffusion 1522 -1903 1522 -1903 0 feedthrough
rlabel pdiffusion 1529 -1903 1529 -1903 0 feedthrough
rlabel pdiffusion 1536 -1903 1536 -1903 0 feedthrough
rlabel pdiffusion 1543 -1903 1543 -1903 0 feedthrough
rlabel pdiffusion 1550 -1903 1550 -1903 0 feedthrough
rlabel pdiffusion 1557 -1903 1557 -1903 0 feedthrough
rlabel pdiffusion 1564 -1903 1564 -1903 0 cellNo=979
rlabel pdiffusion 1571 -1903 1571 -1903 0 feedthrough
rlabel pdiffusion 1578 -1903 1578 -1903 0 feedthrough
rlabel pdiffusion 1585 -1903 1585 -1903 0 feedthrough
rlabel pdiffusion 1592 -1903 1592 -1903 0 feedthrough
rlabel pdiffusion 1599 -1903 1599 -1903 0 feedthrough
rlabel pdiffusion 1606 -1903 1606 -1903 0 feedthrough
rlabel pdiffusion 1613 -1903 1613 -1903 0 feedthrough
rlabel pdiffusion 1620 -1903 1620 -1903 0 feedthrough
rlabel pdiffusion 1627 -1903 1627 -1903 0 feedthrough
rlabel pdiffusion 1634 -1903 1634 -1903 0 feedthrough
rlabel pdiffusion 1641 -1903 1641 -1903 0 feedthrough
rlabel pdiffusion 1648 -1903 1648 -1903 0 feedthrough
rlabel pdiffusion 1655 -1903 1655 -1903 0 feedthrough
rlabel pdiffusion 1662 -1903 1662 -1903 0 feedthrough
rlabel pdiffusion 1669 -1903 1669 -1903 0 feedthrough
rlabel pdiffusion 1676 -1903 1676 -1903 0 feedthrough
rlabel pdiffusion 1683 -1903 1683 -1903 0 feedthrough
rlabel pdiffusion 1690 -1903 1690 -1903 0 feedthrough
rlabel pdiffusion 1697 -1903 1697 -1903 0 feedthrough
rlabel pdiffusion 1704 -1903 1704 -1903 0 feedthrough
rlabel pdiffusion 1711 -1903 1711 -1903 0 feedthrough
rlabel pdiffusion 1718 -1903 1718 -1903 0 feedthrough
rlabel pdiffusion 1725 -1903 1725 -1903 0 feedthrough
rlabel pdiffusion 1732 -1903 1732 -1903 0 feedthrough
rlabel pdiffusion 1739 -1903 1739 -1903 0 feedthrough
rlabel pdiffusion 1746 -1903 1746 -1903 0 feedthrough
rlabel pdiffusion 1753 -1903 1753 -1903 0 feedthrough
rlabel pdiffusion 1760 -1903 1760 -1903 0 feedthrough
rlabel pdiffusion 1767 -1903 1767 -1903 0 feedthrough
rlabel pdiffusion 1774 -1903 1774 -1903 0 feedthrough
rlabel pdiffusion 1781 -1903 1781 -1903 0 feedthrough
rlabel pdiffusion 1788 -1903 1788 -1903 0 feedthrough
rlabel pdiffusion 1795 -1903 1795 -1903 0 feedthrough
rlabel pdiffusion 1802 -1903 1802 -1903 0 feedthrough
rlabel pdiffusion 1809 -1903 1809 -1903 0 feedthrough
rlabel pdiffusion 1816 -1903 1816 -1903 0 feedthrough
rlabel pdiffusion 1823 -1903 1823 -1903 0 feedthrough
rlabel pdiffusion 1830 -1903 1830 -1903 0 feedthrough
rlabel pdiffusion 1837 -1903 1837 -1903 0 feedthrough
rlabel pdiffusion 1844 -1903 1844 -1903 0 feedthrough
rlabel pdiffusion 1851 -1903 1851 -1903 0 feedthrough
rlabel pdiffusion 1858 -1903 1858 -1903 0 feedthrough
rlabel pdiffusion 1865 -1903 1865 -1903 0 feedthrough
rlabel pdiffusion 1872 -1903 1872 -1903 0 feedthrough
rlabel pdiffusion 1879 -1903 1879 -1903 0 feedthrough
rlabel pdiffusion 1886 -1903 1886 -1903 0 feedthrough
rlabel pdiffusion 1893 -1903 1893 -1903 0 feedthrough
rlabel pdiffusion 1900 -1903 1900 -1903 0 feedthrough
rlabel pdiffusion 1907 -1903 1907 -1903 0 feedthrough
rlabel pdiffusion 1914 -1903 1914 -1903 0 feedthrough
rlabel pdiffusion 1921 -1903 1921 -1903 0 feedthrough
rlabel pdiffusion 1928 -1903 1928 -1903 0 feedthrough
rlabel pdiffusion 1935 -1903 1935 -1903 0 feedthrough
rlabel pdiffusion 1942 -1903 1942 -1903 0 feedthrough
rlabel pdiffusion 1949 -1903 1949 -1903 0 feedthrough
rlabel pdiffusion 1956 -1903 1956 -1903 0 feedthrough
rlabel pdiffusion 1963 -1903 1963 -1903 0 feedthrough
rlabel pdiffusion 1970 -1903 1970 -1903 0 feedthrough
rlabel pdiffusion 1977 -1903 1977 -1903 0 feedthrough
rlabel pdiffusion 1984 -1903 1984 -1903 0 feedthrough
rlabel pdiffusion 1991 -1903 1991 -1903 0 feedthrough
rlabel pdiffusion 1998 -1903 1998 -1903 0 feedthrough
rlabel pdiffusion 2005 -1903 2005 -1903 0 feedthrough
rlabel pdiffusion 2012 -1903 2012 -1903 0 cellNo=759
rlabel pdiffusion 2019 -1903 2019 -1903 0 feedthrough
rlabel pdiffusion 2026 -1903 2026 -1903 0 feedthrough
rlabel pdiffusion 3 -2050 3 -2050 0 feedthrough
rlabel pdiffusion 10 -2050 10 -2050 0 feedthrough
rlabel pdiffusion 17 -2050 17 -2050 0 cellNo=388
rlabel pdiffusion 24 -2050 24 -2050 0 feedthrough
rlabel pdiffusion 31 -2050 31 -2050 0 feedthrough
rlabel pdiffusion 38 -2050 38 -2050 0 feedthrough
rlabel pdiffusion 45 -2050 45 -2050 0 feedthrough
rlabel pdiffusion 52 -2050 52 -2050 0 feedthrough
rlabel pdiffusion 59 -2050 59 -2050 0 feedthrough
rlabel pdiffusion 66 -2050 66 -2050 0 cellNo=422
rlabel pdiffusion 73 -2050 73 -2050 0 feedthrough
rlabel pdiffusion 80 -2050 80 -2050 0 feedthrough
rlabel pdiffusion 87 -2050 87 -2050 0 feedthrough
rlabel pdiffusion 94 -2050 94 -2050 0 feedthrough
rlabel pdiffusion 101 -2050 101 -2050 0 feedthrough
rlabel pdiffusion 108 -2050 108 -2050 0 feedthrough
rlabel pdiffusion 115 -2050 115 -2050 0 cellNo=931
rlabel pdiffusion 122 -2050 122 -2050 0 feedthrough
rlabel pdiffusion 129 -2050 129 -2050 0 feedthrough
rlabel pdiffusion 136 -2050 136 -2050 0 feedthrough
rlabel pdiffusion 143 -2050 143 -2050 0 cellNo=166
rlabel pdiffusion 150 -2050 150 -2050 0 feedthrough
rlabel pdiffusion 157 -2050 157 -2050 0 feedthrough
rlabel pdiffusion 164 -2050 164 -2050 0 feedthrough
rlabel pdiffusion 171 -2050 171 -2050 0 feedthrough
rlabel pdiffusion 178 -2050 178 -2050 0 feedthrough
rlabel pdiffusion 185 -2050 185 -2050 0 feedthrough
rlabel pdiffusion 192 -2050 192 -2050 0 feedthrough
rlabel pdiffusion 199 -2050 199 -2050 0 feedthrough
rlabel pdiffusion 206 -2050 206 -2050 0 feedthrough
rlabel pdiffusion 213 -2050 213 -2050 0 feedthrough
rlabel pdiffusion 220 -2050 220 -2050 0 cellNo=385
rlabel pdiffusion 227 -2050 227 -2050 0 feedthrough
rlabel pdiffusion 234 -2050 234 -2050 0 feedthrough
rlabel pdiffusion 241 -2050 241 -2050 0 cellNo=667
rlabel pdiffusion 248 -2050 248 -2050 0 feedthrough
rlabel pdiffusion 255 -2050 255 -2050 0 feedthrough
rlabel pdiffusion 262 -2050 262 -2050 0 feedthrough
rlabel pdiffusion 269 -2050 269 -2050 0 feedthrough
rlabel pdiffusion 276 -2050 276 -2050 0 feedthrough
rlabel pdiffusion 283 -2050 283 -2050 0 feedthrough
rlabel pdiffusion 290 -2050 290 -2050 0 feedthrough
rlabel pdiffusion 297 -2050 297 -2050 0 feedthrough
rlabel pdiffusion 304 -2050 304 -2050 0 feedthrough
rlabel pdiffusion 311 -2050 311 -2050 0 cellNo=100
rlabel pdiffusion 318 -2050 318 -2050 0 feedthrough
rlabel pdiffusion 325 -2050 325 -2050 0 feedthrough
rlabel pdiffusion 332 -2050 332 -2050 0 feedthrough
rlabel pdiffusion 339 -2050 339 -2050 0 cellNo=321
rlabel pdiffusion 346 -2050 346 -2050 0 feedthrough
rlabel pdiffusion 353 -2050 353 -2050 0 feedthrough
rlabel pdiffusion 360 -2050 360 -2050 0 feedthrough
rlabel pdiffusion 367 -2050 367 -2050 0 feedthrough
rlabel pdiffusion 374 -2050 374 -2050 0 feedthrough
rlabel pdiffusion 381 -2050 381 -2050 0 feedthrough
rlabel pdiffusion 388 -2050 388 -2050 0 feedthrough
rlabel pdiffusion 395 -2050 395 -2050 0 feedthrough
rlabel pdiffusion 402 -2050 402 -2050 0 feedthrough
rlabel pdiffusion 409 -2050 409 -2050 0 feedthrough
rlabel pdiffusion 416 -2050 416 -2050 0 feedthrough
rlabel pdiffusion 423 -2050 423 -2050 0 feedthrough
rlabel pdiffusion 430 -2050 430 -2050 0 feedthrough
rlabel pdiffusion 437 -2050 437 -2050 0 feedthrough
rlabel pdiffusion 444 -2050 444 -2050 0 feedthrough
rlabel pdiffusion 451 -2050 451 -2050 0 cellNo=91
rlabel pdiffusion 458 -2050 458 -2050 0 feedthrough
rlabel pdiffusion 465 -2050 465 -2050 0 feedthrough
rlabel pdiffusion 472 -2050 472 -2050 0 feedthrough
rlabel pdiffusion 479 -2050 479 -2050 0 feedthrough
rlabel pdiffusion 486 -2050 486 -2050 0 feedthrough
rlabel pdiffusion 493 -2050 493 -2050 0 feedthrough
rlabel pdiffusion 500 -2050 500 -2050 0 feedthrough
rlabel pdiffusion 507 -2050 507 -2050 0 feedthrough
rlabel pdiffusion 514 -2050 514 -2050 0 feedthrough
rlabel pdiffusion 521 -2050 521 -2050 0 feedthrough
rlabel pdiffusion 528 -2050 528 -2050 0 cellNo=199
rlabel pdiffusion 535 -2050 535 -2050 0 cellNo=10
rlabel pdiffusion 542 -2050 542 -2050 0 feedthrough
rlabel pdiffusion 549 -2050 549 -2050 0 feedthrough
rlabel pdiffusion 556 -2050 556 -2050 0 feedthrough
rlabel pdiffusion 563 -2050 563 -2050 0 feedthrough
rlabel pdiffusion 570 -2050 570 -2050 0 feedthrough
rlabel pdiffusion 577 -2050 577 -2050 0 feedthrough
rlabel pdiffusion 584 -2050 584 -2050 0 feedthrough
rlabel pdiffusion 591 -2050 591 -2050 0 feedthrough
rlabel pdiffusion 598 -2050 598 -2050 0 feedthrough
rlabel pdiffusion 605 -2050 605 -2050 0 feedthrough
rlabel pdiffusion 612 -2050 612 -2050 0 feedthrough
rlabel pdiffusion 619 -2050 619 -2050 0 feedthrough
rlabel pdiffusion 626 -2050 626 -2050 0 feedthrough
rlabel pdiffusion 633 -2050 633 -2050 0 feedthrough
rlabel pdiffusion 640 -2050 640 -2050 0 feedthrough
rlabel pdiffusion 647 -2050 647 -2050 0 feedthrough
rlabel pdiffusion 654 -2050 654 -2050 0 feedthrough
rlabel pdiffusion 661 -2050 661 -2050 0 feedthrough
rlabel pdiffusion 668 -2050 668 -2050 0 feedthrough
rlabel pdiffusion 675 -2050 675 -2050 0 feedthrough
rlabel pdiffusion 682 -2050 682 -2050 0 feedthrough
rlabel pdiffusion 689 -2050 689 -2050 0 feedthrough
rlabel pdiffusion 696 -2050 696 -2050 0 cellNo=971
rlabel pdiffusion 703 -2050 703 -2050 0 feedthrough
rlabel pdiffusion 710 -2050 710 -2050 0 feedthrough
rlabel pdiffusion 717 -2050 717 -2050 0 feedthrough
rlabel pdiffusion 724 -2050 724 -2050 0 cellNo=517
rlabel pdiffusion 731 -2050 731 -2050 0 cellNo=576
rlabel pdiffusion 738 -2050 738 -2050 0 feedthrough
rlabel pdiffusion 745 -2050 745 -2050 0 feedthrough
rlabel pdiffusion 752 -2050 752 -2050 0 cellNo=434
rlabel pdiffusion 759 -2050 759 -2050 0 cellNo=975
rlabel pdiffusion 766 -2050 766 -2050 0 feedthrough
rlabel pdiffusion 773 -2050 773 -2050 0 cellNo=542
rlabel pdiffusion 780 -2050 780 -2050 0 feedthrough
rlabel pdiffusion 787 -2050 787 -2050 0 feedthrough
rlabel pdiffusion 794 -2050 794 -2050 0 feedthrough
rlabel pdiffusion 801 -2050 801 -2050 0 feedthrough
rlabel pdiffusion 808 -2050 808 -2050 0 feedthrough
rlabel pdiffusion 815 -2050 815 -2050 0 cellNo=146
rlabel pdiffusion 822 -2050 822 -2050 0 feedthrough
rlabel pdiffusion 829 -2050 829 -2050 0 feedthrough
rlabel pdiffusion 836 -2050 836 -2050 0 feedthrough
rlabel pdiffusion 843 -2050 843 -2050 0 cellNo=115
rlabel pdiffusion 850 -2050 850 -2050 0 cellNo=177
rlabel pdiffusion 857 -2050 857 -2050 0 feedthrough
rlabel pdiffusion 864 -2050 864 -2050 0 cellNo=51
rlabel pdiffusion 871 -2050 871 -2050 0 feedthrough
rlabel pdiffusion 878 -2050 878 -2050 0 cellNo=69
rlabel pdiffusion 885 -2050 885 -2050 0 feedthrough
rlabel pdiffusion 892 -2050 892 -2050 0 cellNo=213
rlabel pdiffusion 899 -2050 899 -2050 0 feedthrough
rlabel pdiffusion 906 -2050 906 -2050 0 feedthrough
rlabel pdiffusion 913 -2050 913 -2050 0 feedthrough
rlabel pdiffusion 920 -2050 920 -2050 0 cellNo=83
rlabel pdiffusion 927 -2050 927 -2050 0 feedthrough
rlabel pdiffusion 934 -2050 934 -2050 0 feedthrough
rlabel pdiffusion 941 -2050 941 -2050 0 feedthrough
rlabel pdiffusion 948 -2050 948 -2050 0 feedthrough
rlabel pdiffusion 955 -2050 955 -2050 0 feedthrough
rlabel pdiffusion 962 -2050 962 -2050 0 cellNo=66
rlabel pdiffusion 969 -2050 969 -2050 0 cellNo=926
rlabel pdiffusion 976 -2050 976 -2050 0 feedthrough
rlabel pdiffusion 983 -2050 983 -2050 0 feedthrough
rlabel pdiffusion 990 -2050 990 -2050 0 feedthrough
rlabel pdiffusion 997 -2050 997 -2050 0 feedthrough
rlabel pdiffusion 1004 -2050 1004 -2050 0 feedthrough
rlabel pdiffusion 1011 -2050 1011 -2050 0 feedthrough
rlabel pdiffusion 1018 -2050 1018 -2050 0 feedthrough
rlabel pdiffusion 1025 -2050 1025 -2050 0 feedthrough
rlabel pdiffusion 1032 -2050 1032 -2050 0 feedthrough
rlabel pdiffusion 1039 -2050 1039 -2050 0 feedthrough
rlabel pdiffusion 1046 -2050 1046 -2050 0 feedthrough
rlabel pdiffusion 1053 -2050 1053 -2050 0 feedthrough
rlabel pdiffusion 1060 -2050 1060 -2050 0 feedthrough
rlabel pdiffusion 1067 -2050 1067 -2050 0 feedthrough
rlabel pdiffusion 1074 -2050 1074 -2050 0 feedthrough
rlabel pdiffusion 1081 -2050 1081 -2050 0 feedthrough
rlabel pdiffusion 1088 -2050 1088 -2050 0 cellNo=389
rlabel pdiffusion 1095 -2050 1095 -2050 0 feedthrough
rlabel pdiffusion 1102 -2050 1102 -2050 0 feedthrough
rlabel pdiffusion 1109 -2050 1109 -2050 0 cellNo=365
rlabel pdiffusion 1116 -2050 1116 -2050 0 feedthrough
rlabel pdiffusion 1123 -2050 1123 -2050 0 feedthrough
rlabel pdiffusion 1130 -2050 1130 -2050 0 feedthrough
rlabel pdiffusion 1137 -2050 1137 -2050 0 feedthrough
rlabel pdiffusion 1144 -2050 1144 -2050 0 feedthrough
rlabel pdiffusion 1151 -2050 1151 -2050 0 feedthrough
rlabel pdiffusion 1158 -2050 1158 -2050 0 feedthrough
rlabel pdiffusion 1165 -2050 1165 -2050 0 feedthrough
rlabel pdiffusion 1172 -2050 1172 -2050 0 feedthrough
rlabel pdiffusion 1179 -2050 1179 -2050 0 feedthrough
rlabel pdiffusion 1186 -2050 1186 -2050 0 feedthrough
rlabel pdiffusion 1193 -2050 1193 -2050 0 cellNo=290
rlabel pdiffusion 1200 -2050 1200 -2050 0 feedthrough
rlabel pdiffusion 1207 -2050 1207 -2050 0 feedthrough
rlabel pdiffusion 1214 -2050 1214 -2050 0 feedthrough
rlabel pdiffusion 1221 -2050 1221 -2050 0 feedthrough
rlabel pdiffusion 1228 -2050 1228 -2050 0 feedthrough
rlabel pdiffusion 1235 -2050 1235 -2050 0 cellNo=628
rlabel pdiffusion 1242 -2050 1242 -2050 0 feedthrough
rlabel pdiffusion 1249 -2050 1249 -2050 0 feedthrough
rlabel pdiffusion 1256 -2050 1256 -2050 0 cellNo=127
rlabel pdiffusion 1263 -2050 1263 -2050 0 cellNo=836
rlabel pdiffusion 1270 -2050 1270 -2050 0 feedthrough
rlabel pdiffusion 1277 -2050 1277 -2050 0 feedthrough
rlabel pdiffusion 1284 -2050 1284 -2050 0 feedthrough
rlabel pdiffusion 1291 -2050 1291 -2050 0 cellNo=378
rlabel pdiffusion 1298 -2050 1298 -2050 0 feedthrough
rlabel pdiffusion 1305 -2050 1305 -2050 0 feedthrough
rlabel pdiffusion 1312 -2050 1312 -2050 0 feedthrough
rlabel pdiffusion 1319 -2050 1319 -2050 0 feedthrough
rlabel pdiffusion 1326 -2050 1326 -2050 0 feedthrough
rlabel pdiffusion 1333 -2050 1333 -2050 0 feedthrough
rlabel pdiffusion 1340 -2050 1340 -2050 0 feedthrough
rlabel pdiffusion 1347 -2050 1347 -2050 0 feedthrough
rlabel pdiffusion 1354 -2050 1354 -2050 0 feedthrough
rlabel pdiffusion 1361 -2050 1361 -2050 0 feedthrough
rlabel pdiffusion 1368 -2050 1368 -2050 0 feedthrough
rlabel pdiffusion 1375 -2050 1375 -2050 0 feedthrough
rlabel pdiffusion 1382 -2050 1382 -2050 0 feedthrough
rlabel pdiffusion 1389 -2050 1389 -2050 0 feedthrough
rlabel pdiffusion 1396 -2050 1396 -2050 0 feedthrough
rlabel pdiffusion 1403 -2050 1403 -2050 0 feedthrough
rlabel pdiffusion 1410 -2050 1410 -2050 0 feedthrough
rlabel pdiffusion 1417 -2050 1417 -2050 0 feedthrough
rlabel pdiffusion 1424 -2050 1424 -2050 0 feedthrough
rlabel pdiffusion 1431 -2050 1431 -2050 0 feedthrough
rlabel pdiffusion 1438 -2050 1438 -2050 0 feedthrough
rlabel pdiffusion 1445 -2050 1445 -2050 0 feedthrough
rlabel pdiffusion 1452 -2050 1452 -2050 0 cellNo=690
rlabel pdiffusion 1459 -2050 1459 -2050 0 feedthrough
rlabel pdiffusion 1466 -2050 1466 -2050 0 feedthrough
rlabel pdiffusion 1473 -2050 1473 -2050 0 feedthrough
rlabel pdiffusion 1480 -2050 1480 -2050 0 feedthrough
rlabel pdiffusion 1487 -2050 1487 -2050 0 feedthrough
rlabel pdiffusion 1494 -2050 1494 -2050 0 feedthrough
rlabel pdiffusion 1501 -2050 1501 -2050 0 feedthrough
rlabel pdiffusion 1508 -2050 1508 -2050 0 feedthrough
rlabel pdiffusion 1515 -2050 1515 -2050 0 feedthrough
rlabel pdiffusion 1522 -2050 1522 -2050 0 feedthrough
rlabel pdiffusion 1529 -2050 1529 -2050 0 feedthrough
rlabel pdiffusion 1536 -2050 1536 -2050 0 feedthrough
rlabel pdiffusion 1543 -2050 1543 -2050 0 feedthrough
rlabel pdiffusion 1550 -2050 1550 -2050 0 feedthrough
rlabel pdiffusion 1557 -2050 1557 -2050 0 feedthrough
rlabel pdiffusion 1564 -2050 1564 -2050 0 feedthrough
rlabel pdiffusion 1571 -2050 1571 -2050 0 feedthrough
rlabel pdiffusion 1578 -2050 1578 -2050 0 feedthrough
rlabel pdiffusion 1585 -2050 1585 -2050 0 feedthrough
rlabel pdiffusion 1592 -2050 1592 -2050 0 feedthrough
rlabel pdiffusion 1599 -2050 1599 -2050 0 feedthrough
rlabel pdiffusion 1606 -2050 1606 -2050 0 feedthrough
rlabel pdiffusion 1613 -2050 1613 -2050 0 feedthrough
rlabel pdiffusion 1620 -2050 1620 -2050 0 feedthrough
rlabel pdiffusion 1627 -2050 1627 -2050 0 feedthrough
rlabel pdiffusion 1634 -2050 1634 -2050 0 feedthrough
rlabel pdiffusion 1641 -2050 1641 -2050 0 feedthrough
rlabel pdiffusion 1648 -2050 1648 -2050 0 feedthrough
rlabel pdiffusion 1655 -2050 1655 -2050 0 feedthrough
rlabel pdiffusion 1662 -2050 1662 -2050 0 feedthrough
rlabel pdiffusion 1669 -2050 1669 -2050 0 feedthrough
rlabel pdiffusion 1676 -2050 1676 -2050 0 feedthrough
rlabel pdiffusion 1683 -2050 1683 -2050 0 feedthrough
rlabel pdiffusion 1690 -2050 1690 -2050 0 feedthrough
rlabel pdiffusion 1697 -2050 1697 -2050 0 feedthrough
rlabel pdiffusion 1704 -2050 1704 -2050 0 feedthrough
rlabel pdiffusion 1711 -2050 1711 -2050 0 feedthrough
rlabel pdiffusion 1718 -2050 1718 -2050 0 feedthrough
rlabel pdiffusion 1725 -2050 1725 -2050 0 feedthrough
rlabel pdiffusion 1732 -2050 1732 -2050 0 feedthrough
rlabel pdiffusion 1739 -2050 1739 -2050 0 feedthrough
rlabel pdiffusion 1746 -2050 1746 -2050 0 feedthrough
rlabel pdiffusion 1753 -2050 1753 -2050 0 feedthrough
rlabel pdiffusion 1760 -2050 1760 -2050 0 feedthrough
rlabel pdiffusion 1767 -2050 1767 -2050 0 feedthrough
rlabel pdiffusion 1774 -2050 1774 -2050 0 feedthrough
rlabel pdiffusion 1781 -2050 1781 -2050 0 feedthrough
rlabel pdiffusion 1788 -2050 1788 -2050 0 feedthrough
rlabel pdiffusion 1795 -2050 1795 -2050 0 feedthrough
rlabel pdiffusion 1802 -2050 1802 -2050 0 feedthrough
rlabel pdiffusion 1809 -2050 1809 -2050 0 feedthrough
rlabel pdiffusion 1816 -2050 1816 -2050 0 feedthrough
rlabel pdiffusion 1823 -2050 1823 -2050 0 feedthrough
rlabel pdiffusion 1830 -2050 1830 -2050 0 feedthrough
rlabel pdiffusion 1837 -2050 1837 -2050 0 feedthrough
rlabel pdiffusion 1844 -2050 1844 -2050 0 feedthrough
rlabel pdiffusion 1851 -2050 1851 -2050 0 feedthrough
rlabel pdiffusion 1858 -2050 1858 -2050 0 feedthrough
rlabel pdiffusion 1865 -2050 1865 -2050 0 feedthrough
rlabel pdiffusion 1872 -2050 1872 -2050 0 feedthrough
rlabel pdiffusion 1879 -2050 1879 -2050 0 feedthrough
rlabel pdiffusion 1886 -2050 1886 -2050 0 feedthrough
rlabel pdiffusion 1893 -2050 1893 -2050 0 feedthrough
rlabel pdiffusion 1900 -2050 1900 -2050 0 feedthrough
rlabel pdiffusion 1907 -2050 1907 -2050 0 feedthrough
rlabel pdiffusion 1914 -2050 1914 -2050 0 feedthrough
rlabel pdiffusion 1921 -2050 1921 -2050 0 cellNo=726
rlabel pdiffusion 1928 -2050 1928 -2050 0 feedthrough
rlabel pdiffusion 1935 -2050 1935 -2050 0 feedthrough
rlabel pdiffusion 1942 -2050 1942 -2050 0 feedthrough
rlabel pdiffusion 1949 -2050 1949 -2050 0 feedthrough
rlabel pdiffusion 1956 -2050 1956 -2050 0 feedthrough
rlabel pdiffusion 1963 -2050 1963 -2050 0 feedthrough
rlabel pdiffusion 1970 -2050 1970 -2050 0 feedthrough
rlabel pdiffusion 1977 -2050 1977 -2050 0 feedthrough
rlabel pdiffusion 1984 -2050 1984 -2050 0 feedthrough
rlabel pdiffusion 1991 -2050 1991 -2050 0 feedthrough
rlabel pdiffusion 3 -2191 3 -2191 0 feedthrough
rlabel pdiffusion 10 -2191 10 -2191 0 cellNo=547
rlabel pdiffusion 17 -2191 17 -2191 0 feedthrough
rlabel pdiffusion 24 -2191 24 -2191 0 feedthrough
rlabel pdiffusion 31 -2191 31 -2191 0 cellNo=749
rlabel pdiffusion 38 -2191 38 -2191 0 cellNo=526
rlabel pdiffusion 45 -2191 45 -2191 0 feedthrough
rlabel pdiffusion 52 -2191 52 -2191 0 feedthrough
rlabel pdiffusion 59 -2191 59 -2191 0 feedthrough
rlabel pdiffusion 66 -2191 66 -2191 0 feedthrough
rlabel pdiffusion 73 -2191 73 -2191 0 feedthrough
rlabel pdiffusion 80 -2191 80 -2191 0 feedthrough
rlabel pdiffusion 87 -2191 87 -2191 0 cellNo=522
rlabel pdiffusion 94 -2191 94 -2191 0 cellNo=203
rlabel pdiffusion 101 -2191 101 -2191 0 feedthrough
rlabel pdiffusion 108 -2191 108 -2191 0 cellNo=844
rlabel pdiffusion 115 -2191 115 -2191 0 cellNo=1183
rlabel pdiffusion 122 -2191 122 -2191 0 feedthrough
rlabel pdiffusion 129 -2191 129 -2191 0 feedthrough
rlabel pdiffusion 136 -2191 136 -2191 0 feedthrough
rlabel pdiffusion 143 -2191 143 -2191 0 feedthrough
rlabel pdiffusion 150 -2191 150 -2191 0 feedthrough
rlabel pdiffusion 157 -2191 157 -2191 0 feedthrough
rlabel pdiffusion 164 -2191 164 -2191 0 feedthrough
rlabel pdiffusion 171 -2191 171 -2191 0 feedthrough
rlabel pdiffusion 178 -2191 178 -2191 0 feedthrough
rlabel pdiffusion 185 -2191 185 -2191 0 feedthrough
rlabel pdiffusion 192 -2191 192 -2191 0 feedthrough
rlabel pdiffusion 199 -2191 199 -2191 0 feedthrough
rlabel pdiffusion 206 -2191 206 -2191 0 feedthrough
rlabel pdiffusion 213 -2191 213 -2191 0 feedthrough
rlabel pdiffusion 220 -2191 220 -2191 0 feedthrough
rlabel pdiffusion 227 -2191 227 -2191 0 feedthrough
rlabel pdiffusion 234 -2191 234 -2191 0 cellNo=34
rlabel pdiffusion 241 -2191 241 -2191 0 feedthrough
rlabel pdiffusion 248 -2191 248 -2191 0 feedthrough
rlabel pdiffusion 255 -2191 255 -2191 0 feedthrough
rlabel pdiffusion 262 -2191 262 -2191 0 feedthrough
rlabel pdiffusion 269 -2191 269 -2191 0 feedthrough
rlabel pdiffusion 276 -2191 276 -2191 0 feedthrough
rlabel pdiffusion 283 -2191 283 -2191 0 feedthrough
rlabel pdiffusion 290 -2191 290 -2191 0 feedthrough
rlabel pdiffusion 297 -2191 297 -2191 0 feedthrough
rlabel pdiffusion 304 -2191 304 -2191 0 feedthrough
rlabel pdiffusion 311 -2191 311 -2191 0 feedthrough
rlabel pdiffusion 318 -2191 318 -2191 0 feedthrough
rlabel pdiffusion 325 -2191 325 -2191 0 feedthrough
rlabel pdiffusion 332 -2191 332 -2191 0 feedthrough
rlabel pdiffusion 339 -2191 339 -2191 0 cellNo=810
rlabel pdiffusion 346 -2191 346 -2191 0 feedthrough
rlabel pdiffusion 353 -2191 353 -2191 0 feedthrough
rlabel pdiffusion 360 -2191 360 -2191 0 feedthrough
rlabel pdiffusion 367 -2191 367 -2191 0 feedthrough
rlabel pdiffusion 374 -2191 374 -2191 0 feedthrough
rlabel pdiffusion 381 -2191 381 -2191 0 feedthrough
rlabel pdiffusion 388 -2191 388 -2191 0 cellNo=601
rlabel pdiffusion 395 -2191 395 -2191 0 feedthrough
rlabel pdiffusion 402 -2191 402 -2191 0 cellNo=678
rlabel pdiffusion 409 -2191 409 -2191 0 feedthrough
rlabel pdiffusion 416 -2191 416 -2191 0 feedthrough
rlabel pdiffusion 423 -2191 423 -2191 0 feedthrough
rlabel pdiffusion 430 -2191 430 -2191 0 feedthrough
rlabel pdiffusion 437 -2191 437 -2191 0 cellNo=185
rlabel pdiffusion 444 -2191 444 -2191 0 feedthrough
rlabel pdiffusion 451 -2191 451 -2191 0 feedthrough
rlabel pdiffusion 458 -2191 458 -2191 0 feedthrough
rlabel pdiffusion 465 -2191 465 -2191 0 cellNo=79
rlabel pdiffusion 472 -2191 472 -2191 0 feedthrough
rlabel pdiffusion 479 -2191 479 -2191 0 feedthrough
rlabel pdiffusion 486 -2191 486 -2191 0 feedthrough
rlabel pdiffusion 493 -2191 493 -2191 0 feedthrough
rlabel pdiffusion 500 -2191 500 -2191 0 feedthrough
rlabel pdiffusion 507 -2191 507 -2191 0 cellNo=969
rlabel pdiffusion 514 -2191 514 -2191 0 feedthrough
rlabel pdiffusion 521 -2191 521 -2191 0 feedthrough
rlabel pdiffusion 528 -2191 528 -2191 0 feedthrough
rlabel pdiffusion 535 -2191 535 -2191 0 feedthrough
rlabel pdiffusion 542 -2191 542 -2191 0 cellNo=959
rlabel pdiffusion 549 -2191 549 -2191 0 feedthrough
rlabel pdiffusion 556 -2191 556 -2191 0 feedthrough
rlabel pdiffusion 563 -2191 563 -2191 0 feedthrough
rlabel pdiffusion 570 -2191 570 -2191 0 feedthrough
rlabel pdiffusion 577 -2191 577 -2191 0 feedthrough
rlabel pdiffusion 584 -2191 584 -2191 0 feedthrough
rlabel pdiffusion 591 -2191 591 -2191 0 cellNo=231
rlabel pdiffusion 598 -2191 598 -2191 0 feedthrough
rlabel pdiffusion 605 -2191 605 -2191 0 feedthrough
rlabel pdiffusion 612 -2191 612 -2191 0 feedthrough
rlabel pdiffusion 619 -2191 619 -2191 0 feedthrough
rlabel pdiffusion 626 -2191 626 -2191 0 cellNo=483
rlabel pdiffusion 633 -2191 633 -2191 0 feedthrough
rlabel pdiffusion 640 -2191 640 -2191 0 feedthrough
rlabel pdiffusion 647 -2191 647 -2191 0 cellNo=804
rlabel pdiffusion 654 -2191 654 -2191 0 feedthrough
rlabel pdiffusion 661 -2191 661 -2191 0 feedthrough
rlabel pdiffusion 668 -2191 668 -2191 0 feedthrough
rlabel pdiffusion 675 -2191 675 -2191 0 feedthrough
rlabel pdiffusion 682 -2191 682 -2191 0 feedthrough
rlabel pdiffusion 689 -2191 689 -2191 0 feedthrough
rlabel pdiffusion 696 -2191 696 -2191 0 feedthrough
rlabel pdiffusion 703 -2191 703 -2191 0 feedthrough
rlabel pdiffusion 710 -2191 710 -2191 0 feedthrough
rlabel pdiffusion 717 -2191 717 -2191 0 feedthrough
rlabel pdiffusion 724 -2191 724 -2191 0 feedthrough
rlabel pdiffusion 731 -2191 731 -2191 0 feedthrough
rlabel pdiffusion 738 -2191 738 -2191 0 feedthrough
rlabel pdiffusion 745 -2191 745 -2191 0 feedthrough
rlabel pdiffusion 752 -2191 752 -2191 0 feedthrough
rlabel pdiffusion 759 -2191 759 -2191 0 feedthrough
rlabel pdiffusion 766 -2191 766 -2191 0 feedthrough
rlabel pdiffusion 773 -2191 773 -2191 0 feedthrough
rlabel pdiffusion 780 -2191 780 -2191 0 feedthrough
rlabel pdiffusion 787 -2191 787 -2191 0 feedthrough
rlabel pdiffusion 794 -2191 794 -2191 0 feedthrough
rlabel pdiffusion 801 -2191 801 -2191 0 feedthrough
rlabel pdiffusion 808 -2191 808 -2191 0 feedthrough
rlabel pdiffusion 815 -2191 815 -2191 0 feedthrough
rlabel pdiffusion 822 -2191 822 -2191 0 feedthrough
rlabel pdiffusion 829 -2191 829 -2191 0 feedthrough
rlabel pdiffusion 836 -2191 836 -2191 0 cellNo=184
rlabel pdiffusion 843 -2191 843 -2191 0 feedthrough
rlabel pdiffusion 850 -2191 850 -2191 0 feedthrough
rlabel pdiffusion 857 -2191 857 -2191 0 feedthrough
rlabel pdiffusion 864 -2191 864 -2191 0 feedthrough
rlabel pdiffusion 871 -2191 871 -2191 0 feedthrough
rlabel pdiffusion 878 -2191 878 -2191 0 cellNo=117
rlabel pdiffusion 885 -2191 885 -2191 0 feedthrough
rlabel pdiffusion 892 -2191 892 -2191 0 feedthrough
rlabel pdiffusion 899 -2191 899 -2191 0 feedthrough
rlabel pdiffusion 906 -2191 906 -2191 0 feedthrough
rlabel pdiffusion 913 -2191 913 -2191 0 feedthrough
rlabel pdiffusion 920 -2191 920 -2191 0 feedthrough
rlabel pdiffusion 927 -2191 927 -2191 0 feedthrough
rlabel pdiffusion 934 -2191 934 -2191 0 feedthrough
rlabel pdiffusion 941 -2191 941 -2191 0 feedthrough
rlabel pdiffusion 948 -2191 948 -2191 0 feedthrough
rlabel pdiffusion 955 -2191 955 -2191 0 feedthrough
rlabel pdiffusion 962 -2191 962 -2191 0 feedthrough
rlabel pdiffusion 969 -2191 969 -2191 0 cellNo=650
rlabel pdiffusion 976 -2191 976 -2191 0 cellNo=315
rlabel pdiffusion 983 -2191 983 -2191 0 feedthrough
rlabel pdiffusion 990 -2191 990 -2191 0 feedthrough
rlabel pdiffusion 997 -2191 997 -2191 0 feedthrough
rlabel pdiffusion 1004 -2191 1004 -2191 0 feedthrough
rlabel pdiffusion 1011 -2191 1011 -2191 0 feedthrough
rlabel pdiffusion 1018 -2191 1018 -2191 0 feedthrough
rlabel pdiffusion 1025 -2191 1025 -2191 0 feedthrough
rlabel pdiffusion 1032 -2191 1032 -2191 0 feedthrough
rlabel pdiffusion 1039 -2191 1039 -2191 0 feedthrough
rlabel pdiffusion 1046 -2191 1046 -2191 0 feedthrough
rlabel pdiffusion 1053 -2191 1053 -2191 0 cellNo=599
rlabel pdiffusion 1060 -2191 1060 -2191 0 feedthrough
rlabel pdiffusion 1067 -2191 1067 -2191 0 cellNo=653
rlabel pdiffusion 1074 -2191 1074 -2191 0 feedthrough
rlabel pdiffusion 1081 -2191 1081 -2191 0 cellNo=873
rlabel pdiffusion 1088 -2191 1088 -2191 0 feedthrough
rlabel pdiffusion 1095 -2191 1095 -2191 0 feedthrough
rlabel pdiffusion 1102 -2191 1102 -2191 0 feedthrough
rlabel pdiffusion 1109 -2191 1109 -2191 0 cellNo=825
rlabel pdiffusion 1116 -2191 1116 -2191 0 feedthrough
rlabel pdiffusion 1123 -2191 1123 -2191 0 feedthrough
rlabel pdiffusion 1130 -2191 1130 -2191 0 feedthrough
rlabel pdiffusion 1137 -2191 1137 -2191 0 cellNo=908
rlabel pdiffusion 1144 -2191 1144 -2191 0 feedthrough
rlabel pdiffusion 1151 -2191 1151 -2191 0 feedthrough
rlabel pdiffusion 1158 -2191 1158 -2191 0 cellNo=248
rlabel pdiffusion 1165 -2191 1165 -2191 0 feedthrough
rlabel pdiffusion 1172 -2191 1172 -2191 0 feedthrough
rlabel pdiffusion 1179 -2191 1179 -2191 0 feedthrough
rlabel pdiffusion 1186 -2191 1186 -2191 0 feedthrough
rlabel pdiffusion 1193 -2191 1193 -2191 0 feedthrough
rlabel pdiffusion 1200 -2191 1200 -2191 0 feedthrough
rlabel pdiffusion 1207 -2191 1207 -2191 0 feedthrough
rlabel pdiffusion 1214 -2191 1214 -2191 0 feedthrough
rlabel pdiffusion 1221 -2191 1221 -2191 0 feedthrough
rlabel pdiffusion 1228 -2191 1228 -2191 0 feedthrough
rlabel pdiffusion 1235 -2191 1235 -2191 0 feedthrough
rlabel pdiffusion 1242 -2191 1242 -2191 0 feedthrough
rlabel pdiffusion 1249 -2191 1249 -2191 0 feedthrough
rlabel pdiffusion 1256 -2191 1256 -2191 0 feedthrough
rlabel pdiffusion 1263 -2191 1263 -2191 0 feedthrough
rlabel pdiffusion 1270 -2191 1270 -2191 0 feedthrough
rlabel pdiffusion 1277 -2191 1277 -2191 0 cellNo=476
rlabel pdiffusion 1284 -2191 1284 -2191 0 feedthrough
rlabel pdiffusion 1291 -2191 1291 -2191 0 feedthrough
rlabel pdiffusion 1298 -2191 1298 -2191 0 feedthrough
rlabel pdiffusion 1305 -2191 1305 -2191 0 feedthrough
rlabel pdiffusion 1312 -2191 1312 -2191 0 feedthrough
rlabel pdiffusion 1319 -2191 1319 -2191 0 feedthrough
rlabel pdiffusion 1326 -2191 1326 -2191 0 feedthrough
rlabel pdiffusion 1333 -2191 1333 -2191 0 feedthrough
rlabel pdiffusion 1340 -2191 1340 -2191 0 feedthrough
rlabel pdiffusion 1347 -2191 1347 -2191 0 feedthrough
rlabel pdiffusion 1354 -2191 1354 -2191 0 feedthrough
rlabel pdiffusion 1361 -2191 1361 -2191 0 cellNo=212
rlabel pdiffusion 1368 -2191 1368 -2191 0 feedthrough
rlabel pdiffusion 1375 -2191 1375 -2191 0 cellNo=5
rlabel pdiffusion 1382 -2191 1382 -2191 0 feedthrough
rlabel pdiffusion 1389 -2191 1389 -2191 0 feedthrough
rlabel pdiffusion 1396 -2191 1396 -2191 0 cellNo=60
rlabel pdiffusion 1403 -2191 1403 -2191 0 cellNo=635
rlabel pdiffusion 1410 -2191 1410 -2191 0 feedthrough
rlabel pdiffusion 1417 -2191 1417 -2191 0 feedthrough
rlabel pdiffusion 1424 -2191 1424 -2191 0 feedthrough
rlabel pdiffusion 1431 -2191 1431 -2191 0 feedthrough
rlabel pdiffusion 1438 -2191 1438 -2191 0 feedthrough
rlabel pdiffusion 1445 -2191 1445 -2191 0 feedthrough
rlabel pdiffusion 1452 -2191 1452 -2191 0 cellNo=256
rlabel pdiffusion 1459 -2191 1459 -2191 0 feedthrough
rlabel pdiffusion 1466 -2191 1466 -2191 0 feedthrough
rlabel pdiffusion 1473 -2191 1473 -2191 0 cellNo=65
rlabel pdiffusion 1480 -2191 1480 -2191 0 feedthrough
rlabel pdiffusion 1487 -2191 1487 -2191 0 feedthrough
rlabel pdiffusion 1494 -2191 1494 -2191 0 feedthrough
rlabel pdiffusion 1501 -2191 1501 -2191 0 feedthrough
rlabel pdiffusion 1508 -2191 1508 -2191 0 feedthrough
rlabel pdiffusion 1515 -2191 1515 -2191 0 feedthrough
rlabel pdiffusion 1522 -2191 1522 -2191 0 feedthrough
rlabel pdiffusion 1529 -2191 1529 -2191 0 feedthrough
rlabel pdiffusion 1536 -2191 1536 -2191 0 feedthrough
rlabel pdiffusion 1543 -2191 1543 -2191 0 feedthrough
rlabel pdiffusion 1550 -2191 1550 -2191 0 feedthrough
rlabel pdiffusion 1557 -2191 1557 -2191 0 feedthrough
rlabel pdiffusion 1564 -2191 1564 -2191 0 feedthrough
rlabel pdiffusion 1571 -2191 1571 -2191 0 feedthrough
rlabel pdiffusion 1578 -2191 1578 -2191 0 feedthrough
rlabel pdiffusion 1585 -2191 1585 -2191 0 feedthrough
rlabel pdiffusion 1592 -2191 1592 -2191 0 feedthrough
rlabel pdiffusion 1599 -2191 1599 -2191 0 feedthrough
rlabel pdiffusion 1606 -2191 1606 -2191 0 feedthrough
rlabel pdiffusion 1613 -2191 1613 -2191 0 feedthrough
rlabel pdiffusion 1620 -2191 1620 -2191 0 feedthrough
rlabel pdiffusion 1627 -2191 1627 -2191 0 feedthrough
rlabel pdiffusion 1634 -2191 1634 -2191 0 feedthrough
rlabel pdiffusion 1641 -2191 1641 -2191 0 feedthrough
rlabel pdiffusion 1648 -2191 1648 -2191 0 feedthrough
rlabel pdiffusion 1655 -2191 1655 -2191 0 feedthrough
rlabel pdiffusion 1662 -2191 1662 -2191 0 feedthrough
rlabel pdiffusion 1669 -2191 1669 -2191 0 feedthrough
rlabel pdiffusion 1676 -2191 1676 -2191 0 feedthrough
rlabel pdiffusion 1683 -2191 1683 -2191 0 feedthrough
rlabel pdiffusion 1690 -2191 1690 -2191 0 feedthrough
rlabel pdiffusion 1697 -2191 1697 -2191 0 feedthrough
rlabel pdiffusion 1704 -2191 1704 -2191 0 feedthrough
rlabel pdiffusion 1711 -2191 1711 -2191 0 feedthrough
rlabel pdiffusion 1718 -2191 1718 -2191 0 feedthrough
rlabel pdiffusion 1725 -2191 1725 -2191 0 feedthrough
rlabel pdiffusion 1732 -2191 1732 -2191 0 feedthrough
rlabel pdiffusion 1739 -2191 1739 -2191 0 feedthrough
rlabel pdiffusion 1746 -2191 1746 -2191 0 feedthrough
rlabel pdiffusion 1753 -2191 1753 -2191 0 feedthrough
rlabel pdiffusion 1760 -2191 1760 -2191 0 feedthrough
rlabel pdiffusion 1767 -2191 1767 -2191 0 feedthrough
rlabel pdiffusion 1774 -2191 1774 -2191 0 feedthrough
rlabel pdiffusion 1781 -2191 1781 -2191 0 feedthrough
rlabel pdiffusion 1788 -2191 1788 -2191 0 feedthrough
rlabel pdiffusion 1795 -2191 1795 -2191 0 feedthrough
rlabel pdiffusion 1802 -2191 1802 -2191 0 feedthrough
rlabel pdiffusion 1809 -2191 1809 -2191 0 feedthrough
rlabel pdiffusion 1816 -2191 1816 -2191 0 feedthrough
rlabel pdiffusion 1823 -2191 1823 -2191 0 feedthrough
rlabel pdiffusion 1830 -2191 1830 -2191 0 feedthrough
rlabel pdiffusion 1837 -2191 1837 -2191 0 feedthrough
rlabel pdiffusion 1844 -2191 1844 -2191 0 feedthrough
rlabel pdiffusion 1851 -2191 1851 -2191 0 feedthrough
rlabel pdiffusion 1858 -2191 1858 -2191 0 feedthrough
rlabel pdiffusion 1865 -2191 1865 -2191 0 feedthrough
rlabel pdiffusion 1872 -2191 1872 -2191 0 feedthrough
rlabel pdiffusion 1879 -2191 1879 -2191 0 feedthrough
rlabel pdiffusion 1886 -2191 1886 -2191 0 feedthrough
rlabel pdiffusion 1893 -2191 1893 -2191 0 feedthrough
rlabel pdiffusion 1900 -2191 1900 -2191 0 feedthrough
rlabel pdiffusion 1907 -2191 1907 -2191 0 feedthrough
rlabel pdiffusion 1914 -2191 1914 -2191 0 feedthrough
rlabel pdiffusion 3 -2320 3 -2320 0 cellNo=1031
rlabel pdiffusion 10 -2320 10 -2320 0 feedthrough
rlabel pdiffusion 17 -2320 17 -2320 0 cellNo=746
rlabel pdiffusion 24 -2320 24 -2320 0 feedthrough
rlabel pdiffusion 31 -2320 31 -2320 0 feedthrough
rlabel pdiffusion 38 -2320 38 -2320 0 feedthrough
rlabel pdiffusion 45 -2320 45 -2320 0 feedthrough
rlabel pdiffusion 52 -2320 52 -2320 0 feedthrough
rlabel pdiffusion 59 -2320 59 -2320 0 feedthrough
rlabel pdiffusion 66 -2320 66 -2320 0 cellNo=135
rlabel pdiffusion 73 -2320 73 -2320 0 feedthrough
rlabel pdiffusion 80 -2320 80 -2320 0 feedthrough
rlabel pdiffusion 87 -2320 87 -2320 0 feedthrough
rlabel pdiffusion 94 -2320 94 -2320 0 feedthrough
rlabel pdiffusion 101 -2320 101 -2320 0 feedthrough
rlabel pdiffusion 108 -2320 108 -2320 0 feedthrough
rlabel pdiffusion 115 -2320 115 -2320 0 cellNo=13
rlabel pdiffusion 122 -2320 122 -2320 0 cellNo=828
rlabel pdiffusion 129 -2320 129 -2320 0 feedthrough
rlabel pdiffusion 136 -2320 136 -2320 0 feedthrough
rlabel pdiffusion 143 -2320 143 -2320 0 feedthrough
rlabel pdiffusion 150 -2320 150 -2320 0 feedthrough
rlabel pdiffusion 157 -2320 157 -2320 0 cellNo=704
rlabel pdiffusion 164 -2320 164 -2320 0 feedthrough
rlabel pdiffusion 171 -2320 171 -2320 0 cellNo=524
rlabel pdiffusion 178 -2320 178 -2320 0 feedthrough
rlabel pdiffusion 185 -2320 185 -2320 0 feedthrough
rlabel pdiffusion 192 -2320 192 -2320 0 feedthrough
rlabel pdiffusion 199 -2320 199 -2320 0 feedthrough
rlabel pdiffusion 206 -2320 206 -2320 0 cellNo=731
rlabel pdiffusion 213 -2320 213 -2320 0 cellNo=263
rlabel pdiffusion 220 -2320 220 -2320 0 cellNo=137
rlabel pdiffusion 227 -2320 227 -2320 0 feedthrough
rlabel pdiffusion 234 -2320 234 -2320 0 cellNo=35
rlabel pdiffusion 241 -2320 241 -2320 0 cellNo=917
rlabel pdiffusion 248 -2320 248 -2320 0 feedthrough
rlabel pdiffusion 255 -2320 255 -2320 0 feedthrough
rlabel pdiffusion 262 -2320 262 -2320 0 feedthrough
rlabel pdiffusion 269 -2320 269 -2320 0 feedthrough
rlabel pdiffusion 276 -2320 276 -2320 0 feedthrough
rlabel pdiffusion 283 -2320 283 -2320 0 feedthrough
rlabel pdiffusion 290 -2320 290 -2320 0 feedthrough
rlabel pdiffusion 297 -2320 297 -2320 0 feedthrough
rlabel pdiffusion 304 -2320 304 -2320 0 feedthrough
rlabel pdiffusion 311 -2320 311 -2320 0 feedthrough
rlabel pdiffusion 318 -2320 318 -2320 0 feedthrough
rlabel pdiffusion 325 -2320 325 -2320 0 feedthrough
rlabel pdiffusion 332 -2320 332 -2320 0 feedthrough
rlabel pdiffusion 339 -2320 339 -2320 0 feedthrough
rlabel pdiffusion 346 -2320 346 -2320 0 feedthrough
rlabel pdiffusion 353 -2320 353 -2320 0 feedthrough
rlabel pdiffusion 360 -2320 360 -2320 0 feedthrough
rlabel pdiffusion 367 -2320 367 -2320 0 feedthrough
rlabel pdiffusion 374 -2320 374 -2320 0 feedthrough
rlabel pdiffusion 381 -2320 381 -2320 0 feedthrough
rlabel pdiffusion 388 -2320 388 -2320 0 feedthrough
rlabel pdiffusion 395 -2320 395 -2320 0 feedthrough
rlabel pdiffusion 402 -2320 402 -2320 0 feedthrough
rlabel pdiffusion 409 -2320 409 -2320 0 feedthrough
rlabel pdiffusion 416 -2320 416 -2320 0 feedthrough
rlabel pdiffusion 423 -2320 423 -2320 0 feedthrough
rlabel pdiffusion 430 -2320 430 -2320 0 feedthrough
rlabel pdiffusion 437 -2320 437 -2320 0 feedthrough
rlabel pdiffusion 444 -2320 444 -2320 0 feedthrough
rlabel pdiffusion 451 -2320 451 -2320 0 feedthrough
rlabel pdiffusion 458 -2320 458 -2320 0 feedthrough
rlabel pdiffusion 465 -2320 465 -2320 0 cellNo=36
rlabel pdiffusion 472 -2320 472 -2320 0 feedthrough
rlabel pdiffusion 479 -2320 479 -2320 0 feedthrough
rlabel pdiffusion 486 -2320 486 -2320 0 feedthrough
rlabel pdiffusion 493 -2320 493 -2320 0 feedthrough
rlabel pdiffusion 500 -2320 500 -2320 0 feedthrough
rlabel pdiffusion 507 -2320 507 -2320 0 feedthrough
rlabel pdiffusion 514 -2320 514 -2320 0 feedthrough
rlabel pdiffusion 521 -2320 521 -2320 0 feedthrough
rlabel pdiffusion 528 -2320 528 -2320 0 feedthrough
rlabel pdiffusion 535 -2320 535 -2320 0 feedthrough
rlabel pdiffusion 542 -2320 542 -2320 0 feedthrough
rlabel pdiffusion 549 -2320 549 -2320 0 feedthrough
rlabel pdiffusion 556 -2320 556 -2320 0 feedthrough
rlabel pdiffusion 563 -2320 563 -2320 0 feedthrough
rlabel pdiffusion 570 -2320 570 -2320 0 cellNo=333
rlabel pdiffusion 577 -2320 577 -2320 0 feedthrough
rlabel pdiffusion 584 -2320 584 -2320 0 feedthrough
rlabel pdiffusion 591 -2320 591 -2320 0 feedthrough
rlabel pdiffusion 598 -2320 598 -2320 0 feedthrough
rlabel pdiffusion 605 -2320 605 -2320 0 feedthrough
rlabel pdiffusion 612 -2320 612 -2320 0 feedthrough
rlabel pdiffusion 619 -2320 619 -2320 0 feedthrough
rlabel pdiffusion 626 -2320 626 -2320 0 cellNo=622
rlabel pdiffusion 633 -2320 633 -2320 0 feedthrough
rlabel pdiffusion 640 -2320 640 -2320 0 feedthrough
rlabel pdiffusion 647 -2320 647 -2320 0 feedthrough
rlabel pdiffusion 654 -2320 654 -2320 0 cellNo=19
rlabel pdiffusion 661 -2320 661 -2320 0 feedthrough
rlabel pdiffusion 668 -2320 668 -2320 0 cellNo=896
rlabel pdiffusion 675 -2320 675 -2320 0 cellNo=82
rlabel pdiffusion 682 -2320 682 -2320 0 feedthrough
rlabel pdiffusion 689 -2320 689 -2320 0 feedthrough
rlabel pdiffusion 696 -2320 696 -2320 0 feedthrough
rlabel pdiffusion 703 -2320 703 -2320 0 feedthrough
rlabel pdiffusion 710 -2320 710 -2320 0 feedthrough
rlabel pdiffusion 717 -2320 717 -2320 0 feedthrough
rlabel pdiffusion 724 -2320 724 -2320 0 feedthrough
rlabel pdiffusion 731 -2320 731 -2320 0 feedthrough
rlabel pdiffusion 738 -2320 738 -2320 0 feedthrough
rlabel pdiffusion 745 -2320 745 -2320 0 feedthrough
rlabel pdiffusion 752 -2320 752 -2320 0 feedthrough
rlabel pdiffusion 759 -2320 759 -2320 0 cellNo=134
rlabel pdiffusion 766 -2320 766 -2320 0 feedthrough
rlabel pdiffusion 773 -2320 773 -2320 0 feedthrough
rlabel pdiffusion 780 -2320 780 -2320 0 feedthrough
rlabel pdiffusion 787 -2320 787 -2320 0 feedthrough
rlabel pdiffusion 794 -2320 794 -2320 0 cellNo=811
rlabel pdiffusion 801 -2320 801 -2320 0 feedthrough
rlabel pdiffusion 808 -2320 808 -2320 0 feedthrough
rlabel pdiffusion 815 -2320 815 -2320 0 cellNo=548
rlabel pdiffusion 822 -2320 822 -2320 0 cellNo=75
rlabel pdiffusion 829 -2320 829 -2320 0 feedthrough
rlabel pdiffusion 836 -2320 836 -2320 0 feedthrough
rlabel pdiffusion 843 -2320 843 -2320 0 feedthrough
rlabel pdiffusion 850 -2320 850 -2320 0 feedthrough
rlabel pdiffusion 857 -2320 857 -2320 0 feedthrough
rlabel pdiffusion 864 -2320 864 -2320 0 feedthrough
rlabel pdiffusion 871 -2320 871 -2320 0 feedthrough
rlabel pdiffusion 878 -2320 878 -2320 0 feedthrough
rlabel pdiffusion 885 -2320 885 -2320 0 cellNo=328
rlabel pdiffusion 892 -2320 892 -2320 0 feedthrough
rlabel pdiffusion 899 -2320 899 -2320 0 feedthrough
rlabel pdiffusion 906 -2320 906 -2320 0 feedthrough
rlabel pdiffusion 913 -2320 913 -2320 0 feedthrough
rlabel pdiffusion 920 -2320 920 -2320 0 feedthrough
rlabel pdiffusion 927 -2320 927 -2320 0 feedthrough
rlabel pdiffusion 934 -2320 934 -2320 0 feedthrough
rlabel pdiffusion 941 -2320 941 -2320 0 feedthrough
rlabel pdiffusion 948 -2320 948 -2320 0 cellNo=582
rlabel pdiffusion 955 -2320 955 -2320 0 feedthrough
rlabel pdiffusion 962 -2320 962 -2320 0 feedthrough
rlabel pdiffusion 969 -2320 969 -2320 0 feedthrough
rlabel pdiffusion 976 -2320 976 -2320 0 feedthrough
rlabel pdiffusion 983 -2320 983 -2320 0 feedthrough
rlabel pdiffusion 990 -2320 990 -2320 0 feedthrough
rlabel pdiffusion 997 -2320 997 -2320 0 cellNo=977
rlabel pdiffusion 1004 -2320 1004 -2320 0 feedthrough
rlabel pdiffusion 1011 -2320 1011 -2320 0 feedthrough
rlabel pdiffusion 1018 -2320 1018 -2320 0 feedthrough
rlabel pdiffusion 1025 -2320 1025 -2320 0 feedthrough
rlabel pdiffusion 1032 -2320 1032 -2320 0 feedthrough
rlabel pdiffusion 1039 -2320 1039 -2320 0 feedthrough
rlabel pdiffusion 1046 -2320 1046 -2320 0 feedthrough
rlabel pdiffusion 1053 -2320 1053 -2320 0 feedthrough
rlabel pdiffusion 1060 -2320 1060 -2320 0 feedthrough
rlabel pdiffusion 1067 -2320 1067 -2320 0 cellNo=530
rlabel pdiffusion 1074 -2320 1074 -2320 0 feedthrough
rlabel pdiffusion 1081 -2320 1081 -2320 0 feedthrough
rlabel pdiffusion 1088 -2320 1088 -2320 0 feedthrough
rlabel pdiffusion 1095 -2320 1095 -2320 0 feedthrough
rlabel pdiffusion 1102 -2320 1102 -2320 0 feedthrough
rlabel pdiffusion 1109 -2320 1109 -2320 0 feedthrough
rlabel pdiffusion 1116 -2320 1116 -2320 0 cellNo=351
rlabel pdiffusion 1123 -2320 1123 -2320 0 cellNo=600
rlabel pdiffusion 1130 -2320 1130 -2320 0 feedthrough
rlabel pdiffusion 1137 -2320 1137 -2320 0 feedthrough
rlabel pdiffusion 1144 -2320 1144 -2320 0 feedthrough
rlabel pdiffusion 1151 -2320 1151 -2320 0 feedthrough
rlabel pdiffusion 1158 -2320 1158 -2320 0 feedthrough
rlabel pdiffusion 1165 -2320 1165 -2320 0 feedthrough
rlabel pdiffusion 1172 -2320 1172 -2320 0 feedthrough
rlabel pdiffusion 1179 -2320 1179 -2320 0 feedthrough
rlabel pdiffusion 1186 -2320 1186 -2320 0 cellNo=404
rlabel pdiffusion 1193 -2320 1193 -2320 0 feedthrough
rlabel pdiffusion 1200 -2320 1200 -2320 0 feedthrough
rlabel pdiffusion 1207 -2320 1207 -2320 0 feedthrough
rlabel pdiffusion 1214 -2320 1214 -2320 0 feedthrough
rlabel pdiffusion 1221 -2320 1221 -2320 0 feedthrough
rlabel pdiffusion 1228 -2320 1228 -2320 0 feedthrough
rlabel pdiffusion 1235 -2320 1235 -2320 0 feedthrough
rlabel pdiffusion 1242 -2320 1242 -2320 0 feedthrough
rlabel pdiffusion 1249 -2320 1249 -2320 0 feedthrough
rlabel pdiffusion 1256 -2320 1256 -2320 0 feedthrough
rlabel pdiffusion 1263 -2320 1263 -2320 0 feedthrough
rlabel pdiffusion 1270 -2320 1270 -2320 0 feedthrough
rlabel pdiffusion 1277 -2320 1277 -2320 0 feedthrough
rlabel pdiffusion 1284 -2320 1284 -2320 0 feedthrough
rlabel pdiffusion 1291 -2320 1291 -2320 0 cellNo=28
rlabel pdiffusion 1298 -2320 1298 -2320 0 feedthrough
rlabel pdiffusion 1305 -2320 1305 -2320 0 cellNo=489
rlabel pdiffusion 1312 -2320 1312 -2320 0 feedthrough
rlabel pdiffusion 1319 -2320 1319 -2320 0 feedthrough
rlabel pdiffusion 1326 -2320 1326 -2320 0 feedthrough
rlabel pdiffusion 1333 -2320 1333 -2320 0 feedthrough
rlabel pdiffusion 1340 -2320 1340 -2320 0 feedthrough
rlabel pdiffusion 1347 -2320 1347 -2320 0 feedthrough
rlabel pdiffusion 1354 -2320 1354 -2320 0 feedthrough
rlabel pdiffusion 1361 -2320 1361 -2320 0 feedthrough
rlabel pdiffusion 1368 -2320 1368 -2320 0 cellNo=794
rlabel pdiffusion 1375 -2320 1375 -2320 0 feedthrough
rlabel pdiffusion 1382 -2320 1382 -2320 0 feedthrough
rlabel pdiffusion 1389 -2320 1389 -2320 0 feedthrough
rlabel pdiffusion 1396 -2320 1396 -2320 0 feedthrough
rlabel pdiffusion 1403 -2320 1403 -2320 0 feedthrough
rlabel pdiffusion 1410 -2320 1410 -2320 0 feedthrough
rlabel pdiffusion 1417 -2320 1417 -2320 0 feedthrough
rlabel pdiffusion 1424 -2320 1424 -2320 0 feedthrough
rlabel pdiffusion 1431 -2320 1431 -2320 0 feedthrough
rlabel pdiffusion 1438 -2320 1438 -2320 0 feedthrough
rlabel pdiffusion 1445 -2320 1445 -2320 0 feedthrough
rlabel pdiffusion 1452 -2320 1452 -2320 0 feedthrough
rlabel pdiffusion 1459 -2320 1459 -2320 0 feedthrough
rlabel pdiffusion 1466 -2320 1466 -2320 0 feedthrough
rlabel pdiffusion 1473 -2320 1473 -2320 0 feedthrough
rlabel pdiffusion 1480 -2320 1480 -2320 0 feedthrough
rlabel pdiffusion 1487 -2320 1487 -2320 0 feedthrough
rlabel pdiffusion 1494 -2320 1494 -2320 0 feedthrough
rlabel pdiffusion 1501 -2320 1501 -2320 0 feedthrough
rlabel pdiffusion 1508 -2320 1508 -2320 0 feedthrough
rlabel pdiffusion 1515 -2320 1515 -2320 0 feedthrough
rlabel pdiffusion 1522 -2320 1522 -2320 0 feedthrough
rlabel pdiffusion 1529 -2320 1529 -2320 0 feedthrough
rlabel pdiffusion 1536 -2320 1536 -2320 0 feedthrough
rlabel pdiffusion 1543 -2320 1543 -2320 0 feedthrough
rlabel pdiffusion 1550 -2320 1550 -2320 0 feedthrough
rlabel pdiffusion 1557 -2320 1557 -2320 0 feedthrough
rlabel pdiffusion 1564 -2320 1564 -2320 0 feedthrough
rlabel pdiffusion 1571 -2320 1571 -2320 0 feedthrough
rlabel pdiffusion 1578 -2320 1578 -2320 0 feedthrough
rlabel pdiffusion 1585 -2320 1585 -2320 0 feedthrough
rlabel pdiffusion 1592 -2320 1592 -2320 0 feedthrough
rlabel pdiffusion 1599 -2320 1599 -2320 0 feedthrough
rlabel pdiffusion 1606 -2320 1606 -2320 0 feedthrough
rlabel pdiffusion 1613 -2320 1613 -2320 0 feedthrough
rlabel pdiffusion 1620 -2320 1620 -2320 0 feedthrough
rlabel pdiffusion 1627 -2320 1627 -2320 0 feedthrough
rlabel pdiffusion 1634 -2320 1634 -2320 0 feedthrough
rlabel pdiffusion 1641 -2320 1641 -2320 0 feedthrough
rlabel pdiffusion 1648 -2320 1648 -2320 0 feedthrough
rlabel pdiffusion 1655 -2320 1655 -2320 0 feedthrough
rlabel pdiffusion 1662 -2320 1662 -2320 0 feedthrough
rlabel pdiffusion 1669 -2320 1669 -2320 0 feedthrough
rlabel pdiffusion 1676 -2320 1676 -2320 0 feedthrough
rlabel pdiffusion 1683 -2320 1683 -2320 0 feedthrough
rlabel pdiffusion 1690 -2320 1690 -2320 0 feedthrough
rlabel pdiffusion 1697 -2320 1697 -2320 0 feedthrough
rlabel pdiffusion 1704 -2320 1704 -2320 0 feedthrough
rlabel pdiffusion 1711 -2320 1711 -2320 0 cellNo=508
rlabel pdiffusion 1718 -2320 1718 -2320 0 feedthrough
rlabel pdiffusion 1725 -2320 1725 -2320 0 cellNo=282
rlabel pdiffusion 1732 -2320 1732 -2320 0 feedthrough
rlabel pdiffusion 1739 -2320 1739 -2320 0 feedthrough
rlabel pdiffusion 1746 -2320 1746 -2320 0 cellNo=645
rlabel pdiffusion 1753 -2320 1753 -2320 0 feedthrough
rlabel pdiffusion 1760 -2320 1760 -2320 0 feedthrough
rlabel pdiffusion 1767 -2320 1767 -2320 0 feedthrough
rlabel pdiffusion 1774 -2320 1774 -2320 0 feedthrough
rlabel pdiffusion 1781 -2320 1781 -2320 0 feedthrough
rlabel pdiffusion 1788 -2320 1788 -2320 0 feedthrough
rlabel pdiffusion 1795 -2320 1795 -2320 0 feedthrough
rlabel pdiffusion 1823 -2320 1823 -2320 0 feedthrough
rlabel pdiffusion 1830 -2320 1830 -2320 0 feedthrough
rlabel pdiffusion 3 -2445 3 -2445 0 cellNo=1078
rlabel pdiffusion 10 -2445 10 -2445 0 feedthrough
rlabel pdiffusion 17 -2445 17 -2445 0 feedthrough
rlabel pdiffusion 24 -2445 24 -2445 0 cellNo=1150
rlabel pdiffusion 31 -2445 31 -2445 0 feedthrough
rlabel pdiffusion 38 -2445 38 -2445 0 feedthrough
rlabel pdiffusion 45 -2445 45 -2445 0 feedthrough
rlabel pdiffusion 52 -2445 52 -2445 0 feedthrough
rlabel pdiffusion 59 -2445 59 -2445 0 feedthrough
rlabel pdiffusion 66 -2445 66 -2445 0 feedthrough
rlabel pdiffusion 73 -2445 73 -2445 0 feedthrough
rlabel pdiffusion 80 -2445 80 -2445 0 cellNo=691
rlabel pdiffusion 87 -2445 87 -2445 0 feedthrough
rlabel pdiffusion 94 -2445 94 -2445 0 cellNo=138
rlabel pdiffusion 101 -2445 101 -2445 0 feedthrough
rlabel pdiffusion 108 -2445 108 -2445 0 cellNo=98
rlabel pdiffusion 115 -2445 115 -2445 0 feedthrough
rlabel pdiffusion 122 -2445 122 -2445 0 feedthrough
rlabel pdiffusion 129 -2445 129 -2445 0 cellNo=337
rlabel pdiffusion 136 -2445 136 -2445 0 feedthrough
rlabel pdiffusion 143 -2445 143 -2445 0 feedthrough
rlabel pdiffusion 150 -2445 150 -2445 0 feedthrough
rlabel pdiffusion 157 -2445 157 -2445 0 feedthrough
rlabel pdiffusion 164 -2445 164 -2445 0 feedthrough
rlabel pdiffusion 171 -2445 171 -2445 0 feedthrough
rlabel pdiffusion 178 -2445 178 -2445 0 feedthrough
rlabel pdiffusion 185 -2445 185 -2445 0 feedthrough
rlabel pdiffusion 192 -2445 192 -2445 0 cellNo=424
rlabel pdiffusion 199 -2445 199 -2445 0 feedthrough
rlabel pdiffusion 206 -2445 206 -2445 0 feedthrough
rlabel pdiffusion 213 -2445 213 -2445 0 feedthrough
rlabel pdiffusion 220 -2445 220 -2445 0 feedthrough
rlabel pdiffusion 227 -2445 227 -2445 0 feedthrough
rlabel pdiffusion 234 -2445 234 -2445 0 feedthrough
rlabel pdiffusion 241 -2445 241 -2445 0 feedthrough
rlabel pdiffusion 248 -2445 248 -2445 0 feedthrough
rlabel pdiffusion 255 -2445 255 -2445 0 feedthrough
rlabel pdiffusion 262 -2445 262 -2445 0 feedthrough
rlabel pdiffusion 269 -2445 269 -2445 0 feedthrough
rlabel pdiffusion 276 -2445 276 -2445 0 feedthrough
rlabel pdiffusion 283 -2445 283 -2445 0 feedthrough
rlabel pdiffusion 290 -2445 290 -2445 0 feedthrough
rlabel pdiffusion 297 -2445 297 -2445 0 feedthrough
rlabel pdiffusion 304 -2445 304 -2445 0 feedthrough
rlabel pdiffusion 311 -2445 311 -2445 0 feedthrough
rlabel pdiffusion 318 -2445 318 -2445 0 feedthrough
rlabel pdiffusion 325 -2445 325 -2445 0 feedthrough
rlabel pdiffusion 332 -2445 332 -2445 0 feedthrough
rlabel pdiffusion 339 -2445 339 -2445 0 cellNo=420
rlabel pdiffusion 346 -2445 346 -2445 0 feedthrough
rlabel pdiffusion 353 -2445 353 -2445 0 feedthrough
rlabel pdiffusion 360 -2445 360 -2445 0 feedthrough
rlabel pdiffusion 367 -2445 367 -2445 0 feedthrough
rlabel pdiffusion 374 -2445 374 -2445 0 feedthrough
rlabel pdiffusion 381 -2445 381 -2445 0 feedthrough
rlabel pdiffusion 388 -2445 388 -2445 0 cellNo=94
rlabel pdiffusion 395 -2445 395 -2445 0 feedthrough
rlabel pdiffusion 402 -2445 402 -2445 0 cellNo=898
rlabel pdiffusion 409 -2445 409 -2445 0 feedthrough
rlabel pdiffusion 416 -2445 416 -2445 0 feedthrough
rlabel pdiffusion 423 -2445 423 -2445 0 feedthrough
rlabel pdiffusion 430 -2445 430 -2445 0 cellNo=587
rlabel pdiffusion 437 -2445 437 -2445 0 cellNo=304
rlabel pdiffusion 444 -2445 444 -2445 0 cellNo=664
rlabel pdiffusion 451 -2445 451 -2445 0 feedthrough
rlabel pdiffusion 458 -2445 458 -2445 0 cellNo=223
rlabel pdiffusion 465 -2445 465 -2445 0 feedthrough
rlabel pdiffusion 472 -2445 472 -2445 0 feedthrough
rlabel pdiffusion 479 -2445 479 -2445 0 feedthrough
rlabel pdiffusion 486 -2445 486 -2445 0 feedthrough
rlabel pdiffusion 493 -2445 493 -2445 0 feedthrough
rlabel pdiffusion 500 -2445 500 -2445 0 feedthrough
rlabel pdiffusion 507 -2445 507 -2445 0 feedthrough
rlabel pdiffusion 514 -2445 514 -2445 0 cellNo=491
rlabel pdiffusion 521 -2445 521 -2445 0 feedthrough
rlabel pdiffusion 528 -2445 528 -2445 0 cellNo=74
rlabel pdiffusion 535 -2445 535 -2445 0 feedthrough
rlabel pdiffusion 542 -2445 542 -2445 0 cellNo=485
rlabel pdiffusion 549 -2445 549 -2445 0 feedthrough
rlabel pdiffusion 556 -2445 556 -2445 0 feedthrough
rlabel pdiffusion 563 -2445 563 -2445 0 feedthrough
rlabel pdiffusion 570 -2445 570 -2445 0 feedthrough
rlabel pdiffusion 577 -2445 577 -2445 0 feedthrough
rlabel pdiffusion 584 -2445 584 -2445 0 feedthrough
rlabel pdiffusion 591 -2445 591 -2445 0 feedthrough
rlabel pdiffusion 598 -2445 598 -2445 0 cellNo=556
rlabel pdiffusion 605 -2445 605 -2445 0 feedthrough
rlabel pdiffusion 612 -2445 612 -2445 0 feedthrough
rlabel pdiffusion 619 -2445 619 -2445 0 feedthrough
rlabel pdiffusion 626 -2445 626 -2445 0 feedthrough
rlabel pdiffusion 633 -2445 633 -2445 0 feedthrough
rlabel pdiffusion 640 -2445 640 -2445 0 feedthrough
rlabel pdiffusion 647 -2445 647 -2445 0 feedthrough
rlabel pdiffusion 654 -2445 654 -2445 0 feedthrough
rlabel pdiffusion 661 -2445 661 -2445 0 feedthrough
rlabel pdiffusion 668 -2445 668 -2445 0 feedthrough
rlabel pdiffusion 675 -2445 675 -2445 0 cellNo=863
rlabel pdiffusion 682 -2445 682 -2445 0 feedthrough
rlabel pdiffusion 689 -2445 689 -2445 0 feedthrough
rlabel pdiffusion 696 -2445 696 -2445 0 cellNo=793
rlabel pdiffusion 703 -2445 703 -2445 0 feedthrough
rlabel pdiffusion 710 -2445 710 -2445 0 feedthrough
rlabel pdiffusion 717 -2445 717 -2445 0 cellNo=15
rlabel pdiffusion 724 -2445 724 -2445 0 feedthrough
rlabel pdiffusion 731 -2445 731 -2445 0 cellNo=273
rlabel pdiffusion 738 -2445 738 -2445 0 feedthrough
rlabel pdiffusion 745 -2445 745 -2445 0 feedthrough
rlabel pdiffusion 752 -2445 752 -2445 0 feedthrough
rlabel pdiffusion 759 -2445 759 -2445 0 feedthrough
rlabel pdiffusion 766 -2445 766 -2445 0 feedthrough
rlabel pdiffusion 773 -2445 773 -2445 0 feedthrough
rlabel pdiffusion 780 -2445 780 -2445 0 feedthrough
rlabel pdiffusion 787 -2445 787 -2445 0 cellNo=264
rlabel pdiffusion 794 -2445 794 -2445 0 feedthrough
rlabel pdiffusion 801 -2445 801 -2445 0 feedthrough
rlabel pdiffusion 808 -2445 808 -2445 0 feedthrough
rlabel pdiffusion 815 -2445 815 -2445 0 feedthrough
rlabel pdiffusion 822 -2445 822 -2445 0 feedthrough
rlabel pdiffusion 829 -2445 829 -2445 0 cellNo=371
rlabel pdiffusion 836 -2445 836 -2445 0 feedthrough
rlabel pdiffusion 843 -2445 843 -2445 0 feedthrough
rlabel pdiffusion 850 -2445 850 -2445 0 feedthrough
rlabel pdiffusion 857 -2445 857 -2445 0 feedthrough
rlabel pdiffusion 864 -2445 864 -2445 0 feedthrough
rlabel pdiffusion 871 -2445 871 -2445 0 feedthrough
rlabel pdiffusion 878 -2445 878 -2445 0 feedthrough
rlabel pdiffusion 885 -2445 885 -2445 0 cellNo=128
rlabel pdiffusion 892 -2445 892 -2445 0 feedthrough
rlabel pdiffusion 899 -2445 899 -2445 0 feedthrough
rlabel pdiffusion 906 -2445 906 -2445 0 feedthrough
rlabel pdiffusion 913 -2445 913 -2445 0 feedthrough
rlabel pdiffusion 920 -2445 920 -2445 0 feedthrough
rlabel pdiffusion 927 -2445 927 -2445 0 feedthrough
rlabel pdiffusion 934 -2445 934 -2445 0 feedthrough
rlabel pdiffusion 941 -2445 941 -2445 0 feedthrough
rlabel pdiffusion 948 -2445 948 -2445 0 feedthrough
rlabel pdiffusion 955 -2445 955 -2445 0 feedthrough
rlabel pdiffusion 962 -2445 962 -2445 0 feedthrough
rlabel pdiffusion 969 -2445 969 -2445 0 feedthrough
rlabel pdiffusion 976 -2445 976 -2445 0 feedthrough
rlabel pdiffusion 983 -2445 983 -2445 0 feedthrough
rlabel pdiffusion 990 -2445 990 -2445 0 feedthrough
rlabel pdiffusion 997 -2445 997 -2445 0 feedthrough
rlabel pdiffusion 1004 -2445 1004 -2445 0 feedthrough
rlabel pdiffusion 1011 -2445 1011 -2445 0 feedthrough
rlabel pdiffusion 1018 -2445 1018 -2445 0 cellNo=570
rlabel pdiffusion 1025 -2445 1025 -2445 0 feedthrough
rlabel pdiffusion 1032 -2445 1032 -2445 0 feedthrough
rlabel pdiffusion 1039 -2445 1039 -2445 0 feedthrough
rlabel pdiffusion 1046 -2445 1046 -2445 0 feedthrough
rlabel pdiffusion 1053 -2445 1053 -2445 0 cellNo=237
rlabel pdiffusion 1060 -2445 1060 -2445 0 feedthrough
rlabel pdiffusion 1067 -2445 1067 -2445 0 feedthrough
rlabel pdiffusion 1074 -2445 1074 -2445 0 feedthrough
rlabel pdiffusion 1081 -2445 1081 -2445 0 cellNo=838
rlabel pdiffusion 1088 -2445 1088 -2445 0 feedthrough
rlabel pdiffusion 1095 -2445 1095 -2445 0 feedthrough
rlabel pdiffusion 1102 -2445 1102 -2445 0 feedthrough
rlabel pdiffusion 1109 -2445 1109 -2445 0 feedthrough
rlabel pdiffusion 1116 -2445 1116 -2445 0 feedthrough
rlabel pdiffusion 1123 -2445 1123 -2445 0 feedthrough
rlabel pdiffusion 1130 -2445 1130 -2445 0 feedthrough
rlabel pdiffusion 1137 -2445 1137 -2445 0 feedthrough
rlabel pdiffusion 1144 -2445 1144 -2445 0 feedthrough
rlabel pdiffusion 1151 -2445 1151 -2445 0 feedthrough
rlabel pdiffusion 1158 -2445 1158 -2445 0 feedthrough
rlabel pdiffusion 1165 -2445 1165 -2445 0 cellNo=55
rlabel pdiffusion 1172 -2445 1172 -2445 0 feedthrough
rlabel pdiffusion 1179 -2445 1179 -2445 0 feedthrough
rlabel pdiffusion 1186 -2445 1186 -2445 0 feedthrough
rlabel pdiffusion 1193 -2445 1193 -2445 0 feedthrough
rlabel pdiffusion 1200 -2445 1200 -2445 0 feedthrough
rlabel pdiffusion 1207 -2445 1207 -2445 0 feedthrough
rlabel pdiffusion 1214 -2445 1214 -2445 0 cellNo=910
rlabel pdiffusion 1221 -2445 1221 -2445 0 feedthrough
rlabel pdiffusion 1228 -2445 1228 -2445 0 feedthrough
rlabel pdiffusion 1235 -2445 1235 -2445 0 feedthrough
rlabel pdiffusion 1242 -2445 1242 -2445 0 feedthrough
rlabel pdiffusion 1249 -2445 1249 -2445 0 feedthrough
rlabel pdiffusion 1256 -2445 1256 -2445 0 feedthrough
rlabel pdiffusion 1263 -2445 1263 -2445 0 feedthrough
rlabel pdiffusion 1270 -2445 1270 -2445 0 feedthrough
rlabel pdiffusion 1277 -2445 1277 -2445 0 feedthrough
rlabel pdiffusion 1284 -2445 1284 -2445 0 feedthrough
rlabel pdiffusion 1291 -2445 1291 -2445 0 feedthrough
rlabel pdiffusion 1298 -2445 1298 -2445 0 feedthrough
rlabel pdiffusion 1305 -2445 1305 -2445 0 feedthrough
rlabel pdiffusion 1312 -2445 1312 -2445 0 feedthrough
rlabel pdiffusion 1319 -2445 1319 -2445 0 cellNo=573
rlabel pdiffusion 1326 -2445 1326 -2445 0 feedthrough
rlabel pdiffusion 1333 -2445 1333 -2445 0 feedthrough
rlabel pdiffusion 1340 -2445 1340 -2445 0 cellNo=682
rlabel pdiffusion 1347 -2445 1347 -2445 0 feedthrough
rlabel pdiffusion 1354 -2445 1354 -2445 0 feedthrough
rlabel pdiffusion 1361 -2445 1361 -2445 0 feedthrough
rlabel pdiffusion 1368 -2445 1368 -2445 0 feedthrough
rlabel pdiffusion 1375 -2445 1375 -2445 0 feedthrough
rlabel pdiffusion 1382 -2445 1382 -2445 0 feedthrough
rlabel pdiffusion 1389 -2445 1389 -2445 0 cellNo=575
rlabel pdiffusion 1396 -2445 1396 -2445 0 feedthrough
rlabel pdiffusion 1403 -2445 1403 -2445 0 feedthrough
rlabel pdiffusion 1410 -2445 1410 -2445 0 feedthrough
rlabel pdiffusion 1417 -2445 1417 -2445 0 feedthrough
rlabel pdiffusion 1424 -2445 1424 -2445 0 feedthrough
rlabel pdiffusion 1431 -2445 1431 -2445 0 feedthrough
rlabel pdiffusion 1438 -2445 1438 -2445 0 feedthrough
rlabel pdiffusion 1445 -2445 1445 -2445 0 feedthrough
rlabel pdiffusion 1452 -2445 1452 -2445 0 feedthrough
rlabel pdiffusion 1459 -2445 1459 -2445 0 feedthrough
rlabel pdiffusion 1466 -2445 1466 -2445 0 feedthrough
rlabel pdiffusion 1473 -2445 1473 -2445 0 feedthrough
rlabel pdiffusion 1480 -2445 1480 -2445 0 feedthrough
rlabel pdiffusion 1487 -2445 1487 -2445 0 feedthrough
rlabel pdiffusion 1494 -2445 1494 -2445 0 feedthrough
rlabel pdiffusion 1501 -2445 1501 -2445 0 feedthrough
rlabel pdiffusion 1508 -2445 1508 -2445 0 feedthrough
rlabel pdiffusion 1515 -2445 1515 -2445 0 feedthrough
rlabel pdiffusion 1522 -2445 1522 -2445 0 feedthrough
rlabel pdiffusion 1529 -2445 1529 -2445 0 feedthrough
rlabel pdiffusion 1536 -2445 1536 -2445 0 feedthrough
rlabel pdiffusion 1543 -2445 1543 -2445 0 feedthrough
rlabel pdiffusion 1550 -2445 1550 -2445 0 feedthrough
rlabel pdiffusion 1557 -2445 1557 -2445 0 feedthrough
rlabel pdiffusion 1564 -2445 1564 -2445 0 feedthrough
rlabel pdiffusion 1571 -2445 1571 -2445 0 feedthrough
rlabel pdiffusion 1578 -2445 1578 -2445 0 feedthrough
rlabel pdiffusion 1585 -2445 1585 -2445 0 feedthrough
rlabel pdiffusion 1592 -2445 1592 -2445 0 feedthrough
rlabel pdiffusion 1599 -2445 1599 -2445 0 feedthrough
rlabel pdiffusion 1606 -2445 1606 -2445 0 feedthrough
rlabel pdiffusion 1613 -2445 1613 -2445 0 feedthrough
rlabel pdiffusion 1620 -2445 1620 -2445 0 feedthrough
rlabel pdiffusion 1627 -2445 1627 -2445 0 feedthrough
rlabel pdiffusion 1634 -2445 1634 -2445 0 feedthrough
rlabel pdiffusion 1641 -2445 1641 -2445 0 feedthrough
rlabel pdiffusion 1648 -2445 1648 -2445 0 feedthrough
rlabel pdiffusion 1655 -2445 1655 -2445 0 feedthrough
rlabel pdiffusion 1662 -2445 1662 -2445 0 feedthrough
rlabel pdiffusion 1669 -2445 1669 -2445 0 feedthrough
rlabel pdiffusion 1676 -2445 1676 -2445 0 feedthrough
rlabel pdiffusion 1683 -2445 1683 -2445 0 feedthrough
rlabel pdiffusion 1690 -2445 1690 -2445 0 feedthrough
rlabel pdiffusion 1697 -2445 1697 -2445 0 feedthrough
rlabel pdiffusion 1704 -2445 1704 -2445 0 feedthrough
rlabel pdiffusion 1711 -2445 1711 -2445 0 feedthrough
rlabel pdiffusion 1718 -2445 1718 -2445 0 feedthrough
rlabel pdiffusion 1725 -2445 1725 -2445 0 feedthrough
rlabel pdiffusion 1732 -2445 1732 -2445 0 feedthrough
rlabel pdiffusion 1739 -2445 1739 -2445 0 feedthrough
rlabel pdiffusion 1746 -2445 1746 -2445 0 feedthrough
rlabel pdiffusion 1753 -2445 1753 -2445 0 cellNo=564
rlabel pdiffusion 1760 -2445 1760 -2445 0 feedthrough
rlabel pdiffusion 1767 -2445 1767 -2445 0 feedthrough
rlabel pdiffusion 1774 -2445 1774 -2445 0 feedthrough
rlabel pdiffusion 1781 -2445 1781 -2445 0 feedthrough
rlabel pdiffusion 1788 -2445 1788 -2445 0 feedthrough
rlabel pdiffusion 1795 -2445 1795 -2445 0 cellNo=105
rlabel pdiffusion 1802 -2445 1802 -2445 0 feedthrough
rlabel pdiffusion 1809 -2445 1809 -2445 0 feedthrough
rlabel pdiffusion 3 -2580 3 -2580 0 cellNo=1043
rlabel pdiffusion 10 -2580 10 -2580 0 cellNo=1179
rlabel pdiffusion 17 -2580 17 -2580 0 feedthrough
rlabel pdiffusion 24 -2580 24 -2580 0 feedthrough
rlabel pdiffusion 31 -2580 31 -2580 0 feedthrough
rlabel pdiffusion 38 -2580 38 -2580 0 feedthrough
rlabel pdiffusion 45 -2580 45 -2580 0 feedthrough
rlabel pdiffusion 52 -2580 52 -2580 0 feedthrough
rlabel pdiffusion 59 -2580 59 -2580 0 feedthrough
rlabel pdiffusion 66 -2580 66 -2580 0 feedthrough
rlabel pdiffusion 73 -2580 73 -2580 0 feedthrough
rlabel pdiffusion 80 -2580 80 -2580 0 feedthrough
rlabel pdiffusion 87 -2580 87 -2580 0 feedthrough
rlabel pdiffusion 94 -2580 94 -2580 0 feedthrough
rlabel pdiffusion 101 -2580 101 -2580 0 cellNo=869
rlabel pdiffusion 108 -2580 108 -2580 0 cellNo=930
rlabel pdiffusion 115 -2580 115 -2580 0 feedthrough
rlabel pdiffusion 122 -2580 122 -2580 0 feedthrough
rlabel pdiffusion 129 -2580 129 -2580 0 feedthrough
rlabel pdiffusion 136 -2580 136 -2580 0 feedthrough
rlabel pdiffusion 143 -2580 143 -2580 0 feedthrough
rlabel pdiffusion 150 -2580 150 -2580 0 cellNo=308
rlabel pdiffusion 157 -2580 157 -2580 0 cellNo=384
rlabel pdiffusion 164 -2580 164 -2580 0 feedthrough
rlabel pdiffusion 171 -2580 171 -2580 0 cellNo=187
rlabel pdiffusion 178 -2580 178 -2580 0 feedthrough
rlabel pdiffusion 185 -2580 185 -2580 0 feedthrough
rlabel pdiffusion 192 -2580 192 -2580 0 feedthrough
rlabel pdiffusion 199 -2580 199 -2580 0 feedthrough
rlabel pdiffusion 206 -2580 206 -2580 0 feedthrough
rlabel pdiffusion 213 -2580 213 -2580 0 feedthrough
rlabel pdiffusion 220 -2580 220 -2580 0 feedthrough
rlabel pdiffusion 227 -2580 227 -2580 0 feedthrough
rlabel pdiffusion 234 -2580 234 -2580 0 feedthrough
rlabel pdiffusion 241 -2580 241 -2580 0 cellNo=756
rlabel pdiffusion 248 -2580 248 -2580 0 feedthrough
rlabel pdiffusion 255 -2580 255 -2580 0 feedthrough
rlabel pdiffusion 262 -2580 262 -2580 0 feedthrough
rlabel pdiffusion 269 -2580 269 -2580 0 feedthrough
rlabel pdiffusion 276 -2580 276 -2580 0 feedthrough
rlabel pdiffusion 283 -2580 283 -2580 0 feedthrough
rlabel pdiffusion 290 -2580 290 -2580 0 feedthrough
rlabel pdiffusion 297 -2580 297 -2580 0 feedthrough
rlabel pdiffusion 304 -2580 304 -2580 0 feedthrough
rlabel pdiffusion 311 -2580 311 -2580 0 feedthrough
rlabel pdiffusion 318 -2580 318 -2580 0 feedthrough
rlabel pdiffusion 325 -2580 325 -2580 0 feedthrough
rlabel pdiffusion 332 -2580 332 -2580 0 feedthrough
rlabel pdiffusion 339 -2580 339 -2580 0 feedthrough
rlabel pdiffusion 346 -2580 346 -2580 0 feedthrough
rlabel pdiffusion 353 -2580 353 -2580 0 feedthrough
rlabel pdiffusion 360 -2580 360 -2580 0 feedthrough
rlabel pdiffusion 367 -2580 367 -2580 0 feedthrough
rlabel pdiffusion 374 -2580 374 -2580 0 feedthrough
rlabel pdiffusion 381 -2580 381 -2580 0 feedthrough
rlabel pdiffusion 388 -2580 388 -2580 0 feedthrough
rlabel pdiffusion 395 -2580 395 -2580 0 feedthrough
rlabel pdiffusion 402 -2580 402 -2580 0 feedthrough
rlabel pdiffusion 409 -2580 409 -2580 0 feedthrough
rlabel pdiffusion 416 -2580 416 -2580 0 feedthrough
rlabel pdiffusion 423 -2580 423 -2580 0 feedthrough
rlabel pdiffusion 430 -2580 430 -2580 0 feedthrough
rlabel pdiffusion 437 -2580 437 -2580 0 feedthrough
rlabel pdiffusion 444 -2580 444 -2580 0 feedthrough
rlabel pdiffusion 451 -2580 451 -2580 0 cellNo=839
rlabel pdiffusion 458 -2580 458 -2580 0 feedthrough
rlabel pdiffusion 465 -2580 465 -2580 0 feedthrough
rlabel pdiffusion 472 -2580 472 -2580 0 feedthrough
rlabel pdiffusion 479 -2580 479 -2580 0 feedthrough
rlabel pdiffusion 486 -2580 486 -2580 0 feedthrough
rlabel pdiffusion 493 -2580 493 -2580 0 feedthrough
rlabel pdiffusion 500 -2580 500 -2580 0 feedthrough
rlabel pdiffusion 507 -2580 507 -2580 0 feedthrough
rlabel pdiffusion 514 -2580 514 -2580 0 feedthrough
rlabel pdiffusion 521 -2580 521 -2580 0 feedthrough
rlabel pdiffusion 528 -2580 528 -2580 0 feedthrough
rlabel pdiffusion 535 -2580 535 -2580 0 feedthrough
rlabel pdiffusion 542 -2580 542 -2580 0 feedthrough
rlabel pdiffusion 549 -2580 549 -2580 0 feedthrough
rlabel pdiffusion 556 -2580 556 -2580 0 cellNo=961
rlabel pdiffusion 563 -2580 563 -2580 0 feedthrough
rlabel pdiffusion 570 -2580 570 -2580 0 feedthrough
rlabel pdiffusion 577 -2580 577 -2580 0 feedthrough
rlabel pdiffusion 584 -2580 584 -2580 0 feedthrough
rlabel pdiffusion 591 -2580 591 -2580 0 feedthrough
rlabel pdiffusion 598 -2580 598 -2580 0 cellNo=772
rlabel pdiffusion 605 -2580 605 -2580 0 feedthrough
rlabel pdiffusion 612 -2580 612 -2580 0 feedthrough
rlabel pdiffusion 619 -2580 619 -2580 0 feedthrough
rlabel pdiffusion 626 -2580 626 -2580 0 cellNo=67
rlabel pdiffusion 633 -2580 633 -2580 0 feedthrough
rlabel pdiffusion 640 -2580 640 -2580 0 cellNo=626
rlabel pdiffusion 647 -2580 647 -2580 0 feedthrough
rlabel pdiffusion 654 -2580 654 -2580 0 feedthrough
rlabel pdiffusion 661 -2580 661 -2580 0 feedthrough
rlabel pdiffusion 668 -2580 668 -2580 0 cellNo=578
rlabel pdiffusion 675 -2580 675 -2580 0 feedthrough
rlabel pdiffusion 682 -2580 682 -2580 0 feedthrough
rlabel pdiffusion 689 -2580 689 -2580 0 feedthrough
rlabel pdiffusion 696 -2580 696 -2580 0 feedthrough
rlabel pdiffusion 703 -2580 703 -2580 0 feedthrough
rlabel pdiffusion 710 -2580 710 -2580 0 cellNo=217
rlabel pdiffusion 717 -2580 717 -2580 0 feedthrough
rlabel pdiffusion 724 -2580 724 -2580 0 cellNo=610
rlabel pdiffusion 731 -2580 731 -2580 0 feedthrough
rlabel pdiffusion 738 -2580 738 -2580 0 cellNo=171
rlabel pdiffusion 745 -2580 745 -2580 0 feedthrough
rlabel pdiffusion 752 -2580 752 -2580 0 feedthrough
rlabel pdiffusion 759 -2580 759 -2580 0 feedthrough
rlabel pdiffusion 766 -2580 766 -2580 0 feedthrough
rlabel pdiffusion 773 -2580 773 -2580 0 feedthrough
rlabel pdiffusion 780 -2580 780 -2580 0 feedthrough
rlabel pdiffusion 787 -2580 787 -2580 0 feedthrough
rlabel pdiffusion 794 -2580 794 -2580 0 feedthrough
rlabel pdiffusion 801 -2580 801 -2580 0 feedthrough
rlabel pdiffusion 808 -2580 808 -2580 0 feedthrough
rlabel pdiffusion 815 -2580 815 -2580 0 feedthrough
rlabel pdiffusion 822 -2580 822 -2580 0 feedthrough
rlabel pdiffusion 829 -2580 829 -2580 0 feedthrough
rlabel pdiffusion 836 -2580 836 -2580 0 feedthrough
rlabel pdiffusion 843 -2580 843 -2580 0 feedthrough
rlabel pdiffusion 850 -2580 850 -2580 0 cellNo=471
rlabel pdiffusion 857 -2580 857 -2580 0 feedthrough
rlabel pdiffusion 864 -2580 864 -2580 0 feedthrough
rlabel pdiffusion 871 -2580 871 -2580 0 feedthrough
rlabel pdiffusion 878 -2580 878 -2580 0 feedthrough
rlabel pdiffusion 885 -2580 885 -2580 0 feedthrough
rlabel pdiffusion 892 -2580 892 -2580 0 feedthrough
rlabel pdiffusion 899 -2580 899 -2580 0 feedthrough
rlabel pdiffusion 906 -2580 906 -2580 0 feedthrough
rlabel pdiffusion 913 -2580 913 -2580 0 feedthrough
rlabel pdiffusion 920 -2580 920 -2580 0 feedthrough
rlabel pdiffusion 927 -2580 927 -2580 0 feedthrough
rlabel pdiffusion 934 -2580 934 -2580 0 feedthrough
rlabel pdiffusion 941 -2580 941 -2580 0 feedthrough
rlabel pdiffusion 948 -2580 948 -2580 0 cellNo=673
rlabel pdiffusion 955 -2580 955 -2580 0 feedthrough
rlabel pdiffusion 962 -2580 962 -2580 0 feedthrough
rlabel pdiffusion 969 -2580 969 -2580 0 cellNo=955
rlabel pdiffusion 976 -2580 976 -2580 0 feedthrough
rlabel pdiffusion 983 -2580 983 -2580 0 feedthrough
rlabel pdiffusion 990 -2580 990 -2580 0 cellNo=813
rlabel pdiffusion 997 -2580 997 -2580 0 feedthrough
rlabel pdiffusion 1004 -2580 1004 -2580 0 feedthrough
rlabel pdiffusion 1011 -2580 1011 -2580 0 feedthrough
rlabel pdiffusion 1018 -2580 1018 -2580 0 cellNo=202
rlabel pdiffusion 1025 -2580 1025 -2580 0 feedthrough
rlabel pdiffusion 1032 -2580 1032 -2580 0 feedthrough
rlabel pdiffusion 1039 -2580 1039 -2580 0 feedthrough
rlabel pdiffusion 1046 -2580 1046 -2580 0 cellNo=780
rlabel pdiffusion 1053 -2580 1053 -2580 0 cellNo=745
rlabel pdiffusion 1060 -2580 1060 -2580 0 feedthrough
rlabel pdiffusion 1067 -2580 1067 -2580 0 feedthrough
rlabel pdiffusion 1074 -2580 1074 -2580 0 cellNo=877
rlabel pdiffusion 1081 -2580 1081 -2580 0 feedthrough
rlabel pdiffusion 1088 -2580 1088 -2580 0 feedthrough
rlabel pdiffusion 1095 -2580 1095 -2580 0 feedthrough
rlabel pdiffusion 1102 -2580 1102 -2580 0 feedthrough
rlabel pdiffusion 1109 -2580 1109 -2580 0 feedthrough
rlabel pdiffusion 1116 -2580 1116 -2580 0 cellNo=841
rlabel pdiffusion 1123 -2580 1123 -2580 0 feedthrough
rlabel pdiffusion 1130 -2580 1130 -2580 0 cellNo=663
rlabel pdiffusion 1137 -2580 1137 -2580 0 cellNo=467
rlabel pdiffusion 1144 -2580 1144 -2580 0 feedthrough
rlabel pdiffusion 1151 -2580 1151 -2580 0 feedthrough
rlabel pdiffusion 1158 -2580 1158 -2580 0 cellNo=761
rlabel pdiffusion 1165 -2580 1165 -2580 0 feedthrough
rlabel pdiffusion 1172 -2580 1172 -2580 0 cellNo=536
rlabel pdiffusion 1179 -2580 1179 -2580 0 feedthrough
rlabel pdiffusion 1186 -2580 1186 -2580 0 feedthrough
rlabel pdiffusion 1193 -2580 1193 -2580 0 cellNo=269
rlabel pdiffusion 1200 -2580 1200 -2580 0 feedthrough
rlabel pdiffusion 1207 -2580 1207 -2580 0 feedthrough
rlabel pdiffusion 1214 -2580 1214 -2580 0 feedthrough
rlabel pdiffusion 1221 -2580 1221 -2580 0 feedthrough
rlabel pdiffusion 1228 -2580 1228 -2580 0 feedthrough
rlabel pdiffusion 1235 -2580 1235 -2580 0 feedthrough
rlabel pdiffusion 1242 -2580 1242 -2580 0 feedthrough
rlabel pdiffusion 1249 -2580 1249 -2580 0 feedthrough
rlabel pdiffusion 1256 -2580 1256 -2580 0 feedthrough
rlabel pdiffusion 1263 -2580 1263 -2580 0 feedthrough
rlabel pdiffusion 1270 -2580 1270 -2580 0 feedthrough
rlabel pdiffusion 1277 -2580 1277 -2580 0 feedthrough
rlabel pdiffusion 1284 -2580 1284 -2580 0 feedthrough
rlabel pdiffusion 1291 -2580 1291 -2580 0 feedthrough
rlabel pdiffusion 1298 -2580 1298 -2580 0 feedthrough
rlabel pdiffusion 1305 -2580 1305 -2580 0 feedthrough
rlabel pdiffusion 1312 -2580 1312 -2580 0 feedthrough
rlabel pdiffusion 1319 -2580 1319 -2580 0 feedthrough
rlabel pdiffusion 1326 -2580 1326 -2580 0 feedthrough
rlabel pdiffusion 1333 -2580 1333 -2580 0 feedthrough
rlabel pdiffusion 1340 -2580 1340 -2580 0 feedthrough
rlabel pdiffusion 1347 -2580 1347 -2580 0 feedthrough
rlabel pdiffusion 1354 -2580 1354 -2580 0 feedthrough
rlabel pdiffusion 1361 -2580 1361 -2580 0 feedthrough
rlabel pdiffusion 1368 -2580 1368 -2580 0 feedthrough
rlabel pdiffusion 1375 -2580 1375 -2580 0 feedthrough
rlabel pdiffusion 1382 -2580 1382 -2580 0 feedthrough
rlabel pdiffusion 1389 -2580 1389 -2580 0 feedthrough
rlabel pdiffusion 1396 -2580 1396 -2580 0 feedthrough
rlabel pdiffusion 1403 -2580 1403 -2580 0 feedthrough
rlabel pdiffusion 1410 -2580 1410 -2580 0 feedthrough
rlabel pdiffusion 1417 -2580 1417 -2580 0 feedthrough
rlabel pdiffusion 1424 -2580 1424 -2580 0 feedthrough
rlabel pdiffusion 1431 -2580 1431 -2580 0 feedthrough
rlabel pdiffusion 1438 -2580 1438 -2580 0 feedthrough
rlabel pdiffusion 1445 -2580 1445 -2580 0 feedthrough
rlabel pdiffusion 1452 -2580 1452 -2580 0 feedthrough
rlabel pdiffusion 1459 -2580 1459 -2580 0 feedthrough
rlabel pdiffusion 1466 -2580 1466 -2580 0 feedthrough
rlabel pdiffusion 1473 -2580 1473 -2580 0 feedthrough
rlabel pdiffusion 1480 -2580 1480 -2580 0 feedthrough
rlabel pdiffusion 1487 -2580 1487 -2580 0 feedthrough
rlabel pdiffusion 1494 -2580 1494 -2580 0 feedthrough
rlabel pdiffusion 1501 -2580 1501 -2580 0 feedthrough
rlabel pdiffusion 1508 -2580 1508 -2580 0 cellNo=938
rlabel pdiffusion 1515 -2580 1515 -2580 0 feedthrough
rlabel pdiffusion 1522 -2580 1522 -2580 0 feedthrough
rlabel pdiffusion 1529 -2580 1529 -2580 0 feedthrough
rlabel pdiffusion 1536 -2580 1536 -2580 0 feedthrough
rlabel pdiffusion 1543 -2580 1543 -2580 0 feedthrough
rlabel pdiffusion 1550 -2580 1550 -2580 0 feedthrough
rlabel pdiffusion 1557 -2580 1557 -2580 0 feedthrough
rlabel pdiffusion 1564 -2580 1564 -2580 0 feedthrough
rlabel pdiffusion 1571 -2580 1571 -2580 0 feedthrough
rlabel pdiffusion 1578 -2580 1578 -2580 0 feedthrough
rlabel pdiffusion 1585 -2580 1585 -2580 0 feedthrough
rlabel pdiffusion 1592 -2580 1592 -2580 0 feedthrough
rlabel pdiffusion 1599 -2580 1599 -2580 0 feedthrough
rlabel pdiffusion 1606 -2580 1606 -2580 0 feedthrough
rlabel pdiffusion 1613 -2580 1613 -2580 0 feedthrough
rlabel pdiffusion 1620 -2580 1620 -2580 0 feedthrough
rlabel pdiffusion 1627 -2580 1627 -2580 0 feedthrough
rlabel pdiffusion 1634 -2580 1634 -2580 0 feedthrough
rlabel pdiffusion 1641 -2580 1641 -2580 0 feedthrough
rlabel pdiffusion 1648 -2580 1648 -2580 0 feedthrough
rlabel pdiffusion 1655 -2580 1655 -2580 0 feedthrough
rlabel pdiffusion 1662 -2580 1662 -2580 0 feedthrough
rlabel pdiffusion 1669 -2580 1669 -2580 0 feedthrough
rlabel pdiffusion 1676 -2580 1676 -2580 0 feedthrough
rlabel pdiffusion 1683 -2580 1683 -2580 0 feedthrough
rlabel pdiffusion 1690 -2580 1690 -2580 0 feedthrough
rlabel pdiffusion 1697 -2580 1697 -2580 0 cellNo=970
rlabel pdiffusion 1704 -2580 1704 -2580 0 feedthrough
rlabel pdiffusion 1711 -2580 1711 -2580 0 feedthrough
rlabel pdiffusion 1718 -2580 1718 -2580 0 feedthrough
rlabel pdiffusion 1725 -2580 1725 -2580 0 feedthrough
rlabel pdiffusion 1732 -2580 1732 -2580 0 feedthrough
rlabel pdiffusion 1739 -2580 1739 -2580 0 cellNo=911
rlabel pdiffusion 1746 -2580 1746 -2580 0 feedthrough
rlabel pdiffusion 1753 -2580 1753 -2580 0 feedthrough
rlabel pdiffusion 1760 -2580 1760 -2580 0 feedthrough
rlabel pdiffusion 1767 -2580 1767 -2580 0 feedthrough
rlabel pdiffusion 1774 -2580 1774 -2580 0 feedthrough
rlabel pdiffusion 1781 -2580 1781 -2580 0 feedthrough
rlabel pdiffusion 1788 -2580 1788 -2580 0 feedthrough
rlabel pdiffusion 1795 -2580 1795 -2580 0 cellNo=425
rlabel pdiffusion 1802 -2580 1802 -2580 0 feedthrough
rlabel pdiffusion 1809 -2580 1809 -2580 0 feedthrough
rlabel pdiffusion 1816 -2580 1816 -2580 0 feedthrough
rlabel pdiffusion 3 -2713 3 -2713 0 cellNo=1118
rlabel pdiffusion 10 -2713 10 -2713 0 feedthrough
rlabel pdiffusion 17 -2713 17 -2713 0 cellNo=324
rlabel pdiffusion 24 -2713 24 -2713 0 cellNo=1144
rlabel pdiffusion 31 -2713 31 -2713 0 feedthrough
rlabel pdiffusion 38 -2713 38 -2713 0 feedthrough
rlabel pdiffusion 45 -2713 45 -2713 0 feedthrough
rlabel pdiffusion 52 -2713 52 -2713 0 feedthrough
rlabel pdiffusion 59 -2713 59 -2713 0 cellNo=973
rlabel pdiffusion 66 -2713 66 -2713 0 cellNo=912
rlabel pdiffusion 73 -2713 73 -2713 0 feedthrough
rlabel pdiffusion 80 -2713 80 -2713 0 feedthrough
rlabel pdiffusion 87 -2713 87 -2713 0 feedthrough
rlabel pdiffusion 94 -2713 94 -2713 0 feedthrough
rlabel pdiffusion 101 -2713 101 -2713 0 feedthrough
rlabel pdiffusion 108 -2713 108 -2713 0 feedthrough
rlabel pdiffusion 115 -2713 115 -2713 0 feedthrough
rlabel pdiffusion 122 -2713 122 -2713 0 feedthrough
rlabel pdiffusion 129 -2713 129 -2713 0 feedthrough
rlabel pdiffusion 136 -2713 136 -2713 0 feedthrough
rlabel pdiffusion 143 -2713 143 -2713 0 feedthrough
rlabel pdiffusion 150 -2713 150 -2713 0 feedthrough
rlabel pdiffusion 157 -2713 157 -2713 0 feedthrough
rlabel pdiffusion 164 -2713 164 -2713 0 feedthrough
rlabel pdiffusion 171 -2713 171 -2713 0 feedthrough
rlabel pdiffusion 178 -2713 178 -2713 0 feedthrough
rlabel pdiffusion 185 -2713 185 -2713 0 feedthrough
rlabel pdiffusion 192 -2713 192 -2713 0 feedthrough
rlabel pdiffusion 199 -2713 199 -2713 0 cellNo=470
rlabel pdiffusion 206 -2713 206 -2713 0 cellNo=86
rlabel pdiffusion 213 -2713 213 -2713 0 feedthrough
rlabel pdiffusion 220 -2713 220 -2713 0 feedthrough
rlabel pdiffusion 227 -2713 227 -2713 0 feedthrough
rlabel pdiffusion 234 -2713 234 -2713 0 feedthrough
rlabel pdiffusion 241 -2713 241 -2713 0 feedthrough
rlabel pdiffusion 248 -2713 248 -2713 0 feedthrough
rlabel pdiffusion 255 -2713 255 -2713 0 feedthrough
rlabel pdiffusion 262 -2713 262 -2713 0 feedthrough
rlabel pdiffusion 269 -2713 269 -2713 0 feedthrough
rlabel pdiffusion 276 -2713 276 -2713 0 feedthrough
rlabel pdiffusion 283 -2713 283 -2713 0 feedthrough
rlabel pdiffusion 290 -2713 290 -2713 0 cellNo=925
rlabel pdiffusion 297 -2713 297 -2713 0 feedthrough
rlabel pdiffusion 304 -2713 304 -2713 0 feedthrough
rlabel pdiffusion 311 -2713 311 -2713 0 feedthrough
rlabel pdiffusion 318 -2713 318 -2713 0 feedthrough
rlabel pdiffusion 325 -2713 325 -2713 0 feedthrough
rlabel pdiffusion 332 -2713 332 -2713 0 feedthrough
rlabel pdiffusion 339 -2713 339 -2713 0 feedthrough
rlabel pdiffusion 346 -2713 346 -2713 0 feedthrough
rlabel pdiffusion 353 -2713 353 -2713 0 feedthrough
rlabel pdiffusion 360 -2713 360 -2713 0 feedthrough
rlabel pdiffusion 367 -2713 367 -2713 0 feedthrough
rlabel pdiffusion 374 -2713 374 -2713 0 feedthrough
rlabel pdiffusion 381 -2713 381 -2713 0 feedthrough
rlabel pdiffusion 388 -2713 388 -2713 0 feedthrough
rlabel pdiffusion 395 -2713 395 -2713 0 feedthrough
rlabel pdiffusion 402 -2713 402 -2713 0 feedthrough
rlabel pdiffusion 409 -2713 409 -2713 0 feedthrough
rlabel pdiffusion 416 -2713 416 -2713 0 feedthrough
rlabel pdiffusion 423 -2713 423 -2713 0 cellNo=284
rlabel pdiffusion 430 -2713 430 -2713 0 feedthrough
rlabel pdiffusion 437 -2713 437 -2713 0 feedthrough
rlabel pdiffusion 444 -2713 444 -2713 0 feedthrough
rlabel pdiffusion 451 -2713 451 -2713 0 feedthrough
rlabel pdiffusion 458 -2713 458 -2713 0 feedthrough
rlabel pdiffusion 465 -2713 465 -2713 0 feedthrough
rlabel pdiffusion 472 -2713 472 -2713 0 feedthrough
rlabel pdiffusion 479 -2713 479 -2713 0 feedthrough
rlabel pdiffusion 486 -2713 486 -2713 0 feedthrough
rlabel pdiffusion 493 -2713 493 -2713 0 feedthrough
rlabel pdiffusion 500 -2713 500 -2713 0 feedthrough
rlabel pdiffusion 507 -2713 507 -2713 0 feedthrough
rlabel pdiffusion 514 -2713 514 -2713 0 feedthrough
rlabel pdiffusion 521 -2713 521 -2713 0 cellNo=139
rlabel pdiffusion 528 -2713 528 -2713 0 feedthrough
rlabel pdiffusion 535 -2713 535 -2713 0 feedthrough
rlabel pdiffusion 542 -2713 542 -2713 0 feedthrough
rlabel pdiffusion 549 -2713 549 -2713 0 feedthrough
rlabel pdiffusion 556 -2713 556 -2713 0 feedthrough
rlabel pdiffusion 563 -2713 563 -2713 0 feedthrough
rlabel pdiffusion 570 -2713 570 -2713 0 feedthrough
rlabel pdiffusion 577 -2713 577 -2713 0 feedthrough
rlabel pdiffusion 584 -2713 584 -2713 0 cellNo=827
rlabel pdiffusion 591 -2713 591 -2713 0 feedthrough
rlabel pdiffusion 598 -2713 598 -2713 0 feedthrough
rlabel pdiffusion 605 -2713 605 -2713 0 cellNo=344
rlabel pdiffusion 612 -2713 612 -2713 0 feedthrough
rlabel pdiffusion 619 -2713 619 -2713 0 feedthrough
rlabel pdiffusion 626 -2713 626 -2713 0 feedthrough
rlabel pdiffusion 633 -2713 633 -2713 0 cellNo=627
rlabel pdiffusion 640 -2713 640 -2713 0 cellNo=249
rlabel pdiffusion 647 -2713 647 -2713 0 feedthrough
rlabel pdiffusion 654 -2713 654 -2713 0 feedthrough
rlabel pdiffusion 661 -2713 661 -2713 0 feedthrough
rlabel pdiffusion 668 -2713 668 -2713 0 feedthrough
rlabel pdiffusion 675 -2713 675 -2713 0 feedthrough
rlabel pdiffusion 682 -2713 682 -2713 0 feedthrough
rlabel pdiffusion 689 -2713 689 -2713 0 feedthrough
rlabel pdiffusion 696 -2713 696 -2713 0 feedthrough
rlabel pdiffusion 703 -2713 703 -2713 0 feedthrough
rlabel pdiffusion 710 -2713 710 -2713 0 cellNo=419
rlabel pdiffusion 717 -2713 717 -2713 0 feedthrough
rlabel pdiffusion 724 -2713 724 -2713 0 feedthrough
rlabel pdiffusion 731 -2713 731 -2713 0 feedthrough
rlabel pdiffusion 738 -2713 738 -2713 0 feedthrough
rlabel pdiffusion 745 -2713 745 -2713 0 feedthrough
rlabel pdiffusion 752 -2713 752 -2713 0 feedthrough
rlabel pdiffusion 759 -2713 759 -2713 0 feedthrough
rlabel pdiffusion 766 -2713 766 -2713 0 feedthrough
rlabel pdiffusion 773 -2713 773 -2713 0 cellNo=292
rlabel pdiffusion 780 -2713 780 -2713 0 feedthrough
rlabel pdiffusion 787 -2713 787 -2713 0 feedthrough
rlabel pdiffusion 794 -2713 794 -2713 0 feedthrough
rlabel pdiffusion 801 -2713 801 -2713 0 feedthrough
rlabel pdiffusion 808 -2713 808 -2713 0 feedthrough
rlabel pdiffusion 815 -2713 815 -2713 0 feedthrough
rlabel pdiffusion 822 -2713 822 -2713 0 feedthrough
rlabel pdiffusion 829 -2713 829 -2713 0 feedthrough
rlabel pdiffusion 836 -2713 836 -2713 0 feedthrough
rlabel pdiffusion 843 -2713 843 -2713 0 cellNo=267
rlabel pdiffusion 850 -2713 850 -2713 0 cellNo=588
rlabel pdiffusion 857 -2713 857 -2713 0 feedthrough
rlabel pdiffusion 864 -2713 864 -2713 0 cellNo=684
rlabel pdiffusion 871 -2713 871 -2713 0 feedthrough
rlabel pdiffusion 878 -2713 878 -2713 0 feedthrough
rlabel pdiffusion 885 -2713 885 -2713 0 cellNo=510
rlabel pdiffusion 892 -2713 892 -2713 0 feedthrough
rlabel pdiffusion 899 -2713 899 -2713 0 feedthrough
rlabel pdiffusion 906 -2713 906 -2713 0 feedthrough
rlabel pdiffusion 913 -2713 913 -2713 0 cellNo=879
rlabel pdiffusion 920 -2713 920 -2713 0 cellNo=288
rlabel pdiffusion 927 -2713 927 -2713 0 feedthrough
rlabel pdiffusion 934 -2713 934 -2713 0 feedthrough
rlabel pdiffusion 941 -2713 941 -2713 0 feedthrough
rlabel pdiffusion 948 -2713 948 -2713 0 feedthrough
rlabel pdiffusion 955 -2713 955 -2713 0 feedthrough
rlabel pdiffusion 962 -2713 962 -2713 0 feedthrough
rlabel pdiffusion 969 -2713 969 -2713 0 feedthrough
rlabel pdiffusion 976 -2713 976 -2713 0 cellNo=724
rlabel pdiffusion 983 -2713 983 -2713 0 feedthrough
rlabel pdiffusion 990 -2713 990 -2713 0 feedthrough
rlabel pdiffusion 997 -2713 997 -2713 0 feedthrough
rlabel pdiffusion 1004 -2713 1004 -2713 0 feedthrough
rlabel pdiffusion 1011 -2713 1011 -2713 0 feedthrough
rlabel pdiffusion 1018 -2713 1018 -2713 0 cellNo=42
rlabel pdiffusion 1025 -2713 1025 -2713 0 feedthrough
rlabel pdiffusion 1032 -2713 1032 -2713 0 feedthrough
rlabel pdiffusion 1039 -2713 1039 -2713 0 feedthrough
rlabel pdiffusion 1046 -2713 1046 -2713 0 feedthrough
rlabel pdiffusion 1053 -2713 1053 -2713 0 cellNo=597
rlabel pdiffusion 1060 -2713 1060 -2713 0 cellNo=566
rlabel pdiffusion 1067 -2713 1067 -2713 0 feedthrough
rlabel pdiffusion 1074 -2713 1074 -2713 0 feedthrough
rlabel pdiffusion 1081 -2713 1081 -2713 0 feedthrough
rlabel pdiffusion 1088 -2713 1088 -2713 0 feedthrough
rlabel pdiffusion 1095 -2713 1095 -2713 0 feedthrough
rlabel pdiffusion 1102 -2713 1102 -2713 0 feedthrough
rlabel pdiffusion 1109 -2713 1109 -2713 0 feedthrough
rlabel pdiffusion 1116 -2713 1116 -2713 0 feedthrough
rlabel pdiffusion 1123 -2713 1123 -2713 0 feedthrough
rlabel pdiffusion 1130 -2713 1130 -2713 0 feedthrough
rlabel pdiffusion 1137 -2713 1137 -2713 0 feedthrough
rlabel pdiffusion 1144 -2713 1144 -2713 0 feedthrough
rlabel pdiffusion 1151 -2713 1151 -2713 0 cellNo=669
rlabel pdiffusion 1158 -2713 1158 -2713 0 feedthrough
rlabel pdiffusion 1165 -2713 1165 -2713 0 feedthrough
rlabel pdiffusion 1172 -2713 1172 -2713 0 feedthrough
rlabel pdiffusion 1179 -2713 1179 -2713 0 feedthrough
rlabel pdiffusion 1186 -2713 1186 -2713 0 feedthrough
rlabel pdiffusion 1193 -2713 1193 -2713 0 cellNo=702
rlabel pdiffusion 1200 -2713 1200 -2713 0 feedthrough
rlabel pdiffusion 1207 -2713 1207 -2713 0 feedthrough
rlabel pdiffusion 1214 -2713 1214 -2713 0 feedthrough
rlabel pdiffusion 1221 -2713 1221 -2713 0 feedthrough
rlabel pdiffusion 1228 -2713 1228 -2713 0 feedthrough
rlabel pdiffusion 1235 -2713 1235 -2713 0 feedthrough
rlabel pdiffusion 1242 -2713 1242 -2713 0 cellNo=550
rlabel pdiffusion 1249 -2713 1249 -2713 0 feedthrough
rlabel pdiffusion 1256 -2713 1256 -2713 0 feedthrough
rlabel pdiffusion 1263 -2713 1263 -2713 0 feedthrough
rlabel pdiffusion 1270 -2713 1270 -2713 0 feedthrough
rlabel pdiffusion 1277 -2713 1277 -2713 0 feedthrough
rlabel pdiffusion 1284 -2713 1284 -2713 0 feedthrough
rlabel pdiffusion 1291 -2713 1291 -2713 0 cellNo=880
rlabel pdiffusion 1298 -2713 1298 -2713 0 feedthrough
rlabel pdiffusion 1305 -2713 1305 -2713 0 feedthrough
rlabel pdiffusion 1312 -2713 1312 -2713 0 feedthrough
rlabel pdiffusion 1319 -2713 1319 -2713 0 cellNo=939
rlabel pdiffusion 1326 -2713 1326 -2713 0 cellNo=49
rlabel pdiffusion 1333 -2713 1333 -2713 0 feedthrough
rlabel pdiffusion 1340 -2713 1340 -2713 0 feedthrough
rlabel pdiffusion 1347 -2713 1347 -2713 0 feedthrough
rlabel pdiffusion 1354 -2713 1354 -2713 0 feedthrough
rlabel pdiffusion 1361 -2713 1361 -2713 0 feedthrough
rlabel pdiffusion 1368 -2713 1368 -2713 0 feedthrough
rlabel pdiffusion 1375 -2713 1375 -2713 0 feedthrough
rlabel pdiffusion 1382 -2713 1382 -2713 0 feedthrough
rlabel pdiffusion 1389 -2713 1389 -2713 0 feedthrough
rlabel pdiffusion 1396 -2713 1396 -2713 0 feedthrough
rlabel pdiffusion 1403 -2713 1403 -2713 0 feedthrough
rlabel pdiffusion 1410 -2713 1410 -2713 0 feedthrough
rlabel pdiffusion 1417 -2713 1417 -2713 0 feedthrough
rlabel pdiffusion 1424 -2713 1424 -2713 0 feedthrough
rlabel pdiffusion 1431 -2713 1431 -2713 0 feedthrough
rlabel pdiffusion 1438 -2713 1438 -2713 0 feedthrough
rlabel pdiffusion 1445 -2713 1445 -2713 0 feedthrough
rlabel pdiffusion 1452 -2713 1452 -2713 0 feedthrough
rlabel pdiffusion 1459 -2713 1459 -2713 0 feedthrough
rlabel pdiffusion 1466 -2713 1466 -2713 0 feedthrough
rlabel pdiffusion 1473 -2713 1473 -2713 0 feedthrough
rlabel pdiffusion 1480 -2713 1480 -2713 0 feedthrough
rlabel pdiffusion 1487 -2713 1487 -2713 0 feedthrough
rlabel pdiffusion 1494 -2713 1494 -2713 0 feedthrough
rlabel pdiffusion 1501 -2713 1501 -2713 0 feedthrough
rlabel pdiffusion 1508 -2713 1508 -2713 0 feedthrough
rlabel pdiffusion 1515 -2713 1515 -2713 0 feedthrough
rlabel pdiffusion 1522 -2713 1522 -2713 0 feedthrough
rlabel pdiffusion 1529 -2713 1529 -2713 0 feedthrough
rlabel pdiffusion 1536 -2713 1536 -2713 0 feedthrough
rlabel pdiffusion 1543 -2713 1543 -2713 0 feedthrough
rlabel pdiffusion 1550 -2713 1550 -2713 0 feedthrough
rlabel pdiffusion 1557 -2713 1557 -2713 0 feedthrough
rlabel pdiffusion 1564 -2713 1564 -2713 0 feedthrough
rlabel pdiffusion 1571 -2713 1571 -2713 0 feedthrough
rlabel pdiffusion 1578 -2713 1578 -2713 0 feedthrough
rlabel pdiffusion 1585 -2713 1585 -2713 0 feedthrough
rlabel pdiffusion 1592 -2713 1592 -2713 0 feedthrough
rlabel pdiffusion 1599 -2713 1599 -2713 0 feedthrough
rlabel pdiffusion 1606 -2713 1606 -2713 0 feedthrough
rlabel pdiffusion 1613 -2713 1613 -2713 0 feedthrough
rlabel pdiffusion 1620 -2713 1620 -2713 0 feedthrough
rlabel pdiffusion 1627 -2713 1627 -2713 0 feedthrough
rlabel pdiffusion 1634 -2713 1634 -2713 0 feedthrough
rlabel pdiffusion 1641 -2713 1641 -2713 0 feedthrough
rlabel pdiffusion 1648 -2713 1648 -2713 0 feedthrough
rlabel pdiffusion 1655 -2713 1655 -2713 0 feedthrough
rlabel pdiffusion 1662 -2713 1662 -2713 0 feedthrough
rlabel pdiffusion 1669 -2713 1669 -2713 0 feedthrough
rlabel pdiffusion 1676 -2713 1676 -2713 0 feedthrough
rlabel pdiffusion 1683 -2713 1683 -2713 0 feedthrough
rlabel pdiffusion 1690 -2713 1690 -2713 0 feedthrough
rlabel pdiffusion 1697 -2713 1697 -2713 0 feedthrough
rlabel pdiffusion 1704 -2713 1704 -2713 0 feedthrough
rlabel pdiffusion 1711 -2713 1711 -2713 0 feedthrough
rlabel pdiffusion 1718 -2713 1718 -2713 0 feedthrough
rlabel pdiffusion 1725 -2713 1725 -2713 0 feedthrough
rlabel pdiffusion 1732 -2713 1732 -2713 0 feedthrough
rlabel pdiffusion 1739 -2713 1739 -2713 0 feedthrough
rlabel pdiffusion 1746 -2713 1746 -2713 0 feedthrough
rlabel pdiffusion 1753 -2713 1753 -2713 0 feedthrough
rlabel pdiffusion 1760 -2713 1760 -2713 0 feedthrough
rlabel pdiffusion 1767 -2713 1767 -2713 0 cellNo=872
rlabel pdiffusion 1774 -2713 1774 -2713 0 cellNo=251
rlabel pdiffusion 1781 -2713 1781 -2713 0 cellNo=81
rlabel pdiffusion 1788 -2713 1788 -2713 0 feedthrough
rlabel pdiffusion 1795 -2713 1795 -2713 0 feedthrough
rlabel pdiffusion 1802 -2713 1802 -2713 0 feedthrough
rlabel pdiffusion 1809 -2713 1809 -2713 0 feedthrough
rlabel pdiffusion 3 -2834 3 -2834 0 cellNo=1028
rlabel pdiffusion 10 -2834 10 -2834 0 cellNo=1153
rlabel pdiffusion 17 -2834 17 -2834 0 cellNo=1040
rlabel pdiffusion 38 -2834 38 -2834 0 feedthrough
rlabel pdiffusion 45 -2834 45 -2834 0 feedthrough
rlabel pdiffusion 52 -2834 52 -2834 0 feedthrough
rlabel pdiffusion 59 -2834 59 -2834 0 feedthrough
rlabel pdiffusion 66 -2834 66 -2834 0 feedthrough
rlabel pdiffusion 73 -2834 73 -2834 0 feedthrough
rlabel pdiffusion 80 -2834 80 -2834 0 feedthrough
rlabel pdiffusion 87 -2834 87 -2834 0 feedthrough
rlabel pdiffusion 94 -2834 94 -2834 0 cellNo=946
rlabel pdiffusion 101 -2834 101 -2834 0 feedthrough
rlabel pdiffusion 108 -2834 108 -2834 0 feedthrough
rlabel pdiffusion 115 -2834 115 -2834 0 feedthrough
rlabel pdiffusion 122 -2834 122 -2834 0 feedthrough
rlabel pdiffusion 129 -2834 129 -2834 0 feedthrough
rlabel pdiffusion 136 -2834 136 -2834 0 feedthrough
rlabel pdiffusion 143 -2834 143 -2834 0 feedthrough
rlabel pdiffusion 150 -2834 150 -2834 0 feedthrough
rlabel pdiffusion 157 -2834 157 -2834 0 feedthrough
rlabel pdiffusion 164 -2834 164 -2834 0 feedthrough
rlabel pdiffusion 171 -2834 171 -2834 0 feedthrough
rlabel pdiffusion 178 -2834 178 -2834 0 feedthrough
rlabel pdiffusion 185 -2834 185 -2834 0 feedthrough
rlabel pdiffusion 192 -2834 192 -2834 0 feedthrough
rlabel pdiffusion 199 -2834 199 -2834 0 feedthrough
rlabel pdiffusion 206 -2834 206 -2834 0 feedthrough
rlabel pdiffusion 213 -2834 213 -2834 0 feedthrough
rlabel pdiffusion 220 -2834 220 -2834 0 feedthrough
rlabel pdiffusion 227 -2834 227 -2834 0 feedthrough
rlabel pdiffusion 234 -2834 234 -2834 0 feedthrough
rlabel pdiffusion 241 -2834 241 -2834 0 feedthrough
rlabel pdiffusion 248 -2834 248 -2834 0 feedthrough
rlabel pdiffusion 255 -2834 255 -2834 0 feedthrough
rlabel pdiffusion 262 -2834 262 -2834 0 feedthrough
rlabel pdiffusion 269 -2834 269 -2834 0 feedthrough
rlabel pdiffusion 276 -2834 276 -2834 0 feedthrough
rlabel pdiffusion 283 -2834 283 -2834 0 feedthrough
rlabel pdiffusion 290 -2834 290 -2834 0 feedthrough
rlabel pdiffusion 297 -2834 297 -2834 0 feedthrough
rlabel pdiffusion 304 -2834 304 -2834 0 feedthrough
rlabel pdiffusion 311 -2834 311 -2834 0 feedthrough
rlabel pdiffusion 318 -2834 318 -2834 0 feedthrough
rlabel pdiffusion 325 -2834 325 -2834 0 feedthrough
rlabel pdiffusion 332 -2834 332 -2834 0 feedthrough
rlabel pdiffusion 339 -2834 339 -2834 0 feedthrough
rlabel pdiffusion 346 -2834 346 -2834 0 feedthrough
rlabel pdiffusion 353 -2834 353 -2834 0 cellNo=638
rlabel pdiffusion 360 -2834 360 -2834 0 feedthrough
rlabel pdiffusion 367 -2834 367 -2834 0 feedthrough
rlabel pdiffusion 374 -2834 374 -2834 0 feedthrough
rlabel pdiffusion 381 -2834 381 -2834 0 feedthrough
rlabel pdiffusion 388 -2834 388 -2834 0 feedthrough
rlabel pdiffusion 395 -2834 395 -2834 0 feedthrough
rlabel pdiffusion 402 -2834 402 -2834 0 feedthrough
rlabel pdiffusion 409 -2834 409 -2834 0 feedthrough
rlabel pdiffusion 416 -2834 416 -2834 0 feedthrough
rlabel pdiffusion 423 -2834 423 -2834 0 feedthrough
rlabel pdiffusion 430 -2834 430 -2834 0 feedthrough
rlabel pdiffusion 437 -2834 437 -2834 0 feedthrough
rlabel pdiffusion 444 -2834 444 -2834 0 feedthrough
rlabel pdiffusion 451 -2834 451 -2834 0 feedthrough
rlabel pdiffusion 458 -2834 458 -2834 0 feedthrough
rlabel pdiffusion 465 -2834 465 -2834 0 feedthrough
rlabel pdiffusion 472 -2834 472 -2834 0 feedthrough
rlabel pdiffusion 479 -2834 479 -2834 0 cellNo=714
rlabel pdiffusion 486 -2834 486 -2834 0 feedthrough
rlabel pdiffusion 493 -2834 493 -2834 0 feedthrough
rlabel pdiffusion 500 -2834 500 -2834 0 feedthrough
rlabel pdiffusion 507 -2834 507 -2834 0 feedthrough
rlabel pdiffusion 514 -2834 514 -2834 0 feedthrough
rlabel pdiffusion 521 -2834 521 -2834 0 feedthrough
rlabel pdiffusion 528 -2834 528 -2834 0 feedthrough
rlabel pdiffusion 535 -2834 535 -2834 0 feedthrough
rlabel pdiffusion 542 -2834 542 -2834 0 feedthrough
rlabel pdiffusion 549 -2834 549 -2834 0 feedthrough
rlabel pdiffusion 556 -2834 556 -2834 0 cellNo=38
rlabel pdiffusion 563 -2834 563 -2834 0 cellNo=799
rlabel pdiffusion 570 -2834 570 -2834 0 feedthrough
rlabel pdiffusion 577 -2834 577 -2834 0 feedthrough
rlabel pdiffusion 584 -2834 584 -2834 0 cellNo=543
rlabel pdiffusion 591 -2834 591 -2834 0 feedthrough
rlabel pdiffusion 598 -2834 598 -2834 0 feedthrough
rlabel pdiffusion 605 -2834 605 -2834 0 feedthrough
rlabel pdiffusion 612 -2834 612 -2834 0 feedthrough
rlabel pdiffusion 619 -2834 619 -2834 0 cellNo=198
rlabel pdiffusion 626 -2834 626 -2834 0 feedthrough
rlabel pdiffusion 633 -2834 633 -2834 0 feedthrough
rlabel pdiffusion 640 -2834 640 -2834 0 feedthrough
rlabel pdiffusion 647 -2834 647 -2834 0 feedthrough
rlabel pdiffusion 654 -2834 654 -2834 0 feedthrough
rlabel pdiffusion 661 -2834 661 -2834 0 cellNo=182
rlabel pdiffusion 668 -2834 668 -2834 0 feedthrough
rlabel pdiffusion 675 -2834 675 -2834 0 feedthrough
rlabel pdiffusion 682 -2834 682 -2834 0 feedthrough
rlabel pdiffusion 689 -2834 689 -2834 0 feedthrough
rlabel pdiffusion 696 -2834 696 -2834 0 feedthrough
rlabel pdiffusion 703 -2834 703 -2834 0 cellNo=652
rlabel pdiffusion 710 -2834 710 -2834 0 cellNo=821
rlabel pdiffusion 717 -2834 717 -2834 0 feedthrough
rlabel pdiffusion 724 -2834 724 -2834 0 feedthrough
rlabel pdiffusion 731 -2834 731 -2834 0 cellNo=519
rlabel pdiffusion 738 -2834 738 -2834 0 feedthrough
rlabel pdiffusion 745 -2834 745 -2834 0 feedthrough
rlabel pdiffusion 752 -2834 752 -2834 0 feedthrough
rlabel pdiffusion 759 -2834 759 -2834 0 feedthrough
rlabel pdiffusion 766 -2834 766 -2834 0 feedthrough
rlabel pdiffusion 773 -2834 773 -2834 0 feedthrough
rlabel pdiffusion 780 -2834 780 -2834 0 feedthrough
rlabel pdiffusion 787 -2834 787 -2834 0 feedthrough
rlabel pdiffusion 794 -2834 794 -2834 0 feedthrough
rlabel pdiffusion 801 -2834 801 -2834 0 feedthrough
rlabel pdiffusion 808 -2834 808 -2834 0 feedthrough
rlabel pdiffusion 815 -2834 815 -2834 0 feedthrough
rlabel pdiffusion 822 -2834 822 -2834 0 feedthrough
rlabel pdiffusion 829 -2834 829 -2834 0 cellNo=866
rlabel pdiffusion 836 -2834 836 -2834 0 feedthrough
rlabel pdiffusion 843 -2834 843 -2834 0 feedthrough
rlabel pdiffusion 850 -2834 850 -2834 0 cellNo=787
rlabel pdiffusion 857 -2834 857 -2834 0 cellNo=737
rlabel pdiffusion 864 -2834 864 -2834 0 feedthrough
rlabel pdiffusion 871 -2834 871 -2834 0 cellNo=580
rlabel pdiffusion 878 -2834 878 -2834 0 feedthrough
rlabel pdiffusion 885 -2834 885 -2834 0 feedthrough
rlabel pdiffusion 892 -2834 892 -2834 0 feedthrough
rlabel pdiffusion 899 -2834 899 -2834 0 feedthrough
rlabel pdiffusion 906 -2834 906 -2834 0 feedthrough
rlabel pdiffusion 913 -2834 913 -2834 0 feedthrough
rlabel pdiffusion 920 -2834 920 -2834 0 feedthrough
rlabel pdiffusion 927 -2834 927 -2834 0 feedthrough
rlabel pdiffusion 934 -2834 934 -2834 0 feedthrough
rlabel pdiffusion 941 -2834 941 -2834 0 feedthrough
rlabel pdiffusion 948 -2834 948 -2834 0 feedthrough
rlabel pdiffusion 955 -2834 955 -2834 0 feedthrough
rlabel pdiffusion 962 -2834 962 -2834 0 feedthrough
rlabel pdiffusion 969 -2834 969 -2834 0 feedthrough
rlabel pdiffusion 976 -2834 976 -2834 0 feedthrough
rlabel pdiffusion 983 -2834 983 -2834 0 feedthrough
rlabel pdiffusion 990 -2834 990 -2834 0 feedthrough
rlabel pdiffusion 997 -2834 997 -2834 0 cellNo=327
rlabel pdiffusion 1004 -2834 1004 -2834 0 feedthrough
rlabel pdiffusion 1011 -2834 1011 -2834 0 cellNo=954
rlabel pdiffusion 1018 -2834 1018 -2834 0 cellNo=760
rlabel pdiffusion 1025 -2834 1025 -2834 0 feedthrough
rlabel pdiffusion 1032 -2834 1032 -2834 0 feedthrough
rlabel pdiffusion 1039 -2834 1039 -2834 0 feedthrough
rlabel pdiffusion 1046 -2834 1046 -2834 0 feedthrough
rlabel pdiffusion 1053 -2834 1053 -2834 0 feedthrough
rlabel pdiffusion 1060 -2834 1060 -2834 0 feedthrough
rlabel pdiffusion 1067 -2834 1067 -2834 0 cellNo=937
rlabel pdiffusion 1074 -2834 1074 -2834 0 feedthrough
rlabel pdiffusion 1081 -2834 1081 -2834 0 feedthrough
rlabel pdiffusion 1088 -2834 1088 -2834 0 feedthrough
rlabel pdiffusion 1095 -2834 1095 -2834 0 feedthrough
rlabel pdiffusion 1102 -2834 1102 -2834 0 feedthrough
rlabel pdiffusion 1109 -2834 1109 -2834 0 feedthrough
rlabel pdiffusion 1116 -2834 1116 -2834 0 cellNo=593
rlabel pdiffusion 1123 -2834 1123 -2834 0 cellNo=159
rlabel pdiffusion 1130 -2834 1130 -2834 0 cellNo=440
rlabel pdiffusion 1137 -2834 1137 -2834 0 feedthrough
rlabel pdiffusion 1144 -2834 1144 -2834 0 feedthrough
rlabel pdiffusion 1151 -2834 1151 -2834 0 feedthrough
rlabel pdiffusion 1158 -2834 1158 -2834 0 feedthrough
rlabel pdiffusion 1165 -2834 1165 -2834 0 feedthrough
rlabel pdiffusion 1172 -2834 1172 -2834 0 feedthrough
rlabel pdiffusion 1179 -2834 1179 -2834 0 cellNo=935
rlabel pdiffusion 1186 -2834 1186 -2834 0 feedthrough
rlabel pdiffusion 1193 -2834 1193 -2834 0 feedthrough
rlabel pdiffusion 1200 -2834 1200 -2834 0 cellNo=356
rlabel pdiffusion 1207 -2834 1207 -2834 0 feedthrough
rlabel pdiffusion 1214 -2834 1214 -2834 0 feedthrough
rlabel pdiffusion 1221 -2834 1221 -2834 0 feedthrough
rlabel pdiffusion 1228 -2834 1228 -2834 0 feedthrough
rlabel pdiffusion 1235 -2834 1235 -2834 0 cellNo=901
rlabel pdiffusion 1242 -2834 1242 -2834 0 feedthrough
rlabel pdiffusion 1249 -2834 1249 -2834 0 feedthrough
rlabel pdiffusion 1256 -2834 1256 -2834 0 feedthrough
rlabel pdiffusion 1263 -2834 1263 -2834 0 feedthrough
rlabel pdiffusion 1270 -2834 1270 -2834 0 feedthrough
rlabel pdiffusion 1277 -2834 1277 -2834 0 feedthrough
rlabel pdiffusion 1284 -2834 1284 -2834 0 cellNo=414
rlabel pdiffusion 1291 -2834 1291 -2834 0 feedthrough
rlabel pdiffusion 1298 -2834 1298 -2834 0 feedthrough
rlabel pdiffusion 1305 -2834 1305 -2834 0 feedthrough
rlabel pdiffusion 1312 -2834 1312 -2834 0 feedthrough
rlabel pdiffusion 1319 -2834 1319 -2834 0 feedthrough
rlabel pdiffusion 1326 -2834 1326 -2834 0 feedthrough
rlabel pdiffusion 1333 -2834 1333 -2834 0 feedthrough
rlabel pdiffusion 1340 -2834 1340 -2834 0 cellNo=585
rlabel pdiffusion 1347 -2834 1347 -2834 0 feedthrough
rlabel pdiffusion 1354 -2834 1354 -2834 0 cellNo=835
rlabel pdiffusion 1361 -2834 1361 -2834 0 feedthrough
rlabel pdiffusion 1368 -2834 1368 -2834 0 feedthrough
rlabel pdiffusion 1375 -2834 1375 -2834 0 feedthrough
rlabel pdiffusion 1382 -2834 1382 -2834 0 feedthrough
rlabel pdiffusion 1389 -2834 1389 -2834 0 feedthrough
rlabel pdiffusion 1396 -2834 1396 -2834 0 feedthrough
rlabel pdiffusion 1403 -2834 1403 -2834 0 feedthrough
rlabel pdiffusion 1410 -2834 1410 -2834 0 feedthrough
rlabel pdiffusion 1417 -2834 1417 -2834 0 feedthrough
rlabel pdiffusion 1424 -2834 1424 -2834 0 feedthrough
rlabel pdiffusion 1431 -2834 1431 -2834 0 cellNo=395
rlabel pdiffusion 1438 -2834 1438 -2834 0 feedthrough
rlabel pdiffusion 1445 -2834 1445 -2834 0 feedthrough
rlabel pdiffusion 1452 -2834 1452 -2834 0 feedthrough
rlabel pdiffusion 1459 -2834 1459 -2834 0 feedthrough
rlabel pdiffusion 1466 -2834 1466 -2834 0 feedthrough
rlabel pdiffusion 1473 -2834 1473 -2834 0 feedthrough
rlabel pdiffusion 1480 -2834 1480 -2834 0 feedthrough
rlabel pdiffusion 1487 -2834 1487 -2834 0 feedthrough
rlabel pdiffusion 1494 -2834 1494 -2834 0 feedthrough
rlabel pdiffusion 1501 -2834 1501 -2834 0 feedthrough
rlabel pdiffusion 1508 -2834 1508 -2834 0 feedthrough
rlabel pdiffusion 1515 -2834 1515 -2834 0 feedthrough
rlabel pdiffusion 1522 -2834 1522 -2834 0 feedthrough
rlabel pdiffusion 1529 -2834 1529 -2834 0 feedthrough
rlabel pdiffusion 1536 -2834 1536 -2834 0 feedthrough
rlabel pdiffusion 1543 -2834 1543 -2834 0 feedthrough
rlabel pdiffusion 1550 -2834 1550 -2834 0 feedthrough
rlabel pdiffusion 1557 -2834 1557 -2834 0 feedthrough
rlabel pdiffusion 1564 -2834 1564 -2834 0 feedthrough
rlabel pdiffusion 1571 -2834 1571 -2834 0 feedthrough
rlabel pdiffusion 1578 -2834 1578 -2834 0 feedthrough
rlabel pdiffusion 1585 -2834 1585 -2834 0 feedthrough
rlabel pdiffusion 1592 -2834 1592 -2834 0 feedthrough
rlabel pdiffusion 1599 -2834 1599 -2834 0 feedthrough
rlabel pdiffusion 1606 -2834 1606 -2834 0 feedthrough
rlabel pdiffusion 1613 -2834 1613 -2834 0 feedthrough
rlabel pdiffusion 1620 -2834 1620 -2834 0 feedthrough
rlabel pdiffusion 1627 -2834 1627 -2834 0 feedthrough
rlabel pdiffusion 1634 -2834 1634 -2834 0 feedthrough
rlabel pdiffusion 1641 -2834 1641 -2834 0 feedthrough
rlabel pdiffusion 1648 -2834 1648 -2834 0 feedthrough
rlabel pdiffusion 1655 -2834 1655 -2834 0 feedthrough
rlabel pdiffusion 1662 -2834 1662 -2834 0 feedthrough
rlabel pdiffusion 1669 -2834 1669 -2834 0 feedthrough
rlabel pdiffusion 1676 -2834 1676 -2834 0 feedthrough
rlabel pdiffusion 1683 -2834 1683 -2834 0 feedthrough
rlabel pdiffusion 1690 -2834 1690 -2834 0 feedthrough
rlabel pdiffusion 1697 -2834 1697 -2834 0 feedthrough
rlabel pdiffusion 1704 -2834 1704 -2834 0 feedthrough
rlabel pdiffusion 1711 -2834 1711 -2834 0 cellNo=272
rlabel pdiffusion 1718 -2834 1718 -2834 0 cellNo=887
rlabel pdiffusion 1725 -2834 1725 -2834 0 cellNo=57
rlabel pdiffusion 1732 -2834 1732 -2834 0 feedthrough
rlabel pdiffusion 1739 -2834 1739 -2834 0 feedthrough
rlabel pdiffusion 1746 -2834 1746 -2834 0 feedthrough
rlabel pdiffusion 1753 -2834 1753 -2834 0 feedthrough
rlabel pdiffusion 1760 -2834 1760 -2834 0 feedthrough
rlabel pdiffusion 1767 -2834 1767 -2834 0 feedthrough
rlabel pdiffusion 1774 -2834 1774 -2834 0 feedthrough
rlabel pdiffusion 3 -2953 3 -2953 0 cellNo=1032
rlabel pdiffusion 10 -2953 10 -2953 0 cellNo=1172
rlabel pdiffusion 17 -2953 17 -2953 0 cellNo=1036
rlabel pdiffusion 24 -2953 24 -2953 0 feedthrough
rlabel pdiffusion 31 -2953 31 -2953 0 cellNo=1063
rlabel pdiffusion 38 -2953 38 -2953 0 cellNo=1141
rlabel pdiffusion 45 -2953 45 -2953 0 cellNo=1154
rlabel pdiffusion 52 -2953 52 -2953 0 feedthrough
rlabel pdiffusion 59 -2953 59 -2953 0 feedthrough
rlabel pdiffusion 66 -2953 66 -2953 0 feedthrough
rlabel pdiffusion 73 -2953 73 -2953 0 feedthrough
rlabel pdiffusion 80 -2953 80 -2953 0 cellNo=962
rlabel pdiffusion 87 -2953 87 -2953 0 feedthrough
rlabel pdiffusion 94 -2953 94 -2953 0 feedthrough
rlabel pdiffusion 101 -2953 101 -2953 0 feedthrough
rlabel pdiffusion 108 -2953 108 -2953 0 cellNo=421
rlabel pdiffusion 115 -2953 115 -2953 0 feedthrough
rlabel pdiffusion 122 -2953 122 -2953 0 feedthrough
rlabel pdiffusion 129 -2953 129 -2953 0 feedthrough
rlabel pdiffusion 136 -2953 136 -2953 0 cellNo=305
rlabel pdiffusion 143 -2953 143 -2953 0 cellNo=868
rlabel pdiffusion 150 -2953 150 -2953 0 feedthrough
rlabel pdiffusion 157 -2953 157 -2953 0 feedthrough
rlabel pdiffusion 164 -2953 164 -2953 0 cellNo=92
rlabel pdiffusion 171 -2953 171 -2953 0 feedthrough
rlabel pdiffusion 178 -2953 178 -2953 0 feedthrough
rlabel pdiffusion 185 -2953 185 -2953 0 feedthrough
rlabel pdiffusion 192 -2953 192 -2953 0 feedthrough
rlabel pdiffusion 199 -2953 199 -2953 0 feedthrough
rlabel pdiffusion 206 -2953 206 -2953 0 cellNo=656
rlabel pdiffusion 213 -2953 213 -2953 0 feedthrough
rlabel pdiffusion 220 -2953 220 -2953 0 cellNo=603
rlabel pdiffusion 227 -2953 227 -2953 0 cellNo=506
rlabel pdiffusion 234 -2953 234 -2953 0 feedthrough
rlabel pdiffusion 241 -2953 241 -2953 0 feedthrough
rlabel pdiffusion 248 -2953 248 -2953 0 feedthrough
rlabel pdiffusion 255 -2953 255 -2953 0 feedthrough
rlabel pdiffusion 262 -2953 262 -2953 0 feedthrough
rlabel pdiffusion 269 -2953 269 -2953 0 feedthrough
rlabel pdiffusion 276 -2953 276 -2953 0 feedthrough
rlabel pdiffusion 283 -2953 283 -2953 0 feedthrough
rlabel pdiffusion 290 -2953 290 -2953 0 feedthrough
rlabel pdiffusion 297 -2953 297 -2953 0 feedthrough
rlabel pdiffusion 304 -2953 304 -2953 0 feedthrough
rlabel pdiffusion 311 -2953 311 -2953 0 feedthrough
rlabel pdiffusion 318 -2953 318 -2953 0 feedthrough
rlabel pdiffusion 325 -2953 325 -2953 0 feedthrough
rlabel pdiffusion 332 -2953 332 -2953 0 feedthrough
rlabel pdiffusion 339 -2953 339 -2953 0 feedthrough
rlabel pdiffusion 346 -2953 346 -2953 0 feedthrough
rlabel pdiffusion 353 -2953 353 -2953 0 feedthrough
rlabel pdiffusion 360 -2953 360 -2953 0 feedthrough
rlabel pdiffusion 367 -2953 367 -2953 0 feedthrough
rlabel pdiffusion 374 -2953 374 -2953 0 feedthrough
rlabel pdiffusion 381 -2953 381 -2953 0 feedthrough
rlabel pdiffusion 388 -2953 388 -2953 0 feedthrough
rlabel pdiffusion 395 -2953 395 -2953 0 feedthrough
rlabel pdiffusion 402 -2953 402 -2953 0 feedthrough
rlabel pdiffusion 409 -2953 409 -2953 0 cellNo=867
rlabel pdiffusion 416 -2953 416 -2953 0 feedthrough
rlabel pdiffusion 423 -2953 423 -2953 0 feedthrough
rlabel pdiffusion 430 -2953 430 -2953 0 feedthrough
rlabel pdiffusion 437 -2953 437 -2953 0 cellNo=629
rlabel pdiffusion 444 -2953 444 -2953 0 feedthrough
rlabel pdiffusion 451 -2953 451 -2953 0 feedthrough
rlabel pdiffusion 458 -2953 458 -2953 0 feedthrough
rlabel pdiffusion 465 -2953 465 -2953 0 cellNo=162
rlabel pdiffusion 472 -2953 472 -2953 0 feedthrough
rlabel pdiffusion 479 -2953 479 -2953 0 feedthrough
rlabel pdiffusion 486 -2953 486 -2953 0 feedthrough
rlabel pdiffusion 493 -2953 493 -2953 0 feedthrough
rlabel pdiffusion 500 -2953 500 -2953 0 feedthrough
rlabel pdiffusion 507 -2953 507 -2953 0 feedthrough
rlabel pdiffusion 514 -2953 514 -2953 0 feedthrough
rlabel pdiffusion 521 -2953 521 -2953 0 feedthrough
rlabel pdiffusion 528 -2953 528 -2953 0 feedthrough
rlabel pdiffusion 535 -2953 535 -2953 0 cellNo=696
rlabel pdiffusion 542 -2953 542 -2953 0 feedthrough
rlabel pdiffusion 549 -2953 549 -2953 0 feedthrough
rlabel pdiffusion 556 -2953 556 -2953 0 feedthrough
rlabel pdiffusion 563 -2953 563 -2953 0 feedthrough
rlabel pdiffusion 570 -2953 570 -2953 0 feedthrough
rlabel pdiffusion 577 -2953 577 -2953 0 feedthrough
rlabel pdiffusion 584 -2953 584 -2953 0 feedthrough
rlabel pdiffusion 591 -2953 591 -2953 0 feedthrough
rlabel pdiffusion 598 -2953 598 -2953 0 feedthrough
rlabel pdiffusion 605 -2953 605 -2953 0 feedthrough
rlabel pdiffusion 612 -2953 612 -2953 0 feedthrough
rlabel pdiffusion 619 -2953 619 -2953 0 feedthrough
rlabel pdiffusion 626 -2953 626 -2953 0 feedthrough
rlabel pdiffusion 633 -2953 633 -2953 0 feedthrough
rlabel pdiffusion 640 -2953 640 -2953 0 feedthrough
rlabel pdiffusion 647 -2953 647 -2953 0 feedthrough
rlabel pdiffusion 654 -2953 654 -2953 0 cellNo=129
rlabel pdiffusion 661 -2953 661 -2953 0 cellNo=224
rlabel pdiffusion 668 -2953 668 -2953 0 feedthrough
rlabel pdiffusion 675 -2953 675 -2953 0 feedthrough
rlabel pdiffusion 682 -2953 682 -2953 0 feedthrough
rlabel pdiffusion 689 -2953 689 -2953 0 feedthrough
rlabel pdiffusion 696 -2953 696 -2953 0 feedthrough
rlabel pdiffusion 703 -2953 703 -2953 0 feedthrough
rlabel pdiffusion 710 -2953 710 -2953 0 feedthrough
rlabel pdiffusion 717 -2953 717 -2953 0 feedthrough
rlabel pdiffusion 724 -2953 724 -2953 0 feedthrough
rlabel pdiffusion 731 -2953 731 -2953 0 feedthrough
rlabel pdiffusion 738 -2953 738 -2953 0 feedthrough
rlabel pdiffusion 745 -2953 745 -2953 0 feedthrough
rlabel pdiffusion 752 -2953 752 -2953 0 feedthrough
rlabel pdiffusion 759 -2953 759 -2953 0 feedthrough
rlabel pdiffusion 766 -2953 766 -2953 0 feedthrough
rlabel pdiffusion 773 -2953 773 -2953 0 feedthrough
rlabel pdiffusion 780 -2953 780 -2953 0 cellNo=742
rlabel pdiffusion 787 -2953 787 -2953 0 feedthrough
rlabel pdiffusion 794 -2953 794 -2953 0 feedthrough
rlabel pdiffusion 801 -2953 801 -2953 0 feedthrough
rlabel pdiffusion 808 -2953 808 -2953 0 feedthrough
rlabel pdiffusion 815 -2953 815 -2953 0 feedthrough
rlabel pdiffusion 822 -2953 822 -2953 0 cellNo=733
rlabel pdiffusion 829 -2953 829 -2953 0 feedthrough
rlabel pdiffusion 836 -2953 836 -2953 0 feedthrough
rlabel pdiffusion 843 -2953 843 -2953 0 feedthrough
rlabel pdiffusion 850 -2953 850 -2953 0 cellNo=375
rlabel pdiffusion 857 -2953 857 -2953 0 feedthrough
rlabel pdiffusion 864 -2953 864 -2953 0 cellNo=619
rlabel pdiffusion 871 -2953 871 -2953 0 feedthrough
rlabel pdiffusion 878 -2953 878 -2953 0 feedthrough
rlabel pdiffusion 885 -2953 885 -2953 0 feedthrough
rlabel pdiffusion 892 -2953 892 -2953 0 feedthrough
rlabel pdiffusion 899 -2953 899 -2953 0 feedthrough
rlabel pdiffusion 906 -2953 906 -2953 0 feedthrough
rlabel pdiffusion 913 -2953 913 -2953 0 cellNo=768
rlabel pdiffusion 920 -2953 920 -2953 0 feedthrough
rlabel pdiffusion 927 -2953 927 -2953 0 feedthrough
rlabel pdiffusion 934 -2953 934 -2953 0 feedthrough
rlabel pdiffusion 941 -2953 941 -2953 0 cellNo=481
rlabel pdiffusion 948 -2953 948 -2953 0 feedthrough
rlabel pdiffusion 955 -2953 955 -2953 0 feedthrough
rlabel pdiffusion 962 -2953 962 -2953 0 feedthrough
rlabel pdiffusion 969 -2953 969 -2953 0 cellNo=909
rlabel pdiffusion 976 -2953 976 -2953 0 feedthrough
rlabel pdiffusion 983 -2953 983 -2953 0 feedthrough
rlabel pdiffusion 990 -2953 990 -2953 0 feedthrough
rlabel pdiffusion 997 -2953 997 -2953 0 feedthrough
rlabel pdiffusion 1004 -2953 1004 -2953 0 feedthrough
rlabel pdiffusion 1011 -2953 1011 -2953 0 feedthrough
rlabel pdiffusion 1018 -2953 1018 -2953 0 feedthrough
rlabel pdiffusion 1025 -2953 1025 -2953 0 cellNo=899
rlabel pdiffusion 1032 -2953 1032 -2953 0 cellNo=275
rlabel pdiffusion 1039 -2953 1039 -2953 0 feedthrough
rlabel pdiffusion 1046 -2953 1046 -2953 0 feedthrough
rlabel pdiffusion 1053 -2953 1053 -2953 0 cellNo=220
rlabel pdiffusion 1060 -2953 1060 -2953 0 feedthrough
rlabel pdiffusion 1067 -2953 1067 -2953 0 feedthrough
rlabel pdiffusion 1074 -2953 1074 -2953 0 feedthrough
rlabel pdiffusion 1081 -2953 1081 -2953 0 feedthrough
rlabel pdiffusion 1088 -2953 1088 -2953 0 feedthrough
rlabel pdiffusion 1095 -2953 1095 -2953 0 cellNo=949
rlabel pdiffusion 1102 -2953 1102 -2953 0 feedthrough
rlabel pdiffusion 1109 -2953 1109 -2953 0 feedthrough
rlabel pdiffusion 1116 -2953 1116 -2953 0 feedthrough
rlabel pdiffusion 1123 -2953 1123 -2953 0 feedthrough
rlabel pdiffusion 1130 -2953 1130 -2953 0 feedthrough
rlabel pdiffusion 1137 -2953 1137 -2953 0 feedthrough
rlabel pdiffusion 1144 -2953 1144 -2953 0 feedthrough
rlabel pdiffusion 1151 -2953 1151 -2953 0 feedthrough
rlabel pdiffusion 1158 -2953 1158 -2953 0 feedthrough
rlabel pdiffusion 1165 -2953 1165 -2953 0 feedthrough
rlabel pdiffusion 1172 -2953 1172 -2953 0 feedthrough
rlabel pdiffusion 1179 -2953 1179 -2953 0 feedthrough
rlabel pdiffusion 1186 -2953 1186 -2953 0 feedthrough
rlabel pdiffusion 1193 -2953 1193 -2953 0 feedthrough
rlabel pdiffusion 1200 -2953 1200 -2953 0 cellNo=165
rlabel pdiffusion 1207 -2953 1207 -2953 0 feedthrough
rlabel pdiffusion 1214 -2953 1214 -2953 0 feedthrough
rlabel pdiffusion 1221 -2953 1221 -2953 0 feedthrough
rlabel pdiffusion 1228 -2953 1228 -2953 0 feedthrough
rlabel pdiffusion 1235 -2953 1235 -2953 0 feedthrough
rlabel pdiffusion 1242 -2953 1242 -2953 0 feedthrough
rlabel pdiffusion 1249 -2953 1249 -2953 0 feedthrough
rlabel pdiffusion 1256 -2953 1256 -2953 0 feedthrough
rlabel pdiffusion 1263 -2953 1263 -2953 0 feedthrough
rlabel pdiffusion 1270 -2953 1270 -2953 0 feedthrough
rlabel pdiffusion 1277 -2953 1277 -2953 0 feedthrough
rlabel pdiffusion 1284 -2953 1284 -2953 0 feedthrough
rlabel pdiffusion 1291 -2953 1291 -2953 0 feedthrough
rlabel pdiffusion 1298 -2953 1298 -2953 0 feedthrough
rlabel pdiffusion 1305 -2953 1305 -2953 0 feedthrough
rlabel pdiffusion 1312 -2953 1312 -2953 0 feedthrough
rlabel pdiffusion 1319 -2953 1319 -2953 0 feedthrough
rlabel pdiffusion 1326 -2953 1326 -2953 0 feedthrough
rlabel pdiffusion 1333 -2953 1333 -2953 0 cellNo=785
rlabel pdiffusion 1340 -2953 1340 -2953 0 feedthrough
rlabel pdiffusion 1347 -2953 1347 -2953 0 feedthrough
rlabel pdiffusion 1354 -2953 1354 -2953 0 feedthrough
rlabel pdiffusion 1361 -2953 1361 -2953 0 feedthrough
rlabel pdiffusion 1368 -2953 1368 -2953 0 feedthrough
rlabel pdiffusion 1375 -2953 1375 -2953 0 feedthrough
rlabel pdiffusion 1382 -2953 1382 -2953 0 feedthrough
rlabel pdiffusion 1389 -2953 1389 -2953 0 feedthrough
rlabel pdiffusion 1396 -2953 1396 -2953 0 feedthrough
rlabel pdiffusion 1403 -2953 1403 -2953 0 feedthrough
rlabel pdiffusion 1410 -2953 1410 -2953 0 feedthrough
rlabel pdiffusion 1417 -2953 1417 -2953 0 feedthrough
rlabel pdiffusion 1424 -2953 1424 -2953 0 feedthrough
rlabel pdiffusion 1431 -2953 1431 -2953 0 feedthrough
rlabel pdiffusion 1438 -2953 1438 -2953 0 feedthrough
rlabel pdiffusion 1445 -2953 1445 -2953 0 feedthrough
rlabel pdiffusion 1452 -2953 1452 -2953 0 feedthrough
rlabel pdiffusion 1459 -2953 1459 -2953 0 feedthrough
rlabel pdiffusion 1466 -2953 1466 -2953 0 feedthrough
rlabel pdiffusion 1473 -2953 1473 -2953 0 feedthrough
rlabel pdiffusion 1480 -2953 1480 -2953 0 feedthrough
rlabel pdiffusion 1487 -2953 1487 -2953 0 feedthrough
rlabel pdiffusion 1494 -2953 1494 -2953 0 feedthrough
rlabel pdiffusion 1501 -2953 1501 -2953 0 feedthrough
rlabel pdiffusion 1508 -2953 1508 -2953 0 feedthrough
rlabel pdiffusion 1515 -2953 1515 -2953 0 feedthrough
rlabel pdiffusion 1522 -2953 1522 -2953 0 feedthrough
rlabel pdiffusion 1529 -2953 1529 -2953 0 feedthrough
rlabel pdiffusion 1536 -2953 1536 -2953 0 feedthrough
rlabel pdiffusion 1543 -2953 1543 -2953 0 feedthrough
rlabel pdiffusion 1550 -2953 1550 -2953 0 feedthrough
rlabel pdiffusion 1557 -2953 1557 -2953 0 feedthrough
rlabel pdiffusion 1564 -2953 1564 -2953 0 feedthrough
rlabel pdiffusion 1571 -2953 1571 -2953 0 feedthrough
rlabel pdiffusion 1578 -2953 1578 -2953 0 feedthrough
rlabel pdiffusion 1585 -2953 1585 -2953 0 feedthrough
rlabel pdiffusion 1592 -2953 1592 -2953 0 feedthrough
rlabel pdiffusion 1599 -2953 1599 -2953 0 feedthrough
rlabel pdiffusion 1606 -2953 1606 -2953 0 feedthrough
rlabel pdiffusion 1613 -2953 1613 -2953 0 feedthrough
rlabel pdiffusion 1620 -2953 1620 -2953 0 feedthrough
rlabel pdiffusion 1627 -2953 1627 -2953 0 feedthrough
rlabel pdiffusion 1634 -2953 1634 -2953 0 feedthrough
rlabel pdiffusion 1641 -2953 1641 -2953 0 cellNo=174
rlabel pdiffusion 1648 -2953 1648 -2953 0 feedthrough
rlabel pdiffusion 1655 -2953 1655 -2953 0 feedthrough
rlabel pdiffusion 1662 -2953 1662 -2953 0 feedthrough
rlabel pdiffusion 1669 -2953 1669 -2953 0 feedthrough
rlabel pdiffusion 1676 -2953 1676 -2953 0 feedthrough
rlabel pdiffusion 1683 -2953 1683 -2953 0 feedthrough
rlabel pdiffusion 1690 -2953 1690 -2953 0 feedthrough
rlabel pdiffusion 1697 -2953 1697 -2953 0 feedthrough
rlabel pdiffusion 1704 -2953 1704 -2953 0 cellNo=561
rlabel pdiffusion 3 -3080 3 -3080 0 cellNo=1030
rlabel pdiffusion 10 -3080 10 -3080 0 cellNo=1035
rlabel pdiffusion 17 -3080 17 -3080 0 cellNo=1038
rlabel pdiffusion 24 -3080 24 -3080 0 cellNo=1148
rlabel pdiffusion 31 -3080 31 -3080 0 feedthrough
rlabel pdiffusion 38 -3080 38 -3080 0 feedthrough
rlabel pdiffusion 45 -3080 45 -3080 0 feedthrough
rlabel pdiffusion 52 -3080 52 -3080 0 feedthrough
rlabel pdiffusion 59 -3080 59 -3080 0 cellNo=943
rlabel pdiffusion 66 -3080 66 -3080 0 feedthrough
rlabel pdiffusion 73 -3080 73 -3080 0 feedthrough
rlabel pdiffusion 80 -3080 80 -3080 0 cellNo=688
rlabel pdiffusion 87 -3080 87 -3080 0 cellNo=218
rlabel pdiffusion 94 -3080 94 -3080 0 feedthrough
rlabel pdiffusion 101 -3080 101 -3080 0 feedthrough
rlabel pdiffusion 108 -3080 108 -3080 0 feedthrough
rlabel pdiffusion 115 -3080 115 -3080 0 feedthrough
rlabel pdiffusion 122 -3080 122 -3080 0 feedthrough
rlabel pdiffusion 129 -3080 129 -3080 0 feedthrough
rlabel pdiffusion 136 -3080 136 -3080 0 cellNo=608
rlabel pdiffusion 143 -3080 143 -3080 0 cellNo=770
rlabel pdiffusion 150 -3080 150 -3080 0 cellNo=723
rlabel pdiffusion 157 -3080 157 -3080 0 feedthrough
rlabel pdiffusion 164 -3080 164 -3080 0 feedthrough
rlabel pdiffusion 171 -3080 171 -3080 0 feedthrough
rlabel pdiffusion 178 -3080 178 -3080 0 feedthrough
rlabel pdiffusion 185 -3080 185 -3080 0 cellNo=851
rlabel pdiffusion 192 -3080 192 -3080 0 feedthrough
rlabel pdiffusion 199 -3080 199 -3080 0 cellNo=942
rlabel pdiffusion 206 -3080 206 -3080 0 cellNo=415
rlabel pdiffusion 213 -3080 213 -3080 0 cellNo=501
rlabel pdiffusion 220 -3080 220 -3080 0 feedthrough
rlabel pdiffusion 227 -3080 227 -3080 0 feedthrough
rlabel pdiffusion 234 -3080 234 -3080 0 feedthrough
rlabel pdiffusion 241 -3080 241 -3080 0 feedthrough
rlabel pdiffusion 248 -3080 248 -3080 0 feedthrough
rlabel pdiffusion 255 -3080 255 -3080 0 feedthrough
rlabel pdiffusion 262 -3080 262 -3080 0 feedthrough
rlabel pdiffusion 269 -3080 269 -3080 0 feedthrough
rlabel pdiffusion 276 -3080 276 -3080 0 feedthrough
rlabel pdiffusion 283 -3080 283 -3080 0 feedthrough
rlabel pdiffusion 290 -3080 290 -3080 0 feedthrough
rlabel pdiffusion 297 -3080 297 -3080 0 feedthrough
rlabel pdiffusion 304 -3080 304 -3080 0 feedthrough
rlabel pdiffusion 311 -3080 311 -3080 0 feedthrough
rlabel pdiffusion 318 -3080 318 -3080 0 feedthrough
rlabel pdiffusion 325 -3080 325 -3080 0 feedthrough
rlabel pdiffusion 332 -3080 332 -3080 0 feedthrough
rlabel pdiffusion 339 -3080 339 -3080 0 feedthrough
rlabel pdiffusion 346 -3080 346 -3080 0 cellNo=150
rlabel pdiffusion 353 -3080 353 -3080 0 feedthrough
rlabel pdiffusion 360 -3080 360 -3080 0 feedthrough
rlabel pdiffusion 367 -3080 367 -3080 0 cellNo=111
rlabel pdiffusion 374 -3080 374 -3080 0 feedthrough
rlabel pdiffusion 381 -3080 381 -3080 0 feedthrough
rlabel pdiffusion 388 -3080 388 -3080 0 feedthrough
rlabel pdiffusion 395 -3080 395 -3080 0 cellNo=950
rlabel pdiffusion 402 -3080 402 -3080 0 feedthrough
rlabel pdiffusion 409 -3080 409 -3080 0 feedthrough
rlabel pdiffusion 416 -3080 416 -3080 0 feedthrough
rlabel pdiffusion 423 -3080 423 -3080 0 feedthrough
rlabel pdiffusion 430 -3080 430 -3080 0 feedthrough
rlabel pdiffusion 437 -3080 437 -3080 0 feedthrough
rlabel pdiffusion 444 -3080 444 -3080 0 feedthrough
rlabel pdiffusion 451 -3080 451 -3080 0 cellNo=924
rlabel pdiffusion 458 -3080 458 -3080 0 feedthrough
rlabel pdiffusion 465 -3080 465 -3080 0 feedthrough
rlabel pdiffusion 472 -3080 472 -3080 0 feedthrough
rlabel pdiffusion 479 -3080 479 -3080 0 feedthrough
rlabel pdiffusion 486 -3080 486 -3080 0 feedthrough
rlabel pdiffusion 493 -3080 493 -3080 0 feedthrough
rlabel pdiffusion 500 -3080 500 -3080 0 feedthrough
rlabel pdiffusion 507 -3080 507 -3080 0 feedthrough
rlabel pdiffusion 514 -3080 514 -3080 0 feedthrough
rlabel pdiffusion 521 -3080 521 -3080 0 feedthrough
rlabel pdiffusion 528 -3080 528 -3080 0 feedthrough
rlabel pdiffusion 535 -3080 535 -3080 0 feedthrough
rlabel pdiffusion 542 -3080 542 -3080 0 feedthrough
rlabel pdiffusion 549 -3080 549 -3080 0 feedthrough
rlabel pdiffusion 556 -3080 556 -3080 0 feedthrough
rlabel pdiffusion 563 -3080 563 -3080 0 feedthrough
rlabel pdiffusion 570 -3080 570 -3080 0 feedthrough
rlabel pdiffusion 577 -3080 577 -3080 0 feedthrough
rlabel pdiffusion 584 -3080 584 -3080 0 feedthrough
rlabel pdiffusion 591 -3080 591 -3080 0 feedthrough
rlabel pdiffusion 598 -3080 598 -3080 0 feedthrough
rlabel pdiffusion 605 -3080 605 -3080 0 feedthrough
rlabel pdiffusion 612 -3080 612 -3080 0 feedthrough
rlabel pdiffusion 619 -3080 619 -3080 0 cellNo=361
rlabel pdiffusion 626 -3080 626 -3080 0 feedthrough
rlabel pdiffusion 633 -3080 633 -3080 0 cellNo=504
rlabel pdiffusion 640 -3080 640 -3080 0 feedthrough
rlabel pdiffusion 647 -3080 647 -3080 0 feedthrough
rlabel pdiffusion 654 -3080 654 -3080 0 feedthrough
rlabel pdiffusion 661 -3080 661 -3080 0 feedthrough
rlabel pdiffusion 668 -3080 668 -3080 0 feedthrough
rlabel pdiffusion 675 -3080 675 -3080 0 feedthrough
rlabel pdiffusion 682 -3080 682 -3080 0 feedthrough
rlabel pdiffusion 689 -3080 689 -3080 0 cellNo=903
rlabel pdiffusion 696 -3080 696 -3080 0 feedthrough
rlabel pdiffusion 703 -3080 703 -3080 0 feedthrough
rlabel pdiffusion 710 -3080 710 -3080 0 feedthrough
rlabel pdiffusion 717 -3080 717 -3080 0 feedthrough
rlabel pdiffusion 724 -3080 724 -3080 0 feedthrough
rlabel pdiffusion 731 -3080 731 -3080 0 feedthrough
rlabel pdiffusion 738 -3080 738 -3080 0 cellNo=402
rlabel pdiffusion 745 -3080 745 -3080 0 feedthrough
rlabel pdiffusion 752 -3080 752 -3080 0 feedthrough
rlabel pdiffusion 759 -3080 759 -3080 0 cellNo=847
rlabel pdiffusion 766 -3080 766 -3080 0 feedthrough
rlabel pdiffusion 773 -3080 773 -3080 0 feedthrough
rlabel pdiffusion 780 -3080 780 -3080 0 feedthrough
rlabel pdiffusion 787 -3080 787 -3080 0 cellNo=355
rlabel pdiffusion 794 -3080 794 -3080 0 feedthrough
rlabel pdiffusion 801 -3080 801 -3080 0 cellNo=270
rlabel pdiffusion 808 -3080 808 -3080 0 feedthrough
rlabel pdiffusion 815 -3080 815 -3080 0 feedthrough
rlabel pdiffusion 822 -3080 822 -3080 0 feedthrough
rlabel pdiffusion 829 -3080 829 -3080 0 cellNo=796
rlabel pdiffusion 836 -3080 836 -3080 0 cellNo=544
rlabel pdiffusion 843 -3080 843 -3080 0 feedthrough
rlabel pdiffusion 850 -3080 850 -3080 0 feedthrough
rlabel pdiffusion 857 -3080 857 -3080 0 feedthrough
rlabel pdiffusion 864 -3080 864 -3080 0 feedthrough
rlabel pdiffusion 871 -3080 871 -3080 0 feedthrough
rlabel pdiffusion 878 -3080 878 -3080 0 cellNo=621
rlabel pdiffusion 885 -3080 885 -3080 0 feedthrough
rlabel pdiffusion 892 -3080 892 -3080 0 feedthrough
rlabel pdiffusion 899 -3080 899 -3080 0 cellNo=922
rlabel pdiffusion 906 -3080 906 -3080 0 feedthrough
rlabel pdiffusion 913 -3080 913 -3080 0 cellNo=125
rlabel pdiffusion 920 -3080 920 -3080 0 feedthrough
rlabel pdiffusion 927 -3080 927 -3080 0 feedthrough
rlabel pdiffusion 934 -3080 934 -3080 0 feedthrough
rlabel pdiffusion 941 -3080 941 -3080 0 feedthrough
rlabel pdiffusion 948 -3080 948 -3080 0 cellNo=121
rlabel pdiffusion 955 -3080 955 -3080 0 feedthrough
rlabel pdiffusion 962 -3080 962 -3080 0 feedthrough
rlabel pdiffusion 969 -3080 969 -3080 0 feedthrough
rlabel pdiffusion 976 -3080 976 -3080 0 cellNo=403
rlabel pdiffusion 983 -3080 983 -3080 0 feedthrough
rlabel pdiffusion 990 -3080 990 -3080 0 feedthrough
rlabel pdiffusion 997 -3080 997 -3080 0 feedthrough
rlabel pdiffusion 1004 -3080 1004 -3080 0 feedthrough
rlabel pdiffusion 1011 -3080 1011 -3080 0 feedthrough
rlabel pdiffusion 1018 -3080 1018 -3080 0 cellNo=730
rlabel pdiffusion 1025 -3080 1025 -3080 0 feedthrough
rlabel pdiffusion 1032 -3080 1032 -3080 0 feedthrough
rlabel pdiffusion 1039 -3080 1039 -3080 0 feedthrough
rlabel pdiffusion 1046 -3080 1046 -3080 0 feedthrough
rlabel pdiffusion 1053 -3080 1053 -3080 0 feedthrough
rlabel pdiffusion 1060 -3080 1060 -3080 0 feedthrough
rlabel pdiffusion 1067 -3080 1067 -3080 0 feedthrough
rlabel pdiffusion 1074 -3080 1074 -3080 0 feedthrough
rlabel pdiffusion 1081 -3080 1081 -3080 0 cellNo=929
rlabel pdiffusion 1088 -3080 1088 -3080 0 cellNo=211
rlabel pdiffusion 1095 -3080 1095 -3080 0 feedthrough
rlabel pdiffusion 1102 -3080 1102 -3080 0 feedthrough
rlabel pdiffusion 1109 -3080 1109 -3080 0 feedthrough
rlabel pdiffusion 1116 -3080 1116 -3080 0 feedthrough
rlabel pdiffusion 1123 -3080 1123 -3080 0 feedthrough
rlabel pdiffusion 1130 -3080 1130 -3080 0 feedthrough
rlabel pdiffusion 1137 -3080 1137 -3080 0 feedthrough
rlabel pdiffusion 1144 -3080 1144 -3080 0 feedthrough
rlabel pdiffusion 1151 -3080 1151 -3080 0 feedthrough
rlabel pdiffusion 1158 -3080 1158 -3080 0 feedthrough
rlabel pdiffusion 1165 -3080 1165 -3080 0 feedthrough
rlabel pdiffusion 1172 -3080 1172 -3080 0 feedthrough
rlabel pdiffusion 1179 -3080 1179 -3080 0 feedthrough
rlabel pdiffusion 1186 -3080 1186 -3080 0 feedthrough
rlabel pdiffusion 1193 -3080 1193 -3080 0 feedthrough
rlabel pdiffusion 1200 -3080 1200 -3080 0 feedthrough
rlabel pdiffusion 1207 -3080 1207 -3080 0 feedthrough
rlabel pdiffusion 1214 -3080 1214 -3080 0 feedthrough
rlabel pdiffusion 1221 -3080 1221 -3080 0 feedthrough
rlabel pdiffusion 1228 -3080 1228 -3080 0 feedthrough
rlabel pdiffusion 1235 -3080 1235 -3080 0 feedthrough
rlabel pdiffusion 1242 -3080 1242 -3080 0 feedthrough
rlabel pdiffusion 1249 -3080 1249 -3080 0 feedthrough
rlabel pdiffusion 1256 -3080 1256 -3080 0 feedthrough
rlabel pdiffusion 1263 -3080 1263 -3080 0 feedthrough
rlabel pdiffusion 1270 -3080 1270 -3080 0 feedthrough
rlabel pdiffusion 1277 -3080 1277 -3080 0 feedthrough
rlabel pdiffusion 1284 -3080 1284 -3080 0 feedthrough
rlabel pdiffusion 1291 -3080 1291 -3080 0 feedthrough
rlabel pdiffusion 1298 -3080 1298 -3080 0 feedthrough
rlabel pdiffusion 1305 -3080 1305 -3080 0 feedthrough
rlabel pdiffusion 1312 -3080 1312 -3080 0 feedthrough
rlabel pdiffusion 1319 -3080 1319 -3080 0 feedthrough
rlabel pdiffusion 1326 -3080 1326 -3080 0 feedthrough
rlabel pdiffusion 1333 -3080 1333 -3080 0 feedthrough
rlabel pdiffusion 1340 -3080 1340 -3080 0 feedthrough
rlabel pdiffusion 1347 -3080 1347 -3080 0 feedthrough
rlabel pdiffusion 1354 -3080 1354 -3080 0 feedthrough
rlabel pdiffusion 1361 -3080 1361 -3080 0 feedthrough
rlabel pdiffusion 1368 -3080 1368 -3080 0 feedthrough
rlabel pdiffusion 1375 -3080 1375 -3080 0 feedthrough
rlabel pdiffusion 1382 -3080 1382 -3080 0 feedthrough
rlabel pdiffusion 1389 -3080 1389 -3080 0 feedthrough
rlabel pdiffusion 1396 -3080 1396 -3080 0 feedthrough
rlabel pdiffusion 1403 -3080 1403 -3080 0 feedthrough
rlabel pdiffusion 1410 -3080 1410 -3080 0 feedthrough
rlabel pdiffusion 1417 -3080 1417 -3080 0 feedthrough
rlabel pdiffusion 1424 -3080 1424 -3080 0 feedthrough
rlabel pdiffusion 1431 -3080 1431 -3080 0 feedthrough
rlabel pdiffusion 1438 -3080 1438 -3080 0 feedthrough
rlabel pdiffusion 1445 -3080 1445 -3080 0 feedthrough
rlabel pdiffusion 1452 -3080 1452 -3080 0 feedthrough
rlabel pdiffusion 1459 -3080 1459 -3080 0 feedthrough
rlabel pdiffusion 1466 -3080 1466 -3080 0 feedthrough
rlabel pdiffusion 1473 -3080 1473 -3080 0 feedthrough
rlabel pdiffusion 1480 -3080 1480 -3080 0 feedthrough
rlabel pdiffusion 1487 -3080 1487 -3080 0 feedthrough
rlabel pdiffusion 1494 -3080 1494 -3080 0 feedthrough
rlabel pdiffusion 1501 -3080 1501 -3080 0 feedthrough
rlabel pdiffusion 1508 -3080 1508 -3080 0 feedthrough
rlabel pdiffusion 1515 -3080 1515 -3080 0 feedthrough
rlabel pdiffusion 1522 -3080 1522 -3080 0 feedthrough
rlabel pdiffusion 1529 -3080 1529 -3080 0 feedthrough
rlabel pdiffusion 1536 -3080 1536 -3080 0 feedthrough
rlabel pdiffusion 1543 -3080 1543 -3080 0 feedthrough
rlabel pdiffusion 1550 -3080 1550 -3080 0 feedthrough
rlabel pdiffusion 1557 -3080 1557 -3080 0 feedthrough
rlabel pdiffusion 1564 -3080 1564 -3080 0 feedthrough
rlabel pdiffusion 1571 -3080 1571 -3080 0 feedthrough
rlabel pdiffusion 1578 -3080 1578 -3080 0 feedthrough
rlabel pdiffusion 1585 -3080 1585 -3080 0 feedthrough
rlabel pdiffusion 1592 -3080 1592 -3080 0 feedthrough
rlabel pdiffusion 1599 -3080 1599 -3080 0 feedthrough
rlabel pdiffusion 1606 -3080 1606 -3080 0 feedthrough
rlabel pdiffusion 1613 -3080 1613 -3080 0 feedthrough
rlabel pdiffusion 1620 -3080 1620 -3080 0 feedthrough
rlabel pdiffusion 1627 -3080 1627 -3080 0 feedthrough
rlabel pdiffusion 1634 -3080 1634 -3080 0 feedthrough
rlabel pdiffusion 1641 -3080 1641 -3080 0 feedthrough
rlabel pdiffusion 1648 -3080 1648 -3080 0 feedthrough
rlabel pdiffusion 1655 -3080 1655 -3080 0 feedthrough
rlabel pdiffusion 3 -3219 3 -3219 0 cellNo=1034
rlabel pdiffusion 10 -3219 10 -3219 0 cellNo=1045
rlabel pdiffusion 17 -3219 17 -3219 0 cellNo=1044
rlabel pdiffusion 24 -3219 24 -3219 0 cellNo=1048
rlabel pdiffusion 66 -3219 66 -3219 0 cellNo=671
rlabel pdiffusion 73 -3219 73 -3219 0 feedthrough
rlabel pdiffusion 80 -3219 80 -3219 0 feedthrough
rlabel pdiffusion 87 -3219 87 -3219 0 feedthrough
rlabel pdiffusion 94 -3219 94 -3219 0 feedthrough
rlabel pdiffusion 101 -3219 101 -3219 0 feedthrough
rlabel pdiffusion 108 -3219 108 -3219 0 feedthrough
rlabel pdiffusion 115 -3219 115 -3219 0 cellNo=409
rlabel pdiffusion 122 -3219 122 -3219 0 feedthrough
rlabel pdiffusion 129 -3219 129 -3219 0 cellNo=131
rlabel pdiffusion 136 -3219 136 -3219 0 feedthrough
rlabel pdiffusion 143 -3219 143 -3219 0 feedthrough
rlabel pdiffusion 150 -3219 150 -3219 0 cellNo=44
rlabel pdiffusion 157 -3219 157 -3219 0 feedthrough
rlabel pdiffusion 164 -3219 164 -3219 0 feedthrough
rlabel pdiffusion 171 -3219 171 -3219 0 feedthrough
rlabel pdiffusion 178 -3219 178 -3219 0 feedthrough
rlabel pdiffusion 185 -3219 185 -3219 0 feedthrough
rlabel pdiffusion 192 -3219 192 -3219 0 feedthrough
rlabel pdiffusion 199 -3219 199 -3219 0 feedthrough
rlabel pdiffusion 206 -3219 206 -3219 0 feedthrough
rlabel pdiffusion 213 -3219 213 -3219 0 feedthrough
rlabel pdiffusion 220 -3219 220 -3219 0 feedthrough
rlabel pdiffusion 227 -3219 227 -3219 0 feedthrough
rlabel pdiffusion 234 -3219 234 -3219 0 feedthrough
rlabel pdiffusion 241 -3219 241 -3219 0 cellNo=17
rlabel pdiffusion 248 -3219 248 -3219 0 feedthrough
rlabel pdiffusion 255 -3219 255 -3219 0 feedthrough
rlabel pdiffusion 262 -3219 262 -3219 0 feedthrough
rlabel pdiffusion 269 -3219 269 -3219 0 feedthrough
rlabel pdiffusion 276 -3219 276 -3219 0 feedthrough
rlabel pdiffusion 283 -3219 283 -3219 0 feedthrough
rlabel pdiffusion 290 -3219 290 -3219 0 feedthrough
rlabel pdiffusion 297 -3219 297 -3219 0 feedthrough
rlabel pdiffusion 304 -3219 304 -3219 0 feedthrough
rlabel pdiffusion 311 -3219 311 -3219 0 feedthrough
rlabel pdiffusion 318 -3219 318 -3219 0 feedthrough
rlabel pdiffusion 325 -3219 325 -3219 0 feedthrough
rlabel pdiffusion 332 -3219 332 -3219 0 feedthrough
rlabel pdiffusion 339 -3219 339 -3219 0 feedthrough
rlabel pdiffusion 346 -3219 346 -3219 0 feedthrough
rlabel pdiffusion 353 -3219 353 -3219 0 feedthrough
rlabel pdiffusion 360 -3219 360 -3219 0 feedthrough
rlabel pdiffusion 367 -3219 367 -3219 0 feedthrough
rlabel pdiffusion 374 -3219 374 -3219 0 feedthrough
rlabel pdiffusion 381 -3219 381 -3219 0 feedthrough
rlabel pdiffusion 388 -3219 388 -3219 0 feedthrough
rlabel pdiffusion 395 -3219 395 -3219 0 feedthrough
rlabel pdiffusion 402 -3219 402 -3219 0 cellNo=188
rlabel pdiffusion 409 -3219 409 -3219 0 feedthrough
rlabel pdiffusion 416 -3219 416 -3219 0 feedthrough
rlabel pdiffusion 423 -3219 423 -3219 0 feedthrough
rlabel pdiffusion 430 -3219 430 -3219 0 cellNo=462
rlabel pdiffusion 437 -3219 437 -3219 0 feedthrough
rlabel pdiffusion 444 -3219 444 -3219 0 feedthrough
rlabel pdiffusion 451 -3219 451 -3219 0 feedthrough
rlabel pdiffusion 458 -3219 458 -3219 0 feedthrough
rlabel pdiffusion 465 -3219 465 -3219 0 feedthrough
rlabel pdiffusion 472 -3219 472 -3219 0 cellNo=701
rlabel pdiffusion 479 -3219 479 -3219 0 feedthrough
rlabel pdiffusion 486 -3219 486 -3219 0 feedthrough
rlabel pdiffusion 493 -3219 493 -3219 0 cellNo=615
rlabel pdiffusion 500 -3219 500 -3219 0 cellNo=722
rlabel pdiffusion 507 -3219 507 -3219 0 feedthrough
rlabel pdiffusion 514 -3219 514 -3219 0 feedthrough
rlabel pdiffusion 521 -3219 521 -3219 0 feedthrough
rlabel pdiffusion 528 -3219 528 -3219 0 feedthrough
rlabel pdiffusion 535 -3219 535 -3219 0 cellNo=947
rlabel pdiffusion 542 -3219 542 -3219 0 cellNo=855
rlabel pdiffusion 549 -3219 549 -3219 0 feedthrough
rlabel pdiffusion 556 -3219 556 -3219 0 feedthrough
rlabel pdiffusion 563 -3219 563 -3219 0 feedthrough
rlabel pdiffusion 570 -3219 570 -3219 0 feedthrough
rlabel pdiffusion 577 -3219 577 -3219 0 cellNo=944
rlabel pdiffusion 584 -3219 584 -3219 0 feedthrough
rlabel pdiffusion 591 -3219 591 -3219 0 cellNo=648
rlabel pdiffusion 598 -3219 598 -3219 0 feedthrough
rlabel pdiffusion 605 -3219 605 -3219 0 feedthrough
rlabel pdiffusion 612 -3219 612 -3219 0 feedthrough
rlabel pdiffusion 619 -3219 619 -3219 0 feedthrough
rlabel pdiffusion 626 -3219 626 -3219 0 feedthrough
rlabel pdiffusion 633 -3219 633 -3219 0 feedthrough
rlabel pdiffusion 640 -3219 640 -3219 0 feedthrough
rlabel pdiffusion 647 -3219 647 -3219 0 feedthrough
rlabel pdiffusion 654 -3219 654 -3219 0 cellNo=897
rlabel pdiffusion 661 -3219 661 -3219 0 feedthrough
rlabel pdiffusion 668 -3219 668 -3219 0 feedthrough
rlabel pdiffusion 675 -3219 675 -3219 0 feedthrough
rlabel pdiffusion 682 -3219 682 -3219 0 cellNo=4
rlabel pdiffusion 689 -3219 689 -3219 0 feedthrough
rlabel pdiffusion 696 -3219 696 -3219 0 feedthrough
rlabel pdiffusion 703 -3219 703 -3219 0 feedthrough
rlabel pdiffusion 710 -3219 710 -3219 0 feedthrough
rlabel pdiffusion 717 -3219 717 -3219 0 feedthrough
rlabel pdiffusion 724 -3219 724 -3219 0 feedthrough
rlabel pdiffusion 731 -3219 731 -3219 0 feedthrough
rlabel pdiffusion 738 -3219 738 -3219 0 feedthrough
rlabel pdiffusion 745 -3219 745 -3219 0 feedthrough
rlabel pdiffusion 752 -3219 752 -3219 0 feedthrough
rlabel pdiffusion 759 -3219 759 -3219 0 feedthrough
rlabel pdiffusion 766 -3219 766 -3219 0 feedthrough
rlabel pdiffusion 773 -3219 773 -3219 0 feedthrough
rlabel pdiffusion 780 -3219 780 -3219 0 cellNo=803
rlabel pdiffusion 787 -3219 787 -3219 0 feedthrough
rlabel pdiffusion 794 -3219 794 -3219 0 cellNo=776
rlabel pdiffusion 801 -3219 801 -3219 0 feedthrough
rlabel pdiffusion 808 -3219 808 -3219 0 feedthrough
rlabel pdiffusion 815 -3219 815 -3219 0 feedthrough
rlabel pdiffusion 822 -3219 822 -3219 0 cellNo=734
rlabel pdiffusion 829 -3219 829 -3219 0 feedthrough
rlabel pdiffusion 836 -3219 836 -3219 0 cellNo=936
rlabel pdiffusion 843 -3219 843 -3219 0 feedthrough
rlabel pdiffusion 850 -3219 850 -3219 0 feedthrough
rlabel pdiffusion 857 -3219 857 -3219 0 feedthrough
rlabel pdiffusion 864 -3219 864 -3219 0 feedthrough
rlabel pdiffusion 871 -3219 871 -3219 0 feedthrough
rlabel pdiffusion 878 -3219 878 -3219 0 feedthrough
rlabel pdiffusion 885 -3219 885 -3219 0 feedthrough
rlabel pdiffusion 892 -3219 892 -3219 0 cellNo=711
rlabel pdiffusion 899 -3219 899 -3219 0 feedthrough
rlabel pdiffusion 906 -3219 906 -3219 0 feedthrough
rlabel pdiffusion 913 -3219 913 -3219 0 feedthrough
rlabel pdiffusion 920 -3219 920 -3219 0 feedthrough
rlabel pdiffusion 927 -3219 927 -3219 0 feedthrough
rlabel pdiffusion 934 -3219 934 -3219 0 feedthrough
rlabel pdiffusion 941 -3219 941 -3219 0 feedthrough
rlabel pdiffusion 948 -3219 948 -3219 0 cellNo=325
rlabel pdiffusion 955 -3219 955 -3219 0 feedthrough
rlabel pdiffusion 962 -3219 962 -3219 0 feedthrough
rlabel pdiffusion 969 -3219 969 -3219 0 feedthrough
rlabel pdiffusion 976 -3219 976 -3219 0 feedthrough
rlabel pdiffusion 983 -3219 983 -3219 0 feedthrough
rlabel pdiffusion 990 -3219 990 -3219 0 feedthrough
rlabel pdiffusion 997 -3219 997 -3219 0 cellNo=640
rlabel pdiffusion 1004 -3219 1004 -3219 0 feedthrough
rlabel pdiffusion 1011 -3219 1011 -3219 0 cellNo=907
rlabel pdiffusion 1018 -3219 1018 -3219 0 feedthrough
rlabel pdiffusion 1025 -3219 1025 -3219 0 feedthrough
rlabel pdiffusion 1032 -3219 1032 -3219 0 feedthrough
rlabel pdiffusion 1039 -3219 1039 -3219 0 feedthrough
rlabel pdiffusion 1046 -3219 1046 -3219 0 feedthrough
rlabel pdiffusion 1053 -3219 1053 -3219 0 feedthrough
rlabel pdiffusion 1060 -3219 1060 -3219 0 cellNo=123
rlabel pdiffusion 1067 -3219 1067 -3219 0 feedthrough
rlabel pdiffusion 1074 -3219 1074 -3219 0 feedthrough
rlabel pdiffusion 1081 -3219 1081 -3219 0 feedthrough
rlabel pdiffusion 1088 -3219 1088 -3219 0 cellNo=997
rlabel pdiffusion 1095 -3219 1095 -3219 0 feedthrough
rlabel pdiffusion 1102 -3219 1102 -3219 0 feedthrough
rlabel pdiffusion 1109 -3219 1109 -3219 0 feedthrough
rlabel pdiffusion 1116 -3219 1116 -3219 0 feedthrough
rlabel pdiffusion 1123 -3219 1123 -3219 0 feedthrough
rlabel pdiffusion 1130 -3219 1130 -3219 0 feedthrough
rlabel pdiffusion 1137 -3219 1137 -3219 0 feedthrough
rlabel pdiffusion 1144 -3219 1144 -3219 0 feedthrough
rlabel pdiffusion 1151 -3219 1151 -3219 0 feedthrough
rlabel pdiffusion 1158 -3219 1158 -3219 0 feedthrough
rlabel pdiffusion 1165 -3219 1165 -3219 0 feedthrough
rlabel pdiffusion 1172 -3219 1172 -3219 0 feedthrough
rlabel pdiffusion 1179 -3219 1179 -3219 0 feedthrough
rlabel pdiffusion 1186 -3219 1186 -3219 0 feedthrough
rlabel pdiffusion 1193 -3219 1193 -3219 0 feedthrough
rlabel pdiffusion 1200 -3219 1200 -3219 0 feedthrough
rlabel pdiffusion 1207 -3219 1207 -3219 0 feedthrough
rlabel pdiffusion 1214 -3219 1214 -3219 0 feedthrough
rlabel pdiffusion 1221 -3219 1221 -3219 0 feedthrough
rlabel pdiffusion 1228 -3219 1228 -3219 0 feedthrough
rlabel pdiffusion 1235 -3219 1235 -3219 0 feedthrough
rlabel pdiffusion 1242 -3219 1242 -3219 0 feedthrough
rlabel pdiffusion 1249 -3219 1249 -3219 0 feedthrough
rlabel pdiffusion 1256 -3219 1256 -3219 0 feedthrough
rlabel pdiffusion 1263 -3219 1263 -3219 0 feedthrough
rlabel pdiffusion 1270 -3219 1270 -3219 0 feedthrough
rlabel pdiffusion 1277 -3219 1277 -3219 0 feedthrough
rlabel pdiffusion 1284 -3219 1284 -3219 0 feedthrough
rlabel pdiffusion 1291 -3219 1291 -3219 0 feedthrough
rlabel pdiffusion 1298 -3219 1298 -3219 0 cellNo=668
rlabel pdiffusion 1305 -3219 1305 -3219 0 feedthrough
rlabel pdiffusion 1312 -3219 1312 -3219 0 feedthrough
rlabel pdiffusion 1319 -3219 1319 -3219 0 feedthrough
rlabel pdiffusion 1326 -3219 1326 -3219 0 feedthrough
rlabel pdiffusion 1333 -3219 1333 -3219 0 feedthrough
rlabel pdiffusion 1340 -3219 1340 -3219 0 feedthrough
rlabel pdiffusion 1347 -3219 1347 -3219 0 cellNo=805
rlabel pdiffusion 1354 -3219 1354 -3219 0 cellNo=790
rlabel pdiffusion 1361 -3219 1361 -3219 0 feedthrough
rlabel pdiffusion 1368 -3219 1368 -3219 0 feedthrough
rlabel pdiffusion 1375 -3219 1375 -3219 0 feedthrough
rlabel pdiffusion 1382 -3219 1382 -3219 0 feedthrough
rlabel pdiffusion 1389 -3219 1389 -3219 0 feedthrough
rlabel pdiffusion 1396 -3219 1396 -3219 0 feedthrough
rlabel pdiffusion 1403 -3219 1403 -3219 0 feedthrough
rlabel pdiffusion 1410 -3219 1410 -3219 0 cellNo=350
rlabel pdiffusion 1417 -3219 1417 -3219 0 feedthrough
rlabel pdiffusion 1424 -3219 1424 -3219 0 feedthrough
rlabel pdiffusion 1431 -3219 1431 -3219 0 feedthrough
rlabel pdiffusion 1438 -3219 1438 -3219 0 feedthrough
rlabel pdiffusion 1445 -3219 1445 -3219 0 feedthrough
rlabel pdiffusion 1452 -3219 1452 -3219 0 feedthrough
rlabel pdiffusion 1459 -3219 1459 -3219 0 feedthrough
rlabel pdiffusion 1466 -3219 1466 -3219 0 feedthrough
rlabel pdiffusion 1473 -3219 1473 -3219 0 cellNo=238
rlabel pdiffusion 1480 -3219 1480 -3219 0 feedthrough
rlabel pdiffusion 1487 -3219 1487 -3219 0 feedthrough
rlabel pdiffusion 1494 -3219 1494 -3219 0 feedthrough
rlabel pdiffusion 1501 -3219 1501 -3219 0 feedthrough
rlabel pdiffusion 1508 -3219 1508 -3219 0 feedthrough
rlabel pdiffusion 1515 -3219 1515 -3219 0 feedthrough
rlabel pdiffusion 1522 -3219 1522 -3219 0 feedthrough
rlabel pdiffusion 1606 -3219 1606 -3219 0 feedthrough
rlabel pdiffusion 3 -3312 3 -3312 0 cellNo=1037
rlabel pdiffusion 10 -3312 10 -3312 0 cellNo=1042
rlabel pdiffusion 17 -3312 17 -3312 0 cellNo=1098
rlabel pdiffusion 24 -3312 24 -3312 0 cellNo=1054
rlabel pdiffusion 129 -3312 129 -3312 0 cellNo=703
rlabel pdiffusion 136 -3312 136 -3312 0 feedthrough
rlabel pdiffusion 164 -3312 164 -3312 0 feedthrough
rlabel pdiffusion 171 -3312 171 -3312 0 feedthrough
rlabel pdiffusion 178 -3312 178 -3312 0 feedthrough
rlabel pdiffusion 185 -3312 185 -3312 0 feedthrough
rlabel pdiffusion 192 -3312 192 -3312 0 feedthrough
rlabel pdiffusion 199 -3312 199 -3312 0 feedthrough
rlabel pdiffusion 206 -3312 206 -3312 0 feedthrough
rlabel pdiffusion 213 -3312 213 -3312 0 feedthrough
rlabel pdiffusion 220 -3312 220 -3312 0 feedthrough
rlabel pdiffusion 227 -3312 227 -3312 0 feedthrough
rlabel pdiffusion 234 -3312 234 -3312 0 feedthrough
rlabel pdiffusion 241 -3312 241 -3312 0 feedthrough
rlabel pdiffusion 248 -3312 248 -3312 0 feedthrough
rlabel pdiffusion 255 -3312 255 -3312 0 feedthrough
rlabel pdiffusion 262 -3312 262 -3312 0 feedthrough
rlabel pdiffusion 269 -3312 269 -3312 0 feedthrough
rlabel pdiffusion 276 -3312 276 -3312 0 feedthrough
rlabel pdiffusion 283 -3312 283 -3312 0 feedthrough
rlabel pdiffusion 290 -3312 290 -3312 0 feedthrough
rlabel pdiffusion 297 -3312 297 -3312 0 feedthrough
rlabel pdiffusion 304 -3312 304 -3312 0 feedthrough
rlabel pdiffusion 311 -3312 311 -3312 0 feedthrough
rlabel pdiffusion 318 -3312 318 -3312 0 feedthrough
rlabel pdiffusion 325 -3312 325 -3312 0 feedthrough
rlabel pdiffusion 332 -3312 332 -3312 0 feedthrough
rlabel pdiffusion 339 -3312 339 -3312 0 feedthrough
rlabel pdiffusion 346 -3312 346 -3312 0 cellNo=617
rlabel pdiffusion 353 -3312 353 -3312 0 feedthrough
rlabel pdiffusion 360 -3312 360 -3312 0 feedthrough
rlabel pdiffusion 367 -3312 367 -3312 0 feedthrough
rlabel pdiffusion 374 -3312 374 -3312 0 feedthrough
rlabel pdiffusion 381 -3312 381 -3312 0 feedthrough
rlabel pdiffusion 388 -3312 388 -3312 0 feedthrough
rlabel pdiffusion 395 -3312 395 -3312 0 feedthrough
rlabel pdiffusion 402 -3312 402 -3312 0 cellNo=58
rlabel pdiffusion 409 -3312 409 -3312 0 feedthrough
rlabel pdiffusion 416 -3312 416 -3312 0 feedthrough
rlabel pdiffusion 423 -3312 423 -3312 0 feedthrough
rlabel pdiffusion 430 -3312 430 -3312 0 feedthrough
rlabel pdiffusion 437 -3312 437 -3312 0 cellNo=29
rlabel pdiffusion 444 -3312 444 -3312 0 cellNo=914
rlabel pdiffusion 451 -3312 451 -3312 0 feedthrough
rlabel pdiffusion 458 -3312 458 -3312 0 feedthrough
rlabel pdiffusion 465 -3312 465 -3312 0 feedthrough
rlabel pdiffusion 472 -3312 472 -3312 0 feedthrough
rlabel pdiffusion 479 -3312 479 -3312 0 feedthrough
rlabel pdiffusion 486 -3312 486 -3312 0 feedthrough
rlabel pdiffusion 493 -3312 493 -3312 0 cellNo=662
rlabel pdiffusion 500 -3312 500 -3312 0 feedthrough
rlabel pdiffusion 507 -3312 507 -3312 0 feedthrough
rlabel pdiffusion 514 -3312 514 -3312 0 feedthrough
rlabel pdiffusion 521 -3312 521 -3312 0 feedthrough
rlabel pdiffusion 528 -3312 528 -3312 0 cellNo=445
rlabel pdiffusion 535 -3312 535 -3312 0 feedthrough
rlabel pdiffusion 542 -3312 542 -3312 0 cellNo=752
rlabel pdiffusion 549 -3312 549 -3312 0 feedthrough
rlabel pdiffusion 556 -3312 556 -3312 0 feedthrough
rlabel pdiffusion 563 -3312 563 -3312 0 feedthrough
rlabel pdiffusion 570 -3312 570 -3312 0 feedthrough
rlabel pdiffusion 577 -3312 577 -3312 0 feedthrough
rlabel pdiffusion 584 -3312 584 -3312 0 feedthrough
rlabel pdiffusion 591 -3312 591 -3312 0 feedthrough
rlabel pdiffusion 598 -3312 598 -3312 0 feedthrough
rlabel pdiffusion 605 -3312 605 -3312 0 feedthrough
rlabel pdiffusion 612 -3312 612 -3312 0 feedthrough
rlabel pdiffusion 619 -3312 619 -3312 0 cellNo=843
rlabel pdiffusion 626 -3312 626 -3312 0 feedthrough
rlabel pdiffusion 633 -3312 633 -3312 0 feedthrough
rlabel pdiffusion 640 -3312 640 -3312 0 feedthrough
rlabel pdiffusion 647 -3312 647 -3312 0 feedthrough
rlabel pdiffusion 654 -3312 654 -3312 0 feedthrough
rlabel pdiffusion 661 -3312 661 -3312 0 feedthrough
rlabel pdiffusion 668 -3312 668 -3312 0 feedthrough
rlabel pdiffusion 675 -3312 675 -3312 0 cellNo=68
rlabel pdiffusion 682 -3312 682 -3312 0 feedthrough
rlabel pdiffusion 689 -3312 689 -3312 0 cellNo=986
rlabel pdiffusion 696 -3312 696 -3312 0 feedthrough
rlabel pdiffusion 703 -3312 703 -3312 0 cellNo=226
rlabel pdiffusion 710 -3312 710 -3312 0 feedthrough
rlabel pdiffusion 717 -3312 717 -3312 0 feedthrough
rlabel pdiffusion 724 -3312 724 -3312 0 feedthrough
rlabel pdiffusion 731 -3312 731 -3312 0 feedthrough
rlabel pdiffusion 738 -3312 738 -3312 0 feedthrough
rlabel pdiffusion 745 -3312 745 -3312 0 feedthrough
rlabel pdiffusion 752 -3312 752 -3312 0 feedthrough
rlabel pdiffusion 759 -3312 759 -3312 0 feedthrough
rlabel pdiffusion 766 -3312 766 -3312 0 feedthrough
rlabel pdiffusion 773 -3312 773 -3312 0 feedthrough
rlabel pdiffusion 780 -3312 780 -3312 0 feedthrough
rlabel pdiffusion 787 -3312 787 -3312 0 cellNo=457
rlabel pdiffusion 794 -3312 794 -3312 0 feedthrough
rlabel pdiffusion 801 -3312 801 -3312 0 feedthrough
rlabel pdiffusion 808 -3312 808 -3312 0 feedthrough
rlabel pdiffusion 815 -3312 815 -3312 0 feedthrough
rlabel pdiffusion 822 -3312 822 -3312 0 feedthrough
rlabel pdiffusion 829 -3312 829 -3312 0 feedthrough
rlabel pdiffusion 836 -3312 836 -3312 0 feedthrough
rlabel pdiffusion 843 -3312 843 -3312 0 feedthrough
rlabel pdiffusion 850 -3312 850 -3312 0 feedthrough
rlabel pdiffusion 857 -3312 857 -3312 0 feedthrough
rlabel pdiffusion 864 -3312 864 -3312 0 feedthrough
rlabel pdiffusion 871 -3312 871 -3312 0 cellNo=535
rlabel pdiffusion 878 -3312 878 -3312 0 cellNo=456
rlabel pdiffusion 885 -3312 885 -3312 0 feedthrough
rlabel pdiffusion 892 -3312 892 -3312 0 feedthrough
rlabel pdiffusion 899 -3312 899 -3312 0 cellNo=757
rlabel pdiffusion 906 -3312 906 -3312 0 cellNo=594
rlabel pdiffusion 913 -3312 913 -3312 0 cellNo=676
rlabel pdiffusion 920 -3312 920 -3312 0 feedthrough
rlabel pdiffusion 927 -3312 927 -3312 0 feedthrough
rlabel pdiffusion 934 -3312 934 -3312 0 feedthrough
rlabel pdiffusion 941 -3312 941 -3312 0 feedthrough
rlabel pdiffusion 948 -3312 948 -3312 0 feedthrough
rlabel pdiffusion 955 -3312 955 -3312 0 feedthrough
rlabel pdiffusion 962 -3312 962 -3312 0 feedthrough
rlabel pdiffusion 969 -3312 969 -3312 0 feedthrough
rlabel pdiffusion 976 -3312 976 -3312 0 feedthrough
rlabel pdiffusion 983 -3312 983 -3312 0 cellNo=241
rlabel pdiffusion 990 -3312 990 -3312 0 feedthrough
rlabel pdiffusion 997 -3312 997 -3312 0 feedthrough
rlabel pdiffusion 1004 -3312 1004 -3312 0 feedthrough
rlabel pdiffusion 1011 -3312 1011 -3312 0 feedthrough
rlabel pdiffusion 1018 -3312 1018 -3312 0 cellNo=207
rlabel pdiffusion 1025 -3312 1025 -3312 0 feedthrough
rlabel pdiffusion 1032 -3312 1032 -3312 0 feedthrough
rlabel pdiffusion 1039 -3312 1039 -3312 0 feedthrough
rlabel pdiffusion 1046 -3312 1046 -3312 0 feedthrough
rlabel pdiffusion 1053 -3312 1053 -3312 0 feedthrough
rlabel pdiffusion 1060 -3312 1060 -3312 0 feedthrough
rlabel pdiffusion 1067 -3312 1067 -3312 0 feedthrough
rlabel pdiffusion 1074 -3312 1074 -3312 0 feedthrough
rlabel pdiffusion 1081 -3312 1081 -3312 0 feedthrough
rlabel pdiffusion 1088 -3312 1088 -3312 0 feedthrough
rlabel pdiffusion 1095 -3312 1095 -3312 0 feedthrough
rlabel pdiffusion 1102 -3312 1102 -3312 0 feedthrough
rlabel pdiffusion 1109 -3312 1109 -3312 0 cellNo=967
rlabel pdiffusion 1116 -3312 1116 -3312 0 feedthrough
rlabel pdiffusion 1123 -3312 1123 -3312 0 feedthrough
rlabel pdiffusion 1130 -3312 1130 -3312 0 cellNo=709
rlabel pdiffusion 1137 -3312 1137 -3312 0 feedthrough
rlabel pdiffusion 1144 -3312 1144 -3312 0 feedthrough
rlabel pdiffusion 1151 -3312 1151 -3312 0 feedthrough
rlabel pdiffusion 1158 -3312 1158 -3312 0 feedthrough
rlabel pdiffusion 1165 -3312 1165 -3312 0 feedthrough
rlabel pdiffusion 1172 -3312 1172 -3312 0 feedthrough
rlabel pdiffusion 1179 -3312 1179 -3312 0 cellNo=176
rlabel pdiffusion 1186 -3312 1186 -3312 0 cellNo=689
rlabel pdiffusion 1193 -3312 1193 -3312 0 feedthrough
rlabel pdiffusion 1200 -3312 1200 -3312 0 feedthrough
rlabel pdiffusion 1207 -3312 1207 -3312 0 cellNo=871
rlabel pdiffusion 1214 -3312 1214 -3312 0 cellNo=665
rlabel pdiffusion 1221 -3312 1221 -3312 0 feedthrough
rlabel pdiffusion 1228 -3312 1228 -3312 0 feedthrough
rlabel pdiffusion 1235 -3312 1235 -3312 0 feedthrough
rlabel pdiffusion 1242 -3312 1242 -3312 0 feedthrough
rlabel pdiffusion 1249 -3312 1249 -3312 0 cellNo=511
rlabel pdiffusion 1256 -3312 1256 -3312 0 cellNo=394
rlabel pdiffusion 1263 -3312 1263 -3312 0 cellNo=78
rlabel pdiffusion 1270 -3312 1270 -3312 0 feedthrough
rlabel pdiffusion 1277 -3312 1277 -3312 0 feedthrough
rlabel pdiffusion 1284 -3312 1284 -3312 0 feedthrough
rlabel pdiffusion 1291 -3312 1291 -3312 0 feedthrough
rlabel pdiffusion 1298 -3312 1298 -3312 0 feedthrough
rlabel pdiffusion 1305 -3312 1305 -3312 0 feedthrough
rlabel pdiffusion 1312 -3312 1312 -3312 0 feedthrough
rlabel pdiffusion 1319 -3312 1319 -3312 0 feedthrough
rlabel pdiffusion 1326 -3312 1326 -3312 0 feedthrough
rlabel pdiffusion 1333 -3312 1333 -3312 0 feedthrough
rlabel pdiffusion 1340 -3312 1340 -3312 0 feedthrough
rlabel pdiffusion 1347 -3312 1347 -3312 0 feedthrough
rlabel pdiffusion 1354 -3312 1354 -3312 0 feedthrough
rlabel pdiffusion 1361 -3312 1361 -3312 0 feedthrough
rlabel pdiffusion 1382 -3312 1382 -3312 0 feedthrough
rlabel pdiffusion 1389 -3312 1389 -3312 0 feedthrough
rlabel pdiffusion 1529 -3312 1529 -3312 0 cellNo=442
rlabel pdiffusion 1585 -3312 1585 -3312 0 feedthrough
rlabel pdiffusion 3 -3409 3 -3409 0 cellNo=1041
rlabel pdiffusion 10 -3409 10 -3409 0 cellNo=1047
rlabel pdiffusion 17 -3409 17 -3409 0 cellNo=1053
rlabel pdiffusion 24 -3409 24 -3409 0 cellNo=1057
rlabel pdiffusion 31 -3409 31 -3409 0 cellNo=1060
rlabel pdiffusion 38 -3409 38 -3409 0 cellNo=1067
rlabel pdiffusion 45 -3409 45 -3409 0 cellNo=1076
rlabel pdiffusion 52 -3409 52 -3409 0 cellNo=1095
rlabel pdiffusion 59 -3409 59 -3409 0 cellNo=1108
rlabel pdiffusion 241 -3409 241 -3409 0 feedthrough
rlabel pdiffusion 248 -3409 248 -3409 0 feedthrough
rlabel pdiffusion 269 -3409 269 -3409 0 feedthrough
rlabel pdiffusion 283 -3409 283 -3409 0 feedthrough
rlabel pdiffusion 290 -3409 290 -3409 0 cellNo=655
rlabel pdiffusion 297 -3409 297 -3409 0 cellNo=145
rlabel pdiffusion 304 -3409 304 -3409 0 feedthrough
rlabel pdiffusion 311 -3409 311 -3409 0 feedthrough
rlabel pdiffusion 318 -3409 318 -3409 0 feedthrough
rlabel pdiffusion 325 -3409 325 -3409 0 feedthrough
rlabel pdiffusion 332 -3409 332 -3409 0 feedthrough
rlabel pdiffusion 339 -3409 339 -3409 0 feedthrough
rlabel pdiffusion 346 -3409 346 -3409 0 feedthrough
rlabel pdiffusion 353 -3409 353 -3409 0 feedthrough
rlabel pdiffusion 360 -3409 360 -3409 0 feedthrough
rlabel pdiffusion 367 -3409 367 -3409 0 feedthrough
rlabel pdiffusion 374 -3409 374 -3409 0 cellNo=875
rlabel pdiffusion 381 -3409 381 -3409 0 feedthrough
rlabel pdiffusion 388 -3409 388 -3409 0 feedthrough
rlabel pdiffusion 395 -3409 395 -3409 0 feedthrough
rlabel pdiffusion 402 -3409 402 -3409 0 feedthrough
rlabel pdiffusion 409 -3409 409 -3409 0 feedthrough
rlabel pdiffusion 416 -3409 416 -3409 0 feedthrough
rlabel pdiffusion 423 -3409 423 -3409 0 feedthrough
rlabel pdiffusion 430 -3409 430 -3409 0 feedthrough
rlabel pdiffusion 437 -3409 437 -3409 0 feedthrough
rlabel pdiffusion 444 -3409 444 -3409 0 feedthrough
rlabel pdiffusion 451 -3409 451 -3409 0 feedthrough
rlabel pdiffusion 458 -3409 458 -3409 0 feedthrough
rlabel pdiffusion 465 -3409 465 -3409 0 feedthrough
rlabel pdiffusion 472 -3409 472 -3409 0 feedthrough
rlabel pdiffusion 479 -3409 479 -3409 0 feedthrough
rlabel pdiffusion 486 -3409 486 -3409 0 feedthrough
rlabel pdiffusion 493 -3409 493 -3409 0 feedthrough
rlabel pdiffusion 500 -3409 500 -3409 0 cellNo=531
rlabel pdiffusion 507 -3409 507 -3409 0 feedthrough
rlabel pdiffusion 514 -3409 514 -3409 0 feedthrough
rlabel pdiffusion 521 -3409 521 -3409 0 cellNo=687
rlabel pdiffusion 528 -3409 528 -3409 0 feedthrough
rlabel pdiffusion 535 -3409 535 -3409 0 feedthrough
rlabel pdiffusion 542 -3409 542 -3409 0 feedthrough
rlabel pdiffusion 549 -3409 549 -3409 0 feedthrough
rlabel pdiffusion 556 -3409 556 -3409 0 feedthrough
rlabel pdiffusion 563 -3409 563 -3409 0 feedthrough
rlabel pdiffusion 570 -3409 570 -3409 0 feedthrough
rlabel pdiffusion 577 -3409 577 -3409 0 cellNo=797
rlabel pdiffusion 584 -3409 584 -3409 0 feedthrough
rlabel pdiffusion 591 -3409 591 -3409 0 feedthrough
rlabel pdiffusion 598 -3409 598 -3409 0 feedthrough
rlabel pdiffusion 605 -3409 605 -3409 0 feedthrough
rlabel pdiffusion 612 -3409 612 -3409 0 cellNo=192
rlabel pdiffusion 619 -3409 619 -3409 0 feedthrough
rlabel pdiffusion 626 -3409 626 -3409 0 feedthrough
rlabel pdiffusion 633 -3409 633 -3409 0 feedthrough
rlabel pdiffusion 640 -3409 640 -3409 0 feedthrough
rlabel pdiffusion 647 -3409 647 -3409 0 feedthrough
rlabel pdiffusion 654 -3409 654 -3409 0 feedthrough
rlabel pdiffusion 661 -3409 661 -3409 0 feedthrough
rlabel pdiffusion 668 -3409 668 -3409 0 feedthrough
rlabel pdiffusion 675 -3409 675 -3409 0 feedthrough
rlabel pdiffusion 682 -3409 682 -3409 0 feedthrough
rlabel pdiffusion 689 -3409 689 -3409 0 feedthrough
rlabel pdiffusion 696 -3409 696 -3409 0 feedthrough
rlabel pdiffusion 703 -3409 703 -3409 0 feedthrough
rlabel pdiffusion 710 -3409 710 -3409 0 feedthrough
rlabel pdiffusion 717 -3409 717 -3409 0 feedthrough
rlabel pdiffusion 724 -3409 724 -3409 0 feedthrough
rlabel pdiffusion 731 -3409 731 -3409 0 cellNo=630
rlabel pdiffusion 738 -3409 738 -3409 0 feedthrough
rlabel pdiffusion 745 -3409 745 -3409 0 feedthrough
rlabel pdiffusion 752 -3409 752 -3409 0 feedthrough
rlabel pdiffusion 759 -3409 759 -3409 0 feedthrough
rlabel pdiffusion 766 -3409 766 -3409 0 feedthrough
rlabel pdiffusion 773 -3409 773 -3409 0 feedthrough
rlabel pdiffusion 780 -3409 780 -3409 0 feedthrough
rlabel pdiffusion 787 -3409 787 -3409 0 feedthrough
rlabel pdiffusion 794 -3409 794 -3409 0 feedthrough
rlabel pdiffusion 801 -3409 801 -3409 0 cellNo=748
rlabel pdiffusion 808 -3409 808 -3409 0 feedthrough
rlabel pdiffusion 815 -3409 815 -3409 0 feedthrough
rlabel pdiffusion 822 -3409 822 -3409 0 feedthrough
rlabel pdiffusion 829 -3409 829 -3409 0 feedthrough
rlabel pdiffusion 836 -3409 836 -3409 0 feedthrough
rlabel pdiffusion 843 -3409 843 -3409 0 feedthrough
rlabel pdiffusion 850 -3409 850 -3409 0 feedthrough
rlabel pdiffusion 857 -3409 857 -3409 0 feedthrough
rlabel pdiffusion 864 -3409 864 -3409 0 feedthrough
rlabel pdiffusion 871 -3409 871 -3409 0 feedthrough
rlabel pdiffusion 878 -3409 878 -3409 0 cellNo=221
rlabel pdiffusion 885 -3409 885 -3409 0 feedthrough
rlabel pdiffusion 892 -3409 892 -3409 0 cellNo=720
rlabel pdiffusion 899 -3409 899 -3409 0 feedthrough
rlabel pdiffusion 906 -3409 906 -3409 0 feedthrough
rlabel pdiffusion 913 -3409 913 -3409 0 feedthrough
rlabel pdiffusion 920 -3409 920 -3409 0 feedthrough
rlabel pdiffusion 927 -3409 927 -3409 0 feedthrough
rlabel pdiffusion 934 -3409 934 -3409 0 feedthrough
rlabel pdiffusion 941 -3409 941 -3409 0 feedthrough
rlabel pdiffusion 948 -3409 948 -3409 0 cellNo=310
rlabel pdiffusion 955 -3409 955 -3409 0 feedthrough
rlabel pdiffusion 962 -3409 962 -3409 0 feedthrough
rlabel pdiffusion 969 -3409 969 -3409 0 feedthrough
rlabel pdiffusion 976 -3409 976 -3409 0 feedthrough
rlabel pdiffusion 983 -3409 983 -3409 0 feedthrough
rlabel pdiffusion 990 -3409 990 -3409 0 feedthrough
rlabel pdiffusion 997 -3409 997 -3409 0 feedthrough
rlabel pdiffusion 1004 -3409 1004 -3409 0 feedthrough
rlabel pdiffusion 1011 -3409 1011 -3409 0 cellNo=209
rlabel pdiffusion 1018 -3409 1018 -3409 0 cellNo=853
rlabel pdiffusion 1025 -3409 1025 -3409 0 cellNo=495
rlabel pdiffusion 1032 -3409 1032 -3409 0 feedthrough
rlabel pdiffusion 1039 -3409 1039 -3409 0 cellNo=753
rlabel pdiffusion 1046 -3409 1046 -3409 0 feedthrough
rlabel pdiffusion 1053 -3409 1053 -3409 0 cellNo=812
rlabel pdiffusion 1060 -3409 1060 -3409 0 cellNo=989
rlabel pdiffusion 1067 -3409 1067 -3409 0 feedthrough
rlabel pdiffusion 1074 -3409 1074 -3409 0 feedthrough
rlabel pdiffusion 1081 -3409 1081 -3409 0 feedthrough
rlabel pdiffusion 1088 -3409 1088 -3409 0 feedthrough
rlabel pdiffusion 1095 -3409 1095 -3409 0 feedthrough
rlabel pdiffusion 1102 -3409 1102 -3409 0 feedthrough
rlabel pdiffusion 1109 -3409 1109 -3409 0 cellNo=326
rlabel pdiffusion 1116 -3409 1116 -3409 0 feedthrough
rlabel pdiffusion 1123 -3409 1123 -3409 0 feedthrough
rlabel pdiffusion 1130 -3409 1130 -3409 0 feedthrough
rlabel pdiffusion 1137 -3409 1137 -3409 0 feedthrough
rlabel pdiffusion 1144 -3409 1144 -3409 0 feedthrough
rlabel pdiffusion 1151 -3409 1151 -3409 0 cellNo=80
rlabel pdiffusion 1158 -3409 1158 -3409 0 cellNo=940
rlabel pdiffusion 1165 -3409 1165 -3409 0 cellNo=960
rlabel pdiffusion 1172 -3409 1172 -3409 0 feedthrough
rlabel pdiffusion 1186 -3409 1186 -3409 0 feedthrough
rlabel pdiffusion 1193 -3409 1193 -3409 0 feedthrough
rlabel pdiffusion 1200 -3409 1200 -3409 0 feedthrough
rlabel pdiffusion 1207 -3409 1207 -3409 0 feedthrough
rlabel pdiffusion 1214 -3409 1214 -3409 0 cellNo=996
rlabel pdiffusion 1235 -3409 1235 -3409 0 feedthrough
rlabel pdiffusion 1242 -3409 1242 -3409 0 feedthrough
rlabel pdiffusion 1249 -3409 1249 -3409 0 feedthrough
rlabel pdiffusion 1263 -3409 1263 -3409 0 cellNo=985
rlabel pdiffusion 1312 -3409 1312 -3409 0 feedthrough
rlabel pdiffusion 1319 -3409 1319 -3409 0 feedthrough
rlabel pdiffusion 1333 -3409 1333 -3409 0 feedthrough
rlabel pdiffusion 1375 -3409 1375 -3409 0 feedthrough
rlabel pdiffusion 1382 -3409 1382 -3409 0 feedthrough
rlabel pdiffusion 1389 -3409 1389 -3409 0 feedthrough
rlabel pdiffusion 1578 -3409 1578 -3409 0 feedthrough
rlabel pdiffusion 3 -3456 3 -3456 0 cellNo=1051
rlabel pdiffusion 10 -3456 10 -3456 0 cellNo=1052
rlabel pdiffusion 17 -3456 17 -3456 0 cellNo=1056
rlabel pdiffusion 24 -3456 24 -3456 0 cellNo=1059
rlabel pdiffusion 31 -3456 31 -3456 0 cellNo=1066
rlabel pdiffusion 38 -3456 38 -3456 0 cellNo=1073
rlabel pdiffusion 45 -3456 45 -3456 0 cellNo=1094
rlabel pdiffusion 52 -3456 52 -3456 0 cellNo=1101
rlabel pdiffusion 59 -3456 59 -3456 0 cellNo=1106
rlabel pdiffusion 66 -3456 66 -3456 0 cellNo=1112
rlabel pdiffusion 73 -3456 73 -3456 0 cellNo=1130
rlabel pdiffusion 80 -3456 80 -3456 0 cellNo=1134
rlabel pdiffusion 87 -3456 87 -3456 0 cellNo=1146
rlabel pdiffusion 94 -3456 94 -3456 0 cellNo=1168
rlabel pdiffusion 101 -3456 101 -3456 0 cellNo=1174
rlabel pdiffusion 262 -3456 262 -3456 0 feedthrough
rlabel pdiffusion 311 -3456 311 -3456 0 feedthrough
rlabel pdiffusion 318 -3456 318 -3456 0 feedthrough
rlabel pdiffusion 339 -3456 339 -3456 0 feedthrough
rlabel pdiffusion 346 -3456 346 -3456 0 feedthrough
rlabel pdiffusion 353 -3456 353 -3456 0 cellNo=777
rlabel pdiffusion 360 -3456 360 -3456 0 feedthrough
rlabel pdiffusion 367 -3456 367 -3456 0 feedthrough
rlabel pdiffusion 374 -3456 374 -3456 0 feedthrough
rlabel pdiffusion 381 -3456 381 -3456 0 feedthrough
rlabel pdiffusion 388 -3456 388 -3456 0 feedthrough
rlabel pdiffusion 395 -3456 395 -3456 0 feedthrough
rlabel pdiffusion 402 -3456 402 -3456 0 feedthrough
rlabel pdiffusion 409 -3456 409 -3456 0 cellNo=465
rlabel pdiffusion 416 -3456 416 -3456 0 feedthrough
rlabel pdiffusion 423 -3456 423 -3456 0 feedthrough
rlabel pdiffusion 430 -3456 430 -3456 0 feedthrough
rlabel pdiffusion 437 -3456 437 -3456 0 feedthrough
rlabel pdiffusion 444 -3456 444 -3456 0 feedthrough
rlabel pdiffusion 451 -3456 451 -3456 0 feedthrough
rlabel pdiffusion 458 -3456 458 -3456 0 feedthrough
rlabel pdiffusion 465 -3456 465 -3456 0 feedthrough
rlabel pdiffusion 472 -3456 472 -3456 0 cellNo=976
rlabel pdiffusion 479 -3456 479 -3456 0 feedthrough
rlabel pdiffusion 486 -3456 486 -3456 0 feedthrough
rlabel pdiffusion 493 -3456 493 -3456 0 feedthrough
rlabel pdiffusion 500 -3456 500 -3456 0 feedthrough
rlabel pdiffusion 507 -3456 507 -3456 0 cellNo=368
rlabel pdiffusion 514 -3456 514 -3456 0 feedthrough
rlabel pdiffusion 521 -3456 521 -3456 0 feedthrough
rlabel pdiffusion 528 -3456 528 -3456 0 feedthrough
rlabel pdiffusion 535 -3456 535 -3456 0 feedthrough
rlabel pdiffusion 542 -3456 542 -3456 0 feedthrough
rlabel pdiffusion 549 -3456 549 -3456 0 feedthrough
rlabel pdiffusion 556 -3456 556 -3456 0 feedthrough
rlabel pdiffusion 563 -3456 563 -3456 0 feedthrough
rlabel pdiffusion 570 -3456 570 -3456 0 feedthrough
rlabel pdiffusion 577 -3456 577 -3456 0 feedthrough
rlabel pdiffusion 584 -3456 584 -3456 0 cellNo=623
rlabel pdiffusion 591 -3456 591 -3456 0 cellNo=984
rlabel pdiffusion 598 -3456 598 -3456 0 feedthrough
rlabel pdiffusion 605 -3456 605 -3456 0 cellNo=727
rlabel pdiffusion 612 -3456 612 -3456 0 feedthrough
rlabel pdiffusion 619 -3456 619 -3456 0 cellNo=373
rlabel pdiffusion 626 -3456 626 -3456 0 feedthrough
rlabel pdiffusion 633 -3456 633 -3456 0 feedthrough
rlabel pdiffusion 640 -3456 640 -3456 0 feedthrough
rlabel pdiffusion 647 -3456 647 -3456 0 feedthrough
rlabel pdiffusion 654 -3456 654 -3456 0 cellNo=670
rlabel pdiffusion 661 -3456 661 -3456 0 cellNo=352
rlabel pdiffusion 668 -3456 668 -3456 0 feedthrough
rlabel pdiffusion 675 -3456 675 -3456 0 feedthrough
rlabel pdiffusion 682 -3456 682 -3456 0 feedthrough
rlabel pdiffusion 689 -3456 689 -3456 0 feedthrough
rlabel pdiffusion 696 -3456 696 -3456 0 feedthrough
rlabel pdiffusion 703 -3456 703 -3456 0 feedthrough
rlabel pdiffusion 710 -3456 710 -3456 0 feedthrough
rlabel pdiffusion 717 -3456 717 -3456 0 cellNo=562
rlabel pdiffusion 724 -3456 724 -3456 0 feedthrough
rlabel pdiffusion 731 -3456 731 -3456 0 feedthrough
rlabel pdiffusion 738 -3456 738 -3456 0 feedthrough
rlabel pdiffusion 745 -3456 745 -3456 0 feedthrough
rlabel pdiffusion 752 -3456 752 -3456 0 feedthrough
rlabel pdiffusion 759 -3456 759 -3456 0 feedthrough
rlabel pdiffusion 766 -3456 766 -3456 0 feedthrough
rlabel pdiffusion 773 -3456 773 -3456 0 feedthrough
rlabel pdiffusion 780 -3456 780 -3456 0 feedthrough
rlabel pdiffusion 787 -3456 787 -3456 0 feedthrough
rlabel pdiffusion 794 -3456 794 -3456 0 feedthrough
rlabel pdiffusion 801 -3456 801 -3456 0 feedthrough
rlabel pdiffusion 808 -3456 808 -3456 0 cellNo=854
rlabel pdiffusion 815 -3456 815 -3456 0 feedthrough
rlabel pdiffusion 822 -3456 822 -3456 0 cellNo=888
rlabel pdiffusion 829 -3456 829 -3456 0 feedthrough
rlabel pdiffusion 836 -3456 836 -3456 0 feedthrough
rlabel pdiffusion 843 -3456 843 -3456 0 feedthrough
rlabel pdiffusion 850 -3456 850 -3456 0 cellNo=675
rlabel pdiffusion 857 -3456 857 -3456 0 feedthrough
rlabel pdiffusion 864 -3456 864 -3456 0 feedthrough
rlabel pdiffusion 871 -3456 871 -3456 0 feedthrough
rlabel pdiffusion 878 -3456 878 -3456 0 feedthrough
rlabel pdiffusion 885 -3456 885 -3456 0 feedthrough
rlabel pdiffusion 892 -3456 892 -3456 0 feedthrough
rlabel pdiffusion 899 -3456 899 -3456 0 feedthrough
rlabel pdiffusion 906 -3456 906 -3456 0 feedthrough
rlabel pdiffusion 913 -3456 913 -3456 0 feedthrough
rlabel pdiffusion 920 -3456 920 -3456 0 feedthrough
rlabel pdiffusion 927 -3456 927 -3456 0 feedthrough
rlabel pdiffusion 934 -3456 934 -3456 0 feedthrough
rlabel pdiffusion 941 -3456 941 -3456 0 feedthrough
rlabel pdiffusion 948 -3456 948 -3456 0 feedthrough
rlabel pdiffusion 955 -3456 955 -3456 0 feedthrough
rlabel pdiffusion 962 -3456 962 -3456 0 feedthrough
rlabel pdiffusion 969 -3456 969 -3456 0 cellNo=180
rlabel pdiffusion 976 -3456 976 -3456 0 feedthrough
rlabel pdiffusion 983 -3456 983 -3456 0 feedthrough
rlabel pdiffusion 990 -3456 990 -3456 0 feedthrough
rlabel pdiffusion 997 -3456 997 -3456 0 cellNo=964
rlabel pdiffusion 1004 -3456 1004 -3456 0 feedthrough
rlabel pdiffusion 1011 -3456 1011 -3456 0 feedthrough
rlabel pdiffusion 1018 -3456 1018 -3456 0 feedthrough
rlabel pdiffusion 1025 -3456 1025 -3456 0 feedthrough
rlabel pdiffusion 1032 -3456 1032 -3456 0 feedthrough
rlabel pdiffusion 1053 -3456 1053 -3456 0 feedthrough
rlabel pdiffusion 1074 -3456 1074 -3456 0 feedthrough
rlabel pdiffusion 1081 -3456 1081 -3456 0 feedthrough
rlabel pdiffusion 1102 -3456 1102 -3456 0 feedthrough
rlabel pdiffusion 1116 -3456 1116 -3456 0 feedthrough
rlabel pdiffusion 1123 -3456 1123 -3456 0 feedthrough
rlabel pdiffusion 1130 -3456 1130 -3456 0 feedthrough
rlabel pdiffusion 1137 -3456 1137 -3456 0 feedthrough
rlabel pdiffusion 1144 -3456 1144 -3456 0 feedthrough
rlabel pdiffusion 1193 -3456 1193 -3456 0 feedthrough
rlabel pdiffusion 1200 -3456 1200 -3456 0 feedthrough
rlabel pdiffusion 1207 -3456 1207 -3456 0 feedthrough
rlabel pdiffusion 1214 -3456 1214 -3456 0 feedthrough
rlabel pdiffusion 1270 -3456 1270 -3456 0 feedthrough
rlabel pdiffusion 1298 -3456 1298 -3456 0 cellNo=918
rlabel pdiffusion 1305 -3456 1305 -3456 0 feedthrough
rlabel pdiffusion 1319 -3456 1319 -3456 0 feedthrough
rlabel pdiffusion 1347 -3456 1347 -3456 0 feedthrough
rlabel pdiffusion 1382 -3456 1382 -3456 0 feedthrough
rlabel pdiffusion 1389 -3456 1389 -3456 0 feedthrough
rlabel pdiffusion 1396 -3456 1396 -3456 0 feedthrough
rlabel pdiffusion 1578 -3456 1578 -3456 0 feedthrough
rlabel pdiffusion 3 -3497 3 -3497 0 cellNo=1086
rlabel pdiffusion 10 -3497 10 -3497 0 cellNo=1087
rlabel pdiffusion 17 -3497 17 -3497 0 cellNo=1088
rlabel pdiffusion 24 -3497 24 -3497 0 cellNo=1089
rlabel pdiffusion 31 -3497 31 -3497 0 cellNo=1090
rlabel pdiffusion 38 -3497 38 -3497 0 cellNo=1093
rlabel pdiffusion 45 -3497 45 -3497 0 cellNo=1099
rlabel pdiffusion 52 -3497 52 -3497 0 cellNo=1105
rlabel pdiffusion 59 -3497 59 -3497 0 cellNo=1109
rlabel pdiffusion 66 -3497 66 -3497 0 cellNo=1119
rlabel pdiffusion 73 -3497 73 -3497 0 cellNo=1133
rlabel pdiffusion 80 -3497 80 -3497 0 cellNo=1138
rlabel pdiffusion 87 -3497 87 -3497 0 cellNo=1140
rlabel pdiffusion 94 -3497 94 -3497 0 cellNo=1152
rlabel pdiffusion 101 -3497 101 -3497 0 cellNo=1173
rlabel pdiffusion 108 -3497 108 -3497 0 cellNo=1176
rlabel pdiffusion 115 -3497 115 -3497 0 cellNo=1180
rlabel pdiffusion 122 -3497 122 -3497 0 cellNo=1187
rlabel pdiffusion 269 -3497 269 -3497 0 feedthrough
rlabel pdiffusion 283 -3497 283 -3497 0 cellNo=900
rlabel pdiffusion 297 -3497 297 -3497 0 feedthrough
rlabel pdiffusion 367 -3497 367 -3497 0 feedthrough
rlabel pdiffusion 374 -3497 374 -3497 0 feedthrough
rlabel pdiffusion 381 -3497 381 -3497 0 feedthrough
rlabel pdiffusion 388 -3497 388 -3497 0 cellNo=500
rlabel pdiffusion 409 -3497 409 -3497 0 feedthrough
rlabel pdiffusion 423 -3497 423 -3497 0 cellNo=136
rlabel pdiffusion 430 -3497 430 -3497 0 feedthrough
rlabel pdiffusion 437 -3497 437 -3497 0 cellNo=1000
rlabel pdiffusion 444 -3497 444 -3497 0 feedthrough
rlabel pdiffusion 451 -3497 451 -3497 0 feedthrough
rlabel pdiffusion 458 -3497 458 -3497 0 feedthrough
rlabel pdiffusion 472 -3497 472 -3497 0 feedthrough
rlabel pdiffusion 479 -3497 479 -3497 0 feedthrough
rlabel pdiffusion 486 -3497 486 -3497 0 feedthrough
rlabel pdiffusion 493 -3497 493 -3497 0 feedthrough
rlabel pdiffusion 500 -3497 500 -3497 0 feedthrough
rlabel pdiffusion 507 -3497 507 -3497 0 feedthrough
rlabel pdiffusion 514 -3497 514 -3497 0 feedthrough
rlabel pdiffusion 528 -3497 528 -3497 0 feedthrough
rlabel pdiffusion 535 -3497 535 -3497 0 feedthrough
rlabel pdiffusion 542 -3497 542 -3497 0 feedthrough
rlabel pdiffusion 549 -3497 549 -3497 0 feedthrough
rlabel pdiffusion 556 -3497 556 -3497 0 feedthrough
rlabel pdiffusion 563 -3497 563 -3497 0 feedthrough
rlabel pdiffusion 570 -3497 570 -3497 0 feedthrough
rlabel pdiffusion 577 -3497 577 -3497 0 feedthrough
rlabel pdiffusion 584 -3497 584 -3497 0 feedthrough
rlabel pdiffusion 591 -3497 591 -3497 0 feedthrough
rlabel pdiffusion 605 -3497 605 -3497 0 feedthrough
rlabel pdiffusion 619 -3497 619 -3497 0 feedthrough
rlabel pdiffusion 633 -3497 633 -3497 0 feedthrough
rlabel pdiffusion 640 -3497 640 -3497 0 feedthrough
rlabel pdiffusion 647 -3497 647 -3497 0 feedthrough
rlabel pdiffusion 654 -3497 654 -3497 0 cellNo=322
rlabel pdiffusion 689 -3497 689 -3497 0 feedthrough
rlabel pdiffusion 696 -3497 696 -3497 0 feedthrough
rlabel pdiffusion 703 -3497 703 -3497 0 feedthrough
rlabel pdiffusion 710 -3497 710 -3497 0 feedthrough
rlabel pdiffusion 717 -3497 717 -3497 0 feedthrough
rlabel pdiffusion 724 -3497 724 -3497 0 cellNo=699
rlabel pdiffusion 731 -3497 731 -3497 0 cellNo=974
rlabel pdiffusion 738 -3497 738 -3497 0 feedthrough
rlabel pdiffusion 745 -3497 745 -3497 0 feedthrough
rlabel pdiffusion 752 -3497 752 -3497 0 cellNo=87
rlabel pdiffusion 759 -3497 759 -3497 0 feedthrough
rlabel pdiffusion 766 -3497 766 -3497 0 feedthrough
rlabel pdiffusion 773 -3497 773 -3497 0 feedthrough
rlabel pdiffusion 787 -3497 787 -3497 0 feedthrough
rlabel pdiffusion 794 -3497 794 -3497 0 feedthrough
rlabel pdiffusion 801 -3497 801 -3497 0 feedthrough
rlabel pdiffusion 808 -3497 808 -3497 0 feedthrough
rlabel pdiffusion 815 -3497 815 -3497 0 feedthrough
rlabel pdiffusion 822 -3497 822 -3497 0 feedthrough
rlabel pdiffusion 829 -3497 829 -3497 0 feedthrough
rlabel pdiffusion 878 -3497 878 -3497 0 feedthrough
rlabel pdiffusion 885 -3497 885 -3497 0 feedthrough
rlabel pdiffusion 892 -3497 892 -3497 0 feedthrough
rlabel pdiffusion 899 -3497 899 -3497 0 feedthrough
rlabel pdiffusion 906 -3497 906 -3497 0 feedthrough
rlabel pdiffusion 913 -3497 913 -3497 0 cellNo=982
rlabel pdiffusion 920 -3497 920 -3497 0 feedthrough
rlabel pdiffusion 927 -3497 927 -3497 0 feedthrough
rlabel pdiffusion 934 -3497 934 -3497 0 feedthrough
rlabel pdiffusion 941 -3497 941 -3497 0 feedthrough
rlabel pdiffusion 948 -3497 948 -3497 0 feedthrough
rlabel pdiffusion 955 -3497 955 -3497 0 feedthrough
rlabel pdiffusion 962 -3497 962 -3497 0 feedthrough
rlabel pdiffusion 976 -3497 976 -3497 0 feedthrough
rlabel pdiffusion 997 -3497 997 -3497 0 feedthrough
rlabel pdiffusion 1004 -3497 1004 -3497 0 cellNo=253
rlabel pdiffusion 1011 -3497 1011 -3497 0 feedthrough
rlabel pdiffusion 1025 -3497 1025 -3497 0 feedthrough
rlabel pdiffusion 1039 -3497 1039 -3497 0 feedthrough
rlabel pdiffusion 1046 -3497 1046 -3497 0 feedthrough
rlabel pdiffusion 1053 -3497 1053 -3497 0 feedthrough
rlabel pdiffusion 1060 -3497 1060 -3497 0 feedthrough
rlabel pdiffusion 1067 -3497 1067 -3497 0 feedthrough
rlabel pdiffusion 1074 -3497 1074 -3497 0 feedthrough
rlabel pdiffusion 1081 -3497 1081 -3497 0 feedthrough
rlabel pdiffusion 1088 -3497 1088 -3497 0 cellNo=781
rlabel pdiffusion 1116 -3497 1116 -3497 0 feedthrough
rlabel pdiffusion 1123 -3497 1123 -3497 0 feedthrough
rlabel pdiffusion 1137 -3497 1137 -3497 0 feedthrough
rlabel pdiffusion 1158 -3497 1158 -3497 0 feedthrough
rlabel pdiffusion 1179 -3497 1179 -3497 0 cellNo=523
rlabel pdiffusion 1186 -3497 1186 -3497 0 feedthrough
rlabel pdiffusion 1193 -3497 1193 -3497 0 feedthrough
rlabel pdiffusion 1235 -3497 1235 -3497 0 feedthrough
rlabel pdiffusion 1249 -3497 1249 -3497 0 feedthrough
rlabel pdiffusion 1270 -3497 1270 -3497 0 feedthrough
rlabel pdiffusion 1277 -3497 1277 -3497 0 feedthrough
rlabel pdiffusion 1375 -3497 1375 -3497 0 feedthrough
rlabel pdiffusion 1382 -3497 1382 -3497 0 cellNo=427
rlabel pdiffusion 1389 -3497 1389 -3497 0 feedthrough
rlabel pdiffusion 1396 -3497 1396 -3497 0 feedthrough
rlabel pdiffusion 1417 -3497 1417 -3497 0 feedthrough
rlabel pdiffusion 1578 -3497 1578 -3497 0 feedthrough
rlabel pdiffusion 3 -3528 3 -3528 0 cellNo=1121
rlabel pdiffusion 10 -3528 10 -3528 0 cellNo=1122
rlabel pdiffusion 17 -3528 17 -3528 0 cellNo=1123
rlabel pdiffusion 24 -3528 24 -3528 0 cellNo=1124
rlabel pdiffusion 31 -3528 31 -3528 0 cellNo=1125
rlabel pdiffusion 38 -3528 38 -3528 0 cellNo=1126
rlabel pdiffusion 45 -3528 45 -3528 0 cellNo=1127
rlabel pdiffusion 52 -3528 52 -3528 0 cellNo=1128
rlabel pdiffusion 59 -3528 59 -3528 0 cellNo=1129
rlabel pdiffusion 66 -3528 66 -3528 0 cellNo=1131
rlabel pdiffusion 73 -3528 73 -3528 0 cellNo=1135
rlabel pdiffusion 80 -3528 80 -3528 0 cellNo=1139
rlabel pdiffusion 87 -3528 87 -3528 0 cellNo=1151
rlabel pdiffusion 94 -3528 94 -3528 0 cellNo=1171
rlabel pdiffusion 381 -3528 381 -3528 0 feedthrough
rlabel pdiffusion 388 -3528 388 -3528 0 feedthrough
rlabel pdiffusion 395 -3528 395 -3528 0 feedthrough
rlabel pdiffusion 402 -3528 402 -3528 0 feedthrough
rlabel pdiffusion 430 -3528 430 -3528 0 feedthrough
rlabel pdiffusion 444 -3528 444 -3528 0 feedthrough
rlabel pdiffusion 451 -3528 451 -3528 0 feedthrough
rlabel pdiffusion 465 -3528 465 -3528 0 feedthrough
rlabel pdiffusion 479 -3528 479 -3528 0 cellNo=477
rlabel pdiffusion 486 -3528 486 -3528 0 feedthrough
rlabel pdiffusion 493 -3528 493 -3528 0 feedthrough
rlabel pdiffusion 500 -3528 500 -3528 0 feedthrough
rlabel pdiffusion 507 -3528 507 -3528 0 feedthrough
rlabel pdiffusion 514 -3528 514 -3528 0 feedthrough
rlabel pdiffusion 521 -3528 521 -3528 0 cellNo=285
rlabel pdiffusion 528 -3528 528 -3528 0 feedthrough
rlabel pdiffusion 535 -3528 535 -3528 0 feedthrough
rlabel pdiffusion 542 -3528 542 -3528 0 feedthrough
rlabel pdiffusion 549 -3528 549 -3528 0 feedthrough
rlabel pdiffusion 556 -3528 556 -3528 0 cellNo=366
rlabel pdiffusion 563 -3528 563 -3528 0 cellNo=891
rlabel pdiffusion 570 -3528 570 -3528 0 feedthrough
rlabel pdiffusion 577 -3528 577 -3528 0 feedthrough
rlabel pdiffusion 584 -3528 584 -3528 0 feedthrough
rlabel pdiffusion 591 -3528 591 -3528 0 feedthrough
rlabel pdiffusion 598 -3528 598 -3528 0 feedthrough
rlabel pdiffusion 605 -3528 605 -3528 0 feedthrough
rlabel pdiffusion 647 -3528 647 -3528 0 feedthrough
rlabel pdiffusion 654 -3528 654 -3528 0 feedthrough
rlabel pdiffusion 675 -3528 675 -3528 0 feedthrough
rlabel pdiffusion 696 -3528 696 -3528 0 feedthrough
rlabel pdiffusion 703 -3528 703 -3528 0 feedthrough
rlabel pdiffusion 710 -3528 710 -3528 0 feedthrough
rlabel pdiffusion 731 -3528 731 -3528 0 feedthrough
rlabel pdiffusion 759 -3528 759 -3528 0 feedthrough
rlabel pdiffusion 766 -3528 766 -3528 0 feedthrough
rlabel pdiffusion 773 -3528 773 -3528 0 feedthrough
rlabel pdiffusion 780 -3528 780 -3528 0 feedthrough
rlabel pdiffusion 787 -3528 787 -3528 0 feedthrough
rlabel pdiffusion 794 -3528 794 -3528 0 feedthrough
rlabel pdiffusion 801 -3528 801 -3528 0 feedthrough
rlabel pdiffusion 808 -3528 808 -3528 0 feedthrough
rlabel pdiffusion 815 -3528 815 -3528 0 feedthrough
rlabel pdiffusion 822 -3528 822 -3528 0 cellNo=396
rlabel pdiffusion 843 -3528 843 -3528 0 feedthrough
rlabel pdiffusion 864 -3528 864 -3528 0 feedthrough
rlabel pdiffusion 878 -3528 878 -3528 0 feedthrough
rlabel pdiffusion 885 -3528 885 -3528 0 feedthrough
rlabel pdiffusion 892 -3528 892 -3528 0 cellNo=347
rlabel pdiffusion 899 -3528 899 -3528 0 feedthrough
rlabel pdiffusion 906 -3528 906 -3528 0 feedthrough
rlabel pdiffusion 920 -3528 920 -3528 0 feedthrough
rlabel pdiffusion 927 -3528 927 -3528 0 feedthrough
rlabel pdiffusion 934 -3528 934 -3528 0 feedthrough
rlabel pdiffusion 941 -3528 941 -3528 0 feedthrough
rlabel pdiffusion 948 -3528 948 -3528 0 cellNo=154
rlabel pdiffusion 955 -3528 955 -3528 0 cellNo=754
rlabel pdiffusion 962 -3528 962 -3528 0 cellNo=534
rlabel pdiffusion 969 -3528 969 -3528 0 feedthrough
rlabel pdiffusion 1004 -3528 1004 -3528 0 cellNo=233
rlabel pdiffusion 1018 -3528 1018 -3528 0 cellNo=717
rlabel pdiffusion 1032 -3528 1032 -3528 0 cellNo=693
rlabel pdiffusion 1039 -3528 1039 -3528 0 cellNo=644
rlabel pdiffusion 1046 -3528 1046 -3528 0 feedthrough
rlabel pdiffusion 1053 -3528 1053 -3528 0 feedthrough
rlabel pdiffusion 1060 -3528 1060 -3528 0 cellNo=8
rlabel pdiffusion 1074 -3528 1074 -3528 0 feedthrough
rlabel pdiffusion 1116 -3528 1116 -3528 0 feedthrough
rlabel pdiffusion 1130 -3528 1130 -3528 0 feedthrough
rlabel pdiffusion 1137 -3528 1137 -3528 0 feedthrough
rlabel pdiffusion 1144 -3528 1144 -3528 0 feedthrough
rlabel pdiffusion 1158 -3528 1158 -3528 0 cellNo=260
rlabel pdiffusion 1165 -3528 1165 -3528 0 feedthrough
rlabel pdiffusion 1179 -3528 1179 -3528 0 feedthrough
rlabel pdiffusion 1193 -3528 1193 -3528 0 feedthrough
rlabel pdiffusion 1263 -3528 1263 -3528 0 feedthrough
rlabel pdiffusion 1277 -3528 1277 -3528 0 cellNo=817
rlabel pdiffusion 1340 -3528 1340 -3528 0 feedthrough
rlabel pdiffusion 1382 -3528 1382 -3528 0 feedthrough
rlabel pdiffusion 1396 -3528 1396 -3528 0 feedthrough
rlabel pdiffusion 1501 -3528 1501 -3528 0 feedthrough
rlabel pdiffusion 1578 -3528 1578 -3528 0 cellNo=660
rlabel pdiffusion 3 -3557 3 -3557 0 cellNo=1156
rlabel pdiffusion 10 -3557 10 -3557 0 cellNo=1157
rlabel pdiffusion 17 -3557 17 -3557 0 cellNo=1158
rlabel pdiffusion 24 -3557 24 -3557 0 cellNo=1159
rlabel pdiffusion 31 -3557 31 -3557 0 cellNo=1160
rlabel pdiffusion 38 -3557 38 -3557 0 cellNo=1161
rlabel pdiffusion 45 -3557 45 -3557 0 cellNo=1162
rlabel pdiffusion 52 -3557 52 -3557 0 cellNo=1163
rlabel pdiffusion 59 -3557 59 -3557 0 cellNo=1164
rlabel pdiffusion 66 -3557 66 -3557 0 cellNo=1165
rlabel pdiffusion 73 -3557 73 -3557 0 cellNo=1166
rlabel pdiffusion 80 -3557 80 -3557 0 cellNo=1167
rlabel pdiffusion 87 -3557 87 -3557 0 cellNo=1170
rlabel pdiffusion 94 -3557 94 -3557 0 cellNo=1175
rlabel pdiffusion 101 -3557 101 -3557 0 cellNo=1178
rlabel pdiffusion 108 -3557 108 -3557 0 cellNo=1181
rlabel pdiffusion 115 -3557 115 -3557 0 cellNo=1184
rlabel pdiffusion 381 -3557 381 -3557 0 feedthrough
rlabel pdiffusion 388 -3557 388 -3557 0 feedthrough
rlabel pdiffusion 395 -3557 395 -3557 0 feedthrough
rlabel pdiffusion 402 -3557 402 -3557 0 feedthrough
rlabel pdiffusion 409 -3557 409 -3557 0 feedthrough
rlabel pdiffusion 451 -3557 451 -3557 0 feedthrough
rlabel pdiffusion 458 -3557 458 -3557 0 feedthrough
rlabel pdiffusion 472 -3557 472 -3557 0 cellNo=569
rlabel pdiffusion 479 -3557 479 -3557 0 feedthrough
rlabel pdiffusion 493 -3557 493 -3557 0 feedthrough
rlabel pdiffusion 500 -3557 500 -3557 0 cellNo=850
rlabel pdiffusion 507 -3557 507 -3557 0 feedthrough
rlabel pdiffusion 514 -3557 514 -3557 0 feedthrough
rlabel pdiffusion 528 -3557 528 -3557 0 cellNo=932
rlabel pdiffusion 535 -3557 535 -3557 0 feedthrough
rlabel pdiffusion 542 -3557 542 -3557 0 feedthrough
rlabel pdiffusion 549 -3557 549 -3557 0 feedthrough
rlabel pdiffusion 556 -3557 556 -3557 0 feedthrough
rlabel pdiffusion 563 -3557 563 -3557 0 cellNo=713
rlabel pdiffusion 570 -3557 570 -3557 0 feedthrough
rlabel pdiffusion 577 -3557 577 -3557 0 cellNo=893
rlabel pdiffusion 584 -3557 584 -3557 0 feedthrough
rlabel pdiffusion 591 -3557 591 -3557 0 feedthrough
rlabel pdiffusion 598 -3557 598 -3557 0 feedthrough
rlabel pdiffusion 605 -3557 605 -3557 0 cellNo=399
rlabel pdiffusion 661 -3557 661 -3557 0 cellNo=581
rlabel pdiffusion 668 -3557 668 -3557 0 feedthrough
rlabel pdiffusion 703 -3557 703 -3557 0 cellNo=698
rlabel pdiffusion 710 -3557 710 -3557 0 feedthrough
rlabel pdiffusion 738 -3557 738 -3557 0 feedthrough
rlabel pdiffusion 759 -3557 759 -3557 0 feedthrough
rlabel pdiffusion 766 -3557 766 -3557 0 cellNo=557
rlabel pdiffusion 773 -3557 773 -3557 0 feedthrough
rlabel pdiffusion 780 -3557 780 -3557 0 feedthrough
rlabel pdiffusion 787 -3557 787 -3557 0 feedthrough
rlabel pdiffusion 794 -3557 794 -3557 0 cellNo=994
rlabel pdiffusion 801 -3557 801 -3557 0 feedthrough
rlabel pdiffusion 808 -3557 808 -3557 0 feedthrough
rlabel pdiffusion 815 -3557 815 -3557 0 feedthrough
rlabel pdiffusion 878 -3557 878 -3557 0 feedthrough
rlabel pdiffusion 885 -3557 885 -3557 0 feedthrough
rlabel pdiffusion 899 -3557 899 -3557 0 feedthrough
rlabel pdiffusion 906 -3557 906 -3557 0 feedthrough
rlabel pdiffusion 927 -3557 927 -3557 0 feedthrough
rlabel pdiffusion 934 -3557 934 -3557 0 cellNo=113
rlabel pdiffusion 941 -3557 941 -3557 0 feedthrough
rlabel pdiffusion 948 -3557 948 -3557 0 cellNo=801
rlabel pdiffusion 1109 -3557 1109 -3557 0 cellNo=606
rlabel pdiffusion 1116 -3557 1116 -3557 0 feedthrough
rlabel pdiffusion 1130 -3557 1130 -3557 0 feedthrough
rlabel pdiffusion 1137 -3557 1137 -3557 0 feedthrough
rlabel pdiffusion 1165 -3557 1165 -3557 0 feedthrough
rlabel pdiffusion 1179 -3557 1179 -3557 0 feedthrough
rlabel pdiffusion 1193 -3557 1193 -3557 0 feedthrough
rlabel pdiffusion 1361 -3557 1361 -3557 0 feedthrough
rlabel pdiffusion 1389 -3557 1389 -3557 0 feedthrough
rlabel pdiffusion 1396 -3557 1396 -3557 0 feedthrough
rlabel pdiffusion 3 -3572 3 -3572 0 cellNo=1149
rlabel pdiffusion 10 -3572 10 -3572 0 cellNo=1192
rlabel pdiffusion 17 -3572 17 -3572 0 cellNo=1193
rlabel pdiffusion 24 -3572 24 -3572 0 cellNo=1194
rlabel pdiffusion 31 -3572 31 -3572 0 cellNo=1195
rlabel pdiffusion 38 -3572 38 -3572 0 cellNo=1196
rlabel pdiffusion 45 -3572 45 -3572 0 cellNo=1197
rlabel pdiffusion 52 -3572 52 -3572 0 cellNo=1198
rlabel pdiffusion 59 -3572 59 -3572 0 cellNo=1199
rlabel pdiffusion 66 -3572 66 -3572 0 cellNo=1200
rlabel pdiffusion 73 -3572 73 -3572 0 cellNo=1191
rlabel pdiffusion 80 -3572 80 -3572 0 cellNo=1169
rlabel pdiffusion 87 -3572 87 -3572 0 cellNo=1185
rlabel pdiffusion 94 -3572 94 -3572 0 cellNo=1177
rlabel pdiffusion 101 -3572 101 -3572 0 cellNo=1188
rlabel pdiffusion 388 -3572 388 -3572 0 feedthrough
rlabel pdiffusion 395 -3572 395 -3572 0 cellNo=661
rlabel pdiffusion 402 -3572 402 -3572 0 cellNo=983
rlabel pdiffusion 409 -3572 409 -3572 0 feedthrough
rlabel pdiffusion 458 -3572 458 -3572 0 cellNo=2
rlabel pdiffusion 465 -3572 465 -3572 0 feedthrough
rlabel pdiffusion 493 -3572 493 -3572 0 feedthrough
rlabel pdiffusion 500 -3572 500 -3572 0 cellNo=418
rlabel pdiffusion 563 -3572 563 -3572 0 feedthrough
rlabel pdiffusion 577 -3572 577 -3572 0 cellNo=945
rlabel pdiffusion 591 -3572 591 -3572 0 feedthrough
rlabel pdiffusion 598 -3572 598 -3572 0 cellNo=609
rlabel pdiffusion 633 -3572 633 -3572 0 feedthrough
rlabel pdiffusion 745 -3572 745 -3572 0 cellNo=625
rlabel pdiffusion 759 -3572 759 -3572 0 feedthrough
rlabel pdiffusion 801 -3572 801 -3572 0 feedthrough
rlabel pdiffusion 808 -3572 808 -3572 0 cellNo=247
rlabel pdiffusion 885 -3572 885 -3572 0 feedthrough
rlabel pdiffusion 892 -3572 892 -3572 0 cellNo=700
rlabel pdiffusion 899 -3572 899 -3572 0 cellNo=461
rlabel pdiffusion 1130 -3572 1130 -3572 0 cellNo=775
rlabel pdiffusion 1137 -3572 1137 -3572 0 feedthrough
rlabel pdiffusion 1172 -3572 1172 -3572 0 feedthrough
rlabel pdiffusion 1179 -3572 1179 -3572 0 cellNo=972
rlabel pdiffusion 1186 -3572 1186 -3572 0 feedthrough
rlabel pdiffusion 1193 -3572 1193 -3572 0 cellNo=915
rlabel pdiffusion 1200 -3572 1200 -3572 0 feedthrough
rlabel pdiffusion 1389 -3572 1389 -3572 0 cellNo=933
rlabel pdiffusion 1396 -3572 1396 -3572 0 feedthrough
rlabel polysilicon 233 -14 233 -14 0 1
rlabel polysilicon 233 -20 233 -20 0 3
rlabel polysilicon 345 -14 345 -14 0 1
rlabel polysilicon 345 -20 345 -20 0 3
rlabel polysilicon 352 -14 352 -14 0 1
rlabel polysilicon 359 -14 359 -14 0 1
rlabel polysilicon 359 -20 359 -20 0 3
rlabel polysilicon 380 -14 380 -14 0 1
rlabel polysilicon 380 -20 380 -20 0 3
rlabel polysilicon 401 -14 401 -14 0 1
rlabel polysilicon 401 -20 401 -20 0 3
rlabel polysilicon 408 -14 408 -14 0 1
rlabel polysilicon 408 -20 408 -20 0 3
rlabel polysilicon 415 -14 415 -14 0 1
rlabel polysilicon 415 -20 415 -20 0 3
rlabel polysilicon 422 -14 422 -14 0 1
rlabel polysilicon 422 -20 422 -20 0 3
rlabel polysilicon 432 -14 432 -14 0 2
rlabel polysilicon 432 -20 432 -20 0 4
rlabel polysilicon 436 -14 436 -14 0 1
rlabel polysilicon 436 -20 436 -20 0 3
rlabel polysilicon 443 -14 443 -14 0 1
rlabel polysilicon 443 -20 443 -20 0 3
rlabel polysilicon 450 -14 450 -14 0 1
rlabel polysilicon 453 -14 453 -14 0 2
rlabel polysilicon 457 -14 457 -14 0 1
rlabel polysilicon 460 -14 460 -14 0 2
rlabel polysilicon 460 -20 460 -20 0 4
rlabel polysilicon 467 -14 467 -14 0 2
rlabel polysilicon 464 -20 464 -20 0 3
rlabel polysilicon 471 -14 471 -14 0 1
rlabel polysilicon 471 -20 471 -20 0 3
rlabel polysilicon 506 -14 506 -14 0 1
rlabel polysilicon 509 -20 509 -20 0 4
rlabel polysilicon 527 -14 527 -14 0 1
rlabel polysilicon 527 -20 527 -20 0 3
rlabel polysilicon 534 -14 534 -14 0 1
rlabel polysilicon 534 -20 534 -20 0 3
rlabel polysilicon 537 -20 537 -20 0 4
rlabel polysilicon 548 -14 548 -14 0 1
rlabel polysilicon 551 -20 551 -20 0 4
rlabel polysilicon 555 -14 555 -14 0 1
rlabel polysilicon 555 -20 555 -20 0 3
rlabel polysilicon 604 -14 604 -14 0 1
rlabel polysilicon 604 -20 604 -20 0 3
rlabel polysilicon 614 -14 614 -14 0 2
rlabel polysilicon 653 -14 653 -14 0 1
rlabel polysilicon 653 -20 653 -20 0 3
rlabel polysilicon 670 -14 670 -14 0 2
rlabel polysilicon 670 -20 670 -20 0 4
rlabel polysilicon 677 -14 677 -14 0 2
rlabel polysilicon 677 -20 677 -20 0 4
rlabel polysilicon 688 -14 688 -14 0 1
rlabel polysilicon 688 -20 688 -20 0 3
rlabel polysilicon 716 -14 716 -14 0 1
rlabel polysilicon 719 -20 719 -20 0 4
rlabel polysilicon 754 -14 754 -14 0 2
rlabel polysilicon 751 -20 751 -20 0 3
rlabel polysilicon 754 -20 754 -20 0 4
rlabel polysilicon 800 -14 800 -14 0 1
rlabel polysilicon 800 -20 800 -20 0 3
rlabel polysilicon 877 -14 877 -14 0 1
rlabel polysilicon 880 -20 880 -20 0 4
rlabel polysilicon 954 -14 954 -14 0 1
rlabel polysilicon 954 -20 954 -20 0 3
rlabel polysilicon 145 -51 145 -51 0 2
rlabel polysilicon 149 -51 149 -51 0 1
rlabel polysilicon 149 -57 149 -57 0 3
rlabel polysilicon 156 -51 156 -51 0 1
rlabel polysilicon 156 -57 156 -57 0 3
rlabel polysilicon 226 -51 226 -51 0 1
rlabel polysilicon 226 -57 226 -57 0 3
rlabel polysilicon 236 -51 236 -51 0 2
rlabel polysilicon 261 -51 261 -51 0 1
rlabel polysilicon 261 -57 261 -57 0 3
rlabel polysilicon 282 -51 282 -51 0 1
rlabel polysilicon 282 -57 282 -57 0 3
rlabel polysilicon 306 -51 306 -51 0 2
rlabel polysilicon 306 -57 306 -57 0 4
rlabel polysilicon 324 -51 324 -51 0 1
rlabel polysilicon 324 -57 324 -57 0 3
rlabel polysilicon 331 -51 331 -51 0 1
rlabel polysilicon 331 -57 331 -57 0 3
rlabel polysilicon 338 -51 338 -51 0 1
rlabel polysilicon 338 -57 338 -57 0 3
rlabel polysilicon 373 -51 373 -51 0 1
rlabel polysilicon 373 -57 373 -57 0 3
rlabel polysilicon 380 -51 380 -51 0 1
rlabel polysilicon 380 -57 380 -57 0 3
rlabel polysilicon 390 -51 390 -51 0 2
rlabel polysilicon 387 -57 387 -57 0 3
rlabel polysilicon 394 -51 394 -51 0 1
rlabel polysilicon 394 -57 394 -57 0 3
rlabel polysilicon 401 -51 401 -51 0 1
rlabel polysilicon 401 -57 401 -57 0 3
rlabel polysilicon 408 -51 408 -51 0 1
rlabel polysilicon 408 -57 408 -57 0 3
rlabel polysilicon 415 -57 415 -57 0 3
rlabel polysilicon 425 -51 425 -51 0 2
rlabel polysilicon 422 -57 422 -57 0 3
rlabel polysilicon 429 -51 429 -51 0 1
rlabel polysilicon 429 -57 429 -57 0 3
rlabel polysilicon 436 -51 436 -51 0 1
rlabel polysilicon 436 -57 436 -57 0 3
rlabel polysilicon 443 -51 443 -51 0 1
rlabel polysilicon 450 -51 450 -51 0 1
rlabel polysilicon 450 -57 450 -57 0 3
rlabel polysilicon 460 -51 460 -51 0 2
rlabel polysilicon 457 -57 457 -57 0 3
rlabel polysilicon 460 -57 460 -57 0 4
rlabel polysilicon 464 -51 464 -51 0 1
rlabel polysilicon 464 -57 464 -57 0 3
rlabel polysilicon 471 -51 471 -51 0 1
rlabel polysilicon 471 -57 471 -57 0 3
rlabel polysilicon 478 -51 478 -51 0 1
rlabel polysilicon 478 -57 478 -57 0 3
rlabel polysilicon 492 -51 492 -51 0 1
rlabel polysilicon 495 -51 495 -51 0 2
rlabel polysilicon 499 -51 499 -51 0 1
rlabel polysilicon 499 -57 499 -57 0 3
rlabel polysilicon 506 -51 506 -51 0 1
rlabel polysilicon 506 -57 506 -57 0 3
rlabel polysilicon 513 -51 513 -51 0 1
rlabel polysilicon 516 -51 516 -51 0 2
rlabel polysilicon 516 -57 516 -57 0 4
rlabel polysilicon 520 -51 520 -51 0 1
rlabel polysilicon 523 -51 523 -51 0 2
rlabel polysilicon 523 -57 523 -57 0 4
rlabel polysilicon 527 -51 527 -51 0 1
rlabel polysilicon 530 -51 530 -51 0 2
rlabel polysilicon 534 -51 534 -51 0 1
rlabel polysilicon 534 -57 534 -57 0 3
rlabel polysilicon 541 -51 541 -51 0 1
rlabel polysilicon 541 -57 541 -57 0 3
rlabel polysilicon 548 -51 548 -51 0 1
rlabel polysilicon 548 -57 548 -57 0 3
rlabel polysilicon 555 -51 555 -51 0 1
rlabel polysilicon 555 -57 555 -57 0 3
rlabel polysilicon 562 -51 562 -51 0 1
rlabel polysilicon 562 -57 562 -57 0 3
rlabel polysilicon 569 -57 569 -57 0 3
rlabel polysilicon 576 -51 576 -51 0 1
rlabel polysilicon 576 -57 576 -57 0 3
rlabel polysilicon 583 -51 583 -51 0 1
rlabel polysilicon 583 -57 583 -57 0 3
rlabel polysilicon 590 -51 590 -51 0 1
rlabel polysilicon 590 -57 590 -57 0 3
rlabel polysilicon 593 -57 593 -57 0 4
rlabel polysilicon 597 -51 597 -51 0 1
rlabel polysilicon 597 -57 597 -57 0 3
rlabel polysilicon 604 -51 604 -51 0 1
rlabel polysilicon 604 -57 604 -57 0 3
rlabel polysilicon 611 -51 611 -51 0 1
rlabel polysilicon 611 -57 611 -57 0 3
rlabel polysilicon 618 -51 618 -51 0 1
rlabel polysilicon 618 -57 618 -57 0 3
rlabel polysilicon 625 -51 625 -51 0 1
rlabel polysilicon 625 -57 625 -57 0 3
rlabel polysilicon 632 -51 632 -51 0 1
rlabel polysilicon 639 -51 639 -51 0 1
rlabel polysilicon 639 -57 639 -57 0 3
rlabel polysilicon 646 -51 646 -51 0 1
rlabel polysilicon 646 -57 646 -57 0 3
rlabel polysilicon 653 -51 653 -51 0 1
rlabel polysilicon 653 -57 653 -57 0 3
rlabel polysilicon 660 -51 660 -51 0 1
rlabel polysilicon 660 -57 660 -57 0 3
rlabel polysilicon 667 -51 667 -51 0 1
rlabel polysilicon 667 -57 667 -57 0 3
rlabel polysilicon 677 -51 677 -51 0 2
rlabel polysilicon 677 -57 677 -57 0 4
rlabel polysilicon 681 -51 681 -51 0 1
rlabel polysilicon 681 -57 681 -57 0 3
rlabel polysilicon 688 -51 688 -51 0 1
rlabel polysilicon 688 -57 688 -57 0 3
rlabel polysilicon 702 -51 702 -51 0 1
rlabel polysilicon 702 -57 702 -57 0 3
rlabel polysilicon 712 -51 712 -51 0 2
rlabel polysilicon 709 -57 709 -57 0 3
rlabel polysilicon 712 -57 712 -57 0 4
rlabel polysilicon 716 -51 716 -51 0 1
rlabel polysilicon 716 -57 716 -57 0 3
rlabel polysilicon 730 -51 730 -51 0 1
rlabel polysilicon 730 -57 730 -57 0 3
rlabel polysilicon 744 -51 744 -51 0 1
rlabel polysilicon 744 -57 744 -57 0 3
rlabel polysilicon 758 -51 758 -51 0 1
rlabel polysilicon 758 -57 758 -57 0 3
rlabel polysilicon 772 -51 772 -51 0 1
rlabel polysilicon 772 -57 772 -57 0 3
rlabel polysilicon 814 -51 814 -51 0 1
rlabel polysilicon 814 -57 814 -57 0 3
rlabel polysilicon 821 -51 821 -51 0 1
rlabel polysilicon 821 -57 821 -57 0 3
rlabel polysilicon 828 -51 828 -51 0 1
rlabel polysilicon 828 -57 828 -57 0 3
rlabel polysilicon 842 -51 842 -51 0 1
rlabel polysilicon 842 -57 842 -57 0 3
rlabel polysilicon 884 -51 884 -51 0 1
rlabel polysilicon 884 -57 884 -57 0 3
rlabel polysilicon 898 -51 898 -51 0 1
rlabel polysilicon 898 -57 898 -57 0 3
rlabel polysilicon 936 -57 936 -57 0 4
rlabel polysilicon 989 -51 989 -51 0 1
rlabel polysilicon 989 -57 989 -57 0 3
rlabel polysilicon 996 -51 996 -51 0 1
rlabel polysilicon 996 -57 996 -57 0 3
rlabel polysilicon 89 -104 89 -104 0 4
rlabel polysilicon 128 -98 128 -98 0 1
rlabel polysilicon 128 -104 128 -104 0 3
rlabel polysilicon 149 -98 149 -98 0 1
rlabel polysilicon 149 -104 149 -104 0 3
rlabel polysilicon 191 -98 191 -98 0 1
rlabel polysilicon 191 -104 191 -104 0 3
rlabel polysilicon 198 -98 198 -98 0 1
rlabel polysilicon 205 -98 205 -98 0 1
rlabel polysilicon 205 -104 205 -104 0 3
rlabel polysilicon 219 -98 219 -98 0 1
rlabel polysilicon 219 -104 219 -104 0 3
rlabel polysilicon 247 -98 247 -98 0 1
rlabel polysilicon 247 -104 247 -104 0 3
rlabel polysilicon 250 -104 250 -104 0 4
rlabel polysilicon 254 -98 254 -98 0 1
rlabel polysilicon 254 -104 254 -104 0 3
rlabel polysilicon 261 -98 261 -98 0 1
rlabel polysilicon 261 -104 261 -104 0 3
rlabel polysilicon 268 -98 268 -98 0 1
rlabel polysilicon 268 -104 268 -104 0 3
rlabel polysilicon 275 -98 275 -98 0 1
rlabel polysilicon 275 -104 275 -104 0 3
rlabel polysilicon 282 -98 282 -98 0 1
rlabel polysilicon 282 -104 282 -104 0 3
rlabel polysilicon 289 -98 289 -98 0 1
rlabel polysilicon 292 -104 292 -104 0 4
rlabel polysilicon 296 -98 296 -98 0 1
rlabel polysilicon 296 -104 296 -104 0 3
rlabel polysilicon 303 -98 303 -98 0 1
rlabel polysilicon 303 -104 303 -104 0 3
rlabel polysilicon 310 -98 310 -98 0 1
rlabel polysilicon 310 -104 310 -104 0 3
rlabel polysilicon 317 -98 317 -98 0 1
rlabel polysilicon 317 -104 317 -104 0 3
rlabel polysilicon 324 -98 324 -98 0 1
rlabel polysilicon 324 -104 324 -104 0 3
rlabel polysilicon 331 -98 331 -98 0 1
rlabel polysilicon 334 -98 334 -98 0 2
rlabel polysilicon 331 -104 331 -104 0 3
rlabel polysilicon 338 -98 338 -98 0 1
rlabel polysilicon 338 -104 338 -104 0 3
rlabel polysilicon 345 -98 345 -98 0 1
rlabel polysilicon 345 -104 345 -104 0 3
rlabel polysilicon 352 -98 352 -98 0 1
rlabel polysilicon 352 -104 352 -104 0 3
rlabel polysilicon 359 -98 359 -98 0 1
rlabel polysilicon 359 -104 359 -104 0 3
rlabel polysilicon 366 -98 366 -98 0 1
rlabel polysilicon 366 -104 366 -104 0 3
rlabel polysilicon 373 -98 373 -98 0 1
rlabel polysilicon 376 -98 376 -98 0 2
rlabel polysilicon 373 -104 373 -104 0 3
rlabel polysilicon 376 -104 376 -104 0 4
rlabel polysilicon 380 -98 380 -98 0 1
rlabel polysilicon 380 -104 380 -104 0 3
rlabel polysilicon 387 -98 387 -98 0 1
rlabel polysilicon 387 -104 387 -104 0 3
rlabel polysilicon 394 -98 394 -98 0 1
rlabel polysilicon 394 -104 394 -104 0 3
rlabel polysilicon 401 -98 401 -98 0 1
rlabel polysilicon 401 -104 401 -104 0 3
rlabel polysilicon 411 -98 411 -98 0 2
rlabel polysilicon 408 -104 408 -104 0 3
rlabel polysilicon 415 -98 415 -98 0 1
rlabel polysilicon 415 -104 415 -104 0 3
rlabel polysilicon 422 -98 422 -98 0 1
rlabel polysilicon 422 -104 422 -104 0 3
rlabel polysilicon 432 -98 432 -98 0 2
rlabel polysilicon 432 -104 432 -104 0 4
rlabel polysilicon 436 -98 436 -98 0 1
rlabel polysilicon 436 -104 436 -104 0 3
rlabel polysilicon 443 -98 443 -98 0 1
rlabel polysilicon 443 -104 443 -104 0 3
rlabel polysilicon 450 -98 450 -98 0 1
rlabel polysilicon 450 -104 450 -104 0 3
rlabel polysilicon 457 -104 457 -104 0 3
rlabel polysilicon 460 -104 460 -104 0 4
rlabel polysilicon 464 -98 464 -98 0 1
rlabel polysilicon 464 -104 464 -104 0 3
rlabel polysilicon 474 -98 474 -98 0 2
rlabel polysilicon 471 -104 471 -104 0 3
rlabel polysilicon 474 -104 474 -104 0 4
rlabel polysilicon 478 -98 478 -98 0 1
rlabel polysilicon 478 -104 478 -104 0 3
rlabel polysilicon 488 -98 488 -98 0 2
rlabel polysilicon 485 -104 485 -104 0 3
rlabel polysilicon 488 -104 488 -104 0 4
rlabel polysilicon 492 -98 492 -98 0 1
rlabel polysilicon 492 -104 492 -104 0 3
rlabel polysilicon 499 -98 499 -98 0 1
rlabel polysilicon 499 -104 499 -104 0 3
rlabel polysilicon 506 -98 506 -98 0 1
rlabel polysilicon 506 -104 506 -104 0 3
rlabel polysilicon 513 -98 513 -98 0 1
rlabel polysilicon 513 -104 513 -104 0 3
rlabel polysilicon 520 -98 520 -98 0 1
rlabel polysilicon 520 -104 520 -104 0 3
rlabel polysilicon 530 -98 530 -98 0 2
rlabel polysilicon 527 -104 527 -104 0 3
rlabel polysilicon 530 -104 530 -104 0 4
rlabel polysilicon 534 -98 534 -98 0 1
rlabel polysilicon 534 -104 534 -104 0 3
rlabel polysilicon 537 -104 537 -104 0 4
rlabel polysilicon 541 -98 541 -98 0 1
rlabel polysilicon 541 -104 541 -104 0 3
rlabel polysilicon 551 -98 551 -98 0 2
rlabel polysilicon 548 -104 548 -104 0 3
rlabel polysilicon 551 -104 551 -104 0 4
rlabel polysilicon 555 -98 555 -98 0 1
rlabel polysilicon 555 -104 555 -104 0 3
rlabel polysilicon 562 -98 562 -98 0 1
rlabel polysilicon 562 -104 562 -104 0 3
rlabel polysilicon 569 -98 569 -98 0 1
rlabel polysilicon 569 -104 569 -104 0 3
rlabel polysilicon 576 -98 576 -98 0 1
rlabel polysilicon 576 -104 576 -104 0 3
rlabel polysilicon 583 -98 583 -98 0 1
rlabel polysilicon 583 -104 583 -104 0 3
rlabel polysilicon 590 -98 590 -98 0 1
rlabel polysilicon 590 -104 590 -104 0 3
rlabel polysilicon 597 -98 597 -98 0 1
rlabel polysilicon 597 -104 597 -104 0 3
rlabel polysilicon 604 -98 604 -98 0 1
rlabel polysilicon 604 -104 604 -104 0 3
rlabel polysilicon 611 -98 611 -98 0 1
rlabel polysilicon 611 -104 611 -104 0 3
rlabel polysilicon 618 -98 618 -98 0 1
rlabel polysilicon 618 -104 618 -104 0 3
rlabel polysilicon 625 -98 625 -98 0 1
rlabel polysilicon 625 -104 625 -104 0 3
rlabel polysilicon 632 -98 632 -98 0 1
rlabel polysilicon 632 -104 632 -104 0 3
rlabel polysilicon 639 -98 639 -98 0 1
rlabel polysilicon 639 -104 639 -104 0 3
rlabel polysilicon 649 -98 649 -98 0 2
rlabel polysilicon 646 -104 646 -104 0 3
rlabel polysilicon 649 -104 649 -104 0 4
rlabel polysilicon 653 -98 653 -98 0 1
rlabel polysilicon 653 -104 653 -104 0 3
rlabel polysilicon 660 -98 660 -98 0 1
rlabel polysilicon 660 -104 660 -104 0 3
rlabel polysilicon 667 -98 667 -98 0 1
rlabel polysilicon 667 -104 667 -104 0 3
rlabel polysilicon 674 -98 674 -98 0 1
rlabel polysilicon 674 -104 674 -104 0 3
rlabel polysilicon 681 -98 681 -98 0 1
rlabel polysilicon 681 -104 681 -104 0 3
rlabel polysilicon 688 -98 688 -98 0 1
rlabel polysilicon 688 -104 688 -104 0 3
rlabel polysilicon 695 -98 695 -98 0 1
rlabel polysilicon 695 -104 695 -104 0 3
rlabel polysilicon 702 -98 702 -98 0 1
rlabel polysilicon 702 -104 702 -104 0 3
rlabel polysilicon 709 -98 709 -98 0 1
rlabel polysilicon 709 -104 709 -104 0 3
rlabel polysilicon 716 -98 716 -98 0 1
rlabel polysilicon 716 -104 716 -104 0 3
rlabel polysilicon 723 -98 723 -98 0 1
rlabel polysilicon 723 -104 723 -104 0 3
rlabel polysilicon 730 -98 730 -98 0 1
rlabel polysilicon 730 -104 730 -104 0 3
rlabel polysilicon 737 -98 737 -98 0 1
rlabel polysilicon 737 -104 737 -104 0 3
rlabel polysilicon 744 -98 744 -98 0 1
rlabel polysilicon 744 -104 744 -104 0 3
rlabel polysilicon 751 -98 751 -98 0 1
rlabel polysilicon 751 -104 751 -104 0 3
rlabel polysilicon 779 -98 779 -98 0 1
rlabel polysilicon 779 -104 779 -104 0 3
rlabel polysilicon 786 -98 786 -98 0 1
rlabel polysilicon 786 -104 786 -104 0 3
rlabel polysilicon 793 -98 793 -98 0 1
rlabel polysilicon 796 -98 796 -98 0 2
rlabel polysilicon 793 -104 793 -104 0 3
rlabel polysilicon 796 -104 796 -104 0 4
rlabel polysilicon 800 -98 800 -98 0 1
rlabel polysilicon 800 -104 800 -104 0 3
rlabel polysilicon 807 -98 807 -98 0 1
rlabel polysilicon 810 -98 810 -98 0 2
rlabel polysilicon 810 -104 810 -104 0 4
rlabel polysilicon 817 -98 817 -98 0 2
rlabel polysilicon 814 -104 814 -104 0 3
rlabel polysilicon 817 -104 817 -104 0 4
rlabel polysilicon 821 -98 821 -98 0 1
rlabel polysilicon 824 -104 824 -104 0 4
rlabel polysilicon 828 -98 828 -98 0 1
rlabel polysilicon 828 -104 828 -104 0 3
rlabel polysilicon 835 -98 835 -98 0 1
rlabel polysilicon 835 -104 835 -104 0 3
rlabel polysilicon 842 -98 842 -98 0 1
rlabel polysilicon 842 -104 842 -104 0 3
rlabel polysilicon 856 -98 856 -98 0 1
rlabel polysilicon 856 -104 856 -104 0 3
rlabel polysilicon 863 -98 863 -98 0 1
rlabel polysilicon 863 -104 863 -104 0 3
rlabel polysilicon 870 -98 870 -98 0 1
rlabel polysilicon 870 -104 870 -104 0 3
rlabel polysilicon 884 -98 884 -98 0 1
rlabel polysilicon 887 -98 887 -98 0 2
rlabel polysilicon 884 -104 884 -104 0 3
rlabel polysilicon 891 -98 891 -98 0 1
rlabel polysilicon 891 -104 891 -104 0 3
rlabel polysilicon 940 -98 940 -98 0 1
rlabel polysilicon 940 -104 940 -104 0 3
rlabel polysilicon 947 -98 947 -98 0 1
rlabel polysilicon 947 -104 947 -104 0 3
rlabel polysilicon 954 -98 954 -98 0 1
rlabel polysilicon 954 -104 954 -104 0 3
rlabel polysilicon 1010 -98 1010 -98 0 1
rlabel polysilicon 1010 -104 1010 -104 0 3
rlabel polysilicon 1087 -98 1087 -98 0 1
rlabel polysilicon 1087 -104 1087 -104 0 3
rlabel polysilicon 93 -167 93 -167 0 1
rlabel polysilicon 93 -173 93 -173 0 3
rlabel polysilicon 114 -167 114 -167 0 1
rlabel polysilicon 114 -173 114 -173 0 3
rlabel polysilicon 135 -167 135 -167 0 1
rlabel polysilicon 135 -173 135 -173 0 3
rlabel polysilicon 142 -167 142 -167 0 1
rlabel polysilicon 142 -173 142 -173 0 3
rlabel polysilicon 149 -167 149 -167 0 1
rlabel polysilicon 149 -173 149 -173 0 3
rlabel polysilicon 156 -167 156 -167 0 1
rlabel polysilicon 156 -173 156 -173 0 3
rlabel polysilicon 163 -167 163 -167 0 1
rlabel polysilicon 163 -173 163 -173 0 3
rlabel polysilicon 170 -167 170 -167 0 1
rlabel polysilicon 170 -173 170 -173 0 3
rlabel polysilicon 177 -167 177 -167 0 1
rlabel polysilicon 177 -173 177 -173 0 3
rlabel polysilicon 184 -167 184 -167 0 1
rlabel polysilicon 184 -173 184 -173 0 3
rlabel polysilicon 191 -167 191 -167 0 1
rlabel polysilicon 191 -173 191 -173 0 3
rlabel polysilicon 198 -167 198 -167 0 1
rlabel polysilicon 198 -173 198 -173 0 3
rlabel polysilicon 208 -167 208 -167 0 2
rlabel polysilicon 208 -173 208 -173 0 4
rlabel polysilicon 215 -173 215 -173 0 4
rlabel polysilicon 219 -167 219 -167 0 1
rlabel polysilicon 219 -173 219 -173 0 3
rlabel polysilicon 226 -167 226 -167 0 1
rlabel polysilicon 226 -173 226 -173 0 3
rlabel polysilicon 233 -173 233 -173 0 3
rlabel polysilicon 236 -173 236 -173 0 4
rlabel polysilicon 243 -167 243 -167 0 2
rlabel polysilicon 240 -173 240 -173 0 3
rlabel polysilicon 243 -173 243 -173 0 4
rlabel polysilicon 247 -167 247 -167 0 1
rlabel polysilicon 247 -173 247 -173 0 3
rlabel polysilicon 254 -167 254 -167 0 1
rlabel polysilicon 254 -173 254 -173 0 3
rlabel polysilicon 261 -167 261 -167 0 1
rlabel polysilicon 261 -173 261 -173 0 3
rlabel polysilicon 268 -167 268 -167 0 1
rlabel polysilicon 268 -173 268 -173 0 3
rlabel polysilicon 275 -167 275 -167 0 1
rlabel polysilicon 275 -173 275 -173 0 3
rlabel polysilicon 282 -167 282 -167 0 1
rlabel polysilicon 282 -173 282 -173 0 3
rlabel polysilicon 289 -167 289 -167 0 1
rlabel polysilicon 289 -173 289 -173 0 3
rlabel polysilicon 296 -167 296 -167 0 1
rlabel polysilicon 296 -173 296 -173 0 3
rlabel polysilicon 303 -167 303 -167 0 1
rlabel polysilicon 303 -173 303 -173 0 3
rlabel polysilicon 310 -167 310 -167 0 1
rlabel polysilicon 310 -173 310 -173 0 3
rlabel polysilicon 317 -167 317 -167 0 1
rlabel polysilicon 317 -173 317 -173 0 3
rlabel polysilicon 324 -167 324 -167 0 1
rlabel polysilicon 324 -173 324 -173 0 3
rlabel polysilicon 331 -167 331 -167 0 1
rlabel polysilicon 331 -173 331 -173 0 3
rlabel polysilicon 338 -167 338 -167 0 1
rlabel polysilicon 338 -173 338 -173 0 3
rlabel polysilicon 345 -167 345 -167 0 1
rlabel polysilicon 345 -173 345 -173 0 3
rlabel polysilicon 352 -167 352 -167 0 1
rlabel polysilicon 355 -167 355 -167 0 2
rlabel polysilicon 352 -173 352 -173 0 3
rlabel polysilicon 359 -167 359 -167 0 1
rlabel polysilicon 362 -167 362 -167 0 2
rlabel polysilicon 359 -173 359 -173 0 3
rlabel polysilicon 362 -173 362 -173 0 4
rlabel polysilicon 366 -167 366 -167 0 1
rlabel polysilicon 366 -173 366 -173 0 3
rlabel polysilicon 373 -167 373 -167 0 1
rlabel polysilicon 373 -173 373 -173 0 3
rlabel polysilicon 380 -167 380 -167 0 1
rlabel polysilicon 380 -173 380 -173 0 3
rlabel polysilicon 387 -167 387 -167 0 1
rlabel polysilicon 387 -173 387 -173 0 3
rlabel polysilicon 394 -167 394 -167 0 1
rlabel polysilicon 394 -173 394 -173 0 3
rlabel polysilicon 401 -167 401 -167 0 1
rlabel polysilicon 401 -173 401 -173 0 3
rlabel polysilicon 408 -167 408 -167 0 1
rlabel polysilicon 408 -173 408 -173 0 3
rlabel polysilicon 415 -167 415 -167 0 1
rlabel polysilicon 415 -173 415 -173 0 3
rlabel polysilicon 422 -167 422 -167 0 1
rlabel polysilicon 422 -173 422 -173 0 3
rlabel polysilicon 429 -167 429 -167 0 1
rlabel polysilicon 432 -167 432 -167 0 2
rlabel polysilicon 432 -173 432 -173 0 4
rlabel polysilicon 436 -167 436 -167 0 1
rlabel polysilicon 436 -173 436 -173 0 3
rlabel polysilicon 443 -167 443 -167 0 1
rlabel polysilicon 443 -173 443 -173 0 3
rlabel polysilicon 450 -167 450 -167 0 1
rlabel polysilicon 450 -173 450 -173 0 3
rlabel polysilicon 457 -167 457 -167 0 1
rlabel polysilicon 457 -173 457 -173 0 3
rlabel polysilicon 464 -167 464 -167 0 1
rlabel polysilicon 467 -167 467 -167 0 2
rlabel polysilicon 464 -173 464 -173 0 3
rlabel polysilicon 471 -167 471 -167 0 1
rlabel polysilicon 471 -173 471 -173 0 3
rlabel polysilicon 478 -167 478 -167 0 1
rlabel polysilicon 481 -167 481 -167 0 2
rlabel polysilicon 481 -173 481 -173 0 4
rlabel polysilicon 485 -167 485 -167 0 1
rlabel polysilicon 485 -173 485 -173 0 3
rlabel polysilicon 492 -167 492 -167 0 1
rlabel polysilicon 492 -173 492 -173 0 3
rlabel polysilicon 499 -167 499 -167 0 1
rlabel polysilicon 502 -167 502 -167 0 2
rlabel polysilicon 499 -173 499 -173 0 3
rlabel polysilicon 502 -173 502 -173 0 4
rlabel polysilicon 506 -167 506 -167 0 1
rlabel polysilicon 509 -167 509 -167 0 2
rlabel polysilicon 509 -173 509 -173 0 4
rlabel polysilicon 513 -167 513 -167 0 1
rlabel polysilicon 513 -173 513 -173 0 3
rlabel polysilicon 516 -173 516 -173 0 4
rlabel polysilicon 520 -167 520 -167 0 1
rlabel polysilicon 520 -173 520 -173 0 3
rlabel polysilicon 523 -173 523 -173 0 4
rlabel polysilicon 527 -167 527 -167 0 1
rlabel polysilicon 527 -173 527 -173 0 3
rlabel polysilicon 534 -167 534 -167 0 1
rlabel polysilicon 534 -173 534 -173 0 3
rlabel polysilicon 541 -167 541 -167 0 1
rlabel polysilicon 541 -173 541 -173 0 3
rlabel polysilicon 544 -173 544 -173 0 4
rlabel polysilicon 548 -167 548 -167 0 1
rlabel polysilicon 548 -173 548 -173 0 3
rlabel polysilicon 555 -167 555 -167 0 1
rlabel polysilicon 555 -173 555 -173 0 3
rlabel polysilicon 562 -167 562 -167 0 1
rlabel polysilicon 562 -173 562 -173 0 3
rlabel polysilicon 569 -167 569 -167 0 1
rlabel polysilicon 569 -173 569 -173 0 3
rlabel polysilicon 576 -167 576 -167 0 1
rlabel polysilicon 576 -173 576 -173 0 3
rlabel polysilicon 583 -167 583 -167 0 1
rlabel polysilicon 583 -173 583 -173 0 3
rlabel polysilicon 590 -167 590 -167 0 1
rlabel polysilicon 590 -173 590 -173 0 3
rlabel polysilicon 597 -167 597 -167 0 1
rlabel polysilicon 597 -173 597 -173 0 3
rlabel polysilicon 604 -167 604 -167 0 1
rlabel polysilicon 604 -173 604 -173 0 3
rlabel polysilicon 611 -167 611 -167 0 1
rlabel polysilicon 611 -173 611 -173 0 3
rlabel polysilicon 614 -173 614 -173 0 4
rlabel polysilicon 618 -167 618 -167 0 1
rlabel polysilicon 618 -173 618 -173 0 3
rlabel polysilicon 625 -167 625 -167 0 1
rlabel polysilicon 625 -173 625 -173 0 3
rlabel polysilicon 632 -167 632 -167 0 1
rlabel polysilicon 632 -173 632 -173 0 3
rlabel polysilicon 639 -167 639 -167 0 1
rlabel polysilicon 639 -173 639 -173 0 3
rlabel polysilicon 646 -167 646 -167 0 1
rlabel polysilicon 646 -173 646 -173 0 3
rlabel polysilicon 653 -167 653 -167 0 1
rlabel polysilicon 656 -167 656 -167 0 2
rlabel polysilicon 653 -173 653 -173 0 3
rlabel polysilicon 656 -173 656 -173 0 4
rlabel polysilicon 660 -167 660 -167 0 1
rlabel polysilicon 660 -173 660 -173 0 3
rlabel polysilicon 667 -167 667 -167 0 1
rlabel polysilicon 667 -173 667 -173 0 3
rlabel polysilicon 674 -167 674 -167 0 1
rlabel polysilicon 674 -173 674 -173 0 3
rlabel polysilicon 681 -167 681 -167 0 1
rlabel polysilicon 681 -173 681 -173 0 3
rlabel polysilicon 688 -167 688 -167 0 1
rlabel polysilicon 688 -173 688 -173 0 3
rlabel polysilicon 698 -167 698 -167 0 2
rlabel polysilicon 695 -173 695 -173 0 3
rlabel polysilicon 698 -173 698 -173 0 4
rlabel polysilicon 702 -167 702 -167 0 1
rlabel polysilicon 702 -173 702 -173 0 3
rlabel polysilicon 709 -167 709 -167 0 1
rlabel polysilicon 709 -173 709 -173 0 3
rlabel polysilicon 716 -167 716 -167 0 1
rlabel polysilicon 716 -173 716 -173 0 3
rlabel polysilicon 723 -167 723 -167 0 1
rlabel polysilicon 723 -173 723 -173 0 3
rlabel polysilicon 730 -167 730 -167 0 1
rlabel polysilicon 730 -173 730 -173 0 3
rlabel polysilicon 737 -167 737 -167 0 1
rlabel polysilicon 737 -173 737 -173 0 3
rlabel polysilicon 744 -167 744 -167 0 1
rlabel polysilicon 744 -173 744 -173 0 3
rlabel polysilicon 751 -167 751 -167 0 1
rlabel polysilicon 751 -173 751 -173 0 3
rlabel polysilicon 758 -167 758 -167 0 1
rlabel polysilicon 758 -173 758 -173 0 3
rlabel polysilicon 768 -167 768 -167 0 2
rlabel polysilicon 765 -173 765 -173 0 3
rlabel polysilicon 768 -173 768 -173 0 4
rlabel polysilicon 772 -167 772 -167 0 1
rlabel polysilicon 772 -173 772 -173 0 3
rlabel polysilicon 779 -167 779 -167 0 1
rlabel polysilicon 779 -173 779 -173 0 3
rlabel polysilicon 786 -167 786 -167 0 1
rlabel polysilicon 786 -173 786 -173 0 3
rlabel polysilicon 793 -167 793 -167 0 1
rlabel polysilicon 793 -173 793 -173 0 3
rlabel polysilicon 796 -173 796 -173 0 4
rlabel polysilicon 800 -167 800 -167 0 1
rlabel polysilicon 800 -173 800 -173 0 3
rlabel polysilicon 807 -167 807 -167 0 1
rlabel polysilicon 807 -173 807 -173 0 3
rlabel polysilicon 814 -167 814 -167 0 1
rlabel polysilicon 814 -173 814 -173 0 3
rlabel polysilicon 821 -167 821 -167 0 1
rlabel polysilicon 828 -167 828 -167 0 1
rlabel polysilicon 828 -173 828 -173 0 3
rlabel polysilicon 835 -167 835 -167 0 1
rlabel polysilicon 835 -173 835 -173 0 3
rlabel polysilicon 842 -167 842 -167 0 1
rlabel polysilicon 842 -173 842 -173 0 3
rlabel polysilicon 849 -167 849 -167 0 1
rlabel polysilicon 849 -173 849 -173 0 3
rlabel polysilicon 856 -167 856 -167 0 1
rlabel polysilicon 856 -173 856 -173 0 3
rlabel polysilicon 863 -167 863 -167 0 1
rlabel polysilicon 863 -173 863 -173 0 3
rlabel polysilicon 870 -167 870 -167 0 1
rlabel polysilicon 870 -173 870 -173 0 3
rlabel polysilicon 877 -167 877 -167 0 1
rlabel polysilicon 880 -167 880 -167 0 2
rlabel polysilicon 880 -173 880 -173 0 4
rlabel polysilicon 887 -167 887 -167 0 2
rlabel polysilicon 887 -173 887 -173 0 4
rlabel polysilicon 891 -167 891 -167 0 1
rlabel polysilicon 891 -173 891 -173 0 3
rlabel polysilicon 898 -167 898 -167 0 1
rlabel polysilicon 898 -173 898 -173 0 3
rlabel polysilicon 905 -167 905 -167 0 1
rlabel polysilicon 905 -173 905 -173 0 3
rlabel polysilicon 912 -167 912 -167 0 1
rlabel polysilicon 912 -173 912 -173 0 3
rlabel polysilicon 919 -167 919 -167 0 1
rlabel polysilicon 919 -173 919 -173 0 3
rlabel polysilicon 926 -167 926 -167 0 1
rlabel polysilicon 926 -173 926 -173 0 3
rlabel polysilicon 933 -167 933 -167 0 1
rlabel polysilicon 933 -173 933 -173 0 3
rlabel polysilicon 940 -167 940 -167 0 1
rlabel polysilicon 940 -173 940 -173 0 3
rlabel polysilicon 947 -167 947 -167 0 1
rlabel polysilicon 947 -173 947 -173 0 3
rlabel polysilicon 954 -167 954 -167 0 1
rlabel polysilicon 954 -173 954 -173 0 3
rlabel polysilicon 961 -167 961 -167 0 1
rlabel polysilicon 961 -173 961 -173 0 3
rlabel polysilicon 968 -167 968 -167 0 1
rlabel polysilicon 968 -173 968 -173 0 3
rlabel polysilicon 975 -167 975 -167 0 1
rlabel polysilicon 975 -173 975 -173 0 3
rlabel polysilicon 982 -167 982 -167 0 1
rlabel polysilicon 982 -173 982 -173 0 3
rlabel polysilicon 996 -167 996 -167 0 1
rlabel polysilicon 996 -173 996 -173 0 3
rlabel polysilicon 1010 -167 1010 -167 0 1
rlabel polysilicon 1010 -173 1010 -173 0 3
rlabel polysilicon 1038 -167 1038 -167 0 1
rlabel polysilicon 1038 -173 1038 -173 0 3
rlabel polysilicon 1129 -167 1129 -167 0 1
rlabel polysilicon 1129 -173 1129 -173 0 3
rlabel polysilicon 1136 -167 1136 -167 0 1
rlabel polysilicon 1136 -173 1136 -173 0 3
rlabel polysilicon 1195 -167 1195 -167 0 2
rlabel polysilicon 1195 -173 1195 -173 0 4
rlabel polysilicon 1220 -167 1220 -167 0 1
rlabel polysilicon 1220 -173 1220 -173 0 3
rlabel polysilicon 51 -254 51 -254 0 1
rlabel polysilicon 51 -260 51 -260 0 3
rlabel polysilicon 58 -254 58 -254 0 1
rlabel polysilicon 58 -260 58 -260 0 3
rlabel polysilicon 65 -254 65 -254 0 1
rlabel polysilicon 65 -260 65 -260 0 3
rlabel polysilicon 72 -254 72 -254 0 1
rlabel polysilicon 72 -260 72 -260 0 3
rlabel polysilicon 79 -254 79 -254 0 1
rlabel polysilicon 79 -260 79 -260 0 3
rlabel polysilicon 86 -254 86 -254 0 1
rlabel polysilicon 86 -260 86 -260 0 3
rlabel polysilicon 93 -254 93 -254 0 1
rlabel polysilicon 93 -260 93 -260 0 3
rlabel polysilicon 100 -254 100 -254 0 1
rlabel polysilicon 100 -260 100 -260 0 3
rlabel polysilicon 107 -254 107 -254 0 1
rlabel polysilicon 107 -260 107 -260 0 3
rlabel polysilicon 117 -254 117 -254 0 2
rlabel polysilicon 117 -260 117 -260 0 4
rlabel polysilicon 121 -254 121 -254 0 1
rlabel polysilicon 121 -260 121 -260 0 3
rlabel polysilicon 128 -254 128 -254 0 1
rlabel polysilicon 128 -260 128 -260 0 3
rlabel polysilicon 135 -254 135 -254 0 1
rlabel polysilicon 135 -260 135 -260 0 3
rlabel polysilicon 142 -254 142 -254 0 1
rlabel polysilicon 142 -260 142 -260 0 3
rlabel polysilicon 149 -254 149 -254 0 1
rlabel polysilicon 149 -260 149 -260 0 3
rlabel polysilicon 156 -254 156 -254 0 1
rlabel polysilicon 156 -260 156 -260 0 3
rlabel polysilicon 163 -254 163 -254 0 1
rlabel polysilicon 163 -260 163 -260 0 3
rlabel polysilicon 170 -254 170 -254 0 1
rlabel polysilicon 173 -260 173 -260 0 4
rlabel polysilicon 177 -254 177 -254 0 1
rlabel polysilicon 177 -260 177 -260 0 3
rlabel polysilicon 184 -254 184 -254 0 1
rlabel polysilicon 184 -260 184 -260 0 3
rlabel polysilicon 191 -254 191 -254 0 1
rlabel polysilicon 191 -260 191 -260 0 3
rlabel polysilicon 194 -260 194 -260 0 4
rlabel polysilicon 201 -254 201 -254 0 2
rlabel polysilicon 198 -260 198 -260 0 3
rlabel polysilicon 205 -254 205 -254 0 1
rlabel polysilicon 205 -260 205 -260 0 3
rlabel polysilicon 212 -254 212 -254 0 1
rlabel polysilicon 215 -260 215 -260 0 4
rlabel polysilicon 219 -254 219 -254 0 1
rlabel polysilicon 219 -260 219 -260 0 3
rlabel polysilicon 226 -254 226 -254 0 1
rlabel polysilicon 226 -260 226 -260 0 3
rlabel polysilicon 233 -254 233 -254 0 1
rlabel polysilicon 236 -254 236 -254 0 2
rlabel polysilicon 233 -260 233 -260 0 3
rlabel polysilicon 236 -260 236 -260 0 4
rlabel polysilicon 243 -254 243 -254 0 2
rlabel polysilicon 243 -260 243 -260 0 4
rlabel polysilicon 247 -254 247 -254 0 1
rlabel polysilicon 247 -260 247 -260 0 3
rlabel polysilicon 254 -254 254 -254 0 1
rlabel polysilicon 254 -260 254 -260 0 3
rlabel polysilicon 261 -254 261 -254 0 1
rlabel polysilicon 261 -260 261 -260 0 3
rlabel polysilicon 268 -254 268 -254 0 1
rlabel polysilicon 268 -260 268 -260 0 3
rlabel polysilicon 275 -254 275 -254 0 1
rlabel polysilicon 275 -260 275 -260 0 3
rlabel polysilicon 282 -254 282 -254 0 1
rlabel polysilicon 282 -260 282 -260 0 3
rlabel polysilicon 289 -254 289 -254 0 1
rlabel polysilicon 292 -254 292 -254 0 2
rlabel polysilicon 289 -260 289 -260 0 3
rlabel polysilicon 296 -254 296 -254 0 1
rlabel polysilicon 296 -260 296 -260 0 3
rlabel polysilicon 303 -254 303 -254 0 1
rlabel polysilicon 303 -260 303 -260 0 3
rlabel polysilicon 310 -254 310 -254 0 1
rlabel polysilicon 310 -260 310 -260 0 3
rlabel polysilicon 317 -254 317 -254 0 1
rlabel polysilicon 317 -260 317 -260 0 3
rlabel polysilicon 324 -254 324 -254 0 1
rlabel polysilicon 324 -260 324 -260 0 3
rlabel polysilicon 331 -254 331 -254 0 1
rlabel polysilicon 331 -260 331 -260 0 3
rlabel polysilicon 338 -254 338 -254 0 1
rlabel polysilicon 338 -260 338 -260 0 3
rlabel polysilicon 345 -254 345 -254 0 1
rlabel polysilicon 345 -260 345 -260 0 3
rlabel polysilicon 352 -254 352 -254 0 1
rlabel polysilicon 352 -260 352 -260 0 3
rlabel polysilicon 359 -254 359 -254 0 1
rlabel polysilicon 359 -260 359 -260 0 3
rlabel polysilicon 366 -254 366 -254 0 1
rlabel polysilicon 366 -260 366 -260 0 3
rlabel polysilicon 373 -254 373 -254 0 1
rlabel polysilicon 373 -260 373 -260 0 3
rlabel polysilicon 380 -254 380 -254 0 1
rlabel polysilicon 383 -254 383 -254 0 2
rlabel polysilicon 383 -260 383 -260 0 4
rlabel polysilicon 387 -254 387 -254 0 1
rlabel polysilicon 387 -260 387 -260 0 3
rlabel polysilicon 394 -254 394 -254 0 1
rlabel polysilicon 394 -260 394 -260 0 3
rlabel polysilicon 401 -254 401 -254 0 1
rlabel polysilicon 401 -260 401 -260 0 3
rlabel polysilicon 408 -254 408 -254 0 1
rlabel polysilicon 408 -260 408 -260 0 3
rlabel polysilicon 415 -254 415 -254 0 1
rlabel polysilicon 415 -260 415 -260 0 3
rlabel polysilicon 422 -254 422 -254 0 1
rlabel polysilicon 422 -260 422 -260 0 3
rlabel polysilicon 429 -254 429 -254 0 1
rlabel polysilicon 429 -260 429 -260 0 3
rlabel polysilicon 436 -254 436 -254 0 1
rlabel polysilicon 436 -260 436 -260 0 3
rlabel polysilicon 443 -254 443 -254 0 1
rlabel polysilicon 446 -254 446 -254 0 2
rlabel polysilicon 443 -260 443 -260 0 3
rlabel polysilicon 450 -254 450 -254 0 1
rlabel polysilicon 450 -260 450 -260 0 3
rlabel polysilicon 457 -254 457 -254 0 1
rlabel polysilicon 460 -254 460 -254 0 2
rlabel polysilicon 457 -260 457 -260 0 3
rlabel polysilicon 460 -260 460 -260 0 4
rlabel polysilicon 467 -254 467 -254 0 2
rlabel polysilicon 467 -260 467 -260 0 4
rlabel polysilicon 471 -254 471 -254 0 1
rlabel polysilicon 474 -254 474 -254 0 2
rlabel polysilicon 471 -260 471 -260 0 3
rlabel polysilicon 474 -260 474 -260 0 4
rlabel polysilicon 478 -254 478 -254 0 1
rlabel polysilicon 478 -260 478 -260 0 3
rlabel polysilicon 485 -254 485 -254 0 1
rlabel polysilicon 485 -260 485 -260 0 3
rlabel polysilicon 495 -254 495 -254 0 2
rlabel polysilicon 492 -260 492 -260 0 3
rlabel polysilicon 495 -260 495 -260 0 4
rlabel polysilicon 499 -254 499 -254 0 1
rlabel polysilicon 499 -260 499 -260 0 3
rlabel polysilicon 506 -254 506 -254 0 1
rlabel polysilicon 509 -254 509 -254 0 2
rlabel polysilicon 506 -260 506 -260 0 3
rlabel polysilicon 509 -260 509 -260 0 4
rlabel polysilicon 513 -254 513 -254 0 1
rlabel polysilicon 513 -260 513 -260 0 3
rlabel polysilicon 520 -254 520 -254 0 1
rlabel polysilicon 520 -260 520 -260 0 3
rlabel polysilicon 530 -254 530 -254 0 2
rlabel polysilicon 527 -260 527 -260 0 3
rlabel polysilicon 530 -260 530 -260 0 4
rlabel polysilicon 534 -254 534 -254 0 1
rlabel polysilicon 534 -260 534 -260 0 3
rlabel polysilicon 541 -254 541 -254 0 1
rlabel polysilicon 544 -254 544 -254 0 2
rlabel polysilicon 544 -260 544 -260 0 4
rlabel polysilicon 548 -254 548 -254 0 1
rlabel polysilicon 548 -260 548 -260 0 3
rlabel polysilicon 555 -254 555 -254 0 1
rlabel polysilicon 555 -260 555 -260 0 3
rlabel polysilicon 562 -254 562 -254 0 1
rlabel polysilicon 562 -260 562 -260 0 3
rlabel polysilicon 569 -254 569 -254 0 1
rlabel polysilicon 572 -254 572 -254 0 2
rlabel polysilicon 569 -260 569 -260 0 3
rlabel polysilicon 572 -260 572 -260 0 4
rlabel polysilicon 579 -254 579 -254 0 2
rlabel polysilicon 576 -260 576 -260 0 3
rlabel polysilicon 579 -260 579 -260 0 4
rlabel polysilicon 583 -254 583 -254 0 1
rlabel polysilicon 583 -260 583 -260 0 3
rlabel polysilicon 590 -254 590 -254 0 1
rlabel polysilicon 593 -254 593 -254 0 2
rlabel polysilicon 593 -260 593 -260 0 4
rlabel polysilicon 597 -254 597 -254 0 1
rlabel polysilicon 597 -260 597 -260 0 3
rlabel polysilicon 604 -254 604 -254 0 1
rlabel polysilicon 604 -260 604 -260 0 3
rlabel polysilicon 611 -254 611 -254 0 1
rlabel polysilicon 614 -254 614 -254 0 2
rlabel polysilicon 611 -260 611 -260 0 3
rlabel polysilicon 614 -260 614 -260 0 4
rlabel polysilicon 618 -254 618 -254 0 1
rlabel polysilicon 618 -260 618 -260 0 3
rlabel polysilicon 625 -254 625 -254 0 1
rlabel polysilicon 625 -260 625 -260 0 3
rlabel polysilicon 632 -254 632 -254 0 1
rlabel polysilicon 632 -260 632 -260 0 3
rlabel polysilicon 639 -254 639 -254 0 1
rlabel polysilicon 639 -260 639 -260 0 3
rlabel polysilicon 646 -254 646 -254 0 1
rlabel polysilicon 646 -260 646 -260 0 3
rlabel polysilicon 653 -254 653 -254 0 1
rlabel polysilicon 653 -260 653 -260 0 3
rlabel polysilicon 660 -254 660 -254 0 1
rlabel polysilicon 660 -260 660 -260 0 3
rlabel polysilicon 667 -254 667 -254 0 1
rlabel polysilicon 667 -260 667 -260 0 3
rlabel polysilicon 674 -254 674 -254 0 1
rlabel polysilicon 674 -260 674 -260 0 3
rlabel polysilicon 681 -254 681 -254 0 1
rlabel polysilicon 681 -260 681 -260 0 3
rlabel polysilicon 688 -254 688 -254 0 1
rlabel polysilicon 688 -260 688 -260 0 3
rlabel polysilicon 695 -254 695 -254 0 1
rlabel polysilicon 695 -260 695 -260 0 3
rlabel polysilicon 702 -254 702 -254 0 1
rlabel polysilicon 702 -260 702 -260 0 3
rlabel polysilicon 709 -254 709 -254 0 1
rlabel polysilicon 709 -260 709 -260 0 3
rlabel polysilicon 719 -254 719 -254 0 2
rlabel polysilicon 716 -260 716 -260 0 3
rlabel polysilicon 723 -254 723 -254 0 1
rlabel polysilicon 723 -260 723 -260 0 3
rlabel polysilicon 730 -254 730 -254 0 1
rlabel polysilicon 730 -260 730 -260 0 3
rlabel polysilicon 737 -254 737 -254 0 1
rlabel polysilicon 737 -260 737 -260 0 3
rlabel polysilicon 744 -254 744 -254 0 1
rlabel polysilicon 744 -260 744 -260 0 3
rlabel polysilicon 751 -254 751 -254 0 1
rlabel polysilicon 751 -260 751 -260 0 3
rlabel polysilicon 758 -254 758 -254 0 1
rlabel polysilicon 758 -260 758 -260 0 3
rlabel polysilicon 765 -254 765 -254 0 1
rlabel polysilicon 765 -260 765 -260 0 3
rlabel polysilicon 772 -254 772 -254 0 1
rlabel polysilicon 779 -254 779 -254 0 1
rlabel polysilicon 779 -260 779 -260 0 3
rlabel polysilicon 789 -254 789 -254 0 2
rlabel polysilicon 786 -260 786 -260 0 3
rlabel polysilicon 789 -260 789 -260 0 4
rlabel polysilicon 793 -254 793 -254 0 1
rlabel polysilicon 793 -260 793 -260 0 3
rlabel polysilicon 800 -254 800 -254 0 1
rlabel polysilicon 800 -260 800 -260 0 3
rlabel polysilicon 807 -254 807 -254 0 1
rlabel polysilicon 807 -260 807 -260 0 3
rlabel polysilicon 814 -254 814 -254 0 1
rlabel polysilicon 814 -260 814 -260 0 3
rlabel polysilicon 821 -254 821 -254 0 1
rlabel polysilicon 821 -260 821 -260 0 3
rlabel polysilicon 831 -254 831 -254 0 2
rlabel polysilicon 828 -260 828 -260 0 3
rlabel polysilicon 835 -254 835 -254 0 1
rlabel polysilicon 835 -260 835 -260 0 3
rlabel polysilicon 842 -254 842 -254 0 1
rlabel polysilicon 842 -260 842 -260 0 3
rlabel polysilicon 849 -254 849 -254 0 1
rlabel polysilicon 849 -260 849 -260 0 3
rlabel polysilicon 856 -254 856 -254 0 1
rlabel polysilicon 856 -260 856 -260 0 3
rlabel polysilicon 863 -254 863 -254 0 1
rlabel polysilicon 863 -260 863 -260 0 3
rlabel polysilicon 870 -254 870 -254 0 1
rlabel polysilicon 870 -260 870 -260 0 3
rlabel polysilicon 877 -254 877 -254 0 1
rlabel polysilicon 877 -260 877 -260 0 3
rlabel polysilicon 884 -254 884 -254 0 1
rlabel polysilicon 884 -260 884 -260 0 3
rlabel polysilicon 891 -254 891 -254 0 1
rlabel polysilicon 891 -260 891 -260 0 3
rlabel polysilicon 898 -254 898 -254 0 1
rlabel polysilicon 898 -260 898 -260 0 3
rlabel polysilicon 905 -254 905 -254 0 1
rlabel polysilicon 905 -260 905 -260 0 3
rlabel polysilicon 912 -254 912 -254 0 1
rlabel polysilicon 912 -260 912 -260 0 3
rlabel polysilicon 919 -254 919 -254 0 1
rlabel polysilicon 919 -260 919 -260 0 3
rlabel polysilicon 926 -254 926 -254 0 1
rlabel polysilicon 926 -260 926 -260 0 3
rlabel polysilicon 933 -254 933 -254 0 1
rlabel polysilicon 933 -260 933 -260 0 3
rlabel polysilicon 940 -254 940 -254 0 1
rlabel polysilicon 940 -260 940 -260 0 3
rlabel polysilicon 947 -254 947 -254 0 1
rlabel polysilicon 947 -260 947 -260 0 3
rlabel polysilicon 954 -254 954 -254 0 1
rlabel polysilicon 954 -260 954 -260 0 3
rlabel polysilicon 961 -254 961 -254 0 1
rlabel polysilicon 961 -260 961 -260 0 3
rlabel polysilicon 968 -254 968 -254 0 1
rlabel polysilicon 968 -260 968 -260 0 3
rlabel polysilicon 975 -254 975 -254 0 1
rlabel polysilicon 975 -260 975 -260 0 3
rlabel polysilicon 982 -254 982 -254 0 1
rlabel polysilicon 982 -260 982 -260 0 3
rlabel polysilicon 989 -254 989 -254 0 1
rlabel polysilicon 989 -260 989 -260 0 3
rlabel polysilicon 996 -254 996 -254 0 1
rlabel polysilicon 999 -254 999 -254 0 2
rlabel polysilicon 999 -260 999 -260 0 4
rlabel polysilicon 1003 -254 1003 -254 0 1
rlabel polysilicon 1003 -260 1003 -260 0 3
rlabel polysilicon 1010 -254 1010 -254 0 1
rlabel polysilicon 1010 -260 1010 -260 0 3
rlabel polysilicon 1017 -254 1017 -254 0 1
rlabel polysilicon 1017 -260 1017 -260 0 3
rlabel polysilicon 1024 -254 1024 -254 0 1
rlabel polysilicon 1024 -260 1024 -260 0 3
rlabel polysilicon 1031 -254 1031 -254 0 1
rlabel polysilicon 1031 -260 1031 -260 0 3
rlabel polysilicon 1038 -254 1038 -254 0 1
rlabel polysilicon 1038 -260 1038 -260 0 3
rlabel polysilicon 1045 -254 1045 -254 0 1
rlabel polysilicon 1045 -260 1045 -260 0 3
rlabel polysilicon 1052 -254 1052 -254 0 1
rlabel polysilicon 1052 -260 1052 -260 0 3
rlabel polysilicon 1059 -254 1059 -254 0 1
rlabel polysilicon 1059 -260 1059 -260 0 3
rlabel polysilicon 1066 -254 1066 -254 0 1
rlabel polysilicon 1066 -260 1066 -260 0 3
rlabel polysilicon 1073 -254 1073 -254 0 1
rlabel polysilicon 1073 -260 1073 -260 0 3
rlabel polysilicon 1080 -254 1080 -254 0 1
rlabel polysilicon 1080 -260 1080 -260 0 3
rlabel polysilicon 1087 -254 1087 -254 0 1
rlabel polysilicon 1087 -260 1087 -260 0 3
rlabel polysilicon 1097 -254 1097 -254 0 2
rlabel polysilicon 1094 -260 1094 -260 0 3
rlabel polysilicon 1097 -260 1097 -260 0 4
rlabel polysilicon 1101 -254 1101 -254 0 1
rlabel polysilicon 1101 -260 1101 -260 0 3
rlabel polysilicon 1108 -254 1108 -254 0 1
rlabel polysilicon 1108 -260 1108 -260 0 3
rlabel polysilicon 1118 -254 1118 -254 0 2
rlabel polysilicon 1115 -260 1115 -260 0 3
rlabel polysilicon 1118 -260 1118 -260 0 4
rlabel polysilicon 1125 -254 1125 -254 0 2
rlabel polysilicon 1122 -260 1122 -260 0 3
rlabel polysilicon 1129 -254 1129 -254 0 1
rlabel polysilicon 1129 -260 1129 -260 0 3
rlabel polysilicon 1136 -254 1136 -254 0 1
rlabel polysilicon 1136 -260 1136 -260 0 3
rlabel polysilicon 1143 -254 1143 -254 0 1
rlabel polysilicon 1143 -260 1143 -260 0 3
rlabel polysilicon 1150 -254 1150 -254 0 1
rlabel polysilicon 1150 -260 1150 -260 0 3
rlabel polysilicon 1157 -254 1157 -254 0 1
rlabel polysilicon 1157 -260 1157 -260 0 3
rlabel polysilicon 1164 -254 1164 -254 0 1
rlabel polysilicon 1164 -260 1164 -260 0 3
rlabel polysilicon 1171 -254 1171 -254 0 1
rlabel polysilicon 1171 -260 1171 -260 0 3
rlabel polysilicon 1227 -254 1227 -254 0 1
rlabel polysilicon 1227 -260 1227 -260 0 3
rlabel polysilicon 1255 -254 1255 -254 0 1
rlabel polysilicon 1255 -260 1255 -260 0 3
rlabel polysilicon 1283 -254 1283 -254 0 1
rlabel polysilicon 1283 -260 1283 -260 0 3
rlabel polysilicon 44 -385 44 -385 0 1
rlabel polysilicon 44 -391 44 -391 0 3
rlabel polysilicon 51 -385 51 -385 0 1
rlabel polysilicon 51 -391 51 -391 0 3
rlabel polysilicon 58 -385 58 -385 0 1
rlabel polysilicon 61 -385 61 -385 0 2
rlabel polysilicon 65 -385 65 -385 0 1
rlabel polysilicon 65 -391 65 -391 0 3
rlabel polysilicon 72 -385 72 -385 0 1
rlabel polysilicon 72 -391 72 -391 0 3
rlabel polysilicon 79 -385 79 -385 0 1
rlabel polysilicon 79 -391 79 -391 0 3
rlabel polysilicon 86 -385 86 -385 0 1
rlabel polysilicon 86 -391 86 -391 0 3
rlabel polysilicon 93 -385 93 -385 0 1
rlabel polysilicon 96 -385 96 -385 0 2
rlabel polysilicon 96 -391 96 -391 0 4
rlabel polysilicon 100 -385 100 -385 0 1
rlabel polysilicon 100 -391 100 -391 0 3
rlabel polysilicon 107 -385 107 -385 0 1
rlabel polysilicon 107 -391 107 -391 0 3
rlabel polysilicon 114 -385 114 -385 0 1
rlabel polysilicon 117 -385 117 -385 0 2
rlabel polysilicon 117 -391 117 -391 0 4
rlabel polysilicon 121 -385 121 -385 0 1
rlabel polysilicon 121 -391 121 -391 0 3
rlabel polysilicon 124 -391 124 -391 0 4
rlabel polysilicon 128 -385 128 -385 0 1
rlabel polysilicon 128 -391 128 -391 0 3
rlabel polysilicon 138 -385 138 -385 0 2
rlabel polysilicon 135 -391 135 -391 0 3
rlabel polysilicon 138 -391 138 -391 0 4
rlabel polysilicon 142 -385 142 -385 0 1
rlabel polysilicon 142 -391 142 -391 0 3
rlabel polysilicon 149 -385 149 -385 0 1
rlabel polysilicon 149 -391 149 -391 0 3
rlabel polysilicon 156 -385 156 -385 0 1
rlabel polysilicon 156 -391 156 -391 0 3
rlabel polysilicon 163 -385 163 -385 0 1
rlabel polysilicon 163 -391 163 -391 0 3
rlabel polysilicon 170 -385 170 -385 0 1
rlabel polysilicon 170 -391 170 -391 0 3
rlabel polysilicon 177 -385 177 -385 0 1
rlabel polysilicon 177 -391 177 -391 0 3
rlabel polysilicon 184 -385 184 -385 0 1
rlabel polysilicon 184 -391 184 -391 0 3
rlabel polysilicon 191 -385 191 -385 0 1
rlabel polysilicon 191 -391 191 -391 0 3
rlabel polysilicon 198 -385 198 -385 0 1
rlabel polysilicon 201 -385 201 -385 0 2
rlabel polysilicon 198 -391 198 -391 0 3
rlabel polysilicon 205 -385 205 -385 0 1
rlabel polysilicon 208 -385 208 -385 0 2
rlabel polysilicon 205 -391 205 -391 0 3
rlabel polysilicon 212 -391 212 -391 0 3
rlabel polysilicon 215 -391 215 -391 0 4
rlabel polysilicon 219 -385 219 -385 0 1
rlabel polysilicon 219 -391 219 -391 0 3
rlabel polysilicon 226 -385 226 -385 0 1
rlabel polysilicon 226 -391 226 -391 0 3
rlabel polysilicon 240 -385 240 -385 0 1
rlabel polysilicon 240 -391 240 -391 0 3
rlabel polysilicon 254 -385 254 -385 0 1
rlabel polysilicon 254 -391 254 -391 0 3
rlabel polysilicon 261 -385 261 -385 0 1
rlabel polysilicon 261 -391 261 -391 0 3
rlabel polysilicon 268 -385 268 -385 0 1
rlabel polysilicon 268 -391 268 -391 0 3
rlabel polysilicon 275 -385 275 -385 0 1
rlabel polysilicon 275 -391 275 -391 0 3
rlabel polysilicon 282 -385 282 -385 0 1
rlabel polysilicon 285 -385 285 -385 0 2
rlabel polysilicon 282 -391 282 -391 0 3
rlabel polysilicon 285 -391 285 -391 0 4
rlabel polysilicon 289 -385 289 -385 0 1
rlabel polysilicon 289 -391 289 -391 0 3
rlabel polysilicon 296 -385 296 -385 0 1
rlabel polysilicon 296 -391 296 -391 0 3
rlabel polysilicon 303 -385 303 -385 0 1
rlabel polysilicon 303 -391 303 -391 0 3
rlabel polysilicon 310 -385 310 -385 0 1
rlabel polysilicon 310 -391 310 -391 0 3
rlabel polysilicon 320 -391 320 -391 0 4
rlabel polysilicon 324 -385 324 -385 0 1
rlabel polysilicon 324 -391 324 -391 0 3
rlabel polysilicon 331 -385 331 -385 0 1
rlabel polysilicon 331 -391 331 -391 0 3
rlabel polysilicon 338 -385 338 -385 0 1
rlabel polysilicon 341 -385 341 -385 0 2
rlabel polysilicon 338 -391 338 -391 0 3
rlabel polysilicon 345 -385 345 -385 0 1
rlabel polysilicon 345 -391 345 -391 0 3
rlabel polysilicon 352 -385 352 -385 0 1
rlabel polysilicon 352 -391 352 -391 0 3
rlabel polysilicon 359 -385 359 -385 0 1
rlabel polysilicon 359 -391 359 -391 0 3
rlabel polysilicon 366 -385 366 -385 0 1
rlabel polysilicon 366 -391 366 -391 0 3
rlabel polysilicon 373 -385 373 -385 0 1
rlabel polysilicon 373 -391 373 -391 0 3
rlabel polysilicon 380 -385 380 -385 0 1
rlabel polysilicon 380 -391 380 -391 0 3
rlabel polysilicon 387 -385 387 -385 0 1
rlabel polysilicon 387 -391 387 -391 0 3
rlabel polysilicon 394 -385 394 -385 0 1
rlabel polysilicon 394 -391 394 -391 0 3
rlabel polysilicon 401 -385 401 -385 0 1
rlabel polysilicon 401 -391 401 -391 0 3
rlabel polysilicon 408 -385 408 -385 0 1
rlabel polysilicon 411 -385 411 -385 0 2
rlabel polysilicon 408 -391 408 -391 0 3
rlabel polysilicon 415 -385 415 -385 0 1
rlabel polysilicon 415 -391 415 -391 0 3
rlabel polysilicon 422 -385 422 -385 0 1
rlabel polysilicon 422 -391 422 -391 0 3
rlabel polysilicon 429 -385 429 -385 0 1
rlabel polysilicon 429 -391 429 -391 0 3
rlabel polysilicon 436 -385 436 -385 0 1
rlabel polysilicon 439 -385 439 -385 0 2
rlabel polysilicon 436 -391 436 -391 0 3
rlabel polysilicon 439 -391 439 -391 0 4
rlabel polysilicon 443 -385 443 -385 0 1
rlabel polysilicon 443 -391 443 -391 0 3
rlabel polysilicon 450 -385 450 -385 0 1
rlabel polysilicon 453 -385 453 -385 0 2
rlabel polysilicon 450 -391 450 -391 0 3
rlabel polysilicon 457 -385 457 -385 0 1
rlabel polysilicon 457 -391 457 -391 0 3
rlabel polysilicon 464 -385 464 -385 0 1
rlabel polysilicon 464 -391 464 -391 0 3
rlabel polysilicon 471 -385 471 -385 0 1
rlabel polysilicon 474 -385 474 -385 0 2
rlabel polysilicon 474 -391 474 -391 0 4
rlabel polysilicon 478 -385 478 -385 0 1
rlabel polysilicon 478 -391 478 -391 0 3
rlabel polysilicon 485 -385 485 -385 0 1
rlabel polysilicon 485 -391 485 -391 0 3
rlabel polysilicon 492 -385 492 -385 0 1
rlabel polysilicon 492 -391 492 -391 0 3
rlabel polysilicon 499 -385 499 -385 0 1
rlabel polysilicon 499 -391 499 -391 0 3
rlabel polysilicon 506 -385 506 -385 0 1
rlabel polysilicon 509 -385 509 -385 0 2
rlabel polysilicon 506 -391 506 -391 0 3
rlabel polysilicon 509 -391 509 -391 0 4
rlabel polysilicon 513 -385 513 -385 0 1
rlabel polysilicon 513 -391 513 -391 0 3
rlabel polysilicon 520 -385 520 -385 0 1
rlabel polysilicon 520 -391 520 -391 0 3
rlabel polysilicon 527 -385 527 -385 0 1
rlabel polysilicon 527 -391 527 -391 0 3
rlabel polysilicon 534 -385 534 -385 0 1
rlabel polysilicon 534 -391 534 -391 0 3
rlabel polysilicon 541 -385 541 -385 0 1
rlabel polysilicon 541 -391 541 -391 0 3
rlabel polysilicon 548 -385 548 -385 0 1
rlabel polysilicon 548 -391 548 -391 0 3
rlabel polysilicon 555 -385 555 -385 0 1
rlabel polysilicon 555 -391 555 -391 0 3
rlabel polysilicon 562 -385 562 -385 0 1
rlabel polysilicon 562 -391 562 -391 0 3
rlabel polysilicon 569 -385 569 -385 0 1
rlabel polysilicon 569 -391 569 -391 0 3
rlabel polysilicon 576 -385 576 -385 0 1
rlabel polysilicon 576 -391 576 -391 0 3
rlabel polysilicon 583 -385 583 -385 0 1
rlabel polysilicon 583 -391 583 -391 0 3
rlabel polysilicon 590 -385 590 -385 0 1
rlabel polysilicon 590 -391 590 -391 0 3
rlabel polysilicon 597 -385 597 -385 0 1
rlabel polysilicon 597 -391 597 -391 0 3
rlabel polysilicon 604 -385 604 -385 0 1
rlabel polysilicon 607 -385 607 -385 0 2
rlabel polysilicon 604 -391 604 -391 0 3
rlabel polysilicon 607 -391 607 -391 0 4
rlabel polysilicon 611 -385 611 -385 0 1
rlabel polysilicon 614 -385 614 -385 0 2
rlabel polysilicon 611 -391 611 -391 0 3
rlabel polysilicon 614 -391 614 -391 0 4
rlabel polysilicon 618 -385 618 -385 0 1
rlabel polysilicon 618 -391 618 -391 0 3
rlabel polysilicon 625 -385 625 -385 0 1
rlabel polysilicon 625 -391 625 -391 0 3
rlabel polysilicon 632 -385 632 -385 0 1
rlabel polysilicon 632 -391 632 -391 0 3
rlabel polysilicon 639 -385 639 -385 0 1
rlabel polysilicon 639 -391 639 -391 0 3
rlabel polysilicon 646 -385 646 -385 0 1
rlabel polysilicon 646 -391 646 -391 0 3
rlabel polysilicon 653 -385 653 -385 0 1
rlabel polysilicon 653 -391 653 -391 0 3
rlabel polysilicon 660 -385 660 -385 0 1
rlabel polysilicon 660 -391 660 -391 0 3
rlabel polysilicon 667 -385 667 -385 0 1
rlabel polysilicon 670 -385 670 -385 0 2
rlabel polysilicon 670 -391 670 -391 0 4
rlabel polysilicon 674 -385 674 -385 0 1
rlabel polysilicon 674 -391 674 -391 0 3
rlabel polysilicon 681 -385 681 -385 0 1
rlabel polysilicon 681 -391 681 -391 0 3
rlabel polysilicon 688 -385 688 -385 0 1
rlabel polysilicon 688 -391 688 -391 0 3
rlabel polysilicon 695 -385 695 -385 0 1
rlabel polysilicon 695 -391 695 -391 0 3
rlabel polysilicon 702 -385 702 -385 0 1
rlabel polysilicon 705 -385 705 -385 0 2
rlabel polysilicon 702 -391 702 -391 0 3
rlabel polysilicon 709 -385 709 -385 0 1
rlabel polysilicon 712 -385 712 -385 0 2
rlabel polysilicon 712 -391 712 -391 0 4
rlabel polysilicon 716 -385 716 -385 0 1
rlabel polysilicon 716 -391 716 -391 0 3
rlabel polysilicon 723 -385 723 -385 0 1
rlabel polysilicon 723 -391 723 -391 0 3
rlabel polysilicon 730 -385 730 -385 0 1
rlabel polysilicon 733 -385 733 -385 0 2
rlabel polysilicon 730 -391 730 -391 0 3
rlabel polysilicon 733 -391 733 -391 0 4
rlabel polysilicon 737 -385 737 -385 0 1
rlabel polysilicon 737 -391 737 -391 0 3
rlabel polysilicon 747 -385 747 -385 0 2
rlabel polysilicon 744 -391 744 -391 0 3
rlabel polysilicon 747 -391 747 -391 0 4
rlabel polysilicon 751 -385 751 -385 0 1
rlabel polysilicon 754 -385 754 -385 0 2
rlabel polysilicon 751 -391 751 -391 0 3
rlabel polysilicon 758 -385 758 -385 0 1
rlabel polysilicon 758 -391 758 -391 0 3
rlabel polysilicon 765 -385 765 -385 0 1
rlabel polysilicon 765 -391 765 -391 0 3
rlabel polysilicon 772 -385 772 -385 0 1
rlabel polysilicon 772 -391 772 -391 0 3
rlabel polysilicon 779 -385 779 -385 0 1
rlabel polysilicon 779 -391 779 -391 0 3
rlabel polysilicon 786 -385 786 -385 0 1
rlabel polysilicon 786 -391 786 -391 0 3
rlabel polysilicon 793 -385 793 -385 0 1
rlabel polysilicon 793 -391 793 -391 0 3
rlabel polysilicon 800 -385 800 -385 0 1
rlabel polysilicon 800 -391 800 -391 0 3
rlabel polysilicon 807 -385 807 -385 0 1
rlabel polysilicon 807 -391 807 -391 0 3
rlabel polysilicon 814 -385 814 -385 0 1
rlabel polysilicon 814 -391 814 -391 0 3
rlabel polysilicon 821 -385 821 -385 0 1
rlabel polysilicon 821 -391 821 -391 0 3
rlabel polysilicon 828 -385 828 -385 0 1
rlabel polysilicon 828 -391 828 -391 0 3
rlabel polysilicon 835 -385 835 -385 0 1
rlabel polysilicon 835 -391 835 -391 0 3
rlabel polysilicon 842 -385 842 -385 0 1
rlabel polysilicon 842 -391 842 -391 0 3
rlabel polysilicon 849 -385 849 -385 0 1
rlabel polysilicon 849 -391 849 -391 0 3
rlabel polysilicon 856 -385 856 -385 0 1
rlabel polysilicon 856 -391 856 -391 0 3
rlabel polysilicon 863 -385 863 -385 0 1
rlabel polysilicon 863 -391 863 -391 0 3
rlabel polysilicon 870 -385 870 -385 0 1
rlabel polysilicon 870 -391 870 -391 0 3
rlabel polysilicon 877 -385 877 -385 0 1
rlabel polysilicon 877 -391 877 -391 0 3
rlabel polysilicon 884 -385 884 -385 0 1
rlabel polysilicon 884 -391 884 -391 0 3
rlabel polysilicon 891 -385 891 -385 0 1
rlabel polysilicon 891 -391 891 -391 0 3
rlabel polysilicon 898 -385 898 -385 0 1
rlabel polysilicon 898 -391 898 -391 0 3
rlabel polysilicon 905 -385 905 -385 0 1
rlabel polysilicon 905 -391 905 -391 0 3
rlabel polysilicon 912 -385 912 -385 0 1
rlabel polysilicon 912 -391 912 -391 0 3
rlabel polysilicon 919 -385 919 -385 0 1
rlabel polysilicon 919 -391 919 -391 0 3
rlabel polysilicon 926 -385 926 -385 0 1
rlabel polysilicon 926 -391 926 -391 0 3
rlabel polysilicon 933 -385 933 -385 0 1
rlabel polysilicon 933 -391 933 -391 0 3
rlabel polysilicon 940 -385 940 -385 0 1
rlabel polysilicon 940 -391 940 -391 0 3
rlabel polysilicon 947 -385 947 -385 0 1
rlabel polysilicon 947 -391 947 -391 0 3
rlabel polysilicon 954 -385 954 -385 0 1
rlabel polysilicon 954 -391 954 -391 0 3
rlabel polysilicon 961 -385 961 -385 0 1
rlabel polysilicon 961 -391 961 -391 0 3
rlabel polysilicon 968 -385 968 -385 0 1
rlabel polysilicon 968 -391 968 -391 0 3
rlabel polysilicon 975 -385 975 -385 0 1
rlabel polysilicon 975 -391 975 -391 0 3
rlabel polysilicon 982 -385 982 -385 0 1
rlabel polysilicon 982 -391 982 -391 0 3
rlabel polysilicon 989 -385 989 -385 0 1
rlabel polysilicon 989 -391 989 -391 0 3
rlabel polysilicon 996 -385 996 -385 0 1
rlabel polysilicon 996 -391 996 -391 0 3
rlabel polysilicon 1003 -385 1003 -385 0 1
rlabel polysilicon 1003 -391 1003 -391 0 3
rlabel polysilicon 1010 -385 1010 -385 0 1
rlabel polysilicon 1010 -391 1010 -391 0 3
rlabel polysilicon 1017 -385 1017 -385 0 1
rlabel polysilicon 1017 -391 1017 -391 0 3
rlabel polysilicon 1024 -385 1024 -385 0 1
rlabel polysilicon 1024 -391 1024 -391 0 3
rlabel polysilicon 1031 -385 1031 -385 0 1
rlabel polysilicon 1031 -391 1031 -391 0 3
rlabel polysilicon 1038 -385 1038 -385 0 1
rlabel polysilicon 1038 -391 1038 -391 0 3
rlabel polysilicon 1045 -385 1045 -385 0 1
rlabel polysilicon 1045 -391 1045 -391 0 3
rlabel polysilicon 1052 -385 1052 -385 0 1
rlabel polysilicon 1052 -391 1052 -391 0 3
rlabel polysilicon 1059 -385 1059 -385 0 1
rlabel polysilicon 1059 -391 1059 -391 0 3
rlabel polysilicon 1066 -385 1066 -385 0 1
rlabel polysilicon 1066 -391 1066 -391 0 3
rlabel polysilicon 1073 -385 1073 -385 0 1
rlabel polysilicon 1073 -391 1073 -391 0 3
rlabel polysilicon 1080 -385 1080 -385 0 1
rlabel polysilicon 1080 -391 1080 -391 0 3
rlabel polysilicon 1087 -385 1087 -385 0 1
rlabel polysilicon 1087 -391 1087 -391 0 3
rlabel polysilicon 1094 -385 1094 -385 0 1
rlabel polysilicon 1094 -391 1094 -391 0 3
rlabel polysilicon 1101 -385 1101 -385 0 1
rlabel polysilicon 1101 -391 1101 -391 0 3
rlabel polysilicon 1108 -385 1108 -385 0 1
rlabel polysilicon 1108 -391 1108 -391 0 3
rlabel polysilicon 1115 -385 1115 -385 0 1
rlabel polysilicon 1115 -391 1115 -391 0 3
rlabel polysilicon 1122 -385 1122 -385 0 1
rlabel polysilicon 1122 -391 1122 -391 0 3
rlabel polysilicon 1129 -385 1129 -385 0 1
rlabel polysilicon 1129 -391 1129 -391 0 3
rlabel polysilicon 1136 -385 1136 -385 0 1
rlabel polysilicon 1136 -391 1136 -391 0 3
rlabel polysilicon 1143 -385 1143 -385 0 1
rlabel polysilicon 1143 -391 1143 -391 0 3
rlabel polysilicon 1150 -385 1150 -385 0 1
rlabel polysilicon 1150 -391 1150 -391 0 3
rlabel polysilicon 1157 -385 1157 -385 0 1
rlabel polysilicon 1157 -391 1157 -391 0 3
rlabel polysilicon 1164 -385 1164 -385 0 1
rlabel polysilicon 1164 -391 1164 -391 0 3
rlabel polysilicon 1171 -385 1171 -385 0 1
rlabel polysilicon 1171 -391 1171 -391 0 3
rlabel polysilicon 1178 -385 1178 -385 0 1
rlabel polysilicon 1178 -391 1178 -391 0 3
rlabel polysilicon 1185 -385 1185 -385 0 1
rlabel polysilicon 1185 -391 1185 -391 0 3
rlabel polysilicon 1192 -385 1192 -385 0 1
rlabel polysilicon 1192 -391 1192 -391 0 3
rlabel polysilicon 1202 -385 1202 -385 0 2
rlabel polysilicon 1199 -391 1199 -391 0 3
rlabel polysilicon 1206 -385 1206 -385 0 1
rlabel polysilicon 1206 -391 1206 -391 0 3
rlabel polysilicon 1213 -385 1213 -385 0 1
rlabel polysilicon 1213 -391 1213 -391 0 3
rlabel polysilicon 1220 -385 1220 -385 0 1
rlabel polysilicon 1220 -391 1220 -391 0 3
rlabel polysilicon 1227 -385 1227 -385 0 1
rlabel polysilicon 1227 -391 1227 -391 0 3
rlabel polysilicon 1234 -385 1234 -385 0 1
rlabel polysilicon 1234 -391 1234 -391 0 3
rlabel polysilicon 1241 -385 1241 -385 0 1
rlabel polysilicon 1241 -391 1241 -391 0 3
rlabel polysilicon 1248 -385 1248 -385 0 1
rlabel polysilicon 1248 -391 1248 -391 0 3
rlabel polysilicon 1255 -385 1255 -385 0 1
rlabel polysilicon 1255 -391 1255 -391 0 3
rlabel polysilicon 1262 -385 1262 -385 0 1
rlabel polysilicon 1262 -391 1262 -391 0 3
rlabel polysilicon 1269 -385 1269 -385 0 1
rlabel polysilicon 1269 -391 1269 -391 0 3
rlabel polysilicon 1276 -385 1276 -385 0 1
rlabel polysilicon 1276 -391 1276 -391 0 3
rlabel polysilicon 1283 -385 1283 -385 0 1
rlabel polysilicon 1283 -391 1283 -391 0 3
rlabel polysilicon 1290 -385 1290 -385 0 1
rlabel polysilicon 1290 -391 1290 -391 0 3
rlabel polysilicon 1297 -385 1297 -385 0 1
rlabel polysilicon 1297 -391 1297 -391 0 3
rlabel polysilicon 1304 -385 1304 -385 0 1
rlabel polysilicon 1304 -391 1304 -391 0 3
rlabel polysilicon 1311 -385 1311 -385 0 1
rlabel polysilicon 1311 -391 1311 -391 0 3
rlabel polysilicon 1318 -385 1318 -385 0 1
rlabel polysilicon 1318 -391 1318 -391 0 3
rlabel polysilicon 1325 -385 1325 -385 0 1
rlabel polysilicon 1325 -391 1325 -391 0 3
rlabel polysilicon 1332 -385 1332 -385 0 1
rlabel polysilicon 1332 -391 1332 -391 0 3
rlabel polysilicon 1339 -385 1339 -385 0 1
rlabel polysilicon 1339 -391 1339 -391 0 3
rlabel polysilicon 1346 -385 1346 -385 0 1
rlabel polysilicon 1346 -391 1346 -391 0 3
rlabel polysilicon 1353 -385 1353 -385 0 1
rlabel polysilicon 1353 -391 1353 -391 0 3
rlabel polysilicon 1360 -385 1360 -385 0 1
rlabel polysilicon 1360 -391 1360 -391 0 3
rlabel polysilicon 1367 -385 1367 -385 0 1
rlabel polysilicon 1367 -391 1367 -391 0 3
rlabel polysilicon 1374 -385 1374 -385 0 1
rlabel polysilicon 1374 -391 1374 -391 0 3
rlabel polysilicon 1381 -385 1381 -385 0 1
rlabel polysilicon 1381 -391 1381 -391 0 3
rlabel polysilicon 1388 -385 1388 -385 0 1
rlabel polysilicon 1388 -391 1388 -391 0 3
rlabel polysilicon 1395 -385 1395 -385 0 1
rlabel polysilicon 1395 -391 1395 -391 0 3
rlabel polysilicon 1398 -391 1398 -391 0 4
rlabel polysilicon 1591 -385 1591 -385 0 1
rlabel polysilicon 1591 -391 1591 -391 0 3
rlabel polysilicon 23 -496 23 -496 0 1
rlabel polysilicon 26 -496 26 -496 0 2
rlabel polysilicon 30 -496 30 -496 0 1
rlabel polysilicon 30 -502 30 -502 0 3
rlabel polysilicon 37 -496 37 -496 0 1
rlabel polysilicon 37 -502 37 -502 0 3
rlabel polysilicon 44 -496 44 -496 0 1
rlabel polysilicon 44 -502 44 -502 0 3
rlabel polysilicon 51 -496 51 -496 0 1
rlabel polysilicon 51 -502 51 -502 0 3
rlabel polysilicon 58 -496 58 -496 0 1
rlabel polysilicon 58 -502 58 -502 0 3
rlabel polysilicon 65 -496 65 -496 0 1
rlabel polysilicon 65 -502 65 -502 0 3
rlabel polysilicon 72 -496 72 -496 0 1
rlabel polysilicon 72 -502 72 -502 0 3
rlabel polysilicon 79 -496 79 -496 0 1
rlabel polysilicon 82 -496 82 -496 0 2
rlabel polysilicon 79 -502 79 -502 0 3
rlabel polysilicon 86 -496 86 -496 0 1
rlabel polysilicon 89 -496 89 -496 0 2
rlabel polysilicon 86 -502 86 -502 0 3
rlabel polysilicon 93 -496 93 -496 0 1
rlabel polysilicon 93 -502 93 -502 0 3
rlabel polysilicon 100 -496 100 -496 0 1
rlabel polysilicon 103 -496 103 -496 0 2
rlabel polysilicon 100 -502 100 -502 0 3
rlabel polysilicon 103 -502 103 -502 0 4
rlabel polysilicon 107 -496 107 -496 0 1
rlabel polysilicon 110 -496 110 -496 0 2
rlabel polysilicon 110 -502 110 -502 0 4
rlabel polysilicon 114 -496 114 -496 0 1
rlabel polysilicon 114 -502 114 -502 0 3
rlabel polysilicon 121 -496 121 -496 0 1
rlabel polysilicon 121 -502 121 -502 0 3
rlabel polysilicon 128 -496 128 -496 0 1
rlabel polysilicon 128 -502 128 -502 0 3
rlabel polysilicon 135 -496 135 -496 0 1
rlabel polysilicon 138 -496 138 -496 0 2
rlabel polysilicon 135 -502 135 -502 0 3
rlabel polysilicon 138 -502 138 -502 0 4
rlabel polysilicon 142 -496 142 -496 0 1
rlabel polysilicon 142 -502 142 -502 0 3
rlabel polysilicon 149 -496 149 -496 0 1
rlabel polysilicon 149 -502 149 -502 0 3
rlabel polysilicon 156 -496 156 -496 0 1
rlabel polysilicon 156 -502 156 -502 0 3
rlabel polysilicon 163 -496 163 -496 0 1
rlabel polysilicon 163 -502 163 -502 0 3
rlabel polysilicon 170 -496 170 -496 0 1
rlabel polysilicon 170 -502 170 -502 0 3
rlabel polysilicon 177 -496 177 -496 0 1
rlabel polysilicon 180 -496 180 -496 0 2
rlabel polysilicon 180 -502 180 -502 0 4
rlabel polysilicon 187 -496 187 -496 0 2
rlabel polysilicon 187 -502 187 -502 0 4
rlabel polysilicon 191 -496 191 -496 0 1
rlabel polysilicon 194 -496 194 -496 0 2
rlabel polysilicon 194 -502 194 -502 0 4
rlabel polysilicon 198 -496 198 -496 0 1
rlabel polysilicon 198 -502 198 -502 0 3
rlabel polysilicon 205 -496 205 -496 0 1
rlabel polysilicon 205 -502 205 -502 0 3
rlabel polysilicon 212 -496 212 -496 0 1
rlabel polysilicon 212 -502 212 -502 0 3
rlabel polysilicon 219 -496 219 -496 0 1
rlabel polysilicon 222 -502 222 -502 0 4
rlabel polysilicon 226 -496 226 -496 0 1
rlabel polysilicon 226 -502 226 -502 0 3
rlabel polysilicon 233 -496 233 -496 0 1
rlabel polysilicon 233 -502 233 -502 0 3
rlabel polysilicon 240 -496 240 -496 0 1
rlabel polysilicon 240 -502 240 -502 0 3
rlabel polysilicon 247 -496 247 -496 0 1
rlabel polysilicon 247 -502 247 -502 0 3
rlabel polysilicon 254 -496 254 -496 0 1
rlabel polysilicon 254 -502 254 -502 0 3
rlabel polysilicon 261 -496 261 -496 0 1
rlabel polysilicon 261 -502 261 -502 0 3
rlabel polysilicon 268 -496 268 -496 0 1
rlabel polysilicon 268 -502 268 -502 0 3
rlabel polysilicon 275 -496 275 -496 0 1
rlabel polysilicon 275 -502 275 -502 0 3
rlabel polysilicon 282 -496 282 -496 0 1
rlabel polysilicon 282 -502 282 -502 0 3
rlabel polysilicon 289 -496 289 -496 0 1
rlabel polysilicon 289 -502 289 -502 0 3
rlabel polysilicon 299 -496 299 -496 0 2
rlabel polysilicon 299 -502 299 -502 0 4
rlabel polysilicon 303 -496 303 -496 0 1
rlabel polysilicon 303 -502 303 -502 0 3
rlabel polysilicon 310 -496 310 -496 0 1
rlabel polysilicon 310 -502 310 -502 0 3
rlabel polysilicon 317 -496 317 -496 0 1
rlabel polysilicon 317 -502 317 -502 0 3
rlabel polysilicon 324 -496 324 -496 0 1
rlabel polysilicon 324 -502 324 -502 0 3
rlabel polysilicon 331 -496 331 -496 0 1
rlabel polysilicon 331 -502 331 -502 0 3
rlabel polysilicon 338 -496 338 -496 0 1
rlabel polysilicon 338 -502 338 -502 0 3
rlabel polysilicon 345 -496 345 -496 0 1
rlabel polysilicon 345 -502 345 -502 0 3
rlabel polysilicon 352 -496 352 -496 0 1
rlabel polysilicon 352 -502 352 -502 0 3
rlabel polysilicon 359 -496 359 -496 0 1
rlabel polysilicon 362 -496 362 -496 0 2
rlabel polysilicon 359 -502 359 -502 0 3
rlabel polysilicon 362 -502 362 -502 0 4
rlabel polysilicon 366 -496 366 -496 0 1
rlabel polysilicon 366 -502 366 -502 0 3
rlabel polysilicon 373 -496 373 -496 0 1
rlabel polysilicon 373 -502 373 -502 0 3
rlabel polysilicon 380 -496 380 -496 0 1
rlabel polysilicon 380 -502 380 -502 0 3
rlabel polysilicon 387 -496 387 -496 0 1
rlabel polysilicon 387 -502 387 -502 0 3
rlabel polysilicon 394 -496 394 -496 0 1
rlabel polysilicon 394 -502 394 -502 0 3
rlabel polysilicon 401 -496 401 -496 0 1
rlabel polysilicon 401 -502 401 -502 0 3
rlabel polysilicon 408 -496 408 -496 0 1
rlabel polysilicon 408 -502 408 -502 0 3
rlabel polysilicon 418 -496 418 -496 0 2
rlabel polysilicon 418 -502 418 -502 0 4
rlabel polysilicon 422 -496 422 -496 0 1
rlabel polysilicon 422 -502 422 -502 0 3
rlabel polysilicon 429 -496 429 -496 0 1
rlabel polysilicon 429 -502 429 -502 0 3
rlabel polysilicon 436 -496 436 -496 0 1
rlabel polysilicon 436 -502 436 -502 0 3
rlabel polysilicon 443 -496 443 -496 0 1
rlabel polysilicon 443 -502 443 -502 0 3
rlabel polysilicon 453 -496 453 -496 0 2
rlabel polysilicon 450 -502 450 -502 0 3
rlabel polysilicon 453 -502 453 -502 0 4
rlabel polysilicon 457 -496 457 -496 0 1
rlabel polysilicon 457 -502 457 -502 0 3
rlabel polysilicon 464 -496 464 -496 0 1
rlabel polysilicon 464 -502 464 -502 0 3
rlabel polysilicon 471 -496 471 -496 0 1
rlabel polysilicon 474 -496 474 -496 0 2
rlabel polysilicon 474 -502 474 -502 0 4
rlabel polysilicon 478 -496 478 -496 0 1
rlabel polysilicon 481 -496 481 -496 0 2
rlabel polysilicon 478 -502 478 -502 0 3
rlabel polysilicon 481 -502 481 -502 0 4
rlabel polysilicon 485 -496 485 -496 0 1
rlabel polysilicon 485 -502 485 -502 0 3
rlabel polysilicon 492 -496 492 -496 0 1
rlabel polysilicon 495 -496 495 -496 0 2
rlabel polysilicon 492 -502 492 -502 0 3
rlabel polysilicon 495 -502 495 -502 0 4
rlabel polysilicon 499 -496 499 -496 0 1
rlabel polysilicon 499 -502 499 -502 0 3
rlabel polysilicon 506 -496 506 -496 0 1
rlabel polysilicon 506 -502 506 -502 0 3
rlabel polysilicon 513 -496 513 -496 0 1
rlabel polysilicon 516 -502 516 -502 0 4
rlabel polysilicon 520 -496 520 -496 0 1
rlabel polysilicon 523 -496 523 -496 0 2
rlabel polysilicon 520 -502 520 -502 0 3
rlabel polysilicon 523 -502 523 -502 0 4
rlabel polysilicon 527 -496 527 -496 0 1
rlabel polysilicon 530 -496 530 -496 0 2
rlabel polysilicon 527 -502 527 -502 0 3
rlabel polysilicon 530 -502 530 -502 0 4
rlabel polysilicon 534 -496 534 -496 0 1
rlabel polysilicon 534 -502 534 -502 0 3
rlabel polysilicon 537 -502 537 -502 0 4
rlabel polysilicon 541 -496 541 -496 0 1
rlabel polysilicon 541 -502 541 -502 0 3
rlabel polysilicon 548 -496 548 -496 0 1
rlabel polysilicon 548 -502 548 -502 0 3
rlabel polysilicon 555 -496 555 -496 0 1
rlabel polysilicon 555 -502 555 -502 0 3
rlabel polysilicon 562 -496 562 -496 0 1
rlabel polysilicon 562 -502 562 -502 0 3
rlabel polysilicon 569 -496 569 -496 0 1
rlabel polysilicon 569 -502 569 -502 0 3
rlabel polysilicon 576 -496 576 -496 0 1
rlabel polysilicon 576 -502 576 -502 0 3
rlabel polysilicon 583 -496 583 -496 0 1
rlabel polysilicon 583 -502 583 -502 0 3
rlabel polysilicon 590 -496 590 -496 0 1
rlabel polysilicon 593 -496 593 -496 0 2
rlabel polysilicon 593 -502 593 -502 0 4
rlabel polysilicon 597 -496 597 -496 0 1
rlabel polysilicon 597 -502 597 -502 0 3
rlabel polysilicon 600 -502 600 -502 0 4
rlabel polysilicon 604 -496 604 -496 0 1
rlabel polysilicon 604 -502 604 -502 0 3
rlabel polysilicon 611 -496 611 -496 0 1
rlabel polysilicon 611 -502 611 -502 0 3
rlabel polysilicon 618 -496 618 -496 0 1
rlabel polysilicon 618 -502 618 -502 0 3
rlabel polysilicon 625 -496 625 -496 0 1
rlabel polysilicon 625 -502 625 -502 0 3
rlabel polysilicon 632 -496 632 -496 0 1
rlabel polysilicon 635 -496 635 -496 0 2
rlabel polysilicon 635 -502 635 -502 0 4
rlabel polysilicon 639 -496 639 -496 0 1
rlabel polysilicon 639 -502 639 -502 0 3
rlabel polysilicon 646 -496 646 -496 0 1
rlabel polysilicon 649 -496 649 -496 0 2
rlabel polysilicon 649 -502 649 -502 0 4
rlabel polysilicon 653 -496 653 -496 0 1
rlabel polysilicon 653 -502 653 -502 0 3
rlabel polysilicon 660 -496 660 -496 0 1
rlabel polysilicon 660 -502 660 -502 0 3
rlabel polysilicon 667 -496 667 -496 0 1
rlabel polysilicon 667 -502 667 -502 0 3
rlabel polysilicon 674 -496 674 -496 0 1
rlabel polysilicon 674 -502 674 -502 0 3
rlabel polysilicon 681 -496 681 -496 0 1
rlabel polysilicon 681 -502 681 -502 0 3
rlabel polysilicon 688 -496 688 -496 0 1
rlabel polysilicon 688 -502 688 -502 0 3
rlabel polysilicon 695 -496 695 -496 0 1
rlabel polysilicon 695 -502 695 -502 0 3
rlabel polysilicon 698 -502 698 -502 0 4
rlabel polysilicon 702 -496 702 -496 0 1
rlabel polysilicon 702 -502 702 -502 0 3
rlabel polysilicon 709 -496 709 -496 0 1
rlabel polysilicon 709 -502 709 -502 0 3
rlabel polysilicon 712 -502 712 -502 0 4
rlabel polysilicon 716 -496 716 -496 0 1
rlabel polysilicon 716 -502 716 -502 0 3
rlabel polysilicon 723 -496 723 -496 0 1
rlabel polysilicon 723 -502 723 -502 0 3
rlabel polysilicon 730 -496 730 -496 0 1
rlabel polysilicon 730 -502 730 -502 0 3
rlabel polysilicon 737 -496 737 -496 0 1
rlabel polysilicon 737 -502 737 -502 0 3
rlabel polysilicon 744 -496 744 -496 0 1
rlabel polysilicon 744 -502 744 -502 0 3
rlabel polysilicon 751 -496 751 -496 0 1
rlabel polysilicon 751 -502 751 -502 0 3
rlabel polysilicon 758 -496 758 -496 0 1
rlabel polysilicon 758 -502 758 -502 0 3
rlabel polysilicon 761 -502 761 -502 0 4
rlabel polysilicon 765 -496 765 -496 0 1
rlabel polysilicon 765 -502 765 -502 0 3
rlabel polysilicon 772 -496 772 -496 0 1
rlabel polysilicon 772 -502 772 -502 0 3
rlabel polysilicon 779 -496 779 -496 0 1
rlabel polysilicon 779 -502 779 -502 0 3
rlabel polysilicon 786 -496 786 -496 0 1
rlabel polysilicon 786 -502 786 -502 0 3
rlabel polysilicon 793 -496 793 -496 0 1
rlabel polysilicon 793 -502 793 -502 0 3
rlabel polysilicon 800 -496 800 -496 0 1
rlabel polysilicon 800 -502 800 -502 0 3
rlabel polysilicon 807 -496 807 -496 0 1
rlabel polysilicon 807 -502 807 -502 0 3
rlabel polysilicon 814 -496 814 -496 0 1
rlabel polysilicon 814 -502 814 -502 0 3
rlabel polysilicon 821 -496 821 -496 0 1
rlabel polysilicon 821 -502 821 -502 0 3
rlabel polysilicon 828 -496 828 -496 0 1
rlabel polysilicon 828 -502 828 -502 0 3
rlabel polysilicon 831 -502 831 -502 0 4
rlabel polysilicon 835 -496 835 -496 0 1
rlabel polysilicon 835 -502 835 -502 0 3
rlabel polysilicon 842 -496 842 -496 0 1
rlabel polysilicon 842 -502 842 -502 0 3
rlabel polysilicon 849 -496 849 -496 0 1
rlabel polysilicon 849 -502 849 -502 0 3
rlabel polysilicon 856 -496 856 -496 0 1
rlabel polysilicon 856 -502 856 -502 0 3
rlabel polysilicon 863 -496 863 -496 0 1
rlabel polysilicon 863 -502 863 -502 0 3
rlabel polysilicon 870 -496 870 -496 0 1
rlabel polysilicon 870 -502 870 -502 0 3
rlabel polysilicon 877 -496 877 -496 0 1
rlabel polysilicon 877 -502 877 -502 0 3
rlabel polysilicon 884 -496 884 -496 0 1
rlabel polysilicon 884 -502 884 -502 0 3
rlabel polysilicon 891 -496 891 -496 0 1
rlabel polysilicon 891 -502 891 -502 0 3
rlabel polysilicon 898 -496 898 -496 0 1
rlabel polysilicon 901 -502 901 -502 0 4
rlabel polysilicon 905 -496 905 -496 0 1
rlabel polysilicon 905 -502 905 -502 0 3
rlabel polysilicon 912 -496 912 -496 0 1
rlabel polysilicon 912 -502 912 -502 0 3
rlabel polysilicon 919 -496 919 -496 0 1
rlabel polysilicon 919 -502 919 -502 0 3
rlabel polysilicon 926 -496 926 -496 0 1
rlabel polysilicon 926 -502 926 -502 0 3
rlabel polysilicon 933 -496 933 -496 0 1
rlabel polysilicon 933 -502 933 -502 0 3
rlabel polysilicon 940 -496 940 -496 0 1
rlabel polysilicon 940 -502 940 -502 0 3
rlabel polysilicon 947 -496 947 -496 0 1
rlabel polysilicon 947 -502 947 -502 0 3
rlabel polysilicon 954 -496 954 -496 0 1
rlabel polysilicon 954 -502 954 -502 0 3
rlabel polysilicon 961 -496 961 -496 0 1
rlabel polysilicon 961 -502 961 -502 0 3
rlabel polysilicon 968 -496 968 -496 0 1
rlabel polysilicon 968 -502 968 -502 0 3
rlabel polysilicon 975 -496 975 -496 0 1
rlabel polysilicon 975 -502 975 -502 0 3
rlabel polysilicon 982 -496 982 -496 0 1
rlabel polysilicon 982 -502 982 -502 0 3
rlabel polysilicon 989 -496 989 -496 0 1
rlabel polysilicon 996 -496 996 -496 0 1
rlabel polysilicon 996 -502 996 -502 0 3
rlabel polysilicon 1003 -496 1003 -496 0 1
rlabel polysilicon 1003 -502 1003 -502 0 3
rlabel polysilicon 1010 -496 1010 -496 0 1
rlabel polysilicon 1010 -502 1010 -502 0 3
rlabel polysilicon 1017 -496 1017 -496 0 1
rlabel polysilicon 1017 -502 1017 -502 0 3
rlabel polysilicon 1024 -496 1024 -496 0 1
rlabel polysilicon 1024 -502 1024 -502 0 3
rlabel polysilicon 1031 -496 1031 -496 0 1
rlabel polysilicon 1031 -502 1031 -502 0 3
rlabel polysilicon 1038 -496 1038 -496 0 1
rlabel polysilicon 1038 -502 1038 -502 0 3
rlabel polysilicon 1045 -496 1045 -496 0 1
rlabel polysilicon 1045 -502 1045 -502 0 3
rlabel polysilicon 1052 -496 1052 -496 0 1
rlabel polysilicon 1052 -502 1052 -502 0 3
rlabel polysilicon 1059 -496 1059 -496 0 1
rlabel polysilicon 1059 -502 1059 -502 0 3
rlabel polysilicon 1066 -496 1066 -496 0 1
rlabel polysilicon 1066 -502 1066 -502 0 3
rlabel polysilicon 1073 -496 1073 -496 0 1
rlabel polysilicon 1073 -502 1073 -502 0 3
rlabel polysilicon 1080 -496 1080 -496 0 1
rlabel polysilicon 1080 -502 1080 -502 0 3
rlabel polysilicon 1087 -496 1087 -496 0 1
rlabel polysilicon 1087 -502 1087 -502 0 3
rlabel polysilicon 1094 -496 1094 -496 0 1
rlabel polysilicon 1094 -502 1094 -502 0 3
rlabel polysilicon 1101 -496 1101 -496 0 1
rlabel polysilicon 1101 -502 1101 -502 0 3
rlabel polysilicon 1108 -496 1108 -496 0 1
rlabel polysilicon 1108 -502 1108 -502 0 3
rlabel polysilicon 1115 -496 1115 -496 0 1
rlabel polysilicon 1115 -502 1115 -502 0 3
rlabel polysilicon 1122 -496 1122 -496 0 1
rlabel polysilicon 1122 -502 1122 -502 0 3
rlabel polysilicon 1129 -496 1129 -496 0 1
rlabel polysilicon 1129 -502 1129 -502 0 3
rlabel polysilicon 1136 -496 1136 -496 0 1
rlabel polysilicon 1136 -502 1136 -502 0 3
rlabel polysilicon 1143 -496 1143 -496 0 1
rlabel polysilicon 1143 -502 1143 -502 0 3
rlabel polysilicon 1150 -496 1150 -496 0 1
rlabel polysilicon 1150 -502 1150 -502 0 3
rlabel polysilicon 1157 -496 1157 -496 0 1
rlabel polysilicon 1157 -502 1157 -502 0 3
rlabel polysilicon 1164 -496 1164 -496 0 1
rlabel polysilicon 1164 -502 1164 -502 0 3
rlabel polysilicon 1171 -496 1171 -496 0 1
rlabel polysilicon 1171 -502 1171 -502 0 3
rlabel polysilicon 1178 -496 1178 -496 0 1
rlabel polysilicon 1178 -502 1178 -502 0 3
rlabel polysilicon 1185 -496 1185 -496 0 1
rlabel polysilicon 1185 -502 1185 -502 0 3
rlabel polysilicon 1195 -502 1195 -502 0 4
rlabel polysilicon 1199 -496 1199 -496 0 1
rlabel polysilicon 1199 -502 1199 -502 0 3
rlabel polysilicon 1206 -496 1206 -496 0 1
rlabel polysilicon 1206 -502 1206 -502 0 3
rlabel polysilicon 1213 -496 1213 -496 0 1
rlabel polysilicon 1213 -502 1213 -502 0 3
rlabel polysilicon 1220 -496 1220 -496 0 1
rlabel polysilicon 1220 -502 1220 -502 0 3
rlabel polysilicon 1227 -496 1227 -496 0 1
rlabel polysilicon 1227 -502 1227 -502 0 3
rlabel polysilicon 1234 -496 1234 -496 0 1
rlabel polysilicon 1234 -502 1234 -502 0 3
rlabel polysilicon 1241 -496 1241 -496 0 1
rlabel polysilicon 1241 -502 1241 -502 0 3
rlabel polysilicon 1248 -496 1248 -496 0 1
rlabel polysilicon 1248 -502 1248 -502 0 3
rlabel polysilicon 1255 -496 1255 -496 0 1
rlabel polysilicon 1255 -502 1255 -502 0 3
rlabel polysilicon 1262 -496 1262 -496 0 1
rlabel polysilicon 1262 -502 1262 -502 0 3
rlabel polysilicon 1269 -496 1269 -496 0 1
rlabel polysilicon 1269 -502 1269 -502 0 3
rlabel polysilicon 1272 -502 1272 -502 0 4
rlabel polysilicon 1276 -496 1276 -496 0 1
rlabel polysilicon 1276 -502 1276 -502 0 3
rlabel polysilicon 1283 -496 1283 -496 0 1
rlabel polysilicon 1283 -502 1283 -502 0 3
rlabel polysilicon 1290 -496 1290 -496 0 1
rlabel polysilicon 1290 -502 1290 -502 0 3
rlabel polysilicon 1297 -496 1297 -496 0 1
rlabel polysilicon 1297 -502 1297 -502 0 3
rlabel polysilicon 1304 -496 1304 -496 0 1
rlabel polysilicon 1304 -502 1304 -502 0 3
rlabel polysilicon 1311 -496 1311 -496 0 1
rlabel polysilicon 1311 -502 1311 -502 0 3
rlabel polysilicon 1318 -496 1318 -496 0 1
rlabel polysilicon 1318 -502 1318 -502 0 3
rlabel polysilicon 1325 -496 1325 -496 0 1
rlabel polysilicon 1325 -502 1325 -502 0 3
rlabel polysilicon 1332 -496 1332 -496 0 1
rlabel polysilicon 1332 -502 1332 -502 0 3
rlabel polysilicon 1339 -496 1339 -496 0 1
rlabel polysilicon 1339 -502 1339 -502 0 3
rlabel polysilicon 1346 -496 1346 -496 0 1
rlabel polysilicon 1346 -502 1346 -502 0 3
rlabel polysilicon 1353 -496 1353 -496 0 1
rlabel polysilicon 1353 -502 1353 -502 0 3
rlabel polysilicon 1360 -496 1360 -496 0 1
rlabel polysilicon 1360 -502 1360 -502 0 3
rlabel polysilicon 1367 -496 1367 -496 0 1
rlabel polysilicon 1367 -502 1367 -502 0 3
rlabel polysilicon 1374 -496 1374 -496 0 1
rlabel polysilicon 1374 -502 1374 -502 0 3
rlabel polysilicon 1381 -496 1381 -496 0 1
rlabel polysilicon 1381 -502 1381 -502 0 3
rlabel polysilicon 1388 -496 1388 -496 0 1
rlabel polysilicon 1388 -502 1388 -502 0 3
rlabel polysilicon 1395 -496 1395 -496 0 1
rlabel polysilicon 1395 -502 1395 -502 0 3
rlabel polysilicon 1402 -496 1402 -496 0 1
rlabel polysilicon 1402 -502 1402 -502 0 3
rlabel polysilicon 1409 -496 1409 -496 0 1
rlabel polysilicon 1409 -502 1409 -502 0 3
rlabel polysilicon 1416 -496 1416 -496 0 1
rlabel polysilicon 1416 -502 1416 -502 0 3
rlabel polysilicon 1423 -496 1423 -496 0 1
rlabel polysilicon 1423 -502 1423 -502 0 3
rlabel polysilicon 1430 -496 1430 -496 0 1
rlabel polysilicon 1430 -502 1430 -502 0 3
rlabel polysilicon 1437 -496 1437 -496 0 1
rlabel polysilicon 1437 -502 1437 -502 0 3
rlabel polysilicon 1444 -496 1444 -496 0 1
rlabel polysilicon 1444 -502 1444 -502 0 3
rlabel polysilicon 1451 -496 1451 -496 0 1
rlabel polysilicon 1451 -502 1451 -502 0 3
rlabel polysilicon 1458 -496 1458 -496 0 1
rlabel polysilicon 1458 -502 1458 -502 0 3
rlabel polysilicon 1465 -496 1465 -496 0 1
rlabel polysilicon 1465 -502 1465 -502 0 3
rlabel polysilicon 1472 -496 1472 -496 0 1
rlabel polysilicon 1472 -502 1472 -502 0 3
rlabel polysilicon 1479 -496 1479 -496 0 1
rlabel polysilicon 1479 -502 1479 -502 0 3
rlabel polysilicon 1486 -496 1486 -496 0 1
rlabel polysilicon 1486 -502 1486 -502 0 3
rlabel polysilicon 1493 -496 1493 -496 0 1
rlabel polysilicon 1493 -502 1493 -502 0 3
rlabel polysilicon 1500 -496 1500 -496 0 1
rlabel polysilicon 1500 -502 1500 -502 0 3
rlabel polysilicon 1503 -502 1503 -502 0 4
rlabel polysilicon 1507 -496 1507 -496 0 1
rlabel polysilicon 1507 -502 1507 -502 0 3
rlabel polysilicon 1514 -496 1514 -496 0 1
rlabel polysilicon 1514 -502 1514 -502 0 3
rlabel polysilicon 1524 -496 1524 -496 0 2
rlabel polysilicon 1528 -496 1528 -496 0 1
rlabel polysilicon 1528 -502 1528 -502 0 3
rlabel polysilicon 1710 -496 1710 -496 0 1
rlabel polysilicon 1710 -502 1710 -502 0 3
rlabel polysilicon 9 -603 9 -603 0 1
rlabel polysilicon 9 -609 9 -609 0 3
rlabel polysilicon 23 -603 23 -603 0 1
rlabel polysilicon 23 -609 23 -609 0 3
rlabel polysilicon 30 -603 30 -603 0 1
rlabel polysilicon 30 -609 30 -609 0 3
rlabel polysilicon 44 -603 44 -603 0 1
rlabel polysilicon 44 -609 44 -609 0 3
rlabel polysilicon 51 -603 51 -603 0 1
rlabel polysilicon 51 -609 51 -609 0 3
rlabel polysilicon 61 -603 61 -603 0 2
rlabel polysilicon 58 -609 58 -609 0 3
rlabel polysilicon 61 -609 61 -609 0 4
rlabel polysilicon 65 -603 65 -603 0 1
rlabel polysilicon 65 -609 65 -609 0 3
rlabel polysilicon 72 -603 72 -603 0 1
rlabel polysilicon 72 -609 72 -609 0 3
rlabel polysilicon 79 -603 79 -603 0 1
rlabel polysilicon 79 -609 79 -609 0 3
rlabel polysilicon 86 -603 86 -603 0 1
rlabel polysilicon 86 -609 86 -609 0 3
rlabel polysilicon 93 -603 93 -603 0 1
rlabel polysilicon 93 -609 93 -609 0 3
rlabel polysilicon 103 -603 103 -603 0 2
rlabel polysilicon 100 -609 100 -609 0 3
rlabel polysilicon 103 -609 103 -609 0 4
rlabel polysilicon 107 -603 107 -603 0 1
rlabel polysilicon 114 -603 114 -603 0 1
rlabel polysilicon 114 -609 114 -609 0 3
rlabel polysilicon 121 -603 121 -603 0 1
rlabel polysilicon 121 -609 121 -609 0 3
rlabel polysilicon 128 -603 128 -603 0 1
rlabel polysilicon 128 -609 128 -609 0 3
rlabel polysilicon 135 -603 135 -603 0 1
rlabel polysilicon 135 -609 135 -609 0 3
rlabel polysilicon 142 -603 142 -603 0 1
rlabel polysilicon 142 -609 142 -609 0 3
rlabel polysilicon 149 -603 149 -603 0 1
rlabel polysilicon 152 -603 152 -603 0 2
rlabel polysilicon 149 -609 149 -609 0 3
rlabel polysilicon 152 -609 152 -609 0 4
rlabel polysilicon 156 -603 156 -603 0 1
rlabel polysilicon 156 -609 156 -609 0 3
rlabel polysilicon 163 -603 163 -603 0 1
rlabel polysilicon 163 -609 163 -609 0 3
rlabel polysilicon 170 -603 170 -603 0 1
rlabel polysilicon 170 -609 170 -609 0 3
rlabel polysilicon 177 -603 177 -603 0 1
rlabel polysilicon 177 -609 177 -609 0 3
rlabel polysilicon 184 -603 184 -603 0 1
rlabel polysilicon 184 -609 184 -609 0 3
rlabel polysilicon 187 -609 187 -609 0 4
rlabel polysilicon 191 -603 191 -603 0 1
rlabel polysilicon 191 -609 191 -609 0 3
rlabel polysilicon 198 -603 198 -603 0 1
rlabel polysilicon 198 -609 198 -609 0 3
rlabel polysilicon 205 -603 205 -603 0 1
rlabel polysilicon 205 -609 205 -609 0 3
rlabel polysilicon 212 -603 212 -603 0 1
rlabel polysilicon 212 -609 212 -609 0 3
rlabel polysilicon 219 -603 219 -603 0 1
rlabel polysilicon 219 -609 219 -609 0 3
rlabel polysilicon 226 -603 226 -603 0 1
rlabel polysilicon 226 -609 226 -609 0 3
rlabel polysilicon 233 -609 233 -609 0 3
rlabel polysilicon 236 -609 236 -609 0 4
rlabel polysilicon 240 -603 240 -603 0 1
rlabel polysilicon 243 -603 243 -603 0 2
rlabel polysilicon 240 -609 240 -609 0 3
rlabel polysilicon 243 -609 243 -609 0 4
rlabel polysilicon 247 -603 247 -603 0 1
rlabel polysilicon 247 -609 247 -609 0 3
rlabel polysilicon 254 -603 254 -603 0 1
rlabel polysilicon 254 -609 254 -609 0 3
rlabel polysilicon 261 -603 261 -603 0 1
rlabel polysilicon 261 -609 261 -609 0 3
rlabel polysilicon 268 -603 268 -603 0 1
rlabel polysilicon 268 -609 268 -609 0 3
rlabel polysilicon 275 -603 275 -603 0 1
rlabel polysilicon 275 -609 275 -609 0 3
rlabel polysilicon 282 -603 282 -603 0 1
rlabel polysilicon 282 -609 282 -609 0 3
rlabel polysilicon 289 -603 289 -603 0 1
rlabel polysilicon 289 -609 289 -609 0 3
rlabel polysilicon 296 -603 296 -603 0 1
rlabel polysilicon 296 -609 296 -609 0 3
rlabel polysilicon 303 -603 303 -603 0 1
rlabel polysilicon 303 -609 303 -609 0 3
rlabel polysilicon 310 -603 310 -603 0 1
rlabel polysilicon 310 -609 310 -609 0 3
rlabel polysilicon 317 -603 317 -603 0 1
rlabel polysilicon 320 -609 320 -609 0 4
rlabel polysilicon 324 -603 324 -603 0 1
rlabel polysilicon 324 -609 324 -609 0 3
rlabel polysilicon 331 -603 331 -603 0 1
rlabel polysilicon 331 -609 331 -609 0 3
rlabel polysilicon 338 -603 338 -603 0 1
rlabel polysilicon 341 -603 341 -603 0 2
rlabel polysilicon 338 -609 338 -609 0 3
rlabel polysilicon 345 -603 345 -603 0 1
rlabel polysilicon 345 -609 345 -609 0 3
rlabel polysilicon 352 -603 352 -603 0 1
rlabel polysilicon 352 -609 352 -609 0 3
rlabel polysilicon 359 -603 359 -603 0 1
rlabel polysilicon 359 -609 359 -609 0 3
rlabel polysilicon 366 -603 366 -603 0 1
rlabel polysilicon 366 -609 366 -609 0 3
rlabel polysilicon 373 -603 373 -603 0 1
rlabel polysilicon 373 -609 373 -609 0 3
rlabel polysilicon 383 -609 383 -609 0 4
rlabel polysilicon 387 -603 387 -603 0 1
rlabel polysilicon 387 -609 387 -609 0 3
rlabel polysilicon 394 -603 394 -603 0 1
rlabel polysilicon 394 -609 394 -609 0 3
rlabel polysilicon 401 -603 401 -603 0 1
rlabel polysilicon 401 -609 401 -609 0 3
rlabel polysilicon 408 -603 408 -603 0 1
rlabel polysilicon 408 -609 408 -609 0 3
rlabel polysilicon 415 -603 415 -603 0 1
rlabel polysilicon 415 -609 415 -609 0 3
rlabel polysilicon 422 -603 422 -603 0 1
rlabel polysilicon 422 -609 422 -609 0 3
rlabel polysilicon 429 -609 429 -609 0 3
rlabel polysilicon 432 -609 432 -609 0 4
rlabel polysilicon 436 -603 436 -603 0 1
rlabel polysilicon 436 -609 436 -609 0 3
rlabel polysilicon 443 -603 443 -603 0 1
rlabel polysilicon 443 -609 443 -609 0 3
rlabel polysilicon 450 -603 450 -603 0 1
rlabel polysilicon 453 -603 453 -603 0 2
rlabel polysilicon 450 -609 450 -609 0 3
rlabel polysilicon 453 -609 453 -609 0 4
rlabel polysilicon 457 -603 457 -603 0 1
rlabel polysilicon 460 -603 460 -603 0 2
rlabel polysilicon 457 -609 457 -609 0 3
rlabel polysilicon 464 -603 464 -603 0 1
rlabel polysilicon 464 -609 464 -609 0 3
rlabel polysilicon 471 -603 471 -603 0 1
rlabel polysilicon 471 -609 471 -609 0 3
rlabel polysilicon 478 -603 478 -603 0 1
rlabel polysilicon 478 -609 478 -609 0 3
rlabel polysilicon 485 -603 485 -603 0 1
rlabel polysilicon 485 -609 485 -609 0 3
rlabel polysilicon 492 -603 492 -603 0 1
rlabel polysilicon 492 -609 492 -609 0 3
rlabel polysilicon 499 -603 499 -603 0 1
rlabel polysilicon 499 -609 499 -609 0 3
rlabel polysilicon 506 -603 506 -603 0 1
rlabel polysilicon 506 -609 506 -609 0 3
rlabel polysilicon 513 -603 513 -603 0 1
rlabel polysilicon 516 -603 516 -603 0 2
rlabel polysilicon 513 -609 513 -609 0 3
rlabel polysilicon 520 -603 520 -603 0 1
rlabel polysilicon 520 -609 520 -609 0 3
rlabel polysilicon 527 -603 527 -603 0 1
rlabel polysilicon 530 -603 530 -603 0 2
rlabel polysilicon 527 -609 527 -609 0 3
rlabel polysilicon 530 -609 530 -609 0 4
rlabel polysilicon 534 -603 534 -603 0 1
rlabel polysilicon 534 -609 534 -609 0 3
rlabel polysilicon 541 -603 541 -603 0 1
rlabel polysilicon 541 -609 541 -609 0 3
rlabel polysilicon 548 -603 548 -603 0 1
rlabel polysilicon 548 -609 548 -609 0 3
rlabel polysilicon 555 -603 555 -603 0 1
rlabel polysilicon 555 -609 555 -609 0 3
rlabel polysilicon 562 -603 562 -603 0 1
rlabel polysilicon 562 -609 562 -609 0 3
rlabel polysilicon 569 -603 569 -603 0 1
rlabel polysilicon 569 -609 569 -609 0 3
rlabel polysilicon 576 -603 576 -603 0 1
rlabel polysilicon 579 -603 579 -603 0 2
rlabel polysilicon 576 -609 576 -609 0 3
rlabel polysilicon 583 -603 583 -603 0 1
rlabel polysilicon 586 -603 586 -603 0 2
rlabel polysilicon 586 -609 586 -609 0 4
rlabel polysilicon 590 -603 590 -603 0 1
rlabel polysilicon 593 -603 593 -603 0 2
rlabel polysilicon 590 -609 590 -609 0 3
rlabel polysilicon 593 -609 593 -609 0 4
rlabel polysilicon 597 -603 597 -603 0 1
rlabel polysilicon 597 -609 597 -609 0 3
rlabel polysilicon 604 -603 604 -603 0 1
rlabel polysilicon 604 -609 604 -609 0 3
rlabel polysilicon 611 -603 611 -603 0 1
rlabel polysilicon 611 -609 611 -609 0 3
rlabel polysilicon 618 -603 618 -603 0 1
rlabel polysilicon 618 -609 618 -609 0 3
rlabel polysilicon 625 -603 625 -603 0 1
rlabel polysilicon 625 -609 625 -609 0 3
rlabel polysilicon 632 -603 632 -603 0 1
rlabel polysilicon 635 -603 635 -603 0 2
rlabel polysilicon 635 -609 635 -609 0 4
rlabel polysilicon 639 -603 639 -603 0 1
rlabel polysilicon 639 -609 639 -609 0 3
rlabel polysilicon 646 -603 646 -603 0 1
rlabel polysilicon 646 -609 646 -609 0 3
rlabel polysilicon 653 -603 653 -603 0 1
rlabel polysilicon 653 -609 653 -609 0 3
rlabel polysilicon 656 -609 656 -609 0 4
rlabel polysilicon 660 -603 660 -603 0 1
rlabel polysilicon 660 -609 660 -609 0 3
rlabel polysilicon 667 -603 667 -603 0 1
rlabel polysilicon 667 -609 667 -609 0 3
rlabel polysilicon 674 -603 674 -603 0 1
rlabel polysilicon 677 -603 677 -603 0 2
rlabel polysilicon 677 -609 677 -609 0 4
rlabel polysilicon 681 -603 681 -603 0 1
rlabel polysilicon 681 -609 681 -609 0 3
rlabel polysilicon 688 -603 688 -603 0 1
rlabel polysilicon 688 -609 688 -609 0 3
rlabel polysilicon 698 -603 698 -603 0 2
rlabel polysilicon 695 -609 695 -609 0 3
rlabel polysilicon 698 -609 698 -609 0 4
rlabel polysilicon 702 -603 702 -603 0 1
rlabel polysilicon 702 -609 702 -609 0 3
rlabel polysilicon 709 -603 709 -603 0 1
rlabel polysilicon 709 -609 709 -609 0 3
rlabel polysilicon 716 -603 716 -603 0 1
rlabel polysilicon 716 -609 716 -609 0 3
rlabel polysilicon 723 -603 723 -603 0 1
rlabel polysilicon 723 -609 723 -609 0 3
rlabel polysilicon 730 -603 730 -603 0 1
rlabel polysilicon 730 -609 730 -609 0 3
rlabel polysilicon 737 -603 737 -603 0 1
rlabel polysilicon 737 -609 737 -609 0 3
rlabel polysilicon 744 -603 744 -603 0 1
rlabel polysilicon 744 -609 744 -609 0 3
rlabel polysilicon 751 -603 751 -603 0 1
rlabel polysilicon 751 -609 751 -609 0 3
rlabel polysilicon 758 -603 758 -603 0 1
rlabel polysilicon 758 -609 758 -609 0 3
rlabel polysilicon 765 -603 765 -603 0 1
rlabel polysilicon 765 -609 765 -609 0 3
rlabel polysilicon 772 -603 772 -603 0 1
rlabel polysilicon 772 -609 772 -609 0 3
rlabel polysilicon 779 -603 779 -603 0 1
rlabel polysilicon 779 -609 779 -609 0 3
rlabel polysilicon 786 -603 786 -603 0 1
rlabel polysilicon 786 -609 786 -609 0 3
rlabel polysilicon 793 -603 793 -603 0 1
rlabel polysilicon 793 -609 793 -609 0 3
rlabel polysilicon 800 -603 800 -603 0 1
rlabel polysilicon 800 -609 800 -609 0 3
rlabel polysilicon 807 -603 807 -603 0 1
rlabel polysilicon 807 -609 807 -609 0 3
rlabel polysilicon 814 -603 814 -603 0 1
rlabel polysilicon 814 -609 814 -609 0 3
rlabel polysilicon 821 -603 821 -603 0 1
rlabel polysilicon 824 -603 824 -603 0 2
rlabel polysilicon 821 -609 821 -609 0 3
rlabel polysilicon 824 -609 824 -609 0 4
rlabel polysilicon 828 -603 828 -603 0 1
rlabel polysilicon 828 -609 828 -609 0 3
rlabel polysilicon 835 -603 835 -603 0 1
rlabel polysilicon 835 -609 835 -609 0 3
rlabel polysilicon 842 -603 842 -603 0 1
rlabel polysilicon 845 -603 845 -603 0 2
rlabel polysilicon 842 -609 842 -609 0 3
rlabel polysilicon 849 -603 849 -603 0 1
rlabel polysilicon 852 -603 852 -603 0 2
rlabel polysilicon 849 -609 849 -609 0 3
rlabel polysilicon 852 -609 852 -609 0 4
rlabel polysilicon 856 -603 856 -603 0 1
rlabel polysilicon 856 -609 856 -609 0 3
rlabel polysilicon 866 -603 866 -603 0 2
rlabel polysilicon 863 -609 863 -609 0 3
rlabel polysilicon 866 -609 866 -609 0 4
rlabel polysilicon 873 -603 873 -603 0 2
rlabel polysilicon 870 -609 870 -609 0 3
rlabel polysilicon 873 -609 873 -609 0 4
rlabel polysilicon 877 -603 877 -603 0 1
rlabel polysilicon 877 -609 877 -609 0 3
rlabel polysilicon 884 -603 884 -603 0 1
rlabel polysilicon 884 -609 884 -609 0 3
rlabel polysilicon 891 -603 891 -603 0 1
rlabel polysilicon 894 -603 894 -603 0 2
rlabel polysilicon 894 -609 894 -609 0 4
rlabel polysilicon 898 -609 898 -609 0 3
rlabel polysilicon 905 -603 905 -603 0 1
rlabel polysilicon 905 -609 905 -609 0 3
rlabel polysilicon 912 -603 912 -603 0 1
rlabel polysilicon 915 -603 915 -603 0 2
rlabel polysilicon 915 -609 915 -609 0 4
rlabel polysilicon 919 -603 919 -603 0 1
rlabel polysilicon 919 -609 919 -609 0 3
rlabel polysilicon 926 -603 926 -603 0 1
rlabel polysilicon 926 -609 926 -609 0 3
rlabel polysilicon 933 -609 933 -609 0 3
rlabel polysilicon 940 -603 940 -603 0 1
rlabel polysilicon 940 -609 940 -609 0 3
rlabel polysilicon 947 -603 947 -603 0 1
rlabel polysilicon 947 -609 947 -609 0 3
rlabel polysilicon 954 -603 954 -603 0 1
rlabel polysilicon 954 -609 954 -609 0 3
rlabel polysilicon 961 -603 961 -603 0 1
rlabel polysilicon 961 -609 961 -609 0 3
rlabel polysilicon 968 -603 968 -603 0 1
rlabel polysilicon 968 -609 968 -609 0 3
rlabel polysilicon 975 -603 975 -603 0 1
rlabel polysilicon 975 -609 975 -609 0 3
rlabel polysilicon 982 -603 982 -603 0 1
rlabel polysilicon 982 -609 982 -609 0 3
rlabel polysilicon 989 -609 989 -609 0 3
rlabel polysilicon 996 -603 996 -603 0 1
rlabel polysilicon 996 -609 996 -609 0 3
rlabel polysilicon 1003 -603 1003 -603 0 1
rlabel polysilicon 1003 -609 1003 -609 0 3
rlabel polysilicon 1010 -603 1010 -603 0 1
rlabel polysilicon 1010 -609 1010 -609 0 3
rlabel polysilicon 1017 -603 1017 -603 0 1
rlabel polysilicon 1017 -609 1017 -609 0 3
rlabel polysilicon 1024 -603 1024 -603 0 1
rlabel polysilicon 1024 -609 1024 -609 0 3
rlabel polysilicon 1031 -603 1031 -603 0 1
rlabel polysilicon 1031 -609 1031 -609 0 3
rlabel polysilicon 1038 -603 1038 -603 0 1
rlabel polysilicon 1038 -609 1038 -609 0 3
rlabel polysilicon 1045 -603 1045 -603 0 1
rlabel polysilicon 1045 -609 1045 -609 0 3
rlabel polysilicon 1052 -603 1052 -603 0 1
rlabel polysilicon 1055 -603 1055 -603 0 2
rlabel polysilicon 1059 -603 1059 -603 0 1
rlabel polysilicon 1059 -609 1059 -609 0 3
rlabel polysilicon 1066 -603 1066 -603 0 1
rlabel polysilicon 1066 -609 1066 -609 0 3
rlabel polysilicon 1073 -603 1073 -603 0 1
rlabel polysilicon 1073 -609 1073 -609 0 3
rlabel polysilicon 1080 -603 1080 -603 0 1
rlabel polysilicon 1080 -609 1080 -609 0 3
rlabel polysilicon 1087 -603 1087 -603 0 1
rlabel polysilicon 1087 -609 1087 -609 0 3
rlabel polysilicon 1094 -603 1094 -603 0 1
rlabel polysilicon 1094 -609 1094 -609 0 3
rlabel polysilicon 1101 -603 1101 -603 0 1
rlabel polysilicon 1101 -609 1101 -609 0 3
rlabel polysilicon 1108 -603 1108 -603 0 1
rlabel polysilicon 1108 -609 1108 -609 0 3
rlabel polysilicon 1115 -603 1115 -603 0 1
rlabel polysilicon 1115 -609 1115 -609 0 3
rlabel polysilicon 1122 -603 1122 -603 0 1
rlabel polysilicon 1122 -609 1122 -609 0 3
rlabel polysilicon 1129 -603 1129 -603 0 1
rlabel polysilicon 1129 -609 1129 -609 0 3
rlabel polysilicon 1136 -603 1136 -603 0 1
rlabel polysilicon 1136 -609 1136 -609 0 3
rlabel polysilicon 1143 -603 1143 -603 0 1
rlabel polysilicon 1143 -609 1143 -609 0 3
rlabel polysilicon 1150 -603 1150 -603 0 1
rlabel polysilicon 1150 -609 1150 -609 0 3
rlabel polysilicon 1157 -603 1157 -603 0 1
rlabel polysilicon 1157 -609 1157 -609 0 3
rlabel polysilicon 1164 -603 1164 -603 0 1
rlabel polysilicon 1164 -609 1164 -609 0 3
rlabel polysilicon 1171 -603 1171 -603 0 1
rlabel polysilicon 1171 -609 1171 -609 0 3
rlabel polysilicon 1178 -603 1178 -603 0 1
rlabel polysilicon 1178 -609 1178 -609 0 3
rlabel polysilicon 1185 -603 1185 -603 0 1
rlabel polysilicon 1185 -609 1185 -609 0 3
rlabel polysilicon 1192 -603 1192 -603 0 1
rlabel polysilicon 1192 -609 1192 -609 0 3
rlabel polysilicon 1199 -603 1199 -603 0 1
rlabel polysilicon 1199 -609 1199 -609 0 3
rlabel polysilicon 1206 -603 1206 -603 0 1
rlabel polysilicon 1206 -609 1206 -609 0 3
rlabel polysilicon 1213 -603 1213 -603 0 1
rlabel polysilicon 1213 -609 1213 -609 0 3
rlabel polysilicon 1220 -603 1220 -603 0 1
rlabel polysilicon 1220 -609 1220 -609 0 3
rlabel polysilicon 1227 -603 1227 -603 0 1
rlabel polysilicon 1227 -609 1227 -609 0 3
rlabel polysilicon 1234 -603 1234 -603 0 1
rlabel polysilicon 1234 -609 1234 -609 0 3
rlabel polysilicon 1241 -603 1241 -603 0 1
rlabel polysilicon 1241 -609 1241 -609 0 3
rlabel polysilicon 1248 -603 1248 -603 0 1
rlabel polysilicon 1248 -609 1248 -609 0 3
rlabel polysilicon 1255 -603 1255 -603 0 1
rlabel polysilicon 1255 -609 1255 -609 0 3
rlabel polysilicon 1262 -603 1262 -603 0 1
rlabel polysilicon 1262 -609 1262 -609 0 3
rlabel polysilicon 1269 -603 1269 -603 0 1
rlabel polysilicon 1272 -603 1272 -603 0 2
rlabel polysilicon 1269 -609 1269 -609 0 3
rlabel polysilicon 1276 -603 1276 -603 0 1
rlabel polysilicon 1276 -609 1276 -609 0 3
rlabel polysilicon 1283 -603 1283 -603 0 1
rlabel polysilicon 1283 -609 1283 -609 0 3
rlabel polysilicon 1290 -603 1290 -603 0 1
rlabel polysilicon 1290 -609 1290 -609 0 3
rlabel polysilicon 1297 -603 1297 -603 0 1
rlabel polysilicon 1297 -609 1297 -609 0 3
rlabel polysilicon 1304 -603 1304 -603 0 1
rlabel polysilicon 1304 -609 1304 -609 0 3
rlabel polysilicon 1311 -603 1311 -603 0 1
rlabel polysilicon 1311 -609 1311 -609 0 3
rlabel polysilicon 1318 -603 1318 -603 0 1
rlabel polysilicon 1318 -609 1318 -609 0 3
rlabel polysilicon 1325 -603 1325 -603 0 1
rlabel polysilicon 1325 -609 1325 -609 0 3
rlabel polysilicon 1332 -603 1332 -603 0 1
rlabel polysilicon 1332 -609 1332 -609 0 3
rlabel polysilicon 1339 -603 1339 -603 0 1
rlabel polysilicon 1339 -609 1339 -609 0 3
rlabel polysilicon 1346 -603 1346 -603 0 1
rlabel polysilicon 1346 -609 1346 -609 0 3
rlabel polysilicon 1353 -603 1353 -603 0 1
rlabel polysilicon 1353 -609 1353 -609 0 3
rlabel polysilicon 1360 -603 1360 -603 0 1
rlabel polysilicon 1360 -609 1360 -609 0 3
rlabel polysilicon 1367 -603 1367 -603 0 1
rlabel polysilicon 1367 -609 1367 -609 0 3
rlabel polysilicon 1374 -603 1374 -603 0 1
rlabel polysilicon 1374 -609 1374 -609 0 3
rlabel polysilicon 1381 -603 1381 -603 0 1
rlabel polysilicon 1381 -609 1381 -609 0 3
rlabel polysilicon 1388 -603 1388 -603 0 1
rlabel polysilicon 1388 -609 1388 -609 0 3
rlabel polysilicon 1395 -603 1395 -603 0 1
rlabel polysilicon 1395 -609 1395 -609 0 3
rlabel polysilicon 1402 -603 1402 -603 0 1
rlabel polysilicon 1402 -609 1402 -609 0 3
rlabel polysilicon 1409 -603 1409 -603 0 1
rlabel polysilicon 1409 -609 1409 -609 0 3
rlabel polysilicon 1416 -603 1416 -603 0 1
rlabel polysilicon 1416 -609 1416 -609 0 3
rlabel polysilicon 1423 -603 1423 -603 0 1
rlabel polysilicon 1423 -609 1423 -609 0 3
rlabel polysilicon 1430 -603 1430 -603 0 1
rlabel polysilicon 1430 -609 1430 -609 0 3
rlabel polysilicon 1437 -603 1437 -603 0 1
rlabel polysilicon 1437 -609 1437 -609 0 3
rlabel polysilicon 1444 -603 1444 -603 0 1
rlabel polysilicon 1444 -609 1444 -609 0 3
rlabel polysilicon 1451 -603 1451 -603 0 1
rlabel polysilicon 1451 -609 1451 -609 0 3
rlabel polysilicon 1458 -603 1458 -603 0 1
rlabel polysilicon 1458 -609 1458 -609 0 3
rlabel polysilicon 1468 -603 1468 -603 0 2
rlabel polysilicon 1465 -609 1465 -609 0 3
rlabel polysilicon 1468 -609 1468 -609 0 4
rlabel polysilicon 1472 -603 1472 -603 0 1
rlabel polysilicon 1472 -609 1472 -609 0 3
rlabel polysilicon 1479 -603 1479 -603 0 1
rlabel polysilicon 1479 -609 1479 -609 0 3
rlabel polysilicon 1486 -603 1486 -603 0 1
rlabel polysilicon 1486 -609 1486 -609 0 3
rlabel polysilicon 1493 -603 1493 -603 0 1
rlabel polysilicon 1493 -609 1493 -609 0 3
rlabel polysilicon 1500 -603 1500 -603 0 1
rlabel polysilicon 1503 -603 1503 -603 0 2
rlabel polysilicon 1500 -609 1500 -609 0 3
rlabel polysilicon 1507 -603 1507 -603 0 1
rlabel polysilicon 1507 -609 1507 -609 0 3
rlabel polysilicon 1514 -603 1514 -603 0 1
rlabel polysilicon 1514 -609 1514 -609 0 3
rlabel polysilicon 1521 -603 1521 -603 0 1
rlabel polysilicon 1521 -609 1521 -609 0 3
rlabel polysilicon 1535 -603 1535 -603 0 1
rlabel polysilicon 1535 -609 1535 -609 0 3
rlabel polysilicon 1556 -603 1556 -603 0 1
rlabel polysilicon 1556 -609 1556 -609 0 3
rlabel polysilicon 1738 -603 1738 -603 0 1
rlabel polysilicon 1738 -609 1738 -609 0 3
rlabel polysilicon 1759 -603 1759 -603 0 1
rlabel polysilicon 1759 -609 1759 -609 0 3
rlabel polysilicon 1766 -603 1766 -603 0 1
rlabel polysilicon 1766 -609 1766 -609 0 3
rlabel polysilicon 9 -712 9 -712 0 1
rlabel polysilicon 9 -718 9 -718 0 3
rlabel polysilicon 16 -712 16 -712 0 1
rlabel polysilicon 16 -718 16 -718 0 3
rlabel polysilicon 23 -712 23 -712 0 1
rlabel polysilicon 23 -718 23 -718 0 3
rlabel polysilicon 30 -712 30 -712 0 1
rlabel polysilicon 30 -718 30 -718 0 3
rlabel polysilicon 37 -712 37 -712 0 1
rlabel polysilicon 37 -718 37 -718 0 3
rlabel polysilicon 44 -712 44 -712 0 1
rlabel polysilicon 44 -718 44 -718 0 3
rlabel polysilicon 51 -712 51 -712 0 1
rlabel polysilicon 51 -718 51 -718 0 3
rlabel polysilicon 58 -712 58 -712 0 1
rlabel polysilicon 58 -718 58 -718 0 3
rlabel polysilicon 65 -712 65 -712 0 1
rlabel polysilicon 65 -718 65 -718 0 3
rlabel polysilicon 72 -712 72 -712 0 1
rlabel polysilicon 72 -718 72 -718 0 3
rlabel polysilicon 79 -712 79 -712 0 1
rlabel polysilicon 79 -718 79 -718 0 3
rlabel polysilicon 86 -712 86 -712 0 1
rlabel polysilicon 86 -718 86 -718 0 3
rlabel polysilicon 96 -712 96 -712 0 2
rlabel polysilicon 93 -718 93 -718 0 3
rlabel polysilicon 96 -718 96 -718 0 4
rlabel polysilicon 100 -712 100 -712 0 1
rlabel polysilicon 100 -718 100 -718 0 3
rlabel polysilicon 107 -718 107 -718 0 3
rlabel polysilicon 114 -712 114 -712 0 1
rlabel polysilicon 117 -712 117 -712 0 2
rlabel polysilicon 114 -718 114 -718 0 3
rlabel polysilicon 117 -718 117 -718 0 4
rlabel polysilicon 121 -712 121 -712 0 1
rlabel polysilicon 121 -718 121 -718 0 3
rlabel polysilicon 128 -712 128 -712 0 1
rlabel polysilicon 128 -718 128 -718 0 3
rlabel polysilicon 135 -712 135 -712 0 1
rlabel polysilicon 135 -718 135 -718 0 3
rlabel polysilicon 138 -718 138 -718 0 4
rlabel polysilicon 142 -712 142 -712 0 1
rlabel polysilicon 145 -712 145 -712 0 2
rlabel polysilicon 142 -718 142 -718 0 3
rlabel polysilicon 145 -718 145 -718 0 4
rlabel polysilicon 149 -712 149 -712 0 1
rlabel polysilicon 149 -718 149 -718 0 3
rlabel polysilicon 156 -712 156 -712 0 1
rlabel polysilicon 156 -718 156 -718 0 3
rlabel polysilicon 163 -712 163 -712 0 1
rlabel polysilicon 163 -718 163 -718 0 3
rlabel polysilicon 170 -712 170 -712 0 1
rlabel polysilicon 173 -712 173 -712 0 2
rlabel polysilicon 170 -718 170 -718 0 3
rlabel polysilicon 173 -718 173 -718 0 4
rlabel polysilicon 177 -712 177 -712 0 1
rlabel polysilicon 177 -718 177 -718 0 3
rlabel polysilicon 184 -718 184 -718 0 3
rlabel polysilicon 187 -718 187 -718 0 4
rlabel polysilicon 191 -712 191 -712 0 1
rlabel polysilicon 191 -718 191 -718 0 3
rlabel polysilicon 198 -712 198 -712 0 1
rlabel polysilicon 198 -718 198 -718 0 3
rlabel polysilicon 205 -712 205 -712 0 1
rlabel polysilicon 205 -718 205 -718 0 3
rlabel polysilicon 212 -712 212 -712 0 1
rlabel polysilicon 212 -718 212 -718 0 3
rlabel polysilicon 219 -712 219 -712 0 1
rlabel polysilicon 219 -718 219 -718 0 3
rlabel polysilicon 226 -712 226 -712 0 1
rlabel polysilicon 226 -718 226 -718 0 3
rlabel polysilicon 236 -712 236 -712 0 2
rlabel polysilicon 233 -718 233 -718 0 3
rlabel polysilicon 240 -712 240 -712 0 1
rlabel polysilicon 240 -718 240 -718 0 3
rlabel polysilicon 247 -712 247 -712 0 1
rlabel polysilicon 247 -718 247 -718 0 3
rlabel polysilicon 254 -712 254 -712 0 1
rlabel polysilicon 254 -718 254 -718 0 3
rlabel polysilicon 261 -712 261 -712 0 1
rlabel polysilicon 261 -718 261 -718 0 3
rlabel polysilicon 268 -712 268 -712 0 1
rlabel polysilicon 268 -718 268 -718 0 3
rlabel polysilicon 275 -712 275 -712 0 1
rlabel polysilicon 275 -718 275 -718 0 3
rlabel polysilicon 282 -712 282 -712 0 1
rlabel polysilicon 282 -718 282 -718 0 3
rlabel polysilicon 289 -712 289 -712 0 1
rlabel polysilicon 289 -718 289 -718 0 3
rlabel polysilicon 296 -712 296 -712 0 1
rlabel polysilicon 296 -718 296 -718 0 3
rlabel polysilicon 303 -712 303 -712 0 1
rlabel polysilicon 303 -718 303 -718 0 3
rlabel polysilicon 310 -712 310 -712 0 1
rlabel polysilicon 310 -718 310 -718 0 3
rlabel polysilicon 317 -712 317 -712 0 1
rlabel polysilicon 324 -712 324 -712 0 1
rlabel polysilicon 324 -718 324 -718 0 3
rlabel polysilicon 331 -712 331 -712 0 1
rlabel polysilicon 331 -718 331 -718 0 3
rlabel polysilicon 338 -712 338 -712 0 1
rlabel polysilicon 338 -718 338 -718 0 3
rlabel polysilicon 345 -712 345 -712 0 1
rlabel polysilicon 345 -718 345 -718 0 3
rlabel polysilicon 352 -712 352 -712 0 1
rlabel polysilicon 352 -718 352 -718 0 3
rlabel polysilicon 359 -712 359 -712 0 1
rlabel polysilicon 362 -712 362 -712 0 2
rlabel polysilicon 359 -718 359 -718 0 3
rlabel polysilicon 366 -712 366 -712 0 1
rlabel polysilicon 366 -718 366 -718 0 3
rlabel polysilicon 373 -712 373 -712 0 1
rlabel polysilicon 373 -718 373 -718 0 3
rlabel polysilicon 380 -712 380 -712 0 1
rlabel polysilicon 380 -718 380 -718 0 3
rlabel polysilicon 387 -712 387 -712 0 1
rlabel polysilicon 387 -718 387 -718 0 3
rlabel polysilicon 394 -712 394 -712 0 1
rlabel polysilicon 394 -718 394 -718 0 3
rlabel polysilicon 401 -712 401 -712 0 1
rlabel polysilicon 401 -718 401 -718 0 3
rlabel polysilicon 408 -712 408 -712 0 1
rlabel polysilicon 408 -718 408 -718 0 3
rlabel polysilicon 415 -712 415 -712 0 1
rlabel polysilicon 415 -718 415 -718 0 3
rlabel polysilicon 422 -712 422 -712 0 1
rlabel polysilicon 422 -718 422 -718 0 3
rlabel polysilicon 429 -712 429 -712 0 1
rlabel polysilicon 429 -718 429 -718 0 3
rlabel polysilicon 436 -712 436 -712 0 1
rlabel polysilicon 436 -718 436 -718 0 3
rlabel polysilicon 443 -712 443 -712 0 1
rlabel polysilicon 443 -718 443 -718 0 3
rlabel polysilicon 450 -712 450 -712 0 1
rlabel polysilicon 450 -718 450 -718 0 3
rlabel polysilicon 457 -712 457 -712 0 1
rlabel polysilicon 457 -718 457 -718 0 3
rlabel polysilicon 464 -712 464 -712 0 1
rlabel polysilicon 467 -712 467 -712 0 2
rlabel polysilicon 464 -718 464 -718 0 3
rlabel polysilicon 467 -718 467 -718 0 4
rlabel polysilicon 471 -712 471 -712 0 1
rlabel polysilicon 471 -718 471 -718 0 3
rlabel polysilicon 478 -712 478 -712 0 1
rlabel polysilicon 481 -712 481 -712 0 2
rlabel polysilicon 478 -718 478 -718 0 3
rlabel polysilicon 485 -712 485 -712 0 1
rlabel polysilicon 485 -718 485 -718 0 3
rlabel polysilicon 492 -712 492 -712 0 1
rlabel polysilicon 492 -718 492 -718 0 3
rlabel polysilicon 499 -712 499 -712 0 1
rlabel polysilicon 499 -718 499 -718 0 3
rlabel polysilicon 506 -712 506 -712 0 1
rlabel polysilicon 509 -712 509 -712 0 2
rlabel polysilicon 509 -718 509 -718 0 4
rlabel polysilicon 513 -712 513 -712 0 1
rlabel polysilicon 513 -718 513 -718 0 3
rlabel polysilicon 520 -712 520 -712 0 1
rlabel polysilicon 520 -718 520 -718 0 3
rlabel polysilicon 527 -712 527 -712 0 1
rlabel polysilicon 527 -718 527 -718 0 3
rlabel polysilicon 534 -712 534 -712 0 1
rlabel polysilicon 534 -718 534 -718 0 3
rlabel polysilicon 541 -712 541 -712 0 1
rlabel polysilicon 544 -712 544 -712 0 2
rlabel polysilicon 544 -718 544 -718 0 4
rlabel polysilicon 548 -712 548 -712 0 1
rlabel polysilicon 548 -718 548 -718 0 3
rlabel polysilicon 555 -718 555 -718 0 3
rlabel polysilicon 558 -718 558 -718 0 4
rlabel polysilicon 562 -712 562 -712 0 1
rlabel polysilicon 562 -718 562 -718 0 3
rlabel polysilicon 569 -712 569 -712 0 1
rlabel polysilicon 569 -718 569 -718 0 3
rlabel polysilicon 576 -712 576 -712 0 1
rlabel polysilicon 576 -718 576 -718 0 3
rlabel polysilicon 583 -712 583 -712 0 1
rlabel polysilicon 583 -718 583 -718 0 3
rlabel polysilicon 590 -712 590 -712 0 1
rlabel polysilicon 590 -718 590 -718 0 3
rlabel polysilicon 597 -712 597 -712 0 1
rlabel polysilicon 600 -712 600 -712 0 2
rlabel polysilicon 600 -718 600 -718 0 4
rlabel polysilicon 604 -712 604 -712 0 1
rlabel polysilicon 604 -718 604 -718 0 3
rlabel polysilicon 611 -712 611 -712 0 1
rlabel polysilicon 611 -718 611 -718 0 3
rlabel polysilicon 618 -712 618 -712 0 1
rlabel polysilicon 621 -712 621 -712 0 2
rlabel polysilicon 618 -718 618 -718 0 3
rlabel polysilicon 621 -718 621 -718 0 4
rlabel polysilicon 625 -712 625 -712 0 1
rlabel polysilicon 625 -718 625 -718 0 3
rlabel polysilicon 632 -712 632 -712 0 1
rlabel polysilicon 632 -718 632 -718 0 3
rlabel polysilicon 639 -712 639 -712 0 1
rlabel polysilicon 639 -718 639 -718 0 3
rlabel polysilicon 646 -712 646 -712 0 1
rlabel polysilicon 649 -712 649 -712 0 2
rlabel polysilicon 646 -718 646 -718 0 3
rlabel polysilicon 649 -718 649 -718 0 4
rlabel polysilicon 653 -712 653 -712 0 1
rlabel polysilicon 656 -712 656 -712 0 2
rlabel polysilicon 653 -718 653 -718 0 3
rlabel polysilicon 660 -712 660 -712 0 1
rlabel polysilicon 660 -718 660 -718 0 3
rlabel polysilicon 667 -712 667 -712 0 1
rlabel polysilicon 667 -718 667 -718 0 3
rlabel polysilicon 674 -712 674 -712 0 1
rlabel polysilicon 674 -718 674 -718 0 3
rlabel polysilicon 681 -712 681 -712 0 1
rlabel polysilicon 681 -718 681 -718 0 3
rlabel polysilicon 691 -712 691 -712 0 2
rlabel polysilicon 688 -718 688 -718 0 3
rlabel polysilicon 695 -712 695 -712 0 1
rlabel polysilicon 695 -718 695 -718 0 3
rlabel polysilicon 702 -712 702 -712 0 1
rlabel polysilicon 702 -718 702 -718 0 3
rlabel polysilicon 709 -712 709 -712 0 1
rlabel polysilicon 712 -712 712 -712 0 2
rlabel polysilicon 709 -718 709 -718 0 3
rlabel polysilicon 712 -718 712 -718 0 4
rlabel polysilicon 719 -712 719 -712 0 2
rlabel polysilicon 716 -718 716 -718 0 3
rlabel polysilicon 719 -718 719 -718 0 4
rlabel polysilicon 723 -712 723 -712 0 1
rlabel polysilicon 723 -718 723 -718 0 3
rlabel polysilicon 730 -712 730 -712 0 1
rlabel polysilicon 730 -718 730 -718 0 3
rlabel polysilicon 737 -712 737 -712 0 1
rlabel polysilicon 740 -712 740 -712 0 2
rlabel polysilicon 737 -718 737 -718 0 3
rlabel polysilicon 740 -718 740 -718 0 4
rlabel polysilicon 744 -712 744 -712 0 1
rlabel polysilicon 744 -718 744 -718 0 3
rlabel polysilicon 751 -712 751 -712 0 1
rlabel polysilicon 751 -718 751 -718 0 3
rlabel polysilicon 758 -712 758 -712 0 1
rlabel polysilicon 761 -712 761 -712 0 2
rlabel polysilicon 758 -718 758 -718 0 3
rlabel polysilicon 761 -718 761 -718 0 4
rlabel polysilicon 765 -712 765 -712 0 1
rlabel polysilicon 765 -718 765 -718 0 3
rlabel polysilicon 772 -712 772 -712 0 1
rlabel polysilicon 772 -718 772 -718 0 3
rlabel polysilicon 779 -712 779 -712 0 1
rlabel polysilicon 782 -712 782 -712 0 2
rlabel polysilicon 779 -718 779 -718 0 3
rlabel polysilicon 782 -718 782 -718 0 4
rlabel polysilicon 786 -712 786 -712 0 1
rlabel polysilicon 786 -718 786 -718 0 3
rlabel polysilicon 793 -712 793 -712 0 1
rlabel polysilicon 796 -712 796 -712 0 2
rlabel polysilicon 793 -718 793 -718 0 3
rlabel polysilicon 800 -712 800 -712 0 1
rlabel polysilicon 800 -718 800 -718 0 3
rlabel polysilicon 803 -718 803 -718 0 4
rlabel polysilicon 807 -712 807 -712 0 1
rlabel polysilicon 807 -718 807 -718 0 3
rlabel polysilicon 814 -712 814 -712 0 1
rlabel polysilicon 814 -718 814 -718 0 3
rlabel polysilicon 821 -712 821 -712 0 1
rlabel polysilicon 821 -718 821 -718 0 3
rlabel polysilicon 828 -712 828 -712 0 1
rlabel polysilicon 831 -712 831 -712 0 2
rlabel polysilicon 828 -718 828 -718 0 3
rlabel polysilicon 835 -712 835 -712 0 1
rlabel polysilicon 835 -718 835 -718 0 3
rlabel polysilicon 842 -712 842 -712 0 1
rlabel polysilicon 845 -712 845 -712 0 2
rlabel polysilicon 842 -718 842 -718 0 3
rlabel polysilicon 845 -718 845 -718 0 4
rlabel polysilicon 849 -712 849 -712 0 1
rlabel polysilicon 849 -718 849 -718 0 3
rlabel polysilicon 856 -712 856 -712 0 1
rlabel polysilicon 856 -718 856 -718 0 3
rlabel polysilicon 863 -712 863 -712 0 1
rlabel polysilicon 863 -718 863 -718 0 3
rlabel polysilicon 870 -712 870 -712 0 1
rlabel polysilicon 870 -718 870 -718 0 3
rlabel polysilicon 877 -712 877 -712 0 1
rlabel polysilicon 877 -718 877 -718 0 3
rlabel polysilicon 884 -712 884 -712 0 1
rlabel polysilicon 884 -718 884 -718 0 3
rlabel polysilicon 891 -712 891 -712 0 1
rlabel polysilicon 891 -718 891 -718 0 3
rlabel polysilicon 898 -712 898 -712 0 1
rlabel polysilicon 901 -712 901 -712 0 2
rlabel polysilicon 898 -718 898 -718 0 3
rlabel polysilicon 901 -718 901 -718 0 4
rlabel polysilicon 908 -712 908 -712 0 2
rlabel polysilicon 908 -718 908 -718 0 4
rlabel polysilicon 912 -712 912 -712 0 1
rlabel polysilicon 912 -718 912 -718 0 3
rlabel polysilicon 922 -712 922 -712 0 2
rlabel polysilicon 919 -718 919 -718 0 3
rlabel polysilicon 922 -718 922 -718 0 4
rlabel polysilicon 926 -712 926 -712 0 1
rlabel polysilicon 926 -718 926 -718 0 3
rlabel polysilicon 933 -712 933 -712 0 1
rlabel polysilicon 933 -718 933 -718 0 3
rlabel polysilicon 940 -712 940 -712 0 1
rlabel polysilicon 940 -718 940 -718 0 3
rlabel polysilicon 947 -712 947 -712 0 1
rlabel polysilicon 947 -718 947 -718 0 3
rlabel polysilicon 954 -712 954 -712 0 1
rlabel polysilicon 954 -718 954 -718 0 3
rlabel polysilicon 961 -712 961 -712 0 1
rlabel polysilicon 961 -718 961 -718 0 3
rlabel polysilicon 971 -712 971 -712 0 2
rlabel polysilicon 968 -718 968 -718 0 3
rlabel polysilicon 971 -718 971 -718 0 4
rlabel polysilicon 975 -712 975 -712 0 1
rlabel polysilicon 975 -718 975 -718 0 3
rlabel polysilicon 982 -712 982 -712 0 1
rlabel polysilicon 982 -718 982 -718 0 3
rlabel polysilicon 989 -712 989 -712 0 1
rlabel polysilicon 989 -718 989 -718 0 3
rlabel polysilicon 999 -712 999 -712 0 2
rlabel polysilicon 999 -718 999 -718 0 4
rlabel polysilicon 1003 -712 1003 -712 0 1
rlabel polysilicon 1003 -718 1003 -718 0 3
rlabel polysilicon 1010 -712 1010 -712 0 1
rlabel polysilicon 1010 -718 1010 -718 0 3
rlabel polysilicon 1020 -712 1020 -712 0 2
rlabel polysilicon 1017 -718 1017 -718 0 3
rlabel polysilicon 1020 -718 1020 -718 0 4
rlabel polysilicon 1024 -712 1024 -712 0 1
rlabel polysilicon 1024 -718 1024 -718 0 3
rlabel polysilicon 1031 -712 1031 -712 0 1
rlabel polysilicon 1031 -718 1031 -718 0 3
rlabel polysilicon 1038 -712 1038 -712 0 1
rlabel polysilicon 1038 -718 1038 -718 0 3
rlabel polysilicon 1045 -712 1045 -712 0 1
rlabel polysilicon 1045 -718 1045 -718 0 3
rlabel polysilicon 1052 -712 1052 -712 0 1
rlabel polysilicon 1052 -718 1052 -718 0 3
rlabel polysilicon 1059 -712 1059 -712 0 1
rlabel polysilicon 1059 -718 1059 -718 0 3
rlabel polysilicon 1066 -712 1066 -712 0 1
rlabel polysilicon 1066 -718 1066 -718 0 3
rlabel polysilicon 1073 -712 1073 -712 0 1
rlabel polysilicon 1073 -718 1073 -718 0 3
rlabel polysilicon 1080 -712 1080 -712 0 1
rlabel polysilicon 1080 -718 1080 -718 0 3
rlabel polysilicon 1087 -712 1087 -712 0 1
rlabel polysilicon 1087 -718 1087 -718 0 3
rlabel polysilicon 1094 -712 1094 -712 0 1
rlabel polysilicon 1094 -718 1094 -718 0 3
rlabel polysilicon 1101 -712 1101 -712 0 1
rlabel polysilicon 1101 -718 1101 -718 0 3
rlabel polysilicon 1108 -712 1108 -712 0 1
rlabel polysilicon 1108 -718 1108 -718 0 3
rlabel polysilicon 1115 -712 1115 -712 0 1
rlabel polysilicon 1115 -718 1115 -718 0 3
rlabel polysilicon 1122 -712 1122 -712 0 1
rlabel polysilicon 1122 -718 1122 -718 0 3
rlabel polysilicon 1129 -712 1129 -712 0 1
rlabel polysilicon 1129 -718 1129 -718 0 3
rlabel polysilicon 1136 -712 1136 -712 0 1
rlabel polysilicon 1136 -718 1136 -718 0 3
rlabel polysilicon 1143 -712 1143 -712 0 1
rlabel polysilicon 1143 -718 1143 -718 0 3
rlabel polysilicon 1150 -712 1150 -712 0 1
rlabel polysilicon 1150 -718 1150 -718 0 3
rlabel polysilicon 1157 -712 1157 -712 0 1
rlabel polysilicon 1157 -718 1157 -718 0 3
rlabel polysilicon 1164 -712 1164 -712 0 1
rlabel polysilicon 1164 -718 1164 -718 0 3
rlabel polysilicon 1171 -712 1171 -712 0 1
rlabel polysilicon 1171 -718 1171 -718 0 3
rlabel polysilicon 1178 -712 1178 -712 0 1
rlabel polysilicon 1178 -718 1178 -718 0 3
rlabel polysilicon 1185 -712 1185 -712 0 1
rlabel polysilicon 1185 -718 1185 -718 0 3
rlabel polysilicon 1192 -712 1192 -712 0 1
rlabel polysilicon 1192 -718 1192 -718 0 3
rlabel polysilicon 1199 -712 1199 -712 0 1
rlabel polysilicon 1199 -718 1199 -718 0 3
rlabel polysilicon 1206 -712 1206 -712 0 1
rlabel polysilicon 1206 -718 1206 -718 0 3
rlabel polysilicon 1213 -712 1213 -712 0 1
rlabel polysilicon 1213 -718 1213 -718 0 3
rlabel polysilicon 1220 -712 1220 -712 0 1
rlabel polysilicon 1220 -718 1220 -718 0 3
rlabel polysilicon 1227 -712 1227 -712 0 1
rlabel polysilicon 1227 -718 1227 -718 0 3
rlabel polysilicon 1234 -712 1234 -712 0 1
rlabel polysilicon 1234 -718 1234 -718 0 3
rlabel polysilicon 1241 -712 1241 -712 0 1
rlabel polysilicon 1241 -718 1241 -718 0 3
rlabel polysilicon 1248 -712 1248 -712 0 1
rlabel polysilicon 1248 -718 1248 -718 0 3
rlabel polysilicon 1255 -712 1255 -712 0 1
rlabel polysilicon 1255 -718 1255 -718 0 3
rlabel polysilicon 1262 -712 1262 -712 0 1
rlabel polysilicon 1262 -718 1262 -718 0 3
rlabel polysilicon 1269 -712 1269 -712 0 1
rlabel polysilicon 1269 -718 1269 -718 0 3
rlabel polysilicon 1276 -712 1276 -712 0 1
rlabel polysilicon 1276 -718 1276 -718 0 3
rlabel polysilicon 1283 -712 1283 -712 0 1
rlabel polysilicon 1283 -718 1283 -718 0 3
rlabel polysilicon 1290 -712 1290 -712 0 1
rlabel polysilicon 1290 -718 1290 -718 0 3
rlabel polysilicon 1297 -712 1297 -712 0 1
rlabel polysilicon 1297 -718 1297 -718 0 3
rlabel polysilicon 1304 -712 1304 -712 0 1
rlabel polysilicon 1304 -718 1304 -718 0 3
rlabel polysilicon 1311 -712 1311 -712 0 1
rlabel polysilicon 1311 -718 1311 -718 0 3
rlabel polysilicon 1318 -712 1318 -712 0 1
rlabel polysilicon 1318 -718 1318 -718 0 3
rlabel polysilicon 1325 -712 1325 -712 0 1
rlabel polysilicon 1325 -718 1325 -718 0 3
rlabel polysilicon 1332 -712 1332 -712 0 1
rlabel polysilicon 1332 -718 1332 -718 0 3
rlabel polysilicon 1339 -712 1339 -712 0 1
rlabel polysilicon 1339 -718 1339 -718 0 3
rlabel polysilicon 1346 -712 1346 -712 0 1
rlabel polysilicon 1346 -718 1346 -718 0 3
rlabel polysilicon 1353 -712 1353 -712 0 1
rlabel polysilicon 1353 -718 1353 -718 0 3
rlabel polysilicon 1360 -712 1360 -712 0 1
rlabel polysilicon 1360 -718 1360 -718 0 3
rlabel polysilicon 1367 -712 1367 -712 0 1
rlabel polysilicon 1367 -718 1367 -718 0 3
rlabel polysilicon 1374 -712 1374 -712 0 1
rlabel polysilicon 1374 -718 1374 -718 0 3
rlabel polysilicon 1381 -712 1381 -712 0 1
rlabel polysilicon 1381 -718 1381 -718 0 3
rlabel polysilicon 1388 -712 1388 -712 0 1
rlabel polysilicon 1388 -718 1388 -718 0 3
rlabel polysilicon 1395 -712 1395 -712 0 1
rlabel polysilicon 1395 -718 1395 -718 0 3
rlabel polysilicon 1402 -712 1402 -712 0 1
rlabel polysilicon 1402 -718 1402 -718 0 3
rlabel polysilicon 1409 -712 1409 -712 0 1
rlabel polysilicon 1409 -718 1409 -718 0 3
rlabel polysilicon 1416 -712 1416 -712 0 1
rlabel polysilicon 1416 -718 1416 -718 0 3
rlabel polysilicon 1423 -712 1423 -712 0 1
rlabel polysilicon 1423 -718 1423 -718 0 3
rlabel polysilicon 1430 -712 1430 -712 0 1
rlabel polysilicon 1430 -718 1430 -718 0 3
rlabel polysilicon 1437 -712 1437 -712 0 1
rlabel polysilicon 1437 -718 1437 -718 0 3
rlabel polysilicon 1444 -712 1444 -712 0 1
rlabel polysilicon 1444 -718 1444 -718 0 3
rlabel polysilicon 1451 -712 1451 -712 0 1
rlabel polysilicon 1451 -718 1451 -718 0 3
rlabel polysilicon 1458 -712 1458 -712 0 1
rlabel polysilicon 1458 -718 1458 -718 0 3
rlabel polysilicon 1465 -712 1465 -712 0 1
rlabel polysilicon 1465 -718 1465 -718 0 3
rlabel polysilicon 1472 -712 1472 -712 0 1
rlabel polysilicon 1472 -718 1472 -718 0 3
rlabel polysilicon 1479 -712 1479 -712 0 1
rlabel polysilicon 1479 -718 1479 -718 0 3
rlabel polysilicon 1486 -712 1486 -712 0 1
rlabel polysilicon 1486 -718 1486 -718 0 3
rlabel polysilicon 1493 -712 1493 -712 0 1
rlabel polysilicon 1493 -718 1493 -718 0 3
rlabel polysilicon 1500 -712 1500 -712 0 1
rlabel polysilicon 1500 -718 1500 -718 0 3
rlabel polysilicon 1507 -712 1507 -712 0 1
rlabel polysilicon 1507 -718 1507 -718 0 3
rlabel polysilicon 1514 -712 1514 -712 0 1
rlabel polysilicon 1514 -718 1514 -718 0 3
rlabel polysilicon 1521 -712 1521 -712 0 1
rlabel polysilicon 1521 -718 1521 -718 0 3
rlabel polysilicon 1528 -712 1528 -712 0 1
rlabel polysilicon 1528 -718 1528 -718 0 3
rlabel polysilicon 1535 -712 1535 -712 0 1
rlabel polysilicon 1535 -718 1535 -718 0 3
rlabel polysilicon 1542 -712 1542 -712 0 1
rlabel polysilicon 1542 -718 1542 -718 0 3
rlabel polysilicon 1549 -712 1549 -712 0 1
rlabel polysilicon 1549 -718 1549 -718 0 3
rlabel polysilicon 1556 -712 1556 -712 0 1
rlabel polysilicon 1556 -718 1556 -718 0 3
rlabel polysilicon 1563 -712 1563 -712 0 1
rlabel polysilicon 1563 -718 1563 -718 0 3
rlabel polysilicon 1570 -712 1570 -712 0 1
rlabel polysilicon 1570 -718 1570 -718 0 3
rlabel polysilicon 1577 -712 1577 -712 0 1
rlabel polysilicon 1577 -718 1577 -718 0 3
rlabel polysilicon 1584 -712 1584 -712 0 1
rlabel polysilicon 1584 -718 1584 -718 0 3
rlabel polysilicon 1591 -712 1591 -712 0 1
rlabel polysilicon 1591 -718 1591 -718 0 3
rlabel polysilicon 1598 -712 1598 -712 0 1
rlabel polysilicon 1598 -718 1598 -718 0 3
rlabel polysilicon 1605 -712 1605 -712 0 1
rlabel polysilicon 1605 -718 1605 -718 0 3
rlabel polysilicon 1612 -712 1612 -712 0 1
rlabel polysilicon 1612 -718 1612 -718 0 3
rlabel polysilicon 1619 -712 1619 -712 0 1
rlabel polysilicon 1619 -718 1619 -718 0 3
rlabel polysilicon 1626 -712 1626 -712 0 1
rlabel polysilicon 1626 -718 1626 -718 0 3
rlabel polysilicon 1633 -712 1633 -712 0 1
rlabel polysilicon 1633 -718 1633 -718 0 3
rlabel polysilicon 1640 -712 1640 -712 0 1
rlabel polysilicon 1640 -718 1640 -718 0 3
rlabel polysilicon 1647 -712 1647 -712 0 1
rlabel polysilicon 1647 -718 1647 -718 0 3
rlabel polysilicon 1657 -712 1657 -712 0 2
rlabel polysilicon 1654 -718 1654 -718 0 3
rlabel polysilicon 1661 -712 1661 -712 0 1
rlabel polysilicon 1661 -718 1661 -718 0 3
rlabel polysilicon 1668 -712 1668 -712 0 1
rlabel polysilicon 1671 -712 1671 -712 0 2
rlabel polysilicon 1671 -718 1671 -718 0 4
rlabel polysilicon 1787 -712 1787 -712 0 1
rlabel polysilicon 1787 -718 1787 -718 0 3
rlabel polysilicon 1794 -712 1794 -712 0 1
rlabel polysilicon 1794 -718 1794 -718 0 3
rlabel polysilicon 1801 -712 1801 -712 0 1
rlabel polysilicon 1801 -718 1801 -718 0 3
rlabel polysilicon 1822 -712 1822 -712 0 1
rlabel polysilicon 1822 -718 1822 -718 0 3
rlabel polysilicon 1857 -712 1857 -712 0 1
rlabel polysilicon 1857 -718 1857 -718 0 3
rlabel polysilicon 9 -857 9 -857 0 1
rlabel polysilicon 9 -863 9 -863 0 3
rlabel polysilicon 16 -863 16 -863 0 3
rlabel polysilicon 23 -857 23 -857 0 1
rlabel polysilicon 23 -863 23 -863 0 3
rlabel polysilicon 30 -857 30 -857 0 1
rlabel polysilicon 30 -863 30 -863 0 3
rlabel polysilicon 37 -857 37 -857 0 1
rlabel polysilicon 37 -863 37 -863 0 3
rlabel polysilicon 44 -857 44 -857 0 1
rlabel polysilicon 47 -863 47 -863 0 4
rlabel polysilicon 54 -857 54 -857 0 2
rlabel polysilicon 51 -863 51 -863 0 3
rlabel polysilicon 54 -863 54 -863 0 4
rlabel polysilicon 58 -857 58 -857 0 1
rlabel polysilicon 58 -863 58 -863 0 3
rlabel polysilicon 65 -857 65 -857 0 1
rlabel polysilicon 65 -863 65 -863 0 3
rlabel polysilicon 72 -857 72 -857 0 1
rlabel polysilicon 72 -863 72 -863 0 3
rlabel polysilicon 79 -857 79 -857 0 1
rlabel polysilicon 82 -857 82 -857 0 2
rlabel polysilicon 79 -863 79 -863 0 3
rlabel polysilicon 86 -857 86 -857 0 1
rlabel polysilicon 86 -863 86 -863 0 3
rlabel polysilicon 93 -857 93 -857 0 1
rlabel polysilicon 93 -863 93 -863 0 3
rlabel polysilicon 100 -857 100 -857 0 1
rlabel polysilicon 100 -863 100 -863 0 3
rlabel polysilicon 107 -857 107 -857 0 1
rlabel polysilicon 107 -863 107 -863 0 3
rlabel polysilicon 114 -857 114 -857 0 1
rlabel polysilicon 114 -863 114 -863 0 3
rlabel polysilicon 121 -857 121 -857 0 1
rlabel polysilicon 124 -857 124 -857 0 2
rlabel polysilicon 121 -863 121 -863 0 3
rlabel polysilicon 128 -857 128 -857 0 1
rlabel polysilicon 128 -863 128 -863 0 3
rlabel polysilicon 135 -857 135 -857 0 1
rlabel polysilicon 135 -863 135 -863 0 3
rlabel polysilicon 142 -857 142 -857 0 1
rlabel polysilicon 142 -863 142 -863 0 3
rlabel polysilicon 149 -857 149 -857 0 1
rlabel polysilicon 149 -863 149 -863 0 3
rlabel polysilicon 156 -857 156 -857 0 1
rlabel polysilicon 156 -863 156 -863 0 3
rlabel polysilicon 163 -857 163 -857 0 1
rlabel polysilicon 166 -857 166 -857 0 2
rlabel polysilicon 163 -863 163 -863 0 3
rlabel polysilicon 166 -863 166 -863 0 4
rlabel polysilicon 170 -857 170 -857 0 1
rlabel polysilicon 170 -863 170 -863 0 3
rlabel polysilicon 177 -857 177 -857 0 1
rlabel polysilicon 180 -857 180 -857 0 2
rlabel polysilicon 177 -863 177 -863 0 3
rlabel polysilicon 180 -863 180 -863 0 4
rlabel polysilicon 184 -857 184 -857 0 1
rlabel polysilicon 184 -863 184 -863 0 3
rlabel polysilicon 191 -857 191 -857 0 1
rlabel polysilicon 194 -863 194 -863 0 4
rlabel polysilicon 198 -857 198 -857 0 1
rlabel polysilicon 201 -857 201 -857 0 2
rlabel polysilicon 198 -863 198 -863 0 3
rlabel polysilicon 201 -863 201 -863 0 4
rlabel polysilicon 205 -857 205 -857 0 1
rlabel polysilicon 205 -863 205 -863 0 3
rlabel polysilicon 212 -857 212 -857 0 1
rlabel polysilicon 212 -863 212 -863 0 3
rlabel polysilicon 219 -857 219 -857 0 1
rlabel polysilicon 226 -857 226 -857 0 1
rlabel polysilicon 226 -863 226 -863 0 3
rlabel polysilicon 233 -857 233 -857 0 1
rlabel polysilicon 233 -863 233 -863 0 3
rlabel polysilicon 240 -857 240 -857 0 1
rlabel polysilicon 240 -863 240 -863 0 3
rlabel polysilicon 247 -857 247 -857 0 1
rlabel polysilicon 247 -863 247 -863 0 3
rlabel polysilicon 254 -857 254 -857 0 1
rlabel polysilicon 254 -863 254 -863 0 3
rlabel polysilicon 261 -857 261 -857 0 1
rlabel polysilicon 261 -863 261 -863 0 3
rlabel polysilicon 268 -857 268 -857 0 1
rlabel polysilicon 268 -863 268 -863 0 3
rlabel polysilicon 275 -857 275 -857 0 1
rlabel polysilicon 275 -863 275 -863 0 3
rlabel polysilicon 282 -857 282 -857 0 1
rlabel polysilicon 282 -863 282 -863 0 3
rlabel polysilicon 289 -857 289 -857 0 1
rlabel polysilicon 289 -863 289 -863 0 3
rlabel polysilicon 296 -857 296 -857 0 1
rlabel polysilicon 296 -863 296 -863 0 3
rlabel polysilicon 303 -857 303 -857 0 1
rlabel polysilicon 310 -857 310 -857 0 1
rlabel polysilicon 310 -863 310 -863 0 3
rlabel polysilicon 317 -863 317 -863 0 3
rlabel polysilicon 324 -857 324 -857 0 1
rlabel polysilicon 324 -863 324 -863 0 3
rlabel polysilicon 331 -857 331 -857 0 1
rlabel polysilicon 331 -863 331 -863 0 3
rlabel polysilicon 338 -857 338 -857 0 1
rlabel polysilicon 338 -863 338 -863 0 3
rlabel polysilicon 345 -857 345 -857 0 1
rlabel polysilicon 345 -863 345 -863 0 3
rlabel polysilicon 352 -857 352 -857 0 1
rlabel polysilicon 352 -863 352 -863 0 3
rlabel polysilicon 359 -857 359 -857 0 1
rlabel polysilicon 359 -863 359 -863 0 3
rlabel polysilicon 366 -857 366 -857 0 1
rlabel polysilicon 366 -863 366 -863 0 3
rlabel polysilicon 373 -857 373 -857 0 1
rlabel polysilicon 373 -863 373 -863 0 3
rlabel polysilicon 380 -857 380 -857 0 1
rlabel polysilicon 380 -863 380 -863 0 3
rlabel polysilicon 387 -857 387 -857 0 1
rlabel polysilicon 387 -863 387 -863 0 3
rlabel polysilicon 394 -857 394 -857 0 1
rlabel polysilicon 394 -863 394 -863 0 3
rlabel polysilicon 401 -857 401 -857 0 1
rlabel polysilicon 401 -863 401 -863 0 3
rlabel polysilicon 408 -857 408 -857 0 1
rlabel polysilicon 408 -863 408 -863 0 3
rlabel polysilicon 415 -857 415 -857 0 1
rlabel polysilicon 415 -863 415 -863 0 3
rlabel polysilicon 422 -857 422 -857 0 1
rlabel polysilicon 422 -863 422 -863 0 3
rlabel polysilicon 429 -857 429 -857 0 1
rlabel polysilicon 429 -863 429 -863 0 3
rlabel polysilicon 439 -857 439 -857 0 2
rlabel polysilicon 436 -863 436 -863 0 3
rlabel polysilicon 439 -863 439 -863 0 4
rlabel polysilicon 443 -857 443 -857 0 1
rlabel polysilicon 443 -863 443 -863 0 3
rlabel polysilicon 450 -857 450 -857 0 1
rlabel polysilicon 450 -863 450 -863 0 3
rlabel polysilicon 457 -857 457 -857 0 1
rlabel polysilicon 457 -863 457 -863 0 3
rlabel polysilicon 464 -857 464 -857 0 1
rlabel polysilicon 464 -863 464 -863 0 3
rlabel polysilicon 471 -857 471 -857 0 1
rlabel polysilicon 471 -863 471 -863 0 3
rlabel polysilicon 478 -857 478 -857 0 1
rlabel polysilicon 478 -863 478 -863 0 3
rlabel polysilicon 485 -857 485 -857 0 1
rlabel polysilicon 485 -863 485 -863 0 3
rlabel polysilicon 492 -857 492 -857 0 1
rlabel polysilicon 495 -857 495 -857 0 2
rlabel polysilicon 492 -863 492 -863 0 3
rlabel polysilicon 495 -863 495 -863 0 4
rlabel polysilicon 499 -857 499 -857 0 1
rlabel polysilicon 499 -863 499 -863 0 3
rlabel polysilicon 506 -857 506 -857 0 1
rlabel polysilicon 506 -863 506 -863 0 3
rlabel polysilicon 513 -857 513 -857 0 1
rlabel polysilicon 516 -857 516 -857 0 2
rlabel polysilicon 513 -863 513 -863 0 3
rlabel polysilicon 516 -863 516 -863 0 4
rlabel polysilicon 520 -857 520 -857 0 1
rlabel polysilicon 520 -863 520 -863 0 3
rlabel polysilicon 527 -857 527 -857 0 1
rlabel polysilicon 527 -863 527 -863 0 3
rlabel polysilicon 534 -857 534 -857 0 1
rlabel polysilicon 534 -863 534 -863 0 3
rlabel polysilicon 541 -857 541 -857 0 1
rlabel polysilicon 541 -863 541 -863 0 3
rlabel polysilicon 548 -857 548 -857 0 1
rlabel polysilicon 548 -863 548 -863 0 3
rlabel polysilicon 555 -857 555 -857 0 1
rlabel polysilicon 558 -857 558 -857 0 2
rlabel polysilicon 558 -863 558 -863 0 4
rlabel polysilicon 562 -857 562 -857 0 1
rlabel polysilicon 562 -863 562 -863 0 3
rlabel polysilicon 572 -857 572 -857 0 2
rlabel polysilicon 569 -863 569 -863 0 3
rlabel polysilicon 572 -863 572 -863 0 4
rlabel polysilicon 576 -857 576 -857 0 1
rlabel polysilicon 579 -857 579 -857 0 2
rlabel polysilicon 576 -863 576 -863 0 3
rlabel polysilicon 583 -857 583 -857 0 1
rlabel polysilicon 586 -857 586 -857 0 2
rlabel polysilicon 583 -863 583 -863 0 3
rlabel polysilicon 586 -863 586 -863 0 4
rlabel polysilicon 590 -857 590 -857 0 1
rlabel polysilicon 590 -863 590 -863 0 3
rlabel polysilicon 597 -857 597 -857 0 1
rlabel polysilicon 597 -863 597 -863 0 3
rlabel polysilicon 600 -863 600 -863 0 4
rlabel polysilicon 604 -857 604 -857 0 1
rlabel polysilicon 604 -863 604 -863 0 3
rlabel polysilicon 611 -857 611 -857 0 1
rlabel polysilicon 614 -857 614 -857 0 2
rlabel polysilicon 611 -863 611 -863 0 3
rlabel polysilicon 618 -857 618 -857 0 1
rlabel polysilicon 621 -857 621 -857 0 2
rlabel polysilicon 618 -863 618 -863 0 3
rlabel polysilicon 621 -863 621 -863 0 4
rlabel polysilicon 625 -857 625 -857 0 1
rlabel polysilicon 628 -857 628 -857 0 2
rlabel polysilicon 625 -863 625 -863 0 3
rlabel polysilicon 628 -863 628 -863 0 4
rlabel polysilicon 632 -857 632 -857 0 1
rlabel polysilicon 632 -863 632 -863 0 3
rlabel polysilicon 639 -857 639 -857 0 1
rlabel polysilicon 639 -863 639 -863 0 3
rlabel polysilicon 646 -857 646 -857 0 1
rlabel polysilicon 646 -863 646 -863 0 3
rlabel polysilicon 653 -857 653 -857 0 1
rlabel polysilicon 653 -863 653 -863 0 3
rlabel polysilicon 660 -857 660 -857 0 1
rlabel polysilicon 660 -863 660 -863 0 3
rlabel polysilicon 667 -857 667 -857 0 1
rlabel polysilicon 667 -863 667 -863 0 3
rlabel polysilicon 674 -857 674 -857 0 1
rlabel polysilicon 674 -863 674 -863 0 3
rlabel polysilicon 681 -857 681 -857 0 1
rlabel polysilicon 681 -863 681 -863 0 3
rlabel polysilicon 691 -857 691 -857 0 2
rlabel polysilicon 688 -863 688 -863 0 3
rlabel polysilicon 691 -863 691 -863 0 4
rlabel polysilicon 695 -857 695 -857 0 1
rlabel polysilicon 695 -863 695 -863 0 3
rlabel polysilicon 702 -863 702 -863 0 3
rlabel polysilicon 705 -863 705 -863 0 4
rlabel polysilicon 709 -857 709 -857 0 1
rlabel polysilicon 709 -863 709 -863 0 3
rlabel polysilicon 716 -857 716 -857 0 1
rlabel polysilicon 716 -863 716 -863 0 3
rlabel polysilicon 723 -857 723 -857 0 1
rlabel polysilicon 723 -863 723 -863 0 3
rlabel polysilicon 730 -857 730 -857 0 1
rlabel polysilicon 730 -863 730 -863 0 3
rlabel polysilicon 737 -857 737 -857 0 1
rlabel polysilicon 737 -863 737 -863 0 3
rlabel polysilicon 744 -857 744 -857 0 1
rlabel polysilicon 744 -863 744 -863 0 3
rlabel polysilicon 751 -857 751 -857 0 1
rlabel polysilicon 751 -863 751 -863 0 3
rlabel polysilicon 761 -857 761 -857 0 2
rlabel polysilicon 758 -863 758 -863 0 3
rlabel polysilicon 761 -863 761 -863 0 4
rlabel polysilicon 765 -857 765 -857 0 1
rlabel polysilicon 765 -863 765 -863 0 3
rlabel polysilicon 772 -857 772 -857 0 1
rlabel polysilicon 772 -863 772 -863 0 3
rlabel polysilicon 779 -857 779 -857 0 1
rlabel polysilicon 782 -857 782 -857 0 2
rlabel polysilicon 779 -863 779 -863 0 3
rlabel polysilicon 782 -863 782 -863 0 4
rlabel polysilicon 786 -857 786 -857 0 1
rlabel polysilicon 789 -857 789 -857 0 2
rlabel polysilicon 786 -863 786 -863 0 3
rlabel polysilicon 789 -863 789 -863 0 4
rlabel polysilicon 793 -857 793 -857 0 1
rlabel polysilicon 793 -863 793 -863 0 3
rlabel polysilicon 800 -857 800 -857 0 1
rlabel polysilicon 803 -857 803 -857 0 2
rlabel polysilicon 800 -863 800 -863 0 3
rlabel polysilicon 807 -857 807 -857 0 1
rlabel polysilicon 807 -863 807 -863 0 3
rlabel polysilicon 814 -857 814 -857 0 1
rlabel polysilicon 814 -863 814 -863 0 3
rlabel polysilicon 821 -857 821 -857 0 1
rlabel polysilicon 824 -857 824 -857 0 2
rlabel polysilicon 821 -863 821 -863 0 3
rlabel polysilicon 824 -863 824 -863 0 4
rlabel polysilicon 828 -857 828 -857 0 1
rlabel polysilicon 831 -857 831 -857 0 2
rlabel polysilicon 828 -863 828 -863 0 3
rlabel polysilicon 831 -863 831 -863 0 4
rlabel polysilicon 835 -857 835 -857 0 1
rlabel polysilicon 835 -863 835 -863 0 3
rlabel polysilicon 842 -857 842 -857 0 1
rlabel polysilicon 842 -863 842 -863 0 3
rlabel polysilicon 849 -857 849 -857 0 1
rlabel polysilicon 849 -863 849 -863 0 3
rlabel polysilicon 856 -857 856 -857 0 1
rlabel polysilicon 856 -863 856 -863 0 3
rlabel polysilicon 863 -857 863 -857 0 1
rlabel polysilicon 863 -863 863 -863 0 3
rlabel polysilicon 870 -857 870 -857 0 1
rlabel polysilicon 870 -863 870 -863 0 3
rlabel polysilicon 877 -857 877 -857 0 1
rlabel polysilicon 877 -863 877 -863 0 3
rlabel polysilicon 884 -857 884 -857 0 1
rlabel polysilicon 884 -863 884 -863 0 3
rlabel polysilicon 891 -857 891 -857 0 1
rlabel polysilicon 891 -863 891 -863 0 3
rlabel polysilicon 898 -857 898 -857 0 1
rlabel polysilicon 898 -863 898 -863 0 3
rlabel polysilicon 905 -857 905 -857 0 1
rlabel polysilicon 905 -863 905 -863 0 3
rlabel polysilicon 912 -857 912 -857 0 1
rlabel polysilicon 912 -863 912 -863 0 3
rlabel polysilicon 919 -857 919 -857 0 1
rlabel polysilicon 919 -863 919 -863 0 3
rlabel polysilicon 922 -863 922 -863 0 4
rlabel polysilicon 926 -857 926 -857 0 1
rlabel polysilicon 926 -863 926 -863 0 3
rlabel polysilicon 933 -857 933 -857 0 1
rlabel polysilicon 933 -863 933 -863 0 3
rlabel polysilicon 940 -857 940 -857 0 1
rlabel polysilicon 940 -863 940 -863 0 3
rlabel polysilicon 947 -857 947 -857 0 1
rlabel polysilicon 947 -863 947 -863 0 3
rlabel polysilicon 954 -857 954 -857 0 1
rlabel polysilicon 954 -863 954 -863 0 3
rlabel polysilicon 961 -857 961 -857 0 1
rlabel polysilicon 961 -863 961 -863 0 3
rlabel polysilicon 968 -857 968 -857 0 1
rlabel polysilicon 968 -863 968 -863 0 3
rlabel polysilicon 975 -863 975 -863 0 3
rlabel polysilicon 982 -857 982 -857 0 1
rlabel polysilicon 982 -863 982 -863 0 3
rlabel polysilicon 989 -857 989 -857 0 1
rlabel polysilicon 989 -863 989 -863 0 3
rlabel polysilicon 996 -857 996 -857 0 1
rlabel polysilicon 996 -863 996 -863 0 3
rlabel polysilicon 1003 -857 1003 -857 0 1
rlabel polysilicon 1003 -863 1003 -863 0 3
rlabel polysilicon 1010 -857 1010 -857 0 1
rlabel polysilicon 1010 -863 1010 -863 0 3
rlabel polysilicon 1017 -857 1017 -857 0 1
rlabel polysilicon 1017 -863 1017 -863 0 3
rlabel polysilicon 1024 -857 1024 -857 0 1
rlabel polysilicon 1024 -863 1024 -863 0 3
rlabel polysilicon 1031 -857 1031 -857 0 1
rlabel polysilicon 1034 -857 1034 -857 0 2
rlabel polysilicon 1031 -863 1031 -863 0 3
rlabel polysilicon 1034 -863 1034 -863 0 4
rlabel polysilicon 1038 -857 1038 -857 0 1
rlabel polysilicon 1038 -863 1038 -863 0 3
rlabel polysilicon 1045 -857 1045 -857 0 1
rlabel polysilicon 1045 -863 1045 -863 0 3
rlabel polysilicon 1052 -857 1052 -857 0 1
rlabel polysilicon 1052 -863 1052 -863 0 3
rlabel polysilicon 1059 -857 1059 -857 0 1
rlabel polysilicon 1059 -863 1059 -863 0 3
rlabel polysilicon 1066 -857 1066 -857 0 1
rlabel polysilicon 1066 -863 1066 -863 0 3
rlabel polysilicon 1073 -857 1073 -857 0 1
rlabel polysilicon 1073 -863 1073 -863 0 3
rlabel polysilicon 1080 -857 1080 -857 0 1
rlabel polysilicon 1080 -863 1080 -863 0 3
rlabel polysilicon 1087 -857 1087 -857 0 1
rlabel polysilicon 1087 -863 1087 -863 0 3
rlabel polysilicon 1094 -857 1094 -857 0 1
rlabel polysilicon 1094 -863 1094 -863 0 3
rlabel polysilicon 1101 -857 1101 -857 0 1
rlabel polysilicon 1101 -863 1101 -863 0 3
rlabel polysilicon 1108 -857 1108 -857 0 1
rlabel polysilicon 1108 -863 1108 -863 0 3
rlabel polysilicon 1111 -863 1111 -863 0 4
rlabel polysilicon 1115 -857 1115 -857 0 1
rlabel polysilicon 1115 -863 1115 -863 0 3
rlabel polysilicon 1122 -857 1122 -857 0 1
rlabel polysilicon 1122 -863 1122 -863 0 3
rlabel polysilicon 1129 -857 1129 -857 0 1
rlabel polysilicon 1129 -863 1129 -863 0 3
rlabel polysilicon 1136 -857 1136 -857 0 1
rlabel polysilicon 1136 -863 1136 -863 0 3
rlabel polysilicon 1143 -857 1143 -857 0 1
rlabel polysilicon 1143 -863 1143 -863 0 3
rlabel polysilicon 1150 -857 1150 -857 0 1
rlabel polysilicon 1150 -863 1150 -863 0 3
rlabel polysilicon 1157 -857 1157 -857 0 1
rlabel polysilicon 1157 -863 1157 -863 0 3
rlabel polysilicon 1164 -857 1164 -857 0 1
rlabel polysilicon 1164 -863 1164 -863 0 3
rlabel polysilicon 1171 -857 1171 -857 0 1
rlabel polysilicon 1171 -863 1171 -863 0 3
rlabel polysilicon 1178 -857 1178 -857 0 1
rlabel polysilicon 1178 -863 1178 -863 0 3
rlabel polysilicon 1185 -857 1185 -857 0 1
rlabel polysilicon 1185 -863 1185 -863 0 3
rlabel polysilicon 1192 -857 1192 -857 0 1
rlabel polysilicon 1195 -857 1195 -857 0 2
rlabel polysilicon 1192 -863 1192 -863 0 3
rlabel polysilicon 1199 -857 1199 -857 0 1
rlabel polysilicon 1199 -863 1199 -863 0 3
rlabel polysilicon 1206 -857 1206 -857 0 1
rlabel polysilicon 1206 -863 1206 -863 0 3
rlabel polysilicon 1213 -857 1213 -857 0 1
rlabel polysilicon 1213 -863 1213 -863 0 3
rlabel polysilicon 1220 -857 1220 -857 0 1
rlabel polysilicon 1220 -863 1220 -863 0 3
rlabel polysilicon 1227 -857 1227 -857 0 1
rlabel polysilicon 1227 -863 1227 -863 0 3
rlabel polysilicon 1234 -857 1234 -857 0 1
rlabel polysilicon 1234 -863 1234 -863 0 3
rlabel polysilicon 1241 -857 1241 -857 0 1
rlabel polysilicon 1241 -863 1241 -863 0 3
rlabel polysilicon 1248 -857 1248 -857 0 1
rlabel polysilicon 1248 -863 1248 -863 0 3
rlabel polysilicon 1255 -857 1255 -857 0 1
rlabel polysilicon 1255 -863 1255 -863 0 3
rlabel polysilicon 1262 -857 1262 -857 0 1
rlabel polysilicon 1262 -863 1262 -863 0 3
rlabel polysilicon 1269 -857 1269 -857 0 1
rlabel polysilicon 1269 -863 1269 -863 0 3
rlabel polysilicon 1276 -857 1276 -857 0 1
rlabel polysilicon 1276 -863 1276 -863 0 3
rlabel polysilicon 1283 -857 1283 -857 0 1
rlabel polysilicon 1283 -863 1283 -863 0 3
rlabel polysilicon 1290 -857 1290 -857 0 1
rlabel polysilicon 1290 -863 1290 -863 0 3
rlabel polysilicon 1297 -857 1297 -857 0 1
rlabel polysilicon 1297 -863 1297 -863 0 3
rlabel polysilicon 1304 -857 1304 -857 0 1
rlabel polysilicon 1304 -863 1304 -863 0 3
rlabel polysilicon 1311 -857 1311 -857 0 1
rlabel polysilicon 1311 -863 1311 -863 0 3
rlabel polysilicon 1318 -857 1318 -857 0 1
rlabel polysilicon 1318 -863 1318 -863 0 3
rlabel polysilicon 1325 -857 1325 -857 0 1
rlabel polysilicon 1325 -863 1325 -863 0 3
rlabel polysilicon 1332 -857 1332 -857 0 1
rlabel polysilicon 1332 -863 1332 -863 0 3
rlabel polysilicon 1339 -857 1339 -857 0 1
rlabel polysilicon 1339 -863 1339 -863 0 3
rlabel polysilicon 1346 -857 1346 -857 0 1
rlabel polysilicon 1346 -863 1346 -863 0 3
rlabel polysilicon 1353 -857 1353 -857 0 1
rlabel polysilicon 1353 -863 1353 -863 0 3
rlabel polysilicon 1360 -857 1360 -857 0 1
rlabel polysilicon 1360 -863 1360 -863 0 3
rlabel polysilicon 1367 -857 1367 -857 0 1
rlabel polysilicon 1367 -863 1367 -863 0 3
rlabel polysilicon 1374 -857 1374 -857 0 1
rlabel polysilicon 1374 -863 1374 -863 0 3
rlabel polysilicon 1381 -857 1381 -857 0 1
rlabel polysilicon 1381 -863 1381 -863 0 3
rlabel polysilicon 1388 -857 1388 -857 0 1
rlabel polysilicon 1388 -863 1388 -863 0 3
rlabel polysilicon 1395 -857 1395 -857 0 1
rlabel polysilicon 1395 -863 1395 -863 0 3
rlabel polysilicon 1402 -857 1402 -857 0 1
rlabel polysilicon 1402 -863 1402 -863 0 3
rlabel polysilicon 1409 -857 1409 -857 0 1
rlabel polysilicon 1409 -863 1409 -863 0 3
rlabel polysilicon 1416 -857 1416 -857 0 1
rlabel polysilicon 1416 -863 1416 -863 0 3
rlabel polysilicon 1423 -857 1423 -857 0 1
rlabel polysilicon 1423 -863 1423 -863 0 3
rlabel polysilicon 1430 -857 1430 -857 0 1
rlabel polysilicon 1430 -863 1430 -863 0 3
rlabel polysilicon 1437 -857 1437 -857 0 1
rlabel polysilicon 1437 -863 1437 -863 0 3
rlabel polysilicon 1444 -857 1444 -857 0 1
rlabel polysilicon 1444 -863 1444 -863 0 3
rlabel polysilicon 1451 -857 1451 -857 0 1
rlabel polysilicon 1451 -863 1451 -863 0 3
rlabel polysilicon 1458 -857 1458 -857 0 1
rlabel polysilicon 1458 -863 1458 -863 0 3
rlabel polysilicon 1465 -857 1465 -857 0 1
rlabel polysilicon 1465 -863 1465 -863 0 3
rlabel polysilicon 1472 -857 1472 -857 0 1
rlabel polysilicon 1472 -863 1472 -863 0 3
rlabel polysilicon 1479 -857 1479 -857 0 1
rlabel polysilicon 1479 -863 1479 -863 0 3
rlabel polysilicon 1486 -857 1486 -857 0 1
rlabel polysilicon 1486 -863 1486 -863 0 3
rlabel polysilicon 1493 -857 1493 -857 0 1
rlabel polysilicon 1493 -863 1493 -863 0 3
rlabel polysilicon 1500 -857 1500 -857 0 1
rlabel polysilicon 1500 -863 1500 -863 0 3
rlabel polysilicon 1507 -857 1507 -857 0 1
rlabel polysilicon 1507 -863 1507 -863 0 3
rlabel polysilicon 1514 -857 1514 -857 0 1
rlabel polysilicon 1514 -863 1514 -863 0 3
rlabel polysilicon 1521 -857 1521 -857 0 1
rlabel polysilicon 1521 -863 1521 -863 0 3
rlabel polysilicon 1528 -857 1528 -857 0 1
rlabel polysilicon 1528 -863 1528 -863 0 3
rlabel polysilicon 1535 -857 1535 -857 0 1
rlabel polysilicon 1535 -863 1535 -863 0 3
rlabel polysilicon 1542 -857 1542 -857 0 1
rlabel polysilicon 1542 -863 1542 -863 0 3
rlabel polysilicon 1549 -857 1549 -857 0 1
rlabel polysilicon 1549 -863 1549 -863 0 3
rlabel polysilicon 1556 -857 1556 -857 0 1
rlabel polysilicon 1556 -863 1556 -863 0 3
rlabel polysilicon 1563 -857 1563 -857 0 1
rlabel polysilicon 1563 -863 1563 -863 0 3
rlabel polysilicon 1570 -857 1570 -857 0 1
rlabel polysilicon 1570 -863 1570 -863 0 3
rlabel polysilicon 1577 -857 1577 -857 0 1
rlabel polysilicon 1577 -863 1577 -863 0 3
rlabel polysilicon 1584 -857 1584 -857 0 1
rlabel polysilicon 1584 -863 1584 -863 0 3
rlabel polysilicon 1591 -857 1591 -857 0 1
rlabel polysilicon 1591 -863 1591 -863 0 3
rlabel polysilicon 1594 -863 1594 -863 0 4
rlabel polysilicon 1598 -857 1598 -857 0 1
rlabel polysilicon 1598 -863 1598 -863 0 3
rlabel polysilicon 1605 -857 1605 -857 0 1
rlabel polysilicon 1605 -863 1605 -863 0 3
rlabel polysilicon 1612 -857 1612 -857 0 1
rlabel polysilicon 1612 -863 1612 -863 0 3
rlabel polysilicon 1619 -857 1619 -857 0 1
rlabel polysilicon 1619 -863 1619 -863 0 3
rlabel polysilicon 1626 -857 1626 -857 0 1
rlabel polysilicon 1626 -863 1626 -863 0 3
rlabel polysilicon 1633 -857 1633 -857 0 1
rlabel polysilicon 1633 -863 1633 -863 0 3
rlabel polysilicon 1640 -857 1640 -857 0 1
rlabel polysilicon 1640 -863 1640 -863 0 3
rlabel polysilicon 1647 -857 1647 -857 0 1
rlabel polysilicon 1647 -863 1647 -863 0 3
rlabel polysilicon 1654 -857 1654 -857 0 1
rlabel polysilicon 1654 -863 1654 -863 0 3
rlabel polysilicon 1661 -857 1661 -857 0 1
rlabel polysilicon 1661 -863 1661 -863 0 3
rlabel polysilicon 1668 -857 1668 -857 0 1
rlabel polysilicon 1668 -863 1668 -863 0 3
rlabel polysilicon 1675 -857 1675 -857 0 1
rlabel polysilicon 1675 -863 1675 -863 0 3
rlabel polysilicon 1682 -857 1682 -857 0 1
rlabel polysilicon 1682 -863 1682 -863 0 3
rlabel polysilicon 1689 -857 1689 -857 0 1
rlabel polysilicon 1689 -863 1689 -863 0 3
rlabel polysilicon 1696 -857 1696 -857 0 1
rlabel polysilicon 1696 -863 1696 -863 0 3
rlabel polysilicon 1703 -857 1703 -857 0 1
rlabel polysilicon 1703 -863 1703 -863 0 3
rlabel polysilicon 1710 -857 1710 -857 0 1
rlabel polysilicon 1710 -863 1710 -863 0 3
rlabel polysilicon 1717 -857 1717 -857 0 1
rlabel polysilicon 1717 -863 1717 -863 0 3
rlabel polysilicon 1724 -857 1724 -857 0 1
rlabel polysilicon 1724 -863 1724 -863 0 3
rlabel polysilicon 1731 -857 1731 -857 0 1
rlabel polysilicon 1731 -863 1731 -863 0 3
rlabel polysilicon 1738 -857 1738 -857 0 1
rlabel polysilicon 1738 -863 1738 -863 0 3
rlabel polysilicon 1745 -857 1745 -857 0 1
rlabel polysilicon 1745 -863 1745 -863 0 3
rlabel polysilicon 1752 -857 1752 -857 0 1
rlabel polysilicon 1752 -863 1752 -863 0 3
rlabel polysilicon 1759 -857 1759 -857 0 1
rlabel polysilicon 1759 -863 1759 -863 0 3
rlabel polysilicon 1766 -857 1766 -857 0 1
rlabel polysilicon 1766 -863 1766 -863 0 3
rlabel polysilicon 1773 -857 1773 -857 0 1
rlabel polysilicon 1773 -863 1773 -863 0 3
rlabel polysilicon 1780 -857 1780 -857 0 1
rlabel polysilicon 1783 -857 1783 -857 0 2
rlabel polysilicon 1780 -863 1780 -863 0 3
rlabel polysilicon 1783 -863 1783 -863 0 4
rlabel polysilicon 1787 -857 1787 -857 0 1
rlabel polysilicon 1787 -863 1787 -863 0 3
rlabel polysilicon 1794 -857 1794 -857 0 1
rlabel polysilicon 1794 -863 1794 -863 0 3
rlabel polysilicon 1801 -857 1801 -857 0 1
rlabel polysilicon 1801 -863 1801 -863 0 3
rlabel polysilicon 1808 -857 1808 -857 0 1
rlabel polysilicon 1808 -863 1808 -863 0 3
rlabel polysilicon 1818 -863 1818 -863 0 4
rlabel polysilicon 1822 -857 1822 -857 0 1
rlabel polysilicon 1822 -863 1822 -863 0 3
rlabel polysilicon 1829 -857 1829 -857 0 1
rlabel polysilicon 1829 -863 1829 -863 0 3
rlabel polysilicon 1836 -857 1836 -857 0 1
rlabel polysilicon 1836 -863 1836 -863 0 3
rlabel polysilicon 1843 -857 1843 -857 0 1
rlabel polysilicon 1843 -863 1843 -863 0 3
rlabel polysilicon 1850 -857 1850 -857 0 1
rlabel polysilicon 1850 -863 1850 -863 0 3
rlabel polysilicon 1857 -857 1857 -857 0 1
rlabel polysilicon 1857 -863 1857 -863 0 3
rlabel polysilicon 1885 -857 1885 -857 0 1
rlabel polysilicon 1885 -863 1885 -863 0 3
rlabel polysilicon 1892 -857 1892 -857 0 1
rlabel polysilicon 1892 -863 1892 -863 0 3
rlabel polysilicon 2 -978 2 -978 0 1
rlabel polysilicon 2 -984 2 -984 0 3
rlabel polysilicon 9 -978 9 -978 0 1
rlabel polysilicon 9 -984 9 -984 0 3
rlabel polysilicon 16 -978 16 -978 0 1
rlabel polysilicon 16 -984 16 -984 0 3
rlabel polysilicon 23 -978 23 -978 0 1
rlabel polysilicon 23 -984 23 -984 0 3
rlabel polysilicon 30 -978 30 -978 0 1
rlabel polysilicon 30 -984 30 -984 0 3
rlabel polysilicon 37 -978 37 -978 0 1
rlabel polysilicon 37 -984 37 -984 0 3
rlabel polysilicon 44 -978 44 -978 0 1
rlabel polysilicon 44 -984 44 -984 0 3
rlabel polysilicon 51 -978 51 -978 0 1
rlabel polysilicon 51 -984 51 -984 0 3
rlabel polysilicon 58 -978 58 -978 0 1
rlabel polysilicon 58 -984 58 -984 0 3
rlabel polysilicon 65 -978 65 -978 0 1
rlabel polysilicon 68 -978 68 -978 0 2
rlabel polysilicon 65 -984 65 -984 0 3
rlabel polysilicon 68 -984 68 -984 0 4
rlabel polysilicon 72 -978 72 -978 0 1
rlabel polysilicon 72 -984 72 -984 0 3
rlabel polysilicon 79 -978 79 -978 0 1
rlabel polysilicon 79 -984 79 -984 0 3
rlabel polysilicon 86 -978 86 -978 0 1
rlabel polysilicon 86 -984 86 -984 0 3
rlabel polysilicon 93 -978 93 -978 0 1
rlabel polysilicon 96 -984 96 -984 0 4
rlabel polysilicon 100 -978 100 -978 0 1
rlabel polysilicon 100 -984 100 -984 0 3
rlabel polysilicon 107 -978 107 -978 0 1
rlabel polysilicon 110 -978 110 -978 0 2
rlabel polysilicon 110 -984 110 -984 0 4
rlabel polysilicon 114 -978 114 -978 0 1
rlabel polysilicon 114 -984 114 -984 0 3
rlabel polysilicon 121 -978 121 -978 0 1
rlabel polysilicon 121 -984 121 -984 0 3
rlabel polysilicon 128 -978 128 -978 0 1
rlabel polysilicon 128 -984 128 -984 0 3
rlabel polysilicon 135 -978 135 -978 0 1
rlabel polysilicon 135 -984 135 -984 0 3
rlabel polysilicon 142 -978 142 -978 0 1
rlabel polysilicon 142 -984 142 -984 0 3
rlabel polysilicon 145 -984 145 -984 0 4
rlabel polysilicon 149 -978 149 -978 0 1
rlabel polysilicon 149 -984 149 -984 0 3
rlabel polysilicon 156 -978 156 -978 0 1
rlabel polysilicon 156 -984 156 -984 0 3
rlabel polysilicon 159 -984 159 -984 0 4
rlabel polysilicon 163 -978 163 -978 0 1
rlabel polysilicon 163 -984 163 -984 0 3
rlabel polysilicon 170 -978 170 -978 0 1
rlabel polysilicon 170 -984 170 -984 0 3
rlabel polysilicon 177 -978 177 -978 0 1
rlabel polysilicon 177 -984 177 -984 0 3
rlabel polysilicon 184 -978 184 -978 0 1
rlabel polysilicon 187 -978 187 -978 0 2
rlabel polysilicon 184 -984 184 -984 0 3
rlabel polysilicon 191 -978 191 -978 0 1
rlabel polysilicon 191 -984 191 -984 0 3
rlabel polysilicon 198 -978 198 -978 0 1
rlabel polysilicon 198 -984 198 -984 0 3
rlabel polysilicon 205 -978 205 -978 0 1
rlabel polysilicon 205 -984 205 -984 0 3
rlabel polysilicon 212 -978 212 -978 0 1
rlabel polysilicon 212 -984 212 -984 0 3
rlabel polysilicon 219 -984 219 -984 0 3
rlabel polysilicon 226 -978 226 -978 0 1
rlabel polysilicon 226 -984 226 -984 0 3
rlabel polysilicon 233 -978 233 -978 0 1
rlabel polysilicon 236 -978 236 -978 0 2
rlabel polysilicon 236 -984 236 -984 0 4
rlabel polysilicon 240 -978 240 -978 0 1
rlabel polysilicon 240 -984 240 -984 0 3
rlabel polysilicon 247 -978 247 -978 0 1
rlabel polysilicon 247 -984 247 -984 0 3
rlabel polysilicon 254 -978 254 -978 0 1
rlabel polysilicon 254 -984 254 -984 0 3
rlabel polysilicon 261 -978 261 -978 0 1
rlabel polysilicon 261 -984 261 -984 0 3
rlabel polysilicon 268 -978 268 -978 0 1
rlabel polysilicon 268 -984 268 -984 0 3
rlabel polysilicon 275 -978 275 -978 0 1
rlabel polysilicon 275 -984 275 -984 0 3
rlabel polysilicon 282 -978 282 -978 0 1
rlabel polysilicon 282 -984 282 -984 0 3
rlabel polysilicon 289 -978 289 -978 0 1
rlabel polysilicon 289 -984 289 -984 0 3
rlabel polysilicon 296 -978 296 -978 0 1
rlabel polysilicon 296 -984 296 -984 0 3
rlabel polysilicon 303 -984 303 -984 0 3
rlabel polysilicon 310 -978 310 -978 0 1
rlabel polysilicon 310 -984 310 -984 0 3
rlabel polysilicon 317 -978 317 -978 0 1
rlabel polysilicon 317 -984 317 -984 0 3
rlabel polysilicon 324 -978 324 -978 0 1
rlabel polysilicon 324 -984 324 -984 0 3
rlabel polysilicon 331 -978 331 -978 0 1
rlabel polysilicon 331 -984 331 -984 0 3
rlabel polysilicon 338 -978 338 -978 0 1
rlabel polysilicon 338 -984 338 -984 0 3
rlabel polysilicon 345 -978 345 -978 0 1
rlabel polysilicon 345 -984 345 -984 0 3
rlabel polysilicon 352 -978 352 -978 0 1
rlabel polysilicon 352 -984 352 -984 0 3
rlabel polysilicon 359 -978 359 -978 0 1
rlabel polysilicon 359 -984 359 -984 0 3
rlabel polysilicon 366 -978 366 -978 0 1
rlabel polysilicon 366 -984 366 -984 0 3
rlabel polysilicon 373 -978 373 -978 0 1
rlabel polysilicon 373 -984 373 -984 0 3
rlabel polysilicon 380 -978 380 -978 0 1
rlabel polysilicon 380 -984 380 -984 0 3
rlabel polysilicon 390 -978 390 -978 0 2
rlabel polysilicon 387 -984 387 -984 0 3
rlabel polysilicon 390 -984 390 -984 0 4
rlabel polysilicon 394 -978 394 -978 0 1
rlabel polysilicon 394 -984 394 -984 0 3
rlabel polysilicon 401 -978 401 -978 0 1
rlabel polysilicon 401 -984 401 -984 0 3
rlabel polysilicon 408 -978 408 -978 0 1
rlabel polysilicon 408 -984 408 -984 0 3
rlabel polysilicon 415 -978 415 -978 0 1
rlabel polysilicon 415 -984 415 -984 0 3
rlabel polysilicon 422 -978 422 -978 0 1
rlabel polysilicon 422 -984 422 -984 0 3
rlabel polysilicon 429 -978 429 -978 0 1
rlabel polysilicon 429 -984 429 -984 0 3
rlabel polysilicon 436 -978 436 -978 0 1
rlabel polysilicon 436 -984 436 -984 0 3
rlabel polysilicon 443 -978 443 -978 0 1
rlabel polysilicon 443 -984 443 -984 0 3
rlabel polysilicon 450 -978 450 -978 0 1
rlabel polysilicon 450 -984 450 -984 0 3
rlabel polysilicon 457 -978 457 -978 0 1
rlabel polysilicon 460 -978 460 -978 0 2
rlabel polysilicon 457 -984 457 -984 0 3
rlabel polysilicon 464 -978 464 -978 0 1
rlabel polysilicon 464 -984 464 -984 0 3
rlabel polysilicon 471 -978 471 -978 0 1
rlabel polysilicon 471 -984 471 -984 0 3
rlabel polysilicon 478 -978 478 -978 0 1
rlabel polysilicon 478 -984 478 -984 0 3
rlabel polysilicon 485 -978 485 -978 0 1
rlabel polysilicon 485 -984 485 -984 0 3
rlabel polysilicon 492 -978 492 -978 0 1
rlabel polysilicon 492 -984 492 -984 0 3
rlabel polysilicon 499 -978 499 -978 0 1
rlabel polysilicon 499 -984 499 -984 0 3
rlabel polysilicon 506 -978 506 -978 0 1
rlabel polysilicon 506 -984 506 -984 0 3
rlabel polysilicon 513 -978 513 -978 0 1
rlabel polysilicon 513 -984 513 -984 0 3
rlabel polysilicon 520 -978 520 -978 0 1
rlabel polysilicon 520 -984 520 -984 0 3
rlabel polysilicon 527 -978 527 -978 0 1
rlabel polysilicon 527 -984 527 -984 0 3
rlabel polysilicon 534 -978 534 -978 0 1
rlabel polysilicon 537 -978 537 -978 0 2
rlabel polysilicon 534 -984 534 -984 0 3
rlabel polysilicon 537 -984 537 -984 0 4
rlabel polysilicon 541 -978 541 -978 0 1
rlabel polysilicon 544 -978 544 -978 0 2
rlabel polysilicon 548 -978 548 -978 0 1
rlabel polysilicon 548 -984 548 -984 0 3
rlabel polysilicon 555 -978 555 -978 0 1
rlabel polysilicon 555 -984 555 -984 0 3
rlabel polysilicon 562 -978 562 -978 0 1
rlabel polysilicon 562 -984 562 -984 0 3
rlabel polysilicon 569 -978 569 -978 0 1
rlabel polysilicon 569 -984 569 -984 0 3
rlabel polysilicon 576 -978 576 -978 0 1
rlabel polysilicon 576 -984 576 -984 0 3
rlabel polysilicon 583 -978 583 -978 0 1
rlabel polysilicon 583 -984 583 -984 0 3
rlabel polysilicon 590 -978 590 -978 0 1
rlabel polysilicon 590 -984 590 -984 0 3
rlabel polysilicon 597 -978 597 -978 0 1
rlabel polysilicon 597 -984 597 -984 0 3
rlabel polysilicon 604 -978 604 -978 0 1
rlabel polysilicon 604 -984 604 -984 0 3
rlabel polysilicon 607 -984 607 -984 0 4
rlabel polysilicon 611 -978 611 -978 0 1
rlabel polysilicon 611 -984 611 -984 0 3
rlabel polysilicon 618 -978 618 -978 0 1
rlabel polysilicon 618 -984 618 -984 0 3
rlabel polysilicon 625 -978 625 -978 0 1
rlabel polysilicon 625 -984 625 -984 0 3
rlabel polysilicon 632 -978 632 -978 0 1
rlabel polysilicon 632 -984 632 -984 0 3
rlabel polysilicon 639 -978 639 -978 0 1
rlabel polysilicon 639 -984 639 -984 0 3
rlabel polysilicon 646 -978 646 -978 0 1
rlabel polysilicon 646 -984 646 -984 0 3
rlabel polysilicon 653 -978 653 -978 0 1
rlabel polysilicon 653 -984 653 -984 0 3
rlabel polysilicon 660 -978 660 -978 0 1
rlabel polysilicon 660 -984 660 -984 0 3
rlabel polysilicon 667 -978 667 -978 0 1
rlabel polysilicon 667 -984 667 -984 0 3
rlabel polysilicon 674 -978 674 -978 0 1
rlabel polysilicon 674 -984 674 -984 0 3
rlabel polysilicon 684 -978 684 -978 0 2
rlabel polysilicon 681 -984 681 -984 0 3
rlabel polysilicon 684 -984 684 -984 0 4
rlabel polysilicon 688 -978 688 -978 0 1
rlabel polysilicon 688 -984 688 -984 0 3
rlabel polysilicon 695 -978 695 -978 0 1
rlabel polysilicon 695 -984 695 -984 0 3
rlabel polysilicon 702 -978 702 -978 0 1
rlabel polysilicon 702 -984 702 -984 0 3
rlabel polysilicon 709 -978 709 -978 0 1
rlabel polysilicon 709 -984 709 -984 0 3
rlabel polysilicon 716 -978 716 -978 0 1
rlabel polysilicon 716 -984 716 -984 0 3
rlabel polysilicon 726 -978 726 -978 0 2
rlabel polysilicon 723 -984 723 -984 0 3
rlabel polysilicon 726 -984 726 -984 0 4
rlabel polysilicon 730 -978 730 -978 0 1
rlabel polysilicon 730 -984 730 -984 0 3
rlabel polysilicon 740 -978 740 -978 0 2
rlabel polysilicon 737 -984 737 -984 0 3
rlabel polysilicon 740 -984 740 -984 0 4
rlabel polysilicon 744 -978 744 -978 0 1
rlabel polysilicon 747 -978 747 -978 0 2
rlabel polysilicon 744 -984 744 -984 0 3
rlabel polysilicon 747 -984 747 -984 0 4
rlabel polysilicon 754 -978 754 -978 0 2
rlabel polysilicon 751 -984 751 -984 0 3
rlabel polysilicon 754 -984 754 -984 0 4
rlabel polysilicon 758 -978 758 -978 0 1
rlabel polysilicon 758 -984 758 -984 0 3
rlabel polysilicon 765 -978 765 -978 0 1
rlabel polysilicon 765 -984 765 -984 0 3
rlabel polysilicon 772 -978 772 -978 0 1
rlabel polysilicon 775 -978 775 -978 0 2
rlabel polysilicon 772 -984 772 -984 0 3
rlabel polysilicon 775 -984 775 -984 0 4
rlabel polysilicon 779 -978 779 -978 0 1
rlabel polysilicon 779 -984 779 -984 0 3
rlabel polysilicon 786 -978 786 -978 0 1
rlabel polysilicon 786 -984 786 -984 0 3
rlabel polysilicon 793 -978 793 -978 0 1
rlabel polysilicon 793 -984 793 -984 0 3
rlabel polysilicon 800 -978 800 -978 0 1
rlabel polysilicon 800 -984 800 -984 0 3
rlabel polysilicon 807 -978 807 -978 0 1
rlabel polysilicon 807 -984 807 -984 0 3
rlabel polysilicon 814 -978 814 -978 0 1
rlabel polysilicon 814 -984 814 -984 0 3
rlabel polysilicon 821 -978 821 -978 0 1
rlabel polysilicon 821 -984 821 -984 0 3
rlabel polysilicon 828 -978 828 -978 0 1
rlabel polysilicon 828 -984 828 -984 0 3
rlabel polysilicon 835 -978 835 -978 0 1
rlabel polysilicon 835 -984 835 -984 0 3
rlabel polysilicon 842 -978 842 -978 0 1
rlabel polysilicon 842 -984 842 -984 0 3
rlabel polysilicon 849 -978 849 -978 0 1
rlabel polysilicon 849 -984 849 -984 0 3
rlabel polysilicon 856 -978 856 -978 0 1
rlabel polysilicon 856 -984 856 -984 0 3
rlabel polysilicon 863 -978 863 -978 0 1
rlabel polysilicon 863 -984 863 -984 0 3
rlabel polysilicon 870 -978 870 -978 0 1
rlabel polysilicon 870 -984 870 -984 0 3
rlabel polysilicon 877 -978 877 -978 0 1
rlabel polysilicon 877 -984 877 -984 0 3
rlabel polysilicon 884 -978 884 -978 0 1
rlabel polysilicon 884 -984 884 -984 0 3
rlabel polysilicon 891 -978 891 -978 0 1
rlabel polysilicon 891 -984 891 -984 0 3
rlabel polysilicon 898 -978 898 -978 0 1
rlabel polysilicon 898 -984 898 -984 0 3
rlabel polysilicon 905 -978 905 -978 0 1
rlabel polysilicon 905 -984 905 -984 0 3
rlabel polysilicon 915 -978 915 -978 0 2
rlabel polysilicon 912 -984 912 -984 0 3
rlabel polysilicon 915 -984 915 -984 0 4
rlabel polysilicon 922 -978 922 -978 0 2
rlabel polysilicon 919 -984 919 -984 0 3
rlabel polysilicon 922 -984 922 -984 0 4
rlabel polysilicon 926 -978 926 -978 0 1
rlabel polysilicon 926 -984 926 -984 0 3
rlabel polysilicon 933 -978 933 -978 0 1
rlabel polysilicon 933 -984 933 -984 0 3
rlabel polysilicon 940 -978 940 -978 0 1
rlabel polysilicon 943 -978 943 -978 0 2
rlabel polysilicon 940 -984 940 -984 0 3
rlabel polysilicon 943 -984 943 -984 0 4
rlabel polysilicon 947 -978 947 -978 0 1
rlabel polysilicon 947 -984 947 -984 0 3
rlabel polysilicon 954 -978 954 -978 0 1
rlabel polysilicon 954 -984 954 -984 0 3
rlabel polysilicon 961 -978 961 -978 0 1
rlabel polysilicon 961 -984 961 -984 0 3
rlabel polysilicon 968 -978 968 -978 0 1
rlabel polysilicon 968 -984 968 -984 0 3
rlabel polysilicon 975 -978 975 -978 0 1
rlabel polysilicon 975 -984 975 -984 0 3
rlabel polysilicon 982 -978 982 -978 0 1
rlabel polysilicon 985 -978 985 -978 0 2
rlabel polysilicon 982 -984 982 -984 0 3
rlabel polysilicon 985 -984 985 -984 0 4
rlabel polysilicon 989 -978 989 -978 0 1
rlabel polysilicon 989 -984 989 -984 0 3
rlabel polysilicon 996 -978 996 -978 0 1
rlabel polysilicon 996 -984 996 -984 0 3
rlabel polysilicon 1003 -978 1003 -978 0 1
rlabel polysilicon 1006 -978 1006 -978 0 2
rlabel polysilicon 1003 -984 1003 -984 0 3
rlabel polysilicon 1006 -984 1006 -984 0 4
rlabel polysilicon 1010 -978 1010 -978 0 1
rlabel polysilicon 1013 -978 1013 -978 0 2
rlabel polysilicon 1010 -984 1010 -984 0 3
rlabel polysilicon 1013 -984 1013 -984 0 4
rlabel polysilicon 1017 -978 1017 -978 0 1
rlabel polysilicon 1017 -984 1017 -984 0 3
rlabel polysilicon 1024 -978 1024 -978 0 1
rlabel polysilicon 1024 -984 1024 -984 0 3
rlabel polysilicon 1031 -978 1031 -978 0 1
rlabel polysilicon 1034 -978 1034 -978 0 2
rlabel polysilicon 1031 -984 1031 -984 0 3
rlabel polysilicon 1034 -984 1034 -984 0 4
rlabel polysilicon 1038 -978 1038 -978 0 1
rlabel polysilicon 1041 -978 1041 -978 0 2
rlabel polysilicon 1038 -984 1038 -984 0 3
rlabel polysilicon 1041 -984 1041 -984 0 4
rlabel polysilicon 1045 -978 1045 -978 0 1
rlabel polysilicon 1045 -984 1045 -984 0 3
rlabel polysilicon 1052 -978 1052 -978 0 1
rlabel polysilicon 1052 -984 1052 -984 0 3
rlabel polysilicon 1059 -978 1059 -978 0 1
rlabel polysilicon 1062 -978 1062 -978 0 2
rlabel polysilicon 1059 -984 1059 -984 0 3
rlabel polysilicon 1062 -984 1062 -984 0 4
rlabel polysilicon 1066 -978 1066 -978 0 1
rlabel polysilicon 1066 -984 1066 -984 0 3
rlabel polysilicon 1073 -978 1073 -978 0 1
rlabel polysilicon 1073 -984 1073 -984 0 3
rlabel polysilicon 1080 -978 1080 -978 0 1
rlabel polysilicon 1083 -978 1083 -978 0 2
rlabel polysilicon 1080 -984 1080 -984 0 3
rlabel polysilicon 1083 -984 1083 -984 0 4
rlabel polysilicon 1087 -978 1087 -978 0 1
rlabel polysilicon 1087 -984 1087 -984 0 3
rlabel polysilicon 1094 -978 1094 -978 0 1
rlabel polysilicon 1094 -984 1094 -984 0 3
rlabel polysilicon 1101 -978 1101 -978 0 1
rlabel polysilicon 1101 -984 1101 -984 0 3
rlabel polysilicon 1108 -978 1108 -978 0 1
rlabel polysilicon 1111 -978 1111 -978 0 2
rlabel polysilicon 1108 -984 1108 -984 0 3
rlabel polysilicon 1115 -978 1115 -978 0 1
rlabel polysilicon 1115 -984 1115 -984 0 3
rlabel polysilicon 1122 -978 1122 -978 0 1
rlabel polysilicon 1122 -984 1122 -984 0 3
rlabel polysilicon 1129 -978 1129 -978 0 1
rlabel polysilicon 1129 -984 1129 -984 0 3
rlabel polysilicon 1136 -978 1136 -978 0 1
rlabel polysilicon 1136 -984 1136 -984 0 3
rlabel polysilicon 1143 -978 1143 -978 0 1
rlabel polysilicon 1143 -984 1143 -984 0 3
rlabel polysilicon 1153 -978 1153 -978 0 2
rlabel polysilicon 1150 -984 1150 -984 0 3
rlabel polysilicon 1153 -984 1153 -984 0 4
rlabel polysilicon 1157 -978 1157 -978 0 1
rlabel polysilicon 1160 -978 1160 -978 0 2
rlabel polysilicon 1160 -984 1160 -984 0 4
rlabel polysilicon 1164 -978 1164 -978 0 1
rlabel polysilicon 1164 -984 1164 -984 0 3
rlabel polysilicon 1171 -978 1171 -978 0 1
rlabel polysilicon 1171 -984 1171 -984 0 3
rlabel polysilicon 1178 -978 1178 -978 0 1
rlabel polysilicon 1178 -984 1178 -984 0 3
rlabel polysilicon 1185 -978 1185 -978 0 1
rlabel polysilicon 1185 -984 1185 -984 0 3
rlabel polysilicon 1192 -978 1192 -978 0 1
rlabel polysilicon 1192 -984 1192 -984 0 3
rlabel polysilicon 1199 -978 1199 -978 0 1
rlabel polysilicon 1199 -984 1199 -984 0 3
rlabel polysilicon 1206 -978 1206 -978 0 1
rlabel polysilicon 1206 -984 1206 -984 0 3
rlabel polysilicon 1213 -978 1213 -978 0 1
rlabel polysilicon 1213 -984 1213 -984 0 3
rlabel polysilicon 1220 -978 1220 -978 0 1
rlabel polysilicon 1220 -984 1220 -984 0 3
rlabel polysilicon 1227 -984 1227 -984 0 3
rlabel polysilicon 1230 -984 1230 -984 0 4
rlabel polysilicon 1234 -978 1234 -978 0 1
rlabel polysilicon 1234 -984 1234 -984 0 3
rlabel polysilicon 1241 -978 1241 -978 0 1
rlabel polysilicon 1241 -984 1241 -984 0 3
rlabel polysilicon 1248 -978 1248 -978 0 1
rlabel polysilicon 1248 -984 1248 -984 0 3
rlabel polysilicon 1255 -978 1255 -978 0 1
rlabel polysilicon 1255 -984 1255 -984 0 3
rlabel polysilicon 1262 -978 1262 -978 0 1
rlabel polysilicon 1262 -984 1262 -984 0 3
rlabel polysilicon 1269 -978 1269 -978 0 1
rlabel polysilicon 1269 -984 1269 -984 0 3
rlabel polysilicon 1276 -978 1276 -978 0 1
rlabel polysilicon 1276 -984 1276 -984 0 3
rlabel polysilicon 1283 -978 1283 -978 0 1
rlabel polysilicon 1283 -984 1283 -984 0 3
rlabel polysilicon 1290 -978 1290 -978 0 1
rlabel polysilicon 1290 -984 1290 -984 0 3
rlabel polysilicon 1297 -978 1297 -978 0 1
rlabel polysilicon 1297 -984 1297 -984 0 3
rlabel polysilicon 1304 -978 1304 -978 0 1
rlabel polysilicon 1304 -984 1304 -984 0 3
rlabel polysilicon 1311 -978 1311 -978 0 1
rlabel polysilicon 1311 -984 1311 -984 0 3
rlabel polysilicon 1318 -978 1318 -978 0 1
rlabel polysilicon 1318 -984 1318 -984 0 3
rlabel polysilicon 1325 -978 1325 -978 0 1
rlabel polysilicon 1325 -984 1325 -984 0 3
rlabel polysilicon 1332 -978 1332 -978 0 1
rlabel polysilicon 1332 -984 1332 -984 0 3
rlabel polysilicon 1339 -978 1339 -978 0 1
rlabel polysilicon 1339 -984 1339 -984 0 3
rlabel polysilicon 1346 -978 1346 -978 0 1
rlabel polysilicon 1346 -984 1346 -984 0 3
rlabel polysilicon 1353 -978 1353 -978 0 1
rlabel polysilicon 1353 -984 1353 -984 0 3
rlabel polysilicon 1360 -978 1360 -978 0 1
rlabel polysilicon 1360 -984 1360 -984 0 3
rlabel polysilicon 1367 -978 1367 -978 0 1
rlabel polysilicon 1367 -984 1367 -984 0 3
rlabel polysilicon 1374 -978 1374 -978 0 1
rlabel polysilicon 1374 -984 1374 -984 0 3
rlabel polysilicon 1381 -978 1381 -978 0 1
rlabel polysilicon 1381 -984 1381 -984 0 3
rlabel polysilicon 1388 -978 1388 -978 0 1
rlabel polysilicon 1388 -984 1388 -984 0 3
rlabel polysilicon 1395 -978 1395 -978 0 1
rlabel polysilicon 1395 -984 1395 -984 0 3
rlabel polysilicon 1402 -978 1402 -978 0 1
rlabel polysilicon 1402 -984 1402 -984 0 3
rlabel polysilicon 1409 -978 1409 -978 0 1
rlabel polysilicon 1409 -984 1409 -984 0 3
rlabel polysilicon 1416 -978 1416 -978 0 1
rlabel polysilicon 1416 -984 1416 -984 0 3
rlabel polysilicon 1423 -978 1423 -978 0 1
rlabel polysilicon 1423 -984 1423 -984 0 3
rlabel polysilicon 1430 -978 1430 -978 0 1
rlabel polysilicon 1430 -984 1430 -984 0 3
rlabel polysilicon 1437 -978 1437 -978 0 1
rlabel polysilicon 1437 -984 1437 -984 0 3
rlabel polysilicon 1444 -978 1444 -978 0 1
rlabel polysilicon 1444 -984 1444 -984 0 3
rlabel polysilicon 1451 -978 1451 -978 0 1
rlabel polysilicon 1451 -984 1451 -984 0 3
rlabel polysilicon 1458 -978 1458 -978 0 1
rlabel polysilicon 1458 -984 1458 -984 0 3
rlabel polysilicon 1465 -978 1465 -978 0 1
rlabel polysilicon 1465 -984 1465 -984 0 3
rlabel polysilicon 1472 -978 1472 -978 0 1
rlabel polysilicon 1472 -984 1472 -984 0 3
rlabel polysilicon 1479 -978 1479 -978 0 1
rlabel polysilicon 1479 -984 1479 -984 0 3
rlabel polysilicon 1486 -978 1486 -978 0 1
rlabel polysilicon 1486 -984 1486 -984 0 3
rlabel polysilicon 1493 -978 1493 -978 0 1
rlabel polysilicon 1493 -984 1493 -984 0 3
rlabel polysilicon 1500 -978 1500 -978 0 1
rlabel polysilicon 1500 -984 1500 -984 0 3
rlabel polysilicon 1507 -978 1507 -978 0 1
rlabel polysilicon 1507 -984 1507 -984 0 3
rlabel polysilicon 1514 -978 1514 -978 0 1
rlabel polysilicon 1514 -984 1514 -984 0 3
rlabel polysilicon 1521 -978 1521 -978 0 1
rlabel polysilicon 1521 -984 1521 -984 0 3
rlabel polysilicon 1528 -978 1528 -978 0 1
rlabel polysilicon 1528 -984 1528 -984 0 3
rlabel polysilicon 1535 -978 1535 -978 0 1
rlabel polysilicon 1535 -984 1535 -984 0 3
rlabel polysilicon 1542 -978 1542 -978 0 1
rlabel polysilicon 1542 -984 1542 -984 0 3
rlabel polysilicon 1549 -978 1549 -978 0 1
rlabel polysilicon 1549 -984 1549 -984 0 3
rlabel polysilicon 1556 -978 1556 -978 0 1
rlabel polysilicon 1556 -984 1556 -984 0 3
rlabel polysilicon 1563 -978 1563 -978 0 1
rlabel polysilicon 1563 -984 1563 -984 0 3
rlabel polysilicon 1570 -978 1570 -978 0 1
rlabel polysilicon 1570 -984 1570 -984 0 3
rlabel polysilicon 1577 -978 1577 -978 0 1
rlabel polysilicon 1577 -984 1577 -984 0 3
rlabel polysilicon 1584 -978 1584 -978 0 1
rlabel polysilicon 1584 -984 1584 -984 0 3
rlabel polysilicon 1591 -978 1591 -978 0 1
rlabel polysilicon 1594 -978 1594 -978 0 2
rlabel polysilicon 1591 -984 1591 -984 0 3
rlabel polysilicon 1598 -978 1598 -978 0 1
rlabel polysilicon 1598 -984 1598 -984 0 3
rlabel polysilicon 1605 -978 1605 -978 0 1
rlabel polysilicon 1605 -984 1605 -984 0 3
rlabel polysilicon 1612 -978 1612 -978 0 1
rlabel polysilicon 1612 -984 1612 -984 0 3
rlabel polysilicon 1619 -978 1619 -978 0 1
rlabel polysilicon 1619 -984 1619 -984 0 3
rlabel polysilicon 1626 -978 1626 -978 0 1
rlabel polysilicon 1626 -984 1626 -984 0 3
rlabel polysilicon 1633 -978 1633 -978 0 1
rlabel polysilicon 1633 -984 1633 -984 0 3
rlabel polysilicon 1640 -978 1640 -978 0 1
rlabel polysilicon 1640 -984 1640 -984 0 3
rlabel polysilicon 1647 -978 1647 -978 0 1
rlabel polysilicon 1647 -984 1647 -984 0 3
rlabel polysilicon 1654 -978 1654 -978 0 1
rlabel polysilicon 1654 -984 1654 -984 0 3
rlabel polysilicon 1661 -978 1661 -978 0 1
rlabel polysilicon 1661 -984 1661 -984 0 3
rlabel polysilicon 1668 -978 1668 -978 0 1
rlabel polysilicon 1668 -984 1668 -984 0 3
rlabel polysilicon 1675 -978 1675 -978 0 1
rlabel polysilicon 1675 -984 1675 -984 0 3
rlabel polysilicon 1682 -978 1682 -978 0 1
rlabel polysilicon 1682 -984 1682 -984 0 3
rlabel polysilicon 1689 -978 1689 -978 0 1
rlabel polysilicon 1689 -984 1689 -984 0 3
rlabel polysilicon 1696 -978 1696 -978 0 1
rlabel polysilicon 1696 -984 1696 -984 0 3
rlabel polysilicon 1703 -978 1703 -978 0 1
rlabel polysilicon 1703 -984 1703 -984 0 3
rlabel polysilicon 1710 -978 1710 -978 0 1
rlabel polysilicon 1710 -984 1710 -984 0 3
rlabel polysilicon 1717 -978 1717 -978 0 1
rlabel polysilicon 1717 -984 1717 -984 0 3
rlabel polysilicon 1724 -978 1724 -978 0 1
rlabel polysilicon 1724 -984 1724 -984 0 3
rlabel polysilicon 1731 -978 1731 -978 0 1
rlabel polysilicon 1731 -984 1731 -984 0 3
rlabel polysilicon 1738 -978 1738 -978 0 1
rlabel polysilicon 1738 -984 1738 -984 0 3
rlabel polysilicon 1745 -978 1745 -978 0 1
rlabel polysilicon 1745 -984 1745 -984 0 3
rlabel polysilicon 1752 -978 1752 -978 0 1
rlabel polysilicon 1752 -984 1752 -984 0 3
rlabel polysilicon 1759 -978 1759 -978 0 1
rlabel polysilicon 1759 -984 1759 -984 0 3
rlabel polysilicon 1766 -978 1766 -978 0 1
rlabel polysilicon 1766 -984 1766 -984 0 3
rlabel polysilicon 1773 -978 1773 -978 0 1
rlabel polysilicon 1773 -984 1773 -984 0 3
rlabel polysilicon 1780 -978 1780 -978 0 1
rlabel polysilicon 1780 -984 1780 -984 0 3
rlabel polysilicon 1787 -978 1787 -978 0 1
rlabel polysilicon 1787 -984 1787 -984 0 3
rlabel polysilicon 1794 -978 1794 -978 0 1
rlabel polysilicon 1794 -984 1794 -984 0 3
rlabel polysilicon 1801 -978 1801 -978 0 1
rlabel polysilicon 1801 -984 1801 -984 0 3
rlabel polysilicon 1808 -978 1808 -978 0 1
rlabel polysilicon 1808 -984 1808 -984 0 3
rlabel polysilicon 1815 -978 1815 -978 0 1
rlabel polysilicon 1815 -984 1815 -984 0 3
rlabel polysilicon 1822 -978 1822 -978 0 1
rlabel polysilicon 1822 -984 1822 -984 0 3
rlabel polysilicon 1829 -978 1829 -978 0 1
rlabel polysilicon 1829 -984 1829 -984 0 3
rlabel polysilicon 1836 -978 1836 -978 0 1
rlabel polysilicon 1836 -984 1836 -984 0 3
rlabel polysilicon 1843 -978 1843 -978 0 1
rlabel polysilicon 1843 -984 1843 -984 0 3
rlabel polysilicon 1850 -978 1850 -978 0 1
rlabel polysilicon 1850 -984 1850 -984 0 3
rlabel polysilicon 1857 -978 1857 -978 0 1
rlabel polysilicon 1857 -984 1857 -984 0 3
rlabel polysilicon 1864 -978 1864 -978 0 1
rlabel polysilicon 1864 -984 1864 -984 0 3
rlabel polysilicon 1871 -978 1871 -978 0 1
rlabel polysilicon 1871 -984 1871 -984 0 3
rlabel polysilicon 1878 -978 1878 -978 0 1
rlabel polysilicon 1881 -978 1881 -978 0 2
rlabel polysilicon 1878 -984 1878 -984 0 3
rlabel polysilicon 1881 -984 1881 -984 0 4
rlabel polysilicon 1885 -978 1885 -978 0 1
rlabel polysilicon 1885 -984 1885 -984 0 3
rlabel polysilicon 1892 -978 1892 -978 0 1
rlabel polysilicon 1892 -984 1892 -984 0 3
rlabel polysilicon 1899 -978 1899 -978 0 1
rlabel polysilicon 1899 -984 1899 -984 0 3
rlabel polysilicon 1902 -984 1902 -984 0 4
rlabel polysilicon 1906 -978 1906 -978 0 1
rlabel polysilicon 1906 -984 1906 -984 0 3
rlabel polysilicon 1913 -978 1913 -978 0 1
rlabel polysilicon 1916 -978 1916 -978 0 2
rlabel polysilicon 1920 -978 1920 -978 0 1
rlabel polysilicon 1920 -984 1920 -984 0 3
rlabel polysilicon 1927 -978 1927 -978 0 1
rlabel polysilicon 1927 -984 1927 -984 0 3
rlabel polysilicon 1934 -978 1934 -978 0 1
rlabel polysilicon 1934 -984 1934 -984 0 3
rlabel polysilicon 1941 -978 1941 -978 0 1
rlabel polysilicon 1941 -984 1941 -984 0 3
rlabel polysilicon 1948 -978 1948 -978 0 1
rlabel polysilicon 1948 -984 1948 -984 0 3
rlabel polysilicon 1955 -978 1955 -978 0 1
rlabel polysilicon 1955 -984 1955 -984 0 3
rlabel polysilicon 9 -1109 9 -1109 0 1
rlabel polysilicon 9 -1115 9 -1115 0 3
rlabel polysilicon 16 -1109 16 -1109 0 1
rlabel polysilicon 16 -1115 16 -1115 0 3
rlabel polysilicon 23 -1109 23 -1109 0 1
rlabel polysilicon 23 -1115 23 -1115 0 3
rlabel polysilicon 30 -1109 30 -1109 0 1
rlabel polysilicon 30 -1115 30 -1115 0 3
rlabel polysilicon 37 -1109 37 -1109 0 1
rlabel polysilicon 37 -1115 37 -1115 0 3
rlabel polysilicon 47 -1109 47 -1109 0 2
rlabel polysilicon 44 -1115 44 -1115 0 3
rlabel polysilicon 47 -1115 47 -1115 0 4
rlabel polysilicon 51 -1109 51 -1109 0 1
rlabel polysilicon 51 -1115 51 -1115 0 3
rlabel polysilicon 58 -1109 58 -1109 0 1
rlabel polysilicon 58 -1115 58 -1115 0 3
rlabel polysilicon 65 -1109 65 -1109 0 1
rlabel polysilicon 68 -1109 68 -1109 0 2
rlabel polysilicon 65 -1115 65 -1115 0 3
rlabel polysilicon 72 -1109 72 -1109 0 1
rlabel polysilicon 72 -1115 72 -1115 0 3
rlabel polysilicon 79 -1109 79 -1109 0 1
rlabel polysilicon 82 -1109 82 -1109 0 2
rlabel polysilicon 82 -1115 82 -1115 0 4
rlabel polysilicon 86 -1109 86 -1109 0 1
rlabel polysilicon 86 -1115 86 -1115 0 3
rlabel polysilicon 93 -1109 93 -1109 0 1
rlabel polysilicon 93 -1115 93 -1115 0 3
rlabel polysilicon 100 -1109 100 -1109 0 1
rlabel polysilicon 100 -1115 100 -1115 0 3
rlabel polysilicon 107 -1109 107 -1109 0 1
rlabel polysilicon 107 -1115 107 -1115 0 3
rlabel polysilicon 114 -1109 114 -1109 0 1
rlabel polysilicon 114 -1115 114 -1115 0 3
rlabel polysilicon 121 -1109 121 -1109 0 1
rlabel polysilicon 121 -1115 121 -1115 0 3
rlabel polysilicon 128 -1109 128 -1109 0 1
rlabel polysilicon 128 -1115 128 -1115 0 3
rlabel polysilicon 131 -1115 131 -1115 0 4
rlabel polysilicon 135 -1109 135 -1109 0 1
rlabel polysilicon 135 -1115 135 -1115 0 3
rlabel polysilicon 142 -1109 142 -1109 0 1
rlabel polysilicon 142 -1115 142 -1115 0 3
rlabel polysilicon 149 -1109 149 -1109 0 1
rlabel polysilicon 149 -1115 149 -1115 0 3
rlabel polysilicon 156 -1109 156 -1109 0 1
rlabel polysilicon 156 -1115 156 -1115 0 3
rlabel polysilicon 163 -1109 163 -1109 0 1
rlabel polysilicon 163 -1115 163 -1115 0 3
rlabel polysilicon 170 -1109 170 -1109 0 1
rlabel polysilicon 170 -1115 170 -1115 0 3
rlabel polysilicon 177 -1109 177 -1109 0 1
rlabel polysilicon 177 -1115 177 -1115 0 3
rlabel polysilicon 184 -1109 184 -1109 0 1
rlabel polysilicon 184 -1115 184 -1115 0 3
rlabel polysilicon 191 -1109 191 -1109 0 1
rlabel polysilicon 191 -1115 191 -1115 0 3
rlabel polysilicon 198 -1109 198 -1109 0 1
rlabel polysilicon 198 -1115 198 -1115 0 3
rlabel polysilicon 205 -1109 205 -1109 0 1
rlabel polysilicon 205 -1115 205 -1115 0 3
rlabel polysilicon 212 -1109 212 -1109 0 1
rlabel polysilicon 215 -1109 215 -1109 0 2
rlabel polysilicon 212 -1115 212 -1115 0 3
rlabel polysilicon 219 -1109 219 -1109 0 1
rlabel polysilicon 222 -1115 222 -1115 0 4
rlabel polysilicon 226 -1109 226 -1109 0 1
rlabel polysilicon 226 -1115 226 -1115 0 3
rlabel polysilicon 233 -1109 233 -1109 0 1
rlabel polysilicon 233 -1115 233 -1115 0 3
rlabel polysilicon 240 -1109 240 -1109 0 1
rlabel polysilicon 240 -1115 240 -1115 0 3
rlabel polysilicon 247 -1109 247 -1109 0 1
rlabel polysilicon 247 -1115 247 -1115 0 3
rlabel polysilicon 254 -1109 254 -1109 0 1
rlabel polysilicon 254 -1115 254 -1115 0 3
rlabel polysilicon 261 -1109 261 -1109 0 1
rlabel polysilicon 261 -1115 261 -1115 0 3
rlabel polysilicon 268 -1109 268 -1109 0 1
rlabel polysilicon 268 -1115 268 -1115 0 3
rlabel polysilicon 275 -1109 275 -1109 0 1
rlabel polysilicon 275 -1115 275 -1115 0 3
rlabel polysilicon 282 -1109 282 -1109 0 1
rlabel polysilicon 282 -1115 282 -1115 0 3
rlabel polysilicon 289 -1109 289 -1109 0 1
rlabel polysilicon 289 -1115 289 -1115 0 3
rlabel polysilicon 296 -1109 296 -1109 0 1
rlabel polysilicon 296 -1115 296 -1115 0 3
rlabel polysilicon 303 -1109 303 -1109 0 1
rlabel polysilicon 303 -1115 303 -1115 0 3
rlabel polysilicon 310 -1109 310 -1109 0 1
rlabel polysilicon 313 -1115 313 -1115 0 4
rlabel polysilicon 317 -1109 317 -1109 0 1
rlabel polysilicon 317 -1115 317 -1115 0 3
rlabel polysilicon 324 -1109 324 -1109 0 1
rlabel polysilicon 324 -1115 324 -1115 0 3
rlabel polysilicon 331 -1109 331 -1109 0 1
rlabel polysilicon 331 -1115 331 -1115 0 3
rlabel polysilicon 338 -1109 338 -1109 0 1
rlabel polysilicon 338 -1115 338 -1115 0 3
rlabel polysilicon 345 -1109 345 -1109 0 1
rlabel polysilicon 345 -1115 345 -1115 0 3
rlabel polysilicon 352 -1109 352 -1109 0 1
rlabel polysilicon 352 -1115 352 -1115 0 3
rlabel polysilicon 359 -1109 359 -1109 0 1
rlabel polysilicon 359 -1115 359 -1115 0 3
rlabel polysilicon 366 -1109 366 -1109 0 1
rlabel polysilicon 366 -1115 366 -1115 0 3
rlabel polysilicon 373 -1109 373 -1109 0 1
rlabel polysilicon 373 -1115 373 -1115 0 3
rlabel polysilicon 380 -1109 380 -1109 0 1
rlabel polysilicon 380 -1115 380 -1115 0 3
rlabel polysilicon 387 -1109 387 -1109 0 1
rlabel polysilicon 394 -1109 394 -1109 0 1
rlabel polysilicon 397 -1109 397 -1109 0 2
rlabel polysilicon 394 -1115 394 -1115 0 3
rlabel polysilicon 401 -1109 401 -1109 0 1
rlabel polysilicon 401 -1115 401 -1115 0 3
rlabel polysilicon 408 -1109 408 -1109 0 1
rlabel polysilicon 408 -1115 408 -1115 0 3
rlabel polysilicon 415 -1109 415 -1109 0 1
rlabel polysilicon 415 -1115 415 -1115 0 3
rlabel polysilicon 422 -1109 422 -1109 0 1
rlabel polysilicon 422 -1115 422 -1115 0 3
rlabel polysilicon 429 -1109 429 -1109 0 1
rlabel polysilicon 429 -1115 429 -1115 0 3
rlabel polysilicon 436 -1109 436 -1109 0 1
rlabel polysilicon 436 -1115 436 -1115 0 3
rlabel polysilicon 443 -1109 443 -1109 0 1
rlabel polysilicon 443 -1115 443 -1115 0 3
rlabel polysilicon 450 -1109 450 -1109 0 1
rlabel polysilicon 453 -1109 453 -1109 0 2
rlabel polysilicon 450 -1115 450 -1115 0 3
rlabel polysilicon 453 -1115 453 -1115 0 4
rlabel polysilicon 457 -1109 457 -1109 0 1
rlabel polysilicon 457 -1115 457 -1115 0 3
rlabel polysilicon 464 -1109 464 -1109 0 1
rlabel polysilicon 464 -1115 464 -1115 0 3
rlabel polysilicon 471 -1109 471 -1109 0 1
rlabel polysilicon 471 -1115 471 -1115 0 3
rlabel polysilicon 478 -1109 478 -1109 0 1
rlabel polysilicon 478 -1115 478 -1115 0 3
rlabel polysilicon 485 -1109 485 -1109 0 1
rlabel polysilicon 485 -1115 485 -1115 0 3
rlabel polysilicon 492 -1109 492 -1109 0 1
rlabel polysilicon 492 -1115 492 -1115 0 3
rlabel polysilicon 499 -1109 499 -1109 0 1
rlabel polysilicon 499 -1115 499 -1115 0 3
rlabel polysilicon 506 -1109 506 -1109 0 1
rlabel polysilicon 506 -1115 506 -1115 0 3
rlabel polysilicon 513 -1109 513 -1109 0 1
rlabel polysilicon 513 -1115 513 -1115 0 3
rlabel polysilicon 520 -1109 520 -1109 0 1
rlabel polysilicon 520 -1115 520 -1115 0 3
rlabel polysilicon 523 -1115 523 -1115 0 4
rlabel polysilicon 527 -1109 527 -1109 0 1
rlabel polysilicon 527 -1115 527 -1115 0 3
rlabel polysilicon 534 -1109 534 -1109 0 1
rlabel polysilicon 534 -1115 534 -1115 0 3
rlabel polysilicon 541 -1109 541 -1109 0 1
rlabel polysilicon 541 -1115 541 -1115 0 3
rlabel polysilicon 548 -1109 548 -1109 0 1
rlabel polysilicon 548 -1115 548 -1115 0 3
rlabel polysilicon 555 -1109 555 -1109 0 1
rlabel polysilicon 555 -1115 555 -1115 0 3
rlabel polysilicon 565 -1109 565 -1109 0 2
rlabel polysilicon 562 -1115 562 -1115 0 3
rlabel polysilicon 565 -1115 565 -1115 0 4
rlabel polysilicon 569 -1109 569 -1109 0 1
rlabel polysilicon 572 -1109 572 -1109 0 2
rlabel polysilicon 569 -1115 569 -1115 0 3
rlabel polysilicon 572 -1115 572 -1115 0 4
rlabel polysilicon 576 -1109 576 -1109 0 1
rlabel polysilicon 579 -1109 579 -1109 0 2
rlabel polysilicon 576 -1115 576 -1115 0 3
rlabel polysilicon 579 -1115 579 -1115 0 4
rlabel polysilicon 583 -1109 583 -1109 0 1
rlabel polysilicon 583 -1115 583 -1115 0 3
rlabel polysilicon 590 -1109 590 -1109 0 1
rlabel polysilicon 590 -1115 590 -1115 0 3
rlabel polysilicon 597 -1109 597 -1109 0 1
rlabel polysilicon 597 -1115 597 -1115 0 3
rlabel polysilicon 604 -1109 604 -1109 0 1
rlabel polysilicon 604 -1115 604 -1115 0 3
rlabel polysilicon 611 -1109 611 -1109 0 1
rlabel polysilicon 611 -1115 611 -1115 0 3
rlabel polysilicon 618 -1109 618 -1109 0 1
rlabel polysilicon 618 -1115 618 -1115 0 3
rlabel polysilicon 625 -1109 625 -1109 0 1
rlabel polysilicon 628 -1109 628 -1109 0 2
rlabel polysilicon 625 -1115 625 -1115 0 3
rlabel polysilicon 628 -1115 628 -1115 0 4
rlabel polysilicon 632 -1109 632 -1109 0 1
rlabel polysilicon 635 -1109 635 -1109 0 2
rlabel polysilicon 632 -1115 632 -1115 0 3
rlabel polysilicon 639 -1109 639 -1109 0 1
rlabel polysilicon 639 -1115 639 -1115 0 3
rlabel polysilicon 646 -1109 646 -1109 0 1
rlabel polysilicon 649 -1109 649 -1109 0 2
rlabel polysilicon 646 -1115 646 -1115 0 3
rlabel polysilicon 653 -1109 653 -1109 0 1
rlabel polysilicon 656 -1109 656 -1109 0 2
rlabel polysilicon 653 -1115 653 -1115 0 3
rlabel polysilicon 656 -1115 656 -1115 0 4
rlabel polysilicon 660 -1109 660 -1109 0 1
rlabel polysilicon 660 -1115 660 -1115 0 3
rlabel polysilicon 667 -1109 667 -1109 0 1
rlabel polysilicon 667 -1115 667 -1115 0 3
rlabel polysilicon 674 -1109 674 -1109 0 1
rlabel polysilicon 674 -1115 674 -1115 0 3
rlabel polysilicon 681 -1109 681 -1109 0 1
rlabel polysilicon 684 -1109 684 -1109 0 2
rlabel polysilicon 681 -1115 681 -1115 0 3
rlabel polysilicon 684 -1115 684 -1115 0 4
rlabel polysilicon 688 -1109 688 -1109 0 1
rlabel polysilicon 688 -1115 688 -1115 0 3
rlabel polysilicon 695 -1109 695 -1109 0 1
rlabel polysilicon 695 -1115 695 -1115 0 3
rlabel polysilicon 702 -1109 702 -1109 0 1
rlabel polysilicon 702 -1115 702 -1115 0 3
rlabel polysilicon 709 -1109 709 -1109 0 1
rlabel polysilicon 709 -1115 709 -1115 0 3
rlabel polysilicon 716 -1109 716 -1109 0 1
rlabel polysilicon 716 -1115 716 -1115 0 3
rlabel polysilicon 723 -1109 723 -1109 0 1
rlabel polysilicon 723 -1115 723 -1115 0 3
rlabel polysilicon 730 -1109 730 -1109 0 1
rlabel polysilicon 733 -1109 733 -1109 0 2
rlabel polysilicon 730 -1115 730 -1115 0 3
rlabel polysilicon 733 -1115 733 -1115 0 4
rlabel polysilicon 737 -1109 737 -1109 0 1
rlabel polysilicon 740 -1109 740 -1109 0 2
rlabel polysilicon 737 -1115 737 -1115 0 3
rlabel polysilicon 740 -1115 740 -1115 0 4
rlabel polysilicon 744 -1109 744 -1109 0 1
rlabel polysilicon 744 -1115 744 -1115 0 3
rlabel polysilicon 747 -1115 747 -1115 0 4
rlabel polysilicon 751 -1109 751 -1109 0 1
rlabel polysilicon 751 -1115 751 -1115 0 3
rlabel polysilicon 754 -1115 754 -1115 0 4
rlabel polysilicon 758 -1109 758 -1109 0 1
rlabel polysilicon 761 -1109 761 -1109 0 2
rlabel polysilicon 761 -1115 761 -1115 0 4
rlabel polysilicon 765 -1109 765 -1109 0 1
rlabel polysilicon 765 -1115 765 -1115 0 3
rlabel polysilicon 772 -1109 772 -1109 0 1
rlabel polysilicon 772 -1115 772 -1115 0 3
rlabel polysilicon 779 -1109 779 -1109 0 1
rlabel polysilicon 782 -1109 782 -1109 0 2
rlabel polysilicon 779 -1115 779 -1115 0 3
rlabel polysilicon 782 -1115 782 -1115 0 4
rlabel polysilicon 786 -1109 786 -1109 0 1
rlabel polysilicon 789 -1109 789 -1109 0 2
rlabel polysilicon 789 -1115 789 -1115 0 4
rlabel polysilicon 793 -1109 793 -1109 0 1
rlabel polysilicon 793 -1115 793 -1115 0 3
rlabel polysilicon 800 -1109 800 -1109 0 1
rlabel polysilicon 800 -1115 800 -1115 0 3
rlabel polysilicon 807 -1109 807 -1109 0 1
rlabel polysilicon 807 -1115 807 -1115 0 3
rlabel polysilicon 814 -1109 814 -1109 0 1
rlabel polysilicon 814 -1115 814 -1115 0 3
rlabel polysilicon 821 -1109 821 -1109 0 1
rlabel polysilicon 821 -1115 821 -1115 0 3
rlabel polysilicon 828 -1109 828 -1109 0 1
rlabel polysilicon 828 -1115 828 -1115 0 3
rlabel polysilicon 835 -1109 835 -1109 0 1
rlabel polysilicon 835 -1115 835 -1115 0 3
rlabel polysilicon 842 -1109 842 -1109 0 1
rlabel polysilicon 842 -1115 842 -1115 0 3
rlabel polysilicon 849 -1109 849 -1109 0 1
rlabel polysilicon 849 -1115 849 -1115 0 3
rlabel polysilicon 852 -1115 852 -1115 0 4
rlabel polysilicon 856 -1109 856 -1109 0 1
rlabel polysilicon 856 -1115 856 -1115 0 3
rlabel polysilicon 863 -1109 863 -1109 0 1
rlabel polysilicon 866 -1109 866 -1109 0 2
rlabel polysilicon 863 -1115 863 -1115 0 3
rlabel polysilicon 866 -1115 866 -1115 0 4
rlabel polysilicon 870 -1109 870 -1109 0 1
rlabel polysilicon 870 -1115 870 -1115 0 3
rlabel polysilicon 877 -1109 877 -1109 0 1
rlabel polysilicon 877 -1115 877 -1115 0 3
rlabel polysilicon 884 -1109 884 -1109 0 1
rlabel polysilicon 884 -1115 884 -1115 0 3
rlabel polysilicon 891 -1109 891 -1109 0 1
rlabel polysilicon 894 -1109 894 -1109 0 2
rlabel polysilicon 891 -1115 891 -1115 0 3
rlabel polysilicon 894 -1115 894 -1115 0 4
rlabel polysilicon 898 -1109 898 -1109 0 1
rlabel polysilicon 898 -1115 898 -1115 0 3
rlabel polysilicon 905 -1109 905 -1109 0 1
rlabel polysilicon 905 -1115 905 -1115 0 3
rlabel polysilicon 912 -1109 912 -1109 0 1
rlabel polysilicon 912 -1115 912 -1115 0 3
rlabel polysilicon 919 -1109 919 -1109 0 1
rlabel polysilicon 919 -1115 919 -1115 0 3
rlabel polysilicon 926 -1109 926 -1109 0 1
rlabel polysilicon 926 -1115 926 -1115 0 3
rlabel polysilicon 933 -1109 933 -1109 0 1
rlabel polysilicon 933 -1115 933 -1115 0 3
rlabel polysilicon 940 -1109 940 -1109 0 1
rlabel polysilicon 940 -1115 940 -1115 0 3
rlabel polysilicon 947 -1109 947 -1109 0 1
rlabel polysilicon 947 -1115 947 -1115 0 3
rlabel polysilicon 954 -1109 954 -1109 0 1
rlabel polysilicon 957 -1109 957 -1109 0 2
rlabel polysilicon 954 -1115 954 -1115 0 3
rlabel polysilicon 957 -1115 957 -1115 0 4
rlabel polysilicon 961 -1109 961 -1109 0 1
rlabel polysilicon 961 -1115 961 -1115 0 3
rlabel polysilicon 968 -1109 968 -1109 0 1
rlabel polysilicon 968 -1115 968 -1115 0 3
rlabel polysilicon 975 -1109 975 -1109 0 1
rlabel polysilicon 975 -1115 975 -1115 0 3
rlabel polysilicon 982 -1109 982 -1109 0 1
rlabel polysilicon 982 -1115 982 -1115 0 3
rlabel polysilicon 989 -1109 989 -1109 0 1
rlabel polysilicon 989 -1115 989 -1115 0 3
rlabel polysilicon 996 -1109 996 -1109 0 1
rlabel polysilicon 996 -1115 996 -1115 0 3
rlabel polysilicon 1003 -1109 1003 -1109 0 1
rlabel polysilicon 1003 -1115 1003 -1115 0 3
rlabel polysilicon 1010 -1109 1010 -1109 0 1
rlabel polysilicon 1010 -1115 1010 -1115 0 3
rlabel polysilicon 1017 -1109 1017 -1109 0 1
rlabel polysilicon 1020 -1109 1020 -1109 0 2
rlabel polysilicon 1017 -1115 1017 -1115 0 3
rlabel polysilicon 1020 -1115 1020 -1115 0 4
rlabel polysilicon 1024 -1109 1024 -1109 0 1
rlabel polysilicon 1024 -1115 1024 -1115 0 3
rlabel polysilicon 1031 -1109 1031 -1109 0 1
rlabel polysilicon 1031 -1115 1031 -1115 0 3
rlabel polysilicon 1038 -1109 1038 -1109 0 1
rlabel polysilicon 1038 -1115 1038 -1115 0 3
rlabel polysilicon 1045 -1109 1045 -1109 0 1
rlabel polysilicon 1048 -1109 1048 -1109 0 2
rlabel polysilicon 1045 -1115 1045 -1115 0 3
rlabel polysilicon 1048 -1115 1048 -1115 0 4
rlabel polysilicon 1052 -1109 1052 -1109 0 1
rlabel polysilicon 1052 -1115 1052 -1115 0 3
rlabel polysilicon 1059 -1109 1059 -1109 0 1
rlabel polysilicon 1059 -1115 1059 -1115 0 3
rlabel polysilicon 1066 -1109 1066 -1109 0 1
rlabel polysilicon 1066 -1115 1066 -1115 0 3
rlabel polysilicon 1073 -1109 1073 -1109 0 1
rlabel polysilicon 1073 -1115 1073 -1115 0 3
rlabel polysilicon 1080 -1109 1080 -1109 0 1
rlabel polysilicon 1080 -1115 1080 -1115 0 3
rlabel polysilicon 1087 -1109 1087 -1109 0 1
rlabel polysilicon 1087 -1115 1087 -1115 0 3
rlabel polysilicon 1094 -1109 1094 -1109 0 1
rlabel polysilicon 1094 -1115 1094 -1115 0 3
rlabel polysilicon 1101 -1109 1101 -1109 0 1
rlabel polysilicon 1101 -1115 1101 -1115 0 3
rlabel polysilicon 1108 -1109 1108 -1109 0 1
rlabel polysilicon 1108 -1115 1108 -1115 0 3
rlabel polysilicon 1115 -1109 1115 -1109 0 1
rlabel polysilicon 1115 -1115 1115 -1115 0 3
rlabel polysilicon 1122 -1109 1122 -1109 0 1
rlabel polysilicon 1122 -1115 1122 -1115 0 3
rlabel polysilicon 1129 -1109 1129 -1109 0 1
rlabel polysilicon 1129 -1115 1129 -1115 0 3
rlabel polysilicon 1136 -1109 1136 -1109 0 1
rlabel polysilicon 1139 -1109 1139 -1109 0 2
rlabel polysilicon 1136 -1115 1136 -1115 0 3
rlabel polysilicon 1139 -1115 1139 -1115 0 4
rlabel polysilicon 1143 -1109 1143 -1109 0 1
rlabel polysilicon 1143 -1115 1143 -1115 0 3
rlabel polysilicon 1150 -1109 1150 -1109 0 1
rlabel polysilicon 1153 -1109 1153 -1109 0 2
rlabel polysilicon 1153 -1115 1153 -1115 0 4
rlabel polysilicon 1157 -1109 1157 -1109 0 1
rlabel polysilicon 1157 -1115 1157 -1115 0 3
rlabel polysilicon 1164 -1109 1164 -1109 0 1
rlabel polysilicon 1164 -1115 1164 -1115 0 3
rlabel polysilicon 1171 -1109 1171 -1109 0 1
rlabel polysilicon 1171 -1115 1171 -1115 0 3
rlabel polysilicon 1178 -1109 1178 -1109 0 1
rlabel polysilicon 1178 -1115 1178 -1115 0 3
rlabel polysilicon 1185 -1109 1185 -1109 0 1
rlabel polysilicon 1185 -1115 1185 -1115 0 3
rlabel polysilicon 1192 -1109 1192 -1109 0 1
rlabel polysilicon 1192 -1115 1192 -1115 0 3
rlabel polysilicon 1199 -1109 1199 -1109 0 1
rlabel polysilicon 1199 -1115 1199 -1115 0 3
rlabel polysilicon 1206 -1109 1206 -1109 0 1
rlabel polysilicon 1206 -1115 1206 -1115 0 3
rlabel polysilicon 1213 -1109 1213 -1109 0 1
rlabel polysilicon 1213 -1115 1213 -1115 0 3
rlabel polysilicon 1220 -1109 1220 -1109 0 1
rlabel polysilicon 1220 -1115 1220 -1115 0 3
rlabel polysilicon 1227 -1109 1227 -1109 0 1
rlabel polysilicon 1230 -1109 1230 -1109 0 2
rlabel polysilicon 1230 -1115 1230 -1115 0 4
rlabel polysilicon 1234 -1109 1234 -1109 0 1
rlabel polysilicon 1234 -1115 1234 -1115 0 3
rlabel polysilicon 1241 -1109 1241 -1109 0 1
rlabel polysilicon 1241 -1115 1241 -1115 0 3
rlabel polysilicon 1248 -1109 1248 -1109 0 1
rlabel polysilicon 1248 -1115 1248 -1115 0 3
rlabel polysilicon 1255 -1109 1255 -1109 0 1
rlabel polysilicon 1255 -1115 1255 -1115 0 3
rlabel polysilicon 1262 -1109 1262 -1109 0 1
rlabel polysilicon 1262 -1115 1262 -1115 0 3
rlabel polysilicon 1269 -1109 1269 -1109 0 1
rlabel polysilicon 1269 -1115 1269 -1115 0 3
rlabel polysilicon 1276 -1109 1276 -1109 0 1
rlabel polysilicon 1276 -1115 1276 -1115 0 3
rlabel polysilicon 1283 -1109 1283 -1109 0 1
rlabel polysilicon 1283 -1115 1283 -1115 0 3
rlabel polysilicon 1290 -1109 1290 -1109 0 1
rlabel polysilicon 1290 -1115 1290 -1115 0 3
rlabel polysilicon 1297 -1109 1297 -1109 0 1
rlabel polysilicon 1297 -1115 1297 -1115 0 3
rlabel polysilicon 1304 -1109 1304 -1109 0 1
rlabel polysilicon 1304 -1115 1304 -1115 0 3
rlabel polysilicon 1311 -1109 1311 -1109 0 1
rlabel polysilicon 1311 -1115 1311 -1115 0 3
rlabel polysilicon 1318 -1109 1318 -1109 0 1
rlabel polysilicon 1318 -1115 1318 -1115 0 3
rlabel polysilicon 1325 -1109 1325 -1109 0 1
rlabel polysilicon 1325 -1115 1325 -1115 0 3
rlabel polysilicon 1332 -1109 1332 -1109 0 1
rlabel polysilicon 1332 -1115 1332 -1115 0 3
rlabel polysilicon 1339 -1109 1339 -1109 0 1
rlabel polysilicon 1339 -1115 1339 -1115 0 3
rlabel polysilicon 1346 -1109 1346 -1109 0 1
rlabel polysilicon 1346 -1115 1346 -1115 0 3
rlabel polysilicon 1353 -1109 1353 -1109 0 1
rlabel polysilicon 1353 -1115 1353 -1115 0 3
rlabel polysilicon 1360 -1109 1360 -1109 0 1
rlabel polysilicon 1360 -1115 1360 -1115 0 3
rlabel polysilicon 1367 -1109 1367 -1109 0 1
rlabel polysilicon 1367 -1115 1367 -1115 0 3
rlabel polysilicon 1374 -1109 1374 -1109 0 1
rlabel polysilicon 1374 -1115 1374 -1115 0 3
rlabel polysilicon 1381 -1109 1381 -1109 0 1
rlabel polysilicon 1381 -1115 1381 -1115 0 3
rlabel polysilicon 1388 -1109 1388 -1109 0 1
rlabel polysilicon 1388 -1115 1388 -1115 0 3
rlabel polysilicon 1395 -1109 1395 -1109 0 1
rlabel polysilicon 1395 -1115 1395 -1115 0 3
rlabel polysilicon 1402 -1109 1402 -1109 0 1
rlabel polysilicon 1402 -1115 1402 -1115 0 3
rlabel polysilicon 1409 -1109 1409 -1109 0 1
rlabel polysilicon 1409 -1115 1409 -1115 0 3
rlabel polysilicon 1416 -1109 1416 -1109 0 1
rlabel polysilicon 1416 -1115 1416 -1115 0 3
rlabel polysilicon 1423 -1109 1423 -1109 0 1
rlabel polysilicon 1423 -1115 1423 -1115 0 3
rlabel polysilicon 1430 -1109 1430 -1109 0 1
rlabel polysilicon 1430 -1115 1430 -1115 0 3
rlabel polysilicon 1437 -1109 1437 -1109 0 1
rlabel polysilicon 1437 -1115 1437 -1115 0 3
rlabel polysilicon 1444 -1109 1444 -1109 0 1
rlabel polysilicon 1444 -1115 1444 -1115 0 3
rlabel polysilicon 1451 -1109 1451 -1109 0 1
rlabel polysilicon 1451 -1115 1451 -1115 0 3
rlabel polysilicon 1458 -1109 1458 -1109 0 1
rlabel polysilicon 1458 -1115 1458 -1115 0 3
rlabel polysilicon 1465 -1109 1465 -1109 0 1
rlabel polysilicon 1465 -1115 1465 -1115 0 3
rlabel polysilicon 1472 -1109 1472 -1109 0 1
rlabel polysilicon 1472 -1115 1472 -1115 0 3
rlabel polysilicon 1479 -1109 1479 -1109 0 1
rlabel polysilicon 1479 -1115 1479 -1115 0 3
rlabel polysilicon 1486 -1109 1486 -1109 0 1
rlabel polysilicon 1486 -1115 1486 -1115 0 3
rlabel polysilicon 1493 -1109 1493 -1109 0 1
rlabel polysilicon 1493 -1115 1493 -1115 0 3
rlabel polysilicon 1500 -1109 1500 -1109 0 1
rlabel polysilicon 1500 -1115 1500 -1115 0 3
rlabel polysilicon 1507 -1109 1507 -1109 0 1
rlabel polysilicon 1507 -1115 1507 -1115 0 3
rlabel polysilicon 1514 -1109 1514 -1109 0 1
rlabel polysilicon 1514 -1115 1514 -1115 0 3
rlabel polysilicon 1521 -1109 1521 -1109 0 1
rlabel polysilicon 1521 -1115 1521 -1115 0 3
rlabel polysilicon 1528 -1109 1528 -1109 0 1
rlabel polysilicon 1528 -1115 1528 -1115 0 3
rlabel polysilicon 1535 -1109 1535 -1109 0 1
rlabel polysilicon 1535 -1115 1535 -1115 0 3
rlabel polysilicon 1542 -1109 1542 -1109 0 1
rlabel polysilicon 1542 -1115 1542 -1115 0 3
rlabel polysilicon 1549 -1109 1549 -1109 0 1
rlabel polysilicon 1549 -1115 1549 -1115 0 3
rlabel polysilicon 1556 -1109 1556 -1109 0 1
rlabel polysilicon 1556 -1115 1556 -1115 0 3
rlabel polysilicon 1563 -1109 1563 -1109 0 1
rlabel polysilicon 1563 -1115 1563 -1115 0 3
rlabel polysilicon 1570 -1109 1570 -1109 0 1
rlabel polysilicon 1570 -1115 1570 -1115 0 3
rlabel polysilicon 1577 -1109 1577 -1109 0 1
rlabel polysilicon 1577 -1115 1577 -1115 0 3
rlabel polysilicon 1584 -1109 1584 -1109 0 1
rlabel polysilicon 1584 -1115 1584 -1115 0 3
rlabel polysilicon 1591 -1109 1591 -1109 0 1
rlabel polysilicon 1591 -1115 1591 -1115 0 3
rlabel polysilicon 1598 -1109 1598 -1109 0 1
rlabel polysilicon 1598 -1115 1598 -1115 0 3
rlabel polysilicon 1605 -1109 1605 -1109 0 1
rlabel polysilicon 1605 -1115 1605 -1115 0 3
rlabel polysilicon 1612 -1109 1612 -1109 0 1
rlabel polysilicon 1612 -1115 1612 -1115 0 3
rlabel polysilicon 1619 -1109 1619 -1109 0 1
rlabel polysilicon 1619 -1115 1619 -1115 0 3
rlabel polysilicon 1626 -1109 1626 -1109 0 1
rlabel polysilicon 1626 -1115 1626 -1115 0 3
rlabel polysilicon 1633 -1109 1633 -1109 0 1
rlabel polysilicon 1633 -1115 1633 -1115 0 3
rlabel polysilicon 1640 -1109 1640 -1109 0 1
rlabel polysilicon 1640 -1115 1640 -1115 0 3
rlabel polysilicon 1647 -1109 1647 -1109 0 1
rlabel polysilicon 1647 -1115 1647 -1115 0 3
rlabel polysilicon 1654 -1109 1654 -1109 0 1
rlabel polysilicon 1654 -1115 1654 -1115 0 3
rlabel polysilicon 1661 -1109 1661 -1109 0 1
rlabel polysilicon 1661 -1115 1661 -1115 0 3
rlabel polysilicon 1668 -1109 1668 -1109 0 1
rlabel polysilicon 1668 -1115 1668 -1115 0 3
rlabel polysilicon 1675 -1109 1675 -1109 0 1
rlabel polysilicon 1675 -1115 1675 -1115 0 3
rlabel polysilicon 1682 -1109 1682 -1109 0 1
rlabel polysilicon 1682 -1115 1682 -1115 0 3
rlabel polysilicon 1689 -1109 1689 -1109 0 1
rlabel polysilicon 1689 -1115 1689 -1115 0 3
rlabel polysilicon 1696 -1109 1696 -1109 0 1
rlabel polysilicon 1696 -1115 1696 -1115 0 3
rlabel polysilicon 1703 -1109 1703 -1109 0 1
rlabel polysilicon 1703 -1115 1703 -1115 0 3
rlabel polysilicon 1710 -1109 1710 -1109 0 1
rlabel polysilicon 1710 -1115 1710 -1115 0 3
rlabel polysilicon 1717 -1109 1717 -1109 0 1
rlabel polysilicon 1717 -1115 1717 -1115 0 3
rlabel polysilicon 1724 -1109 1724 -1109 0 1
rlabel polysilicon 1724 -1115 1724 -1115 0 3
rlabel polysilicon 1731 -1109 1731 -1109 0 1
rlabel polysilicon 1731 -1115 1731 -1115 0 3
rlabel polysilicon 1738 -1109 1738 -1109 0 1
rlabel polysilicon 1738 -1115 1738 -1115 0 3
rlabel polysilicon 1745 -1109 1745 -1109 0 1
rlabel polysilicon 1745 -1115 1745 -1115 0 3
rlabel polysilicon 1752 -1109 1752 -1109 0 1
rlabel polysilicon 1752 -1115 1752 -1115 0 3
rlabel polysilicon 1759 -1109 1759 -1109 0 1
rlabel polysilicon 1759 -1115 1759 -1115 0 3
rlabel polysilicon 1766 -1109 1766 -1109 0 1
rlabel polysilicon 1766 -1115 1766 -1115 0 3
rlabel polysilicon 1773 -1109 1773 -1109 0 1
rlabel polysilicon 1773 -1115 1773 -1115 0 3
rlabel polysilicon 1780 -1109 1780 -1109 0 1
rlabel polysilicon 1780 -1115 1780 -1115 0 3
rlabel polysilicon 1787 -1109 1787 -1109 0 1
rlabel polysilicon 1787 -1115 1787 -1115 0 3
rlabel polysilicon 1794 -1109 1794 -1109 0 1
rlabel polysilicon 1794 -1115 1794 -1115 0 3
rlabel polysilicon 1801 -1109 1801 -1109 0 1
rlabel polysilicon 1801 -1115 1801 -1115 0 3
rlabel polysilicon 1808 -1109 1808 -1109 0 1
rlabel polysilicon 1808 -1115 1808 -1115 0 3
rlabel polysilicon 1815 -1109 1815 -1109 0 1
rlabel polysilicon 1815 -1115 1815 -1115 0 3
rlabel polysilicon 1822 -1109 1822 -1109 0 1
rlabel polysilicon 1822 -1115 1822 -1115 0 3
rlabel polysilicon 1829 -1109 1829 -1109 0 1
rlabel polysilicon 1829 -1115 1829 -1115 0 3
rlabel polysilicon 1836 -1109 1836 -1109 0 1
rlabel polysilicon 1836 -1115 1836 -1115 0 3
rlabel polysilicon 1843 -1109 1843 -1109 0 1
rlabel polysilicon 1843 -1115 1843 -1115 0 3
rlabel polysilicon 1850 -1109 1850 -1109 0 1
rlabel polysilicon 1850 -1115 1850 -1115 0 3
rlabel polysilicon 1857 -1109 1857 -1109 0 1
rlabel polysilicon 1857 -1115 1857 -1115 0 3
rlabel polysilicon 1867 -1109 1867 -1109 0 2
rlabel polysilicon 1864 -1115 1864 -1115 0 3
rlabel polysilicon 1867 -1115 1867 -1115 0 4
rlabel polysilicon 1871 -1109 1871 -1109 0 1
rlabel polysilicon 1871 -1115 1871 -1115 0 3
rlabel polysilicon 1878 -1109 1878 -1109 0 1
rlabel polysilicon 1878 -1115 1878 -1115 0 3
rlabel polysilicon 1927 -1109 1927 -1109 0 1
rlabel polysilicon 1927 -1115 1927 -1115 0 3
rlabel polysilicon 1948 -1109 1948 -1109 0 1
rlabel polysilicon 1948 -1115 1948 -1115 0 3
rlabel polysilicon 1962 -1109 1962 -1109 0 1
rlabel polysilicon 1962 -1115 1962 -1115 0 3
rlabel polysilicon 1969 -1109 1969 -1109 0 1
rlabel polysilicon 1969 -1115 1969 -1115 0 3
rlabel polysilicon 1976 -1109 1976 -1109 0 1
rlabel polysilicon 1976 -1115 1976 -1115 0 3
rlabel polysilicon 2 -1244 2 -1244 0 1
rlabel polysilicon 2 -1250 2 -1250 0 3
rlabel polysilicon 9 -1244 9 -1244 0 1
rlabel polysilicon 9 -1250 9 -1250 0 3
rlabel polysilicon 16 -1244 16 -1244 0 1
rlabel polysilicon 16 -1250 16 -1250 0 3
rlabel polysilicon 30 -1244 30 -1244 0 1
rlabel polysilicon 30 -1250 30 -1250 0 3
rlabel polysilicon 37 -1244 37 -1244 0 1
rlabel polysilicon 40 -1244 40 -1244 0 2
rlabel polysilicon 40 -1250 40 -1250 0 4
rlabel polysilicon 44 -1244 44 -1244 0 1
rlabel polysilicon 44 -1250 44 -1250 0 3
rlabel polysilicon 51 -1244 51 -1244 0 1
rlabel polysilicon 51 -1250 51 -1250 0 3
rlabel polysilicon 58 -1244 58 -1244 0 1
rlabel polysilicon 61 -1244 61 -1244 0 2
rlabel polysilicon 58 -1250 58 -1250 0 3
rlabel polysilicon 61 -1250 61 -1250 0 4
rlabel polysilicon 65 -1244 65 -1244 0 1
rlabel polysilicon 65 -1250 65 -1250 0 3
rlabel polysilicon 72 -1244 72 -1244 0 1
rlabel polysilicon 72 -1250 72 -1250 0 3
rlabel polysilicon 79 -1244 79 -1244 0 1
rlabel polysilicon 82 -1244 82 -1244 0 2
rlabel polysilicon 79 -1250 79 -1250 0 3
rlabel polysilicon 82 -1250 82 -1250 0 4
rlabel polysilicon 86 -1244 86 -1244 0 1
rlabel polysilicon 86 -1250 86 -1250 0 3
rlabel polysilicon 93 -1244 93 -1244 0 1
rlabel polysilicon 93 -1250 93 -1250 0 3
rlabel polysilicon 100 -1244 100 -1244 0 1
rlabel polysilicon 100 -1250 100 -1250 0 3
rlabel polysilicon 107 -1244 107 -1244 0 1
rlabel polysilicon 107 -1250 107 -1250 0 3
rlabel polysilicon 114 -1244 114 -1244 0 1
rlabel polysilicon 114 -1250 114 -1250 0 3
rlabel polysilicon 121 -1244 121 -1244 0 1
rlabel polysilicon 124 -1244 124 -1244 0 2
rlabel polysilicon 124 -1250 124 -1250 0 4
rlabel polysilicon 128 -1244 128 -1244 0 1
rlabel polysilicon 128 -1250 128 -1250 0 3
rlabel polysilicon 135 -1244 135 -1244 0 1
rlabel polysilicon 135 -1250 135 -1250 0 3
rlabel polysilicon 142 -1244 142 -1244 0 1
rlabel polysilicon 142 -1250 142 -1250 0 3
rlabel polysilicon 149 -1244 149 -1244 0 1
rlabel polysilicon 149 -1250 149 -1250 0 3
rlabel polysilicon 159 -1244 159 -1244 0 2
rlabel polysilicon 156 -1250 156 -1250 0 3
rlabel polysilicon 159 -1250 159 -1250 0 4
rlabel polysilicon 163 -1244 163 -1244 0 1
rlabel polysilicon 163 -1250 163 -1250 0 3
rlabel polysilicon 170 -1244 170 -1244 0 1
rlabel polysilicon 170 -1250 170 -1250 0 3
rlabel polysilicon 173 -1250 173 -1250 0 4
rlabel polysilicon 177 -1244 177 -1244 0 1
rlabel polysilicon 180 -1244 180 -1244 0 2
rlabel polysilicon 177 -1250 177 -1250 0 3
rlabel polysilicon 180 -1250 180 -1250 0 4
rlabel polysilicon 184 -1244 184 -1244 0 1
rlabel polysilicon 184 -1250 184 -1250 0 3
rlabel polysilicon 191 -1244 191 -1244 0 1
rlabel polysilicon 191 -1250 191 -1250 0 3
rlabel polysilicon 198 -1244 198 -1244 0 1
rlabel polysilicon 198 -1250 198 -1250 0 3
rlabel polysilicon 205 -1244 205 -1244 0 1
rlabel polysilicon 205 -1250 205 -1250 0 3
rlabel polysilicon 212 -1244 212 -1244 0 1
rlabel polysilicon 212 -1250 212 -1250 0 3
rlabel polysilicon 219 -1244 219 -1244 0 1
rlabel polysilicon 219 -1250 219 -1250 0 3
rlabel polysilicon 229 -1244 229 -1244 0 2
rlabel polysilicon 226 -1250 226 -1250 0 3
rlabel polysilicon 229 -1250 229 -1250 0 4
rlabel polysilicon 233 -1244 233 -1244 0 1
rlabel polysilicon 233 -1250 233 -1250 0 3
rlabel polysilicon 240 -1244 240 -1244 0 1
rlabel polysilicon 240 -1250 240 -1250 0 3
rlabel polysilicon 247 -1244 247 -1244 0 1
rlabel polysilicon 247 -1250 247 -1250 0 3
rlabel polysilicon 254 -1244 254 -1244 0 1
rlabel polysilicon 254 -1250 254 -1250 0 3
rlabel polysilicon 261 -1250 261 -1250 0 3
rlabel polysilicon 264 -1250 264 -1250 0 4
rlabel polysilicon 268 -1244 268 -1244 0 1
rlabel polysilicon 268 -1250 268 -1250 0 3
rlabel polysilicon 275 -1244 275 -1244 0 1
rlabel polysilicon 275 -1250 275 -1250 0 3
rlabel polysilicon 282 -1244 282 -1244 0 1
rlabel polysilicon 282 -1250 282 -1250 0 3
rlabel polysilicon 289 -1244 289 -1244 0 1
rlabel polysilicon 292 -1244 292 -1244 0 2
rlabel polysilicon 296 -1244 296 -1244 0 1
rlabel polysilicon 296 -1250 296 -1250 0 3
rlabel polysilicon 303 -1244 303 -1244 0 1
rlabel polysilicon 303 -1250 303 -1250 0 3
rlabel polysilicon 310 -1244 310 -1244 0 1
rlabel polysilicon 310 -1250 310 -1250 0 3
rlabel polysilicon 317 -1244 317 -1244 0 1
rlabel polysilicon 317 -1250 317 -1250 0 3
rlabel polysilicon 324 -1244 324 -1244 0 1
rlabel polysilicon 324 -1250 324 -1250 0 3
rlabel polysilicon 331 -1244 331 -1244 0 1
rlabel polysilicon 338 -1244 338 -1244 0 1
rlabel polysilicon 338 -1250 338 -1250 0 3
rlabel polysilicon 345 -1244 345 -1244 0 1
rlabel polysilicon 345 -1250 345 -1250 0 3
rlabel polysilicon 352 -1244 352 -1244 0 1
rlabel polysilicon 352 -1250 352 -1250 0 3
rlabel polysilicon 359 -1244 359 -1244 0 1
rlabel polysilicon 359 -1250 359 -1250 0 3
rlabel polysilicon 366 -1244 366 -1244 0 1
rlabel polysilicon 366 -1250 366 -1250 0 3
rlabel polysilicon 373 -1244 373 -1244 0 1
rlabel polysilicon 373 -1250 373 -1250 0 3
rlabel polysilicon 380 -1244 380 -1244 0 1
rlabel polysilicon 380 -1250 380 -1250 0 3
rlabel polysilicon 387 -1250 387 -1250 0 3
rlabel polysilicon 394 -1244 394 -1244 0 1
rlabel polysilicon 394 -1250 394 -1250 0 3
rlabel polysilicon 401 -1244 401 -1244 0 1
rlabel polysilicon 401 -1250 401 -1250 0 3
rlabel polysilicon 408 -1244 408 -1244 0 1
rlabel polysilicon 408 -1250 408 -1250 0 3
rlabel polysilicon 415 -1244 415 -1244 0 1
rlabel polysilicon 415 -1250 415 -1250 0 3
rlabel polysilicon 422 -1244 422 -1244 0 1
rlabel polysilicon 425 -1244 425 -1244 0 2
rlabel polysilicon 422 -1250 422 -1250 0 3
rlabel polysilicon 425 -1250 425 -1250 0 4
rlabel polysilicon 429 -1244 429 -1244 0 1
rlabel polysilicon 429 -1250 429 -1250 0 3
rlabel polysilicon 436 -1244 436 -1244 0 1
rlabel polysilicon 436 -1250 436 -1250 0 3
rlabel polysilicon 443 -1244 443 -1244 0 1
rlabel polysilicon 446 -1244 446 -1244 0 2
rlabel polysilicon 443 -1250 443 -1250 0 3
rlabel polysilicon 446 -1250 446 -1250 0 4
rlabel polysilicon 450 -1244 450 -1244 0 1
rlabel polysilicon 453 -1244 453 -1244 0 2
rlabel polysilicon 450 -1250 450 -1250 0 3
rlabel polysilicon 453 -1250 453 -1250 0 4
rlabel polysilicon 457 -1244 457 -1244 0 1
rlabel polysilicon 457 -1250 457 -1250 0 3
rlabel polysilicon 464 -1244 464 -1244 0 1
rlabel polysilicon 464 -1250 464 -1250 0 3
rlabel polysilicon 471 -1244 471 -1244 0 1
rlabel polysilicon 474 -1244 474 -1244 0 2
rlabel polysilicon 474 -1250 474 -1250 0 4
rlabel polysilicon 478 -1244 478 -1244 0 1
rlabel polysilicon 478 -1250 478 -1250 0 3
rlabel polysilicon 485 -1244 485 -1244 0 1
rlabel polysilicon 485 -1250 485 -1250 0 3
rlabel polysilicon 492 -1244 492 -1244 0 1
rlabel polysilicon 492 -1250 492 -1250 0 3
rlabel polysilicon 499 -1244 499 -1244 0 1
rlabel polysilicon 499 -1250 499 -1250 0 3
rlabel polysilicon 506 -1244 506 -1244 0 1
rlabel polysilicon 506 -1250 506 -1250 0 3
rlabel polysilicon 516 -1244 516 -1244 0 2
rlabel polysilicon 513 -1250 513 -1250 0 3
rlabel polysilicon 516 -1250 516 -1250 0 4
rlabel polysilicon 520 -1244 520 -1244 0 1
rlabel polysilicon 520 -1250 520 -1250 0 3
rlabel polysilicon 527 -1244 527 -1244 0 1
rlabel polysilicon 527 -1250 527 -1250 0 3
rlabel polysilicon 534 -1244 534 -1244 0 1
rlabel polysilicon 534 -1250 534 -1250 0 3
rlabel polysilicon 541 -1244 541 -1244 0 1
rlabel polysilicon 541 -1250 541 -1250 0 3
rlabel polysilicon 548 -1244 548 -1244 0 1
rlabel polysilicon 548 -1250 548 -1250 0 3
rlabel polysilicon 555 -1244 555 -1244 0 1
rlabel polysilicon 555 -1250 555 -1250 0 3
rlabel polysilicon 562 -1244 562 -1244 0 1
rlabel polysilicon 562 -1250 562 -1250 0 3
rlabel polysilicon 565 -1250 565 -1250 0 4
rlabel polysilicon 569 -1244 569 -1244 0 1
rlabel polysilicon 569 -1250 569 -1250 0 3
rlabel polysilicon 576 -1244 576 -1244 0 1
rlabel polysilicon 576 -1250 576 -1250 0 3
rlabel polysilicon 583 -1244 583 -1244 0 1
rlabel polysilicon 586 -1244 586 -1244 0 2
rlabel polysilicon 583 -1250 583 -1250 0 3
rlabel polysilicon 586 -1250 586 -1250 0 4
rlabel polysilicon 590 -1244 590 -1244 0 1
rlabel polysilicon 590 -1250 590 -1250 0 3
rlabel polysilicon 597 -1244 597 -1244 0 1
rlabel polysilicon 597 -1250 597 -1250 0 3
rlabel polysilicon 604 -1244 604 -1244 0 1
rlabel polysilicon 604 -1250 604 -1250 0 3
rlabel polysilicon 611 -1244 611 -1244 0 1
rlabel polysilicon 611 -1250 611 -1250 0 3
rlabel polysilicon 618 -1244 618 -1244 0 1
rlabel polysilicon 618 -1250 618 -1250 0 3
rlabel polysilicon 625 -1244 625 -1244 0 1
rlabel polysilicon 625 -1250 625 -1250 0 3
rlabel polysilicon 632 -1244 632 -1244 0 1
rlabel polysilicon 632 -1250 632 -1250 0 3
rlabel polysilicon 639 -1244 639 -1244 0 1
rlabel polysilicon 639 -1250 639 -1250 0 3
rlabel polysilicon 646 -1244 646 -1244 0 1
rlabel polysilicon 646 -1250 646 -1250 0 3
rlabel polysilicon 653 -1244 653 -1244 0 1
rlabel polysilicon 653 -1250 653 -1250 0 3
rlabel polysilicon 660 -1244 660 -1244 0 1
rlabel polysilicon 660 -1250 660 -1250 0 3
rlabel polysilicon 667 -1244 667 -1244 0 1
rlabel polysilicon 670 -1244 670 -1244 0 2
rlabel polysilicon 667 -1250 667 -1250 0 3
rlabel polysilicon 670 -1250 670 -1250 0 4
rlabel polysilicon 674 -1244 674 -1244 0 1
rlabel polysilicon 674 -1250 674 -1250 0 3
rlabel polysilicon 681 -1244 681 -1244 0 1
rlabel polysilicon 681 -1250 681 -1250 0 3
rlabel polysilicon 688 -1244 688 -1244 0 1
rlabel polysilicon 688 -1250 688 -1250 0 3
rlabel polysilicon 695 -1244 695 -1244 0 1
rlabel polysilicon 695 -1250 695 -1250 0 3
rlabel polysilicon 702 -1244 702 -1244 0 1
rlabel polysilicon 702 -1250 702 -1250 0 3
rlabel polysilicon 709 -1244 709 -1244 0 1
rlabel polysilicon 709 -1250 709 -1250 0 3
rlabel polysilicon 716 -1244 716 -1244 0 1
rlabel polysilicon 716 -1250 716 -1250 0 3
rlabel polysilicon 723 -1244 723 -1244 0 1
rlabel polysilicon 723 -1250 723 -1250 0 3
rlabel polysilicon 730 -1244 730 -1244 0 1
rlabel polysilicon 730 -1250 730 -1250 0 3
rlabel polysilicon 737 -1244 737 -1244 0 1
rlabel polysilicon 737 -1250 737 -1250 0 3
rlabel polysilicon 744 -1244 744 -1244 0 1
rlabel polysilicon 747 -1244 747 -1244 0 2
rlabel polysilicon 744 -1250 744 -1250 0 3
rlabel polysilicon 751 -1244 751 -1244 0 1
rlabel polysilicon 751 -1250 751 -1250 0 3
rlabel polysilicon 758 -1244 758 -1244 0 1
rlabel polysilicon 758 -1250 758 -1250 0 3
rlabel polysilicon 765 -1244 765 -1244 0 1
rlabel polysilicon 765 -1250 765 -1250 0 3
rlabel polysilicon 772 -1244 772 -1244 0 1
rlabel polysilicon 775 -1244 775 -1244 0 2
rlabel polysilicon 772 -1250 772 -1250 0 3
rlabel polysilicon 775 -1250 775 -1250 0 4
rlabel polysilicon 779 -1244 779 -1244 0 1
rlabel polysilicon 782 -1244 782 -1244 0 2
rlabel polysilicon 779 -1250 779 -1250 0 3
rlabel polysilicon 786 -1244 786 -1244 0 1
rlabel polysilicon 786 -1250 786 -1250 0 3
rlabel polysilicon 793 -1244 793 -1244 0 1
rlabel polysilicon 793 -1250 793 -1250 0 3
rlabel polysilicon 800 -1244 800 -1244 0 1
rlabel polysilicon 800 -1250 800 -1250 0 3
rlabel polysilicon 807 -1244 807 -1244 0 1
rlabel polysilicon 810 -1244 810 -1244 0 2
rlabel polysilicon 807 -1250 807 -1250 0 3
rlabel polysilicon 810 -1250 810 -1250 0 4
rlabel polysilicon 814 -1244 814 -1244 0 1
rlabel polysilicon 814 -1250 814 -1250 0 3
rlabel polysilicon 821 -1244 821 -1244 0 1
rlabel polysilicon 821 -1250 821 -1250 0 3
rlabel polysilicon 824 -1250 824 -1250 0 4
rlabel polysilicon 828 -1244 828 -1244 0 1
rlabel polysilicon 828 -1250 828 -1250 0 3
rlabel polysilicon 835 -1244 835 -1244 0 1
rlabel polysilicon 835 -1250 835 -1250 0 3
rlabel polysilicon 842 -1244 842 -1244 0 1
rlabel polysilicon 842 -1250 842 -1250 0 3
rlabel polysilicon 849 -1244 849 -1244 0 1
rlabel polysilicon 849 -1250 849 -1250 0 3
rlabel polysilicon 856 -1244 856 -1244 0 1
rlabel polysilicon 859 -1244 859 -1244 0 2
rlabel polysilicon 856 -1250 856 -1250 0 3
rlabel polysilicon 859 -1250 859 -1250 0 4
rlabel polysilicon 863 -1244 863 -1244 0 1
rlabel polysilicon 863 -1250 863 -1250 0 3
rlabel polysilicon 870 -1244 870 -1244 0 1
rlabel polysilicon 873 -1244 873 -1244 0 2
rlabel polysilicon 873 -1250 873 -1250 0 4
rlabel polysilicon 877 -1244 877 -1244 0 1
rlabel polysilicon 880 -1244 880 -1244 0 2
rlabel polysilicon 877 -1250 877 -1250 0 3
rlabel polysilicon 884 -1244 884 -1244 0 1
rlabel polysilicon 884 -1250 884 -1250 0 3
rlabel polysilicon 891 -1244 891 -1244 0 1
rlabel polysilicon 891 -1250 891 -1250 0 3
rlabel polysilicon 898 -1244 898 -1244 0 1
rlabel polysilicon 898 -1250 898 -1250 0 3
rlabel polysilicon 905 -1244 905 -1244 0 1
rlabel polysilicon 908 -1244 908 -1244 0 2
rlabel polysilicon 905 -1250 905 -1250 0 3
rlabel polysilicon 908 -1250 908 -1250 0 4
rlabel polysilicon 912 -1244 912 -1244 0 1
rlabel polysilicon 912 -1250 912 -1250 0 3
rlabel polysilicon 919 -1244 919 -1244 0 1
rlabel polysilicon 919 -1250 919 -1250 0 3
rlabel polysilicon 926 -1244 926 -1244 0 1
rlabel polysilicon 929 -1244 929 -1244 0 2
rlabel polysilicon 926 -1250 926 -1250 0 3
rlabel polysilicon 929 -1250 929 -1250 0 4
rlabel polysilicon 933 -1244 933 -1244 0 1
rlabel polysilicon 933 -1250 933 -1250 0 3
rlabel polysilicon 940 -1244 940 -1244 0 1
rlabel polysilicon 940 -1250 940 -1250 0 3
rlabel polysilicon 947 -1244 947 -1244 0 1
rlabel polysilicon 947 -1250 947 -1250 0 3
rlabel polysilicon 954 -1244 954 -1244 0 1
rlabel polysilicon 954 -1250 954 -1250 0 3
rlabel polysilicon 964 -1244 964 -1244 0 2
rlabel polysilicon 961 -1250 961 -1250 0 3
rlabel polysilicon 964 -1250 964 -1250 0 4
rlabel polysilicon 968 -1244 968 -1244 0 1
rlabel polysilicon 968 -1250 968 -1250 0 3
rlabel polysilicon 975 -1244 975 -1244 0 1
rlabel polysilicon 975 -1250 975 -1250 0 3
rlabel polysilicon 982 -1244 982 -1244 0 1
rlabel polysilicon 982 -1250 982 -1250 0 3
rlabel polysilicon 989 -1244 989 -1244 0 1
rlabel polysilicon 989 -1250 989 -1250 0 3
rlabel polysilicon 996 -1244 996 -1244 0 1
rlabel polysilicon 996 -1250 996 -1250 0 3
rlabel polysilicon 1003 -1244 1003 -1244 0 1
rlabel polysilicon 1003 -1250 1003 -1250 0 3
rlabel polysilicon 1010 -1244 1010 -1244 0 1
rlabel polysilicon 1010 -1250 1010 -1250 0 3
rlabel polysilicon 1017 -1244 1017 -1244 0 1
rlabel polysilicon 1017 -1250 1017 -1250 0 3
rlabel polysilicon 1020 -1250 1020 -1250 0 4
rlabel polysilicon 1024 -1244 1024 -1244 0 1
rlabel polysilicon 1024 -1250 1024 -1250 0 3
rlabel polysilicon 1031 -1244 1031 -1244 0 1
rlabel polysilicon 1031 -1250 1031 -1250 0 3
rlabel polysilicon 1038 -1244 1038 -1244 0 1
rlabel polysilicon 1038 -1250 1038 -1250 0 3
rlabel polysilicon 1045 -1244 1045 -1244 0 1
rlabel polysilicon 1048 -1244 1048 -1244 0 2
rlabel polysilicon 1052 -1244 1052 -1244 0 1
rlabel polysilicon 1052 -1250 1052 -1250 0 3
rlabel polysilicon 1059 -1244 1059 -1244 0 1
rlabel polysilicon 1059 -1250 1059 -1250 0 3
rlabel polysilicon 1066 -1244 1066 -1244 0 1
rlabel polysilicon 1066 -1250 1066 -1250 0 3
rlabel polysilicon 1073 -1244 1073 -1244 0 1
rlabel polysilicon 1073 -1250 1073 -1250 0 3
rlabel polysilicon 1080 -1244 1080 -1244 0 1
rlabel polysilicon 1080 -1250 1080 -1250 0 3
rlabel polysilicon 1087 -1244 1087 -1244 0 1
rlabel polysilicon 1087 -1250 1087 -1250 0 3
rlabel polysilicon 1094 -1244 1094 -1244 0 1
rlabel polysilicon 1094 -1250 1094 -1250 0 3
rlabel polysilicon 1101 -1244 1101 -1244 0 1
rlabel polysilicon 1101 -1250 1101 -1250 0 3
rlabel polysilicon 1108 -1244 1108 -1244 0 1
rlabel polysilicon 1108 -1250 1108 -1250 0 3
rlabel polysilicon 1115 -1244 1115 -1244 0 1
rlabel polysilicon 1115 -1250 1115 -1250 0 3
rlabel polysilicon 1122 -1244 1122 -1244 0 1
rlabel polysilicon 1122 -1250 1122 -1250 0 3
rlabel polysilicon 1129 -1244 1129 -1244 0 1
rlabel polysilicon 1132 -1244 1132 -1244 0 2
rlabel polysilicon 1129 -1250 1129 -1250 0 3
rlabel polysilicon 1132 -1250 1132 -1250 0 4
rlabel polysilicon 1136 -1244 1136 -1244 0 1
rlabel polysilicon 1136 -1250 1136 -1250 0 3
rlabel polysilicon 1143 -1244 1143 -1244 0 1
rlabel polysilicon 1143 -1250 1143 -1250 0 3
rlabel polysilicon 1150 -1244 1150 -1244 0 1
rlabel polysilicon 1150 -1250 1150 -1250 0 3
rlabel polysilicon 1157 -1244 1157 -1244 0 1
rlabel polysilicon 1160 -1244 1160 -1244 0 2
rlabel polysilicon 1164 -1244 1164 -1244 0 1
rlabel polysilicon 1164 -1250 1164 -1250 0 3
rlabel polysilicon 1171 -1244 1171 -1244 0 1
rlabel polysilicon 1171 -1250 1171 -1250 0 3
rlabel polysilicon 1178 -1244 1178 -1244 0 1
rlabel polysilicon 1181 -1244 1181 -1244 0 2
rlabel polysilicon 1178 -1250 1178 -1250 0 3
rlabel polysilicon 1181 -1250 1181 -1250 0 4
rlabel polysilicon 1185 -1244 1185 -1244 0 1
rlabel polysilicon 1185 -1250 1185 -1250 0 3
rlabel polysilicon 1192 -1244 1192 -1244 0 1
rlabel polysilicon 1192 -1250 1192 -1250 0 3
rlabel polysilicon 1199 -1244 1199 -1244 0 1
rlabel polysilicon 1199 -1250 1199 -1250 0 3
rlabel polysilicon 1206 -1244 1206 -1244 0 1
rlabel polysilicon 1206 -1250 1206 -1250 0 3
rlabel polysilicon 1213 -1244 1213 -1244 0 1
rlabel polysilicon 1213 -1250 1213 -1250 0 3
rlabel polysilicon 1220 -1244 1220 -1244 0 1
rlabel polysilicon 1220 -1250 1220 -1250 0 3
rlabel polysilicon 1227 -1244 1227 -1244 0 1
rlabel polysilicon 1227 -1250 1227 -1250 0 3
rlabel polysilicon 1234 -1244 1234 -1244 0 1
rlabel polysilicon 1234 -1250 1234 -1250 0 3
rlabel polysilicon 1241 -1244 1241 -1244 0 1
rlabel polysilicon 1241 -1250 1241 -1250 0 3
rlabel polysilicon 1248 -1244 1248 -1244 0 1
rlabel polysilicon 1248 -1250 1248 -1250 0 3
rlabel polysilicon 1255 -1244 1255 -1244 0 1
rlabel polysilicon 1255 -1250 1255 -1250 0 3
rlabel polysilicon 1262 -1244 1262 -1244 0 1
rlabel polysilicon 1262 -1250 1262 -1250 0 3
rlabel polysilicon 1269 -1244 1269 -1244 0 1
rlabel polysilicon 1269 -1250 1269 -1250 0 3
rlabel polysilicon 1276 -1244 1276 -1244 0 1
rlabel polysilicon 1276 -1250 1276 -1250 0 3
rlabel polysilicon 1283 -1244 1283 -1244 0 1
rlabel polysilicon 1283 -1250 1283 -1250 0 3
rlabel polysilicon 1290 -1244 1290 -1244 0 1
rlabel polysilicon 1290 -1250 1290 -1250 0 3
rlabel polysilicon 1297 -1244 1297 -1244 0 1
rlabel polysilicon 1297 -1250 1297 -1250 0 3
rlabel polysilicon 1304 -1244 1304 -1244 0 1
rlabel polysilicon 1304 -1250 1304 -1250 0 3
rlabel polysilicon 1311 -1244 1311 -1244 0 1
rlabel polysilicon 1311 -1250 1311 -1250 0 3
rlabel polysilicon 1318 -1244 1318 -1244 0 1
rlabel polysilicon 1318 -1250 1318 -1250 0 3
rlabel polysilicon 1325 -1244 1325 -1244 0 1
rlabel polysilicon 1325 -1250 1325 -1250 0 3
rlabel polysilicon 1332 -1244 1332 -1244 0 1
rlabel polysilicon 1332 -1250 1332 -1250 0 3
rlabel polysilicon 1339 -1244 1339 -1244 0 1
rlabel polysilicon 1339 -1250 1339 -1250 0 3
rlabel polysilicon 1346 -1244 1346 -1244 0 1
rlabel polysilicon 1346 -1250 1346 -1250 0 3
rlabel polysilicon 1353 -1244 1353 -1244 0 1
rlabel polysilicon 1353 -1250 1353 -1250 0 3
rlabel polysilicon 1360 -1244 1360 -1244 0 1
rlabel polysilicon 1360 -1250 1360 -1250 0 3
rlabel polysilicon 1367 -1244 1367 -1244 0 1
rlabel polysilicon 1367 -1250 1367 -1250 0 3
rlabel polysilicon 1374 -1244 1374 -1244 0 1
rlabel polysilicon 1374 -1250 1374 -1250 0 3
rlabel polysilicon 1381 -1244 1381 -1244 0 1
rlabel polysilicon 1381 -1250 1381 -1250 0 3
rlabel polysilicon 1388 -1244 1388 -1244 0 1
rlabel polysilicon 1388 -1250 1388 -1250 0 3
rlabel polysilicon 1391 -1250 1391 -1250 0 4
rlabel polysilicon 1395 -1244 1395 -1244 0 1
rlabel polysilicon 1395 -1250 1395 -1250 0 3
rlabel polysilicon 1402 -1244 1402 -1244 0 1
rlabel polysilicon 1402 -1250 1402 -1250 0 3
rlabel polysilicon 1409 -1244 1409 -1244 0 1
rlabel polysilicon 1409 -1250 1409 -1250 0 3
rlabel polysilicon 1416 -1244 1416 -1244 0 1
rlabel polysilicon 1416 -1250 1416 -1250 0 3
rlabel polysilicon 1423 -1244 1423 -1244 0 1
rlabel polysilicon 1423 -1250 1423 -1250 0 3
rlabel polysilicon 1430 -1244 1430 -1244 0 1
rlabel polysilicon 1430 -1250 1430 -1250 0 3
rlabel polysilicon 1437 -1244 1437 -1244 0 1
rlabel polysilicon 1437 -1250 1437 -1250 0 3
rlabel polysilicon 1444 -1244 1444 -1244 0 1
rlabel polysilicon 1444 -1250 1444 -1250 0 3
rlabel polysilicon 1451 -1244 1451 -1244 0 1
rlabel polysilicon 1451 -1250 1451 -1250 0 3
rlabel polysilicon 1458 -1244 1458 -1244 0 1
rlabel polysilicon 1458 -1250 1458 -1250 0 3
rlabel polysilicon 1465 -1244 1465 -1244 0 1
rlabel polysilicon 1465 -1250 1465 -1250 0 3
rlabel polysilicon 1472 -1244 1472 -1244 0 1
rlabel polysilicon 1472 -1250 1472 -1250 0 3
rlabel polysilicon 1479 -1244 1479 -1244 0 1
rlabel polysilicon 1479 -1250 1479 -1250 0 3
rlabel polysilicon 1486 -1244 1486 -1244 0 1
rlabel polysilicon 1486 -1250 1486 -1250 0 3
rlabel polysilicon 1493 -1244 1493 -1244 0 1
rlabel polysilicon 1493 -1250 1493 -1250 0 3
rlabel polysilicon 1500 -1244 1500 -1244 0 1
rlabel polysilicon 1500 -1250 1500 -1250 0 3
rlabel polysilicon 1507 -1244 1507 -1244 0 1
rlabel polysilicon 1507 -1250 1507 -1250 0 3
rlabel polysilicon 1514 -1244 1514 -1244 0 1
rlabel polysilicon 1514 -1250 1514 -1250 0 3
rlabel polysilicon 1521 -1244 1521 -1244 0 1
rlabel polysilicon 1521 -1250 1521 -1250 0 3
rlabel polysilicon 1528 -1244 1528 -1244 0 1
rlabel polysilicon 1528 -1250 1528 -1250 0 3
rlabel polysilicon 1535 -1244 1535 -1244 0 1
rlabel polysilicon 1535 -1250 1535 -1250 0 3
rlabel polysilicon 1542 -1244 1542 -1244 0 1
rlabel polysilicon 1542 -1250 1542 -1250 0 3
rlabel polysilicon 1549 -1244 1549 -1244 0 1
rlabel polysilicon 1549 -1250 1549 -1250 0 3
rlabel polysilicon 1556 -1244 1556 -1244 0 1
rlabel polysilicon 1556 -1250 1556 -1250 0 3
rlabel polysilicon 1563 -1244 1563 -1244 0 1
rlabel polysilicon 1563 -1250 1563 -1250 0 3
rlabel polysilicon 1570 -1244 1570 -1244 0 1
rlabel polysilicon 1570 -1250 1570 -1250 0 3
rlabel polysilicon 1577 -1244 1577 -1244 0 1
rlabel polysilicon 1577 -1250 1577 -1250 0 3
rlabel polysilicon 1584 -1244 1584 -1244 0 1
rlabel polysilicon 1584 -1250 1584 -1250 0 3
rlabel polysilicon 1591 -1244 1591 -1244 0 1
rlabel polysilicon 1591 -1250 1591 -1250 0 3
rlabel polysilicon 1598 -1244 1598 -1244 0 1
rlabel polysilicon 1598 -1250 1598 -1250 0 3
rlabel polysilicon 1605 -1244 1605 -1244 0 1
rlabel polysilicon 1605 -1250 1605 -1250 0 3
rlabel polysilicon 1612 -1244 1612 -1244 0 1
rlabel polysilicon 1612 -1250 1612 -1250 0 3
rlabel polysilicon 1619 -1244 1619 -1244 0 1
rlabel polysilicon 1619 -1250 1619 -1250 0 3
rlabel polysilicon 1626 -1244 1626 -1244 0 1
rlabel polysilicon 1626 -1250 1626 -1250 0 3
rlabel polysilicon 1633 -1244 1633 -1244 0 1
rlabel polysilicon 1633 -1250 1633 -1250 0 3
rlabel polysilicon 1640 -1244 1640 -1244 0 1
rlabel polysilicon 1640 -1250 1640 -1250 0 3
rlabel polysilicon 1647 -1244 1647 -1244 0 1
rlabel polysilicon 1647 -1250 1647 -1250 0 3
rlabel polysilicon 1654 -1244 1654 -1244 0 1
rlabel polysilicon 1654 -1250 1654 -1250 0 3
rlabel polysilicon 1661 -1244 1661 -1244 0 1
rlabel polysilicon 1661 -1250 1661 -1250 0 3
rlabel polysilicon 1668 -1244 1668 -1244 0 1
rlabel polysilicon 1668 -1250 1668 -1250 0 3
rlabel polysilicon 1675 -1244 1675 -1244 0 1
rlabel polysilicon 1675 -1250 1675 -1250 0 3
rlabel polysilicon 1682 -1244 1682 -1244 0 1
rlabel polysilicon 1682 -1250 1682 -1250 0 3
rlabel polysilicon 1689 -1244 1689 -1244 0 1
rlabel polysilicon 1689 -1250 1689 -1250 0 3
rlabel polysilicon 1696 -1244 1696 -1244 0 1
rlabel polysilicon 1696 -1250 1696 -1250 0 3
rlabel polysilicon 1703 -1244 1703 -1244 0 1
rlabel polysilicon 1703 -1250 1703 -1250 0 3
rlabel polysilicon 1710 -1244 1710 -1244 0 1
rlabel polysilicon 1710 -1250 1710 -1250 0 3
rlabel polysilicon 1717 -1244 1717 -1244 0 1
rlabel polysilicon 1717 -1250 1717 -1250 0 3
rlabel polysilicon 1724 -1244 1724 -1244 0 1
rlabel polysilicon 1724 -1250 1724 -1250 0 3
rlabel polysilicon 1731 -1244 1731 -1244 0 1
rlabel polysilicon 1731 -1250 1731 -1250 0 3
rlabel polysilicon 1738 -1244 1738 -1244 0 1
rlabel polysilicon 1738 -1250 1738 -1250 0 3
rlabel polysilicon 1745 -1244 1745 -1244 0 1
rlabel polysilicon 1745 -1250 1745 -1250 0 3
rlabel polysilicon 1752 -1244 1752 -1244 0 1
rlabel polysilicon 1752 -1250 1752 -1250 0 3
rlabel polysilicon 1759 -1244 1759 -1244 0 1
rlabel polysilicon 1759 -1250 1759 -1250 0 3
rlabel polysilicon 1766 -1244 1766 -1244 0 1
rlabel polysilicon 1766 -1250 1766 -1250 0 3
rlabel polysilicon 1773 -1244 1773 -1244 0 1
rlabel polysilicon 1773 -1250 1773 -1250 0 3
rlabel polysilicon 1780 -1244 1780 -1244 0 1
rlabel polysilicon 1780 -1250 1780 -1250 0 3
rlabel polysilicon 1787 -1244 1787 -1244 0 1
rlabel polysilicon 1787 -1250 1787 -1250 0 3
rlabel polysilicon 1794 -1244 1794 -1244 0 1
rlabel polysilicon 1794 -1250 1794 -1250 0 3
rlabel polysilicon 1801 -1244 1801 -1244 0 1
rlabel polysilicon 1801 -1250 1801 -1250 0 3
rlabel polysilicon 1808 -1244 1808 -1244 0 1
rlabel polysilicon 1808 -1250 1808 -1250 0 3
rlabel polysilicon 1815 -1244 1815 -1244 0 1
rlabel polysilicon 1815 -1250 1815 -1250 0 3
rlabel polysilicon 1822 -1244 1822 -1244 0 1
rlabel polysilicon 1822 -1250 1822 -1250 0 3
rlabel polysilicon 1829 -1244 1829 -1244 0 1
rlabel polysilicon 1829 -1250 1829 -1250 0 3
rlabel polysilicon 1836 -1244 1836 -1244 0 1
rlabel polysilicon 1836 -1250 1836 -1250 0 3
rlabel polysilicon 1843 -1244 1843 -1244 0 1
rlabel polysilicon 1843 -1250 1843 -1250 0 3
rlabel polysilicon 1850 -1244 1850 -1244 0 1
rlabel polysilicon 1850 -1250 1850 -1250 0 3
rlabel polysilicon 1857 -1244 1857 -1244 0 1
rlabel polysilicon 1857 -1250 1857 -1250 0 3
rlabel polysilicon 1864 -1244 1864 -1244 0 1
rlabel polysilicon 1864 -1250 1864 -1250 0 3
rlabel polysilicon 1871 -1244 1871 -1244 0 1
rlabel polysilicon 1871 -1250 1871 -1250 0 3
rlabel polysilicon 1878 -1244 1878 -1244 0 1
rlabel polysilicon 1878 -1250 1878 -1250 0 3
rlabel polysilicon 1885 -1244 1885 -1244 0 1
rlabel polysilicon 1885 -1250 1885 -1250 0 3
rlabel polysilicon 1892 -1244 1892 -1244 0 1
rlabel polysilicon 1892 -1250 1892 -1250 0 3
rlabel polysilicon 1899 -1244 1899 -1244 0 1
rlabel polysilicon 1899 -1250 1899 -1250 0 3
rlabel polysilicon 1906 -1244 1906 -1244 0 1
rlabel polysilicon 1906 -1250 1906 -1250 0 3
rlabel polysilicon 1913 -1244 1913 -1244 0 1
rlabel polysilicon 1913 -1250 1913 -1250 0 3
rlabel polysilicon 1920 -1244 1920 -1244 0 1
rlabel polysilicon 1920 -1250 1920 -1250 0 3
rlabel polysilicon 1927 -1244 1927 -1244 0 1
rlabel polysilicon 1927 -1250 1927 -1250 0 3
rlabel polysilicon 1955 -1244 1955 -1244 0 1
rlabel polysilicon 1955 -1250 1955 -1250 0 3
rlabel polysilicon 1962 -1244 1962 -1244 0 1
rlabel polysilicon 1962 -1250 1962 -1250 0 3
rlabel polysilicon 1969 -1244 1969 -1244 0 1
rlabel polysilicon 1969 -1250 1969 -1250 0 3
rlabel polysilicon 1976 -1244 1976 -1244 0 1
rlabel polysilicon 1976 -1250 1976 -1250 0 3
rlabel polysilicon 1990 -1244 1990 -1244 0 1
rlabel polysilicon 1990 -1250 1990 -1250 0 3
rlabel polysilicon 9 -1387 9 -1387 0 1
rlabel polysilicon 9 -1393 9 -1393 0 3
rlabel polysilicon 16 -1387 16 -1387 0 1
rlabel polysilicon 16 -1393 16 -1393 0 3
rlabel polysilicon 23 -1387 23 -1387 0 1
rlabel polysilicon 23 -1393 23 -1393 0 3
rlabel polysilicon 30 -1387 30 -1387 0 1
rlabel polysilicon 30 -1393 30 -1393 0 3
rlabel polysilicon 37 -1387 37 -1387 0 1
rlabel polysilicon 37 -1393 37 -1393 0 3
rlabel polysilicon 44 -1387 44 -1387 0 1
rlabel polysilicon 44 -1393 44 -1393 0 3
rlabel polysilicon 51 -1387 51 -1387 0 1
rlabel polysilicon 54 -1387 54 -1387 0 2
rlabel polysilicon 51 -1393 51 -1393 0 3
rlabel polysilicon 58 -1387 58 -1387 0 1
rlabel polysilicon 58 -1393 58 -1393 0 3
rlabel polysilicon 61 -1393 61 -1393 0 4
rlabel polysilicon 65 -1387 65 -1387 0 1
rlabel polysilicon 65 -1393 65 -1393 0 3
rlabel polysilicon 72 -1387 72 -1387 0 1
rlabel polysilicon 75 -1387 75 -1387 0 2
rlabel polysilicon 75 -1393 75 -1393 0 4
rlabel polysilicon 79 -1387 79 -1387 0 1
rlabel polysilicon 79 -1393 79 -1393 0 3
rlabel polysilicon 86 -1387 86 -1387 0 1
rlabel polysilicon 86 -1393 86 -1393 0 3
rlabel polysilicon 93 -1387 93 -1387 0 1
rlabel polysilicon 93 -1393 93 -1393 0 3
rlabel polysilicon 100 -1387 100 -1387 0 1
rlabel polysilicon 100 -1393 100 -1393 0 3
rlabel polysilicon 107 -1387 107 -1387 0 1
rlabel polysilicon 110 -1387 110 -1387 0 2
rlabel polysilicon 110 -1393 110 -1393 0 4
rlabel polysilicon 114 -1387 114 -1387 0 1
rlabel polysilicon 114 -1393 114 -1393 0 3
rlabel polysilicon 121 -1387 121 -1387 0 1
rlabel polysilicon 121 -1393 121 -1393 0 3
rlabel polysilicon 128 -1387 128 -1387 0 1
rlabel polysilicon 128 -1393 128 -1393 0 3
rlabel polysilicon 131 -1393 131 -1393 0 4
rlabel polysilicon 135 -1387 135 -1387 0 1
rlabel polysilicon 135 -1393 135 -1393 0 3
rlabel polysilicon 142 -1387 142 -1387 0 1
rlabel polysilicon 145 -1387 145 -1387 0 2
rlabel polysilicon 145 -1393 145 -1393 0 4
rlabel polysilicon 152 -1387 152 -1387 0 2
rlabel polysilicon 149 -1393 149 -1393 0 3
rlabel polysilicon 152 -1393 152 -1393 0 4
rlabel polysilicon 156 -1387 156 -1387 0 1
rlabel polysilicon 156 -1393 156 -1393 0 3
rlabel polysilicon 163 -1387 163 -1387 0 1
rlabel polysilicon 163 -1393 163 -1393 0 3
rlabel polysilicon 166 -1393 166 -1393 0 4
rlabel polysilicon 170 -1387 170 -1387 0 1
rlabel polysilicon 170 -1393 170 -1393 0 3
rlabel polysilicon 177 -1387 177 -1387 0 1
rlabel polysilicon 177 -1393 177 -1393 0 3
rlabel polysilicon 184 -1387 184 -1387 0 1
rlabel polysilicon 184 -1393 184 -1393 0 3
rlabel polysilicon 191 -1387 191 -1387 0 1
rlabel polysilicon 191 -1393 191 -1393 0 3
rlabel polysilicon 198 -1387 198 -1387 0 1
rlabel polysilicon 198 -1393 198 -1393 0 3
rlabel polysilicon 205 -1387 205 -1387 0 1
rlabel polysilicon 208 -1387 208 -1387 0 2
rlabel polysilicon 208 -1393 208 -1393 0 4
rlabel polysilicon 212 -1387 212 -1387 0 1
rlabel polysilicon 212 -1393 212 -1393 0 3
rlabel polysilicon 219 -1387 219 -1387 0 1
rlabel polysilicon 219 -1393 219 -1393 0 3
rlabel polysilicon 226 -1387 226 -1387 0 1
rlabel polysilicon 226 -1393 226 -1393 0 3
rlabel polysilicon 233 -1387 233 -1387 0 1
rlabel polysilicon 233 -1393 233 -1393 0 3
rlabel polysilicon 240 -1387 240 -1387 0 1
rlabel polysilicon 240 -1393 240 -1393 0 3
rlabel polysilicon 247 -1387 247 -1387 0 1
rlabel polysilicon 247 -1393 247 -1393 0 3
rlabel polysilicon 254 -1387 254 -1387 0 1
rlabel polysilicon 254 -1393 254 -1393 0 3
rlabel polysilicon 261 -1387 261 -1387 0 1
rlabel polysilicon 261 -1393 261 -1393 0 3
rlabel polysilicon 268 -1387 268 -1387 0 1
rlabel polysilicon 268 -1393 268 -1393 0 3
rlabel polysilicon 275 -1387 275 -1387 0 1
rlabel polysilicon 275 -1393 275 -1393 0 3
rlabel polysilicon 282 -1387 282 -1387 0 1
rlabel polysilicon 282 -1393 282 -1393 0 3
rlabel polysilicon 289 -1387 289 -1387 0 1
rlabel polysilicon 289 -1393 289 -1393 0 3
rlabel polysilicon 296 -1387 296 -1387 0 1
rlabel polysilicon 296 -1393 296 -1393 0 3
rlabel polysilicon 303 -1387 303 -1387 0 1
rlabel polysilicon 303 -1393 303 -1393 0 3
rlabel polysilicon 310 -1387 310 -1387 0 1
rlabel polysilicon 310 -1393 310 -1393 0 3
rlabel polysilicon 317 -1387 317 -1387 0 1
rlabel polysilicon 317 -1393 317 -1393 0 3
rlabel polysilicon 324 -1387 324 -1387 0 1
rlabel polysilicon 324 -1393 324 -1393 0 3
rlabel polysilicon 331 -1393 331 -1393 0 3
rlabel polysilicon 338 -1387 338 -1387 0 1
rlabel polysilicon 338 -1393 338 -1393 0 3
rlabel polysilicon 345 -1387 345 -1387 0 1
rlabel polysilicon 345 -1393 345 -1393 0 3
rlabel polysilicon 352 -1387 352 -1387 0 1
rlabel polysilicon 352 -1393 352 -1393 0 3
rlabel polysilicon 359 -1387 359 -1387 0 1
rlabel polysilicon 359 -1393 359 -1393 0 3
rlabel polysilicon 366 -1387 366 -1387 0 1
rlabel polysilicon 366 -1393 366 -1393 0 3
rlabel polysilicon 373 -1387 373 -1387 0 1
rlabel polysilicon 373 -1393 373 -1393 0 3
rlabel polysilicon 380 -1387 380 -1387 0 1
rlabel polysilicon 380 -1393 380 -1393 0 3
rlabel polysilicon 387 -1387 387 -1387 0 1
rlabel polysilicon 387 -1393 387 -1393 0 3
rlabel polysilicon 394 -1387 394 -1387 0 1
rlabel polysilicon 394 -1393 394 -1393 0 3
rlabel polysilicon 401 -1387 401 -1387 0 1
rlabel polysilicon 401 -1393 401 -1393 0 3
rlabel polysilicon 408 -1387 408 -1387 0 1
rlabel polysilicon 408 -1393 408 -1393 0 3
rlabel polysilicon 415 -1387 415 -1387 0 1
rlabel polysilicon 415 -1393 415 -1393 0 3
rlabel polysilicon 422 -1387 422 -1387 0 1
rlabel polysilicon 422 -1393 422 -1393 0 3
rlabel polysilicon 429 -1387 429 -1387 0 1
rlabel polysilicon 432 -1387 432 -1387 0 2
rlabel polysilicon 429 -1393 429 -1393 0 3
rlabel polysilicon 432 -1393 432 -1393 0 4
rlabel polysilicon 436 -1387 436 -1387 0 1
rlabel polysilicon 436 -1393 436 -1393 0 3
rlabel polysilicon 443 -1387 443 -1387 0 1
rlabel polysilicon 443 -1393 443 -1393 0 3
rlabel polysilicon 450 -1387 450 -1387 0 1
rlabel polysilicon 450 -1393 450 -1393 0 3
rlabel polysilicon 457 -1387 457 -1387 0 1
rlabel polysilicon 457 -1393 457 -1393 0 3
rlabel polysilicon 464 -1387 464 -1387 0 1
rlabel polysilicon 464 -1393 464 -1393 0 3
rlabel polysilicon 471 -1387 471 -1387 0 1
rlabel polysilicon 471 -1393 471 -1393 0 3
rlabel polysilicon 478 -1387 478 -1387 0 1
rlabel polysilicon 478 -1393 478 -1393 0 3
rlabel polysilicon 485 -1387 485 -1387 0 1
rlabel polysilicon 485 -1393 485 -1393 0 3
rlabel polysilicon 492 -1387 492 -1387 0 1
rlabel polysilicon 492 -1393 492 -1393 0 3
rlabel polysilicon 499 -1387 499 -1387 0 1
rlabel polysilicon 499 -1393 499 -1393 0 3
rlabel polysilicon 506 -1387 506 -1387 0 1
rlabel polysilicon 506 -1393 506 -1393 0 3
rlabel polysilicon 513 -1387 513 -1387 0 1
rlabel polysilicon 513 -1393 513 -1393 0 3
rlabel polysilicon 520 -1387 520 -1387 0 1
rlabel polysilicon 520 -1393 520 -1393 0 3
rlabel polysilicon 527 -1387 527 -1387 0 1
rlabel polysilicon 530 -1387 530 -1387 0 2
rlabel polysilicon 527 -1393 527 -1393 0 3
rlabel polysilicon 530 -1393 530 -1393 0 4
rlabel polysilicon 534 -1387 534 -1387 0 1
rlabel polysilicon 534 -1393 534 -1393 0 3
rlabel polysilicon 541 -1387 541 -1387 0 1
rlabel polysilicon 541 -1393 541 -1393 0 3
rlabel polysilicon 548 -1387 548 -1387 0 1
rlabel polysilicon 548 -1393 548 -1393 0 3
rlabel polysilicon 555 -1387 555 -1387 0 1
rlabel polysilicon 555 -1393 555 -1393 0 3
rlabel polysilicon 562 -1387 562 -1387 0 1
rlabel polysilicon 562 -1393 562 -1393 0 3
rlabel polysilicon 569 -1387 569 -1387 0 1
rlabel polysilicon 569 -1393 569 -1393 0 3
rlabel polysilicon 579 -1387 579 -1387 0 2
rlabel polysilicon 576 -1393 576 -1393 0 3
rlabel polysilicon 579 -1393 579 -1393 0 4
rlabel polysilicon 583 -1387 583 -1387 0 1
rlabel polysilicon 583 -1393 583 -1393 0 3
rlabel polysilicon 590 -1387 590 -1387 0 1
rlabel polysilicon 590 -1393 590 -1393 0 3
rlabel polysilicon 597 -1387 597 -1387 0 1
rlabel polysilicon 597 -1393 597 -1393 0 3
rlabel polysilicon 604 -1387 604 -1387 0 1
rlabel polysilicon 604 -1393 604 -1393 0 3
rlabel polysilicon 611 -1387 611 -1387 0 1
rlabel polysilicon 611 -1393 611 -1393 0 3
rlabel polysilicon 618 -1387 618 -1387 0 1
rlabel polysilicon 618 -1393 618 -1393 0 3
rlabel polysilicon 625 -1387 625 -1387 0 1
rlabel polysilicon 628 -1387 628 -1387 0 2
rlabel polysilicon 625 -1393 625 -1393 0 3
rlabel polysilicon 628 -1393 628 -1393 0 4
rlabel polysilicon 632 -1387 632 -1387 0 1
rlabel polysilicon 632 -1393 632 -1393 0 3
rlabel polysilicon 639 -1387 639 -1387 0 1
rlabel polysilicon 639 -1393 639 -1393 0 3
rlabel polysilicon 646 -1387 646 -1387 0 1
rlabel polysilicon 646 -1393 646 -1393 0 3
rlabel polysilicon 653 -1387 653 -1387 0 1
rlabel polysilicon 656 -1387 656 -1387 0 2
rlabel polysilicon 653 -1393 653 -1393 0 3
rlabel polysilicon 656 -1393 656 -1393 0 4
rlabel polysilicon 660 -1387 660 -1387 0 1
rlabel polysilicon 660 -1393 660 -1393 0 3
rlabel polysilicon 667 -1387 667 -1387 0 1
rlabel polysilicon 670 -1387 670 -1387 0 2
rlabel polysilicon 667 -1393 667 -1393 0 3
rlabel polysilicon 674 -1387 674 -1387 0 1
rlabel polysilicon 677 -1387 677 -1387 0 2
rlabel polysilicon 677 -1393 677 -1393 0 4
rlabel polysilicon 681 -1387 681 -1387 0 1
rlabel polysilicon 681 -1393 681 -1393 0 3
rlabel polysilicon 688 -1387 688 -1387 0 1
rlabel polysilicon 688 -1393 688 -1393 0 3
rlabel polysilicon 695 -1387 695 -1387 0 1
rlabel polysilicon 695 -1393 695 -1393 0 3
rlabel polysilicon 702 -1387 702 -1387 0 1
rlabel polysilicon 702 -1393 702 -1393 0 3
rlabel polysilicon 709 -1387 709 -1387 0 1
rlabel polysilicon 712 -1387 712 -1387 0 2
rlabel polysilicon 709 -1393 709 -1393 0 3
rlabel polysilicon 712 -1393 712 -1393 0 4
rlabel polysilicon 716 -1387 716 -1387 0 1
rlabel polysilicon 716 -1393 716 -1393 0 3
rlabel polysilicon 723 -1387 723 -1387 0 1
rlabel polysilicon 723 -1393 723 -1393 0 3
rlabel polysilicon 730 -1387 730 -1387 0 1
rlabel polysilicon 730 -1393 730 -1393 0 3
rlabel polysilicon 737 -1387 737 -1387 0 1
rlabel polysilicon 737 -1393 737 -1393 0 3
rlabel polysilicon 744 -1387 744 -1387 0 1
rlabel polysilicon 744 -1393 744 -1393 0 3
rlabel polysilicon 751 -1387 751 -1387 0 1
rlabel polysilicon 751 -1393 751 -1393 0 3
rlabel polysilicon 758 -1387 758 -1387 0 1
rlabel polysilicon 758 -1393 758 -1393 0 3
rlabel polysilicon 765 -1387 765 -1387 0 1
rlabel polysilicon 765 -1393 765 -1393 0 3
rlabel polysilicon 772 -1387 772 -1387 0 1
rlabel polysilicon 772 -1393 772 -1393 0 3
rlabel polysilicon 779 -1387 779 -1387 0 1
rlabel polysilicon 779 -1393 779 -1393 0 3
rlabel polysilicon 786 -1387 786 -1387 0 1
rlabel polysilicon 786 -1393 786 -1393 0 3
rlabel polysilicon 793 -1387 793 -1387 0 1
rlabel polysilicon 793 -1393 793 -1393 0 3
rlabel polysilicon 800 -1387 800 -1387 0 1
rlabel polysilicon 800 -1393 800 -1393 0 3
rlabel polysilicon 807 -1387 807 -1387 0 1
rlabel polysilicon 807 -1393 807 -1393 0 3
rlabel polysilicon 814 -1387 814 -1387 0 1
rlabel polysilicon 814 -1393 814 -1393 0 3
rlabel polysilicon 821 -1387 821 -1387 0 1
rlabel polysilicon 821 -1393 821 -1393 0 3
rlabel polysilicon 828 -1387 828 -1387 0 1
rlabel polysilicon 828 -1393 828 -1393 0 3
rlabel polysilicon 835 -1387 835 -1387 0 1
rlabel polysilicon 838 -1387 838 -1387 0 2
rlabel polysilicon 835 -1393 835 -1393 0 3
rlabel polysilicon 842 -1387 842 -1387 0 1
rlabel polysilicon 842 -1393 842 -1393 0 3
rlabel polysilicon 849 -1387 849 -1387 0 1
rlabel polysilicon 849 -1393 849 -1393 0 3
rlabel polysilicon 856 -1387 856 -1387 0 1
rlabel polysilicon 859 -1387 859 -1387 0 2
rlabel polysilicon 856 -1393 856 -1393 0 3
rlabel polysilicon 859 -1393 859 -1393 0 4
rlabel polysilicon 863 -1387 863 -1387 0 1
rlabel polysilicon 863 -1393 863 -1393 0 3
rlabel polysilicon 870 -1387 870 -1387 0 1
rlabel polysilicon 870 -1393 870 -1393 0 3
rlabel polysilicon 877 -1387 877 -1387 0 1
rlabel polysilicon 877 -1393 877 -1393 0 3
rlabel polysilicon 884 -1387 884 -1387 0 1
rlabel polysilicon 884 -1393 884 -1393 0 3
rlabel polysilicon 891 -1387 891 -1387 0 1
rlabel polysilicon 891 -1393 891 -1393 0 3
rlabel polysilicon 898 -1387 898 -1387 0 1
rlabel polysilicon 898 -1393 898 -1393 0 3
rlabel polysilicon 905 -1387 905 -1387 0 1
rlabel polysilicon 905 -1393 905 -1393 0 3
rlabel polysilicon 912 -1387 912 -1387 0 1
rlabel polysilicon 912 -1393 912 -1393 0 3
rlabel polysilicon 919 -1387 919 -1387 0 1
rlabel polysilicon 922 -1387 922 -1387 0 2
rlabel polysilicon 919 -1393 919 -1393 0 3
rlabel polysilicon 922 -1393 922 -1393 0 4
rlabel polysilicon 929 -1387 929 -1387 0 2
rlabel polysilicon 926 -1393 926 -1393 0 3
rlabel polysilicon 929 -1393 929 -1393 0 4
rlabel polysilicon 933 -1387 933 -1387 0 1
rlabel polysilicon 933 -1393 933 -1393 0 3
rlabel polysilicon 943 -1387 943 -1387 0 2
rlabel polysilicon 940 -1393 940 -1393 0 3
rlabel polysilicon 943 -1393 943 -1393 0 4
rlabel polysilicon 947 -1387 947 -1387 0 1
rlabel polysilicon 947 -1393 947 -1393 0 3
rlabel polysilicon 954 -1387 954 -1387 0 1
rlabel polysilicon 954 -1393 954 -1393 0 3
rlabel polysilicon 961 -1387 961 -1387 0 1
rlabel polysilicon 961 -1393 961 -1393 0 3
rlabel polysilicon 968 -1387 968 -1387 0 1
rlabel polysilicon 968 -1393 968 -1393 0 3
rlabel polysilicon 975 -1387 975 -1387 0 1
rlabel polysilicon 975 -1393 975 -1393 0 3
rlabel polysilicon 982 -1387 982 -1387 0 1
rlabel polysilicon 982 -1393 982 -1393 0 3
rlabel polysilicon 989 -1387 989 -1387 0 1
rlabel polysilicon 989 -1393 989 -1393 0 3
rlabel polysilicon 996 -1387 996 -1387 0 1
rlabel polysilicon 999 -1387 999 -1387 0 2
rlabel polysilicon 996 -1393 996 -1393 0 3
rlabel polysilicon 999 -1393 999 -1393 0 4
rlabel polysilicon 1003 -1387 1003 -1387 0 1
rlabel polysilicon 1003 -1393 1003 -1393 0 3
rlabel polysilicon 1010 -1387 1010 -1387 0 1
rlabel polysilicon 1010 -1393 1010 -1393 0 3
rlabel polysilicon 1017 -1387 1017 -1387 0 1
rlabel polysilicon 1017 -1393 1017 -1393 0 3
rlabel polysilicon 1024 -1387 1024 -1387 0 1
rlabel polysilicon 1024 -1393 1024 -1393 0 3
rlabel polysilicon 1031 -1387 1031 -1387 0 1
rlabel polysilicon 1031 -1393 1031 -1393 0 3
rlabel polysilicon 1034 -1393 1034 -1393 0 4
rlabel polysilicon 1038 -1387 1038 -1387 0 1
rlabel polysilicon 1038 -1393 1038 -1393 0 3
rlabel polysilicon 1045 -1387 1045 -1387 0 1
rlabel polysilicon 1052 -1387 1052 -1387 0 1
rlabel polysilicon 1055 -1387 1055 -1387 0 2
rlabel polysilicon 1052 -1393 1052 -1393 0 3
rlabel polysilicon 1055 -1393 1055 -1393 0 4
rlabel polysilicon 1059 -1387 1059 -1387 0 1
rlabel polysilicon 1059 -1393 1059 -1393 0 3
rlabel polysilicon 1066 -1387 1066 -1387 0 1
rlabel polysilicon 1069 -1387 1069 -1387 0 2
rlabel polysilicon 1066 -1393 1066 -1393 0 3
rlabel polysilicon 1069 -1393 1069 -1393 0 4
rlabel polysilicon 1073 -1387 1073 -1387 0 1
rlabel polysilicon 1076 -1387 1076 -1387 0 2
rlabel polysilicon 1076 -1393 1076 -1393 0 4
rlabel polysilicon 1080 -1387 1080 -1387 0 1
rlabel polysilicon 1080 -1393 1080 -1393 0 3
rlabel polysilicon 1087 -1387 1087 -1387 0 1
rlabel polysilicon 1087 -1393 1087 -1393 0 3
rlabel polysilicon 1094 -1387 1094 -1387 0 1
rlabel polysilicon 1094 -1393 1094 -1393 0 3
rlabel polysilicon 1101 -1387 1101 -1387 0 1
rlabel polysilicon 1101 -1393 1101 -1393 0 3
rlabel polysilicon 1108 -1387 1108 -1387 0 1
rlabel polysilicon 1111 -1387 1111 -1387 0 2
rlabel polysilicon 1108 -1393 1108 -1393 0 3
rlabel polysilicon 1111 -1393 1111 -1393 0 4
rlabel polysilicon 1115 -1387 1115 -1387 0 1
rlabel polysilicon 1115 -1393 1115 -1393 0 3
rlabel polysilicon 1122 -1387 1122 -1387 0 1
rlabel polysilicon 1122 -1393 1122 -1393 0 3
rlabel polysilicon 1129 -1387 1129 -1387 0 1
rlabel polysilicon 1129 -1393 1129 -1393 0 3
rlabel polysilicon 1136 -1387 1136 -1387 0 1
rlabel polysilicon 1136 -1393 1136 -1393 0 3
rlabel polysilicon 1143 -1387 1143 -1387 0 1
rlabel polysilicon 1143 -1393 1143 -1393 0 3
rlabel polysilicon 1150 -1387 1150 -1387 0 1
rlabel polysilicon 1150 -1393 1150 -1393 0 3
rlabel polysilicon 1157 -1387 1157 -1387 0 1
rlabel polysilicon 1157 -1393 1157 -1393 0 3
rlabel polysilicon 1164 -1387 1164 -1387 0 1
rlabel polysilicon 1164 -1393 1164 -1393 0 3
rlabel polysilicon 1171 -1387 1171 -1387 0 1
rlabel polysilicon 1171 -1393 1171 -1393 0 3
rlabel polysilicon 1178 -1387 1178 -1387 0 1
rlabel polysilicon 1178 -1393 1178 -1393 0 3
rlabel polysilicon 1185 -1387 1185 -1387 0 1
rlabel polysilicon 1185 -1393 1185 -1393 0 3
rlabel polysilicon 1192 -1387 1192 -1387 0 1
rlabel polysilicon 1192 -1393 1192 -1393 0 3
rlabel polysilicon 1199 -1387 1199 -1387 0 1
rlabel polysilicon 1199 -1393 1199 -1393 0 3
rlabel polysilicon 1206 -1387 1206 -1387 0 1
rlabel polysilicon 1206 -1393 1206 -1393 0 3
rlabel polysilicon 1213 -1387 1213 -1387 0 1
rlabel polysilicon 1213 -1393 1213 -1393 0 3
rlabel polysilicon 1220 -1387 1220 -1387 0 1
rlabel polysilicon 1220 -1393 1220 -1393 0 3
rlabel polysilicon 1227 -1387 1227 -1387 0 1
rlabel polysilicon 1227 -1393 1227 -1393 0 3
rlabel polysilicon 1234 -1387 1234 -1387 0 1
rlabel polysilicon 1234 -1393 1234 -1393 0 3
rlabel polysilicon 1241 -1387 1241 -1387 0 1
rlabel polysilicon 1244 -1387 1244 -1387 0 2
rlabel polysilicon 1241 -1393 1241 -1393 0 3
rlabel polysilicon 1244 -1393 1244 -1393 0 4
rlabel polysilicon 1248 -1387 1248 -1387 0 1
rlabel polysilicon 1248 -1393 1248 -1393 0 3
rlabel polysilicon 1255 -1387 1255 -1387 0 1
rlabel polysilicon 1255 -1393 1255 -1393 0 3
rlabel polysilicon 1262 -1387 1262 -1387 0 1
rlabel polysilicon 1262 -1393 1262 -1393 0 3
rlabel polysilicon 1269 -1387 1269 -1387 0 1
rlabel polysilicon 1269 -1393 1269 -1393 0 3
rlabel polysilicon 1276 -1387 1276 -1387 0 1
rlabel polysilicon 1276 -1393 1276 -1393 0 3
rlabel polysilicon 1283 -1387 1283 -1387 0 1
rlabel polysilicon 1283 -1393 1283 -1393 0 3
rlabel polysilicon 1286 -1393 1286 -1393 0 4
rlabel polysilicon 1290 -1387 1290 -1387 0 1
rlabel polysilicon 1290 -1393 1290 -1393 0 3
rlabel polysilicon 1297 -1387 1297 -1387 0 1
rlabel polysilicon 1297 -1393 1297 -1393 0 3
rlabel polysilicon 1304 -1387 1304 -1387 0 1
rlabel polysilicon 1304 -1393 1304 -1393 0 3
rlabel polysilicon 1311 -1387 1311 -1387 0 1
rlabel polysilicon 1311 -1393 1311 -1393 0 3
rlabel polysilicon 1318 -1387 1318 -1387 0 1
rlabel polysilicon 1318 -1393 1318 -1393 0 3
rlabel polysilicon 1325 -1387 1325 -1387 0 1
rlabel polysilicon 1325 -1393 1325 -1393 0 3
rlabel polysilicon 1332 -1387 1332 -1387 0 1
rlabel polysilicon 1332 -1393 1332 -1393 0 3
rlabel polysilicon 1339 -1387 1339 -1387 0 1
rlabel polysilicon 1339 -1393 1339 -1393 0 3
rlabel polysilicon 1346 -1387 1346 -1387 0 1
rlabel polysilicon 1346 -1393 1346 -1393 0 3
rlabel polysilicon 1353 -1387 1353 -1387 0 1
rlabel polysilicon 1353 -1393 1353 -1393 0 3
rlabel polysilicon 1360 -1387 1360 -1387 0 1
rlabel polysilicon 1360 -1393 1360 -1393 0 3
rlabel polysilicon 1367 -1387 1367 -1387 0 1
rlabel polysilicon 1367 -1393 1367 -1393 0 3
rlabel polysilicon 1374 -1387 1374 -1387 0 1
rlabel polysilicon 1374 -1393 1374 -1393 0 3
rlabel polysilicon 1381 -1387 1381 -1387 0 1
rlabel polysilicon 1381 -1393 1381 -1393 0 3
rlabel polysilicon 1388 -1387 1388 -1387 0 1
rlabel polysilicon 1391 -1387 1391 -1387 0 2
rlabel polysilicon 1388 -1393 1388 -1393 0 3
rlabel polysilicon 1395 -1387 1395 -1387 0 1
rlabel polysilicon 1395 -1393 1395 -1393 0 3
rlabel polysilicon 1402 -1387 1402 -1387 0 1
rlabel polysilicon 1402 -1393 1402 -1393 0 3
rlabel polysilicon 1409 -1387 1409 -1387 0 1
rlabel polysilicon 1409 -1393 1409 -1393 0 3
rlabel polysilicon 1416 -1387 1416 -1387 0 1
rlabel polysilicon 1416 -1393 1416 -1393 0 3
rlabel polysilicon 1423 -1387 1423 -1387 0 1
rlabel polysilicon 1423 -1393 1423 -1393 0 3
rlabel polysilicon 1430 -1387 1430 -1387 0 1
rlabel polysilicon 1430 -1393 1430 -1393 0 3
rlabel polysilicon 1437 -1387 1437 -1387 0 1
rlabel polysilicon 1437 -1393 1437 -1393 0 3
rlabel polysilicon 1444 -1387 1444 -1387 0 1
rlabel polysilicon 1444 -1393 1444 -1393 0 3
rlabel polysilicon 1451 -1387 1451 -1387 0 1
rlabel polysilicon 1451 -1393 1451 -1393 0 3
rlabel polysilicon 1458 -1387 1458 -1387 0 1
rlabel polysilicon 1458 -1393 1458 -1393 0 3
rlabel polysilicon 1465 -1387 1465 -1387 0 1
rlabel polysilicon 1465 -1393 1465 -1393 0 3
rlabel polysilicon 1472 -1387 1472 -1387 0 1
rlabel polysilicon 1472 -1393 1472 -1393 0 3
rlabel polysilicon 1479 -1387 1479 -1387 0 1
rlabel polysilicon 1479 -1393 1479 -1393 0 3
rlabel polysilicon 1486 -1387 1486 -1387 0 1
rlabel polysilicon 1486 -1393 1486 -1393 0 3
rlabel polysilicon 1493 -1387 1493 -1387 0 1
rlabel polysilicon 1493 -1393 1493 -1393 0 3
rlabel polysilicon 1500 -1387 1500 -1387 0 1
rlabel polysilicon 1500 -1393 1500 -1393 0 3
rlabel polysilicon 1507 -1387 1507 -1387 0 1
rlabel polysilicon 1507 -1393 1507 -1393 0 3
rlabel polysilicon 1514 -1387 1514 -1387 0 1
rlabel polysilicon 1514 -1393 1514 -1393 0 3
rlabel polysilicon 1521 -1387 1521 -1387 0 1
rlabel polysilicon 1521 -1393 1521 -1393 0 3
rlabel polysilicon 1528 -1387 1528 -1387 0 1
rlabel polysilicon 1528 -1393 1528 -1393 0 3
rlabel polysilicon 1535 -1387 1535 -1387 0 1
rlabel polysilicon 1535 -1393 1535 -1393 0 3
rlabel polysilicon 1542 -1387 1542 -1387 0 1
rlabel polysilicon 1542 -1393 1542 -1393 0 3
rlabel polysilicon 1549 -1387 1549 -1387 0 1
rlabel polysilicon 1549 -1393 1549 -1393 0 3
rlabel polysilicon 1556 -1387 1556 -1387 0 1
rlabel polysilicon 1556 -1393 1556 -1393 0 3
rlabel polysilicon 1563 -1387 1563 -1387 0 1
rlabel polysilicon 1563 -1393 1563 -1393 0 3
rlabel polysilicon 1570 -1387 1570 -1387 0 1
rlabel polysilicon 1570 -1393 1570 -1393 0 3
rlabel polysilicon 1577 -1387 1577 -1387 0 1
rlabel polysilicon 1577 -1393 1577 -1393 0 3
rlabel polysilicon 1584 -1387 1584 -1387 0 1
rlabel polysilicon 1584 -1393 1584 -1393 0 3
rlabel polysilicon 1591 -1387 1591 -1387 0 1
rlabel polysilicon 1591 -1393 1591 -1393 0 3
rlabel polysilicon 1598 -1387 1598 -1387 0 1
rlabel polysilicon 1598 -1393 1598 -1393 0 3
rlabel polysilicon 1605 -1387 1605 -1387 0 1
rlabel polysilicon 1605 -1393 1605 -1393 0 3
rlabel polysilicon 1612 -1387 1612 -1387 0 1
rlabel polysilicon 1612 -1393 1612 -1393 0 3
rlabel polysilicon 1619 -1387 1619 -1387 0 1
rlabel polysilicon 1619 -1393 1619 -1393 0 3
rlabel polysilicon 1626 -1387 1626 -1387 0 1
rlabel polysilicon 1626 -1393 1626 -1393 0 3
rlabel polysilicon 1633 -1387 1633 -1387 0 1
rlabel polysilicon 1633 -1393 1633 -1393 0 3
rlabel polysilicon 1640 -1387 1640 -1387 0 1
rlabel polysilicon 1640 -1393 1640 -1393 0 3
rlabel polysilicon 1647 -1387 1647 -1387 0 1
rlabel polysilicon 1647 -1393 1647 -1393 0 3
rlabel polysilicon 1654 -1387 1654 -1387 0 1
rlabel polysilicon 1654 -1393 1654 -1393 0 3
rlabel polysilicon 1661 -1387 1661 -1387 0 1
rlabel polysilicon 1661 -1393 1661 -1393 0 3
rlabel polysilicon 1668 -1387 1668 -1387 0 1
rlabel polysilicon 1668 -1393 1668 -1393 0 3
rlabel polysilicon 1675 -1387 1675 -1387 0 1
rlabel polysilicon 1675 -1393 1675 -1393 0 3
rlabel polysilicon 1682 -1387 1682 -1387 0 1
rlabel polysilicon 1682 -1393 1682 -1393 0 3
rlabel polysilicon 1689 -1387 1689 -1387 0 1
rlabel polysilicon 1689 -1393 1689 -1393 0 3
rlabel polysilicon 1696 -1387 1696 -1387 0 1
rlabel polysilicon 1696 -1393 1696 -1393 0 3
rlabel polysilicon 1703 -1387 1703 -1387 0 1
rlabel polysilicon 1703 -1393 1703 -1393 0 3
rlabel polysilicon 1710 -1387 1710 -1387 0 1
rlabel polysilicon 1710 -1393 1710 -1393 0 3
rlabel polysilicon 1717 -1387 1717 -1387 0 1
rlabel polysilicon 1717 -1393 1717 -1393 0 3
rlabel polysilicon 1724 -1387 1724 -1387 0 1
rlabel polysilicon 1724 -1393 1724 -1393 0 3
rlabel polysilicon 1731 -1387 1731 -1387 0 1
rlabel polysilicon 1731 -1393 1731 -1393 0 3
rlabel polysilicon 1738 -1387 1738 -1387 0 1
rlabel polysilicon 1738 -1393 1738 -1393 0 3
rlabel polysilicon 1745 -1387 1745 -1387 0 1
rlabel polysilicon 1745 -1393 1745 -1393 0 3
rlabel polysilicon 1752 -1387 1752 -1387 0 1
rlabel polysilicon 1752 -1393 1752 -1393 0 3
rlabel polysilicon 1759 -1387 1759 -1387 0 1
rlabel polysilicon 1759 -1393 1759 -1393 0 3
rlabel polysilicon 1766 -1387 1766 -1387 0 1
rlabel polysilicon 1766 -1393 1766 -1393 0 3
rlabel polysilicon 1773 -1387 1773 -1387 0 1
rlabel polysilicon 1773 -1393 1773 -1393 0 3
rlabel polysilicon 1780 -1387 1780 -1387 0 1
rlabel polysilicon 1780 -1393 1780 -1393 0 3
rlabel polysilicon 1787 -1387 1787 -1387 0 1
rlabel polysilicon 1787 -1393 1787 -1393 0 3
rlabel polysilicon 1794 -1387 1794 -1387 0 1
rlabel polysilicon 1794 -1393 1794 -1393 0 3
rlabel polysilicon 1801 -1387 1801 -1387 0 1
rlabel polysilicon 1801 -1393 1801 -1393 0 3
rlabel polysilicon 1808 -1387 1808 -1387 0 1
rlabel polysilicon 1808 -1393 1808 -1393 0 3
rlabel polysilicon 1815 -1387 1815 -1387 0 1
rlabel polysilicon 1815 -1393 1815 -1393 0 3
rlabel polysilicon 1822 -1387 1822 -1387 0 1
rlabel polysilicon 1822 -1393 1822 -1393 0 3
rlabel polysilicon 1829 -1387 1829 -1387 0 1
rlabel polysilicon 1829 -1393 1829 -1393 0 3
rlabel polysilicon 1836 -1387 1836 -1387 0 1
rlabel polysilicon 1836 -1393 1836 -1393 0 3
rlabel polysilicon 1843 -1387 1843 -1387 0 1
rlabel polysilicon 1843 -1393 1843 -1393 0 3
rlabel polysilicon 1850 -1387 1850 -1387 0 1
rlabel polysilicon 1850 -1393 1850 -1393 0 3
rlabel polysilicon 1857 -1387 1857 -1387 0 1
rlabel polysilicon 1857 -1393 1857 -1393 0 3
rlabel polysilicon 1864 -1387 1864 -1387 0 1
rlabel polysilicon 1864 -1393 1864 -1393 0 3
rlabel polysilicon 1871 -1387 1871 -1387 0 1
rlabel polysilicon 1871 -1393 1871 -1393 0 3
rlabel polysilicon 1878 -1387 1878 -1387 0 1
rlabel polysilicon 1878 -1393 1878 -1393 0 3
rlabel polysilicon 1885 -1387 1885 -1387 0 1
rlabel polysilicon 1885 -1393 1885 -1393 0 3
rlabel polysilicon 1892 -1387 1892 -1387 0 1
rlabel polysilicon 1892 -1393 1892 -1393 0 3
rlabel polysilicon 1899 -1387 1899 -1387 0 1
rlabel polysilicon 1899 -1393 1899 -1393 0 3
rlabel polysilicon 1906 -1387 1906 -1387 0 1
rlabel polysilicon 1906 -1393 1906 -1393 0 3
rlabel polysilicon 1913 -1387 1913 -1387 0 1
rlabel polysilicon 1916 -1387 1916 -1387 0 2
rlabel polysilicon 1913 -1393 1913 -1393 0 3
rlabel polysilicon 1916 -1393 1916 -1393 0 4
rlabel polysilicon 1920 -1387 1920 -1387 0 1
rlabel polysilicon 1920 -1393 1920 -1393 0 3
rlabel polysilicon 1927 -1387 1927 -1387 0 1
rlabel polysilicon 1927 -1393 1927 -1393 0 3
rlabel polysilicon 1934 -1387 1934 -1387 0 1
rlabel polysilicon 1934 -1393 1934 -1393 0 3
rlabel polysilicon 1941 -1387 1941 -1387 0 1
rlabel polysilicon 1941 -1393 1941 -1393 0 3
rlabel polysilicon 1948 -1387 1948 -1387 0 1
rlabel polysilicon 1948 -1393 1948 -1393 0 3
rlabel polysilicon 1969 -1387 1969 -1387 0 1
rlabel polysilicon 1969 -1393 1969 -1393 0 3
rlabel polysilicon 1976 -1387 1976 -1387 0 1
rlabel polysilicon 1976 -1393 1976 -1393 0 3
rlabel polysilicon 1983 -1387 1983 -1387 0 1
rlabel polysilicon 1983 -1393 1983 -1393 0 3
rlabel polysilicon 1986 -1393 1986 -1393 0 4
rlabel polysilicon 1990 -1387 1990 -1387 0 1
rlabel polysilicon 1990 -1393 1990 -1393 0 3
rlabel polysilicon 1997 -1387 1997 -1387 0 1
rlabel polysilicon 1997 -1393 1997 -1393 0 3
rlabel polysilicon 2 -1518 2 -1518 0 1
rlabel polysilicon 2 -1524 2 -1524 0 3
rlabel polysilicon 9 -1518 9 -1518 0 1
rlabel polysilicon 9 -1524 9 -1524 0 3
rlabel polysilicon 16 -1518 16 -1518 0 1
rlabel polysilicon 16 -1524 16 -1524 0 3
rlabel polysilicon 23 -1518 23 -1518 0 1
rlabel polysilicon 23 -1524 23 -1524 0 3
rlabel polysilicon 30 -1518 30 -1518 0 1
rlabel polysilicon 30 -1524 30 -1524 0 3
rlabel polysilicon 37 -1518 37 -1518 0 1
rlabel polysilicon 37 -1524 37 -1524 0 3
rlabel polysilicon 44 -1518 44 -1518 0 1
rlabel polysilicon 47 -1518 47 -1518 0 2
rlabel polysilicon 44 -1524 44 -1524 0 3
rlabel polysilicon 47 -1524 47 -1524 0 4
rlabel polysilicon 51 -1518 51 -1518 0 1
rlabel polysilicon 51 -1524 51 -1524 0 3
rlabel polysilicon 58 -1518 58 -1518 0 1
rlabel polysilicon 61 -1518 61 -1518 0 2
rlabel polysilicon 58 -1524 58 -1524 0 3
rlabel polysilicon 65 -1518 65 -1518 0 1
rlabel polysilicon 65 -1524 65 -1524 0 3
rlabel polysilicon 72 -1518 72 -1518 0 1
rlabel polysilicon 72 -1524 72 -1524 0 3
rlabel polysilicon 79 -1518 79 -1518 0 1
rlabel polysilicon 82 -1518 82 -1518 0 2
rlabel polysilicon 79 -1524 79 -1524 0 3
rlabel polysilicon 82 -1524 82 -1524 0 4
rlabel polysilicon 86 -1518 86 -1518 0 1
rlabel polysilicon 86 -1524 86 -1524 0 3
rlabel polysilicon 93 -1518 93 -1518 0 1
rlabel polysilicon 93 -1524 93 -1524 0 3
rlabel polysilicon 100 -1518 100 -1518 0 1
rlabel polysilicon 100 -1524 100 -1524 0 3
rlabel polysilicon 107 -1518 107 -1518 0 1
rlabel polysilicon 107 -1524 107 -1524 0 3
rlabel polysilicon 114 -1518 114 -1518 0 1
rlabel polysilicon 114 -1524 114 -1524 0 3
rlabel polysilicon 121 -1518 121 -1518 0 1
rlabel polysilicon 121 -1524 121 -1524 0 3
rlabel polysilicon 128 -1518 128 -1518 0 1
rlabel polysilicon 128 -1524 128 -1524 0 3
rlabel polysilicon 135 -1518 135 -1518 0 1
rlabel polysilicon 135 -1524 135 -1524 0 3
rlabel polysilicon 142 -1518 142 -1518 0 1
rlabel polysilicon 145 -1518 145 -1518 0 2
rlabel polysilicon 142 -1524 142 -1524 0 3
rlabel polysilicon 145 -1524 145 -1524 0 4
rlabel polysilicon 149 -1518 149 -1518 0 1
rlabel polysilicon 149 -1524 149 -1524 0 3
rlabel polysilicon 156 -1518 156 -1518 0 1
rlabel polysilicon 156 -1524 156 -1524 0 3
rlabel polysilicon 163 -1518 163 -1518 0 1
rlabel polysilicon 163 -1524 163 -1524 0 3
rlabel polysilicon 170 -1518 170 -1518 0 1
rlabel polysilicon 170 -1524 170 -1524 0 3
rlabel polysilicon 177 -1518 177 -1518 0 1
rlabel polysilicon 177 -1524 177 -1524 0 3
rlabel polysilicon 184 -1518 184 -1518 0 1
rlabel polysilicon 184 -1524 184 -1524 0 3
rlabel polysilicon 191 -1518 191 -1518 0 1
rlabel polysilicon 194 -1518 194 -1518 0 2
rlabel polysilicon 191 -1524 191 -1524 0 3
rlabel polysilicon 194 -1524 194 -1524 0 4
rlabel polysilicon 198 -1518 198 -1518 0 1
rlabel polysilicon 198 -1524 198 -1524 0 3
rlabel polysilicon 205 -1518 205 -1518 0 1
rlabel polysilicon 205 -1524 205 -1524 0 3
rlabel polysilicon 212 -1518 212 -1518 0 1
rlabel polysilicon 215 -1518 215 -1518 0 2
rlabel polysilicon 212 -1524 212 -1524 0 3
rlabel polysilicon 219 -1518 219 -1518 0 1
rlabel polysilicon 219 -1524 219 -1524 0 3
rlabel polysilicon 226 -1518 226 -1518 0 1
rlabel polysilicon 226 -1524 226 -1524 0 3
rlabel polysilicon 233 -1518 233 -1518 0 1
rlabel polysilicon 233 -1524 233 -1524 0 3
rlabel polysilicon 240 -1518 240 -1518 0 1
rlabel polysilicon 243 -1518 243 -1518 0 2
rlabel polysilicon 240 -1524 240 -1524 0 3
rlabel polysilicon 247 -1518 247 -1518 0 1
rlabel polysilicon 247 -1524 247 -1524 0 3
rlabel polysilicon 254 -1518 254 -1518 0 1
rlabel polysilicon 254 -1524 254 -1524 0 3
rlabel polysilicon 261 -1518 261 -1518 0 1
rlabel polysilicon 261 -1524 261 -1524 0 3
rlabel polysilicon 268 -1518 268 -1518 0 1
rlabel polysilicon 268 -1524 268 -1524 0 3
rlabel polysilicon 275 -1518 275 -1518 0 1
rlabel polysilicon 275 -1524 275 -1524 0 3
rlabel polysilicon 282 -1518 282 -1518 0 1
rlabel polysilicon 282 -1524 282 -1524 0 3
rlabel polysilicon 289 -1518 289 -1518 0 1
rlabel polysilicon 289 -1524 289 -1524 0 3
rlabel polysilicon 296 -1518 296 -1518 0 1
rlabel polysilicon 296 -1524 296 -1524 0 3
rlabel polysilicon 303 -1518 303 -1518 0 1
rlabel polysilicon 303 -1524 303 -1524 0 3
rlabel polysilicon 310 -1518 310 -1518 0 1
rlabel polysilicon 310 -1524 310 -1524 0 3
rlabel polysilicon 317 -1518 317 -1518 0 1
rlabel polysilicon 317 -1524 317 -1524 0 3
rlabel polysilicon 324 -1518 324 -1518 0 1
rlabel polysilicon 324 -1524 324 -1524 0 3
rlabel polysilicon 331 -1518 331 -1518 0 1
rlabel polysilicon 331 -1524 331 -1524 0 3
rlabel polysilicon 338 -1518 338 -1518 0 1
rlabel polysilicon 338 -1524 338 -1524 0 3
rlabel polysilicon 345 -1518 345 -1518 0 1
rlabel polysilicon 345 -1524 345 -1524 0 3
rlabel polysilicon 352 -1518 352 -1518 0 1
rlabel polysilicon 352 -1524 352 -1524 0 3
rlabel polysilicon 359 -1518 359 -1518 0 1
rlabel polysilicon 359 -1524 359 -1524 0 3
rlabel polysilicon 366 -1518 366 -1518 0 1
rlabel polysilicon 366 -1524 366 -1524 0 3
rlabel polysilicon 373 -1518 373 -1518 0 1
rlabel polysilicon 373 -1524 373 -1524 0 3
rlabel polysilicon 380 -1518 380 -1518 0 1
rlabel polysilicon 380 -1524 380 -1524 0 3
rlabel polysilicon 387 -1518 387 -1518 0 1
rlabel polysilicon 387 -1524 387 -1524 0 3
rlabel polysilicon 394 -1518 394 -1518 0 1
rlabel polysilicon 394 -1524 394 -1524 0 3
rlabel polysilicon 401 -1518 401 -1518 0 1
rlabel polysilicon 401 -1524 401 -1524 0 3
rlabel polysilicon 408 -1518 408 -1518 0 1
rlabel polysilicon 408 -1524 408 -1524 0 3
rlabel polysilicon 415 -1518 415 -1518 0 1
rlabel polysilicon 415 -1524 415 -1524 0 3
rlabel polysilicon 422 -1518 422 -1518 0 1
rlabel polysilicon 422 -1524 422 -1524 0 3
rlabel polysilicon 429 -1518 429 -1518 0 1
rlabel polysilicon 429 -1524 429 -1524 0 3
rlabel polysilicon 436 -1518 436 -1518 0 1
rlabel polysilicon 436 -1524 436 -1524 0 3
rlabel polysilicon 443 -1518 443 -1518 0 1
rlabel polysilicon 443 -1524 443 -1524 0 3
rlabel polysilicon 450 -1518 450 -1518 0 1
rlabel polysilicon 450 -1524 450 -1524 0 3
rlabel polysilicon 457 -1518 457 -1518 0 1
rlabel polysilicon 457 -1524 457 -1524 0 3
rlabel polysilicon 464 -1518 464 -1518 0 1
rlabel polysilicon 464 -1524 464 -1524 0 3
rlabel polysilicon 471 -1518 471 -1518 0 1
rlabel polysilicon 471 -1524 471 -1524 0 3
rlabel polysilicon 478 -1518 478 -1518 0 1
rlabel polysilicon 478 -1524 478 -1524 0 3
rlabel polysilicon 485 -1518 485 -1518 0 1
rlabel polysilicon 485 -1524 485 -1524 0 3
rlabel polysilicon 492 -1518 492 -1518 0 1
rlabel polysilicon 492 -1524 492 -1524 0 3
rlabel polysilicon 502 -1518 502 -1518 0 2
rlabel polysilicon 499 -1524 499 -1524 0 3
rlabel polysilicon 502 -1524 502 -1524 0 4
rlabel polysilicon 506 -1518 506 -1518 0 1
rlabel polysilicon 506 -1524 506 -1524 0 3
rlabel polysilicon 513 -1518 513 -1518 0 1
rlabel polysilicon 513 -1524 513 -1524 0 3
rlabel polysilicon 520 -1518 520 -1518 0 1
rlabel polysilicon 520 -1524 520 -1524 0 3
rlabel polysilicon 527 -1518 527 -1518 0 1
rlabel polysilicon 527 -1524 527 -1524 0 3
rlabel polysilicon 534 -1518 534 -1518 0 1
rlabel polysilicon 534 -1524 534 -1524 0 3
rlabel polysilicon 541 -1518 541 -1518 0 1
rlabel polysilicon 541 -1524 541 -1524 0 3
rlabel polysilicon 548 -1518 548 -1518 0 1
rlabel polysilicon 548 -1524 548 -1524 0 3
rlabel polysilicon 555 -1518 555 -1518 0 1
rlabel polysilicon 555 -1524 555 -1524 0 3
rlabel polysilicon 562 -1518 562 -1518 0 1
rlabel polysilicon 562 -1524 562 -1524 0 3
rlabel polysilicon 569 -1518 569 -1518 0 1
rlabel polysilicon 569 -1524 569 -1524 0 3
rlabel polysilicon 576 -1518 576 -1518 0 1
rlabel polysilicon 576 -1524 576 -1524 0 3
rlabel polysilicon 583 -1518 583 -1518 0 1
rlabel polysilicon 583 -1524 583 -1524 0 3
rlabel polysilicon 590 -1518 590 -1518 0 1
rlabel polysilicon 590 -1524 590 -1524 0 3
rlabel polysilicon 593 -1524 593 -1524 0 4
rlabel polysilicon 597 -1518 597 -1518 0 1
rlabel polysilicon 597 -1524 597 -1524 0 3
rlabel polysilicon 604 -1518 604 -1518 0 1
rlabel polysilicon 604 -1524 604 -1524 0 3
rlabel polysilicon 611 -1518 611 -1518 0 1
rlabel polysilicon 611 -1524 611 -1524 0 3
rlabel polysilicon 618 -1518 618 -1518 0 1
rlabel polysilicon 618 -1524 618 -1524 0 3
rlabel polysilicon 625 -1518 625 -1518 0 1
rlabel polysilicon 628 -1518 628 -1518 0 2
rlabel polysilicon 625 -1524 625 -1524 0 3
rlabel polysilicon 628 -1524 628 -1524 0 4
rlabel polysilicon 632 -1518 632 -1518 0 1
rlabel polysilicon 632 -1524 632 -1524 0 3
rlabel polysilicon 639 -1518 639 -1518 0 1
rlabel polysilicon 639 -1524 639 -1524 0 3
rlabel polysilicon 646 -1518 646 -1518 0 1
rlabel polysilicon 646 -1524 646 -1524 0 3
rlabel polysilicon 653 -1518 653 -1518 0 1
rlabel polysilicon 653 -1524 653 -1524 0 3
rlabel polysilicon 660 -1518 660 -1518 0 1
rlabel polysilicon 663 -1518 663 -1518 0 2
rlabel polysilicon 660 -1524 660 -1524 0 3
rlabel polysilicon 663 -1524 663 -1524 0 4
rlabel polysilicon 667 -1518 667 -1518 0 1
rlabel polysilicon 670 -1518 670 -1518 0 2
rlabel polysilicon 667 -1524 667 -1524 0 3
rlabel polysilicon 670 -1524 670 -1524 0 4
rlabel polysilicon 674 -1518 674 -1518 0 1
rlabel polysilicon 674 -1524 674 -1524 0 3
rlabel polysilicon 681 -1518 681 -1518 0 1
rlabel polysilicon 681 -1524 681 -1524 0 3
rlabel polysilicon 688 -1518 688 -1518 0 1
rlabel polysilicon 688 -1524 688 -1524 0 3
rlabel polysilicon 695 -1518 695 -1518 0 1
rlabel polysilicon 695 -1524 695 -1524 0 3
rlabel polysilicon 702 -1518 702 -1518 0 1
rlabel polysilicon 702 -1524 702 -1524 0 3
rlabel polysilicon 709 -1518 709 -1518 0 1
rlabel polysilicon 712 -1518 712 -1518 0 2
rlabel polysilicon 709 -1524 709 -1524 0 3
rlabel polysilicon 712 -1524 712 -1524 0 4
rlabel polysilicon 716 -1518 716 -1518 0 1
rlabel polysilicon 716 -1524 716 -1524 0 3
rlabel polysilicon 723 -1518 723 -1518 0 1
rlabel polysilicon 723 -1524 723 -1524 0 3
rlabel polysilicon 730 -1518 730 -1518 0 1
rlabel polysilicon 730 -1524 730 -1524 0 3
rlabel polysilicon 737 -1518 737 -1518 0 1
rlabel polysilicon 737 -1524 737 -1524 0 3
rlabel polysilicon 744 -1518 744 -1518 0 1
rlabel polysilicon 744 -1524 744 -1524 0 3
rlabel polysilicon 751 -1518 751 -1518 0 1
rlabel polysilicon 754 -1518 754 -1518 0 2
rlabel polysilicon 751 -1524 751 -1524 0 3
rlabel polysilicon 754 -1524 754 -1524 0 4
rlabel polysilicon 758 -1518 758 -1518 0 1
rlabel polysilicon 758 -1524 758 -1524 0 3
rlabel polysilicon 765 -1518 765 -1518 0 1
rlabel polysilicon 765 -1524 765 -1524 0 3
rlabel polysilicon 772 -1518 772 -1518 0 1
rlabel polysilicon 772 -1524 772 -1524 0 3
rlabel polysilicon 779 -1518 779 -1518 0 1
rlabel polysilicon 779 -1524 779 -1524 0 3
rlabel polysilicon 786 -1518 786 -1518 0 1
rlabel polysilicon 786 -1524 786 -1524 0 3
rlabel polysilicon 793 -1518 793 -1518 0 1
rlabel polysilicon 793 -1524 793 -1524 0 3
rlabel polysilicon 800 -1518 800 -1518 0 1
rlabel polysilicon 800 -1524 800 -1524 0 3
rlabel polysilicon 807 -1518 807 -1518 0 1
rlabel polysilicon 807 -1524 807 -1524 0 3
rlabel polysilicon 814 -1518 814 -1518 0 1
rlabel polysilicon 814 -1524 814 -1524 0 3
rlabel polysilicon 821 -1518 821 -1518 0 1
rlabel polysilicon 821 -1524 821 -1524 0 3
rlabel polysilicon 828 -1518 828 -1518 0 1
rlabel polysilicon 828 -1524 828 -1524 0 3
rlabel polysilicon 835 -1518 835 -1518 0 1
rlabel polysilicon 835 -1524 835 -1524 0 3
rlabel polysilicon 842 -1518 842 -1518 0 1
rlabel polysilicon 842 -1524 842 -1524 0 3
rlabel polysilicon 849 -1518 849 -1518 0 1
rlabel polysilicon 849 -1524 849 -1524 0 3
rlabel polysilicon 856 -1518 856 -1518 0 1
rlabel polysilicon 856 -1524 856 -1524 0 3
rlabel polysilicon 863 -1518 863 -1518 0 1
rlabel polysilicon 863 -1524 863 -1524 0 3
rlabel polysilicon 870 -1518 870 -1518 0 1
rlabel polysilicon 870 -1524 870 -1524 0 3
rlabel polysilicon 877 -1518 877 -1518 0 1
rlabel polysilicon 877 -1524 877 -1524 0 3
rlabel polysilicon 884 -1518 884 -1518 0 1
rlabel polysilicon 884 -1524 884 -1524 0 3
rlabel polysilicon 891 -1518 891 -1518 0 1
rlabel polysilicon 891 -1524 891 -1524 0 3
rlabel polysilicon 898 -1518 898 -1518 0 1
rlabel polysilicon 898 -1524 898 -1524 0 3
rlabel polysilicon 905 -1518 905 -1518 0 1
rlabel polysilicon 905 -1524 905 -1524 0 3
rlabel polysilicon 912 -1518 912 -1518 0 1
rlabel polysilicon 912 -1524 912 -1524 0 3
rlabel polysilicon 922 -1518 922 -1518 0 2
rlabel polysilicon 919 -1524 919 -1524 0 3
rlabel polysilicon 922 -1524 922 -1524 0 4
rlabel polysilicon 926 -1518 926 -1518 0 1
rlabel polysilicon 926 -1524 926 -1524 0 3
rlabel polysilicon 933 -1518 933 -1518 0 1
rlabel polysilicon 933 -1524 933 -1524 0 3
rlabel polysilicon 940 -1518 940 -1518 0 1
rlabel polysilicon 940 -1524 940 -1524 0 3
rlabel polysilicon 947 -1518 947 -1518 0 1
rlabel polysilicon 950 -1518 950 -1518 0 2
rlabel polysilicon 950 -1524 950 -1524 0 4
rlabel polysilicon 954 -1518 954 -1518 0 1
rlabel polysilicon 957 -1518 957 -1518 0 2
rlabel polysilicon 954 -1524 954 -1524 0 3
rlabel polysilicon 957 -1524 957 -1524 0 4
rlabel polysilicon 961 -1518 961 -1518 0 1
rlabel polysilicon 968 -1518 968 -1518 0 1
rlabel polysilicon 968 -1524 968 -1524 0 3
rlabel polysilicon 975 -1518 975 -1518 0 1
rlabel polysilicon 975 -1524 975 -1524 0 3
rlabel polysilicon 982 -1518 982 -1518 0 1
rlabel polysilicon 985 -1518 985 -1518 0 2
rlabel polysilicon 982 -1524 982 -1524 0 3
rlabel polysilicon 985 -1524 985 -1524 0 4
rlabel polysilicon 989 -1518 989 -1518 0 1
rlabel polysilicon 989 -1524 989 -1524 0 3
rlabel polysilicon 996 -1518 996 -1518 0 1
rlabel polysilicon 996 -1524 996 -1524 0 3
rlabel polysilicon 1003 -1518 1003 -1518 0 1
rlabel polysilicon 1006 -1518 1006 -1518 0 2
rlabel polysilicon 1003 -1524 1003 -1524 0 3
rlabel polysilicon 1006 -1524 1006 -1524 0 4
rlabel polysilicon 1010 -1518 1010 -1518 0 1
rlabel polysilicon 1010 -1524 1010 -1524 0 3
rlabel polysilicon 1017 -1518 1017 -1518 0 1
rlabel polysilicon 1017 -1524 1017 -1524 0 3
rlabel polysilicon 1024 -1518 1024 -1518 0 1
rlabel polysilicon 1024 -1524 1024 -1524 0 3
rlabel polysilicon 1031 -1518 1031 -1518 0 1
rlabel polysilicon 1031 -1524 1031 -1524 0 3
rlabel polysilicon 1038 -1518 1038 -1518 0 1
rlabel polysilicon 1038 -1524 1038 -1524 0 3
rlabel polysilicon 1045 -1524 1045 -1524 0 3
rlabel polysilicon 1052 -1518 1052 -1518 0 1
rlabel polysilicon 1052 -1524 1052 -1524 0 3
rlabel polysilicon 1059 -1518 1059 -1518 0 1
rlabel polysilicon 1059 -1524 1059 -1524 0 3
rlabel polysilicon 1069 -1518 1069 -1518 0 2
rlabel polysilicon 1066 -1524 1066 -1524 0 3
rlabel polysilicon 1069 -1524 1069 -1524 0 4
rlabel polysilicon 1073 -1518 1073 -1518 0 1
rlabel polysilicon 1073 -1524 1073 -1524 0 3
rlabel polysilicon 1080 -1518 1080 -1518 0 1
rlabel polysilicon 1080 -1524 1080 -1524 0 3
rlabel polysilicon 1087 -1518 1087 -1518 0 1
rlabel polysilicon 1087 -1524 1087 -1524 0 3
rlabel polysilicon 1094 -1518 1094 -1518 0 1
rlabel polysilicon 1094 -1524 1094 -1524 0 3
rlabel polysilicon 1101 -1518 1101 -1518 0 1
rlabel polysilicon 1104 -1518 1104 -1518 0 2
rlabel polysilicon 1101 -1524 1101 -1524 0 3
rlabel polysilicon 1104 -1524 1104 -1524 0 4
rlabel polysilicon 1108 -1518 1108 -1518 0 1
rlabel polysilicon 1111 -1518 1111 -1518 0 2
rlabel polysilicon 1108 -1524 1108 -1524 0 3
rlabel polysilicon 1111 -1524 1111 -1524 0 4
rlabel polysilicon 1115 -1518 1115 -1518 0 1
rlabel polysilicon 1118 -1518 1118 -1518 0 2
rlabel polysilicon 1115 -1524 1115 -1524 0 3
rlabel polysilicon 1118 -1524 1118 -1524 0 4
rlabel polysilicon 1122 -1518 1122 -1518 0 1
rlabel polysilicon 1122 -1524 1122 -1524 0 3
rlabel polysilicon 1129 -1518 1129 -1518 0 1
rlabel polysilicon 1132 -1518 1132 -1518 0 2
rlabel polysilicon 1129 -1524 1129 -1524 0 3
rlabel polysilicon 1132 -1524 1132 -1524 0 4
rlabel polysilicon 1136 -1518 1136 -1518 0 1
rlabel polysilicon 1136 -1524 1136 -1524 0 3
rlabel polysilicon 1143 -1518 1143 -1518 0 1
rlabel polysilicon 1143 -1524 1143 -1524 0 3
rlabel polysilicon 1150 -1518 1150 -1518 0 1
rlabel polysilicon 1150 -1524 1150 -1524 0 3
rlabel polysilicon 1157 -1518 1157 -1518 0 1
rlabel polysilicon 1160 -1518 1160 -1518 0 2
rlabel polysilicon 1157 -1524 1157 -1524 0 3
rlabel polysilicon 1160 -1524 1160 -1524 0 4
rlabel polysilicon 1164 -1518 1164 -1518 0 1
rlabel polysilicon 1164 -1524 1164 -1524 0 3
rlabel polysilicon 1171 -1518 1171 -1518 0 1
rlabel polysilicon 1171 -1524 1171 -1524 0 3
rlabel polysilicon 1178 -1518 1178 -1518 0 1
rlabel polysilicon 1178 -1524 1178 -1524 0 3
rlabel polysilicon 1185 -1518 1185 -1518 0 1
rlabel polysilicon 1185 -1524 1185 -1524 0 3
rlabel polysilicon 1192 -1518 1192 -1518 0 1
rlabel polysilicon 1192 -1524 1192 -1524 0 3
rlabel polysilicon 1195 -1524 1195 -1524 0 4
rlabel polysilicon 1199 -1518 1199 -1518 0 1
rlabel polysilicon 1199 -1524 1199 -1524 0 3
rlabel polysilicon 1206 -1518 1206 -1518 0 1
rlabel polysilicon 1206 -1524 1206 -1524 0 3
rlabel polysilicon 1213 -1518 1213 -1518 0 1
rlabel polysilicon 1213 -1524 1213 -1524 0 3
rlabel polysilicon 1220 -1518 1220 -1518 0 1
rlabel polysilicon 1220 -1524 1220 -1524 0 3
rlabel polysilicon 1227 -1518 1227 -1518 0 1
rlabel polysilicon 1227 -1524 1227 -1524 0 3
rlabel polysilicon 1234 -1518 1234 -1518 0 1
rlabel polysilicon 1234 -1524 1234 -1524 0 3
rlabel polysilicon 1241 -1518 1241 -1518 0 1
rlabel polysilicon 1241 -1524 1241 -1524 0 3
rlabel polysilicon 1248 -1518 1248 -1518 0 1
rlabel polysilicon 1248 -1524 1248 -1524 0 3
rlabel polysilicon 1255 -1518 1255 -1518 0 1
rlabel polysilicon 1255 -1524 1255 -1524 0 3
rlabel polysilicon 1262 -1518 1262 -1518 0 1
rlabel polysilicon 1265 -1518 1265 -1518 0 2
rlabel polysilicon 1262 -1524 1262 -1524 0 3
rlabel polysilicon 1265 -1524 1265 -1524 0 4
rlabel polysilicon 1269 -1518 1269 -1518 0 1
rlabel polysilicon 1269 -1524 1269 -1524 0 3
rlabel polysilicon 1276 -1518 1276 -1518 0 1
rlabel polysilicon 1276 -1524 1276 -1524 0 3
rlabel polysilicon 1283 -1518 1283 -1518 0 1
rlabel polysilicon 1283 -1524 1283 -1524 0 3
rlabel polysilicon 1290 -1518 1290 -1518 0 1
rlabel polysilicon 1290 -1524 1290 -1524 0 3
rlabel polysilicon 1297 -1518 1297 -1518 0 1
rlabel polysilicon 1297 -1524 1297 -1524 0 3
rlabel polysilicon 1304 -1518 1304 -1518 0 1
rlabel polysilicon 1307 -1518 1307 -1518 0 2
rlabel polysilicon 1307 -1524 1307 -1524 0 4
rlabel polysilicon 1311 -1518 1311 -1518 0 1
rlabel polysilicon 1311 -1524 1311 -1524 0 3
rlabel polysilicon 1318 -1518 1318 -1518 0 1
rlabel polysilicon 1318 -1524 1318 -1524 0 3
rlabel polysilicon 1325 -1518 1325 -1518 0 1
rlabel polysilicon 1325 -1524 1325 -1524 0 3
rlabel polysilicon 1332 -1518 1332 -1518 0 1
rlabel polysilicon 1335 -1518 1335 -1518 0 2
rlabel polysilicon 1332 -1524 1332 -1524 0 3
rlabel polysilicon 1335 -1524 1335 -1524 0 4
rlabel polysilicon 1339 -1518 1339 -1518 0 1
rlabel polysilicon 1339 -1524 1339 -1524 0 3
rlabel polysilicon 1346 -1518 1346 -1518 0 1
rlabel polysilicon 1346 -1524 1346 -1524 0 3
rlabel polysilicon 1353 -1518 1353 -1518 0 1
rlabel polysilicon 1353 -1524 1353 -1524 0 3
rlabel polysilicon 1360 -1518 1360 -1518 0 1
rlabel polysilicon 1360 -1524 1360 -1524 0 3
rlabel polysilicon 1367 -1518 1367 -1518 0 1
rlabel polysilicon 1367 -1524 1367 -1524 0 3
rlabel polysilicon 1374 -1518 1374 -1518 0 1
rlabel polysilicon 1374 -1524 1374 -1524 0 3
rlabel polysilicon 1381 -1518 1381 -1518 0 1
rlabel polysilicon 1381 -1524 1381 -1524 0 3
rlabel polysilicon 1388 -1518 1388 -1518 0 1
rlabel polysilicon 1388 -1524 1388 -1524 0 3
rlabel polysilicon 1395 -1518 1395 -1518 0 1
rlabel polysilicon 1395 -1524 1395 -1524 0 3
rlabel polysilicon 1402 -1518 1402 -1518 0 1
rlabel polysilicon 1402 -1524 1402 -1524 0 3
rlabel polysilicon 1409 -1518 1409 -1518 0 1
rlabel polysilicon 1409 -1524 1409 -1524 0 3
rlabel polysilicon 1416 -1518 1416 -1518 0 1
rlabel polysilicon 1416 -1524 1416 -1524 0 3
rlabel polysilicon 1423 -1518 1423 -1518 0 1
rlabel polysilicon 1423 -1524 1423 -1524 0 3
rlabel polysilicon 1430 -1518 1430 -1518 0 1
rlabel polysilicon 1430 -1524 1430 -1524 0 3
rlabel polysilicon 1437 -1518 1437 -1518 0 1
rlabel polysilicon 1437 -1524 1437 -1524 0 3
rlabel polysilicon 1444 -1518 1444 -1518 0 1
rlabel polysilicon 1444 -1524 1444 -1524 0 3
rlabel polysilicon 1451 -1518 1451 -1518 0 1
rlabel polysilicon 1451 -1524 1451 -1524 0 3
rlabel polysilicon 1458 -1518 1458 -1518 0 1
rlabel polysilicon 1458 -1524 1458 -1524 0 3
rlabel polysilicon 1465 -1518 1465 -1518 0 1
rlabel polysilicon 1465 -1524 1465 -1524 0 3
rlabel polysilicon 1472 -1518 1472 -1518 0 1
rlabel polysilicon 1472 -1524 1472 -1524 0 3
rlabel polysilicon 1479 -1518 1479 -1518 0 1
rlabel polysilicon 1479 -1524 1479 -1524 0 3
rlabel polysilicon 1486 -1518 1486 -1518 0 1
rlabel polysilicon 1486 -1524 1486 -1524 0 3
rlabel polysilicon 1493 -1518 1493 -1518 0 1
rlabel polysilicon 1493 -1524 1493 -1524 0 3
rlabel polysilicon 1500 -1518 1500 -1518 0 1
rlabel polysilicon 1500 -1524 1500 -1524 0 3
rlabel polysilicon 1507 -1518 1507 -1518 0 1
rlabel polysilicon 1507 -1524 1507 -1524 0 3
rlabel polysilicon 1514 -1518 1514 -1518 0 1
rlabel polysilicon 1514 -1524 1514 -1524 0 3
rlabel polysilicon 1521 -1518 1521 -1518 0 1
rlabel polysilicon 1521 -1524 1521 -1524 0 3
rlabel polysilicon 1528 -1518 1528 -1518 0 1
rlabel polysilicon 1528 -1524 1528 -1524 0 3
rlabel polysilicon 1535 -1518 1535 -1518 0 1
rlabel polysilicon 1535 -1524 1535 -1524 0 3
rlabel polysilicon 1542 -1518 1542 -1518 0 1
rlabel polysilicon 1542 -1524 1542 -1524 0 3
rlabel polysilicon 1549 -1518 1549 -1518 0 1
rlabel polysilicon 1549 -1524 1549 -1524 0 3
rlabel polysilicon 1556 -1518 1556 -1518 0 1
rlabel polysilicon 1556 -1524 1556 -1524 0 3
rlabel polysilicon 1563 -1518 1563 -1518 0 1
rlabel polysilicon 1563 -1524 1563 -1524 0 3
rlabel polysilicon 1570 -1518 1570 -1518 0 1
rlabel polysilicon 1570 -1524 1570 -1524 0 3
rlabel polysilicon 1577 -1518 1577 -1518 0 1
rlabel polysilicon 1577 -1524 1577 -1524 0 3
rlabel polysilicon 1584 -1518 1584 -1518 0 1
rlabel polysilicon 1584 -1524 1584 -1524 0 3
rlabel polysilicon 1591 -1518 1591 -1518 0 1
rlabel polysilicon 1591 -1524 1591 -1524 0 3
rlabel polysilicon 1598 -1518 1598 -1518 0 1
rlabel polysilicon 1598 -1524 1598 -1524 0 3
rlabel polysilicon 1605 -1518 1605 -1518 0 1
rlabel polysilicon 1605 -1524 1605 -1524 0 3
rlabel polysilicon 1612 -1518 1612 -1518 0 1
rlabel polysilicon 1612 -1524 1612 -1524 0 3
rlabel polysilicon 1619 -1518 1619 -1518 0 1
rlabel polysilicon 1619 -1524 1619 -1524 0 3
rlabel polysilicon 1626 -1518 1626 -1518 0 1
rlabel polysilicon 1626 -1524 1626 -1524 0 3
rlabel polysilicon 1633 -1518 1633 -1518 0 1
rlabel polysilicon 1633 -1524 1633 -1524 0 3
rlabel polysilicon 1640 -1518 1640 -1518 0 1
rlabel polysilicon 1640 -1524 1640 -1524 0 3
rlabel polysilicon 1647 -1518 1647 -1518 0 1
rlabel polysilicon 1647 -1524 1647 -1524 0 3
rlabel polysilicon 1654 -1518 1654 -1518 0 1
rlabel polysilicon 1654 -1524 1654 -1524 0 3
rlabel polysilicon 1661 -1518 1661 -1518 0 1
rlabel polysilicon 1661 -1524 1661 -1524 0 3
rlabel polysilicon 1668 -1518 1668 -1518 0 1
rlabel polysilicon 1668 -1524 1668 -1524 0 3
rlabel polysilicon 1675 -1518 1675 -1518 0 1
rlabel polysilicon 1675 -1524 1675 -1524 0 3
rlabel polysilicon 1682 -1518 1682 -1518 0 1
rlabel polysilicon 1682 -1524 1682 -1524 0 3
rlabel polysilicon 1689 -1518 1689 -1518 0 1
rlabel polysilicon 1689 -1524 1689 -1524 0 3
rlabel polysilicon 1696 -1518 1696 -1518 0 1
rlabel polysilicon 1696 -1524 1696 -1524 0 3
rlabel polysilicon 1703 -1518 1703 -1518 0 1
rlabel polysilicon 1703 -1524 1703 -1524 0 3
rlabel polysilicon 1710 -1518 1710 -1518 0 1
rlabel polysilicon 1710 -1524 1710 -1524 0 3
rlabel polysilicon 1717 -1518 1717 -1518 0 1
rlabel polysilicon 1717 -1524 1717 -1524 0 3
rlabel polysilicon 1724 -1518 1724 -1518 0 1
rlabel polysilicon 1724 -1524 1724 -1524 0 3
rlabel polysilicon 1731 -1518 1731 -1518 0 1
rlabel polysilicon 1731 -1524 1731 -1524 0 3
rlabel polysilicon 1738 -1518 1738 -1518 0 1
rlabel polysilicon 1738 -1524 1738 -1524 0 3
rlabel polysilicon 1745 -1518 1745 -1518 0 1
rlabel polysilicon 1745 -1524 1745 -1524 0 3
rlabel polysilicon 1752 -1518 1752 -1518 0 1
rlabel polysilicon 1752 -1524 1752 -1524 0 3
rlabel polysilicon 1759 -1518 1759 -1518 0 1
rlabel polysilicon 1759 -1524 1759 -1524 0 3
rlabel polysilicon 1766 -1518 1766 -1518 0 1
rlabel polysilicon 1766 -1524 1766 -1524 0 3
rlabel polysilicon 1773 -1518 1773 -1518 0 1
rlabel polysilicon 1773 -1524 1773 -1524 0 3
rlabel polysilicon 1780 -1518 1780 -1518 0 1
rlabel polysilicon 1780 -1524 1780 -1524 0 3
rlabel polysilicon 1787 -1518 1787 -1518 0 1
rlabel polysilicon 1787 -1524 1787 -1524 0 3
rlabel polysilicon 1794 -1518 1794 -1518 0 1
rlabel polysilicon 1794 -1524 1794 -1524 0 3
rlabel polysilicon 1801 -1518 1801 -1518 0 1
rlabel polysilicon 1801 -1524 1801 -1524 0 3
rlabel polysilicon 1808 -1518 1808 -1518 0 1
rlabel polysilicon 1808 -1524 1808 -1524 0 3
rlabel polysilicon 1815 -1518 1815 -1518 0 1
rlabel polysilicon 1815 -1524 1815 -1524 0 3
rlabel polysilicon 1822 -1518 1822 -1518 0 1
rlabel polysilicon 1822 -1524 1822 -1524 0 3
rlabel polysilicon 1829 -1518 1829 -1518 0 1
rlabel polysilicon 1829 -1524 1829 -1524 0 3
rlabel polysilicon 1836 -1518 1836 -1518 0 1
rlabel polysilicon 1836 -1524 1836 -1524 0 3
rlabel polysilicon 1843 -1518 1843 -1518 0 1
rlabel polysilicon 1843 -1524 1843 -1524 0 3
rlabel polysilicon 1850 -1518 1850 -1518 0 1
rlabel polysilicon 1850 -1524 1850 -1524 0 3
rlabel polysilicon 1857 -1518 1857 -1518 0 1
rlabel polysilicon 1857 -1524 1857 -1524 0 3
rlabel polysilicon 1864 -1518 1864 -1518 0 1
rlabel polysilicon 1864 -1524 1864 -1524 0 3
rlabel polysilicon 1871 -1518 1871 -1518 0 1
rlabel polysilicon 1871 -1524 1871 -1524 0 3
rlabel polysilicon 1878 -1518 1878 -1518 0 1
rlabel polysilicon 1878 -1524 1878 -1524 0 3
rlabel polysilicon 1885 -1518 1885 -1518 0 1
rlabel polysilicon 1885 -1524 1885 -1524 0 3
rlabel polysilicon 1892 -1518 1892 -1518 0 1
rlabel polysilicon 1892 -1524 1892 -1524 0 3
rlabel polysilicon 1899 -1518 1899 -1518 0 1
rlabel polysilicon 1899 -1524 1899 -1524 0 3
rlabel polysilicon 1906 -1518 1906 -1518 0 1
rlabel polysilicon 1906 -1524 1906 -1524 0 3
rlabel polysilicon 1913 -1518 1913 -1518 0 1
rlabel polysilicon 1913 -1524 1913 -1524 0 3
rlabel polysilicon 1920 -1518 1920 -1518 0 1
rlabel polysilicon 1920 -1524 1920 -1524 0 3
rlabel polysilicon 1927 -1518 1927 -1518 0 1
rlabel polysilicon 1927 -1524 1927 -1524 0 3
rlabel polysilicon 1934 -1518 1934 -1518 0 1
rlabel polysilicon 1934 -1524 1934 -1524 0 3
rlabel polysilicon 1941 -1518 1941 -1518 0 1
rlabel polysilicon 1941 -1524 1941 -1524 0 3
rlabel polysilicon 1948 -1518 1948 -1518 0 1
rlabel polysilicon 1948 -1524 1948 -1524 0 3
rlabel polysilicon 1955 -1518 1955 -1518 0 1
rlabel polysilicon 1955 -1524 1955 -1524 0 3
rlabel polysilicon 1962 -1518 1962 -1518 0 1
rlabel polysilicon 1962 -1524 1962 -1524 0 3
rlabel polysilicon 1969 -1518 1969 -1518 0 1
rlabel polysilicon 1969 -1524 1969 -1524 0 3
rlabel polysilicon 1972 -1524 1972 -1524 0 4
rlabel polysilicon 1976 -1524 1976 -1524 0 3
rlabel polysilicon 1979 -1524 1979 -1524 0 4
rlabel polysilicon 1983 -1518 1983 -1518 0 1
rlabel polysilicon 1986 -1518 1986 -1518 0 2
rlabel polysilicon 1983 -1524 1983 -1524 0 3
rlabel polysilicon 1990 -1518 1990 -1518 0 1
rlabel polysilicon 1990 -1524 1990 -1524 0 3
rlabel polysilicon 1997 -1518 1997 -1518 0 1
rlabel polysilicon 2000 -1524 2000 -1524 0 4
rlabel polysilicon 2007 -1518 2007 -1518 0 2
rlabel polysilicon 2004 -1524 2004 -1524 0 3
rlabel polysilicon 2007 -1524 2007 -1524 0 4
rlabel polysilicon 2011 -1518 2011 -1518 0 1
rlabel polysilicon 2011 -1524 2011 -1524 0 3
rlabel polysilicon 2018 -1518 2018 -1518 0 1
rlabel polysilicon 2018 -1524 2018 -1524 0 3
rlabel polysilicon 2025 -1518 2025 -1518 0 1
rlabel polysilicon 2025 -1524 2025 -1524 0 3
rlabel polysilicon 2 -1645 2 -1645 0 1
rlabel polysilicon 2 -1651 2 -1651 0 3
rlabel polysilicon 9 -1645 9 -1645 0 1
rlabel polysilicon 9 -1651 9 -1651 0 3
rlabel polysilicon 16 -1645 16 -1645 0 1
rlabel polysilicon 16 -1651 16 -1651 0 3
rlabel polysilicon 23 -1645 23 -1645 0 1
rlabel polysilicon 23 -1651 23 -1651 0 3
rlabel polysilicon 30 -1645 30 -1645 0 1
rlabel polysilicon 30 -1651 30 -1651 0 3
rlabel polysilicon 37 -1645 37 -1645 0 1
rlabel polysilicon 37 -1651 37 -1651 0 3
rlabel polysilicon 44 -1645 44 -1645 0 1
rlabel polysilicon 44 -1651 44 -1651 0 3
rlabel polysilicon 51 -1645 51 -1645 0 1
rlabel polysilicon 51 -1651 51 -1651 0 3
rlabel polysilicon 58 -1645 58 -1645 0 1
rlabel polysilicon 58 -1651 58 -1651 0 3
rlabel polysilicon 65 -1645 65 -1645 0 1
rlabel polysilicon 68 -1645 68 -1645 0 2
rlabel polysilicon 65 -1651 65 -1651 0 3
rlabel polysilicon 72 -1645 72 -1645 0 1
rlabel polysilicon 72 -1651 72 -1651 0 3
rlabel polysilicon 79 -1645 79 -1645 0 1
rlabel polysilicon 82 -1645 82 -1645 0 2
rlabel polysilicon 82 -1651 82 -1651 0 4
rlabel polysilicon 86 -1645 86 -1645 0 1
rlabel polysilicon 89 -1645 89 -1645 0 2
rlabel polysilicon 89 -1651 89 -1651 0 4
rlabel polysilicon 93 -1645 93 -1645 0 1
rlabel polysilicon 93 -1651 93 -1651 0 3
rlabel polysilicon 100 -1645 100 -1645 0 1
rlabel polysilicon 100 -1651 100 -1651 0 3
rlabel polysilicon 107 -1645 107 -1645 0 1
rlabel polysilicon 107 -1651 107 -1651 0 3
rlabel polysilicon 114 -1645 114 -1645 0 1
rlabel polysilicon 117 -1645 117 -1645 0 2
rlabel polysilicon 114 -1651 114 -1651 0 3
rlabel polysilicon 117 -1651 117 -1651 0 4
rlabel polysilicon 121 -1645 121 -1645 0 1
rlabel polysilicon 121 -1651 121 -1651 0 3
rlabel polysilicon 128 -1645 128 -1645 0 1
rlabel polysilicon 128 -1651 128 -1651 0 3
rlabel polysilicon 135 -1645 135 -1645 0 1
rlabel polysilicon 135 -1651 135 -1651 0 3
rlabel polysilicon 142 -1645 142 -1645 0 1
rlabel polysilicon 145 -1645 145 -1645 0 2
rlabel polysilicon 142 -1651 142 -1651 0 3
rlabel polysilicon 149 -1645 149 -1645 0 1
rlabel polysilicon 149 -1651 149 -1651 0 3
rlabel polysilicon 156 -1645 156 -1645 0 1
rlabel polysilicon 156 -1651 156 -1651 0 3
rlabel polysilicon 163 -1645 163 -1645 0 1
rlabel polysilicon 163 -1651 163 -1651 0 3
rlabel polysilicon 170 -1645 170 -1645 0 1
rlabel polysilicon 173 -1645 173 -1645 0 2
rlabel polysilicon 170 -1651 170 -1651 0 3
rlabel polysilicon 177 -1645 177 -1645 0 1
rlabel polysilicon 180 -1645 180 -1645 0 2
rlabel polysilicon 180 -1651 180 -1651 0 4
rlabel polysilicon 184 -1645 184 -1645 0 1
rlabel polysilicon 184 -1651 184 -1651 0 3
rlabel polysilicon 191 -1645 191 -1645 0 1
rlabel polysilicon 191 -1651 191 -1651 0 3
rlabel polysilicon 198 -1645 198 -1645 0 1
rlabel polysilicon 198 -1651 198 -1651 0 3
rlabel polysilicon 205 -1645 205 -1645 0 1
rlabel polysilicon 205 -1651 205 -1651 0 3
rlabel polysilicon 212 -1645 212 -1645 0 1
rlabel polysilicon 212 -1651 212 -1651 0 3
rlabel polysilicon 219 -1645 219 -1645 0 1
rlabel polysilicon 219 -1651 219 -1651 0 3
rlabel polysilicon 226 -1645 226 -1645 0 1
rlabel polysilicon 226 -1651 226 -1651 0 3
rlabel polysilicon 233 -1645 233 -1645 0 1
rlabel polysilicon 233 -1651 233 -1651 0 3
rlabel polysilicon 240 -1645 240 -1645 0 1
rlabel polysilicon 240 -1651 240 -1651 0 3
rlabel polysilicon 247 -1645 247 -1645 0 1
rlabel polysilicon 247 -1651 247 -1651 0 3
rlabel polysilicon 254 -1645 254 -1645 0 1
rlabel polysilicon 254 -1651 254 -1651 0 3
rlabel polysilicon 261 -1645 261 -1645 0 1
rlabel polysilicon 261 -1651 261 -1651 0 3
rlabel polysilicon 268 -1645 268 -1645 0 1
rlabel polysilicon 268 -1651 268 -1651 0 3
rlabel polysilicon 275 -1645 275 -1645 0 1
rlabel polysilicon 275 -1651 275 -1651 0 3
rlabel polysilicon 282 -1645 282 -1645 0 1
rlabel polysilicon 282 -1651 282 -1651 0 3
rlabel polysilicon 289 -1645 289 -1645 0 1
rlabel polysilicon 289 -1651 289 -1651 0 3
rlabel polysilicon 296 -1645 296 -1645 0 1
rlabel polysilicon 296 -1651 296 -1651 0 3
rlabel polysilicon 303 -1645 303 -1645 0 1
rlabel polysilicon 303 -1651 303 -1651 0 3
rlabel polysilicon 310 -1645 310 -1645 0 1
rlabel polysilicon 310 -1651 310 -1651 0 3
rlabel polysilicon 317 -1645 317 -1645 0 1
rlabel polysilicon 317 -1651 317 -1651 0 3
rlabel polysilicon 324 -1645 324 -1645 0 1
rlabel polysilicon 324 -1651 324 -1651 0 3
rlabel polysilicon 331 -1645 331 -1645 0 1
rlabel polysilicon 331 -1651 331 -1651 0 3
rlabel polysilicon 338 -1645 338 -1645 0 1
rlabel polysilicon 338 -1651 338 -1651 0 3
rlabel polysilicon 345 -1645 345 -1645 0 1
rlabel polysilicon 345 -1651 345 -1651 0 3
rlabel polysilicon 352 -1645 352 -1645 0 1
rlabel polysilicon 352 -1651 352 -1651 0 3
rlabel polysilicon 359 -1645 359 -1645 0 1
rlabel polysilicon 359 -1651 359 -1651 0 3
rlabel polysilicon 366 -1645 366 -1645 0 1
rlabel polysilicon 366 -1651 366 -1651 0 3
rlabel polysilicon 373 -1645 373 -1645 0 1
rlabel polysilicon 373 -1651 373 -1651 0 3
rlabel polysilicon 380 -1645 380 -1645 0 1
rlabel polysilicon 380 -1651 380 -1651 0 3
rlabel polysilicon 387 -1645 387 -1645 0 1
rlabel polysilicon 387 -1651 387 -1651 0 3
rlabel polysilicon 394 -1645 394 -1645 0 1
rlabel polysilicon 397 -1645 397 -1645 0 2
rlabel polysilicon 394 -1651 394 -1651 0 3
rlabel polysilicon 397 -1651 397 -1651 0 4
rlabel polysilicon 401 -1645 401 -1645 0 1
rlabel polysilicon 401 -1651 401 -1651 0 3
rlabel polysilicon 408 -1645 408 -1645 0 1
rlabel polysilicon 408 -1651 408 -1651 0 3
rlabel polysilicon 418 -1645 418 -1645 0 2
rlabel polysilicon 418 -1651 418 -1651 0 4
rlabel polysilicon 422 -1645 422 -1645 0 1
rlabel polysilicon 422 -1651 422 -1651 0 3
rlabel polysilicon 429 -1645 429 -1645 0 1
rlabel polysilicon 429 -1651 429 -1651 0 3
rlabel polysilicon 436 -1645 436 -1645 0 1
rlabel polysilicon 436 -1651 436 -1651 0 3
rlabel polysilicon 443 -1645 443 -1645 0 1
rlabel polysilicon 443 -1651 443 -1651 0 3
rlabel polysilicon 450 -1645 450 -1645 0 1
rlabel polysilicon 450 -1651 450 -1651 0 3
rlabel polysilicon 457 -1645 457 -1645 0 1
rlabel polysilicon 457 -1651 457 -1651 0 3
rlabel polysilicon 464 -1645 464 -1645 0 1
rlabel polysilicon 464 -1651 464 -1651 0 3
rlabel polysilicon 471 -1645 471 -1645 0 1
rlabel polysilicon 471 -1651 471 -1651 0 3
rlabel polysilicon 478 -1645 478 -1645 0 1
rlabel polysilicon 478 -1651 478 -1651 0 3
rlabel polysilicon 485 -1645 485 -1645 0 1
rlabel polysilicon 485 -1651 485 -1651 0 3
rlabel polysilicon 492 -1645 492 -1645 0 1
rlabel polysilicon 492 -1651 492 -1651 0 3
rlabel polysilicon 499 -1645 499 -1645 0 1
rlabel polysilicon 499 -1651 499 -1651 0 3
rlabel polysilicon 506 -1645 506 -1645 0 1
rlabel polysilicon 506 -1651 506 -1651 0 3
rlabel polysilicon 513 -1645 513 -1645 0 1
rlabel polysilicon 513 -1651 513 -1651 0 3
rlabel polysilicon 520 -1645 520 -1645 0 1
rlabel polysilicon 520 -1651 520 -1651 0 3
rlabel polysilicon 527 -1645 527 -1645 0 1
rlabel polysilicon 527 -1651 527 -1651 0 3
rlabel polysilicon 534 -1645 534 -1645 0 1
rlabel polysilicon 534 -1651 534 -1651 0 3
rlabel polysilicon 541 -1645 541 -1645 0 1
rlabel polysilicon 544 -1645 544 -1645 0 2
rlabel polysilicon 541 -1651 541 -1651 0 3
rlabel polysilicon 544 -1651 544 -1651 0 4
rlabel polysilicon 548 -1645 548 -1645 0 1
rlabel polysilicon 548 -1651 548 -1651 0 3
rlabel polysilicon 555 -1645 555 -1645 0 1
rlabel polysilicon 555 -1651 555 -1651 0 3
rlabel polysilicon 562 -1645 562 -1645 0 1
rlabel polysilicon 562 -1651 562 -1651 0 3
rlabel polysilicon 569 -1645 569 -1645 0 1
rlabel polysilicon 569 -1651 569 -1651 0 3
rlabel polysilicon 576 -1645 576 -1645 0 1
rlabel polysilicon 576 -1651 576 -1651 0 3
rlabel polysilicon 583 -1645 583 -1645 0 1
rlabel polysilicon 583 -1651 583 -1651 0 3
rlabel polysilicon 590 -1645 590 -1645 0 1
rlabel polysilicon 590 -1651 590 -1651 0 3
rlabel polysilicon 597 -1645 597 -1645 0 1
rlabel polysilicon 597 -1651 597 -1651 0 3
rlabel polysilicon 604 -1645 604 -1645 0 1
rlabel polysilicon 604 -1651 604 -1651 0 3
rlabel polysilicon 611 -1645 611 -1645 0 1
rlabel polysilicon 611 -1651 611 -1651 0 3
rlabel polysilicon 618 -1645 618 -1645 0 1
rlabel polysilicon 618 -1651 618 -1651 0 3
rlabel polysilicon 625 -1645 625 -1645 0 1
rlabel polysilicon 625 -1651 625 -1651 0 3
rlabel polysilicon 632 -1645 632 -1645 0 1
rlabel polysilicon 632 -1651 632 -1651 0 3
rlabel polysilicon 639 -1645 639 -1645 0 1
rlabel polysilicon 639 -1651 639 -1651 0 3
rlabel polysilicon 646 -1645 646 -1645 0 1
rlabel polysilicon 646 -1651 646 -1651 0 3
rlabel polysilicon 653 -1645 653 -1645 0 1
rlabel polysilicon 653 -1651 653 -1651 0 3
rlabel polysilicon 660 -1645 660 -1645 0 1
rlabel polysilicon 663 -1645 663 -1645 0 2
rlabel polysilicon 660 -1651 660 -1651 0 3
rlabel polysilicon 663 -1651 663 -1651 0 4
rlabel polysilicon 667 -1645 667 -1645 0 1
rlabel polysilicon 670 -1645 670 -1645 0 2
rlabel polysilicon 667 -1651 667 -1651 0 3
rlabel polysilicon 670 -1651 670 -1651 0 4
rlabel polysilicon 674 -1645 674 -1645 0 1
rlabel polysilicon 674 -1651 674 -1651 0 3
rlabel polysilicon 681 -1645 681 -1645 0 1
rlabel polysilicon 681 -1651 681 -1651 0 3
rlabel polysilicon 688 -1645 688 -1645 0 1
rlabel polysilicon 688 -1651 688 -1651 0 3
rlabel polysilicon 698 -1645 698 -1645 0 2
rlabel polysilicon 695 -1651 695 -1651 0 3
rlabel polysilicon 702 -1645 702 -1645 0 1
rlabel polysilicon 702 -1651 702 -1651 0 3
rlabel polysilicon 712 -1645 712 -1645 0 2
rlabel polysilicon 709 -1651 709 -1651 0 3
rlabel polysilicon 712 -1651 712 -1651 0 4
rlabel polysilicon 716 -1645 716 -1645 0 1
rlabel polysilicon 716 -1651 716 -1651 0 3
rlabel polysilicon 723 -1645 723 -1645 0 1
rlabel polysilicon 723 -1651 723 -1651 0 3
rlabel polysilicon 730 -1645 730 -1645 0 1
rlabel polysilicon 730 -1651 730 -1651 0 3
rlabel polysilicon 737 -1645 737 -1645 0 1
rlabel polysilicon 740 -1645 740 -1645 0 2
rlabel polysilicon 737 -1651 737 -1651 0 3
rlabel polysilicon 740 -1651 740 -1651 0 4
rlabel polysilicon 744 -1645 744 -1645 0 1
rlabel polysilicon 744 -1651 744 -1651 0 3
rlabel polysilicon 751 -1645 751 -1645 0 1
rlabel polysilicon 751 -1651 751 -1651 0 3
rlabel polysilicon 758 -1645 758 -1645 0 1
rlabel polysilicon 758 -1651 758 -1651 0 3
rlabel polysilicon 768 -1645 768 -1645 0 2
rlabel polysilicon 768 -1651 768 -1651 0 4
rlabel polysilicon 772 -1645 772 -1645 0 1
rlabel polysilicon 772 -1651 772 -1651 0 3
rlabel polysilicon 779 -1645 779 -1645 0 1
rlabel polysilicon 779 -1651 779 -1651 0 3
rlabel polysilicon 786 -1645 786 -1645 0 1
rlabel polysilicon 786 -1651 786 -1651 0 3
rlabel polysilicon 793 -1645 793 -1645 0 1
rlabel polysilicon 793 -1651 793 -1651 0 3
rlabel polysilicon 800 -1645 800 -1645 0 1
rlabel polysilicon 800 -1651 800 -1651 0 3
rlabel polysilicon 807 -1645 807 -1645 0 1
rlabel polysilicon 807 -1651 807 -1651 0 3
rlabel polysilicon 814 -1645 814 -1645 0 1
rlabel polysilicon 817 -1645 817 -1645 0 2
rlabel polysilicon 814 -1651 814 -1651 0 3
rlabel polysilicon 821 -1645 821 -1645 0 1
rlabel polysilicon 821 -1651 821 -1651 0 3
rlabel polysilicon 828 -1645 828 -1645 0 1
rlabel polysilicon 831 -1645 831 -1645 0 2
rlabel polysilicon 828 -1651 828 -1651 0 3
rlabel polysilicon 831 -1651 831 -1651 0 4
rlabel polysilicon 835 -1645 835 -1645 0 1
rlabel polysilicon 835 -1651 835 -1651 0 3
rlabel polysilicon 842 -1645 842 -1645 0 1
rlabel polysilicon 842 -1651 842 -1651 0 3
rlabel polysilicon 849 -1645 849 -1645 0 1
rlabel polysilicon 849 -1651 849 -1651 0 3
rlabel polysilicon 856 -1645 856 -1645 0 1
rlabel polysilicon 856 -1651 856 -1651 0 3
rlabel polysilicon 863 -1645 863 -1645 0 1
rlabel polysilicon 863 -1651 863 -1651 0 3
rlabel polysilicon 870 -1645 870 -1645 0 1
rlabel polysilicon 870 -1651 870 -1651 0 3
rlabel polysilicon 877 -1645 877 -1645 0 1
rlabel polysilicon 877 -1651 877 -1651 0 3
rlabel polysilicon 884 -1645 884 -1645 0 1
rlabel polysilicon 884 -1651 884 -1651 0 3
rlabel polysilicon 891 -1645 891 -1645 0 1
rlabel polysilicon 891 -1651 891 -1651 0 3
rlabel polysilicon 898 -1645 898 -1645 0 1
rlabel polysilicon 898 -1651 898 -1651 0 3
rlabel polysilicon 905 -1645 905 -1645 0 1
rlabel polysilicon 905 -1651 905 -1651 0 3
rlabel polysilicon 912 -1645 912 -1645 0 1
rlabel polysilicon 912 -1651 912 -1651 0 3
rlabel polysilicon 919 -1645 919 -1645 0 1
rlabel polysilicon 922 -1645 922 -1645 0 2
rlabel polysilicon 919 -1651 919 -1651 0 3
rlabel polysilicon 922 -1651 922 -1651 0 4
rlabel polysilicon 926 -1645 926 -1645 0 1
rlabel polysilicon 926 -1651 926 -1651 0 3
rlabel polysilicon 933 -1645 933 -1645 0 1
rlabel polysilicon 933 -1651 933 -1651 0 3
rlabel polysilicon 940 -1645 940 -1645 0 1
rlabel polysilicon 940 -1651 940 -1651 0 3
rlabel polysilicon 943 -1651 943 -1651 0 4
rlabel polysilicon 947 -1645 947 -1645 0 1
rlabel polysilicon 947 -1651 947 -1651 0 3
rlabel polysilicon 954 -1645 954 -1645 0 1
rlabel polysilicon 954 -1651 954 -1651 0 3
rlabel polysilicon 961 -1645 961 -1645 0 1
rlabel polysilicon 961 -1651 961 -1651 0 3
rlabel polysilicon 968 -1645 968 -1645 0 1
rlabel polysilicon 971 -1645 971 -1645 0 2
rlabel polysilicon 968 -1651 968 -1651 0 3
rlabel polysilicon 971 -1651 971 -1651 0 4
rlabel polysilicon 975 -1645 975 -1645 0 1
rlabel polysilicon 975 -1651 975 -1651 0 3
rlabel polysilicon 982 -1645 982 -1645 0 1
rlabel polysilicon 982 -1651 982 -1651 0 3
rlabel polysilicon 989 -1645 989 -1645 0 1
rlabel polysilicon 989 -1651 989 -1651 0 3
rlabel polysilicon 996 -1645 996 -1645 0 1
rlabel polysilicon 996 -1651 996 -1651 0 3
rlabel polysilicon 1003 -1645 1003 -1645 0 1
rlabel polysilicon 1003 -1651 1003 -1651 0 3
rlabel polysilicon 1010 -1645 1010 -1645 0 1
rlabel polysilicon 1010 -1651 1010 -1651 0 3
rlabel polysilicon 1017 -1645 1017 -1645 0 1
rlabel polysilicon 1017 -1651 1017 -1651 0 3
rlabel polysilicon 1024 -1645 1024 -1645 0 1
rlabel polysilicon 1024 -1651 1024 -1651 0 3
rlabel polysilicon 1031 -1645 1031 -1645 0 1
rlabel polysilicon 1031 -1651 1031 -1651 0 3
rlabel polysilicon 1038 -1645 1038 -1645 0 1
rlabel polysilicon 1038 -1651 1038 -1651 0 3
rlabel polysilicon 1041 -1651 1041 -1651 0 4
rlabel polysilicon 1045 -1645 1045 -1645 0 1
rlabel polysilicon 1045 -1651 1045 -1651 0 3
rlabel polysilicon 1052 -1645 1052 -1645 0 1
rlabel polysilicon 1055 -1645 1055 -1645 0 2
rlabel polysilicon 1052 -1651 1052 -1651 0 3
rlabel polysilicon 1055 -1651 1055 -1651 0 4
rlabel polysilicon 1059 -1645 1059 -1645 0 1
rlabel polysilicon 1059 -1651 1059 -1651 0 3
rlabel polysilicon 1066 -1645 1066 -1645 0 1
rlabel polysilicon 1066 -1651 1066 -1651 0 3
rlabel polysilicon 1073 -1645 1073 -1645 0 1
rlabel polysilicon 1073 -1651 1073 -1651 0 3
rlabel polysilicon 1080 -1645 1080 -1645 0 1
rlabel polysilicon 1080 -1651 1080 -1651 0 3
rlabel polysilicon 1087 -1645 1087 -1645 0 1
rlabel polysilicon 1090 -1645 1090 -1645 0 2
rlabel polysilicon 1087 -1651 1087 -1651 0 3
rlabel polysilicon 1094 -1645 1094 -1645 0 1
rlabel polysilicon 1094 -1651 1094 -1651 0 3
rlabel polysilicon 1101 -1645 1101 -1645 0 1
rlabel polysilicon 1101 -1651 1101 -1651 0 3
rlabel polysilicon 1108 -1645 1108 -1645 0 1
rlabel polysilicon 1108 -1651 1108 -1651 0 3
rlabel polysilicon 1115 -1645 1115 -1645 0 1
rlabel polysilicon 1115 -1651 1115 -1651 0 3
rlabel polysilicon 1122 -1645 1122 -1645 0 1
rlabel polysilicon 1122 -1651 1122 -1651 0 3
rlabel polysilicon 1129 -1645 1129 -1645 0 1
rlabel polysilicon 1132 -1645 1132 -1645 0 2
rlabel polysilicon 1129 -1651 1129 -1651 0 3
rlabel polysilicon 1132 -1651 1132 -1651 0 4
rlabel polysilicon 1136 -1645 1136 -1645 0 1
rlabel polysilicon 1136 -1651 1136 -1651 0 3
rlabel polysilicon 1143 -1645 1143 -1645 0 1
rlabel polysilicon 1143 -1651 1143 -1651 0 3
rlabel polysilicon 1150 -1645 1150 -1645 0 1
rlabel polysilicon 1150 -1651 1150 -1651 0 3
rlabel polysilicon 1157 -1645 1157 -1645 0 1
rlabel polysilicon 1157 -1651 1157 -1651 0 3
rlabel polysilicon 1164 -1645 1164 -1645 0 1
rlabel polysilicon 1164 -1651 1164 -1651 0 3
rlabel polysilicon 1171 -1645 1171 -1645 0 1
rlabel polysilicon 1171 -1651 1171 -1651 0 3
rlabel polysilicon 1178 -1645 1178 -1645 0 1
rlabel polysilicon 1178 -1651 1178 -1651 0 3
rlabel polysilicon 1185 -1645 1185 -1645 0 1
rlabel polysilicon 1185 -1651 1185 -1651 0 3
rlabel polysilicon 1192 -1645 1192 -1645 0 1
rlabel polysilicon 1192 -1651 1192 -1651 0 3
rlabel polysilicon 1199 -1645 1199 -1645 0 1
rlabel polysilicon 1199 -1651 1199 -1651 0 3
rlabel polysilicon 1206 -1645 1206 -1645 0 1
rlabel polysilicon 1209 -1645 1209 -1645 0 2
rlabel polysilicon 1206 -1651 1206 -1651 0 3
rlabel polysilicon 1209 -1651 1209 -1651 0 4
rlabel polysilicon 1213 -1645 1213 -1645 0 1
rlabel polysilicon 1213 -1651 1213 -1651 0 3
rlabel polysilicon 1220 -1645 1220 -1645 0 1
rlabel polysilicon 1220 -1651 1220 -1651 0 3
rlabel polysilicon 1227 -1645 1227 -1645 0 1
rlabel polysilicon 1227 -1651 1227 -1651 0 3
rlabel polysilicon 1234 -1645 1234 -1645 0 1
rlabel polysilicon 1234 -1651 1234 -1651 0 3
rlabel polysilicon 1241 -1645 1241 -1645 0 1
rlabel polysilicon 1244 -1645 1244 -1645 0 2
rlabel polysilicon 1241 -1651 1241 -1651 0 3
rlabel polysilicon 1244 -1651 1244 -1651 0 4
rlabel polysilicon 1248 -1645 1248 -1645 0 1
rlabel polysilicon 1248 -1651 1248 -1651 0 3
rlabel polysilicon 1255 -1645 1255 -1645 0 1
rlabel polysilicon 1255 -1651 1255 -1651 0 3
rlabel polysilicon 1262 -1645 1262 -1645 0 1
rlabel polysilicon 1262 -1651 1262 -1651 0 3
rlabel polysilicon 1269 -1645 1269 -1645 0 1
rlabel polysilicon 1269 -1651 1269 -1651 0 3
rlabel polysilicon 1276 -1645 1276 -1645 0 1
rlabel polysilicon 1276 -1651 1276 -1651 0 3
rlabel polysilicon 1283 -1645 1283 -1645 0 1
rlabel polysilicon 1286 -1645 1286 -1645 0 2
rlabel polysilicon 1283 -1651 1283 -1651 0 3
rlabel polysilicon 1286 -1651 1286 -1651 0 4
rlabel polysilicon 1290 -1645 1290 -1645 0 1
rlabel polysilicon 1290 -1651 1290 -1651 0 3
rlabel polysilicon 1297 -1645 1297 -1645 0 1
rlabel polysilicon 1297 -1651 1297 -1651 0 3
rlabel polysilicon 1304 -1645 1304 -1645 0 1
rlabel polysilicon 1307 -1645 1307 -1645 0 2
rlabel polysilicon 1304 -1651 1304 -1651 0 3
rlabel polysilicon 1307 -1651 1307 -1651 0 4
rlabel polysilicon 1311 -1645 1311 -1645 0 1
rlabel polysilicon 1311 -1651 1311 -1651 0 3
rlabel polysilicon 1318 -1645 1318 -1645 0 1
rlabel polysilicon 1318 -1651 1318 -1651 0 3
rlabel polysilicon 1325 -1645 1325 -1645 0 1
rlabel polysilicon 1325 -1651 1325 -1651 0 3
rlabel polysilicon 1332 -1645 1332 -1645 0 1
rlabel polysilicon 1335 -1645 1335 -1645 0 2
rlabel polysilicon 1332 -1651 1332 -1651 0 3
rlabel polysilicon 1335 -1651 1335 -1651 0 4
rlabel polysilicon 1339 -1645 1339 -1645 0 1
rlabel polysilicon 1339 -1651 1339 -1651 0 3
rlabel polysilicon 1346 -1645 1346 -1645 0 1
rlabel polysilicon 1346 -1651 1346 -1651 0 3
rlabel polysilicon 1353 -1645 1353 -1645 0 1
rlabel polysilicon 1356 -1645 1356 -1645 0 2
rlabel polysilicon 1353 -1651 1353 -1651 0 3
rlabel polysilicon 1356 -1651 1356 -1651 0 4
rlabel polysilicon 1360 -1645 1360 -1645 0 1
rlabel polysilicon 1360 -1651 1360 -1651 0 3
rlabel polysilicon 1367 -1645 1367 -1645 0 1
rlabel polysilicon 1367 -1651 1367 -1651 0 3
rlabel polysilicon 1374 -1645 1374 -1645 0 1
rlabel polysilicon 1374 -1651 1374 -1651 0 3
rlabel polysilicon 1381 -1645 1381 -1645 0 1
rlabel polysilicon 1381 -1651 1381 -1651 0 3
rlabel polysilicon 1388 -1645 1388 -1645 0 1
rlabel polysilicon 1388 -1651 1388 -1651 0 3
rlabel polysilicon 1395 -1645 1395 -1645 0 1
rlabel polysilicon 1395 -1651 1395 -1651 0 3
rlabel polysilicon 1402 -1645 1402 -1645 0 1
rlabel polysilicon 1402 -1651 1402 -1651 0 3
rlabel polysilicon 1409 -1645 1409 -1645 0 1
rlabel polysilicon 1409 -1651 1409 -1651 0 3
rlabel polysilicon 1416 -1645 1416 -1645 0 1
rlabel polysilicon 1416 -1651 1416 -1651 0 3
rlabel polysilicon 1423 -1645 1423 -1645 0 1
rlabel polysilicon 1423 -1651 1423 -1651 0 3
rlabel polysilicon 1430 -1645 1430 -1645 0 1
rlabel polysilicon 1430 -1651 1430 -1651 0 3
rlabel polysilicon 1437 -1645 1437 -1645 0 1
rlabel polysilicon 1437 -1651 1437 -1651 0 3
rlabel polysilicon 1444 -1645 1444 -1645 0 1
rlabel polysilicon 1444 -1651 1444 -1651 0 3
rlabel polysilicon 1451 -1645 1451 -1645 0 1
rlabel polysilicon 1451 -1651 1451 -1651 0 3
rlabel polysilicon 1458 -1645 1458 -1645 0 1
rlabel polysilicon 1458 -1651 1458 -1651 0 3
rlabel polysilicon 1465 -1645 1465 -1645 0 1
rlabel polysilicon 1465 -1651 1465 -1651 0 3
rlabel polysilicon 1468 -1651 1468 -1651 0 4
rlabel polysilicon 1472 -1645 1472 -1645 0 1
rlabel polysilicon 1472 -1651 1472 -1651 0 3
rlabel polysilicon 1479 -1645 1479 -1645 0 1
rlabel polysilicon 1479 -1651 1479 -1651 0 3
rlabel polysilicon 1486 -1645 1486 -1645 0 1
rlabel polysilicon 1486 -1651 1486 -1651 0 3
rlabel polysilicon 1493 -1645 1493 -1645 0 1
rlabel polysilicon 1493 -1651 1493 -1651 0 3
rlabel polysilicon 1500 -1645 1500 -1645 0 1
rlabel polysilicon 1503 -1645 1503 -1645 0 2
rlabel polysilicon 1500 -1651 1500 -1651 0 3
rlabel polysilicon 1507 -1645 1507 -1645 0 1
rlabel polysilicon 1507 -1651 1507 -1651 0 3
rlabel polysilicon 1514 -1645 1514 -1645 0 1
rlabel polysilicon 1514 -1651 1514 -1651 0 3
rlabel polysilicon 1521 -1645 1521 -1645 0 1
rlabel polysilicon 1521 -1651 1521 -1651 0 3
rlabel polysilicon 1528 -1645 1528 -1645 0 1
rlabel polysilicon 1528 -1651 1528 -1651 0 3
rlabel polysilicon 1535 -1645 1535 -1645 0 1
rlabel polysilicon 1535 -1651 1535 -1651 0 3
rlabel polysilicon 1542 -1645 1542 -1645 0 1
rlabel polysilicon 1542 -1651 1542 -1651 0 3
rlabel polysilicon 1549 -1645 1549 -1645 0 1
rlabel polysilicon 1549 -1651 1549 -1651 0 3
rlabel polysilicon 1556 -1645 1556 -1645 0 1
rlabel polysilicon 1556 -1651 1556 -1651 0 3
rlabel polysilicon 1563 -1645 1563 -1645 0 1
rlabel polysilicon 1563 -1651 1563 -1651 0 3
rlabel polysilicon 1570 -1645 1570 -1645 0 1
rlabel polysilicon 1570 -1651 1570 -1651 0 3
rlabel polysilicon 1577 -1645 1577 -1645 0 1
rlabel polysilicon 1577 -1651 1577 -1651 0 3
rlabel polysilicon 1584 -1645 1584 -1645 0 1
rlabel polysilicon 1584 -1651 1584 -1651 0 3
rlabel polysilicon 1591 -1645 1591 -1645 0 1
rlabel polysilicon 1591 -1651 1591 -1651 0 3
rlabel polysilicon 1598 -1645 1598 -1645 0 1
rlabel polysilicon 1598 -1651 1598 -1651 0 3
rlabel polysilicon 1605 -1645 1605 -1645 0 1
rlabel polysilicon 1605 -1651 1605 -1651 0 3
rlabel polysilicon 1612 -1645 1612 -1645 0 1
rlabel polysilicon 1612 -1651 1612 -1651 0 3
rlabel polysilicon 1619 -1645 1619 -1645 0 1
rlabel polysilicon 1619 -1651 1619 -1651 0 3
rlabel polysilicon 1626 -1645 1626 -1645 0 1
rlabel polysilicon 1626 -1651 1626 -1651 0 3
rlabel polysilicon 1633 -1645 1633 -1645 0 1
rlabel polysilicon 1633 -1651 1633 -1651 0 3
rlabel polysilicon 1640 -1645 1640 -1645 0 1
rlabel polysilicon 1640 -1651 1640 -1651 0 3
rlabel polysilicon 1647 -1645 1647 -1645 0 1
rlabel polysilicon 1647 -1651 1647 -1651 0 3
rlabel polysilicon 1654 -1645 1654 -1645 0 1
rlabel polysilicon 1654 -1651 1654 -1651 0 3
rlabel polysilicon 1661 -1645 1661 -1645 0 1
rlabel polysilicon 1661 -1651 1661 -1651 0 3
rlabel polysilicon 1668 -1645 1668 -1645 0 1
rlabel polysilicon 1668 -1651 1668 -1651 0 3
rlabel polysilicon 1675 -1645 1675 -1645 0 1
rlabel polysilicon 1675 -1651 1675 -1651 0 3
rlabel polysilicon 1682 -1645 1682 -1645 0 1
rlabel polysilicon 1682 -1651 1682 -1651 0 3
rlabel polysilicon 1689 -1645 1689 -1645 0 1
rlabel polysilicon 1689 -1651 1689 -1651 0 3
rlabel polysilicon 1696 -1645 1696 -1645 0 1
rlabel polysilicon 1696 -1651 1696 -1651 0 3
rlabel polysilicon 1703 -1645 1703 -1645 0 1
rlabel polysilicon 1703 -1651 1703 -1651 0 3
rlabel polysilicon 1710 -1645 1710 -1645 0 1
rlabel polysilicon 1710 -1651 1710 -1651 0 3
rlabel polysilicon 1717 -1645 1717 -1645 0 1
rlabel polysilicon 1717 -1651 1717 -1651 0 3
rlabel polysilicon 1724 -1645 1724 -1645 0 1
rlabel polysilicon 1724 -1651 1724 -1651 0 3
rlabel polysilicon 1731 -1645 1731 -1645 0 1
rlabel polysilicon 1731 -1651 1731 -1651 0 3
rlabel polysilicon 1738 -1645 1738 -1645 0 1
rlabel polysilicon 1738 -1651 1738 -1651 0 3
rlabel polysilicon 1745 -1645 1745 -1645 0 1
rlabel polysilicon 1745 -1651 1745 -1651 0 3
rlabel polysilicon 1752 -1645 1752 -1645 0 1
rlabel polysilicon 1752 -1651 1752 -1651 0 3
rlabel polysilicon 1759 -1645 1759 -1645 0 1
rlabel polysilicon 1759 -1651 1759 -1651 0 3
rlabel polysilicon 1766 -1645 1766 -1645 0 1
rlabel polysilicon 1766 -1651 1766 -1651 0 3
rlabel polysilicon 1773 -1645 1773 -1645 0 1
rlabel polysilicon 1773 -1651 1773 -1651 0 3
rlabel polysilicon 1780 -1645 1780 -1645 0 1
rlabel polysilicon 1780 -1651 1780 -1651 0 3
rlabel polysilicon 1787 -1645 1787 -1645 0 1
rlabel polysilicon 1787 -1651 1787 -1651 0 3
rlabel polysilicon 1794 -1645 1794 -1645 0 1
rlabel polysilicon 1794 -1651 1794 -1651 0 3
rlabel polysilicon 1801 -1645 1801 -1645 0 1
rlabel polysilicon 1801 -1651 1801 -1651 0 3
rlabel polysilicon 1808 -1645 1808 -1645 0 1
rlabel polysilicon 1808 -1651 1808 -1651 0 3
rlabel polysilicon 1815 -1645 1815 -1645 0 1
rlabel polysilicon 1815 -1651 1815 -1651 0 3
rlabel polysilicon 1822 -1645 1822 -1645 0 1
rlabel polysilicon 1822 -1651 1822 -1651 0 3
rlabel polysilicon 1829 -1645 1829 -1645 0 1
rlabel polysilicon 1829 -1651 1829 -1651 0 3
rlabel polysilicon 1836 -1645 1836 -1645 0 1
rlabel polysilicon 1836 -1651 1836 -1651 0 3
rlabel polysilicon 1843 -1645 1843 -1645 0 1
rlabel polysilicon 1843 -1651 1843 -1651 0 3
rlabel polysilicon 1846 -1651 1846 -1651 0 4
rlabel polysilicon 1850 -1645 1850 -1645 0 1
rlabel polysilicon 1850 -1651 1850 -1651 0 3
rlabel polysilicon 1857 -1645 1857 -1645 0 1
rlabel polysilicon 1857 -1651 1857 -1651 0 3
rlabel polysilicon 1864 -1645 1864 -1645 0 1
rlabel polysilicon 1864 -1651 1864 -1651 0 3
rlabel polysilicon 1871 -1645 1871 -1645 0 1
rlabel polysilicon 1871 -1651 1871 -1651 0 3
rlabel polysilicon 1878 -1645 1878 -1645 0 1
rlabel polysilicon 1881 -1645 1881 -1645 0 2
rlabel polysilicon 1878 -1651 1878 -1651 0 3
rlabel polysilicon 1885 -1645 1885 -1645 0 1
rlabel polysilicon 1885 -1651 1885 -1651 0 3
rlabel polysilicon 1892 -1645 1892 -1645 0 1
rlabel polysilicon 1892 -1651 1892 -1651 0 3
rlabel polysilicon 1899 -1645 1899 -1645 0 1
rlabel polysilicon 1899 -1651 1899 -1651 0 3
rlabel polysilicon 1906 -1645 1906 -1645 0 1
rlabel polysilicon 1906 -1651 1906 -1651 0 3
rlabel polysilicon 1913 -1645 1913 -1645 0 1
rlabel polysilicon 1913 -1651 1913 -1651 0 3
rlabel polysilicon 1920 -1645 1920 -1645 0 1
rlabel polysilicon 1920 -1651 1920 -1651 0 3
rlabel polysilicon 1927 -1645 1927 -1645 0 1
rlabel polysilicon 1927 -1651 1927 -1651 0 3
rlabel polysilicon 1934 -1645 1934 -1645 0 1
rlabel polysilicon 1934 -1651 1934 -1651 0 3
rlabel polysilicon 1941 -1645 1941 -1645 0 1
rlabel polysilicon 1941 -1651 1941 -1651 0 3
rlabel polysilicon 1948 -1645 1948 -1645 0 1
rlabel polysilicon 1948 -1651 1948 -1651 0 3
rlabel polysilicon 1976 -1645 1976 -1645 0 1
rlabel polysilicon 1976 -1651 1976 -1651 0 3
rlabel polysilicon 2018 -1645 2018 -1645 0 1
rlabel polysilicon 2018 -1651 2018 -1651 0 3
rlabel polysilicon 9 -1774 9 -1774 0 1
rlabel polysilicon 9 -1780 9 -1780 0 3
rlabel polysilicon 16 -1774 16 -1774 0 1
rlabel polysilicon 16 -1780 16 -1780 0 3
rlabel polysilicon 23 -1774 23 -1774 0 1
rlabel polysilicon 23 -1780 23 -1780 0 3
rlabel polysilicon 30 -1774 30 -1774 0 1
rlabel polysilicon 30 -1780 30 -1780 0 3
rlabel polysilicon 37 -1774 37 -1774 0 1
rlabel polysilicon 37 -1780 37 -1780 0 3
rlabel polysilicon 44 -1774 44 -1774 0 1
rlabel polysilicon 44 -1780 44 -1780 0 3
rlabel polysilicon 51 -1774 51 -1774 0 1
rlabel polysilicon 51 -1780 51 -1780 0 3
rlabel polysilicon 58 -1774 58 -1774 0 1
rlabel polysilicon 58 -1780 58 -1780 0 3
rlabel polysilicon 68 -1774 68 -1774 0 2
rlabel polysilicon 65 -1780 65 -1780 0 3
rlabel polysilicon 68 -1780 68 -1780 0 4
rlabel polysilicon 72 -1774 72 -1774 0 1
rlabel polysilicon 72 -1780 72 -1780 0 3
rlabel polysilicon 79 -1774 79 -1774 0 1
rlabel polysilicon 79 -1780 79 -1780 0 3
rlabel polysilicon 86 -1774 86 -1774 0 1
rlabel polysilicon 86 -1780 86 -1780 0 3
rlabel polysilicon 93 -1774 93 -1774 0 1
rlabel polysilicon 93 -1780 93 -1780 0 3
rlabel polysilicon 100 -1774 100 -1774 0 1
rlabel polysilicon 100 -1780 100 -1780 0 3
rlabel polysilicon 107 -1774 107 -1774 0 1
rlabel polysilicon 107 -1780 107 -1780 0 3
rlabel polysilicon 114 -1774 114 -1774 0 1
rlabel polysilicon 114 -1780 114 -1780 0 3
rlabel polysilicon 121 -1774 121 -1774 0 1
rlabel polysilicon 121 -1780 121 -1780 0 3
rlabel polysilicon 128 -1774 128 -1774 0 1
rlabel polysilicon 131 -1774 131 -1774 0 2
rlabel polysilicon 131 -1780 131 -1780 0 4
rlabel polysilicon 135 -1774 135 -1774 0 1
rlabel polysilicon 135 -1780 135 -1780 0 3
rlabel polysilicon 142 -1774 142 -1774 0 1
rlabel polysilicon 142 -1780 142 -1780 0 3
rlabel polysilicon 149 -1774 149 -1774 0 1
rlabel polysilicon 149 -1780 149 -1780 0 3
rlabel polysilicon 156 -1774 156 -1774 0 1
rlabel polysilicon 156 -1780 156 -1780 0 3
rlabel polysilicon 163 -1774 163 -1774 0 1
rlabel polysilicon 163 -1780 163 -1780 0 3
rlabel polysilicon 170 -1774 170 -1774 0 1
rlabel polysilicon 170 -1780 170 -1780 0 3
rlabel polysilicon 177 -1774 177 -1774 0 1
rlabel polysilicon 177 -1780 177 -1780 0 3
rlabel polysilicon 184 -1774 184 -1774 0 1
rlabel polysilicon 187 -1774 187 -1774 0 2
rlabel polysilicon 184 -1780 184 -1780 0 3
rlabel polysilicon 187 -1780 187 -1780 0 4
rlabel polysilicon 191 -1774 191 -1774 0 1
rlabel polysilicon 194 -1774 194 -1774 0 2
rlabel polysilicon 191 -1780 191 -1780 0 3
rlabel polysilicon 198 -1774 198 -1774 0 1
rlabel polysilicon 201 -1774 201 -1774 0 2
rlabel polysilicon 198 -1780 198 -1780 0 3
rlabel polysilicon 205 -1774 205 -1774 0 1
rlabel polysilicon 205 -1780 205 -1780 0 3
rlabel polysilicon 212 -1774 212 -1774 0 1
rlabel polysilicon 212 -1780 212 -1780 0 3
rlabel polysilicon 219 -1774 219 -1774 0 1
rlabel polysilicon 219 -1780 219 -1780 0 3
rlabel polysilicon 226 -1774 226 -1774 0 1
rlabel polysilicon 226 -1780 226 -1780 0 3
rlabel polysilicon 233 -1774 233 -1774 0 1
rlabel polysilicon 233 -1780 233 -1780 0 3
rlabel polysilicon 240 -1774 240 -1774 0 1
rlabel polysilicon 240 -1780 240 -1780 0 3
rlabel polysilicon 247 -1774 247 -1774 0 1
rlabel polysilicon 247 -1780 247 -1780 0 3
rlabel polysilicon 254 -1774 254 -1774 0 1
rlabel polysilicon 254 -1780 254 -1780 0 3
rlabel polysilicon 261 -1774 261 -1774 0 1
rlabel polysilicon 261 -1780 261 -1780 0 3
rlabel polysilicon 268 -1774 268 -1774 0 1
rlabel polysilicon 268 -1780 268 -1780 0 3
rlabel polysilicon 275 -1774 275 -1774 0 1
rlabel polysilicon 275 -1780 275 -1780 0 3
rlabel polysilicon 282 -1774 282 -1774 0 1
rlabel polysilicon 282 -1780 282 -1780 0 3
rlabel polysilicon 289 -1774 289 -1774 0 1
rlabel polysilicon 289 -1780 289 -1780 0 3
rlabel polysilicon 296 -1774 296 -1774 0 1
rlabel polysilicon 296 -1780 296 -1780 0 3
rlabel polysilicon 303 -1774 303 -1774 0 1
rlabel polysilicon 303 -1780 303 -1780 0 3
rlabel polysilicon 310 -1774 310 -1774 0 1
rlabel polysilicon 310 -1780 310 -1780 0 3
rlabel polysilicon 317 -1774 317 -1774 0 1
rlabel polysilicon 317 -1780 317 -1780 0 3
rlabel polysilicon 324 -1774 324 -1774 0 1
rlabel polysilicon 324 -1780 324 -1780 0 3
rlabel polysilicon 331 -1774 331 -1774 0 1
rlabel polysilicon 331 -1780 331 -1780 0 3
rlabel polysilicon 338 -1774 338 -1774 0 1
rlabel polysilicon 345 -1774 345 -1774 0 1
rlabel polysilicon 345 -1780 345 -1780 0 3
rlabel polysilicon 352 -1774 352 -1774 0 1
rlabel polysilicon 352 -1780 352 -1780 0 3
rlabel polysilicon 359 -1774 359 -1774 0 1
rlabel polysilicon 359 -1780 359 -1780 0 3
rlabel polysilicon 366 -1774 366 -1774 0 1
rlabel polysilicon 366 -1780 366 -1780 0 3
rlabel polysilicon 373 -1774 373 -1774 0 1
rlabel polysilicon 373 -1780 373 -1780 0 3
rlabel polysilicon 380 -1774 380 -1774 0 1
rlabel polysilicon 380 -1780 380 -1780 0 3
rlabel polysilicon 387 -1774 387 -1774 0 1
rlabel polysilicon 387 -1780 387 -1780 0 3
rlabel polysilicon 394 -1774 394 -1774 0 1
rlabel polysilicon 397 -1774 397 -1774 0 2
rlabel polysilicon 394 -1780 394 -1780 0 3
rlabel polysilicon 397 -1780 397 -1780 0 4
rlabel polysilicon 401 -1774 401 -1774 0 1
rlabel polysilicon 401 -1780 401 -1780 0 3
rlabel polysilicon 408 -1774 408 -1774 0 1
rlabel polysilicon 408 -1780 408 -1780 0 3
rlabel polysilicon 415 -1774 415 -1774 0 1
rlabel polysilicon 418 -1774 418 -1774 0 2
rlabel polysilicon 415 -1780 415 -1780 0 3
rlabel polysilicon 418 -1780 418 -1780 0 4
rlabel polysilicon 422 -1774 422 -1774 0 1
rlabel polysilicon 422 -1780 422 -1780 0 3
rlabel polysilicon 429 -1774 429 -1774 0 1
rlabel polysilicon 429 -1780 429 -1780 0 3
rlabel polysilicon 436 -1774 436 -1774 0 1
rlabel polysilicon 436 -1780 436 -1780 0 3
rlabel polysilicon 443 -1774 443 -1774 0 1
rlabel polysilicon 443 -1780 443 -1780 0 3
rlabel polysilicon 450 -1774 450 -1774 0 1
rlabel polysilicon 450 -1780 450 -1780 0 3
rlabel polysilicon 457 -1774 457 -1774 0 1
rlabel polysilicon 457 -1780 457 -1780 0 3
rlabel polysilicon 464 -1774 464 -1774 0 1
rlabel polysilicon 464 -1780 464 -1780 0 3
rlabel polysilicon 471 -1774 471 -1774 0 1
rlabel polysilicon 471 -1780 471 -1780 0 3
rlabel polysilicon 481 -1774 481 -1774 0 2
rlabel polysilicon 478 -1780 478 -1780 0 3
rlabel polysilicon 481 -1780 481 -1780 0 4
rlabel polysilicon 485 -1774 485 -1774 0 1
rlabel polysilicon 485 -1780 485 -1780 0 3
rlabel polysilicon 492 -1774 492 -1774 0 1
rlabel polysilicon 492 -1780 492 -1780 0 3
rlabel polysilicon 499 -1774 499 -1774 0 1
rlabel polysilicon 499 -1780 499 -1780 0 3
rlabel polysilicon 506 -1774 506 -1774 0 1
rlabel polysilicon 506 -1780 506 -1780 0 3
rlabel polysilicon 513 -1774 513 -1774 0 1
rlabel polysilicon 516 -1774 516 -1774 0 2
rlabel polysilicon 513 -1780 513 -1780 0 3
rlabel polysilicon 516 -1780 516 -1780 0 4
rlabel polysilicon 523 -1774 523 -1774 0 2
rlabel polysilicon 520 -1780 520 -1780 0 3
rlabel polysilicon 523 -1780 523 -1780 0 4
rlabel polysilicon 527 -1774 527 -1774 0 1
rlabel polysilicon 527 -1780 527 -1780 0 3
rlabel polysilicon 530 -1780 530 -1780 0 4
rlabel polysilicon 534 -1774 534 -1774 0 1
rlabel polysilicon 534 -1780 534 -1780 0 3
rlabel polysilicon 541 -1774 541 -1774 0 1
rlabel polysilicon 541 -1780 541 -1780 0 3
rlabel polysilicon 548 -1774 548 -1774 0 1
rlabel polysilicon 548 -1780 548 -1780 0 3
rlabel polysilicon 555 -1774 555 -1774 0 1
rlabel polysilicon 558 -1774 558 -1774 0 2
rlabel polysilicon 555 -1780 555 -1780 0 3
rlabel polysilicon 558 -1780 558 -1780 0 4
rlabel polysilicon 565 -1774 565 -1774 0 2
rlabel polysilicon 562 -1780 562 -1780 0 3
rlabel polysilicon 565 -1780 565 -1780 0 4
rlabel polysilicon 569 -1774 569 -1774 0 1
rlabel polysilicon 569 -1780 569 -1780 0 3
rlabel polysilicon 576 -1774 576 -1774 0 1
rlabel polysilicon 576 -1780 576 -1780 0 3
rlabel polysilicon 583 -1774 583 -1774 0 1
rlabel polysilicon 583 -1780 583 -1780 0 3
rlabel polysilicon 590 -1774 590 -1774 0 1
rlabel polysilicon 590 -1780 590 -1780 0 3
rlabel polysilicon 597 -1774 597 -1774 0 1
rlabel polysilicon 600 -1774 600 -1774 0 2
rlabel polysilicon 597 -1780 597 -1780 0 3
rlabel polysilicon 600 -1780 600 -1780 0 4
rlabel polysilicon 604 -1774 604 -1774 0 1
rlabel polysilicon 604 -1780 604 -1780 0 3
rlabel polysilicon 611 -1774 611 -1774 0 1
rlabel polysilicon 611 -1780 611 -1780 0 3
rlabel polysilicon 618 -1774 618 -1774 0 1
rlabel polysilicon 618 -1780 618 -1780 0 3
rlabel polysilicon 625 -1774 625 -1774 0 1
rlabel polysilicon 625 -1780 625 -1780 0 3
rlabel polysilicon 632 -1774 632 -1774 0 1
rlabel polysilicon 632 -1780 632 -1780 0 3
rlabel polysilicon 639 -1774 639 -1774 0 1
rlabel polysilicon 639 -1780 639 -1780 0 3
rlabel polysilicon 646 -1774 646 -1774 0 1
rlabel polysilicon 649 -1774 649 -1774 0 2
rlabel polysilicon 646 -1780 646 -1780 0 3
rlabel polysilicon 649 -1780 649 -1780 0 4
rlabel polysilicon 653 -1774 653 -1774 0 1
rlabel polysilicon 653 -1780 653 -1780 0 3
rlabel polysilicon 660 -1774 660 -1774 0 1
rlabel polysilicon 660 -1780 660 -1780 0 3
rlabel polysilicon 667 -1774 667 -1774 0 1
rlabel polysilicon 667 -1780 667 -1780 0 3
rlabel polysilicon 674 -1774 674 -1774 0 1
rlabel polysilicon 674 -1780 674 -1780 0 3
rlabel polysilicon 681 -1774 681 -1774 0 1
rlabel polysilicon 684 -1774 684 -1774 0 2
rlabel polysilicon 681 -1780 681 -1780 0 3
rlabel polysilicon 684 -1780 684 -1780 0 4
rlabel polysilicon 688 -1774 688 -1774 0 1
rlabel polysilicon 688 -1780 688 -1780 0 3
rlabel polysilicon 695 -1774 695 -1774 0 1
rlabel polysilicon 698 -1774 698 -1774 0 2
rlabel polysilicon 695 -1780 695 -1780 0 3
rlabel polysilicon 702 -1774 702 -1774 0 1
rlabel polysilicon 702 -1780 702 -1780 0 3
rlabel polysilicon 709 -1774 709 -1774 0 1
rlabel polysilicon 709 -1780 709 -1780 0 3
rlabel polysilicon 716 -1774 716 -1774 0 1
rlabel polysilicon 716 -1780 716 -1780 0 3
rlabel polysilicon 723 -1774 723 -1774 0 1
rlabel polysilicon 723 -1780 723 -1780 0 3
rlabel polysilicon 730 -1774 730 -1774 0 1
rlabel polysilicon 730 -1780 730 -1780 0 3
rlabel polysilicon 737 -1774 737 -1774 0 1
rlabel polysilicon 740 -1774 740 -1774 0 2
rlabel polysilicon 737 -1780 737 -1780 0 3
rlabel polysilicon 744 -1774 744 -1774 0 1
rlabel polysilicon 744 -1780 744 -1780 0 3
rlabel polysilicon 751 -1774 751 -1774 0 1
rlabel polysilicon 751 -1780 751 -1780 0 3
rlabel polysilicon 758 -1774 758 -1774 0 1
rlabel polysilicon 758 -1780 758 -1780 0 3
rlabel polysilicon 765 -1774 765 -1774 0 1
rlabel polysilicon 765 -1780 765 -1780 0 3
rlabel polysilicon 772 -1774 772 -1774 0 1
rlabel polysilicon 772 -1780 772 -1780 0 3
rlabel polysilicon 779 -1774 779 -1774 0 1
rlabel polysilicon 779 -1780 779 -1780 0 3
rlabel polysilicon 786 -1774 786 -1774 0 1
rlabel polysilicon 786 -1780 786 -1780 0 3
rlabel polysilicon 793 -1774 793 -1774 0 1
rlabel polysilicon 793 -1780 793 -1780 0 3
rlabel polysilicon 800 -1774 800 -1774 0 1
rlabel polysilicon 800 -1780 800 -1780 0 3
rlabel polysilicon 810 -1774 810 -1774 0 2
rlabel polysilicon 810 -1780 810 -1780 0 4
rlabel polysilicon 814 -1774 814 -1774 0 1
rlabel polysilicon 814 -1780 814 -1780 0 3
rlabel polysilicon 821 -1774 821 -1774 0 1
rlabel polysilicon 821 -1780 821 -1780 0 3
rlabel polysilicon 831 -1774 831 -1774 0 2
rlabel polysilicon 828 -1780 828 -1780 0 3
rlabel polysilicon 831 -1780 831 -1780 0 4
rlabel polysilicon 835 -1774 835 -1774 0 1
rlabel polysilicon 835 -1780 835 -1780 0 3
rlabel polysilicon 842 -1774 842 -1774 0 1
rlabel polysilicon 842 -1780 842 -1780 0 3
rlabel polysilicon 849 -1774 849 -1774 0 1
rlabel polysilicon 849 -1780 849 -1780 0 3
rlabel polysilicon 856 -1774 856 -1774 0 1
rlabel polysilicon 856 -1780 856 -1780 0 3
rlabel polysilicon 863 -1774 863 -1774 0 1
rlabel polysilicon 863 -1780 863 -1780 0 3
rlabel polysilicon 870 -1774 870 -1774 0 1
rlabel polysilicon 870 -1780 870 -1780 0 3
rlabel polysilicon 877 -1774 877 -1774 0 1
rlabel polysilicon 877 -1780 877 -1780 0 3
rlabel polysilicon 887 -1774 887 -1774 0 2
rlabel polysilicon 884 -1780 884 -1780 0 3
rlabel polysilicon 887 -1780 887 -1780 0 4
rlabel polysilicon 891 -1774 891 -1774 0 1
rlabel polysilicon 891 -1780 891 -1780 0 3
rlabel polysilicon 898 -1774 898 -1774 0 1
rlabel polysilicon 901 -1774 901 -1774 0 2
rlabel polysilicon 905 -1774 905 -1774 0 1
rlabel polysilicon 905 -1780 905 -1780 0 3
rlabel polysilicon 912 -1774 912 -1774 0 1
rlabel polysilicon 912 -1780 912 -1780 0 3
rlabel polysilicon 919 -1774 919 -1774 0 1
rlabel polysilicon 919 -1780 919 -1780 0 3
rlabel polysilicon 926 -1774 926 -1774 0 1
rlabel polysilicon 926 -1780 926 -1780 0 3
rlabel polysilicon 933 -1774 933 -1774 0 1
rlabel polysilicon 933 -1780 933 -1780 0 3
rlabel polysilicon 943 -1774 943 -1774 0 2
rlabel polysilicon 940 -1780 940 -1780 0 3
rlabel polysilicon 943 -1780 943 -1780 0 4
rlabel polysilicon 947 -1774 947 -1774 0 1
rlabel polysilicon 947 -1780 947 -1780 0 3
rlabel polysilicon 954 -1774 954 -1774 0 1
rlabel polysilicon 954 -1780 954 -1780 0 3
rlabel polysilicon 961 -1774 961 -1774 0 1
rlabel polysilicon 961 -1780 961 -1780 0 3
rlabel polysilicon 968 -1774 968 -1774 0 1
rlabel polysilicon 968 -1780 968 -1780 0 3
rlabel polysilicon 975 -1774 975 -1774 0 1
rlabel polysilicon 975 -1780 975 -1780 0 3
rlabel polysilicon 982 -1774 982 -1774 0 1
rlabel polysilicon 985 -1774 985 -1774 0 2
rlabel polysilicon 989 -1774 989 -1774 0 1
rlabel polysilicon 989 -1780 989 -1780 0 3
rlabel polysilicon 996 -1774 996 -1774 0 1
rlabel polysilicon 996 -1780 996 -1780 0 3
rlabel polysilicon 1003 -1774 1003 -1774 0 1
rlabel polysilicon 1003 -1780 1003 -1780 0 3
rlabel polysilicon 1010 -1774 1010 -1774 0 1
rlabel polysilicon 1010 -1780 1010 -1780 0 3
rlabel polysilicon 1017 -1774 1017 -1774 0 1
rlabel polysilicon 1017 -1780 1017 -1780 0 3
rlabel polysilicon 1024 -1774 1024 -1774 0 1
rlabel polysilicon 1024 -1780 1024 -1780 0 3
rlabel polysilicon 1031 -1774 1031 -1774 0 1
rlabel polysilicon 1031 -1780 1031 -1780 0 3
rlabel polysilicon 1038 -1774 1038 -1774 0 1
rlabel polysilicon 1038 -1780 1038 -1780 0 3
rlabel polysilicon 1045 -1774 1045 -1774 0 1
rlabel polysilicon 1045 -1780 1045 -1780 0 3
rlabel polysilicon 1052 -1774 1052 -1774 0 1
rlabel polysilicon 1052 -1780 1052 -1780 0 3
rlabel polysilicon 1059 -1774 1059 -1774 0 1
rlabel polysilicon 1059 -1780 1059 -1780 0 3
rlabel polysilicon 1066 -1774 1066 -1774 0 1
rlabel polysilicon 1066 -1780 1066 -1780 0 3
rlabel polysilicon 1073 -1774 1073 -1774 0 1
rlabel polysilicon 1076 -1774 1076 -1774 0 2
rlabel polysilicon 1073 -1780 1073 -1780 0 3
rlabel polysilicon 1076 -1780 1076 -1780 0 4
rlabel polysilicon 1080 -1774 1080 -1774 0 1
rlabel polysilicon 1083 -1774 1083 -1774 0 2
rlabel polysilicon 1080 -1780 1080 -1780 0 3
rlabel polysilicon 1083 -1780 1083 -1780 0 4
rlabel polysilicon 1087 -1774 1087 -1774 0 1
rlabel polysilicon 1087 -1780 1087 -1780 0 3
rlabel polysilicon 1094 -1774 1094 -1774 0 1
rlabel polysilicon 1094 -1780 1094 -1780 0 3
rlabel polysilicon 1101 -1774 1101 -1774 0 1
rlabel polysilicon 1104 -1774 1104 -1774 0 2
rlabel polysilicon 1104 -1780 1104 -1780 0 4
rlabel polysilicon 1111 -1774 1111 -1774 0 2
rlabel polysilicon 1108 -1780 1108 -1780 0 3
rlabel polysilicon 1111 -1780 1111 -1780 0 4
rlabel polysilicon 1115 -1774 1115 -1774 0 1
rlabel polysilicon 1115 -1780 1115 -1780 0 3
rlabel polysilicon 1122 -1774 1122 -1774 0 1
rlabel polysilicon 1122 -1780 1122 -1780 0 3
rlabel polysilicon 1129 -1774 1129 -1774 0 1
rlabel polysilicon 1129 -1780 1129 -1780 0 3
rlabel polysilicon 1136 -1774 1136 -1774 0 1
rlabel polysilicon 1136 -1780 1136 -1780 0 3
rlabel polysilicon 1143 -1774 1143 -1774 0 1
rlabel polysilicon 1143 -1780 1143 -1780 0 3
rlabel polysilicon 1150 -1774 1150 -1774 0 1
rlabel polysilicon 1150 -1780 1150 -1780 0 3
rlabel polysilicon 1157 -1774 1157 -1774 0 1
rlabel polysilicon 1157 -1780 1157 -1780 0 3
rlabel polysilicon 1164 -1774 1164 -1774 0 1
rlabel polysilicon 1164 -1780 1164 -1780 0 3
rlabel polysilicon 1171 -1774 1171 -1774 0 1
rlabel polysilicon 1171 -1780 1171 -1780 0 3
rlabel polysilicon 1178 -1774 1178 -1774 0 1
rlabel polysilicon 1178 -1780 1178 -1780 0 3
rlabel polysilicon 1185 -1774 1185 -1774 0 1
rlabel polysilicon 1185 -1780 1185 -1780 0 3
rlabel polysilicon 1192 -1774 1192 -1774 0 1
rlabel polysilicon 1192 -1780 1192 -1780 0 3
rlabel polysilicon 1199 -1774 1199 -1774 0 1
rlabel polysilicon 1199 -1780 1199 -1780 0 3
rlabel polysilicon 1206 -1774 1206 -1774 0 1
rlabel polysilicon 1206 -1780 1206 -1780 0 3
rlabel polysilicon 1213 -1774 1213 -1774 0 1
rlabel polysilicon 1213 -1780 1213 -1780 0 3
rlabel polysilicon 1220 -1774 1220 -1774 0 1
rlabel polysilicon 1220 -1780 1220 -1780 0 3
rlabel polysilicon 1227 -1774 1227 -1774 0 1
rlabel polysilicon 1227 -1780 1227 -1780 0 3
rlabel polysilicon 1234 -1774 1234 -1774 0 1
rlabel polysilicon 1234 -1780 1234 -1780 0 3
rlabel polysilicon 1241 -1774 1241 -1774 0 1
rlabel polysilicon 1244 -1774 1244 -1774 0 2
rlabel polysilicon 1241 -1780 1241 -1780 0 3
rlabel polysilicon 1244 -1780 1244 -1780 0 4
rlabel polysilicon 1248 -1774 1248 -1774 0 1
rlabel polysilicon 1248 -1780 1248 -1780 0 3
rlabel polysilicon 1255 -1774 1255 -1774 0 1
rlabel polysilicon 1255 -1780 1255 -1780 0 3
rlabel polysilicon 1262 -1774 1262 -1774 0 1
rlabel polysilicon 1262 -1780 1262 -1780 0 3
rlabel polysilicon 1269 -1774 1269 -1774 0 1
rlabel polysilicon 1269 -1780 1269 -1780 0 3
rlabel polysilicon 1276 -1774 1276 -1774 0 1
rlabel polysilicon 1276 -1780 1276 -1780 0 3
rlabel polysilicon 1283 -1774 1283 -1774 0 1
rlabel polysilicon 1283 -1780 1283 -1780 0 3
rlabel polysilicon 1290 -1774 1290 -1774 0 1
rlabel polysilicon 1290 -1780 1290 -1780 0 3
rlabel polysilicon 1297 -1774 1297 -1774 0 1
rlabel polysilicon 1297 -1780 1297 -1780 0 3
rlabel polysilicon 1304 -1774 1304 -1774 0 1
rlabel polysilicon 1307 -1774 1307 -1774 0 2
rlabel polysilicon 1304 -1780 1304 -1780 0 3
rlabel polysilicon 1307 -1780 1307 -1780 0 4
rlabel polysilicon 1311 -1774 1311 -1774 0 1
rlabel polysilicon 1311 -1780 1311 -1780 0 3
rlabel polysilicon 1318 -1774 1318 -1774 0 1
rlabel polysilicon 1318 -1780 1318 -1780 0 3
rlabel polysilicon 1321 -1780 1321 -1780 0 4
rlabel polysilicon 1325 -1774 1325 -1774 0 1
rlabel polysilicon 1325 -1780 1325 -1780 0 3
rlabel polysilicon 1332 -1774 1332 -1774 0 1
rlabel polysilicon 1332 -1780 1332 -1780 0 3
rlabel polysilicon 1339 -1774 1339 -1774 0 1
rlabel polysilicon 1339 -1780 1339 -1780 0 3
rlabel polysilicon 1346 -1774 1346 -1774 0 1
rlabel polysilicon 1346 -1780 1346 -1780 0 3
rlabel polysilicon 1353 -1774 1353 -1774 0 1
rlabel polysilicon 1356 -1774 1356 -1774 0 2
rlabel polysilicon 1360 -1774 1360 -1774 0 1
rlabel polysilicon 1363 -1774 1363 -1774 0 2
rlabel polysilicon 1360 -1780 1360 -1780 0 3
rlabel polysilicon 1363 -1780 1363 -1780 0 4
rlabel polysilicon 1367 -1774 1367 -1774 0 1
rlabel polysilicon 1367 -1780 1367 -1780 0 3
rlabel polysilicon 1374 -1774 1374 -1774 0 1
rlabel polysilicon 1374 -1780 1374 -1780 0 3
rlabel polysilicon 1381 -1774 1381 -1774 0 1
rlabel polysilicon 1381 -1780 1381 -1780 0 3
rlabel polysilicon 1388 -1774 1388 -1774 0 1
rlabel polysilicon 1388 -1780 1388 -1780 0 3
rlabel polysilicon 1395 -1774 1395 -1774 0 1
rlabel polysilicon 1395 -1780 1395 -1780 0 3
rlabel polysilicon 1402 -1774 1402 -1774 0 1
rlabel polysilicon 1402 -1780 1402 -1780 0 3
rlabel polysilicon 1409 -1774 1409 -1774 0 1
rlabel polysilicon 1409 -1780 1409 -1780 0 3
rlabel polysilicon 1416 -1774 1416 -1774 0 1
rlabel polysilicon 1416 -1780 1416 -1780 0 3
rlabel polysilicon 1423 -1774 1423 -1774 0 1
rlabel polysilicon 1423 -1780 1423 -1780 0 3
rlabel polysilicon 1430 -1774 1430 -1774 0 1
rlabel polysilicon 1430 -1780 1430 -1780 0 3
rlabel polysilicon 1437 -1774 1437 -1774 0 1
rlabel polysilicon 1437 -1780 1437 -1780 0 3
rlabel polysilicon 1444 -1774 1444 -1774 0 1
rlabel polysilicon 1444 -1780 1444 -1780 0 3
rlabel polysilicon 1451 -1774 1451 -1774 0 1
rlabel polysilicon 1451 -1780 1451 -1780 0 3
rlabel polysilicon 1458 -1774 1458 -1774 0 1
rlabel polysilicon 1458 -1780 1458 -1780 0 3
rlabel polysilicon 1465 -1774 1465 -1774 0 1
rlabel polysilicon 1468 -1774 1468 -1774 0 2
rlabel polysilicon 1465 -1780 1465 -1780 0 3
rlabel polysilicon 1468 -1780 1468 -1780 0 4
rlabel polysilicon 1472 -1774 1472 -1774 0 1
rlabel polysilicon 1472 -1780 1472 -1780 0 3
rlabel polysilicon 1479 -1774 1479 -1774 0 1
rlabel polysilicon 1479 -1780 1479 -1780 0 3
rlabel polysilicon 1486 -1774 1486 -1774 0 1
rlabel polysilicon 1486 -1780 1486 -1780 0 3
rlabel polysilicon 1493 -1774 1493 -1774 0 1
rlabel polysilicon 1493 -1780 1493 -1780 0 3
rlabel polysilicon 1500 -1774 1500 -1774 0 1
rlabel polysilicon 1500 -1780 1500 -1780 0 3
rlabel polysilicon 1507 -1774 1507 -1774 0 1
rlabel polysilicon 1507 -1780 1507 -1780 0 3
rlabel polysilicon 1514 -1774 1514 -1774 0 1
rlabel polysilicon 1514 -1780 1514 -1780 0 3
rlabel polysilicon 1521 -1774 1521 -1774 0 1
rlabel polysilicon 1521 -1780 1521 -1780 0 3
rlabel polysilicon 1528 -1774 1528 -1774 0 1
rlabel polysilicon 1528 -1780 1528 -1780 0 3
rlabel polysilicon 1535 -1774 1535 -1774 0 1
rlabel polysilicon 1535 -1780 1535 -1780 0 3
rlabel polysilicon 1542 -1774 1542 -1774 0 1
rlabel polysilicon 1542 -1780 1542 -1780 0 3
rlabel polysilicon 1549 -1774 1549 -1774 0 1
rlabel polysilicon 1549 -1780 1549 -1780 0 3
rlabel polysilicon 1556 -1774 1556 -1774 0 1
rlabel polysilicon 1556 -1780 1556 -1780 0 3
rlabel polysilicon 1563 -1774 1563 -1774 0 1
rlabel polysilicon 1563 -1780 1563 -1780 0 3
rlabel polysilicon 1570 -1774 1570 -1774 0 1
rlabel polysilicon 1570 -1780 1570 -1780 0 3
rlabel polysilicon 1577 -1774 1577 -1774 0 1
rlabel polysilicon 1577 -1780 1577 -1780 0 3
rlabel polysilicon 1584 -1774 1584 -1774 0 1
rlabel polysilicon 1584 -1780 1584 -1780 0 3
rlabel polysilicon 1591 -1774 1591 -1774 0 1
rlabel polysilicon 1591 -1780 1591 -1780 0 3
rlabel polysilicon 1598 -1774 1598 -1774 0 1
rlabel polysilicon 1598 -1780 1598 -1780 0 3
rlabel polysilicon 1605 -1774 1605 -1774 0 1
rlabel polysilicon 1605 -1780 1605 -1780 0 3
rlabel polysilicon 1612 -1774 1612 -1774 0 1
rlabel polysilicon 1612 -1780 1612 -1780 0 3
rlabel polysilicon 1619 -1774 1619 -1774 0 1
rlabel polysilicon 1619 -1780 1619 -1780 0 3
rlabel polysilicon 1626 -1774 1626 -1774 0 1
rlabel polysilicon 1626 -1780 1626 -1780 0 3
rlabel polysilicon 1633 -1774 1633 -1774 0 1
rlabel polysilicon 1633 -1780 1633 -1780 0 3
rlabel polysilicon 1640 -1774 1640 -1774 0 1
rlabel polysilicon 1640 -1780 1640 -1780 0 3
rlabel polysilicon 1647 -1774 1647 -1774 0 1
rlabel polysilicon 1647 -1780 1647 -1780 0 3
rlabel polysilicon 1654 -1774 1654 -1774 0 1
rlabel polysilicon 1654 -1780 1654 -1780 0 3
rlabel polysilicon 1661 -1774 1661 -1774 0 1
rlabel polysilicon 1661 -1780 1661 -1780 0 3
rlabel polysilicon 1668 -1774 1668 -1774 0 1
rlabel polysilicon 1668 -1780 1668 -1780 0 3
rlabel polysilicon 1675 -1774 1675 -1774 0 1
rlabel polysilicon 1675 -1780 1675 -1780 0 3
rlabel polysilicon 1682 -1774 1682 -1774 0 1
rlabel polysilicon 1682 -1780 1682 -1780 0 3
rlabel polysilicon 1689 -1774 1689 -1774 0 1
rlabel polysilicon 1689 -1780 1689 -1780 0 3
rlabel polysilicon 1696 -1774 1696 -1774 0 1
rlabel polysilicon 1696 -1780 1696 -1780 0 3
rlabel polysilicon 1703 -1774 1703 -1774 0 1
rlabel polysilicon 1703 -1780 1703 -1780 0 3
rlabel polysilicon 1710 -1774 1710 -1774 0 1
rlabel polysilicon 1710 -1780 1710 -1780 0 3
rlabel polysilicon 1717 -1774 1717 -1774 0 1
rlabel polysilicon 1717 -1780 1717 -1780 0 3
rlabel polysilicon 1724 -1774 1724 -1774 0 1
rlabel polysilicon 1724 -1780 1724 -1780 0 3
rlabel polysilicon 1731 -1774 1731 -1774 0 1
rlabel polysilicon 1731 -1780 1731 -1780 0 3
rlabel polysilicon 1738 -1774 1738 -1774 0 1
rlabel polysilicon 1738 -1780 1738 -1780 0 3
rlabel polysilicon 1745 -1774 1745 -1774 0 1
rlabel polysilicon 1745 -1780 1745 -1780 0 3
rlabel polysilicon 1752 -1774 1752 -1774 0 1
rlabel polysilicon 1752 -1780 1752 -1780 0 3
rlabel polysilicon 1759 -1774 1759 -1774 0 1
rlabel polysilicon 1759 -1780 1759 -1780 0 3
rlabel polysilicon 1766 -1774 1766 -1774 0 1
rlabel polysilicon 1766 -1780 1766 -1780 0 3
rlabel polysilicon 1773 -1774 1773 -1774 0 1
rlabel polysilicon 1773 -1780 1773 -1780 0 3
rlabel polysilicon 1780 -1774 1780 -1774 0 1
rlabel polysilicon 1780 -1780 1780 -1780 0 3
rlabel polysilicon 1787 -1774 1787 -1774 0 1
rlabel polysilicon 1787 -1780 1787 -1780 0 3
rlabel polysilicon 1794 -1774 1794 -1774 0 1
rlabel polysilicon 1794 -1780 1794 -1780 0 3
rlabel polysilicon 1801 -1774 1801 -1774 0 1
rlabel polysilicon 1801 -1780 1801 -1780 0 3
rlabel polysilicon 1808 -1774 1808 -1774 0 1
rlabel polysilicon 1808 -1780 1808 -1780 0 3
rlabel polysilicon 1815 -1774 1815 -1774 0 1
rlabel polysilicon 1815 -1780 1815 -1780 0 3
rlabel polysilicon 1822 -1774 1822 -1774 0 1
rlabel polysilicon 1822 -1780 1822 -1780 0 3
rlabel polysilicon 1829 -1774 1829 -1774 0 1
rlabel polysilicon 1829 -1780 1829 -1780 0 3
rlabel polysilicon 1836 -1774 1836 -1774 0 1
rlabel polysilicon 1836 -1780 1836 -1780 0 3
rlabel polysilicon 1843 -1774 1843 -1774 0 1
rlabel polysilicon 1843 -1780 1843 -1780 0 3
rlabel polysilicon 1850 -1774 1850 -1774 0 1
rlabel polysilicon 1850 -1780 1850 -1780 0 3
rlabel polysilicon 1857 -1774 1857 -1774 0 1
rlabel polysilicon 1857 -1780 1857 -1780 0 3
rlabel polysilicon 1864 -1774 1864 -1774 0 1
rlabel polysilicon 1864 -1780 1864 -1780 0 3
rlabel polysilicon 1871 -1774 1871 -1774 0 1
rlabel polysilicon 1871 -1780 1871 -1780 0 3
rlabel polysilicon 1878 -1774 1878 -1774 0 1
rlabel polysilicon 1878 -1780 1878 -1780 0 3
rlabel polysilicon 1885 -1774 1885 -1774 0 1
rlabel polysilicon 1885 -1780 1885 -1780 0 3
rlabel polysilicon 1892 -1774 1892 -1774 0 1
rlabel polysilicon 1892 -1780 1892 -1780 0 3
rlabel polysilicon 1899 -1774 1899 -1774 0 1
rlabel polysilicon 1899 -1780 1899 -1780 0 3
rlabel polysilicon 1906 -1774 1906 -1774 0 1
rlabel polysilicon 1906 -1780 1906 -1780 0 3
rlabel polysilicon 1913 -1774 1913 -1774 0 1
rlabel polysilicon 1913 -1780 1913 -1780 0 3
rlabel polysilicon 1920 -1774 1920 -1774 0 1
rlabel polysilicon 1920 -1780 1920 -1780 0 3
rlabel polysilicon 1927 -1774 1927 -1774 0 1
rlabel polysilicon 1927 -1780 1927 -1780 0 3
rlabel polysilicon 1934 -1774 1934 -1774 0 1
rlabel polysilicon 1937 -1774 1937 -1774 0 2
rlabel polysilicon 1934 -1780 1934 -1780 0 3
rlabel polysilicon 1941 -1774 1941 -1774 0 1
rlabel polysilicon 1944 -1774 1944 -1774 0 2
rlabel polysilicon 1941 -1780 1941 -1780 0 3
rlabel polysilicon 1944 -1780 1944 -1780 0 4
rlabel polysilicon 1948 -1774 1948 -1774 0 1
rlabel polysilicon 1948 -1780 1948 -1780 0 3
rlabel polysilicon 1955 -1774 1955 -1774 0 1
rlabel polysilicon 1955 -1780 1955 -1780 0 3
rlabel polysilicon 1962 -1774 1962 -1774 0 1
rlabel polysilicon 1962 -1780 1962 -1780 0 3
rlabel polysilicon 1969 -1774 1969 -1774 0 1
rlabel polysilicon 1969 -1780 1969 -1780 0 3
rlabel polysilicon 2018 -1774 2018 -1774 0 1
rlabel polysilicon 2018 -1780 2018 -1780 0 3
rlabel polysilicon 5 -1905 5 -1905 0 4
rlabel polysilicon 16 -1899 16 -1899 0 1
rlabel polysilicon 16 -1905 16 -1905 0 3
rlabel polysilicon 23 -1899 23 -1899 0 1
rlabel polysilicon 23 -1905 23 -1905 0 3
rlabel polysilicon 30 -1899 30 -1899 0 1
rlabel polysilicon 30 -1905 30 -1905 0 3
rlabel polysilicon 37 -1899 37 -1899 0 1
rlabel polysilicon 37 -1905 37 -1905 0 3
rlabel polysilicon 44 -1899 44 -1899 0 1
rlabel polysilicon 44 -1905 44 -1905 0 3
rlabel polysilicon 51 -1899 51 -1899 0 1
rlabel polysilicon 51 -1905 51 -1905 0 3
rlabel polysilicon 58 -1899 58 -1899 0 1
rlabel polysilicon 61 -1899 61 -1899 0 2
rlabel polysilicon 61 -1905 61 -1905 0 4
rlabel polysilicon 65 -1899 65 -1899 0 1
rlabel polysilicon 65 -1905 65 -1905 0 3
rlabel polysilicon 72 -1899 72 -1899 0 1
rlabel polysilicon 72 -1905 72 -1905 0 3
rlabel polysilicon 79 -1899 79 -1899 0 1
rlabel polysilicon 79 -1905 79 -1905 0 3
rlabel polysilicon 86 -1899 86 -1899 0 1
rlabel polysilicon 86 -1905 86 -1905 0 3
rlabel polysilicon 93 -1899 93 -1899 0 1
rlabel polysilicon 93 -1905 93 -1905 0 3
rlabel polysilicon 103 -1899 103 -1899 0 2
rlabel polysilicon 100 -1905 100 -1905 0 3
rlabel polysilicon 103 -1905 103 -1905 0 4
rlabel polysilicon 107 -1899 107 -1899 0 1
rlabel polysilicon 107 -1905 107 -1905 0 3
rlabel polysilicon 114 -1899 114 -1899 0 1
rlabel polysilicon 114 -1905 114 -1905 0 3
rlabel polysilicon 121 -1899 121 -1899 0 1
rlabel polysilicon 121 -1905 121 -1905 0 3
rlabel polysilicon 128 -1899 128 -1899 0 1
rlabel polysilicon 128 -1905 128 -1905 0 3
rlabel polysilicon 135 -1899 135 -1899 0 1
rlabel polysilicon 138 -1899 138 -1899 0 2
rlabel polysilicon 135 -1905 135 -1905 0 3
rlabel polysilicon 138 -1905 138 -1905 0 4
rlabel polysilicon 142 -1899 142 -1899 0 1
rlabel polysilicon 145 -1899 145 -1899 0 2
rlabel polysilicon 142 -1905 142 -1905 0 3
rlabel polysilicon 145 -1905 145 -1905 0 4
rlabel polysilicon 149 -1899 149 -1899 0 1
rlabel polysilicon 149 -1905 149 -1905 0 3
rlabel polysilicon 156 -1899 156 -1899 0 1
rlabel polysilicon 156 -1905 156 -1905 0 3
rlabel polysilicon 163 -1899 163 -1899 0 1
rlabel polysilicon 163 -1905 163 -1905 0 3
rlabel polysilicon 170 -1899 170 -1899 0 1
rlabel polysilicon 170 -1905 170 -1905 0 3
rlabel polysilicon 177 -1899 177 -1899 0 1
rlabel polysilicon 177 -1905 177 -1905 0 3
rlabel polysilicon 184 -1899 184 -1899 0 1
rlabel polysilicon 184 -1905 184 -1905 0 3
rlabel polysilicon 191 -1899 191 -1899 0 1
rlabel polysilicon 191 -1905 191 -1905 0 3
rlabel polysilicon 198 -1899 198 -1899 0 1
rlabel polysilicon 201 -1899 201 -1899 0 2
rlabel polysilicon 198 -1905 198 -1905 0 3
rlabel polysilicon 205 -1899 205 -1899 0 1
rlabel polysilicon 205 -1905 205 -1905 0 3
rlabel polysilicon 212 -1899 212 -1899 0 1
rlabel polysilicon 212 -1905 212 -1905 0 3
rlabel polysilicon 219 -1899 219 -1899 0 1
rlabel polysilicon 219 -1905 219 -1905 0 3
rlabel polysilicon 226 -1899 226 -1899 0 1
rlabel polysilicon 226 -1905 226 -1905 0 3
rlabel polysilicon 233 -1899 233 -1899 0 1
rlabel polysilicon 233 -1905 233 -1905 0 3
rlabel polysilicon 240 -1899 240 -1899 0 1
rlabel polysilicon 240 -1905 240 -1905 0 3
rlabel polysilicon 247 -1899 247 -1899 0 1
rlabel polysilicon 247 -1905 247 -1905 0 3
rlabel polysilicon 254 -1899 254 -1899 0 1
rlabel polysilicon 254 -1905 254 -1905 0 3
rlabel polysilicon 261 -1899 261 -1899 0 1
rlabel polysilicon 261 -1905 261 -1905 0 3
rlabel polysilicon 268 -1899 268 -1899 0 1
rlabel polysilicon 268 -1905 268 -1905 0 3
rlabel polysilicon 275 -1899 275 -1899 0 1
rlabel polysilicon 275 -1905 275 -1905 0 3
rlabel polysilicon 282 -1899 282 -1899 0 1
rlabel polysilicon 282 -1905 282 -1905 0 3
rlabel polysilicon 289 -1899 289 -1899 0 1
rlabel polysilicon 289 -1905 289 -1905 0 3
rlabel polysilicon 296 -1899 296 -1899 0 1
rlabel polysilicon 296 -1905 296 -1905 0 3
rlabel polysilicon 303 -1899 303 -1899 0 1
rlabel polysilicon 303 -1905 303 -1905 0 3
rlabel polysilicon 310 -1899 310 -1899 0 1
rlabel polysilicon 310 -1905 310 -1905 0 3
rlabel polysilicon 317 -1899 317 -1899 0 1
rlabel polysilicon 317 -1905 317 -1905 0 3
rlabel polysilicon 324 -1899 324 -1899 0 1
rlabel polysilicon 324 -1905 324 -1905 0 3
rlabel polysilicon 331 -1899 331 -1899 0 1
rlabel polysilicon 331 -1905 331 -1905 0 3
rlabel polysilicon 338 -1905 338 -1905 0 3
rlabel polysilicon 345 -1899 345 -1899 0 1
rlabel polysilicon 345 -1905 345 -1905 0 3
rlabel polysilicon 352 -1899 352 -1899 0 1
rlabel polysilicon 352 -1905 352 -1905 0 3
rlabel polysilicon 359 -1899 359 -1899 0 1
rlabel polysilicon 359 -1905 359 -1905 0 3
rlabel polysilicon 366 -1899 366 -1899 0 1
rlabel polysilicon 366 -1905 366 -1905 0 3
rlabel polysilicon 373 -1899 373 -1899 0 1
rlabel polysilicon 373 -1905 373 -1905 0 3
rlabel polysilicon 380 -1899 380 -1899 0 1
rlabel polysilicon 380 -1905 380 -1905 0 3
rlabel polysilicon 387 -1899 387 -1899 0 1
rlabel polysilicon 387 -1905 387 -1905 0 3
rlabel polysilicon 394 -1899 394 -1899 0 1
rlabel polysilicon 394 -1905 394 -1905 0 3
rlabel polysilicon 401 -1899 401 -1899 0 1
rlabel polysilicon 404 -1899 404 -1899 0 2
rlabel polysilicon 408 -1899 408 -1899 0 1
rlabel polysilicon 408 -1905 408 -1905 0 3
rlabel polysilicon 415 -1899 415 -1899 0 1
rlabel polysilicon 415 -1905 415 -1905 0 3
rlabel polysilicon 422 -1899 422 -1899 0 1
rlabel polysilicon 422 -1905 422 -1905 0 3
rlabel polysilicon 429 -1899 429 -1899 0 1
rlabel polysilicon 429 -1905 429 -1905 0 3
rlabel polysilicon 436 -1899 436 -1899 0 1
rlabel polysilicon 436 -1905 436 -1905 0 3
rlabel polysilicon 443 -1899 443 -1899 0 1
rlabel polysilicon 443 -1905 443 -1905 0 3
rlabel polysilicon 450 -1899 450 -1899 0 1
rlabel polysilicon 450 -1905 450 -1905 0 3
rlabel polysilicon 457 -1899 457 -1899 0 1
rlabel polysilicon 457 -1905 457 -1905 0 3
rlabel polysilicon 464 -1899 464 -1899 0 1
rlabel polysilicon 464 -1905 464 -1905 0 3
rlabel polysilicon 471 -1899 471 -1899 0 1
rlabel polysilicon 471 -1905 471 -1905 0 3
rlabel polysilicon 478 -1899 478 -1899 0 1
rlabel polysilicon 481 -1905 481 -1905 0 4
rlabel polysilicon 485 -1899 485 -1899 0 1
rlabel polysilicon 488 -1899 488 -1899 0 2
rlabel polysilicon 485 -1905 485 -1905 0 3
rlabel polysilicon 488 -1905 488 -1905 0 4
rlabel polysilicon 492 -1899 492 -1899 0 1
rlabel polysilicon 492 -1905 492 -1905 0 3
rlabel polysilicon 499 -1899 499 -1899 0 1
rlabel polysilicon 499 -1905 499 -1905 0 3
rlabel polysilicon 509 -1899 509 -1899 0 2
rlabel polysilicon 506 -1905 506 -1905 0 3
rlabel polysilicon 509 -1905 509 -1905 0 4
rlabel polysilicon 513 -1899 513 -1899 0 1
rlabel polysilicon 513 -1905 513 -1905 0 3
rlabel polysilicon 520 -1899 520 -1899 0 1
rlabel polysilicon 520 -1905 520 -1905 0 3
rlabel polysilicon 527 -1899 527 -1899 0 1
rlabel polysilicon 530 -1899 530 -1899 0 2
rlabel polysilicon 527 -1905 527 -1905 0 3
rlabel polysilicon 534 -1899 534 -1899 0 1
rlabel polysilicon 534 -1905 534 -1905 0 3
rlabel polysilicon 541 -1899 541 -1899 0 1
rlabel polysilicon 541 -1905 541 -1905 0 3
rlabel polysilicon 548 -1899 548 -1899 0 1
rlabel polysilicon 548 -1905 548 -1905 0 3
rlabel polysilicon 555 -1899 555 -1899 0 1
rlabel polysilicon 555 -1905 555 -1905 0 3
rlabel polysilicon 562 -1899 562 -1899 0 1
rlabel polysilicon 562 -1905 562 -1905 0 3
rlabel polysilicon 569 -1899 569 -1899 0 1
rlabel polysilicon 569 -1905 569 -1905 0 3
rlabel polysilicon 579 -1899 579 -1899 0 2
rlabel polysilicon 579 -1905 579 -1905 0 4
rlabel polysilicon 583 -1899 583 -1899 0 1
rlabel polysilicon 583 -1905 583 -1905 0 3
rlabel polysilicon 590 -1899 590 -1899 0 1
rlabel polysilicon 590 -1905 590 -1905 0 3
rlabel polysilicon 597 -1899 597 -1899 0 1
rlabel polysilicon 597 -1905 597 -1905 0 3
rlabel polysilicon 604 -1899 604 -1899 0 1
rlabel polysilicon 604 -1905 604 -1905 0 3
rlabel polysilicon 611 -1899 611 -1899 0 1
rlabel polysilicon 614 -1899 614 -1899 0 2
rlabel polysilicon 611 -1905 611 -1905 0 3
rlabel polysilicon 614 -1905 614 -1905 0 4
rlabel polysilicon 618 -1899 618 -1899 0 1
rlabel polysilicon 618 -1905 618 -1905 0 3
rlabel polysilicon 625 -1899 625 -1899 0 1
rlabel polysilicon 625 -1905 625 -1905 0 3
rlabel polysilicon 632 -1899 632 -1899 0 1
rlabel polysilicon 632 -1905 632 -1905 0 3
rlabel polysilicon 639 -1899 639 -1899 0 1
rlabel polysilicon 639 -1905 639 -1905 0 3
rlabel polysilicon 646 -1899 646 -1899 0 1
rlabel polysilicon 646 -1905 646 -1905 0 3
rlabel polysilicon 653 -1899 653 -1899 0 1
rlabel polysilicon 653 -1905 653 -1905 0 3
rlabel polysilicon 660 -1899 660 -1899 0 1
rlabel polysilicon 660 -1905 660 -1905 0 3
rlabel polysilicon 667 -1899 667 -1899 0 1
rlabel polysilicon 674 -1899 674 -1899 0 1
rlabel polysilicon 674 -1905 674 -1905 0 3
rlabel polysilicon 681 -1899 681 -1899 0 1
rlabel polysilicon 681 -1905 681 -1905 0 3
rlabel polysilicon 691 -1899 691 -1899 0 2
rlabel polysilicon 688 -1905 688 -1905 0 3
rlabel polysilicon 691 -1905 691 -1905 0 4
rlabel polysilicon 695 -1899 695 -1899 0 1
rlabel polysilicon 695 -1905 695 -1905 0 3
rlabel polysilicon 702 -1899 702 -1899 0 1
rlabel polysilicon 702 -1905 702 -1905 0 3
rlabel polysilicon 709 -1899 709 -1899 0 1
rlabel polysilicon 709 -1905 709 -1905 0 3
rlabel polysilicon 716 -1899 716 -1899 0 1
rlabel polysilicon 719 -1899 719 -1899 0 2
rlabel polysilicon 716 -1905 716 -1905 0 3
rlabel polysilicon 719 -1905 719 -1905 0 4
rlabel polysilicon 723 -1899 723 -1899 0 1
rlabel polysilicon 723 -1905 723 -1905 0 3
rlabel polysilicon 726 -1905 726 -1905 0 4
rlabel polysilicon 730 -1899 730 -1899 0 1
rlabel polysilicon 730 -1905 730 -1905 0 3
rlabel polysilicon 737 -1899 737 -1899 0 1
rlabel polysilicon 737 -1905 737 -1905 0 3
rlabel polysilicon 744 -1899 744 -1899 0 1
rlabel polysilicon 744 -1905 744 -1905 0 3
rlabel polysilicon 751 -1899 751 -1899 0 1
rlabel polysilicon 751 -1905 751 -1905 0 3
rlabel polysilicon 758 -1899 758 -1899 0 1
rlabel polysilicon 758 -1905 758 -1905 0 3
rlabel polysilicon 765 -1899 765 -1899 0 1
rlabel polysilicon 768 -1899 768 -1899 0 2
rlabel polysilicon 765 -1905 765 -1905 0 3
rlabel polysilicon 768 -1905 768 -1905 0 4
rlabel polysilicon 772 -1899 772 -1899 0 1
rlabel polysilicon 772 -1905 772 -1905 0 3
rlabel polysilicon 775 -1905 775 -1905 0 4
rlabel polysilicon 779 -1899 779 -1899 0 1
rlabel polysilicon 779 -1905 779 -1905 0 3
rlabel polysilicon 786 -1899 786 -1899 0 1
rlabel polysilicon 786 -1905 786 -1905 0 3
rlabel polysilicon 793 -1899 793 -1899 0 1
rlabel polysilicon 793 -1905 793 -1905 0 3
rlabel polysilicon 800 -1899 800 -1899 0 1
rlabel polysilicon 800 -1905 800 -1905 0 3
rlabel polysilicon 807 -1899 807 -1899 0 1
rlabel polysilicon 807 -1905 807 -1905 0 3
rlabel polysilicon 814 -1899 814 -1899 0 1
rlabel polysilicon 814 -1905 814 -1905 0 3
rlabel polysilicon 821 -1899 821 -1899 0 1
rlabel polysilicon 821 -1905 821 -1905 0 3
rlabel polysilicon 828 -1899 828 -1899 0 1
rlabel polysilicon 828 -1905 828 -1905 0 3
rlabel polysilicon 835 -1899 835 -1899 0 1
rlabel polysilicon 835 -1905 835 -1905 0 3
rlabel polysilicon 842 -1899 842 -1899 0 1
rlabel polysilicon 842 -1905 842 -1905 0 3
rlabel polysilicon 849 -1899 849 -1899 0 1
rlabel polysilicon 849 -1905 849 -1905 0 3
rlabel polysilicon 856 -1899 856 -1899 0 1
rlabel polysilicon 856 -1905 856 -1905 0 3
rlabel polysilicon 863 -1899 863 -1899 0 1
rlabel polysilicon 863 -1905 863 -1905 0 3
rlabel polysilicon 870 -1899 870 -1899 0 1
rlabel polysilicon 870 -1905 870 -1905 0 3
rlabel polysilicon 877 -1899 877 -1899 0 1
rlabel polysilicon 877 -1905 877 -1905 0 3
rlabel polysilicon 884 -1899 884 -1899 0 1
rlabel polysilicon 887 -1899 887 -1899 0 2
rlabel polysilicon 884 -1905 884 -1905 0 3
rlabel polysilicon 887 -1905 887 -1905 0 4
rlabel polysilicon 891 -1899 891 -1899 0 1
rlabel polysilicon 891 -1905 891 -1905 0 3
rlabel polysilicon 898 -1899 898 -1899 0 1
rlabel polysilicon 898 -1905 898 -1905 0 3
rlabel polysilicon 905 -1899 905 -1899 0 1
rlabel polysilicon 908 -1899 908 -1899 0 2
rlabel polysilicon 905 -1905 905 -1905 0 3
rlabel polysilicon 908 -1905 908 -1905 0 4
rlabel polysilicon 912 -1899 912 -1899 0 1
rlabel polysilicon 912 -1905 912 -1905 0 3
rlabel polysilicon 919 -1899 919 -1899 0 1
rlabel polysilicon 919 -1905 919 -1905 0 3
rlabel polysilicon 926 -1899 926 -1899 0 1
rlabel polysilicon 926 -1905 926 -1905 0 3
rlabel polysilicon 933 -1899 933 -1899 0 1
rlabel polysilicon 936 -1899 936 -1899 0 2
rlabel polysilicon 933 -1905 933 -1905 0 3
rlabel polysilicon 936 -1905 936 -1905 0 4
rlabel polysilicon 940 -1899 940 -1899 0 1
rlabel polysilicon 940 -1905 940 -1905 0 3
rlabel polysilicon 947 -1899 947 -1899 0 1
rlabel polysilicon 947 -1905 947 -1905 0 3
rlabel polysilicon 954 -1899 954 -1899 0 1
rlabel polysilicon 954 -1905 954 -1905 0 3
rlabel polysilicon 961 -1899 961 -1899 0 1
rlabel polysilicon 961 -1905 961 -1905 0 3
rlabel polysilicon 968 -1899 968 -1899 0 1
rlabel polysilicon 968 -1905 968 -1905 0 3
rlabel polysilicon 975 -1899 975 -1899 0 1
rlabel polysilicon 975 -1905 975 -1905 0 3
rlabel polysilicon 982 -1899 982 -1899 0 1
rlabel polysilicon 985 -1899 985 -1899 0 2
rlabel polysilicon 982 -1905 982 -1905 0 3
rlabel polysilicon 985 -1905 985 -1905 0 4
rlabel polysilicon 989 -1899 989 -1899 0 1
rlabel polysilicon 989 -1905 989 -1905 0 3
rlabel polysilicon 996 -1899 996 -1899 0 1
rlabel polysilicon 996 -1905 996 -1905 0 3
rlabel polysilicon 1003 -1899 1003 -1899 0 1
rlabel polysilicon 1003 -1905 1003 -1905 0 3
rlabel polysilicon 1010 -1899 1010 -1899 0 1
rlabel polysilicon 1010 -1905 1010 -1905 0 3
rlabel polysilicon 1017 -1899 1017 -1899 0 1
rlabel polysilicon 1017 -1905 1017 -1905 0 3
rlabel polysilicon 1024 -1899 1024 -1899 0 1
rlabel polysilicon 1024 -1905 1024 -1905 0 3
rlabel polysilicon 1027 -1905 1027 -1905 0 4
rlabel polysilicon 1031 -1899 1031 -1899 0 1
rlabel polysilicon 1031 -1905 1031 -1905 0 3
rlabel polysilicon 1038 -1899 1038 -1899 0 1
rlabel polysilicon 1038 -1905 1038 -1905 0 3
rlabel polysilicon 1045 -1899 1045 -1899 0 1
rlabel polysilicon 1045 -1905 1045 -1905 0 3
rlabel polysilicon 1052 -1899 1052 -1899 0 1
rlabel polysilicon 1052 -1905 1052 -1905 0 3
rlabel polysilicon 1059 -1899 1059 -1899 0 1
rlabel polysilicon 1059 -1905 1059 -1905 0 3
rlabel polysilicon 1066 -1899 1066 -1899 0 1
rlabel polysilicon 1066 -1905 1066 -1905 0 3
rlabel polysilicon 1073 -1899 1073 -1899 0 1
rlabel polysilicon 1073 -1905 1073 -1905 0 3
rlabel polysilicon 1080 -1899 1080 -1899 0 1
rlabel polysilicon 1080 -1905 1080 -1905 0 3
rlabel polysilicon 1090 -1899 1090 -1899 0 2
rlabel polysilicon 1087 -1905 1087 -1905 0 3
rlabel polysilicon 1090 -1905 1090 -1905 0 4
rlabel polysilicon 1094 -1899 1094 -1899 0 1
rlabel polysilicon 1094 -1905 1094 -1905 0 3
rlabel polysilicon 1101 -1899 1101 -1899 0 1
rlabel polysilicon 1104 -1899 1104 -1899 0 2
rlabel polysilicon 1104 -1905 1104 -1905 0 4
rlabel polysilicon 1108 -1899 1108 -1899 0 1
rlabel polysilicon 1111 -1899 1111 -1899 0 2
rlabel polysilicon 1108 -1905 1108 -1905 0 3
rlabel polysilicon 1111 -1905 1111 -1905 0 4
rlabel polysilicon 1115 -1899 1115 -1899 0 1
rlabel polysilicon 1115 -1905 1115 -1905 0 3
rlabel polysilicon 1122 -1899 1122 -1899 0 1
rlabel polysilicon 1125 -1899 1125 -1899 0 2
rlabel polysilicon 1122 -1905 1122 -1905 0 3
rlabel polysilicon 1129 -1899 1129 -1899 0 1
rlabel polysilicon 1129 -1905 1129 -1905 0 3
rlabel polysilicon 1136 -1899 1136 -1899 0 1
rlabel polysilicon 1136 -1905 1136 -1905 0 3
rlabel polysilicon 1143 -1899 1143 -1899 0 1
rlabel polysilicon 1143 -1905 1143 -1905 0 3
rlabel polysilicon 1150 -1899 1150 -1899 0 1
rlabel polysilicon 1153 -1899 1153 -1899 0 2
rlabel polysilicon 1150 -1905 1150 -1905 0 3
rlabel polysilicon 1153 -1905 1153 -1905 0 4
rlabel polysilicon 1157 -1899 1157 -1899 0 1
rlabel polysilicon 1157 -1905 1157 -1905 0 3
rlabel polysilicon 1164 -1899 1164 -1899 0 1
rlabel polysilicon 1164 -1905 1164 -1905 0 3
rlabel polysilicon 1171 -1899 1171 -1899 0 1
rlabel polysilicon 1171 -1905 1171 -1905 0 3
rlabel polysilicon 1178 -1899 1178 -1899 0 1
rlabel polysilicon 1178 -1905 1178 -1905 0 3
rlabel polysilicon 1185 -1899 1185 -1899 0 1
rlabel polysilicon 1185 -1905 1185 -1905 0 3
rlabel polysilicon 1192 -1899 1192 -1899 0 1
rlabel polysilicon 1192 -1905 1192 -1905 0 3
rlabel polysilicon 1199 -1899 1199 -1899 0 1
rlabel polysilicon 1199 -1905 1199 -1905 0 3
rlabel polysilicon 1209 -1899 1209 -1899 0 2
rlabel polysilicon 1206 -1905 1206 -1905 0 3
rlabel polysilicon 1209 -1905 1209 -1905 0 4
rlabel polysilicon 1213 -1899 1213 -1899 0 1
rlabel polysilicon 1213 -1905 1213 -1905 0 3
rlabel polysilicon 1216 -1905 1216 -1905 0 4
rlabel polysilicon 1220 -1899 1220 -1899 0 1
rlabel polysilicon 1223 -1899 1223 -1899 0 2
rlabel polysilicon 1220 -1905 1220 -1905 0 3
rlabel polysilicon 1223 -1905 1223 -1905 0 4
rlabel polysilicon 1227 -1899 1227 -1899 0 1
rlabel polysilicon 1227 -1905 1227 -1905 0 3
rlabel polysilicon 1234 -1899 1234 -1899 0 1
rlabel polysilicon 1234 -1905 1234 -1905 0 3
rlabel polysilicon 1241 -1899 1241 -1899 0 1
rlabel polysilicon 1241 -1905 1241 -1905 0 3
rlabel polysilicon 1248 -1899 1248 -1899 0 1
rlabel polysilicon 1248 -1905 1248 -1905 0 3
rlabel polysilicon 1255 -1899 1255 -1899 0 1
rlabel polysilicon 1255 -1905 1255 -1905 0 3
rlabel polysilicon 1262 -1899 1262 -1899 0 1
rlabel polysilicon 1262 -1905 1262 -1905 0 3
rlabel polysilicon 1269 -1899 1269 -1899 0 1
rlabel polysilicon 1269 -1905 1269 -1905 0 3
rlabel polysilicon 1276 -1905 1276 -1905 0 3
rlabel polysilicon 1279 -1905 1279 -1905 0 4
rlabel polysilicon 1283 -1899 1283 -1899 0 1
rlabel polysilicon 1283 -1905 1283 -1905 0 3
rlabel polysilicon 1290 -1899 1290 -1899 0 1
rlabel polysilicon 1290 -1905 1290 -1905 0 3
rlabel polysilicon 1297 -1899 1297 -1899 0 1
rlabel polysilicon 1297 -1905 1297 -1905 0 3
rlabel polysilicon 1304 -1899 1304 -1899 0 1
rlabel polysilicon 1304 -1905 1304 -1905 0 3
rlabel polysilicon 1311 -1899 1311 -1899 0 1
rlabel polysilicon 1311 -1905 1311 -1905 0 3
rlabel polysilicon 1318 -1899 1318 -1899 0 1
rlabel polysilicon 1318 -1905 1318 -1905 0 3
rlabel polysilicon 1325 -1899 1325 -1899 0 1
rlabel polysilicon 1325 -1905 1325 -1905 0 3
rlabel polysilicon 1332 -1899 1332 -1899 0 1
rlabel polysilicon 1332 -1905 1332 -1905 0 3
rlabel polysilicon 1339 -1899 1339 -1899 0 1
rlabel polysilicon 1339 -1905 1339 -1905 0 3
rlabel polysilicon 1346 -1899 1346 -1899 0 1
rlabel polysilicon 1346 -1905 1346 -1905 0 3
rlabel polysilicon 1353 -1899 1353 -1899 0 1
rlabel polysilicon 1353 -1905 1353 -1905 0 3
rlabel polysilicon 1360 -1899 1360 -1899 0 1
rlabel polysilicon 1360 -1905 1360 -1905 0 3
rlabel polysilicon 1367 -1899 1367 -1899 0 1
rlabel polysilicon 1367 -1905 1367 -1905 0 3
rlabel polysilicon 1374 -1899 1374 -1899 0 1
rlabel polysilicon 1374 -1905 1374 -1905 0 3
rlabel polysilicon 1381 -1899 1381 -1899 0 1
rlabel polysilicon 1381 -1905 1381 -1905 0 3
rlabel polysilicon 1388 -1899 1388 -1899 0 1
rlabel polysilicon 1388 -1905 1388 -1905 0 3
rlabel polysilicon 1395 -1899 1395 -1899 0 1
rlabel polysilicon 1395 -1905 1395 -1905 0 3
rlabel polysilicon 1402 -1899 1402 -1899 0 1
rlabel polysilicon 1402 -1905 1402 -1905 0 3
rlabel polysilicon 1409 -1899 1409 -1899 0 1
rlabel polysilicon 1409 -1905 1409 -1905 0 3
rlabel polysilicon 1416 -1899 1416 -1899 0 1
rlabel polysilicon 1416 -1905 1416 -1905 0 3
rlabel polysilicon 1423 -1899 1423 -1899 0 1
rlabel polysilicon 1423 -1905 1423 -1905 0 3
rlabel polysilicon 1430 -1899 1430 -1899 0 1
rlabel polysilicon 1430 -1905 1430 -1905 0 3
rlabel polysilicon 1437 -1899 1437 -1899 0 1
rlabel polysilicon 1437 -1905 1437 -1905 0 3
rlabel polysilicon 1444 -1899 1444 -1899 0 1
rlabel polysilicon 1444 -1905 1444 -1905 0 3
rlabel polysilicon 1451 -1899 1451 -1899 0 1
rlabel polysilicon 1451 -1905 1451 -1905 0 3
rlabel polysilicon 1458 -1899 1458 -1899 0 1
rlabel polysilicon 1458 -1905 1458 -1905 0 3
rlabel polysilicon 1465 -1899 1465 -1899 0 1
rlabel polysilicon 1465 -1905 1465 -1905 0 3
rlabel polysilicon 1472 -1899 1472 -1899 0 1
rlabel polysilicon 1472 -1905 1472 -1905 0 3
rlabel polysilicon 1479 -1899 1479 -1899 0 1
rlabel polysilicon 1479 -1905 1479 -1905 0 3
rlabel polysilicon 1486 -1899 1486 -1899 0 1
rlabel polysilicon 1486 -1905 1486 -1905 0 3
rlabel polysilicon 1493 -1899 1493 -1899 0 1
rlabel polysilicon 1493 -1905 1493 -1905 0 3
rlabel polysilicon 1500 -1899 1500 -1899 0 1
rlabel polysilicon 1500 -1905 1500 -1905 0 3
rlabel polysilicon 1507 -1899 1507 -1899 0 1
rlabel polysilicon 1507 -1905 1507 -1905 0 3
rlabel polysilicon 1514 -1899 1514 -1899 0 1
rlabel polysilicon 1514 -1905 1514 -1905 0 3
rlabel polysilicon 1521 -1899 1521 -1899 0 1
rlabel polysilicon 1521 -1905 1521 -1905 0 3
rlabel polysilicon 1528 -1899 1528 -1899 0 1
rlabel polysilicon 1528 -1905 1528 -1905 0 3
rlabel polysilicon 1535 -1899 1535 -1899 0 1
rlabel polysilicon 1535 -1905 1535 -1905 0 3
rlabel polysilicon 1542 -1899 1542 -1899 0 1
rlabel polysilicon 1542 -1905 1542 -1905 0 3
rlabel polysilicon 1549 -1899 1549 -1899 0 1
rlabel polysilicon 1549 -1905 1549 -1905 0 3
rlabel polysilicon 1556 -1899 1556 -1899 0 1
rlabel polysilicon 1556 -1905 1556 -1905 0 3
rlabel polysilicon 1563 -1899 1563 -1899 0 1
rlabel polysilicon 1566 -1899 1566 -1899 0 2
rlabel polysilicon 1566 -1905 1566 -1905 0 4
rlabel polysilicon 1570 -1899 1570 -1899 0 1
rlabel polysilicon 1570 -1905 1570 -1905 0 3
rlabel polysilicon 1577 -1899 1577 -1899 0 1
rlabel polysilicon 1577 -1905 1577 -1905 0 3
rlabel polysilicon 1584 -1899 1584 -1899 0 1
rlabel polysilicon 1584 -1905 1584 -1905 0 3
rlabel polysilicon 1591 -1899 1591 -1899 0 1
rlabel polysilicon 1591 -1905 1591 -1905 0 3
rlabel polysilicon 1598 -1899 1598 -1899 0 1
rlabel polysilicon 1598 -1905 1598 -1905 0 3
rlabel polysilicon 1605 -1899 1605 -1899 0 1
rlabel polysilicon 1605 -1905 1605 -1905 0 3
rlabel polysilicon 1612 -1899 1612 -1899 0 1
rlabel polysilicon 1612 -1905 1612 -1905 0 3
rlabel polysilicon 1619 -1899 1619 -1899 0 1
rlabel polysilicon 1619 -1905 1619 -1905 0 3
rlabel polysilicon 1626 -1899 1626 -1899 0 1
rlabel polysilicon 1626 -1905 1626 -1905 0 3
rlabel polysilicon 1633 -1899 1633 -1899 0 1
rlabel polysilicon 1633 -1905 1633 -1905 0 3
rlabel polysilicon 1640 -1899 1640 -1899 0 1
rlabel polysilicon 1640 -1905 1640 -1905 0 3
rlabel polysilicon 1647 -1899 1647 -1899 0 1
rlabel polysilicon 1647 -1905 1647 -1905 0 3
rlabel polysilicon 1654 -1899 1654 -1899 0 1
rlabel polysilicon 1654 -1905 1654 -1905 0 3
rlabel polysilicon 1661 -1899 1661 -1899 0 1
rlabel polysilicon 1661 -1905 1661 -1905 0 3
rlabel polysilicon 1668 -1899 1668 -1899 0 1
rlabel polysilicon 1668 -1905 1668 -1905 0 3
rlabel polysilicon 1675 -1899 1675 -1899 0 1
rlabel polysilicon 1675 -1905 1675 -1905 0 3
rlabel polysilicon 1682 -1899 1682 -1899 0 1
rlabel polysilicon 1682 -1905 1682 -1905 0 3
rlabel polysilicon 1689 -1899 1689 -1899 0 1
rlabel polysilicon 1689 -1905 1689 -1905 0 3
rlabel polysilicon 1696 -1899 1696 -1899 0 1
rlabel polysilicon 1696 -1905 1696 -1905 0 3
rlabel polysilicon 1703 -1899 1703 -1899 0 1
rlabel polysilicon 1703 -1905 1703 -1905 0 3
rlabel polysilicon 1710 -1899 1710 -1899 0 1
rlabel polysilicon 1710 -1905 1710 -1905 0 3
rlabel polysilicon 1717 -1899 1717 -1899 0 1
rlabel polysilicon 1717 -1905 1717 -1905 0 3
rlabel polysilicon 1724 -1899 1724 -1899 0 1
rlabel polysilicon 1724 -1905 1724 -1905 0 3
rlabel polysilicon 1731 -1899 1731 -1899 0 1
rlabel polysilicon 1731 -1905 1731 -1905 0 3
rlabel polysilicon 1738 -1899 1738 -1899 0 1
rlabel polysilicon 1738 -1905 1738 -1905 0 3
rlabel polysilicon 1745 -1899 1745 -1899 0 1
rlabel polysilicon 1745 -1905 1745 -1905 0 3
rlabel polysilicon 1752 -1899 1752 -1899 0 1
rlabel polysilicon 1752 -1905 1752 -1905 0 3
rlabel polysilicon 1759 -1899 1759 -1899 0 1
rlabel polysilicon 1759 -1905 1759 -1905 0 3
rlabel polysilicon 1766 -1899 1766 -1899 0 1
rlabel polysilicon 1766 -1905 1766 -1905 0 3
rlabel polysilicon 1773 -1899 1773 -1899 0 1
rlabel polysilicon 1773 -1905 1773 -1905 0 3
rlabel polysilicon 1780 -1899 1780 -1899 0 1
rlabel polysilicon 1780 -1905 1780 -1905 0 3
rlabel polysilicon 1787 -1899 1787 -1899 0 1
rlabel polysilicon 1787 -1905 1787 -1905 0 3
rlabel polysilicon 1794 -1899 1794 -1899 0 1
rlabel polysilicon 1794 -1905 1794 -1905 0 3
rlabel polysilicon 1801 -1899 1801 -1899 0 1
rlabel polysilicon 1801 -1905 1801 -1905 0 3
rlabel polysilicon 1808 -1899 1808 -1899 0 1
rlabel polysilicon 1808 -1905 1808 -1905 0 3
rlabel polysilicon 1815 -1899 1815 -1899 0 1
rlabel polysilicon 1815 -1905 1815 -1905 0 3
rlabel polysilicon 1822 -1899 1822 -1899 0 1
rlabel polysilicon 1822 -1905 1822 -1905 0 3
rlabel polysilicon 1829 -1899 1829 -1899 0 1
rlabel polysilicon 1829 -1905 1829 -1905 0 3
rlabel polysilicon 1836 -1899 1836 -1899 0 1
rlabel polysilicon 1836 -1905 1836 -1905 0 3
rlabel polysilicon 1843 -1899 1843 -1899 0 1
rlabel polysilicon 1843 -1905 1843 -1905 0 3
rlabel polysilicon 1850 -1899 1850 -1899 0 1
rlabel polysilicon 1850 -1905 1850 -1905 0 3
rlabel polysilicon 1857 -1899 1857 -1899 0 1
rlabel polysilicon 1857 -1905 1857 -1905 0 3
rlabel polysilicon 1864 -1899 1864 -1899 0 1
rlabel polysilicon 1864 -1905 1864 -1905 0 3
rlabel polysilicon 1871 -1899 1871 -1899 0 1
rlabel polysilicon 1871 -1905 1871 -1905 0 3
rlabel polysilicon 1878 -1899 1878 -1899 0 1
rlabel polysilicon 1878 -1905 1878 -1905 0 3
rlabel polysilicon 1885 -1899 1885 -1899 0 1
rlabel polysilicon 1885 -1905 1885 -1905 0 3
rlabel polysilicon 1892 -1899 1892 -1899 0 1
rlabel polysilicon 1892 -1905 1892 -1905 0 3
rlabel polysilicon 1899 -1899 1899 -1899 0 1
rlabel polysilicon 1899 -1905 1899 -1905 0 3
rlabel polysilicon 1906 -1899 1906 -1899 0 1
rlabel polysilicon 1906 -1905 1906 -1905 0 3
rlabel polysilicon 1913 -1899 1913 -1899 0 1
rlabel polysilicon 1913 -1905 1913 -1905 0 3
rlabel polysilicon 1920 -1899 1920 -1899 0 1
rlabel polysilicon 1920 -1905 1920 -1905 0 3
rlabel polysilicon 1927 -1899 1927 -1899 0 1
rlabel polysilicon 1927 -1905 1927 -1905 0 3
rlabel polysilicon 1934 -1899 1934 -1899 0 1
rlabel polysilicon 1934 -1905 1934 -1905 0 3
rlabel polysilicon 1941 -1899 1941 -1899 0 1
rlabel polysilicon 1941 -1905 1941 -1905 0 3
rlabel polysilicon 1948 -1899 1948 -1899 0 1
rlabel polysilicon 1948 -1905 1948 -1905 0 3
rlabel polysilicon 1955 -1899 1955 -1899 0 1
rlabel polysilicon 1955 -1905 1955 -1905 0 3
rlabel polysilicon 1962 -1899 1962 -1899 0 1
rlabel polysilicon 1962 -1905 1962 -1905 0 3
rlabel polysilicon 1969 -1899 1969 -1899 0 1
rlabel polysilicon 1969 -1905 1969 -1905 0 3
rlabel polysilicon 1976 -1899 1976 -1899 0 1
rlabel polysilicon 1976 -1905 1976 -1905 0 3
rlabel polysilicon 1983 -1899 1983 -1899 0 1
rlabel polysilicon 1983 -1905 1983 -1905 0 3
rlabel polysilicon 1990 -1899 1990 -1899 0 1
rlabel polysilicon 1990 -1905 1990 -1905 0 3
rlabel polysilicon 1997 -1899 1997 -1899 0 1
rlabel polysilicon 1997 -1905 1997 -1905 0 3
rlabel polysilicon 2004 -1899 2004 -1899 0 1
rlabel polysilicon 2004 -1905 2004 -1905 0 3
rlabel polysilicon 2011 -1899 2011 -1899 0 1
rlabel polysilicon 2014 -1899 2014 -1899 0 2
rlabel polysilicon 2011 -1905 2011 -1905 0 3
rlabel polysilicon 2018 -1899 2018 -1899 0 1
rlabel polysilicon 2018 -1905 2018 -1905 0 3
rlabel polysilicon 2025 -1899 2025 -1899 0 1
rlabel polysilicon 2025 -1905 2025 -1905 0 3
rlabel polysilicon 2 -2046 2 -2046 0 1
rlabel polysilicon 2 -2052 2 -2052 0 3
rlabel polysilicon 9 -2046 9 -2046 0 1
rlabel polysilicon 9 -2052 9 -2052 0 3
rlabel polysilicon 16 -2046 16 -2046 0 1
rlabel polysilicon 16 -2052 16 -2052 0 3
rlabel polysilicon 23 -2046 23 -2046 0 1
rlabel polysilicon 23 -2052 23 -2052 0 3
rlabel polysilicon 30 -2046 30 -2046 0 1
rlabel polysilicon 30 -2052 30 -2052 0 3
rlabel polysilicon 37 -2046 37 -2046 0 1
rlabel polysilicon 37 -2052 37 -2052 0 3
rlabel polysilicon 44 -2046 44 -2046 0 1
rlabel polysilicon 44 -2052 44 -2052 0 3
rlabel polysilicon 51 -2046 51 -2046 0 1
rlabel polysilicon 51 -2052 51 -2052 0 3
rlabel polysilicon 58 -2046 58 -2046 0 1
rlabel polysilicon 58 -2052 58 -2052 0 3
rlabel polysilicon 68 -2046 68 -2046 0 2
rlabel polysilicon 65 -2052 65 -2052 0 3
rlabel polysilicon 68 -2052 68 -2052 0 4
rlabel polysilicon 72 -2046 72 -2046 0 1
rlabel polysilicon 72 -2052 72 -2052 0 3
rlabel polysilicon 79 -2046 79 -2046 0 1
rlabel polysilicon 79 -2052 79 -2052 0 3
rlabel polysilicon 86 -2046 86 -2046 0 1
rlabel polysilicon 86 -2052 86 -2052 0 3
rlabel polysilicon 93 -2046 93 -2046 0 1
rlabel polysilicon 93 -2052 93 -2052 0 3
rlabel polysilicon 100 -2046 100 -2046 0 1
rlabel polysilicon 100 -2052 100 -2052 0 3
rlabel polysilicon 107 -2046 107 -2046 0 1
rlabel polysilicon 107 -2052 107 -2052 0 3
rlabel polysilicon 114 -2046 114 -2046 0 1
rlabel polysilicon 114 -2052 114 -2052 0 3
rlabel polysilicon 117 -2052 117 -2052 0 4
rlabel polysilicon 121 -2046 121 -2046 0 1
rlabel polysilicon 121 -2052 121 -2052 0 3
rlabel polysilicon 128 -2046 128 -2046 0 1
rlabel polysilicon 128 -2052 128 -2052 0 3
rlabel polysilicon 135 -2046 135 -2046 0 1
rlabel polysilicon 135 -2052 135 -2052 0 3
rlabel polysilicon 142 -2046 142 -2046 0 1
rlabel polysilicon 145 -2046 145 -2046 0 2
rlabel polysilicon 142 -2052 142 -2052 0 3
rlabel polysilicon 145 -2052 145 -2052 0 4
rlabel polysilicon 149 -2046 149 -2046 0 1
rlabel polysilicon 149 -2052 149 -2052 0 3
rlabel polysilicon 156 -2046 156 -2046 0 1
rlabel polysilicon 156 -2052 156 -2052 0 3
rlabel polysilicon 163 -2046 163 -2046 0 1
rlabel polysilicon 163 -2052 163 -2052 0 3
rlabel polysilicon 170 -2046 170 -2046 0 1
rlabel polysilicon 170 -2052 170 -2052 0 3
rlabel polysilicon 177 -2046 177 -2046 0 1
rlabel polysilicon 177 -2052 177 -2052 0 3
rlabel polysilicon 184 -2046 184 -2046 0 1
rlabel polysilicon 184 -2052 184 -2052 0 3
rlabel polysilicon 191 -2046 191 -2046 0 1
rlabel polysilicon 191 -2052 191 -2052 0 3
rlabel polysilicon 198 -2046 198 -2046 0 1
rlabel polysilicon 198 -2052 198 -2052 0 3
rlabel polysilicon 205 -2046 205 -2046 0 1
rlabel polysilicon 205 -2052 205 -2052 0 3
rlabel polysilicon 212 -2046 212 -2046 0 1
rlabel polysilicon 212 -2052 212 -2052 0 3
rlabel polysilicon 219 -2046 219 -2046 0 1
rlabel polysilicon 222 -2046 222 -2046 0 2
rlabel polysilicon 219 -2052 219 -2052 0 3
rlabel polysilicon 222 -2052 222 -2052 0 4
rlabel polysilicon 226 -2046 226 -2046 0 1
rlabel polysilicon 226 -2052 226 -2052 0 3
rlabel polysilicon 233 -2046 233 -2046 0 1
rlabel polysilicon 233 -2052 233 -2052 0 3
rlabel polysilicon 243 -2046 243 -2046 0 2
rlabel polysilicon 243 -2052 243 -2052 0 4
rlabel polysilicon 247 -2046 247 -2046 0 1
rlabel polysilicon 247 -2052 247 -2052 0 3
rlabel polysilicon 254 -2046 254 -2046 0 1
rlabel polysilicon 254 -2052 254 -2052 0 3
rlabel polysilicon 261 -2046 261 -2046 0 1
rlabel polysilicon 261 -2052 261 -2052 0 3
rlabel polysilicon 268 -2046 268 -2046 0 1
rlabel polysilicon 268 -2052 268 -2052 0 3
rlabel polysilicon 275 -2046 275 -2046 0 1
rlabel polysilicon 275 -2052 275 -2052 0 3
rlabel polysilicon 282 -2046 282 -2046 0 1
rlabel polysilicon 282 -2052 282 -2052 0 3
rlabel polysilicon 289 -2046 289 -2046 0 1
rlabel polysilicon 289 -2052 289 -2052 0 3
rlabel polysilicon 296 -2046 296 -2046 0 1
rlabel polysilicon 296 -2052 296 -2052 0 3
rlabel polysilicon 303 -2046 303 -2046 0 1
rlabel polysilicon 303 -2052 303 -2052 0 3
rlabel polysilicon 310 -2046 310 -2046 0 1
rlabel polysilicon 313 -2046 313 -2046 0 2
rlabel polysilicon 310 -2052 310 -2052 0 3
rlabel polysilicon 313 -2052 313 -2052 0 4
rlabel polysilicon 317 -2046 317 -2046 0 1
rlabel polysilicon 317 -2052 317 -2052 0 3
rlabel polysilicon 324 -2046 324 -2046 0 1
rlabel polysilicon 324 -2052 324 -2052 0 3
rlabel polysilicon 331 -2046 331 -2046 0 1
rlabel polysilicon 331 -2052 331 -2052 0 3
rlabel polysilicon 341 -2046 341 -2046 0 2
rlabel polysilicon 338 -2052 338 -2052 0 3
rlabel polysilicon 345 -2046 345 -2046 0 1
rlabel polysilicon 345 -2052 345 -2052 0 3
rlabel polysilicon 352 -2046 352 -2046 0 1
rlabel polysilicon 352 -2052 352 -2052 0 3
rlabel polysilicon 359 -2046 359 -2046 0 1
rlabel polysilicon 359 -2052 359 -2052 0 3
rlabel polysilicon 366 -2046 366 -2046 0 1
rlabel polysilicon 366 -2052 366 -2052 0 3
rlabel polysilicon 373 -2046 373 -2046 0 1
rlabel polysilicon 373 -2052 373 -2052 0 3
rlabel polysilicon 380 -2046 380 -2046 0 1
rlabel polysilicon 380 -2052 380 -2052 0 3
rlabel polysilicon 387 -2046 387 -2046 0 1
rlabel polysilicon 387 -2052 387 -2052 0 3
rlabel polysilicon 394 -2046 394 -2046 0 1
rlabel polysilicon 394 -2052 394 -2052 0 3
rlabel polysilicon 401 -2046 401 -2046 0 1
rlabel polysilicon 401 -2052 401 -2052 0 3
rlabel polysilicon 408 -2046 408 -2046 0 1
rlabel polysilicon 408 -2052 408 -2052 0 3
rlabel polysilicon 415 -2046 415 -2046 0 1
rlabel polysilicon 415 -2052 415 -2052 0 3
rlabel polysilicon 422 -2046 422 -2046 0 1
rlabel polysilicon 422 -2052 422 -2052 0 3
rlabel polysilicon 429 -2046 429 -2046 0 1
rlabel polysilicon 429 -2052 429 -2052 0 3
rlabel polysilicon 436 -2046 436 -2046 0 1
rlabel polysilicon 436 -2052 436 -2052 0 3
rlabel polysilicon 443 -2046 443 -2046 0 1
rlabel polysilicon 443 -2052 443 -2052 0 3
rlabel polysilicon 450 -2052 450 -2052 0 3
rlabel polysilicon 453 -2052 453 -2052 0 4
rlabel polysilicon 457 -2046 457 -2046 0 1
rlabel polysilicon 457 -2052 457 -2052 0 3
rlabel polysilicon 464 -2046 464 -2046 0 1
rlabel polysilicon 464 -2052 464 -2052 0 3
rlabel polysilicon 471 -2046 471 -2046 0 1
rlabel polysilicon 471 -2052 471 -2052 0 3
rlabel polysilicon 478 -2046 478 -2046 0 1
rlabel polysilicon 478 -2052 478 -2052 0 3
rlabel polysilicon 485 -2046 485 -2046 0 1
rlabel polysilicon 485 -2052 485 -2052 0 3
rlabel polysilicon 492 -2046 492 -2046 0 1
rlabel polysilicon 492 -2052 492 -2052 0 3
rlabel polysilicon 499 -2046 499 -2046 0 1
rlabel polysilicon 499 -2052 499 -2052 0 3
rlabel polysilicon 506 -2046 506 -2046 0 1
rlabel polysilicon 506 -2052 506 -2052 0 3
rlabel polysilicon 513 -2046 513 -2046 0 1
rlabel polysilicon 513 -2052 513 -2052 0 3
rlabel polysilicon 520 -2046 520 -2046 0 1
rlabel polysilicon 520 -2052 520 -2052 0 3
rlabel polysilicon 527 -2046 527 -2046 0 1
rlabel polysilicon 530 -2046 530 -2046 0 2
rlabel polysilicon 527 -2052 527 -2052 0 3
rlabel polysilicon 530 -2052 530 -2052 0 4
rlabel polysilicon 534 -2046 534 -2046 0 1
rlabel polysilicon 537 -2046 537 -2046 0 2
rlabel polysilicon 534 -2052 534 -2052 0 3
rlabel polysilicon 537 -2052 537 -2052 0 4
rlabel polysilicon 541 -2046 541 -2046 0 1
rlabel polysilicon 541 -2052 541 -2052 0 3
rlabel polysilicon 548 -2046 548 -2046 0 1
rlabel polysilicon 548 -2052 548 -2052 0 3
rlabel polysilicon 555 -2046 555 -2046 0 1
rlabel polysilicon 555 -2052 555 -2052 0 3
rlabel polysilicon 562 -2046 562 -2046 0 1
rlabel polysilicon 562 -2052 562 -2052 0 3
rlabel polysilicon 569 -2046 569 -2046 0 1
rlabel polysilicon 569 -2052 569 -2052 0 3
rlabel polysilicon 576 -2046 576 -2046 0 1
rlabel polysilicon 576 -2052 576 -2052 0 3
rlabel polysilicon 583 -2046 583 -2046 0 1
rlabel polysilicon 583 -2052 583 -2052 0 3
rlabel polysilicon 590 -2046 590 -2046 0 1
rlabel polysilicon 590 -2052 590 -2052 0 3
rlabel polysilicon 597 -2046 597 -2046 0 1
rlabel polysilicon 597 -2052 597 -2052 0 3
rlabel polysilicon 604 -2046 604 -2046 0 1
rlabel polysilicon 604 -2052 604 -2052 0 3
rlabel polysilicon 611 -2046 611 -2046 0 1
rlabel polysilicon 611 -2052 611 -2052 0 3
rlabel polysilicon 618 -2046 618 -2046 0 1
rlabel polysilicon 618 -2052 618 -2052 0 3
rlabel polysilicon 625 -2046 625 -2046 0 1
rlabel polysilicon 625 -2052 625 -2052 0 3
rlabel polysilicon 632 -2046 632 -2046 0 1
rlabel polysilicon 632 -2052 632 -2052 0 3
rlabel polysilicon 639 -2046 639 -2046 0 1
rlabel polysilicon 639 -2052 639 -2052 0 3
rlabel polysilicon 646 -2046 646 -2046 0 1
rlabel polysilicon 646 -2052 646 -2052 0 3
rlabel polysilicon 653 -2046 653 -2046 0 1
rlabel polysilicon 653 -2052 653 -2052 0 3
rlabel polysilicon 660 -2046 660 -2046 0 1
rlabel polysilicon 660 -2052 660 -2052 0 3
rlabel polysilicon 667 -2052 667 -2052 0 3
rlabel polysilicon 674 -2046 674 -2046 0 1
rlabel polysilicon 674 -2052 674 -2052 0 3
rlabel polysilicon 681 -2046 681 -2046 0 1
rlabel polysilicon 681 -2052 681 -2052 0 3
rlabel polysilicon 688 -2046 688 -2046 0 1
rlabel polysilicon 688 -2052 688 -2052 0 3
rlabel polysilicon 698 -2046 698 -2046 0 2
rlabel polysilicon 695 -2052 695 -2052 0 3
rlabel polysilicon 698 -2052 698 -2052 0 4
rlabel polysilicon 702 -2046 702 -2046 0 1
rlabel polysilicon 702 -2052 702 -2052 0 3
rlabel polysilicon 709 -2046 709 -2046 0 1
rlabel polysilicon 709 -2052 709 -2052 0 3
rlabel polysilicon 716 -2046 716 -2046 0 1
rlabel polysilicon 716 -2052 716 -2052 0 3
rlabel polysilicon 723 -2046 723 -2046 0 1
rlabel polysilicon 723 -2052 723 -2052 0 3
rlabel polysilicon 726 -2052 726 -2052 0 4
rlabel polysilicon 730 -2046 730 -2046 0 1
rlabel polysilicon 733 -2046 733 -2046 0 2
rlabel polysilicon 730 -2052 730 -2052 0 3
rlabel polysilicon 733 -2052 733 -2052 0 4
rlabel polysilicon 737 -2046 737 -2046 0 1
rlabel polysilicon 737 -2052 737 -2052 0 3
rlabel polysilicon 744 -2046 744 -2046 0 1
rlabel polysilicon 744 -2052 744 -2052 0 3
rlabel polysilicon 751 -2046 751 -2046 0 1
rlabel polysilicon 754 -2046 754 -2046 0 2
rlabel polysilicon 751 -2052 751 -2052 0 3
rlabel polysilicon 754 -2052 754 -2052 0 4
rlabel polysilicon 758 -2046 758 -2046 0 1
rlabel polysilicon 761 -2046 761 -2046 0 2
rlabel polysilicon 758 -2052 758 -2052 0 3
rlabel polysilicon 761 -2052 761 -2052 0 4
rlabel polysilicon 765 -2046 765 -2046 0 1
rlabel polysilicon 765 -2052 765 -2052 0 3
rlabel polysilicon 772 -2046 772 -2046 0 1
rlabel polysilicon 775 -2046 775 -2046 0 2
rlabel polysilicon 772 -2052 772 -2052 0 3
rlabel polysilicon 779 -2046 779 -2046 0 1
rlabel polysilicon 779 -2052 779 -2052 0 3
rlabel polysilicon 786 -2046 786 -2046 0 1
rlabel polysilicon 786 -2052 786 -2052 0 3
rlabel polysilicon 793 -2046 793 -2046 0 1
rlabel polysilicon 793 -2052 793 -2052 0 3
rlabel polysilicon 800 -2046 800 -2046 0 1
rlabel polysilicon 800 -2052 800 -2052 0 3
rlabel polysilicon 807 -2046 807 -2046 0 1
rlabel polysilicon 807 -2052 807 -2052 0 3
rlabel polysilicon 814 -2046 814 -2046 0 1
rlabel polysilicon 817 -2046 817 -2046 0 2
rlabel polysilicon 814 -2052 814 -2052 0 3
rlabel polysilicon 817 -2052 817 -2052 0 4
rlabel polysilicon 821 -2046 821 -2046 0 1
rlabel polysilicon 821 -2052 821 -2052 0 3
rlabel polysilicon 828 -2046 828 -2046 0 1
rlabel polysilicon 828 -2052 828 -2052 0 3
rlabel polysilicon 835 -2046 835 -2046 0 1
rlabel polysilicon 835 -2052 835 -2052 0 3
rlabel polysilicon 842 -2046 842 -2046 0 1
rlabel polysilicon 845 -2046 845 -2046 0 2
rlabel polysilicon 842 -2052 842 -2052 0 3
rlabel polysilicon 845 -2052 845 -2052 0 4
rlabel polysilicon 849 -2046 849 -2046 0 1
rlabel polysilicon 849 -2052 849 -2052 0 3
rlabel polysilicon 852 -2052 852 -2052 0 4
rlabel polysilicon 856 -2046 856 -2046 0 1
rlabel polysilicon 856 -2052 856 -2052 0 3
rlabel polysilicon 863 -2046 863 -2046 0 1
rlabel polysilicon 866 -2046 866 -2046 0 2
rlabel polysilicon 863 -2052 863 -2052 0 3
rlabel polysilicon 866 -2052 866 -2052 0 4
rlabel polysilicon 870 -2046 870 -2046 0 1
rlabel polysilicon 870 -2052 870 -2052 0 3
rlabel polysilicon 877 -2046 877 -2046 0 1
rlabel polysilicon 880 -2046 880 -2046 0 2
rlabel polysilicon 877 -2052 877 -2052 0 3
rlabel polysilicon 880 -2052 880 -2052 0 4
rlabel polysilicon 884 -2046 884 -2046 0 1
rlabel polysilicon 884 -2052 884 -2052 0 3
rlabel polysilicon 891 -2046 891 -2046 0 1
rlabel polysilicon 894 -2046 894 -2046 0 2
rlabel polysilicon 891 -2052 891 -2052 0 3
rlabel polysilicon 894 -2052 894 -2052 0 4
rlabel polysilicon 898 -2046 898 -2046 0 1
rlabel polysilicon 898 -2052 898 -2052 0 3
rlabel polysilicon 905 -2046 905 -2046 0 1
rlabel polysilicon 905 -2052 905 -2052 0 3
rlabel polysilicon 912 -2046 912 -2046 0 1
rlabel polysilicon 912 -2052 912 -2052 0 3
rlabel polysilicon 919 -2046 919 -2046 0 1
rlabel polysilicon 922 -2046 922 -2046 0 2
rlabel polysilicon 919 -2052 919 -2052 0 3
rlabel polysilicon 922 -2052 922 -2052 0 4
rlabel polysilicon 926 -2046 926 -2046 0 1
rlabel polysilicon 926 -2052 926 -2052 0 3
rlabel polysilicon 933 -2046 933 -2046 0 1
rlabel polysilicon 933 -2052 933 -2052 0 3
rlabel polysilicon 940 -2046 940 -2046 0 1
rlabel polysilicon 940 -2052 940 -2052 0 3
rlabel polysilicon 947 -2046 947 -2046 0 1
rlabel polysilicon 947 -2052 947 -2052 0 3
rlabel polysilicon 954 -2046 954 -2046 0 1
rlabel polysilicon 954 -2052 954 -2052 0 3
rlabel polysilicon 961 -2046 961 -2046 0 1
rlabel polysilicon 964 -2046 964 -2046 0 2
rlabel polysilicon 961 -2052 961 -2052 0 3
rlabel polysilicon 964 -2052 964 -2052 0 4
rlabel polysilicon 968 -2046 968 -2046 0 1
rlabel polysilicon 968 -2052 968 -2052 0 3
rlabel polysilicon 971 -2052 971 -2052 0 4
rlabel polysilicon 975 -2046 975 -2046 0 1
rlabel polysilicon 975 -2052 975 -2052 0 3
rlabel polysilicon 982 -2046 982 -2046 0 1
rlabel polysilicon 982 -2052 982 -2052 0 3
rlabel polysilicon 989 -2046 989 -2046 0 1
rlabel polysilicon 989 -2052 989 -2052 0 3
rlabel polysilicon 996 -2046 996 -2046 0 1
rlabel polysilicon 996 -2052 996 -2052 0 3
rlabel polysilicon 1003 -2046 1003 -2046 0 1
rlabel polysilicon 1003 -2052 1003 -2052 0 3
rlabel polysilicon 1010 -2046 1010 -2046 0 1
rlabel polysilicon 1010 -2052 1010 -2052 0 3
rlabel polysilicon 1017 -2046 1017 -2046 0 1
rlabel polysilicon 1017 -2052 1017 -2052 0 3
rlabel polysilicon 1024 -2046 1024 -2046 0 1
rlabel polysilicon 1024 -2052 1024 -2052 0 3
rlabel polysilicon 1031 -2046 1031 -2046 0 1
rlabel polysilicon 1031 -2052 1031 -2052 0 3
rlabel polysilicon 1038 -2046 1038 -2046 0 1
rlabel polysilicon 1038 -2052 1038 -2052 0 3
rlabel polysilicon 1045 -2046 1045 -2046 0 1
rlabel polysilicon 1045 -2052 1045 -2052 0 3
rlabel polysilicon 1052 -2046 1052 -2046 0 1
rlabel polysilicon 1052 -2052 1052 -2052 0 3
rlabel polysilicon 1059 -2046 1059 -2046 0 1
rlabel polysilicon 1059 -2052 1059 -2052 0 3
rlabel polysilicon 1066 -2046 1066 -2046 0 1
rlabel polysilicon 1066 -2052 1066 -2052 0 3
rlabel polysilicon 1073 -2046 1073 -2046 0 1
rlabel polysilicon 1073 -2052 1073 -2052 0 3
rlabel polysilicon 1080 -2046 1080 -2046 0 1
rlabel polysilicon 1080 -2052 1080 -2052 0 3
rlabel polysilicon 1087 -2046 1087 -2046 0 1
rlabel polysilicon 1087 -2052 1087 -2052 0 3
rlabel polysilicon 1090 -2052 1090 -2052 0 4
rlabel polysilicon 1094 -2046 1094 -2046 0 1
rlabel polysilicon 1094 -2052 1094 -2052 0 3
rlabel polysilicon 1101 -2046 1101 -2046 0 1
rlabel polysilicon 1101 -2052 1101 -2052 0 3
rlabel polysilicon 1108 -2046 1108 -2046 0 1
rlabel polysilicon 1111 -2046 1111 -2046 0 2
rlabel polysilicon 1108 -2052 1108 -2052 0 3
rlabel polysilicon 1111 -2052 1111 -2052 0 4
rlabel polysilicon 1115 -2046 1115 -2046 0 1
rlabel polysilicon 1115 -2052 1115 -2052 0 3
rlabel polysilicon 1122 -2046 1122 -2046 0 1
rlabel polysilicon 1122 -2052 1122 -2052 0 3
rlabel polysilicon 1129 -2046 1129 -2046 0 1
rlabel polysilicon 1129 -2052 1129 -2052 0 3
rlabel polysilicon 1136 -2046 1136 -2046 0 1
rlabel polysilicon 1136 -2052 1136 -2052 0 3
rlabel polysilicon 1143 -2046 1143 -2046 0 1
rlabel polysilicon 1143 -2052 1143 -2052 0 3
rlabel polysilicon 1150 -2046 1150 -2046 0 1
rlabel polysilicon 1150 -2052 1150 -2052 0 3
rlabel polysilicon 1157 -2046 1157 -2046 0 1
rlabel polysilicon 1157 -2052 1157 -2052 0 3
rlabel polysilicon 1164 -2046 1164 -2046 0 1
rlabel polysilicon 1164 -2052 1164 -2052 0 3
rlabel polysilicon 1171 -2046 1171 -2046 0 1
rlabel polysilicon 1171 -2052 1171 -2052 0 3
rlabel polysilicon 1178 -2046 1178 -2046 0 1
rlabel polysilicon 1178 -2052 1178 -2052 0 3
rlabel polysilicon 1185 -2046 1185 -2046 0 1
rlabel polysilicon 1185 -2052 1185 -2052 0 3
rlabel polysilicon 1192 -2046 1192 -2046 0 1
rlabel polysilicon 1192 -2052 1192 -2052 0 3
rlabel polysilicon 1199 -2046 1199 -2046 0 1
rlabel polysilicon 1199 -2052 1199 -2052 0 3
rlabel polysilicon 1206 -2046 1206 -2046 0 1
rlabel polysilicon 1206 -2052 1206 -2052 0 3
rlabel polysilicon 1213 -2046 1213 -2046 0 1
rlabel polysilicon 1216 -2046 1216 -2046 0 2
rlabel polysilicon 1213 -2052 1213 -2052 0 3
rlabel polysilicon 1220 -2046 1220 -2046 0 1
rlabel polysilicon 1220 -2052 1220 -2052 0 3
rlabel polysilicon 1227 -2046 1227 -2046 0 1
rlabel polysilicon 1227 -2052 1227 -2052 0 3
rlabel polysilicon 1237 -2046 1237 -2046 0 2
rlabel polysilicon 1237 -2052 1237 -2052 0 4
rlabel polysilicon 1241 -2046 1241 -2046 0 1
rlabel polysilicon 1241 -2052 1241 -2052 0 3
rlabel polysilicon 1248 -2046 1248 -2046 0 1
rlabel polysilicon 1248 -2052 1248 -2052 0 3
rlabel polysilicon 1255 -2046 1255 -2046 0 1
rlabel polysilicon 1255 -2052 1255 -2052 0 3
rlabel polysilicon 1262 -2046 1262 -2046 0 1
rlabel polysilicon 1265 -2046 1265 -2046 0 2
rlabel polysilicon 1262 -2052 1262 -2052 0 3
rlabel polysilicon 1265 -2052 1265 -2052 0 4
rlabel polysilicon 1269 -2046 1269 -2046 0 1
rlabel polysilicon 1269 -2052 1269 -2052 0 3
rlabel polysilicon 1276 -2046 1276 -2046 0 1
rlabel polysilicon 1276 -2052 1276 -2052 0 3
rlabel polysilicon 1283 -2046 1283 -2046 0 1
rlabel polysilicon 1283 -2052 1283 -2052 0 3
rlabel polysilicon 1290 -2046 1290 -2046 0 1
rlabel polysilicon 1293 -2046 1293 -2046 0 2
rlabel polysilicon 1293 -2052 1293 -2052 0 4
rlabel polysilicon 1297 -2046 1297 -2046 0 1
rlabel polysilicon 1297 -2052 1297 -2052 0 3
rlabel polysilicon 1304 -2046 1304 -2046 0 1
rlabel polysilicon 1304 -2052 1304 -2052 0 3
rlabel polysilicon 1311 -2046 1311 -2046 0 1
rlabel polysilicon 1311 -2052 1311 -2052 0 3
rlabel polysilicon 1318 -2046 1318 -2046 0 1
rlabel polysilicon 1318 -2052 1318 -2052 0 3
rlabel polysilicon 1325 -2046 1325 -2046 0 1
rlabel polysilicon 1325 -2052 1325 -2052 0 3
rlabel polysilicon 1332 -2046 1332 -2046 0 1
rlabel polysilicon 1332 -2052 1332 -2052 0 3
rlabel polysilicon 1339 -2046 1339 -2046 0 1
rlabel polysilicon 1339 -2052 1339 -2052 0 3
rlabel polysilicon 1346 -2046 1346 -2046 0 1
rlabel polysilicon 1346 -2052 1346 -2052 0 3
rlabel polysilicon 1353 -2046 1353 -2046 0 1
rlabel polysilicon 1353 -2052 1353 -2052 0 3
rlabel polysilicon 1360 -2046 1360 -2046 0 1
rlabel polysilicon 1360 -2052 1360 -2052 0 3
rlabel polysilicon 1367 -2046 1367 -2046 0 1
rlabel polysilicon 1367 -2052 1367 -2052 0 3
rlabel polysilicon 1374 -2046 1374 -2046 0 1
rlabel polysilicon 1374 -2052 1374 -2052 0 3
rlabel polysilicon 1381 -2046 1381 -2046 0 1
rlabel polysilicon 1381 -2052 1381 -2052 0 3
rlabel polysilicon 1388 -2046 1388 -2046 0 1
rlabel polysilicon 1388 -2052 1388 -2052 0 3
rlabel polysilicon 1395 -2046 1395 -2046 0 1
rlabel polysilicon 1395 -2052 1395 -2052 0 3
rlabel polysilicon 1402 -2046 1402 -2046 0 1
rlabel polysilicon 1402 -2052 1402 -2052 0 3
rlabel polysilicon 1409 -2046 1409 -2046 0 1
rlabel polysilicon 1409 -2052 1409 -2052 0 3
rlabel polysilicon 1416 -2046 1416 -2046 0 1
rlabel polysilicon 1416 -2052 1416 -2052 0 3
rlabel polysilicon 1423 -2046 1423 -2046 0 1
rlabel polysilicon 1423 -2052 1423 -2052 0 3
rlabel polysilicon 1430 -2046 1430 -2046 0 1
rlabel polysilicon 1430 -2052 1430 -2052 0 3
rlabel polysilicon 1437 -2046 1437 -2046 0 1
rlabel polysilicon 1437 -2052 1437 -2052 0 3
rlabel polysilicon 1444 -2046 1444 -2046 0 1
rlabel polysilicon 1444 -2052 1444 -2052 0 3
rlabel polysilicon 1451 -2046 1451 -2046 0 1
rlabel polysilicon 1454 -2046 1454 -2046 0 2
rlabel polysilicon 1451 -2052 1451 -2052 0 3
rlabel polysilicon 1458 -2046 1458 -2046 0 1
rlabel polysilicon 1458 -2052 1458 -2052 0 3
rlabel polysilicon 1465 -2046 1465 -2046 0 1
rlabel polysilicon 1465 -2052 1465 -2052 0 3
rlabel polysilicon 1472 -2046 1472 -2046 0 1
rlabel polysilicon 1472 -2052 1472 -2052 0 3
rlabel polysilicon 1479 -2046 1479 -2046 0 1
rlabel polysilicon 1479 -2052 1479 -2052 0 3
rlabel polysilicon 1486 -2046 1486 -2046 0 1
rlabel polysilicon 1486 -2052 1486 -2052 0 3
rlabel polysilicon 1493 -2046 1493 -2046 0 1
rlabel polysilicon 1493 -2052 1493 -2052 0 3
rlabel polysilicon 1500 -2046 1500 -2046 0 1
rlabel polysilicon 1500 -2052 1500 -2052 0 3
rlabel polysilicon 1507 -2046 1507 -2046 0 1
rlabel polysilicon 1507 -2052 1507 -2052 0 3
rlabel polysilicon 1514 -2046 1514 -2046 0 1
rlabel polysilicon 1514 -2052 1514 -2052 0 3
rlabel polysilicon 1521 -2046 1521 -2046 0 1
rlabel polysilicon 1521 -2052 1521 -2052 0 3
rlabel polysilicon 1528 -2046 1528 -2046 0 1
rlabel polysilicon 1528 -2052 1528 -2052 0 3
rlabel polysilicon 1535 -2046 1535 -2046 0 1
rlabel polysilicon 1535 -2052 1535 -2052 0 3
rlabel polysilicon 1542 -2046 1542 -2046 0 1
rlabel polysilicon 1542 -2052 1542 -2052 0 3
rlabel polysilicon 1549 -2046 1549 -2046 0 1
rlabel polysilicon 1549 -2052 1549 -2052 0 3
rlabel polysilicon 1556 -2046 1556 -2046 0 1
rlabel polysilicon 1556 -2052 1556 -2052 0 3
rlabel polysilicon 1563 -2046 1563 -2046 0 1
rlabel polysilicon 1563 -2052 1563 -2052 0 3
rlabel polysilicon 1570 -2046 1570 -2046 0 1
rlabel polysilicon 1570 -2052 1570 -2052 0 3
rlabel polysilicon 1577 -2046 1577 -2046 0 1
rlabel polysilicon 1577 -2052 1577 -2052 0 3
rlabel polysilicon 1584 -2046 1584 -2046 0 1
rlabel polysilicon 1584 -2052 1584 -2052 0 3
rlabel polysilicon 1591 -2046 1591 -2046 0 1
rlabel polysilicon 1591 -2052 1591 -2052 0 3
rlabel polysilicon 1598 -2046 1598 -2046 0 1
rlabel polysilicon 1598 -2052 1598 -2052 0 3
rlabel polysilicon 1605 -2046 1605 -2046 0 1
rlabel polysilicon 1605 -2052 1605 -2052 0 3
rlabel polysilicon 1612 -2046 1612 -2046 0 1
rlabel polysilicon 1612 -2052 1612 -2052 0 3
rlabel polysilicon 1619 -2046 1619 -2046 0 1
rlabel polysilicon 1619 -2052 1619 -2052 0 3
rlabel polysilicon 1626 -2046 1626 -2046 0 1
rlabel polysilicon 1626 -2052 1626 -2052 0 3
rlabel polysilicon 1633 -2046 1633 -2046 0 1
rlabel polysilicon 1633 -2052 1633 -2052 0 3
rlabel polysilicon 1640 -2046 1640 -2046 0 1
rlabel polysilicon 1640 -2052 1640 -2052 0 3
rlabel polysilicon 1647 -2046 1647 -2046 0 1
rlabel polysilicon 1647 -2052 1647 -2052 0 3
rlabel polysilicon 1654 -2046 1654 -2046 0 1
rlabel polysilicon 1654 -2052 1654 -2052 0 3
rlabel polysilicon 1661 -2046 1661 -2046 0 1
rlabel polysilicon 1661 -2052 1661 -2052 0 3
rlabel polysilicon 1668 -2046 1668 -2046 0 1
rlabel polysilicon 1668 -2052 1668 -2052 0 3
rlabel polysilicon 1675 -2046 1675 -2046 0 1
rlabel polysilicon 1675 -2052 1675 -2052 0 3
rlabel polysilicon 1682 -2046 1682 -2046 0 1
rlabel polysilicon 1682 -2052 1682 -2052 0 3
rlabel polysilicon 1689 -2046 1689 -2046 0 1
rlabel polysilicon 1689 -2052 1689 -2052 0 3
rlabel polysilicon 1696 -2046 1696 -2046 0 1
rlabel polysilicon 1696 -2052 1696 -2052 0 3
rlabel polysilicon 1703 -2046 1703 -2046 0 1
rlabel polysilicon 1703 -2052 1703 -2052 0 3
rlabel polysilicon 1710 -2046 1710 -2046 0 1
rlabel polysilicon 1710 -2052 1710 -2052 0 3
rlabel polysilicon 1717 -2046 1717 -2046 0 1
rlabel polysilicon 1717 -2052 1717 -2052 0 3
rlabel polysilicon 1724 -2046 1724 -2046 0 1
rlabel polysilicon 1724 -2052 1724 -2052 0 3
rlabel polysilicon 1731 -2046 1731 -2046 0 1
rlabel polysilicon 1731 -2052 1731 -2052 0 3
rlabel polysilicon 1738 -2046 1738 -2046 0 1
rlabel polysilicon 1738 -2052 1738 -2052 0 3
rlabel polysilicon 1745 -2046 1745 -2046 0 1
rlabel polysilicon 1745 -2052 1745 -2052 0 3
rlabel polysilicon 1752 -2046 1752 -2046 0 1
rlabel polysilicon 1752 -2052 1752 -2052 0 3
rlabel polysilicon 1759 -2046 1759 -2046 0 1
rlabel polysilicon 1759 -2052 1759 -2052 0 3
rlabel polysilicon 1766 -2046 1766 -2046 0 1
rlabel polysilicon 1766 -2052 1766 -2052 0 3
rlabel polysilicon 1773 -2046 1773 -2046 0 1
rlabel polysilicon 1773 -2052 1773 -2052 0 3
rlabel polysilicon 1780 -2046 1780 -2046 0 1
rlabel polysilicon 1780 -2052 1780 -2052 0 3
rlabel polysilicon 1787 -2046 1787 -2046 0 1
rlabel polysilicon 1787 -2052 1787 -2052 0 3
rlabel polysilicon 1794 -2046 1794 -2046 0 1
rlabel polysilicon 1794 -2052 1794 -2052 0 3
rlabel polysilicon 1801 -2046 1801 -2046 0 1
rlabel polysilicon 1801 -2052 1801 -2052 0 3
rlabel polysilicon 1808 -2046 1808 -2046 0 1
rlabel polysilicon 1808 -2052 1808 -2052 0 3
rlabel polysilicon 1815 -2046 1815 -2046 0 1
rlabel polysilicon 1815 -2052 1815 -2052 0 3
rlabel polysilicon 1822 -2046 1822 -2046 0 1
rlabel polysilicon 1822 -2052 1822 -2052 0 3
rlabel polysilicon 1829 -2046 1829 -2046 0 1
rlabel polysilicon 1829 -2052 1829 -2052 0 3
rlabel polysilicon 1836 -2046 1836 -2046 0 1
rlabel polysilicon 1836 -2052 1836 -2052 0 3
rlabel polysilicon 1843 -2046 1843 -2046 0 1
rlabel polysilicon 1843 -2052 1843 -2052 0 3
rlabel polysilicon 1850 -2046 1850 -2046 0 1
rlabel polysilicon 1850 -2052 1850 -2052 0 3
rlabel polysilicon 1857 -2046 1857 -2046 0 1
rlabel polysilicon 1857 -2052 1857 -2052 0 3
rlabel polysilicon 1864 -2046 1864 -2046 0 1
rlabel polysilicon 1864 -2052 1864 -2052 0 3
rlabel polysilicon 1871 -2046 1871 -2046 0 1
rlabel polysilicon 1871 -2052 1871 -2052 0 3
rlabel polysilicon 1878 -2046 1878 -2046 0 1
rlabel polysilicon 1878 -2052 1878 -2052 0 3
rlabel polysilicon 1885 -2046 1885 -2046 0 1
rlabel polysilicon 1885 -2052 1885 -2052 0 3
rlabel polysilicon 1892 -2046 1892 -2046 0 1
rlabel polysilicon 1892 -2052 1892 -2052 0 3
rlabel polysilicon 1899 -2046 1899 -2046 0 1
rlabel polysilicon 1899 -2052 1899 -2052 0 3
rlabel polysilicon 1906 -2046 1906 -2046 0 1
rlabel polysilicon 1906 -2052 1906 -2052 0 3
rlabel polysilicon 1913 -2046 1913 -2046 0 1
rlabel polysilicon 1913 -2052 1913 -2052 0 3
rlabel polysilicon 1920 -2046 1920 -2046 0 1
rlabel polysilicon 1920 -2052 1920 -2052 0 3
rlabel polysilicon 1923 -2052 1923 -2052 0 4
rlabel polysilicon 1927 -2046 1927 -2046 0 1
rlabel polysilicon 1927 -2052 1927 -2052 0 3
rlabel polysilicon 1934 -2046 1934 -2046 0 1
rlabel polysilicon 1934 -2052 1934 -2052 0 3
rlabel polysilicon 1941 -2046 1941 -2046 0 1
rlabel polysilicon 1941 -2052 1941 -2052 0 3
rlabel polysilicon 1948 -2046 1948 -2046 0 1
rlabel polysilicon 1948 -2052 1948 -2052 0 3
rlabel polysilicon 1955 -2046 1955 -2046 0 1
rlabel polysilicon 1955 -2052 1955 -2052 0 3
rlabel polysilicon 1962 -2046 1962 -2046 0 1
rlabel polysilicon 1962 -2052 1962 -2052 0 3
rlabel polysilicon 1969 -2046 1969 -2046 0 1
rlabel polysilicon 1969 -2052 1969 -2052 0 3
rlabel polysilicon 1976 -2046 1976 -2046 0 1
rlabel polysilicon 1976 -2052 1976 -2052 0 3
rlabel polysilicon 1983 -2046 1983 -2046 0 1
rlabel polysilicon 1983 -2052 1983 -2052 0 3
rlabel polysilicon 1990 -2046 1990 -2046 0 1
rlabel polysilicon 1990 -2052 1990 -2052 0 3
rlabel polysilicon 2 -2187 2 -2187 0 1
rlabel polysilicon 2 -2193 2 -2193 0 3
rlabel polysilicon 12 -2193 12 -2193 0 4
rlabel polysilicon 16 -2187 16 -2187 0 1
rlabel polysilicon 16 -2193 16 -2193 0 3
rlabel polysilicon 23 -2187 23 -2187 0 1
rlabel polysilicon 23 -2193 23 -2193 0 3
rlabel polysilicon 30 -2187 30 -2187 0 1
rlabel polysilicon 33 -2187 33 -2187 0 2
rlabel polysilicon 30 -2193 30 -2193 0 3
rlabel polysilicon 33 -2193 33 -2193 0 4
rlabel polysilicon 40 -2187 40 -2187 0 2
rlabel polysilicon 37 -2193 37 -2193 0 3
rlabel polysilicon 40 -2193 40 -2193 0 4
rlabel polysilicon 44 -2187 44 -2187 0 1
rlabel polysilicon 44 -2193 44 -2193 0 3
rlabel polysilicon 51 -2187 51 -2187 0 1
rlabel polysilicon 51 -2193 51 -2193 0 3
rlabel polysilicon 58 -2187 58 -2187 0 1
rlabel polysilicon 58 -2193 58 -2193 0 3
rlabel polysilicon 65 -2187 65 -2187 0 1
rlabel polysilicon 65 -2193 65 -2193 0 3
rlabel polysilicon 72 -2187 72 -2187 0 1
rlabel polysilicon 72 -2193 72 -2193 0 3
rlabel polysilicon 79 -2187 79 -2187 0 1
rlabel polysilicon 79 -2193 79 -2193 0 3
rlabel polysilicon 86 -2187 86 -2187 0 1
rlabel polysilicon 89 -2187 89 -2187 0 2
rlabel polysilicon 86 -2193 86 -2193 0 3
rlabel polysilicon 89 -2193 89 -2193 0 4
rlabel polysilicon 93 -2187 93 -2187 0 1
rlabel polysilicon 96 -2187 96 -2187 0 2
rlabel polysilicon 93 -2193 93 -2193 0 3
rlabel polysilicon 100 -2187 100 -2187 0 1
rlabel polysilicon 100 -2193 100 -2193 0 3
rlabel polysilicon 110 -2187 110 -2187 0 2
rlabel polysilicon 107 -2193 107 -2193 0 3
rlabel polysilicon 110 -2193 110 -2193 0 4
rlabel polysilicon 121 -2187 121 -2187 0 1
rlabel polysilicon 121 -2193 121 -2193 0 3
rlabel polysilicon 128 -2187 128 -2187 0 1
rlabel polysilicon 128 -2193 128 -2193 0 3
rlabel polysilicon 135 -2187 135 -2187 0 1
rlabel polysilicon 135 -2193 135 -2193 0 3
rlabel polysilicon 142 -2187 142 -2187 0 1
rlabel polysilicon 142 -2193 142 -2193 0 3
rlabel polysilicon 149 -2187 149 -2187 0 1
rlabel polysilicon 149 -2193 149 -2193 0 3
rlabel polysilicon 156 -2187 156 -2187 0 1
rlabel polysilicon 156 -2193 156 -2193 0 3
rlabel polysilicon 163 -2187 163 -2187 0 1
rlabel polysilicon 163 -2193 163 -2193 0 3
rlabel polysilicon 170 -2187 170 -2187 0 1
rlabel polysilicon 170 -2193 170 -2193 0 3
rlabel polysilicon 177 -2187 177 -2187 0 1
rlabel polysilicon 177 -2193 177 -2193 0 3
rlabel polysilicon 184 -2187 184 -2187 0 1
rlabel polysilicon 184 -2193 184 -2193 0 3
rlabel polysilicon 191 -2187 191 -2187 0 1
rlabel polysilicon 191 -2193 191 -2193 0 3
rlabel polysilicon 198 -2187 198 -2187 0 1
rlabel polysilicon 198 -2193 198 -2193 0 3
rlabel polysilicon 205 -2187 205 -2187 0 1
rlabel polysilicon 205 -2193 205 -2193 0 3
rlabel polysilicon 212 -2187 212 -2187 0 1
rlabel polysilicon 212 -2193 212 -2193 0 3
rlabel polysilicon 219 -2187 219 -2187 0 1
rlabel polysilicon 219 -2193 219 -2193 0 3
rlabel polysilicon 226 -2187 226 -2187 0 1
rlabel polysilicon 226 -2193 226 -2193 0 3
rlabel polysilicon 233 -2187 233 -2187 0 1
rlabel polysilicon 236 -2187 236 -2187 0 2
rlabel polysilicon 240 -2187 240 -2187 0 1
rlabel polysilicon 240 -2193 240 -2193 0 3
rlabel polysilicon 247 -2187 247 -2187 0 1
rlabel polysilicon 247 -2193 247 -2193 0 3
rlabel polysilicon 254 -2187 254 -2187 0 1
rlabel polysilicon 254 -2193 254 -2193 0 3
rlabel polysilicon 261 -2187 261 -2187 0 1
rlabel polysilicon 261 -2193 261 -2193 0 3
rlabel polysilicon 268 -2187 268 -2187 0 1
rlabel polysilicon 268 -2193 268 -2193 0 3
rlabel polysilicon 275 -2187 275 -2187 0 1
rlabel polysilicon 275 -2193 275 -2193 0 3
rlabel polysilicon 282 -2187 282 -2187 0 1
rlabel polysilicon 282 -2193 282 -2193 0 3
rlabel polysilicon 289 -2187 289 -2187 0 1
rlabel polysilicon 289 -2193 289 -2193 0 3
rlabel polysilicon 296 -2187 296 -2187 0 1
rlabel polysilicon 296 -2193 296 -2193 0 3
rlabel polysilicon 303 -2187 303 -2187 0 1
rlabel polysilicon 303 -2193 303 -2193 0 3
rlabel polysilicon 310 -2187 310 -2187 0 1
rlabel polysilicon 310 -2193 310 -2193 0 3
rlabel polysilicon 317 -2187 317 -2187 0 1
rlabel polysilicon 317 -2193 317 -2193 0 3
rlabel polysilicon 324 -2187 324 -2187 0 1
rlabel polysilicon 324 -2193 324 -2193 0 3
rlabel polysilicon 331 -2187 331 -2187 0 1
rlabel polysilicon 331 -2193 331 -2193 0 3
rlabel polysilicon 341 -2187 341 -2187 0 2
rlabel polysilicon 341 -2193 341 -2193 0 4
rlabel polysilicon 345 -2187 345 -2187 0 1
rlabel polysilicon 345 -2193 345 -2193 0 3
rlabel polysilicon 352 -2187 352 -2187 0 1
rlabel polysilicon 352 -2193 352 -2193 0 3
rlabel polysilicon 359 -2187 359 -2187 0 1
rlabel polysilicon 359 -2193 359 -2193 0 3
rlabel polysilicon 366 -2187 366 -2187 0 1
rlabel polysilicon 366 -2193 366 -2193 0 3
rlabel polysilicon 373 -2187 373 -2187 0 1
rlabel polysilicon 373 -2193 373 -2193 0 3
rlabel polysilicon 380 -2187 380 -2187 0 1
rlabel polysilicon 380 -2193 380 -2193 0 3
rlabel polysilicon 387 -2187 387 -2187 0 1
rlabel polysilicon 390 -2187 390 -2187 0 2
rlabel polysilicon 387 -2193 387 -2193 0 3
rlabel polysilicon 390 -2193 390 -2193 0 4
rlabel polysilicon 394 -2187 394 -2187 0 1
rlabel polysilicon 394 -2193 394 -2193 0 3
rlabel polysilicon 401 -2187 401 -2187 0 1
rlabel polysilicon 404 -2187 404 -2187 0 2
rlabel polysilicon 401 -2193 401 -2193 0 3
rlabel polysilicon 408 -2187 408 -2187 0 1
rlabel polysilicon 408 -2193 408 -2193 0 3
rlabel polysilicon 415 -2187 415 -2187 0 1
rlabel polysilicon 415 -2193 415 -2193 0 3
rlabel polysilicon 422 -2187 422 -2187 0 1
rlabel polysilicon 422 -2193 422 -2193 0 3
rlabel polysilicon 429 -2187 429 -2187 0 1
rlabel polysilicon 429 -2193 429 -2193 0 3
rlabel polysilicon 436 -2187 436 -2187 0 1
rlabel polysilicon 439 -2187 439 -2187 0 2
rlabel polysilicon 436 -2193 436 -2193 0 3
rlabel polysilicon 443 -2187 443 -2187 0 1
rlabel polysilicon 443 -2193 443 -2193 0 3
rlabel polysilicon 450 -2187 450 -2187 0 1
rlabel polysilicon 450 -2193 450 -2193 0 3
rlabel polysilicon 457 -2187 457 -2187 0 1
rlabel polysilicon 457 -2193 457 -2193 0 3
rlabel polysilicon 464 -2187 464 -2187 0 1
rlabel polysilicon 467 -2187 467 -2187 0 2
rlabel polysilicon 464 -2193 464 -2193 0 3
rlabel polysilicon 471 -2187 471 -2187 0 1
rlabel polysilicon 471 -2193 471 -2193 0 3
rlabel polysilicon 478 -2187 478 -2187 0 1
rlabel polysilicon 478 -2193 478 -2193 0 3
rlabel polysilicon 485 -2187 485 -2187 0 1
rlabel polysilicon 485 -2193 485 -2193 0 3
rlabel polysilicon 492 -2187 492 -2187 0 1
rlabel polysilicon 492 -2193 492 -2193 0 3
rlabel polysilicon 499 -2187 499 -2187 0 1
rlabel polysilicon 499 -2193 499 -2193 0 3
rlabel polysilicon 506 -2187 506 -2187 0 1
rlabel polysilicon 509 -2187 509 -2187 0 2
rlabel polysilicon 506 -2193 506 -2193 0 3
rlabel polysilicon 509 -2193 509 -2193 0 4
rlabel polysilicon 513 -2187 513 -2187 0 1
rlabel polysilicon 513 -2193 513 -2193 0 3
rlabel polysilicon 520 -2187 520 -2187 0 1
rlabel polysilicon 520 -2193 520 -2193 0 3
rlabel polysilicon 527 -2187 527 -2187 0 1
rlabel polysilicon 527 -2193 527 -2193 0 3
rlabel polysilicon 534 -2187 534 -2187 0 1
rlabel polysilicon 534 -2193 534 -2193 0 3
rlabel polysilicon 541 -2193 541 -2193 0 3
rlabel polysilicon 544 -2193 544 -2193 0 4
rlabel polysilicon 548 -2187 548 -2187 0 1
rlabel polysilicon 548 -2193 548 -2193 0 3
rlabel polysilicon 555 -2187 555 -2187 0 1
rlabel polysilicon 555 -2193 555 -2193 0 3
rlabel polysilicon 562 -2187 562 -2187 0 1
rlabel polysilicon 562 -2193 562 -2193 0 3
rlabel polysilicon 569 -2187 569 -2187 0 1
rlabel polysilicon 569 -2193 569 -2193 0 3
rlabel polysilicon 576 -2187 576 -2187 0 1
rlabel polysilicon 576 -2193 576 -2193 0 3
rlabel polysilicon 583 -2187 583 -2187 0 1
rlabel polysilicon 583 -2193 583 -2193 0 3
rlabel polysilicon 590 -2187 590 -2187 0 1
rlabel polysilicon 593 -2187 593 -2187 0 2
rlabel polysilicon 590 -2193 590 -2193 0 3
rlabel polysilicon 597 -2187 597 -2187 0 1
rlabel polysilicon 597 -2193 597 -2193 0 3
rlabel polysilicon 604 -2187 604 -2187 0 1
rlabel polysilicon 604 -2193 604 -2193 0 3
rlabel polysilicon 611 -2187 611 -2187 0 1
rlabel polysilicon 611 -2193 611 -2193 0 3
rlabel polysilicon 618 -2187 618 -2187 0 1
rlabel polysilicon 618 -2193 618 -2193 0 3
rlabel polysilicon 625 -2187 625 -2187 0 1
rlabel polysilicon 628 -2187 628 -2187 0 2
rlabel polysilicon 632 -2187 632 -2187 0 1
rlabel polysilicon 632 -2193 632 -2193 0 3
rlabel polysilicon 639 -2187 639 -2187 0 1
rlabel polysilicon 639 -2193 639 -2193 0 3
rlabel polysilicon 646 -2187 646 -2187 0 1
rlabel polysilicon 649 -2187 649 -2187 0 2
rlabel polysilicon 649 -2193 649 -2193 0 4
rlabel polysilicon 653 -2187 653 -2187 0 1
rlabel polysilicon 653 -2193 653 -2193 0 3
rlabel polysilicon 660 -2187 660 -2187 0 1
rlabel polysilicon 660 -2193 660 -2193 0 3
rlabel polysilicon 667 -2187 667 -2187 0 1
rlabel polysilicon 667 -2193 667 -2193 0 3
rlabel polysilicon 674 -2187 674 -2187 0 1
rlabel polysilicon 674 -2193 674 -2193 0 3
rlabel polysilicon 681 -2187 681 -2187 0 1
rlabel polysilicon 681 -2193 681 -2193 0 3
rlabel polysilicon 688 -2187 688 -2187 0 1
rlabel polysilicon 688 -2193 688 -2193 0 3
rlabel polysilicon 695 -2187 695 -2187 0 1
rlabel polysilicon 695 -2193 695 -2193 0 3
rlabel polysilicon 702 -2187 702 -2187 0 1
rlabel polysilicon 702 -2193 702 -2193 0 3
rlabel polysilicon 709 -2187 709 -2187 0 1
rlabel polysilicon 709 -2193 709 -2193 0 3
rlabel polysilicon 716 -2187 716 -2187 0 1
rlabel polysilicon 716 -2193 716 -2193 0 3
rlabel polysilicon 723 -2187 723 -2187 0 1
rlabel polysilicon 723 -2193 723 -2193 0 3
rlabel polysilicon 730 -2187 730 -2187 0 1
rlabel polysilicon 730 -2193 730 -2193 0 3
rlabel polysilicon 737 -2187 737 -2187 0 1
rlabel polysilicon 737 -2193 737 -2193 0 3
rlabel polysilicon 744 -2187 744 -2187 0 1
rlabel polysilicon 744 -2193 744 -2193 0 3
rlabel polysilicon 751 -2187 751 -2187 0 1
rlabel polysilicon 751 -2193 751 -2193 0 3
rlabel polysilicon 758 -2187 758 -2187 0 1
rlabel polysilicon 758 -2193 758 -2193 0 3
rlabel polysilicon 765 -2187 765 -2187 0 1
rlabel polysilicon 765 -2193 765 -2193 0 3
rlabel polysilicon 772 -2187 772 -2187 0 1
rlabel polysilicon 772 -2193 772 -2193 0 3
rlabel polysilicon 779 -2187 779 -2187 0 1
rlabel polysilicon 779 -2193 779 -2193 0 3
rlabel polysilicon 786 -2187 786 -2187 0 1
rlabel polysilicon 786 -2193 786 -2193 0 3
rlabel polysilicon 793 -2187 793 -2187 0 1
rlabel polysilicon 793 -2193 793 -2193 0 3
rlabel polysilicon 800 -2187 800 -2187 0 1
rlabel polysilicon 800 -2193 800 -2193 0 3
rlabel polysilicon 807 -2187 807 -2187 0 1
rlabel polysilicon 807 -2193 807 -2193 0 3
rlabel polysilicon 814 -2187 814 -2187 0 1
rlabel polysilicon 814 -2193 814 -2193 0 3
rlabel polysilicon 821 -2187 821 -2187 0 1
rlabel polysilicon 821 -2193 821 -2193 0 3
rlabel polysilicon 828 -2187 828 -2187 0 1
rlabel polysilicon 828 -2193 828 -2193 0 3
rlabel polysilicon 835 -2187 835 -2187 0 1
rlabel polysilicon 838 -2187 838 -2187 0 2
rlabel polysilicon 835 -2193 835 -2193 0 3
rlabel polysilicon 842 -2187 842 -2187 0 1
rlabel polysilicon 842 -2193 842 -2193 0 3
rlabel polysilicon 849 -2187 849 -2187 0 1
rlabel polysilicon 849 -2193 849 -2193 0 3
rlabel polysilicon 856 -2187 856 -2187 0 1
rlabel polysilicon 856 -2193 856 -2193 0 3
rlabel polysilicon 863 -2187 863 -2187 0 1
rlabel polysilicon 863 -2193 863 -2193 0 3
rlabel polysilicon 870 -2187 870 -2187 0 1
rlabel polysilicon 870 -2193 870 -2193 0 3
rlabel polysilicon 877 -2187 877 -2187 0 1
rlabel polysilicon 880 -2187 880 -2187 0 2
rlabel polysilicon 877 -2193 877 -2193 0 3
rlabel polysilicon 880 -2193 880 -2193 0 4
rlabel polysilicon 884 -2187 884 -2187 0 1
rlabel polysilicon 884 -2193 884 -2193 0 3
rlabel polysilicon 891 -2187 891 -2187 0 1
rlabel polysilicon 891 -2193 891 -2193 0 3
rlabel polysilicon 898 -2187 898 -2187 0 1
rlabel polysilicon 898 -2193 898 -2193 0 3
rlabel polysilicon 905 -2187 905 -2187 0 1
rlabel polysilicon 905 -2193 905 -2193 0 3
rlabel polysilicon 912 -2187 912 -2187 0 1
rlabel polysilicon 912 -2193 912 -2193 0 3
rlabel polysilicon 919 -2187 919 -2187 0 1
rlabel polysilicon 919 -2193 919 -2193 0 3
rlabel polysilicon 926 -2187 926 -2187 0 1
rlabel polysilicon 926 -2193 926 -2193 0 3
rlabel polysilicon 933 -2187 933 -2187 0 1
rlabel polysilicon 933 -2193 933 -2193 0 3
rlabel polysilicon 940 -2187 940 -2187 0 1
rlabel polysilicon 940 -2193 940 -2193 0 3
rlabel polysilicon 947 -2187 947 -2187 0 1
rlabel polysilicon 947 -2193 947 -2193 0 3
rlabel polysilicon 954 -2187 954 -2187 0 1
rlabel polysilicon 954 -2193 954 -2193 0 3
rlabel polysilicon 961 -2187 961 -2187 0 1
rlabel polysilicon 961 -2193 961 -2193 0 3
rlabel polysilicon 968 -2187 968 -2187 0 1
rlabel polysilicon 971 -2187 971 -2187 0 2
rlabel polysilicon 968 -2193 968 -2193 0 3
rlabel polysilicon 971 -2193 971 -2193 0 4
rlabel polysilicon 975 -2187 975 -2187 0 1
rlabel polysilicon 978 -2187 978 -2187 0 2
rlabel polysilicon 975 -2193 975 -2193 0 3
rlabel polysilicon 978 -2193 978 -2193 0 4
rlabel polysilicon 982 -2187 982 -2187 0 1
rlabel polysilicon 982 -2193 982 -2193 0 3
rlabel polysilicon 989 -2187 989 -2187 0 1
rlabel polysilicon 989 -2193 989 -2193 0 3
rlabel polysilicon 996 -2187 996 -2187 0 1
rlabel polysilicon 996 -2193 996 -2193 0 3
rlabel polysilicon 1003 -2187 1003 -2187 0 1
rlabel polysilicon 1003 -2193 1003 -2193 0 3
rlabel polysilicon 1010 -2187 1010 -2187 0 1
rlabel polysilicon 1010 -2193 1010 -2193 0 3
rlabel polysilicon 1017 -2187 1017 -2187 0 1
rlabel polysilicon 1017 -2193 1017 -2193 0 3
rlabel polysilicon 1024 -2187 1024 -2187 0 1
rlabel polysilicon 1024 -2193 1024 -2193 0 3
rlabel polysilicon 1031 -2187 1031 -2187 0 1
rlabel polysilicon 1031 -2193 1031 -2193 0 3
rlabel polysilicon 1038 -2187 1038 -2187 0 1
rlabel polysilicon 1038 -2193 1038 -2193 0 3
rlabel polysilicon 1045 -2187 1045 -2187 0 1
rlabel polysilicon 1045 -2193 1045 -2193 0 3
rlabel polysilicon 1052 -2187 1052 -2187 0 1
rlabel polysilicon 1052 -2193 1052 -2193 0 3
rlabel polysilicon 1055 -2193 1055 -2193 0 4
rlabel polysilicon 1059 -2187 1059 -2187 0 1
rlabel polysilicon 1059 -2193 1059 -2193 0 3
rlabel polysilicon 1066 -2187 1066 -2187 0 1
rlabel polysilicon 1069 -2187 1069 -2187 0 2
rlabel polysilicon 1066 -2193 1066 -2193 0 3
rlabel polysilicon 1069 -2193 1069 -2193 0 4
rlabel polysilicon 1073 -2187 1073 -2187 0 1
rlabel polysilicon 1073 -2193 1073 -2193 0 3
rlabel polysilicon 1080 -2187 1080 -2187 0 1
rlabel polysilicon 1083 -2187 1083 -2187 0 2
rlabel polysilicon 1083 -2193 1083 -2193 0 4
rlabel polysilicon 1087 -2187 1087 -2187 0 1
rlabel polysilicon 1087 -2193 1087 -2193 0 3
rlabel polysilicon 1094 -2187 1094 -2187 0 1
rlabel polysilicon 1094 -2193 1094 -2193 0 3
rlabel polysilicon 1101 -2187 1101 -2187 0 1
rlabel polysilicon 1101 -2193 1101 -2193 0 3
rlabel polysilicon 1108 -2187 1108 -2187 0 1
rlabel polysilicon 1111 -2187 1111 -2187 0 2
rlabel polysilicon 1108 -2193 1108 -2193 0 3
rlabel polysilicon 1111 -2193 1111 -2193 0 4
rlabel polysilicon 1115 -2187 1115 -2187 0 1
rlabel polysilicon 1115 -2193 1115 -2193 0 3
rlabel polysilicon 1122 -2187 1122 -2187 0 1
rlabel polysilicon 1122 -2193 1122 -2193 0 3
rlabel polysilicon 1129 -2187 1129 -2187 0 1
rlabel polysilicon 1129 -2193 1129 -2193 0 3
rlabel polysilicon 1139 -2187 1139 -2187 0 2
rlabel polysilicon 1139 -2193 1139 -2193 0 4
rlabel polysilicon 1143 -2187 1143 -2187 0 1
rlabel polysilicon 1143 -2193 1143 -2193 0 3
rlabel polysilicon 1150 -2187 1150 -2187 0 1
rlabel polysilicon 1150 -2193 1150 -2193 0 3
rlabel polysilicon 1157 -2187 1157 -2187 0 1
rlabel polysilicon 1160 -2187 1160 -2187 0 2
rlabel polysilicon 1157 -2193 1157 -2193 0 3
rlabel polysilicon 1160 -2193 1160 -2193 0 4
rlabel polysilicon 1164 -2187 1164 -2187 0 1
rlabel polysilicon 1164 -2193 1164 -2193 0 3
rlabel polysilicon 1171 -2187 1171 -2187 0 1
rlabel polysilicon 1171 -2193 1171 -2193 0 3
rlabel polysilicon 1178 -2187 1178 -2187 0 1
rlabel polysilicon 1178 -2193 1178 -2193 0 3
rlabel polysilicon 1185 -2187 1185 -2187 0 1
rlabel polysilicon 1185 -2193 1185 -2193 0 3
rlabel polysilicon 1192 -2187 1192 -2187 0 1
rlabel polysilicon 1192 -2193 1192 -2193 0 3
rlabel polysilicon 1199 -2187 1199 -2187 0 1
rlabel polysilicon 1199 -2193 1199 -2193 0 3
rlabel polysilicon 1206 -2187 1206 -2187 0 1
rlabel polysilicon 1206 -2193 1206 -2193 0 3
rlabel polysilicon 1213 -2187 1213 -2187 0 1
rlabel polysilicon 1213 -2193 1213 -2193 0 3
rlabel polysilicon 1220 -2187 1220 -2187 0 1
rlabel polysilicon 1220 -2193 1220 -2193 0 3
rlabel polysilicon 1227 -2187 1227 -2187 0 1
rlabel polysilicon 1227 -2193 1227 -2193 0 3
rlabel polysilicon 1234 -2187 1234 -2187 0 1
rlabel polysilicon 1234 -2193 1234 -2193 0 3
rlabel polysilicon 1241 -2187 1241 -2187 0 1
rlabel polysilicon 1241 -2193 1241 -2193 0 3
rlabel polysilicon 1248 -2187 1248 -2187 0 1
rlabel polysilicon 1248 -2193 1248 -2193 0 3
rlabel polysilicon 1255 -2187 1255 -2187 0 1
rlabel polysilicon 1255 -2193 1255 -2193 0 3
rlabel polysilicon 1262 -2187 1262 -2187 0 1
rlabel polysilicon 1262 -2193 1262 -2193 0 3
rlabel polysilicon 1269 -2187 1269 -2187 0 1
rlabel polysilicon 1269 -2193 1269 -2193 0 3
rlabel polysilicon 1276 -2187 1276 -2187 0 1
rlabel polysilicon 1276 -2193 1276 -2193 0 3
rlabel polysilicon 1279 -2193 1279 -2193 0 4
rlabel polysilicon 1283 -2187 1283 -2187 0 1
rlabel polysilicon 1283 -2193 1283 -2193 0 3
rlabel polysilicon 1290 -2187 1290 -2187 0 1
rlabel polysilicon 1290 -2193 1290 -2193 0 3
rlabel polysilicon 1297 -2187 1297 -2187 0 1
rlabel polysilicon 1297 -2193 1297 -2193 0 3
rlabel polysilicon 1304 -2187 1304 -2187 0 1
rlabel polysilicon 1304 -2193 1304 -2193 0 3
rlabel polysilicon 1311 -2187 1311 -2187 0 1
rlabel polysilicon 1311 -2193 1311 -2193 0 3
rlabel polysilicon 1318 -2187 1318 -2187 0 1
rlabel polysilicon 1318 -2193 1318 -2193 0 3
rlabel polysilicon 1325 -2187 1325 -2187 0 1
rlabel polysilicon 1325 -2193 1325 -2193 0 3
rlabel polysilicon 1332 -2187 1332 -2187 0 1
rlabel polysilicon 1332 -2193 1332 -2193 0 3
rlabel polysilicon 1339 -2187 1339 -2187 0 1
rlabel polysilicon 1339 -2193 1339 -2193 0 3
rlabel polysilicon 1346 -2187 1346 -2187 0 1
rlabel polysilicon 1346 -2193 1346 -2193 0 3
rlabel polysilicon 1353 -2187 1353 -2187 0 1
rlabel polysilicon 1353 -2193 1353 -2193 0 3
rlabel polysilicon 1360 -2187 1360 -2187 0 1
rlabel polysilicon 1363 -2187 1363 -2187 0 2
rlabel polysilicon 1360 -2193 1360 -2193 0 3
rlabel polysilicon 1367 -2187 1367 -2187 0 1
rlabel polysilicon 1367 -2193 1367 -2193 0 3
rlabel polysilicon 1374 -2187 1374 -2187 0 1
rlabel polysilicon 1377 -2187 1377 -2187 0 2
rlabel polysilicon 1374 -2193 1374 -2193 0 3
rlabel polysilicon 1381 -2187 1381 -2187 0 1
rlabel polysilicon 1381 -2193 1381 -2193 0 3
rlabel polysilicon 1388 -2187 1388 -2187 0 1
rlabel polysilicon 1388 -2193 1388 -2193 0 3
rlabel polysilicon 1395 -2187 1395 -2187 0 1
rlabel polysilicon 1398 -2187 1398 -2187 0 2
rlabel polysilicon 1395 -2193 1395 -2193 0 3
rlabel polysilicon 1398 -2193 1398 -2193 0 4
rlabel polysilicon 1402 -2187 1402 -2187 0 1
rlabel polysilicon 1402 -2193 1402 -2193 0 3
rlabel polysilicon 1409 -2187 1409 -2187 0 1
rlabel polysilicon 1409 -2193 1409 -2193 0 3
rlabel polysilicon 1416 -2187 1416 -2187 0 1
rlabel polysilicon 1416 -2193 1416 -2193 0 3
rlabel polysilicon 1423 -2187 1423 -2187 0 1
rlabel polysilicon 1423 -2193 1423 -2193 0 3
rlabel polysilicon 1430 -2187 1430 -2187 0 1
rlabel polysilicon 1430 -2193 1430 -2193 0 3
rlabel polysilicon 1437 -2187 1437 -2187 0 1
rlabel polysilicon 1437 -2193 1437 -2193 0 3
rlabel polysilicon 1444 -2187 1444 -2187 0 1
rlabel polysilicon 1444 -2193 1444 -2193 0 3
rlabel polysilicon 1451 -2187 1451 -2187 0 1
rlabel polysilicon 1454 -2187 1454 -2187 0 2
rlabel polysilicon 1454 -2193 1454 -2193 0 4
rlabel polysilicon 1458 -2187 1458 -2187 0 1
rlabel polysilicon 1458 -2193 1458 -2193 0 3
rlabel polysilicon 1465 -2187 1465 -2187 0 1
rlabel polysilicon 1465 -2193 1465 -2193 0 3
rlabel polysilicon 1475 -2187 1475 -2187 0 2
rlabel polysilicon 1472 -2193 1472 -2193 0 3
rlabel polysilicon 1475 -2193 1475 -2193 0 4
rlabel polysilicon 1479 -2187 1479 -2187 0 1
rlabel polysilicon 1479 -2193 1479 -2193 0 3
rlabel polysilicon 1486 -2187 1486 -2187 0 1
rlabel polysilicon 1486 -2193 1486 -2193 0 3
rlabel polysilicon 1493 -2187 1493 -2187 0 1
rlabel polysilicon 1493 -2193 1493 -2193 0 3
rlabel polysilicon 1500 -2187 1500 -2187 0 1
rlabel polysilicon 1500 -2193 1500 -2193 0 3
rlabel polysilicon 1507 -2187 1507 -2187 0 1
rlabel polysilicon 1507 -2193 1507 -2193 0 3
rlabel polysilicon 1514 -2187 1514 -2187 0 1
rlabel polysilicon 1514 -2193 1514 -2193 0 3
rlabel polysilicon 1521 -2187 1521 -2187 0 1
rlabel polysilicon 1521 -2193 1521 -2193 0 3
rlabel polysilicon 1528 -2187 1528 -2187 0 1
rlabel polysilicon 1528 -2193 1528 -2193 0 3
rlabel polysilicon 1535 -2187 1535 -2187 0 1
rlabel polysilicon 1535 -2193 1535 -2193 0 3
rlabel polysilicon 1542 -2187 1542 -2187 0 1
rlabel polysilicon 1542 -2193 1542 -2193 0 3
rlabel polysilicon 1549 -2187 1549 -2187 0 1
rlabel polysilicon 1549 -2193 1549 -2193 0 3
rlabel polysilicon 1556 -2187 1556 -2187 0 1
rlabel polysilicon 1556 -2193 1556 -2193 0 3
rlabel polysilicon 1563 -2187 1563 -2187 0 1
rlabel polysilicon 1563 -2193 1563 -2193 0 3
rlabel polysilicon 1570 -2187 1570 -2187 0 1
rlabel polysilicon 1570 -2193 1570 -2193 0 3
rlabel polysilicon 1577 -2187 1577 -2187 0 1
rlabel polysilicon 1577 -2193 1577 -2193 0 3
rlabel polysilicon 1584 -2187 1584 -2187 0 1
rlabel polysilicon 1584 -2193 1584 -2193 0 3
rlabel polysilicon 1591 -2187 1591 -2187 0 1
rlabel polysilicon 1591 -2193 1591 -2193 0 3
rlabel polysilicon 1598 -2187 1598 -2187 0 1
rlabel polysilicon 1598 -2193 1598 -2193 0 3
rlabel polysilicon 1605 -2187 1605 -2187 0 1
rlabel polysilicon 1605 -2193 1605 -2193 0 3
rlabel polysilicon 1612 -2187 1612 -2187 0 1
rlabel polysilicon 1612 -2193 1612 -2193 0 3
rlabel polysilicon 1619 -2187 1619 -2187 0 1
rlabel polysilicon 1619 -2193 1619 -2193 0 3
rlabel polysilicon 1626 -2187 1626 -2187 0 1
rlabel polysilicon 1626 -2193 1626 -2193 0 3
rlabel polysilicon 1633 -2187 1633 -2187 0 1
rlabel polysilicon 1633 -2193 1633 -2193 0 3
rlabel polysilicon 1640 -2187 1640 -2187 0 1
rlabel polysilicon 1640 -2193 1640 -2193 0 3
rlabel polysilicon 1647 -2187 1647 -2187 0 1
rlabel polysilicon 1647 -2193 1647 -2193 0 3
rlabel polysilicon 1654 -2187 1654 -2187 0 1
rlabel polysilicon 1654 -2193 1654 -2193 0 3
rlabel polysilicon 1661 -2187 1661 -2187 0 1
rlabel polysilicon 1661 -2193 1661 -2193 0 3
rlabel polysilicon 1668 -2187 1668 -2187 0 1
rlabel polysilicon 1668 -2193 1668 -2193 0 3
rlabel polysilicon 1675 -2187 1675 -2187 0 1
rlabel polysilicon 1675 -2193 1675 -2193 0 3
rlabel polysilicon 1682 -2187 1682 -2187 0 1
rlabel polysilicon 1682 -2193 1682 -2193 0 3
rlabel polysilicon 1689 -2187 1689 -2187 0 1
rlabel polysilicon 1689 -2193 1689 -2193 0 3
rlabel polysilicon 1696 -2187 1696 -2187 0 1
rlabel polysilicon 1696 -2193 1696 -2193 0 3
rlabel polysilicon 1703 -2187 1703 -2187 0 1
rlabel polysilicon 1703 -2193 1703 -2193 0 3
rlabel polysilicon 1710 -2187 1710 -2187 0 1
rlabel polysilicon 1710 -2193 1710 -2193 0 3
rlabel polysilicon 1717 -2187 1717 -2187 0 1
rlabel polysilicon 1717 -2193 1717 -2193 0 3
rlabel polysilicon 1724 -2187 1724 -2187 0 1
rlabel polysilicon 1724 -2193 1724 -2193 0 3
rlabel polysilicon 1731 -2187 1731 -2187 0 1
rlabel polysilicon 1731 -2193 1731 -2193 0 3
rlabel polysilicon 1738 -2187 1738 -2187 0 1
rlabel polysilicon 1738 -2193 1738 -2193 0 3
rlabel polysilicon 1745 -2187 1745 -2187 0 1
rlabel polysilicon 1745 -2193 1745 -2193 0 3
rlabel polysilicon 1752 -2187 1752 -2187 0 1
rlabel polysilicon 1752 -2193 1752 -2193 0 3
rlabel polysilicon 1759 -2187 1759 -2187 0 1
rlabel polysilicon 1759 -2193 1759 -2193 0 3
rlabel polysilicon 1766 -2187 1766 -2187 0 1
rlabel polysilicon 1766 -2193 1766 -2193 0 3
rlabel polysilicon 1773 -2187 1773 -2187 0 1
rlabel polysilicon 1773 -2193 1773 -2193 0 3
rlabel polysilicon 1780 -2187 1780 -2187 0 1
rlabel polysilicon 1780 -2193 1780 -2193 0 3
rlabel polysilicon 1787 -2187 1787 -2187 0 1
rlabel polysilicon 1787 -2193 1787 -2193 0 3
rlabel polysilicon 1794 -2187 1794 -2187 0 1
rlabel polysilicon 1794 -2193 1794 -2193 0 3
rlabel polysilicon 1801 -2187 1801 -2187 0 1
rlabel polysilicon 1801 -2193 1801 -2193 0 3
rlabel polysilicon 1808 -2187 1808 -2187 0 1
rlabel polysilicon 1808 -2193 1808 -2193 0 3
rlabel polysilicon 1815 -2187 1815 -2187 0 1
rlabel polysilicon 1815 -2193 1815 -2193 0 3
rlabel polysilicon 1822 -2187 1822 -2187 0 1
rlabel polysilicon 1822 -2193 1822 -2193 0 3
rlabel polysilicon 1829 -2187 1829 -2187 0 1
rlabel polysilicon 1829 -2193 1829 -2193 0 3
rlabel polysilicon 1836 -2187 1836 -2187 0 1
rlabel polysilicon 1836 -2193 1836 -2193 0 3
rlabel polysilicon 1843 -2187 1843 -2187 0 1
rlabel polysilicon 1843 -2193 1843 -2193 0 3
rlabel polysilicon 1850 -2187 1850 -2187 0 1
rlabel polysilicon 1850 -2193 1850 -2193 0 3
rlabel polysilicon 1857 -2187 1857 -2187 0 1
rlabel polysilicon 1857 -2193 1857 -2193 0 3
rlabel polysilicon 1864 -2187 1864 -2187 0 1
rlabel polysilicon 1864 -2193 1864 -2193 0 3
rlabel polysilicon 1871 -2187 1871 -2187 0 1
rlabel polysilicon 1871 -2193 1871 -2193 0 3
rlabel polysilicon 1878 -2187 1878 -2187 0 1
rlabel polysilicon 1878 -2193 1878 -2193 0 3
rlabel polysilicon 1885 -2187 1885 -2187 0 1
rlabel polysilicon 1885 -2193 1885 -2193 0 3
rlabel polysilicon 1892 -2187 1892 -2187 0 1
rlabel polysilicon 1892 -2193 1892 -2193 0 3
rlabel polysilicon 1899 -2187 1899 -2187 0 1
rlabel polysilicon 1899 -2193 1899 -2193 0 3
rlabel polysilicon 1906 -2187 1906 -2187 0 1
rlabel polysilicon 1906 -2193 1906 -2193 0 3
rlabel polysilicon 1913 -2187 1913 -2187 0 1
rlabel polysilicon 1913 -2193 1913 -2193 0 3
rlabel polysilicon 9 -2316 9 -2316 0 1
rlabel polysilicon 9 -2322 9 -2322 0 3
rlabel polysilicon 16 -2316 16 -2316 0 1
rlabel polysilicon 16 -2322 16 -2322 0 3
rlabel polysilicon 23 -2316 23 -2316 0 1
rlabel polysilicon 23 -2322 23 -2322 0 3
rlabel polysilicon 30 -2316 30 -2316 0 1
rlabel polysilicon 30 -2322 30 -2322 0 3
rlabel polysilicon 37 -2316 37 -2316 0 1
rlabel polysilicon 37 -2322 37 -2322 0 3
rlabel polysilicon 44 -2316 44 -2316 0 1
rlabel polysilicon 44 -2322 44 -2322 0 3
rlabel polysilicon 51 -2316 51 -2316 0 1
rlabel polysilicon 51 -2322 51 -2322 0 3
rlabel polysilicon 58 -2316 58 -2316 0 1
rlabel polysilicon 58 -2322 58 -2322 0 3
rlabel polysilicon 65 -2316 65 -2316 0 1
rlabel polysilicon 68 -2316 68 -2316 0 2
rlabel polysilicon 72 -2316 72 -2316 0 1
rlabel polysilicon 72 -2322 72 -2322 0 3
rlabel polysilicon 79 -2316 79 -2316 0 1
rlabel polysilicon 79 -2322 79 -2322 0 3
rlabel polysilicon 86 -2316 86 -2316 0 1
rlabel polysilicon 86 -2322 86 -2322 0 3
rlabel polysilicon 93 -2316 93 -2316 0 1
rlabel polysilicon 93 -2322 93 -2322 0 3
rlabel polysilicon 100 -2316 100 -2316 0 1
rlabel polysilicon 100 -2322 100 -2322 0 3
rlabel polysilicon 107 -2316 107 -2316 0 1
rlabel polysilicon 107 -2322 107 -2322 0 3
rlabel polysilicon 117 -2316 117 -2316 0 2
rlabel polysilicon 114 -2322 114 -2322 0 3
rlabel polysilicon 117 -2322 117 -2322 0 4
rlabel polysilicon 121 -2316 121 -2316 0 1
rlabel polysilicon 124 -2316 124 -2316 0 2
rlabel polysilicon 124 -2322 124 -2322 0 4
rlabel polysilicon 128 -2316 128 -2316 0 1
rlabel polysilicon 128 -2322 128 -2322 0 3
rlabel polysilicon 135 -2316 135 -2316 0 1
rlabel polysilicon 135 -2322 135 -2322 0 3
rlabel polysilicon 142 -2316 142 -2316 0 1
rlabel polysilicon 142 -2322 142 -2322 0 3
rlabel polysilicon 149 -2316 149 -2316 0 1
rlabel polysilicon 149 -2322 149 -2322 0 3
rlabel polysilicon 156 -2316 156 -2316 0 1
rlabel polysilicon 159 -2316 159 -2316 0 2
rlabel polysilicon 156 -2322 156 -2322 0 3
rlabel polysilicon 159 -2322 159 -2322 0 4
rlabel polysilicon 163 -2316 163 -2316 0 1
rlabel polysilicon 163 -2322 163 -2322 0 3
rlabel polysilicon 170 -2316 170 -2316 0 1
rlabel polysilicon 173 -2316 173 -2316 0 2
rlabel polysilicon 170 -2322 170 -2322 0 3
rlabel polysilicon 177 -2316 177 -2316 0 1
rlabel polysilicon 177 -2322 177 -2322 0 3
rlabel polysilicon 184 -2316 184 -2316 0 1
rlabel polysilicon 184 -2322 184 -2322 0 3
rlabel polysilicon 191 -2316 191 -2316 0 1
rlabel polysilicon 191 -2322 191 -2322 0 3
rlabel polysilicon 198 -2316 198 -2316 0 1
rlabel polysilicon 198 -2322 198 -2322 0 3
rlabel polysilicon 205 -2316 205 -2316 0 1
rlabel polysilicon 208 -2316 208 -2316 0 2
rlabel polysilicon 205 -2322 205 -2322 0 3
rlabel polysilicon 212 -2316 212 -2316 0 1
rlabel polysilicon 215 -2316 215 -2316 0 2
rlabel polysilicon 212 -2322 212 -2322 0 3
rlabel polysilicon 215 -2322 215 -2322 0 4
rlabel polysilicon 219 -2316 219 -2316 0 1
rlabel polysilicon 222 -2316 222 -2316 0 2
rlabel polysilicon 219 -2322 219 -2322 0 3
rlabel polysilicon 226 -2316 226 -2316 0 1
rlabel polysilicon 226 -2322 226 -2322 0 3
rlabel polysilicon 236 -2316 236 -2316 0 2
rlabel polysilicon 236 -2322 236 -2322 0 4
rlabel polysilicon 240 -2316 240 -2316 0 1
rlabel polysilicon 240 -2322 240 -2322 0 3
rlabel polysilicon 243 -2322 243 -2322 0 4
rlabel polysilicon 247 -2316 247 -2316 0 1
rlabel polysilicon 247 -2322 247 -2322 0 3
rlabel polysilicon 254 -2316 254 -2316 0 1
rlabel polysilicon 254 -2322 254 -2322 0 3
rlabel polysilicon 261 -2316 261 -2316 0 1
rlabel polysilicon 261 -2322 261 -2322 0 3
rlabel polysilicon 268 -2316 268 -2316 0 1
rlabel polysilicon 268 -2322 268 -2322 0 3
rlabel polysilicon 275 -2316 275 -2316 0 1
rlabel polysilicon 275 -2322 275 -2322 0 3
rlabel polysilicon 282 -2316 282 -2316 0 1
rlabel polysilicon 282 -2322 282 -2322 0 3
rlabel polysilicon 289 -2316 289 -2316 0 1
rlabel polysilicon 289 -2322 289 -2322 0 3
rlabel polysilicon 296 -2316 296 -2316 0 1
rlabel polysilicon 296 -2322 296 -2322 0 3
rlabel polysilicon 303 -2316 303 -2316 0 1
rlabel polysilicon 303 -2322 303 -2322 0 3
rlabel polysilicon 310 -2316 310 -2316 0 1
rlabel polysilicon 310 -2322 310 -2322 0 3
rlabel polysilicon 317 -2316 317 -2316 0 1
rlabel polysilicon 317 -2322 317 -2322 0 3
rlabel polysilicon 324 -2316 324 -2316 0 1
rlabel polysilicon 324 -2322 324 -2322 0 3
rlabel polysilicon 331 -2316 331 -2316 0 1
rlabel polysilicon 331 -2322 331 -2322 0 3
rlabel polysilicon 338 -2316 338 -2316 0 1
rlabel polysilicon 338 -2322 338 -2322 0 3
rlabel polysilicon 345 -2316 345 -2316 0 1
rlabel polysilicon 345 -2322 345 -2322 0 3
rlabel polysilicon 352 -2316 352 -2316 0 1
rlabel polysilicon 352 -2322 352 -2322 0 3
rlabel polysilicon 359 -2316 359 -2316 0 1
rlabel polysilicon 359 -2322 359 -2322 0 3
rlabel polysilicon 366 -2316 366 -2316 0 1
rlabel polysilicon 366 -2322 366 -2322 0 3
rlabel polysilicon 373 -2316 373 -2316 0 1
rlabel polysilicon 373 -2322 373 -2322 0 3
rlabel polysilicon 380 -2316 380 -2316 0 1
rlabel polysilicon 380 -2322 380 -2322 0 3
rlabel polysilicon 387 -2316 387 -2316 0 1
rlabel polysilicon 387 -2322 387 -2322 0 3
rlabel polysilicon 394 -2316 394 -2316 0 1
rlabel polysilicon 394 -2322 394 -2322 0 3
rlabel polysilicon 401 -2316 401 -2316 0 1
rlabel polysilicon 401 -2322 401 -2322 0 3
rlabel polysilicon 408 -2316 408 -2316 0 1
rlabel polysilicon 408 -2322 408 -2322 0 3
rlabel polysilicon 415 -2316 415 -2316 0 1
rlabel polysilicon 415 -2322 415 -2322 0 3
rlabel polysilicon 422 -2316 422 -2316 0 1
rlabel polysilicon 422 -2322 422 -2322 0 3
rlabel polysilicon 429 -2316 429 -2316 0 1
rlabel polysilicon 429 -2322 429 -2322 0 3
rlabel polysilicon 436 -2316 436 -2316 0 1
rlabel polysilicon 436 -2322 436 -2322 0 3
rlabel polysilicon 443 -2316 443 -2316 0 1
rlabel polysilicon 443 -2322 443 -2322 0 3
rlabel polysilicon 450 -2316 450 -2316 0 1
rlabel polysilicon 450 -2322 450 -2322 0 3
rlabel polysilicon 457 -2316 457 -2316 0 1
rlabel polysilicon 457 -2322 457 -2322 0 3
rlabel polysilicon 467 -2316 467 -2316 0 2
rlabel polysilicon 464 -2322 464 -2322 0 3
rlabel polysilicon 467 -2322 467 -2322 0 4
rlabel polysilicon 471 -2316 471 -2316 0 1
rlabel polysilicon 471 -2322 471 -2322 0 3
rlabel polysilicon 478 -2316 478 -2316 0 1
rlabel polysilicon 478 -2322 478 -2322 0 3
rlabel polysilicon 485 -2316 485 -2316 0 1
rlabel polysilicon 485 -2322 485 -2322 0 3
rlabel polysilicon 492 -2316 492 -2316 0 1
rlabel polysilicon 492 -2322 492 -2322 0 3
rlabel polysilicon 499 -2316 499 -2316 0 1
rlabel polysilicon 499 -2322 499 -2322 0 3
rlabel polysilicon 506 -2316 506 -2316 0 1
rlabel polysilicon 506 -2322 506 -2322 0 3
rlabel polysilicon 513 -2316 513 -2316 0 1
rlabel polysilicon 513 -2322 513 -2322 0 3
rlabel polysilicon 520 -2316 520 -2316 0 1
rlabel polysilicon 520 -2322 520 -2322 0 3
rlabel polysilicon 527 -2316 527 -2316 0 1
rlabel polysilicon 527 -2322 527 -2322 0 3
rlabel polysilicon 534 -2316 534 -2316 0 1
rlabel polysilicon 534 -2322 534 -2322 0 3
rlabel polysilicon 541 -2316 541 -2316 0 1
rlabel polysilicon 541 -2322 541 -2322 0 3
rlabel polysilicon 548 -2316 548 -2316 0 1
rlabel polysilicon 548 -2322 548 -2322 0 3
rlabel polysilicon 555 -2316 555 -2316 0 1
rlabel polysilicon 555 -2322 555 -2322 0 3
rlabel polysilicon 562 -2316 562 -2316 0 1
rlabel polysilicon 562 -2322 562 -2322 0 3
rlabel polysilicon 569 -2316 569 -2316 0 1
rlabel polysilicon 572 -2316 572 -2316 0 2
rlabel polysilicon 569 -2322 569 -2322 0 3
rlabel polysilicon 572 -2322 572 -2322 0 4
rlabel polysilicon 576 -2316 576 -2316 0 1
rlabel polysilicon 576 -2322 576 -2322 0 3
rlabel polysilicon 583 -2316 583 -2316 0 1
rlabel polysilicon 583 -2322 583 -2322 0 3
rlabel polysilicon 590 -2316 590 -2316 0 1
rlabel polysilicon 590 -2322 590 -2322 0 3
rlabel polysilicon 597 -2316 597 -2316 0 1
rlabel polysilicon 597 -2322 597 -2322 0 3
rlabel polysilicon 604 -2316 604 -2316 0 1
rlabel polysilicon 604 -2322 604 -2322 0 3
rlabel polysilicon 611 -2316 611 -2316 0 1
rlabel polysilicon 611 -2322 611 -2322 0 3
rlabel polysilicon 618 -2316 618 -2316 0 1
rlabel polysilicon 618 -2322 618 -2322 0 3
rlabel polysilicon 625 -2316 625 -2316 0 1
rlabel polysilicon 628 -2316 628 -2316 0 2
rlabel polysilicon 625 -2322 625 -2322 0 3
rlabel polysilicon 632 -2316 632 -2316 0 1
rlabel polysilicon 632 -2322 632 -2322 0 3
rlabel polysilicon 639 -2316 639 -2316 0 1
rlabel polysilicon 639 -2322 639 -2322 0 3
rlabel polysilicon 646 -2316 646 -2316 0 1
rlabel polysilicon 646 -2322 646 -2322 0 3
rlabel polysilicon 653 -2316 653 -2316 0 1
rlabel polysilicon 656 -2316 656 -2316 0 2
rlabel polysilicon 656 -2322 656 -2322 0 4
rlabel polysilicon 660 -2316 660 -2316 0 1
rlabel polysilicon 660 -2322 660 -2322 0 3
rlabel polysilicon 670 -2316 670 -2316 0 2
rlabel polysilicon 667 -2322 667 -2322 0 3
rlabel polysilicon 674 -2316 674 -2316 0 1
rlabel polysilicon 677 -2316 677 -2316 0 2
rlabel polysilicon 674 -2322 674 -2322 0 3
rlabel polysilicon 677 -2322 677 -2322 0 4
rlabel polysilicon 681 -2316 681 -2316 0 1
rlabel polysilicon 681 -2322 681 -2322 0 3
rlabel polysilicon 688 -2316 688 -2316 0 1
rlabel polysilicon 688 -2322 688 -2322 0 3
rlabel polysilicon 695 -2316 695 -2316 0 1
rlabel polysilicon 695 -2322 695 -2322 0 3
rlabel polysilicon 702 -2316 702 -2316 0 1
rlabel polysilicon 702 -2322 702 -2322 0 3
rlabel polysilicon 709 -2316 709 -2316 0 1
rlabel polysilicon 709 -2322 709 -2322 0 3
rlabel polysilicon 716 -2316 716 -2316 0 1
rlabel polysilicon 716 -2322 716 -2322 0 3
rlabel polysilicon 723 -2316 723 -2316 0 1
rlabel polysilicon 723 -2322 723 -2322 0 3
rlabel polysilicon 730 -2316 730 -2316 0 1
rlabel polysilicon 730 -2322 730 -2322 0 3
rlabel polysilicon 737 -2316 737 -2316 0 1
rlabel polysilicon 737 -2322 737 -2322 0 3
rlabel polysilicon 744 -2316 744 -2316 0 1
rlabel polysilicon 744 -2322 744 -2322 0 3
rlabel polysilicon 751 -2316 751 -2316 0 1
rlabel polysilicon 751 -2322 751 -2322 0 3
rlabel polysilicon 758 -2316 758 -2316 0 1
rlabel polysilicon 761 -2316 761 -2316 0 2
rlabel polysilicon 758 -2322 758 -2322 0 3
rlabel polysilicon 765 -2316 765 -2316 0 1
rlabel polysilicon 765 -2322 765 -2322 0 3
rlabel polysilicon 772 -2316 772 -2316 0 1
rlabel polysilicon 772 -2322 772 -2322 0 3
rlabel polysilicon 779 -2316 779 -2316 0 1
rlabel polysilicon 779 -2322 779 -2322 0 3
rlabel polysilicon 786 -2316 786 -2316 0 1
rlabel polysilicon 786 -2322 786 -2322 0 3
rlabel polysilicon 793 -2316 793 -2316 0 1
rlabel polysilicon 796 -2316 796 -2316 0 2
rlabel polysilicon 796 -2322 796 -2322 0 4
rlabel polysilicon 800 -2316 800 -2316 0 1
rlabel polysilicon 800 -2322 800 -2322 0 3
rlabel polysilicon 807 -2316 807 -2316 0 1
rlabel polysilicon 807 -2322 807 -2322 0 3
rlabel polysilicon 817 -2316 817 -2316 0 2
rlabel polysilicon 817 -2322 817 -2322 0 4
rlabel polysilicon 821 -2316 821 -2316 0 1
rlabel polysilicon 824 -2316 824 -2316 0 2
rlabel polysilicon 821 -2322 821 -2322 0 3
rlabel polysilicon 824 -2322 824 -2322 0 4
rlabel polysilicon 828 -2316 828 -2316 0 1
rlabel polysilicon 828 -2322 828 -2322 0 3
rlabel polysilicon 835 -2316 835 -2316 0 1
rlabel polysilicon 835 -2322 835 -2322 0 3
rlabel polysilicon 842 -2316 842 -2316 0 1
rlabel polysilicon 842 -2322 842 -2322 0 3
rlabel polysilicon 849 -2316 849 -2316 0 1
rlabel polysilicon 849 -2322 849 -2322 0 3
rlabel polysilicon 856 -2316 856 -2316 0 1
rlabel polysilicon 856 -2322 856 -2322 0 3
rlabel polysilicon 863 -2316 863 -2316 0 1
rlabel polysilicon 863 -2322 863 -2322 0 3
rlabel polysilicon 870 -2316 870 -2316 0 1
rlabel polysilicon 870 -2322 870 -2322 0 3
rlabel polysilicon 877 -2316 877 -2316 0 1
rlabel polysilicon 877 -2322 877 -2322 0 3
rlabel polysilicon 887 -2316 887 -2316 0 2
rlabel polysilicon 884 -2322 884 -2322 0 3
rlabel polysilicon 887 -2322 887 -2322 0 4
rlabel polysilicon 891 -2316 891 -2316 0 1
rlabel polysilicon 891 -2322 891 -2322 0 3
rlabel polysilicon 898 -2316 898 -2316 0 1
rlabel polysilicon 898 -2322 898 -2322 0 3
rlabel polysilicon 905 -2316 905 -2316 0 1
rlabel polysilicon 905 -2322 905 -2322 0 3
rlabel polysilicon 912 -2316 912 -2316 0 1
rlabel polysilicon 912 -2322 912 -2322 0 3
rlabel polysilicon 919 -2316 919 -2316 0 1
rlabel polysilicon 919 -2322 919 -2322 0 3
rlabel polysilicon 926 -2316 926 -2316 0 1
rlabel polysilicon 926 -2322 926 -2322 0 3
rlabel polysilicon 933 -2316 933 -2316 0 1
rlabel polysilicon 933 -2322 933 -2322 0 3
rlabel polysilicon 940 -2316 940 -2316 0 1
rlabel polysilicon 940 -2322 940 -2322 0 3
rlabel polysilicon 947 -2316 947 -2316 0 1
rlabel polysilicon 950 -2316 950 -2316 0 2
rlabel polysilicon 947 -2322 947 -2322 0 3
rlabel polysilicon 950 -2322 950 -2322 0 4
rlabel polysilicon 954 -2316 954 -2316 0 1
rlabel polysilicon 954 -2322 954 -2322 0 3
rlabel polysilicon 961 -2316 961 -2316 0 1
rlabel polysilicon 961 -2322 961 -2322 0 3
rlabel polysilicon 968 -2316 968 -2316 0 1
rlabel polysilicon 968 -2322 968 -2322 0 3
rlabel polysilicon 975 -2316 975 -2316 0 1
rlabel polysilicon 975 -2322 975 -2322 0 3
rlabel polysilicon 982 -2316 982 -2316 0 1
rlabel polysilicon 982 -2322 982 -2322 0 3
rlabel polysilicon 989 -2316 989 -2316 0 1
rlabel polysilicon 989 -2322 989 -2322 0 3
rlabel polysilicon 996 -2316 996 -2316 0 1
rlabel polysilicon 999 -2316 999 -2316 0 2
rlabel polysilicon 996 -2322 996 -2322 0 3
rlabel polysilicon 999 -2322 999 -2322 0 4
rlabel polysilicon 1003 -2316 1003 -2316 0 1
rlabel polysilicon 1003 -2322 1003 -2322 0 3
rlabel polysilicon 1010 -2316 1010 -2316 0 1
rlabel polysilicon 1010 -2322 1010 -2322 0 3
rlabel polysilicon 1017 -2316 1017 -2316 0 1
rlabel polysilicon 1017 -2322 1017 -2322 0 3
rlabel polysilicon 1024 -2316 1024 -2316 0 1
rlabel polysilicon 1024 -2322 1024 -2322 0 3
rlabel polysilicon 1031 -2316 1031 -2316 0 1
rlabel polysilicon 1031 -2322 1031 -2322 0 3
rlabel polysilicon 1038 -2316 1038 -2316 0 1
rlabel polysilicon 1038 -2322 1038 -2322 0 3
rlabel polysilicon 1045 -2316 1045 -2316 0 1
rlabel polysilicon 1045 -2322 1045 -2322 0 3
rlabel polysilicon 1052 -2316 1052 -2316 0 1
rlabel polysilicon 1052 -2322 1052 -2322 0 3
rlabel polysilicon 1059 -2316 1059 -2316 0 1
rlabel polysilicon 1059 -2322 1059 -2322 0 3
rlabel polysilicon 1069 -2316 1069 -2316 0 2
rlabel polysilicon 1066 -2322 1066 -2322 0 3
rlabel polysilicon 1069 -2322 1069 -2322 0 4
rlabel polysilicon 1073 -2316 1073 -2316 0 1
rlabel polysilicon 1073 -2322 1073 -2322 0 3
rlabel polysilicon 1080 -2316 1080 -2316 0 1
rlabel polysilicon 1080 -2322 1080 -2322 0 3
rlabel polysilicon 1087 -2316 1087 -2316 0 1
rlabel polysilicon 1087 -2322 1087 -2322 0 3
rlabel polysilicon 1094 -2316 1094 -2316 0 1
rlabel polysilicon 1094 -2322 1094 -2322 0 3
rlabel polysilicon 1101 -2316 1101 -2316 0 1
rlabel polysilicon 1101 -2322 1101 -2322 0 3
rlabel polysilicon 1108 -2316 1108 -2316 0 1
rlabel polysilicon 1108 -2322 1108 -2322 0 3
rlabel polysilicon 1115 -2316 1115 -2316 0 1
rlabel polysilicon 1115 -2322 1115 -2322 0 3
rlabel polysilicon 1118 -2322 1118 -2322 0 4
rlabel polysilicon 1122 -2316 1122 -2316 0 1
rlabel polysilicon 1125 -2316 1125 -2316 0 2
rlabel polysilicon 1122 -2322 1122 -2322 0 3
rlabel polysilicon 1129 -2316 1129 -2316 0 1
rlabel polysilicon 1129 -2322 1129 -2322 0 3
rlabel polysilicon 1136 -2316 1136 -2316 0 1
rlabel polysilicon 1136 -2322 1136 -2322 0 3
rlabel polysilicon 1143 -2316 1143 -2316 0 1
rlabel polysilicon 1143 -2322 1143 -2322 0 3
rlabel polysilicon 1150 -2316 1150 -2316 0 1
rlabel polysilicon 1150 -2322 1150 -2322 0 3
rlabel polysilicon 1157 -2316 1157 -2316 0 1
rlabel polysilicon 1157 -2322 1157 -2322 0 3
rlabel polysilicon 1164 -2316 1164 -2316 0 1
rlabel polysilicon 1164 -2322 1164 -2322 0 3
rlabel polysilicon 1171 -2316 1171 -2316 0 1
rlabel polysilicon 1171 -2322 1171 -2322 0 3
rlabel polysilicon 1178 -2316 1178 -2316 0 1
rlabel polysilicon 1178 -2322 1178 -2322 0 3
rlabel polysilicon 1185 -2316 1185 -2316 0 1
rlabel polysilicon 1188 -2316 1188 -2316 0 2
rlabel polysilicon 1185 -2322 1185 -2322 0 3
rlabel polysilicon 1188 -2322 1188 -2322 0 4
rlabel polysilicon 1192 -2316 1192 -2316 0 1
rlabel polysilicon 1192 -2322 1192 -2322 0 3
rlabel polysilicon 1199 -2316 1199 -2316 0 1
rlabel polysilicon 1199 -2322 1199 -2322 0 3
rlabel polysilicon 1206 -2316 1206 -2316 0 1
rlabel polysilicon 1206 -2322 1206 -2322 0 3
rlabel polysilicon 1213 -2316 1213 -2316 0 1
rlabel polysilicon 1213 -2322 1213 -2322 0 3
rlabel polysilicon 1220 -2316 1220 -2316 0 1
rlabel polysilicon 1220 -2322 1220 -2322 0 3
rlabel polysilicon 1227 -2316 1227 -2316 0 1
rlabel polysilicon 1227 -2322 1227 -2322 0 3
rlabel polysilicon 1234 -2316 1234 -2316 0 1
rlabel polysilicon 1234 -2322 1234 -2322 0 3
rlabel polysilicon 1241 -2316 1241 -2316 0 1
rlabel polysilicon 1241 -2322 1241 -2322 0 3
rlabel polysilicon 1248 -2316 1248 -2316 0 1
rlabel polysilicon 1248 -2322 1248 -2322 0 3
rlabel polysilicon 1255 -2316 1255 -2316 0 1
rlabel polysilicon 1255 -2322 1255 -2322 0 3
rlabel polysilicon 1262 -2316 1262 -2316 0 1
rlabel polysilicon 1262 -2322 1262 -2322 0 3
rlabel polysilicon 1269 -2316 1269 -2316 0 1
rlabel polysilicon 1269 -2322 1269 -2322 0 3
rlabel polysilicon 1276 -2316 1276 -2316 0 1
rlabel polysilicon 1276 -2322 1276 -2322 0 3
rlabel polysilicon 1283 -2316 1283 -2316 0 1
rlabel polysilicon 1283 -2322 1283 -2322 0 3
rlabel polysilicon 1290 -2316 1290 -2316 0 1
rlabel polysilicon 1293 -2316 1293 -2316 0 2
rlabel polysilicon 1290 -2322 1290 -2322 0 3
rlabel polysilicon 1293 -2322 1293 -2322 0 4
rlabel polysilicon 1297 -2316 1297 -2316 0 1
rlabel polysilicon 1297 -2322 1297 -2322 0 3
rlabel polysilicon 1304 -2316 1304 -2316 0 1
rlabel polysilicon 1304 -2322 1304 -2322 0 3
rlabel polysilicon 1307 -2322 1307 -2322 0 4
rlabel polysilicon 1311 -2316 1311 -2316 0 1
rlabel polysilicon 1311 -2322 1311 -2322 0 3
rlabel polysilicon 1318 -2316 1318 -2316 0 1
rlabel polysilicon 1318 -2322 1318 -2322 0 3
rlabel polysilicon 1325 -2316 1325 -2316 0 1
rlabel polysilicon 1325 -2322 1325 -2322 0 3
rlabel polysilicon 1332 -2316 1332 -2316 0 1
rlabel polysilicon 1332 -2322 1332 -2322 0 3
rlabel polysilicon 1339 -2316 1339 -2316 0 1
rlabel polysilicon 1339 -2322 1339 -2322 0 3
rlabel polysilicon 1346 -2316 1346 -2316 0 1
rlabel polysilicon 1346 -2322 1346 -2322 0 3
rlabel polysilicon 1353 -2316 1353 -2316 0 1
rlabel polysilicon 1353 -2322 1353 -2322 0 3
rlabel polysilicon 1360 -2316 1360 -2316 0 1
rlabel polysilicon 1360 -2322 1360 -2322 0 3
rlabel polysilicon 1367 -2316 1367 -2316 0 1
rlabel polysilicon 1367 -2322 1367 -2322 0 3
rlabel polysilicon 1370 -2322 1370 -2322 0 4
rlabel polysilicon 1374 -2316 1374 -2316 0 1
rlabel polysilicon 1374 -2322 1374 -2322 0 3
rlabel polysilicon 1381 -2316 1381 -2316 0 1
rlabel polysilicon 1381 -2322 1381 -2322 0 3
rlabel polysilicon 1388 -2316 1388 -2316 0 1
rlabel polysilicon 1388 -2322 1388 -2322 0 3
rlabel polysilicon 1395 -2316 1395 -2316 0 1
rlabel polysilicon 1395 -2322 1395 -2322 0 3
rlabel polysilicon 1402 -2316 1402 -2316 0 1
rlabel polysilicon 1402 -2322 1402 -2322 0 3
rlabel polysilicon 1409 -2316 1409 -2316 0 1
rlabel polysilicon 1409 -2322 1409 -2322 0 3
rlabel polysilicon 1416 -2316 1416 -2316 0 1
rlabel polysilicon 1416 -2322 1416 -2322 0 3
rlabel polysilicon 1423 -2316 1423 -2316 0 1
rlabel polysilicon 1423 -2322 1423 -2322 0 3
rlabel polysilicon 1430 -2316 1430 -2316 0 1
rlabel polysilicon 1430 -2322 1430 -2322 0 3
rlabel polysilicon 1437 -2316 1437 -2316 0 1
rlabel polysilicon 1437 -2322 1437 -2322 0 3
rlabel polysilicon 1444 -2316 1444 -2316 0 1
rlabel polysilicon 1444 -2322 1444 -2322 0 3
rlabel polysilicon 1451 -2316 1451 -2316 0 1
rlabel polysilicon 1451 -2322 1451 -2322 0 3
rlabel polysilicon 1458 -2316 1458 -2316 0 1
rlabel polysilicon 1458 -2322 1458 -2322 0 3
rlabel polysilicon 1465 -2316 1465 -2316 0 1
rlabel polysilicon 1465 -2322 1465 -2322 0 3
rlabel polysilicon 1472 -2316 1472 -2316 0 1
rlabel polysilicon 1472 -2322 1472 -2322 0 3
rlabel polysilicon 1479 -2316 1479 -2316 0 1
rlabel polysilicon 1479 -2322 1479 -2322 0 3
rlabel polysilicon 1486 -2316 1486 -2316 0 1
rlabel polysilicon 1486 -2322 1486 -2322 0 3
rlabel polysilicon 1493 -2316 1493 -2316 0 1
rlabel polysilicon 1493 -2322 1493 -2322 0 3
rlabel polysilicon 1500 -2316 1500 -2316 0 1
rlabel polysilicon 1500 -2322 1500 -2322 0 3
rlabel polysilicon 1507 -2316 1507 -2316 0 1
rlabel polysilicon 1507 -2322 1507 -2322 0 3
rlabel polysilicon 1514 -2316 1514 -2316 0 1
rlabel polysilicon 1514 -2322 1514 -2322 0 3
rlabel polysilicon 1521 -2316 1521 -2316 0 1
rlabel polysilicon 1521 -2322 1521 -2322 0 3
rlabel polysilicon 1528 -2316 1528 -2316 0 1
rlabel polysilicon 1528 -2322 1528 -2322 0 3
rlabel polysilicon 1535 -2316 1535 -2316 0 1
rlabel polysilicon 1535 -2322 1535 -2322 0 3
rlabel polysilicon 1542 -2316 1542 -2316 0 1
rlabel polysilicon 1542 -2322 1542 -2322 0 3
rlabel polysilicon 1549 -2316 1549 -2316 0 1
rlabel polysilicon 1549 -2322 1549 -2322 0 3
rlabel polysilicon 1556 -2316 1556 -2316 0 1
rlabel polysilicon 1556 -2322 1556 -2322 0 3
rlabel polysilicon 1563 -2316 1563 -2316 0 1
rlabel polysilicon 1563 -2322 1563 -2322 0 3
rlabel polysilicon 1570 -2316 1570 -2316 0 1
rlabel polysilicon 1570 -2322 1570 -2322 0 3
rlabel polysilicon 1577 -2316 1577 -2316 0 1
rlabel polysilicon 1577 -2322 1577 -2322 0 3
rlabel polysilicon 1584 -2316 1584 -2316 0 1
rlabel polysilicon 1584 -2322 1584 -2322 0 3
rlabel polysilicon 1591 -2316 1591 -2316 0 1
rlabel polysilicon 1591 -2322 1591 -2322 0 3
rlabel polysilicon 1598 -2316 1598 -2316 0 1
rlabel polysilicon 1598 -2322 1598 -2322 0 3
rlabel polysilicon 1605 -2316 1605 -2316 0 1
rlabel polysilicon 1605 -2322 1605 -2322 0 3
rlabel polysilicon 1612 -2316 1612 -2316 0 1
rlabel polysilicon 1612 -2322 1612 -2322 0 3
rlabel polysilicon 1619 -2316 1619 -2316 0 1
rlabel polysilicon 1619 -2322 1619 -2322 0 3
rlabel polysilicon 1626 -2316 1626 -2316 0 1
rlabel polysilicon 1626 -2322 1626 -2322 0 3
rlabel polysilicon 1633 -2316 1633 -2316 0 1
rlabel polysilicon 1633 -2322 1633 -2322 0 3
rlabel polysilicon 1640 -2316 1640 -2316 0 1
rlabel polysilicon 1640 -2322 1640 -2322 0 3
rlabel polysilicon 1647 -2316 1647 -2316 0 1
rlabel polysilicon 1647 -2322 1647 -2322 0 3
rlabel polysilicon 1654 -2316 1654 -2316 0 1
rlabel polysilicon 1654 -2322 1654 -2322 0 3
rlabel polysilicon 1661 -2316 1661 -2316 0 1
rlabel polysilicon 1661 -2322 1661 -2322 0 3
rlabel polysilicon 1668 -2316 1668 -2316 0 1
rlabel polysilicon 1668 -2322 1668 -2322 0 3
rlabel polysilicon 1675 -2316 1675 -2316 0 1
rlabel polysilicon 1675 -2322 1675 -2322 0 3
rlabel polysilicon 1682 -2316 1682 -2316 0 1
rlabel polysilicon 1682 -2322 1682 -2322 0 3
rlabel polysilicon 1689 -2316 1689 -2316 0 1
rlabel polysilicon 1689 -2322 1689 -2322 0 3
rlabel polysilicon 1696 -2316 1696 -2316 0 1
rlabel polysilicon 1696 -2322 1696 -2322 0 3
rlabel polysilicon 1703 -2316 1703 -2316 0 1
rlabel polysilicon 1703 -2322 1703 -2322 0 3
rlabel polysilicon 1710 -2316 1710 -2316 0 1
rlabel polysilicon 1713 -2316 1713 -2316 0 2
rlabel polysilicon 1713 -2322 1713 -2322 0 4
rlabel polysilicon 1717 -2316 1717 -2316 0 1
rlabel polysilicon 1717 -2322 1717 -2322 0 3
rlabel polysilicon 1727 -2316 1727 -2316 0 2
rlabel polysilicon 1727 -2322 1727 -2322 0 4
rlabel polysilicon 1731 -2316 1731 -2316 0 1
rlabel polysilicon 1731 -2322 1731 -2322 0 3
rlabel polysilicon 1738 -2316 1738 -2316 0 1
rlabel polysilicon 1738 -2322 1738 -2322 0 3
rlabel polysilicon 1745 -2316 1745 -2316 0 1
rlabel polysilicon 1748 -2322 1748 -2322 0 4
rlabel polysilicon 1752 -2316 1752 -2316 0 1
rlabel polysilicon 1752 -2322 1752 -2322 0 3
rlabel polysilicon 1759 -2316 1759 -2316 0 1
rlabel polysilicon 1759 -2322 1759 -2322 0 3
rlabel polysilicon 1766 -2316 1766 -2316 0 1
rlabel polysilicon 1766 -2322 1766 -2322 0 3
rlabel polysilicon 1773 -2316 1773 -2316 0 1
rlabel polysilicon 1773 -2322 1773 -2322 0 3
rlabel polysilicon 1780 -2316 1780 -2316 0 1
rlabel polysilicon 1780 -2322 1780 -2322 0 3
rlabel polysilicon 1787 -2316 1787 -2316 0 1
rlabel polysilicon 1787 -2322 1787 -2322 0 3
rlabel polysilicon 1794 -2316 1794 -2316 0 1
rlabel polysilicon 1794 -2322 1794 -2322 0 3
rlabel polysilicon 1822 -2316 1822 -2316 0 1
rlabel polysilicon 1822 -2322 1822 -2322 0 3
rlabel polysilicon 1829 -2316 1829 -2316 0 1
rlabel polysilicon 1829 -2322 1829 -2322 0 3
rlabel polysilicon 9 -2441 9 -2441 0 1
rlabel polysilicon 9 -2447 9 -2447 0 3
rlabel polysilicon 16 -2441 16 -2441 0 1
rlabel polysilicon 16 -2447 16 -2447 0 3
rlabel polysilicon 30 -2441 30 -2441 0 1
rlabel polysilicon 30 -2447 30 -2447 0 3
rlabel polysilicon 37 -2441 37 -2441 0 1
rlabel polysilicon 37 -2447 37 -2447 0 3
rlabel polysilicon 44 -2441 44 -2441 0 1
rlabel polysilicon 44 -2447 44 -2447 0 3
rlabel polysilicon 51 -2441 51 -2441 0 1
rlabel polysilicon 51 -2447 51 -2447 0 3
rlabel polysilicon 58 -2441 58 -2441 0 1
rlabel polysilicon 58 -2447 58 -2447 0 3
rlabel polysilicon 65 -2441 65 -2441 0 1
rlabel polysilicon 65 -2447 65 -2447 0 3
rlabel polysilicon 72 -2441 72 -2441 0 1
rlabel polysilicon 72 -2447 72 -2447 0 3
rlabel polysilicon 82 -2441 82 -2441 0 2
rlabel polysilicon 79 -2447 79 -2447 0 3
rlabel polysilicon 82 -2447 82 -2447 0 4
rlabel polysilicon 86 -2441 86 -2441 0 1
rlabel polysilicon 86 -2447 86 -2447 0 3
rlabel polysilicon 93 -2441 93 -2441 0 1
rlabel polysilicon 96 -2441 96 -2441 0 2
rlabel polysilicon 93 -2447 93 -2447 0 3
rlabel polysilicon 96 -2447 96 -2447 0 4
rlabel polysilicon 100 -2441 100 -2441 0 1
rlabel polysilicon 100 -2447 100 -2447 0 3
rlabel polysilicon 107 -2441 107 -2441 0 1
rlabel polysilicon 110 -2441 110 -2441 0 2
rlabel polysilicon 107 -2447 107 -2447 0 3
rlabel polysilicon 110 -2447 110 -2447 0 4
rlabel polysilicon 114 -2441 114 -2441 0 1
rlabel polysilicon 114 -2447 114 -2447 0 3
rlabel polysilicon 121 -2441 121 -2441 0 1
rlabel polysilicon 121 -2447 121 -2447 0 3
rlabel polysilicon 128 -2441 128 -2441 0 1
rlabel polysilicon 131 -2441 131 -2441 0 2
rlabel polysilicon 128 -2447 128 -2447 0 3
rlabel polysilicon 131 -2447 131 -2447 0 4
rlabel polysilicon 135 -2441 135 -2441 0 1
rlabel polysilicon 135 -2447 135 -2447 0 3
rlabel polysilicon 142 -2441 142 -2441 0 1
rlabel polysilicon 142 -2447 142 -2447 0 3
rlabel polysilicon 149 -2441 149 -2441 0 1
rlabel polysilicon 149 -2447 149 -2447 0 3
rlabel polysilicon 156 -2441 156 -2441 0 1
rlabel polysilicon 156 -2447 156 -2447 0 3
rlabel polysilicon 163 -2441 163 -2441 0 1
rlabel polysilicon 163 -2447 163 -2447 0 3
rlabel polysilicon 170 -2441 170 -2441 0 1
rlabel polysilicon 170 -2447 170 -2447 0 3
rlabel polysilicon 177 -2441 177 -2441 0 1
rlabel polysilicon 177 -2447 177 -2447 0 3
rlabel polysilicon 184 -2441 184 -2441 0 1
rlabel polysilicon 184 -2447 184 -2447 0 3
rlabel polysilicon 191 -2441 191 -2441 0 1
rlabel polysilicon 191 -2447 191 -2447 0 3
rlabel polysilicon 194 -2447 194 -2447 0 4
rlabel polysilicon 198 -2441 198 -2441 0 1
rlabel polysilicon 198 -2447 198 -2447 0 3
rlabel polysilicon 205 -2441 205 -2441 0 1
rlabel polysilicon 205 -2447 205 -2447 0 3
rlabel polysilicon 212 -2441 212 -2441 0 1
rlabel polysilicon 212 -2447 212 -2447 0 3
rlabel polysilicon 219 -2441 219 -2441 0 1
rlabel polysilicon 219 -2447 219 -2447 0 3
rlabel polysilicon 226 -2441 226 -2441 0 1
rlabel polysilicon 226 -2447 226 -2447 0 3
rlabel polysilicon 233 -2441 233 -2441 0 1
rlabel polysilicon 233 -2447 233 -2447 0 3
rlabel polysilicon 240 -2441 240 -2441 0 1
rlabel polysilicon 240 -2447 240 -2447 0 3
rlabel polysilicon 247 -2441 247 -2441 0 1
rlabel polysilicon 247 -2447 247 -2447 0 3
rlabel polysilicon 254 -2441 254 -2441 0 1
rlabel polysilicon 254 -2447 254 -2447 0 3
rlabel polysilicon 261 -2441 261 -2441 0 1
rlabel polysilicon 261 -2447 261 -2447 0 3
rlabel polysilicon 268 -2441 268 -2441 0 1
rlabel polysilicon 268 -2447 268 -2447 0 3
rlabel polysilicon 275 -2441 275 -2441 0 1
rlabel polysilicon 275 -2447 275 -2447 0 3
rlabel polysilicon 282 -2441 282 -2441 0 1
rlabel polysilicon 282 -2447 282 -2447 0 3
rlabel polysilicon 289 -2441 289 -2441 0 1
rlabel polysilicon 289 -2447 289 -2447 0 3
rlabel polysilicon 296 -2441 296 -2441 0 1
rlabel polysilicon 296 -2447 296 -2447 0 3
rlabel polysilicon 303 -2441 303 -2441 0 1
rlabel polysilicon 303 -2447 303 -2447 0 3
rlabel polysilicon 310 -2441 310 -2441 0 1
rlabel polysilicon 310 -2447 310 -2447 0 3
rlabel polysilicon 317 -2441 317 -2441 0 1
rlabel polysilicon 317 -2447 317 -2447 0 3
rlabel polysilicon 324 -2441 324 -2441 0 1
rlabel polysilicon 324 -2447 324 -2447 0 3
rlabel polysilicon 331 -2441 331 -2441 0 1
rlabel polysilicon 331 -2447 331 -2447 0 3
rlabel polysilicon 338 -2441 338 -2441 0 1
rlabel polysilicon 341 -2441 341 -2441 0 2
rlabel polysilicon 338 -2447 338 -2447 0 3
rlabel polysilicon 341 -2447 341 -2447 0 4
rlabel polysilicon 345 -2441 345 -2441 0 1
rlabel polysilicon 345 -2447 345 -2447 0 3
rlabel polysilicon 352 -2441 352 -2441 0 1
rlabel polysilicon 352 -2447 352 -2447 0 3
rlabel polysilicon 359 -2441 359 -2441 0 1
rlabel polysilicon 359 -2447 359 -2447 0 3
rlabel polysilicon 366 -2441 366 -2441 0 1
rlabel polysilicon 366 -2447 366 -2447 0 3
rlabel polysilicon 373 -2441 373 -2441 0 1
rlabel polysilicon 373 -2447 373 -2447 0 3
rlabel polysilicon 380 -2441 380 -2441 0 1
rlabel polysilicon 380 -2447 380 -2447 0 3
rlabel polysilicon 387 -2441 387 -2441 0 1
rlabel polysilicon 390 -2441 390 -2441 0 2
rlabel polysilicon 387 -2447 387 -2447 0 3
rlabel polysilicon 390 -2447 390 -2447 0 4
rlabel polysilicon 394 -2441 394 -2441 0 1
rlabel polysilicon 394 -2447 394 -2447 0 3
rlabel polysilicon 401 -2441 401 -2441 0 1
rlabel polysilicon 404 -2441 404 -2441 0 2
rlabel polysilicon 401 -2447 401 -2447 0 3
rlabel polysilicon 404 -2447 404 -2447 0 4
rlabel polysilicon 408 -2441 408 -2441 0 1
rlabel polysilicon 408 -2447 408 -2447 0 3
rlabel polysilicon 415 -2441 415 -2441 0 1
rlabel polysilicon 415 -2447 415 -2447 0 3
rlabel polysilicon 422 -2441 422 -2441 0 1
rlabel polysilicon 422 -2447 422 -2447 0 3
rlabel polysilicon 429 -2441 429 -2441 0 1
rlabel polysilicon 432 -2441 432 -2441 0 2
rlabel polysilicon 432 -2447 432 -2447 0 4
rlabel polysilicon 436 -2441 436 -2441 0 1
rlabel polysilicon 439 -2441 439 -2441 0 2
rlabel polysilicon 436 -2447 436 -2447 0 3
rlabel polysilicon 439 -2447 439 -2447 0 4
rlabel polysilicon 443 -2441 443 -2441 0 1
rlabel polysilicon 446 -2441 446 -2441 0 2
rlabel polysilicon 443 -2447 443 -2447 0 3
rlabel polysilicon 450 -2441 450 -2441 0 1
rlabel polysilicon 450 -2447 450 -2447 0 3
rlabel polysilicon 457 -2441 457 -2441 0 1
rlabel polysilicon 460 -2441 460 -2441 0 2
rlabel polysilicon 457 -2447 457 -2447 0 3
rlabel polysilicon 460 -2447 460 -2447 0 4
rlabel polysilicon 464 -2441 464 -2441 0 1
rlabel polysilicon 464 -2447 464 -2447 0 3
rlabel polysilicon 471 -2441 471 -2441 0 1
rlabel polysilicon 471 -2447 471 -2447 0 3
rlabel polysilicon 478 -2441 478 -2441 0 1
rlabel polysilicon 478 -2447 478 -2447 0 3
rlabel polysilicon 485 -2441 485 -2441 0 1
rlabel polysilicon 485 -2447 485 -2447 0 3
rlabel polysilicon 492 -2441 492 -2441 0 1
rlabel polysilicon 492 -2447 492 -2447 0 3
rlabel polysilicon 499 -2441 499 -2441 0 1
rlabel polysilicon 499 -2447 499 -2447 0 3
rlabel polysilicon 506 -2441 506 -2441 0 1
rlabel polysilicon 506 -2447 506 -2447 0 3
rlabel polysilicon 513 -2441 513 -2441 0 1
rlabel polysilicon 513 -2447 513 -2447 0 3
rlabel polysilicon 516 -2447 516 -2447 0 4
rlabel polysilicon 520 -2441 520 -2441 0 1
rlabel polysilicon 520 -2447 520 -2447 0 3
rlabel polysilicon 527 -2441 527 -2441 0 1
rlabel polysilicon 530 -2441 530 -2441 0 2
rlabel polysilicon 527 -2447 527 -2447 0 3
rlabel polysilicon 530 -2447 530 -2447 0 4
rlabel polysilicon 534 -2441 534 -2441 0 1
rlabel polysilicon 534 -2447 534 -2447 0 3
rlabel polysilicon 541 -2441 541 -2441 0 1
rlabel polysilicon 544 -2441 544 -2441 0 2
rlabel polysilicon 544 -2447 544 -2447 0 4
rlabel polysilicon 548 -2441 548 -2441 0 1
rlabel polysilicon 548 -2447 548 -2447 0 3
rlabel polysilicon 555 -2441 555 -2441 0 1
rlabel polysilicon 555 -2447 555 -2447 0 3
rlabel polysilicon 562 -2441 562 -2441 0 1
rlabel polysilicon 562 -2447 562 -2447 0 3
rlabel polysilicon 569 -2441 569 -2441 0 1
rlabel polysilicon 569 -2447 569 -2447 0 3
rlabel polysilicon 576 -2441 576 -2441 0 1
rlabel polysilicon 576 -2447 576 -2447 0 3
rlabel polysilicon 583 -2441 583 -2441 0 1
rlabel polysilicon 583 -2447 583 -2447 0 3
rlabel polysilicon 590 -2441 590 -2441 0 1
rlabel polysilicon 590 -2447 590 -2447 0 3
rlabel polysilicon 597 -2441 597 -2441 0 1
rlabel polysilicon 597 -2447 597 -2447 0 3
rlabel polysilicon 600 -2447 600 -2447 0 4
rlabel polysilicon 604 -2441 604 -2441 0 1
rlabel polysilicon 604 -2447 604 -2447 0 3
rlabel polysilicon 611 -2441 611 -2441 0 1
rlabel polysilicon 611 -2447 611 -2447 0 3
rlabel polysilicon 618 -2441 618 -2441 0 1
rlabel polysilicon 618 -2447 618 -2447 0 3
rlabel polysilicon 625 -2441 625 -2441 0 1
rlabel polysilicon 625 -2447 625 -2447 0 3
rlabel polysilicon 632 -2441 632 -2441 0 1
rlabel polysilicon 632 -2447 632 -2447 0 3
rlabel polysilicon 639 -2441 639 -2441 0 1
rlabel polysilicon 639 -2447 639 -2447 0 3
rlabel polysilicon 646 -2441 646 -2441 0 1
rlabel polysilicon 646 -2447 646 -2447 0 3
rlabel polysilicon 653 -2441 653 -2441 0 1
rlabel polysilicon 653 -2447 653 -2447 0 3
rlabel polysilicon 660 -2441 660 -2441 0 1
rlabel polysilicon 660 -2447 660 -2447 0 3
rlabel polysilicon 667 -2441 667 -2441 0 1
rlabel polysilicon 667 -2447 667 -2447 0 3
rlabel polysilicon 674 -2441 674 -2441 0 1
rlabel polysilicon 677 -2441 677 -2441 0 2
rlabel polysilicon 674 -2447 674 -2447 0 3
rlabel polysilicon 677 -2447 677 -2447 0 4
rlabel polysilicon 681 -2441 681 -2441 0 1
rlabel polysilicon 681 -2447 681 -2447 0 3
rlabel polysilicon 688 -2441 688 -2441 0 1
rlabel polysilicon 688 -2447 688 -2447 0 3
rlabel polysilicon 695 -2441 695 -2441 0 1
rlabel polysilicon 698 -2441 698 -2441 0 2
rlabel polysilicon 695 -2447 695 -2447 0 3
rlabel polysilicon 702 -2441 702 -2441 0 1
rlabel polysilicon 702 -2447 702 -2447 0 3
rlabel polysilicon 709 -2441 709 -2441 0 1
rlabel polysilicon 709 -2447 709 -2447 0 3
rlabel polysilicon 716 -2447 716 -2447 0 3
rlabel polysilicon 719 -2447 719 -2447 0 4
rlabel polysilicon 723 -2441 723 -2441 0 1
rlabel polysilicon 723 -2447 723 -2447 0 3
rlabel polysilicon 730 -2441 730 -2441 0 1
rlabel polysilicon 733 -2441 733 -2441 0 2
rlabel polysilicon 730 -2447 730 -2447 0 3
rlabel polysilicon 737 -2441 737 -2441 0 1
rlabel polysilicon 737 -2447 737 -2447 0 3
rlabel polysilicon 744 -2441 744 -2441 0 1
rlabel polysilicon 744 -2447 744 -2447 0 3
rlabel polysilicon 751 -2441 751 -2441 0 1
rlabel polysilicon 751 -2447 751 -2447 0 3
rlabel polysilicon 758 -2441 758 -2441 0 1
rlabel polysilicon 758 -2447 758 -2447 0 3
rlabel polysilicon 765 -2441 765 -2441 0 1
rlabel polysilicon 765 -2447 765 -2447 0 3
rlabel polysilicon 772 -2441 772 -2441 0 1
rlabel polysilicon 772 -2447 772 -2447 0 3
rlabel polysilicon 779 -2441 779 -2441 0 1
rlabel polysilicon 779 -2447 779 -2447 0 3
rlabel polysilicon 786 -2441 786 -2441 0 1
rlabel polysilicon 786 -2447 786 -2447 0 3
rlabel polysilicon 789 -2447 789 -2447 0 4
rlabel polysilicon 793 -2441 793 -2441 0 1
rlabel polysilicon 793 -2447 793 -2447 0 3
rlabel polysilicon 800 -2441 800 -2441 0 1
rlabel polysilicon 800 -2447 800 -2447 0 3
rlabel polysilicon 807 -2441 807 -2441 0 1
rlabel polysilicon 807 -2447 807 -2447 0 3
rlabel polysilicon 814 -2441 814 -2441 0 1
rlabel polysilicon 814 -2447 814 -2447 0 3
rlabel polysilicon 821 -2441 821 -2441 0 1
rlabel polysilicon 821 -2447 821 -2447 0 3
rlabel polysilicon 828 -2441 828 -2441 0 1
rlabel polysilicon 831 -2441 831 -2441 0 2
rlabel polysilicon 828 -2447 828 -2447 0 3
rlabel polysilicon 831 -2447 831 -2447 0 4
rlabel polysilicon 835 -2441 835 -2441 0 1
rlabel polysilicon 835 -2447 835 -2447 0 3
rlabel polysilicon 842 -2441 842 -2441 0 1
rlabel polysilicon 842 -2447 842 -2447 0 3
rlabel polysilicon 849 -2441 849 -2441 0 1
rlabel polysilicon 849 -2447 849 -2447 0 3
rlabel polysilicon 856 -2441 856 -2441 0 1
rlabel polysilicon 856 -2447 856 -2447 0 3
rlabel polysilicon 863 -2441 863 -2441 0 1
rlabel polysilicon 863 -2447 863 -2447 0 3
rlabel polysilicon 870 -2441 870 -2441 0 1
rlabel polysilicon 870 -2447 870 -2447 0 3
rlabel polysilicon 877 -2441 877 -2441 0 1
rlabel polysilicon 877 -2447 877 -2447 0 3
rlabel polysilicon 884 -2441 884 -2441 0 1
rlabel polysilicon 887 -2441 887 -2441 0 2
rlabel polysilicon 884 -2447 884 -2447 0 3
rlabel polysilicon 887 -2447 887 -2447 0 4
rlabel polysilicon 891 -2441 891 -2441 0 1
rlabel polysilicon 891 -2447 891 -2447 0 3
rlabel polysilicon 898 -2441 898 -2441 0 1
rlabel polysilicon 898 -2447 898 -2447 0 3
rlabel polysilicon 905 -2441 905 -2441 0 1
rlabel polysilicon 905 -2447 905 -2447 0 3
rlabel polysilicon 912 -2441 912 -2441 0 1
rlabel polysilicon 912 -2447 912 -2447 0 3
rlabel polysilicon 919 -2441 919 -2441 0 1
rlabel polysilicon 919 -2447 919 -2447 0 3
rlabel polysilicon 926 -2441 926 -2441 0 1
rlabel polysilicon 926 -2447 926 -2447 0 3
rlabel polysilicon 933 -2441 933 -2441 0 1
rlabel polysilicon 933 -2447 933 -2447 0 3
rlabel polysilicon 940 -2441 940 -2441 0 1
rlabel polysilicon 940 -2447 940 -2447 0 3
rlabel polysilicon 947 -2441 947 -2441 0 1
rlabel polysilicon 947 -2447 947 -2447 0 3
rlabel polysilicon 954 -2441 954 -2441 0 1
rlabel polysilicon 954 -2447 954 -2447 0 3
rlabel polysilicon 961 -2441 961 -2441 0 1
rlabel polysilicon 961 -2447 961 -2447 0 3
rlabel polysilicon 968 -2441 968 -2441 0 1
rlabel polysilicon 968 -2447 968 -2447 0 3
rlabel polysilicon 975 -2441 975 -2441 0 1
rlabel polysilicon 975 -2447 975 -2447 0 3
rlabel polysilicon 982 -2441 982 -2441 0 1
rlabel polysilicon 982 -2447 982 -2447 0 3
rlabel polysilicon 989 -2441 989 -2441 0 1
rlabel polysilicon 989 -2447 989 -2447 0 3
rlabel polysilicon 996 -2441 996 -2441 0 1
rlabel polysilicon 996 -2447 996 -2447 0 3
rlabel polysilicon 1003 -2441 1003 -2441 0 1
rlabel polysilicon 1003 -2447 1003 -2447 0 3
rlabel polysilicon 1010 -2441 1010 -2441 0 1
rlabel polysilicon 1010 -2447 1010 -2447 0 3
rlabel polysilicon 1017 -2441 1017 -2441 0 1
rlabel polysilicon 1020 -2441 1020 -2441 0 2
rlabel polysilicon 1017 -2447 1017 -2447 0 3
rlabel polysilicon 1020 -2447 1020 -2447 0 4
rlabel polysilicon 1024 -2441 1024 -2441 0 1
rlabel polysilicon 1024 -2447 1024 -2447 0 3
rlabel polysilicon 1031 -2441 1031 -2441 0 1
rlabel polysilicon 1031 -2447 1031 -2447 0 3
rlabel polysilicon 1038 -2441 1038 -2441 0 1
rlabel polysilicon 1038 -2447 1038 -2447 0 3
rlabel polysilicon 1045 -2441 1045 -2441 0 1
rlabel polysilicon 1045 -2447 1045 -2447 0 3
rlabel polysilicon 1052 -2441 1052 -2441 0 1
rlabel polysilicon 1055 -2441 1055 -2441 0 2
rlabel polysilicon 1059 -2441 1059 -2441 0 1
rlabel polysilicon 1059 -2447 1059 -2447 0 3
rlabel polysilicon 1066 -2441 1066 -2441 0 1
rlabel polysilicon 1066 -2447 1066 -2447 0 3
rlabel polysilicon 1073 -2441 1073 -2441 0 1
rlabel polysilicon 1073 -2447 1073 -2447 0 3
rlabel polysilicon 1080 -2441 1080 -2441 0 1
rlabel polysilicon 1083 -2441 1083 -2441 0 2
rlabel polysilicon 1080 -2447 1080 -2447 0 3
rlabel polysilicon 1087 -2441 1087 -2441 0 1
rlabel polysilicon 1087 -2447 1087 -2447 0 3
rlabel polysilicon 1094 -2441 1094 -2441 0 1
rlabel polysilicon 1094 -2447 1094 -2447 0 3
rlabel polysilicon 1101 -2441 1101 -2441 0 1
rlabel polysilicon 1101 -2447 1101 -2447 0 3
rlabel polysilicon 1108 -2441 1108 -2441 0 1
rlabel polysilicon 1108 -2447 1108 -2447 0 3
rlabel polysilicon 1115 -2441 1115 -2441 0 1
rlabel polysilicon 1115 -2447 1115 -2447 0 3
rlabel polysilicon 1122 -2441 1122 -2441 0 1
rlabel polysilicon 1122 -2447 1122 -2447 0 3
rlabel polysilicon 1129 -2441 1129 -2441 0 1
rlabel polysilicon 1129 -2447 1129 -2447 0 3
rlabel polysilicon 1136 -2441 1136 -2441 0 1
rlabel polysilicon 1136 -2447 1136 -2447 0 3
rlabel polysilicon 1143 -2441 1143 -2441 0 1
rlabel polysilicon 1143 -2447 1143 -2447 0 3
rlabel polysilicon 1150 -2441 1150 -2441 0 1
rlabel polysilicon 1150 -2447 1150 -2447 0 3
rlabel polysilicon 1157 -2441 1157 -2441 0 1
rlabel polysilicon 1157 -2447 1157 -2447 0 3
rlabel polysilicon 1164 -2441 1164 -2441 0 1
rlabel polysilicon 1167 -2441 1167 -2441 0 2
rlabel polysilicon 1164 -2447 1164 -2447 0 3
rlabel polysilicon 1167 -2447 1167 -2447 0 4
rlabel polysilicon 1171 -2441 1171 -2441 0 1
rlabel polysilicon 1171 -2447 1171 -2447 0 3
rlabel polysilicon 1178 -2441 1178 -2441 0 1
rlabel polysilicon 1178 -2447 1178 -2447 0 3
rlabel polysilicon 1185 -2441 1185 -2441 0 1
rlabel polysilicon 1185 -2447 1185 -2447 0 3
rlabel polysilicon 1192 -2441 1192 -2441 0 1
rlabel polysilicon 1192 -2447 1192 -2447 0 3
rlabel polysilicon 1199 -2441 1199 -2441 0 1
rlabel polysilicon 1199 -2447 1199 -2447 0 3
rlabel polysilicon 1206 -2441 1206 -2441 0 1
rlabel polysilicon 1206 -2447 1206 -2447 0 3
rlabel polysilicon 1213 -2441 1213 -2441 0 1
rlabel polysilicon 1216 -2441 1216 -2441 0 2
rlabel polysilicon 1213 -2447 1213 -2447 0 3
rlabel polysilicon 1220 -2441 1220 -2441 0 1
rlabel polysilicon 1220 -2447 1220 -2447 0 3
rlabel polysilicon 1227 -2441 1227 -2441 0 1
rlabel polysilicon 1227 -2447 1227 -2447 0 3
rlabel polysilicon 1234 -2441 1234 -2441 0 1
rlabel polysilicon 1234 -2447 1234 -2447 0 3
rlabel polysilicon 1241 -2441 1241 -2441 0 1
rlabel polysilicon 1241 -2447 1241 -2447 0 3
rlabel polysilicon 1248 -2441 1248 -2441 0 1
rlabel polysilicon 1248 -2447 1248 -2447 0 3
rlabel polysilicon 1255 -2441 1255 -2441 0 1
rlabel polysilicon 1255 -2447 1255 -2447 0 3
rlabel polysilicon 1262 -2441 1262 -2441 0 1
rlabel polysilicon 1262 -2447 1262 -2447 0 3
rlabel polysilicon 1269 -2441 1269 -2441 0 1
rlabel polysilicon 1269 -2447 1269 -2447 0 3
rlabel polysilicon 1276 -2441 1276 -2441 0 1
rlabel polysilicon 1276 -2447 1276 -2447 0 3
rlabel polysilicon 1283 -2441 1283 -2441 0 1
rlabel polysilicon 1283 -2447 1283 -2447 0 3
rlabel polysilicon 1290 -2441 1290 -2441 0 1
rlabel polysilicon 1290 -2447 1290 -2447 0 3
rlabel polysilicon 1297 -2441 1297 -2441 0 1
rlabel polysilicon 1297 -2447 1297 -2447 0 3
rlabel polysilicon 1304 -2441 1304 -2441 0 1
rlabel polysilicon 1304 -2447 1304 -2447 0 3
rlabel polysilicon 1311 -2441 1311 -2441 0 1
rlabel polysilicon 1311 -2447 1311 -2447 0 3
rlabel polysilicon 1321 -2441 1321 -2441 0 2
rlabel polysilicon 1318 -2447 1318 -2447 0 3
rlabel polysilicon 1321 -2447 1321 -2447 0 4
rlabel polysilicon 1325 -2441 1325 -2441 0 1
rlabel polysilicon 1325 -2447 1325 -2447 0 3
rlabel polysilicon 1332 -2441 1332 -2441 0 1
rlabel polysilicon 1332 -2447 1332 -2447 0 3
rlabel polysilicon 1339 -2441 1339 -2441 0 1
rlabel polysilicon 1342 -2441 1342 -2441 0 2
rlabel polysilicon 1346 -2441 1346 -2441 0 1
rlabel polysilicon 1346 -2447 1346 -2447 0 3
rlabel polysilicon 1353 -2441 1353 -2441 0 1
rlabel polysilicon 1353 -2447 1353 -2447 0 3
rlabel polysilicon 1360 -2441 1360 -2441 0 1
rlabel polysilicon 1360 -2447 1360 -2447 0 3
rlabel polysilicon 1367 -2441 1367 -2441 0 1
rlabel polysilicon 1367 -2447 1367 -2447 0 3
rlabel polysilicon 1374 -2441 1374 -2441 0 1
rlabel polysilicon 1374 -2447 1374 -2447 0 3
rlabel polysilicon 1381 -2441 1381 -2441 0 1
rlabel polysilicon 1381 -2447 1381 -2447 0 3
rlabel polysilicon 1388 -2441 1388 -2441 0 1
rlabel polysilicon 1391 -2441 1391 -2441 0 2
rlabel polysilicon 1388 -2447 1388 -2447 0 3
rlabel polysilicon 1395 -2441 1395 -2441 0 1
rlabel polysilicon 1395 -2447 1395 -2447 0 3
rlabel polysilicon 1402 -2441 1402 -2441 0 1
rlabel polysilicon 1402 -2447 1402 -2447 0 3
rlabel polysilicon 1409 -2441 1409 -2441 0 1
rlabel polysilicon 1409 -2447 1409 -2447 0 3
rlabel polysilicon 1416 -2441 1416 -2441 0 1
rlabel polysilicon 1416 -2447 1416 -2447 0 3
rlabel polysilicon 1423 -2441 1423 -2441 0 1
rlabel polysilicon 1423 -2447 1423 -2447 0 3
rlabel polysilicon 1430 -2441 1430 -2441 0 1
rlabel polysilicon 1430 -2447 1430 -2447 0 3
rlabel polysilicon 1437 -2441 1437 -2441 0 1
rlabel polysilicon 1437 -2447 1437 -2447 0 3
rlabel polysilicon 1444 -2441 1444 -2441 0 1
rlabel polysilicon 1444 -2447 1444 -2447 0 3
rlabel polysilicon 1451 -2441 1451 -2441 0 1
rlabel polysilicon 1451 -2447 1451 -2447 0 3
rlabel polysilicon 1458 -2441 1458 -2441 0 1
rlabel polysilicon 1458 -2447 1458 -2447 0 3
rlabel polysilicon 1465 -2441 1465 -2441 0 1
rlabel polysilicon 1465 -2447 1465 -2447 0 3
rlabel polysilicon 1472 -2441 1472 -2441 0 1
rlabel polysilicon 1472 -2447 1472 -2447 0 3
rlabel polysilicon 1479 -2441 1479 -2441 0 1
rlabel polysilicon 1479 -2447 1479 -2447 0 3
rlabel polysilicon 1486 -2441 1486 -2441 0 1
rlabel polysilicon 1486 -2447 1486 -2447 0 3
rlabel polysilicon 1493 -2441 1493 -2441 0 1
rlabel polysilicon 1493 -2447 1493 -2447 0 3
rlabel polysilicon 1500 -2441 1500 -2441 0 1
rlabel polysilicon 1500 -2447 1500 -2447 0 3
rlabel polysilicon 1507 -2441 1507 -2441 0 1
rlabel polysilicon 1507 -2447 1507 -2447 0 3
rlabel polysilicon 1514 -2441 1514 -2441 0 1
rlabel polysilicon 1514 -2447 1514 -2447 0 3
rlabel polysilicon 1521 -2441 1521 -2441 0 1
rlabel polysilicon 1521 -2447 1521 -2447 0 3
rlabel polysilicon 1528 -2441 1528 -2441 0 1
rlabel polysilicon 1528 -2447 1528 -2447 0 3
rlabel polysilicon 1535 -2441 1535 -2441 0 1
rlabel polysilicon 1535 -2447 1535 -2447 0 3
rlabel polysilicon 1542 -2441 1542 -2441 0 1
rlabel polysilicon 1542 -2447 1542 -2447 0 3
rlabel polysilicon 1549 -2441 1549 -2441 0 1
rlabel polysilicon 1549 -2447 1549 -2447 0 3
rlabel polysilicon 1556 -2441 1556 -2441 0 1
rlabel polysilicon 1556 -2447 1556 -2447 0 3
rlabel polysilicon 1563 -2441 1563 -2441 0 1
rlabel polysilicon 1563 -2447 1563 -2447 0 3
rlabel polysilicon 1570 -2441 1570 -2441 0 1
rlabel polysilicon 1570 -2447 1570 -2447 0 3
rlabel polysilicon 1577 -2441 1577 -2441 0 1
rlabel polysilicon 1577 -2447 1577 -2447 0 3
rlabel polysilicon 1584 -2441 1584 -2441 0 1
rlabel polysilicon 1584 -2447 1584 -2447 0 3
rlabel polysilicon 1591 -2441 1591 -2441 0 1
rlabel polysilicon 1591 -2447 1591 -2447 0 3
rlabel polysilicon 1598 -2441 1598 -2441 0 1
rlabel polysilicon 1598 -2447 1598 -2447 0 3
rlabel polysilicon 1605 -2441 1605 -2441 0 1
rlabel polysilicon 1605 -2447 1605 -2447 0 3
rlabel polysilicon 1612 -2441 1612 -2441 0 1
rlabel polysilicon 1612 -2447 1612 -2447 0 3
rlabel polysilicon 1619 -2441 1619 -2441 0 1
rlabel polysilicon 1619 -2447 1619 -2447 0 3
rlabel polysilicon 1626 -2441 1626 -2441 0 1
rlabel polysilicon 1626 -2447 1626 -2447 0 3
rlabel polysilicon 1633 -2441 1633 -2441 0 1
rlabel polysilicon 1633 -2447 1633 -2447 0 3
rlabel polysilicon 1640 -2441 1640 -2441 0 1
rlabel polysilicon 1640 -2447 1640 -2447 0 3
rlabel polysilicon 1647 -2441 1647 -2441 0 1
rlabel polysilicon 1647 -2447 1647 -2447 0 3
rlabel polysilicon 1654 -2441 1654 -2441 0 1
rlabel polysilicon 1654 -2447 1654 -2447 0 3
rlabel polysilicon 1661 -2441 1661 -2441 0 1
rlabel polysilicon 1661 -2447 1661 -2447 0 3
rlabel polysilicon 1668 -2441 1668 -2441 0 1
rlabel polysilicon 1668 -2447 1668 -2447 0 3
rlabel polysilicon 1675 -2441 1675 -2441 0 1
rlabel polysilicon 1675 -2447 1675 -2447 0 3
rlabel polysilicon 1682 -2441 1682 -2441 0 1
rlabel polysilicon 1682 -2447 1682 -2447 0 3
rlabel polysilicon 1689 -2441 1689 -2441 0 1
rlabel polysilicon 1689 -2447 1689 -2447 0 3
rlabel polysilicon 1696 -2441 1696 -2441 0 1
rlabel polysilicon 1696 -2447 1696 -2447 0 3
rlabel polysilicon 1703 -2441 1703 -2441 0 1
rlabel polysilicon 1703 -2447 1703 -2447 0 3
rlabel polysilicon 1710 -2441 1710 -2441 0 1
rlabel polysilicon 1710 -2447 1710 -2447 0 3
rlabel polysilicon 1717 -2441 1717 -2441 0 1
rlabel polysilicon 1717 -2447 1717 -2447 0 3
rlabel polysilicon 1724 -2441 1724 -2441 0 1
rlabel polysilicon 1724 -2447 1724 -2447 0 3
rlabel polysilicon 1731 -2441 1731 -2441 0 1
rlabel polysilicon 1731 -2447 1731 -2447 0 3
rlabel polysilicon 1738 -2441 1738 -2441 0 1
rlabel polysilicon 1738 -2447 1738 -2447 0 3
rlabel polysilicon 1745 -2441 1745 -2441 0 1
rlabel polysilicon 1745 -2447 1745 -2447 0 3
rlabel polysilicon 1752 -2441 1752 -2441 0 1
rlabel polysilicon 1755 -2441 1755 -2441 0 2
rlabel polysilicon 1759 -2441 1759 -2441 0 1
rlabel polysilicon 1759 -2447 1759 -2447 0 3
rlabel polysilicon 1766 -2441 1766 -2441 0 1
rlabel polysilicon 1766 -2447 1766 -2447 0 3
rlabel polysilicon 1773 -2441 1773 -2441 0 1
rlabel polysilicon 1773 -2447 1773 -2447 0 3
rlabel polysilicon 1780 -2441 1780 -2441 0 1
rlabel polysilicon 1780 -2447 1780 -2447 0 3
rlabel polysilicon 1787 -2441 1787 -2441 0 1
rlabel polysilicon 1787 -2447 1787 -2447 0 3
rlabel polysilicon 1794 -2441 1794 -2441 0 1
rlabel polysilicon 1797 -2441 1797 -2441 0 2
rlabel polysilicon 1794 -2447 1794 -2447 0 3
rlabel polysilicon 1801 -2441 1801 -2441 0 1
rlabel polysilicon 1801 -2447 1801 -2447 0 3
rlabel polysilicon 1808 -2441 1808 -2441 0 1
rlabel polysilicon 1808 -2447 1808 -2447 0 3
rlabel polysilicon 16 -2576 16 -2576 0 1
rlabel polysilicon 16 -2582 16 -2582 0 3
rlabel polysilicon 23 -2576 23 -2576 0 1
rlabel polysilicon 23 -2582 23 -2582 0 3
rlabel polysilicon 30 -2576 30 -2576 0 1
rlabel polysilicon 30 -2582 30 -2582 0 3
rlabel polysilicon 37 -2576 37 -2576 0 1
rlabel polysilicon 37 -2582 37 -2582 0 3
rlabel polysilicon 44 -2576 44 -2576 0 1
rlabel polysilicon 44 -2582 44 -2582 0 3
rlabel polysilicon 51 -2576 51 -2576 0 1
rlabel polysilicon 51 -2582 51 -2582 0 3
rlabel polysilicon 58 -2576 58 -2576 0 1
rlabel polysilicon 58 -2582 58 -2582 0 3
rlabel polysilicon 65 -2576 65 -2576 0 1
rlabel polysilicon 65 -2582 65 -2582 0 3
rlabel polysilicon 72 -2576 72 -2576 0 1
rlabel polysilicon 72 -2582 72 -2582 0 3
rlabel polysilicon 79 -2576 79 -2576 0 1
rlabel polysilicon 79 -2582 79 -2582 0 3
rlabel polysilicon 86 -2576 86 -2576 0 1
rlabel polysilicon 86 -2582 86 -2582 0 3
rlabel polysilicon 93 -2576 93 -2576 0 1
rlabel polysilicon 93 -2582 93 -2582 0 3
rlabel polysilicon 100 -2576 100 -2576 0 1
rlabel polysilicon 103 -2576 103 -2576 0 2
rlabel polysilicon 100 -2582 100 -2582 0 3
rlabel polysilicon 103 -2582 103 -2582 0 4
rlabel polysilicon 107 -2576 107 -2576 0 1
rlabel polysilicon 110 -2576 110 -2576 0 2
rlabel polysilicon 107 -2582 107 -2582 0 3
rlabel polysilicon 110 -2582 110 -2582 0 4
rlabel polysilicon 114 -2576 114 -2576 0 1
rlabel polysilicon 114 -2582 114 -2582 0 3
rlabel polysilicon 121 -2576 121 -2576 0 1
rlabel polysilicon 121 -2582 121 -2582 0 3
rlabel polysilicon 128 -2576 128 -2576 0 1
rlabel polysilicon 128 -2582 128 -2582 0 3
rlabel polysilicon 135 -2576 135 -2576 0 1
rlabel polysilicon 135 -2582 135 -2582 0 3
rlabel polysilicon 142 -2576 142 -2576 0 1
rlabel polysilicon 142 -2582 142 -2582 0 3
rlabel polysilicon 149 -2576 149 -2576 0 1
rlabel polysilicon 152 -2576 152 -2576 0 2
rlabel polysilicon 149 -2582 149 -2582 0 3
rlabel polysilicon 152 -2582 152 -2582 0 4
rlabel polysilicon 156 -2576 156 -2576 0 1
rlabel polysilicon 159 -2576 159 -2576 0 2
rlabel polysilicon 156 -2582 156 -2582 0 3
rlabel polysilicon 159 -2582 159 -2582 0 4
rlabel polysilicon 163 -2576 163 -2576 0 1
rlabel polysilicon 163 -2582 163 -2582 0 3
rlabel polysilicon 170 -2576 170 -2576 0 1
rlabel polysilicon 173 -2576 173 -2576 0 2
rlabel polysilicon 170 -2582 170 -2582 0 3
rlabel polysilicon 173 -2582 173 -2582 0 4
rlabel polysilicon 177 -2576 177 -2576 0 1
rlabel polysilicon 177 -2582 177 -2582 0 3
rlabel polysilicon 184 -2576 184 -2576 0 1
rlabel polysilicon 184 -2582 184 -2582 0 3
rlabel polysilicon 191 -2576 191 -2576 0 1
rlabel polysilicon 191 -2582 191 -2582 0 3
rlabel polysilicon 198 -2576 198 -2576 0 1
rlabel polysilicon 198 -2582 198 -2582 0 3
rlabel polysilicon 205 -2576 205 -2576 0 1
rlabel polysilicon 205 -2582 205 -2582 0 3
rlabel polysilicon 212 -2576 212 -2576 0 1
rlabel polysilicon 212 -2582 212 -2582 0 3
rlabel polysilicon 219 -2576 219 -2576 0 1
rlabel polysilicon 219 -2582 219 -2582 0 3
rlabel polysilicon 226 -2576 226 -2576 0 1
rlabel polysilicon 226 -2582 226 -2582 0 3
rlabel polysilicon 233 -2576 233 -2576 0 1
rlabel polysilicon 233 -2582 233 -2582 0 3
rlabel polysilicon 243 -2576 243 -2576 0 2
rlabel polysilicon 243 -2582 243 -2582 0 4
rlabel polysilicon 247 -2576 247 -2576 0 1
rlabel polysilicon 247 -2582 247 -2582 0 3
rlabel polysilicon 254 -2576 254 -2576 0 1
rlabel polysilicon 254 -2582 254 -2582 0 3
rlabel polysilicon 261 -2576 261 -2576 0 1
rlabel polysilicon 261 -2582 261 -2582 0 3
rlabel polysilicon 268 -2576 268 -2576 0 1
rlabel polysilicon 268 -2582 268 -2582 0 3
rlabel polysilicon 275 -2576 275 -2576 0 1
rlabel polysilicon 275 -2582 275 -2582 0 3
rlabel polysilicon 282 -2576 282 -2576 0 1
rlabel polysilicon 282 -2582 282 -2582 0 3
rlabel polysilicon 289 -2576 289 -2576 0 1
rlabel polysilicon 289 -2582 289 -2582 0 3
rlabel polysilicon 296 -2576 296 -2576 0 1
rlabel polysilicon 296 -2582 296 -2582 0 3
rlabel polysilicon 303 -2576 303 -2576 0 1
rlabel polysilicon 303 -2582 303 -2582 0 3
rlabel polysilicon 310 -2576 310 -2576 0 1
rlabel polysilicon 310 -2582 310 -2582 0 3
rlabel polysilicon 317 -2576 317 -2576 0 1
rlabel polysilicon 317 -2582 317 -2582 0 3
rlabel polysilicon 324 -2576 324 -2576 0 1
rlabel polysilicon 324 -2582 324 -2582 0 3
rlabel polysilicon 331 -2576 331 -2576 0 1
rlabel polysilicon 331 -2582 331 -2582 0 3
rlabel polysilicon 338 -2576 338 -2576 0 1
rlabel polysilicon 338 -2582 338 -2582 0 3
rlabel polysilicon 345 -2576 345 -2576 0 1
rlabel polysilicon 345 -2582 345 -2582 0 3
rlabel polysilicon 352 -2576 352 -2576 0 1
rlabel polysilicon 352 -2582 352 -2582 0 3
rlabel polysilicon 359 -2576 359 -2576 0 1
rlabel polysilicon 359 -2582 359 -2582 0 3
rlabel polysilicon 366 -2576 366 -2576 0 1
rlabel polysilicon 366 -2582 366 -2582 0 3
rlabel polysilicon 373 -2576 373 -2576 0 1
rlabel polysilicon 373 -2582 373 -2582 0 3
rlabel polysilicon 380 -2576 380 -2576 0 1
rlabel polysilicon 380 -2582 380 -2582 0 3
rlabel polysilicon 387 -2576 387 -2576 0 1
rlabel polysilicon 387 -2582 387 -2582 0 3
rlabel polysilicon 394 -2576 394 -2576 0 1
rlabel polysilicon 394 -2582 394 -2582 0 3
rlabel polysilicon 401 -2576 401 -2576 0 1
rlabel polysilicon 401 -2582 401 -2582 0 3
rlabel polysilicon 408 -2576 408 -2576 0 1
rlabel polysilicon 408 -2582 408 -2582 0 3
rlabel polysilicon 415 -2576 415 -2576 0 1
rlabel polysilicon 415 -2582 415 -2582 0 3
rlabel polysilicon 422 -2576 422 -2576 0 1
rlabel polysilicon 422 -2582 422 -2582 0 3
rlabel polysilicon 429 -2576 429 -2576 0 1
rlabel polysilicon 429 -2582 429 -2582 0 3
rlabel polysilicon 436 -2576 436 -2576 0 1
rlabel polysilicon 436 -2582 436 -2582 0 3
rlabel polysilicon 443 -2576 443 -2576 0 1
rlabel polysilicon 443 -2582 443 -2582 0 3
rlabel polysilicon 450 -2576 450 -2576 0 1
rlabel polysilicon 453 -2576 453 -2576 0 2
rlabel polysilicon 450 -2582 450 -2582 0 3
rlabel polysilicon 453 -2582 453 -2582 0 4
rlabel polysilicon 457 -2576 457 -2576 0 1
rlabel polysilicon 457 -2582 457 -2582 0 3
rlabel polysilicon 464 -2576 464 -2576 0 1
rlabel polysilicon 464 -2582 464 -2582 0 3
rlabel polysilicon 471 -2576 471 -2576 0 1
rlabel polysilicon 471 -2582 471 -2582 0 3
rlabel polysilicon 478 -2576 478 -2576 0 1
rlabel polysilicon 478 -2582 478 -2582 0 3
rlabel polysilicon 485 -2576 485 -2576 0 1
rlabel polysilicon 485 -2582 485 -2582 0 3
rlabel polysilicon 492 -2576 492 -2576 0 1
rlabel polysilicon 492 -2582 492 -2582 0 3
rlabel polysilicon 499 -2576 499 -2576 0 1
rlabel polysilicon 499 -2582 499 -2582 0 3
rlabel polysilicon 506 -2576 506 -2576 0 1
rlabel polysilicon 506 -2582 506 -2582 0 3
rlabel polysilicon 513 -2576 513 -2576 0 1
rlabel polysilicon 513 -2582 513 -2582 0 3
rlabel polysilicon 520 -2576 520 -2576 0 1
rlabel polysilicon 520 -2582 520 -2582 0 3
rlabel polysilicon 527 -2576 527 -2576 0 1
rlabel polysilicon 527 -2582 527 -2582 0 3
rlabel polysilicon 534 -2576 534 -2576 0 1
rlabel polysilicon 534 -2582 534 -2582 0 3
rlabel polysilicon 541 -2576 541 -2576 0 1
rlabel polysilicon 541 -2582 541 -2582 0 3
rlabel polysilicon 548 -2576 548 -2576 0 1
rlabel polysilicon 548 -2582 548 -2582 0 3
rlabel polysilicon 555 -2576 555 -2576 0 1
rlabel polysilicon 558 -2576 558 -2576 0 2
rlabel polysilicon 555 -2582 555 -2582 0 3
rlabel polysilicon 558 -2582 558 -2582 0 4
rlabel polysilicon 562 -2576 562 -2576 0 1
rlabel polysilicon 562 -2582 562 -2582 0 3
rlabel polysilicon 569 -2576 569 -2576 0 1
rlabel polysilicon 569 -2582 569 -2582 0 3
rlabel polysilicon 576 -2576 576 -2576 0 1
rlabel polysilicon 576 -2582 576 -2582 0 3
rlabel polysilicon 583 -2576 583 -2576 0 1
rlabel polysilicon 583 -2582 583 -2582 0 3
rlabel polysilicon 590 -2576 590 -2576 0 1
rlabel polysilicon 590 -2582 590 -2582 0 3
rlabel polysilicon 597 -2576 597 -2576 0 1
rlabel polysilicon 600 -2576 600 -2576 0 2
rlabel polysilicon 597 -2582 597 -2582 0 3
rlabel polysilicon 604 -2576 604 -2576 0 1
rlabel polysilicon 604 -2582 604 -2582 0 3
rlabel polysilicon 611 -2576 611 -2576 0 1
rlabel polysilicon 611 -2582 611 -2582 0 3
rlabel polysilicon 618 -2576 618 -2576 0 1
rlabel polysilicon 618 -2582 618 -2582 0 3
rlabel polysilicon 625 -2576 625 -2576 0 1
rlabel polysilicon 628 -2576 628 -2576 0 2
rlabel polysilicon 625 -2582 625 -2582 0 3
rlabel polysilicon 628 -2582 628 -2582 0 4
rlabel polysilicon 632 -2576 632 -2576 0 1
rlabel polysilicon 632 -2582 632 -2582 0 3
rlabel polysilicon 639 -2576 639 -2576 0 1
rlabel polysilicon 639 -2582 639 -2582 0 3
rlabel polysilicon 646 -2576 646 -2576 0 1
rlabel polysilicon 646 -2582 646 -2582 0 3
rlabel polysilicon 653 -2576 653 -2576 0 1
rlabel polysilicon 653 -2582 653 -2582 0 3
rlabel polysilicon 660 -2576 660 -2576 0 1
rlabel polysilicon 660 -2582 660 -2582 0 3
rlabel polysilicon 670 -2576 670 -2576 0 2
rlabel polysilicon 667 -2582 667 -2582 0 3
rlabel polysilicon 670 -2582 670 -2582 0 4
rlabel polysilicon 674 -2576 674 -2576 0 1
rlabel polysilicon 674 -2582 674 -2582 0 3
rlabel polysilicon 681 -2576 681 -2576 0 1
rlabel polysilicon 681 -2582 681 -2582 0 3
rlabel polysilicon 688 -2576 688 -2576 0 1
rlabel polysilicon 688 -2582 688 -2582 0 3
rlabel polysilicon 695 -2576 695 -2576 0 1
rlabel polysilicon 695 -2582 695 -2582 0 3
rlabel polysilicon 702 -2576 702 -2576 0 1
rlabel polysilicon 702 -2582 702 -2582 0 3
rlabel polysilicon 709 -2576 709 -2576 0 1
rlabel polysilicon 712 -2576 712 -2576 0 2
rlabel polysilicon 709 -2582 709 -2582 0 3
rlabel polysilicon 712 -2582 712 -2582 0 4
rlabel polysilicon 716 -2576 716 -2576 0 1
rlabel polysilicon 716 -2582 716 -2582 0 3
rlabel polysilicon 723 -2576 723 -2576 0 1
rlabel polysilicon 726 -2576 726 -2576 0 2
rlabel polysilicon 723 -2582 723 -2582 0 3
rlabel polysilicon 726 -2582 726 -2582 0 4
rlabel polysilicon 730 -2576 730 -2576 0 1
rlabel polysilicon 730 -2582 730 -2582 0 3
rlabel polysilicon 737 -2576 737 -2576 0 1
rlabel polysilicon 740 -2576 740 -2576 0 2
rlabel polysilicon 737 -2582 737 -2582 0 3
rlabel polysilicon 740 -2582 740 -2582 0 4
rlabel polysilicon 744 -2576 744 -2576 0 1
rlabel polysilicon 744 -2582 744 -2582 0 3
rlabel polysilicon 751 -2576 751 -2576 0 1
rlabel polysilicon 751 -2582 751 -2582 0 3
rlabel polysilicon 758 -2576 758 -2576 0 1
rlabel polysilicon 758 -2582 758 -2582 0 3
rlabel polysilicon 765 -2576 765 -2576 0 1
rlabel polysilicon 765 -2582 765 -2582 0 3
rlabel polysilicon 772 -2576 772 -2576 0 1
rlabel polysilicon 772 -2582 772 -2582 0 3
rlabel polysilicon 779 -2576 779 -2576 0 1
rlabel polysilicon 779 -2582 779 -2582 0 3
rlabel polysilicon 786 -2576 786 -2576 0 1
rlabel polysilicon 786 -2582 786 -2582 0 3
rlabel polysilicon 793 -2576 793 -2576 0 1
rlabel polysilicon 793 -2582 793 -2582 0 3
rlabel polysilicon 800 -2576 800 -2576 0 1
rlabel polysilicon 800 -2582 800 -2582 0 3
rlabel polysilicon 807 -2576 807 -2576 0 1
rlabel polysilicon 807 -2582 807 -2582 0 3
rlabel polysilicon 814 -2576 814 -2576 0 1
rlabel polysilicon 814 -2582 814 -2582 0 3
rlabel polysilicon 821 -2576 821 -2576 0 1
rlabel polysilicon 821 -2582 821 -2582 0 3
rlabel polysilicon 828 -2576 828 -2576 0 1
rlabel polysilicon 828 -2582 828 -2582 0 3
rlabel polysilicon 835 -2576 835 -2576 0 1
rlabel polysilicon 835 -2582 835 -2582 0 3
rlabel polysilicon 842 -2576 842 -2576 0 1
rlabel polysilicon 842 -2582 842 -2582 0 3
rlabel polysilicon 849 -2576 849 -2576 0 1
rlabel polysilicon 852 -2576 852 -2576 0 2
rlabel polysilicon 849 -2582 849 -2582 0 3
rlabel polysilicon 852 -2582 852 -2582 0 4
rlabel polysilicon 856 -2576 856 -2576 0 1
rlabel polysilicon 856 -2582 856 -2582 0 3
rlabel polysilicon 863 -2576 863 -2576 0 1
rlabel polysilicon 863 -2582 863 -2582 0 3
rlabel polysilicon 870 -2576 870 -2576 0 1
rlabel polysilicon 870 -2582 870 -2582 0 3
rlabel polysilicon 877 -2576 877 -2576 0 1
rlabel polysilicon 877 -2582 877 -2582 0 3
rlabel polysilicon 884 -2576 884 -2576 0 1
rlabel polysilicon 884 -2582 884 -2582 0 3
rlabel polysilicon 891 -2576 891 -2576 0 1
rlabel polysilicon 891 -2582 891 -2582 0 3
rlabel polysilicon 898 -2576 898 -2576 0 1
rlabel polysilicon 898 -2582 898 -2582 0 3
rlabel polysilicon 905 -2576 905 -2576 0 1
rlabel polysilicon 905 -2582 905 -2582 0 3
rlabel polysilicon 912 -2576 912 -2576 0 1
rlabel polysilicon 912 -2582 912 -2582 0 3
rlabel polysilicon 919 -2576 919 -2576 0 1
rlabel polysilicon 919 -2582 919 -2582 0 3
rlabel polysilicon 926 -2576 926 -2576 0 1
rlabel polysilicon 926 -2582 926 -2582 0 3
rlabel polysilicon 933 -2576 933 -2576 0 1
rlabel polysilicon 933 -2582 933 -2582 0 3
rlabel polysilicon 940 -2576 940 -2576 0 1
rlabel polysilicon 940 -2582 940 -2582 0 3
rlabel polysilicon 947 -2576 947 -2576 0 1
rlabel polysilicon 950 -2576 950 -2576 0 2
rlabel polysilicon 950 -2582 950 -2582 0 4
rlabel polysilicon 954 -2576 954 -2576 0 1
rlabel polysilicon 954 -2582 954 -2582 0 3
rlabel polysilicon 961 -2576 961 -2576 0 1
rlabel polysilicon 961 -2582 961 -2582 0 3
rlabel polysilicon 968 -2576 968 -2576 0 1
rlabel polysilicon 971 -2576 971 -2576 0 2
rlabel polysilicon 968 -2582 968 -2582 0 3
rlabel polysilicon 971 -2582 971 -2582 0 4
rlabel polysilicon 975 -2576 975 -2576 0 1
rlabel polysilicon 975 -2582 975 -2582 0 3
rlabel polysilicon 982 -2576 982 -2576 0 1
rlabel polysilicon 982 -2582 982 -2582 0 3
rlabel polysilicon 989 -2576 989 -2576 0 1
rlabel polysilicon 992 -2576 992 -2576 0 2
rlabel polysilicon 989 -2582 989 -2582 0 3
rlabel polysilicon 996 -2576 996 -2576 0 1
rlabel polysilicon 996 -2582 996 -2582 0 3
rlabel polysilicon 1003 -2576 1003 -2576 0 1
rlabel polysilicon 1003 -2582 1003 -2582 0 3
rlabel polysilicon 1010 -2576 1010 -2576 0 1
rlabel polysilicon 1010 -2582 1010 -2582 0 3
rlabel polysilicon 1017 -2576 1017 -2576 0 1
rlabel polysilicon 1020 -2576 1020 -2576 0 2
rlabel polysilicon 1017 -2582 1017 -2582 0 3
rlabel polysilicon 1020 -2582 1020 -2582 0 4
rlabel polysilicon 1024 -2576 1024 -2576 0 1
rlabel polysilicon 1024 -2582 1024 -2582 0 3
rlabel polysilicon 1031 -2576 1031 -2576 0 1
rlabel polysilicon 1031 -2582 1031 -2582 0 3
rlabel polysilicon 1038 -2576 1038 -2576 0 1
rlabel polysilicon 1038 -2582 1038 -2582 0 3
rlabel polysilicon 1045 -2576 1045 -2576 0 1
rlabel polysilicon 1048 -2576 1048 -2576 0 2
rlabel polysilicon 1045 -2582 1045 -2582 0 3
rlabel polysilicon 1048 -2582 1048 -2582 0 4
rlabel polysilicon 1052 -2576 1052 -2576 0 1
rlabel polysilicon 1055 -2576 1055 -2576 0 2
rlabel polysilicon 1052 -2582 1052 -2582 0 3
rlabel polysilicon 1055 -2582 1055 -2582 0 4
rlabel polysilicon 1059 -2576 1059 -2576 0 1
rlabel polysilicon 1059 -2582 1059 -2582 0 3
rlabel polysilicon 1066 -2576 1066 -2576 0 1
rlabel polysilicon 1066 -2582 1066 -2582 0 3
rlabel polysilicon 1076 -2576 1076 -2576 0 2
rlabel polysilicon 1076 -2582 1076 -2582 0 4
rlabel polysilicon 1080 -2576 1080 -2576 0 1
rlabel polysilicon 1080 -2582 1080 -2582 0 3
rlabel polysilicon 1087 -2576 1087 -2576 0 1
rlabel polysilicon 1087 -2582 1087 -2582 0 3
rlabel polysilicon 1094 -2576 1094 -2576 0 1
rlabel polysilicon 1094 -2582 1094 -2582 0 3
rlabel polysilicon 1101 -2576 1101 -2576 0 1
rlabel polysilicon 1101 -2582 1101 -2582 0 3
rlabel polysilicon 1108 -2576 1108 -2576 0 1
rlabel polysilicon 1108 -2582 1108 -2582 0 3
rlabel polysilicon 1115 -2576 1115 -2576 0 1
rlabel polysilicon 1118 -2576 1118 -2576 0 2
rlabel polysilicon 1118 -2582 1118 -2582 0 4
rlabel polysilicon 1122 -2576 1122 -2576 0 1
rlabel polysilicon 1122 -2582 1122 -2582 0 3
rlabel polysilicon 1129 -2576 1129 -2576 0 1
rlabel polysilicon 1132 -2576 1132 -2576 0 2
rlabel polysilicon 1129 -2582 1129 -2582 0 3
rlabel polysilicon 1132 -2582 1132 -2582 0 4
rlabel polysilicon 1136 -2582 1136 -2582 0 3
rlabel polysilicon 1139 -2582 1139 -2582 0 4
rlabel polysilicon 1143 -2576 1143 -2576 0 1
rlabel polysilicon 1143 -2582 1143 -2582 0 3
rlabel polysilicon 1150 -2576 1150 -2576 0 1
rlabel polysilicon 1150 -2582 1150 -2582 0 3
rlabel polysilicon 1157 -2576 1157 -2576 0 1
rlabel polysilicon 1160 -2576 1160 -2576 0 2
rlabel polysilicon 1160 -2582 1160 -2582 0 4
rlabel polysilicon 1164 -2576 1164 -2576 0 1
rlabel polysilicon 1164 -2582 1164 -2582 0 3
rlabel polysilicon 1171 -2576 1171 -2576 0 1
rlabel polysilicon 1174 -2576 1174 -2576 0 2
rlabel polysilicon 1171 -2582 1171 -2582 0 3
rlabel polysilicon 1174 -2582 1174 -2582 0 4
rlabel polysilicon 1178 -2576 1178 -2576 0 1
rlabel polysilicon 1178 -2582 1178 -2582 0 3
rlabel polysilicon 1185 -2576 1185 -2576 0 1
rlabel polysilicon 1185 -2582 1185 -2582 0 3
rlabel polysilicon 1192 -2576 1192 -2576 0 1
rlabel polysilicon 1195 -2576 1195 -2576 0 2
rlabel polysilicon 1192 -2582 1192 -2582 0 3
rlabel polysilicon 1195 -2582 1195 -2582 0 4
rlabel polysilicon 1199 -2576 1199 -2576 0 1
rlabel polysilicon 1199 -2582 1199 -2582 0 3
rlabel polysilicon 1206 -2576 1206 -2576 0 1
rlabel polysilicon 1206 -2582 1206 -2582 0 3
rlabel polysilicon 1213 -2576 1213 -2576 0 1
rlabel polysilicon 1213 -2582 1213 -2582 0 3
rlabel polysilicon 1220 -2576 1220 -2576 0 1
rlabel polysilicon 1220 -2582 1220 -2582 0 3
rlabel polysilicon 1227 -2576 1227 -2576 0 1
rlabel polysilicon 1227 -2582 1227 -2582 0 3
rlabel polysilicon 1234 -2576 1234 -2576 0 1
rlabel polysilicon 1234 -2582 1234 -2582 0 3
rlabel polysilicon 1241 -2576 1241 -2576 0 1
rlabel polysilicon 1241 -2582 1241 -2582 0 3
rlabel polysilicon 1248 -2576 1248 -2576 0 1
rlabel polysilicon 1248 -2582 1248 -2582 0 3
rlabel polysilicon 1255 -2576 1255 -2576 0 1
rlabel polysilicon 1255 -2582 1255 -2582 0 3
rlabel polysilicon 1262 -2576 1262 -2576 0 1
rlabel polysilicon 1262 -2582 1262 -2582 0 3
rlabel polysilicon 1269 -2576 1269 -2576 0 1
rlabel polysilicon 1269 -2582 1269 -2582 0 3
rlabel polysilicon 1276 -2576 1276 -2576 0 1
rlabel polysilicon 1276 -2582 1276 -2582 0 3
rlabel polysilicon 1283 -2576 1283 -2576 0 1
rlabel polysilicon 1283 -2582 1283 -2582 0 3
rlabel polysilicon 1290 -2576 1290 -2576 0 1
rlabel polysilicon 1290 -2582 1290 -2582 0 3
rlabel polysilicon 1297 -2576 1297 -2576 0 1
rlabel polysilicon 1297 -2582 1297 -2582 0 3
rlabel polysilicon 1304 -2576 1304 -2576 0 1
rlabel polysilicon 1304 -2582 1304 -2582 0 3
rlabel polysilicon 1311 -2576 1311 -2576 0 1
rlabel polysilicon 1311 -2582 1311 -2582 0 3
rlabel polysilicon 1318 -2576 1318 -2576 0 1
rlabel polysilicon 1318 -2582 1318 -2582 0 3
rlabel polysilicon 1325 -2576 1325 -2576 0 1
rlabel polysilicon 1325 -2582 1325 -2582 0 3
rlabel polysilicon 1332 -2576 1332 -2576 0 1
rlabel polysilicon 1332 -2582 1332 -2582 0 3
rlabel polysilicon 1339 -2576 1339 -2576 0 1
rlabel polysilicon 1339 -2582 1339 -2582 0 3
rlabel polysilicon 1346 -2576 1346 -2576 0 1
rlabel polysilicon 1346 -2582 1346 -2582 0 3
rlabel polysilicon 1353 -2576 1353 -2576 0 1
rlabel polysilicon 1353 -2582 1353 -2582 0 3
rlabel polysilicon 1360 -2576 1360 -2576 0 1
rlabel polysilicon 1360 -2582 1360 -2582 0 3
rlabel polysilicon 1367 -2576 1367 -2576 0 1
rlabel polysilicon 1367 -2582 1367 -2582 0 3
rlabel polysilicon 1374 -2576 1374 -2576 0 1
rlabel polysilicon 1374 -2582 1374 -2582 0 3
rlabel polysilicon 1381 -2576 1381 -2576 0 1
rlabel polysilicon 1381 -2582 1381 -2582 0 3
rlabel polysilicon 1388 -2576 1388 -2576 0 1
rlabel polysilicon 1388 -2582 1388 -2582 0 3
rlabel polysilicon 1395 -2576 1395 -2576 0 1
rlabel polysilicon 1395 -2582 1395 -2582 0 3
rlabel polysilicon 1402 -2576 1402 -2576 0 1
rlabel polysilicon 1402 -2582 1402 -2582 0 3
rlabel polysilicon 1409 -2576 1409 -2576 0 1
rlabel polysilicon 1409 -2582 1409 -2582 0 3
rlabel polysilicon 1416 -2576 1416 -2576 0 1
rlabel polysilicon 1416 -2582 1416 -2582 0 3
rlabel polysilicon 1423 -2576 1423 -2576 0 1
rlabel polysilicon 1423 -2582 1423 -2582 0 3
rlabel polysilicon 1430 -2576 1430 -2576 0 1
rlabel polysilicon 1430 -2582 1430 -2582 0 3
rlabel polysilicon 1437 -2576 1437 -2576 0 1
rlabel polysilicon 1437 -2582 1437 -2582 0 3
rlabel polysilicon 1444 -2576 1444 -2576 0 1
rlabel polysilicon 1444 -2582 1444 -2582 0 3
rlabel polysilicon 1451 -2576 1451 -2576 0 1
rlabel polysilicon 1451 -2582 1451 -2582 0 3
rlabel polysilicon 1458 -2576 1458 -2576 0 1
rlabel polysilicon 1458 -2582 1458 -2582 0 3
rlabel polysilicon 1465 -2576 1465 -2576 0 1
rlabel polysilicon 1465 -2582 1465 -2582 0 3
rlabel polysilicon 1472 -2576 1472 -2576 0 1
rlabel polysilicon 1472 -2582 1472 -2582 0 3
rlabel polysilicon 1479 -2576 1479 -2576 0 1
rlabel polysilicon 1479 -2582 1479 -2582 0 3
rlabel polysilicon 1486 -2576 1486 -2576 0 1
rlabel polysilicon 1486 -2582 1486 -2582 0 3
rlabel polysilicon 1493 -2576 1493 -2576 0 1
rlabel polysilicon 1493 -2582 1493 -2582 0 3
rlabel polysilicon 1500 -2576 1500 -2576 0 1
rlabel polysilicon 1500 -2582 1500 -2582 0 3
rlabel polysilicon 1507 -2582 1507 -2582 0 3
rlabel polysilicon 1510 -2582 1510 -2582 0 4
rlabel polysilicon 1514 -2576 1514 -2576 0 1
rlabel polysilicon 1514 -2582 1514 -2582 0 3
rlabel polysilicon 1521 -2576 1521 -2576 0 1
rlabel polysilicon 1521 -2582 1521 -2582 0 3
rlabel polysilicon 1528 -2576 1528 -2576 0 1
rlabel polysilicon 1528 -2582 1528 -2582 0 3
rlabel polysilicon 1535 -2576 1535 -2576 0 1
rlabel polysilicon 1535 -2582 1535 -2582 0 3
rlabel polysilicon 1542 -2576 1542 -2576 0 1
rlabel polysilicon 1542 -2582 1542 -2582 0 3
rlabel polysilicon 1549 -2576 1549 -2576 0 1
rlabel polysilicon 1549 -2582 1549 -2582 0 3
rlabel polysilicon 1556 -2576 1556 -2576 0 1
rlabel polysilicon 1556 -2582 1556 -2582 0 3
rlabel polysilicon 1563 -2576 1563 -2576 0 1
rlabel polysilicon 1563 -2582 1563 -2582 0 3
rlabel polysilicon 1570 -2576 1570 -2576 0 1
rlabel polysilicon 1570 -2582 1570 -2582 0 3
rlabel polysilicon 1577 -2576 1577 -2576 0 1
rlabel polysilicon 1577 -2582 1577 -2582 0 3
rlabel polysilicon 1584 -2576 1584 -2576 0 1
rlabel polysilicon 1584 -2582 1584 -2582 0 3
rlabel polysilicon 1591 -2576 1591 -2576 0 1
rlabel polysilicon 1591 -2582 1591 -2582 0 3
rlabel polysilicon 1598 -2576 1598 -2576 0 1
rlabel polysilicon 1598 -2582 1598 -2582 0 3
rlabel polysilicon 1605 -2576 1605 -2576 0 1
rlabel polysilicon 1605 -2582 1605 -2582 0 3
rlabel polysilicon 1612 -2576 1612 -2576 0 1
rlabel polysilicon 1612 -2582 1612 -2582 0 3
rlabel polysilicon 1619 -2576 1619 -2576 0 1
rlabel polysilicon 1619 -2582 1619 -2582 0 3
rlabel polysilicon 1626 -2576 1626 -2576 0 1
rlabel polysilicon 1626 -2582 1626 -2582 0 3
rlabel polysilicon 1633 -2576 1633 -2576 0 1
rlabel polysilicon 1633 -2582 1633 -2582 0 3
rlabel polysilicon 1640 -2576 1640 -2576 0 1
rlabel polysilicon 1640 -2582 1640 -2582 0 3
rlabel polysilicon 1647 -2576 1647 -2576 0 1
rlabel polysilicon 1647 -2582 1647 -2582 0 3
rlabel polysilicon 1654 -2576 1654 -2576 0 1
rlabel polysilicon 1654 -2582 1654 -2582 0 3
rlabel polysilicon 1661 -2576 1661 -2576 0 1
rlabel polysilicon 1661 -2582 1661 -2582 0 3
rlabel polysilicon 1668 -2576 1668 -2576 0 1
rlabel polysilicon 1668 -2582 1668 -2582 0 3
rlabel polysilicon 1675 -2576 1675 -2576 0 1
rlabel polysilicon 1675 -2582 1675 -2582 0 3
rlabel polysilicon 1682 -2576 1682 -2576 0 1
rlabel polysilicon 1682 -2582 1682 -2582 0 3
rlabel polysilicon 1689 -2576 1689 -2576 0 1
rlabel polysilicon 1689 -2582 1689 -2582 0 3
rlabel polysilicon 1696 -2576 1696 -2576 0 1
rlabel polysilicon 1699 -2576 1699 -2576 0 2
rlabel polysilicon 1696 -2582 1696 -2582 0 3
rlabel polysilicon 1699 -2582 1699 -2582 0 4
rlabel polysilicon 1703 -2576 1703 -2576 0 1
rlabel polysilicon 1703 -2582 1703 -2582 0 3
rlabel polysilicon 1710 -2576 1710 -2576 0 1
rlabel polysilicon 1710 -2582 1710 -2582 0 3
rlabel polysilicon 1717 -2576 1717 -2576 0 1
rlabel polysilicon 1717 -2582 1717 -2582 0 3
rlabel polysilicon 1724 -2576 1724 -2576 0 1
rlabel polysilicon 1724 -2582 1724 -2582 0 3
rlabel polysilicon 1731 -2576 1731 -2576 0 1
rlabel polysilicon 1731 -2582 1731 -2582 0 3
rlabel polysilicon 1738 -2576 1738 -2576 0 1
rlabel polysilicon 1741 -2576 1741 -2576 0 2
rlabel polysilicon 1738 -2582 1738 -2582 0 3
rlabel polysilicon 1741 -2582 1741 -2582 0 4
rlabel polysilicon 1745 -2576 1745 -2576 0 1
rlabel polysilicon 1745 -2582 1745 -2582 0 3
rlabel polysilicon 1752 -2576 1752 -2576 0 1
rlabel polysilicon 1752 -2582 1752 -2582 0 3
rlabel polysilicon 1759 -2576 1759 -2576 0 1
rlabel polysilicon 1759 -2582 1759 -2582 0 3
rlabel polysilicon 1766 -2576 1766 -2576 0 1
rlabel polysilicon 1766 -2582 1766 -2582 0 3
rlabel polysilicon 1773 -2576 1773 -2576 0 1
rlabel polysilicon 1773 -2582 1773 -2582 0 3
rlabel polysilicon 1780 -2576 1780 -2576 0 1
rlabel polysilicon 1780 -2582 1780 -2582 0 3
rlabel polysilicon 1787 -2576 1787 -2576 0 1
rlabel polysilicon 1787 -2582 1787 -2582 0 3
rlabel polysilicon 1794 -2582 1794 -2582 0 3
rlabel polysilicon 1801 -2576 1801 -2576 0 1
rlabel polysilicon 1801 -2582 1801 -2582 0 3
rlabel polysilicon 1808 -2576 1808 -2576 0 1
rlabel polysilicon 1808 -2582 1808 -2582 0 3
rlabel polysilicon 1815 -2576 1815 -2576 0 1
rlabel polysilicon 1815 -2582 1815 -2582 0 3
rlabel polysilicon 9 -2709 9 -2709 0 1
rlabel polysilicon 9 -2715 9 -2715 0 3
rlabel polysilicon 16 -2709 16 -2709 0 1
rlabel polysilicon 30 -2709 30 -2709 0 1
rlabel polysilicon 30 -2715 30 -2715 0 3
rlabel polysilicon 37 -2709 37 -2709 0 1
rlabel polysilicon 37 -2715 37 -2715 0 3
rlabel polysilicon 44 -2709 44 -2709 0 1
rlabel polysilicon 44 -2715 44 -2715 0 3
rlabel polysilicon 51 -2709 51 -2709 0 1
rlabel polysilicon 51 -2715 51 -2715 0 3
rlabel polysilicon 58 -2709 58 -2709 0 1
rlabel polysilicon 58 -2715 58 -2715 0 3
rlabel polysilicon 61 -2715 61 -2715 0 4
rlabel polysilicon 68 -2709 68 -2709 0 2
rlabel polysilicon 68 -2715 68 -2715 0 4
rlabel polysilicon 72 -2709 72 -2709 0 1
rlabel polysilicon 72 -2715 72 -2715 0 3
rlabel polysilicon 79 -2709 79 -2709 0 1
rlabel polysilicon 79 -2715 79 -2715 0 3
rlabel polysilicon 86 -2709 86 -2709 0 1
rlabel polysilicon 86 -2715 86 -2715 0 3
rlabel polysilicon 93 -2709 93 -2709 0 1
rlabel polysilicon 93 -2715 93 -2715 0 3
rlabel polysilicon 100 -2709 100 -2709 0 1
rlabel polysilicon 100 -2715 100 -2715 0 3
rlabel polysilicon 107 -2709 107 -2709 0 1
rlabel polysilicon 107 -2715 107 -2715 0 3
rlabel polysilicon 114 -2709 114 -2709 0 1
rlabel polysilicon 114 -2715 114 -2715 0 3
rlabel polysilicon 121 -2709 121 -2709 0 1
rlabel polysilicon 121 -2715 121 -2715 0 3
rlabel polysilicon 128 -2709 128 -2709 0 1
rlabel polysilicon 128 -2715 128 -2715 0 3
rlabel polysilicon 135 -2709 135 -2709 0 1
rlabel polysilicon 135 -2715 135 -2715 0 3
rlabel polysilicon 142 -2709 142 -2709 0 1
rlabel polysilicon 142 -2715 142 -2715 0 3
rlabel polysilicon 149 -2709 149 -2709 0 1
rlabel polysilicon 149 -2715 149 -2715 0 3
rlabel polysilicon 156 -2709 156 -2709 0 1
rlabel polysilicon 156 -2715 156 -2715 0 3
rlabel polysilicon 163 -2709 163 -2709 0 1
rlabel polysilicon 163 -2715 163 -2715 0 3
rlabel polysilicon 170 -2709 170 -2709 0 1
rlabel polysilicon 170 -2715 170 -2715 0 3
rlabel polysilicon 177 -2709 177 -2709 0 1
rlabel polysilicon 177 -2715 177 -2715 0 3
rlabel polysilicon 184 -2709 184 -2709 0 1
rlabel polysilicon 184 -2715 184 -2715 0 3
rlabel polysilicon 191 -2709 191 -2709 0 1
rlabel polysilicon 191 -2715 191 -2715 0 3
rlabel polysilicon 198 -2709 198 -2709 0 1
rlabel polysilicon 201 -2709 201 -2709 0 2
rlabel polysilicon 198 -2715 198 -2715 0 3
rlabel polysilicon 201 -2715 201 -2715 0 4
rlabel polysilicon 205 -2709 205 -2709 0 1
rlabel polysilicon 208 -2709 208 -2709 0 2
rlabel polysilicon 208 -2715 208 -2715 0 4
rlabel polysilicon 212 -2709 212 -2709 0 1
rlabel polysilicon 212 -2715 212 -2715 0 3
rlabel polysilicon 219 -2709 219 -2709 0 1
rlabel polysilicon 219 -2715 219 -2715 0 3
rlabel polysilicon 226 -2709 226 -2709 0 1
rlabel polysilicon 226 -2715 226 -2715 0 3
rlabel polysilicon 233 -2709 233 -2709 0 1
rlabel polysilicon 233 -2715 233 -2715 0 3
rlabel polysilicon 240 -2709 240 -2709 0 1
rlabel polysilicon 240 -2715 240 -2715 0 3
rlabel polysilicon 247 -2709 247 -2709 0 1
rlabel polysilicon 247 -2715 247 -2715 0 3
rlabel polysilicon 254 -2709 254 -2709 0 1
rlabel polysilicon 254 -2715 254 -2715 0 3
rlabel polysilicon 261 -2709 261 -2709 0 1
rlabel polysilicon 261 -2715 261 -2715 0 3
rlabel polysilicon 268 -2709 268 -2709 0 1
rlabel polysilicon 268 -2715 268 -2715 0 3
rlabel polysilicon 275 -2709 275 -2709 0 1
rlabel polysilicon 275 -2715 275 -2715 0 3
rlabel polysilicon 282 -2709 282 -2709 0 1
rlabel polysilicon 282 -2715 282 -2715 0 3
rlabel polysilicon 289 -2709 289 -2709 0 1
rlabel polysilicon 292 -2709 292 -2709 0 2
rlabel polysilicon 292 -2715 292 -2715 0 4
rlabel polysilicon 296 -2709 296 -2709 0 1
rlabel polysilicon 296 -2715 296 -2715 0 3
rlabel polysilicon 303 -2709 303 -2709 0 1
rlabel polysilicon 303 -2715 303 -2715 0 3
rlabel polysilicon 310 -2709 310 -2709 0 1
rlabel polysilicon 310 -2715 310 -2715 0 3
rlabel polysilicon 317 -2709 317 -2709 0 1
rlabel polysilicon 317 -2715 317 -2715 0 3
rlabel polysilicon 324 -2709 324 -2709 0 1
rlabel polysilicon 324 -2715 324 -2715 0 3
rlabel polysilicon 331 -2709 331 -2709 0 1
rlabel polysilicon 331 -2715 331 -2715 0 3
rlabel polysilicon 338 -2709 338 -2709 0 1
rlabel polysilicon 338 -2715 338 -2715 0 3
rlabel polysilicon 345 -2709 345 -2709 0 1
rlabel polysilicon 345 -2715 345 -2715 0 3
rlabel polysilicon 352 -2709 352 -2709 0 1
rlabel polysilicon 352 -2715 352 -2715 0 3
rlabel polysilicon 359 -2709 359 -2709 0 1
rlabel polysilicon 359 -2715 359 -2715 0 3
rlabel polysilicon 366 -2709 366 -2709 0 1
rlabel polysilicon 366 -2715 366 -2715 0 3
rlabel polysilicon 373 -2709 373 -2709 0 1
rlabel polysilicon 373 -2715 373 -2715 0 3
rlabel polysilicon 380 -2709 380 -2709 0 1
rlabel polysilicon 380 -2715 380 -2715 0 3
rlabel polysilicon 387 -2709 387 -2709 0 1
rlabel polysilicon 387 -2715 387 -2715 0 3
rlabel polysilicon 394 -2709 394 -2709 0 1
rlabel polysilicon 394 -2715 394 -2715 0 3
rlabel polysilicon 401 -2709 401 -2709 0 1
rlabel polysilicon 401 -2715 401 -2715 0 3
rlabel polysilicon 408 -2709 408 -2709 0 1
rlabel polysilicon 408 -2715 408 -2715 0 3
rlabel polysilicon 415 -2709 415 -2709 0 1
rlabel polysilicon 415 -2715 415 -2715 0 3
rlabel polysilicon 422 -2709 422 -2709 0 1
rlabel polysilicon 425 -2709 425 -2709 0 2
rlabel polysilicon 422 -2715 422 -2715 0 3
rlabel polysilicon 425 -2715 425 -2715 0 4
rlabel polysilicon 429 -2709 429 -2709 0 1
rlabel polysilicon 429 -2715 429 -2715 0 3
rlabel polysilicon 436 -2709 436 -2709 0 1
rlabel polysilicon 436 -2715 436 -2715 0 3
rlabel polysilicon 443 -2709 443 -2709 0 1
rlabel polysilicon 443 -2715 443 -2715 0 3
rlabel polysilicon 450 -2709 450 -2709 0 1
rlabel polysilicon 450 -2715 450 -2715 0 3
rlabel polysilicon 457 -2709 457 -2709 0 1
rlabel polysilicon 457 -2715 457 -2715 0 3
rlabel polysilicon 464 -2709 464 -2709 0 1
rlabel polysilicon 464 -2715 464 -2715 0 3
rlabel polysilicon 471 -2709 471 -2709 0 1
rlabel polysilicon 471 -2715 471 -2715 0 3
rlabel polysilicon 478 -2709 478 -2709 0 1
rlabel polysilicon 478 -2715 478 -2715 0 3
rlabel polysilicon 485 -2709 485 -2709 0 1
rlabel polysilicon 485 -2715 485 -2715 0 3
rlabel polysilicon 492 -2709 492 -2709 0 1
rlabel polysilicon 492 -2715 492 -2715 0 3
rlabel polysilicon 499 -2709 499 -2709 0 1
rlabel polysilicon 499 -2715 499 -2715 0 3
rlabel polysilicon 506 -2709 506 -2709 0 1
rlabel polysilicon 506 -2715 506 -2715 0 3
rlabel polysilicon 513 -2709 513 -2709 0 1
rlabel polysilicon 513 -2715 513 -2715 0 3
rlabel polysilicon 520 -2709 520 -2709 0 1
rlabel polysilicon 523 -2709 523 -2709 0 2
rlabel polysilicon 520 -2715 520 -2715 0 3
rlabel polysilicon 523 -2715 523 -2715 0 4
rlabel polysilicon 527 -2709 527 -2709 0 1
rlabel polysilicon 527 -2715 527 -2715 0 3
rlabel polysilicon 534 -2709 534 -2709 0 1
rlabel polysilicon 534 -2715 534 -2715 0 3
rlabel polysilicon 541 -2709 541 -2709 0 1
rlabel polysilicon 541 -2715 541 -2715 0 3
rlabel polysilicon 548 -2709 548 -2709 0 1
rlabel polysilicon 548 -2715 548 -2715 0 3
rlabel polysilicon 555 -2709 555 -2709 0 1
rlabel polysilicon 555 -2715 555 -2715 0 3
rlabel polysilicon 562 -2709 562 -2709 0 1
rlabel polysilicon 562 -2715 562 -2715 0 3
rlabel polysilicon 569 -2709 569 -2709 0 1
rlabel polysilicon 569 -2715 569 -2715 0 3
rlabel polysilicon 576 -2709 576 -2709 0 1
rlabel polysilicon 576 -2715 576 -2715 0 3
rlabel polysilicon 583 -2709 583 -2709 0 1
rlabel polysilicon 586 -2709 586 -2709 0 2
rlabel polysilicon 583 -2715 583 -2715 0 3
rlabel polysilicon 590 -2709 590 -2709 0 1
rlabel polysilicon 590 -2715 590 -2715 0 3
rlabel polysilicon 597 -2709 597 -2709 0 1
rlabel polysilicon 597 -2715 597 -2715 0 3
rlabel polysilicon 604 -2709 604 -2709 0 1
rlabel polysilicon 607 -2715 607 -2715 0 4
rlabel polysilicon 611 -2709 611 -2709 0 1
rlabel polysilicon 611 -2715 611 -2715 0 3
rlabel polysilicon 618 -2709 618 -2709 0 1
rlabel polysilicon 618 -2715 618 -2715 0 3
rlabel polysilicon 625 -2709 625 -2709 0 1
rlabel polysilicon 625 -2715 625 -2715 0 3
rlabel polysilicon 632 -2709 632 -2709 0 1
rlabel polysilicon 635 -2709 635 -2709 0 2
rlabel polysilicon 632 -2715 632 -2715 0 3
rlabel polysilicon 635 -2715 635 -2715 0 4
rlabel polysilicon 642 -2709 642 -2709 0 2
rlabel polysilicon 639 -2715 639 -2715 0 3
rlabel polysilicon 642 -2715 642 -2715 0 4
rlabel polysilicon 646 -2709 646 -2709 0 1
rlabel polysilicon 646 -2715 646 -2715 0 3
rlabel polysilicon 653 -2709 653 -2709 0 1
rlabel polysilicon 653 -2715 653 -2715 0 3
rlabel polysilicon 660 -2709 660 -2709 0 1
rlabel polysilicon 660 -2715 660 -2715 0 3
rlabel polysilicon 667 -2709 667 -2709 0 1
rlabel polysilicon 667 -2715 667 -2715 0 3
rlabel polysilicon 674 -2709 674 -2709 0 1
rlabel polysilicon 674 -2715 674 -2715 0 3
rlabel polysilicon 681 -2709 681 -2709 0 1
rlabel polysilicon 681 -2715 681 -2715 0 3
rlabel polysilicon 688 -2709 688 -2709 0 1
rlabel polysilicon 688 -2715 688 -2715 0 3
rlabel polysilicon 695 -2709 695 -2709 0 1
rlabel polysilicon 695 -2715 695 -2715 0 3
rlabel polysilicon 702 -2709 702 -2709 0 1
rlabel polysilicon 702 -2715 702 -2715 0 3
rlabel polysilicon 709 -2709 709 -2709 0 1
rlabel polysilicon 712 -2709 712 -2709 0 2
rlabel polysilicon 709 -2715 709 -2715 0 3
rlabel polysilicon 712 -2715 712 -2715 0 4
rlabel polysilicon 716 -2709 716 -2709 0 1
rlabel polysilicon 716 -2715 716 -2715 0 3
rlabel polysilicon 723 -2709 723 -2709 0 1
rlabel polysilicon 723 -2715 723 -2715 0 3
rlabel polysilicon 730 -2709 730 -2709 0 1
rlabel polysilicon 730 -2715 730 -2715 0 3
rlabel polysilicon 737 -2709 737 -2709 0 1
rlabel polysilicon 737 -2715 737 -2715 0 3
rlabel polysilicon 744 -2709 744 -2709 0 1
rlabel polysilicon 744 -2715 744 -2715 0 3
rlabel polysilicon 751 -2709 751 -2709 0 1
rlabel polysilicon 751 -2715 751 -2715 0 3
rlabel polysilicon 758 -2709 758 -2709 0 1
rlabel polysilicon 758 -2715 758 -2715 0 3
rlabel polysilicon 765 -2709 765 -2709 0 1
rlabel polysilicon 765 -2715 765 -2715 0 3
rlabel polysilicon 772 -2709 772 -2709 0 1
rlabel polysilicon 775 -2709 775 -2709 0 2
rlabel polysilicon 775 -2715 775 -2715 0 4
rlabel polysilicon 779 -2709 779 -2709 0 1
rlabel polysilicon 779 -2715 779 -2715 0 3
rlabel polysilicon 786 -2709 786 -2709 0 1
rlabel polysilicon 786 -2715 786 -2715 0 3
rlabel polysilicon 793 -2709 793 -2709 0 1
rlabel polysilicon 793 -2715 793 -2715 0 3
rlabel polysilicon 800 -2709 800 -2709 0 1
rlabel polysilicon 800 -2715 800 -2715 0 3
rlabel polysilicon 807 -2709 807 -2709 0 1
rlabel polysilicon 807 -2715 807 -2715 0 3
rlabel polysilicon 814 -2709 814 -2709 0 1
rlabel polysilicon 814 -2715 814 -2715 0 3
rlabel polysilicon 821 -2709 821 -2709 0 1
rlabel polysilicon 821 -2715 821 -2715 0 3
rlabel polysilicon 828 -2709 828 -2709 0 1
rlabel polysilicon 828 -2715 828 -2715 0 3
rlabel polysilicon 835 -2709 835 -2709 0 1
rlabel polysilicon 835 -2715 835 -2715 0 3
rlabel polysilicon 842 -2709 842 -2709 0 1
rlabel polysilicon 845 -2709 845 -2709 0 2
rlabel polysilicon 842 -2715 842 -2715 0 3
rlabel polysilicon 845 -2715 845 -2715 0 4
rlabel polysilicon 849 -2709 849 -2709 0 1
rlabel polysilicon 852 -2709 852 -2709 0 2
rlabel polysilicon 856 -2709 856 -2709 0 1
rlabel polysilicon 856 -2715 856 -2715 0 3
rlabel polysilicon 866 -2709 866 -2709 0 2
rlabel polysilicon 863 -2715 863 -2715 0 3
rlabel polysilicon 866 -2715 866 -2715 0 4
rlabel polysilicon 870 -2709 870 -2709 0 1
rlabel polysilicon 870 -2715 870 -2715 0 3
rlabel polysilicon 877 -2709 877 -2709 0 1
rlabel polysilicon 877 -2715 877 -2715 0 3
rlabel polysilicon 884 -2715 884 -2715 0 3
rlabel polysilicon 887 -2715 887 -2715 0 4
rlabel polysilicon 891 -2709 891 -2709 0 1
rlabel polysilicon 891 -2715 891 -2715 0 3
rlabel polysilicon 898 -2709 898 -2709 0 1
rlabel polysilicon 898 -2715 898 -2715 0 3
rlabel polysilicon 905 -2709 905 -2709 0 1
rlabel polysilicon 905 -2715 905 -2715 0 3
rlabel polysilicon 912 -2709 912 -2709 0 1
rlabel polysilicon 915 -2709 915 -2709 0 2
rlabel polysilicon 912 -2715 912 -2715 0 3
rlabel polysilicon 915 -2715 915 -2715 0 4
rlabel polysilicon 919 -2715 919 -2715 0 3
rlabel polysilicon 926 -2709 926 -2709 0 1
rlabel polysilicon 926 -2715 926 -2715 0 3
rlabel polysilicon 933 -2709 933 -2709 0 1
rlabel polysilicon 933 -2715 933 -2715 0 3
rlabel polysilicon 940 -2709 940 -2709 0 1
rlabel polysilicon 940 -2715 940 -2715 0 3
rlabel polysilicon 947 -2709 947 -2709 0 1
rlabel polysilicon 947 -2715 947 -2715 0 3
rlabel polysilicon 954 -2709 954 -2709 0 1
rlabel polysilicon 954 -2715 954 -2715 0 3
rlabel polysilicon 961 -2709 961 -2709 0 1
rlabel polysilicon 961 -2715 961 -2715 0 3
rlabel polysilicon 968 -2709 968 -2709 0 1
rlabel polysilicon 968 -2715 968 -2715 0 3
rlabel polysilicon 975 -2709 975 -2709 0 1
rlabel polysilicon 978 -2709 978 -2709 0 2
rlabel polysilicon 975 -2715 975 -2715 0 3
rlabel polysilicon 978 -2715 978 -2715 0 4
rlabel polysilicon 982 -2709 982 -2709 0 1
rlabel polysilicon 982 -2715 982 -2715 0 3
rlabel polysilicon 989 -2709 989 -2709 0 1
rlabel polysilicon 989 -2715 989 -2715 0 3
rlabel polysilicon 996 -2709 996 -2709 0 1
rlabel polysilicon 996 -2715 996 -2715 0 3
rlabel polysilicon 1003 -2709 1003 -2709 0 1
rlabel polysilicon 1003 -2715 1003 -2715 0 3
rlabel polysilicon 1010 -2709 1010 -2709 0 1
rlabel polysilicon 1010 -2715 1010 -2715 0 3
rlabel polysilicon 1017 -2709 1017 -2709 0 1
rlabel polysilicon 1020 -2709 1020 -2709 0 2
rlabel polysilicon 1020 -2715 1020 -2715 0 4
rlabel polysilicon 1024 -2709 1024 -2709 0 1
rlabel polysilicon 1024 -2715 1024 -2715 0 3
rlabel polysilicon 1031 -2709 1031 -2709 0 1
rlabel polysilicon 1031 -2715 1031 -2715 0 3
rlabel polysilicon 1038 -2709 1038 -2709 0 1
rlabel polysilicon 1038 -2715 1038 -2715 0 3
rlabel polysilicon 1045 -2709 1045 -2709 0 1
rlabel polysilicon 1045 -2715 1045 -2715 0 3
rlabel polysilicon 1052 -2709 1052 -2709 0 1
rlabel polysilicon 1055 -2709 1055 -2709 0 2
rlabel polysilicon 1052 -2715 1052 -2715 0 3
rlabel polysilicon 1059 -2709 1059 -2709 0 1
rlabel polysilicon 1062 -2709 1062 -2709 0 2
rlabel polysilicon 1059 -2715 1059 -2715 0 3
rlabel polysilicon 1062 -2715 1062 -2715 0 4
rlabel polysilicon 1066 -2709 1066 -2709 0 1
rlabel polysilicon 1066 -2715 1066 -2715 0 3
rlabel polysilicon 1073 -2709 1073 -2709 0 1
rlabel polysilicon 1073 -2715 1073 -2715 0 3
rlabel polysilicon 1080 -2709 1080 -2709 0 1
rlabel polysilicon 1080 -2715 1080 -2715 0 3
rlabel polysilicon 1087 -2709 1087 -2709 0 1
rlabel polysilicon 1087 -2715 1087 -2715 0 3
rlabel polysilicon 1094 -2709 1094 -2709 0 1
rlabel polysilicon 1094 -2715 1094 -2715 0 3
rlabel polysilicon 1101 -2709 1101 -2709 0 1
rlabel polysilicon 1101 -2715 1101 -2715 0 3
rlabel polysilicon 1108 -2709 1108 -2709 0 1
rlabel polysilicon 1108 -2715 1108 -2715 0 3
rlabel polysilicon 1115 -2709 1115 -2709 0 1
rlabel polysilicon 1115 -2715 1115 -2715 0 3
rlabel polysilicon 1122 -2709 1122 -2709 0 1
rlabel polysilicon 1122 -2715 1122 -2715 0 3
rlabel polysilicon 1129 -2709 1129 -2709 0 1
rlabel polysilicon 1129 -2715 1129 -2715 0 3
rlabel polysilicon 1136 -2709 1136 -2709 0 1
rlabel polysilicon 1136 -2715 1136 -2715 0 3
rlabel polysilicon 1143 -2709 1143 -2709 0 1
rlabel polysilicon 1143 -2715 1143 -2715 0 3
rlabel polysilicon 1150 -2709 1150 -2709 0 1
rlabel polysilicon 1150 -2715 1150 -2715 0 3
rlabel polysilicon 1153 -2715 1153 -2715 0 4
rlabel polysilicon 1157 -2709 1157 -2709 0 1
rlabel polysilicon 1157 -2715 1157 -2715 0 3
rlabel polysilicon 1164 -2709 1164 -2709 0 1
rlabel polysilicon 1164 -2715 1164 -2715 0 3
rlabel polysilicon 1171 -2709 1171 -2709 0 1
rlabel polysilicon 1171 -2715 1171 -2715 0 3
rlabel polysilicon 1178 -2709 1178 -2709 0 1
rlabel polysilicon 1178 -2715 1178 -2715 0 3
rlabel polysilicon 1185 -2709 1185 -2709 0 1
rlabel polysilicon 1185 -2715 1185 -2715 0 3
rlabel polysilicon 1192 -2709 1192 -2709 0 1
rlabel polysilicon 1195 -2709 1195 -2709 0 2
rlabel polysilicon 1192 -2715 1192 -2715 0 3
rlabel polysilicon 1195 -2715 1195 -2715 0 4
rlabel polysilicon 1199 -2709 1199 -2709 0 1
rlabel polysilicon 1199 -2715 1199 -2715 0 3
rlabel polysilicon 1206 -2709 1206 -2709 0 1
rlabel polysilicon 1206 -2715 1206 -2715 0 3
rlabel polysilicon 1213 -2709 1213 -2709 0 1
rlabel polysilicon 1213 -2715 1213 -2715 0 3
rlabel polysilicon 1220 -2709 1220 -2709 0 1
rlabel polysilicon 1220 -2715 1220 -2715 0 3
rlabel polysilicon 1227 -2709 1227 -2709 0 1
rlabel polysilicon 1227 -2715 1227 -2715 0 3
rlabel polysilicon 1234 -2709 1234 -2709 0 1
rlabel polysilicon 1234 -2715 1234 -2715 0 3
rlabel polysilicon 1241 -2709 1241 -2709 0 1
rlabel polysilicon 1244 -2709 1244 -2709 0 2
rlabel polysilicon 1241 -2715 1241 -2715 0 3
rlabel polysilicon 1244 -2715 1244 -2715 0 4
rlabel polysilicon 1248 -2709 1248 -2709 0 1
rlabel polysilicon 1248 -2715 1248 -2715 0 3
rlabel polysilicon 1255 -2709 1255 -2709 0 1
rlabel polysilicon 1255 -2715 1255 -2715 0 3
rlabel polysilicon 1262 -2709 1262 -2709 0 1
rlabel polysilicon 1262 -2715 1262 -2715 0 3
rlabel polysilicon 1269 -2709 1269 -2709 0 1
rlabel polysilicon 1269 -2715 1269 -2715 0 3
rlabel polysilicon 1276 -2709 1276 -2709 0 1
rlabel polysilicon 1276 -2715 1276 -2715 0 3
rlabel polysilicon 1283 -2709 1283 -2709 0 1
rlabel polysilicon 1283 -2715 1283 -2715 0 3
rlabel polysilicon 1293 -2709 1293 -2709 0 2
rlabel polysilicon 1297 -2709 1297 -2709 0 1
rlabel polysilicon 1297 -2715 1297 -2715 0 3
rlabel polysilicon 1304 -2709 1304 -2709 0 1
rlabel polysilicon 1304 -2715 1304 -2715 0 3
rlabel polysilicon 1311 -2709 1311 -2709 0 1
rlabel polysilicon 1311 -2715 1311 -2715 0 3
rlabel polysilicon 1318 -2709 1318 -2709 0 1
rlabel polysilicon 1321 -2709 1321 -2709 0 2
rlabel polysilicon 1318 -2715 1318 -2715 0 3
rlabel polysilicon 1321 -2715 1321 -2715 0 4
rlabel polysilicon 1325 -2709 1325 -2709 0 1
rlabel polysilicon 1325 -2715 1325 -2715 0 3
rlabel polysilicon 1328 -2715 1328 -2715 0 4
rlabel polysilicon 1332 -2709 1332 -2709 0 1
rlabel polysilicon 1332 -2715 1332 -2715 0 3
rlabel polysilicon 1339 -2709 1339 -2709 0 1
rlabel polysilicon 1339 -2715 1339 -2715 0 3
rlabel polysilicon 1346 -2709 1346 -2709 0 1
rlabel polysilicon 1346 -2715 1346 -2715 0 3
rlabel polysilicon 1353 -2709 1353 -2709 0 1
rlabel polysilicon 1353 -2715 1353 -2715 0 3
rlabel polysilicon 1360 -2709 1360 -2709 0 1
rlabel polysilicon 1360 -2715 1360 -2715 0 3
rlabel polysilicon 1367 -2709 1367 -2709 0 1
rlabel polysilicon 1367 -2715 1367 -2715 0 3
rlabel polysilicon 1374 -2709 1374 -2709 0 1
rlabel polysilicon 1374 -2715 1374 -2715 0 3
rlabel polysilicon 1381 -2709 1381 -2709 0 1
rlabel polysilicon 1381 -2715 1381 -2715 0 3
rlabel polysilicon 1388 -2709 1388 -2709 0 1
rlabel polysilicon 1388 -2715 1388 -2715 0 3
rlabel polysilicon 1395 -2709 1395 -2709 0 1
rlabel polysilicon 1395 -2715 1395 -2715 0 3
rlabel polysilicon 1402 -2709 1402 -2709 0 1
rlabel polysilicon 1402 -2715 1402 -2715 0 3
rlabel polysilicon 1409 -2709 1409 -2709 0 1
rlabel polysilicon 1409 -2715 1409 -2715 0 3
rlabel polysilicon 1416 -2709 1416 -2709 0 1
rlabel polysilicon 1416 -2715 1416 -2715 0 3
rlabel polysilicon 1423 -2709 1423 -2709 0 1
rlabel polysilicon 1423 -2715 1423 -2715 0 3
rlabel polysilicon 1430 -2709 1430 -2709 0 1
rlabel polysilicon 1430 -2715 1430 -2715 0 3
rlabel polysilicon 1437 -2709 1437 -2709 0 1
rlabel polysilicon 1437 -2715 1437 -2715 0 3
rlabel polysilicon 1444 -2709 1444 -2709 0 1
rlabel polysilicon 1444 -2715 1444 -2715 0 3
rlabel polysilicon 1451 -2709 1451 -2709 0 1
rlabel polysilicon 1451 -2715 1451 -2715 0 3
rlabel polysilicon 1458 -2709 1458 -2709 0 1
rlabel polysilicon 1458 -2715 1458 -2715 0 3
rlabel polysilicon 1465 -2709 1465 -2709 0 1
rlabel polysilicon 1465 -2715 1465 -2715 0 3
rlabel polysilicon 1472 -2709 1472 -2709 0 1
rlabel polysilicon 1472 -2715 1472 -2715 0 3
rlabel polysilicon 1479 -2709 1479 -2709 0 1
rlabel polysilicon 1479 -2715 1479 -2715 0 3
rlabel polysilicon 1486 -2709 1486 -2709 0 1
rlabel polysilicon 1486 -2715 1486 -2715 0 3
rlabel polysilicon 1493 -2709 1493 -2709 0 1
rlabel polysilicon 1493 -2715 1493 -2715 0 3
rlabel polysilicon 1500 -2709 1500 -2709 0 1
rlabel polysilicon 1500 -2715 1500 -2715 0 3
rlabel polysilicon 1507 -2709 1507 -2709 0 1
rlabel polysilicon 1507 -2715 1507 -2715 0 3
rlabel polysilicon 1514 -2709 1514 -2709 0 1
rlabel polysilicon 1514 -2715 1514 -2715 0 3
rlabel polysilicon 1521 -2709 1521 -2709 0 1
rlabel polysilicon 1521 -2715 1521 -2715 0 3
rlabel polysilicon 1528 -2709 1528 -2709 0 1
rlabel polysilicon 1528 -2715 1528 -2715 0 3
rlabel polysilicon 1535 -2709 1535 -2709 0 1
rlabel polysilicon 1535 -2715 1535 -2715 0 3
rlabel polysilicon 1542 -2709 1542 -2709 0 1
rlabel polysilicon 1542 -2715 1542 -2715 0 3
rlabel polysilicon 1549 -2709 1549 -2709 0 1
rlabel polysilicon 1549 -2715 1549 -2715 0 3
rlabel polysilicon 1556 -2709 1556 -2709 0 1
rlabel polysilicon 1556 -2715 1556 -2715 0 3
rlabel polysilicon 1563 -2709 1563 -2709 0 1
rlabel polysilicon 1563 -2715 1563 -2715 0 3
rlabel polysilicon 1570 -2709 1570 -2709 0 1
rlabel polysilicon 1570 -2715 1570 -2715 0 3
rlabel polysilicon 1577 -2709 1577 -2709 0 1
rlabel polysilicon 1577 -2715 1577 -2715 0 3
rlabel polysilicon 1584 -2709 1584 -2709 0 1
rlabel polysilicon 1584 -2715 1584 -2715 0 3
rlabel polysilicon 1591 -2709 1591 -2709 0 1
rlabel polysilicon 1591 -2715 1591 -2715 0 3
rlabel polysilicon 1598 -2709 1598 -2709 0 1
rlabel polysilicon 1598 -2715 1598 -2715 0 3
rlabel polysilicon 1605 -2709 1605 -2709 0 1
rlabel polysilicon 1605 -2715 1605 -2715 0 3
rlabel polysilicon 1612 -2709 1612 -2709 0 1
rlabel polysilicon 1612 -2715 1612 -2715 0 3
rlabel polysilicon 1619 -2709 1619 -2709 0 1
rlabel polysilicon 1619 -2715 1619 -2715 0 3
rlabel polysilicon 1626 -2709 1626 -2709 0 1
rlabel polysilicon 1626 -2715 1626 -2715 0 3
rlabel polysilicon 1633 -2709 1633 -2709 0 1
rlabel polysilicon 1633 -2715 1633 -2715 0 3
rlabel polysilicon 1640 -2709 1640 -2709 0 1
rlabel polysilicon 1640 -2715 1640 -2715 0 3
rlabel polysilicon 1647 -2709 1647 -2709 0 1
rlabel polysilicon 1647 -2715 1647 -2715 0 3
rlabel polysilicon 1654 -2709 1654 -2709 0 1
rlabel polysilicon 1654 -2715 1654 -2715 0 3
rlabel polysilicon 1661 -2709 1661 -2709 0 1
rlabel polysilicon 1661 -2715 1661 -2715 0 3
rlabel polysilicon 1668 -2709 1668 -2709 0 1
rlabel polysilicon 1668 -2715 1668 -2715 0 3
rlabel polysilicon 1675 -2709 1675 -2709 0 1
rlabel polysilicon 1675 -2715 1675 -2715 0 3
rlabel polysilicon 1682 -2709 1682 -2709 0 1
rlabel polysilicon 1682 -2715 1682 -2715 0 3
rlabel polysilicon 1689 -2709 1689 -2709 0 1
rlabel polysilicon 1689 -2715 1689 -2715 0 3
rlabel polysilicon 1696 -2709 1696 -2709 0 1
rlabel polysilicon 1696 -2715 1696 -2715 0 3
rlabel polysilicon 1703 -2709 1703 -2709 0 1
rlabel polysilicon 1703 -2715 1703 -2715 0 3
rlabel polysilicon 1710 -2709 1710 -2709 0 1
rlabel polysilicon 1710 -2715 1710 -2715 0 3
rlabel polysilicon 1717 -2709 1717 -2709 0 1
rlabel polysilicon 1717 -2715 1717 -2715 0 3
rlabel polysilicon 1724 -2709 1724 -2709 0 1
rlabel polysilicon 1724 -2715 1724 -2715 0 3
rlabel polysilicon 1731 -2709 1731 -2709 0 1
rlabel polysilicon 1731 -2715 1731 -2715 0 3
rlabel polysilicon 1738 -2709 1738 -2709 0 1
rlabel polysilicon 1738 -2715 1738 -2715 0 3
rlabel polysilicon 1745 -2709 1745 -2709 0 1
rlabel polysilicon 1745 -2715 1745 -2715 0 3
rlabel polysilicon 1752 -2709 1752 -2709 0 1
rlabel polysilicon 1752 -2715 1752 -2715 0 3
rlabel polysilicon 1759 -2709 1759 -2709 0 1
rlabel polysilicon 1759 -2715 1759 -2715 0 3
rlabel polysilicon 1766 -2709 1766 -2709 0 1
rlabel polysilicon 1769 -2709 1769 -2709 0 2
rlabel polysilicon 1766 -2715 1766 -2715 0 3
rlabel polysilicon 1769 -2715 1769 -2715 0 4
rlabel polysilicon 1773 -2709 1773 -2709 0 1
rlabel polysilicon 1776 -2709 1776 -2709 0 2
rlabel polysilicon 1773 -2715 1773 -2715 0 3
rlabel polysilicon 1776 -2715 1776 -2715 0 4
rlabel polysilicon 1783 -2709 1783 -2709 0 2
rlabel polysilicon 1780 -2715 1780 -2715 0 3
rlabel polysilicon 1783 -2715 1783 -2715 0 4
rlabel polysilicon 1787 -2709 1787 -2709 0 1
rlabel polysilicon 1787 -2715 1787 -2715 0 3
rlabel polysilicon 1794 -2709 1794 -2709 0 1
rlabel polysilicon 1794 -2715 1794 -2715 0 3
rlabel polysilicon 1801 -2709 1801 -2709 0 1
rlabel polysilicon 1801 -2715 1801 -2715 0 3
rlabel polysilicon 1808 -2709 1808 -2709 0 1
rlabel polysilicon 1808 -2715 1808 -2715 0 3
rlabel polysilicon 37 -2830 37 -2830 0 1
rlabel polysilicon 37 -2836 37 -2836 0 3
rlabel polysilicon 44 -2830 44 -2830 0 1
rlabel polysilicon 44 -2836 44 -2836 0 3
rlabel polysilicon 51 -2830 51 -2830 0 1
rlabel polysilicon 51 -2836 51 -2836 0 3
rlabel polysilicon 58 -2830 58 -2830 0 1
rlabel polysilicon 58 -2836 58 -2836 0 3
rlabel polysilicon 65 -2830 65 -2830 0 1
rlabel polysilicon 65 -2836 65 -2836 0 3
rlabel polysilicon 72 -2830 72 -2830 0 1
rlabel polysilicon 72 -2836 72 -2836 0 3
rlabel polysilicon 79 -2830 79 -2830 0 1
rlabel polysilicon 79 -2836 79 -2836 0 3
rlabel polysilicon 86 -2830 86 -2830 0 1
rlabel polysilicon 86 -2836 86 -2836 0 3
rlabel polysilicon 93 -2830 93 -2830 0 1
rlabel polysilicon 96 -2830 96 -2830 0 2
rlabel polysilicon 93 -2836 93 -2836 0 3
rlabel polysilicon 96 -2836 96 -2836 0 4
rlabel polysilicon 100 -2830 100 -2830 0 1
rlabel polysilicon 100 -2836 100 -2836 0 3
rlabel polysilicon 107 -2830 107 -2830 0 1
rlabel polysilicon 107 -2836 107 -2836 0 3
rlabel polysilicon 114 -2830 114 -2830 0 1
rlabel polysilicon 114 -2836 114 -2836 0 3
rlabel polysilicon 121 -2830 121 -2830 0 1
rlabel polysilicon 121 -2836 121 -2836 0 3
rlabel polysilicon 128 -2830 128 -2830 0 1
rlabel polysilicon 128 -2836 128 -2836 0 3
rlabel polysilicon 135 -2830 135 -2830 0 1
rlabel polysilicon 135 -2836 135 -2836 0 3
rlabel polysilicon 142 -2830 142 -2830 0 1
rlabel polysilicon 142 -2836 142 -2836 0 3
rlabel polysilicon 149 -2830 149 -2830 0 1
rlabel polysilicon 149 -2836 149 -2836 0 3
rlabel polysilicon 156 -2830 156 -2830 0 1
rlabel polysilicon 156 -2836 156 -2836 0 3
rlabel polysilicon 163 -2830 163 -2830 0 1
rlabel polysilicon 163 -2836 163 -2836 0 3
rlabel polysilicon 170 -2830 170 -2830 0 1
rlabel polysilicon 170 -2836 170 -2836 0 3
rlabel polysilicon 177 -2830 177 -2830 0 1
rlabel polysilicon 177 -2836 177 -2836 0 3
rlabel polysilicon 184 -2830 184 -2830 0 1
rlabel polysilicon 184 -2836 184 -2836 0 3
rlabel polysilicon 191 -2830 191 -2830 0 1
rlabel polysilicon 191 -2836 191 -2836 0 3
rlabel polysilicon 198 -2830 198 -2830 0 1
rlabel polysilicon 198 -2836 198 -2836 0 3
rlabel polysilicon 205 -2830 205 -2830 0 1
rlabel polysilicon 205 -2836 205 -2836 0 3
rlabel polysilicon 212 -2830 212 -2830 0 1
rlabel polysilicon 212 -2836 212 -2836 0 3
rlabel polysilicon 219 -2830 219 -2830 0 1
rlabel polysilicon 219 -2836 219 -2836 0 3
rlabel polysilicon 226 -2830 226 -2830 0 1
rlabel polysilicon 226 -2836 226 -2836 0 3
rlabel polysilicon 233 -2830 233 -2830 0 1
rlabel polysilicon 233 -2836 233 -2836 0 3
rlabel polysilicon 240 -2830 240 -2830 0 1
rlabel polysilicon 240 -2836 240 -2836 0 3
rlabel polysilicon 247 -2830 247 -2830 0 1
rlabel polysilicon 247 -2836 247 -2836 0 3
rlabel polysilicon 254 -2830 254 -2830 0 1
rlabel polysilicon 254 -2836 254 -2836 0 3
rlabel polysilicon 261 -2830 261 -2830 0 1
rlabel polysilicon 261 -2836 261 -2836 0 3
rlabel polysilicon 268 -2830 268 -2830 0 1
rlabel polysilicon 268 -2836 268 -2836 0 3
rlabel polysilicon 275 -2830 275 -2830 0 1
rlabel polysilicon 275 -2836 275 -2836 0 3
rlabel polysilicon 282 -2830 282 -2830 0 1
rlabel polysilicon 282 -2836 282 -2836 0 3
rlabel polysilicon 289 -2830 289 -2830 0 1
rlabel polysilicon 289 -2836 289 -2836 0 3
rlabel polysilicon 296 -2830 296 -2830 0 1
rlabel polysilicon 296 -2836 296 -2836 0 3
rlabel polysilicon 303 -2830 303 -2830 0 1
rlabel polysilicon 303 -2836 303 -2836 0 3
rlabel polysilicon 310 -2830 310 -2830 0 1
rlabel polysilicon 310 -2836 310 -2836 0 3
rlabel polysilicon 317 -2830 317 -2830 0 1
rlabel polysilicon 317 -2836 317 -2836 0 3
rlabel polysilicon 324 -2830 324 -2830 0 1
rlabel polysilicon 324 -2836 324 -2836 0 3
rlabel polysilicon 331 -2830 331 -2830 0 1
rlabel polysilicon 331 -2836 331 -2836 0 3
rlabel polysilicon 338 -2830 338 -2830 0 1
rlabel polysilicon 338 -2836 338 -2836 0 3
rlabel polysilicon 345 -2830 345 -2830 0 1
rlabel polysilicon 345 -2836 345 -2836 0 3
rlabel polysilicon 355 -2830 355 -2830 0 2
rlabel polysilicon 355 -2836 355 -2836 0 4
rlabel polysilicon 359 -2830 359 -2830 0 1
rlabel polysilicon 359 -2836 359 -2836 0 3
rlabel polysilicon 366 -2830 366 -2830 0 1
rlabel polysilicon 366 -2836 366 -2836 0 3
rlabel polysilicon 373 -2830 373 -2830 0 1
rlabel polysilicon 373 -2836 373 -2836 0 3
rlabel polysilicon 380 -2830 380 -2830 0 1
rlabel polysilicon 380 -2836 380 -2836 0 3
rlabel polysilicon 387 -2830 387 -2830 0 1
rlabel polysilicon 387 -2836 387 -2836 0 3
rlabel polysilicon 394 -2830 394 -2830 0 1
rlabel polysilicon 394 -2836 394 -2836 0 3
rlabel polysilicon 401 -2830 401 -2830 0 1
rlabel polysilicon 401 -2836 401 -2836 0 3
rlabel polysilicon 408 -2830 408 -2830 0 1
rlabel polysilicon 408 -2836 408 -2836 0 3
rlabel polysilicon 415 -2830 415 -2830 0 1
rlabel polysilicon 415 -2836 415 -2836 0 3
rlabel polysilicon 422 -2830 422 -2830 0 1
rlabel polysilicon 422 -2836 422 -2836 0 3
rlabel polysilicon 429 -2830 429 -2830 0 1
rlabel polysilicon 429 -2836 429 -2836 0 3
rlabel polysilicon 436 -2830 436 -2830 0 1
rlabel polysilicon 436 -2836 436 -2836 0 3
rlabel polysilicon 443 -2830 443 -2830 0 1
rlabel polysilicon 443 -2836 443 -2836 0 3
rlabel polysilicon 450 -2830 450 -2830 0 1
rlabel polysilicon 450 -2836 450 -2836 0 3
rlabel polysilicon 457 -2830 457 -2830 0 1
rlabel polysilicon 457 -2836 457 -2836 0 3
rlabel polysilicon 464 -2830 464 -2830 0 1
rlabel polysilicon 464 -2836 464 -2836 0 3
rlabel polysilicon 471 -2830 471 -2830 0 1
rlabel polysilicon 471 -2836 471 -2836 0 3
rlabel polysilicon 478 -2830 478 -2830 0 1
rlabel polysilicon 481 -2830 481 -2830 0 2
rlabel polysilicon 478 -2836 478 -2836 0 3
rlabel polysilicon 481 -2836 481 -2836 0 4
rlabel polysilicon 485 -2830 485 -2830 0 1
rlabel polysilicon 485 -2836 485 -2836 0 3
rlabel polysilicon 492 -2830 492 -2830 0 1
rlabel polysilicon 492 -2836 492 -2836 0 3
rlabel polysilicon 499 -2830 499 -2830 0 1
rlabel polysilicon 499 -2836 499 -2836 0 3
rlabel polysilicon 506 -2830 506 -2830 0 1
rlabel polysilicon 506 -2836 506 -2836 0 3
rlabel polysilicon 513 -2830 513 -2830 0 1
rlabel polysilicon 513 -2836 513 -2836 0 3
rlabel polysilicon 520 -2830 520 -2830 0 1
rlabel polysilicon 520 -2836 520 -2836 0 3
rlabel polysilicon 527 -2830 527 -2830 0 1
rlabel polysilicon 527 -2836 527 -2836 0 3
rlabel polysilicon 534 -2830 534 -2830 0 1
rlabel polysilicon 534 -2836 534 -2836 0 3
rlabel polysilicon 541 -2830 541 -2830 0 1
rlabel polysilicon 541 -2836 541 -2836 0 3
rlabel polysilicon 548 -2830 548 -2830 0 1
rlabel polysilicon 548 -2836 548 -2836 0 3
rlabel polysilicon 555 -2830 555 -2830 0 1
rlabel polysilicon 555 -2836 555 -2836 0 3
rlabel polysilicon 558 -2836 558 -2836 0 4
rlabel polysilicon 562 -2830 562 -2830 0 1
rlabel polysilicon 565 -2830 565 -2830 0 2
rlabel polysilicon 562 -2836 562 -2836 0 3
rlabel polysilicon 565 -2836 565 -2836 0 4
rlabel polysilicon 569 -2830 569 -2830 0 1
rlabel polysilicon 569 -2836 569 -2836 0 3
rlabel polysilicon 576 -2830 576 -2830 0 1
rlabel polysilicon 576 -2836 576 -2836 0 3
rlabel polysilicon 583 -2830 583 -2830 0 1
rlabel polysilicon 583 -2836 583 -2836 0 3
rlabel polysilicon 586 -2836 586 -2836 0 4
rlabel polysilicon 590 -2830 590 -2830 0 1
rlabel polysilicon 590 -2836 590 -2836 0 3
rlabel polysilicon 597 -2830 597 -2830 0 1
rlabel polysilicon 597 -2836 597 -2836 0 3
rlabel polysilicon 604 -2830 604 -2830 0 1
rlabel polysilicon 604 -2836 604 -2836 0 3
rlabel polysilicon 611 -2830 611 -2830 0 1
rlabel polysilicon 611 -2836 611 -2836 0 3
rlabel polysilicon 618 -2830 618 -2830 0 1
rlabel polysilicon 621 -2830 621 -2830 0 2
rlabel polysilicon 618 -2836 618 -2836 0 3
rlabel polysilicon 621 -2836 621 -2836 0 4
rlabel polysilicon 625 -2830 625 -2830 0 1
rlabel polysilicon 625 -2836 625 -2836 0 3
rlabel polysilicon 632 -2830 632 -2830 0 1
rlabel polysilicon 632 -2836 632 -2836 0 3
rlabel polysilicon 639 -2830 639 -2830 0 1
rlabel polysilicon 639 -2836 639 -2836 0 3
rlabel polysilicon 646 -2830 646 -2830 0 1
rlabel polysilicon 646 -2836 646 -2836 0 3
rlabel polysilicon 653 -2830 653 -2830 0 1
rlabel polysilicon 653 -2836 653 -2836 0 3
rlabel polysilicon 660 -2830 660 -2830 0 1
rlabel polysilicon 663 -2830 663 -2830 0 2
rlabel polysilicon 660 -2836 660 -2836 0 3
rlabel polysilicon 663 -2836 663 -2836 0 4
rlabel polysilicon 667 -2830 667 -2830 0 1
rlabel polysilicon 667 -2836 667 -2836 0 3
rlabel polysilicon 674 -2830 674 -2830 0 1
rlabel polysilicon 674 -2836 674 -2836 0 3
rlabel polysilicon 681 -2830 681 -2830 0 1
rlabel polysilicon 681 -2836 681 -2836 0 3
rlabel polysilicon 688 -2830 688 -2830 0 1
rlabel polysilicon 688 -2836 688 -2836 0 3
rlabel polysilicon 695 -2830 695 -2830 0 1
rlabel polysilicon 695 -2836 695 -2836 0 3
rlabel polysilicon 702 -2830 702 -2830 0 1
rlabel polysilicon 705 -2830 705 -2830 0 2
rlabel polysilicon 705 -2836 705 -2836 0 4
rlabel polysilicon 709 -2830 709 -2830 0 1
rlabel polysilicon 712 -2830 712 -2830 0 2
rlabel polysilicon 712 -2836 712 -2836 0 4
rlabel polysilicon 716 -2830 716 -2830 0 1
rlabel polysilicon 716 -2836 716 -2836 0 3
rlabel polysilicon 723 -2830 723 -2830 0 1
rlabel polysilicon 723 -2836 723 -2836 0 3
rlabel polysilicon 730 -2830 730 -2830 0 1
rlabel polysilicon 733 -2830 733 -2830 0 2
rlabel polysilicon 733 -2836 733 -2836 0 4
rlabel polysilicon 737 -2830 737 -2830 0 1
rlabel polysilicon 737 -2836 737 -2836 0 3
rlabel polysilicon 744 -2830 744 -2830 0 1
rlabel polysilicon 744 -2836 744 -2836 0 3
rlabel polysilicon 751 -2830 751 -2830 0 1
rlabel polysilicon 751 -2836 751 -2836 0 3
rlabel polysilicon 758 -2830 758 -2830 0 1
rlabel polysilicon 758 -2836 758 -2836 0 3
rlabel polysilicon 765 -2830 765 -2830 0 1
rlabel polysilicon 765 -2836 765 -2836 0 3
rlabel polysilicon 772 -2830 772 -2830 0 1
rlabel polysilicon 772 -2836 772 -2836 0 3
rlabel polysilicon 779 -2830 779 -2830 0 1
rlabel polysilicon 779 -2836 779 -2836 0 3
rlabel polysilicon 786 -2830 786 -2830 0 1
rlabel polysilicon 786 -2836 786 -2836 0 3
rlabel polysilicon 793 -2830 793 -2830 0 1
rlabel polysilicon 793 -2836 793 -2836 0 3
rlabel polysilicon 800 -2830 800 -2830 0 1
rlabel polysilicon 800 -2836 800 -2836 0 3
rlabel polysilicon 807 -2830 807 -2830 0 1
rlabel polysilicon 807 -2836 807 -2836 0 3
rlabel polysilicon 814 -2830 814 -2830 0 1
rlabel polysilicon 814 -2836 814 -2836 0 3
rlabel polysilicon 821 -2830 821 -2830 0 1
rlabel polysilicon 821 -2836 821 -2836 0 3
rlabel polysilicon 831 -2830 831 -2830 0 2
rlabel polysilicon 828 -2836 828 -2836 0 3
rlabel polysilicon 835 -2830 835 -2830 0 1
rlabel polysilicon 835 -2836 835 -2836 0 3
rlabel polysilicon 842 -2830 842 -2830 0 1
rlabel polysilicon 842 -2836 842 -2836 0 3
rlabel polysilicon 849 -2830 849 -2830 0 1
rlabel polysilicon 852 -2830 852 -2830 0 2
rlabel polysilicon 849 -2836 849 -2836 0 3
rlabel polysilicon 852 -2836 852 -2836 0 4
rlabel polysilicon 856 -2830 856 -2830 0 1
rlabel polysilicon 859 -2830 859 -2830 0 2
rlabel polysilicon 856 -2836 856 -2836 0 3
rlabel polysilicon 859 -2836 859 -2836 0 4
rlabel polysilicon 863 -2830 863 -2830 0 1
rlabel polysilicon 863 -2836 863 -2836 0 3
rlabel polysilicon 870 -2836 870 -2836 0 3
rlabel polysilicon 873 -2836 873 -2836 0 4
rlabel polysilicon 877 -2830 877 -2830 0 1
rlabel polysilicon 877 -2836 877 -2836 0 3
rlabel polysilicon 884 -2830 884 -2830 0 1
rlabel polysilicon 884 -2836 884 -2836 0 3
rlabel polysilicon 891 -2830 891 -2830 0 1
rlabel polysilicon 891 -2836 891 -2836 0 3
rlabel polysilicon 898 -2830 898 -2830 0 1
rlabel polysilicon 898 -2836 898 -2836 0 3
rlabel polysilicon 905 -2830 905 -2830 0 1
rlabel polysilicon 905 -2836 905 -2836 0 3
rlabel polysilicon 912 -2830 912 -2830 0 1
rlabel polysilicon 912 -2836 912 -2836 0 3
rlabel polysilicon 919 -2830 919 -2830 0 1
rlabel polysilicon 919 -2836 919 -2836 0 3
rlabel polysilicon 926 -2830 926 -2830 0 1
rlabel polysilicon 926 -2836 926 -2836 0 3
rlabel polysilicon 933 -2830 933 -2830 0 1
rlabel polysilicon 933 -2836 933 -2836 0 3
rlabel polysilicon 940 -2830 940 -2830 0 1
rlabel polysilicon 940 -2836 940 -2836 0 3
rlabel polysilicon 947 -2830 947 -2830 0 1
rlabel polysilicon 947 -2836 947 -2836 0 3
rlabel polysilicon 954 -2830 954 -2830 0 1
rlabel polysilicon 954 -2836 954 -2836 0 3
rlabel polysilicon 961 -2830 961 -2830 0 1
rlabel polysilicon 961 -2836 961 -2836 0 3
rlabel polysilicon 968 -2830 968 -2830 0 1
rlabel polysilicon 968 -2836 968 -2836 0 3
rlabel polysilicon 975 -2830 975 -2830 0 1
rlabel polysilicon 975 -2836 975 -2836 0 3
rlabel polysilicon 982 -2830 982 -2830 0 1
rlabel polysilicon 982 -2836 982 -2836 0 3
rlabel polysilicon 989 -2830 989 -2830 0 1
rlabel polysilicon 989 -2836 989 -2836 0 3
rlabel polysilicon 996 -2830 996 -2830 0 1
rlabel polysilicon 999 -2836 999 -2836 0 4
rlabel polysilicon 1003 -2830 1003 -2830 0 1
rlabel polysilicon 1003 -2836 1003 -2836 0 3
rlabel polysilicon 1010 -2830 1010 -2830 0 1
rlabel polysilicon 1013 -2830 1013 -2830 0 2
rlabel polysilicon 1010 -2836 1010 -2836 0 3
rlabel polysilicon 1013 -2836 1013 -2836 0 4
rlabel polysilicon 1017 -2830 1017 -2830 0 1
rlabel polysilicon 1020 -2830 1020 -2830 0 2
rlabel polysilicon 1020 -2836 1020 -2836 0 4
rlabel polysilicon 1024 -2830 1024 -2830 0 1
rlabel polysilicon 1024 -2836 1024 -2836 0 3
rlabel polysilicon 1031 -2830 1031 -2830 0 1
rlabel polysilicon 1031 -2836 1031 -2836 0 3
rlabel polysilicon 1038 -2830 1038 -2830 0 1
rlabel polysilicon 1038 -2836 1038 -2836 0 3
rlabel polysilicon 1045 -2830 1045 -2830 0 1
rlabel polysilicon 1045 -2836 1045 -2836 0 3
rlabel polysilicon 1052 -2830 1052 -2830 0 1
rlabel polysilicon 1052 -2836 1052 -2836 0 3
rlabel polysilicon 1059 -2830 1059 -2830 0 1
rlabel polysilicon 1059 -2836 1059 -2836 0 3
rlabel polysilicon 1066 -2830 1066 -2830 0 1
rlabel polysilicon 1069 -2830 1069 -2830 0 2
rlabel polysilicon 1066 -2836 1066 -2836 0 3
rlabel polysilicon 1069 -2836 1069 -2836 0 4
rlabel polysilicon 1073 -2830 1073 -2830 0 1
rlabel polysilicon 1073 -2836 1073 -2836 0 3
rlabel polysilicon 1080 -2830 1080 -2830 0 1
rlabel polysilicon 1080 -2836 1080 -2836 0 3
rlabel polysilicon 1087 -2830 1087 -2830 0 1
rlabel polysilicon 1087 -2836 1087 -2836 0 3
rlabel polysilicon 1094 -2830 1094 -2830 0 1
rlabel polysilicon 1094 -2836 1094 -2836 0 3
rlabel polysilicon 1101 -2830 1101 -2830 0 1
rlabel polysilicon 1101 -2836 1101 -2836 0 3
rlabel polysilicon 1108 -2830 1108 -2830 0 1
rlabel polysilicon 1108 -2836 1108 -2836 0 3
rlabel polysilicon 1115 -2830 1115 -2830 0 1
rlabel polysilicon 1118 -2830 1118 -2830 0 2
rlabel polysilicon 1115 -2836 1115 -2836 0 3
rlabel polysilicon 1125 -2830 1125 -2830 0 2
rlabel polysilicon 1122 -2836 1122 -2836 0 3
rlabel polysilicon 1125 -2836 1125 -2836 0 4
rlabel polysilicon 1129 -2830 1129 -2830 0 1
rlabel polysilicon 1129 -2836 1129 -2836 0 3
rlabel polysilicon 1136 -2830 1136 -2830 0 1
rlabel polysilicon 1136 -2836 1136 -2836 0 3
rlabel polysilicon 1143 -2830 1143 -2830 0 1
rlabel polysilicon 1143 -2836 1143 -2836 0 3
rlabel polysilicon 1150 -2830 1150 -2830 0 1
rlabel polysilicon 1150 -2836 1150 -2836 0 3
rlabel polysilicon 1157 -2830 1157 -2830 0 1
rlabel polysilicon 1157 -2836 1157 -2836 0 3
rlabel polysilicon 1164 -2830 1164 -2830 0 1
rlabel polysilicon 1164 -2836 1164 -2836 0 3
rlabel polysilicon 1171 -2830 1171 -2830 0 1
rlabel polysilicon 1171 -2836 1171 -2836 0 3
rlabel polysilicon 1178 -2830 1178 -2830 0 1
rlabel polysilicon 1181 -2830 1181 -2830 0 2
rlabel polysilicon 1178 -2836 1178 -2836 0 3
rlabel polysilicon 1185 -2830 1185 -2830 0 1
rlabel polysilicon 1185 -2836 1185 -2836 0 3
rlabel polysilicon 1192 -2830 1192 -2830 0 1
rlabel polysilicon 1192 -2836 1192 -2836 0 3
rlabel polysilicon 1199 -2830 1199 -2830 0 1
rlabel polysilicon 1202 -2830 1202 -2830 0 2
rlabel polysilicon 1199 -2836 1199 -2836 0 3
rlabel polysilicon 1202 -2836 1202 -2836 0 4
rlabel polysilicon 1206 -2830 1206 -2830 0 1
rlabel polysilicon 1206 -2836 1206 -2836 0 3
rlabel polysilicon 1213 -2830 1213 -2830 0 1
rlabel polysilicon 1213 -2836 1213 -2836 0 3
rlabel polysilicon 1220 -2830 1220 -2830 0 1
rlabel polysilicon 1220 -2836 1220 -2836 0 3
rlabel polysilicon 1227 -2830 1227 -2830 0 1
rlabel polysilicon 1227 -2836 1227 -2836 0 3
rlabel polysilicon 1237 -2830 1237 -2830 0 2
rlabel polysilicon 1234 -2836 1234 -2836 0 3
rlabel polysilicon 1237 -2836 1237 -2836 0 4
rlabel polysilicon 1241 -2830 1241 -2830 0 1
rlabel polysilicon 1241 -2836 1241 -2836 0 3
rlabel polysilicon 1248 -2830 1248 -2830 0 1
rlabel polysilicon 1248 -2836 1248 -2836 0 3
rlabel polysilicon 1255 -2830 1255 -2830 0 1
rlabel polysilicon 1255 -2836 1255 -2836 0 3
rlabel polysilicon 1262 -2830 1262 -2830 0 1
rlabel polysilicon 1262 -2836 1262 -2836 0 3
rlabel polysilicon 1269 -2830 1269 -2830 0 1
rlabel polysilicon 1269 -2836 1269 -2836 0 3
rlabel polysilicon 1276 -2830 1276 -2830 0 1
rlabel polysilicon 1276 -2836 1276 -2836 0 3
rlabel polysilicon 1283 -2830 1283 -2830 0 1
rlabel polysilicon 1283 -2836 1283 -2836 0 3
rlabel polysilicon 1286 -2836 1286 -2836 0 4
rlabel polysilicon 1290 -2830 1290 -2830 0 1
rlabel polysilicon 1290 -2836 1290 -2836 0 3
rlabel polysilicon 1297 -2830 1297 -2830 0 1
rlabel polysilicon 1297 -2836 1297 -2836 0 3
rlabel polysilicon 1304 -2830 1304 -2830 0 1
rlabel polysilicon 1304 -2836 1304 -2836 0 3
rlabel polysilicon 1311 -2830 1311 -2830 0 1
rlabel polysilicon 1311 -2836 1311 -2836 0 3
rlabel polysilicon 1318 -2830 1318 -2830 0 1
rlabel polysilicon 1318 -2836 1318 -2836 0 3
rlabel polysilicon 1325 -2830 1325 -2830 0 1
rlabel polysilicon 1325 -2836 1325 -2836 0 3
rlabel polysilicon 1332 -2830 1332 -2830 0 1
rlabel polysilicon 1332 -2836 1332 -2836 0 3
rlabel polysilicon 1342 -2830 1342 -2830 0 2
rlabel polysilicon 1342 -2836 1342 -2836 0 4
rlabel polysilicon 1346 -2830 1346 -2830 0 1
rlabel polysilicon 1346 -2836 1346 -2836 0 3
rlabel polysilicon 1353 -2830 1353 -2830 0 1
rlabel polysilicon 1353 -2836 1353 -2836 0 3
rlabel polysilicon 1356 -2836 1356 -2836 0 4
rlabel polysilicon 1360 -2830 1360 -2830 0 1
rlabel polysilicon 1360 -2836 1360 -2836 0 3
rlabel polysilicon 1367 -2830 1367 -2830 0 1
rlabel polysilicon 1367 -2836 1367 -2836 0 3
rlabel polysilicon 1374 -2830 1374 -2830 0 1
rlabel polysilicon 1374 -2836 1374 -2836 0 3
rlabel polysilicon 1381 -2830 1381 -2830 0 1
rlabel polysilicon 1381 -2836 1381 -2836 0 3
rlabel polysilicon 1388 -2830 1388 -2830 0 1
rlabel polysilicon 1388 -2836 1388 -2836 0 3
rlabel polysilicon 1395 -2830 1395 -2830 0 1
rlabel polysilicon 1395 -2836 1395 -2836 0 3
rlabel polysilicon 1402 -2830 1402 -2830 0 1
rlabel polysilicon 1402 -2836 1402 -2836 0 3
rlabel polysilicon 1409 -2830 1409 -2830 0 1
rlabel polysilicon 1409 -2836 1409 -2836 0 3
rlabel polysilicon 1416 -2830 1416 -2830 0 1
rlabel polysilicon 1416 -2836 1416 -2836 0 3
rlabel polysilicon 1423 -2830 1423 -2830 0 1
rlabel polysilicon 1423 -2836 1423 -2836 0 3
rlabel polysilicon 1430 -2830 1430 -2830 0 1
rlabel polysilicon 1433 -2830 1433 -2830 0 2
rlabel polysilicon 1430 -2836 1430 -2836 0 3
rlabel polysilicon 1433 -2836 1433 -2836 0 4
rlabel polysilicon 1437 -2830 1437 -2830 0 1
rlabel polysilicon 1437 -2836 1437 -2836 0 3
rlabel polysilicon 1444 -2830 1444 -2830 0 1
rlabel polysilicon 1444 -2836 1444 -2836 0 3
rlabel polysilicon 1451 -2830 1451 -2830 0 1
rlabel polysilicon 1451 -2836 1451 -2836 0 3
rlabel polysilicon 1458 -2830 1458 -2830 0 1
rlabel polysilicon 1458 -2836 1458 -2836 0 3
rlabel polysilicon 1465 -2830 1465 -2830 0 1
rlabel polysilicon 1465 -2836 1465 -2836 0 3
rlabel polysilicon 1472 -2830 1472 -2830 0 1
rlabel polysilicon 1472 -2836 1472 -2836 0 3
rlabel polysilicon 1479 -2830 1479 -2830 0 1
rlabel polysilicon 1479 -2836 1479 -2836 0 3
rlabel polysilicon 1486 -2830 1486 -2830 0 1
rlabel polysilicon 1486 -2836 1486 -2836 0 3
rlabel polysilicon 1493 -2830 1493 -2830 0 1
rlabel polysilicon 1493 -2836 1493 -2836 0 3
rlabel polysilicon 1500 -2830 1500 -2830 0 1
rlabel polysilicon 1500 -2836 1500 -2836 0 3
rlabel polysilicon 1507 -2830 1507 -2830 0 1
rlabel polysilicon 1507 -2836 1507 -2836 0 3
rlabel polysilicon 1514 -2830 1514 -2830 0 1
rlabel polysilicon 1514 -2836 1514 -2836 0 3
rlabel polysilicon 1521 -2830 1521 -2830 0 1
rlabel polysilicon 1521 -2836 1521 -2836 0 3
rlabel polysilicon 1528 -2830 1528 -2830 0 1
rlabel polysilicon 1528 -2836 1528 -2836 0 3
rlabel polysilicon 1535 -2830 1535 -2830 0 1
rlabel polysilicon 1535 -2836 1535 -2836 0 3
rlabel polysilicon 1542 -2830 1542 -2830 0 1
rlabel polysilicon 1542 -2836 1542 -2836 0 3
rlabel polysilicon 1549 -2830 1549 -2830 0 1
rlabel polysilicon 1549 -2836 1549 -2836 0 3
rlabel polysilicon 1556 -2830 1556 -2830 0 1
rlabel polysilicon 1556 -2836 1556 -2836 0 3
rlabel polysilicon 1563 -2830 1563 -2830 0 1
rlabel polysilicon 1563 -2836 1563 -2836 0 3
rlabel polysilicon 1570 -2830 1570 -2830 0 1
rlabel polysilicon 1570 -2836 1570 -2836 0 3
rlabel polysilicon 1577 -2830 1577 -2830 0 1
rlabel polysilicon 1577 -2836 1577 -2836 0 3
rlabel polysilicon 1584 -2830 1584 -2830 0 1
rlabel polysilicon 1584 -2836 1584 -2836 0 3
rlabel polysilicon 1591 -2830 1591 -2830 0 1
rlabel polysilicon 1591 -2836 1591 -2836 0 3
rlabel polysilicon 1598 -2830 1598 -2830 0 1
rlabel polysilicon 1598 -2836 1598 -2836 0 3
rlabel polysilicon 1605 -2830 1605 -2830 0 1
rlabel polysilicon 1605 -2836 1605 -2836 0 3
rlabel polysilicon 1612 -2830 1612 -2830 0 1
rlabel polysilicon 1612 -2836 1612 -2836 0 3
rlabel polysilicon 1619 -2830 1619 -2830 0 1
rlabel polysilicon 1619 -2836 1619 -2836 0 3
rlabel polysilicon 1626 -2830 1626 -2830 0 1
rlabel polysilicon 1626 -2836 1626 -2836 0 3
rlabel polysilicon 1633 -2830 1633 -2830 0 1
rlabel polysilicon 1633 -2836 1633 -2836 0 3
rlabel polysilicon 1640 -2830 1640 -2830 0 1
rlabel polysilicon 1640 -2836 1640 -2836 0 3
rlabel polysilicon 1647 -2830 1647 -2830 0 1
rlabel polysilicon 1647 -2836 1647 -2836 0 3
rlabel polysilicon 1654 -2830 1654 -2830 0 1
rlabel polysilicon 1654 -2836 1654 -2836 0 3
rlabel polysilicon 1661 -2830 1661 -2830 0 1
rlabel polysilicon 1661 -2836 1661 -2836 0 3
rlabel polysilicon 1668 -2830 1668 -2830 0 1
rlabel polysilicon 1668 -2836 1668 -2836 0 3
rlabel polysilicon 1675 -2830 1675 -2830 0 1
rlabel polysilicon 1675 -2836 1675 -2836 0 3
rlabel polysilicon 1682 -2830 1682 -2830 0 1
rlabel polysilicon 1682 -2836 1682 -2836 0 3
rlabel polysilicon 1689 -2830 1689 -2830 0 1
rlabel polysilicon 1689 -2836 1689 -2836 0 3
rlabel polysilicon 1696 -2830 1696 -2830 0 1
rlabel polysilicon 1696 -2836 1696 -2836 0 3
rlabel polysilicon 1703 -2830 1703 -2830 0 1
rlabel polysilicon 1703 -2836 1703 -2836 0 3
rlabel polysilicon 1710 -2830 1710 -2830 0 1
rlabel polysilicon 1713 -2830 1713 -2830 0 2
rlabel polysilicon 1710 -2836 1710 -2836 0 3
rlabel polysilicon 1713 -2836 1713 -2836 0 4
rlabel polysilicon 1717 -2830 1717 -2830 0 1
rlabel polysilicon 1720 -2830 1720 -2830 0 2
rlabel polysilicon 1717 -2836 1717 -2836 0 3
rlabel polysilicon 1720 -2836 1720 -2836 0 4
rlabel polysilicon 1724 -2830 1724 -2830 0 1
rlabel polysilicon 1724 -2836 1724 -2836 0 3
rlabel polysilicon 1727 -2836 1727 -2836 0 4
rlabel polysilicon 1731 -2830 1731 -2830 0 1
rlabel polysilicon 1731 -2836 1731 -2836 0 3
rlabel polysilicon 1738 -2830 1738 -2830 0 1
rlabel polysilicon 1738 -2836 1738 -2836 0 3
rlabel polysilicon 1745 -2830 1745 -2830 0 1
rlabel polysilicon 1745 -2836 1745 -2836 0 3
rlabel polysilicon 1752 -2830 1752 -2830 0 1
rlabel polysilicon 1752 -2836 1752 -2836 0 3
rlabel polysilicon 1759 -2830 1759 -2830 0 1
rlabel polysilicon 1759 -2836 1759 -2836 0 3
rlabel polysilicon 1766 -2830 1766 -2830 0 1
rlabel polysilicon 1766 -2836 1766 -2836 0 3
rlabel polysilicon 1773 -2830 1773 -2830 0 1
rlabel polysilicon 1773 -2836 1773 -2836 0 3
rlabel polysilicon 23 -2949 23 -2949 0 1
rlabel polysilicon 23 -2955 23 -2955 0 3
rlabel polysilicon 51 -2949 51 -2949 0 1
rlabel polysilicon 51 -2955 51 -2955 0 3
rlabel polysilicon 58 -2949 58 -2949 0 1
rlabel polysilicon 58 -2955 58 -2955 0 3
rlabel polysilicon 65 -2949 65 -2949 0 1
rlabel polysilicon 65 -2955 65 -2955 0 3
rlabel polysilicon 72 -2949 72 -2949 0 1
rlabel polysilicon 72 -2955 72 -2955 0 3
rlabel polysilicon 82 -2949 82 -2949 0 2
rlabel polysilicon 79 -2955 79 -2955 0 3
rlabel polysilicon 82 -2955 82 -2955 0 4
rlabel polysilicon 86 -2949 86 -2949 0 1
rlabel polysilicon 86 -2955 86 -2955 0 3
rlabel polysilicon 93 -2949 93 -2949 0 1
rlabel polysilicon 93 -2955 93 -2955 0 3
rlabel polysilicon 100 -2949 100 -2949 0 1
rlabel polysilicon 100 -2955 100 -2955 0 3
rlabel polysilicon 107 -2949 107 -2949 0 1
rlabel polysilicon 110 -2949 110 -2949 0 2
rlabel polysilicon 107 -2955 107 -2955 0 3
rlabel polysilicon 110 -2955 110 -2955 0 4
rlabel polysilicon 114 -2949 114 -2949 0 1
rlabel polysilicon 114 -2955 114 -2955 0 3
rlabel polysilicon 121 -2949 121 -2949 0 1
rlabel polysilicon 121 -2955 121 -2955 0 3
rlabel polysilicon 128 -2949 128 -2949 0 1
rlabel polysilicon 128 -2955 128 -2955 0 3
rlabel polysilicon 135 -2955 135 -2955 0 3
rlabel polysilicon 138 -2955 138 -2955 0 4
rlabel polysilicon 142 -2949 142 -2949 0 1
rlabel polysilicon 145 -2949 145 -2949 0 2
rlabel polysilicon 142 -2955 142 -2955 0 3
rlabel polysilicon 149 -2949 149 -2949 0 1
rlabel polysilicon 149 -2955 149 -2955 0 3
rlabel polysilicon 156 -2949 156 -2949 0 1
rlabel polysilicon 156 -2955 156 -2955 0 3
rlabel polysilicon 163 -2949 163 -2949 0 1
rlabel polysilicon 166 -2949 166 -2949 0 2
rlabel polysilicon 163 -2955 163 -2955 0 3
rlabel polysilicon 170 -2949 170 -2949 0 1
rlabel polysilicon 170 -2955 170 -2955 0 3
rlabel polysilicon 177 -2949 177 -2949 0 1
rlabel polysilicon 177 -2955 177 -2955 0 3
rlabel polysilicon 184 -2949 184 -2949 0 1
rlabel polysilicon 184 -2955 184 -2955 0 3
rlabel polysilicon 191 -2949 191 -2949 0 1
rlabel polysilicon 191 -2955 191 -2955 0 3
rlabel polysilicon 198 -2949 198 -2949 0 1
rlabel polysilicon 198 -2955 198 -2955 0 3
rlabel polysilicon 205 -2949 205 -2949 0 1
rlabel polysilicon 208 -2949 208 -2949 0 2
rlabel polysilicon 205 -2955 205 -2955 0 3
rlabel polysilicon 212 -2949 212 -2949 0 1
rlabel polysilicon 212 -2955 212 -2955 0 3
rlabel polysilicon 219 -2949 219 -2949 0 1
rlabel polysilicon 219 -2955 219 -2955 0 3
rlabel polysilicon 226 -2949 226 -2949 0 1
rlabel polysilicon 229 -2949 229 -2949 0 2
rlabel polysilicon 226 -2955 226 -2955 0 3
rlabel polysilicon 233 -2949 233 -2949 0 1
rlabel polysilicon 233 -2955 233 -2955 0 3
rlabel polysilicon 240 -2949 240 -2949 0 1
rlabel polysilicon 240 -2955 240 -2955 0 3
rlabel polysilicon 247 -2949 247 -2949 0 1
rlabel polysilicon 247 -2955 247 -2955 0 3
rlabel polysilicon 254 -2949 254 -2949 0 1
rlabel polysilicon 254 -2955 254 -2955 0 3
rlabel polysilicon 261 -2949 261 -2949 0 1
rlabel polysilicon 261 -2955 261 -2955 0 3
rlabel polysilicon 268 -2949 268 -2949 0 1
rlabel polysilicon 268 -2955 268 -2955 0 3
rlabel polysilicon 275 -2949 275 -2949 0 1
rlabel polysilicon 275 -2955 275 -2955 0 3
rlabel polysilicon 282 -2949 282 -2949 0 1
rlabel polysilicon 282 -2955 282 -2955 0 3
rlabel polysilicon 289 -2949 289 -2949 0 1
rlabel polysilicon 289 -2955 289 -2955 0 3
rlabel polysilicon 296 -2949 296 -2949 0 1
rlabel polysilicon 296 -2955 296 -2955 0 3
rlabel polysilicon 303 -2949 303 -2949 0 1
rlabel polysilicon 303 -2955 303 -2955 0 3
rlabel polysilicon 310 -2949 310 -2949 0 1
rlabel polysilicon 310 -2955 310 -2955 0 3
rlabel polysilicon 317 -2949 317 -2949 0 1
rlabel polysilicon 317 -2955 317 -2955 0 3
rlabel polysilicon 324 -2949 324 -2949 0 1
rlabel polysilicon 324 -2955 324 -2955 0 3
rlabel polysilicon 331 -2949 331 -2949 0 1
rlabel polysilicon 331 -2955 331 -2955 0 3
rlabel polysilicon 338 -2949 338 -2949 0 1
rlabel polysilicon 338 -2955 338 -2955 0 3
rlabel polysilicon 345 -2949 345 -2949 0 1
rlabel polysilicon 345 -2955 345 -2955 0 3
rlabel polysilicon 352 -2949 352 -2949 0 1
rlabel polysilicon 352 -2955 352 -2955 0 3
rlabel polysilicon 359 -2949 359 -2949 0 1
rlabel polysilicon 359 -2955 359 -2955 0 3
rlabel polysilicon 366 -2949 366 -2949 0 1
rlabel polysilicon 366 -2955 366 -2955 0 3
rlabel polysilicon 373 -2949 373 -2949 0 1
rlabel polysilicon 373 -2955 373 -2955 0 3
rlabel polysilicon 380 -2949 380 -2949 0 1
rlabel polysilicon 380 -2955 380 -2955 0 3
rlabel polysilicon 387 -2949 387 -2949 0 1
rlabel polysilicon 387 -2955 387 -2955 0 3
rlabel polysilicon 394 -2949 394 -2949 0 1
rlabel polysilicon 394 -2955 394 -2955 0 3
rlabel polysilicon 401 -2949 401 -2949 0 1
rlabel polysilicon 401 -2955 401 -2955 0 3
rlabel polysilicon 411 -2949 411 -2949 0 2
rlabel polysilicon 408 -2955 408 -2955 0 3
rlabel polysilicon 411 -2955 411 -2955 0 4
rlabel polysilicon 415 -2949 415 -2949 0 1
rlabel polysilicon 415 -2955 415 -2955 0 3
rlabel polysilicon 422 -2949 422 -2949 0 1
rlabel polysilicon 422 -2955 422 -2955 0 3
rlabel polysilicon 429 -2949 429 -2949 0 1
rlabel polysilicon 429 -2955 429 -2955 0 3
rlabel polysilicon 436 -2949 436 -2949 0 1
rlabel polysilicon 439 -2949 439 -2949 0 2
rlabel polysilicon 439 -2955 439 -2955 0 4
rlabel polysilicon 443 -2949 443 -2949 0 1
rlabel polysilicon 443 -2955 443 -2955 0 3
rlabel polysilicon 450 -2949 450 -2949 0 1
rlabel polysilicon 450 -2955 450 -2955 0 3
rlabel polysilicon 457 -2949 457 -2949 0 1
rlabel polysilicon 457 -2955 457 -2955 0 3
rlabel polysilicon 464 -2949 464 -2949 0 1
rlabel polysilicon 467 -2949 467 -2949 0 2
rlabel polysilicon 464 -2955 464 -2955 0 3
rlabel polysilicon 471 -2949 471 -2949 0 1
rlabel polysilicon 471 -2955 471 -2955 0 3
rlabel polysilicon 478 -2949 478 -2949 0 1
rlabel polysilicon 478 -2955 478 -2955 0 3
rlabel polysilicon 485 -2949 485 -2949 0 1
rlabel polysilicon 485 -2955 485 -2955 0 3
rlabel polysilicon 492 -2949 492 -2949 0 1
rlabel polysilicon 492 -2955 492 -2955 0 3
rlabel polysilicon 499 -2949 499 -2949 0 1
rlabel polysilicon 499 -2955 499 -2955 0 3
rlabel polysilicon 506 -2949 506 -2949 0 1
rlabel polysilicon 506 -2955 506 -2955 0 3
rlabel polysilicon 513 -2949 513 -2949 0 1
rlabel polysilicon 513 -2955 513 -2955 0 3
rlabel polysilicon 520 -2949 520 -2949 0 1
rlabel polysilicon 520 -2955 520 -2955 0 3
rlabel polysilicon 527 -2949 527 -2949 0 1
rlabel polysilicon 527 -2955 527 -2955 0 3
rlabel polysilicon 534 -2949 534 -2949 0 1
rlabel polysilicon 537 -2949 537 -2949 0 2
rlabel polysilicon 534 -2955 534 -2955 0 3
rlabel polysilicon 537 -2955 537 -2955 0 4
rlabel polysilicon 541 -2949 541 -2949 0 1
rlabel polysilicon 541 -2955 541 -2955 0 3
rlabel polysilicon 548 -2949 548 -2949 0 1
rlabel polysilicon 548 -2955 548 -2955 0 3
rlabel polysilicon 555 -2949 555 -2949 0 1
rlabel polysilicon 555 -2955 555 -2955 0 3
rlabel polysilicon 562 -2949 562 -2949 0 1
rlabel polysilicon 562 -2955 562 -2955 0 3
rlabel polysilicon 569 -2949 569 -2949 0 1
rlabel polysilicon 569 -2955 569 -2955 0 3
rlabel polysilicon 576 -2949 576 -2949 0 1
rlabel polysilicon 576 -2955 576 -2955 0 3
rlabel polysilicon 583 -2949 583 -2949 0 1
rlabel polysilicon 583 -2955 583 -2955 0 3
rlabel polysilicon 590 -2949 590 -2949 0 1
rlabel polysilicon 590 -2955 590 -2955 0 3
rlabel polysilicon 597 -2949 597 -2949 0 1
rlabel polysilicon 597 -2955 597 -2955 0 3
rlabel polysilicon 604 -2949 604 -2949 0 1
rlabel polysilicon 604 -2955 604 -2955 0 3
rlabel polysilicon 611 -2949 611 -2949 0 1
rlabel polysilicon 611 -2955 611 -2955 0 3
rlabel polysilicon 618 -2949 618 -2949 0 1
rlabel polysilicon 618 -2955 618 -2955 0 3
rlabel polysilicon 625 -2949 625 -2949 0 1
rlabel polysilicon 625 -2955 625 -2955 0 3
rlabel polysilicon 632 -2949 632 -2949 0 1
rlabel polysilicon 632 -2955 632 -2955 0 3
rlabel polysilicon 639 -2949 639 -2949 0 1
rlabel polysilicon 639 -2955 639 -2955 0 3
rlabel polysilicon 646 -2949 646 -2949 0 1
rlabel polysilicon 646 -2955 646 -2955 0 3
rlabel polysilicon 653 -2949 653 -2949 0 1
rlabel polysilicon 656 -2949 656 -2949 0 2
rlabel polysilicon 653 -2955 653 -2955 0 3
rlabel polysilicon 656 -2955 656 -2955 0 4
rlabel polysilicon 660 -2949 660 -2949 0 1
rlabel polysilicon 663 -2949 663 -2949 0 2
rlabel polysilicon 660 -2955 660 -2955 0 3
rlabel polysilicon 663 -2955 663 -2955 0 4
rlabel polysilicon 667 -2949 667 -2949 0 1
rlabel polysilicon 667 -2955 667 -2955 0 3
rlabel polysilicon 674 -2949 674 -2949 0 1
rlabel polysilicon 674 -2955 674 -2955 0 3
rlabel polysilicon 681 -2949 681 -2949 0 1
rlabel polysilicon 681 -2955 681 -2955 0 3
rlabel polysilicon 688 -2949 688 -2949 0 1
rlabel polysilicon 688 -2955 688 -2955 0 3
rlabel polysilicon 695 -2949 695 -2949 0 1
rlabel polysilicon 695 -2955 695 -2955 0 3
rlabel polysilicon 702 -2949 702 -2949 0 1
rlabel polysilicon 702 -2955 702 -2955 0 3
rlabel polysilicon 709 -2949 709 -2949 0 1
rlabel polysilicon 709 -2955 709 -2955 0 3
rlabel polysilicon 716 -2949 716 -2949 0 1
rlabel polysilicon 716 -2955 716 -2955 0 3
rlabel polysilicon 723 -2949 723 -2949 0 1
rlabel polysilicon 723 -2955 723 -2955 0 3
rlabel polysilicon 730 -2949 730 -2949 0 1
rlabel polysilicon 730 -2955 730 -2955 0 3
rlabel polysilicon 737 -2949 737 -2949 0 1
rlabel polysilicon 737 -2955 737 -2955 0 3
rlabel polysilicon 744 -2949 744 -2949 0 1
rlabel polysilicon 744 -2955 744 -2955 0 3
rlabel polysilicon 751 -2949 751 -2949 0 1
rlabel polysilicon 751 -2955 751 -2955 0 3
rlabel polysilicon 758 -2949 758 -2949 0 1
rlabel polysilicon 758 -2955 758 -2955 0 3
rlabel polysilicon 765 -2949 765 -2949 0 1
rlabel polysilicon 765 -2955 765 -2955 0 3
rlabel polysilicon 772 -2949 772 -2949 0 1
rlabel polysilicon 772 -2955 772 -2955 0 3
rlabel polysilicon 782 -2949 782 -2949 0 2
rlabel polysilicon 779 -2955 779 -2955 0 3
rlabel polysilicon 782 -2955 782 -2955 0 4
rlabel polysilicon 786 -2949 786 -2949 0 1
rlabel polysilicon 786 -2955 786 -2955 0 3
rlabel polysilicon 793 -2949 793 -2949 0 1
rlabel polysilicon 793 -2955 793 -2955 0 3
rlabel polysilicon 800 -2949 800 -2949 0 1
rlabel polysilicon 800 -2955 800 -2955 0 3
rlabel polysilicon 807 -2949 807 -2949 0 1
rlabel polysilicon 807 -2955 807 -2955 0 3
rlabel polysilicon 814 -2949 814 -2949 0 1
rlabel polysilicon 814 -2955 814 -2955 0 3
rlabel polysilicon 824 -2949 824 -2949 0 2
rlabel polysilicon 828 -2949 828 -2949 0 1
rlabel polysilicon 828 -2955 828 -2955 0 3
rlabel polysilicon 835 -2949 835 -2949 0 1
rlabel polysilicon 835 -2955 835 -2955 0 3
rlabel polysilicon 842 -2949 842 -2949 0 1
rlabel polysilicon 842 -2955 842 -2955 0 3
rlabel polysilicon 849 -2949 849 -2949 0 1
rlabel polysilicon 852 -2949 852 -2949 0 2
rlabel polysilicon 849 -2955 849 -2955 0 3
rlabel polysilicon 852 -2955 852 -2955 0 4
rlabel polysilicon 856 -2949 856 -2949 0 1
rlabel polysilicon 856 -2955 856 -2955 0 3
rlabel polysilicon 863 -2949 863 -2949 0 1
rlabel polysilicon 866 -2949 866 -2949 0 2
rlabel polysilicon 863 -2955 863 -2955 0 3
rlabel polysilicon 866 -2955 866 -2955 0 4
rlabel polysilicon 870 -2949 870 -2949 0 1
rlabel polysilicon 870 -2955 870 -2955 0 3
rlabel polysilicon 877 -2949 877 -2949 0 1
rlabel polysilicon 877 -2955 877 -2955 0 3
rlabel polysilicon 884 -2949 884 -2949 0 1
rlabel polysilicon 884 -2955 884 -2955 0 3
rlabel polysilicon 891 -2949 891 -2949 0 1
rlabel polysilicon 891 -2955 891 -2955 0 3
rlabel polysilicon 898 -2949 898 -2949 0 1
rlabel polysilicon 898 -2955 898 -2955 0 3
rlabel polysilicon 905 -2949 905 -2949 0 1
rlabel polysilicon 905 -2955 905 -2955 0 3
rlabel polysilicon 912 -2949 912 -2949 0 1
rlabel polysilicon 915 -2949 915 -2949 0 2
rlabel polysilicon 912 -2955 912 -2955 0 3
rlabel polysilicon 915 -2955 915 -2955 0 4
rlabel polysilicon 919 -2949 919 -2949 0 1
rlabel polysilicon 919 -2955 919 -2955 0 3
rlabel polysilicon 926 -2949 926 -2949 0 1
rlabel polysilicon 926 -2955 926 -2955 0 3
rlabel polysilicon 933 -2949 933 -2949 0 1
rlabel polysilicon 933 -2955 933 -2955 0 3
rlabel polysilicon 943 -2949 943 -2949 0 2
rlabel polysilicon 940 -2955 940 -2955 0 3
rlabel polysilicon 943 -2955 943 -2955 0 4
rlabel polysilicon 947 -2949 947 -2949 0 1
rlabel polysilicon 947 -2955 947 -2955 0 3
rlabel polysilicon 954 -2949 954 -2949 0 1
rlabel polysilicon 954 -2955 954 -2955 0 3
rlabel polysilicon 961 -2949 961 -2949 0 1
rlabel polysilicon 961 -2955 961 -2955 0 3
rlabel polysilicon 968 -2949 968 -2949 0 1
rlabel polysilicon 971 -2949 971 -2949 0 2
rlabel polysilicon 968 -2955 968 -2955 0 3
rlabel polysilicon 975 -2949 975 -2949 0 1
rlabel polysilicon 975 -2955 975 -2955 0 3
rlabel polysilicon 982 -2949 982 -2949 0 1
rlabel polysilicon 982 -2955 982 -2955 0 3
rlabel polysilicon 989 -2949 989 -2949 0 1
rlabel polysilicon 989 -2955 989 -2955 0 3
rlabel polysilicon 996 -2949 996 -2949 0 1
rlabel polysilicon 996 -2955 996 -2955 0 3
rlabel polysilicon 1003 -2949 1003 -2949 0 1
rlabel polysilicon 1003 -2955 1003 -2955 0 3
rlabel polysilicon 1010 -2949 1010 -2949 0 1
rlabel polysilicon 1010 -2955 1010 -2955 0 3
rlabel polysilicon 1017 -2949 1017 -2949 0 1
rlabel polysilicon 1017 -2955 1017 -2955 0 3
rlabel polysilicon 1024 -2949 1024 -2949 0 1
rlabel polysilicon 1027 -2949 1027 -2949 0 2
rlabel polysilicon 1024 -2955 1024 -2955 0 3
rlabel polysilicon 1027 -2955 1027 -2955 0 4
rlabel polysilicon 1031 -2949 1031 -2949 0 1
rlabel polysilicon 1031 -2955 1031 -2955 0 3
rlabel polysilicon 1034 -2955 1034 -2955 0 4
rlabel polysilicon 1038 -2949 1038 -2949 0 1
rlabel polysilicon 1038 -2955 1038 -2955 0 3
rlabel polysilicon 1045 -2949 1045 -2949 0 1
rlabel polysilicon 1045 -2955 1045 -2955 0 3
rlabel polysilicon 1052 -2949 1052 -2949 0 1
rlabel polysilicon 1055 -2949 1055 -2949 0 2
rlabel polysilicon 1055 -2955 1055 -2955 0 4
rlabel polysilicon 1059 -2949 1059 -2949 0 1
rlabel polysilicon 1059 -2955 1059 -2955 0 3
rlabel polysilicon 1066 -2949 1066 -2949 0 1
rlabel polysilicon 1066 -2955 1066 -2955 0 3
rlabel polysilicon 1073 -2949 1073 -2949 0 1
rlabel polysilicon 1073 -2955 1073 -2955 0 3
rlabel polysilicon 1080 -2949 1080 -2949 0 1
rlabel polysilicon 1080 -2955 1080 -2955 0 3
rlabel polysilicon 1087 -2949 1087 -2949 0 1
rlabel polysilicon 1087 -2955 1087 -2955 0 3
rlabel polysilicon 1097 -2949 1097 -2949 0 2
rlabel polysilicon 1097 -2955 1097 -2955 0 4
rlabel polysilicon 1101 -2949 1101 -2949 0 1
rlabel polysilicon 1101 -2955 1101 -2955 0 3
rlabel polysilicon 1108 -2949 1108 -2949 0 1
rlabel polysilicon 1108 -2955 1108 -2955 0 3
rlabel polysilicon 1115 -2949 1115 -2949 0 1
rlabel polysilicon 1115 -2955 1115 -2955 0 3
rlabel polysilicon 1122 -2949 1122 -2949 0 1
rlabel polysilicon 1122 -2955 1122 -2955 0 3
rlabel polysilicon 1129 -2949 1129 -2949 0 1
rlabel polysilicon 1129 -2955 1129 -2955 0 3
rlabel polysilicon 1136 -2949 1136 -2949 0 1
rlabel polysilicon 1136 -2955 1136 -2955 0 3
rlabel polysilicon 1143 -2949 1143 -2949 0 1
rlabel polysilicon 1143 -2955 1143 -2955 0 3
rlabel polysilicon 1150 -2949 1150 -2949 0 1
rlabel polysilicon 1150 -2955 1150 -2955 0 3
rlabel polysilicon 1157 -2949 1157 -2949 0 1
rlabel polysilicon 1157 -2955 1157 -2955 0 3
rlabel polysilicon 1164 -2949 1164 -2949 0 1
rlabel polysilicon 1164 -2955 1164 -2955 0 3
rlabel polysilicon 1171 -2949 1171 -2949 0 1
rlabel polysilicon 1171 -2955 1171 -2955 0 3
rlabel polysilicon 1178 -2949 1178 -2949 0 1
rlabel polysilicon 1178 -2955 1178 -2955 0 3
rlabel polysilicon 1185 -2949 1185 -2949 0 1
rlabel polysilicon 1185 -2955 1185 -2955 0 3
rlabel polysilicon 1192 -2949 1192 -2949 0 1
rlabel polysilicon 1192 -2955 1192 -2955 0 3
rlabel polysilicon 1202 -2949 1202 -2949 0 2
rlabel polysilicon 1199 -2955 1199 -2955 0 3
rlabel polysilicon 1202 -2955 1202 -2955 0 4
rlabel polysilicon 1206 -2949 1206 -2949 0 1
rlabel polysilicon 1206 -2955 1206 -2955 0 3
rlabel polysilicon 1213 -2949 1213 -2949 0 1
rlabel polysilicon 1213 -2955 1213 -2955 0 3
rlabel polysilicon 1220 -2949 1220 -2949 0 1
rlabel polysilicon 1220 -2955 1220 -2955 0 3
rlabel polysilicon 1227 -2949 1227 -2949 0 1
rlabel polysilicon 1227 -2955 1227 -2955 0 3
rlabel polysilicon 1234 -2949 1234 -2949 0 1
rlabel polysilicon 1234 -2955 1234 -2955 0 3
rlabel polysilicon 1241 -2949 1241 -2949 0 1
rlabel polysilicon 1241 -2955 1241 -2955 0 3
rlabel polysilicon 1248 -2949 1248 -2949 0 1
rlabel polysilicon 1248 -2955 1248 -2955 0 3
rlabel polysilicon 1255 -2949 1255 -2949 0 1
rlabel polysilicon 1255 -2955 1255 -2955 0 3
rlabel polysilicon 1262 -2949 1262 -2949 0 1
rlabel polysilicon 1262 -2955 1262 -2955 0 3
rlabel polysilicon 1269 -2949 1269 -2949 0 1
rlabel polysilicon 1269 -2955 1269 -2955 0 3
rlabel polysilicon 1276 -2949 1276 -2949 0 1
rlabel polysilicon 1276 -2955 1276 -2955 0 3
rlabel polysilicon 1283 -2949 1283 -2949 0 1
rlabel polysilicon 1283 -2955 1283 -2955 0 3
rlabel polysilicon 1290 -2949 1290 -2949 0 1
rlabel polysilicon 1290 -2955 1290 -2955 0 3
rlabel polysilicon 1297 -2949 1297 -2949 0 1
rlabel polysilicon 1297 -2955 1297 -2955 0 3
rlabel polysilicon 1304 -2949 1304 -2949 0 1
rlabel polysilicon 1304 -2955 1304 -2955 0 3
rlabel polysilicon 1311 -2949 1311 -2949 0 1
rlabel polysilicon 1311 -2955 1311 -2955 0 3
rlabel polysilicon 1318 -2949 1318 -2949 0 1
rlabel polysilicon 1318 -2955 1318 -2955 0 3
rlabel polysilicon 1325 -2949 1325 -2949 0 1
rlabel polysilicon 1325 -2955 1325 -2955 0 3
rlabel polysilicon 1332 -2955 1332 -2955 0 3
rlabel polysilicon 1335 -2955 1335 -2955 0 4
rlabel polysilicon 1339 -2949 1339 -2949 0 1
rlabel polysilicon 1339 -2955 1339 -2955 0 3
rlabel polysilicon 1346 -2949 1346 -2949 0 1
rlabel polysilicon 1346 -2955 1346 -2955 0 3
rlabel polysilicon 1353 -2949 1353 -2949 0 1
rlabel polysilicon 1353 -2955 1353 -2955 0 3
rlabel polysilicon 1360 -2949 1360 -2949 0 1
rlabel polysilicon 1360 -2955 1360 -2955 0 3
rlabel polysilicon 1367 -2949 1367 -2949 0 1
rlabel polysilicon 1367 -2955 1367 -2955 0 3
rlabel polysilicon 1374 -2949 1374 -2949 0 1
rlabel polysilicon 1374 -2955 1374 -2955 0 3
rlabel polysilicon 1381 -2949 1381 -2949 0 1
rlabel polysilicon 1381 -2955 1381 -2955 0 3
rlabel polysilicon 1388 -2949 1388 -2949 0 1
rlabel polysilicon 1388 -2955 1388 -2955 0 3
rlabel polysilicon 1395 -2949 1395 -2949 0 1
rlabel polysilicon 1395 -2955 1395 -2955 0 3
rlabel polysilicon 1402 -2949 1402 -2949 0 1
rlabel polysilicon 1402 -2955 1402 -2955 0 3
rlabel polysilicon 1409 -2949 1409 -2949 0 1
rlabel polysilicon 1409 -2955 1409 -2955 0 3
rlabel polysilicon 1416 -2949 1416 -2949 0 1
rlabel polysilicon 1416 -2955 1416 -2955 0 3
rlabel polysilicon 1423 -2949 1423 -2949 0 1
rlabel polysilicon 1423 -2955 1423 -2955 0 3
rlabel polysilicon 1430 -2949 1430 -2949 0 1
rlabel polysilicon 1430 -2955 1430 -2955 0 3
rlabel polysilicon 1437 -2949 1437 -2949 0 1
rlabel polysilicon 1437 -2955 1437 -2955 0 3
rlabel polysilicon 1444 -2949 1444 -2949 0 1
rlabel polysilicon 1444 -2955 1444 -2955 0 3
rlabel polysilicon 1451 -2949 1451 -2949 0 1
rlabel polysilicon 1451 -2955 1451 -2955 0 3
rlabel polysilicon 1458 -2949 1458 -2949 0 1
rlabel polysilicon 1458 -2955 1458 -2955 0 3
rlabel polysilicon 1465 -2949 1465 -2949 0 1
rlabel polysilicon 1465 -2955 1465 -2955 0 3
rlabel polysilicon 1472 -2949 1472 -2949 0 1
rlabel polysilicon 1472 -2955 1472 -2955 0 3
rlabel polysilicon 1479 -2949 1479 -2949 0 1
rlabel polysilicon 1479 -2955 1479 -2955 0 3
rlabel polysilicon 1486 -2949 1486 -2949 0 1
rlabel polysilicon 1486 -2955 1486 -2955 0 3
rlabel polysilicon 1493 -2949 1493 -2949 0 1
rlabel polysilicon 1493 -2955 1493 -2955 0 3
rlabel polysilicon 1500 -2949 1500 -2949 0 1
rlabel polysilicon 1500 -2955 1500 -2955 0 3
rlabel polysilicon 1507 -2949 1507 -2949 0 1
rlabel polysilicon 1507 -2955 1507 -2955 0 3
rlabel polysilicon 1514 -2949 1514 -2949 0 1
rlabel polysilicon 1514 -2955 1514 -2955 0 3
rlabel polysilicon 1521 -2949 1521 -2949 0 1
rlabel polysilicon 1521 -2955 1521 -2955 0 3
rlabel polysilicon 1528 -2949 1528 -2949 0 1
rlabel polysilicon 1528 -2955 1528 -2955 0 3
rlabel polysilicon 1535 -2949 1535 -2949 0 1
rlabel polysilicon 1535 -2955 1535 -2955 0 3
rlabel polysilicon 1542 -2949 1542 -2949 0 1
rlabel polysilicon 1542 -2955 1542 -2955 0 3
rlabel polysilicon 1549 -2949 1549 -2949 0 1
rlabel polysilicon 1549 -2955 1549 -2955 0 3
rlabel polysilicon 1556 -2949 1556 -2949 0 1
rlabel polysilicon 1556 -2955 1556 -2955 0 3
rlabel polysilicon 1563 -2949 1563 -2949 0 1
rlabel polysilicon 1563 -2955 1563 -2955 0 3
rlabel polysilicon 1570 -2949 1570 -2949 0 1
rlabel polysilicon 1570 -2955 1570 -2955 0 3
rlabel polysilicon 1577 -2949 1577 -2949 0 1
rlabel polysilicon 1577 -2955 1577 -2955 0 3
rlabel polysilicon 1584 -2949 1584 -2949 0 1
rlabel polysilicon 1584 -2955 1584 -2955 0 3
rlabel polysilicon 1591 -2949 1591 -2949 0 1
rlabel polysilicon 1591 -2955 1591 -2955 0 3
rlabel polysilicon 1598 -2949 1598 -2949 0 1
rlabel polysilicon 1598 -2955 1598 -2955 0 3
rlabel polysilicon 1605 -2949 1605 -2949 0 1
rlabel polysilicon 1605 -2955 1605 -2955 0 3
rlabel polysilicon 1612 -2949 1612 -2949 0 1
rlabel polysilicon 1612 -2955 1612 -2955 0 3
rlabel polysilicon 1619 -2949 1619 -2949 0 1
rlabel polysilicon 1619 -2955 1619 -2955 0 3
rlabel polysilicon 1626 -2949 1626 -2949 0 1
rlabel polysilicon 1626 -2955 1626 -2955 0 3
rlabel polysilicon 1633 -2949 1633 -2949 0 1
rlabel polysilicon 1633 -2955 1633 -2955 0 3
rlabel polysilicon 1640 -2949 1640 -2949 0 1
rlabel polysilicon 1640 -2955 1640 -2955 0 3
rlabel polysilicon 1647 -2949 1647 -2949 0 1
rlabel polysilicon 1647 -2955 1647 -2955 0 3
rlabel polysilicon 1654 -2949 1654 -2949 0 1
rlabel polysilicon 1654 -2955 1654 -2955 0 3
rlabel polysilicon 1661 -2949 1661 -2949 0 1
rlabel polysilicon 1661 -2955 1661 -2955 0 3
rlabel polysilicon 1668 -2949 1668 -2949 0 1
rlabel polysilicon 1668 -2955 1668 -2955 0 3
rlabel polysilicon 1675 -2949 1675 -2949 0 1
rlabel polysilicon 1675 -2955 1675 -2955 0 3
rlabel polysilicon 1682 -2949 1682 -2949 0 1
rlabel polysilicon 1682 -2955 1682 -2955 0 3
rlabel polysilicon 1689 -2949 1689 -2949 0 1
rlabel polysilicon 1689 -2955 1689 -2955 0 3
rlabel polysilicon 1696 -2949 1696 -2949 0 1
rlabel polysilicon 1696 -2955 1696 -2955 0 3
rlabel polysilicon 1703 -2949 1703 -2949 0 1
rlabel polysilicon 1703 -2955 1703 -2955 0 3
rlabel polysilicon 1706 -2955 1706 -2955 0 4
rlabel polysilicon 30 -3076 30 -3076 0 1
rlabel polysilicon 30 -3082 30 -3082 0 3
rlabel polysilicon 37 -3076 37 -3076 0 1
rlabel polysilicon 37 -3082 37 -3082 0 3
rlabel polysilicon 44 -3076 44 -3076 0 1
rlabel polysilicon 44 -3082 44 -3082 0 3
rlabel polysilicon 51 -3076 51 -3076 0 1
rlabel polysilicon 51 -3082 51 -3082 0 3
rlabel polysilicon 58 -3076 58 -3076 0 1
rlabel polysilicon 61 -3076 61 -3076 0 2
rlabel polysilicon 61 -3082 61 -3082 0 4
rlabel polysilicon 65 -3076 65 -3076 0 1
rlabel polysilicon 65 -3082 65 -3082 0 3
rlabel polysilicon 72 -3076 72 -3076 0 1
rlabel polysilicon 72 -3082 72 -3082 0 3
rlabel polysilicon 79 -3076 79 -3076 0 1
rlabel polysilicon 82 -3076 82 -3076 0 2
rlabel polysilicon 79 -3082 79 -3082 0 3
rlabel polysilicon 82 -3082 82 -3082 0 4
rlabel polysilicon 86 -3076 86 -3076 0 1
rlabel polysilicon 89 -3076 89 -3076 0 2
rlabel polysilicon 86 -3082 86 -3082 0 3
rlabel polysilicon 89 -3082 89 -3082 0 4
rlabel polysilicon 93 -3076 93 -3076 0 1
rlabel polysilicon 93 -3082 93 -3082 0 3
rlabel polysilicon 100 -3076 100 -3076 0 1
rlabel polysilicon 100 -3082 100 -3082 0 3
rlabel polysilicon 107 -3076 107 -3076 0 1
rlabel polysilicon 107 -3082 107 -3082 0 3
rlabel polysilicon 114 -3076 114 -3076 0 1
rlabel polysilicon 114 -3082 114 -3082 0 3
rlabel polysilicon 121 -3076 121 -3076 0 1
rlabel polysilicon 121 -3082 121 -3082 0 3
rlabel polysilicon 128 -3076 128 -3076 0 1
rlabel polysilicon 128 -3082 128 -3082 0 3
rlabel polysilicon 135 -3082 135 -3082 0 3
rlabel polysilicon 145 -3076 145 -3076 0 2
rlabel polysilicon 142 -3082 142 -3082 0 3
rlabel polysilicon 145 -3082 145 -3082 0 4
rlabel polysilicon 149 -3076 149 -3076 0 1
rlabel polysilicon 152 -3076 152 -3076 0 2
rlabel polysilicon 149 -3082 149 -3082 0 3
rlabel polysilicon 152 -3082 152 -3082 0 4
rlabel polysilicon 156 -3076 156 -3076 0 1
rlabel polysilicon 156 -3082 156 -3082 0 3
rlabel polysilicon 163 -3076 163 -3076 0 1
rlabel polysilicon 163 -3082 163 -3082 0 3
rlabel polysilicon 170 -3076 170 -3076 0 1
rlabel polysilicon 170 -3082 170 -3082 0 3
rlabel polysilicon 177 -3076 177 -3076 0 1
rlabel polysilicon 177 -3082 177 -3082 0 3
rlabel polysilicon 184 -3076 184 -3076 0 1
rlabel polysilicon 187 -3076 187 -3076 0 2
rlabel polysilicon 184 -3082 184 -3082 0 3
rlabel polysilicon 191 -3076 191 -3076 0 1
rlabel polysilicon 191 -3082 191 -3082 0 3
rlabel polysilicon 198 -3082 198 -3082 0 3
rlabel polysilicon 201 -3082 201 -3082 0 4
rlabel polysilicon 205 -3076 205 -3076 0 1
rlabel polysilicon 208 -3076 208 -3076 0 2
rlabel polysilicon 215 -3082 215 -3082 0 4
rlabel polysilicon 219 -3076 219 -3076 0 1
rlabel polysilicon 219 -3082 219 -3082 0 3
rlabel polysilicon 226 -3076 226 -3076 0 1
rlabel polysilicon 226 -3082 226 -3082 0 3
rlabel polysilicon 233 -3076 233 -3076 0 1
rlabel polysilicon 233 -3082 233 -3082 0 3
rlabel polysilicon 240 -3076 240 -3076 0 1
rlabel polysilicon 240 -3082 240 -3082 0 3
rlabel polysilicon 247 -3076 247 -3076 0 1
rlabel polysilicon 247 -3082 247 -3082 0 3
rlabel polysilicon 254 -3076 254 -3076 0 1
rlabel polysilicon 254 -3082 254 -3082 0 3
rlabel polysilicon 261 -3076 261 -3076 0 1
rlabel polysilicon 261 -3082 261 -3082 0 3
rlabel polysilicon 268 -3076 268 -3076 0 1
rlabel polysilicon 268 -3082 268 -3082 0 3
rlabel polysilicon 275 -3076 275 -3076 0 1
rlabel polysilicon 275 -3082 275 -3082 0 3
rlabel polysilicon 282 -3076 282 -3076 0 1
rlabel polysilicon 282 -3082 282 -3082 0 3
rlabel polysilicon 289 -3076 289 -3076 0 1
rlabel polysilicon 289 -3082 289 -3082 0 3
rlabel polysilicon 296 -3076 296 -3076 0 1
rlabel polysilicon 296 -3082 296 -3082 0 3
rlabel polysilicon 303 -3076 303 -3076 0 1
rlabel polysilicon 303 -3082 303 -3082 0 3
rlabel polysilicon 310 -3076 310 -3076 0 1
rlabel polysilicon 310 -3082 310 -3082 0 3
rlabel polysilicon 317 -3076 317 -3076 0 1
rlabel polysilicon 317 -3082 317 -3082 0 3
rlabel polysilicon 324 -3076 324 -3076 0 1
rlabel polysilicon 324 -3082 324 -3082 0 3
rlabel polysilicon 331 -3076 331 -3076 0 1
rlabel polysilicon 331 -3082 331 -3082 0 3
rlabel polysilicon 338 -3076 338 -3076 0 1
rlabel polysilicon 338 -3082 338 -3082 0 3
rlabel polysilicon 345 -3076 345 -3076 0 1
rlabel polysilicon 348 -3082 348 -3082 0 4
rlabel polysilicon 352 -3076 352 -3076 0 1
rlabel polysilicon 352 -3082 352 -3082 0 3
rlabel polysilicon 359 -3076 359 -3076 0 1
rlabel polysilicon 359 -3082 359 -3082 0 3
rlabel polysilicon 366 -3076 366 -3076 0 1
rlabel polysilicon 369 -3076 369 -3076 0 2
rlabel polysilicon 366 -3082 366 -3082 0 3
rlabel polysilicon 369 -3082 369 -3082 0 4
rlabel polysilicon 373 -3076 373 -3076 0 1
rlabel polysilicon 373 -3082 373 -3082 0 3
rlabel polysilicon 380 -3076 380 -3076 0 1
rlabel polysilicon 380 -3082 380 -3082 0 3
rlabel polysilicon 387 -3076 387 -3076 0 1
rlabel polysilicon 387 -3082 387 -3082 0 3
rlabel polysilicon 394 -3076 394 -3076 0 1
rlabel polysilicon 394 -3082 394 -3082 0 3
rlabel polysilicon 401 -3076 401 -3076 0 1
rlabel polysilicon 401 -3082 401 -3082 0 3
rlabel polysilicon 408 -3076 408 -3076 0 1
rlabel polysilicon 408 -3082 408 -3082 0 3
rlabel polysilicon 415 -3076 415 -3076 0 1
rlabel polysilicon 415 -3082 415 -3082 0 3
rlabel polysilicon 422 -3076 422 -3076 0 1
rlabel polysilicon 422 -3082 422 -3082 0 3
rlabel polysilicon 429 -3076 429 -3076 0 1
rlabel polysilicon 429 -3082 429 -3082 0 3
rlabel polysilicon 436 -3076 436 -3076 0 1
rlabel polysilicon 436 -3082 436 -3082 0 3
rlabel polysilicon 443 -3076 443 -3076 0 1
rlabel polysilicon 443 -3082 443 -3082 0 3
rlabel polysilicon 450 -3076 450 -3076 0 1
rlabel polysilicon 453 -3076 453 -3076 0 2
rlabel polysilicon 450 -3082 450 -3082 0 3
rlabel polysilicon 453 -3082 453 -3082 0 4
rlabel polysilicon 457 -3076 457 -3076 0 1
rlabel polysilicon 457 -3082 457 -3082 0 3
rlabel polysilicon 464 -3076 464 -3076 0 1
rlabel polysilicon 464 -3082 464 -3082 0 3
rlabel polysilicon 471 -3076 471 -3076 0 1
rlabel polysilicon 471 -3082 471 -3082 0 3
rlabel polysilicon 478 -3076 478 -3076 0 1
rlabel polysilicon 478 -3082 478 -3082 0 3
rlabel polysilicon 485 -3076 485 -3076 0 1
rlabel polysilicon 485 -3082 485 -3082 0 3
rlabel polysilicon 492 -3076 492 -3076 0 1
rlabel polysilicon 492 -3082 492 -3082 0 3
rlabel polysilicon 499 -3076 499 -3076 0 1
rlabel polysilicon 499 -3082 499 -3082 0 3
rlabel polysilicon 506 -3076 506 -3076 0 1
rlabel polysilicon 506 -3082 506 -3082 0 3
rlabel polysilicon 513 -3076 513 -3076 0 1
rlabel polysilicon 513 -3082 513 -3082 0 3
rlabel polysilicon 520 -3076 520 -3076 0 1
rlabel polysilicon 520 -3082 520 -3082 0 3
rlabel polysilicon 527 -3076 527 -3076 0 1
rlabel polysilicon 527 -3082 527 -3082 0 3
rlabel polysilicon 534 -3076 534 -3076 0 1
rlabel polysilicon 534 -3082 534 -3082 0 3
rlabel polysilicon 541 -3076 541 -3076 0 1
rlabel polysilicon 541 -3082 541 -3082 0 3
rlabel polysilicon 548 -3076 548 -3076 0 1
rlabel polysilicon 548 -3082 548 -3082 0 3
rlabel polysilicon 555 -3076 555 -3076 0 1
rlabel polysilicon 555 -3082 555 -3082 0 3
rlabel polysilicon 562 -3076 562 -3076 0 1
rlabel polysilicon 562 -3082 562 -3082 0 3
rlabel polysilicon 569 -3076 569 -3076 0 1
rlabel polysilicon 569 -3082 569 -3082 0 3
rlabel polysilicon 576 -3076 576 -3076 0 1
rlabel polysilicon 576 -3082 576 -3082 0 3
rlabel polysilicon 583 -3076 583 -3076 0 1
rlabel polysilicon 583 -3082 583 -3082 0 3
rlabel polysilicon 590 -3076 590 -3076 0 1
rlabel polysilicon 590 -3082 590 -3082 0 3
rlabel polysilicon 597 -3076 597 -3076 0 1
rlabel polysilicon 597 -3082 597 -3082 0 3
rlabel polysilicon 604 -3076 604 -3076 0 1
rlabel polysilicon 604 -3082 604 -3082 0 3
rlabel polysilicon 611 -3076 611 -3076 0 1
rlabel polysilicon 611 -3082 611 -3082 0 3
rlabel polysilicon 618 -3076 618 -3076 0 1
rlabel polysilicon 621 -3076 621 -3076 0 2
rlabel polysilicon 621 -3082 621 -3082 0 4
rlabel polysilicon 625 -3076 625 -3076 0 1
rlabel polysilicon 625 -3082 625 -3082 0 3
rlabel polysilicon 632 -3076 632 -3076 0 1
rlabel polysilicon 635 -3076 635 -3076 0 2
rlabel polysilicon 632 -3082 632 -3082 0 3
rlabel polysilicon 635 -3082 635 -3082 0 4
rlabel polysilicon 639 -3076 639 -3076 0 1
rlabel polysilicon 639 -3082 639 -3082 0 3
rlabel polysilicon 646 -3076 646 -3076 0 1
rlabel polysilicon 646 -3082 646 -3082 0 3
rlabel polysilicon 653 -3076 653 -3076 0 1
rlabel polysilicon 653 -3082 653 -3082 0 3
rlabel polysilicon 660 -3076 660 -3076 0 1
rlabel polysilicon 660 -3082 660 -3082 0 3
rlabel polysilicon 667 -3076 667 -3076 0 1
rlabel polysilicon 667 -3082 667 -3082 0 3
rlabel polysilicon 674 -3076 674 -3076 0 1
rlabel polysilicon 674 -3082 674 -3082 0 3
rlabel polysilicon 681 -3076 681 -3076 0 1
rlabel polysilicon 681 -3082 681 -3082 0 3
rlabel polysilicon 688 -3076 688 -3076 0 1
rlabel polysilicon 691 -3076 691 -3076 0 2
rlabel polysilicon 688 -3082 688 -3082 0 3
rlabel polysilicon 691 -3082 691 -3082 0 4
rlabel polysilicon 695 -3076 695 -3076 0 1
rlabel polysilicon 695 -3082 695 -3082 0 3
rlabel polysilicon 702 -3076 702 -3076 0 1
rlabel polysilicon 702 -3082 702 -3082 0 3
rlabel polysilicon 709 -3076 709 -3076 0 1
rlabel polysilicon 709 -3082 709 -3082 0 3
rlabel polysilicon 716 -3076 716 -3076 0 1
rlabel polysilicon 716 -3082 716 -3082 0 3
rlabel polysilicon 723 -3076 723 -3076 0 1
rlabel polysilicon 723 -3082 723 -3082 0 3
rlabel polysilicon 730 -3076 730 -3076 0 1
rlabel polysilicon 730 -3082 730 -3082 0 3
rlabel polysilicon 737 -3076 737 -3076 0 1
rlabel polysilicon 740 -3076 740 -3076 0 2
rlabel polysilicon 737 -3082 737 -3082 0 3
rlabel polysilicon 740 -3082 740 -3082 0 4
rlabel polysilicon 744 -3076 744 -3076 0 1
rlabel polysilicon 744 -3082 744 -3082 0 3
rlabel polysilicon 751 -3076 751 -3076 0 1
rlabel polysilicon 751 -3082 751 -3082 0 3
rlabel polysilicon 758 -3076 758 -3076 0 1
rlabel polysilicon 761 -3082 761 -3082 0 4
rlabel polysilicon 765 -3076 765 -3076 0 1
rlabel polysilicon 765 -3082 765 -3082 0 3
rlabel polysilicon 772 -3076 772 -3076 0 1
rlabel polysilicon 772 -3082 772 -3082 0 3
rlabel polysilicon 779 -3076 779 -3076 0 1
rlabel polysilicon 779 -3082 779 -3082 0 3
rlabel polysilicon 786 -3076 786 -3076 0 1
rlabel polysilicon 789 -3076 789 -3076 0 2
rlabel polysilicon 786 -3082 786 -3082 0 3
rlabel polysilicon 789 -3082 789 -3082 0 4
rlabel polysilicon 793 -3076 793 -3076 0 1
rlabel polysilicon 793 -3082 793 -3082 0 3
rlabel polysilicon 800 -3076 800 -3076 0 1
rlabel polysilicon 800 -3082 800 -3082 0 3
rlabel polysilicon 803 -3082 803 -3082 0 4
rlabel polysilicon 807 -3076 807 -3076 0 1
rlabel polysilicon 807 -3082 807 -3082 0 3
rlabel polysilicon 814 -3076 814 -3076 0 1
rlabel polysilicon 814 -3082 814 -3082 0 3
rlabel polysilicon 821 -3076 821 -3076 0 1
rlabel polysilicon 821 -3082 821 -3082 0 3
rlabel polysilicon 828 -3076 828 -3076 0 1
rlabel polysilicon 831 -3076 831 -3076 0 2
rlabel polysilicon 828 -3082 828 -3082 0 3
rlabel polysilicon 835 -3076 835 -3076 0 1
rlabel polysilicon 835 -3082 835 -3082 0 3
rlabel polysilicon 838 -3082 838 -3082 0 4
rlabel polysilicon 842 -3076 842 -3076 0 1
rlabel polysilicon 842 -3082 842 -3082 0 3
rlabel polysilicon 849 -3076 849 -3076 0 1
rlabel polysilicon 849 -3082 849 -3082 0 3
rlabel polysilicon 856 -3076 856 -3076 0 1
rlabel polysilicon 856 -3082 856 -3082 0 3
rlabel polysilicon 863 -3076 863 -3076 0 1
rlabel polysilicon 863 -3082 863 -3082 0 3
rlabel polysilicon 870 -3076 870 -3076 0 1
rlabel polysilicon 870 -3082 870 -3082 0 3
rlabel polysilicon 877 -3076 877 -3076 0 1
rlabel polysilicon 880 -3076 880 -3076 0 2
rlabel polysilicon 877 -3082 877 -3082 0 3
rlabel polysilicon 884 -3076 884 -3076 0 1
rlabel polysilicon 884 -3082 884 -3082 0 3
rlabel polysilicon 891 -3076 891 -3076 0 1
rlabel polysilicon 891 -3082 891 -3082 0 3
rlabel polysilicon 898 -3076 898 -3076 0 1
rlabel polysilicon 901 -3076 901 -3076 0 2
rlabel polysilicon 898 -3082 898 -3082 0 3
rlabel polysilicon 905 -3076 905 -3076 0 1
rlabel polysilicon 905 -3082 905 -3082 0 3
rlabel polysilicon 915 -3076 915 -3076 0 2
rlabel polysilicon 912 -3082 912 -3082 0 3
rlabel polysilicon 915 -3082 915 -3082 0 4
rlabel polysilicon 919 -3076 919 -3076 0 1
rlabel polysilicon 919 -3082 919 -3082 0 3
rlabel polysilicon 926 -3076 926 -3076 0 1
rlabel polysilicon 926 -3082 926 -3082 0 3
rlabel polysilicon 933 -3076 933 -3076 0 1
rlabel polysilicon 933 -3082 933 -3082 0 3
rlabel polysilicon 940 -3076 940 -3076 0 1
rlabel polysilicon 940 -3082 940 -3082 0 3
rlabel polysilicon 947 -3076 947 -3076 0 1
rlabel polysilicon 947 -3082 947 -3082 0 3
rlabel polysilicon 950 -3082 950 -3082 0 4
rlabel polysilicon 954 -3076 954 -3076 0 1
rlabel polysilicon 954 -3082 954 -3082 0 3
rlabel polysilicon 961 -3076 961 -3076 0 1
rlabel polysilicon 961 -3082 961 -3082 0 3
rlabel polysilicon 968 -3076 968 -3076 0 1
rlabel polysilicon 968 -3082 968 -3082 0 3
rlabel polysilicon 978 -3076 978 -3076 0 2
rlabel polysilicon 975 -3082 975 -3082 0 3
rlabel polysilicon 978 -3082 978 -3082 0 4
rlabel polysilicon 982 -3076 982 -3076 0 1
rlabel polysilicon 982 -3082 982 -3082 0 3
rlabel polysilicon 989 -3076 989 -3076 0 1
rlabel polysilicon 989 -3082 989 -3082 0 3
rlabel polysilicon 996 -3076 996 -3076 0 1
rlabel polysilicon 996 -3082 996 -3082 0 3
rlabel polysilicon 1003 -3076 1003 -3076 0 1
rlabel polysilicon 1003 -3082 1003 -3082 0 3
rlabel polysilicon 1010 -3076 1010 -3076 0 1
rlabel polysilicon 1010 -3082 1010 -3082 0 3
rlabel polysilicon 1017 -3076 1017 -3076 0 1
rlabel polysilicon 1020 -3076 1020 -3076 0 2
rlabel polysilicon 1017 -3082 1017 -3082 0 3
rlabel polysilicon 1020 -3082 1020 -3082 0 4
rlabel polysilicon 1024 -3076 1024 -3076 0 1
rlabel polysilicon 1024 -3082 1024 -3082 0 3
rlabel polysilicon 1031 -3076 1031 -3076 0 1
rlabel polysilicon 1031 -3082 1031 -3082 0 3
rlabel polysilicon 1038 -3076 1038 -3076 0 1
rlabel polysilicon 1038 -3082 1038 -3082 0 3
rlabel polysilicon 1045 -3076 1045 -3076 0 1
rlabel polysilicon 1045 -3082 1045 -3082 0 3
rlabel polysilicon 1052 -3076 1052 -3076 0 1
rlabel polysilicon 1052 -3082 1052 -3082 0 3
rlabel polysilicon 1059 -3076 1059 -3076 0 1
rlabel polysilicon 1059 -3082 1059 -3082 0 3
rlabel polysilicon 1066 -3076 1066 -3076 0 1
rlabel polysilicon 1066 -3082 1066 -3082 0 3
rlabel polysilicon 1073 -3076 1073 -3076 0 1
rlabel polysilicon 1073 -3082 1073 -3082 0 3
rlabel polysilicon 1080 -3076 1080 -3076 0 1
rlabel polysilicon 1080 -3082 1080 -3082 0 3
rlabel polysilicon 1083 -3082 1083 -3082 0 4
rlabel polysilicon 1087 -3082 1087 -3082 0 3
rlabel polysilicon 1090 -3082 1090 -3082 0 4
rlabel polysilicon 1094 -3076 1094 -3076 0 1
rlabel polysilicon 1094 -3082 1094 -3082 0 3
rlabel polysilicon 1101 -3076 1101 -3076 0 1
rlabel polysilicon 1101 -3082 1101 -3082 0 3
rlabel polysilicon 1108 -3076 1108 -3076 0 1
rlabel polysilicon 1108 -3082 1108 -3082 0 3
rlabel polysilicon 1115 -3076 1115 -3076 0 1
rlabel polysilicon 1115 -3082 1115 -3082 0 3
rlabel polysilicon 1122 -3076 1122 -3076 0 1
rlabel polysilicon 1122 -3082 1122 -3082 0 3
rlabel polysilicon 1129 -3076 1129 -3076 0 1
rlabel polysilicon 1129 -3082 1129 -3082 0 3
rlabel polysilicon 1136 -3076 1136 -3076 0 1
rlabel polysilicon 1136 -3082 1136 -3082 0 3
rlabel polysilicon 1143 -3076 1143 -3076 0 1
rlabel polysilicon 1143 -3082 1143 -3082 0 3
rlabel polysilicon 1150 -3076 1150 -3076 0 1
rlabel polysilicon 1150 -3082 1150 -3082 0 3
rlabel polysilicon 1157 -3076 1157 -3076 0 1
rlabel polysilicon 1157 -3082 1157 -3082 0 3
rlabel polysilicon 1164 -3076 1164 -3076 0 1
rlabel polysilicon 1164 -3082 1164 -3082 0 3
rlabel polysilicon 1171 -3076 1171 -3076 0 1
rlabel polysilicon 1171 -3082 1171 -3082 0 3
rlabel polysilicon 1178 -3076 1178 -3076 0 1
rlabel polysilicon 1178 -3082 1178 -3082 0 3
rlabel polysilicon 1185 -3076 1185 -3076 0 1
rlabel polysilicon 1185 -3082 1185 -3082 0 3
rlabel polysilicon 1192 -3076 1192 -3076 0 1
rlabel polysilicon 1192 -3082 1192 -3082 0 3
rlabel polysilicon 1199 -3076 1199 -3076 0 1
rlabel polysilicon 1199 -3082 1199 -3082 0 3
rlabel polysilicon 1206 -3076 1206 -3076 0 1
rlabel polysilicon 1206 -3082 1206 -3082 0 3
rlabel polysilicon 1213 -3076 1213 -3076 0 1
rlabel polysilicon 1213 -3082 1213 -3082 0 3
rlabel polysilicon 1220 -3076 1220 -3076 0 1
rlabel polysilicon 1220 -3082 1220 -3082 0 3
rlabel polysilicon 1227 -3076 1227 -3076 0 1
rlabel polysilicon 1227 -3082 1227 -3082 0 3
rlabel polysilicon 1234 -3076 1234 -3076 0 1
rlabel polysilicon 1234 -3082 1234 -3082 0 3
rlabel polysilicon 1241 -3076 1241 -3076 0 1
rlabel polysilicon 1241 -3082 1241 -3082 0 3
rlabel polysilicon 1248 -3076 1248 -3076 0 1
rlabel polysilicon 1248 -3082 1248 -3082 0 3
rlabel polysilicon 1255 -3076 1255 -3076 0 1
rlabel polysilicon 1255 -3082 1255 -3082 0 3
rlabel polysilicon 1262 -3076 1262 -3076 0 1
rlabel polysilicon 1262 -3082 1262 -3082 0 3
rlabel polysilicon 1269 -3076 1269 -3076 0 1
rlabel polysilicon 1269 -3082 1269 -3082 0 3
rlabel polysilicon 1276 -3076 1276 -3076 0 1
rlabel polysilicon 1276 -3082 1276 -3082 0 3
rlabel polysilicon 1283 -3076 1283 -3076 0 1
rlabel polysilicon 1283 -3082 1283 -3082 0 3
rlabel polysilicon 1290 -3076 1290 -3076 0 1
rlabel polysilicon 1290 -3082 1290 -3082 0 3
rlabel polysilicon 1297 -3076 1297 -3076 0 1
rlabel polysilicon 1297 -3082 1297 -3082 0 3
rlabel polysilicon 1304 -3076 1304 -3076 0 1
rlabel polysilicon 1304 -3082 1304 -3082 0 3
rlabel polysilicon 1311 -3076 1311 -3076 0 1
rlabel polysilicon 1311 -3082 1311 -3082 0 3
rlabel polysilicon 1318 -3076 1318 -3076 0 1
rlabel polysilicon 1318 -3082 1318 -3082 0 3
rlabel polysilicon 1325 -3076 1325 -3076 0 1
rlabel polysilicon 1325 -3082 1325 -3082 0 3
rlabel polysilicon 1332 -3076 1332 -3076 0 1
rlabel polysilicon 1332 -3082 1332 -3082 0 3
rlabel polysilicon 1339 -3076 1339 -3076 0 1
rlabel polysilicon 1339 -3082 1339 -3082 0 3
rlabel polysilicon 1346 -3076 1346 -3076 0 1
rlabel polysilicon 1346 -3082 1346 -3082 0 3
rlabel polysilicon 1353 -3076 1353 -3076 0 1
rlabel polysilicon 1353 -3082 1353 -3082 0 3
rlabel polysilicon 1360 -3076 1360 -3076 0 1
rlabel polysilicon 1360 -3082 1360 -3082 0 3
rlabel polysilicon 1367 -3076 1367 -3076 0 1
rlabel polysilicon 1367 -3082 1367 -3082 0 3
rlabel polysilicon 1374 -3076 1374 -3076 0 1
rlabel polysilicon 1374 -3082 1374 -3082 0 3
rlabel polysilicon 1381 -3076 1381 -3076 0 1
rlabel polysilicon 1381 -3082 1381 -3082 0 3
rlabel polysilicon 1388 -3076 1388 -3076 0 1
rlabel polysilicon 1388 -3082 1388 -3082 0 3
rlabel polysilicon 1395 -3076 1395 -3076 0 1
rlabel polysilicon 1395 -3082 1395 -3082 0 3
rlabel polysilicon 1402 -3076 1402 -3076 0 1
rlabel polysilicon 1402 -3082 1402 -3082 0 3
rlabel polysilicon 1409 -3076 1409 -3076 0 1
rlabel polysilicon 1409 -3082 1409 -3082 0 3
rlabel polysilicon 1416 -3076 1416 -3076 0 1
rlabel polysilicon 1416 -3082 1416 -3082 0 3
rlabel polysilicon 1423 -3076 1423 -3076 0 1
rlabel polysilicon 1423 -3082 1423 -3082 0 3
rlabel polysilicon 1430 -3076 1430 -3076 0 1
rlabel polysilicon 1430 -3082 1430 -3082 0 3
rlabel polysilicon 1437 -3076 1437 -3076 0 1
rlabel polysilicon 1437 -3082 1437 -3082 0 3
rlabel polysilicon 1444 -3076 1444 -3076 0 1
rlabel polysilicon 1444 -3082 1444 -3082 0 3
rlabel polysilicon 1451 -3076 1451 -3076 0 1
rlabel polysilicon 1451 -3082 1451 -3082 0 3
rlabel polysilicon 1458 -3076 1458 -3076 0 1
rlabel polysilicon 1458 -3082 1458 -3082 0 3
rlabel polysilicon 1465 -3076 1465 -3076 0 1
rlabel polysilicon 1465 -3082 1465 -3082 0 3
rlabel polysilicon 1472 -3076 1472 -3076 0 1
rlabel polysilicon 1472 -3082 1472 -3082 0 3
rlabel polysilicon 1479 -3076 1479 -3076 0 1
rlabel polysilicon 1479 -3082 1479 -3082 0 3
rlabel polysilicon 1486 -3076 1486 -3076 0 1
rlabel polysilicon 1486 -3082 1486 -3082 0 3
rlabel polysilicon 1493 -3076 1493 -3076 0 1
rlabel polysilicon 1493 -3082 1493 -3082 0 3
rlabel polysilicon 1500 -3076 1500 -3076 0 1
rlabel polysilicon 1500 -3082 1500 -3082 0 3
rlabel polysilicon 1507 -3076 1507 -3076 0 1
rlabel polysilicon 1507 -3082 1507 -3082 0 3
rlabel polysilicon 1514 -3076 1514 -3076 0 1
rlabel polysilicon 1514 -3082 1514 -3082 0 3
rlabel polysilicon 1521 -3076 1521 -3076 0 1
rlabel polysilicon 1521 -3082 1521 -3082 0 3
rlabel polysilicon 1528 -3076 1528 -3076 0 1
rlabel polysilicon 1528 -3082 1528 -3082 0 3
rlabel polysilicon 1535 -3076 1535 -3076 0 1
rlabel polysilicon 1535 -3082 1535 -3082 0 3
rlabel polysilicon 1542 -3076 1542 -3076 0 1
rlabel polysilicon 1542 -3082 1542 -3082 0 3
rlabel polysilicon 1549 -3076 1549 -3076 0 1
rlabel polysilicon 1549 -3082 1549 -3082 0 3
rlabel polysilicon 1556 -3076 1556 -3076 0 1
rlabel polysilicon 1556 -3082 1556 -3082 0 3
rlabel polysilicon 1563 -3076 1563 -3076 0 1
rlabel polysilicon 1563 -3082 1563 -3082 0 3
rlabel polysilicon 1570 -3076 1570 -3076 0 1
rlabel polysilicon 1570 -3082 1570 -3082 0 3
rlabel polysilicon 1577 -3076 1577 -3076 0 1
rlabel polysilicon 1577 -3082 1577 -3082 0 3
rlabel polysilicon 1584 -3076 1584 -3076 0 1
rlabel polysilicon 1584 -3082 1584 -3082 0 3
rlabel polysilicon 1591 -3076 1591 -3076 0 1
rlabel polysilicon 1591 -3082 1591 -3082 0 3
rlabel polysilicon 1598 -3076 1598 -3076 0 1
rlabel polysilicon 1598 -3082 1598 -3082 0 3
rlabel polysilicon 1605 -3076 1605 -3076 0 1
rlabel polysilicon 1605 -3082 1605 -3082 0 3
rlabel polysilicon 1612 -3076 1612 -3076 0 1
rlabel polysilicon 1612 -3082 1612 -3082 0 3
rlabel polysilicon 1619 -3076 1619 -3076 0 1
rlabel polysilicon 1619 -3082 1619 -3082 0 3
rlabel polysilicon 1626 -3076 1626 -3076 0 1
rlabel polysilicon 1626 -3082 1626 -3082 0 3
rlabel polysilicon 1633 -3076 1633 -3076 0 1
rlabel polysilicon 1633 -3082 1633 -3082 0 3
rlabel polysilicon 1640 -3076 1640 -3076 0 1
rlabel polysilicon 1640 -3082 1640 -3082 0 3
rlabel polysilicon 1647 -3076 1647 -3076 0 1
rlabel polysilicon 1647 -3082 1647 -3082 0 3
rlabel polysilicon 1654 -3076 1654 -3076 0 1
rlabel polysilicon 1654 -3082 1654 -3082 0 3
rlabel polysilicon 65 -3221 65 -3221 0 3
rlabel polysilicon 72 -3215 72 -3215 0 1
rlabel polysilicon 72 -3221 72 -3221 0 3
rlabel polysilicon 79 -3215 79 -3215 0 1
rlabel polysilicon 79 -3221 79 -3221 0 3
rlabel polysilicon 86 -3215 86 -3215 0 1
rlabel polysilicon 86 -3221 86 -3221 0 3
rlabel polysilicon 93 -3215 93 -3215 0 1
rlabel polysilicon 93 -3221 93 -3221 0 3
rlabel polysilicon 100 -3215 100 -3215 0 1
rlabel polysilicon 100 -3221 100 -3221 0 3
rlabel polysilicon 107 -3215 107 -3215 0 1
rlabel polysilicon 107 -3221 107 -3221 0 3
rlabel polysilicon 114 -3215 114 -3215 0 1
rlabel polysilicon 117 -3215 117 -3215 0 2
rlabel polysilicon 114 -3221 114 -3221 0 3
rlabel polysilicon 121 -3215 121 -3215 0 1
rlabel polysilicon 121 -3221 121 -3221 0 3
rlabel polysilicon 128 -3215 128 -3215 0 1
rlabel polysilicon 131 -3215 131 -3215 0 2
rlabel polysilicon 128 -3221 128 -3221 0 3
rlabel polysilicon 135 -3215 135 -3215 0 1
rlabel polysilicon 135 -3221 135 -3221 0 3
rlabel polysilicon 142 -3215 142 -3215 0 1
rlabel polysilicon 142 -3221 142 -3221 0 3
rlabel polysilicon 149 -3215 149 -3215 0 1
rlabel polysilicon 152 -3215 152 -3215 0 2
rlabel polysilicon 149 -3221 149 -3221 0 3
rlabel polysilicon 152 -3221 152 -3221 0 4
rlabel polysilicon 156 -3215 156 -3215 0 1
rlabel polysilicon 156 -3221 156 -3221 0 3
rlabel polysilicon 163 -3215 163 -3215 0 1
rlabel polysilicon 163 -3221 163 -3221 0 3
rlabel polysilicon 170 -3215 170 -3215 0 1
rlabel polysilicon 170 -3221 170 -3221 0 3
rlabel polysilicon 177 -3215 177 -3215 0 1
rlabel polysilicon 177 -3221 177 -3221 0 3
rlabel polysilicon 184 -3215 184 -3215 0 1
rlabel polysilicon 184 -3221 184 -3221 0 3
rlabel polysilicon 191 -3215 191 -3215 0 1
rlabel polysilicon 191 -3221 191 -3221 0 3
rlabel polysilicon 198 -3215 198 -3215 0 1
rlabel polysilicon 198 -3221 198 -3221 0 3
rlabel polysilicon 205 -3215 205 -3215 0 1
rlabel polysilicon 205 -3221 205 -3221 0 3
rlabel polysilicon 212 -3215 212 -3215 0 1
rlabel polysilicon 212 -3221 212 -3221 0 3
rlabel polysilicon 219 -3215 219 -3215 0 1
rlabel polysilicon 219 -3221 219 -3221 0 3
rlabel polysilicon 226 -3215 226 -3215 0 1
rlabel polysilicon 226 -3221 226 -3221 0 3
rlabel polysilicon 233 -3215 233 -3215 0 1
rlabel polysilicon 233 -3221 233 -3221 0 3
rlabel polysilicon 243 -3221 243 -3221 0 4
rlabel polysilicon 247 -3215 247 -3215 0 1
rlabel polysilicon 247 -3221 247 -3221 0 3
rlabel polysilicon 254 -3215 254 -3215 0 1
rlabel polysilicon 254 -3221 254 -3221 0 3
rlabel polysilicon 261 -3215 261 -3215 0 1
rlabel polysilicon 261 -3221 261 -3221 0 3
rlabel polysilicon 268 -3215 268 -3215 0 1
rlabel polysilicon 268 -3221 268 -3221 0 3
rlabel polysilicon 275 -3215 275 -3215 0 1
rlabel polysilicon 275 -3221 275 -3221 0 3
rlabel polysilicon 282 -3215 282 -3215 0 1
rlabel polysilicon 282 -3221 282 -3221 0 3
rlabel polysilicon 289 -3215 289 -3215 0 1
rlabel polysilicon 289 -3221 289 -3221 0 3
rlabel polysilicon 296 -3215 296 -3215 0 1
rlabel polysilicon 296 -3221 296 -3221 0 3
rlabel polysilicon 303 -3215 303 -3215 0 1
rlabel polysilicon 303 -3221 303 -3221 0 3
rlabel polysilicon 310 -3215 310 -3215 0 1
rlabel polysilicon 310 -3221 310 -3221 0 3
rlabel polysilicon 317 -3215 317 -3215 0 1
rlabel polysilicon 317 -3221 317 -3221 0 3
rlabel polysilicon 324 -3215 324 -3215 0 1
rlabel polysilicon 324 -3221 324 -3221 0 3
rlabel polysilicon 331 -3215 331 -3215 0 1
rlabel polysilicon 331 -3221 331 -3221 0 3
rlabel polysilicon 338 -3215 338 -3215 0 1
rlabel polysilicon 338 -3221 338 -3221 0 3
rlabel polysilicon 345 -3215 345 -3215 0 1
rlabel polysilicon 345 -3221 345 -3221 0 3
rlabel polysilicon 352 -3215 352 -3215 0 1
rlabel polysilicon 352 -3221 352 -3221 0 3
rlabel polysilicon 359 -3215 359 -3215 0 1
rlabel polysilicon 359 -3221 359 -3221 0 3
rlabel polysilicon 366 -3215 366 -3215 0 1
rlabel polysilicon 366 -3221 366 -3221 0 3
rlabel polysilicon 373 -3215 373 -3215 0 1
rlabel polysilicon 373 -3221 373 -3221 0 3
rlabel polysilicon 380 -3215 380 -3215 0 1
rlabel polysilicon 380 -3221 380 -3221 0 3
rlabel polysilicon 387 -3215 387 -3215 0 1
rlabel polysilicon 387 -3221 387 -3221 0 3
rlabel polysilicon 394 -3215 394 -3215 0 1
rlabel polysilicon 394 -3221 394 -3221 0 3
rlabel polysilicon 401 -3215 401 -3215 0 1
rlabel polysilicon 404 -3215 404 -3215 0 2
rlabel polysilicon 401 -3221 401 -3221 0 3
rlabel polysilicon 404 -3221 404 -3221 0 4
rlabel polysilicon 408 -3215 408 -3215 0 1
rlabel polysilicon 408 -3221 408 -3221 0 3
rlabel polysilicon 415 -3215 415 -3215 0 1
rlabel polysilicon 415 -3221 415 -3221 0 3
rlabel polysilicon 422 -3215 422 -3215 0 1
rlabel polysilicon 422 -3221 422 -3221 0 3
rlabel polysilicon 429 -3215 429 -3215 0 1
rlabel polysilicon 432 -3215 432 -3215 0 2
rlabel polysilicon 429 -3221 429 -3221 0 3
rlabel polysilicon 436 -3215 436 -3215 0 1
rlabel polysilicon 436 -3221 436 -3221 0 3
rlabel polysilicon 443 -3215 443 -3215 0 1
rlabel polysilicon 443 -3221 443 -3221 0 3
rlabel polysilicon 450 -3215 450 -3215 0 1
rlabel polysilicon 450 -3221 450 -3221 0 3
rlabel polysilicon 457 -3215 457 -3215 0 1
rlabel polysilicon 457 -3221 457 -3221 0 3
rlabel polysilicon 464 -3215 464 -3215 0 1
rlabel polysilicon 464 -3221 464 -3221 0 3
rlabel polysilicon 471 -3215 471 -3215 0 1
rlabel polysilicon 474 -3215 474 -3215 0 2
rlabel polysilicon 471 -3221 471 -3221 0 3
rlabel polysilicon 478 -3215 478 -3215 0 1
rlabel polysilicon 478 -3221 478 -3221 0 3
rlabel polysilicon 485 -3215 485 -3215 0 1
rlabel polysilicon 485 -3221 485 -3221 0 3
rlabel polysilicon 492 -3215 492 -3215 0 1
rlabel polysilicon 492 -3221 492 -3221 0 3
rlabel polysilicon 495 -3221 495 -3221 0 4
rlabel polysilicon 499 -3215 499 -3215 0 1
rlabel polysilicon 502 -3215 502 -3215 0 2
rlabel polysilicon 499 -3221 499 -3221 0 3
rlabel polysilicon 502 -3221 502 -3221 0 4
rlabel polysilicon 506 -3215 506 -3215 0 1
rlabel polysilicon 506 -3221 506 -3221 0 3
rlabel polysilicon 513 -3215 513 -3215 0 1
rlabel polysilicon 513 -3221 513 -3221 0 3
rlabel polysilicon 520 -3215 520 -3215 0 1
rlabel polysilicon 520 -3221 520 -3221 0 3
rlabel polysilicon 527 -3215 527 -3215 0 1
rlabel polysilicon 527 -3221 527 -3221 0 3
rlabel polysilicon 534 -3215 534 -3215 0 1
rlabel polysilicon 537 -3215 537 -3215 0 2
rlabel polysilicon 534 -3221 534 -3221 0 3
rlabel polysilicon 541 -3221 541 -3221 0 3
rlabel polysilicon 544 -3221 544 -3221 0 4
rlabel polysilicon 548 -3215 548 -3215 0 1
rlabel polysilicon 548 -3221 548 -3221 0 3
rlabel polysilicon 555 -3215 555 -3215 0 1
rlabel polysilicon 555 -3221 555 -3221 0 3
rlabel polysilicon 562 -3215 562 -3215 0 1
rlabel polysilicon 562 -3221 562 -3221 0 3
rlabel polysilicon 569 -3215 569 -3215 0 1
rlabel polysilicon 569 -3221 569 -3221 0 3
rlabel polysilicon 576 -3215 576 -3215 0 1
rlabel polysilicon 579 -3215 579 -3215 0 2
rlabel polysilicon 576 -3221 576 -3221 0 3
rlabel polysilicon 579 -3221 579 -3221 0 4
rlabel polysilicon 583 -3215 583 -3215 0 1
rlabel polysilicon 583 -3221 583 -3221 0 3
rlabel polysilicon 590 -3215 590 -3215 0 1
rlabel polysilicon 593 -3215 593 -3215 0 2
rlabel polysilicon 593 -3221 593 -3221 0 4
rlabel polysilicon 597 -3215 597 -3215 0 1
rlabel polysilicon 597 -3221 597 -3221 0 3
rlabel polysilicon 604 -3215 604 -3215 0 1
rlabel polysilicon 604 -3221 604 -3221 0 3
rlabel polysilicon 611 -3215 611 -3215 0 1
rlabel polysilicon 611 -3221 611 -3221 0 3
rlabel polysilicon 618 -3215 618 -3215 0 1
rlabel polysilicon 618 -3221 618 -3221 0 3
rlabel polysilicon 625 -3215 625 -3215 0 1
rlabel polysilicon 625 -3221 625 -3221 0 3
rlabel polysilicon 632 -3215 632 -3215 0 1
rlabel polysilicon 632 -3221 632 -3221 0 3
rlabel polysilicon 639 -3215 639 -3215 0 1
rlabel polysilicon 639 -3221 639 -3221 0 3
rlabel polysilicon 646 -3215 646 -3215 0 1
rlabel polysilicon 653 -3215 653 -3215 0 1
rlabel polysilicon 656 -3215 656 -3215 0 2
rlabel polysilicon 656 -3221 656 -3221 0 4
rlabel polysilicon 660 -3215 660 -3215 0 1
rlabel polysilicon 660 -3221 660 -3221 0 3
rlabel polysilicon 667 -3215 667 -3215 0 1
rlabel polysilicon 667 -3221 667 -3221 0 3
rlabel polysilicon 674 -3215 674 -3215 0 1
rlabel polysilicon 674 -3221 674 -3221 0 3
rlabel polysilicon 681 -3215 681 -3215 0 1
rlabel polysilicon 684 -3215 684 -3215 0 2
rlabel polysilicon 681 -3221 681 -3221 0 3
rlabel polysilicon 684 -3221 684 -3221 0 4
rlabel polysilicon 688 -3215 688 -3215 0 1
rlabel polysilicon 688 -3221 688 -3221 0 3
rlabel polysilicon 695 -3215 695 -3215 0 1
rlabel polysilicon 695 -3221 695 -3221 0 3
rlabel polysilicon 702 -3215 702 -3215 0 1
rlabel polysilicon 702 -3221 702 -3221 0 3
rlabel polysilicon 709 -3215 709 -3215 0 1
rlabel polysilicon 709 -3221 709 -3221 0 3
rlabel polysilicon 716 -3215 716 -3215 0 1
rlabel polysilicon 716 -3221 716 -3221 0 3
rlabel polysilicon 723 -3215 723 -3215 0 1
rlabel polysilicon 723 -3221 723 -3221 0 3
rlabel polysilicon 730 -3215 730 -3215 0 1
rlabel polysilicon 730 -3221 730 -3221 0 3
rlabel polysilicon 737 -3215 737 -3215 0 1
rlabel polysilicon 737 -3221 737 -3221 0 3
rlabel polysilicon 744 -3215 744 -3215 0 1
rlabel polysilicon 744 -3221 744 -3221 0 3
rlabel polysilicon 751 -3215 751 -3215 0 1
rlabel polysilicon 751 -3221 751 -3221 0 3
rlabel polysilicon 758 -3215 758 -3215 0 1
rlabel polysilicon 758 -3221 758 -3221 0 3
rlabel polysilicon 765 -3215 765 -3215 0 1
rlabel polysilicon 765 -3221 765 -3221 0 3
rlabel polysilicon 772 -3215 772 -3215 0 1
rlabel polysilicon 772 -3221 772 -3221 0 3
rlabel polysilicon 779 -3215 779 -3215 0 1
rlabel polysilicon 782 -3215 782 -3215 0 2
rlabel polysilicon 779 -3221 779 -3221 0 3
rlabel polysilicon 786 -3215 786 -3215 0 1
rlabel polysilicon 786 -3221 786 -3221 0 3
rlabel polysilicon 793 -3215 793 -3215 0 1
rlabel polysilicon 796 -3215 796 -3215 0 2
rlabel polysilicon 793 -3221 793 -3221 0 3
rlabel polysilicon 796 -3221 796 -3221 0 4
rlabel polysilicon 800 -3215 800 -3215 0 1
rlabel polysilicon 800 -3221 800 -3221 0 3
rlabel polysilicon 807 -3215 807 -3215 0 1
rlabel polysilicon 807 -3221 807 -3221 0 3
rlabel polysilicon 814 -3215 814 -3215 0 1
rlabel polysilicon 814 -3221 814 -3221 0 3
rlabel polysilicon 821 -3215 821 -3215 0 1
rlabel polysilicon 824 -3215 824 -3215 0 2
rlabel polysilicon 821 -3221 821 -3221 0 3
rlabel polysilicon 824 -3221 824 -3221 0 4
rlabel polysilicon 828 -3215 828 -3215 0 1
rlabel polysilicon 828 -3221 828 -3221 0 3
rlabel polysilicon 835 -3215 835 -3215 0 1
rlabel polysilicon 838 -3215 838 -3215 0 2
rlabel polysilicon 835 -3221 835 -3221 0 3
rlabel polysilicon 838 -3221 838 -3221 0 4
rlabel polysilicon 842 -3215 842 -3215 0 1
rlabel polysilicon 842 -3221 842 -3221 0 3
rlabel polysilicon 849 -3215 849 -3215 0 1
rlabel polysilicon 849 -3221 849 -3221 0 3
rlabel polysilicon 856 -3215 856 -3215 0 1
rlabel polysilicon 856 -3221 856 -3221 0 3
rlabel polysilicon 863 -3215 863 -3215 0 1
rlabel polysilicon 863 -3221 863 -3221 0 3
rlabel polysilicon 870 -3215 870 -3215 0 1
rlabel polysilicon 870 -3221 870 -3221 0 3
rlabel polysilicon 877 -3215 877 -3215 0 1
rlabel polysilicon 877 -3221 877 -3221 0 3
rlabel polysilicon 884 -3215 884 -3215 0 1
rlabel polysilicon 884 -3221 884 -3221 0 3
rlabel polysilicon 891 -3221 891 -3221 0 3
rlabel polysilicon 894 -3221 894 -3221 0 4
rlabel polysilicon 898 -3215 898 -3215 0 1
rlabel polysilicon 898 -3221 898 -3221 0 3
rlabel polysilicon 905 -3215 905 -3215 0 1
rlabel polysilicon 905 -3221 905 -3221 0 3
rlabel polysilicon 912 -3215 912 -3215 0 1
rlabel polysilicon 912 -3221 912 -3221 0 3
rlabel polysilicon 919 -3215 919 -3215 0 1
rlabel polysilicon 919 -3221 919 -3221 0 3
rlabel polysilicon 926 -3215 926 -3215 0 1
rlabel polysilicon 926 -3221 926 -3221 0 3
rlabel polysilicon 933 -3215 933 -3215 0 1
rlabel polysilicon 933 -3221 933 -3221 0 3
rlabel polysilicon 940 -3215 940 -3215 0 1
rlabel polysilicon 940 -3221 940 -3221 0 3
rlabel polysilicon 947 -3215 947 -3215 0 1
rlabel polysilicon 947 -3221 947 -3221 0 3
rlabel polysilicon 950 -3221 950 -3221 0 4
rlabel polysilicon 954 -3215 954 -3215 0 1
rlabel polysilicon 954 -3221 954 -3221 0 3
rlabel polysilicon 961 -3215 961 -3215 0 1
rlabel polysilicon 961 -3221 961 -3221 0 3
rlabel polysilicon 968 -3215 968 -3215 0 1
rlabel polysilicon 968 -3221 968 -3221 0 3
rlabel polysilicon 975 -3215 975 -3215 0 1
rlabel polysilicon 975 -3221 975 -3221 0 3
rlabel polysilicon 982 -3215 982 -3215 0 1
rlabel polysilicon 982 -3221 982 -3221 0 3
rlabel polysilicon 989 -3215 989 -3215 0 1
rlabel polysilicon 989 -3221 989 -3221 0 3
rlabel polysilicon 996 -3215 996 -3215 0 1
rlabel polysilicon 999 -3215 999 -3215 0 2
rlabel polysilicon 996 -3221 996 -3221 0 3
rlabel polysilicon 999 -3221 999 -3221 0 4
rlabel polysilicon 1003 -3215 1003 -3215 0 1
rlabel polysilicon 1003 -3221 1003 -3221 0 3
rlabel polysilicon 1013 -3215 1013 -3215 0 2
rlabel polysilicon 1010 -3221 1010 -3221 0 3
rlabel polysilicon 1013 -3221 1013 -3221 0 4
rlabel polysilicon 1017 -3215 1017 -3215 0 1
rlabel polysilicon 1017 -3221 1017 -3221 0 3
rlabel polysilicon 1024 -3215 1024 -3215 0 1
rlabel polysilicon 1024 -3221 1024 -3221 0 3
rlabel polysilicon 1031 -3215 1031 -3215 0 1
rlabel polysilicon 1031 -3221 1031 -3221 0 3
rlabel polysilicon 1038 -3215 1038 -3215 0 1
rlabel polysilicon 1038 -3221 1038 -3221 0 3
rlabel polysilicon 1045 -3215 1045 -3215 0 1
rlabel polysilicon 1045 -3221 1045 -3221 0 3
rlabel polysilicon 1052 -3215 1052 -3215 0 1
rlabel polysilicon 1052 -3221 1052 -3221 0 3
rlabel polysilicon 1059 -3215 1059 -3215 0 1
rlabel polysilicon 1062 -3215 1062 -3215 0 2
rlabel polysilicon 1066 -3215 1066 -3215 0 1
rlabel polysilicon 1066 -3221 1066 -3221 0 3
rlabel polysilicon 1073 -3215 1073 -3215 0 1
rlabel polysilicon 1073 -3221 1073 -3221 0 3
rlabel polysilicon 1080 -3215 1080 -3215 0 1
rlabel polysilicon 1080 -3221 1080 -3221 0 3
rlabel polysilicon 1087 -3215 1087 -3215 0 1
rlabel polysilicon 1090 -3215 1090 -3215 0 2
rlabel polysilicon 1090 -3221 1090 -3221 0 4
rlabel polysilicon 1094 -3215 1094 -3215 0 1
rlabel polysilicon 1094 -3221 1094 -3221 0 3
rlabel polysilicon 1101 -3215 1101 -3215 0 1
rlabel polysilicon 1101 -3221 1101 -3221 0 3
rlabel polysilicon 1108 -3215 1108 -3215 0 1
rlabel polysilicon 1108 -3221 1108 -3221 0 3
rlabel polysilicon 1115 -3215 1115 -3215 0 1
rlabel polysilicon 1115 -3221 1115 -3221 0 3
rlabel polysilicon 1122 -3215 1122 -3215 0 1
rlabel polysilicon 1122 -3221 1122 -3221 0 3
rlabel polysilicon 1129 -3215 1129 -3215 0 1
rlabel polysilicon 1129 -3221 1129 -3221 0 3
rlabel polysilicon 1136 -3215 1136 -3215 0 1
rlabel polysilicon 1136 -3221 1136 -3221 0 3
rlabel polysilicon 1143 -3215 1143 -3215 0 1
rlabel polysilicon 1143 -3221 1143 -3221 0 3
rlabel polysilicon 1150 -3215 1150 -3215 0 1
rlabel polysilicon 1150 -3221 1150 -3221 0 3
rlabel polysilicon 1157 -3215 1157 -3215 0 1
rlabel polysilicon 1157 -3221 1157 -3221 0 3
rlabel polysilicon 1164 -3215 1164 -3215 0 1
rlabel polysilicon 1164 -3221 1164 -3221 0 3
rlabel polysilicon 1171 -3215 1171 -3215 0 1
rlabel polysilicon 1171 -3221 1171 -3221 0 3
rlabel polysilicon 1178 -3215 1178 -3215 0 1
rlabel polysilicon 1178 -3221 1178 -3221 0 3
rlabel polysilicon 1185 -3215 1185 -3215 0 1
rlabel polysilicon 1185 -3221 1185 -3221 0 3
rlabel polysilicon 1192 -3215 1192 -3215 0 1
rlabel polysilicon 1192 -3221 1192 -3221 0 3
rlabel polysilicon 1199 -3215 1199 -3215 0 1
rlabel polysilicon 1199 -3221 1199 -3221 0 3
rlabel polysilicon 1206 -3215 1206 -3215 0 1
rlabel polysilicon 1206 -3221 1206 -3221 0 3
rlabel polysilicon 1213 -3215 1213 -3215 0 1
rlabel polysilicon 1213 -3221 1213 -3221 0 3
rlabel polysilicon 1220 -3215 1220 -3215 0 1
rlabel polysilicon 1220 -3221 1220 -3221 0 3
rlabel polysilicon 1227 -3215 1227 -3215 0 1
rlabel polysilicon 1227 -3221 1227 -3221 0 3
rlabel polysilicon 1234 -3215 1234 -3215 0 1
rlabel polysilicon 1234 -3221 1234 -3221 0 3
rlabel polysilicon 1241 -3215 1241 -3215 0 1
rlabel polysilicon 1241 -3221 1241 -3221 0 3
rlabel polysilicon 1248 -3215 1248 -3215 0 1
rlabel polysilicon 1248 -3221 1248 -3221 0 3
rlabel polysilicon 1255 -3215 1255 -3215 0 1
rlabel polysilicon 1255 -3221 1255 -3221 0 3
rlabel polysilicon 1262 -3215 1262 -3215 0 1
rlabel polysilicon 1262 -3221 1262 -3221 0 3
rlabel polysilicon 1269 -3215 1269 -3215 0 1
rlabel polysilicon 1269 -3221 1269 -3221 0 3
rlabel polysilicon 1276 -3215 1276 -3215 0 1
rlabel polysilicon 1276 -3221 1276 -3221 0 3
rlabel polysilicon 1283 -3215 1283 -3215 0 1
rlabel polysilicon 1283 -3221 1283 -3221 0 3
rlabel polysilicon 1290 -3215 1290 -3215 0 1
rlabel polysilicon 1290 -3221 1290 -3221 0 3
rlabel polysilicon 1297 -3215 1297 -3215 0 1
rlabel polysilicon 1300 -3221 1300 -3221 0 4
rlabel polysilicon 1304 -3215 1304 -3215 0 1
rlabel polysilicon 1304 -3221 1304 -3221 0 3
rlabel polysilicon 1311 -3215 1311 -3215 0 1
rlabel polysilicon 1311 -3221 1311 -3221 0 3
rlabel polysilicon 1318 -3215 1318 -3215 0 1
rlabel polysilicon 1318 -3221 1318 -3221 0 3
rlabel polysilicon 1325 -3215 1325 -3215 0 1
rlabel polysilicon 1325 -3221 1325 -3221 0 3
rlabel polysilicon 1328 -3221 1328 -3221 0 4
rlabel polysilicon 1332 -3215 1332 -3215 0 1
rlabel polysilicon 1332 -3221 1332 -3221 0 3
rlabel polysilicon 1339 -3215 1339 -3215 0 1
rlabel polysilicon 1339 -3221 1339 -3221 0 3
rlabel polysilicon 1346 -3215 1346 -3215 0 1
rlabel polysilicon 1346 -3221 1346 -3221 0 3
rlabel polysilicon 1349 -3221 1349 -3221 0 4
rlabel polysilicon 1353 -3221 1353 -3221 0 3
rlabel polysilicon 1356 -3221 1356 -3221 0 4
rlabel polysilicon 1360 -3215 1360 -3215 0 1
rlabel polysilicon 1360 -3221 1360 -3221 0 3
rlabel polysilicon 1367 -3215 1367 -3215 0 1
rlabel polysilicon 1367 -3221 1367 -3221 0 3
rlabel polysilicon 1374 -3215 1374 -3215 0 1
rlabel polysilicon 1374 -3221 1374 -3221 0 3
rlabel polysilicon 1381 -3215 1381 -3215 0 1
rlabel polysilicon 1381 -3221 1381 -3221 0 3
rlabel polysilicon 1388 -3215 1388 -3215 0 1
rlabel polysilicon 1388 -3221 1388 -3221 0 3
rlabel polysilicon 1395 -3215 1395 -3215 0 1
rlabel polysilicon 1395 -3221 1395 -3221 0 3
rlabel polysilicon 1402 -3215 1402 -3215 0 1
rlabel polysilicon 1402 -3221 1402 -3221 0 3
rlabel polysilicon 1409 -3215 1409 -3215 0 1
rlabel polysilicon 1412 -3215 1412 -3215 0 2
rlabel polysilicon 1409 -3221 1409 -3221 0 3
rlabel polysilicon 1416 -3215 1416 -3215 0 1
rlabel polysilicon 1416 -3221 1416 -3221 0 3
rlabel polysilicon 1423 -3215 1423 -3215 0 1
rlabel polysilicon 1423 -3221 1423 -3221 0 3
rlabel polysilicon 1430 -3215 1430 -3215 0 1
rlabel polysilicon 1430 -3221 1430 -3221 0 3
rlabel polysilicon 1437 -3215 1437 -3215 0 1
rlabel polysilicon 1437 -3221 1437 -3221 0 3
rlabel polysilicon 1444 -3215 1444 -3215 0 1
rlabel polysilicon 1444 -3221 1444 -3221 0 3
rlabel polysilicon 1451 -3215 1451 -3215 0 1
rlabel polysilicon 1451 -3221 1451 -3221 0 3
rlabel polysilicon 1458 -3215 1458 -3215 0 1
rlabel polysilicon 1458 -3221 1458 -3221 0 3
rlabel polysilicon 1465 -3215 1465 -3215 0 1
rlabel polysilicon 1465 -3221 1465 -3221 0 3
rlabel polysilicon 1475 -3215 1475 -3215 0 2
rlabel polysilicon 1475 -3221 1475 -3221 0 4
rlabel polysilicon 1479 -3215 1479 -3215 0 1
rlabel polysilicon 1479 -3221 1479 -3221 0 3
rlabel polysilicon 1486 -3215 1486 -3215 0 1
rlabel polysilicon 1486 -3221 1486 -3221 0 3
rlabel polysilicon 1493 -3215 1493 -3215 0 1
rlabel polysilicon 1493 -3221 1493 -3221 0 3
rlabel polysilicon 1500 -3215 1500 -3215 0 1
rlabel polysilicon 1500 -3221 1500 -3221 0 3
rlabel polysilicon 1507 -3215 1507 -3215 0 1
rlabel polysilicon 1507 -3221 1507 -3221 0 3
rlabel polysilicon 1514 -3215 1514 -3215 0 1
rlabel polysilicon 1514 -3221 1514 -3221 0 3
rlabel polysilicon 1521 -3215 1521 -3215 0 1
rlabel polysilicon 1521 -3221 1521 -3221 0 3
rlabel polysilicon 1605 -3215 1605 -3215 0 1
rlabel polysilicon 1605 -3221 1605 -3221 0 3
rlabel polysilicon 131 -3314 131 -3314 0 4
rlabel polysilicon 135 -3308 135 -3308 0 1
rlabel polysilicon 135 -3314 135 -3314 0 3
rlabel polysilicon 163 -3308 163 -3308 0 1
rlabel polysilicon 163 -3314 163 -3314 0 3
rlabel polysilicon 170 -3308 170 -3308 0 1
rlabel polysilicon 170 -3314 170 -3314 0 3
rlabel polysilicon 177 -3308 177 -3308 0 1
rlabel polysilicon 177 -3314 177 -3314 0 3
rlabel polysilicon 184 -3308 184 -3308 0 1
rlabel polysilicon 184 -3314 184 -3314 0 3
rlabel polysilicon 191 -3308 191 -3308 0 1
rlabel polysilicon 191 -3314 191 -3314 0 3
rlabel polysilicon 198 -3308 198 -3308 0 1
rlabel polysilicon 198 -3314 198 -3314 0 3
rlabel polysilicon 205 -3308 205 -3308 0 1
rlabel polysilicon 205 -3314 205 -3314 0 3
rlabel polysilicon 212 -3308 212 -3308 0 1
rlabel polysilicon 212 -3314 212 -3314 0 3
rlabel polysilicon 219 -3308 219 -3308 0 1
rlabel polysilicon 219 -3314 219 -3314 0 3
rlabel polysilicon 226 -3308 226 -3308 0 1
rlabel polysilicon 226 -3314 226 -3314 0 3
rlabel polysilicon 233 -3308 233 -3308 0 1
rlabel polysilicon 233 -3314 233 -3314 0 3
rlabel polysilicon 240 -3308 240 -3308 0 1
rlabel polysilicon 240 -3314 240 -3314 0 3
rlabel polysilicon 247 -3308 247 -3308 0 1
rlabel polysilicon 247 -3314 247 -3314 0 3
rlabel polysilicon 254 -3308 254 -3308 0 1
rlabel polysilicon 254 -3314 254 -3314 0 3
rlabel polysilicon 261 -3308 261 -3308 0 1
rlabel polysilicon 261 -3314 261 -3314 0 3
rlabel polysilicon 268 -3308 268 -3308 0 1
rlabel polysilicon 268 -3314 268 -3314 0 3
rlabel polysilicon 275 -3308 275 -3308 0 1
rlabel polysilicon 275 -3314 275 -3314 0 3
rlabel polysilicon 282 -3308 282 -3308 0 1
rlabel polysilicon 282 -3314 282 -3314 0 3
rlabel polysilicon 289 -3308 289 -3308 0 1
rlabel polysilicon 289 -3314 289 -3314 0 3
rlabel polysilicon 296 -3308 296 -3308 0 1
rlabel polysilicon 296 -3314 296 -3314 0 3
rlabel polysilicon 303 -3308 303 -3308 0 1
rlabel polysilicon 303 -3314 303 -3314 0 3
rlabel polysilicon 310 -3308 310 -3308 0 1
rlabel polysilicon 310 -3314 310 -3314 0 3
rlabel polysilicon 317 -3308 317 -3308 0 1
rlabel polysilicon 317 -3314 317 -3314 0 3
rlabel polysilicon 324 -3308 324 -3308 0 1
rlabel polysilicon 324 -3314 324 -3314 0 3
rlabel polysilicon 331 -3308 331 -3308 0 1
rlabel polysilicon 331 -3314 331 -3314 0 3
rlabel polysilicon 338 -3308 338 -3308 0 1
rlabel polysilicon 338 -3314 338 -3314 0 3
rlabel polysilicon 345 -3308 345 -3308 0 1
rlabel polysilicon 348 -3308 348 -3308 0 2
rlabel polysilicon 345 -3314 345 -3314 0 3
rlabel polysilicon 352 -3308 352 -3308 0 1
rlabel polysilicon 352 -3314 352 -3314 0 3
rlabel polysilicon 359 -3308 359 -3308 0 1
rlabel polysilicon 359 -3314 359 -3314 0 3
rlabel polysilicon 366 -3308 366 -3308 0 1
rlabel polysilicon 366 -3314 366 -3314 0 3
rlabel polysilicon 373 -3308 373 -3308 0 1
rlabel polysilicon 373 -3314 373 -3314 0 3
rlabel polysilicon 380 -3308 380 -3308 0 1
rlabel polysilicon 380 -3314 380 -3314 0 3
rlabel polysilicon 387 -3308 387 -3308 0 1
rlabel polysilicon 387 -3314 387 -3314 0 3
rlabel polysilicon 394 -3308 394 -3308 0 1
rlabel polysilicon 394 -3314 394 -3314 0 3
rlabel polysilicon 401 -3314 401 -3314 0 3
rlabel polysilicon 408 -3308 408 -3308 0 1
rlabel polysilicon 408 -3314 408 -3314 0 3
rlabel polysilicon 415 -3308 415 -3308 0 1
rlabel polysilicon 415 -3314 415 -3314 0 3
rlabel polysilicon 422 -3308 422 -3308 0 1
rlabel polysilicon 422 -3314 422 -3314 0 3
rlabel polysilicon 429 -3308 429 -3308 0 1
rlabel polysilicon 429 -3314 429 -3314 0 3
rlabel polysilicon 436 -3308 436 -3308 0 1
rlabel polysilicon 439 -3308 439 -3308 0 2
rlabel polysilicon 443 -3308 443 -3308 0 1
rlabel polysilicon 443 -3314 443 -3314 0 3
rlabel polysilicon 446 -3314 446 -3314 0 4
rlabel polysilicon 450 -3308 450 -3308 0 1
rlabel polysilicon 450 -3314 450 -3314 0 3
rlabel polysilicon 457 -3308 457 -3308 0 1
rlabel polysilicon 457 -3314 457 -3314 0 3
rlabel polysilicon 464 -3308 464 -3308 0 1
rlabel polysilicon 464 -3314 464 -3314 0 3
rlabel polysilicon 471 -3308 471 -3308 0 1
rlabel polysilicon 471 -3314 471 -3314 0 3
rlabel polysilicon 478 -3308 478 -3308 0 1
rlabel polysilicon 478 -3314 478 -3314 0 3
rlabel polysilicon 485 -3308 485 -3308 0 1
rlabel polysilicon 485 -3314 485 -3314 0 3
rlabel polysilicon 492 -3308 492 -3308 0 1
rlabel polysilicon 499 -3308 499 -3308 0 1
rlabel polysilicon 499 -3314 499 -3314 0 3
rlabel polysilicon 506 -3308 506 -3308 0 1
rlabel polysilicon 506 -3314 506 -3314 0 3
rlabel polysilicon 513 -3308 513 -3308 0 1
rlabel polysilicon 513 -3314 513 -3314 0 3
rlabel polysilicon 520 -3308 520 -3308 0 1
rlabel polysilicon 520 -3314 520 -3314 0 3
rlabel polysilicon 527 -3308 527 -3308 0 1
rlabel polysilicon 530 -3308 530 -3308 0 2
rlabel polysilicon 527 -3314 527 -3314 0 3
rlabel polysilicon 530 -3314 530 -3314 0 4
rlabel polysilicon 534 -3308 534 -3308 0 1
rlabel polysilicon 534 -3314 534 -3314 0 3
rlabel polysilicon 541 -3308 541 -3308 0 1
rlabel polysilicon 544 -3308 544 -3308 0 2
rlabel polysilicon 544 -3314 544 -3314 0 4
rlabel polysilicon 548 -3308 548 -3308 0 1
rlabel polysilicon 548 -3314 548 -3314 0 3
rlabel polysilicon 555 -3308 555 -3308 0 1
rlabel polysilicon 555 -3314 555 -3314 0 3
rlabel polysilicon 562 -3308 562 -3308 0 1
rlabel polysilicon 562 -3314 562 -3314 0 3
rlabel polysilicon 569 -3308 569 -3308 0 1
rlabel polysilicon 569 -3314 569 -3314 0 3
rlabel polysilicon 576 -3308 576 -3308 0 1
rlabel polysilicon 576 -3314 576 -3314 0 3
rlabel polysilicon 583 -3308 583 -3308 0 1
rlabel polysilicon 583 -3314 583 -3314 0 3
rlabel polysilicon 590 -3308 590 -3308 0 1
rlabel polysilicon 590 -3314 590 -3314 0 3
rlabel polysilicon 597 -3308 597 -3308 0 1
rlabel polysilicon 597 -3314 597 -3314 0 3
rlabel polysilicon 604 -3308 604 -3308 0 1
rlabel polysilicon 604 -3314 604 -3314 0 3
rlabel polysilicon 611 -3308 611 -3308 0 1
rlabel polysilicon 611 -3314 611 -3314 0 3
rlabel polysilicon 618 -3308 618 -3308 0 1
rlabel polysilicon 618 -3314 618 -3314 0 3
rlabel polysilicon 621 -3314 621 -3314 0 4
rlabel polysilicon 625 -3308 625 -3308 0 1
rlabel polysilicon 625 -3314 625 -3314 0 3
rlabel polysilicon 632 -3308 632 -3308 0 1
rlabel polysilicon 632 -3314 632 -3314 0 3
rlabel polysilicon 639 -3308 639 -3308 0 1
rlabel polysilicon 639 -3314 639 -3314 0 3
rlabel polysilicon 646 -3314 646 -3314 0 3
rlabel polysilicon 653 -3308 653 -3308 0 1
rlabel polysilicon 653 -3314 653 -3314 0 3
rlabel polysilicon 660 -3308 660 -3308 0 1
rlabel polysilicon 660 -3314 660 -3314 0 3
rlabel polysilicon 667 -3308 667 -3308 0 1
rlabel polysilicon 667 -3314 667 -3314 0 3
rlabel polysilicon 677 -3308 677 -3308 0 2
rlabel polysilicon 674 -3314 674 -3314 0 3
rlabel polysilicon 681 -3308 681 -3308 0 1
rlabel polysilicon 681 -3314 681 -3314 0 3
rlabel polysilicon 688 -3314 688 -3314 0 3
rlabel polysilicon 691 -3314 691 -3314 0 4
rlabel polysilicon 695 -3308 695 -3308 0 1
rlabel polysilicon 695 -3314 695 -3314 0 3
rlabel polysilicon 702 -3308 702 -3308 0 1
rlabel polysilicon 705 -3308 705 -3308 0 2
rlabel polysilicon 702 -3314 702 -3314 0 3
rlabel polysilicon 705 -3314 705 -3314 0 4
rlabel polysilicon 709 -3308 709 -3308 0 1
rlabel polysilicon 709 -3314 709 -3314 0 3
rlabel polysilicon 716 -3308 716 -3308 0 1
rlabel polysilicon 716 -3314 716 -3314 0 3
rlabel polysilicon 723 -3308 723 -3308 0 1
rlabel polysilicon 723 -3314 723 -3314 0 3
rlabel polysilicon 730 -3308 730 -3308 0 1
rlabel polysilicon 730 -3314 730 -3314 0 3
rlabel polysilicon 737 -3308 737 -3308 0 1
rlabel polysilicon 737 -3314 737 -3314 0 3
rlabel polysilicon 744 -3308 744 -3308 0 1
rlabel polysilicon 744 -3314 744 -3314 0 3
rlabel polysilicon 751 -3308 751 -3308 0 1
rlabel polysilicon 751 -3314 751 -3314 0 3
rlabel polysilicon 758 -3308 758 -3308 0 1
rlabel polysilicon 758 -3314 758 -3314 0 3
rlabel polysilicon 765 -3308 765 -3308 0 1
rlabel polysilicon 765 -3314 765 -3314 0 3
rlabel polysilicon 772 -3308 772 -3308 0 1
rlabel polysilicon 772 -3314 772 -3314 0 3
rlabel polysilicon 779 -3308 779 -3308 0 1
rlabel polysilicon 779 -3314 779 -3314 0 3
rlabel polysilicon 789 -3308 789 -3308 0 2
rlabel polysilicon 786 -3314 786 -3314 0 3
rlabel polysilicon 789 -3314 789 -3314 0 4
rlabel polysilicon 793 -3308 793 -3308 0 1
rlabel polysilicon 793 -3314 793 -3314 0 3
rlabel polysilicon 800 -3308 800 -3308 0 1
rlabel polysilicon 800 -3314 800 -3314 0 3
rlabel polysilicon 807 -3308 807 -3308 0 1
rlabel polysilicon 807 -3314 807 -3314 0 3
rlabel polysilicon 814 -3308 814 -3308 0 1
rlabel polysilicon 814 -3314 814 -3314 0 3
rlabel polysilicon 821 -3308 821 -3308 0 1
rlabel polysilicon 821 -3314 821 -3314 0 3
rlabel polysilicon 828 -3308 828 -3308 0 1
rlabel polysilicon 828 -3314 828 -3314 0 3
rlabel polysilicon 835 -3308 835 -3308 0 1
rlabel polysilicon 835 -3314 835 -3314 0 3
rlabel polysilicon 842 -3308 842 -3308 0 1
rlabel polysilicon 842 -3314 842 -3314 0 3
rlabel polysilicon 849 -3308 849 -3308 0 1
rlabel polysilicon 849 -3314 849 -3314 0 3
rlabel polysilicon 856 -3308 856 -3308 0 1
rlabel polysilicon 856 -3314 856 -3314 0 3
rlabel polysilicon 863 -3308 863 -3308 0 1
rlabel polysilicon 863 -3314 863 -3314 0 3
rlabel polysilicon 870 -3314 870 -3314 0 3
rlabel polysilicon 873 -3314 873 -3314 0 4
rlabel polysilicon 877 -3308 877 -3308 0 1
rlabel polysilicon 880 -3308 880 -3308 0 2
rlabel polysilicon 877 -3314 877 -3314 0 3
rlabel polysilicon 880 -3314 880 -3314 0 4
rlabel polysilicon 884 -3308 884 -3308 0 1
rlabel polysilicon 884 -3314 884 -3314 0 3
rlabel polysilicon 891 -3308 891 -3308 0 1
rlabel polysilicon 891 -3314 891 -3314 0 3
rlabel polysilicon 901 -3308 901 -3308 0 2
rlabel polysilicon 898 -3314 898 -3314 0 3
rlabel polysilicon 901 -3314 901 -3314 0 4
rlabel polysilicon 905 -3308 905 -3308 0 1
rlabel polysilicon 905 -3314 905 -3314 0 3
rlabel polysilicon 908 -3314 908 -3314 0 4
rlabel polysilicon 912 -3308 912 -3308 0 1
rlabel polysilicon 915 -3308 915 -3308 0 2
rlabel polysilicon 912 -3314 912 -3314 0 3
rlabel polysilicon 915 -3314 915 -3314 0 4
rlabel polysilicon 919 -3308 919 -3308 0 1
rlabel polysilicon 919 -3314 919 -3314 0 3
rlabel polysilicon 926 -3308 926 -3308 0 1
rlabel polysilicon 926 -3314 926 -3314 0 3
rlabel polysilicon 933 -3308 933 -3308 0 1
rlabel polysilicon 933 -3314 933 -3314 0 3
rlabel polysilicon 940 -3308 940 -3308 0 1
rlabel polysilicon 940 -3314 940 -3314 0 3
rlabel polysilicon 947 -3308 947 -3308 0 1
rlabel polysilicon 947 -3314 947 -3314 0 3
rlabel polysilicon 954 -3308 954 -3308 0 1
rlabel polysilicon 954 -3314 954 -3314 0 3
rlabel polysilicon 961 -3308 961 -3308 0 1
rlabel polysilicon 961 -3314 961 -3314 0 3
rlabel polysilicon 968 -3308 968 -3308 0 1
rlabel polysilicon 968 -3314 968 -3314 0 3
rlabel polysilicon 975 -3308 975 -3308 0 1
rlabel polysilicon 975 -3314 975 -3314 0 3
rlabel polysilicon 982 -3308 982 -3308 0 1
rlabel polysilicon 985 -3308 985 -3308 0 2
rlabel polysilicon 982 -3314 982 -3314 0 3
rlabel polysilicon 985 -3314 985 -3314 0 4
rlabel polysilicon 989 -3308 989 -3308 0 1
rlabel polysilicon 989 -3314 989 -3314 0 3
rlabel polysilicon 996 -3308 996 -3308 0 1
rlabel polysilicon 996 -3314 996 -3314 0 3
rlabel polysilicon 1003 -3308 1003 -3308 0 1
rlabel polysilicon 1003 -3314 1003 -3314 0 3
rlabel polysilicon 1010 -3308 1010 -3308 0 1
rlabel polysilicon 1010 -3314 1010 -3314 0 3
rlabel polysilicon 1020 -3308 1020 -3308 0 2
rlabel polysilicon 1020 -3314 1020 -3314 0 4
rlabel polysilicon 1024 -3308 1024 -3308 0 1
rlabel polysilicon 1024 -3314 1024 -3314 0 3
rlabel polysilicon 1031 -3308 1031 -3308 0 1
rlabel polysilicon 1031 -3314 1031 -3314 0 3
rlabel polysilicon 1038 -3308 1038 -3308 0 1
rlabel polysilicon 1038 -3314 1038 -3314 0 3
rlabel polysilicon 1045 -3308 1045 -3308 0 1
rlabel polysilicon 1045 -3314 1045 -3314 0 3
rlabel polysilicon 1052 -3308 1052 -3308 0 1
rlabel polysilicon 1052 -3314 1052 -3314 0 3
rlabel polysilicon 1059 -3308 1059 -3308 0 1
rlabel polysilicon 1059 -3314 1059 -3314 0 3
rlabel polysilicon 1066 -3308 1066 -3308 0 1
rlabel polysilicon 1066 -3314 1066 -3314 0 3
rlabel polysilicon 1073 -3308 1073 -3308 0 1
rlabel polysilicon 1073 -3314 1073 -3314 0 3
rlabel polysilicon 1080 -3308 1080 -3308 0 1
rlabel polysilicon 1080 -3314 1080 -3314 0 3
rlabel polysilicon 1087 -3308 1087 -3308 0 1
rlabel polysilicon 1087 -3314 1087 -3314 0 3
rlabel polysilicon 1094 -3308 1094 -3308 0 1
rlabel polysilicon 1094 -3314 1094 -3314 0 3
rlabel polysilicon 1101 -3308 1101 -3308 0 1
rlabel polysilicon 1101 -3314 1101 -3314 0 3
rlabel polysilicon 1108 -3308 1108 -3308 0 1
rlabel polysilicon 1108 -3314 1108 -3314 0 3
rlabel polysilicon 1111 -3314 1111 -3314 0 4
rlabel polysilicon 1115 -3308 1115 -3308 0 1
rlabel polysilicon 1115 -3314 1115 -3314 0 3
rlabel polysilicon 1122 -3308 1122 -3308 0 1
rlabel polysilicon 1122 -3314 1122 -3314 0 3
rlabel polysilicon 1129 -3308 1129 -3308 0 1
rlabel polysilicon 1129 -3314 1129 -3314 0 3
rlabel polysilicon 1136 -3308 1136 -3308 0 1
rlabel polysilicon 1136 -3314 1136 -3314 0 3
rlabel polysilicon 1143 -3308 1143 -3308 0 1
rlabel polysilicon 1143 -3314 1143 -3314 0 3
rlabel polysilicon 1150 -3308 1150 -3308 0 1
rlabel polysilicon 1150 -3314 1150 -3314 0 3
rlabel polysilicon 1157 -3308 1157 -3308 0 1
rlabel polysilicon 1157 -3314 1157 -3314 0 3
rlabel polysilicon 1164 -3308 1164 -3308 0 1
rlabel polysilicon 1164 -3314 1164 -3314 0 3
rlabel polysilicon 1171 -3308 1171 -3308 0 1
rlabel polysilicon 1171 -3314 1171 -3314 0 3
rlabel polysilicon 1178 -3308 1178 -3308 0 1
rlabel polysilicon 1178 -3314 1178 -3314 0 3
rlabel polysilicon 1188 -3308 1188 -3308 0 2
rlabel polysilicon 1185 -3314 1185 -3314 0 3
rlabel polysilicon 1192 -3308 1192 -3308 0 1
rlabel polysilicon 1192 -3314 1192 -3314 0 3
rlabel polysilicon 1199 -3308 1199 -3308 0 1
rlabel polysilicon 1199 -3314 1199 -3314 0 3
rlabel polysilicon 1209 -3308 1209 -3308 0 2
rlabel polysilicon 1206 -3314 1206 -3314 0 3
rlabel polysilicon 1209 -3314 1209 -3314 0 4
rlabel polysilicon 1213 -3308 1213 -3308 0 1
rlabel polysilicon 1213 -3314 1213 -3314 0 3
rlabel polysilicon 1216 -3314 1216 -3314 0 4
rlabel polysilicon 1220 -3308 1220 -3308 0 1
rlabel polysilicon 1220 -3314 1220 -3314 0 3
rlabel polysilicon 1227 -3308 1227 -3308 0 1
rlabel polysilicon 1227 -3314 1227 -3314 0 3
rlabel polysilicon 1234 -3308 1234 -3308 0 1
rlabel polysilicon 1234 -3314 1234 -3314 0 3
rlabel polysilicon 1241 -3308 1241 -3308 0 1
rlabel polysilicon 1241 -3314 1241 -3314 0 3
rlabel polysilicon 1248 -3314 1248 -3314 0 3
rlabel polysilicon 1251 -3314 1251 -3314 0 4
rlabel polysilicon 1255 -3308 1255 -3308 0 1
rlabel polysilicon 1258 -3308 1258 -3308 0 2
rlabel polysilicon 1262 -3308 1262 -3308 0 1
rlabel polysilicon 1265 -3308 1265 -3308 0 2
rlabel polysilicon 1262 -3314 1262 -3314 0 3
rlabel polysilicon 1265 -3314 1265 -3314 0 4
rlabel polysilicon 1269 -3308 1269 -3308 0 1
rlabel polysilicon 1269 -3314 1269 -3314 0 3
rlabel polysilicon 1276 -3308 1276 -3308 0 1
rlabel polysilicon 1276 -3314 1276 -3314 0 3
rlabel polysilicon 1283 -3308 1283 -3308 0 1
rlabel polysilicon 1283 -3314 1283 -3314 0 3
rlabel polysilicon 1290 -3308 1290 -3308 0 1
rlabel polysilicon 1290 -3314 1290 -3314 0 3
rlabel polysilicon 1297 -3308 1297 -3308 0 1
rlabel polysilicon 1297 -3314 1297 -3314 0 3
rlabel polysilicon 1304 -3308 1304 -3308 0 1
rlabel polysilicon 1304 -3314 1304 -3314 0 3
rlabel polysilicon 1311 -3308 1311 -3308 0 1
rlabel polysilicon 1311 -3314 1311 -3314 0 3
rlabel polysilicon 1318 -3308 1318 -3308 0 1
rlabel polysilicon 1318 -3314 1318 -3314 0 3
rlabel polysilicon 1325 -3308 1325 -3308 0 1
rlabel polysilicon 1328 -3308 1328 -3308 0 2
rlabel polysilicon 1325 -3314 1325 -3314 0 3
rlabel polysilicon 1332 -3308 1332 -3308 0 1
rlabel polysilicon 1332 -3314 1332 -3314 0 3
rlabel polysilicon 1339 -3308 1339 -3308 0 1
rlabel polysilicon 1339 -3314 1339 -3314 0 3
rlabel polysilicon 1346 -3308 1346 -3308 0 1
rlabel polysilicon 1346 -3314 1346 -3314 0 3
rlabel polysilicon 1353 -3308 1353 -3308 0 1
rlabel polysilicon 1353 -3314 1353 -3314 0 3
rlabel polysilicon 1360 -3308 1360 -3308 0 1
rlabel polysilicon 1360 -3314 1360 -3314 0 3
rlabel polysilicon 1381 -3308 1381 -3308 0 1
rlabel polysilicon 1381 -3314 1381 -3314 0 3
rlabel polysilicon 1388 -3308 1388 -3308 0 1
rlabel polysilicon 1388 -3314 1388 -3314 0 3
rlabel polysilicon 1531 -3308 1531 -3308 0 2
rlabel polysilicon 1528 -3314 1528 -3314 0 3
rlabel polysilicon 1584 -3308 1584 -3308 0 1
rlabel polysilicon 1584 -3314 1584 -3314 0 3
rlabel polysilicon 240 -3405 240 -3405 0 1
rlabel polysilicon 240 -3411 240 -3411 0 3
rlabel polysilicon 247 -3405 247 -3405 0 1
rlabel polysilicon 247 -3411 247 -3411 0 3
rlabel polysilicon 268 -3405 268 -3405 0 1
rlabel polysilicon 268 -3411 268 -3411 0 3
rlabel polysilicon 282 -3405 282 -3405 0 1
rlabel polysilicon 282 -3411 282 -3411 0 3
rlabel polysilicon 289 -3405 289 -3405 0 1
rlabel polysilicon 289 -3411 289 -3411 0 3
rlabel polysilicon 292 -3411 292 -3411 0 4
rlabel polysilicon 296 -3405 296 -3405 0 1
rlabel polysilicon 299 -3411 299 -3411 0 4
rlabel polysilicon 303 -3405 303 -3405 0 1
rlabel polysilicon 303 -3411 303 -3411 0 3
rlabel polysilicon 310 -3405 310 -3405 0 1
rlabel polysilicon 310 -3411 310 -3411 0 3
rlabel polysilicon 317 -3405 317 -3405 0 1
rlabel polysilicon 317 -3411 317 -3411 0 3
rlabel polysilicon 324 -3405 324 -3405 0 1
rlabel polysilicon 324 -3411 324 -3411 0 3
rlabel polysilicon 331 -3405 331 -3405 0 1
rlabel polysilicon 331 -3411 331 -3411 0 3
rlabel polysilicon 338 -3405 338 -3405 0 1
rlabel polysilicon 338 -3411 338 -3411 0 3
rlabel polysilicon 345 -3405 345 -3405 0 1
rlabel polysilicon 345 -3411 345 -3411 0 3
rlabel polysilicon 352 -3405 352 -3405 0 1
rlabel polysilicon 352 -3411 352 -3411 0 3
rlabel polysilicon 359 -3405 359 -3405 0 1
rlabel polysilicon 359 -3411 359 -3411 0 3
rlabel polysilicon 366 -3405 366 -3405 0 1
rlabel polysilicon 366 -3411 366 -3411 0 3
rlabel polysilicon 373 -3405 373 -3405 0 1
rlabel polysilicon 376 -3411 376 -3411 0 4
rlabel polysilicon 380 -3405 380 -3405 0 1
rlabel polysilicon 380 -3411 380 -3411 0 3
rlabel polysilicon 387 -3405 387 -3405 0 1
rlabel polysilicon 387 -3411 387 -3411 0 3
rlabel polysilicon 394 -3405 394 -3405 0 1
rlabel polysilicon 394 -3411 394 -3411 0 3
rlabel polysilicon 401 -3405 401 -3405 0 1
rlabel polysilicon 401 -3411 401 -3411 0 3
rlabel polysilicon 408 -3405 408 -3405 0 1
rlabel polysilicon 408 -3411 408 -3411 0 3
rlabel polysilicon 415 -3405 415 -3405 0 1
rlabel polysilicon 415 -3411 415 -3411 0 3
rlabel polysilicon 422 -3405 422 -3405 0 1
rlabel polysilicon 422 -3411 422 -3411 0 3
rlabel polysilicon 429 -3405 429 -3405 0 1
rlabel polysilicon 429 -3411 429 -3411 0 3
rlabel polysilicon 436 -3405 436 -3405 0 1
rlabel polysilicon 436 -3411 436 -3411 0 3
rlabel polysilicon 443 -3405 443 -3405 0 1
rlabel polysilicon 443 -3411 443 -3411 0 3
rlabel polysilicon 450 -3405 450 -3405 0 1
rlabel polysilicon 450 -3411 450 -3411 0 3
rlabel polysilicon 457 -3405 457 -3405 0 1
rlabel polysilicon 457 -3411 457 -3411 0 3
rlabel polysilicon 464 -3405 464 -3405 0 1
rlabel polysilicon 464 -3411 464 -3411 0 3
rlabel polysilicon 471 -3405 471 -3405 0 1
rlabel polysilicon 471 -3411 471 -3411 0 3
rlabel polysilicon 478 -3405 478 -3405 0 1
rlabel polysilicon 478 -3411 478 -3411 0 3
rlabel polysilicon 485 -3405 485 -3405 0 1
rlabel polysilicon 485 -3411 485 -3411 0 3
rlabel polysilicon 492 -3405 492 -3405 0 1
rlabel polysilicon 492 -3411 492 -3411 0 3
rlabel polysilicon 499 -3405 499 -3405 0 1
rlabel polysilicon 499 -3411 499 -3411 0 3
rlabel polysilicon 506 -3405 506 -3405 0 1
rlabel polysilicon 506 -3411 506 -3411 0 3
rlabel polysilicon 513 -3405 513 -3405 0 1
rlabel polysilicon 513 -3411 513 -3411 0 3
rlabel polysilicon 523 -3405 523 -3405 0 2
rlabel polysilicon 520 -3411 520 -3411 0 3
rlabel polysilicon 523 -3411 523 -3411 0 4
rlabel polysilicon 527 -3405 527 -3405 0 1
rlabel polysilicon 527 -3411 527 -3411 0 3
rlabel polysilicon 534 -3405 534 -3405 0 1
rlabel polysilicon 534 -3411 534 -3411 0 3
rlabel polysilicon 541 -3405 541 -3405 0 1
rlabel polysilicon 541 -3411 541 -3411 0 3
rlabel polysilicon 548 -3405 548 -3405 0 1
rlabel polysilicon 548 -3411 548 -3411 0 3
rlabel polysilicon 555 -3405 555 -3405 0 1
rlabel polysilicon 555 -3411 555 -3411 0 3
rlabel polysilicon 562 -3405 562 -3405 0 1
rlabel polysilicon 562 -3411 562 -3411 0 3
rlabel polysilicon 569 -3405 569 -3405 0 1
rlabel polysilicon 569 -3411 569 -3411 0 3
rlabel polysilicon 576 -3405 576 -3405 0 1
rlabel polysilicon 579 -3405 579 -3405 0 2
rlabel polysilicon 579 -3411 579 -3411 0 4
rlabel polysilicon 583 -3405 583 -3405 0 1
rlabel polysilicon 583 -3411 583 -3411 0 3
rlabel polysilicon 590 -3405 590 -3405 0 1
rlabel polysilicon 590 -3411 590 -3411 0 3
rlabel polysilicon 597 -3405 597 -3405 0 1
rlabel polysilicon 597 -3411 597 -3411 0 3
rlabel polysilicon 604 -3405 604 -3405 0 1
rlabel polysilicon 604 -3411 604 -3411 0 3
rlabel polysilicon 611 -3405 611 -3405 0 1
rlabel polysilicon 614 -3405 614 -3405 0 2
rlabel polysilicon 614 -3411 614 -3411 0 4
rlabel polysilicon 618 -3405 618 -3405 0 1
rlabel polysilicon 618 -3411 618 -3411 0 3
rlabel polysilicon 625 -3405 625 -3405 0 1
rlabel polysilicon 625 -3411 625 -3411 0 3
rlabel polysilicon 632 -3405 632 -3405 0 1
rlabel polysilicon 632 -3411 632 -3411 0 3
rlabel polysilicon 639 -3405 639 -3405 0 1
rlabel polysilicon 639 -3411 639 -3411 0 3
rlabel polysilicon 646 -3405 646 -3405 0 1
rlabel polysilicon 646 -3411 646 -3411 0 3
rlabel polysilicon 653 -3405 653 -3405 0 1
rlabel polysilicon 653 -3411 653 -3411 0 3
rlabel polysilicon 660 -3405 660 -3405 0 1
rlabel polysilicon 660 -3411 660 -3411 0 3
rlabel polysilicon 667 -3405 667 -3405 0 1
rlabel polysilicon 667 -3411 667 -3411 0 3
rlabel polysilicon 674 -3405 674 -3405 0 1
rlabel polysilicon 674 -3411 674 -3411 0 3
rlabel polysilicon 681 -3405 681 -3405 0 1
rlabel polysilicon 681 -3411 681 -3411 0 3
rlabel polysilicon 688 -3405 688 -3405 0 1
rlabel polysilicon 688 -3411 688 -3411 0 3
rlabel polysilicon 695 -3405 695 -3405 0 1
rlabel polysilicon 695 -3411 695 -3411 0 3
rlabel polysilicon 702 -3405 702 -3405 0 1
rlabel polysilicon 702 -3411 702 -3411 0 3
rlabel polysilicon 709 -3405 709 -3405 0 1
rlabel polysilicon 709 -3411 709 -3411 0 3
rlabel polysilicon 716 -3405 716 -3405 0 1
rlabel polysilicon 716 -3411 716 -3411 0 3
rlabel polysilicon 723 -3405 723 -3405 0 1
rlabel polysilicon 723 -3411 723 -3411 0 3
rlabel polysilicon 730 -3411 730 -3411 0 3
rlabel polysilicon 733 -3411 733 -3411 0 4
rlabel polysilicon 737 -3405 737 -3405 0 1
rlabel polysilicon 737 -3411 737 -3411 0 3
rlabel polysilicon 744 -3405 744 -3405 0 1
rlabel polysilicon 744 -3411 744 -3411 0 3
rlabel polysilicon 751 -3405 751 -3405 0 1
rlabel polysilicon 751 -3411 751 -3411 0 3
rlabel polysilicon 758 -3405 758 -3405 0 1
rlabel polysilicon 758 -3411 758 -3411 0 3
rlabel polysilicon 765 -3405 765 -3405 0 1
rlabel polysilicon 765 -3411 765 -3411 0 3
rlabel polysilicon 772 -3405 772 -3405 0 1
rlabel polysilicon 772 -3411 772 -3411 0 3
rlabel polysilicon 779 -3405 779 -3405 0 1
rlabel polysilicon 779 -3411 779 -3411 0 3
rlabel polysilicon 786 -3405 786 -3405 0 1
rlabel polysilicon 786 -3411 786 -3411 0 3
rlabel polysilicon 793 -3405 793 -3405 0 1
rlabel polysilicon 793 -3411 793 -3411 0 3
rlabel polysilicon 800 -3405 800 -3405 0 1
rlabel polysilicon 803 -3405 803 -3405 0 2
rlabel polysilicon 803 -3411 803 -3411 0 4
rlabel polysilicon 807 -3405 807 -3405 0 1
rlabel polysilicon 807 -3411 807 -3411 0 3
rlabel polysilicon 814 -3405 814 -3405 0 1
rlabel polysilicon 814 -3411 814 -3411 0 3
rlabel polysilicon 821 -3405 821 -3405 0 1
rlabel polysilicon 821 -3411 821 -3411 0 3
rlabel polysilicon 828 -3405 828 -3405 0 1
rlabel polysilicon 828 -3411 828 -3411 0 3
rlabel polysilicon 835 -3405 835 -3405 0 1
rlabel polysilicon 835 -3411 835 -3411 0 3
rlabel polysilicon 842 -3405 842 -3405 0 1
rlabel polysilicon 842 -3411 842 -3411 0 3
rlabel polysilicon 849 -3405 849 -3405 0 1
rlabel polysilicon 849 -3411 849 -3411 0 3
rlabel polysilicon 856 -3405 856 -3405 0 1
rlabel polysilicon 856 -3411 856 -3411 0 3
rlabel polysilicon 863 -3405 863 -3405 0 1
rlabel polysilicon 863 -3411 863 -3411 0 3
rlabel polysilicon 870 -3405 870 -3405 0 1
rlabel polysilicon 870 -3411 870 -3411 0 3
rlabel polysilicon 877 -3405 877 -3405 0 1
rlabel polysilicon 877 -3411 877 -3411 0 3
rlabel polysilicon 884 -3405 884 -3405 0 1
rlabel polysilicon 884 -3411 884 -3411 0 3
rlabel polysilicon 894 -3405 894 -3405 0 2
rlabel polysilicon 891 -3411 891 -3411 0 3
rlabel polysilicon 894 -3411 894 -3411 0 4
rlabel polysilicon 898 -3405 898 -3405 0 1
rlabel polysilicon 898 -3411 898 -3411 0 3
rlabel polysilicon 905 -3405 905 -3405 0 1
rlabel polysilicon 905 -3411 905 -3411 0 3
rlabel polysilicon 912 -3405 912 -3405 0 1
rlabel polysilicon 912 -3411 912 -3411 0 3
rlabel polysilicon 919 -3405 919 -3405 0 1
rlabel polysilicon 919 -3411 919 -3411 0 3
rlabel polysilicon 926 -3405 926 -3405 0 1
rlabel polysilicon 926 -3411 926 -3411 0 3
rlabel polysilicon 933 -3405 933 -3405 0 1
rlabel polysilicon 933 -3411 933 -3411 0 3
rlabel polysilicon 940 -3405 940 -3405 0 1
rlabel polysilicon 940 -3411 940 -3411 0 3
rlabel polysilicon 947 -3405 947 -3405 0 1
rlabel polysilicon 950 -3405 950 -3405 0 2
rlabel polysilicon 947 -3411 947 -3411 0 3
rlabel polysilicon 954 -3405 954 -3405 0 1
rlabel polysilicon 954 -3411 954 -3411 0 3
rlabel polysilicon 961 -3405 961 -3405 0 1
rlabel polysilicon 961 -3411 961 -3411 0 3
rlabel polysilicon 968 -3405 968 -3405 0 1
rlabel polysilicon 968 -3411 968 -3411 0 3
rlabel polysilicon 975 -3405 975 -3405 0 1
rlabel polysilicon 975 -3411 975 -3411 0 3
rlabel polysilicon 982 -3405 982 -3405 0 1
rlabel polysilicon 982 -3411 982 -3411 0 3
rlabel polysilicon 989 -3405 989 -3405 0 1
rlabel polysilicon 989 -3411 989 -3411 0 3
rlabel polysilicon 996 -3405 996 -3405 0 1
rlabel polysilicon 996 -3411 996 -3411 0 3
rlabel polysilicon 1003 -3405 1003 -3405 0 1
rlabel polysilicon 1003 -3411 1003 -3411 0 3
rlabel polysilicon 1013 -3405 1013 -3405 0 2
rlabel polysilicon 1010 -3411 1010 -3411 0 3
rlabel polysilicon 1017 -3405 1017 -3405 0 1
rlabel polysilicon 1020 -3405 1020 -3405 0 2
rlabel polysilicon 1017 -3411 1017 -3411 0 3
rlabel polysilicon 1020 -3411 1020 -3411 0 4
rlabel polysilicon 1024 -3405 1024 -3405 0 1
rlabel polysilicon 1024 -3411 1024 -3411 0 3
rlabel polysilicon 1031 -3405 1031 -3405 0 1
rlabel polysilicon 1031 -3411 1031 -3411 0 3
rlabel polysilicon 1038 -3405 1038 -3405 0 1
rlabel polysilicon 1038 -3411 1038 -3411 0 3
rlabel polysilicon 1041 -3411 1041 -3411 0 4
rlabel polysilicon 1045 -3405 1045 -3405 0 1
rlabel polysilicon 1045 -3411 1045 -3411 0 3
rlabel polysilicon 1055 -3411 1055 -3411 0 4
rlabel polysilicon 1059 -3405 1059 -3405 0 1
rlabel polysilicon 1062 -3405 1062 -3405 0 2
rlabel polysilicon 1066 -3405 1066 -3405 0 1
rlabel polysilicon 1066 -3411 1066 -3411 0 3
rlabel polysilicon 1073 -3405 1073 -3405 0 1
rlabel polysilicon 1073 -3411 1073 -3411 0 3
rlabel polysilicon 1080 -3405 1080 -3405 0 1
rlabel polysilicon 1080 -3411 1080 -3411 0 3
rlabel polysilicon 1087 -3405 1087 -3405 0 1
rlabel polysilicon 1087 -3411 1087 -3411 0 3
rlabel polysilicon 1094 -3405 1094 -3405 0 1
rlabel polysilicon 1094 -3411 1094 -3411 0 3
rlabel polysilicon 1101 -3405 1101 -3405 0 1
rlabel polysilicon 1101 -3411 1101 -3411 0 3
rlabel polysilicon 1108 -3405 1108 -3405 0 1
rlabel polysilicon 1111 -3411 1111 -3411 0 4
rlabel polysilicon 1115 -3405 1115 -3405 0 1
rlabel polysilicon 1115 -3411 1115 -3411 0 3
rlabel polysilicon 1122 -3405 1122 -3405 0 1
rlabel polysilicon 1122 -3411 1122 -3411 0 3
rlabel polysilicon 1129 -3405 1129 -3405 0 1
rlabel polysilicon 1129 -3411 1129 -3411 0 3
rlabel polysilicon 1136 -3405 1136 -3405 0 1
rlabel polysilicon 1136 -3411 1136 -3411 0 3
rlabel polysilicon 1143 -3405 1143 -3405 0 1
rlabel polysilicon 1153 -3405 1153 -3405 0 2
rlabel polysilicon 1150 -3411 1150 -3411 0 3
rlabel polysilicon 1153 -3411 1153 -3411 0 4
rlabel polysilicon 1157 -3405 1157 -3405 0 1
rlabel polysilicon 1157 -3411 1157 -3411 0 3
rlabel polysilicon 1160 -3411 1160 -3411 0 4
rlabel polysilicon 1164 -3405 1164 -3405 0 1
rlabel polysilicon 1167 -3405 1167 -3405 0 2
rlabel polysilicon 1167 -3411 1167 -3411 0 4
rlabel polysilicon 1171 -3405 1171 -3405 0 1
rlabel polysilicon 1171 -3411 1171 -3411 0 3
rlabel polysilicon 1185 -3405 1185 -3405 0 1
rlabel polysilicon 1185 -3411 1185 -3411 0 3
rlabel polysilicon 1192 -3405 1192 -3405 0 1
rlabel polysilicon 1192 -3411 1192 -3411 0 3
rlabel polysilicon 1199 -3405 1199 -3405 0 1
rlabel polysilicon 1199 -3411 1199 -3411 0 3
rlabel polysilicon 1206 -3405 1206 -3405 0 1
rlabel polysilicon 1206 -3411 1206 -3411 0 3
rlabel polysilicon 1213 -3405 1213 -3405 0 1
rlabel polysilicon 1213 -3411 1213 -3411 0 3
rlabel polysilicon 1216 -3411 1216 -3411 0 4
rlabel polysilicon 1234 -3405 1234 -3405 0 1
rlabel polysilicon 1234 -3411 1234 -3411 0 3
rlabel polysilicon 1241 -3405 1241 -3405 0 1
rlabel polysilicon 1241 -3411 1241 -3411 0 3
rlabel polysilicon 1248 -3405 1248 -3405 0 1
rlabel polysilicon 1248 -3411 1248 -3411 0 3
rlabel polysilicon 1265 -3405 1265 -3405 0 2
rlabel polysilicon 1265 -3411 1265 -3411 0 4
rlabel polysilicon 1311 -3405 1311 -3405 0 1
rlabel polysilicon 1311 -3411 1311 -3411 0 3
rlabel polysilicon 1318 -3405 1318 -3405 0 1
rlabel polysilicon 1318 -3411 1318 -3411 0 3
rlabel polysilicon 1332 -3405 1332 -3405 0 1
rlabel polysilicon 1332 -3411 1332 -3411 0 3
rlabel polysilicon 1374 -3405 1374 -3405 0 1
rlabel polysilicon 1374 -3411 1374 -3411 0 3
rlabel polysilicon 1381 -3405 1381 -3405 0 1
rlabel polysilicon 1381 -3411 1381 -3411 0 3
rlabel polysilicon 1384 -3411 1384 -3411 0 4
rlabel polysilicon 1388 -3405 1388 -3405 0 1
rlabel polysilicon 1388 -3411 1388 -3411 0 3
rlabel polysilicon 1577 -3405 1577 -3405 0 1
rlabel polysilicon 1577 -3411 1577 -3411 0 3
rlabel polysilicon 261 -3452 261 -3452 0 1
rlabel polysilicon 261 -3458 261 -3458 0 3
rlabel polysilicon 310 -3452 310 -3452 0 1
rlabel polysilicon 310 -3458 310 -3458 0 3
rlabel polysilicon 317 -3452 317 -3452 0 1
rlabel polysilicon 317 -3458 317 -3458 0 3
rlabel polysilicon 338 -3452 338 -3452 0 1
rlabel polysilicon 338 -3458 338 -3458 0 3
rlabel polysilicon 345 -3452 345 -3452 0 1
rlabel polysilicon 345 -3458 345 -3458 0 3
rlabel polysilicon 352 -3452 352 -3452 0 1
rlabel polysilicon 355 -3452 355 -3452 0 2
rlabel polysilicon 355 -3458 355 -3458 0 4
rlabel polysilicon 359 -3452 359 -3452 0 1
rlabel polysilicon 359 -3458 359 -3458 0 3
rlabel polysilicon 366 -3452 366 -3452 0 1
rlabel polysilicon 366 -3458 366 -3458 0 3
rlabel polysilicon 373 -3452 373 -3452 0 1
rlabel polysilicon 373 -3458 373 -3458 0 3
rlabel polysilicon 380 -3452 380 -3452 0 1
rlabel polysilicon 380 -3458 380 -3458 0 3
rlabel polysilicon 387 -3452 387 -3452 0 1
rlabel polysilicon 387 -3458 387 -3458 0 3
rlabel polysilicon 394 -3452 394 -3452 0 1
rlabel polysilicon 394 -3458 394 -3458 0 3
rlabel polysilicon 401 -3452 401 -3452 0 1
rlabel polysilicon 401 -3458 401 -3458 0 3
rlabel polysilicon 411 -3458 411 -3458 0 4
rlabel polysilicon 415 -3452 415 -3452 0 1
rlabel polysilicon 415 -3458 415 -3458 0 3
rlabel polysilicon 422 -3452 422 -3452 0 1
rlabel polysilicon 422 -3458 422 -3458 0 3
rlabel polysilicon 429 -3452 429 -3452 0 1
rlabel polysilicon 429 -3458 429 -3458 0 3
rlabel polysilicon 436 -3452 436 -3452 0 1
rlabel polysilicon 436 -3458 436 -3458 0 3
rlabel polysilicon 443 -3452 443 -3452 0 1
rlabel polysilicon 443 -3458 443 -3458 0 3
rlabel polysilicon 450 -3452 450 -3452 0 1
rlabel polysilicon 450 -3458 450 -3458 0 3
rlabel polysilicon 457 -3452 457 -3452 0 1
rlabel polysilicon 457 -3458 457 -3458 0 3
rlabel polysilicon 464 -3452 464 -3452 0 1
rlabel polysilicon 464 -3458 464 -3458 0 3
rlabel polysilicon 471 -3452 471 -3452 0 1
rlabel polysilicon 474 -3452 474 -3452 0 2
rlabel polysilicon 478 -3452 478 -3452 0 1
rlabel polysilicon 478 -3458 478 -3458 0 3
rlabel polysilicon 485 -3452 485 -3452 0 1
rlabel polysilicon 485 -3458 485 -3458 0 3
rlabel polysilicon 492 -3452 492 -3452 0 1
rlabel polysilicon 492 -3458 492 -3458 0 3
rlabel polysilicon 499 -3452 499 -3452 0 1
rlabel polysilicon 499 -3458 499 -3458 0 3
rlabel polysilicon 506 -3452 506 -3452 0 1
rlabel polysilicon 509 -3452 509 -3452 0 2
rlabel polysilicon 506 -3458 506 -3458 0 3
rlabel polysilicon 513 -3452 513 -3452 0 1
rlabel polysilicon 513 -3458 513 -3458 0 3
rlabel polysilicon 520 -3452 520 -3452 0 1
rlabel polysilicon 520 -3458 520 -3458 0 3
rlabel polysilicon 527 -3452 527 -3452 0 1
rlabel polysilicon 527 -3458 527 -3458 0 3
rlabel polysilicon 534 -3452 534 -3452 0 1
rlabel polysilicon 534 -3458 534 -3458 0 3
rlabel polysilicon 541 -3452 541 -3452 0 1
rlabel polysilicon 541 -3458 541 -3458 0 3
rlabel polysilicon 548 -3452 548 -3452 0 1
rlabel polysilicon 548 -3458 548 -3458 0 3
rlabel polysilicon 555 -3452 555 -3452 0 1
rlabel polysilicon 555 -3458 555 -3458 0 3
rlabel polysilicon 562 -3452 562 -3452 0 1
rlabel polysilicon 562 -3458 562 -3458 0 3
rlabel polysilicon 569 -3452 569 -3452 0 1
rlabel polysilicon 569 -3458 569 -3458 0 3
rlabel polysilicon 576 -3452 576 -3452 0 1
rlabel polysilicon 576 -3458 576 -3458 0 3
rlabel polysilicon 583 -3452 583 -3452 0 1
rlabel polysilicon 586 -3452 586 -3452 0 2
rlabel polysilicon 583 -3458 583 -3458 0 3
rlabel polysilicon 586 -3458 586 -3458 0 4
rlabel polysilicon 590 -3458 590 -3458 0 3
rlabel polysilicon 593 -3458 593 -3458 0 4
rlabel polysilicon 597 -3452 597 -3452 0 1
rlabel polysilicon 597 -3458 597 -3458 0 3
rlabel polysilicon 604 -3452 604 -3452 0 1
rlabel polysilicon 604 -3458 604 -3458 0 3
rlabel polysilicon 607 -3458 607 -3458 0 4
rlabel polysilicon 611 -3452 611 -3452 0 1
rlabel polysilicon 611 -3458 611 -3458 0 3
rlabel polysilicon 621 -3452 621 -3452 0 2
rlabel polysilicon 618 -3458 618 -3458 0 3
rlabel polysilicon 621 -3458 621 -3458 0 4
rlabel polysilicon 625 -3452 625 -3452 0 1
rlabel polysilicon 625 -3458 625 -3458 0 3
rlabel polysilicon 632 -3452 632 -3452 0 1
rlabel polysilicon 632 -3458 632 -3458 0 3
rlabel polysilicon 639 -3452 639 -3452 0 1
rlabel polysilicon 639 -3458 639 -3458 0 3
rlabel polysilicon 646 -3452 646 -3452 0 1
rlabel polysilicon 646 -3458 646 -3458 0 3
rlabel polysilicon 656 -3452 656 -3452 0 2
rlabel polysilicon 653 -3458 653 -3458 0 3
rlabel polysilicon 660 -3452 660 -3452 0 1
rlabel polysilicon 663 -3452 663 -3452 0 2
rlabel polysilicon 660 -3458 660 -3458 0 3
rlabel polysilicon 663 -3458 663 -3458 0 4
rlabel polysilicon 667 -3452 667 -3452 0 1
rlabel polysilicon 667 -3458 667 -3458 0 3
rlabel polysilicon 674 -3452 674 -3452 0 1
rlabel polysilicon 674 -3458 674 -3458 0 3
rlabel polysilicon 681 -3452 681 -3452 0 1
rlabel polysilicon 681 -3458 681 -3458 0 3
rlabel polysilicon 688 -3452 688 -3452 0 1
rlabel polysilicon 688 -3458 688 -3458 0 3
rlabel polysilicon 695 -3452 695 -3452 0 1
rlabel polysilicon 695 -3458 695 -3458 0 3
rlabel polysilicon 702 -3452 702 -3452 0 1
rlabel polysilicon 702 -3458 702 -3458 0 3
rlabel polysilicon 709 -3452 709 -3452 0 1
rlabel polysilicon 709 -3458 709 -3458 0 3
rlabel polysilicon 716 -3452 716 -3452 0 1
rlabel polysilicon 719 -3458 719 -3458 0 4
rlabel polysilicon 723 -3452 723 -3452 0 1
rlabel polysilicon 723 -3458 723 -3458 0 3
rlabel polysilicon 730 -3452 730 -3452 0 1
rlabel polysilicon 730 -3458 730 -3458 0 3
rlabel polysilicon 737 -3452 737 -3452 0 1
rlabel polysilicon 737 -3458 737 -3458 0 3
rlabel polysilicon 744 -3452 744 -3452 0 1
rlabel polysilicon 744 -3458 744 -3458 0 3
rlabel polysilicon 751 -3452 751 -3452 0 1
rlabel polysilicon 751 -3458 751 -3458 0 3
rlabel polysilicon 758 -3452 758 -3452 0 1
rlabel polysilicon 758 -3458 758 -3458 0 3
rlabel polysilicon 765 -3452 765 -3452 0 1
rlabel polysilicon 765 -3458 765 -3458 0 3
rlabel polysilicon 772 -3452 772 -3452 0 1
rlabel polysilicon 772 -3458 772 -3458 0 3
rlabel polysilicon 779 -3452 779 -3452 0 1
rlabel polysilicon 779 -3458 779 -3458 0 3
rlabel polysilicon 786 -3452 786 -3452 0 1
rlabel polysilicon 786 -3458 786 -3458 0 3
rlabel polysilicon 793 -3452 793 -3452 0 1
rlabel polysilicon 793 -3458 793 -3458 0 3
rlabel polysilicon 800 -3452 800 -3452 0 1
rlabel polysilicon 800 -3458 800 -3458 0 3
rlabel polysilicon 807 -3452 807 -3452 0 1
rlabel polysilicon 810 -3452 810 -3452 0 2
rlabel polysilicon 807 -3458 807 -3458 0 3
rlabel polysilicon 814 -3452 814 -3452 0 1
rlabel polysilicon 814 -3458 814 -3458 0 3
rlabel polysilicon 821 -3452 821 -3452 0 1
rlabel polysilicon 824 -3452 824 -3452 0 2
rlabel polysilicon 821 -3458 821 -3458 0 3
rlabel polysilicon 828 -3452 828 -3452 0 1
rlabel polysilicon 828 -3458 828 -3458 0 3
rlabel polysilicon 835 -3452 835 -3452 0 1
rlabel polysilicon 835 -3458 835 -3458 0 3
rlabel polysilicon 842 -3452 842 -3452 0 1
rlabel polysilicon 842 -3458 842 -3458 0 3
rlabel polysilicon 849 -3452 849 -3452 0 1
rlabel polysilicon 852 -3452 852 -3452 0 2
rlabel polysilicon 852 -3458 852 -3458 0 4
rlabel polysilicon 856 -3452 856 -3452 0 1
rlabel polysilicon 856 -3458 856 -3458 0 3
rlabel polysilicon 863 -3452 863 -3452 0 1
rlabel polysilicon 863 -3458 863 -3458 0 3
rlabel polysilicon 870 -3452 870 -3452 0 1
rlabel polysilicon 870 -3458 870 -3458 0 3
rlabel polysilicon 877 -3452 877 -3452 0 1
rlabel polysilicon 877 -3458 877 -3458 0 3
rlabel polysilicon 884 -3452 884 -3452 0 1
rlabel polysilicon 884 -3458 884 -3458 0 3
rlabel polysilicon 891 -3452 891 -3452 0 1
rlabel polysilicon 891 -3458 891 -3458 0 3
rlabel polysilicon 898 -3452 898 -3452 0 1
rlabel polysilicon 898 -3458 898 -3458 0 3
rlabel polysilicon 905 -3452 905 -3452 0 1
rlabel polysilicon 905 -3458 905 -3458 0 3
rlabel polysilicon 912 -3452 912 -3452 0 1
rlabel polysilicon 912 -3458 912 -3458 0 3
rlabel polysilicon 919 -3452 919 -3452 0 1
rlabel polysilicon 919 -3458 919 -3458 0 3
rlabel polysilicon 926 -3452 926 -3452 0 1
rlabel polysilicon 926 -3458 926 -3458 0 3
rlabel polysilicon 933 -3452 933 -3452 0 1
rlabel polysilicon 933 -3458 933 -3458 0 3
rlabel polysilicon 940 -3452 940 -3452 0 1
rlabel polysilicon 940 -3458 940 -3458 0 3
rlabel polysilicon 947 -3452 947 -3452 0 1
rlabel polysilicon 947 -3458 947 -3458 0 3
rlabel polysilicon 954 -3452 954 -3452 0 1
rlabel polysilicon 961 -3452 961 -3452 0 1
rlabel polysilicon 961 -3458 961 -3458 0 3
rlabel polysilicon 968 -3458 968 -3458 0 3
rlabel polysilicon 975 -3452 975 -3452 0 1
rlabel polysilicon 975 -3458 975 -3458 0 3
rlabel polysilicon 982 -3452 982 -3452 0 1
rlabel polysilicon 982 -3458 982 -3458 0 3
rlabel polysilicon 989 -3452 989 -3452 0 1
rlabel polysilicon 989 -3458 989 -3458 0 3
rlabel polysilicon 996 -3452 996 -3452 0 1
rlabel polysilicon 999 -3452 999 -3452 0 2
rlabel polysilicon 996 -3458 996 -3458 0 3
rlabel polysilicon 1003 -3452 1003 -3452 0 1
rlabel polysilicon 1003 -3458 1003 -3458 0 3
rlabel polysilicon 1010 -3452 1010 -3452 0 1
rlabel polysilicon 1010 -3458 1010 -3458 0 3
rlabel polysilicon 1017 -3452 1017 -3452 0 1
rlabel polysilicon 1017 -3458 1017 -3458 0 3
rlabel polysilicon 1024 -3452 1024 -3452 0 1
rlabel polysilicon 1024 -3458 1024 -3458 0 3
rlabel polysilicon 1031 -3452 1031 -3452 0 1
rlabel polysilicon 1031 -3458 1031 -3458 0 3
rlabel polysilicon 1052 -3452 1052 -3452 0 1
rlabel polysilicon 1052 -3458 1052 -3458 0 3
rlabel polysilicon 1073 -3452 1073 -3452 0 1
rlabel polysilicon 1073 -3458 1073 -3458 0 3
rlabel polysilicon 1080 -3452 1080 -3452 0 1
rlabel polysilicon 1080 -3458 1080 -3458 0 3
rlabel polysilicon 1101 -3452 1101 -3452 0 1
rlabel polysilicon 1101 -3458 1101 -3458 0 3
rlabel polysilicon 1115 -3452 1115 -3452 0 1
rlabel polysilicon 1115 -3458 1115 -3458 0 3
rlabel polysilicon 1118 -3458 1118 -3458 0 4
rlabel polysilicon 1122 -3452 1122 -3452 0 1
rlabel polysilicon 1122 -3458 1122 -3458 0 3
rlabel polysilicon 1129 -3452 1129 -3452 0 1
rlabel polysilicon 1129 -3458 1129 -3458 0 3
rlabel polysilicon 1136 -3452 1136 -3452 0 1
rlabel polysilicon 1136 -3458 1136 -3458 0 3
rlabel polysilicon 1143 -3458 1143 -3458 0 3
rlabel polysilicon 1192 -3452 1192 -3452 0 1
rlabel polysilicon 1192 -3458 1192 -3458 0 3
rlabel polysilicon 1199 -3452 1199 -3452 0 1
rlabel polysilicon 1199 -3458 1199 -3458 0 3
rlabel polysilicon 1206 -3452 1206 -3452 0 1
rlabel polysilicon 1206 -3458 1206 -3458 0 3
rlabel polysilicon 1213 -3452 1213 -3452 0 1
rlabel polysilicon 1213 -3458 1213 -3458 0 3
rlabel polysilicon 1269 -3452 1269 -3452 0 1
rlabel polysilicon 1269 -3458 1269 -3458 0 3
rlabel polysilicon 1300 -3452 1300 -3452 0 2
rlabel polysilicon 1297 -3458 1297 -3458 0 3
rlabel polysilicon 1300 -3458 1300 -3458 0 4
rlabel polysilicon 1304 -3452 1304 -3452 0 1
rlabel polysilicon 1304 -3458 1304 -3458 0 3
rlabel polysilicon 1318 -3452 1318 -3452 0 1
rlabel polysilicon 1318 -3458 1318 -3458 0 3
rlabel polysilicon 1346 -3452 1346 -3452 0 1
rlabel polysilicon 1346 -3458 1346 -3458 0 3
rlabel polysilicon 1381 -3452 1381 -3452 0 1
rlabel polysilicon 1384 -3452 1384 -3452 0 2
rlabel polysilicon 1381 -3458 1381 -3458 0 3
rlabel polysilicon 1388 -3452 1388 -3452 0 1
rlabel polysilicon 1388 -3458 1388 -3458 0 3
rlabel polysilicon 1395 -3452 1395 -3452 0 1
rlabel polysilicon 1395 -3458 1395 -3458 0 3
rlabel polysilicon 1577 -3452 1577 -3452 0 1
rlabel polysilicon 1577 -3458 1577 -3458 0 3
rlabel polysilicon 268 -3493 268 -3493 0 1
rlabel polysilicon 268 -3499 268 -3499 0 3
rlabel polysilicon 282 -3499 282 -3499 0 3
rlabel polysilicon 285 -3499 285 -3499 0 4
rlabel polysilicon 296 -3493 296 -3493 0 1
rlabel polysilicon 296 -3499 296 -3499 0 3
rlabel polysilicon 366 -3493 366 -3493 0 1
rlabel polysilicon 366 -3499 366 -3499 0 3
rlabel polysilicon 373 -3493 373 -3493 0 1
rlabel polysilicon 373 -3499 373 -3499 0 3
rlabel polysilicon 380 -3493 380 -3493 0 1
rlabel polysilicon 380 -3499 380 -3499 0 3
rlabel polysilicon 390 -3493 390 -3493 0 2
rlabel polysilicon 390 -3499 390 -3499 0 4
rlabel polysilicon 408 -3493 408 -3493 0 1
rlabel polysilicon 408 -3499 408 -3499 0 3
rlabel polysilicon 422 -3493 422 -3493 0 1
rlabel polysilicon 425 -3493 425 -3493 0 2
rlabel polysilicon 429 -3493 429 -3493 0 1
rlabel polysilicon 429 -3499 429 -3499 0 3
rlabel polysilicon 439 -3493 439 -3493 0 2
rlabel polysilicon 439 -3499 439 -3499 0 4
rlabel polysilicon 443 -3493 443 -3493 0 1
rlabel polysilicon 443 -3499 443 -3499 0 3
rlabel polysilicon 450 -3493 450 -3493 0 1
rlabel polysilicon 450 -3499 450 -3499 0 3
rlabel polysilicon 457 -3493 457 -3493 0 1
rlabel polysilicon 457 -3499 457 -3499 0 3
rlabel polysilicon 471 -3493 471 -3493 0 1
rlabel polysilicon 471 -3499 471 -3499 0 3
rlabel polysilicon 478 -3493 478 -3493 0 1
rlabel polysilicon 478 -3499 478 -3499 0 3
rlabel polysilicon 485 -3493 485 -3493 0 1
rlabel polysilicon 485 -3499 485 -3499 0 3
rlabel polysilicon 492 -3493 492 -3493 0 1
rlabel polysilicon 492 -3499 492 -3499 0 3
rlabel polysilicon 499 -3493 499 -3493 0 1
rlabel polysilicon 499 -3499 499 -3499 0 3
rlabel polysilicon 506 -3493 506 -3493 0 1
rlabel polysilicon 506 -3499 506 -3499 0 3
rlabel polysilicon 513 -3493 513 -3493 0 1
rlabel polysilicon 513 -3499 513 -3499 0 3
rlabel polysilicon 527 -3493 527 -3493 0 1
rlabel polysilicon 527 -3499 527 -3499 0 3
rlabel polysilicon 534 -3493 534 -3493 0 1
rlabel polysilicon 534 -3499 534 -3499 0 3
rlabel polysilicon 541 -3493 541 -3493 0 1
rlabel polysilicon 541 -3499 541 -3499 0 3
rlabel polysilicon 548 -3493 548 -3493 0 1
rlabel polysilicon 548 -3499 548 -3499 0 3
rlabel polysilicon 555 -3493 555 -3493 0 1
rlabel polysilicon 555 -3499 555 -3499 0 3
rlabel polysilicon 562 -3493 562 -3493 0 1
rlabel polysilicon 562 -3499 562 -3499 0 3
rlabel polysilicon 569 -3493 569 -3493 0 1
rlabel polysilicon 569 -3499 569 -3499 0 3
rlabel polysilicon 576 -3493 576 -3493 0 1
rlabel polysilicon 576 -3499 576 -3499 0 3
rlabel polysilicon 583 -3493 583 -3493 0 1
rlabel polysilicon 583 -3499 583 -3499 0 3
rlabel polysilicon 590 -3493 590 -3493 0 1
rlabel polysilicon 590 -3499 590 -3499 0 3
rlabel polysilicon 604 -3493 604 -3493 0 1
rlabel polysilicon 604 -3499 604 -3499 0 3
rlabel polysilicon 618 -3493 618 -3493 0 1
rlabel polysilicon 618 -3499 618 -3499 0 3
rlabel polysilicon 632 -3493 632 -3493 0 1
rlabel polysilicon 632 -3499 632 -3499 0 3
rlabel polysilicon 639 -3493 639 -3493 0 1
rlabel polysilicon 639 -3499 639 -3499 0 3
rlabel polysilicon 646 -3493 646 -3493 0 1
rlabel polysilicon 646 -3499 646 -3499 0 3
rlabel polysilicon 653 -3493 653 -3493 0 1
rlabel polysilicon 656 -3493 656 -3493 0 2
rlabel polysilicon 656 -3499 656 -3499 0 4
rlabel polysilicon 688 -3493 688 -3493 0 1
rlabel polysilicon 688 -3499 688 -3499 0 3
rlabel polysilicon 695 -3493 695 -3493 0 1
rlabel polysilicon 695 -3499 695 -3499 0 3
rlabel polysilicon 702 -3493 702 -3493 0 1
rlabel polysilicon 702 -3499 702 -3499 0 3
rlabel polysilicon 709 -3493 709 -3493 0 1
rlabel polysilicon 709 -3499 709 -3499 0 3
rlabel polysilicon 716 -3493 716 -3493 0 1
rlabel polysilicon 716 -3499 716 -3499 0 3
rlabel polysilicon 723 -3493 723 -3493 0 1
rlabel polysilicon 726 -3499 726 -3499 0 4
rlabel polysilicon 730 -3493 730 -3493 0 1
rlabel polysilicon 733 -3493 733 -3493 0 2
rlabel polysilicon 730 -3499 730 -3499 0 3
rlabel polysilicon 733 -3499 733 -3499 0 4
rlabel polysilicon 737 -3493 737 -3493 0 1
rlabel polysilicon 737 -3499 737 -3499 0 3
rlabel polysilicon 744 -3493 744 -3493 0 1
rlabel polysilicon 744 -3499 744 -3499 0 3
rlabel polysilicon 754 -3493 754 -3493 0 2
rlabel polysilicon 754 -3499 754 -3499 0 4
rlabel polysilicon 758 -3493 758 -3493 0 1
rlabel polysilicon 758 -3499 758 -3499 0 3
rlabel polysilicon 765 -3493 765 -3493 0 1
rlabel polysilicon 765 -3499 765 -3499 0 3
rlabel polysilicon 772 -3493 772 -3493 0 1
rlabel polysilicon 772 -3499 772 -3499 0 3
rlabel polysilicon 786 -3493 786 -3493 0 1
rlabel polysilicon 786 -3499 786 -3499 0 3
rlabel polysilicon 793 -3493 793 -3493 0 1
rlabel polysilicon 800 -3493 800 -3493 0 1
rlabel polysilicon 800 -3499 800 -3499 0 3
rlabel polysilicon 807 -3493 807 -3493 0 1
rlabel polysilicon 807 -3499 807 -3499 0 3
rlabel polysilicon 814 -3493 814 -3493 0 1
rlabel polysilicon 814 -3499 814 -3499 0 3
rlabel polysilicon 821 -3493 821 -3493 0 1
rlabel polysilicon 821 -3499 821 -3499 0 3
rlabel polysilicon 828 -3493 828 -3493 0 1
rlabel polysilicon 828 -3499 828 -3499 0 3
rlabel polysilicon 877 -3493 877 -3493 0 1
rlabel polysilicon 877 -3499 877 -3499 0 3
rlabel polysilicon 884 -3493 884 -3493 0 1
rlabel polysilicon 884 -3499 884 -3499 0 3
rlabel polysilicon 891 -3493 891 -3493 0 1
rlabel polysilicon 891 -3499 891 -3499 0 3
rlabel polysilicon 898 -3493 898 -3493 0 1
rlabel polysilicon 898 -3499 898 -3499 0 3
rlabel polysilicon 905 -3493 905 -3493 0 1
rlabel polysilicon 905 -3499 905 -3499 0 3
rlabel polysilicon 912 -3493 912 -3493 0 1
rlabel polysilicon 915 -3493 915 -3493 0 2
rlabel polysilicon 912 -3499 912 -3499 0 3
rlabel polysilicon 919 -3493 919 -3493 0 1
rlabel polysilicon 919 -3499 919 -3499 0 3
rlabel polysilicon 926 -3493 926 -3493 0 1
rlabel polysilicon 926 -3499 926 -3499 0 3
rlabel polysilicon 933 -3493 933 -3493 0 1
rlabel polysilicon 933 -3499 933 -3499 0 3
rlabel polysilicon 940 -3493 940 -3493 0 1
rlabel polysilicon 940 -3499 940 -3499 0 3
rlabel polysilicon 947 -3493 947 -3493 0 1
rlabel polysilicon 947 -3499 947 -3499 0 3
rlabel polysilicon 954 -3499 954 -3499 0 3
rlabel polysilicon 961 -3493 961 -3493 0 1
rlabel polysilicon 961 -3499 961 -3499 0 3
rlabel polysilicon 975 -3493 975 -3493 0 1
rlabel polysilicon 975 -3499 975 -3499 0 3
rlabel polysilicon 996 -3493 996 -3493 0 1
rlabel polysilicon 996 -3499 996 -3499 0 3
rlabel polysilicon 1003 -3493 1003 -3493 0 1
rlabel polysilicon 1006 -3493 1006 -3493 0 2
rlabel polysilicon 1003 -3499 1003 -3499 0 3
rlabel polysilicon 1010 -3493 1010 -3493 0 1
rlabel polysilicon 1010 -3499 1010 -3499 0 3
rlabel polysilicon 1024 -3493 1024 -3493 0 1
rlabel polysilicon 1024 -3499 1024 -3499 0 3
rlabel polysilicon 1038 -3493 1038 -3493 0 1
rlabel polysilicon 1038 -3499 1038 -3499 0 3
rlabel polysilicon 1045 -3493 1045 -3493 0 1
rlabel polysilicon 1045 -3499 1045 -3499 0 3
rlabel polysilicon 1048 -3499 1048 -3499 0 4
rlabel polysilicon 1052 -3493 1052 -3493 0 1
rlabel polysilicon 1052 -3499 1052 -3499 0 3
rlabel polysilicon 1059 -3493 1059 -3493 0 1
rlabel polysilicon 1059 -3499 1059 -3499 0 3
rlabel polysilicon 1066 -3493 1066 -3493 0 1
rlabel polysilicon 1066 -3499 1066 -3499 0 3
rlabel polysilicon 1073 -3493 1073 -3493 0 1
rlabel polysilicon 1073 -3499 1073 -3499 0 3
rlabel polysilicon 1080 -3493 1080 -3493 0 1
rlabel polysilicon 1080 -3499 1080 -3499 0 3
rlabel polysilicon 1087 -3493 1087 -3493 0 1
rlabel polysilicon 1090 -3493 1090 -3493 0 2
rlabel polysilicon 1090 -3499 1090 -3499 0 4
rlabel polysilicon 1115 -3493 1115 -3493 0 1
rlabel polysilicon 1118 -3493 1118 -3493 0 2
rlabel polysilicon 1115 -3499 1115 -3499 0 3
rlabel polysilicon 1122 -3493 1122 -3493 0 1
rlabel polysilicon 1122 -3499 1122 -3499 0 3
rlabel polysilicon 1136 -3493 1136 -3493 0 1
rlabel polysilicon 1136 -3499 1136 -3499 0 3
rlabel polysilicon 1157 -3493 1157 -3493 0 1
rlabel polysilicon 1157 -3499 1157 -3499 0 3
rlabel polysilicon 1178 -3493 1178 -3493 0 1
rlabel polysilicon 1181 -3493 1181 -3493 0 2
rlabel polysilicon 1181 -3499 1181 -3499 0 4
rlabel polysilicon 1185 -3493 1185 -3493 0 1
rlabel polysilicon 1185 -3499 1185 -3499 0 3
rlabel polysilicon 1192 -3493 1192 -3493 0 1
rlabel polysilicon 1192 -3499 1192 -3499 0 3
rlabel polysilicon 1234 -3493 1234 -3493 0 1
rlabel polysilicon 1234 -3499 1234 -3499 0 3
rlabel polysilicon 1248 -3493 1248 -3493 0 1
rlabel polysilicon 1248 -3499 1248 -3499 0 3
rlabel polysilicon 1269 -3493 1269 -3493 0 1
rlabel polysilicon 1269 -3499 1269 -3499 0 3
rlabel polysilicon 1276 -3493 1276 -3493 0 1
rlabel polysilicon 1276 -3499 1276 -3499 0 3
rlabel polysilicon 1374 -3493 1374 -3493 0 1
rlabel polysilicon 1374 -3499 1374 -3499 0 3
rlabel polysilicon 1381 -3493 1381 -3493 0 1
rlabel polysilicon 1384 -3499 1384 -3499 0 4
rlabel polysilicon 1388 -3493 1388 -3493 0 1
rlabel polysilicon 1388 -3499 1388 -3499 0 3
rlabel polysilicon 1395 -3493 1395 -3493 0 1
rlabel polysilicon 1395 -3499 1395 -3499 0 3
rlabel polysilicon 1416 -3493 1416 -3493 0 1
rlabel polysilicon 1416 -3499 1416 -3499 0 3
rlabel polysilicon 1577 -3493 1577 -3493 0 1
rlabel polysilicon 1577 -3499 1577 -3499 0 3
rlabel polysilicon 380 -3524 380 -3524 0 1
rlabel polysilicon 380 -3530 380 -3530 0 3
rlabel polysilicon 387 -3524 387 -3524 0 1
rlabel polysilicon 387 -3530 387 -3530 0 3
rlabel polysilicon 394 -3524 394 -3524 0 1
rlabel polysilicon 394 -3530 394 -3530 0 3
rlabel polysilicon 401 -3524 401 -3524 0 1
rlabel polysilicon 401 -3530 401 -3530 0 3
rlabel polysilicon 429 -3524 429 -3524 0 1
rlabel polysilicon 429 -3530 429 -3530 0 3
rlabel polysilicon 443 -3524 443 -3524 0 1
rlabel polysilicon 443 -3530 443 -3530 0 3
rlabel polysilicon 450 -3524 450 -3524 0 1
rlabel polysilicon 450 -3530 450 -3530 0 3
rlabel polysilicon 464 -3524 464 -3524 0 1
rlabel polysilicon 464 -3530 464 -3530 0 3
rlabel polysilicon 478 -3524 478 -3524 0 1
rlabel polysilicon 481 -3524 481 -3524 0 2
rlabel polysilicon 478 -3530 478 -3530 0 3
rlabel polysilicon 485 -3524 485 -3524 0 1
rlabel polysilicon 485 -3530 485 -3530 0 3
rlabel polysilicon 492 -3524 492 -3524 0 1
rlabel polysilicon 492 -3530 492 -3530 0 3
rlabel polysilicon 499 -3524 499 -3524 0 1
rlabel polysilicon 499 -3530 499 -3530 0 3
rlabel polysilicon 506 -3524 506 -3524 0 1
rlabel polysilicon 506 -3530 506 -3530 0 3
rlabel polysilicon 513 -3524 513 -3524 0 1
rlabel polysilicon 513 -3530 513 -3530 0 3
rlabel polysilicon 520 -3524 520 -3524 0 1
rlabel polysilicon 520 -3530 520 -3530 0 3
rlabel polysilicon 527 -3524 527 -3524 0 1
rlabel polysilicon 527 -3530 527 -3530 0 3
rlabel polysilicon 534 -3524 534 -3524 0 1
rlabel polysilicon 534 -3530 534 -3530 0 3
rlabel polysilicon 541 -3524 541 -3524 0 1
rlabel polysilicon 541 -3530 541 -3530 0 3
rlabel polysilicon 548 -3524 548 -3524 0 1
rlabel polysilicon 548 -3530 548 -3530 0 3
rlabel polysilicon 558 -3524 558 -3524 0 2
rlabel polysilicon 555 -3530 555 -3530 0 3
rlabel polysilicon 558 -3530 558 -3530 0 4
rlabel polysilicon 565 -3524 565 -3524 0 2
rlabel polysilicon 562 -3530 562 -3530 0 3
rlabel polysilicon 565 -3530 565 -3530 0 4
rlabel polysilicon 569 -3524 569 -3524 0 1
rlabel polysilicon 569 -3530 569 -3530 0 3
rlabel polysilicon 576 -3524 576 -3524 0 1
rlabel polysilicon 576 -3530 576 -3530 0 3
rlabel polysilicon 583 -3524 583 -3524 0 1
rlabel polysilicon 583 -3530 583 -3530 0 3
rlabel polysilicon 590 -3524 590 -3524 0 1
rlabel polysilicon 590 -3530 590 -3530 0 3
rlabel polysilicon 597 -3524 597 -3524 0 1
rlabel polysilicon 597 -3530 597 -3530 0 3
rlabel polysilicon 604 -3524 604 -3524 0 1
rlabel polysilicon 604 -3530 604 -3530 0 3
rlabel polysilicon 646 -3524 646 -3524 0 1
rlabel polysilicon 646 -3530 646 -3530 0 3
rlabel polysilicon 653 -3524 653 -3524 0 1
rlabel polysilicon 653 -3530 653 -3530 0 3
rlabel polysilicon 674 -3524 674 -3524 0 1
rlabel polysilicon 674 -3530 674 -3530 0 3
rlabel polysilicon 695 -3524 695 -3524 0 1
rlabel polysilicon 695 -3530 695 -3530 0 3
rlabel polysilicon 702 -3524 702 -3524 0 1
rlabel polysilicon 702 -3530 702 -3530 0 3
rlabel polysilicon 709 -3524 709 -3524 0 1
rlabel polysilicon 709 -3530 709 -3530 0 3
rlabel polysilicon 730 -3524 730 -3524 0 1
rlabel polysilicon 730 -3530 730 -3530 0 3
rlabel polysilicon 758 -3524 758 -3524 0 1
rlabel polysilicon 758 -3530 758 -3530 0 3
rlabel polysilicon 765 -3524 765 -3524 0 1
rlabel polysilicon 765 -3530 765 -3530 0 3
rlabel polysilicon 772 -3524 772 -3524 0 1
rlabel polysilicon 772 -3530 772 -3530 0 3
rlabel polysilicon 779 -3524 779 -3524 0 1
rlabel polysilicon 779 -3530 779 -3530 0 3
rlabel polysilicon 786 -3524 786 -3524 0 1
rlabel polysilicon 786 -3530 786 -3530 0 3
rlabel polysilicon 793 -3530 793 -3530 0 3
rlabel polysilicon 800 -3524 800 -3524 0 1
rlabel polysilicon 800 -3530 800 -3530 0 3
rlabel polysilicon 807 -3524 807 -3524 0 1
rlabel polysilicon 807 -3530 807 -3530 0 3
rlabel polysilicon 814 -3524 814 -3524 0 1
rlabel polysilicon 814 -3530 814 -3530 0 3
rlabel polysilicon 821 -3524 821 -3524 0 1
rlabel polysilicon 824 -3530 824 -3530 0 4
rlabel polysilicon 842 -3524 842 -3524 0 1
rlabel polysilicon 842 -3530 842 -3530 0 3
rlabel polysilicon 863 -3524 863 -3524 0 1
rlabel polysilicon 863 -3530 863 -3530 0 3
rlabel polysilicon 877 -3524 877 -3524 0 1
rlabel polysilicon 877 -3530 877 -3530 0 3
rlabel polysilicon 884 -3524 884 -3524 0 1
rlabel polysilicon 884 -3530 884 -3530 0 3
rlabel polysilicon 891 -3530 891 -3530 0 3
rlabel polysilicon 898 -3524 898 -3524 0 1
rlabel polysilicon 898 -3530 898 -3530 0 3
rlabel polysilicon 905 -3524 905 -3524 0 1
rlabel polysilicon 905 -3530 905 -3530 0 3
rlabel polysilicon 919 -3524 919 -3524 0 1
rlabel polysilicon 919 -3530 919 -3530 0 3
rlabel polysilicon 926 -3524 926 -3524 0 1
rlabel polysilicon 926 -3530 926 -3530 0 3
rlabel polysilicon 933 -3524 933 -3524 0 1
rlabel polysilicon 933 -3530 933 -3530 0 3
rlabel polysilicon 940 -3524 940 -3524 0 1
rlabel polysilicon 940 -3530 940 -3530 0 3
rlabel polysilicon 947 -3524 947 -3524 0 1
rlabel polysilicon 950 -3530 950 -3530 0 4
rlabel polysilicon 954 -3524 954 -3524 0 1
rlabel polysilicon 957 -3524 957 -3524 0 2
rlabel polysilicon 957 -3530 957 -3530 0 4
rlabel polysilicon 961 -3524 961 -3524 0 1
rlabel polysilicon 964 -3524 964 -3524 0 2
rlabel polysilicon 968 -3524 968 -3524 0 1
rlabel polysilicon 968 -3530 968 -3530 0 3
rlabel polysilicon 1003 -3524 1003 -3524 0 1
rlabel polysilicon 1017 -3524 1017 -3524 0 1
rlabel polysilicon 1020 -3524 1020 -3524 0 2
rlabel polysilicon 1031 -3524 1031 -3524 0 1
rlabel polysilicon 1034 -3524 1034 -3524 0 2
rlabel polysilicon 1038 -3524 1038 -3524 0 1
rlabel polysilicon 1041 -3524 1041 -3524 0 2
rlabel polysilicon 1038 -3530 1038 -3530 0 3
rlabel polysilicon 1045 -3524 1045 -3524 0 1
rlabel polysilicon 1048 -3524 1048 -3524 0 2
rlabel polysilicon 1045 -3530 1045 -3530 0 3
rlabel polysilicon 1052 -3524 1052 -3524 0 1
rlabel polysilicon 1052 -3530 1052 -3530 0 3
rlabel polysilicon 1062 -3524 1062 -3524 0 2
rlabel polysilicon 1059 -3530 1059 -3530 0 3
rlabel polysilicon 1073 -3524 1073 -3524 0 1
rlabel polysilicon 1073 -3530 1073 -3530 0 3
rlabel polysilicon 1115 -3524 1115 -3524 0 1
rlabel polysilicon 1115 -3530 1115 -3530 0 3
rlabel polysilicon 1129 -3524 1129 -3524 0 1
rlabel polysilicon 1129 -3530 1129 -3530 0 3
rlabel polysilicon 1136 -3524 1136 -3524 0 1
rlabel polysilicon 1136 -3530 1136 -3530 0 3
rlabel polysilicon 1143 -3524 1143 -3524 0 1
rlabel polysilicon 1143 -3530 1143 -3530 0 3
rlabel polysilicon 1157 -3530 1157 -3530 0 3
rlabel polysilicon 1164 -3524 1164 -3524 0 1
rlabel polysilicon 1164 -3530 1164 -3530 0 3
rlabel polysilicon 1178 -3524 1178 -3524 0 1
rlabel polysilicon 1178 -3530 1178 -3530 0 3
rlabel polysilicon 1192 -3524 1192 -3524 0 1
rlabel polysilicon 1192 -3530 1192 -3530 0 3
rlabel polysilicon 1262 -3524 1262 -3524 0 1
rlabel polysilicon 1262 -3530 1262 -3530 0 3
rlabel polysilicon 1276 -3524 1276 -3524 0 1
rlabel polysilicon 1279 -3524 1279 -3524 0 2
rlabel polysilicon 1279 -3530 1279 -3530 0 4
rlabel polysilicon 1339 -3524 1339 -3524 0 1
rlabel polysilicon 1339 -3530 1339 -3530 0 3
rlabel polysilicon 1381 -3524 1381 -3524 0 1
rlabel polysilicon 1381 -3530 1381 -3530 0 3
rlabel polysilicon 1395 -3524 1395 -3524 0 1
rlabel polysilicon 1395 -3530 1395 -3530 0 3
rlabel polysilicon 1500 -3524 1500 -3524 0 1
rlabel polysilicon 1500 -3530 1500 -3530 0 3
rlabel polysilicon 1577 -3524 1577 -3524 0 1
rlabel polysilicon 1580 -3530 1580 -3530 0 4
rlabel polysilicon 380 -3553 380 -3553 0 1
rlabel polysilicon 380 -3559 380 -3559 0 3
rlabel polysilicon 387 -3553 387 -3553 0 1
rlabel polysilicon 387 -3559 387 -3559 0 3
rlabel polysilicon 394 -3553 394 -3553 0 1
rlabel polysilicon 394 -3559 394 -3559 0 3
rlabel polysilicon 401 -3553 401 -3553 0 1
rlabel polysilicon 401 -3559 401 -3559 0 3
rlabel polysilicon 408 -3553 408 -3553 0 1
rlabel polysilicon 408 -3559 408 -3559 0 3
rlabel polysilicon 450 -3553 450 -3553 0 1
rlabel polysilicon 450 -3559 450 -3559 0 3
rlabel polysilicon 457 -3553 457 -3553 0 1
rlabel polysilicon 457 -3559 457 -3559 0 3
rlabel polysilicon 474 -3553 474 -3553 0 2
rlabel polysilicon 474 -3559 474 -3559 0 4
rlabel polysilicon 478 -3553 478 -3553 0 1
rlabel polysilicon 478 -3559 478 -3559 0 3
rlabel polysilicon 492 -3553 492 -3553 0 1
rlabel polysilicon 492 -3559 492 -3559 0 3
rlabel polysilicon 499 -3553 499 -3553 0 1
rlabel polysilicon 502 -3559 502 -3559 0 4
rlabel polysilicon 506 -3553 506 -3553 0 1
rlabel polysilicon 506 -3559 506 -3559 0 3
rlabel polysilicon 513 -3553 513 -3553 0 1
rlabel polysilicon 513 -3559 513 -3559 0 3
rlabel polysilicon 527 -3553 527 -3553 0 1
rlabel polysilicon 527 -3559 527 -3559 0 3
rlabel polysilicon 530 -3559 530 -3559 0 4
rlabel polysilicon 534 -3553 534 -3553 0 1
rlabel polysilicon 534 -3559 534 -3559 0 3
rlabel polysilicon 541 -3553 541 -3553 0 1
rlabel polysilicon 541 -3559 541 -3559 0 3
rlabel polysilicon 548 -3553 548 -3553 0 1
rlabel polysilicon 548 -3559 548 -3559 0 3
rlabel polysilicon 555 -3553 555 -3553 0 1
rlabel polysilicon 555 -3559 555 -3559 0 3
rlabel polysilicon 565 -3553 565 -3553 0 2
rlabel polysilicon 562 -3559 562 -3559 0 3
rlabel polysilicon 569 -3553 569 -3553 0 1
rlabel polysilicon 569 -3559 569 -3559 0 3
rlabel polysilicon 576 -3553 576 -3553 0 1
rlabel polysilicon 576 -3559 576 -3559 0 3
rlabel polysilicon 579 -3559 579 -3559 0 4
rlabel polysilicon 583 -3553 583 -3553 0 1
rlabel polysilicon 583 -3559 583 -3559 0 3
rlabel polysilicon 590 -3553 590 -3553 0 1
rlabel polysilicon 590 -3559 590 -3559 0 3
rlabel polysilicon 597 -3553 597 -3553 0 1
rlabel polysilicon 597 -3559 597 -3559 0 3
rlabel polysilicon 607 -3553 607 -3553 0 2
rlabel polysilicon 660 -3553 660 -3553 0 1
rlabel polysilicon 663 -3553 663 -3553 0 2
rlabel polysilicon 667 -3553 667 -3553 0 1
rlabel polysilicon 667 -3559 667 -3559 0 3
rlabel polysilicon 702 -3553 702 -3553 0 1
rlabel polysilicon 705 -3553 705 -3553 0 2
rlabel polysilicon 702 -3559 702 -3559 0 3
rlabel polysilicon 709 -3553 709 -3553 0 1
rlabel polysilicon 709 -3559 709 -3559 0 3
rlabel polysilicon 737 -3553 737 -3553 0 1
rlabel polysilicon 737 -3559 737 -3559 0 3
rlabel polysilicon 758 -3553 758 -3553 0 1
rlabel polysilicon 758 -3559 758 -3559 0 3
rlabel polysilicon 765 -3559 765 -3559 0 3
rlabel polysilicon 768 -3559 768 -3559 0 4
rlabel polysilicon 772 -3553 772 -3553 0 1
rlabel polysilicon 772 -3559 772 -3559 0 3
rlabel polysilicon 779 -3553 779 -3553 0 1
rlabel polysilicon 779 -3559 779 -3559 0 3
rlabel polysilicon 786 -3553 786 -3553 0 1
rlabel polysilicon 786 -3559 786 -3559 0 3
rlabel polysilicon 796 -3553 796 -3553 0 2
rlabel polysilicon 793 -3559 793 -3559 0 3
rlabel polysilicon 796 -3559 796 -3559 0 4
rlabel polysilicon 800 -3553 800 -3553 0 1
rlabel polysilicon 800 -3559 800 -3559 0 3
rlabel polysilicon 807 -3553 807 -3553 0 1
rlabel polysilicon 807 -3559 807 -3559 0 3
rlabel polysilicon 814 -3553 814 -3553 0 1
rlabel polysilicon 814 -3559 814 -3559 0 3
rlabel polysilicon 877 -3553 877 -3553 0 1
rlabel polysilicon 877 -3559 877 -3559 0 3
rlabel polysilicon 884 -3553 884 -3553 0 1
rlabel polysilicon 884 -3559 884 -3559 0 3
rlabel polysilicon 898 -3553 898 -3553 0 1
rlabel polysilicon 898 -3559 898 -3559 0 3
rlabel polysilicon 905 -3553 905 -3553 0 1
rlabel polysilicon 905 -3559 905 -3559 0 3
rlabel polysilicon 926 -3553 926 -3553 0 1
rlabel polysilicon 926 -3559 926 -3559 0 3
rlabel polysilicon 936 -3553 936 -3553 0 2
rlabel polysilicon 933 -3559 933 -3559 0 3
rlabel polysilicon 940 -3553 940 -3553 0 1
rlabel polysilicon 940 -3559 940 -3559 0 3
rlabel polysilicon 950 -3559 950 -3559 0 4
rlabel polysilicon 1108 -3553 1108 -3553 0 1
rlabel polysilicon 1111 -3553 1111 -3553 0 2
rlabel polysilicon 1111 -3559 1111 -3559 0 4
rlabel polysilicon 1115 -3553 1115 -3553 0 1
rlabel polysilicon 1115 -3559 1115 -3559 0 3
rlabel polysilicon 1129 -3553 1129 -3553 0 1
rlabel polysilicon 1129 -3559 1129 -3559 0 3
rlabel polysilicon 1136 -3553 1136 -3553 0 1
rlabel polysilicon 1136 -3559 1136 -3559 0 3
rlabel polysilicon 1164 -3553 1164 -3553 0 1
rlabel polysilicon 1164 -3559 1164 -3559 0 3
rlabel polysilicon 1178 -3553 1178 -3553 0 1
rlabel polysilicon 1178 -3559 1178 -3559 0 3
rlabel polysilicon 1192 -3553 1192 -3553 0 1
rlabel polysilicon 1192 -3559 1192 -3559 0 3
rlabel polysilicon 1360 -3553 1360 -3553 0 1
rlabel polysilicon 1360 -3559 1360 -3559 0 3
rlabel polysilicon 1388 -3553 1388 -3553 0 1
rlabel polysilicon 1388 -3559 1388 -3559 0 3
rlabel polysilicon 1395 -3553 1395 -3553 0 1
rlabel polysilicon 1395 -3559 1395 -3559 0 3
rlabel polysilicon 387 -3568 387 -3568 0 1
rlabel polysilicon 387 -3574 387 -3574 0 3
rlabel polysilicon 394 -3568 394 -3568 0 1
rlabel polysilicon 397 -3574 397 -3574 0 4
rlabel polysilicon 401 -3568 401 -3568 0 1
rlabel polysilicon 404 -3568 404 -3568 0 2
rlabel polysilicon 401 -3574 401 -3574 0 3
rlabel polysilicon 408 -3568 408 -3568 0 1
rlabel polysilicon 408 -3574 408 -3574 0 3
rlabel polysilicon 457 -3568 457 -3568 0 1
rlabel polysilicon 457 -3574 457 -3574 0 3
rlabel polysilicon 464 -3568 464 -3568 0 1
rlabel polysilicon 464 -3574 464 -3574 0 3
rlabel polysilicon 492 -3568 492 -3568 0 1
rlabel polysilicon 492 -3574 492 -3574 0 3
rlabel polysilicon 499 -3568 499 -3568 0 1
rlabel polysilicon 502 -3574 502 -3574 0 4
rlabel polysilicon 562 -3568 562 -3568 0 1
rlabel polysilicon 562 -3574 562 -3574 0 3
rlabel polysilicon 576 -3568 576 -3568 0 1
rlabel polysilicon 579 -3574 579 -3574 0 4
rlabel polysilicon 590 -3568 590 -3568 0 1
rlabel polysilicon 590 -3574 590 -3574 0 3
rlabel polysilicon 597 -3574 597 -3574 0 3
rlabel polysilicon 600 -3574 600 -3574 0 4
rlabel polysilicon 632 -3568 632 -3568 0 1
rlabel polysilicon 632 -3574 632 -3574 0 3
rlabel polysilicon 747 -3568 747 -3568 0 2
rlabel polysilicon 747 -3574 747 -3574 0 4
rlabel polysilicon 758 -3568 758 -3568 0 1
rlabel polysilicon 758 -3574 758 -3574 0 3
rlabel polysilicon 800 -3568 800 -3568 0 1
rlabel polysilicon 800 -3574 800 -3574 0 3
rlabel polysilicon 807 -3568 807 -3568 0 1
rlabel polysilicon 810 -3574 810 -3574 0 4
rlabel polysilicon 884 -3568 884 -3568 0 1
rlabel polysilicon 884 -3574 884 -3574 0 3
rlabel polysilicon 891 -3568 891 -3568 0 1
rlabel polysilicon 894 -3568 894 -3568 0 2
rlabel polysilicon 901 -3568 901 -3568 0 2
rlabel polysilicon 898 -3574 898 -3574 0 3
rlabel polysilicon 1132 -3568 1132 -3568 0 2
rlabel polysilicon 1129 -3574 1129 -3574 0 3
rlabel polysilicon 1136 -3568 1136 -3568 0 1
rlabel polysilicon 1136 -3574 1136 -3574 0 3
rlabel polysilicon 1171 -3568 1171 -3568 0 1
rlabel polysilicon 1171 -3574 1171 -3574 0 3
rlabel polysilicon 1178 -3574 1178 -3574 0 3
rlabel polysilicon 1181 -3574 1181 -3574 0 4
rlabel polysilicon 1185 -3568 1185 -3568 0 1
rlabel polysilicon 1185 -3574 1185 -3574 0 3
rlabel polysilicon 1195 -3574 1195 -3574 0 4
rlabel polysilicon 1199 -3568 1199 -3568 0 1
rlabel polysilicon 1199 -3574 1199 -3574 0 3
rlabel polysilicon 1388 -3568 1388 -3568 0 1
rlabel polysilicon 1391 -3568 1391 -3568 0 2
rlabel polysilicon 1388 -3574 1388 -3574 0 3
rlabel polysilicon 1395 -3568 1395 -3568 0 1
rlabel polysilicon 1395 -3574 1395 -3574 0 3
rlabel metal2 233 1 233 1 0 net=6363
rlabel metal2 443 1 443 1 0 net=12455
rlabel metal2 527 1 527 1 0 net=9869
rlabel metal2 555 1 555 1 0 net=4491
rlabel metal2 877 1 877 1 0 net=12963
rlabel metal2 345 -1 345 -1 0 net=5349
rlabel metal2 359 -1 359 -1 0 net=5635
rlabel metal2 604 -1 604 -1 0 net=11041
rlabel metal2 653 -1 653 -1 0 net=6065
rlabel metal2 716 -1 716 -1 0 net=9775
rlabel metal2 380 -3 380 -3 0 net=3243
rlabel metal2 670 -3 670 -3 0 net=9439
rlabel metal2 401 -5 401 -5 0 net=8281
rlabel metal2 408 -7 408 -7 0 net=2517
rlabel metal2 453 -7 453 -7 0 net=3903
rlabel metal2 415 -9 415 -9 0 net=3831
rlabel metal2 422 -11 422 -11 0 net=3501
rlabel metal2 145 -22 145 -22 0 net=4839
rlabel metal2 156 -22 156 -22 0 net=6365
rlabel metal2 261 -22 261 -22 0 net=5097
rlabel metal2 324 -22 324 -22 0 net=5637
rlabel metal2 373 -22 373 -22 0 net=2519
rlabel metal2 425 -22 425 -22 0 net=12456
rlabel metal2 450 -22 450 -22 0 net=4493
rlabel metal2 590 -22 590 -22 0 net=9117
rlabel metal2 842 -22 842 -22 0 net=11633
rlabel metal2 954 -22 954 -22 0 net=12965
rlabel metal2 226 -24 226 -24 0 net=11269
rlabel metal2 282 -24 282 -24 0 net=4413
rlabel metal2 394 -24 394 -24 0 net=3833
rlabel metal2 429 -24 429 -24 0 net=4973
rlabel metal2 460 -24 460 -24 0 net=11815
rlabel metal2 604 -24 604 -24 0 net=11043
rlabel metal2 604 -24 604 -24 0 net=11043
rlabel metal2 618 -24 618 -24 0 net=8603
rlabel metal2 653 -24 653 -24 0 net=6067
rlabel metal2 677 -24 677 -24 0 net=5825
rlabel metal2 688 -24 688 -24 0 net=9441
rlabel metal2 712 -24 712 -24 0 net=7591
rlabel metal2 800 -24 800 -24 0 net=9777
rlabel metal2 331 -26 331 -26 0 net=3245
rlabel metal2 408 -26 408 -26 0 net=13167
rlabel metal2 653 -26 653 -26 0 net=2315
rlabel metal2 677 -26 677 -26 0 net=12895
rlabel metal2 751 -26 751 -26 0 net=12531
rlabel metal2 338 -28 338 -28 0 net=5351
rlabel metal2 380 -28 380 -28 0 net=8283
rlabel metal2 436 -28 436 -28 0 net=9003
rlabel metal2 688 -28 688 -28 0 net=7263
rlabel metal2 758 -28 758 -28 0 net=10167
rlabel metal2 401 -30 401 -30 0 net=3503
rlabel metal2 432 -30 432 -30 0 net=4789
rlabel metal2 460 -30 460 -30 0 net=13351
rlabel metal2 814 -30 814 -30 0 net=5993
rlabel metal2 464 -32 464 -32 0 net=13631
rlabel metal2 716 -32 716 -32 0 net=12237
rlabel metal2 471 -34 471 -34 0 net=3905
rlabel metal2 492 -34 492 -34 0 net=1571
rlabel metal2 509 -34 509 -34 0 net=9935
rlabel metal2 471 -36 471 -36 0 net=12331
rlabel metal2 520 -36 520 -36 0 net=9509
rlabel metal2 495 -38 495 -38 0 net=1975
rlabel metal2 513 -38 513 -38 0 net=4613
rlabel metal2 523 -40 523 -40 0 net=9087
rlabel metal2 551 -40 551 -40 0 net=6157
rlabel metal2 530 -42 530 -42 0 net=8645
rlabel metal2 534 -44 534 -44 0 net=11777
rlabel metal2 527 -46 527 -46 0 net=9871
rlabel metal2 537 -46 537 -46 0 net=13233
rlabel metal2 464 -48 464 -48 0 net=4869
rlabel metal2 128 -59 128 -59 0 net=6367
rlabel metal2 191 -59 191 -59 0 net=10271
rlabel metal2 205 -59 205 -59 0 net=11271
rlabel metal2 254 -59 254 -59 0 net=8875
rlabel metal2 474 -59 474 -59 0 net=13081
rlabel metal2 744 -59 744 -59 0 net=13353
rlabel metal2 884 -59 884 -59 0 net=13557
rlabel metal2 989 -59 989 -59 0 net=12967
rlabel metal2 149 -61 149 -61 0 net=4841
rlabel metal2 149 -61 149 -61 0 net=4841
rlabel metal2 219 -61 219 -61 0 net=4415
rlabel metal2 289 -61 289 -61 0 net=5638
rlabel metal2 345 -61 345 -61 0 net=4271
rlabel metal2 478 -61 478 -61 0 net=3906
rlabel metal2 492 -61 492 -61 0 net=7471
rlabel metal2 716 -61 716 -61 0 net=12239
rlabel metal2 751 -61 751 -61 0 net=7445
rlabel metal2 898 -61 898 -61 0 net=10169
rlabel metal2 996 -61 996 -61 0 net=12533
rlabel metal2 261 -63 261 -63 0 net=5099
rlabel metal2 275 -63 275 -63 0 net=3105
rlabel metal2 478 -63 478 -63 0 net=8117
rlabel metal2 625 -63 625 -63 0 net=4615
rlabel metal2 730 -63 730 -63 0 net=12897
rlabel metal2 796 -63 796 -63 0 net=13189
rlabel metal2 936 -63 936 -63 0 net=9895
rlabel metal2 247 -65 247 -65 0 net=10483
rlabel metal2 282 -65 282 -65 0 net=2481
rlabel metal2 506 -65 506 -65 0 net=1573
rlabel metal2 551 -65 551 -65 0 net=45
rlabel metal2 688 -65 688 -65 0 net=7265
rlabel metal2 772 -65 772 -65 0 net=7593
rlabel metal2 296 -67 296 -67 0 net=8857
rlabel metal2 422 -67 422 -67 0 net=4791
rlabel metal2 506 -67 506 -67 0 net=6259
rlabel metal2 625 -67 625 -67 0 net=11463
rlabel metal2 817 -67 817 -67 0 net=12929
rlabel metal2 303 -69 303 -69 0 net=5353
rlabel metal2 352 -69 352 -69 0 net=9661
rlabel metal2 555 -69 555 -69 0 net=11817
rlabel metal2 702 -69 702 -69 0 net=9443
rlabel metal2 779 -69 779 -69 0 net=8629
rlabel metal2 306 -71 306 -71 0 net=7819
rlabel metal2 366 -71 366 -71 0 net=3505
rlabel metal2 415 -71 415 -71 0 net=8639
rlabel metal2 555 -71 555 -71 0 net=6159
rlabel metal2 583 -71 583 -71 0 net=13235
rlabel metal2 800 -71 800 -71 0 net=9779
rlabel metal2 310 -73 310 -73 0 net=4495
rlabel metal2 530 -73 530 -73 0 net=7381
rlabel metal2 590 -73 590 -73 0 net=8605
rlabel metal2 646 -73 646 -73 0 net=11779
rlabel metal2 807 -73 807 -73 0 net=11634
rlabel metal2 317 -75 317 -75 0 net=3247
rlabel metal2 338 -75 338 -75 0 net=4871
rlabel metal2 541 -75 541 -75 0 net=9089
rlabel metal2 597 -75 597 -75 0 net=13633
rlabel metal2 712 -75 712 -75 0 net=9567
rlabel metal2 324 -77 324 -77 0 net=2521
rlabel metal2 376 -77 376 -77 0 net=8284
rlabel metal2 387 -77 387 -77 0 net=2435
rlabel metal2 464 -77 464 -77 0 net=12333
rlabel metal2 499 -77 499 -77 0 net=1977
rlabel metal2 604 -77 604 -77 0 net=11045
rlabel metal2 649 -77 649 -77 0 net=410
rlabel metal2 814 -77 814 -77 0 net=5995
rlabel metal2 331 -79 331 -79 0 net=12351
rlabel metal2 534 -79 534 -79 0 net=9873
rlabel metal2 660 -79 660 -79 0 net=9005
rlabel metal2 821 -79 821 -79 0 net=9119
rlabel metal2 334 -81 334 -81 0 net=7891
rlabel metal2 513 -81 513 -81 0 net=8235
rlabel metal2 569 -81 569 -81 0 net=9507
rlabel metal2 611 -81 611 -81 0 net=9937
rlabel metal2 373 -83 373 -83 0 net=5171
rlabel metal2 387 -83 387 -83 0 net=2337
rlabel metal2 548 -83 548 -83 0 net=8647
rlabel metal2 632 -83 632 -83 0 net=2427
rlabel metal2 394 -85 394 -85 0 net=3835
rlabel metal2 394 -85 394 -85 0 net=3835
rlabel metal2 401 -85 401 -85 0 net=4975
rlabel metal2 562 -85 562 -85 0 net=13169
rlabel metal2 411 -87 411 -87 0 net=10015
rlabel metal2 562 -87 562 -87 0 net=2317
rlabel metal2 653 -89 653 -89 0 net=6069
rlabel metal2 667 -91 667 -91 0 net=5827
rlabel metal2 639 -93 639 -93 0 net=9511
rlabel metal2 639 -95 639 -95 0 net=3049
rlabel metal2 89 -106 89 -106 0 net=2011
rlabel metal2 114 -106 114 -106 0 net=6369
rlabel metal2 135 -106 135 -106 0 net=4417
rlabel metal2 226 -106 226 -106 0 net=3413
rlabel metal2 324 -106 324 -106 0 net=2523
rlabel metal2 324 -106 324 -106 0 net=2523
rlabel metal2 345 -106 345 -106 0 net=4272
rlabel metal2 373 -106 373 -106 0 net=3836
rlabel metal2 408 -106 408 -106 0 net=722
rlabel metal2 471 -106 471 -106 0 net=1252
rlabel metal2 513 -106 513 -106 0 net=8236
rlabel metal2 583 -106 583 -106 0 net=7383
rlabel metal2 583 -106 583 -106 0 net=7383
rlabel metal2 611 -106 611 -106 0 net=13170
rlabel metal2 656 -106 656 -106 0 net=12240
rlabel metal2 793 -106 793 -106 0 net=1108
rlabel metal2 828 -106 828 -106 0 net=5997
rlabel metal2 940 -106 940 -106 0 net=13559
rlabel metal2 1010 -106 1010 -106 0 net=12969
rlabel metal2 1087 -106 1087 -106 0 net=12535
rlabel metal2 1195 -106 1195 -106 0 net=11327
rlabel metal2 142 -108 142 -108 0 net=8877
rlabel metal2 261 -108 261 -108 0 net=10485
rlabel metal2 481 -108 481 -108 0 net=479
rlabel metal2 646 -108 646 -108 0 net=7267
rlabel metal2 723 -108 723 -108 0 net=9007
rlabel metal2 856 -108 856 -108 0 net=12931
rlabel metal2 947 -108 947 -108 0 net=9897
rlabel metal2 149 -110 149 -110 0 net=4843
rlabel metal2 149 -110 149 -110 0 net=4843
rlabel metal2 156 -110 156 -110 0 net=7883
rlabel metal2 380 -110 380 -110 0 net=5173
rlabel metal2 394 -110 394 -110 0 net=3051
rlabel metal2 674 -110 674 -110 0 net=11819
rlabel metal2 810 -110 810 -110 0 net=8817
rlabel metal2 954 -110 954 -110 0 net=10171
rlabel metal2 163 -112 163 -112 0 net=11273
rlabel metal2 219 -112 219 -112 0 net=5355
rlabel metal2 310 -112 310 -112 0 net=4497
rlabel metal2 380 -112 380 -112 0 net=12353
rlabel metal2 450 -112 450 -112 0 net=10016
rlabel metal2 485 -112 485 -112 0 net=850
rlabel metal2 513 -112 513 -112 0 net=8885
rlabel metal2 170 -114 170 -114 0 net=5369
rlabel metal2 376 -114 376 -114 0 net=7725
rlabel metal2 530 -114 530 -114 0 net=8085
rlabel metal2 576 -114 576 -114 0 net=9091
rlabel metal2 681 -114 681 -114 0 net=9513
rlabel metal2 744 -114 744 -114 0 net=9781
rlabel metal2 817 -114 817 -114 0 net=4095
rlabel metal2 835 -114 835 -114 0 net=7595
rlabel metal2 177 -116 177 -116 0 net=4873
rlabel metal2 352 -116 352 -116 0 net=9663
rlabel metal2 537 -116 537 -116 0 net=11464
rlabel metal2 660 -116 660 -116 0 net=9939
rlabel metal2 824 -116 824 -116 0 net=12911
rlabel metal2 184 -118 184 -118 0 net=10273
rlabel metal2 198 -118 198 -118 0 net=1883
rlabel metal2 250 -118 250 -118 0 net=2857
rlabel metal2 317 -118 317 -118 0 net=3249
rlabel metal2 338 -118 338 -118 0 net=2429
rlabel metal2 698 -118 698 -118 0 net=10681
rlabel metal2 191 -120 191 -120 0 net=3107
rlabel metal2 289 -120 289 -120 0 net=8159
rlabel metal2 450 -120 450 -120 0 net=5551
rlabel metal2 576 -120 576 -120 0 net=6071
rlabel metal2 709 -120 709 -120 0 net=11781
rlabel metal2 842 -120 842 -120 0 net=9569
rlabel metal2 208 -122 208 -122 0 net=2641
rlabel metal2 460 -122 460 -122 0 net=8601
rlabel metal2 716 -122 716 -122 0 net=12861
rlabel metal2 779 -122 779 -122 0 net=8631
rlabel metal2 856 -122 856 -122 0 net=7741
rlabel metal2 880 -122 880 -122 0 net=8683
rlabel metal2 243 -124 243 -124 0 net=3391
rlabel metal2 408 -124 408 -124 0 net=4793
rlabel metal2 590 -124 590 -124 0 net=8607
rlabel metal2 796 -124 796 -124 0 net=9335
rlabel metal2 863 -124 863 -124 0 net=13191
rlabel metal2 247 -126 247 -126 0 net=1575
rlabel metal2 569 -126 569 -126 0 net=8649
rlabel metal2 597 -126 597 -126 0 net=9875
rlabel metal2 814 -126 814 -126 0 net=12815
rlabel metal2 870 -126 870 -126 0 net=13355
rlabel metal2 254 -128 254 -128 0 net=2483
rlabel metal2 296 -128 296 -128 0 net=8859
rlabel metal2 432 -128 432 -128 0 net=9423
rlabel metal2 611 -128 611 -128 0 net=9435
rlabel metal2 737 -128 737 -128 0 net=13083
rlabel metal2 884 -128 884 -128 0 net=13745
rlabel metal2 261 -130 261 -130 0 net=3875
rlabel metal2 520 -130 520 -130 0 net=9223
rlabel metal2 268 -132 268 -132 0 net=5101
rlabel metal2 432 -132 432 -132 0 net=12334
rlabel metal2 618 -132 618 -132 0 net=11047
rlabel metal2 786 -132 786 -132 0 net=12899
rlabel metal2 891 -132 891 -132 0 net=9121
rlabel metal2 891 -132 891 -132 0 net=9121
rlabel metal2 268 -134 268 -134 0 net=3507
rlabel metal2 415 -134 415 -134 0 net=8640
rlabel metal2 618 -134 618 -134 0 net=7447
rlabel metal2 275 -136 275 -136 0 net=2319
rlabel metal2 625 -136 625 -136 0 net=5829
rlabel metal2 688 -136 688 -136 0 net=13237
rlabel metal2 282 -138 282 -138 0 net=2339
rlabel metal2 401 -138 401 -138 0 net=4977
rlabel metal2 534 -138 534 -138 0 net=7577
rlabel metal2 649 -138 649 -138 0 net=10633
rlabel metal2 296 -140 296 -140 0 net=8119
rlabel metal2 534 -140 534 -140 0 net=6161
rlabel metal2 667 -140 667 -140 0 net=7113
rlabel metal2 366 -142 366 -142 0 net=3229
rlabel metal2 702 -142 702 -142 0 net=13635
rlabel metal2 352 -144 352 -144 0 net=9711
rlabel metal2 730 -144 730 -144 0 net=9445
rlabel metal2 387 -146 387 -146 0 net=2437
rlabel metal2 478 -146 478 -146 0 net=12703
rlabel metal2 695 -146 695 -146 0 net=4617
rlabel metal2 401 -148 401 -148 0 net=6393
rlabel metal2 359 -150 359 -150 0 net=7821
rlabel metal2 359 -152 359 -152 0 net=11933
rlabel metal2 436 -154 436 -154 0 net=1979
rlabel metal2 492 -156 492 -156 0 net=7473
rlabel metal2 492 -158 492 -158 0 net=6261
rlabel metal2 541 -158 541 -158 0 net=9508
rlabel metal2 499 -160 499 -160 0 net=7893
rlabel metal2 499 -162 499 -162 0 net=174
rlabel metal2 506 -164 506 -164 0 net=9469
rlabel metal2 51 -175 51 -175 0 net=11275
rlabel metal2 177 -175 177 -175 0 net=4874
rlabel metal2 516 -175 516 -175 0 net=9729
rlabel metal2 1220 -175 1220 -175 0 net=11329
rlabel metal2 58 -177 58 -177 0 net=3877
rlabel metal2 296 -177 296 -177 0 net=8120
rlabel metal2 530 -177 530 -177 0 net=4096
rlabel metal2 849 -177 849 -177 0 net=9009
rlabel metal2 887 -177 887 -177 0 net=13669
rlabel metal2 1097 -177 1097 -177 0 net=6299
rlabel metal2 65 -179 65 -179 0 net=5553
rlabel metal2 457 -179 457 -179 0 net=9664
rlabel metal2 544 -179 544 -179 0 net=9514
rlabel metal2 737 -179 737 -179 0 net=13637
rlabel metal2 1038 -179 1038 -179 0 net=12971
rlabel metal2 1118 -179 1118 -179 0 net=609
rlabel metal2 72 -181 72 -181 0 net=7885
rlabel metal2 163 -181 163 -181 0 net=5301
rlabel metal2 443 -181 443 -181 0 net=5175
rlabel metal2 541 -181 541 -181 0 net=9163
rlabel metal2 772 -181 772 -181 0 net=11935
rlabel metal2 1129 -181 1129 -181 0 net=12537
rlabel metal2 79 -183 79 -183 0 net=10029
rlabel metal2 474 -183 474 -183 0 net=11727
rlabel metal2 86 -185 86 -185 0 net=6061
rlabel metal2 261 -185 261 -185 0 net=2037
rlabel metal2 366 -185 366 -185 0 net=3230
rlabel metal2 548 -185 548 -185 0 net=8087
rlabel metal2 772 -185 772 -185 0 net=6487
rlabel metal2 863 -185 863 -185 0 net=12817
rlabel metal2 1125 -185 1125 -185 0 net=8435
rlabel metal2 1136 -185 1136 -185 0 net=13747
rlabel metal2 93 -187 93 -187 0 net=2013
rlabel metal2 107 -187 107 -187 0 net=6371
rlabel metal2 121 -187 121 -187 0 net=4729
rlabel metal2 548 -187 548 -187 0 net=7229
rlabel metal2 639 -187 639 -187 0 net=9093
rlabel metal2 639 -187 639 -187 0 net=9093
rlabel metal2 646 -187 646 -187 0 net=7269
rlabel metal2 646 -187 646 -187 0 net=7269
rlabel metal2 653 -187 653 -187 0 net=8632
rlabel metal2 870 -187 870 -187 0 net=12901
rlabel metal2 93 -189 93 -189 0 net=5371
rlabel metal2 177 -189 177 -189 0 net=3109
rlabel metal2 212 -189 212 -189 0 net=5102
rlabel metal2 317 -189 317 -189 0 net=2643
rlabel metal2 380 -189 380 -189 0 net=12354
rlabel metal2 614 -189 614 -189 0 net=11820
rlabel metal2 789 -189 789 -189 0 net=9336
rlabel metal2 877 -189 877 -189 0 net=9123
rlabel metal2 905 -189 905 -189 0 net=10683
rlabel metal2 117 -191 117 -191 0 net=1495
rlabel metal2 184 -191 184 -191 0 net=10274
rlabel metal2 219 -191 219 -191 0 net=5356
rlabel metal2 380 -191 380 -191 0 net=7822
rlabel metal2 569 -191 569 -191 0 net=12705
rlabel metal2 880 -191 880 -191 0 net=12932
rlabel metal2 905 -191 905 -191 0 net=9899
rlabel metal2 975 -191 975 -191 0 net=13357
rlabel metal2 128 -193 128 -193 0 net=3509
rlabel metal2 292 -193 292 -193 0 net=3317
rlabel metal2 383 -193 383 -193 0 net=5167
rlabel metal2 656 -193 656 -193 0 net=11097
rlabel metal2 996 -193 996 -193 0 net=13561
rlabel metal2 142 -195 142 -195 0 net=8878
rlabel metal2 219 -195 219 -195 0 net=2341
rlabel metal2 296 -195 296 -195 0 net=7385
rlabel metal2 688 -195 688 -195 0 net=9471
rlabel metal2 898 -195 898 -195 0 net=8819
rlabel metal2 954 -195 954 -195 0 net=13193
rlabel metal2 142 -197 142 -197 0 net=4845
rlabel metal2 156 -197 156 -197 0 net=8599
rlabel metal2 688 -197 688 -197 0 net=7743
rlabel metal2 933 -197 933 -197 0 net=8887
rlabel metal2 149 -199 149 -199 0 net=4795
rlabel metal2 415 -199 415 -199 0 net=4978
rlabel metal2 457 -199 457 -199 0 net=8602
rlabel metal2 681 -199 681 -199 0 net=9877
rlabel metal2 940 -199 940 -199 0 net=9571
rlabel metal2 968 -199 968 -199 0 net=10173
rlabel metal2 996 -199 996 -199 0 net=11111
rlabel metal2 184 -201 184 -201 0 net=1885
rlabel metal2 254 -201 254 -201 0 net=2485
rlabel metal2 303 -201 303 -201 0 net=1751
rlabel metal2 632 -201 632 -201 0 net=8609
rlabel metal2 681 -201 681 -201 0 net=7597
rlabel metal2 999 -201 999 -201 0 net=12161
rlabel metal2 191 -203 191 -203 0 net=2169
rlabel metal2 254 -203 254 -203 0 net=2525
rlabel metal2 345 -203 345 -203 0 net=3393
rlabel metal2 429 -203 429 -203 0 net=6163
rlabel metal2 562 -203 562 -203 0 net=7579
rlabel metal2 698 -203 698 -203 0 net=13491
rlabel metal2 1010 -203 1010 -203 0 net=12913
rlabel metal2 268 -205 268 -205 0 net=2439
rlabel metal2 394 -205 394 -205 0 net=3053
rlabel metal2 492 -205 492 -205 0 net=6263
rlabel metal2 709 -205 709 -205 0 net=11049
rlabel metal2 947 -205 947 -205 0 net=9225
rlabel metal2 275 -207 275 -207 0 net=2321
rlabel metal2 509 -207 509 -207 0 net=5807
rlabel metal2 716 -207 716 -207 0 net=12863
rlabel metal2 208 -209 208 -209 0 net=1947
rlabel metal2 289 -209 289 -209 0 net=8161
rlabel metal2 345 -209 345 -209 0 net=2625
rlabel metal2 387 -209 387 -209 0 net=4759
rlabel metal2 534 -209 534 -209 0 net=4619
rlabel metal2 744 -209 744 -209 0 net=9783
rlabel metal2 243 -211 243 -211 0 net=1116
rlabel metal2 310 -211 310 -211 0 net=2859
rlabel metal2 422 -211 422 -211 0 net=8861
rlabel metal2 751 -211 751 -211 0 net=13239
rlabel metal2 135 -213 135 -213 0 net=4418
rlabel metal2 310 -213 310 -213 0 net=3251
rlabel metal2 359 -213 359 -213 0 net=4121
rlabel metal2 135 -215 135 -215 0 net=13103
rlabel metal2 317 -215 317 -215 0 net=2431
rlabel metal2 422 -215 422 -215 0 net=3099
rlabel metal2 604 -215 604 -215 0 net=7895
rlabel metal2 765 -215 765 -215 0 net=8415
rlabel metal2 233 -217 233 -217 0 net=10199
rlabel metal2 765 -217 765 -217 0 net=8685
rlabel metal2 247 -219 247 -219 0 net=1577
rlabel metal2 471 -219 471 -219 0 net=10487
rlabel metal2 247 -221 247 -221 0 net=1561
rlabel metal2 562 -221 562 -221 0 net=8651
rlabel metal2 604 -221 604 -221 0 net=5831
rlabel metal2 660 -221 660 -221 0 net=9437
rlabel metal2 768 -221 768 -221 0 net=9955
rlabel metal2 331 -223 331 -223 0 net=4395
rlabel metal2 702 -223 702 -223 0 net=9713
rlabel metal2 779 -223 779 -223 0 net=10635
rlabel metal2 436 -225 436 -225 0 net=1980
rlabel metal2 478 -225 478 -225 0 net=4951
rlabel metal2 611 -225 611 -225 0 net=6975
rlabel metal2 793 -225 793 -225 0 net=10879
rlabel metal2 236 -227 236 -227 0 net=4171
rlabel metal2 520 -227 520 -227 0 net=6073
rlabel metal2 611 -227 611 -227 0 net=10089
rlabel metal2 226 -229 226 -229 0 net=3414
rlabel metal2 541 -229 541 -229 0 net=7169
rlabel metal2 793 -229 793 -229 0 net=5999
rlabel metal2 226 -231 226 -231 0 net=4499
rlabel metal2 555 -231 555 -231 0 net=7475
rlabel metal2 719 -231 719 -231 0 net=12425
rlabel metal2 373 -233 373 -233 0 net=4103
rlabel metal2 555 -233 555 -233 0 net=5605
rlabel metal2 796 -233 796 -233 0 net=13725
rlabel metal2 572 -235 572 -235 0 net=8715
rlabel metal2 800 -235 800 -235 0 net=9941
rlabel metal2 502 -237 502 -237 0 net=9611
rlabel metal2 807 -237 807 -237 0 net=11783
rlabel metal2 618 -239 618 -239 0 net=7449
rlabel metal2 786 -239 786 -239 0 net=9447
rlabel metal2 814 -239 814 -239 0 net=13085
rlabel metal2 460 -241 460 -241 0 net=4775
rlabel metal2 597 -243 597 -243 0 net=9425
rlabel metal2 597 -245 597 -245 0 net=7115
rlabel metal2 485 -247 485 -247 0 net=7727
rlabel metal2 401 -249 401 -249 0 net=6395
rlabel metal2 401 -251 401 -251 0 net=4295
rlabel metal2 44 -262 44 -262 0 net=7387
rlabel metal2 383 -262 383 -262 0 net=5049
rlabel metal2 548 -262 548 -262 0 net=7231
rlabel metal2 593 -262 593 -262 0 net=10090
rlabel metal2 989 -262 989 -262 0 net=11785
rlabel metal2 51 -264 51 -264 0 net=11276
rlabel metal2 285 -264 285 -264 0 net=6300
rlabel metal2 1164 -264 1164 -264 0 net=13727
rlabel metal2 51 -266 51 -266 0 net=6165
rlabel metal2 460 -266 460 -266 0 net=7728
rlabel metal2 681 -266 681 -266 0 net=7599
rlabel metal2 996 -266 996 -266 0 net=9731
rlabel metal2 1202 -266 1202 -266 0 net=13429
rlabel metal2 58 -268 58 -268 0 net=3878
rlabel metal2 415 -268 415 -268 0 net=2323
rlabel metal2 471 -268 471 -268 0 net=9438
rlabel metal2 772 -268 772 -268 0 net=6489
rlabel metal2 828 -268 828 -268 0 net=12345
rlabel metal2 1227 -268 1227 -268 0 net=11331
rlabel metal2 1227 -268 1227 -268 0 net=11331
rlabel metal2 1255 -268 1255 -268 0 net=13749
rlabel metal2 61 -270 61 -270 0 net=7886
rlabel metal2 86 -270 86 -270 0 net=6062
rlabel metal2 474 -270 474 -270 0 net=9472
rlabel metal2 842 -270 842 -270 0 net=12707
rlabel metal2 72 -272 72 -272 0 net=5373
rlabel metal2 96 -272 96 -272 0 net=4730
rlabel metal2 142 -272 142 -272 0 net=4847
rlabel metal2 474 -272 474 -272 0 net=13099
rlabel metal2 65 -274 65 -274 0 net=5555
rlabel metal2 156 -274 156 -274 0 net=8600
rlabel metal2 338 -274 338 -274 0 net=1579
rlabel metal2 506 -274 506 -274 0 net=11021
rlabel metal2 1283 -274 1283 -274 0 net=11729
rlabel metal2 65 -276 65 -276 0 net=2249
rlabel metal2 509 -276 509 -276 0 net=9878
rlabel metal2 863 -276 863 -276 0 net=11051
rlabel metal2 86 -278 86 -278 0 net=6295
rlabel metal2 163 -278 163 -278 0 net=5302
rlabel metal2 513 -278 513 -278 0 net=5169
rlabel metal2 107 -280 107 -280 0 net=6373
rlabel metal2 387 -280 387 -280 0 net=4761
rlabel metal2 527 -280 527 -280 0 net=11129
rlabel metal2 107 -282 107 -282 0 net=1927
rlabel metal2 527 -282 527 -282 0 net=6265
rlabel metal2 614 -282 614 -282 0 net=13240
rlabel metal2 1024 -282 1024 -282 0 net=11937
rlabel metal2 93 -284 93 -284 0 net=4551
rlabel metal2 499 -284 499 -284 0 net=5177
rlabel metal2 632 -284 632 -284 0 net=8611
rlabel metal2 863 -284 863 -284 0 net=8641
rlabel metal2 1101 -284 1101 -284 0 net=13563
rlabel metal2 121 -286 121 -286 0 net=5079
rlabel metal2 163 -286 163 -286 0 net=2171
rlabel metal2 215 -286 215 -286 0 net=12555
rlabel metal2 170 -288 170 -288 0 net=2487
rlabel metal2 352 -288 352 -288 0 net=2645
rlabel metal2 450 -288 450 -288 0 net=3054
rlabel metal2 509 -288 509 -288 0 net=5941
rlabel metal2 667 -288 667 -288 0 net=12781
rlabel metal2 184 -290 184 -290 0 net=1887
rlabel metal2 184 -290 184 -290 0 net=1887
rlabel metal2 198 -290 198 -290 0 net=8127
rlabel metal2 576 -290 576 -290 0 net=8055
rlabel metal2 891 -290 891 -290 0 net=8417
rlabel metal2 905 -290 905 -290 0 net=9901
rlabel metal2 1038 -290 1038 -290 0 net=12819
rlabel metal2 135 -292 135 -292 0 net=13105
rlabel metal2 579 -292 579 -292 0 net=9094
rlabel metal2 681 -292 681 -292 0 net=6243
rlabel metal2 723 -292 723 -292 0 net=8089
rlabel metal2 891 -292 891 -292 0 net=8821
rlabel metal2 912 -292 912 -292 0 net=12427
rlabel metal2 201 -294 201 -294 0 net=1581
rlabel metal2 408 -294 408 -294 0 net=3394
rlabel metal2 478 -294 478 -294 0 net=4953
rlabel metal2 688 -294 688 -294 0 net=7745
rlabel metal2 933 -294 933 -294 0 net=10637
rlabel metal2 1101 -294 1101 -294 0 net=8889
rlabel metal2 1171 -294 1171 -294 0 net=12539
rlabel metal2 114 -296 114 -296 0 net=9061
rlabel metal2 1045 -296 1045 -296 0 net=12865
rlabel metal2 205 -298 205 -298 0 net=440
rlabel metal2 544 -298 544 -298 0 net=7245
rlabel metal2 744 -298 744 -298 0 net=9715
rlabel metal2 1052 -298 1052 -298 0 net=12903
rlabel metal2 282 -300 282 -300 0 net=2626
rlabel metal2 359 -300 359 -300 0 net=4123
rlabel metal2 499 -300 499 -300 0 net=4403
rlabel metal2 275 -302 275 -302 0 net=1949
rlabel metal2 359 -302 359 -302 0 net=4105
rlabel metal2 443 -302 443 -302 0 net=11841
rlabel metal2 198 -304 198 -304 0 net=3725
rlabel metal2 611 -304 611 -304 0 net=10123
rlabel metal2 1059 -304 1059 -304 0 net=11113
rlabel metal2 317 -306 317 -306 0 net=2433
rlabel metal2 373 -306 373 -306 0 net=3101
rlabel metal2 611 -306 611 -306 0 net=13638
rlabel metal2 1073 -306 1073 -306 0 net=13195
rlabel metal2 58 -308 58 -308 0 net=9973
rlabel metal2 1073 -308 1073 -308 0 net=10349
rlabel metal2 1108 -308 1108 -308 0 net=12973
rlabel metal2 324 -310 324 -310 0 net=8162
rlabel metal2 422 -310 422 -310 0 net=5607
rlabel metal2 614 -310 614 -310 0 net=6915
rlabel metal2 747 -310 747 -310 0 net=13492
rlabel metal2 1017 -310 1017 -310 0 net=10685
rlabel metal2 1115 -310 1115 -310 0 net=8436
rlabel metal2 1136 -310 1136 -310 0 net=12915
rlabel metal2 173 -312 173 -312 0 net=10747
rlabel metal2 1118 -312 1118 -312 0 net=12329
rlabel metal2 324 -314 324 -314 0 net=2969
rlabel metal2 751 -314 751 -314 0 net=11409
rlabel metal2 492 -316 492 -316 0 net=9999
rlabel metal2 226 -318 226 -318 0 net=4501
rlabel metal2 555 -318 555 -318 0 net=6001
rlabel metal2 800 -318 800 -318 0 net=9613
rlabel metal2 968 -318 968 -318 0 net=10175
rlabel metal2 1066 -318 1066 -318 0 net=12163
rlabel metal2 149 -320 149 -320 0 net=4797
rlabel metal2 495 -320 495 -320 0 net=7729
rlabel metal2 807 -320 807 -320 0 net=9449
rlabel metal2 807 -320 807 -320 0 net=9449
rlabel metal2 814 -320 814 -320 0 net=9427
rlabel metal2 1080 -320 1080 -320 0 net=13359
rlabel metal2 149 -322 149 -322 0 net=2557
rlabel metal2 618 -322 618 -322 0 net=4777
rlabel metal2 695 -322 695 -322 0 net=8717
rlabel metal2 919 -322 919 -322 0 net=9957
rlabel metal2 975 -322 975 -322 0 net=11099
rlabel metal2 1087 -322 1087 -322 0 net=13671
rlabel metal2 607 -324 607 -324 0 net=6267
rlabel metal2 625 -324 625 -324 0 net=7171
rlabel metal2 705 -324 705 -324 0 net=11355
rlabel metal2 520 -326 520 -326 0 net=6075
rlabel metal2 670 -326 670 -326 0 net=10163
rlabel metal2 1122 -326 1122 -326 0 net=11671
rlabel metal2 520 -328 520 -328 0 net=4621
rlabel metal2 674 -328 674 -328 0 net=7581
rlabel metal2 870 -328 870 -328 0 net=9785
rlabel metal2 366 -330 366 -330 0 net=3319
rlabel metal2 562 -330 562 -330 0 net=8653
rlabel metal2 926 -330 926 -330 0 net=10489
rlabel metal2 191 -332 191 -332 0 net=5459
rlabel metal2 653 -332 653 -332 0 net=5809
rlabel metal2 709 -332 709 -332 0 net=7897
rlabel metal2 884 -332 884 -332 0 net=9011
rlabel metal2 961 -332 961 -332 0 net=10881
rlabel metal2 79 -334 79 -334 0 net=10030
rlabel metal2 712 -334 712 -334 0 net=12669
rlabel metal2 79 -336 79 -336 0 net=4397
rlabel metal2 439 -336 439 -336 0 net=8779
rlabel metal2 730 -336 730 -336 0 net=8863
rlabel metal2 975 -336 975 -336 0 net=9227
rlabel metal2 177 -338 177 -338 0 net=3111
rlabel metal2 254 -338 254 -338 0 net=2527
rlabel metal2 730 -338 730 -338 0 net=10503
rlabel metal2 177 -340 177 -340 0 net=1563
rlabel metal2 331 -340 331 -340 0 net=2727
rlabel metal2 754 -340 754 -340 0 net=11605
rlabel metal2 999 -340 999 -340 0 net=10387
rlabel metal2 208 -342 208 -342 0 net=1651
rlabel metal2 758 -342 758 -342 0 net=10201
rlabel metal2 646 -344 646 -344 0 net=7271
rlabel metal2 779 -344 779 -344 0 net=6977
rlabel metal2 877 -344 877 -344 0 net=9125
rlabel metal2 194 -346 194 -346 0 net=6009
rlabel metal2 660 -346 660 -346 0 net=7477
rlabel metal2 786 -346 786 -346 0 net=13177
rlabel metal2 117 -348 117 -348 0 net=7583
rlabel metal2 789 -348 789 -348 0 net=13086
rlabel metal2 117 -350 117 -350 0 net=2115
rlabel metal2 569 -350 569 -350 0 net=8783
rlabel metal2 940 -350 940 -350 0 net=9573
rlabel metal2 569 -352 569 -352 0 net=11169
rlabel metal2 604 -354 604 -354 0 net=5833
rlabel metal2 737 -354 737 -354 0 net=9165
rlabel metal2 485 -356 485 -356 0 net=6397
rlabel metal2 849 -356 849 -356 0 net=9943
rlabel metal2 401 -358 401 -358 0 net=4297
rlabel metal2 597 -358 597 -358 0 net=7116
rlabel metal2 765 -358 765 -358 0 net=8687
rlabel metal2 289 -360 289 -360 0 net=6057
rlabel metal2 702 -360 702 -360 0 net=7451
rlabel metal2 275 -362 275 -362 0 net=5503
rlabel metal2 289 -364 289 -364 0 net=1753
rlabel metal2 338 -364 338 -364 0 net=3653
rlabel metal2 303 -366 303 -366 0 net=2861
rlabel metal2 268 -368 268 -368 0 net=2441
rlabel metal2 268 -370 268 -370 0 net=3253
rlabel metal2 261 -372 261 -372 0 net=2039
rlabel metal2 219 -374 219 -374 0 net=2343
rlabel metal2 219 -376 219 -376 0 net=4173
rlabel metal2 128 -378 128 -378 0 net=3510
rlabel metal2 100 -380 100 -380 0 net=2015
rlabel metal2 100 -382 100 -382 0 net=3683
rlabel metal2 23 -393 23 -393 0 net=2007
rlabel metal2 247 -393 247 -393 0 net=1511
rlabel metal2 506 -393 506 -393 0 net=12708
rlabel metal2 1297 -393 1297 -393 0 net=12867
rlabel metal2 1591 -393 1591 -393 0 net=11731
rlabel metal2 30 -395 30 -395 0 net=3727
rlabel metal2 450 -395 450 -395 0 net=13465
rlabel metal2 37 -397 37 -397 0 net=3685
rlabel metal2 107 -397 107 -397 0 net=1928
rlabel metal2 408 -397 408 -397 0 net=5178
rlabel metal2 597 -397 597 -397 0 net=6058
rlabel metal2 772 -397 772 -397 0 net=6491
rlabel metal2 772 -397 772 -397 0 net=6491
rlabel metal2 1143 -397 1143 -397 0 net=13179
rlabel metal2 58 -399 58 -399 0 net=5505
rlabel metal2 317 -399 317 -399 0 net=2647
rlabel metal2 429 -399 429 -399 0 net=1580
rlabel metal2 530 -399 530 -399 0 net=608
rlabel metal2 1031 -399 1031 -399 0 net=9975
rlabel metal2 1164 -399 1164 -399 0 net=13361
rlabel metal2 72 -401 72 -401 0 net=5375
rlabel metal2 72 -401 72 -401 0 net=5375
rlabel metal2 82 -401 82 -401 0 net=13106
rlabel metal2 607 -401 607 -401 0 net=11052
rlabel metal2 1346 -401 1346 -401 0 net=13729
rlabel metal2 86 -403 86 -403 0 net=6297
rlabel metal2 429 -403 429 -403 0 net=7273
rlabel metal2 933 -403 933 -403 0 net=9063
rlabel metal2 1052 -403 1052 -403 0 net=10165
rlabel metal2 1171 -403 1171 -403 0 net=11843
rlabel metal2 1353 -403 1353 -403 0 net=13431
rlabel metal2 86 -405 86 -405 0 net=7917
rlabel metal2 611 -405 611 -405 0 net=7582
rlabel metal2 807 -405 807 -405 0 net=9451
rlabel metal2 1066 -405 1066 -405 0 net=10203
rlabel metal2 1178 -405 1178 -405 0 net=11357
rlabel metal2 1304 -405 1304 -405 0 net=12905
rlabel metal2 89 -407 89 -407 0 net=2016
rlabel metal2 135 -407 135 -407 0 net=8487
rlabel metal2 982 -407 982 -407 0 net=9717
rlabel metal2 1073 -407 1073 -407 0 net=10351
rlabel metal2 1220 -407 1220 -407 0 net=13673
rlabel metal2 93 -409 93 -409 0 net=7531
rlabel metal2 110 -409 110 -409 0 net=8864
rlabel metal2 982 -409 982 -409 0 net=10389
rlabel metal2 1094 -409 1094 -409 0 net=10639
rlabel metal2 1227 -409 1227 -409 0 net=11333
rlabel metal2 1311 -409 1311 -409 0 net=12917
rlabel metal2 96 -411 96 -411 0 net=6244
rlabel metal2 695 -411 695 -411 0 net=7173
rlabel metal2 905 -411 905 -411 0 net=9615
rlabel metal2 1115 -411 1115 -411 0 net=10749
rlabel metal2 1269 -411 1269 -411 0 net=12671
rlabel metal2 100 -413 100 -413 0 net=12330
rlabel metal2 1269 -413 1269 -413 0 net=11295
rlabel metal2 114 -415 114 -415 0 net=2345
rlabel metal2 268 -415 268 -415 0 net=3254
rlabel metal2 324 -415 324 -415 0 net=2970
rlabel metal2 481 -415 481 -415 0 net=10467
rlabel metal2 1136 -415 1136 -415 0 net=12165
rlabel metal2 1353 -415 1353 -415 0 net=12113
rlabel metal2 65 -417 65 -417 0 net=2251
rlabel metal2 324 -417 324 -417 0 net=4461
rlabel metal2 576 -417 576 -417 0 net=4779
rlabel metal2 695 -417 695 -417 0 net=6398
rlabel metal2 747 -417 747 -417 0 net=11365
rlabel metal2 1318 -417 1318 -417 0 net=12975
rlabel metal2 65 -419 65 -419 0 net=4107
rlabel metal2 366 -419 366 -419 0 net=2529
rlabel metal2 436 -419 436 -419 0 net=6266
rlabel metal2 534 -419 534 -419 0 net=3320
rlabel metal2 618 -419 618 -419 0 net=6269
rlabel metal2 733 -419 733 -419 0 net=11385
rlabel metal2 1325 -419 1325 -419 0 net=13101
rlabel metal2 79 -421 79 -421 0 net=4399
rlabel metal2 401 -421 401 -421 0 net=3655
rlabel metal2 439 -421 439 -421 0 net=6325
rlabel metal2 758 -421 758 -421 0 net=8090
rlabel metal2 884 -421 884 -421 0 net=11607
rlabel metal2 1332 -421 1332 -421 0 net=13197
rlabel metal2 79 -423 79 -423 0 net=233
rlabel metal2 474 -423 474 -423 0 net=10119
rlabel metal2 1192 -423 1192 -423 0 net=11673
rlabel metal2 1374 -423 1374 -423 0 net=13751
rlabel metal2 121 -425 121 -425 0 net=764
rlabel metal2 331 -425 331 -425 0 net=2729
rlabel metal2 485 -425 485 -425 0 net=4299
rlabel metal2 534 -425 534 -425 0 net=11515
rlabel metal2 121 -427 121 -427 0 net=4405
rlabel metal2 541 -427 541 -427 0 net=5051
rlabel metal2 639 -427 639 -427 0 net=4954
rlabel metal2 842 -427 842 -427 0 net=10883
rlabel metal2 1206 -427 1206 -427 0 net=11939
rlabel metal2 124 -429 124 -429 0 net=10000
rlabel metal2 1276 -429 1276 -429 0 net=12783
rlabel metal2 128 -431 128 -431 0 net=2801
rlabel metal2 156 -431 156 -431 0 net=5081
rlabel metal2 156 -431 156 -431 0 net=5081
rlabel metal2 163 -431 163 -431 0 net=2173
rlabel metal2 170 -431 170 -431 0 net=2488
rlabel metal2 464 -431 464 -431 0 net=2325
rlabel metal2 492 -431 492 -431 0 net=4503
rlabel metal2 653 -431 653 -431 0 net=8781
rlabel metal2 856 -431 856 -431 0 net=6979
rlabel metal2 919 -431 919 -431 0 net=9013
rlabel metal2 954 -431 954 -431 0 net=9575
rlabel metal2 1283 -431 1283 -431 0 net=12821
rlabel metal2 51 -433 51 -433 0 net=6167
rlabel metal2 660 -433 660 -433 0 net=5835
rlabel metal2 670 -433 670 -433 0 net=5170
rlabel metal2 51 -435 51 -435 0 net=2863
rlabel metal2 331 -435 331 -435 0 net=2819
rlabel metal2 478 -435 478 -435 0 net=4125
rlabel metal2 509 -435 509 -435 0 net=7765
rlabel metal2 898 -435 898 -435 0 net=8419
rlabel metal2 968 -435 968 -435 0 net=9959
rlabel metal2 1255 -435 1255 -435 0 net=12541
rlabel metal2 163 -437 163 -437 0 net=1755
rlabel metal2 303 -437 303 -437 0 net=2443
rlabel metal2 443 -437 443 -437 0 net=3279
rlabel metal2 604 -437 604 -437 0 net=8203
rlabel metal2 989 -437 989 -437 0 net=9903
rlabel metal2 1150 -437 1150 -437 0 net=11115
rlabel metal2 1283 -437 1283 -437 0 net=13565
rlabel metal2 352 -439 352 -439 0 net=2434
rlabel metal2 562 -439 562 -439 0 net=5461
rlabel metal2 625 -439 625 -439 0 net=6077
rlabel metal2 674 -439 674 -439 0 net=5811
rlabel metal2 702 -439 702 -439 0 net=11786
rlabel metal2 26 -441 26 -441 0 net=4625
rlabel metal2 632 -441 632 -441 0 net=5943
rlabel metal2 712 -441 712 -441 0 net=11277
rlabel metal2 142 -443 142 -443 0 net=5557
rlabel metal2 632 -443 632 -443 0 net=6381
rlabel metal2 142 -445 142 -445 0 net=6375
rlabel metal2 352 -445 352 -445 0 net=6003
rlabel metal2 716 -445 716 -445 0 net=7247
rlabel metal2 863 -445 863 -445 0 net=8643
rlabel metal2 1010 -445 1010 -445 0 net=9945
rlabel metal2 1213 -445 1213 -445 0 net=12347
rlabel metal2 117 -447 117 -447 0 net=6189
rlabel metal2 800 -447 800 -447 0 net=7731
rlabel metal2 877 -447 877 -447 0 net=8785
rlabel metal2 1017 -447 1017 -447 0 net=10505
rlabel metal2 1241 -447 1241 -447 0 net=12429
rlabel metal2 170 -449 170 -449 0 net=5609
rlabel metal2 464 -449 464 -449 0 net=7233
rlabel metal2 649 -449 649 -449 0 net=7955
rlabel metal2 891 -449 891 -449 0 net=8823
rlabel metal2 1017 -449 1017 -449 0 net=8891
rlabel metal2 1108 -449 1108 -449 0 net=10687
rlabel metal2 180 -451 180 -451 0 net=6127
rlabel metal2 709 -451 709 -451 0 net=10925
rlabel metal2 187 -453 187 -453 0 net=2893
rlabel metal2 478 -453 478 -453 0 net=11130
rlabel metal2 194 -455 194 -455 0 net=5365
rlabel metal2 779 -455 779 -455 0 net=7479
rlabel metal2 898 -455 898 -455 0 net=9515
rlabel metal2 198 -457 198 -457 0 net=8033
rlabel metal2 996 -457 996 -457 0 net=9733
rlabel metal2 1199 -457 1199 -457 0 net=11755
rlabel metal2 184 -459 184 -459 0 net=1889
rlabel metal2 205 -459 205 -459 0 net=3631
rlabel metal2 282 -459 282 -459 0 net=6311
rlabel metal2 870 -459 870 -459 0 net=8655
rlabel metal2 1003 -459 1003 -459 0 net=9787
rlabel metal2 1185 -459 1185 -459 0 net=11411
rlabel metal2 205 -461 205 -461 0 net=4763
rlabel metal2 520 -461 520 -461 0 net=4623
rlabel metal2 590 -461 590 -461 0 net=7746
rlabel metal2 870 -461 870 -461 0 net=7601
rlabel metal2 1003 -461 1003 -461 0 net=6345
rlabel metal2 44 -463 44 -463 0 net=7389
rlabel metal2 849 -463 849 -463 0 net=8689
rlabel metal2 1038 -463 1038 -463 0 net=10125
rlabel metal2 1262 -463 1262 -463 0 net=12557
rlabel metal2 44 -465 44 -465 0 net=4799
rlabel metal2 254 -465 254 -465 0 net=1653
rlabel metal2 282 -465 282 -465 0 net=5749
rlabel metal2 520 -465 520 -465 0 net=9428
rlabel metal2 1045 -465 1045 -465 0 net=11101
rlabel metal2 1087 -465 1087 -465 0 net=10491
rlabel metal2 191 -467 191 -467 0 net=3113
rlabel metal2 254 -467 254 -467 0 net=1917
rlabel metal2 635 -467 635 -467 0 net=9577
rlabel metal2 191 -469 191 -469 0 net=1273
rlabel metal2 723 -469 723 -469 0 net=6917
rlabel metal2 786 -469 786 -469 0 net=7585
rlabel metal2 940 -469 940 -469 0 net=9167
rlabel metal2 1087 -469 1087 -469 0 net=11171
rlabel metal2 138 -471 138 -471 0 net=7841
rlabel metal2 961 -471 961 -471 0 net=9127
rlabel metal2 1059 -471 1059 -471 0 net=10177
rlabel metal2 138 -473 138 -473 0 net=8657
rlabel metal2 723 -473 723 -473 0 net=7899
rlabel metal2 828 -473 828 -473 0 net=8057
rlabel metal2 215 -475 215 -475 0 net=3651
rlabel metal2 828 -475 828 -475 0 net=11022
rlabel metal2 107 -477 107 -477 0 net=10807
rlabel metal2 219 -479 219 -479 0 net=4175
rlabel metal2 835 -479 835 -479 0 net=8613
rlabel metal2 975 -479 975 -479 0 net=9229
rlabel metal2 338 -481 338 -481 0 net=7361
rlabel metal2 912 -481 912 -481 0 net=8719
rlabel metal2 338 -483 338 -483 0 net=1951
rlabel metal2 380 -483 380 -483 0 net=1583
rlabel metal2 548 -483 548 -483 0 net=8129
rlabel metal2 149 -485 149 -485 0 net=2559
rlabel metal2 457 -485 457 -485 0 net=4553
rlabel metal2 597 -485 597 -485 0 net=8521
rlabel metal2 149 -487 149 -487 0 net=1565
rlabel metal2 310 -487 310 -487 0 net=2041
rlabel metal2 457 -487 457 -487 0 net=6011
rlabel metal2 765 -487 765 -487 0 net=7453
rlabel metal2 177 -489 177 -489 0 net=1440
rlabel metal2 310 -489 310 -489 0 net=4849
rlabel metal2 646 -489 646 -489 0 net=3701
rlabel metal2 212 -491 212 -491 0 net=2117
rlabel metal2 373 -491 373 -491 0 net=3103
rlabel metal2 219 -493 219 -493 0 net=2279
rlabel metal2 320 -493 320 -493 0 net=1869
rlabel metal2 9 -504 9 -504 0 net=5751
rlabel metal2 317 -504 317 -504 0 net=2649
rlabel metal2 450 -504 450 -504 0 net=7732
rlabel metal2 873 -504 873 -504 0 net=10390
rlabel metal2 1045 -504 1045 -504 0 net=9169
rlabel metal2 1045 -504 1045 -504 0 net=9169
rlabel metal2 1136 -504 1136 -504 0 net=10121
rlabel metal2 1269 -504 1269 -504 0 net=11297
rlabel metal2 1468 -504 1468 -504 0 net=6561
rlabel metal2 1710 -504 1710 -504 0 net=11733
rlabel metal2 23 -506 23 -506 0 net=2865
rlabel metal2 58 -506 58 -506 0 net=5506
rlabel metal2 103 -506 103 -506 0 net=4462
rlabel metal2 345 -506 345 -506 0 net=2043
rlabel metal2 345 -506 345 -506 0 net=2043
rlabel metal2 359 -506 359 -506 0 net=6298
rlabel metal2 450 -506 450 -506 0 net=5052
rlabel metal2 583 -506 583 -506 0 net=7919
rlabel metal2 618 -506 618 -506 0 net=8659
rlabel metal2 1129 -506 1129 -506 0 net=9961
rlabel metal2 1171 -506 1171 -506 0 net=10205
rlabel metal2 1171 -506 1171 -506 0 net=10205
rlabel metal2 1269 -506 1269 -506 0 net=11387
rlabel metal2 1486 -506 1486 -506 0 net=13467
rlabel metal2 1528 -506 1528 -506 0 net=9517
rlabel metal2 37 -508 37 -508 0 net=3686
rlabel metal2 194 -508 194 -508 0 net=10166
rlabel metal2 1493 -508 1493 -508 0 net=13675
rlabel metal2 1493 -508 1493 -508 0 net=13675
rlabel metal2 1500 -508 1500 -508 0 net=13731
rlabel metal2 1514 -508 1514 -508 0 net=6383
rlabel metal2 61 -510 61 -510 0 net=9578
rlabel metal2 1458 -510 1458 -510 0 net=13199
rlabel metal2 79 -512 79 -512 0 net=2243
rlabel metal2 362 -512 362 -512 0 net=8782
rlabel metal2 758 -512 758 -512 0 net=11756
rlabel metal2 1451 -512 1451 -512 0 net=13181
rlabel metal2 1500 -512 1500 -512 0 net=13753
rlabel metal2 72 -514 72 -514 0 net=5377
rlabel metal2 103 -514 103 -514 0 net=7609
rlabel metal2 453 -514 453 -514 0 net=1157
rlabel metal2 604 -514 604 -514 0 net=5463
rlabel metal2 604 -514 604 -514 0 net=5463
rlabel metal2 618 -514 618 -514 0 net=10469
rlabel metal2 1122 -514 1122 -514 0 net=9947
rlabel metal2 1150 -514 1150 -514 0 net=10127
rlabel metal2 1325 -514 1325 -514 0 net=11609
rlabel metal2 1430 -514 1430 -514 0 net=12977
rlabel metal2 72 -516 72 -516 0 net=2347
rlabel metal2 128 -516 128 -516 0 net=2803
rlabel metal2 222 -516 222 -516 0 net=3652
rlabel metal2 709 -516 709 -516 0 net=10640
rlabel metal2 1402 -516 1402 -516 0 net=12785
rlabel metal2 107 -518 107 -518 0 net=4407
rlabel metal2 128 -518 128 -518 0 net=1585
rlabel metal2 401 -518 401 -518 0 net=2730
rlabel metal2 481 -518 481 -518 0 net=3702
rlabel metal2 824 -518 824 -518 0 net=9576
rlabel metal2 114 -520 114 -520 0 net=6055
rlabel metal2 541 -520 541 -520 0 net=4505
rlabel metal2 541 -520 541 -520 0 net=4505
rlabel metal2 548 -520 548 -520 0 net=4555
rlabel metal2 583 -520 583 -520 0 net=8614
rlabel metal2 1052 -520 1052 -520 0 net=9453
rlabel metal2 1185 -520 1185 -520 0 net=10493
rlabel metal2 121 -522 121 -522 0 net=1953
rlabel metal2 341 -522 341 -522 0 net=4517
rlabel metal2 590 -522 590 -522 0 net=80
rlabel metal2 831 -522 831 -522 0 net=10049
rlabel metal2 1199 -522 1199 -522 0 net=11413
rlabel metal2 138 -524 138 -524 0 net=12868
rlabel metal2 152 -526 152 -526 0 net=1364
rlabel metal2 593 -526 593 -526 0 net=9277
rlabel metal2 1080 -526 1080 -526 0 net=11103
rlabel metal2 1416 -526 1416 -526 0 net=12919
rlabel metal2 156 -528 156 -528 0 net=5082
rlabel metal2 243 -528 243 -528 0 net=7551
rlabel metal2 373 -528 373 -528 0 net=1870
rlabel metal2 593 -528 593 -528 0 net=10439
rlabel metal2 1213 -528 1213 -528 0 net=10689
rlabel metal2 1395 -528 1395 -528 0 net=12559
rlabel metal2 44 -530 44 -530 0 net=4801
rlabel metal2 597 -530 597 -530 0 net=7363
rlabel metal2 828 -530 828 -530 0 net=7455
rlabel metal2 842 -530 842 -530 0 net=10885
rlabel metal2 1367 -530 1367 -530 0 net=12349
rlabel metal2 44 -532 44 -532 0 net=6059
rlabel metal2 905 -532 905 -532 0 net=8035
rlabel metal2 905 -532 905 -532 0 net=8035
rlabel metal2 947 -532 947 -532 0 net=8691
rlabel metal2 961 -532 961 -532 0 net=9719
rlabel metal2 1178 -532 1178 -532 0 net=10353
rlabel metal2 1332 -532 1332 -532 0 net=11675
rlabel metal2 93 -534 93 -534 0 net=7533
rlabel metal2 177 -534 177 -534 0 net=1891
rlabel metal2 268 -534 268 -534 0 net=2253
rlabel metal2 317 -534 317 -534 0 net=3104
rlabel metal2 779 -534 779 -534 0 net=6919
rlabel metal2 842 -534 842 -534 0 net=12822
rlabel metal2 93 -536 93 -536 0 net=6377
rlabel metal2 180 -536 180 -536 0 net=4764
rlabel metal2 268 -536 268 -536 0 net=4341
rlabel metal2 530 -536 530 -536 0 net=6270
rlabel metal2 761 -536 761 -536 0 net=10187
rlabel metal2 1318 -536 1318 -536 0 net=11517
rlabel metal2 1409 -536 1409 -536 0 net=12907
rlabel metal2 65 -538 65 -538 0 net=4109
rlabel metal2 530 -538 530 -538 0 net=5963
rlabel metal2 667 -538 667 -538 0 net=5836
rlabel metal2 716 -538 716 -538 0 net=6191
rlabel metal2 765 -538 765 -538 0 net=11845
rlabel metal2 1388 -538 1388 -538 0 net=12543
rlabel metal2 65 -540 65 -540 0 net=6291
rlabel metal2 142 -540 142 -540 0 net=6013
rlabel metal2 460 -540 460 -540 0 net=12672
rlabel metal2 135 -542 135 -542 0 net=1567
rlabel metal2 191 -542 191 -542 0 net=2209
rlabel metal2 464 -542 464 -542 0 net=7234
rlabel metal2 653 -542 653 -542 0 net=6169
rlabel metal2 677 -542 677 -542 0 net=6657
rlabel metal2 723 -542 723 -542 0 net=7901
rlabel metal2 915 -542 915 -542 0 net=12219
rlabel metal2 149 -544 149 -544 0 net=4850
rlabel metal2 352 -544 352 -544 0 net=6005
rlabel metal2 681 -544 681 -544 0 net=5813
rlabel metal2 730 -544 730 -544 0 net=7175
rlabel metal2 947 -544 947 -544 0 net=8787
rlabel metal2 1017 -544 1017 -544 0 net=8893
rlabel metal2 1157 -544 1157 -544 0 net=10179
rlabel metal2 1297 -544 1297 -544 0 net=11359
rlabel metal2 1339 -544 1339 -544 0 net=12431
rlabel metal2 198 -546 198 -546 0 net=1919
rlabel metal2 275 -546 275 -546 0 net=1655
rlabel metal2 310 -546 310 -546 0 net=4301
rlabel metal2 516 -546 516 -546 0 net=6277
rlabel metal2 779 -546 779 -546 0 net=13102
rlabel metal2 30 -548 30 -548 0 net=3729
rlabel metal2 516 -548 516 -548 0 net=10069
rlabel metal2 1297 -548 1297 -548 0 net=12167
rlabel metal2 1472 -548 1472 -548 0 net=13433
rlabel metal2 163 -550 163 -550 0 net=1757
rlabel metal2 366 -550 366 -550 0 net=4401
rlabel metal2 380 -550 380 -550 0 net=2561
rlabel metal2 464 -550 464 -550 0 net=2357
rlabel metal2 786 -550 786 -550 0 net=7843
rlabel metal2 954 -550 954 -550 0 net=8421
rlabel metal2 1038 -550 1038 -550 0 net=9129
rlabel metal2 1283 -550 1283 -550 0 net=13567
rlabel metal2 163 -552 163 -552 0 net=3633
rlabel metal2 366 -552 366 -552 0 net=2327
rlabel metal2 492 -552 492 -552 0 net=7480
rlabel metal2 919 -552 919 -552 0 net=9015
rlabel metal2 1052 -552 1052 -552 0 net=11366
rlabel metal2 1346 -552 1346 -552 0 net=13363
rlabel metal2 205 -554 205 -554 0 net=1513
rlabel metal2 254 -554 254 -554 0 net=4781
rlabel metal2 625 -554 625 -554 0 net=5558
rlabel metal2 891 -554 891 -554 0 net=11367
rlabel metal2 30 -556 30 -556 0 net=6703
rlabel metal2 261 -556 261 -556 0 net=1509
rlabel metal2 485 -556 485 -556 0 net=5367
rlabel metal2 625 -556 625 -556 0 net=6313
rlabel metal2 786 -556 786 -556 0 net=6347
rlabel metal2 1241 -556 1241 -556 0 net=10927
rlabel metal2 1290 -556 1290 -556 0 net=11335
rlabel metal2 170 -558 170 -558 0 net=5611
rlabel metal2 632 -558 632 -558 0 net=8656
rlabel metal2 1087 -558 1087 -558 0 net=11173
rlabel metal2 170 -560 170 -560 0 net=7275
rlabel metal2 436 -560 436 -560 0 net=3657
rlabel metal2 492 -560 492 -560 0 net=7767
rlabel metal2 919 -560 919 -560 0 net=8059
rlabel metal2 1087 -560 1087 -560 0 net=10751
rlabel metal2 226 -562 226 -562 0 net=3115
rlabel metal2 387 -562 387 -562 0 net=2531
rlabel metal2 418 -562 418 -562 0 net=10655
rlabel metal2 226 -564 226 -564 0 net=3281
rlabel metal2 471 -564 471 -564 0 net=4627
rlabel metal2 576 -564 576 -564 0 net=9734
rlabel metal2 1195 -564 1195 -564 0 net=10589
rlabel metal2 233 -566 233 -566 0 net=2009
rlabel metal2 495 -566 495 -566 0 net=8644
rlabel metal2 1055 -566 1055 -566 0 net=9019
rlabel metal2 303 -568 303 -568 0 net=2445
rlabel metal2 499 -568 499 -568 0 net=4127
rlabel metal2 499 -568 499 -568 0 net=4127
rlabel metal2 523 -568 523 -568 0 net=12143
rlabel metal2 240 -570 240 -570 0 net=2281
rlabel metal2 331 -570 331 -570 0 net=2821
rlabel metal2 527 -570 527 -570 0 net=12655
rlabel metal2 212 -572 212 -572 0 net=2119
rlabel metal2 527 -572 527 -572 0 net=11278
rlabel metal2 212 -574 212 -574 0 net=2895
rlabel metal2 562 -574 562 -574 0 net=6493
rlabel metal2 793 -574 793 -574 0 net=6981
rlabel metal2 1255 -574 1255 -574 0 net=11117
rlabel metal2 240 -576 240 -576 0 net=2174
rlabel metal2 338 -576 338 -576 0 net=3443
rlabel metal2 635 -576 635 -576 0 net=9616
rlabel metal2 1234 -576 1234 -576 0 net=10809
rlabel metal2 1503 -576 1503 -576 0 net=1
rlabel metal2 289 -578 289 -578 0 net=1823
rlabel metal2 579 -578 579 -578 0 net=256
rlabel metal2 639 -578 639 -578 0 net=4177
rlabel metal2 772 -578 772 -578 0 net=7587
rlabel metal2 856 -578 856 -578 0 net=8489
rlabel metal2 968 -578 968 -578 0 net=8721
rlabel metal2 1094 -578 1094 -578 0 net=9905
rlabel metal2 1206 -578 1206 -578 0 net=10507
rlabel metal2 639 -580 639 -580 0 net=5945
rlabel metal2 688 -580 688 -580 0 net=7249
rlabel metal2 849 -580 849 -580 0 net=8941
rlabel metal2 1101 -580 1101 -580 0 net=9789
rlabel metal2 1143 -580 1143 -580 0 net=9977
rlabel metal2 555 -582 555 -582 0 net=4624
rlabel metal2 698 -582 698 -582 0 net=8791
rlabel metal2 1031 -582 1031 -582 0 net=9065
rlabel metal2 51 -584 51 -584 0 net=8405
rlabel metal2 702 -584 702 -584 0 net=6129
rlabel metal2 866 -584 866 -584 0 net=10211
rlabel metal2 513 -586 513 -586 0 net=4657
rlabel metal2 660 -586 660 -586 0 net=6079
rlabel metal2 702 -586 702 -586 0 net=5857
rlabel metal2 877 -586 877 -586 0 net=7957
rlabel metal2 1024 -586 1024 -586 0 net=9231
rlabel metal2 86 -588 86 -588 0 net=7539
rlabel metal2 737 -588 737 -588 0 net=6327
rlabel metal2 870 -588 870 -588 0 net=7603
rlabel metal2 884 -588 884 -588 0 net=7635
rlabel metal2 926 -588 926 -588 0 net=8205
rlabel metal2 1010 -588 1010 -588 0 net=8825
rlabel metal2 86 -590 86 -590 0 net=3559
rlabel metal2 744 -590 744 -590 0 net=7391
rlabel metal2 912 -590 912 -590 0 net=8131
rlabel metal2 940 -590 940 -590 0 net=8523
rlabel metal2 453 -592 453 -592 0 net=8333
rlabel metal2 821 -594 821 -594 0 net=13611
rlabel metal2 912 -596 912 -596 0 net=11940
rlabel metal2 1353 -598 1353 -598 0 net=12115
rlabel metal2 110 -600 110 -600 0 net=11563
rlabel metal2 9 -611 9 -611 0 net=5752
rlabel metal2 492 -611 492 -611 0 net=7768
rlabel metal2 604 -611 604 -611 0 net=5465
rlabel metal2 653 -611 653 -611 0 net=6007
rlabel metal2 674 -611 674 -611 0 net=6279
rlabel metal2 761 -611 761 -611 0 net=8788
rlabel metal2 1017 -611 1017 -611 0 net=8423
rlabel metal2 1332 -611 1332 -611 0 net=11519
rlabel metal2 1332 -611 1332 -611 0 net=11519
rlabel metal2 1339 -611 1339 -611 0 net=12433
rlabel metal2 1535 -611 1535 -611 0 net=11369
rlabel metal2 9 -613 9 -613 0 net=4343
rlabel metal2 282 -613 282 -613 0 net=1657
rlabel metal2 282 -613 282 -613 0 net=1657
rlabel metal2 303 -613 303 -613 0 net=2283
rlabel metal2 320 -613 320 -613 0 net=5499
rlabel metal2 408 -613 408 -613 0 net=7610
rlabel metal2 786 -613 786 -613 0 net=6348
rlabel metal2 824 -613 824 -613 0 net=9720
rlabel metal2 1241 -613 1241 -613 0 net=10657
rlabel metal2 1346 -613 1346 -613 0 net=13365
rlabel metal2 1668 -613 1668 -613 0 net=6463
rlabel metal2 16 -615 16 -615 0 net=6379
rlabel metal2 114 -615 114 -615 0 net=6056
rlabel metal2 205 -615 205 -615 0 net=1515
rlabel metal2 205 -615 205 -615 0 net=1515
rlabel metal2 233 -615 233 -615 0 net=1510
rlabel metal2 303 -615 303 -615 0 net=2245
rlabel metal2 362 -615 362 -615 0 net=714
rlabel metal2 653 -615 653 -615 0 net=6171
rlabel metal2 677 -615 677 -615 0 net=12786
rlabel metal2 1437 -615 1437 -615 0 net=12909
rlabel metal2 1738 -615 1738 -615 0 net=6385
rlabel metal2 30 -617 30 -617 0 net=1461
rlabel metal2 72 -617 72 -617 0 net=2348
rlabel metal2 534 -617 534 -617 0 net=4803
rlabel metal2 534 -617 534 -617 0 net=4803
rlabel metal2 544 -617 544 -617 0 net=5612
rlabel metal2 660 -617 660 -617 0 net=7541
rlabel metal2 1087 -617 1087 -617 0 net=10753
rlabel metal2 1388 -617 1388 -617 0 net=12221
rlabel metal2 1556 -617 1556 -617 0 net=6562
rlabel metal2 1759 -617 1759 -617 0 net=11735
rlabel metal2 30 -619 30 -619 0 net=2367
rlabel metal2 145 -619 145 -619 0 net=3455
rlabel metal2 352 -619 352 -619 0 net=3117
rlabel metal2 569 -619 569 -619 0 net=4557
rlabel metal2 604 -619 604 -619 0 net=6659
rlabel metal2 786 -619 786 -619 0 net=6285
rlabel metal2 1157 -619 1157 -619 0 net=10071
rlabel metal2 1325 -619 1325 -619 0 net=11415
rlabel metal2 1444 -619 1444 -619 0 net=12921
rlabel metal2 1766 -619 1766 -619 0 net=9519
rlabel metal2 37 -621 37 -621 0 net=7379
rlabel metal2 873 -621 873 -621 0 net=11279
rlabel metal2 1409 -621 1409 -621 0 net=12545
rlabel metal2 44 -623 44 -623 0 net=6060
rlabel metal2 114 -623 114 -623 0 net=10886
rlabel metal2 1290 -623 1290 -623 0 net=11175
rlabel metal2 1416 -623 1416 -623 0 net=12561
rlabel metal2 44 -625 44 -625 0 net=4129
rlabel metal2 667 -625 667 -625 0 net=5859
rlabel metal2 709 -625 709 -625 0 net=12855
rlabel metal2 51 -627 51 -627 0 net=8407
rlabel metal2 79 -627 79 -627 0 net=5379
rlabel metal2 128 -627 128 -627 0 net=1587
rlabel metal2 373 -627 373 -627 0 net=4402
rlabel metal2 436 -627 436 -627 0 net=2823
rlabel metal2 436 -627 436 -627 0 net=2823
rlabel metal2 499 -627 499 -627 0 net=3731
rlabel metal2 681 -627 681 -627 0 net=6081
rlabel metal2 793 -627 793 -627 0 net=6983
rlabel metal2 933 -627 933 -627 0 net=10122
rlabel metal2 1206 -627 1206 -627 0 net=9979
rlabel metal2 1269 -627 1269 -627 0 net=11389
rlabel metal2 1423 -627 1423 -627 0 net=12657
rlabel metal2 51 -629 51 -629 0 net=6085
rlabel metal2 128 -629 128 -629 0 net=1569
rlabel metal2 149 -629 149 -629 0 net=5315
rlabel metal2 373 -629 373 -629 0 net=3813
rlabel metal2 408 -629 408 -629 0 net=3445
rlabel metal2 429 -629 429 -629 0 net=4629
rlabel metal2 509 -629 509 -629 0 net=8881
rlabel metal2 1227 -629 1227 -629 0 net=10591
rlabel metal2 1451 -629 1451 -629 0 net=12979
rlabel metal2 58 -631 58 -631 0 net=6293
rlabel metal2 79 -631 79 -631 0 net=4409
rlabel metal2 135 -631 135 -631 0 net=13645
rlabel metal2 65 -633 65 -633 0 net=6015
rlabel metal2 149 -633 149 -633 0 net=2897
rlabel metal2 243 -633 243 -633 0 net=2010
rlabel metal2 681 -633 681 -633 0 net=4179
rlabel metal2 796 -633 796 -633 0 net=678
rlabel metal2 1472 -633 1472 -633 0 net=13435
rlabel metal2 142 -635 142 -635 0 net=11846
rlabel metal2 800 -635 800 -635 0 net=6921
rlabel metal2 842 -635 842 -635 0 net=9066
rlabel metal2 1108 -635 1108 -635 0 net=9021
rlabel metal2 1178 -635 1178 -635 0 net=10181
rlabel metal2 1353 -635 1353 -635 0 net=11565
rlabel metal2 1479 -635 1479 -635 0 net=13569
rlabel metal2 100 -637 100 -637 0 net=9113
rlabel metal2 1129 -637 1129 -637 0 net=9949
rlabel metal2 1360 -637 1360 -637 0 net=11611
rlabel metal2 1468 -637 1468 -637 0 net=11941
rlabel metal2 1486 -637 1486 -637 0 net=13613
rlabel metal2 100 -639 100 -639 0 net=2211
rlabel metal2 212 -639 212 -639 0 net=7491
rlabel metal2 562 -639 562 -639 0 net=6495
rlabel metal2 849 -639 849 -639 0 net=13200
rlabel metal2 156 -641 156 -641 0 net=7535
rlabel metal2 894 -641 894 -641 0 net=11104
rlabel metal2 1458 -641 1458 -641 0 net=13183
rlabel metal2 156 -643 156 -643 0 net=2563
rlabel metal2 415 -643 415 -643 0 net=2650
rlabel metal2 562 -643 562 -643 0 net=7177
rlabel metal2 737 -643 737 -643 0 net=6329
rlabel metal2 782 -643 782 -643 0 net=11589
rlabel metal2 1493 -643 1493 -643 0 net=13677
rlabel metal2 163 -645 163 -645 0 net=3635
rlabel metal2 513 -645 513 -645 0 net=4519
rlabel metal2 569 -645 569 -645 0 net=6929
rlabel metal2 845 -645 845 -645 0 net=11775
rlabel metal2 163 -647 163 -647 0 net=5965
rlabel metal2 660 -647 660 -647 0 net=7357
rlabel metal2 852 -647 852 -647 0 net=10354
rlabel metal2 1255 -647 1255 -647 0 net=10811
rlabel metal2 1374 -647 1374 -647 0 net=12117
rlabel metal2 1500 -647 1500 -647 0 net=13755
rlabel metal2 170 -649 170 -649 0 net=7276
rlabel metal2 593 -649 593 -649 0 net=6673
rlabel metal2 863 -649 863 -649 0 net=10319
rlabel metal2 1507 -649 1507 -649 0 net=13733
rlabel metal2 170 -651 170 -651 0 net=10257
rlabel metal2 1297 -651 1297 -651 0 net=12169
rlabel metal2 173 -653 173 -653 0 net=10470
rlabel metal2 646 -653 646 -653 0 net=1333
rlabel metal2 723 -653 723 -653 0 net=5815
rlabel metal2 870 -653 870 -653 0 net=5591
rlabel metal2 989 -653 989 -653 0 net=8693
rlabel metal2 1115 -653 1115 -653 0 net=9791
rlabel metal2 1248 -653 1248 -653 0 net=10691
rlabel metal2 1311 -653 1311 -653 0 net=11337
rlabel metal2 1381 -653 1381 -653 0 net=12145
rlabel metal2 177 -655 177 -655 0 net=1893
rlabel metal2 177 -655 177 -655 0 net=1893
rlabel metal2 187 -655 187 -655 0 net=11583
rlabel metal2 191 -657 191 -657 0 net=1921
rlabel metal2 236 -657 236 -657 0 net=1699
rlabel metal2 422 -657 422 -657 0 net=4821
rlabel metal2 635 -657 635 -657 0 net=7981
rlabel metal2 996 -657 996 -657 0 net=8943
rlabel metal2 1136 -657 1136 -657 0 net=9963
rlabel metal2 1367 -657 1367 -657 0 net=11677
rlabel metal2 198 -659 198 -659 0 net=1709
rlabel metal2 366 -659 366 -659 0 net=2329
rlabel metal2 520 -659 520 -659 0 net=4111
rlabel metal2 656 -659 656 -659 0 net=1
rlabel metal2 730 -659 730 -659 0 net=7393
rlabel metal2 877 -659 877 -659 0 net=7605
rlabel metal2 1024 -659 1024 -659 0 net=8827
rlabel metal2 1164 -659 1164 -659 0 net=10129
rlabel metal2 1276 -659 1276 -659 0 net=11119
rlabel metal2 61 -661 61 -661 0 net=8953
rlabel metal2 1031 -661 1031 -661 0 net=9233
rlabel metal2 1185 -661 1185 -661 0 net=10189
rlabel metal2 1283 -661 1283 -661 0 net=10929
rlabel metal2 236 -663 236 -663 0 net=5237
rlabel metal2 625 -663 625 -663 0 net=6315
rlabel metal2 828 -663 828 -663 0 net=7457
rlabel metal2 898 -663 898 -663 0 net=7921
rlabel metal2 1038 -663 1038 -663 0 net=9017
rlabel metal2 1318 -663 1318 -663 0 net=11361
rlabel metal2 240 -665 240 -665 0 net=2031
rlabel metal2 387 -665 387 -665 0 net=2446
rlabel metal2 625 -665 625 -665 0 net=5727
rlabel metal2 1059 -665 1059 -665 0 net=9737
rlabel metal2 1199 -665 1199 -665 0 net=10441
rlabel metal2 240 -667 240 -667 0 net=7425
rlabel metal2 856 -667 856 -667 0 net=8491
rlabel metal2 1066 -667 1066 -667 0 net=9131
rlabel metal2 1171 -667 1171 -667 0 net=10207
rlabel metal2 152 -669 152 -669 0 net=7237
rlabel metal2 908 -669 908 -669 0 net=13313
rlabel metal2 254 -671 254 -671 0 net=4782
rlabel metal2 926 -671 926 -671 0 net=8133
rlabel metal2 1045 -671 1045 -671 0 net=9171
rlabel metal2 1234 -671 1234 -671 0 net=10509
rlabel metal2 261 -673 261 -673 0 net=2045
rlabel metal2 387 -673 387 -673 0 net=2349
rlabel metal2 688 -673 688 -673 0 net=7251
rlabel metal2 884 -673 884 -673 0 net=7637
rlabel metal2 954 -673 954 -673 0 net=8207
rlabel metal2 1073 -673 1073 -673 0 net=9279
rlabel metal2 331 -675 331 -675 0 net=2121
rlabel metal2 345 -675 345 -675 0 net=2195
rlabel metal2 520 -675 520 -675 0 net=4507
rlabel metal2 586 -675 586 -675 0 net=827
rlabel metal2 940 -675 940 -675 0 net=8335
rlabel metal2 1080 -675 1080 -675 0 net=8895
rlabel metal2 1143 -675 1143 -675 0 net=10213
rlabel metal2 275 -677 275 -677 0 net=1759
rlabel metal2 401 -677 401 -677 0 net=5947
rlabel metal2 691 -677 691 -677 0 net=570
rlabel metal2 975 -677 975 -677 0 net=7959
rlabel metal2 1150 -677 1150 -677 0 net=10051
rlabel metal2 275 -679 275 -679 0 net=2533
rlabel metal2 432 -679 432 -679 0 net=10705
rlabel metal2 394 -681 394 -681 0 net=2919
rlabel metal2 793 -681 793 -681 0 net=7629
rlabel metal2 982 -681 982 -681 0 net=8661
rlabel metal2 247 -683 247 -683 0 net=6704
rlabel metal2 814 -683 814 -683 0 net=7903
rlabel metal2 1003 -683 1003 -683 0 net=8793
rlabel metal2 247 -685 247 -685 0 net=1825
rlabel metal2 443 -685 443 -685 0 net=3403
rlabel metal2 597 -685 597 -685 0 net=7365
rlabel metal2 695 -685 695 -685 0 net=9454
rlabel metal2 289 -687 289 -687 0 net=2255
rlabel metal2 464 -687 464 -687 0 net=2359
rlabel metal2 541 -687 541 -687 0 net=5187
rlabel metal2 695 -687 695 -687 0 net=6121
rlabel metal2 1010 -687 1010 -687 0 net=8525
rlabel metal2 1122 -687 1122 -687 0 net=12350
rlabel metal2 23 -689 23 -689 0 net=2866
rlabel metal2 555 -689 555 -689 0 net=4659
rlabel metal2 597 -689 597 -689 0 net=12617
rlabel metal2 1304 -689 1304 -689 0 net=11299
rlabel metal2 23 -691 23 -691 0 net=4303
rlabel metal2 698 -691 698 -691 0 net=12205
rlabel metal2 121 -693 121 -693 0 net=1955
rlabel metal2 740 -693 740 -693 0 net=8287
rlabel metal2 1220 -693 1220 -693 0 net=10495
rlabel metal2 121 -695 121 -695 0 net=3287
rlabel metal2 772 -695 772 -695 0 net=7589
rlabel metal2 1094 -695 1094 -695 0 net=9907
rlabel metal2 219 -697 219 -697 0 net=2805
rlabel metal2 450 -697 450 -697 0 net=3659
rlabel metal2 758 -697 758 -697 0 net=6193
rlabel metal2 807 -697 807 -697 0 net=6131
rlabel metal2 828 -697 828 -697 0 net=13468
rlabel metal2 86 -699 86 -699 0 net=3561
rlabel metal2 254 -699 254 -699 0 net=4585
rlabel metal2 506 -699 506 -699 0 net=12223
rlabel metal2 86 -701 86 -701 0 net=3283
rlabel metal2 621 -701 621 -701 0 net=7159
rlabel metal2 835 -701 835 -701 0 net=7845
rlabel metal2 968 -701 968 -701 0 net=8723
rlabel metal2 226 -703 226 -703 0 net=5759
rlabel metal2 884 -703 884 -703 0 net=12207
rlabel metal2 905 -703 905 -703 0 net=8037
rlabel metal2 359 -705 359 -705 0 net=7553
rlabel metal2 919 -705 919 -705 0 net=8061
rlabel metal2 359 -707 359 -707 0 net=5368
rlabel metal2 485 -709 485 -709 0 net=2449
rlabel metal2 9 -720 9 -720 0 net=4344
rlabel metal2 114 -720 114 -720 0 net=779
rlabel metal2 1787 -720 1787 -720 0 net=11371
rlabel metal2 9 -722 9 -722 0 net=4823
rlabel metal2 439 -722 439 -722 0 net=696
rlabel metal2 562 -722 562 -722 0 net=7178
rlabel metal2 709 -722 709 -722 0 net=9018
rlabel metal2 1458 -722 1458 -722 0 net=11591
rlabel metal2 1857 -722 1857 -722 0 net=9521
rlabel metal2 16 -724 16 -724 0 net=6380
rlabel metal2 121 -724 121 -724 0 net=3288
rlabel metal2 128 -724 128 -724 0 net=1570
rlabel metal2 170 -724 170 -724 0 net=865
rlabel metal2 254 -724 254 -724 0 net=4587
rlabel metal2 303 -724 303 -724 0 net=2247
rlabel metal2 422 -724 422 -724 0 net=7065
rlabel metal2 723 -724 723 -724 0 net=6008
rlabel metal2 740 -724 740 -724 0 net=12910
rlabel metal2 1605 -724 1605 -724 0 net=13315
rlabel metal2 1801 -724 1801 -724 0 net=6465
rlabel metal2 37 -726 37 -726 0 net=7380
rlabel metal2 254 -726 254 -726 0 net=2361
rlabel metal2 548 -726 548 -726 0 net=4113
rlabel metal2 586 -726 586 -726 0 net=7343
rlabel metal2 999 -726 999 -726 0 net=12562
rlabel metal2 1577 -726 1577 -726 0 net=12923
rlabel metal2 1822 -726 1822 -726 0 net=6387
rlabel metal2 37 -728 37 -728 0 net=6473
rlabel metal2 597 -728 597 -728 0 net=10442
rlabel metal2 1486 -728 1486 -728 0 net=12119
rlabel metal2 1794 -728 1794 -728 0 net=11737
rlabel metal2 58 -730 58 -730 0 net=6294
rlabel metal2 555 -730 555 -730 0 net=12033
rlabel metal2 1612 -730 1612 -730 0 net=13571
rlabel metal2 30 -732 30 -732 0 net=2369
rlabel metal2 79 -732 79 -732 0 net=4411
rlabel metal2 121 -732 121 -732 0 net=4077
rlabel metal2 268 -732 268 -732 0 net=3457
rlabel metal2 618 -732 618 -732 0 net=9403
rlabel metal2 1360 -732 1360 -732 0 net=10813
rlabel metal2 1493 -732 1493 -732 0 net=12147
rlabel metal2 1626 -732 1626 -732 0 net=13615
rlabel metal2 30 -734 30 -734 0 net=2213
rlabel metal2 135 -734 135 -734 0 net=278
rlabel metal2 170 -734 170 -734 0 net=1895
rlabel metal2 201 -734 201 -734 0 net=10587
rlabel metal2 1570 -734 1570 -734 0 net=12857
rlabel metal2 1584 -734 1584 -734 0 net=12981
rlabel metal2 93 -736 93 -736 0 net=1873
rlabel metal2 268 -736 268 -736 0 net=1701
rlabel metal2 443 -736 443 -736 0 net=3405
rlabel metal2 520 -736 520 -736 0 net=4509
rlabel metal2 614 -736 614 -736 0 net=346
rlabel metal2 621 -736 621 -736 0 net=11105
rlabel metal2 1542 -736 1542 -736 0 net=12547
rlabel metal2 65 -738 65 -738 0 net=6017
rlabel metal2 628 -738 628 -738 0 net=7394
rlabel metal2 779 -738 779 -738 0 net=11566
rlabel metal2 1479 -738 1479 -738 0 net=11943
rlabel metal2 1633 -738 1633 -738 0 net=13647
rlabel metal2 65 -740 65 -740 0 net=3963
rlabel metal2 632 -740 632 -740 0 net=5467
rlabel metal2 758 -740 758 -740 0 net=10947
rlabel metal2 1549 -740 1549 -740 0 net=13437
rlabel metal2 100 -742 100 -742 0 net=2257
rlabel metal2 303 -742 303 -742 0 net=2351
rlabel metal2 443 -742 443 -742 0 net=2451
rlabel metal2 495 -742 495 -742 0 net=219
rlabel metal2 831 -742 831 -742 0 net=12081
rlabel metal2 1671 -742 1671 -742 0 net=13123
rlabel metal2 107 -744 107 -744 0 net=5381
rlabel metal2 275 -744 275 -744 0 net=2535
rlabel metal2 450 -744 450 -744 0 net=3661
rlabel metal2 590 -744 590 -744 0 net=4559
rlabel metal2 674 -744 674 -744 0 net=6281
rlabel metal2 712 -744 712 -744 0 net=6763
rlabel metal2 107 -746 107 -746 0 net=2331
rlabel metal2 478 -746 478 -746 0 net=7590
rlabel metal2 1034 -746 1034 -746 0 net=8705
rlabel metal2 135 -748 135 -748 0 net=3733
rlabel metal2 653 -748 653 -748 0 net=6173
rlabel metal2 681 -748 681 -748 0 net=4181
rlabel metal2 779 -748 779 -748 0 net=13059
rlabel metal2 173 -750 173 -750 0 net=3118
rlabel metal2 464 -750 464 -750 0 net=8336
rlabel metal2 1143 -750 1143 -750 0 net=12619
rlabel metal2 96 -752 96 -752 0 net=5279
rlabel metal2 478 -752 478 -752 0 net=5861
rlabel metal2 716 -752 716 -752 0 net=9172
rlabel metal2 1234 -752 1234 -752 0 net=10053
rlabel metal2 1367 -752 1367 -752 0 net=10931
rlabel metal2 1465 -752 1465 -752 0 net=11613
rlabel metal2 1549 -752 1549 -752 0 net=13185
rlabel metal2 1633 -752 1633 -752 0 net=13757
rlabel metal2 156 -754 156 -754 0 net=2565
rlabel metal2 467 -754 467 -754 0 net=4865
rlabel metal2 723 -754 723 -754 0 net=7631
rlabel metal2 1045 -754 1045 -754 0 net=8209
rlabel metal2 1178 -754 1178 -754 0 net=9235
rlabel metal2 1234 -754 1234 -754 0 net=10497
rlabel metal2 1339 -754 1339 -754 0 net=10659
rlabel metal2 1556 -754 1556 -754 0 net=12659
rlabel metal2 51 -756 51 -756 0 net=6087
rlabel metal2 275 -756 275 -756 0 net=1659
rlabel metal2 289 -756 289 -756 0 net=1717
rlabel metal2 639 -756 639 -756 0 net=7367
rlabel metal2 782 -756 782 -756 0 net=6667
rlabel metal2 919 -756 919 -756 0 net=7542
rlabel metal2 1073 -756 1073 -756 0 net=9909
rlabel metal2 1241 -756 1241 -756 0 net=10073
rlabel metal2 1381 -756 1381 -756 0 net=11121
rlabel metal2 1556 -756 1556 -756 0 net=11823
rlabel metal2 282 -758 282 -758 0 net=2285
rlabel metal2 324 -758 324 -758 0 net=5317
rlabel metal2 793 -758 793 -758 0 net=11176
rlabel metal2 1444 -758 1444 -758 0 net=11585
rlabel metal2 1640 -758 1640 -758 0 net=13679
rlabel metal2 296 -760 296 -760 0 net=2806
rlabel metal2 835 -760 835 -760 0 net=7555
rlabel metal2 1080 -760 1080 -760 0 net=8663
rlabel metal2 1195 -760 1195 -760 0 net=12403
rlabel metal2 324 -762 324 -762 0 net=3435
rlabel metal2 922 -762 922 -762 0 net=13449
rlabel metal2 345 -764 345 -764 0 net=2196
rlabel metal2 772 -764 772 -764 0 net=6195
rlabel metal2 800 -764 800 -764 0 net=6497
rlabel metal2 807 -764 807 -764 0 net=7161
rlabel metal2 1052 -764 1052 -764 0 net=8425
rlabel metal2 1094 -764 1094 -764 0 net=8725
rlabel metal2 1262 -764 1262 -764 0 net=9981
rlabel metal2 1388 -764 1388 -764 0 net=11281
rlabel metal2 1647 -764 1647 -764 0 net=13735
rlabel metal2 345 -766 345 -766 0 net=2033
rlabel metal2 373 -766 373 -766 0 net=3815
rlabel metal2 1136 -766 1136 -766 0 net=8829
rlabel metal2 1269 -766 1269 -766 0 net=10183
rlabel metal2 1402 -766 1402 -766 0 net=11363
rlabel metal2 310 -768 310 -768 0 net=1957
rlabel metal2 373 -768 373 -768 0 net=5949
rlabel metal2 436 -768 436 -768 0 net=2825
rlabel metal2 492 -768 492 -768 0 net=3637
rlabel metal2 569 -768 569 -768 0 net=6931
rlabel metal2 695 -768 695 -768 0 net=6123
rlabel metal2 800 -768 800 -768 0 net=5593
rlabel metal2 884 -768 884 -768 0 net=12209
rlabel metal2 54 -770 54 -770 0 net=2153
rlabel metal2 401 -770 401 -770 0 net=3447
rlabel metal2 450 -770 450 -770 0 net=2955
rlabel metal2 933 -770 933 -770 0 net=7923
rlabel metal2 1157 -770 1157 -770 0 net=9023
rlabel metal2 1276 -770 1276 -770 0 net=10191
rlabel metal2 1430 -770 1430 -770 0 net=10321
rlabel metal2 142 -772 142 -772 0 net=7123
rlabel metal2 954 -772 954 -772 0 net=7847
rlabel metal2 1101 -772 1101 -772 0 net=8945
rlabel metal2 1283 -772 1283 -772 0 net=10209
rlabel metal2 1465 -772 1465 -772 0 net=12435
rlabel metal2 142 -774 142 -774 0 net=1711
rlabel metal2 359 -774 359 -774 0 net=2311
rlabel metal2 492 -774 492 -774 0 net=4804
rlabel metal2 576 -774 576 -774 0 net=4661
rlabel metal2 803 -774 803 -774 0 net=1
rlabel metal2 898 -774 898 -774 0 net=9537
rlabel metal2 1318 -774 1318 -774 0 net=10511
rlabel metal2 1521 -774 1521 -774 0 net=12225
rlabel metal2 44 -776 44 -776 0 net=4130
rlabel metal2 604 -776 604 -776 0 net=6661
rlabel metal2 814 -776 814 -776 0 net=6133
rlabel metal2 842 -776 842 -776 0 net=9964
rlabel metal2 1437 -776 1437 -776 0 net=11417
rlabel metal2 177 -778 177 -778 0 net=6541
rlabel metal2 901 -778 901 -778 0 net=13366
rlabel metal2 198 -780 198 -780 0 net=4905
rlabel metal2 534 -780 534 -780 0 net=5473
rlabel metal2 824 -780 824 -780 0 net=11776
rlabel metal2 548 -782 548 -782 0 net=6239
rlabel metal2 845 -782 845 -782 0 net=13201
rlabel metal2 583 -784 583 -784 0 net=5239
rlabel metal2 611 -784 611 -784 0 net=5189
rlabel metal2 782 -784 782 -784 0 net=10877
rlabel metal2 163 -786 163 -786 0 net=5966
rlabel metal2 625 -786 625 -786 0 net=5729
rlabel metal2 849 -786 849 -786 0 net=6674
rlabel metal2 1020 -786 1020 -786 0 net=11847
rlabel metal2 1507 -786 1507 -786 0 net=12171
rlabel metal2 163 -788 163 -788 0 net=12206
rlabel metal2 583 -790 583 -790 0 net=3783
rlabel metal2 625 -790 625 -790 0 net=12355
rlabel metal2 646 -792 646 -792 0 net=6503
rlabel metal2 912 -792 912 -792 0 net=6985
rlabel metal2 1010 -792 1010 -792 0 net=8063
rlabel metal2 1290 -792 1290 -792 0 net=10259
rlabel metal2 212 -794 212 -794 0 net=7493
rlabel metal2 1031 -794 1031 -794 0 net=8135
rlabel metal2 1185 -794 1185 -794 0 net=9281
rlabel metal2 1311 -794 1311 -794 0 net=10707
rlabel metal2 296 -796 296 -796 0 net=2931
rlabel metal2 1038 -796 1038 -796 0 net=7961
rlabel metal2 1108 -796 1108 -796 0 net=9115
rlabel metal2 1325 -796 1325 -796 0 net=10593
rlabel metal2 1416 -796 1416 -796 0 net=11391
rlabel metal2 166 -798 166 -798 0 net=13037
rlabel metal2 1332 -798 1332 -798 0 net=11521
rlabel metal2 1374 -798 1374 -798 0 net=11339
rlabel metal2 429 -800 429 -800 0 net=4631
rlabel metal2 744 -800 744 -800 0 net=6317
rlabel metal2 926 -800 926 -800 0 net=7639
rlabel metal2 1087 -800 1087 -800 0 net=8695
rlabel metal2 1192 -800 1192 -800 0 net=9739
rlabel metal2 1346 -800 1346 -800 0 net=10755
rlabel metal2 79 -802 79 -802 0 net=7877
rlabel metal2 1115 -802 1115 -802 0 net=9133
rlabel metal2 352 -804 352 -804 0 net=1589
rlabel metal2 509 -804 509 -804 0 net=7755
rlabel metal2 1066 -804 1066 -804 0 net=8527
rlabel metal2 1213 -804 1213 -804 0 net=9793
rlabel metal2 338 -806 338 -806 0 net=2123
rlabel metal2 691 -806 691 -806 0 net=6957
rlabel metal2 947 -806 947 -806 0 net=7607
rlabel metal2 1227 -806 1227 -806 0 net=9951
rlabel metal2 82 -808 82 -808 0 net=1997
rlabel metal2 744 -808 744 -808 0 net=5817
rlabel metal2 761 -808 761 -808 0 net=8701
rlabel metal2 1248 -808 1248 -808 0 net=10131
rlabel metal2 702 -810 702 -810 0 net=6083
rlabel metal2 761 -810 761 -810 0 net=8882
rlabel metal2 1255 -810 1255 -810 0 net=10693
rlabel metal2 789 -812 789 -812 0 net=7187
rlabel metal2 971 -812 971 -812 0 net=10041
rlabel metal2 821 -814 821 -814 0 net=6923
rlabel metal2 982 -814 982 -814 0 net=7905
rlabel metal2 821 -816 821 -816 0 net=11678
rlabel metal2 863 -818 863 -818 0 net=7253
rlabel metal2 989 -818 989 -818 0 net=7983
rlabel metal2 1129 -818 1129 -818 0 net=8897
rlabel metal2 1395 -818 1395 -818 0 net=11301
rlabel metal2 765 -820 765 -820 0 net=6331
rlabel metal2 989 -820 989 -820 0 net=7035
rlabel metal2 226 -822 226 -822 0 net=5761
rlabel metal2 1003 -822 1003 -822 0 net=8039
rlabel metal2 1150 -822 1150 -822 0 net=8795
rlabel metal2 226 -824 226 -824 0 net=2047
rlabel metal2 1024 -824 1024 -824 0 net=8955
rlabel metal2 240 -826 240 -826 0 net=7427
rlabel metal2 1150 -826 1150 -826 0 net=8289
rlabel metal2 1171 -826 1171 -826 0 net=10215
rlabel metal2 72 -828 72 -828 0 net=8409
rlabel metal2 1192 -828 1192 -828 0 net=12233
rlabel metal2 72 -830 72 -830 0 net=2899
rlabel metal2 240 -830 240 -830 0 net=1827
rlabel metal2 261 -830 261 -830 0 net=1761
rlabel metal2 891 -830 891 -830 0 net=7537
rlabel metal2 1059 -830 1059 -830 0 net=8493
rlabel metal2 44 -832 44 -832 0 net=2225
rlabel metal2 205 -832 205 -832 0 net=1517
rlabel metal2 331 -832 331 -832 0 net=5501
rlabel metal2 877 -832 877 -832 0 net=7459
rlabel metal2 968 -832 968 -832 0 net=10429
rlabel metal2 191 -834 191 -834 0 net=1923
rlabel metal2 380 -834 380 -834 0 net=4521
rlabel metal2 660 -834 660 -834 0 net=7359
rlabel metal2 128 -836 128 -836 0 net=1665
rlabel metal2 212 -836 212 -836 0 net=4983
rlabel metal2 579 -836 579 -836 0 net=4731
rlabel metal2 856 -836 856 -836 0 net=7239
rlabel metal2 786 -838 786 -838 0 net=6287
rlabel metal2 786 -840 786 -840 0 net=12222
rlabel metal2 1122 -842 1122 -842 0 net=11529
rlabel metal2 558 -844 558 -844 0 net=8023
rlabel metal2 86 -846 86 -846 0 net=3284
rlabel metal2 86 -848 86 -848 0 net=3563
rlabel metal2 23 -850 23 -850 0 net=4305
rlabel metal2 23 -852 23 -852 0 net=2921
rlabel metal2 187 -854 187 -854 0 net=2719
rlabel metal2 2 -865 2 -865 0 net=5059
rlabel metal2 86 -865 86 -865 0 net=3565
rlabel metal2 110 -865 110 -865 0 net=10498
rlabel metal2 1339 -865 1339 -865 0 net=9983
rlabel metal2 1339 -865 1339 -865 0 net=9983
rlabel metal2 1591 -865 1591 -865 0 net=12035
rlabel metal2 1724 -865 1724 -865 0 net=13203
rlabel metal2 1885 -865 1885 -865 0 net=9522
rlabel metal2 16 -867 16 -867 0 net=8107
rlabel metal2 16 -867 16 -867 0 net=8107
rlabel metal2 37 -867 37 -867 0 net=6474
rlabel metal2 86 -867 86 -867 0 net=1925
rlabel metal2 261 -867 261 -867 0 net=1763
rlabel metal2 310 -867 310 -867 0 net=2154
rlabel metal2 968 -867 968 -867 0 net=7241
rlabel metal2 968 -867 968 -867 0 net=7241
rlabel metal2 1006 -867 1006 -867 0 net=12982
rlabel metal2 1780 -867 1780 -867 0 net=11738
rlabel metal2 1829 -867 1829 -867 0 net=8707
rlabel metal2 30 -869 30 -869 0 net=2215
rlabel metal2 114 -869 114 -869 0 net=4412
rlabel metal2 135 -869 135 -869 0 net=3734
rlabel metal2 516 -869 516 -869 0 net=12082
rlabel metal2 1703 -869 1703 -869 0 net=12661
rlabel metal2 1787 -869 1787 -869 0 net=13617
rlabel metal2 1836 -869 1836 -869 0 net=10261
rlabel metal2 30 -871 30 -871 0 net=2049
rlabel metal2 261 -871 261 -871 0 net=1661
rlabel metal2 310 -871 310 -871 0 net=2957
rlabel metal2 460 -871 460 -871 0 net=166
rlabel metal2 37 -873 37 -873 0 net=2901
rlabel metal2 121 -873 121 -873 0 net=1667
rlabel metal2 156 -873 156 -873 0 net=6088
rlabel metal2 828 -873 828 -873 0 net=11586
rlabel metal2 1633 -873 1633 -873 0 net=13759
rlabel metal2 1892 -873 1892 -873 0 net=11373
rlabel metal2 51 -875 51 -875 0 net=1639
rlabel metal2 163 -875 163 -875 0 net=1518
rlabel metal2 275 -875 275 -875 0 net=2353
rlabel metal2 338 -875 338 -875 0 net=1998
rlabel metal2 450 -875 450 -875 0 net=2991
rlabel metal2 779 -875 779 -875 0 net=7608
rlabel metal2 1083 -875 1083 -875 0 net=12924
rlabel metal2 1759 -875 1759 -875 0 net=13573
rlabel metal2 47 -877 47 -877 0 net=7557
rlabel metal2 1108 -877 1108 -877 0 net=7985
rlabel metal2 1136 -877 1136 -877 0 net=8137
rlabel metal2 1136 -877 1136 -877 0 net=8137
rlabel metal2 1153 -877 1153 -877 0 net=12120
rlabel metal2 1717 -877 1717 -877 0 net=13125
rlabel metal2 1801 -877 1801 -877 0 net=6765
rlabel metal2 51 -879 51 -879 0 net=1875
rlabel metal2 177 -879 177 -879 0 net=7538
rlabel metal2 1031 -879 1031 -879 0 net=11282
rlabel metal2 1619 -879 1619 -879 0 net=12173
rlabel metal2 1752 -879 1752 -879 0 net=13451
rlabel metal2 1843 -879 1843 -879 0 net=11593
rlabel metal2 65 -881 65 -881 0 net=3964
rlabel metal2 572 -881 572 -881 0 net=13038
rlabel metal2 1353 -881 1353 -881 0 net=11523
rlabel metal2 1633 -881 1633 -881 0 net=11919
rlabel metal2 65 -883 65 -883 0 net=301
rlabel metal2 1031 -883 1031 -883 0 net=10694
rlabel metal2 1556 -883 1556 -883 0 net=11825
rlabel metal2 1654 -883 1654 -883 0 net=12235
rlabel metal2 1794 -883 1794 -883 0 net=13649
rlabel metal2 1850 -883 1850 -883 0 net=6388
rlabel metal2 72 -885 72 -885 0 net=4079
rlabel metal2 247 -885 247 -885 0 net=1591
rlabel metal2 492 -885 492 -885 0 net=4662
rlabel metal2 684 -885 684 -885 0 net=7907
rlabel metal2 915 -885 915 -885 0 net=9177
rlabel metal2 1360 -885 1360 -885 0 net=10055
rlabel metal2 1661 -885 1661 -885 0 net=12357
rlabel metal2 1738 -885 1738 -885 0 net=13317
rlabel metal2 1857 -885 1857 -885 0 net=6467
rlabel metal2 93 -887 93 -887 0 net=1685
rlabel metal2 177 -887 177 -887 0 net=7369
rlabel metal2 688 -887 688 -887 0 net=10660
rlabel metal2 1500 -887 1500 -887 0 net=11303
rlabel metal2 1577 -887 1577 -887 0 net=12859
rlabel metal2 128 -889 128 -889 0 net=2457
rlabel metal2 268 -889 268 -889 0 net=1703
rlabel metal2 492 -889 492 -889 0 net=4115
rlabel metal2 576 -889 576 -889 0 net=7360
rlabel metal2 919 -889 919 -889 0 net=9910
rlabel metal2 1108 -889 1108 -889 0 net=8665
rlabel metal2 1220 -889 1220 -889 0 net=8727
rlabel metal2 1220 -889 1220 -889 0 net=8727
rlabel metal2 1297 -889 1297 -889 0 net=9405
rlabel metal2 1381 -889 1381 -889 0 net=10185
rlabel metal2 1668 -889 1668 -889 0 net=13439
rlabel metal2 1808 -889 1808 -889 0 net=13737
rlabel metal2 156 -891 156 -891 0 net=9493
rlabel metal2 1430 -891 1430 -891 0 net=10757
rlabel metal2 1521 -891 1521 -891 0 net=11419
rlabel metal2 1591 -891 1591 -891 0 net=13061
rlabel metal2 180 -893 180 -893 0 net=4522
rlabel metal2 387 -893 387 -893 0 net=2248
rlabel metal2 705 -893 705 -893 0 net=3816
rlabel metal2 985 -893 985 -893 0 net=12837
rlabel metal2 58 -895 58 -895 0 net=2371
rlabel metal2 429 -895 429 -895 0 net=3785
rlabel metal2 604 -895 604 -895 0 net=5241
rlabel metal2 688 -895 688 -895 0 net=7037
rlabel metal2 1003 -895 1003 -895 0 net=7429
rlabel metal2 1034 -895 1034 -895 0 net=10210
rlabel metal2 1451 -895 1451 -895 0 net=10815
rlabel metal2 1521 -895 1521 -895 0 net=11945
rlabel metal2 1605 -895 1605 -895 0 net=12149
rlabel metal2 1689 -895 1689 -895 0 net=12549
rlabel metal2 187 -897 187 -897 0 net=749
rlabel metal2 604 -897 604 -897 0 net=10588
rlabel metal2 1640 -897 1640 -897 0 net=12227
rlabel metal2 1696 -897 1696 -897 0 net=12621
rlabel metal2 191 -899 191 -899 0 net=6333
rlabel metal2 877 -899 877 -899 0 net=6349
rlabel metal2 1374 -899 1374 -899 0 net=10133
rlabel metal2 1465 -899 1465 -899 0 net=12437
rlabel metal2 198 -901 198 -901 0 net=5653
rlabel metal2 583 -901 583 -901 0 net=6174
rlabel metal2 723 -901 723 -901 0 net=7633
rlabel metal2 1402 -901 1402 -901 0 net=10513
rlabel metal2 1465 -901 1465 -901 0 net=11615
rlabel metal2 1549 -901 1549 -901 0 net=13187
rlabel metal2 170 -903 170 -903 0 net=1897
rlabel metal2 201 -903 201 -903 0 net=2286
rlabel metal2 338 -903 338 -903 0 net=2453
rlabel metal2 478 -903 478 -903 0 net=5863
rlabel metal2 618 -903 618 -903 0 net=5318
rlabel metal2 726 -903 726 -903 0 net=12263
rlabel metal2 170 -905 170 -905 0 net=3437
rlabel metal2 366 -905 366 -905 0 net=1959
rlabel metal2 366 -905 366 -905 0 net=1959
rlabel metal2 394 -905 394 -905 0 net=2721
rlabel metal2 485 -905 485 -905 0 net=3663
rlabel metal2 586 -905 586 -905 0 net=7556
rlabel metal2 1059 -905 1059 -905 0 net=10431
rlabel metal2 1535 -905 1535 -905 0 net=11531
rlabel metal2 1647 -905 1647 -905 0 net=10323
rlabel metal2 184 -907 184 -907 0 net=5383
rlabel metal2 408 -907 408 -907 0 net=2313
rlabel metal2 495 -907 495 -907 0 net=10091
rlabel metal2 782 -907 782 -907 0 net=12267
rlabel metal2 184 -909 184 -909 0 net=5502
rlabel metal2 506 -909 506 -909 0 net=3407
rlabel metal2 590 -909 590 -909 0 net=4633
rlabel metal2 674 -909 674 -909 0 net=7757
rlabel metal2 1041 -909 1041 -909 0 net=11364
rlabel metal2 205 -911 205 -911 0 net=4307
rlabel metal2 240 -911 240 -911 0 net=1829
rlabel metal2 422 -911 422 -911 0 net=7067
rlabel metal2 513 -911 513 -911 0 net=6319
rlabel metal2 856 -911 856 -911 0 net=6289
rlabel metal2 1409 -911 1409 -911 0 net=10595
rlabel metal2 1472 -911 1472 -911 0 net=10949
rlabel metal2 212 -913 212 -913 0 net=4985
rlabel metal2 527 -913 527 -913 0 net=3458
rlabel metal2 618 -913 618 -913 0 net=2789
rlabel metal2 831 -913 831 -913 0 net=9579
rlabel metal2 1395 -913 1395 -913 0 net=10217
rlabel metal2 1416 -913 1416 -913 0 net=11341
rlabel metal2 142 -915 142 -915 0 net=1713
rlabel metal2 240 -915 240 -915 0 net=2035
rlabel metal2 415 -915 415 -915 0 net=2537
rlabel metal2 499 -915 499 -915 0 net=3639
rlabel metal2 534 -915 534 -915 0 net=5475
rlabel metal2 621 -915 621 -915 0 net=13533
rlabel metal2 226 -917 226 -917 0 net=5899
rlabel metal2 537 -917 537 -917 0 net=7906
rlabel metal2 1255 -917 1255 -917 0 net=8957
rlabel metal2 1423 -917 1423 -917 0 net=10709
rlabel metal2 1563 -917 1563 -917 0 net=12567
rlabel metal2 268 -919 268 -919 0 net=3179
rlabel metal2 625 -919 625 -919 0 net=6084
rlabel metal2 758 -919 758 -919 0 net=7435
rlabel metal2 1059 -919 1059 -919 0 net=8931
rlabel metal2 1318 -919 1318 -919 0 net=9795
rlabel metal2 1486 -919 1486 -919 0 net=11107
rlabel metal2 282 -921 282 -921 0 net=4907
rlabel metal2 415 -921 415 -921 0 net=7925
rlabel metal2 1115 -921 1115 -921 0 net=8529
rlabel metal2 1276 -921 1276 -921 0 net=9135
rlabel metal2 1346 -921 1346 -921 0 net=10043
rlabel metal2 1486 -921 1486 -921 0 net=10017
rlabel metal2 289 -923 289 -923 0 net=1719
rlabel metal2 359 -923 359 -923 0 net=4567
rlabel metal2 289 -925 289 -925 0 net=2125
rlabel metal2 499 -925 499 -925 0 net=5029
rlabel metal2 758 -925 758 -925 0 net=6125
rlabel metal2 775 -925 775 -925 0 net=9529
rlabel metal2 254 -927 254 -927 0 net=2363
rlabel metal2 541 -927 541 -927 0 net=4511
rlabel metal2 625 -927 625 -927 0 net=4733
rlabel metal2 709 -927 709 -927 0 net=6283
rlabel metal2 856 -927 856 -927 0 net=11631
rlabel metal2 1017 -927 1017 -927 0 net=7641
rlabel metal2 1087 -927 1087 -927 0 net=7879
rlabel metal2 1129 -927 1129 -927 0 net=8041
rlabel metal2 1276 -927 1276 -927 0 net=10193
rlabel metal2 1493 -927 1493 -927 0 net=11123
rlabel metal2 58 -929 58 -929 0 net=7167
rlabel metal2 632 -929 632 -929 0 net=4561
rlabel metal2 632 -929 632 -929 0 net=4561
rlabel metal2 639 -929 639 -929 0 net=6933
rlabel metal2 1052 -929 1052 -929 0 net=7849
rlabel metal2 1094 -929 1094 -929 0 net=7963
rlabel metal2 1122 -929 1122 -929 0 net=8025
rlabel metal2 1164 -929 1164 -929 0 net=8411
rlabel metal2 1283 -929 1283 -929 0 net=9283
rlabel metal2 1367 -929 1367 -929 0 net=10075
rlabel metal2 1493 -929 1493 -929 0 net=12405
rlabel metal2 254 -931 254 -931 0 net=1929
rlabel metal2 639 -931 639 -931 0 net=5595
rlabel metal2 814 -931 814 -931 0 net=5731
rlabel metal2 1171 -931 1171 -931 0 net=8495
rlabel metal2 1241 -931 1241 -931 0 net=8831
rlabel metal2 1304 -931 1304 -931 0 net=9539
rlabel metal2 1507 -931 1507 -931 0 net=11393
rlabel metal2 1682 -931 1682 -931 0 net=12097
rlabel metal2 142 -933 142 -933 0 net=6359
rlabel metal2 821 -933 821 -933 0 net=6241
rlabel metal2 863 -933 863 -933 0 net=6925
rlabel metal2 922 -933 922 -933 0 net=12465
rlabel metal2 296 -935 296 -935 0 net=2933
rlabel metal2 520 -935 520 -935 0 net=6019
rlabel metal2 716 -935 716 -935 0 net=5469
rlabel metal2 740 -935 740 -935 0 net=10961
rlabel metal2 296 -937 296 -937 0 net=2827
rlabel metal2 544 -937 544 -937 0 net=3699
rlabel metal2 646 -937 646 -937 0 net=6669
rlabel metal2 922 -937 922 -937 0 net=6689
rlabel metal2 166 -939 166 -939 0 net=13367
rlabel metal2 926 -939 926 -939 0 net=6959
rlabel metal2 926 -939 926 -939 0 net=6959
rlabel metal2 933 -939 933 -939 0 net=7125
rlabel metal2 933 -939 933 -939 0 net=7125
rlabel metal2 947 -939 947 -939 0 net=7189
rlabel metal2 1003 -939 1003 -939 0 net=8185
rlabel metal2 1311 -939 1311 -939 0 net=9741
rlabel metal2 1458 -939 1458 -939 0 net=10933
rlabel metal2 1594 -939 1594 -939 0 net=1
rlabel metal2 317 -941 317 -941 0 net=4589
rlabel metal2 401 -941 401 -941 0 net=3449
rlabel metal2 660 -941 660 -941 0 net=7163
rlabel metal2 947 -941 947 -941 0 net=7255
rlabel metal2 1062 -941 1062 -941 0 net=10878
rlabel metal2 149 -943 149 -943 0 net=2227
rlabel metal2 401 -943 401 -943 0 net=2567
rlabel metal2 464 -943 464 -943 0 net=5281
rlabel metal2 702 -943 702 -943 0 net=8761
rlabel metal2 1262 -943 1262 -943 0 net=9025
rlabel metal2 100 -945 100 -945 0 net=2259
rlabel metal2 373 -945 373 -945 0 net=5951
rlabel metal2 730 -945 730 -945 0 net=7495
rlabel metal2 1143 -945 1143 -945 0 net=8211
rlabel metal2 1213 -945 1213 -945 0 net=8703
rlabel metal2 9 -947 9 -947 0 net=4825
rlabel metal2 107 -947 107 -947 0 net=2333
rlabel metal2 390 -947 390 -947 0 net=4377
rlabel metal2 744 -947 744 -947 0 net=5818
rlabel metal2 789 -947 789 -947 0 net=12335
rlabel metal2 891 -947 891 -947 0 net=7461
rlabel metal2 1080 -947 1080 -947 0 net=8427
rlabel metal2 1157 -947 1157 -947 0 net=8947
rlabel metal2 9 -949 9 -949 0 net=2923
rlabel metal2 44 -949 44 -949 0 net=4995
rlabel metal2 135 -949 135 -949 0 net=2591
rlabel metal2 611 -949 611 -949 0 net=5763
rlabel metal2 800 -949 800 -949 0 net=5061
rlabel metal2 954 -949 954 -949 0 net=6987
rlabel metal2 1010 -949 1010 -949 0 net=13680
rlabel metal2 23 -951 23 -951 0 net=4217
rlabel metal2 611 -951 611 -951 0 net=5191
rlabel metal2 744 -951 744 -951 0 net=9116
rlabel metal2 667 -953 667 -953 0 net=4867
rlabel metal2 761 -953 761 -953 0 net=10997
rlabel metal2 667 -955 667 -955 0 net=6499
rlabel metal2 884 -955 884 -955 0 net=6505
rlabel metal2 961 -955 961 -955 0 net=7345
rlabel metal2 1034 -955 1034 -955 0 net=10763
rlabel metal2 765 -957 765 -957 0 net=5762
rlabel metal2 996 -957 996 -957 0 net=7017
rlabel metal2 1080 -957 1080 -957 0 net=13371
rlabel metal2 737 -959 737 -959 0 net=4183
rlabel metal2 772 -959 772 -959 0 net=8064
rlabel metal2 807 -961 807 -961 0 net=6663
rlabel metal2 1157 -961 1157 -961 0 net=9911
rlabel metal2 793 -963 793 -963 0 net=6197
rlabel metal2 835 -963 835 -963 0 net=6135
rlabel metal2 884 -963 884 -963 0 net=6543
rlabel metal2 1185 -963 1185 -963 0 net=8697
rlabel metal2 1227 -963 1227 -963 0 net=8797
rlabel metal2 54 -965 54 -965 0 net=6413
rlabel metal2 1150 -965 1150 -965 0 net=8291
rlabel metal2 1248 -965 1248 -965 0 net=8899
rlabel metal2 236 -967 236 -967 0 net=8513
rlabel metal2 1262 -967 1262 -967 0 net=12211
rlabel metal2 439 -969 439 -969 0 net=6461
rlabel metal2 1437 -969 1437 -969 0 net=11849
rlabel metal2 793 -971 793 -971 0 net=7043
rlabel metal2 1332 -971 1332 -971 0 net=9953
rlabel metal2 1199 -973 1199 -973 0 net=9237
rlabel metal2 628 -975 628 -975 0 net=8459
rlabel metal2 47 -986 47 -986 0 net=5952
rlabel metal2 733 -986 733 -986 0 net=968
rlabel metal2 775 -986 775 -986 0 net=6242
rlabel metal2 866 -986 866 -986 0 net=9796
rlabel metal2 1444 -986 1444 -986 0 net=10515
rlabel metal2 1444 -986 1444 -986 0 net=10515
rlabel metal2 1745 -986 1745 -986 0 net=10950
rlabel metal2 1927 -986 1927 -986 0 net=6691
rlabel metal2 58 -988 58 -988 0 net=7168
rlabel metal2 457 -988 457 -988 0 net=529
rlabel metal2 541 -988 541 -988 0 net=4735
rlabel metal2 656 -988 656 -988 0 net=8958
rlabel metal2 1710 -988 1710 -988 0 net=10325
rlabel metal2 1867 -988 1867 -988 0 net=6468
rlabel metal2 1927 -988 1927 -988 0 net=6767
rlabel metal2 1941 -988 1941 -988 0 net=8709
rlabel metal2 58 -990 58 -990 0 net=3439
rlabel metal2 240 -990 240 -990 0 net=2036
rlabel metal2 709 -990 709 -990 0 net=6021
rlabel metal2 870 -990 870 -990 0 net=6136
rlabel metal2 919 -990 919 -990 0 net=10134
rlabel metal2 1710 -990 1710 -990 0 net=12663
rlabel metal2 1878 -990 1878 -990 0 net=11594
rlabel metal2 1948 -990 1948 -990 0 net=10263
rlabel metal2 68 -992 68 -992 0 net=5384
rlabel metal2 443 -992 443 -992 0 net=2723
rlabel metal2 485 -992 485 -992 0 net=2314
rlabel metal2 625 -992 625 -992 0 net=9954
rlabel metal2 1584 -992 1584 -992 0 net=9531
rlabel metal2 1948 -992 1948 -992 0 net=11375
rlabel metal2 30 -994 30 -994 0 net=2050
rlabel metal2 485 -994 485 -994 0 net=2791
rlabel metal2 674 -994 674 -994 0 net=7759
rlabel metal2 716 -994 716 -994 0 net=5471
rlabel metal2 779 -994 779 -994 0 net=10093
rlabel metal2 1493 -994 1493 -994 0 net=12407
rlabel metal2 30 -996 30 -996 0 net=1877
rlabel metal2 72 -996 72 -996 0 net=4080
rlabel metal2 513 -996 513 -996 0 net=6321
rlabel metal2 667 -996 667 -996 0 net=6501
rlabel metal2 737 -996 737 -996 0 net=6126
rlabel metal2 761 -996 761 -996 0 net=12236
rlabel metal2 51 -998 51 -998 0 net=2935
rlabel metal2 478 -998 478 -998 0 net=4987
rlabel metal2 674 -998 674 -998 0 net=8413
rlabel metal2 1241 -998 1241 -998 0 net=8763
rlabel metal2 1276 -998 1276 -998 0 net=10195
rlabel metal2 1493 -998 1493 -998 0 net=10817
rlabel metal2 1724 -998 1724 -998 0 net=13761
rlabel metal2 72 -1000 72 -1000 0 net=5143
rlabel metal2 681 -1000 681 -1000 0 net=8042
rlabel metal2 1241 -1000 1241 -1000 0 net=8799
rlabel metal2 1276 -1000 1276 -1000 0 net=8901
rlabel metal2 1346 -1000 1346 -1000 0 net=9285
rlabel metal2 1346 -1000 1346 -1000 0 net=9285
rlabel metal2 1374 -1000 1374 -1000 0 net=9581
rlabel metal2 1374 -1000 1374 -1000 0 net=9581
rlabel metal2 1409 -1000 1409 -1000 0 net=10219
rlabel metal2 1500 -1000 1500 -1000 0 net=10935
rlabel metal2 82 -1002 82 -1002 0 net=6934
rlabel metal2 1020 -1002 1020 -1002 0 net=8530
rlabel metal2 1367 -1002 1367 -1002 0 net=9541
rlabel metal2 1507 -1002 1507 -1002 0 net=10999
rlabel metal2 86 -1004 86 -1004 0 net=1926
rlabel metal2 149 -1004 149 -1004 0 net=2261
rlabel metal2 240 -1004 240 -1004 0 net=2569
rlabel metal2 408 -1004 408 -1004 0 net=4117
rlabel metal2 513 -1004 513 -1004 0 net=5193
rlabel metal2 646 -1004 646 -1004 0 net=6671
rlabel metal2 1514 -1004 1514 -1004 0 net=11343
rlabel metal2 9 -1006 9 -1006 0 net=2925
rlabel metal2 93 -1006 93 -1006 0 net=3567
rlabel metal2 261 -1006 261 -1006 0 net=1663
rlabel metal2 261 -1006 261 -1006 0 net=1663
rlabel metal2 282 -1006 282 -1006 0 net=4908
rlabel metal2 737 -1006 737 -1006 0 net=10459
rlabel metal2 1535 -1006 1535 -1006 0 net=11109
rlabel metal2 9 -1008 9 -1008 0 net=5901
rlabel metal2 282 -1008 282 -1008 0 net=1705
rlabel metal2 478 -1008 478 -1008 0 net=5529
rlabel metal2 786 -1008 786 -1008 0 net=5764
rlabel metal2 968 -1008 968 -1008 0 net=7243
rlabel metal2 1535 -1008 1535 -1008 0 net=11525
rlabel metal2 79 -1010 79 -1010 0 net=2217
rlabel metal2 156 -1010 156 -1010 0 net=7949
rlabel metal2 492 -1010 492 -1010 0 net=7497
rlabel metal2 747 -1010 747 -1010 0 net=8704
rlabel metal2 1598 -1010 1598 -1010 0 net=11921
rlabel metal2 79 -1012 79 -1012 0 net=7634
rlabel metal2 1255 -1012 1255 -1012 0 net=8933
rlabel metal2 1451 -1012 1451 -1012 0 net=10597
rlabel metal2 68 -1014 68 -1014 0 net=11539
rlabel metal2 96 -1016 96 -1016 0 net=525
rlabel metal2 863 -1016 863 -1016 0 net=6927
rlabel metal2 891 -1016 891 -1016 0 net=6665
rlabel metal2 107 -1018 107 -1018 0 net=2459
rlabel metal2 142 -1018 142 -1018 0 net=304
rlabel metal2 226 -1018 226 -1018 0 net=7165
rlabel metal2 681 -1018 681 -1018 0 net=10432
rlabel metal2 128 -1020 128 -1020 0 net=2958
rlabel metal2 345 -1020 345 -1020 0 net=4591
rlabel metal2 506 -1020 506 -1020 0 net=7069
rlabel metal2 982 -1020 982 -1020 0 net=13204
rlabel metal2 142 -1022 142 -1022 0 net=6335
rlabel metal2 268 -1022 268 -1022 0 net=3180
rlabel metal2 842 -1022 842 -1022 0 net=12336
rlabel metal2 894 -1022 894 -1022 0 net=6462
rlabel metal2 912 -1022 912 -1022 0 net=10076
rlabel metal2 37 -1024 37 -1024 0 net=2903
rlabel metal2 296 -1024 296 -1024 0 net=2828
rlabel metal2 548 -1024 548 -1024 0 net=3409
rlabel metal2 548 -1024 548 -1024 0 net=3409
rlabel metal2 565 -1024 565 -1024 0 net=4901
rlabel metal2 632 -1024 632 -1024 0 net=4563
rlabel metal2 702 -1024 702 -1024 0 net=4829
rlabel metal2 751 -1024 751 -1024 0 net=10764
rlabel metal2 37 -1026 37 -1026 0 net=3451
rlabel metal2 499 -1026 499 -1026 0 net=5031
rlabel metal2 569 -1026 569 -1026 0 net=3700
rlabel metal2 1108 -1026 1108 -1026 0 net=8667
rlabel metal2 1160 -1026 1160 -1026 0 net=13188
rlabel metal2 156 -1028 156 -1028 0 net=3749
rlabel metal2 1108 -1028 1108 -1028 0 net=7987
rlabel metal2 1136 -1028 1136 -1028 0 net=8139
rlabel metal2 1773 -1028 1773 -1028 0 net=13281
rlabel metal2 191 -1030 191 -1030 0 net=2867
rlabel metal2 303 -1030 303 -1030 0 net=1765
rlabel metal2 387 -1030 387 -1030 0 net=3664
rlabel metal2 579 -1030 579 -1030 0 net=12049
rlabel metal2 198 -1032 198 -1032 0 net=1899
rlabel metal2 380 -1032 380 -1032 0 net=2373
rlabel metal2 397 -1032 397 -1032 0 net=6645
rlabel metal2 919 -1032 919 -1032 0 net=6961
rlabel metal2 940 -1032 940 -1032 0 net=13574
rlabel metal2 121 -1034 121 -1034 0 net=1669
rlabel metal2 205 -1034 205 -1034 0 net=4309
rlabel metal2 499 -1034 499 -1034 0 net=3641
rlabel metal2 583 -1034 583 -1034 0 net=5477
rlabel metal2 583 -1034 583 -1034 0 net=5477
rlabel metal2 618 -1034 618 -1034 0 net=4219
rlabel metal2 1139 -1034 1139 -1034 0 net=10962
rlabel metal2 100 -1036 100 -1036 0 net=4827
rlabel metal2 646 -1036 646 -1036 0 net=6284
rlabel metal2 877 -1036 877 -1036 0 net=6351
rlabel metal2 905 -1036 905 -1036 0 net=13369
rlabel metal2 44 -1038 44 -1038 0 net=4997
rlabel metal2 114 -1038 114 -1038 0 net=1641
rlabel metal2 219 -1038 219 -1038 0 net=9351
rlabel metal2 954 -1038 954 -1038 0 net=6506
rlabel metal2 1010 -1038 1010 -1038 0 net=12983
rlabel metal2 1808 -1038 1808 -1038 0 net=13619
rlabel metal2 114 -1040 114 -1040 0 net=7371
rlabel metal2 205 -1040 205 -1040 0 net=2085
rlabel metal2 982 -1040 982 -1040 0 net=7019
rlabel metal2 1010 -1040 1010 -1040 0 net=7463
rlabel metal2 1059 -1040 1059 -1040 0 net=10710
rlabel metal2 1591 -1040 1591 -1040 0 net=13063
rlabel metal2 177 -1042 177 -1042 0 net=3787
rlabel metal2 450 -1042 450 -1042 0 net=2993
rlabel metal2 520 -1042 520 -1042 0 net=5282
rlabel metal2 688 -1042 688 -1042 0 net=7039
rlabel metal2 961 -1042 961 -1042 0 net=7347
rlabel metal2 1013 -1042 1013 -1042 0 net=6063
rlabel metal2 1220 -1042 1220 -1042 0 net=8729
rlabel metal2 1297 -1042 1297 -1042 0 net=8949
rlabel metal2 1360 -1042 1360 -1042 0 net=9495
rlabel metal2 233 -1044 233 -1044 0 net=1813
rlabel metal2 520 -1044 520 -1044 0 net=925
rlabel metal2 985 -1044 985 -1044 0 net=10186
rlabel metal2 254 -1046 254 -1046 0 net=1931
rlabel metal2 352 -1046 352 -1046 0 net=2365
rlabel metal2 688 -1046 688 -1046 0 net=2197
rlabel metal2 1206 -1046 1206 -1046 0 net=8497
rlabel metal2 1262 -1046 1262 -1046 0 net=12213
rlabel metal2 254 -1048 254 -1048 0 net=1831
rlabel metal2 352 -1048 352 -1048 0 net=3321
rlabel metal2 695 -1048 695 -1048 0 net=4868
rlabel metal2 1199 -1048 1199 -1048 0 net=8461
rlabel metal2 1213 -1048 1213 -1048 0 net=8699
rlabel metal2 1304 -1048 1304 -1048 0 net=9027
rlabel metal2 1353 -1048 1353 -1048 0 net=9407
rlabel metal2 1472 -1048 1472 -1048 0 net=10759
rlabel metal2 1549 -1048 1549 -1048 0 net=13127
rlabel metal2 366 -1050 366 -1050 0 net=1961
rlabel metal2 401 -1050 401 -1050 0 net=2539
rlabel metal2 607 -1050 607 -1050 0 net=3897
rlabel metal2 723 -1050 723 -1050 0 net=8163
rlabel metal2 1213 -1050 1213 -1050 0 net=8833
rlabel metal2 1479 -1050 1479 -1050 0 net=11305
rlabel metal2 1591 -1050 1591 -1050 0 net=12229
rlabel metal2 1787 -1050 1787 -1050 0 net=13373
rlabel metal2 275 -1052 275 -1052 0 net=2355
rlabel metal2 653 -1052 653 -1052 0 net=5243
rlabel metal2 751 -1052 751 -1052 0 net=11632
rlabel metal2 877 -1052 877 -1052 0 net=6545
rlabel metal2 989 -1052 989 -1052 0 net=7191
rlabel metal2 989 -1052 989 -1052 0 net=7191
rlabel metal2 1003 -1052 1003 -1052 0 net=9357
rlabel metal2 1465 -1052 1465 -1052 0 net=11617
rlabel metal2 1563 -1052 1563 -1052 0 net=12569
rlabel metal2 1815 -1052 1815 -1052 0 net=13651
rlabel metal2 16 -1054 16 -1054 0 net=8109
rlabel metal2 1003 -1054 1003 -1054 0 net=7437
rlabel metal2 1048 -1054 1048 -1054 0 net=12438
rlabel metal2 16 -1056 16 -1056 0 net=2929
rlabel metal2 275 -1056 275 -1056 0 net=2229
rlabel metal2 324 -1056 324 -1056 0 net=4533
rlabel metal2 1052 -1056 1052 -1056 0 net=7643
rlabel metal2 1122 -1056 1122 -1056 0 net=8027
rlabel metal2 1150 -1056 1150 -1056 0 net=12098
rlabel metal2 1696 -1056 1696 -1056 0 net=12265
rlabel metal2 317 -1058 317 -1058 0 net=1815
rlabel metal2 782 -1058 782 -1058 0 net=8925
rlabel metal2 1563 -1058 1563 -1058 0 net=11851
rlabel metal2 1682 -1058 1682 -1058 0 net=12551
rlabel metal2 1759 -1058 1759 -1058 0 net=13453
rlabel metal2 338 -1060 338 -1060 0 net=2455
rlabel metal2 1150 -1060 1150 -1060 0 net=10733
rlabel metal2 1626 -1060 1626 -1060 0 net=12037
rlabel metal2 1696 -1060 1696 -1060 0 net=12623
rlabel metal2 331 -1062 331 -1062 0 net=1721
rlabel metal2 366 -1062 366 -1062 0 net=2293
rlabel metal2 744 -1062 744 -1062 0 net=5063
rlabel metal2 807 -1062 807 -1062 0 net=6199
rlabel metal2 1017 -1062 1017 -1062 0 net=12787
rlabel metal2 135 -1064 135 -1064 0 net=2593
rlabel metal2 765 -1064 765 -1064 0 net=4185
rlabel metal2 835 -1064 835 -1064 0 net=6415
rlabel metal2 1031 -1064 1031 -1064 0 net=12925
rlabel metal2 135 -1066 135 -1066 0 net=7927
rlabel metal2 597 -1066 597 -1066 0 net=5865
rlabel metal2 793 -1066 793 -1066 0 net=7045
rlabel metal2 1038 -1066 1038 -1066 0 net=5732
rlabel metal2 1227 -1066 1227 -1066 0 net=9067
rlabel metal2 1612 -1066 1612 -1066 0 net=11827
rlabel metal2 359 -1068 359 -1068 0 net=4569
rlabel metal2 628 -1068 628 -1068 0 net=6425
rlabel metal2 842 -1068 842 -1068 0 net=7881
rlabel metal2 1227 -1068 1227 -1068 0 net=12860
rlabel metal2 359 -1070 359 -1070 0 net=2335
rlabel metal2 415 -1070 415 -1070 0 net=4379
rlabel metal2 639 -1070 639 -1070 0 net=5597
rlabel metal2 800 -1070 800 -1070 0 net=4909
rlabel metal2 1041 -1070 1041 -1070 0 net=11394
rlabel metal2 1836 -1070 1836 -1070 0 net=13739
rlabel metal2 247 -1072 247 -1072 0 net=1593
rlabel metal2 639 -1072 639 -1072 0 net=1999
rlabel metal2 828 -1072 828 -1072 0 net=7909
rlabel metal2 1115 -1072 1115 -1072 0 net=8187
rlabel metal2 1521 -1072 1521 -1072 0 net=11947
rlabel metal2 1640 -1072 1640 -1072 0 net=12151
rlabel metal2 1822 -1072 1822 -1072 0 net=13535
rlabel metal2 184 -1074 184 -1074 0 net=3019
rlabel metal2 289 -1074 289 -1074 0 net=2127
rlabel metal2 653 -1074 653 -1074 0 net=11423
rlabel metal2 1661 -1074 1661 -1074 0 net=12269
rlabel metal2 163 -1076 163 -1076 0 net=1687
rlabel metal2 212 -1076 212 -1076 0 net=1715
rlabel metal2 684 -1076 684 -1076 0 net=10875
rlabel metal2 23 -1078 23 -1078 0 net=4218
rlabel metal2 849 -1078 849 -1078 0 net=6290
rlabel metal2 1675 -1078 1675 -1078 0 net=12175
rlabel metal2 23 -1080 23 -1080 0 net=4345
rlabel metal2 947 -1080 947 -1080 0 net=7257
rlabel metal2 1059 -1080 1059 -1080 0 net=7965
rlabel metal2 1143 -1080 1143 -1080 0 net=8429
rlabel metal2 1381 -1080 1381 -1080 0 net=9743
rlabel metal2 1675 -1080 1675 -1080 0 net=12467
rlabel metal2 163 -1082 163 -1082 0 net=4635
rlabel metal2 947 -1082 947 -1082 0 net=6989
rlabel metal2 1024 -1082 1024 -1082 0 net=7431
rlabel metal2 1066 -1082 1066 -1082 0 net=7559
rlabel metal2 1143 -1082 1143 -1082 0 net=8293
rlabel metal2 1388 -1082 1388 -1082 0 net=9913
rlabel metal2 1577 -1082 1577 -1082 0 net=11421
rlabel metal2 555 -1084 555 -1084 0 net=5655
rlabel metal2 863 -1084 863 -1084 0 net=7795
rlabel metal2 1073 -1084 1073 -1084 0 net=7851
rlabel metal2 1185 -1084 1185 -1084 0 net=10783
rlabel metal2 1339 -1084 1339 -1084 0 net=9985
rlabel metal2 1542 -1084 1542 -1084 0 net=11125
rlabel metal2 555 -1086 555 -1086 0 net=4513
rlabel metal2 740 -1086 740 -1086 0 net=7887
rlabel metal2 1332 -1086 1332 -1086 0 net=9239
rlabel metal2 1542 -1086 1542 -1086 0 net=11533
rlabel metal2 576 -1088 576 -1088 0 net=8514
rlabel metal2 1325 -1088 1325 -1088 0 net=9179
rlabel metal2 1605 -1088 1605 -1088 0 net=12359
rlabel metal2 740 -1090 740 -1090 0 net=10056
rlabel metal2 1717 -1090 1717 -1090 0 net=12839
rlabel metal2 65 -1092 65 -1092 0 net=12023
rlabel metal2 1780 -1092 1780 -1092 0 net=13319
rlabel metal2 2 -1094 2 -1094 0 net=5060
rlabel metal2 828 -1094 828 -1094 0 net=6097
rlabel metal2 1248 -1094 1248 -1094 0 net=10045
rlabel metal2 1668 -1094 1668 -1094 0 net=13441
rlabel metal2 110 -1096 110 -1096 0 net=12457
rlabel metal2 933 -1098 933 -1098 0 net=7127
rlabel metal2 1024 -1098 1024 -1098 0 net=8213
rlabel metal2 1318 -1098 1318 -1098 0 net=9137
rlabel metal2 1402 -1098 1402 -1098 0 net=10019
rlabel metal2 572 -1100 572 -1100 0 net=8149
rlabel metal2 1080 -1100 1080 -1100 0 net=12869
rlabel metal2 789 -1102 789 -1102 0 net=8009
rlabel metal2 1486 -1102 1486 -1102 0 net=10339
rlabel metal2 814 -1104 814 -1104 0 net=6361
rlabel metal2 814 -1106 814 -1106 0 net=5981
rlabel metal2 1080 -1106 1080 -1106 0 net=5765
rlabel metal2 2 -1117 2 -1117 0 net=5145
rlabel metal2 86 -1117 86 -1117 0 net=2927
rlabel metal2 86 -1117 86 -1117 0 net=2927
rlabel metal2 128 -1117 128 -1117 0 net=8414
rlabel metal2 716 -1117 716 -1117 0 net=6502
rlabel metal2 933 -1117 933 -1117 0 net=8151
rlabel metal2 1153 -1117 1153 -1117 0 net=13064
rlabel metal2 1843 -1117 1843 -1117 0 net=12266
rlabel metal2 1878 -1117 1878 -1117 0 net=9533
rlabel metal2 1927 -1117 1927 -1117 0 net=6769
rlabel metal2 1927 -1117 1927 -1117 0 net=6769
rlabel metal2 1948 -1117 1948 -1117 0 net=11377
rlabel metal2 1976 -1117 1976 -1117 0 net=6693
rlabel metal2 16 -1119 16 -1119 0 net=2930
rlabel metal2 233 -1119 233 -1119 0 net=1814
rlabel metal2 656 -1119 656 -1119 0 net=5472
rlabel metal2 775 -1119 775 -1119 0 net=6928
rlabel metal2 880 -1119 880 -1119 0 net=6666
rlabel metal2 1549 -1119 1549 -1119 0 net=13129
rlabel metal2 1969 -1119 1969 -1119 0 net=10265
rlabel metal2 16 -1121 16 -1121 0 net=7373
rlabel metal2 135 -1121 135 -1121 0 net=7928
rlabel metal2 779 -1121 779 -1121 0 net=6200
rlabel metal2 866 -1121 866 -1121 0 net=8214
rlabel metal2 1045 -1121 1045 -1121 0 net=8164
rlabel metal2 1206 -1121 1206 -1121 0 net=8463
rlabel metal2 1206 -1121 1206 -1121 0 net=8463
rlabel metal2 1269 -1121 1269 -1121 0 net=8765
rlabel metal2 1269 -1121 1269 -1121 0 net=8765
rlabel metal2 1276 -1121 1276 -1121 0 net=8903
rlabel metal2 1276 -1121 1276 -1121 0 net=8903
rlabel metal2 1318 -1121 1318 -1121 0 net=8011
rlabel metal2 1962 -1121 1962 -1121 0 net=8711
rlabel metal2 23 -1123 23 -1123 0 net=4346
rlabel metal2 572 -1123 572 -1123 0 net=4564
rlabel metal2 674 -1123 674 -1123 0 net=4831
rlabel metal2 716 -1123 716 -1123 0 net=5767
rlabel metal2 1122 -1123 1122 -1123 0 net=8029
rlabel metal2 1122 -1123 1122 -1123 0 net=8029
rlabel metal2 1132 -1123 1132 -1123 0 net=11110
rlabel metal2 1584 -1123 1584 -1123 0 net=12409
rlabel metal2 30 -1125 30 -1125 0 net=1878
rlabel metal2 44 -1125 44 -1125 0 net=6807
rlabel metal2 957 -1125 957 -1125 0 net=12176
rlabel metal2 1759 -1125 1759 -1125 0 net=12927
rlabel metal2 30 -1127 30 -1127 0 net=1671
rlabel metal2 219 -1127 219 -1127 0 net=5033
rlabel metal2 562 -1127 562 -1127 0 net=7882
rlabel metal2 870 -1127 870 -1127 0 net=7244
rlabel metal2 1311 -1127 1311 -1127 0 net=9069
rlabel metal2 1367 -1127 1367 -1127 0 net=9915
rlabel metal2 1451 -1127 1451 -1127 0 net=11541
rlabel metal2 1591 -1127 1591 -1127 0 net=12231
rlabel metal2 1766 -1127 1766 -1127 0 net=12985
rlabel metal2 1766 -1127 1766 -1127 0 net=12985
rlabel metal2 1773 -1127 1773 -1127 0 net=13283
rlabel metal2 1773 -1127 1773 -1127 0 net=13283
rlabel metal2 1780 -1127 1780 -1127 0 net=13321
rlabel metal2 61 -1129 61 -1129 0 net=2904
rlabel metal2 282 -1129 282 -1129 0 net=1706
rlabel metal2 758 -1129 758 -1129 0 net=7439
rlabel metal2 1010 -1129 1010 -1129 0 net=7465
rlabel metal2 1045 -1129 1045 -1129 0 net=11422
rlabel metal2 1780 -1129 1780 -1129 0 net=13375
rlabel metal2 1808 -1129 1808 -1129 0 net=13621
rlabel metal2 1836 -1129 1836 -1129 0 net=13741
rlabel metal2 1871 -1129 1871 -1129 0 net=9497
rlabel metal2 65 -1131 65 -1131 0 net=4828
rlabel metal2 562 -1131 562 -1131 0 net=1423
rlabel metal2 1360 -1131 1360 -1131 0 net=9409
rlabel metal2 1500 -1131 1500 -1131 0 net=10937
rlabel metal2 1591 -1131 1591 -1131 0 net=11923
rlabel metal2 1689 -1131 1689 -1131 0 net=12571
rlabel metal2 1787 -1131 1787 -1131 0 net=13455
rlabel metal2 1822 -1131 1822 -1131 0 net=10876
rlabel metal2 65 -1133 65 -1133 0 net=4381
rlabel metal2 422 -1133 422 -1133 0 net=2356
rlabel metal2 464 -1133 464 -1133 0 net=1594
rlabel metal2 695 -1133 695 -1133 0 net=3899
rlabel metal2 730 -1133 730 -1133 0 net=4765
rlabel metal2 751 -1133 751 -1133 0 net=10305
rlabel metal2 1458 -1133 1458 -1133 0 net=10599
rlabel metal2 1542 -1133 1542 -1133 0 net=11535
rlabel metal2 72 -1135 72 -1135 0 net=8515
rlabel metal2 401 -1135 401 -1135 0 net=2541
rlabel metal2 401 -1135 401 -1135 0 net=2541
rlabel metal2 415 -1135 415 -1135 0 net=3255
rlabel metal2 625 -1135 625 -1135 0 net=4699
rlabel metal2 660 -1135 660 -1135 0 net=7129
rlabel metal2 996 -1135 996 -1135 0 net=7349
rlabel metal2 1017 -1135 1017 -1135 0 net=11126
rlabel metal2 1598 -1135 1598 -1135 0 net=11949
rlabel metal2 1682 -1135 1682 -1135 0 net=12553
rlabel metal2 100 -1137 100 -1137 0 net=4999
rlabel metal2 131 -1137 131 -1137 0 net=4851
rlabel metal2 695 -1137 695 -1137 0 net=5245
rlabel metal2 730 -1137 730 -1137 0 net=5867
rlabel metal2 782 -1137 782 -1137 0 net=8700
rlabel metal2 1423 -1137 1423 -1137 0 net=10197
rlabel metal2 1696 -1137 1696 -1137 0 net=12625
rlabel metal2 9 -1139 9 -1139 0 net=5903
rlabel metal2 114 -1139 114 -1139 0 net=5247
rlabel metal2 810 -1139 810 -1139 0 net=7258
rlabel metal2 1080 -1139 1080 -1139 0 net=7911
rlabel metal2 1139 -1139 1139 -1139 0 net=6064
rlabel metal2 1402 -1139 1402 -1139 0 net=10021
rlabel metal2 1458 -1139 1458 -1139 0 net=10341
rlabel metal2 1493 -1139 1493 -1139 0 net=10819
rlabel metal2 1563 -1139 1563 -1139 0 net=11853
rlabel metal2 1605 -1139 1605 -1139 0 net=12361
rlabel metal2 1724 -1139 1724 -1139 0 net=13763
rlabel metal2 9 -1141 9 -1141 0 net=3879
rlabel metal2 429 -1141 429 -1141 0 net=2366
rlabel metal2 859 -1141 859 -1141 0 net=8865
rlabel metal2 1381 -1141 1381 -1141 0 net=9745
rlabel metal2 1444 -1141 1444 -1141 0 net=10517
rlabel metal2 1521 -1141 1521 -1141 0 net=11425
rlabel metal2 1794 -1141 1794 -1141 0 net=13443
rlabel metal2 79 -1143 79 -1143 0 net=11233
rlabel metal2 1605 -1143 1605 -1143 0 net=12039
rlabel metal2 1668 -1143 1668 -1143 0 net=12459
rlabel metal2 1752 -1143 1752 -1143 0 net=12871
rlabel metal2 121 -1145 121 -1145 0 net=1643
rlabel metal2 159 -1145 159 -1145 0 net=3799
rlabel metal2 331 -1145 331 -1145 0 net=2595
rlabel metal2 555 -1145 555 -1145 0 net=4515
rlabel metal2 723 -1145 723 -1145 0 net=5065
rlabel metal2 761 -1145 761 -1145 0 net=7073
rlabel metal2 1444 -1145 1444 -1145 0 net=11307
rlabel metal2 1486 -1145 1486 -1145 0 net=11619
rlabel metal2 1612 -1145 1612 -1145 0 net=12051
rlabel metal2 1668 -1145 1668 -1145 0 net=13653
rlabel metal2 121 -1147 121 -1147 0 net=331
rlabel metal2 814 -1147 814 -1147 0 net=5983
rlabel metal2 863 -1147 863 -1147 0 net=9373
rlabel metal2 1437 -1147 1437 -1147 0 net=10461
rlabel metal2 1507 -1147 1507 -1147 0 net=11001
rlabel metal2 1626 -1147 1626 -1147 0 net=12153
rlabel metal2 1745 -1147 1745 -1147 0 net=10327
rlabel metal2 180 -1149 180 -1149 0 net=1006
rlabel metal2 863 -1149 863 -1149 0 net=6547
rlabel metal2 894 -1149 894 -1149 0 net=11828
rlabel metal2 1717 -1149 1717 -1149 0 net=12841
rlabel metal2 184 -1151 184 -1151 0 net=1689
rlabel metal2 184 -1151 184 -1151 0 net=1689
rlabel metal2 198 -1151 198 -1151 0 net=1817
rlabel metal2 359 -1151 359 -1151 0 net=2336
rlabel metal2 670 -1151 670 -1151 0 net=10607
rlabel metal2 1514 -1151 1514 -1151 0 net=11345
rlabel metal2 1647 -1151 1647 -1151 0 net=12469
rlabel metal2 1717 -1151 1717 -1151 0 net=12789
rlabel metal2 82 -1153 82 -1153 0 net=3527
rlabel metal2 359 -1153 359 -1153 0 net=1963
rlabel metal2 422 -1153 422 -1153 0 net=2456
rlabel metal2 1136 -1153 1136 -1153 0 net=12027
rlabel metal2 1710 -1153 1710 -1153 0 net=12665
rlabel metal2 233 -1155 233 -1155 0 net=3021
rlabel metal2 261 -1155 261 -1155 0 net=1664
rlabel metal2 303 -1155 303 -1155 0 net=1933
rlabel metal2 366 -1155 366 -1155 0 net=2295
rlabel metal2 373 -1155 373 -1155 0 net=2129
rlabel metal2 436 -1155 436 -1155 0 net=4592
rlabel metal2 555 -1155 555 -1155 0 net=4989
rlabel metal2 684 -1155 684 -1155 0 net=13497
rlabel metal2 51 -1157 51 -1157 0 net=2937
rlabel metal2 380 -1157 380 -1157 0 net=4911
rlabel metal2 873 -1157 873 -1157 0 net=11667
rlabel metal2 1633 -1157 1633 -1157 0 net=12271
rlabel metal2 51 -1159 51 -1159 0 net=2055
rlabel metal2 779 -1159 779 -1159 0 net=10297
rlabel metal2 1465 -1159 1465 -1159 0 net=10735
rlabel metal2 1521 -1159 1521 -1159 0 net=12215
rlabel metal2 240 -1161 240 -1161 0 net=2571
rlabel metal2 268 -1161 268 -1161 0 net=2231
rlabel metal2 282 -1161 282 -1161 0 net=1767
rlabel metal2 366 -1161 366 -1161 0 net=2375
rlabel metal2 436 -1161 436 -1161 0 net=6647
rlabel metal2 926 -1161 926 -1161 0 net=9353
rlabel metal2 1472 -1161 1472 -1161 0 net=10761
rlabel metal2 163 -1163 163 -1163 0 net=4637
rlabel metal2 352 -1163 352 -1163 0 net=3322
rlabel metal2 975 -1163 975 -1163 0 net=7021
rlabel metal2 989 -1163 989 -1163 0 net=7193
rlabel metal2 1003 -1163 1003 -1163 0 net=8499
rlabel metal2 1248 -1163 1248 -1163 0 net=10047
rlabel metal2 1535 -1163 1535 -1163 0 net=11527
rlabel metal2 58 -1165 58 -1165 0 net=3441
rlabel metal2 446 -1165 446 -1165 0 net=12375
rlabel metal2 163 -1167 163 -1167 0 net=2725
rlabel metal2 464 -1167 464 -1167 0 net=4737
rlabel metal2 583 -1167 583 -1167 0 net=5479
rlabel metal2 912 -1167 912 -1167 0 net=6201
rlabel metal2 1160 -1167 1160 -1167 0 net=8165
rlabel metal2 142 -1169 142 -1169 0 net=6337
rlabel metal2 583 -1169 583 -1169 0 net=7675
rlabel metal2 1038 -1169 1038 -1169 0 net=7433
rlabel metal2 1241 -1169 1241 -1169 0 net=8801
rlabel metal2 142 -1171 142 -1171 0 net=1519
rlabel metal2 240 -1171 240 -1171 0 net=1901
rlabel metal2 303 -1171 303 -1171 0 net=1879
rlabel metal2 961 -1171 961 -1171 0 net=7047
rlabel metal2 1017 -1171 1017 -1171 0 net=10443
rlabel metal2 254 -1173 254 -1173 0 net=1833
rlabel metal2 313 -1173 313 -1173 0 net=8141
rlabel metal2 1164 -1173 1164 -1173 0 net=8431
rlabel metal2 1234 -1173 1234 -1173 0 net=8731
rlabel metal2 212 -1175 212 -1175 0 net=6701
rlabel metal2 275 -1175 275 -1175 0 net=1723
rlabel metal2 450 -1175 450 -1175 0 net=12443
rlabel metal2 37 -1177 37 -1177 0 net=3452
rlabel metal2 453 -1177 453 -1177 0 net=11027
rlabel metal2 1213 -1177 1213 -1177 0 net=8835
rlabel metal2 289 -1179 289 -1179 0 net=1716
rlabel metal2 590 -1179 590 -1179 0 net=5657
rlabel metal2 849 -1179 849 -1179 0 net=8441
rlabel metal2 1048 -1179 1048 -1179 0 net=12419
rlabel metal2 107 -1181 107 -1181 0 net=2460
rlabel metal2 1087 -1181 1087 -1181 0 net=7889
rlabel metal2 107 -1183 107 -1183 0 net=5299
rlabel metal2 982 -1183 982 -1183 0 net=7645
rlabel metal2 1059 -1183 1059 -1183 0 net=7967
rlabel metal2 1094 -1183 1094 -1183 0 net=7561
rlabel metal2 1115 -1183 1115 -1183 0 net=8189
rlabel metal2 156 -1185 156 -1185 0 net=3751
rlabel metal2 632 -1185 632 -1185 0 net=10791
rlabel metal2 324 -1187 324 -1187 0 net=4535
rlabel metal2 667 -1187 667 -1187 0 net=8140
rlabel metal2 324 -1189 324 -1189 0 net=2793
rlabel metal2 516 -1189 516 -1189 0 net=9649
rlabel metal2 338 -1191 338 -1191 0 net=6323
rlabel metal2 709 -1191 709 -1191 0 net=7761
rlabel metal2 821 -1191 821 -1191 0 net=6023
rlabel metal2 877 -1191 877 -1191 0 net=8807
rlabel metal2 1108 -1191 1108 -1191 0 net=7989
rlabel metal2 1157 -1191 1157 -1191 0 net=8669
rlabel metal2 37 -1193 37 -1193 0 net=6245
rlabel metal2 709 -1193 709 -1193 0 net=4187
rlabel metal2 891 -1193 891 -1193 0 net=6353
rlabel metal2 1052 -1193 1052 -1193 0 net=7797
rlabel metal2 1108 -1193 1108 -1193 0 net=8927
rlabel metal2 408 -1195 408 -1195 0 net=4119
rlabel metal2 408 -1197 408 -1197 0 net=2199
rlabel metal2 733 -1197 733 -1197 0 net=13370
rlabel metal2 443 -1199 443 -1199 0 net=7951
rlabel metal2 1157 -1199 1157 -1199 0 net=9542
rlabel metal2 212 -1201 212 -1201 0 net=3069
rlabel metal2 457 -1201 457 -1201 0 net=2995
rlabel metal2 576 -1201 576 -1201 0 net=4221
rlabel metal2 737 -1201 737 -1201 0 net=6672
rlabel metal2 1181 -1201 1181 -1201 0 net=12709
rlabel metal2 44 -1203 44 -1203 0 net=5199
rlabel metal2 1185 -1203 1185 -1203 0 net=10785
rlabel metal2 289 -1205 289 -1205 0 net=4473
rlabel metal2 744 -1205 744 -1205 0 net=5443
rlabel metal2 898 -1205 898 -1205 0 net=6417
rlabel metal2 1066 -1205 1066 -1205 0 net=7853
rlabel metal2 1143 -1205 1143 -1205 0 net=8295
rlabel metal2 1395 -1205 1395 -1205 0 net=9987
rlabel metal2 471 -1207 471 -1207 0 net=4311
rlabel metal2 611 -1207 611 -1207 0 net=4903
rlabel metal2 747 -1207 747 -1207 0 net=1
rlabel metal2 807 -1207 807 -1207 0 net=337
rlabel metal2 1143 -1207 1143 -1207 0 net=8935
rlabel metal2 1374 -1207 1374 -1207 0 net=9583
rlabel metal2 429 -1209 429 -1209 0 net=5385
rlabel metal2 474 -1209 474 -1209 0 net=3642
rlabel metal2 506 -1209 506 -1209 0 net=2001
rlabel metal2 905 -1209 905 -1209 0 net=13536
rlabel metal2 124 -1211 124 -1211 0 net=3485
rlabel metal2 513 -1211 513 -1211 0 net=5195
rlabel metal2 940 -1211 940 -1211 0 net=7041
rlabel metal2 1255 -1211 1255 -1211 0 net=9241
rlabel metal2 1353 -1211 1353 -1211 0 net=9359
rlabel metal2 1619 -1211 1619 -1211 0 net=12025
rlabel metal2 82 -1213 82 -1213 0 net=8285
rlabel metal2 478 -1215 478 -1215 0 net=5531
rlabel metal2 940 -1215 940 -1215 0 net=3907
rlabel metal2 1325 -1215 1325 -1215 0 net=9139
rlabel metal2 1346 -1215 1346 -1215 0 net=9287
rlabel metal2 177 -1217 177 -1217 0 net=3789
rlabel metal2 485 -1217 485 -1217 0 net=3411
rlabel metal2 579 -1217 579 -1217 0 net=4471
rlabel metal2 947 -1217 947 -1217 0 net=6991
rlabel metal2 1297 -1217 1297 -1217 0 net=8951
rlabel metal2 1332 -1217 1332 -1217 0 net=9181
rlabel metal2 177 -1219 177 -1219 0 net=6362
rlabel metal2 1297 -1219 1297 -1219 0 net=9029
rlabel metal2 520 -1221 520 -1221 0 net=8215
rlabel metal2 1304 -1221 1304 -1221 0 net=10221
rlabel metal2 93 -1223 93 -1223 0 net=3569
rlabel metal2 548 -1223 548 -1223 0 net=7071
rlabel metal2 1416 -1223 1416 -1223 0 net=10095
rlabel metal2 47 -1225 47 -1225 0 net=10001
rlabel metal2 93 -1227 93 -1227 0 net=2219
rlabel metal2 569 -1227 569 -1227 0 net=9097
rlabel metal2 149 -1229 149 -1229 0 net=2087
rlabel metal2 492 -1229 492 -1229 0 net=7499
rlabel metal2 597 -1229 597 -1229 0 net=4571
rlabel metal2 828 -1229 828 -1229 0 net=6099
rlabel metal2 58 -1231 58 -1231 0 net=4333
rlabel metal2 828 -1231 828 -1231 0 net=8111
rlabel metal2 919 -1231 919 -1231 0 net=6963
rlabel metal2 191 -1233 191 -1233 0 net=2869
rlabel metal2 492 -1233 492 -1233 0 net=3543
rlabel metal2 170 -1235 170 -1235 0 net=2263
rlabel metal2 646 -1235 646 -1235 0 net=6633
rlabel metal2 170 -1237 170 -1237 0 net=5573
rlabel metal2 835 -1237 835 -1237 0 net=6427
rlabel metal2 793 -1239 793 -1239 0 net=5599
rlabel metal2 226 -1241 226 -1241 0 net=7166
rlabel metal2 16 -1252 16 -1252 0 net=7375
rlabel metal2 16 -1252 16 -1252 0 net=7375
rlabel metal2 23 -1252 23 -1252 0 net=2221
rlabel metal2 107 -1252 107 -1252 0 net=5300
rlabel metal2 163 -1252 163 -1252 0 net=2726
rlabel metal2 247 -1252 247 -1252 0 net=2572
rlabel metal2 282 -1252 282 -1252 0 net=1768
rlabel metal2 457 -1252 457 -1252 0 net=2996
rlabel metal2 688 -1252 688 -1252 0 net=4904
rlabel metal2 793 -1252 793 -1252 0 net=352
rlabel metal2 1101 -1252 1101 -1252 0 net=7563
rlabel metal2 1101 -1252 1101 -1252 0 net=7563
rlabel metal2 1111 -1252 1111 -1252 0 net=12928
rlabel metal2 1906 -1252 1906 -1252 0 net=8013
rlabel metal2 1962 -1252 1962 -1252 0 net=9499
rlabel metal2 30 -1254 30 -1254 0 net=1672
rlabel metal2 457 -1254 457 -1254 0 net=4335
rlabel metal2 628 -1254 628 -1254 0 net=5480
rlabel metal2 821 -1254 821 -1254 0 net=7854
rlabel metal2 1129 -1254 1129 -1254 0 net=12554
rlabel metal2 1843 -1254 1843 -1254 0 net=13743
rlabel metal2 1913 -1254 1913 -1254 0 net=8167
rlabel metal2 1969 -1254 1969 -1254 0 net=8713
rlabel metal2 1969 -1254 1969 -1254 0 net=8713
rlabel metal2 1976 -1254 1976 -1254 0 net=10267
rlabel metal2 1990 -1254 1990 -1254 0 net=6695
rlabel metal2 1990 -1254 1990 -1254 0 net=6695
rlabel metal2 30 -1256 30 -1256 0 net=3747
rlabel metal2 226 -1256 226 -1256 0 net=3323
rlabel metal2 541 -1256 541 -1256 0 net=6339
rlabel metal2 604 -1256 604 -1256 0 net=6247
rlabel metal2 838 -1256 838 -1256 0 net=10048
rlabel metal2 1675 -1256 1675 -1256 0 net=12029
rlabel metal2 1920 -1256 1920 -1256 0 net=9535
rlabel metal2 1955 -1256 1955 -1256 0 net=11379
rlabel metal2 37 -1258 37 -1258 0 net=5201
rlabel metal2 58 -1258 58 -1258 0 net=6563
rlabel metal2 856 -1258 856 -1258 0 net=12232
rlabel metal2 1927 -1258 1927 -1258 0 net=6771
rlabel metal2 1927 -1258 1927 -1258 0 net=6771
rlabel metal2 40 -1260 40 -1260 0 net=10762
rlabel metal2 1689 -1260 1689 -1260 0 net=12363
rlabel metal2 1689 -1260 1689 -1260 0 net=12363
rlabel metal2 1759 -1260 1759 -1260 0 net=12563
rlabel metal2 44 -1262 44 -1262 0 net=4223
rlabel metal2 586 -1262 586 -1262 0 net=6024
rlabel metal2 856 -1262 856 -1262 0 net=200
rlabel metal2 908 -1262 908 -1262 0 net=7434
rlabel metal2 1269 -1262 1269 -1262 0 net=8767
rlabel metal2 1290 -1262 1290 -1262 0 net=7075
rlabel metal2 58 -1264 58 -1264 0 net=12026
rlabel metal2 61 -1266 61 -1266 0 net=12216
rlabel metal2 1612 -1266 1612 -1266 0 net=12053
rlabel metal2 1787 -1266 1787 -1266 0 net=13457
rlabel metal2 65 -1268 65 -1268 0 net=4383
rlabel metal2 289 -1268 289 -1268 0 net=2543
rlabel metal2 415 -1268 415 -1268 0 net=3257
rlabel metal2 562 -1268 562 -1268 0 net=7042
rlabel metal2 1129 -1268 1129 -1268 0 net=8143
rlabel metal2 1150 -1268 1150 -1268 0 net=8153
rlabel metal2 1150 -1268 1150 -1268 0 net=8153
rlabel metal2 1178 -1268 1178 -1268 0 net=12410
rlabel metal2 51 -1270 51 -1270 0 net=2057
rlabel metal2 79 -1270 79 -1270 0 net=6324
rlabel metal2 352 -1270 352 -1270 0 net=3442
rlabel metal2 688 -1270 688 -1270 0 net=5067
rlabel metal2 730 -1270 730 -1270 0 net=5869
rlabel metal2 730 -1270 730 -1270 0 net=5869
rlabel metal2 775 -1270 775 -1270 0 net=12710
rlabel metal2 9 -1272 9 -1272 0 net=3881
rlabel metal2 82 -1272 82 -1272 0 net=4391
rlabel metal2 646 -1272 646 -1272 0 net=5574
rlabel metal2 1171 -1272 1171 -1272 0 net=8217
rlabel metal2 1220 -1272 1220 -1272 0 net=8837
rlabel metal2 1269 -1272 1269 -1272 0 net=8905
rlabel metal2 1290 -1272 1290 -1272 0 net=9031
rlabel metal2 1388 -1272 1388 -1272 0 net=9411
rlabel metal2 1430 -1272 1430 -1272 0 net=10097
rlabel metal2 1430 -1272 1430 -1272 0 net=10097
rlabel metal2 1458 -1272 1458 -1272 0 net=10343
rlabel metal2 1542 -1272 1542 -1272 0 net=10821
rlabel metal2 1626 -1272 1626 -1272 0 net=12155
rlabel metal2 1787 -1272 1787 -1272 0 net=13087
rlabel metal2 9 -1274 9 -1274 0 net=7763
rlabel metal2 824 -1274 824 -1274 0 net=6683
rlabel metal2 870 -1274 870 -1274 0 net=6203
rlabel metal2 922 -1274 922 -1274 0 net=13130
rlabel metal2 2 -1276 2 -1276 0 net=5147
rlabel metal2 912 -1276 912 -1276 0 net=8929
rlabel metal2 1122 -1276 1122 -1276 0 net=8031
rlabel metal2 1171 -1276 1171 -1276 0 net=10711
rlabel metal2 1808 -1276 1808 -1276 0 net=13445
rlabel metal2 86 -1278 86 -1278 0 net=2928
rlabel metal2 177 -1278 177 -1278 0 net=4472
rlabel metal2 681 -1278 681 -1278 0 net=4853
rlabel metal2 779 -1278 779 -1278 0 net=3365
rlabel metal2 1073 -1278 1073 -1278 0 net=11528
rlabel metal2 1829 -1278 1829 -1278 0 net=13623
rlabel metal2 54 -1280 54 -1280 0 net=3415
rlabel metal2 93 -1280 93 -1280 0 net=1521
rlabel metal2 149 -1280 149 -1280 0 net=2089
rlabel metal2 247 -1280 247 -1280 0 net=7953
rlabel metal2 1234 -1280 1234 -1280 0 net=8867
rlabel metal2 1297 -1280 1297 -1280 0 net=9099
rlabel metal2 1388 -1280 1388 -1280 0 net=9989
rlabel metal2 1437 -1280 1437 -1280 0 net=10299
rlabel metal2 1486 -1280 1486 -1280 0 net=11621
rlabel metal2 1773 -1280 1773 -1280 0 net=13285
rlabel metal2 107 -1282 107 -1282 0 net=7072
rlabel metal2 611 -1282 611 -1282 0 net=4475
rlabel metal2 653 -1282 653 -1282 0 net=4701
rlabel metal2 877 -1282 877 -1282 0 net=10855
rlabel metal2 1143 -1282 1143 -1282 0 net=8937
rlabel metal2 1416 -1282 1416 -1282 0 net=10003
rlabel metal2 1479 -1282 1479 -1282 0 net=10463
rlabel metal2 1493 -1282 1493 -1282 0 net=10519
rlabel metal2 1591 -1282 1591 -1282 0 net=11925
rlabel metal2 1745 -1282 1745 -1282 0 net=12843
rlabel metal2 110 -1284 110 -1284 0 net=13255
rlabel metal2 121 -1286 121 -1286 0 net=5415
rlabel metal2 254 -1286 254 -1286 0 net=6702
rlabel metal2 618 -1286 618 -1286 0 net=6355
rlabel metal2 926 -1286 926 -1286 0 net=13575
rlabel metal2 135 -1288 135 -1288 0 net=1645
rlabel metal2 135 -1288 135 -1288 0 net=1645
rlabel metal2 152 -1288 152 -1288 0 net=6475
rlabel metal2 296 -1288 296 -1288 0 net=1835
rlabel metal2 317 -1288 317 -1288 0 net=3529
rlabel metal2 548 -1288 548 -1288 0 net=3909
rlabel metal2 964 -1288 964 -1288 0 net=10198
rlabel metal2 156 -1290 156 -1290 0 net=13711
rlabel metal2 156 -1292 156 -1292 0 net=7131
rlabel metal2 712 -1292 712 -1292 0 net=11481
rlabel metal2 128 -1294 128 -1294 0 net=5001
rlabel metal2 877 -1294 877 -1294 0 net=7467
rlabel metal2 1038 -1294 1038 -1294 0 net=8443
rlabel metal2 1244 -1294 1244 -1294 0 net=12631
rlabel metal2 1563 -1294 1563 -1294 0 net=11235
rlabel metal2 1605 -1294 1605 -1294 0 net=12041
rlabel metal2 75 -1296 75 -1296 0 net=13135
rlabel metal2 1045 -1296 1045 -1296 0 net=7969
rlabel metal2 1094 -1296 1094 -1296 0 net=7991
rlabel metal2 1143 -1296 1143 -1296 0 net=8297
rlabel metal2 1255 -1296 1255 -1296 0 net=9243
rlabel metal2 1416 -1296 1416 -1296 0 net=10023
rlabel metal2 1465 -1296 1465 -1296 0 net=10445
rlabel metal2 124 -1298 124 -1298 0 net=10641
rlabel metal2 1185 -1298 1185 -1298 0 net=12626
rlabel metal2 128 -1300 128 -1300 0 net=5984
rlabel metal2 891 -1300 891 -1300 0 net=6965
rlabel metal2 961 -1300 961 -1300 0 net=7321
rlabel metal2 1055 -1300 1055 -1300 0 net=12585
rlabel metal2 163 -1302 163 -1302 0 net=1902
rlabel metal2 254 -1302 254 -1302 0 net=1611
rlabel metal2 842 -1302 842 -1302 0 net=6419
rlabel metal2 929 -1302 929 -1302 0 net=11503
rlabel metal2 1780 -1302 1780 -1302 0 net=13377
rlabel metal2 170 -1304 170 -1304 0 net=4913
rlabel metal2 394 -1304 394 -1304 0 net=2130
rlabel metal2 443 -1304 443 -1304 0 net=7890
rlabel metal2 1423 -1304 1423 -1304 0 net=10609
rlabel metal2 1766 -1304 1766 -1304 0 net=12987
rlabel metal2 205 -1306 205 -1306 0 net=2871
rlabel metal2 268 -1306 268 -1306 0 net=2233
rlabel metal2 401 -1306 401 -1306 0 net=4991
rlabel metal2 807 -1306 807 -1306 0 net=7079
rlabel metal2 929 -1306 929 -1306 0 net=10891
rlabel metal2 1752 -1306 1752 -1306 0 net=10329
rlabel metal2 184 -1308 184 -1308 0 net=1690
rlabel metal2 233 -1308 233 -1308 0 net=3023
rlabel metal2 296 -1308 296 -1308 0 net=1935
rlabel metal2 338 -1308 338 -1308 0 net=2201
rlabel metal2 422 -1308 422 -1308 0 net=12444
rlabel metal2 184 -1310 184 -1310 0 net=1881
rlabel metal2 310 -1310 310 -1310 0 net=3801
rlabel metal2 807 -1310 807 -1310 0 net=7913
rlabel metal2 1108 -1310 1108 -1310 0 net=10577
rlabel metal2 1696 -1310 1696 -1310 0 net=11427
rlabel metal2 100 -1312 100 -1312 0 net=5905
rlabel metal2 317 -1312 317 -1312 0 net=2297
rlabel metal2 408 -1312 408 -1312 0 net=3571
rlabel metal2 534 -1312 534 -1312 0 net=2597
rlabel metal2 810 -1312 810 -1312 0 net=13159
rlabel metal2 72 -1314 72 -1314 0 net=8517
rlabel metal2 422 -1314 422 -1314 0 net=3677
rlabel metal2 947 -1314 947 -1314 0 net=6993
rlabel metal2 961 -1314 961 -1314 0 net=7049
rlabel metal2 1017 -1314 1017 -1314 0 net=11536
rlabel metal2 51 -1316 51 -1316 0 net=910
rlabel metal2 954 -1316 954 -1316 0 net=7023
rlabel metal2 989 -1316 989 -1316 0 net=7677
rlabel metal2 1066 -1316 1066 -1316 0 net=8749
rlabel metal2 1391 -1316 1391 -1316 0 net=1
rlabel metal2 1451 -1316 1451 -1316 0 net=10307
rlabel metal2 1668 -1316 1668 -1316 0 net=13655
rlabel metal2 72 -1318 72 -1318 0 net=7500
rlabel metal2 968 -1318 968 -1318 0 net=6101
rlabel metal2 1255 -1318 1255 -1318 0 net=9361
rlabel metal2 1598 -1318 1598 -1318 0 net=11951
rlabel metal2 1696 -1318 1696 -1318 0 net=12377
rlabel metal2 100 -1320 100 -1320 0 net=2101
rlabel metal2 352 -1320 352 -1320 0 net=1965
rlabel metal2 366 -1320 366 -1320 0 net=2377
rlabel metal2 443 -1320 443 -1320 0 net=3939
rlabel metal2 968 -1320 968 -1320 0 net=815
rlabel metal2 1031 -1320 1031 -1320 0 net=8952
rlabel metal2 1360 -1320 1360 -1320 0 net=9355
rlabel metal2 142 -1322 142 -1322 0 net=2781
rlabel metal2 324 -1322 324 -1322 0 net=2795
rlabel metal2 366 -1322 366 -1322 0 net=6773
rlabel metal2 534 -1322 534 -1322 0 net=4767
rlabel metal2 772 -1322 772 -1322 0 net=5659
rlabel metal2 975 -1322 975 -1322 0 net=7647
rlabel metal2 996 -1322 996 -1322 0 net=7195
rlabel metal2 1080 -1322 1080 -1322 0 net=8191
rlabel metal2 1304 -1322 1304 -1322 0 net=10223
rlabel metal2 1374 -1322 1374 -1322 0 net=9585
rlabel metal2 1444 -1322 1444 -1322 0 net=11309
rlabel metal2 233 -1324 233 -1324 0 net=3545
rlabel metal2 530 -1324 530 -1324 0 net=9111
rlabel metal2 275 -1326 275 -1326 0 net=1725
rlabel metal2 373 -1326 373 -1326 0 net=2939
rlabel metal2 450 -1326 450 -1326 0 net=6823
rlabel metal2 859 -1326 859 -1326 0 net=8883
rlabel metal2 1325 -1326 1325 -1326 0 net=9141
rlabel metal2 212 -1328 212 -1328 0 net=3071
rlabel metal2 373 -1328 373 -1328 0 net=3305
rlabel metal2 765 -1328 765 -1328 0 net=5601
rlabel metal2 859 -1328 859 -1328 0 net=12399
rlabel metal2 198 -1330 198 -1330 0 net=1819
rlabel metal2 436 -1330 436 -1330 0 net=6649
rlabel metal2 464 -1330 464 -1330 0 net=4739
rlabel metal2 905 -1330 905 -1330 0 net=7669
rlabel metal2 996 -1330 996 -1330 0 net=13322
rlabel metal2 198 -1332 198 -1332 0 net=4573
rlabel metal2 884 -1332 884 -1332 0 net=6429
rlabel metal2 1164 -1332 1164 -1332 0 net=8671
rlabel metal2 1227 -1332 1227 -1332 0 net=9651
rlabel metal2 1864 -1332 1864 -1332 0 net=13765
rlabel metal2 436 -1334 436 -1334 0 net=7441
rlabel metal2 884 -1334 884 -1334 0 net=6635
rlabel metal2 1059 -1334 1059 -1334 0 net=8809
rlabel metal2 1227 -1334 1227 -1334 0 net=8803
rlabel metal2 1318 -1334 1318 -1334 0 net=9071
rlabel metal2 1815 -1334 1815 -1334 0 net=13499
rlabel metal2 464 -1336 464 -1336 0 net=5769
rlabel metal2 751 -1336 751 -1336 0 net=5533
rlabel metal2 1052 -1336 1052 -1336 0 net=7799
rlabel metal2 1248 -1336 1248 -1336 0 net=9183
rlabel metal2 1794 -1336 1794 -1336 0 net=12873
rlabel metal2 471 -1338 471 -1338 0 net=8501
rlabel metal2 1318 -1338 1318 -1338 0 net=9747
rlabel metal2 1647 -1338 1647 -1338 0 net=12471
rlabel metal2 474 -1340 474 -1340 0 net=4516
rlabel metal2 639 -1340 639 -1340 0 net=4833
rlabel metal2 716 -1340 716 -1340 0 net=5197
rlabel metal2 744 -1340 744 -1340 0 net=5445
rlabel metal2 1003 -1340 1003 -1340 0 net=7277
rlabel metal2 1346 -1340 1346 -1340 0 net=9289
rlabel metal2 1647 -1340 1647 -1340 0 net=12667
rlabel metal2 114 -1342 114 -1342 0 net=5248
rlabel metal2 737 -1342 737 -1342 0 net=7351
rlabel metal2 1052 -1342 1052 -1342 0 net=9855
rlabel metal2 1717 -1342 1717 -1342 0 net=12791
rlabel metal2 114 -1344 114 -1344 0 net=4639
rlabel metal2 478 -1344 478 -1344 0 net=3791
rlabel metal2 569 -1344 569 -1344 0 net=4189
rlabel metal2 943 -1344 943 -1344 0 net=12743
rlabel metal2 159 -1346 159 -1346 0 net=2973
rlabel metal2 478 -1346 478 -1346 0 net=3487
rlabel metal2 590 -1346 590 -1346 0 net=3752
rlabel metal2 1353 -1346 1353 -1346 0 net=9917
rlabel metal2 173 -1348 173 -1348 0 net=7711
rlabel metal2 1367 -1348 1367 -1348 0 net=9375
rlabel metal2 485 -1350 485 -1350 0 net=3412
rlabel metal2 625 -1350 625 -1350 0 net=5246
rlabel metal2 709 -1350 709 -1350 0 net=6141
rlabel metal2 1241 -1350 1241 -1350 0 net=8733
rlabel metal2 219 -1352 219 -1352 0 net=5035
rlabel metal2 1241 -1352 1241 -1352 0 net=11346
rlabel metal2 191 -1354 191 -1354 0 net=2265
rlabel metal2 432 -1354 432 -1354 0 net=7407
rlabel metal2 1556 -1354 1556 -1354 0 net=11003
rlabel metal2 191 -1356 191 -1356 0 net=3965
rlabel metal2 1535 -1356 1535 -1356 0 net=10793
rlabel metal2 485 -1358 485 -1358 0 net=3901
rlabel metal2 1528 -1358 1528 -1358 0 net=10787
rlabel metal2 429 -1360 429 -1360 0 net=5387
rlabel metal2 1514 -1360 1514 -1360 0 net=10737
rlabel metal2 429 -1362 429 -1362 0 net=8286
rlabel metal2 492 -1364 492 -1364 0 net=2003
rlabel metal2 527 -1364 527 -1364 0 net=4313
rlabel metal2 1500 -1364 1500 -1364 0 net=10601
rlabel metal2 1570 -1364 1570 -1364 0 net=11543
rlabel metal2 499 -1366 499 -1366 0 net=6809
rlabel metal2 1500 -1366 1500 -1366 0 net=12273
rlabel metal2 506 -1368 506 -1368 0 net=4537
rlabel metal2 933 -1368 933 -1368 0 net=6705
rlabel metal2 1549 -1368 1549 -1368 0 net=10939
rlabel metal2 1577 -1368 1577 -1368 0 net=11855
rlabel metal2 527 -1370 527 -1370 0 net=4120
rlabel metal2 1549 -1370 1549 -1370 0 net=12573
rlabel metal2 632 -1372 632 -1372 0 net=8113
rlabel metal2 919 -1372 919 -1372 0 net=8391
rlabel metal2 1724 -1372 1724 -1372 0 net=12461
rlabel metal2 744 -1374 744 -1374 0 net=5507
rlabel metal2 1710 -1374 1710 -1374 0 net=12421
rlabel metal2 828 -1376 828 -1376 0 net=6549
rlabel metal2 1584 -1376 1584 -1376 0 net=11669
rlabel metal2 653 -1378 653 -1378 0 net=7133
rlabel metal2 1199 -1378 1199 -1378 0 net=11029
rlabel metal2 1192 -1380 1192 -1380 0 net=8433
rlabel metal2 1192 -1382 1192 -1382 0 net=8465
rlabel metal2 180 -1384 180 -1384 0 net=8439
rlabel metal2 2 -1395 2 -1395 0 net=2051
rlabel metal2 485 -1395 485 -1395 0 net=3902
rlabel metal2 940 -1395 940 -1395 0 net=12668
rlabel metal2 1766 -1395 1766 -1395 0 net=10331
rlabel metal2 1766 -1395 1766 -1395 0 net=10331
rlabel metal2 1892 -1395 1892 -1395 0 net=13713
rlabel metal2 1892 -1395 1892 -1395 0 net=13713
rlabel metal2 1899 -1395 1899 -1395 0 net=13767
rlabel metal2 1969 -1395 1969 -1395 0 net=8714
rlabel metal2 1969 -1395 1969 -1395 0 net=8714
rlabel metal2 1976 -1395 1976 -1395 0 net=11381
rlabel metal2 9 -1397 9 -1397 0 net=7764
rlabel metal2 485 -1397 485 -1397 0 net=2005
rlabel metal2 527 -1397 527 -1397 0 net=4740
rlabel metal2 674 -1397 674 -1397 0 net=4703
rlabel metal2 712 -1397 712 -1397 0 net=8930
rlabel metal2 947 -1397 947 -1397 0 net=6994
rlabel metal2 1003 -1397 1003 -1397 0 net=7279
rlabel metal2 1038 -1397 1038 -1397 0 net=7323
rlabel metal2 1104 -1397 1104 -1397 0 net=10520
rlabel metal2 1647 -1397 1647 -1397 0 net=13257
rlabel metal2 1913 -1397 1913 -1397 0 net=6772
rlabel metal2 1941 -1397 1941 -1397 0 net=8169
rlabel metal2 9 -1399 9 -1399 0 net=6477
rlabel metal2 527 -1399 527 -1399 0 net=3007
rlabel metal2 926 -1399 926 -1399 0 net=7747
rlabel metal2 1052 -1399 1052 -1399 0 net=12586
rlabel metal2 1822 -1399 1822 -1399 0 net=7077
rlabel metal2 1948 -1399 1948 -1399 0 net=8015
rlabel metal2 1983 -1399 1983 -1399 0 net=10269
rlabel metal2 1997 -1399 1997 -1399 0 net=9501
rlabel metal2 16 -1401 16 -1401 0 net=7376
rlabel metal2 184 -1401 184 -1401 0 net=1882
rlabel metal2 1241 -1401 1241 -1401 0 net=12472
rlabel metal2 1843 -1401 1843 -1401 0 net=12031
rlabel metal2 1983 -1401 1983 -1401 0 net=6697
rlabel metal2 16 -1403 16 -1403 0 net=5417
rlabel metal2 142 -1403 142 -1403 0 net=11482
rlabel metal2 1780 -1403 1780 -1403 0 net=12989
rlabel metal2 1864 -1403 1864 -1403 0 net=13501
rlabel metal2 23 -1405 23 -1405 0 net=2223
rlabel metal2 23 -1405 23 -1405 0 net=2223
rlabel metal2 30 -1405 30 -1405 0 net=3748
rlabel metal2 968 -1405 968 -1405 0 net=9112
rlabel metal2 1577 -1405 1577 -1405 0 net=8393
rlabel metal2 1864 -1405 1864 -1405 0 net=13577
rlabel metal2 1916 -1405 1916 -1405 0 net=9536
rlabel metal2 30 -1407 30 -1407 0 net=6357
rlabel metal2 632 -1407 632 -1407 0 net=8114
rlabel metal2 677 -1407 677 -1407 0 net=7050
rlabel metal2 975 -1407 975 -1407 0 net=7649
rlabel metal2 1055 -1407 1055 -1407 0 net=8734
rlabel metal2 1444 -1407 1444 -1407 0 net=11237
rlabel metal2 1605 -1407 1605 -1407 0 net=11505
rlabel metal2 1738 -1407 1738 -1407 0 net=12793
rlabel metal2 1787 -1407 1787 -1407 0 net=13089
rlabel metal2 1885 -1407 1885 -1407 0 net=13625
rlabel metal2 47 -1409 47 -1409 0 net=10725
rlabel metal2 1556 -1409 1556 -1409 0 net=10795
rlabel metal2 1661 -1409 1661 -1409 0 net=11927
rlabel metal2 1794 -1409 1794 -1409 0 net=13459
rlabel metal2 51 -1411 51 -1411 0 net=13141
rlabel metal2 51 -1413 51 -1413 0 net=2103
rlabel metal2 107 -1413 107 -1413 0 net=3547
rlabel metal2 450 -1413 450 -1413 0 net=6651
rlabel metal2 814 -1413 814 -1413 0 net=6825
rlabel metal2 975 -1413 975 -1413 0 net=5343
rlabel metal2 1335 -1413 1335 -1413 0 net=13744
rlabel metal2 58 -1415 58 -1415 0 net=6810
rlabel metal2 548 -1415 548 -1415 0 net=3911
rlabel metal2 814 -1415 814 -1415 0 net=6551
rlabel metal2 849 -1415 849 -1415 0 net=6685
rlabel metal2 947 -1415 947 -1415 0 net=10224
rlabel metal2 1437 -1415 1437 -1415 0 net=10005
rlabel metal2 1801 -1415 1801 -1415 0 net=13161
rlabel metal2 58 -1417 58 -1417 0 net=7954
rlabel metal2 408 -1417 408 -1417 0 net=3573
rlabel metal2 562 -1417 562 -1417 0 net=2598
rlabel metal2 744 -1417 744 -1417 0 net=5509
rlabel metal2 877 -1417 877 -1417 0 net=7469
rlabel metal2 877 -1417 877 -1417 0 net=7469
rlabel metal2 905 -1417 905 -1417 0 net=6431
rlabel metal2 922 -1417 922 -1417 0 net=13657
rlabel metal2 65 -1419 65 -1419 0 net=2059
rlabel metal2 79 -1419 79 -1419 0 net=3883
rlabel metal2 408 -1419 408 -1419 0 net=4539
rlabel metal2 562 -1419 562 -1419 0 net=3761
rlabel metal2 744 -1419 744 -1419 0 net=9473
rlabel metal2 842 -1419 842 -1419 0 net=6421
rlabel metal2 926 -1419 926 -1419 0 net=6707
rlabel metal2 961 -1419 961 -1419 0 net=8218
rlabel metal2 1185 -1419 1185 -1419 0 net=8939
rlabel metal2 1283 -1419 1283 -1419 0 net=13378
rlabel metal2 1850 -1419 1850 -1419 0 net=13447
rlabel metal2 79 -1421 79 -1421 0 net=5953
rlabel metal2 884 -1421 884 -1421 0 net=6637
rlabel metal2 985 -1421 985 -1421 0 net=9412
rlabel metal2 1521 -1421 1521 -1421 0 net=10713
rlabel metal2 1577 -1421 1577 -1421 0 net=12055
rlabel metal2 1703 -1421 1703 -1421 0 net=12401
rlabel metal2 82 -1423 82 -1423 0 net=8032
rlabel metal2 1164 -1423 1164 -1423 0 net=8673
rlabel metal2 1283 -1423 1283 -1423 0 net=9143
rlabel metal2 1346 -1423 1346 -1423 0 net=9291
rlabel metal2 1374 -1423 1374 -1423 0 net=9587
rlabel metal2 1507 -1423 1507 -1423 0 net=10579
rlabel metal2 1535 -1423 1535 -1423 0 net=10789
rlabel metal2 1703 -1423 1703 -1423 0 net=12845
rlabel metal2 86 -1425 86 -1425 0 net=3417
rlabel metal2 194 -1425 194 -1425 0 net=5036
rlabel metal2 751 -1425 751 -1425 0 net=5447
rlabel metal2 982 -1425 982 -1425 0 net=7671
rlabel metal2 1150 -1425 1150 -1425 0 net=8155
rlabel metal2 1171 -1425 1171 -1425 0 net=9356
rlabel metal2 1479 -1425 1479 -1425 0 net=10447
rlabel metal2 1549 -1425 1549 -1425 0 net=12575
rlabel metal2 93 -1427 93 -1427 0 net=1523
rlabel metal2 114 -1427 114 -1427 0 net=4640
rlabel metal2 450 -1427 450 -1427 0 net=8091
rlabel metal2 583 -1427 583 -1427 0 net=7409
rlabel metal2 786 -1427 786 -1427 0 net=6143
rlabel metal2 982 -1427 982 -1427 0 net=11004
rlabel metal2 1717 -1427 1717 -1427 0 net=12745
rlabel metal2 93 -1429 93 -1429 0 net=2913
rlabel metal2 198 -1429 198 -1429 0 net=4574
rlabel metal2 247 -1429 247 -1429 0 net=4191
rlabel metal2 996 -1429 996 -1429 0 net=9327
rlabel metal2 1388 -1429 1388 -1429 0 net=9991
rlabel metal2 1549 -1429 1549 -1429 0 net=11623
rlabel metal2 1640 -1429 1640 -1429 0 net=10823
rlabel metal2 114 -1431 114 -1431 0 net=7443
rlabel metal2 492 -1431 492 -1431 0 net=2489
rlabel metal2 807 -1431 807 -1431 0 net=7915
rlabel metal2 1178 -1431 1178 -1431 0 net=9653
rlabel metal2 1759 -1431 1759 -1431 0 net=12565
rlabel metal2 121 -1433 121 -1433 0 net=8879
rlabel metal2 145 -1433 145 -1433 0 net=13303
rlabel metal2 145 -1435 145 -1435 0 net=8440
rlabel metal2 1248 -1435 1248 -1435 0 net=9185
rlabel metal2 1346 -1435 1346 -1435 0 net=10345
rlabel metal2 1752 -1435 1752 -1435 0 net=11429
rlabel metal2 149 -1437 149 -1437 0 net=3955
rlabel metal2 1111 -1437 1111 -1437 0 net=10822
rlabel metal2 198 -1439 198 -1439 0 net=4385
rlabel metal2 310 -1439 310 -1439 0 net=5907
rlabel metal2 793 -1439 793 -1439 0 net=6565
rlabel metal2 929 -1439 929 -1439 0 net=10225
rlabel metal2 1493 -1439 1493 -1439 0 net=12633
rlabel metal2 37 -1441 37 -1441 0 net=5203
rlabel metal2 303 -1441 303 -1441 0 net=2783
rlabel metal2 373 -1441 373 -1441 0 net=3307
rlabel metal2 506 -1441 506 -1441 0 net=3259
rlabel metal2 569 -1441 569 -1441 0 net=4190
rlabel metal2 954 -1441 954 -1441 0 net=7025
rlabel metal2 1003 -1441 1003 -1441 0 net=7970
rlabel metal2 1066 -1441 1066 -1441 0 net=11670
rlabel metal2 37 -1443 37 -1443 0 net=1801
rlabel metal2 86 -1443 86 -1443 0 net=4693
rlabel metal2 1006 -1443 1006 -1443 0 net=8434
rlabel metal2 1248 -1443 1248 -1443 0 net=9033
rlabel metal2 1367 -1443 1367 -1443 0 net=9377
rlabel metal2 1493 -1443 1493 -1443 0 net=10941
rlabel metal2 1633 -1443 1633 -1443 0 net=11857
rlabel metal2 1986 -1443 1986 -1443 0 net=1
rlabel metal2 110 -1445 110 -1445 0 net=7529
rlabel metal2 338 -1445 338 -1445 0 net=2203
rlabel metal2 387 -1445 387 -1445 0 net=8519
rlabel metal2 1255 -1445 1255 -1445 0 net=9363
rlabel metal2 1528 -1445 1528 -1445 0 net=10739
rlabel metal2 128 -1447 128 -1447 0 net=10963
rlabel metal2 128 -1449 128 -1449 0 net=1647
rlabel metal2 205 -1449 205 -1449 0 net=3325
rlabel metal2 233 -1449 233 -1449 0 net=8884
rlabel metal2 1367 -1449 1367 -1449 0 net=10611
rlabel metal2 1486 -1449 1486 -1449 0 net=10465
rlabel metal2 1563 -1449 1563 -1449 0 net=10893
rlabel metal2 135 -1451 135 -1451 0 net=2091
rlabel metal2 226 -1451 226 -1451 0 net=1837
rlabel metal2 338 -1451 338 -1451 0 net=3793
rlabel metal2 555 -1451 555 -1451 0 net=3803
rlabel metal2 576 -1451 576 -1451 0 net=992
rlabel metal2 1010 -1451 1010 -1451 0 net=7713
rlabel metal2 296 -1453 296 -1453 0 net=1937
rlabel metal2 387 -1453 387 -1453 0 net=2235
rlabel metal2 422 -1453 422 -1453 0 net=3679
rlabel metal2 590 -1453 590 -1453 0 net=4315
rlabel metal2 663 -1453 663 -1453 0 net=9965
rlabel metal2 163 -1455 163 -1455 0 net=3077
rlabel metal2 415 -1455 415 -1455 0 net=2941
rlabel metal2 513 -1455 513 -1455 0 net=4477
rlabel metal2 618 -1455 618 -1455 0 net=7211
rlabel metal2 793 -1455 793 -1455 0 net=5149
rlabel metal2 898 -1455 898 -1455 0 net=7081
rlabel metal2 1024 -1455 1024 -1455 0 net=13137
rlabel metal2 163 -1457 163 -1457 0 net=1613
rlabel metal2 415 -1457 415 -1457 0 net=4337
rlabel metal2 478 -1457 478 -1457 0 net=3489
rlabel metal2 821 -1457 821 -1457 0 net=6249
rlabel metal2 1031 -1457 1031 -1457 0 net=11261
rlabel metal2 212 -1459 212 -1459 0 net=1821
rlabel metal2 520 -1459 520 -1459 0 net=5069
rlabel metal2 702 -1459 702 -1459 0 net=5389
rlabel metal2 989 -1459 989 -1459 0 net=7679
rlabel metal2 1034 -1459 1034 -1459 0 net=11215
rlabel metal2 177 -1461 177 -1461 0 net=6729
rlabel metal2 219 -1461 219 -1461 0 net=2267
rlabel metal2 443 -1461 443 -1461 0 net=3941
rlabel metal2 534 -1461 534 -1461 0 net=4769
rlabel metal2 751 -1461 751 -1461 0 net=7215
rlabel metal2 1087 -1461 1087 -1461 0 net=10643
rlabel metal2 191 -1463 191 -1463 0 net=3967
rlabel metal2 555 -1463 555 -1463 0 net=3597
rlabel metal2 191 -1465 191 -1465 0 net=5660
rlabel metal2 989 -1465 989 -1465 0 net=7197
rlabel metal2 1087 -1465 1087 -1465 0 net=7993
rlabel metal2 1108 -1465 1108 -1465 0 net=10247
rlabel metal2 219 -1467 219 -1467 0 net=2545
rlabel metal2 359 -1467 359 -1467 0 net=2797
rlabel metal2 576 -1467 576 -1467 0 net=3367
rlabel metal2 863 -1467 863 -1467 0 net=7135
rlabel metal2 1080 -1467 1080 -1467 0 net=8193
rlabel metal2 1111 -1467 1111 -1467 0 net=4459
rlabel metal2 1304 -1467 1304 -1467 0 net=13286
rlabel metal2 254 -1469 254 -1469 0 net=3025
rlabel metal2 275 -1469 275 -1469 0 net=3073
rlabel metal2 324 -1469 324 -1469 0 net=1727
rlabel metal2 590 -1469 590 -1469 0 net=1306
rlabel metal2 1080 -1469 1080 -1469 0 net=7665
rlabel metal2 1286 -1469 1286 -1469 0 net=9072
rlabel metal2 1402 -1469 1402 -1469 0 net=9857
rlabel metal2 1731 -1469 1731 -1469 0 net=12463
rlabel metal2 240 -1471 240 -1471 0 net=2873
rlabel metal2 275 -1471 275 -1471 0 net=1967
rlabel metal2 597 -1471 597 -1471 0 net=6340
rlabel metal2 670 -1471 670 -1471 0 net=9483
rlabel metal2 1724 -1471 1724 -1471 0 net=12423
rlabel metal2 324 -1473 324 -1473 0 net=4993
rlabel metal2 464 -1473 464 -1473 0 net=5771
rlabel metal2 604 -1473 604 -1473 0 net=4393
rlabel metal2 1115 -1473 1115 -1473 0 net=6102
rlabel metal2 1339 -1473 1339 -1473 0 net=10301
rlabel metal2 1696 -1473 1696 -1473 0 net=12379
rlabel metal2 352 -1475 352 -1475 0 net=4835
rlabel metal2 653 -1475 653 -1475 0 net=12605
rlabel metal2 1118 -1475 1118 -1475 0 net=12042
rlabel metal2 401 -1477 401 -1477 0 net=2017
rlabel metal2 541 -1477 541 -1477 0 net=3531
rlabel metal2 653 -1477 653 -1477 0 net=4069
rlabel metal2 1143 -1477 1143 -1477 0 net=8299
rlabel metal2 1160 -1477 1160 -1477 0 net=10289
rlabel metal2 1675 -1477 1675 -1477 0 net=12157
rlabel metal2 44 -1479 44 -1479 0 net=4225
rlabel metal2 604 -1479 604 -1479 0 net=4043
rlabel metal2 758 -1479 758 -1479 0 net=5535
rlabel metal2 779 -1479 779 -1479 0 net=6967
rlabel metal2 1059 -1479 1059 -1479 0 net=7801
rlabel metal2 1199 -1479 1199 -1479 0 net=8811
rlabel metal2 1220 -1479 1220 -1479 0 net=8839
rlabel metal2 1416 -1479 1416 -1479 0 net=10025
rlabel metal2 1584 -1479 1584 -1479 0 net=11031
rlabel metal2 44 -1481 44 -1481 0 net=13331
rlabel metal2 170 -1483 170 -1483 0 net=4915
rlabel metal2 856 -1483 856 -1483 0 net=6389
rlabel metal2 1122 -1483 1122 -1483 0 net=10857
rlabel metal2 61 -1485 61 -1485 0 net=2627
rlabel metal2 464 -1485 464 -1485 0 net=4667
rlabel metal2 611 -1485 611 -1485 0 net=1535
rlabel metal2 1101 -1485 1101 -1485 0 net=7565
rlabel metal2 1157 -1485 1157 -1485 0 net=8445
rlabel metal2 1244 -1485 1244 -1485 0 net=11787
rlabel metal2 61 -1487 61 -1487 0 net=5013
rlabel metal2 628 -1487 628 -1487 0 net=5198
rlabel metal2 870 -1487 870 -1487 0 net=6205
rlabel metal2 1059 -1487 1059 -1487 0 net=8145
rlabel metal2 1157 -1487 1157 -1487 0 net=13656
rlabel metal2 471 -1489 471 -1489 0 net=8503
rlabel metal2 1101 -1489 1101 -1489 0 net=8750
rlabel metal2 1318 -1489 1318 -1489 0 net=9749
rlabel metal2 1815 -1489 1815 -1489 0 net=12875
rlabel metal2 366 -1491 366 -1491 0 net=6775
rlabel metal2 688 -1491 688 -1491 0 net=5871
rlabel metal2 1129 -1491 1129 -1491 0 net=9665
rlabel metal2 1668 -1491 1668 -1491 0 net=11953
rlabel metal2 366 -1493 366 -1493 0 net=2379
rlabel metal2 716 -1493 716 -1493 0 net=7353
rlabel metal2 1192 -1493 1192 -1493 0 net=8467
rlabel metal2 1297 -1493 1297 -1493 0 net=9101
rlabel metal2 1598 -1493 1598 -1493 0 net=11311
rlabel metal2 380 -1495 380 -1495 0 net=5603
rlabel metal2 1192 -1495 1192 -1495 0 net=12933
rlabel metal2 660 -1497 660 -1497 0 net=5003
rlabel metal2 1269 -1497 1269 -1497 0 net=8907
rlabel metal2 1311 -1497 1311 -1497 0 net=10603
rlabel metal2 1598 -1497 1598 -1497 0 net=12365
rlabel metal2 156 -1499 156 -1499 0 net=7132
rlabel metal2 723 -1499 723 -1499 0 net=4855
rlabel metal2 1269 -1499 1269 -1499 0 net=8769
rlabel metal2 1619 -1499 1619 -1499 0 net=11545
rlabel metal2 156 -1501 156 -1501 0 net=1501
rlabel metal2 730 -1501 730 -1501 0 net=3737
rlabel metal2 1069 -1501 1069 -1501 0 net=10951
rlabel metal2 240 -1503 240 -1503 0 net=5181
rlabel metal2 1069 -1503 1069 -1503 0 net=12274
rlabel metal2 317 -1505 317 -1505 0 net=2299
rlabel metal2 1234 -1505 1234 -1505 0 net=8869
rlabel metal2 1465 -1505 1465 -1505 0 net=10309
rlabel metal2 317 -1507 317 -1507 0 net=2975
rlabel metal2 1227 -1507 1227 -1507 0 net=8805
rlabel metal2 1430 -1507 1430 -1507 0 net=10099
rlabel metal2 166 -1509 166 -1509 0 net=2053
rlabel metal2 625 -1509 625 -1509 0 net=8575
rlabel metal2 1353 -1509 1353 -1509 0 net=9919
rlabel metal2 625 -1511 625 -1511 0 net=10765
rlabel metal2 1332 -1513 1332 -1513 0 net=9245
rlabel metal2 1332 -1515 1332 -1515 0 net=10521
rlabel metal2 2 -1526 2 -1526 0 net=2052
rlabel metal2 58 -1526 58 -1526 0 net=12380
rlabel metal2 1780 -1526 1780 -1526 0 net=12795
rlabel metal2 1780 -1526 1780 -1526 0 net=12795
rlabel metal2 1808 -1526 1808 -1526 0 net=8394
rlabel metal2 1948 -1526 1948 -1526 0 net=12032
rlabel metal2 1979 -1526 1979 -1526 0 net=10270
rlabel metal2 2018 -1526 2018 -1526 0 net=9503
rlabel metal2 2018 -1526 2018 -1526 0 net=9503
rlabel metal2 2 -1528 2 -1528 0 net=6731
rlabel metal2 180 -1528 180 -1528 0 net=3026
rlabel metal2 338 -1528 338 -1528 0 net=3794
rlabel metal2 754 -1528 754 -1528 0 net=10790
rlabel metal2 1689 -1528 1689 -1528 0 net=11547
rlabel metal2 1766 -1528 1766 -1528 0 net=10333
rlabel metal2 1955 -1528 1955 -1528 0 net=8016
rlabel metal2 1983 -1528 1983 -1528 0 net=6698
rlabel metal2 23 -1530 23 -1530 0 net=2224
rlabel metal2 72 -1530 72 -1530 0 net=2061
rlabel metal2 72 -1530 72 -1530 0 net=2061
rlabel metal2 82 -1530 82 -1530 0 net=52
rlabel metal2 1108 -1530 1108 -1530 0 net=12464
rlabel metal2 23 -1532 23 -1532 0 net=4387
rlabel metal2 233 -1532 233 -1532 0 net=4994
rlabel metal2 338 -1532 338 -1532 0 net=1729
rlabel metal2 485 -1532 485 -1532 0 net=2006
rlabel metal2 663 -1532 663 -1532 0 net=9765
rlabel metal2 768 -1532 768 -1532 0 net=6552
rlabel metal2 884 -1532 884 -1532 0 net=4394
rlabel metal2 1192 -1532 1192 -1532 0 net=8806
rlabel metal2 1262 -1532 1262 -1532 0 net=10346
rlabel metal2 1356 -1532 1356 -1532 0 net=12424
rlabel metal2 1808 -1532 1808 -1532 0 net=13091
rlabel metal2 30 -1534 30 -1534 0 net=6358
rlabel metal2 954 -1534 954 -1534 0 net=12576
rlabel metal2 30 -1536 30 -1536 0 net=4193
rlabel metal2 254 -1536 254 -1536 0 net=5639
rlabel metal2 1101 -1536 1101 -1536 0 net=10302
rlabel metal2 1346 -1536 1346 -1536 0 net=9293
rlabel metal2 1437 -1536 1437 -1536 0 net=9967
rlabel metal2 1437 -1536 1437 -1536 0 net=9967
rlabel metal2 1503 -1536 1503 -1536 0 net=12566
rlabel metal2 37 -1538 37 -1538 0 net=1802
rlabel metal2 502 -1538 502 -1538 0 net=7748
rlabel metal2 1108 -1538 1108 -1538 0 net=7481
rlabel metal2 1339 -1538 1339 -1538 0 net=9247
rlabel metal2 1360 -1538 1360 -1538 0 net=9329
rlabel metal2 1514 -1538 1514 -1538 0 net=10523
rlabel metal2 1514 -1538 1514 -1538 0 net=10523
rlabel metal2 1591 -1538 1591 -1538 0 net=10006
rlabel metal2 37 -1540 37 -1540 0 net=2105
rlabel metal2 58 -1540 58 -1540 0 net=3549
rlabel metal2 117 -1540 117 -1540 0 net=8880
rlabel metal2 135 -1540 135 -1540 0 net=2093
rlabel metal2 135 -1540 135 -1540 0 net=2093
rlabel metal2 142 -1540 142 -1540 0 net=7530
rlabel metal2 324 -1540 324 -1540 0 net=2799
rlabel metal2 499 -1540 499 -1540 0 net=3599
rlabel metal2 593 -1540 593 -1540 0 net=5872
rlabel metal2 709 -1540 709 -1540 0 net=7470
rlabel metal2 905 -1540 905 -1540 0 net=6423
rlabel metal2 957 -1540 957 -1540 0 net=10117
rlabel metal2 1703 -1540 1703 -1540 0 net=12847
rlabel metal2 9 -1542 9 -1542 0 net=6479
rlabel metal2 86 -1542 86 -1542 0 net=4695
rlabel metal2 121 -1542 121 -1542 0 net=3419
rlabel metal2 194 -1542 194 -1542 0 net=8520
rlabel metal2 1234 -1542 1234 -1542 0 net=8841
rlabel metal2 1262 -1542 1262 -1542 0 net=7179
rlabel metal2 1325 -1542 1325 -1542 0 net=9187
rlabel metal2 1325 -1542 1325 -1542 0 net=9187
rlabel metal2 1353 -1542 1353 -1542 0 net=10466
rlabel metal2 1577 -1542 1577 -1542 0 net=12057
rlabel metal2 1717 -1542 1717 -1542 0 net=7715
rlabel metal2 9 -1544 9 -1544 0 net=1503
rlabel metal2 184 -1544 184 -1544 0 net=1915
rlabel metal2 548 -1544 548 -1544 0 net=3575
rlabel metal2 548 -1544 548 -1544 0 net=3575
rlabel metal2 555 -1544 555 -1544 0 net=4771
rlabel metal2 712 -1544 712 -1544 0 net=10726
rlabel metal2 1577 -1544 1577 -1544 0 net=10895
rlabel metal2 1661 -1544 1661 -1544 0 net=11567
rlabel metal2 44 -1546 44 -1546 0 net=1524
rlabel metal2 142 -1546 142 -1546 0 net=987
rlabel metal2 667 -1546 667 -1546 0 net=7916
rlabel metal2 1199 -1546 1199 -1546 0 net=8813
rlabel metal2 1265 -1546 1265 -1546 0 net=13768
rlabel metal2 1976 -1546 1976 -1546 0 net=11383
rlabel metal2 16 -1548 16 -1548 0 net=5419
rlabel metal2 79 -1548 79 -1548 0 net=10727
rlabel metal2 114 -1548 114 -1548 0 net=7444
rlabel metal2 674 -1548 674 -1548 0 net=4704
rlabel metal2 1111 -1548 1111 -1548 0 net=7078
rlabel metal2 1829 -1548 1829 -1548 0 net=13139
rlabel metal2 16 -1550 16 -1550 0 net=3129
rlabel metal2 145 -1550 145 -1550 0 net=5229
rlabel metal2 226 -1550 226 -1550 0 net=1839
rlabel metal2 289 -1550 289 -1550 0 net=3075
rlabel metal2 506 -1550 506 -1550 0 net=3261
rlabel metal2 506 -1550 506 -1550 0 net=3261
rlabel metal2 618 -1550 618 -1550 0 net=7213
rlabel metal2 1118 -1550 1118 -1550 0 net=8940
rlabel metal2 1199 -1550 1199 -1550 0 net=8447
rlabel metal2 1269 -1550 1269 -1550 0 net=8771
rlabel metal2 1269 -1550 1269 -1550 0 net=8771
rlabel metal2 1374 -1550 1374 -1550 0 net=9667
rlabel metal2 1493 -1550 1493 -1550 0 net=10943
rlabel metal2 1612 -1550 1612 -1550 0 net=10953
rlabel metal2 1731 -1550 1731 -1550 0 net=12635
rlabel metal2 1794 -1550 1794 -1550 0 net=13461
rlabel metal2 86 -1552 86 -1552 0 net=882
rlabel metal2 702 -1552 702 -1552 0 net=5391
rlabel metal2 835 -1552 835 -1552 0 net=5955
rlabel metal2 961 -1552 961 -1552 0 net=6575
rlabel metal2 1374 -1552 1374 -1552 0 net=9379
rlabel metal2 1493 -1552 1493 -1552 0 net=11313
rlabel metal2 1822 -1552 1822 -1552 0 net=13163
rlabel metal2 128 -1554 128 -1554 0 net=1648
rlabel metal2 156 -1554 156 -1554 0 net=2547
rlabel metal2 226 -1554 226 -1554 0 net=4351
rlabel metal2 1122 -1554 1122 -1554 0 net=7567
rlabel metal2 1122 -1554 1122 -1554 0 net=7567
rlabel metal2 1129 -1554 1129 -1554 0 net=1264
rlabel metal2 1906 -1554 1906 -1554 0 net=13627
rlabel metal2 93 -1556 93 -1556 0 net=2915
rlabel metal2 191 -1556 191 -1556 0 net=10031
rlabel metal2 233 -1556 233 -1556 0 net=2785
rlabel metal2 345 -1556 345 -1556 0 net=2054
rlabel metal2 681 -1556 681 -1556 0 net=3912
rlabel metal2 1307 -1556 1307 -1556 0 net=12765
rlabel metal2 1871 -1556 1871 -1556 0 net=12877
rlabel metal2 65 -1558 65 -1558 0 net=5015
rlabel metal2 163 -1558 163 -1558 0 net=1615
rlabel metal2 205 -1558 205 -1558 0 net=3327
rlabel metal2 415 -1558 415 -1558 0 net=4339
rlabel metal2 849 -1558 849 -1558 0 net=6145
rlabel metal2 971 -1558 971 -1558 0 net=9144
rlabel metal2 1307 -1558 1307 -1558 0 net=13448
rlabel metal2 1871 -1558 1871 -1558 0 net=13333
rlabel metal2 163 -1560 163 -1560 0 net=1847
rlabel metal2 663 -1560 663 -1560 0 net=13065
rlabel metal2 205 -1562 205 -1562 0 net=5071
rlabel metal2 646 -1562 646 -1562 0 net=4317
rlabel metal2 681 -1562 681 -1562 0 net=5511
rlabel metal2 863 -1562 863 -1562 0 net=12607
rlabel metal2 268 -1564 268 -1564 0 net=2875
rlabel metal2 397 -1564 397 -1564 0 net=4419
rlabel metal2 670 -1564 670 -1564 0 net=5448
rlabel metal2 996 -1564 996 -1564 0 net=7027
rlabel metal2 996 -1564 996 -1564 0 net=7027
rlabel metal2 1003 -1564 1003 -1564 0 net=12402
rlabel metal2 268 -1566 268 -1566 0 net=3805
rlabel metal2 583 -1566 583 -1566 0 net=3681
rlabel metal2 968 -1566 968 -1566 0 net=6827
rlabel metal2 1073 -1566 1073 -1566 0 net=7325
rlabel metal2 1132 -1566 1132 -1566 0 net=10604
rlabel metal2 1332 -1566 1332 -1566 0 net=13578
rlabel metal2 282 -1568 282 -1568 0 net=5205
rlabel metal2 569 -1568 569 -1568 0 net=3369
rlabel metal2 583 -1568 583 -1568 0 net=3739
rlabel metal2 800 -1568 800 -1568 0 net=3490
rlabel metal2 1132 -1568 1132 -1568 0 net=11624
rlabel metal2 1619 -1568 1619 -1568 0 net=10965
rlabel metal2 1647 -1568 1647 -1568 0 net=13259
rlabel metal2 1864 -1568 1864 -1568 0 net=13305
rlabel metal2 282 -1570 282 -1570 0 net=8093
rlabel metal2 457 -1570 457 -1570 0 net=1822
rlabel metal2 723 -1570 723 -1570 0 net=5182
rlabel metal2 1213 -1570 1213 -1570 0 net=11239
rlabel metal2 1507 -1570 1507 -1570 0 net=10449
rlabel metal2 1647 -1570 1647 -1570 0 net=11217
rlabel metal2 1668 -1570 1668 -1570 0 net=11789
rlabel metal2 1787 -1570 1787 -1570 0 net=12935
rlabel metal2 1913 -1570 1913 -1570 0 net=13659
rlabel metal2 261 -1572 261 -1572 0 net=3885
rlabel metal2 464 -1572 464 -1572 0 net=4669
rlabel metal2 723 -1572 723 -1572 0 net=2829
rlabel metal2 1024 -1572 1024 -1572 0 net=7217
rlabel metal2 1150 -1572 1150 -1572 0 net=8301
rlabel metal2 1283 -1572 1283 -1572 0 net=11262
rlabel metal2 1654 -1572 1654 -1572 0 net=11507
rlabel metal2 1696 -1572 1696 -1572 0 net=12991
rlabel metal2 1941 -1572 1941 -1572 0 net=8171
rlabel metal2 261 -1574 261 -1574 0 net=2573
rlabel metal2 1171 -1574 1171 -1574 0 net=8675
rlabel metal2 1311 -1574 1311 -1574 0 net=9103
rlabel metal2 1395 -1574 1395 -1574 0 net=9485
rlabel metal2 1444 -1574 1444 -1574 0 net=10101
rlabel metal2 1521 -1574 1521 -1574 0 net=10581
rlabel metal2 1542 -1574 1542 -1574 0 net=10859
rlabel metal2 1626 -1574 1626 -1574 0 net=11859
rlabel metal2 1787 -1574 1787 -1574 0 net=13503
rlabel metal2 65 -1576 65 -1576 0 net=11487
rlabel metal2 1843 -1576 1843 -1576 0 net=5961
rlabel metal2 289 -1578 289 -1578 0 net=2381
rlabel metal2 418 -1578 418 -1578 0 net=5577
rlabel metal2 919 -1578 919 -1578 0 net=10451
rlabel metal2 1521 -1578 1521 -1578 0 net=10797
rlabel metal2 296 -1580 296 -1580 0 net=2269
rlabel metal2 366 -1580 366 -1580 0 net=2301
rlabel metal2 443 -1580 443 -1580 0 net=4071
rlabel metal2 730 -1580 730 -1580 0 net=5345
rlabel metal2 1006 -1580 1006 -1580 0 net=12369
rlabel metal2 114 -1582 114 -1582 0 net=6885
rlabel metal2 772 -1582 772 -1582 0 net=5537
rlabel metal2 807 -1582 807 -1582 0 net=6567
rlabel metal2 968 -1582 968 -1582 0 net=7198
rlabel metal2 1024 -1582 1024 -1582 0 net=7673
rlabel metal2 1185 -1582 1185 -1582 0 net=9035
rlabel metal2 1290 -1582 1290 -1582 0 net=4460
rlabel metal2 1549 -1582 1549 -1582 0 net=10715
rlabel metal2 1563 -1582 1563 -1582 0 net=10767
rlabel metal2 1598 -1582 1598 -1582 0 net=12367
rlabel metal2 296 -1584 296 -1584 0 net=4287
rlabel metal2 989 -1584 989 -1584 0 net=6755
rlabel metal2 1220 -1584 1220 -1584 0 net=8469
rlabel metal2 1290 -1584 1290 -1584 0 net=8909
rlabel metal2 1402 -1584 1402 -1584 0 net=9751
rlabel metal2 1535 -1584 1535 -1584 0 net=10645
rlabel metal2 1598 -1584 1598 -1584 0 net=10825
rlabel metal2 303 -1586 303 -1586 0 net=1939
rlabel metal2 422 -1586 422 -1586 0 net=2943
rlabel metal2 478 -1586 478 -1586 0 net=3943
rlabel metal2 765 -1586 765 -1586 0 net=5005
rlabel metal2 793 -1586 793 -1586 0 net=5151
rlabel metal2 817 -1586 817 -1586 0 net=13205
rlabel metal2 212 -1588 212 -1588 0 net=9159
rlabel metal2 429 -1588 429 -1588 0 net=6877
rlabel metal2 1031 -1588 1031 -1588 0 net=7681
rlabel metal2 1164 -1588 1164 -1588 0 net=8157
rlabel metal2 1367 -1588 1367 -1588 0 net=10613
rlabel metal2 1570 -1588 1570 -1588 0 net=10741
rlabel metal2 170 -1590 170 -1590 0 net=2629
rlabel metal2 317 -1590 317 -1590 0 net=2977
rlabel metal2 478 -1590 478 -1590 0 net=4479
rlabel metal2 597 -1590 597 -1590 0 net=5773
rlabel metal2 922 -1590 922 -1590 0 net=11033
rlabel metal2 317 -1592 317 -1592 0 net=1537
rlabel metal2 793 -1592 793 -1592 0 net=6391
rlabel metal2 884 -1592 884 -1592 0 net=5975
rlabel metal2 926 -1592 926 -1592 0 net=6709
rlabel metal2 1010 -1592 1010 -1592 0 net=7083
rlabel metal2 1059 -1592 1059 -1592 0 net=8147
rlabel metal2 1367 -1592 1367 -1592 0 net=9365
rlabel metal2 1416 -1592 1416 -1592 0 net=9859
rlabel metal2 79 -1594 79 -1594 0 net=10377
rlabel metal2 1080 -1594 1080 -1594 0 net=7667
rlabel metal2 1195 -1594 1195 -1594 0 net=10887
rlabel metal2 331 -1596 331 -1596 0 net=2237
rlabel metal2 513 -1596 513 -1596 0 net=4227
rlabel metal2 611 -1596 611 -1596 0 net=1805
rlabel metal2 828 -1596 828 -1596 0 net=8237
rlabel metal2 1220 -1596 1220 -1596 0 net=8871
rlabel metal2 1388 -1596 1388 -1596 0 net=9993
rlabel metal2 387 -1598 387 -1598 0 net=2509
rlabel metal2 856 -1598 856 -1598 0 net=6207
rlabel metal2 912 -1598 912 -1598 0 net=6433
rlabel metal2 933 -1598 933 -1598 0 net=6639
rlabel metal2 1080 -1598 1080 -1598 0 net=8577
rlabel metal2 1241 -1598 1241 -1598 0 net=11954
rlabel metal2 177 -1600 177 -1600 0 net=10543
rlabel metal2 940 -1600 940 -1600 0 net=6687
rlabel metal2 1227 -1600 1227 -1600 0 net=9589
rlabel metal2 1423 -1600 1423 -1600 0 net=9921
rlabel metal2 1451 -1600 1451 -1600 0 net=10227
rlabel metal2 1815 -1600 1815 -1600 0 net=13143
rlabel metal2 352 -1602 352 -1602 0 net=4837
rlabel metal2 1458 -1602 1458 -1602 0 net=10027
rlabel metal2 352 -1604 352 -1604 0 net=3763
rlabel metal2 870 -1604 870 -1604 0 net=8505
rlabel metal2 1458 -1604 1458 -1604 0 net=10249
rlabel metal2 380 -1606 380 -1606 0 net=5604
rlabel metal2 1094 -1606 1094 -1606 0 net=8195
rlabel metal2 1479 -1606 1479 -1606 0 net=10291
rlabel metal2 380 -1608 380 -1608 0 net=2491
rlabel metal2 534 -1608 534 -1608 0 net=3969
rlabel metal2 786 -1608 786 -1608 0 net=5909
rlabel metal2 891 -1608 891 -1608 0 net=9655
rlabel metal2 1206 -1608 1206 -1608 0 net=13601
rlabel metal2 394 -1610 394 -1610 0 net=3079
rlabel metal2 541 -1610 541 -1610 0 net=4593
rlabel metal2 744 -1610 744 -1610 0 net=9475
rlabel metal2 898 -1610 898 -1610 0 net=6251
rlabel metal2 1045 -1610 1045 -1610 0 net=7281
rlabel metal2 1244 -1610 1244 -1610 0 net=6275
rlabel metal2 173 -1612 173 -1612 0 net=7149
rlabel metal2 898 -1612 898 -1612 0 net=6107
rlabel metal2 1087 -1612 1087 -1612 0 net=7995
rlabel metal2 1486 -1612 1486 -1612 0 net=10311
rlabel metal2 82 -1614 82 -1614 0 net=1321
rlabel metal2 1500 -1614 1500 -1614 0 net=11032
rlabel metal2 394 -1616 394 -1616 0 net=5677
rlabel metal2 1017 -1616 1017 -1616 0 net=7137
rlabel metal2 1675 -1616 1675 -1616 0 net=11929
rlabel metal2 471 -1618 471 -1618 0 net=6777
rlabel metal2 562 -1618 562 -1618 0 net=4011
rlabel metal2 1738 -1618 1738 -1618 0 net=12159
rlabel metal2 471 -1620 471 -1620 0 net=3009
rlabel metal2 779 -1620 779 -1620 0 net=6969
rlabel metal2 1045 -1620 1045 -1620 0 net=6865
rlabel metal2 1745 -1620 1745 -1620 0 net=12747
rlabel metal2 408 -1622 408 -1622 0 net=4541
rlabel metal2 695 -1622 695 -1622 0 net=7411
rlabel metal2 1143 -1622 1143 -1622 0 net=7803
rlabel metal2 1759 -1622 1759 -1622 0 net=11431
rlabel metal2 408 -1624 408 -1624 0 net=2881
rlabel metal2 1052 -1624 1052 -1624 0 net=7651
rlabel metal2 1759 -1624 1759 -1624 0 net=10773
rlabel metal2 590 -1626 590 -1626 0 net=7355
rlabel metal2 1052 -1626 1052 -1626 0 net=13714
rlabel metal2 240 -1628 240 -1628 0 net=13513
rlabel metal2 240 -1630 240 -1630 0 net=2019
rlabel metal2 716 -1630 716 -1630 0 net=4917
rlabel metal2 401 -1632 401 -1632 0 net=3309
rlabel metal2 737 -1632 737 -1632 0 net=4857
rlabel metal2 373 -1634 373 -1634 0 net=2205
rlabel metal2 625 -1634 625 -1634 0 net=1316
rlabel metal2 275 -1636 275 -1636 0 net=1969
rlabel metal2 604 -1636 604 -1636 0 net=4045
rlabel metal2 149 -1638 149 -1638 0 net=3957
rlabel metal2 604 -1638 604 -1638 0 net=3533
rlabel metal2 149 -1640 149 -1640 0 net=3153
rlabel metal2 632 -1640 632 -1640 0 net=6653
rlabel metal2 632 -1642 632 -1642 0 net=3579
rlabel metal2 9 -1653 9 -1653 0 net=1504
rlabel metal2 670 -1653 670 -1653 0 net=4918
rlabel metal2 737 -1653 737 -1653 0 net=6276
rlabel metal2 1570 -1653 1570 -1653 0 net=10889
rlabel metal2 1570 -1653 1570 -1653 0 net=10889
rlabel metal2 1801 -1653 1801 -1653 0 net=12937
rlabel metal2 1801 -1653 1801 -1653 0 net=12937
rlabel metal2 1843 -1653 1843 -1653 0 net=12878
rlabel metal2 1937 -1653 1937 -1653 0 net=11384
rlabel metal2 2018 -1653 2018 -1653 0 net=9505
rlabel metal2 2018 -1653 2018 -1653 0 net=9505
rlabel metal2 9 -1655 9 -1655 0 net=2917
rlabel metal2 131 -1655 131 -1655 0 net=7214
rlabel metal2 1206 -1655 1206 -1655 0 net=12058
rlabel metal2 1815 -1655 1815 -1655 0 net=13145
rlabel metal2 1850 -1655 1850 -1655 0 net=7716
rlabel metal2 1941 -1655 1941 -1655 0 net=8173
rlabel metal2 44 -1657 44 -1657 0 net=5421
rlabel metal2 86 -1657 86 -1657 0 net=3959
rlabel metal2 324 -1657 324 -1657 0 net=2800
rlabel metal2 590 -1657 590 -1657 0 net=7356
rlabel metal2 842 -1657 842 -1657 0 net=3682
rlabel metal2 1206 -1657 1206 -1657 0 net=8911
rlabel metal2 1332 -1657 1332 -1657 0 net=13039
rlabel metal2 1850 -1657 1850 -1657 0 net=13261
rlabel metal2 1871 -1657 1871 -1657 0 net=13335
rlabel metal2 1871 -1657 1871 -1657 0 net=13335
rlabel metal2 1885 -1657 1885 -1657 0 net=13463
rlabel metal2 1885 -1657 1885 -1657 0 net=13463
rlabel metal2 1913 -1657 1913 -1657 0 net=13661
rlabel metal2 1913 -1657 1913 -1657 0 net=13661
rlabel metal2 1944 -1657 1944 -1657 0 net=2613
rlabel metal2 37 -1659 37 -1659 0 net=2107
rlabel metal2 51 -1659 51 -1659 0 net=6481
rlabel metal2 51 -1659 51 -1659 0 net=6481
rlabel metal2 65 -1659 65 -1659 0 net=4319
rlabel metal2 180 -1659 180 -1659 0 net=2270
rlabel metal2 422 -1659 422 -1659 0 net=9161
rlabel metal2 485 -1659 485 -1659 0 net=3076
rlabel metal2 709 -1659 709 -1659 0 net=9486
rlabel metal2 1451 -1659 1451 -1659 0 net=10229
rlabel metal2 1451 -1659 1451 -1659 0 net=10229
rlabel metal2 1468 -1659 1468 -1659 0 net=12992
rlabel metal2 1857 -1659 1857 -1659 0 net=13307
rlabel metal2 1948 -1659 1948 -1659 0 net=10335
rlabel metal2 37 -1661 37 -1661 0 net=3551
rlabel metal2 68 -1661 68 -1661 0 net=6778
rlabel metal2 541 -1661 541 -1661 0 net=5006
rlabel metal2 793 -1661 793 -1661 0 net=6392
rlabel metal2 1055 -1661 1055 -1661 0 net=8158
rlabel metal2 1332 -1661 1332 -1661 0 net=9861
rlabel metal2 1468 -1661 1468 -1661 0 net=11488
rlabel metal2 1822 -1661 1822 -1661 0 net=13165
rlabel metal2 1941 -1661 1941 -1661 0 net=1677
rlabel metal2 58 -1663 58 -1663 0 net=6879
rlabel metal2 478 -1663 478 -1663 0 net=4481
rlabel metal2 534 -1663 534 -1663 0 net=4047
rlabel metal2 688 -1663 688 -1663 0 net=4671
rlabel metal2 712 -1663 712 -1663 0 net=7419
rlabel metal2 1076 -1663 1076 -1663 0 net=969
rlabel metal2 1395 -1663 1395 -1663 0 net=9753
rlabel metal2 1416 -1663 1416 -1663 0 net=9923
rlabel metal2 1500 -1663 1500 -1663 0 net=12796
rlabel metal2 1794 -1663 1794 -1663 0 net=13067
rlabel metal2 72 -1665 72 -1665 0 net=2062
rlabel metal2 89 -1665 89 -1665 0 net=10118
rlabel metal2 1696 -1665 1696 -1665 0 net=10775
rlabel metal2 1766 -1665 1766 -1665 0 net=12849
rlabel metal2 72 -1667 72 -1667 0 net=5303
rlabel metal2 688 -1667 688 -1667 0 net=6757
rlabel metal2 1083 -1667 1083 -1667 0 net=5962
rlabel metal2 117 -1669 117 -1669 0 net=7668
rlabel metal2 1220 -1669 1220 -1669 0 net=8873
rlabel metal2 1297 -1669 1297 -1669 0 net=9383
rlabel metal2 1556 -1669 1556 -1669 0 net=10769
rlabel metal2 1640 -1669 1640 -1669 0 net=11035
rlabel metal2 1731 -1669 1731 -1669 0 net=12637
rlabel metal2 1906 -1669 1906 -1669 0 net=13629
rlabel metal2 128 -1671 128 -1671 0 net=689
rlabel metal2 985 -1671 985 -1671 0 net=11240
rlabel metal2 1262 -1671 1262 -1671 0 net=7181
rlabel metal2 1262 -1671 1262 -1671 0 net=7181
rlabel metal2 1286 -1671 1286 -1671 0 net=12368
rlabel metal2 156 -1673 156 -1673 0 net=2548
rlabel metal2 422 -1673 422 -1673 0 net=3601
rlabel metal2 523 -1673 523 -1673 0 net=12823
rlabel metal2 1899 -1673 1899 -1673 0 net=13603
rlabel metal2 114 -1675 114 -1675 0 net=778
rlabel metal2 429 -1675 429 -1675 0 net=2207
rlabel metal2 499 -1675 499 -1675 0 net=5183
rlabel metal2 1335 -1675 1335 -1675 0 net=12160
rlabel metal2 1752 -1675 1752 -1675 0 net=12767
rlabel metal2 1892 -1675 1892 -1675 0 net=13515
rlabel metal2 114 -1677 114 -1677 0 net=4073
rlabel metal2 541 -1677 541 -1677 0 net=3619
rlabel metal2 751 -1677 751 -1677 0 net=9767
rlabel metal2 1423 -1677 1423 -1677 0 net=9969
rlabel metal2 1521 -1677 1521 -1677 0 net=10799
rlabel metal2 1619 -1677 1619 -1677 0 net=10967
rlabel metal2 1654 -1677 1654 -1677 0 net=11509
rlabel metal2 1717 -1677 1717 -1677 0 net=12609
rlabel metal2 1752 -1677 1752 -1677 0 net=11433
rlabel metal2 1787 -1677 1787 -1677 0 net=13505
rlabel metal2 149 -1679 149 -1679 0 net=3155
rlabel metal2 443 -1679 443 -1679 0 net=4421
rlabel metal2 660 -1679 660 -1679 0 net=6579
rlabel metal2 943 -1679 943 -1679 0 net=11548
rlabel metal2 121 -1681 121 -1681 0 net=3421
rlabel metal2 156 -1681 156 -1681 0 net=1539
rlabel metal2 324 -1681 324 -1681 0 net=2883
rlabel metal2 481 -1681 481 -1681 0 net=6845
rlabel metal2 765 -1681 765 -1681 0 net=5775
rlabel metal2 901 -1681 901 -1681 0 net=7674
rlabel metal2 1087 -1681 1087 -1681 0 net=10028
rlabel metal2 1493 -1681 1493 -1681 0 net=11315
rlabel metal2 1626 -1681 1626 -1681 0 net=11861
rlabel metal2 121 -1683 121 -1683 0 net=7333
rlabel metal2 828 -1683 828 -1683 0 net=527
rlabel metal2 1185 -1683 1185 -1683 0 net=9037
rlabel metal2 1241 -1683 1241 -1683 0 net=11829
rlabel metal2 1675 -1683 1675 -1683 0 net=11931
rlabel metal2 184 -1685 184 -1685 0 net=1916
rlabel metal2 702 -1685 702 -1685 0 net=5393
rlabel metal2 800 -1685 800 -1685 0 net=5539
rlabel metal2 800 -1685 800 -1685 0 net=5539
rlabel metal2 831 -1685 831 -1685 0 net=8148
rlabel metal2 1339 -1685 1339 -1685 0 net=9249
rlabel metal2 1472 -1685 1472 -1685 0 net=10293
rlabel metal2 1591 -1685 1591 -1685 0 net=10945
rlabel metal2 1682 -1685 1682 -1685 0 net=12371
rlabel metal2 187 -1687 187 -1687 0 net=8506
rlabel metal2 1311 -1687 1311 -1687 0 net=9105
rlabel metal2 1542 -1687 1542 -1687 0 net=10861
rlabel metal2 1668 -1687 1668 -1687 0 net=11791
rlabel metal2 100 -1689 100 -1689 0 net=10729
rlabel metal2 1661 -1689 1661 -1689 0 net=11569
rlabel metal2 2 -1691 2 -1691 0 net=6733
rlabel metal2 201 -1691 201 -1691 0 net=1148
rlabel metal2 716 -1691 716 -1691 0 net=7219
rlabel metal2 1101 -1691 1101 -1691 0 net=11687
rlabel metal2 205 -1693 205 -1693 0 net=5073
rlabel metal2 254 -1693 254 -1693 0 net=5640
rlabel metal2 408 -1693 408 -1693 0 net=4013
rlabel metal2 583 -1693 583 -1693 0 net=3741
rlabel metal2 639 -1693 639 -1693 0 net=6655
rlabel metal2 842 -1693 842 -1693 0 net=5957
rlabel metal2 919 -1693 919 -1693 0 net=10646
rlabel metal2 1661 -1693 1661 -1693 0 net=12749
rlabel metal2 191 -1695 191 -1695 0 net=1617
rlabel metal2 275 -1695 275 -1695 0 net=3887
rlabel metal2 520 -1695 520 -1695 0 net=5207
rlabel metal2 737 -1695 737 -1695 0 net=1354
rlabel metal2 856 -1695 856 -1695 0 net=6209
rlabel metal2 856 -1695 856 -1695 0 net=6209
rlabel metal2 863 -1695 863 -1695 0 net=6253
rlabel metal2 919 -1695 919 -1695 0 net=4583
rlabel metal2 1241 -1695 1241 -1695 0 net=10413
rlabel metal2 1584 -1695 1584 -1695 0 net=10827
rlabel metal2 1745 -1695 1745 -1695 0 net=13207
rlabel metal2 191 -1697 191 -1697 0 net=1393
rlabel metal2 576 -1697 576 -1697 0 net=4595
rlabel metal2 740 -1697 740 -1697 0 net=4838
rlabel metal2 1479 -1697 1479 -1697 0 net=10313
rlabel metal2 1598 -1697 1598 -1697 0 net=10955
rlabel metal2 1808 -1697 1808 -1697 0 net=13093
rlabel metal2 198 -1699 198 -1699 0 net=5231
rlabel metal2 527 -1699 527 -1699 0 net=4543
rlabel metal2 583 -1699 583 -1699 0 net=5513
rlabel metal2 768 -1699 768 -1699 0 net=7005
rlabel metal2 1024 -1699 1024 -1699 0 net=8239
rlabel metal2 1185 -1699 1185 -1699 0 net=8449
rlabel metal2 1244 -1699 1244 -1699 0 net=12577
rlabel metal2 198 -1701 198 -1701 0 net=5578
rlabel metal2 877 -1701 877 -1701 0 net=6577
rlabel metal2 968 -1701 968 -1701 0 net=6867
rlabel metal2 1073 -1701 1073 -1701 0 net=13140
rlabel metal2 205 -1703 205 -1703 0 net=3081
rlabel metal2 527 -1703 527 -1703 0 net=3581
rlabel metal2 681 -1703 681 -1703 0 net=12509
rlabel metal2 219 -1705 219 -1705 0 net=10033
rlabel metal2 1129 -1705 1129 -1705 0 net=13019
rlabel metal2 219 -1707 219 -1707 0 net=2575
rlabel metal2 317 -1707 317 -1707 0 net=1731
rlabel metal2 359 -1707 359 -1707 0 net=2945
rlabel metal2 492 -1707 492 -1707 0 net=5347
rlabel metal2 772 -1707 772 -1707 0 net=7139
rlabel metal2 1122 -1707 1122 -1707 0 net=7569
rlabel metal2 1132 -1707 1132 -1707 0 net=13071
rlabel metal2 261 -1709 261 -1709 0 net=3263
rlabel metal2 590 -1709 590 -1709 0 net=3971
rlabel metal2 604 -1709 604 -1709 0 net=3535
rlabel metal2 786 -1709 786 -1709 0 net=9477
rlabel metal2 1311 -1709 1311 -1709 0 net=10399
rlabel metal2 1612 -1709 1612 -1709 0 net=11219
rlabel metal2 310 -1711 310 -1711 0 net=2877
rlabel metal2 373 -1711 373 -1711 0 net=1970
rlabel metal2 849 -1711 849 -1711 0 net=6109
rlabel metal2 912 -1711 912 -1711 0 net=6435
rlabel metal2 933 -1711 933 -1711 0 net=10545
rlabel metal2 282 -1713 282 -1713 0 net=8095
rlabel metal2 373 -1713 373 -1713 0 net=3311
rlabel metal2 457 -1713 457 -1713 0 net=2979
rlabel metal2 506 -1713 506 -1713 0 net=2831
rlabel metal2 922 -1713 922 -1713 0 net=6424
rlabel metal2 961 -1713 961 -1713 0 net=6829
rlabel metal2 1041 -1713 1041 -1713 0 net=7659
rlabel metal2 1136 -1713 1136 -1713 0 net=7805
rlabel metal2 1199 -1713 1199 -1713 0 net=8471
rlabel metal2 1269 -1713 1269 -1713 0 net=8773
rlabel metal2 1318 -1713 1318 -1713 0 net=13769
rlabel metal2 142 -1715 142 -1715 0 net=8789
rlabel metal2 569 -1715 569 -1715 0 net=3371
rlabel metal2 632 -1715 632 -1715 0 net=4257
rlabel metal2 723 -1715 723 -1715 0 net=5911
rlabel metal2 943 -1715 943 -1715 0 net=7509
rlabel metal2 1157 -1715 1157 -1715 0 net=8303
rlabel metal2 1244 -1715 1244 -1715 0 net=10742
rlabel metal2 93 -1717 93 -1717 0 net=5017
rlabel metal2 194 -1717 194 -1717 0 net=11177
rlabel metal2 93 -1719 93 -1719 0 net=3515
rlabel metal2 653 -1719 653 -1719 0 net=6887
rlabel metal2 947 -1719 947 -1719 0 net=6711
rlabel metal2 996 -1719 996 -1719 0 net=7029
rlabel metal2 1066 -1719 1066 -1719 0 net=7683
rlabel metal2 1192 -1719 1192 -1719 0 net=9295
rlabel metal2 1353 -1719 1353 -1719 0 net=10450
rlabel metal2 16 -1721 16 -1721 0 net=3130
rlabel metal2 1010 -1721 1010 -1721 0 net=10379
rlabel metal2 16 -1723 16 -1723 0 net=6593
rlabel metal2 184 -1723 184 -1723 0 net=7091
rlabel metal2 1150 -1723 1150 -1723 0 net=7997
rlabel metal2 1248 -1723 1248 -1723 0 net=9189
rlabel metal2 1339 -1723 1339 -1723 0 net=10525
rlabel metal2 170 -1725 170 -1725 0 net=3807
rlabel metal2 397 -1725 397 -1725 0 net=4340
rlabel metal2 870 -1725 870 -1725 0 net=6147
rlabel metal2 971 -1725 971 -1725 0 net=12293
rlabel metal2 1507 -1725 1507 -1725 0 net=10453
rlabel metal2 233 -1727 233 -1727 0 net=2787
rlabel metal2 569 -1727 569 -1727 0 net=1807
rlabel metal2 646 -1727 646 -1727 0 net=7319
rlabel metal2 1171 -1727 1171 -1727 0 net=8677
rlabel metal2 1227 -1727 1227 -1727 0 net=9591
rlabel metal2 1356 -1727 1356 -1727 0 net=12587
rlabel metal2 233 -1729 233 -1729 0 net=1941
rlabel metal2 597 -1729 597 -1729 0 net=8337
rlabel metal2 1220 -1729 1220 -1729 0 net=8395
rlabel metal2 1388 -1729 1388 -1729 0 net=9995
rlabel metal2 1507 -1729 1507 -1729 0 net=10897
rlabel metal2 240 -1731 240 -1731 0 net=2021
rlabel metal2 611 -1731 611 -1731 0 net=3945
rlabel metal2 653 -1731 653 -1731 0 net=4653
rlabel metal2 1388 -1731 1388 -1731 0 net=10103
rlabel metal2 226 -1733 226 -1733 0 net=4353
rlabel metal2 821 -1733 821 -1733 0 net=5679
rlabel metal2 891 -1733 891 -1733 0 net=9657
rlabel metal2 1444 -1733 1444 -1733 0 net=10615
rlabel metal2 226 -1735 226 -1735 0 net=2239
rlabel metal2 807 -1735 807 -1735 0 net=5153
rlabel metal2 891 -1735 891 -1735 0 net=6569
rlabel metal2 1080 -1735 1080 -1735 0 net=8579
rlabel metal2 1227 -1735 1227 -1735 0 net=8843
rlabel metal2 1269 -1735 1269 -1735 0 net=9331
rlabel metal2 1528 -1735 1528 -1735 0 net=10583
rlabel metal2 240 -1737 240 -1737 0 net=2619
rlabel metal2 898 -1737 898 -1737 0 net=11991
rlabel metal2 247 -1739 247 -1739 0 net=1841
rlabel metal2 331 -1739 331 -1739 0 net=3765
rlabel metal2 905 -1739 905 -1739 0 net=6641
rlabel metal2 1234 -1739 1234 -1739 0 net=9367
rlabel metal2 1528 -1739 1528 -1739 0 net=10717
rlabel metal2 247 -1741 247 -1741 0 net=3329
rlabel metal2 352 -1741 352 -1741 0 net=3577
rlabel metal2 933 -1741 933 -1741 0 net=5873
rlabel metal2 1304 -1741 1304 -1741 0 net=11395
rlabel metal2 268 -1743 268 -1743 0 net=2303
rlabel metal2 513 -1743 513 -1743 0 net=4229
rlabel metal2 954 -1743 954 -1743 0 net=6841
rlabel metal2 23 -1745 23 -1745 0 net=4389
rlabel metal2 513 -1745 513 -1745 0 net=4318
rlabel metal2 975 -1745 975 -1745 0 net=6971
rlabel metal2 1307 -1745 1307 -1745 0 net=13481
rlabel metal2 23 -1747 23 -1747 0 net=10425
rlabel metal2 674 -1747 674 -1747 0 net=7413
rlabel metal2 1052 -1747 1052 -1747 0 net=907
rlabel metal2 1360 -1747 1360 -1747 0 net=1068
rlabel metal2 1367 -1747 1367 -1747 0 net=10251
rlabel metal2 289 -1749 289 -1749 0 net=2383
rlabel metal2 744 -1749 744 -1749 0 net=7151
rlabel metal2 1052 -1749 1052 -1749 0 net=7483
rlabel metal2 1374 -1749 1374 -1749 0 net=9381
rlabel metal2 289 -1751 289 -1751 0 net=2493
rlabel metal2 744 -1751 744 -1751 0 net=4859
rlabel metal2 779 -1751 779 -1751 0 net=7085
rlabel metal2 1374 -1751 1374 -1751 0 net=9669
rlabel metal2 1409 -1751 1409 -1751 0 net=8197
rlabel metal2 107 -1753 107 -1753 0 net=4697
rlabel metal2 758 -1753 758 -1753 0 net=5977
rlabel metal2 1031 -1753 1031 -1753 0 net=7283
rlabel metal2 1115 -1753 1115 -1753 0 net=7327
rlabel metal2 107 -1755 107 -1755 0 net=2095
rlabel metal2 695 -1755 695 -1755 0 net=7331
rlabel metal2 1115 -1755 1115 -1755 0 net=7653
rlabel metal2 1381 -1755 1381 -1755 0 net=9725
rlabel metal2 135 -1757 135 -1757 0 net=1849
rlabel metal2 565 -1757 565 -1757 0 net=7941
rlabel metal2 163 -1759 163 -1759 0 net=2631
rlabel metal2 695 -1759 695 -1759 0 net=6688
rlabel metal2 212 -1761 212 -1761 0 net=2511
rlabel metal2 1059 -1761 1059 -1761 0 net=8815
rlabel metal2 296 -1763 296 -1763 0 net=4289
rlabel metal2 516 -1763 516 -1763 0 net=9297
rlabel metal2 296 -1765 296 -1765 0 net=3011
rlabel metal2 30 -1767 30 -1767 0 net=4195
rlabel metal2 30 -1769 30 -1769 0 net=4773
rlabel metal2 555 -1771 555 -1771 0 net=145
rlabel metal2 65 -1782 65 -1782 0 net=5753
rlabel metal2 93 -1782 93 -1782 0 net=3516
rlabel metal2 170 -1782 170 -1782 0 net=3808
rlabel metal2 527 -1782 527 -1782 0 net=3583
rlabel metal2 555 -1782 555 -1782 0 net=5394
rlabel metal2 810 -1782 810 -1782 0 net=13770
rlabel metal2 1955 -1782 1955 -1782 0 net=10337
rlabel metal2 2011 -1782 2011 -1782 0 net=9506
rlabel metal2 65 -1784 65 -1784 0 net=3889
rlabel metal2 282 -1784 282 -1784 0 net=1842
rlabel metal2 506 -1784 506 -1784 0 net=2833
rlabel metal2 590 -1784 590 -1784 0 net=3973
rlabel metal2 590 -1784 590 -1784 0 net=3973
rlabel metal2 597 -1784 597 -1784 0 net=6148
rlabel metal2 884 -1784 884 -1784 0 net=11036
rlabel metal2 1878 -1784 1878 -1784 0 net=13483
rlabel metal2 1962 -1784 1962 -1784 0 net=2615
rlabel metal2 93 -1786 93 -1786 0 net=2097
rlabel metal2 114 -1786 114 -1786 0 net=4074
rlabel metal2 198 -1786 198 -1786 0 net=6578
rlabel metal2 884 -1786 884 -1786 0 net=13709
rlabel metal2 107 -1788 107 -1788 0 net=5185
rlabel metal2 527 -1788 527 -1788 0 net=2659
rlabel metal2 1080 -1788 1080 -1788 0 net=11651
rlabel metal2 1878 -1788 1878 -1788 0 net=12853
rlabel metal2 1969 -1788 1969 -1788 0 net=8175
rlabel metal2 114 -1790 114 -1790 0 net=2513
rlabel metal2 254 -1790 254 -1790 0 net=1618
rlabel metal2 695 -1790 695 -1790 0 net=6888
rlabel metal2 943 -1790 943 -1790 0 net=9106
rlabel metal2 1500 -1790 1500 -1790 0 net=10415
rlabel metal2 1500 -1790 1500 -1790 0 net=10415
rlabel metal2 1521 -1790 1521 -1790 0 net=10547
rlabel metal2 1521 -1790 1521 -1790 0 net=10547
rlabel metal2 1566 -1790 1566 -1790 0 net=13464
rlabel metal2 1892 -1790 1892 -1790 0 net=13507
rlabel metal2 58 -1792 58 -1792 0 net=6881
rlabel metal2 254 -1792 254 -1792 0 net=2495
rlabel metal2 303 -1792 303 -1792 0 net=2023
rlabel metal2 303 -1792 303 -1792 0 net=2023
rlabel metal2 310 -1792 310 -1792 0 net=8097
rlabel metal2 870 -1792 870 -1792 0 net=5875
rlabel metal2 947 -1792 947 -1792 0 net=6713
rlabel metal2 947 -1792 947 -1792 0 net=6713
rlabel metal2 968 -1792 968 -1792 0 net=6869
rlabel metal2 968 -1792 968 -1792 0 net=6869
rlabel metal2 985 -1792 985 -1792 0 net=10890
rlabel metal2 1584 -1792 1584 -1792 0 net=10829
rlabel metal2 1584 -1792 1584 -1792 0 net=10829
rlabel metal2 1619 -1792 1619 -1792 0 net=11317
rlabel metal2 1619 -1792 1619 -1792 0 net=11317
rlabel metal2 1829 -1792 1829 -1792 0 net=13073
rlabel metal2 1899 -1792 1899 -1792 0 net=13517
rlabel metal2 16 -1794 16 -1794 0 net=6594
rlabel metal2 128 -1794 128 -1794 0 net=1851
rlabel metal2 138 -1794 138 -1794 0 net=1909
rlabel metal2 352 -1794 352 -1794 0 net=3578
rlabel metal2 499 -1794 499 -1794 0 net=3743
rlabel metal2 649 -1794 649 -1794 0 net=6656
rlabel metal2 898 -1794 898 -1794 0 net=7421
rlabel metal2 1059 -1794 1059 -1794 0 net=8816
rlabel metal2 1080 -1794 1080 -1794 0 net=7511
rlabel metal2 1090 -1794 1090 -1794 0 net=8912
rlabel metal2 1209 -1794 1209 -1794 0 net=10946
rlabel metal2 1731 -1794 1731 -1794 0 net=12611
rlabel metal2 1843 -1794 1843 -1794 0 net=13147
rlabel metal2 1906 -1794 1906 -1794 0 net=13605
rlabel metal2 9 -1796 9 -1796 0 net=2918
rlabel metal2 142 -1796 142 -1796 0 net=5019
rlabel metal2 352 -1796 352 -1796 0 net=2947
rlabel metal2 366 -1796 366 -1796 0 net=4390
rlabel metal2 583 -1796 583 -1796 0 net=5515
rlabel metal2 600 -1796 600 -1796 0 net=5208
rlabel metal2 719 -1796 719 -1796 0 net=5074
rlabel metal2 744 -1796 744 -1796 0 net=4861
rlabel metal2 744 -1796 744 -1796 0 net=4861
rlabel metal2 751 -1796 751 -1796 0 net=6847
rlabel metal2 908 -1796 908 -1796 0 net=7332
rlabel metal2 1104 -1796 1104 -1796 0 net=10616
rlabel metal2 1468 -1796 1468 -1796 0 net=13630
rlabel metal2 16 -1798 16 -1798 0 net=6483
rlabel metal2 121 -1798 121 -1798 0 net=7335
rlabel metal2 639 -1798 639 -1798 0 net=4597
rlabel metal2 730 -1798 730 -1798 0 net=9727
rlabel metal2 1409 -1798 1409 -1798 0 net=7329
rlabel metal2 37 -1800 37 -1800 0 net=3553
rlabel metal2 79 -1800 79 -1800 0 net=5423
rlabel metal2 131 -1800 131 -1800 0 net=2401
rlabel metal2 387 -1800 387 -1800 0 net=4291
rlabel metal2 660 -1800 660 -1800 0 net=6581
rlabel metal2 660 -1800 660 -1800 0 net=6581
rlabel metal2 681 -1800 681 -1800 0 net=7395
rlabel metal2 814 -1800 814 -1800 0 net=5959
rlabel metal2 954 -1800 954 -1800 0 net=6843
rlabel metal2 1059 -1800 1059 -1800 0 net=8874
rlabel metal2 1304 -1800 1304 -1800 0 net=12510
rlabel metal2 1850 -1800 1850 -1800 0 net=13263
rlabel metal2 1913 -1800 1913 -1800 0 net=13663
rlabel metal2 37 -1802 37 -1802 0 net=4875
rlabel metal2 156 -1802 156 -1802 0 net=1541
rlabel metal2 387 -1802 387 -1802 0 net=2063
rlabel metal2 562 -1802 562 -1802 0 net=3373
rlabel metal2 632 -1802 632 -1802 0 net=4259
rlabel metal2 684 -1802 684 -1802 0 net=1025
rlabel metal2 1010 -1802 1010 -1802 0 net=7093
rlabel metal2 1010 -1802 1010 -1802 0 net=7093
rlabel metal2 1017 -1802 1017 -1802 0 net=7153
rlabel metal2 1104 -1802 1104 -1802 0 net=9038
rlabel metal2 1244 -1802 1244 -1802 0 net=10968
rlabel metal2 1717 -1802 1717 -1802 0 net=12579
rlabel metal2 1815 -1802 1815 -1802 0 net=13041
rlabel metal2 1871 -1802 1871 -1802 0 net=13337
rlabel metal2 79 -1804 79 -1804 0 net=4655
rlabel metal2 765 -1804 765 -1804 0 net=5777
rlabel metal2 1073 -1804 1073 -1804 0 net=8581
rlabel metal2 1248 -1804 1248 -1804 0 net=9191
rlabel metal2 1304 -1804 1304 -1804 0 net=9251
rlabel metal2 1535 -1804 1535 -1804 0 net=10585
rlabel metal2 156 -1806 156 -1806 0 net=4015
rlabel metal2 415 -1806 415 -1806 0 net=4584
rlabel metal2 1108 -1806 1108 -1806 0 net=13585
rlabel metal2 170 -1808 170 -1808 0 net=2181
rlabel metal2 1111 -1808 1111 -1808 0 net=9296
rlabel metal2 1269 -1808 1269 -1808 0 net=9333
rlabel metal2 1360 -1808 1360 -1808 0 net=11862
rlabel metal2 1745 -1808 1745 -1808 0 net=13209
rlabel metal2 177 -1810 177 -1810 0 net=4321
rlabel metal2 401 -1810 401 -1810 0 net=8790
rlabel metal2 1129 -1810 1129 -1810 0 net=7571
rlabel metal2 1129 -1810 1129 -1810 0 net=7571
rlabel metal2 1136 -1810 1136 -1810 0 net=7807
rlabel metal2 1185 -1810 1185 -1810 0 net=8451
rlabel metal2 1262 -1810 1262 -1810 0 net=7183
rlabel metal2 1283 -1810 1283 -1810 0 net=9479
rlabel metal2 1363 -1810 1363 -1810 0 net=13287
rlabel metal2 177 -1812 177 -1812 0 net=8847
rlabel metal2 404 -1812 404 -1812 0 net=3491
rlabel metal2 429 -1812 429 -1812 0 net=2208
rlabel metal2 583 -1812 583 -1812 0 net=3841
rlabel metal2 1115 -1812 1115 -1812 0 net=7655
rlabel metal2 1150 -1812 1150 -1812 0 net=7999
rlabel metal2 1276 -1812 1276 -1812 0 net=8775
rlabel metal2 1307 -1812 1307 -1812 0 net=11932
rlabel metal2 1794 -1812 1794 -1812 0 net=12851
rlabel metal2 191 -1814 191 -1814 0 net=2577
rlabel metal2 240 -1814 240 -1814 0 net=2621
rlabel metal2 408 -1814 408 -1814 0 net=5783
rlabel metal2 1150 -1814 1150 -1814 0 net=9879
rlabel metal2 1535 -1814 1535 -1814 0 net=12825
rlabel metal2 1822 -1814 1822 -1814 0 net=13069
rlabel metal2 201 -1816 201 -1816 0 net=3012
rlabel metal2 380 -1816 380 -1816 0 net=4698
rlabel metal2 429 -1816 429 -1816 0 net=4231
rlabel metal2 604 -1816 604 -1816 0 net=5913
rlabel metal2 751 -1816 751 -1816 0 net=5219
rlabel metal2 1157 -1816 1157 -1816 0 net=8305
rlabel metal2 1311 -1816 1311 -1816 0 net=10401
rlabel metal2 1563 -1816 1563 -1816 0 net=10801
rlabel metal2 1577 -1816 1577 -1816 0 net=11993
rlabel metal2 1759 -1816 1759 -1816 0 net=12639
rlabel metal2 1801 -1816 1801 -1816 0 net=12939
rlabel metal2 187 -1818 187 -1818 0 net=12343
rlabel metal2 219 -1820 219 -1820 0 net=4423
rlabel metal2 450 -1820 450 -1820 0 net=5233
rlabel metal2 723 -1820 723 -1820 0 net=315
rlabel metal2 831 -1820 831 -1820 0 net=10081
rlabel metal2 1598 -1820 1598 -1820 0 net=10957
rlabel metal2 23 -1822 23 -1822 0 net=10427
rlabel metal2 863 -1822 863 -1822 0 net=6255
rlabel metal2 1318 -1822 1318 -1822 0 net=11510
rlabel metal2 1738 -1822 1738 -1822 0 net=11435
rlabel metal2 1766 -1822 1766 -1822 0 net=12769
rlabel metal2 23 -1824 23 -1824 0 net=6137
rlabel metal2 632 -1824 632 -1824 0 net=3537
rlabel metal2 765 -1824 765 -1824 0 net=6891
rlabel metal2 891 -1824 891 -1824 0 net=6571
rlabel metal2 975 -1824 975 -1824 0 net=6973
rlabel metal2 1164 -1824 1164 -1824 0 net=8339
rlabel metal2 1321 -1824 1321 -1824 0 net=11661
rlabel metal2 1654 -1824 1654 -1824 0 net=11831
rlabel metal2 72 -1826 72 -1826 0 net=5305
rlabel metal2 464 -1826 464 -1826 0 net=2788
rlabel metal2 541 -1826 541 -1826 0 net=3621
rlabel metal2 576 -1826 576 -1826 0 net=4545
rlabel metal2 768 -1826 768 -1826 0 net=9382
rlabel metal2 1486 -1826 1486 -1826 0 net=12295
rlabel metal2 44 -1828 44 -1828 0 net=2109
rlabel metal2 100 -1828 100 -1828 0 net=6735
rlabel metal2 1024 -1828 1024 -1828 0 net=8241
rlabel metal2 1178 -1828 1178 -1828 0 net=8679
rlabel metal2 1325 -1828 1325 -1828 0 net=9593
rlabel metal2 1409 -1828 1409 -1828 0 net=8199
rlabel metal2 1598 -1828 1598 -1828 0 net=12751
rlabel metal2 1696 -1828 1696 -1828 0 net=10777
rlabel metal2 30 -1830 30 -1830 0 net=4774
rlabel metal2 1083 -1830 1083 -1830 0 net=12003
rlabel metal2 30 -1832 30 -1832 0 net=2241
rlabel metal2 240 -1832 240 -1832 0 net=2879
rlabel metal2 373 -1832 373 -1832 0 net=3313
rlabel metal2 464 -1832 464 -1832 0 net=3947
rlabel metal2 772 -1832 772 -1832 0 net=7141
rlabel metal2 1143 -1832 1143 -1832 0 net=7943
rlabel metal2 1255 -1832 1255 -1832 0 net=9299
rlabel metal2 1339 -1832 1339 -1832 0 net=10527
rlabel metal2 1605 -1832 1605 -1832 0 net=11179
rlabel metal2 1661 -1832 1661 -1832 0 net=13095
rlabel metal2 44 -1834 44 -1834 0 net=2971
rlabel metal2 436 -1834 436 -1834 0 net=3157
rlabel metal2 772 -1834 772 -1834 0 net=7320
rlabel metal2 1122 -1834 1122 -1834 0 net=7661
rlabel metal2 1199 -1834 1199 -1834 0 net=8473
rlabel metal2 1430 -1834 1430 -1834 0 net=9997
rlabel metal2 1808 -1834 1808 -1834 0 net=13021
rlabel metal2 184 -1836 184 -1836 0 net=9267
rlabel metal2 1451 -1836 1451 -1836 0 net=10231
rlabel metal2 1479 -1836 1479 -1836 0 net=10315
rlabel metal2 1633 -1836 1633 -1836 0 net=10381
rlabel metal2 1682 -1836 1682 -1836 0 net=11793
rlabel metal2 1710 -1836 1710 -1836 0 net=12373
rlabel metal2 163 -1838 163 -1838 0 net=2633
rlabel metal2 205 -1838 205 -1838 0 net=3083
rlabel metal2 380 -1838 380 -1838 0 net=3603
rlabel metal2 485 -1838 485 -1838 0 net=4483
rlabel metal2 558 -1838 558 -1838 0 net=9617
rlabel metal2 1234 -1838 1234 -1838 0 net=9369
rlabel metal2 1367 -1838 1367 -1838 0 net=10253
rlabel metal2 1542 -1838 1542 -1838 0 net=10731
rlabel metal2 163 -1840 163 -1840 0 net=8583
rlabel metal2 520 -1840 520 -1840 0 net=6759
rlabel metal2 891 -1840 891 -1840 0 net=5357
rlabel metal2 1367 -1840 1367 -1840 0 net=9671
rlabel metal2 1388 -1840 1388 -1840 0 net=10105
rlabel metal2 1556 -1840 1556 -1840 0 net=10771
rlabel metal2 1668 -1840 1668 -1840 0 net=11571
rlabel metal2 205 -1842 205 -1842 0 net=1943
rlabel metal2 261 -1842 261 -1842 0 net=3265
rlabel metal2 478 -1842 478 -1842 0 net=10561
rlabel metal2 1556 -1842 1556 -1842 0 net=10661
rlabel metal2 149 -1844 149 -1844 0 net=3423
rlabel metal2 296 -1844 296 -1844 0 net=1551
rlabel metal2 485 -1844 485 -1844 0 net=12739
rlabel metal2 149 -1846 149 -1846 0 net=2287
rlabel metal2 912 -1846 912 -1846 0 net=6437
rlabel metal2 933 -1846 933 -1846 0 net=12017
rlabel metal2 226 -1848 226 -1848 0 net=2385
rlabel metal2 492 -1848 492 -1848 0 net=5348
rlabel metal2 912 -1848 912 -1848 0 net=6831
rlabel metal2 996 -1848 996 -1848 0 net=7031
rlabel metal2 1045 -1848 1045 -1848 0 net=10035
rlabel metal2 1647 -1848 1647 -1848 0 net=11397
rlabel metal2 233 -1850 233 -1850 0 net=2305
rlabel metal2 331 -1850 331 -1850 0 net=3767
rlabel metal2 492 -1850 492 -1850 0 net=4355
rlabel metal2 779 -1850 779 -1850 0 net=7087
rlabel metal2 1031 -1850 1031 -1850 0 net=7285
rlabel metal2 1122 -1850 1122 -1850 0 net=13166
rlabel metal2 86 -1852 86 -1852 0 net=3961
rlabel metal2 324 -1852 324 -1852 0 net=2885
rlabel metal2 513 -1852 513 -1852 0 net=3779
rlabel metal2 1220 -1852 1220 -1852 0 net=8397
rlabel metal2 1241 -1852 1241 -1852 0 net=9853
rlabel metal2 1612 -1852 1612 -1852 0 net=11221
rlabel metal2 86 -1854 86 -1854 0 net=4641
rlabel metal2 1374 -1854 1374 -1854 0 net=9755
rlabel metal2 1423 -1854 1423 -1854 0 net=9971
rlabel metal2 247 -1856 247 -1856 0 net=3331
rlabel metal2 530 -1856 530 -1856 0 net=1
rlabel metal2 1346 -1856 1346 -1856 0 net=9659
rlabel metal2 1416 -1856 1416 -1856 0 net=9925
rlabel metal2 1465 -1856 1465 -1856 0 net=10719
rlabel metal2 247 -1858 247 -1858 0 net=4059
rlabel metal2 317 -1860 317 -1860 0 net=1733
rlabel metal2 579 -1860 579 -1860 0 net=10647
rlabel metal2 317 -1862 317 -1862 0 net=2981
rlabel metal2 611 -1862 611 -1862 0 net=11065
rlabel metal2 198 -1864 198 -1864 0 net=4139
rlabel metal2 618 -1864 618 -1864 0 net=9162
rlabel metal2 905 -1864 905 -1864 0 net=6643
rlabel metal2 1031 -1864 1031 -1864 0 net=7685
rlabel metal2 1111 -1864 1111 -1864 0 net=13051
rlabel metal2 422 -1866 422 -1866 0 net=3673
rlabel metal2 954 -1866 954 -1866 0 net=4955
rlabel metal2 1297 -1866 1297 -1866 0 net=9385
rlabel metal2 1388 -1866 1388 -1866 0 net=9769
rlabel metal2 1416 -1866 1416 -1866 0 net=9881
rlabel metal2 779 -1868 779 -1868 0 net=6211
rlabel metal2 1052 -1868 1052 -1868 0 net=7485
rlabel metal2 1227 -1868 1227 -1868 0 net=8845
rlabel metal2 1332 -1868 1332 -1868 0 net=9863
rlabel metal2 1528 -1868 1528 -1868 0 net=10863
rlabel metal2 1857 -1868 1857 -1868 0 net=13309
rlabel metal2 61 -1870 61 -1870 0 net=8371
rlabel metal2 1507 -1870 1507 -1870 0 net=10899
rlabel metal2 68 -1872 68 -1872 0 net=10347
rlabel metal2 103 -1874 103 -1874 0 net=5843
rlabel metal2 989 -1874 989 -1874 0 net=7007
rlabel metal2 1507 -1874 1507 -1874 0 net=10455
rlabel metal2 534 -1876 534 -1876 0 net=4049
rlabel metal2 1472 -1876 1472 -1876 0 net=10295
rlabel metal2 534 -1878 534 -1878 0 net=5979
rlabel metal2 786 -1878 786 -1878 0 net=6111
rlabel metal2 1472 -1878 1472 -1878 0 net=11689
rlabel metal2 674 -1880 674 -1880 0 net=7415
rlabel metal2 1675 -1880 1675 -1880 0 net=12589
rlabel metal2 418 -1882 418 -1882 0 net=11871
rlabel metal2 674 -1884 674 -1884 0 net=4673
rlabel metal2 737 -1884 737 -1884 0 net=9259
rlabel metal2 565 -1886 565 -1886 0 net=4705
rlabel metal2 758 -1886 758 -1886 0 net=5681
rlabel metal2 646 -1888 646 -1888 0 net=4717
rlabel metal2 821 -1888 821 -1888 0 net=5155
rlabel metal2 569 -1890 569 -1890 0 net=1809
rlabel metal2 800 -1890 800 -1890 0 net=5541
rlabel metal2 471 -1892 471 -1892 0 net=4197
rlabel metal2 716 -1892 716 -1892 0 net=7221
rlabel metal2 471 -1894 471 -1894 0 net=1679
rlabel metal2 716 -1896 716 -1896 0 net=9203
rlabel metal2 1563 -1896 1563 -1896 0 net=13389
rlabel metal2 2 -1907 2 -1907 0 net=2387
rlabel metal2 313 -1907 313 -1907 0 net=5306
rlabel metal2 478 -1907 478 -1907 0 net=2835
rlabel metal2 562 -1907 562 -1907 0 net=3375
rlabel metal2 614 -1907 614 -1907 0 net=4050
rlabel metal2 1024 -1907 1024 -1907 0 net=9594
rlabel metal2 1430 -1907 1430 -1907 0 net=10037
rlabel metal2 1430 -1907 1430 -1907 0 net=10037
rlabel metal2 1454 -1907 1454 -1907 0 net=12852
rlabel metal2 5 -1909 5 -1909 0 net=484
rlabel metal2 79 -1909 79 -1909 0 net=4656
rlabel metal2 537 -1909 537 -1909 0 net=3584
rlabel metal2 1153 -1909 1153 -1909 0 net=12374
rlabel metal2 1871 -1909 1871 -1909 0 net=13211
rlabel metal2 9 -1911 9 -1911 0 net=4877
rlabel metal2 44 -1911 44 -1911 0 net=2972
rlabel metal2 142 -1911 142 -1911 0 net=9880
rlabel metal2 1458 -1911 1458 -1911 0 net=10233
rlabel metal2 1458 -1911 1458 -1911 0 net=10233
rlabel metal2 1535 -1911 1535 -1911 0 net=12827
rlabel metal2 1899 -1911 1899 -1911 0 net=13391
rlabel metal2 37 -1913 37 -1913 0 net=4485
rlabel metal2 555 -1913 555 -1913 0 net=4719
rlabel metal2 744 -1913 744 -1913 0 net=4863
rlabel metal2 1108 -1913 1108 -1913 0 net=8846
rlabel metal2 1367 -1913 1367 -1913 0 net=9673
rlabel metal2 1444 -1913 1444 -1913 0 net=10107
rlabel metal2 1535 -1913 1535 -1913 0 net=10627
rlabel metal2 44 -1915 44 -1915 0 net=1911
rlabel metal2 317 -1915 317 -1915 0 net=2983
rlabel metal2 828 -1915 828 -1915 0 net=10428
rlabel metal2 947 -1915 947 -1915 0 net=6715
rlabel metal2 947 -1915 947 -1915 0 net=6715
rlabel metal2 964 -1915 964 -1915 0 net=6256
rlabel metal2 1451 -1915 1451 -1915 0 net=10864
rlabel metal2 1563 -1915 1563 -1915 0 net=10803
rlabel metal2 1745 -1915 1745 -1915 0 net=11995
rlabel metal2 1745 -1915 1745 -1915 0 net=11995
rlabel metal2 1948 -1915 1948 -1915 0 net=13587
rlabel metal2 58 -1917 58 -1917 0 net=5235
rlabel metal2 716 -1917 716 -1917 0 net=5025
rlabel metal2 772 -1917 772 -1917 0 net=12193
rlabel metal2 1976 -1917 1976 -1917 0 net=2617
rlabel metal2 79 -1919 79 -1919 0 net=1681
rlabel metal2 481 -1919 481 -1919 0 net=9854
rlabel metal2 1283 -1919 1283 -1919 0 net=8777
rlabel metal2 1528 -1919 1528 -1919 0 net=12005
rlabel metal2 23 -1921 23 -1921 0 net=6139
rlabel metal2 485 -1921 485 -1921 0 net=1338
rlabel metal2 919 -1921 919 -1921 0 net=6439
rlabel metal2 982 -1921 982 -1921 0 net=10772
rlabel metal2 23 -1923 23 -1923 0 net=2515
rlabel metal2 128 -1923 128 -1923 0 net=1853
rlabel metal2 128 -1923 128 -1923 0 net=1853
rlabel metal2 135 -1923 135 -1923 0 net=1376
rlabel metal2 730 -1923 730 -1923 0 net=9728
rlabel metal2 905 -1923 905 -1923 0 net=10958
rlabel metal2 86 -1925 86 -1925 0 net=4643
rlabel metal2 317 -1925 317 -1925 0 net=5683
rlabel metal2 779 -1925 779 -1925 0 net=6213
rlabel metal2 982 -1925 982 -1925 0 net=7657
rlabel metal2 1143 -1925 1143 -1925 0 net=7663
rlabel metal2 1293 -1925 1293 -1925 0 net=10586
rlabel metal2 100 -1927 100 -1927 0 net=3962
rlabel metal2 338 -1927 338 -1927 0 net=5755
rlabel metal2 845 -1927 845 -1927 0 net=6974
rlabel metal2 1199 -1927 1199 -1927 0 net=9619
rlabel metal2 1566 -1927 1566 -1927 0 net=10830
rlabel metal2 1633 -1927 1633 -1927 0 net=10383
rlabel metal2 1815 -1927 1815 -1927 0 net=12941
rlabel metal2 1843 -1927 1843 -1927 0 net=13075
rlabel metal2 100 -1929 100 -1929 0 net=2661
rlabel metal2 562 -1929 562 -1929 0 net=3843
rlabel metal2 632 -1929 632 -1929 0 net=3538
rlabel metal2 779 -1929 779 -1929 0 net=5845
rlabel metal2 880 -1929 880 -1929 0 net=6844
rlabel metal2 1090 -1929 1090 -1929 0 net=7330
rlabel metal2 30 -1931 30 -1931 0 net=2242
rlabel metal2 583 -1931 583 -1931 0 net=5517
rlabel metal2 660 -1931 660 -1931 0 net=6583
rlabel metal2 688 -1931 688 -1931 0 net=9660
rlabel metal2 1472 -1931 1472 -1931 0 net=11691
rlabel metal2 1822 -1931 1822 -1931 0 net=13023
rlabel metal2 1885 -1931 1885 -1931 0 net=13289
rlabel metal2 1990 -1931 1990 -1931 0 net=8177
rlabel metal2 30 -1933 30 -1933 0 net=3781
rlabel metal2 660 -1933 660 -1933 0 net=4547
rlabel metal2 681 -1933 681 -1933 0 net=4261
rlabel metal2 698 -1933 698 -1933 0 net=8967
rlabel metal2 1297 -1933 1297 -1933 0 net=10403
rlabel metal2 1584 -1933 1584 -1933 0 net=11067
rlabel metal2 1836 -1933 1836 -1933 0 net=13043
rlabel metal2 1927 -1933 1927 -1933 0 net=13485
rlabel metal2 16 -1935 16 -1935 0 net=6485
rlabel metal2 674 -1935 674 -1935 0 net=4675
rlabel metal2 709 -1935 709 -1935 0 net=4707
rlabel metal2 719 -1935 719 -1935 0 net=5960
rlabel metal2 856 -1935 856 -1935 0 net=7513
rlabel metal2 1094 -1935 1094 -1935 0 net=7155
rlabel metal2 1129 -1935 1129 -1935 0 net=7573
rlabel metal2 1157 -1935 1157 -1935 0 net=7809
rlabel metal2 1206 -1935 1206 -1935 0 net=10695
rlabel metal2 1220 -1935 1220 -1935 0 net=9998
rlabel metal2 1955 -1935 1955 -1935 0 net=13607
rlabel metal2 65 -1937 65 -1937 0 net=3891
rlabel metal2 674 -1937 674 -1937 0 net=4599
rlabel metal2 709 -1937 709 -1937 0 net=2807
rlabel metal2 1066 -1937 1066 -1937 0 net=7487
rlabel metal2 1094 -1937 1094 -1937 0 net=9269
rlabel metal2 1395 -1937 1395 -1937 0 net=10417
rlabel metal2 1661 -1937 1661 -1937 0 net=13097
rlabel metal2 103 -1939 103 -1939 0 net=6736
rlabel metal2 989 -1939 989 -1939 0 net=7687
rlabel metal2 1052 -1939 1052 -1939 0 net=7009
rlabel metal2 1108 -1939 1108 -1939 0 net=10296
rlabel metal2 16 -1941 16 -1941 0 net=6801
rlabel metal2 1136 -1941 1136 -1941 0 net=7945
rlabel metal2 1206 -1941 1206 -1941 0 net=10549
rlabel metal2 107 -1943 107 -1943 0 net=5186
rlabel metal2 135 -1943 135 -1943 0 net=2065
rlabel metal2 401 -1943 401 -1943 0 net=5037
rlabel metal2 1213 -1943 1213 -1943 0 net=8341
rlabel metal2 1213 -1943 1213 -1943 0 net=8341
rlabel metal2 1220 -1943 1220 -1943 0 net=9883
rlabel metal2 1472 -1943 1472 -1943 0 net=10563
rlabel metal2 93 -1945 93 -1945 0 net=2099
rlabel metal2 415 -1945 415 -1945 0 net=3493
rlabel metal2 639 -1945 639 -1945 0 net=4293
rlabel metal2 730 -1945 730 -1945 0 net=12854
rlabel metal2 51 -1947 51 -1947 0 net=3555
rlabel metal2 107 -1947 107 -1947 0 net=3359
rlabel metal2 1003 -1947 1003 -1947 0 net=7089
rlabel metal2 1164 -1947 1164 -1947 0 net=8243
rlabel metal2 1223 -1947 1223 -1947 0 net=13664
rlabel metal2 51 -1949 51 -1949 0 net=3521
rlabel metal2 733 -1949 733 -1949 0 net=12501
rlabel metal2 1878 -1949 1878 -1949 0 net=13265
rlabel metal2 1920 -1949 1920 -1949 0 net=10338
rlabel metal2 142 -1951 142 -1951 0 net=12612
rlabel metal2 1906 -1951 1906 -1951 0 net=13311
rlabel metal2 145 -1953 145 -1953 0 net=2880
rlabel metal2 408 -1953 408 -1953 0 net=5785
rlabel metal2 464 -1953 464 -1953 0 net=3949
rlabel metal2 758 -1953 758 -1953 0 net=6644
rlabel metal2 1010 -1953 1010 -1953 0 net=7095
rlabel metal2 1027 -1953 1027 -1953 0 net=12344
rlabel metal2 1934 -1953 1934 -1953 0 net=13509
rlabel metal2 86 -1955 86 -1955 0 net=6149
rlabel metal2 156 -1955 156 -1955 0 net=4017
rlabel metal2 156 -1955 156 -1955 0 net=4017
rlabel metal2 198 -1955 198 -1955 0 net=3424
rlabel metal2 408 -1955 408 -1955 0 net=5221
rlabel metal2 800 -1955 800 -1955 0 net=7223
rlabel metal2 1164 -1955 1164 -1955 0 net=8453
rlabel metal2 1262 -1955 1262 -1955 0 net=8681
rlabel metal2 1521 -1955 1521 -1955 0 net=10649
rlabel metal2 1787 -1955 1787 -1955 0 net=12741
rlabel metal2 170 -1957 170 -1957 0 net=2183
rlabel metal2 464 -1957 464 -1957 0 net=2735
rlabel metal2 807 -1957 807 -1957 0 net=8099
rlabel metal2 1171 -1957 1171 -1957 0 net=8475
rlabel metal2 1265 -1957 1265 -1957 0 net=12381
rlabel metal2 1794 -1957 1794 -1957 0 net=12771
rlabel metal2 170 -1959 170 -1959 0 net=3131
rlabel metal2 807 -1959 807 -1959 0 net=5543
rlabel metal2 849 -1959 849 -1959 0 net=7417
rlabel metal2 1178 -1959 1178 -1959 0 net=8001
rlabel metal2 1216 -1959 1216 -1959 0 net=1
rlabel metal2 1598 -1959 1598 -1959 0 net=12753
rlabel metal2 198 -1961 198 -1961 0 net=2461
rlabel metal2 1290 -1961 1290 -1961 0 net=9193
rlabel metal2 1416 -1961 1416 -1961 0 net=9927
rlabel metal2 1479 -1961 1479 -1961 0 net=10255
rlabel metal2 1542 -1961 1542 -1961 0 net=10663
rlabel metal2 212 -1963 212 -1963 0 net=6882
rlabel metal2 268 -1963 268 -1963 0 net=3395
rlabel metal2 1409 -1963 1409 -1963 0 net=8201
rlabel metal2 1465 -1963 1465 -1963 0 net=10721
rlabel metal2 184 -1965 184 -1965 0 net=2635
rlabel metal2 226 -1965 226 -1965 0 net=2025
rlabel metal2 485 -1965 485 -1965 0 net=3159
rlabel metal2 814 -1965 814 -1965 0 net=9260
rlabel metal2 1388 -1965 1388 -1965 0 net=9771
rlabel metal2 1486 -1965 1486 -1965 0 net=10317
rlabel metal2 1507 -1965 1507 -1965 0 net=10457
rlabel metal2 184 -1967 184 -1967 0 net=2579
rlabel metal2 205 -1967 205 -1967 0 net=1945
rlabel metal2 457 -1967 457 -1967 0 net=4141
rlabel metal2 821 -1967 821 -1967 0 net=5157
rlabel metal2 849 -1967 849 -1967 0 net=8582
rlabel metal2 1087 -1967 1087 -1967 0 net=10355
rlabel metal2 1486 -1967 1486 -1967 0 net=11223
rlabel metal2 163 -1969 163 -1969 0 net=8585
rlabel metal2 205 -1969 205 -1969 0 net=3539
rlabel metal2 618 -1969 618 -1969 0 net=548
rlabel metal2 793 -1969 793 -1969 0 net=7397
rlabel metal2 1087 -1969 1087 -1969 0 net=9334
rlabel metal2 1360 -1969 1360 -1969 0 net=9481
rlabel metal2 1647 -1969 1647 -1969 0 net=11653
rlabel metal2 72 -1971 72 -1971 0 net=2111
rlabel metal2 341 -1971 341 -1971 0 net=5123
rlabel metal2 793 -1971 793 -1971 0 net=4957
rlabel metal2 961 -1971 961 -1971 0 net=12681
rlabel metal2 61 -1973 61 -1973 0 net=6091
rlabel metal2 380 -1973 380 -1973 0 net=3605
rlabel metal2 499 -1973 499 -1973 0 net=3745
rlabel metal2 821 -1973 821 -1973 0 net=8307
rlabel metal2 1227 -1973 1227 -1973 0 net=8373
rlabel metal2 1227 -1973 1227 -1973 0 net=8373
rlabel metal2 1237 -1973 1237 -1973 0 net=15
rlabel metal2 1325 -1973 1325 -1973 0 net=9301
rlabel metal2 1374 -1973 1374 -1973 0 net=9757
rlabel metal2 1689 -1973 1689 -1973 0 net=12019
rlabel metal2 380 -1975 380 -1975 0 net=3769
rlabel metal2 443 -1975 443 -1975 0 net=3315
rlabel metal2 506 -1975 506 -1975 0 net=8479
rlabel metal2 1269 -1975 1269 -1975 0 net=7185
rlabel metal2 247 -1977 247 -1977 0 net=4061
rlabel metal2 754 -1977 754 -1977 0 net=8737
rlabel metal2 1276 -1977 1276 -1977 0 net=11325
rlabel metal2 177 -1979 177 -1979 0 net=8849
rlabel metal2 1304 -1979 1304 -1979 0 net=9253
rlabel metal2 1339 -1979 1339 -1979 0 net=9371
rlabel metal2 177 -1981 177 -1981 0 net=2403
rlabel metal2 863 -1981 863 -1981 0 net=6893
rlabel metal2 1150 -1981 1150 -1981 0 net=12527
rlabel metal2 247 -1983 247 -1983 0 net=1735
rlabel metal2 352 -1983 352 -1983 0 net=2949
rlabel metal2 611 -1983 611 -1983 0 net=6883
rlabel metal2 1192 -1983 1192 -1983 0 net=13070
rlabel metal2 254 -1985 254 -1985 0 net=2497
rlabel metal2 611 -1985 611 -1985 0 net=8533
rlabel metal2 863 -1985 863 -1985 0 net=13710
rlabel metal2 254 -1987 254 -1987 0 net=5021
rlabel metal2 324 -1987 324 -1987 0 net=3675
rlabel metal2 866 -1987 866 -1987 0 net=13665
rlabel metal2 275 -1989 275 -1989 0 net=4323
rlabel metal2 877 -1989 877 -1989 0 net=6849
rlabel metal2 996 -1989 996 -1989 0 net=7033
rlabel metal2 1255 -1989 1255 -1989 0 net=13417
rlabel metal2 275 -1991 275 -1991 0 net=5877
rlabel metal2 877 -1991 877 -1991 0 net=10528
rlabel metal2 296 -1993 296 -1993 0 net=1552
rlabel metal2 345 -1993 345 -1993 0 net=3333
rlabel metal2 842 -1993 842 -1993 0 net=5779
rlabel metal2 884 -1993 884 -1993 0 net=9972
rlabel metal2 121 -1995 121 -1995 0 net=5425
rlabel metal2 345 -1995 345 -1995 0 net=4023
rlabel metal2 604 -1995 604 -1995 0 net=5915
rlabel metal2 887 -1995 887 -1995 0 net=2959
rlabel metal2 121 -1997 121 -1997 0 net=4233
rlabel metal2 604 -1997 604 -1997 0 net=7287
rlabel metal2 1339 -1997 1339 -1997 0 net=9387
rlabel metal2 1577 -1997 1577 -1997 0 net=10901
rlabel metal2 1612 -1997 1612 -1997 0 net=12591
rlabel metal2 219 -1999 219 -1999 0 net=4425
rlabel metal2 842 -1999 842 -1999 0 net=10732
rlabel metal2 219 -2001 219 -2001 0 net=5980
rlabel metal2 912 -2001 912 -2001 0 net=6833
rlabel metal2 968 -2001 968 -2001 0 net=6871
rlabel metal2 1017 -2001 1017 -2001 0 net=7143
rlabel metal2 1111 -2001 1111 -2001 0 net=12065
rlabel metal2 352 -2003 352 -2003 0 net=4199
rlabel metal2 800 -2003 800 -2003 0 net=3043
rlabel metal2 1017 -2003 1017 -2003 0 net=10083
rlabel metal2 1591 -2003 1591 -2003 0 net=11399
rlabel metal2 1675 -2003 1675 -2003 0 net=10779
rlabel metal2 492 -2005 492 -2005 0 net=4357
rlabel metal2 912 -2005 912 -2005 0 net=4979
rlabel metal2 1111 -2005 1111 -2005 0 net=9393
rlabel metal2 1402 -2005 1402 -2005 0 net=9865
rlabel metal2 1668 -2005 1668 -2005 0 net=11795
rlabel metal2 1703 -2005 1703 -2005 0 net=11437
rlabel metal2 359 -2007 359 -2007 0 net=3267
rlabel metal2 520 -2007 520 -2007 0 net=6760
rlabel metal2 723 -2007 723 -2007 0 net=9527
rlabel metal2 1640 -2007 1640 -2007 0 net=11181
rlabel metal2 331 -2009 331 -2009 0 net=2887
rlabel metal2 394 -2009 394 -2009 0 net=2623
rlabel metal2 530 -2009 530 -2009 0 net=12415
rlabel metal2 149 -2011 149 -2011 0 net=2289
rlabel metal2 723 -2011 723 -2011 0 net=11739
rlabel metal2 149 -2013 149 -2013 0 net=3461
rlabel metal2 233 -2013 233 -2013 0 net=2307
rlabel metal2 919 -2013 919 -2013 0 net=8989
rlabel metal2 1640 -2013 1640 -2013 0 net=11573
rlabel metal2 233 -2015 233 -2015 0 net=1543
rlabel metal2 922 -2015 922 -2015 0 net=11489
rlabel metal2 1682 -2015 1682 -2015 0 net=11873
rlabel metal2 282 -2017 282 -2017 0 net=3085
rlabel metal2 926 -2017 926 -2017 0 net=9205
rlabel metal2 1234 -2017 1234 -2017 0 net=8399
rlabel metal2 1724 -2017 1724 -2017 0 net=12297
rlabel metal2 373 -2019 373 -2019 0 net=5163
rlabel metal2 1766 -2019 1766 -2019 0 net=12581
rlabel metal2 898 -2021 898 -2021 0 net=7423
rlabel metal2 940 -2021 940 -2021 0 net=6573
rlabel metal2 1773 -2021 1773 -2021 0 net=12641
rlabel metal2 625 -2023 625 -2023 0 net=7337
rlabel metal2 1619 -2023 1619 -2023 0 net=11319
rlabel metal2 548 -2025 548 -2025 0 net=3623
rlabel metal2 786 -2025 786 -2025 0 net=6113
rlabel metal2 1619 -2025 1619 -2025 0 net=11833
rlabel metal2 548 -2027 548 -2027 0 net=1811
rlabel metal2 772 -2027 772 -2027 0 net=3829
rlabel metal2 1626 -2027 1626 -2027 0 net=11663
rlabel metal2 590 -2029 590 -2029 0 net=3975
rlabel metal2 1626 -2029 1626 -2029 0 net=13053
rlabel metal2 590 -2031 590 -2031 0 net=3715
rlabel metal2 1104 -2031 1104 -2031 0 net=13153
rlabel metal2 765 -2033 765 -2033 0 net=5359
rlabel metal2 891 -2035 891 -2035 0 net=10348
rlabel metal2 1857 -2037 1857 -2037 0 net=13149
rlabel metal2 1892 -2039 1892 -2039 0 net=13339
rlabel metal2 1941 -2041 1941 -2041 0 net=13519
rlabel metal2 761 -2043 761 -2043 0 net=13681
rlabel metal2 2 -2054 2 -2054 0 net=2388
rlabel metal2 352 -2054 352 -2054 0 net=4200
rlabel metal2 733 -2054 733 -2054 0 net=4864
rlabel metal2 1108 -2054 1108 -2054 0 net=10256
rlabel metal2 1920 -2054 1920 -2054 0 net=2618
rlabel metal2 2 -2056 2 -2056 0 net=3541
rlabel metal2 219 -2056 219 -2056 0 net=367
rlabel metal2 548 -2056 548 -2056 0 net=1812
rlabel metal2 817 -2056 817 -2056 0 net=7658
rlabel metal2 1087 -2056 1087 -2056 0 net=9271
rlabel metal2 1237 -2056 1237 -2056 0 net=10318
rlabel metal2 23 -2058 23 -2058 0 net=2516
rlabel metal2 149 -2058 149 -2058 0 net=3463
rlabel metal2 222 -2058 222 -2058 0 net=4294
rlabel metal2 723 -2058 723 -2058 0 net=7424
rlabel metal2 947 -2058 947 -2058 0 net=6717
rlabel metal2 947 -2058 947 -2058 0 net=6717
rlabel metal2 961 -2058 961 -2058 0 net=8682
rlabel metal2 9 -2060 9 -2060 0 net=4879
rlabel metal2 177 -2060 177 -2060 0 net=2405
rlabel metal2 352 -2060 352 -2060 0 net=2309
rlabel metal2 401 -2060 401 -2060 0 net=5039
rlabel metal2 723 -2060 723 -2060 0 net=6873
rlabel metal2 1087 -2060 1087 -2060 0 net=9207
rlabel metal2 1241 -2060 1241 -2060 0 net=7664
rlabel metal2 1265 -2060 1265 -2060 0 net=13098
rlabel metal2 23 -2062 23 -2062 0 net=9107
rlabel metal2 117 -2062 117 -2062 0 net=9482
rlabel metal2 1850 -2062 1850 -2062 0 net=13487
rlabel metal2 30 -2064 30 -2064 0 net=3782
rlabel metal2 394 -2064 394 -2064 0 net=2809
rlabel metal2 751 -2064 751 -2064 0 net=7418
rlabel metal2 1139 -2064 1139 -2064 0 net=9866
rlabel metal2 1493 -2064 1493 -2064 0 net=11491
rlabel metal2 30 -2066 30 -2066 0 net=483
rlabel metal2 520 -2066 520 -2066 0 net=2624
rlabel metal2 695 -2066 695 -2066 0 net=8100
rlabel metal2 1101 -2066 1101 -2066 0 net=8003
rlabel metal2 1241 -2066 1241 -2066 0 net=8991
rlabel metal2 1360 -2066 1360 -2066 0 net=7186
rlabel metal2 1500 -2066 1500 -2066 0 net=12529
rlabel metal2 37 -2068 37 -2068 0 net=4486
rlabel metal2 450 -2068 450 -2068 0 net=3316
rlabel metal2 530 -2068 530 -2068 0 net=9528
rlabel metal2 1437 -2068 1437 -2068 0 net=10565
rlabel metal2 1507 -2068 1507 -2068 0 net=12067
rlabel metal2 1759 -2068 1759 -2068 0 net=13151
rlabel metal2 51 -2070 51 -2070 0 net=3522
rlabel metal2 751 -2070 751 -2070 0 net=7971
rlabel metal2 1129 -2070 1129 -2070 0 net=7947
rlabel metal2 1143 -2070 1143 -2070 0 net=7575
rlabel metal2 1290 -2070 1290 -2070 0 net=9395
rlabel metal2 1363 -2070 1363 -2070 0 net=12742
rlabel metal2 1857 -2070 1857 -2070 0 net=13521
rlabel metal2 51 -2072 51 -2072 0 net=2185
rlabel metal2 303 -2072 303 -2072 0 net=1946
rlabel metal2 408 -2072 408 -2072 0 net=5222
rlabel metal2 845 -2072 845 -2072 0 net=11203
rlabel metal2 1605 -2072 1605 -2072 0 net=12643
rlabel metal2 1829 -2072 1829 -2072 0 net=13393
rlabel metal2 65 -2074 65 -2074 0 net=446
rlabel metal2 1710 -2074 1710 -2074 0 net=13045
rlabel metal2 1899 -2074 1899 -2074 0 net=8179
rlabel metal2 65 -2076 65 -2076 0 net=3771
rlabel metal2 415 -2076 415 -2076 0 net=5786
rlabel metal2 761 -2076 761 -2076 0 net=3830
rlabel metal2 807 -2076 807 -2076 0 net=5545
rlabel metal2 891 -2076 891 -2076 0 net=6802
rlabel metal2 1038 -2076 1038 -2076 0 net=7225
rlabel metal2 1143 -2076 1143 -2076 0 net=8343
rlabel metal2 1255 -2076 1255 -2076 0 net=8778
rlabel metal2 1353 -2076 1353 -2076 0 net=12195
rlabel metal2 1773 -2076 1773 -2076 0 net=13077
rlabel metal2 44 -2078 44 -2078 0 net=1913
rlabel metal2 422 -2078 422 -2078 0 net=3335
rlabel metal2 492 -2078 492 -2078 0 net=3269
rlabel metal2 548 -2078 548 -2078 0 net=3845
rlabel metal2 583 -2078 583 -2078 0 net=5519
rlabel metal2 919 -2078 919 -2078 0 net=10458
rlabel metal2 1843 -2078 1843 -2078 0 net=13419
rlabel metal2 44 -2080 44 -2080 0 net=6151
rlabel metal2 89 -2080 89 -2080 0 net=3676
rlabel metal2 422 -2080 422 -2080 0 net=6851
rlabel metal2 978 -2080 978 -2080 0 net=9372
rlabel metal2 1475 -2080 1475 -2080 0 net=13405
rlabel metal2 68 -2082 68 -2082 0 net=6140
rlabel metal2 492 -2082 492 -2082 0 net=3495
rlabel metal2 562 -2082 562 -2082 0 net=3951
rlabel metal2 1160 -2082 1160 -2082 0 net=9463
rlabel metal2 1311 -2082 1311 -2082 0 net=9759
rlabel metal2 1570 -2082 1570 -2082 0 net=11741
rlabel metal2 1717 -2082 1717 -2082 0 net=11665
rlabel metal2 79 -2084 79 -2084 0 net=1683
rlabel metal2 86 -2084 86 -2084 0 net=6486
rlabel metal2 583 -2084 583 -2084 0 net=3977
rlabel metal2 695 -2084 695 -2084 0 net=4709
rlabel metal2 730 -2084 730 -2084 0 net=5103
rlabel metal2 968 -2084 968 -2084 0 net=11326
rlabel metal2 1661 -2084 1661 -2084 0 net=12299
rlabel metal2 79 -2086 79 -2086 0 net=2067
rlabel metal2 163 -2086 163 -2086 0 net=2113
rlabel metal2 436 -2086 436 -2086 0 net=4063
rlabel metal2 590 -2086 590 -2086 0 net=3716
rlabel metal2 1479 -2086 1479 -2086 0 net=11069
rlabel metal2 1633 -2086 1633 -2086 0 net=10385
rlabel metal2 93 -2088 93 -2088 0 net=3557
rlabel metal2 593 -2088 593 -2088 0 net=2984
rlabel metal2 772 -2088 772 -2088 0 net=7090
rlabel metal2 1171 -2088 1171 -2088 0 net=8477
rlabel metal2 1213 -2088 1213 -2088 0 net=9389
rlabel metal2 1374 -2088 1374 -2088 0 net=13312
rlabel metal2 33 -2090 33 -2090 0 net=9561
rlabel metal2 772 -2090 772 -2090 0 net=4941
rlabel metal2 1171 -2090 1171 -2090 0 net=8401
rlabel metal2 1388 -2090 1388 -2090 0 net=10235
rlabel metal2 1584 -2090 1584 -2090 0 net=11797
rlabel metal2 1675 -2090 1675 -2090 0 net=10781
rlabel metal2 93 -2092 93 -2092 0 net=2100
rlabel metal2 467 -2092 467 -2092 0 net=11
rlabel metal2 971 -2092 971 -2092 0 net=8202
rlabel metal2 1458 -2092 1458 -2092 0 net=10665
rlabel metal2 1675 -2092 1675 -2092 0 net=12383
rlabel metal2 96 -2094 96 -2094 0 net=1245
rlabel metal2 597 -2094 597 -2094 0 net=3746
rlabel metal2 852 -2094 852 -2094 0 net=12131
rlabel metal2 1703 -2094 1703 -2094 0 net=11439
rlabel metal2 16 -2096 16 -2096 0 net=5575
rlabel metal2 905 -2096 905 -2096 0 net=6215
rlabel metal2 922 -2096 922 -2096 0 net=6574
rlabel metal2 1178 -2096 1178 -2096 0 net=9929
rlabel metal2 1542 -2096 1542 -2096 0 net=11835
rlabel metal2 1703 -2096 1703 -2096 0 net=12755
rlabel metal2 16 -2098 16 -2098 0 net=5265
rlabel metal2 247 -2098 247 -2098 0 net=1737
rlabel metal2 268 -2098 268 -2098 0 net=3397
rlabel metal2 506 -2098 506 -2098 0 net=4325
rlabel metal2 604 -2098 604 -2098 0 net=7289
rlabel metal2 779 -2098 779 -2098 0 net=5847
rlabel metal2 926 -2098 926 -2098 0 net=6441
rlabel metal2 954 -2098 954 -2098 0 net=6835
rlabel metal2 975 -2098 975 -2098 0 net=7034
rlabel metal2 1031 -2098 1031 -2098 0 net=10551
rlabel metal2 1220 -2098 1220 -2098 0 net=9885
rlabel metal2 1346 -2098 1346 -2098 0 net=10077
rlabel metal2 128 -2100 128 -2100 0 net=1855
rlabel metal2 163 -2100 163 -2100 0 net=2599
rlabel metal2 324 -2100 324 -2100 0 net=9173
rlabel metal2 618 -2100 618 -2100 0 net=5125
rlabel metal2 786 -2100 786 -2100 0 net=8455
rlabel metal2 1192 -2100 1192 -2100 0 net=8751
rlabel metal2 1220 -2100 1220 -2100 0 net=8969
rlabel metal2 1395 -2100 1395 -2100 0 net=10419
rlabel metal2 1619 -2100 1619 -2100 0 net=12583
rlabel metal2 1794 -2100 1794 -2100 0 net=12943
rlabel metal2 107 -2102 107 -2102 0 net=3361
rlabel metal2 135 -2102 135 -2102 0 net=4019
rlabel metal2 177 -2102 177 -2102 0 net=4645
rlabel metal2 341 -2102 341 -2102 0 net=5967
rlabel metal2 639 -2102 639 -2102 0 net=3950
rlabel metal2 884 -2102 884 -2102 0 net=5917
rlabel metal2 933 -2102 933 -2102 0 net=10085
rlabel metal2 1052 -2102 1052 -2102 0 net=11182
rlabel metal2 1717 -2102 1717 -2102 0 net=11997
rlabel metal2 1766 -2102 1766 -2102 0 net=13025
rlabel metal2 156 -2104 156 -2104 0 net=2581
rlabel metal2 191 -2104 191 -2104 0 net=8587
rlabel metal2 506 -2104 506 -2104 0 net=5307
rlabel metal2 870 -2104 870 -2104 0 net=5781
rlabel metal2 954 -2104 954 -2104 0 net=10405
rlabel metal2 1409 -2104 1409 -2104 0 net=9773
rlabel metal2 1696 -2104 1696 -2104 0 net=13683
rlabel metal2 184 -2106 184 -2106 0 net=1785
rlabel metal2 982 -2106 982 -2106 0 net=6895
rlabel metal2 1010 -2106 1010 -2106 0 net=7011
rlabel metal2 1066 -2106 1066 -2106 0 net=12993
rlabel metal2 1815 -2106 1815 -2106 0 net=13341
rlabel metal2 191 -2108 191 -2108 0 net=2889
rlabel metal2 485 -2108 485 -2108 0 net=3161
rlabel metal2 989 -2108 989 -2108 0 net=7689
rlabel metal2 1059 -2108 1059 -2108 0 net=7811
rlabel metal2 1192 -2108 1192 -2108 0 net=9255
rlabel metal2 1409 -2108 1409 -2108 0 net=10357
rlabel metal2 1822 -2108 1822 -2108 0 net=13589
rlabel metal2 198 -2110 198 -2110 0 net=2463
rlabel metal2 485 -2110 485 -2110 0 net=4359
rlabel metal2 576 -2110 576 -2110 0 net=3377
rlabel metal2 611 -2110 611 -2110 0 net=8535
rlabel metal2 1248 -2110 1248 -2110 0 net=8481
rlabel metal2 1465 -2110 1465 -2110 0 net=10903
rlabel metal2 1892 -2110 1892 -2110 0 net=2961
rlabel metal2 198 -2112 198 -2112 0 net=2027
rlabel metal2 236 -2112 236 -2112 0 net=295
rlabel metal2 989 -2112 989 -2112 0 net=7145
rlabel metal2 1115 -2112 1115 -2112 0 net=7157
rlabel metal2 1157 -2112 1157 -2112 0 net=13266
rlabel metal2 205 -2114 205 -2114 0 net=2411
rlabel metal2 996 -2114 996 -2114 0 net=7097
rlabel metal2 1045 -2114 1045 -2114 0 net=7227
rlabel metal2 1577 -2114 1577 -2114 0 net=12829
rlabel metal2 226 -2116 226 -2116 0 net=1545
rlabel metal2 247 -2116 247 -2116 0 net=4025
rlabel metal2 527 -2116 527 -2116 0 net=9337
rlabel metal2 1325 -2116 1325 -2116 0 net=9675
rlabel metal2 1738 -2116 1738 -2116 0 net=12417
rlabel metal2 212 -2118 212 -2118 0 net=2636
rlabel metal2 268 -2118 268 -2118 0 net=5165
rlabel metal2 527 -2118 527 -2118 0 net=6699
rlabel metal2 1003 -2118 1003 -2118 0 net=7399
rlabel metal2 1115 -2118 1115 -2118 0 net=8245
rlabel metal2 1248 -2118 1248 -2118 0 net=9621
rlabel metal2 1381 -2118 1381 -2118 0 net=11401
rlabel metal2 1738 -2118 1738 -2118 0 net=12773
rlabel metal2 1808 -2118 1808 -2118 0 net=13511
rlabel metal2 145 -2120 145 -2120 0 net=10155
rlabel metal2 1591 -2120 1591 -2120 0 net=11875
rlabel metal2 1801 -2120 1801 -2120 0 net=13291
rlabel metal2 170 -2122 170 -2122 0 net=3133
rlabel metal2 415 -2122 415 -2122 0 net=4201
rlabel metal2 1024 -2122 1024 -2122 0 net=10651
rlabel metal2 1682 -2122 1682 -2122 0 net=12503
rlabel metal2 1885 -2122 1885 -2122 0 net=13667
rlabel metal2 40 -2124 40 -2124 0 net=4783
rlabel metal2 212 -2124 212 -2124 0 net=2499
rlabel metal2 576 -2124 576 -2124 0 net=4143
rlabel metal2 737 -2124 737 -2124 0 net=5027
rlabel metal2 863 -2124 863 -2124 0 net=5715
rlabel metal2 1073 -2124 1073 -2124 0 net=7489
rlabel metal2 1199 -2124 1199 -2124 0 net=8851
rlabel metal2 1486 -2124 1486 -2124 0 net=11225
rlabel metal2 1689 -2124 1689 -2124 0 net=12021
rlabel metal2 114 -2126 114 -2126 0 net=3913
rlabel metal2 611 -2126 611 -2126 0 net=3625
rlabel metal2 628 -2126 628 -2126 0 net=5787
rlabel metal2 894 -2126 894 -2126 0 net=57
rlabel metal2 1486 -2126 1486 -2126 0 net=10697
rlabel metal2 1689 -2126 1689 -2126 0 net=12683
rlabel metal2 282 -2128 282 -2128 0 net=3087
rlabel metal2 625 -2128 625 -2128 0 net=3044
rlabel metal2 1080 -2128 1080 -2128 0 net=11320
rlabel metal2 1787 -2128 1787 -2128 0 net=13213
rlabel metal2 100 -2130 100 -2130 0 net=2663
rlabel metal2 289 -2130 289 -2130 0 net=4347
rlabel metal2 1255 -2130 1255 -2130 0 net=9829
rlabel metal2 1549 -2130 1549 -2130 0 net=10723
rlabel metal2 1780 -2130 1780 -2130 0 net=13155
rlabel metal2 1871 -2130 1871 -2130 0 net=13609
rlabel metal2 100 -2132 100 -2132 0 net=2757
rlabel metal2 1556 -2132 1556 -2132 0 net=11655
rlabel metal2 296 -2134 296 -2134 0 net=5427
rlabel metal2 639 -2134 639 -2134 0 net=7515
rlabel metal2 1269 -2134 1269 -2134 0 net=8739
rlabel metal2 1451 -2134 1451 -2134 0 net=11905
rlabel metal2 1612 -2134 1612 -2134 0 net=12593
rlabel metal2 254 -2136 254 -2136 0 net=5023
rlabel metal2 317 -2136 317 -2136 0 net=5685
rlabel metal2 1269 -2136 1269 -2136 0 net=9303
rlabel metal2 317 -2138 317 -2138 0 net=2291
rlabel metal2 345 -2138 345 -2138 0 net=2951
rlabel metal2 646 -2138 646 -2138 0 net=9270
rlabel metal2 1293 -2138 1293 -2138 0 net=12121
rlabel metal2 331 -2140 331 -2140 0 net=2837
rlabel metal2 653 -2140 653 -2140 0 net=4601
rlabel metal2 737 -2140 737 -2140 0 net=4959
rlabel metal2 800 -2140 800 -2140 0 net=8309
rlabel metal2 940 -2140 940 -2140 0 net=7339
rlabel metal2 1332 -2140 1332 -2140 0 net=10109
rlabel metal2 443 -2142 443 -2142 0 net=5361
rlabel metal2 793 -2142 793 -2142 0 net=6115
rlabel metal2 1444 -2142 1444 -2142 0 net=10629
rlabel metal2 275 -2144 275 -2144 0 net=5879
rlabel metal2 1430 -2144 1430 -2144 0 net=10039
rlabel metal2 275 -2146 275 -2146 0 net=5757
rlabel metal2 1430 -2146 1430 -2146 0 net=12007
rlabel metal2 453 -2148 453 -2148 0 net=5661
rlabel metal2 1528 -2148 1528 -2148 0 net=11575
rlabel metal2 457 -2150 457 -2150 0 net=3607
rlabel metal2 667 -2150 667 -2150 0 net=6585
rlabel metal2 1626 -2150 1626 -2150 0 net=13055
rlabel metal2 457 -2152 457 -2152 0 net=4549
rlabel metal2 667 -2152 667 -2152 0 net=4263
rlabel metal2 754 -2152 754 -2152 0 net=13715
rlabel metal2 555 -2154 555 -2154 0 net=4721
rlabel metal2 765 -2154 765 -2154 0 net=7855
rlabel metal2 1563 -2154 1563 -2154 0 net=10805
rlabel metal2 555 -2156 555 -2156 0 net=3893
rlabel metal2 660 -2156 660 -2156 0 net=4439
rlabel metal2 1563 -2156 1563 -2156 0 net=11693
rlabel metal2 404 -2158 404 -2158 0 net=12187
rlabel metal2 429 -2160 429 -2160 0 net=4427
rlabel metal2 674 -2160 674 -2160 0 net=4677
rlabel metal2 821 -2160 821 -2160 0 net=5159
rlabel metal2 429 -2162 429 -2162 0 net=4741
rlabel metal2 534 -2162 534 -2162 0 net=293
rlabel metal2 534 -2164 534 -2164 0 net=3523
rlabel metal2 681 -2166 681 -2166 0 net=5559
rlabel metal2 880 -2168 880 -2168 0 net=6884
rlabel metal2 1150 -2170 1150 -2170 0 net=8375
rlabel metal2 1227 -2172 1227 -2172 0 net=9195
rlabel metal2 912 -2174 912 -2174 0 net=4981
rlabel metal2 121 -2176 121 -2176 0 net=4235
rlabel metal2 72 -2178 72 -2178 0 net=6093
rlabel metal2 72 -2180 72 -2180 0 net=2737
rlabel metal2 58 -2182 58 -2182 0 net=5236
rlabel metal2 58 -2184 58 -2184 0 net=2425
rlabel metal2 2 -2195 2 -2195 0 net=3542
rlabel metal2 58 -2195 58 -2195 0 net=2426
rlabel metal2 222 -2195 222 -2195 0 net=964
rlabel metal2 1178 -2195 1178 -2195 0 net=9931
rlabel metal2 1454 -2195 1454 -2195 0 net=13512
rlabel metal2 12 -2197 12 -2197 0 net=5266
rlabel metal2 33 -2197 33 -2197 0 net=3558
rlabel metal2 527 -2197 527 -2197 0 net=6700
rlabel metal2 779 -2197 779 -2197 0 net=5309
rlabel metal2 779 -2197 779 -2197 0 net=5309
rlabel metal2 817 -2197 817 -2197 0 net=7226
rlabel metal2 1055 -2197 1055 -2197 0 net=4982
rlabel metal2 1360 -2197 1360 -2197 0 net=10698
rlabel metal2 1713 -2197 1713 -2197 0 net=10386
rlabel metal2 1727 -2197 1727 -2197 0 net=10782
rlabel metal2 16 -2199 16 -2199 0 net=2114
rlabel metal2 317 -2199 317 -2199 0 net=2292
rlabel metal2 352 -2199 352 -2199 0 net=2310
rlabel metal2 646 -2199 646 -2199 0 net=5849
rlabel metal2 950 -2199 950 -2199 0 net=12418
rlabel metal2 37 -2201 37 -2201 0 net=5576
rlabel metal2 877 -2201 877 -2201 0 net=8740
rlabel metal2 1318 -2201 1318 -2201 0 net=10667
rlabel metal2 1475 -2201 1475 -2201 0 net=13152
rlabel metal2 23 -2203 23 -2203 0 net=9109
rlabel metal2 44 -2203 44 -2203 0 net=6153
rlabel metal2 68 -2203 68 -2203 0 net=5024
rlabel metal2 303 -2203 303 -2203 0 net=3953
rlabel metal2 572 -2203 572 -2203 0 net=5782
rlabel metal2 891 -2203 891 -2203 0 net=9465
rlabel metal2 1395 -2203 1395 -2203 0 net=13214
rlabel metal2 23 -2205 23 -2205 0 net=2891
rlabel metal2 254 -2205 254 -2205 0 net=1684
rlabel metal2 1108 -2205 1108 -2205 0 net=7576
rlabel metal2 1276 -2205 1276 -2205 0 net=13215
rlabel metal2 1304 -2205 1304 -2205 0 net=13590
rlabel metal2 44 -2207 44 -2207 0 net=3363
rlabel metal2 163 -2207 163 -2207 0 net=2600
rlabel metal2 1136 -2207 1136 -2207 0 net=8971
rlabel metal2 1248 -2207 1248 -2207 0 net=9623
rlabel metal2 1248 -2207 1248 -2207 0 net=9623
rlabel metal2 1255 -2207 1255 -2207 0 net=9831
rlabel metal2 1276 -2207 1276 -2207 0 net=9677
rlabel metal2 1395 -2207 1395 -2207 0 net=12645
rlabel metal2 1717 -2207 1717 -2207 0 net=11999
rlabel metal2 1717 -2207 1717 -2207 0 net=11999
rlabel metal2 1787 -2207 1787 -2207 0 net=12945
rlabel metal2 1822 -2207 1822 -2207 0 net=2963
rlabel metal2 107 -2209 107 -2209 0 net=5758
rlabel metal2 282 -2209 282 -2209 0 net=2665
rlabel metal2 352 -2209 352 -2209 0 net=4327
rlabel metal2 670 -2209 670 -2209 0 net=13668
rlabel metal2 107 -2211 107 -2211 0 net=5547
rlabel metal2 877 -2211 877 -2211 0 net=6217
rlabel metal2 954 -2211 954 -2211 0 net=10407
rlabel metal2 1325 -2211 1325 -2211 0 net=10631
rlabel metal2 1458 -2211 1458 -2211 0 net=11071
rlabel metal2 1605 -2211 1605 -2211 0 net=12595
rlabel metal2 1794 -2211 1794 -2211 0 net=8181
rlabel metal2 110 -2213 110 -2213 0 net=9174
rlabel metal2 387 -2213 387 -2213 0 net=3608
rlabel metal2 520 -2213 520 -2213 0 net=5127
rlabel metal2 730 -2213 730 -2213 0 net=5105
rlabel metal2 730 -2213 730 -2213 0 net=5105
rlabel metal2 786 -2213 786 -2213 0 net=8457
rlabel metal2 1640 -2213 1640 -2213 0 net=13057
rlabel metal2 117 -2215 117 -2215 0 net=1856
rlabel metal2 163 -2215 163 -2215 0 net=4027
rlabel metal2 254 -2215 254 -2215 0 net=2839
rlabel metal2 408 -2215 408 -2215 0 net=3399
rlabel metal2 527 -2215 527 -2215 0 net=3627
rlabel metal2 695 -2215 695 -2215 0 net=4711
rlabel metal2 695 -2215 695 -2215 0 net=4711
rlabel metal2 737 -2215 737 -2215 0 net=4961
rlabel metal2 793 -2215 793 -2215 0 net=6117
rlabel metal2 880 -2215 880 -2215 0 net=12530
rlabel metal2 1640 -2215 1640 -2215 0 net=12995
rlabel metal2 128 -2217 128 -2217 0 net=4021
rlabel metal2 170 -2217 170 -2217 0 net=4785
rlabel metal2 408 -2217 408 -2217 0 net=4361
rlabel metal2 544 -2217 544 -2217 0 net=4236
rlabel metal2 919 -2217 919 -2217 0 net=6719
rlabel metal2 968 -2217 968 -2217 0 net=12830
rlabel metal2 1745 -2217 1745 -2217 0 net=11666
rlabel metal2 135 -2219 135 -2219 0 net=1787
rlabel metal2 191 -2219 191 -2219 0 net=1595
rlabel metal2 999 -2219 999 -2219 0 net=10040
rlabel metal2 170 -2221 170 -2221 0 net=5166
rlabel metal2 289 -2221 289 -2221 0 net=4349
rlabel metal2 331 -2221 331 -2221 0 net=2077
rlabel metal2 471 -2221 471 -2221 0 net=8589
rlabel metal2 1108 -2221 1108 -2221 0 net=9339
rlabel metal2 1353 -2221 1353 -2221 0 net=12197
rlabel metal2 79 -2223 79 -2223 0 net=2069
rlabel metal2 296 -2223 296 -2223 0 net=5363
rlabel metal2 457 -2223 457 -2223 0 net=4550
rlabel metal2 562 -2223 562 -2223 0 net=6875
rlabel metal2 737 -2223 737 -2223 0 net=5717
rlabel metal2 912 -2223 912 -2223 0 net=6443
rlabel metal2 968 -2223 968 -2223 0 net=7401
rlabel metal2 1038 -2223 1038 -2223 0 net=8005
rlabel metal2 1111 -2223 1111 -2223 0 net=10806
rlabel metal2 51 -2225 51 -2225 0 net=2187
rlabel metal2 485 -2225 485 -2225 0 net=3497
rlabel metal2 569 -2225 569 -2225 0 net=5429
rlabel metal2 796 -2225 796 -2225 0 net=6935
rlabel metal2 971 -2225 971 -2225 0 net=7340
rlabel metal2 1101 -2225 1101 -2225 0 net=8377
rlabel metal2 1178 -2225 1178 -2225 0 net=9887
rlabel metal2 1353 -2225 1353 -2225 0 net=8483
rlabel metal2 1444 -2225 1444 -2225 0 net=11493
rlabel metal2 1500 -2225 1500 -2225 0 net=11877
rlabel metal2 1626 -2225 1626 -2225 0 net=12775
rlabel metal2 30 -2227 30 -2227 0 net=10617
rlabel metal2 79 -2227 79 -2227 0 net=2759
rlabel metal2 142 -2227 142 -2227 0 net=4881
rlabel metal2 380 -2227 380 -2227 0 net=1914
rlabel metal2 590 -2227 590 -2227 0 net=8992
rlabel metal2 1279 -2227 1279 -2227 0 net=10724
rlabel metal2 1591 -2227 1591 -2227 0 net=12385
rlabel metal2 1696 -2227 1696 -2227 0 net=13685
rlabel metal2 30 -2229 30 -2229 0 net=10653
rlabel metal2 1031 -2229 1031 -2229 0 net=10553
rlabel metal2 1398 -2229 1398 -2229 0 net=13610
rlabel metal2 65 -2231 65 -2231 0 net=3773
rlabel metal2 177 -2231 177 -2231 0 net=4647
rlabel metal2 576 -2231 576 -2231 0 net=4145
rlabel metal2 597 -2231 597 -2231 0 net=4429
rlabel metal2 639 -2231 639 -2231 0 net=7516
rlabel metal2 926 -2231 926 -2231 0 net=6837
rlabel metal2 989 -2231 989 -2231 0 net=7147
rlabel metal2 1010 -2231 1010 -2231 0 net=7013
rlabel metal2 1052 -2231 1052 -2231 0 net=10865
rlabel metal2 1402 -2231 1402 -2231 0 net=12584
rlabel metal2 1675 -2231 1675 -2231 0 net=13395
rlabel metal2 86 -2233 86 -2233 0 net=6089
rlabel metal2 184 -2233 184 -2233 0 net=3465
rlabel metal2 226 -2233 226 -2233 0 net=1547
rlabel metal2 261 -2233 261 -2233 0 net=1739
rlabel metal2 415 -2233 415 -2233 0 net=4203
rlabel metal2 506 -2233 506 -2233 0 net=6995
rlabel metal2 989 -2233 989 -2233 0 net=7691
rlabel metal2 1024 -2233 1024 -2233 0 net=7813
rlabel metal2 1066 -2233 1066 -2233 0 net=8478
rlabel metal2 1188 -2233 1188 -2233 0 net=10110
rlabel metal2 1402 -2233 1402 -2233 0 net=12009
rlabel metal2 1479 -2233 1479 -2233 0 net=11695
rlabel metal2 1619 -2233 1619 -2233 0 net=12757
rlabel metal2 1829 -2233 1829 -2233 0 net=13489
rlabel metal2 86 -2235 86 -2235 0 net=2811
rlabel metal2 415 -2235 415 -2235 0 net=1627
rlabel metal2 506 -2235 506 -2235 0 net=4943
rlabel metal2 800 -2235 800 -2235 0 net=8311
rlabel metal2 1087 -2235 1087 -2235 0 net=9209
rlabel metal2 1192 -2235 1192 -2235 0 net=9257
rlabel metal2 1283 -2235 1283 -2235 0 net=10237
rlabel metal2 1430 -2235 1430 -2235 0 net=11205
rlabel metal2 1535 -2235 1535 -2235 0 net=12685
rlabel metal2 1696 -2235 1696 -2235 0 net=13343
rlabel metal2 173 -2237 173 -2237 0 net=9145
rlabel metal2 1010 -2237 1010 -2237 0 net=8537
rlabel metal2 1192 -2237 1192 -2237 0 net=9397
rlabel metal2 1332 -2237 1332 -2237 0 net=10421
rlabel metal2 1493 -2237 1493 -2237 0 net=11837
rlabel metal2 1549 -2237 1549 -2237 0 net=13079
rlabel metal2 93 -2239 93 -2239 0 net=11187
rlabel metal2 1514 -2239 1514 -2239 0 net=11743
rlabel metal2 1689 -2239 1689 -2239 0 net=13421
rlabel metal2 93 -2241 93 -2241 0 net=3181
rlabel metal2 198 -2241 198 -2241 0 net=2029
rlabel metal2 394 -2241 394 -2241 0 net=4051
rlabel metal2 576 -2241 576 -2241 0 net=2907
rlabel metal2 975 -2241 975 -2241 0 net=5733
rlabel metal2 1542 -2241 1542 -2241 0 net=11799
rlabel metal2 1703 -2241 1703 -2241 0 net=13523
rlabel metal2 198 -2243 198 -2243 0 net=2745
rlabel metal2 429 -2243 429 -2243 0 net=4743
rlabel metal2 649 -2243 649 -2243 0 net=11153
rlabel metal2 1563 -2243 1563 -2243 0 net=12133
rlabel metal2 1773 -2243 1773 -2243 0 net=13293
rlabel metal2 205 -2245 205 -2245 0 net=2413
rlabel metal2 345 -2245 345 -2245 0 net=2953
rlabel metal2 429 -2245 429 -2245 0 net=3163
rlabel metal2 1052 -2245 1052 -2245 0 net=10079
rlabel metal2 1570 -2245 1570 -2245 0 net=12189
rlabel metal2 72 -2247 72 -2247 0 net=2739
rlabel metal2 366 -2247 366 -2247 0 net=3915
rlabel metal2 611 -2247 611 -2247 0 net=4603
rlabel metal2 656 -2247 656 -2247 0 net=8633
rlabel metal2 1122 -2247 1122 -2247 0 net=7158
rlabel metal2 1164 -2247 1164 -2247 0 net=9273
rlabel metal2 1346 -2247 1346 -2247 0 net=10567
rlabel metal2 1584 -2247 1584 -2247 0 net=12301
rlabel metal2 72 -2249 72 -2249 0 net=6095
rlabel metal2 156 -2249 156 -2249 0 net=2582
rlabel metal2 208 -2249 208 -2249 0 net=7769
rlabel metal2 744 -2249 744 -2249 0 net=9563
rlabel metal2 121 -2251 121 -2251 0 net=9809
rlabel metal2 156 -2251 156 -2251 0 net=9774
rlabel metal2 212 -2253 212 -2253 0 net=2501
rlabel metal2 443 -2253 443 -2253 0 net=3337
rlabel metal2 618 -2253 618 -2253 0 net=5969
rlabel metal2 842 -2253 842 -2253 0 net=5919
rlabel metal2 1087 -2253 1087 -2253 0 net=8247
rlabel metal2 1122 -2253 1122 -2253 0 net=13046
rlabel metal2 212 -2255 212 -2255 0 net=5028
rlabel metal2 765 -2255 765 -2255 0 net=7857
rlabel metal2 1115 -2255 1115 -2255 0 net=7948
rlabel metal2 1213 -2255 1213 -2255 0 net=9391
rlabel metal2 1293 -2255 1293 -2255 0 net=13471
rlabel metal2 1710 -2255 1710 -2255 0 net=3193
rlabel metal2 219 -2257 219 -2257 0 net=569
rlabel metal2 450 -2257 450 -2257 0 net=3271
rlabel metal2 618 -2257 618 -2257 0 net=10087
rlabel metal2 1129 -2257 1129 -2257 0 net=8753
rlabel metal2 1220 -2257 1220 -2257 0 net=10359
rlabel metal2 1437 -2257 1437 -2257 0 net=11227
rlabel metal2 1633 -2257 1633 -2257 0 net=13407
rlabel metal2 226 -2259 226 -2259 0 net=2407
rlabel metal2 261 -2259 261 -2259 0 net=3089
rlabel metal2 366 -2259 366 -2259 0 net=3895
rlabel metal2 628 -2259 628 -2259 0 net=6175
rlabel metal2 1409 -2259 1409 -2259 0 net=11657
rlabel metal2 236 -2261 236 -2261 0 net=13047
rlabel metal2 240 -2263 240 -2263 0 net=12022
rlabel metal2 310 -2265 310 -2265 0 net=2465
rlabel metal2 422 -2265 422 -2265 0 net=6853
rlabel metal2 1521 -2265 1521 -2265 0 net=12505
rlabel metal2 1752 -2265 1752 -2265 0 net=13717
rlabel metal2 159 -2267 159 -2267 0 net=8735
rlabel metal2 373 -2267 373 -2267 0 net=3135
rlabel metal2 436 -2267 436 -2267 0 net=5789
rlabel metal2 905 -2267 905 -2267 0 net=6587
rlabel metal2 1556 -2267 1556 -2267 0 net=12123
rlabel metal2 1682 -2267 1682 -2267 0 net=13157
rlabel metal2 373 -2269 373 -2269 0 net=3847
rlabel metal2 555 -2269 555 -2269 0 net=5561
rlabel metal2 709 -2269 709 -2269 0 net=7291
rlabel metal2 870 -2269 870 -2269 0 net=5881
rlabel metal2 940 -2269 940 -2269 0 net=6897
rlabel metal2 1612 -2269 1612 -2269 0 net=13027
rlabel metal2 390 -2271 390 -2271 0 net=7501
rlabel metal2 499 -2273 499 -2273 0 net=3525
rlabel metal2 548 -2273 548 -2273 0 net=3379
rlabel metal2 639 -2273 639 -2273 0 net=2905
rlabel metal2 765 -2273 765 -2273 0 net=5687
rlabel metal2 898 -2273 898 -2273 0 net=6471
rlabel metal2 1731 -2273 1731 -2273 0 net=11441
rlabel metal2 89 -2275 89 -2275 0 net=7117
rlabel metal2 604 -2275 604 -2275 0 net=4679
rlabel metal2 677 -2275 677 -2275 0 net=11005
rlabel metal2 1472 -2275 1472 -2275 0 net=13537
rlabel metal2 653 -2277 653 -2277 0 net=7228
rlabel metal2 1157 -2277 1157 -2277 0 net=9197
rlabel metal2 660 -2279 660 -2279 0 net=4441
rlabel metal2 702 -2279 702 -2279 0 net=5041
rlabel metal2 744 -2279 744 -2279 0 net=5521
rlabel metal2 821 -2279 821 -2279 0 net=5161
rlabel metal2 982 -2279 982 -2279 0 net=7099
rlabel metal2 1185 -2279 1185 -2279 0 net=11635
rlabel metal2 9 -2281 9 -2281 0 net=11537
rlabel metal2 1227 -2281 1227 -2281 0 net=9761
rlabel metal2 660 -2283 660 -2283 0 net=4265
rlabel metal2 674 -2283 674 -2283 0 net=7490
rlabel metal2 1311 -2283 1311 -2283 0 net=11403
rlabel metal2 688 -2285 688 -2285 0 net=4723
rlabel metal2 751 -2285 751 -2285 0 net=7973
rlabel metal2 1073 -2285 1073 -2285 0 net=8345
rlabel metal2 583 -2287 583 -2287 0 net=3979
rlabel metal2 751 -2287 751 -2287 0 net=5325
rlabel metal2 835 -2287 835 -2287 0 net=10969
rlabel metal2 513 -2289 513 -2289 0 net=4065
rlabel metal2 807 -2289 807 -2289 0 net=5663
rlabel metal2 835 -2289 835 -2289 0 net=7059
rlabel metal2 978 -2289 978 -2289 0 net=10135
rlabel metal2 65 -2291 65 -2291 0 net=3703
rlabel metal2 821 -2291 821 -2291 0 net=9555
rlabel metal2 828 -2293 828 -2293 0 net=8853
rlabel metal2 1199 -2295 1199 -2295 0 net=9595
rlabel metal2 1374 -2297 1374 -2297 0 net=10905
rlabel metal2 1465 -2299 1465 -2299 0 net=11577
rlabel metal2 1507 -2301 1507 -2301 0 net=12069
rlabel metal2 1507 -2303 1507 -2303 0 net=11907
rlabel metal2 1069 -2305 1069 -2305 0 net=12675
rlabel metal2 1069 -2307 1069 -2307 0 net=8402
rlabel metal2 1171 -2309 1171 -2309 0 net=9305
rlabel metal2 1269 -2311 1269 -2311 0 net=10157
rlabel metal2 149 -2313 149 -2313 0 net=5985
rlabel metal2 9 -2324 9 -2324 0 net=11538
rlabel metal2 177 -2324 177 -2324 0 net=6090
rlabel metal2 1731 -2324 1731 -2324 0 net=13539
rlabel metal2 1748 -2324 1748 -2324 0 net=2964
rlabel metal2 9 -2326 9 -2326 0 net=4205
rlabel metal2 499 -2326 499 -2326 0 net=3526
rlabel metal2 821 -2326 821 -2326 0 net=6176
rlabel metal2 1216 -2326 1216 -2326 0 net=9932
rlabel metal2 1577 -2326 1577 -2326 0 net=12199
rlabel metal2 1755 -2326 1755 -2326 0 net=11442
rlabel metal2 1780 -2326 1780 -2326 0 net=7503
rlabel metal2 16 -2328 16 -2328 0 net=10088
rlabel metal2 625 -2328 625 -2328 0 net=10080
rlabel metal2 1069 -2328 1069 -2328 0 net=9392
rlabel metal2 1276 -2328 1276 -2328 0 net=9678
rlabel metal2 1307 -2328 1307 -2328 0 net=11072
rlabel metal2 1738 -2328 1738 -2328 0 net=13687
rlabel metal2 1787 -2328 1787 -2328 0 net=12947
rlabel metal2 16 -2330 16 -2330 0 net=5481
rlabel metal2 439 -2330 439 -2330 0 net=2188
rlabel metal2 460 -2330 460 -2330 0 net=4146
rlabel metal2 625 -2330 625 -2330 0 net=6589
rlabel metal2 947 -2330 947 -2330 0 net=8006
rlabel metal2 1052 -2330 1052 -2330 0 net=8458
rlabel metal2 1675 -2330 1675 -2330 0 net=13397
rlabel metal2 1759 -2330 1759 -2330 0 net=3195
rlabel metal2 1787 -2330 1787 -2330 0 net=8183
rlabel metal2 1797 -2330 1797 -2330 0 net=13490
rlabel metal2 30 -2332 30 -2332 0 net=10654
rlabel metal2 128 -2332 128 -2332 0 net=4022
rlabel metal2 128 -2332 128 -2332 0 net=4022
rlabel metal2 142 -2332 142 -2332 0 net=9810
rlabel metal2 233 -2332 233 -2332 0 net=4787
rlabel metal2 401 -2332 401 -2332 0 net=2954
rlabel metal2 401 -2332 401 -2332 0 net=2954
rlabel metal2 408 -2332 408 -2332 0 net=4362
rlabel metal2 793 -2332 793 -2332 0 net=5665
rlabel metal2 814 -2332 814 -2332 0 net=5735
rlabel metal2 989 -2332 989 -2332 0 net=7693
rlabel metal2 989 -2332 989 -2332 0 net=7693
rlabel metal2 996 -2332 996 -2332 0 net=11959
rlabel metal2 1619 -2332 1619 -2332 0 net=12759
rlabel metal2 1759 -2332 1759 -2332 0 net=13295
rlabel metal2 30 -2334 30 -2334 0 net=5987
rlabel metal2 159 -2334 159 -2334 0 net=4350
rlabel metal2 352 -2334 352 -2334 0 net=4328
rlabel metal2 698 -2334 698 -2334 0 net=5920
rlabel metal2 863 -2334 863 -2334 0 net=7293
rlabel metal2 1020 -2334 1020 -2334 0 net=9258
rlabel metal2 1248 -2334 1248 -2334 0 net=9625
rlabel metal2 1290 -2334 1290 -2334 0 net=13080
rlabel metal2 1619 -2334 1619 -2334 0 net=13423
rlabel metal2 1717 -2334 1717 -2334 0 net=12001
rlabel metal2 44 -2336 44 -2336 0 net=3364
rlabel metal2 247 -2336 247 -2336 0 net=1549
rlabel metal2 247 -2336 247 -2336 0 net=1549
rlabel metal2 282 -2336 282 -2336 0 net=2030
rlabel metal2 471 -2336 471 -2336 0 net=4649
rlabel metal2 632 -2336 632 -2336 0 net=4745
rlabel metal2 632 -2336 632 -2336 0 net=4745
rlabel metal2 646 -2336 646 -2336 0 net=5851
rlabel metal2 884 -2336 884 -2336 0 net=7148
rlabel metal2 1017 -2336 1017 -2336 0 net=7859
rlabel metal2 1321 -2336 1321 -2336 0 net=10632
rlabel metal2 1342 -2336 1342 -2336 0 net=13271
rlabel metal2 44 -2338 44 -2338 0 net=2409
rlabel metal2 303 -2338 303 -2338 0 net=3954
rlabel metal2 544 -2338 544 -2338 0 net=2906
rlabel metal2 646 -2338 646 -2338 0 net=4891
rlabel metal2 905 -2338 905 -2338 0 net=6445
rlabel metal2 947 -2338 947 -2338 0 net=6997
rlabel metal2 1024 -2338 1024 -2338 0 net=7815
rlabel metal2 1024 -2338 1024 -2338 0 net=7815
rlabel metal2 1038 -2338 1038 -2338 0 net=8313
rlabel metal2 1066 -2338 1066 -2338 0 net=9811
rlabel metal2 1370 -2338 1370 -2338 0 net=12646
rlabel metal2 1423 -2338 1423 -2338 0 net=11189
rlabel metal2 1486 -2338 1486 -2338 0 net=11839
rlabel metal2 1542 -2338 1542 -2338 0 net=11801
rlabel metal2 1633 -2338 1633 -2338 0 net=13409
rlabel metal2 51 -2340 51 -2340 0 net=10619
rlabel metal2 1010 -2340 1010 -2340 0 net=8539
rlabel metal2 1066 -2340 1066 -2340 0 net=8591
rlabel metal2 1087 -2340 1087 -2340 0 net=8249
rlabel metal2 1087 -2340 1087 -2340 0 net=8249
rlabel metal2 1101 -2340 1101 -2340 0 net=8379
rlabel metal2 1101 -2340 1101 -2340 0 net=8379
rlabel metal2 1115 -2340 1115 -2340 0 net=11744
rlabel metal2 1521 -2340 1521 -2340 0 net=12507
rlabel metal2 37 -2342 37 -2342 0 net=9110
rlabel metal2 1115 -2342 1115 -2342 0 net=9889
rlabel metal2 1188 -2342 1188 -2342 0 net=13158
rlabel metal2 37 -2344 37 -2344 0 net=4609
rlabel metal2 310 -2344 310 -2344 0 net=8736
rlabel metal2 467 -2344 467 -2344 0 net=11089
rlabel metal2 1430 -2344 1430 -2344 0 net=11207
rlabel metal2 1465 -2344 1465 -2344 0 net=11579
rlabel metal2 1521 -2344 1521 -2344 0 net=12125
rlabel metal2 1640 -2344 1640 -2344 0 net=12997
rlabel metal2 51 -2346 51 -2346 0 net=11095
rlabel metal2 310 -2346 310 -2346 0 net=1871
rlabel metal2 450 -2346 450 -2346 0 net=3273
rlabel metal2 478 -2346 478 -2346 0 net=3401
rlabel metal2 534 -2346 534 -2346 0 net=7119
rlabel metal2 1010 -2346 1010 -2346 0 net=8635
rlabel metal2 1129 -2346 1129 -2346 0 net=8755
rlabel metal2 1129 -2346 1129 -2346 0 net=8755
rlabel metal2 1136 -2346 1136 -2346 0 net=8973
rlabel metal2 1136 -2346 1136 -2346 0 net=8973
rlabel metal2 1157 -2346 1157 -2346 0 net=9199
rlabel metal2 1171 -2346 1171 -2346 0 net=9307
rlabel metal2 1213 -2346 1213 -2346 0 net=9557
rlabel metal2 1283 -2346 1283 -2346 0 net=10239
rlabel metal2 1360 -2346 1360 -2346 0 net=10867
rlabel metal2 1437 -2346 1437 -2346 0 net=11229
rlabel metal2 1479 -2346 1479 -2346 0 net=11697
rlabel metal2 1640 -2346 1640 -2346 0 net=13525
rlabel metal2 58 -2348 58 -2348 0 net=6154
rlabel metal2 86 -2348 86 -2348 0 net=2812
rlabel metal2 723 -2348 723 -2348 0 net=7771
rlabel metal2 1017 -2348 1017 -2348 0 net=9039
rlabel metal2 1227 -2348 1227 -2348 0 net=9763
rlabel metal2 1339 -2348 1339 -2348 0 net=10555
rlabel metal2 1416 -2348 1416 -2348 0 net=11155
rlabel metal2 1444 -2348 1444 -2348 0 net=11495
rlabel metal2 1500 -2348 1500 -2348 0 net=11879
rlabel metal2 1661 -2348 1661 -2348 0 net=13217
rlabel metal2 58 -2350 58 -2350 0 net=3735
rlabel metal2 296 -2350 296 -2350 0 net=5364
rlabel metal2 772 -2350 772 -2350 0 net=9147
rlabel metal2 1227 -2350 1227 -2350 0 net=9455
rlabel metal2 65 -2352 65 -2352 0 net=3499
rlabel metal2 513 -2352 513 -2352 0 net=3705
rlabel metal2 562 -2352 562 -2352 0 net=6876
rlabel metal2 831 -2352 831 -2352 0 net=11717
rlabel metal2 1626 -2352 1626 -2352 0 net=12777
rlabel metal2 72 -2354 72 -2354 0 net=6096
rlabel metal2 114 -2354 114 -2354 0 net=2747
rlabel metal2 205 -2354 205 -2354 0 net=7831
rlabel metal2 541 -2354 541 -2354 0 net=3917
rlabel metal2 583 -2354 583 -2354 0 net=4067
rlabel metal2 604 -2354 604 -2354 0 net=4681
rlabel metal2 667 -2354 667 -2354 0 net=4725
rlabel metal2 772 -2354 772 -2354 0 net=4963
rlabel metal2 856 -2354 856 -2354 0 net=5162
rlabel metal2 912 -2354 912 -2354 0 net=6839
rlabel metal2 1055 -2354 1055 -2354 0 net=9707
rlabel metal2 1332 -2354 1332 -2354 0 net=10423
rlabel metal2 1591 -2354 1591 -2354 0 net=12387
rlabel metal2 72 -2356 72 -2356 0 net=3775
rlabel metal2 107 -2356 107 -2356 0 net=5549
rlabel metal2 415 -2356 415 -2356 0 net=1629
rlabel metal2 478 -2356 478 -2356 0 net=4443
rlabel metal2 786 -2356 786 -2356 0 net=8103
rlabel metal2 856 -2356 856 -2356 0 net=5883
rlabel metal2 926 -2356 926 -2356 0 net=10159
rlabel metal2 1339 -2356 1339 -2356 0 net=13058
rlabel metal2 79 -2358 79 -2358 0 net=2761
rlabel metal2 289 -2358 289 -2358 0 net=2071
rlabel metal2 324 -2358 324 -2358 0 net=3629
rlabel metal2 541 -2358 541 -2358 0 net=3980
rlabel metal2 863 -2358 863 -2358 0 net=6029
rlabel metal2 1094 -2358 1094 -2358 0 net=9275
rlabel metal2 1199 -2358 1199 -2358 0 net=9597
rlabel metal2 1388 -2358 1388 -2358 0 net=11007
rlabel metal2 1528 -2358 1528 -2358 0 net=12071
rlabel metal2 1605 -2358 1605 -2358 0 net=12597
rlabel metal2 86 -2360 86 -2360 0 net=3183
rlabel metal2 96 -2360 96 -2360 0 net=13639
rlabel metal2 93 -2362 93 -2362 0 net=1126
rlabel metal2 135 -2362 135 -2362 0 net=1789
rlabel metal2 352 -2362 352 -2362 0 net=10915
rlabel metal2 1150 -2362 1150 -2362 0 net=9211
rlabel metal2 1269 -2362 1269 -2362 0 net=10669
rlabel metal2 1388 -2362 1388 -2362 0 net=13344
rlabel metal2 100 -2364 100 -2364 0 net=4029
rlabel metal2 170 -2364 170 -2364 0 net=3137
rlabel metal2 429 -2364 429 -2364 0 net=3165
rlabel metal2 870 -2364 870 -2364 0 net=6219
rlabel metal2 1150 -2364 1150 -2364 0 net=11321
rlabel metal2 1563 -2364 1563 -2364 0 net=12135
rlabel metal2 1654 -2364 1654 -2364 0 net=13049
rlabel metal2 121 -2366 121 -2366 0 net=1631
rlabel metal2 520 -2366 520 -2366 0 net=5129
rlabel metal2 877 -2366 877 -2366 0 net=6899
rlabel metal2 1157 -2366 1157 -2366 0 net=10361
rlabel metal2 1507 -2366 1507 -2366 0 net=11909
rlabel metal2 1598 -2366 1598 -2366 0 net=12677
rlabel metal2 107 -2368 107 -2368 0 net=6947
rlabel metal2 1083 -2368 1083 -2368 0 net=11625
rlabel metal2 1598 -2368 1598 -2368 0 net=13473
rlabel metal2 131 -2370 131 -2370 0 net=3357
rlabel metal2 142 -2370 142 -2370 0 net=3055
rlabel metal2 1164 -2370 1164 -2370 0 net=13028
rlabel metal2 149 -2372 149 -2372 0 net=2909
rlabel metal2 583 -2372 583 -2372 0 net=7403
rlabel metal2 1192 -2372 1192 -2372 0 net=9399
rlabel metal2 1535 -2372 1535 -2372 0 net=12687
rlabel metal2 156 -2374 156 -2374 0 net=2271
rlabel metal2 212 -2374 212 -2374 0 net=3425
rlabel metal2 219 -2374 219 -2374 0 net=5791
rlabel metal2 450 -2374 450 -2374 0 net=5719
rlabel metal2 968 -2374 968 -2374 0 net=7101
rlabel metal2 1535 -2374 1535 -2374 0 net=12191
rlabel metal2 1584 -2374 1584 -2374 0 net=12303
rlabel metal2 156 -2376 156 -2376 0 net=2141
rlabel metal2 1402 -2376 1402 -2376 0 net=12011
rlabel metal2 163 -2378 163 -2378 0 net=5107
rlabel metal2 737 -2378 737 -2378 0 net=5311
rlabel metal2 891 -2378 891 -2378 0 net=9467
rlabel metal2 1374 -2378 1374 -2378 0 net=10907
rlabel metal2 1570 -2378 1570 -2378 0 net=13719
rlabel metal2 177 -2380 177 -2380 0 net=2415
rlabel metal2 366 -2380 366 -2380 0 net=3896
rlabel metal2 436 -2380 436 -2380 0 net=4805
rlabel metal2 681 -2380 681 -2380 0 net=4713
rlabel metal2 730 -2380 730 -2380 0 net=11595
rlabel metal2 184 -2382 184 -2382 0 net=3467
rlabel metal2 366 -2382 366 -2382 0 net=2503
rlabel metal2 387 -2382 387 -2382 0 net=7405
rlabel metal2 891 -2382 891 -2382 0 net=6721
rlabel metal2 982 -2382 982 -2382 0 net=7015
rlabel metal2 1346 -2382 1346 -2382 0 net=10569
rlabel metal2 184 -2384 184 -2384 0 net=2467
rlabel metal2 390 -2384 390 -2384 0 net=7611
rlabel metal2 828 -2384 828 -2384 0 net=8855
rlabel metal2 191 -2386 191 -2386 0 net=1597
rlabel metal2 261 -2386 261 -2386 0 net=3091
rlabel metal2 485 -2386 485 -2386 0 net=3381
rlabel metal2 572 -2386 572 -2386 0 net=5613
rlabel metal2 828 -2386 828 -2386 0 net=13323
rlabel metal2 23 -2388 23 -2388 0 net=2892
rlabel metal2 205 -2388 205 -2388 0 net=2389
rlabel metal2 261 -2390 261 -2390 0 net=3339
rlabel metal2 520 -2390 520 -2390 0 net=6119
rlabel metal2 919 -2390 919 -2390 0 net=6855
rlabel metal2 1031 -2390 1031 -2390 0 net=7975
rlabel metal2 275 -2392 275 -2392 0 net=1741
rlabel metal2 338 -2392 338 -2392 0 net=2667
rlabel metal2 394 -2392 394 -2392 0 net=4053
rlabel metal2 527 -2392 527 -2392 0 net=11131
rlabel metal2 289 -2394 289 -2394 0 net=1803
rlabel metal2 548 -2394 548 -2394 0 net=5043
rlabel metal2 800 -2394 800 -2394 0 net=5971
rlabel metal2 933 -2394 933 -2394 0 net=6937
rlabel metal2 1045 -2394 1045 -2394 0 net=8913
rlabel metal2 317 -2396 317 -2396 0 net=4945
rlabel metal2 569 -2396 569 -2396 0 net=5267
rlabel metal2 765 -2396 765 -2396 0 net=5689
rlabel metal2 835 -2396 835 -2396 0 net=7061
rlabel metal2 1262 -2396 1262 -2396 0 net=9833
rlabel metal2 268 -2398 268 -2398 0 net=4883
rlabel metal2 555 -2398 555 -2398 0 net=5563
rlabel metal2 835 -2398 835 -2398 0 net=1903
rlabel metal2 268 -2400 268 -2400 0 net=2079
rlabel metal2 338 -2400 338 -2400 0 net=6472
rlabel metal2 1143 -2400 1143 -2400 0 net=10137
rlabel metal2 331 -2402 331 -2402 0 net=3517
rlabel metal2 695 -2402 695 -2402 0 net=1088
rlabel metal2 254 -2404 254 -2404 0 net=2840
rlabel metal2 898 -2404 898 -2404 0 net=5819
rlabel metal2 117 -2406 117 -2406 0 net=3197
rlabel metal2 341 -2406 341 -2406 0 net=9867
rlabel metal2 404 -2406 404 -2406 0 net=11701
rlabel metal2 345 -2408 345 -2408 0 net=2741
rlabel metal2 569 -2408 569 -2408 0 net=4605
rlabel metal2 656 -2408 656 -2408 0 net=9085
rlabel metal2 373 -2410 373 -2410 0 net=3849
rlabel metal2 576 -2410 576 -2410 0 net=4363
rlabel metal2 373 -2412 373 -2412 0 net=2601
rlabel metal2 1108 -2412 1108 -2412 0 net=9341
rlabel metal2 597 -2414 597 -2414 0 net=4431
rlabel metal2 1073 -2414 1073 -2414 0 net=8347
rlabel metal2 345 -2416 345 -2416 0 net=8403
rlabel metal2 604 -2416 604 -2416 0 net=4267
rlabel metal2 1073 -2416 1073 -2416 0 net=6341
rlabel metal2 660 -2418 660 -2418 0 net=3981
rlabel metal2 1367 -2418 1367 -2418 0 net=11637
rlabel metal2 1311 -2420 1311 -2420 0 net=11405
rlabel metal2 1311 -2422 1311 -2422 0 net=8485
rlabel metal2 1297 -2424 1297 -2424 0 net=10409
rlabel metal2 1297 -2426 1297 -2426 0 net=11659
rlabel metal2 1381 -2428 1381 -2428 0 net=10971
rlabel metal2 1234 -2430 1234 -2430 0 net=9565
rlabel metal2 758 -2432 758 -2432 0 net=9523
rlabel metal2 744 -2434 744 -2434 0 net=5523
rlabel metal2 744 -2436 744 -2436 0 net=5327
rlabel metal2 716 -2438 716 -2438 0 net=5431
rlabel metal2 9 -2449 9 -2449 0 net=4206
rlabel metal2 632 -2449 632 -2449 0 net=4747
rlabel metal2 632 -2449 632 -2449 0 net=4747
rlabel metal2 646 -2449 646 -2449 0 net=4893
rlabel metal2 646 -2449 646 -2449 0 net=4893
rlabel metal2 723 -2449 723 -2449 0 net=3166
rlabel metal2 1020 -2449 1020 -2449 0 net=11840
rlabel metal2 1741 -2449 1741 -2449 0 net=12002
rlabel metal2 1808 -2449 1808 -2449 0 net=12949
rlabel metal2 16 -2451 16 -2451 0 net=5483
rlabel metal2 44 -2451 44 -2451 0 net=2410
rlabel metal2 408 -2451 408 -2451 0 net=5550
rlabel metal2 726 -2451 726 -2451 0 net=13640
rlabel metal2 1745 -2451 1745 -2451 0 net=13541
rlabel metal2 1745 -2451 1745 -2451 0 net=13541
rlabel metal2 1752 -2451 1752 -2451 0 net=13297
rlabel metal2 1773 -2451 1773 -2451 0 net=13771
rlabel metal2 1801 -2451 1801 -2451 0 net=7505
rlabel metal2 16 -2453 16 -2453 0 net=12217
rlabel metal2 807 -2453 807 -2453 0 net=8105
rlabel metal2 814 -2453 814 -2453 0 net=5737
rlabel metal2 814 -2453 814 -2453 0 net=5737
rlabel metal2 828 -2453 828 -2453 0 net=1355
rlabel metal2 856 -2453 856 -2453 0 net=5885
rlabel metal2 856 -2453 856 -2453 0 net=5885
rlabel metal2 884 -2453 884 -2453 0 net=6840
rlabel metal2 919 -2453 919 -2453 0 net=6857
rlabel metal2 919 -2453 919 -2453 0 net=6857
rlabel metal2 950 -2453 950 -2453 0 net=9566
rlabel metal2 1423 -2453 1423 -2453 0 net=11091
rlabel metal2 1423 -2453 1423 -2453 0 net=11091
rlabel metal2 1619 -2453 1619 -2453 0 net=13425
rlabel metal2 1759 -2453 1759 -2453 0 net=13689
rlabel metal2 44 -2455 44 -2455 0 net=2911
rlabel metal2 159 -2455 159 -2455 0 net=554
rlabel metal2 439 -2455 439 -2455 0 net=9276
rlabel metal2 1132 -2455 1132 -2455 0 net=12126
rlabel metal2 1570 -2455 1570 -2455 0 net=13721
rlabel metal2 51 -2457 51 -2457 0 net=11096
rlabel metal2 583 -2457 583 -2457 0 net=7404
rlabel metal2 807 -2457 807 -2457 0 net=7063
rlabel metal2 982 -2457 982 -2457 0 net=7016
rlabel metal2 1150 -2457 1150 -2457 0 net=11323
rlabel metal2 1521 -2457 1521 -2457 0 net=11719
rlabel metal2 1619 -2457 1619 -2457 0 net=12689
rlabel metal2 51 -2459 51 -2459 0 net=4365
rlabel metal2 597 -2459 597 -2459 0 net=7406
rlabel metal2 828 -2459 828 -2459 0 net=6031
rlabel metal2 884 -2459 884 -2459 0 net=10161
rlabel metal2 940 -2459 940 -2459 0 net=6949
rlabel metal2 968 -2459 968 -2459 0 net=7103
rlabel metal2 1038 -2459 1038 -2459 0 net=8315
rlabel metal2 1038 -2459 1038 -2459 0 net=8315
rlabel metal2 1055 -2459 1055 -2459 0 net=9764
rlabel metal2 1325 -2459 1325 -2459 0 net=10241
rlabel metal2 1353 -2459 1353 -2459 0 net=10411
rlabel metal2 1353 -2459 1353 -2459 0 net=10411
rlabel metal2 1381 -2459 1381 -2459 0 net=10869
rlabel metal2 1542 -2459 1542 -2459 0 net=11881
rlabel metal2 1668 -2459 1668 -2459 0 net=13273
rlabel metal2 58 -2461 58 -2461 0 net=3736
rlabel metal2 408 -2461 408 -2461 0 net=7299
rlabel metal2 786 -2461 786 -2461 0 net=5853
rlabel metal2 887 -2461 887 -2461 0 net=12200
rlabel metal2 58 -2463 58 -2463 0 net=3341
rlabel metal2 324 -2463 324 -2463 0 net=3630
rlabel metal2 821 -2463 821 -2463 0 net=8915
rlabel metal2 1076 -2463 1076 -2463 0 net=13050
rlabel metal2 30 -2465 30 -2465 0 net=5989
rlabel metal2 275 -2465 275 -2465 0 net=1743
rlabel metal2 352 -2465 352 -2465 0 net=10917
rlabel metal2 1556 -2465 1556 -2465 0 net=12761
rlabel metal2 1689 -2465 1689 -2465 0 net=13411
rlabel metal2 30 -2467 30 -2467 0 net=3427
rlabel metal2 226 -2467 226 -2467 0 net=2763
rlabel metal2 429 -2467 429 -2467 0 net=4433
rlabel metal2 842 -2467 842 -2467 0 net=8593
rlabel metal2 1087 -2467 1087 -2467 0 net=8251
rlabel metal2 1150 -2467 1150 -2467 0 net=9149
rlabel metal2 1195 -2467 1195 -2467 0 net=12508
rlabel metal2 1640 -2467 1640 -2467 0 net=13527
rlabel metal2 65 -2469 65 -2469 0 net=3500
rlabel metal2 450 -2469 450 -2469 0 net=5720
rlabel metal2 530 -2469 530 -2469 0 net=4606
rlabel metal2 600 -2469 600 -2469 0 net=9261
rlabel metal2 1325 -2469 1325 -2469 0 net=10571
rlabel metal2 1640 -2469 1640 -2469 0 net=12679
rlabel metal2 1675 -2469 1675 -2469 0 net=13325
rlabel metal2 65 -2471 65 -2471 0 net=4947
rlabel metal2 352 -2471 352 -2471 0 net=2155
rlabel metal2 1332 -2471 1332 -2471 0 net=9599
rlabel metal2 72 -2473 72 -2473 0 net=3777
rlabel metal2 457 -2473 457 -2473 0 net=3013
rlabel metal2 600 -2473 600 -2473 0 net=357
rlabel metal2 905 -2473 905 -2473 0 net=6447
rlabel metal2 940 -2473 940 -2473 0 net=8541
rlabel metal2 1066 -2473 1066 -2473 0 net=8757
rlabel metal2 1160 -2473 1160 -2473 0 net=12778
rlabel metal2 1689 -2473 1689 -2473 0 net=13399
rlabel metal2 72 -2475 72 -2475 0 net=10275
rlabel metal2 198 -2475 198 -2475 0 net=2273
rlabel metal2 226 -2475 226 -2475 0 net=6999
rlabel metal2 971 -2475 971 -2475 0 net=10699
rlabel metal2 1598 -2475 1598 -2475 0 net=13475
rlabel metal2 1738 -2475 1738 -2475 0 net=3196
rlabel metal2 82 -2477 82 -2477 0 net=4788
rlabel metal2 243 -2477 243 -2477 0 net=8636
rlabel metal2 1048 -2477 1048 -2477 0 net=12779
rlabel metal2 1696 -2477 1696 -2477 0 net=8184
rlabel metal2 86 -2479 86 -2479 0 net=3185
rlabel metal2 86 -2479 86 -2479 0 net=3185
rlabel metal2 93 -2479 93 -2479 0 net=9868
rlabel metal2 443 -2479 443 -2479 0 net=12177
rlabel metal2 1654 -2479 1654 -2479 0 net=12999
rlabel metal2 93 -2481 93 -2481 0 net=2081
rlabel metal2 275 -2481 275 -2481 0 net=2743
rlabel metal2 443 -2481 443 -2481 0 net=4885
rlabel metal2 513 -2481 513 -2481 0 net=4068
rlabel metal2 681 -2481 681 -2481 0 net=4715
rlabel metal2 740 -2481 740 -2481 0 net=75
rlabel metal2 996 -2481 996 -2481 0 net=7773
rlabel metal2 1087 -2481 1087 -2481 0 net=9317
rlabel metal2 96 -2483 96 -2483 0 net=8404
rlabel metal2 366 -2483 366 -2483 0 net=2505
rlabel metal2 457 -2483 457 -2483 0 net=5973
rlabel metal2 877 -2483 877 -2483 0 net=6901
rlabel metal2 989 -2483 989 -2483 0 net=7695
rlabel metal2 1129 -2483 1129 -2483 0 net=10303
rlabel metal2 1255 -2483 1255 -2483 0 net=9559
rlabel metal2 37 -2485 37 -2485 0 net=4611
rlabel metal2 366 -2485 366 -2485 0 net=4651
rlabel metal2 653 -2485 653 -2485 0 net=4807
rlabel metal2 1115 -2485 1115 -2485 0 net=9891
rlabel metal2 1321 -2485 1321 -2485 0 net=1553
rlabel metal2 37 -2487 37 -2487 0 net=2749
rlabel metal2 128 -2487 128 -2487 0 net=1804
rlabel metal2 317 -2487 317 -2487 0 net=1989
rlabel metal2 471 -2487 471 -2487 0 net=1630
rlabel metal2 541 -2487 541 -2487 0 net=3983
rlabel metal2 849 -2487 849 -2487 0 net=3285
rlabel metal2 989 -2487 989 -2487 0 net=307
rlabel metal2 1332 -2487 1332 -2487 0 net=11581
rlabel metal2 100 -2489 100 -2489 0 net=4031
rlabel metal2 128 -2489 128 -2489 0 net=3469
rlabel metal2 289 -2489 289 -2489 0 net=1791
rlabel metal2 415 -2489 415 -2489 0 net=4055
rlabel metal2 478 -2489 478 -2489 0 net=4445
rlabel metal2 604 -2489 604 -2489 0 net=4269
rlabel metal2 1115 -2489 1115 -2489 0 net=11660
rlabel metal2 1318 -2489 1318 -2489 0 net=10557
rlabel metal2 1367 -2489 1367 -2489 0 net=11639
rlabel metal2 100 -2491 100 -2491 0 net=8856
rlabel metal2 1367 -2491 1367 -2491 0 net=11231
rlabel metal2 107 -2493 107 -2493 0 net=1466
rlabel metal2 478 -2493 478 -2493 0 net=5313
rlabel metal2 1003 -2493 1003 -2493 0 net=10621
rlabel metal2 1388 -2493 1388 -2493 0 net=10909
rlabel metal2 1465 -2493 1465 -2493 0 net=11497
rlabel metal2 107 -2495 107 -2495 0 net=9468
rlabel metal2 1241 -2495 1241 -2495 0 net=7861
rlabel metal2 110 -2497 110 -2497 0 net=739
rlabel metal2 1101 -2497 1101 -2497 0 net=8381
rlabel metal2 1241 -2497 1241 -2497 0 net=9813
rlabel metal2 1402 -2497 1402 -2497 0 net=10973
rlabel metal2 1479 -2497 1479 -2497 0 net=11627
rlabel metal2 103 -2499 103 -2499 0 net=7057
rlabel metal2 1157 -2499 1157 -2499 0 net=10363
rlabel metal2 1409 -2499 1409 -2499 0 net=11009
rlabel metal2 131 -2501 131 -2501 0 net=6743
rlabel metal2 1164 -2501 1164 -2501 0 net=8486
rlabel metal2 1416 -2501 1416 -2501 0 net=11157
rlabel metal2 135 -2503 135 -2503 0 net=3358
rlabel metal2 485 -2503 485 -2503 0 net=3383
rlabel metal2 604 -2503 604 -2503 0 net=7733
rlabel metal2 1164 -2503 1164 -2503 0 net=9213
rlabel metal2 1269 -2503 1269 -2503 0 net=10671
rlabel metal2 1437 -2503 1437 -2503 0 net=11191
rlabel metal2 135 -2505 135 -2505 0 net=1971
rlabel metal2 1080 -2505 1080 -2505 0 net=12953
rlabel metal2 1290 -2505 1290 -2505 0 net=11699
rlabel metal2 142 -2507 142 -2507 0 net=3057
rlabel metal2 436 -2507 436 -2507 0 net=7977
rlabel metal2 1080 -2507 1080 -2507 0 net=8975
rlabel metal2 1311 -2507 1311 -2507 0 net=8065
rlabel metal2 121 -2509 121 -2509 0 net=1633
rlabel metal2 149 -2509 149 -2509 0 net=12797
rlabel metal2 121 -2511 121 -2511 0 net=2143
rlabel metal2 163 -2511 163 -2511 0 net=5109
rlabel metal2 485 -2511 485 -2511 0 net=1905
rlabel metal2 1024 -2511 1024 -2511 0 net=7817
rlabel metal2 1122 -2511 1122 -2511 0 net=9343
rlabel metal2 1514 -2511 1514 -2511 0 net=11703
rlabel metal2 152 -2513 152 -2513 0 net=8121
rlabel metal2 639 -2513 639 -2513 0 net=4683
rlabel metal2 674 -2513 674 -2513 0 net=11241
rlabel metal2 1528 -2513 1528 -2513 0 net=13219
rlabel metal2 163 -2515 163 -2515 0 net=3665
rlabel metal2 1073 -2515 1073 -2515 0 net=6343
rlabel metal2 170 -2517 170 -2517 0 net=3139
rlabel metal2 492 -2517 492 -2517 0 net=3402
rlabel metal2 1108 -2517 1108 -2517 0 net=8349
rlabel metal2 170 -2519 170 -2519 0 net=9086
rlabel metal2 173 -2521 173 -2521 0 net=1872
rlabel metal2 492 -2521 492 -2521 0 net=7833
rlabel metal2 506 -2521 506 -2521 0 net=5131
rlabel metal2 702 -2521 702 -2521 0 net=7613
rlabel metal2 1108 -2521 1108 -2521 0 net=9201
rlabel metal2 191 -2523 191 -2523 0 net=6811
rlabel metal2 1143 -2523 1143 -2523 0 net=9309
rlabel metal2 191 -2525 191 -2525 0 net=6221
rlabel metal2 1192 -2525 1192 -2525 0 net=10424
rlabel metal2 198 -2527 198 -2527 0 net=1555
rlabel metal2 569 -2527 569 -2527 0 net=7121
rlabel metal2 1206 -2527 1206 -2527 0 net=9401
rlabel metal2 1444 -2527 1444 -2527 0 net=11209
rlabel metal2 219 -2529 219 -2529 0 net=5793
rlabel metal2 667 -2529 667 -2529 0 net=4727
rlabel metal2 737 -2529 737 -2529 0 net=12059
rlabel metal2 219 -2531 219 -2531 0 net=3275
rlabel metal2 499 -2531 499 -2531 0 net=3707
rlabel metal2 674 -2531 674 -2531 0 net=5269
rlabel metal2 789 -2531 789 -2531 0 net=6619
rlabel metal2 870 -2531 870 -2531 0 net=6939
rlabel metal2 961 -2531 961 -2531 0 net=7295
rlabel metal2 1220 -2531 1220 -2531 0 net=9627
rlabel metal2 233 -2533 233 -2533 0 net=1599
rlabel metal2 247 -2533 247 -2533 0 net=1550
rlabel metal2 464 -2533 464 -2533 0 net=5045
rlabel metal2 688 -2533 688 -2533 0 net=5433
rlabel metal2 975 -2533 975 -2533 0 net=9041
rlabel metal2 1276 -2533 1276 -2533 0 net=11407
rlabel metal2 247 -2535 247 -2535 0 net=1525
rlabel metal2 1171 -2535 1171 -2535 0 net=12192
rlabel metal2 254 -2537 254 -2537 0 net=3199
rlabel metal2 310 -2537 310 -2537 0 net=9095
rlabel metal2 709 -2537 709 -2537 0 net=8017
rlabel metal2 1472 -2537 1472 -2537 0 net=11597
rlabel metal2 1535 -2537 1535 -2537 0 net=11803
rlabel metal2 254 -2539 254 -2539 0 net=2603
rlabel metal2 513 -2539 513 -2539 0 net=3851
rlabel metal2 730 -2539 730 -2539 0 net=8051
rlabel metal2 1500 -2539 1500 -2539 0 net=11911
rlabel metal2 268 -2541 268 -2541 0 net=5053
rlabel metal2 730 -2541 730 -2541 0 net=2605
rlabel metal2 1549 -2541 1549 -2541 0 net=11961
rlabel metal2 282 -2543 282 -2543 0 net=3519
rlabel metal2 359 -2543 359 -2543 0 net=2669
rlabel metal2 520 -2543 520 -2543 0 net=6120
rlabel metal2 716 -2543 716 -2543 0 net=5525
rlabel metal2 1563 -2543 1563 -2543 0 net=12013
rlabel metal2 177 -2545 177 -2545 0 net=2417
rlabel metal2 520 -2545 520 -2545 0 net=5691
rlabel metal2 1577 -2545 1577 -2545 0 net=12073
rlabel metal2 177 -2547 177 -2547 0 net=2391
rlabel metal2 527 -2547 527 -2547 0 net=3919
rlabel metal2 625 -2547 625 -2547 0 net=6591
rlabel metal2 1584 -2547 1584 -2547 0 net=12137
rlabel metal2 184 -2549 184 -2549 0 net=2469
rlabel metal2 534 -2549 534 -2549 0 net=5329
rlabel metal2 751 -2549 751 -2549 0 net=3209
rlabel metal2 1591 -2549 1591 -2549 0 net=12599
rlabel metal2 184 -2551 184 -2551 0 net=7717
rlabel metal2 548 -2551 548 -2551 0 net=3669
rlabel metal2 1213 -2551 1213 -2551 0 net=9457
rlabel metal2 1283 -2551 1283 -2551 0 net=9709
rlabel metal2 205 -2553 205 -2553 0 net=3093
rlabel metal2 562 -2553 562 -2553 0 net=3293
rlabel metal2 744 -2553 744 -2553 0 net=5565
rlabel metal2 968 -2553 968 -2553 0 net=9721
rlabel metal2 1262 -2553 1262 -2553 0 net=10139
rlabel metal2 1605 -2553 1605 -2553 0 net=12305
rlabel metal2 156 -2555 156 -2555 0 net=3609
rlabel metal2 625 -2555 625 -2555 0 net=11447
rlabel metal2 1612 -2555 1612 -2555 0 net=12389
rlabel metal2 79 -2557 79 -2557 0 net=12711
rlabel metal2 79 -2559 79 -2559 0 net=2073
rlabel metal2 758 -2559 758 -2559 0 net=4965
rlabel metal2 1262 -2559 1262 -2559 0 net=11133
rlabel metal2 296 -2561 296 -2561 0 net=2447
rlabel metal2 765 -2561 765 -2561 0 net=5615
rlabel metal2 1234 -2561 1234 -2561 0 net=9525
rlabel metal2 772 -2563 772 -2563 0 net=5667
rlabel metal2 1234 -2563 1234 -2563 0 net=9835
rlabel metal2 110 -2565 110 -2565 0 net=10471
rlabel metal2 670 -2567 670 -2567 0 net=6271
rlabel metal2 779 -2569 779 -2569 0 net=5821
rlabel metal2 891 -2571 891 -2571 0 net=6723
rlabel metal2 453 -2573 453 -2573 0 net=6953
rlabel metal2 9 -2584 9 -2584 0 net=4887
rlabel metal2 450 -2584 450 -2584 0 net=8106
rlabel metal2 1062 -2584 1062 -2584 0 net=11408
rlabel metal2 1293 -2584 1293 -2584 0 net=10242
rlabel metal2 1465 -2584 1465 -2584 0 net=11499
rlabel metal2 1465 -2584 1465 -2584 0 net=11499
rlabel metal2 1510 -2584 1510 -2584 0 net=12600
rlabel metal2 1724 -2584 1724 -2584 0 net=13477
rlabel metal2 1724 -2584 1724 -2584 0 net=13477
rlabel metal2 1738 -2584 1738 -2584 0 net=1554
rlabel metal2 16 -2586 16 -2586 0 net=12218
rlabel metal2 16 -2586 16 -2586 0 net=12218
rlabel metal2 44 -2586 44 -2586 0 net=2912
rlabel metal2 639 -2586 639 -2586 0 net=7064
rlabel metal2 852 -2586 852 -2586 0 net=7696
rlabel metal2 1020 -2586 1020 -2586 0 net=9202
rlabel metal2 1115 -2586 1115 -2586 0 net=8067
rlabel metal2 1339 -2586 1339 -2586 0 net=10701
rlabel metal2 1563 -2586 1563 -2586 0 net=12015
rlabel metal2 1563 -2586 1563 -2586 0 net=12015
rlabel metal2 1769 -2586 1769 -2586 0 net=1147
rlabel metal2 44 -2588 44 -2588 0 net=5823
rlabel metal2 807 -2588 807 -2588 0 net=6033
rlabel metal2 866 -2588 866 -2588 0 net=1462
rlabel metal2 107 -2590 107 -2590 0 net=4652
rlabel metal2 443 -2590 443 -2590 0 net=3015
rlabel metal2 660 -2590 660 -2590 0 net=4270
rlabel metal2 726 -2590 726 -2590 0 net=9710
rlabel metal2 79 -2592 79 -2592 0 net=2075
rlabel metal2 121 -2592 121 -2592 0 net=2145
rlabel metal2 243 -2592 243 -2592 0 net=3520
rlabel metal2 292 -2592 292 -2592 0 net=121
rlabel metal2 660 -2592 660 -2592 0 net=6941
rlabel metal2 898 -2592 898 -2592 0 net=6725
rlabel metal2 898 -2592 898 -2592 0 net=6725
rlabel metal2 915 -2592 915 -2592 0 net=10412
rlabel metal2 1507 -2592 1507 -2592 0 net=11805
rlabel metal2 1647 -2592 1647 -2592 0 net=13001
rlabel metal2 79 -2594 79 -2594 0 net=8595
rlabel metal2 947 -2594 947 -2594 0 net=6601
rlabel metal2 1276 -2594 1276 -2594 0 net=10473
rlabel metal2 1311 -2594 1311 -2594 0 net=10911
rlabel metal2 1654 -2594 1654 -2594 0 net=13029
rlabel metal2 121 -2596 121 -2596 0 net=3471
rlabel metal2 149 -2596 149 -2596 0 net=3778
rlabel metal2 457 -2596 457 -2596 0 net=5974
rlabel metal2 695 -2596 695 -2596 0 net=4716
rlabel metal2 737 -2596 737 -2596 0 net=11324
rlabel metal2 68 -2598 68 -2598 0 net=2189
rlabel metal2 156 -2598 156 -2598 0 net=2604
rlabel metal2 261 -2598 261 -2598 0 net=5991
rlabel metal2 261 -2598 261 -2598 0 net=5991
rlabel metal2 275 -2598 275 -2598 0 net=2744
rlabel metal2 642 -2598 642 -2598 0 net=12043
rlabel metal2 86 -2600 86 -2600 0 net=3187
rlabel metal2 142 -2600 142 -2600 0 net=1635
rlabel metal2 282 -2600 282 -2600 0 net=1793
rlabel metal2 296 -2600 296 -2600 0 net=2448
rlabel metal2 681 -2600 681 -2600 0 net=4809
rlabel metal2 758 -2600 758 -2600 0 net=4967
rlabel metal2 758 -2600 758 -2600 0 net=4967
rlabel metal2 765 -2600 765 -2600 0 net=5617
rlabel metal2 842 -2600 842 -2600 0 net=10162
rlabel metal2 968 -2600 968 -2600 0 net=9526
rlabel metal2 1486 -2600 1486 -2600 0 net=11883
rlabel metal2 86 -2602 86 -2602 0 net=8383
rlabel metal2 103 -2602 103 -2602 0 net=464
rlabel metal2 296 -2602 296 -2602 0 net=5395
rlabel metal2 1048 -2602 1048 -2602 0 net=11700
rlabel metal2 1304 -2602 1304 -2602 0 net=10673
rlabel metal2 1430 -2602 1430 -2602 0 net=11211
rlabel metal2 1542 -2602 1542 -2602 0 net=12061
rlabel metal2 37 -2604 37 -2604 0 net=2751
rlabel metal2 142 -2604 142 -2604 0 net=7979
rlabel metal2 453 -2604 453 -2604 0 net=1857
rlabel metal2 695 -2604 695 -2604 0 net=6813
rlabel metal2 905 -2604 905 -2604 0 net=6903
rlabel metal2 971 -2604 971 -2604 0 net=6344
rlabel metal2 37 -2606 37 -2606 0 net=6401
rlabel metal2 856 -2606 856 -2606 0 net=5887
rlabel metal2 905 -2606 905 -2606 0 net=10743
rlabel metal2 989 -2606 989 -2606 0 net=8316
rlabel metal2 1073 -2606 1073 -2606 0 net=8253
rlabel metal2 1108 -2606 1108 -2606 0 net=9311
rlabel metal2 1157 -2606 1157 -2606 0 net=9629
rlabel metal2 1262 -2606 1262 -2606 0 net=11135
rlabel metal2 1444 -2606 1444 -2606 0 net=11449
rlabel metal2 1570 -2606 1570 -2606 0 net=12179
rlabel metal2 1675 -2606 1675 -2606 0 net=13327
rlabel metal2 156 -2608 156 -2608 0 net=1557
rlabel metal2 205 -2608 205 -2608 0 net=3095
rlabel metal2 492 -2608 492 -2608 0 net=7835
rlabel metal2 775 -2608 775 -2608 0 net=6599
rlabel metal2 1458 -2608 1458 -2608 0 net=11705
rlabel metal2 1598 -2608 1598 -2608 0 net=12691
rlabel metal2 1675 -2608 1675 -2608 0 net=13427
rlabel metal2 159 -2610 159 -2610 0 net=3286
rlabel metal2 940 -2610 940 -2610 0 net=8543
rlabel metal2 1174 -2610 1174 -2610 0 net=11582
rlabel metal2 1353 -2610 1353 -2610 0 net=11011
rlabel metal2 1514 -2610 1514 -2610 0 net=11127
rlabel metal2 1710 -2610 1710 -2610 0 net=13413
rlabel metal2 170 -2612 170 -2612 0 net=10304
rlabel metal2 1409 -2612 1409 -2612 0 net=12307
rlabel metal2 1689 -2612 1689 -2612 0 net=13401
rlabel metal2 170 -2614 170 -2614 0 net=7735
rlabel metal2 702 -2614 702 -2614 0 net=4728
rlabel metal2 856 -2614 856 -2614 0 net=6519
rlabel metal2 1066 -2614 1066 -2614 0 net=8759
rlabel metal2 1556 -2614 1556 -2614 0 net=12763
rlabel metal2 1689 -2614 1689 -2614 0 net=13723
rlabel metal2 173 -2616 173 -2616 0 net=7058
rlabel metal2 1118 -2616 1118 -2616 0 net=12445
rlabel metal2 177 -2618 177 -2618 0 net=2393
rlabel metal2 303 -2618 303 -2618 0 net=3201
rlabel metal2 492 -2618 492 -2618 0 net=2607
rlabel metal2 828 -2618 828 -2618 0 net=4273
rlabel metal2 23 -2620 23 -2620 0 net=5485
rlabel metal2 184 -2620 184 -2620 0 net=7718
rlabel metal2 702 -2620 702 -2620 0 net=5855
rlabel metal2 870 -2620 870 -2620 0 net=6103
rlabel metal2 1076 -2620 1076 -2620 0 net=8382
rlabel metal2 1220 -2620 1220 -2620 0 net=10559
rlabel metal2 1556 -2620 1556 -2620 0 net=12139
rlabel metal2 184 -2622 184 -2622 0 net=1619
rlabel metal2 205 -2622 205 -2622 0 net=4612
rlabel metal2 387 -2622 387 -2622 0 net=5435
rlabel metal2 709 -2622 709 -2622 0 net=9402
rlabel metal2 1241 -2622 1241 -2622 0 net=9815
rlabel metal2 1584 -2622 1584 -2622 0 net=12391
rlabel metal2 226 -2624 226 -2624 0 net=7000
rlabel metal2 1024 -2624 1024 -2624 0 net=7615
rlabel metal2 1094 -2624 1094 -2624 0 net=9151
rlabel metal2 1241 -2624 1241 -2624 0 net=11232
rlabel metal2 1612 -2624 1612 -2624 0 net=12713
rlabel metal2 30 -2626 30 -2626 0 net=3429
rlabel metal2 303 -2626 303 -2626 0 net=1907
rlabel metal2 513 -2626 513 -2626 0 net=3852
rlabel metal2 646 -2626 646 -2626 0 net=4895
rlabel metal2 723 -2626 723 -2626 0 net=11053
rlabel metal2 1367 -2626 1367 -2626 0 net=11641
rlabel metal2 1626 -2626 1626 -2626 0 net=12799
rlabel metal2 30 -2628 30 -2628 0 net=4949
rlabel metal2 310 -2628 310 -2628 0 net=9096
rlabel metal2 436 -2628 436 -2628 0 net=5527
rlabel metal2 730 -2628 730 -2628 0 net=5567
rlabel metal2 786 -2628 786 -2628 0 net=8961
rlabel metal2 1248 -2628 1248 -2628 0 net=9797
rlabel metal2 1479 -2628 1479 -2628 0 net=11629
rlabel metal2 1633 -2628 1633 -2628 0 net=13529
rlabel metal2 58 -2630 58 -2630 0 net=3343
rlabel metal2 520 -2630 520 -2630 0 net=5692
rlabel metal2 912 -2630 912 -2630 0 net=6449
rlabel metal2 933 -2630 933 -2630 0 net=8053
rlabel metal2 1731 -2630 1731 -2630 0 net=13543
rlabel metal2 58 -2632 58 -2632 0 net=6592
rlabel metal2 835 -2632 835 -2632 0 net=6621
rlabel metal2 940 -2632 940 -2632 0 net=10919
rlabel metal2 1745 -2632 1745 -2632 0 net=13299
rlabel metal2 110 -2634 110 -2634 0 net=6025
rlabel metal2 317 -2634 317 -2634 0 net=1991
rlabel metal2 317 -2634 317 -2634 0 net=1991
rlabel metal2 338 -2634 338 -2634 0 net=3141
rlabel metal2 380 -2634 380 -2634 0 net=5111
rlabel metal2 716 -2634 716 -2634 0 net=2711
rlabel metal2 1395 -2634 1395 -2634 0 net=11159
rlabel metal2 1752 -2634 1752 -2634 0 net=13691
rlabel metal2 135 -2636 135 -2636 0 net=1973
rlabel metal2 919 -2636 919 -2636 0 net=6859
rlabel metal2 1416 -2636 1416 -2636 0 net=11599
rlabel metal2 1759 -2636 1759 -2636 0 net=13773
rlabel metal2 135 -2638 135 -2638 0 net=1601
rlabel metal2 338 -2638 338 -2638 0 net=2765
rlabel metal2 408 -2638 408 -2638 0 net=7301
rlabel metal2 996 -2638 996 -2638 0 net=7775
rlabel metal2 1017 -2638 1017 -2638 0 net=9560
rlabel metal2 72 -2640 72 -2640 0 net=10277
rlabel metal2 345 -2640 345 -2640 0 net=2157
rlabel metal2 359 -2640 359 -2640 0 net=2471
rlabel metal2 394 -2640 394 -2640 0 net=2507
rlabel metal2 422 -2640 422 -2640 0 net=3611
rlabel metal2 520 -2640 520 -2640 0 net=12780
rlabel metal2 72 -2642 72 -2642 0 net=5047
rlabel metal2 523 -2642 523 -2642 0 net=7122
rlabel metal2 646 -2642 646 -2642 0 net=4685
rlabel metal2 674 -2642 674 -2642 0 net=5271
rlabel metal2 800 -2642 800 -2642 0 net=5249
rlabel metal2 1003 -2642 1003 -2642 0 net=8019
rlabel metal2 1101 -2642 1101 -2642 0 net=9215
rlabel metal2 1171 -2642 1171 -2642 0 net=10365
rlabel metal2 1472 -2642 1472 -2642 0 net=11721
rlabel metal2 152 -2644 152 -2644 0 net=12961
rlabel metal2 201 -2646 201 -2646 0 net=11867
rlabel metal2 1521 -2646 1521 -2646 0 net=11963
rlabel metal2 268 -2648 268 -2648 0 net=5055
rlabel metal2 891 -2648 891 -2648 0 net=6955
rlabel metal2 1024 -2648 1024 -2648 0 net=8977
rlabel metal2 1122 -2648 1122 -2648 0 net=8350
rlabel metal2 1139 -2648 1139 -2648 0 net=13641
rlabel metal2 268 -2650 268 -2650 0 net=2637
rlabel metal2 1297 -2650 1297 -2650 0 net=10573
rlabel metal2 1549 -2650 1549 -2650 0 net=12075
rlabel metal2 324 -2652 324 -2652 0 net=1745
rlabel metal2 359 -2652 359 -2652 0 net=4435
rlabel metal2 464 -2652 464 -2652 0 net=6273
rlabel metal2 821 -2652 821 -2652 0 net=8917
rlabel metal2 1325 -2652 1325 -2652 0 net=12731
rlabel metal2 324 -2654 324 -2654 0 net=3671
rlabel metal2 569 -2654 569 -2654 0 net=4447
rlabel metal2 625 -2654 625 -2654 0 net=6155
rlabel metal2 912 -2654 912 -2654 0 net=7341
rlabel metal2 1122 -2654 1122 -2654 0 net=9263
rlabel metal2 1577 -2654 1577 -2654 0 net=12275
rlabel metal2 163 -2656 163 -2656 0 net=3667
rlabel metal2 590 -2656 590 -2656 0 net=5795
rlabel metal2 625 -2656 625 -2656 0 net=4237
rlabel metal2 954 -2656 954 -2656 0 net=6951
rlabel metal2 1087 -2656 1087 -2656 0 net=9319
rlabel metal2 163 -2658 163 -2658 0 net=3277
rlabel metal2 373 -2658 373 -2658 0 net=2671
rlabel metal2 415 -2658 415 -2658 0 net=3059
rlabel metal2 506 -2658 506 -2658 0 net=5133
rlabel metal2 632 -2658 632 -2658 0 net=4749
rlabel metal2 772 -2658 772 -2658 0 net=5669
rlabel metal2 814 -2658 814 -2658 0 net=5739
rlabel metal2 849 -2658 849 -2658 0 net=13241
rlabel metal2 219 -2660 219 -2660 0 net=1527
rlabel metal2 331 -2660 331 -2660 0 net=2419
rlabel metal2 394 -2660 394 -2660 0 net=3211
rlabel metal2 814 -2660 814 -2660 0 net=9345
rlabel metal2 93 -2662 93 -2662 0 net=2083
rlabel metal2 415 -2662 415 -2662 0 net=2693
rlabel metal2 1199 -2662 1199 -2662 0 net=9459
rlabel metal2 93 -2664 93 -2664 0 net=4033
rlabel metal2 191 -2664 191 -2664 0 net=6223
rlabel metal2 478 -2664 478 -2664 0 net=5314
rlabel metal2 863 -2664 863 -2664 0 net=6745
rlabel metal2 961 -2664 961 -2664 0 net=7297
rlabel metal2 1195 -2664 1195 -2664 0 net=11912
rlabel metal2 114 -2666 114 -2666 0 net=3717
rlabel metal2 471 -2666 471 -2666 0 net=4057
rlabel metal2 506 -2666 506 -2666 0 net=3295
rlabel metal2 597 -2666 597 -2666 0 net=4449
rlabel metal2 635 -2666 635 -2666 0 net=10243
rlabel metal2 961 -2666 961 -2666 0 net=7105
rlabel metal2 1045 -2666 1045 -2666 0 net=5449
rlabel metal2 1132 -2666 1132 -2666 0 net=13274
rlabel metal2 191 -2668 191 -2668 0 net=2275
rlabel metal2 471 -2668 471 -2668 0 net=4663
rlabel metal2 1213 -2668 1213 -2668 0 net=9601
rlabel metal2 51 -2670 51 -2670 0 net=4367
rlabel metal2 499 -2670 499 -2670 0 net=3709
rlabel metal2 975 -2670 975 -2670 0 net=9043
rlabel metal2 1045 -2670 1045 -2670 0 net=10623
rlabel metal2 1500 -2670 1500 -2670 0 net=7863
rlabel metal2 1801 -2670 1801 -2670 0 net=7507
rlabel metal2 51 -2672 51 -2672 0 net=7749
rlabel metal2 499 -2672 499 -2672 0 net=5405
rlabel metal2 975 -2672 975 -2672 0 net=7818
rlabel metal2 1346 -2672 1346 -2672 0 net=10871
rlabel metal2 1528 -2672 1528 -2672 0 net=13221
rlabel metal2 1787 -2672 1787 -2672 0 net=12613
rlabel metal2 1808 -2672 1808 -2672 0 net=12951
rlabel metal2 527 -2674 527 -2674 0 net=3921
rlabel metal2 534 -2674 534 -2674 0 net=5331
rlabel metal2 1381 -2674 1381 -2674 0 net=10975
rlabel metal2 1696 -2674 1696 -2674 0 net=11955
rlabel metal2 527 -2676 527 -2676 0 net=3985
rlabel metal2 555 -2676 555 -2676 0 net=13267
rlabel metal2 555 -2678 555 -2678 0 net=3385
rlabel metal2 611 -2678 611 -2678 0 net=8123
rlabel metal2 1192 -2678 1192 -2678 0 net=11183
rlabel metal2 534 -2680 534 -2680 0 net=6257
rlabel metal2 576 -2682 576 -2682 0 net=3795
rlabel metal2 611 -2684 611 -2684 0 net=4523
rlabel metal2 709 -2686 709 -2686 0 net=11985
rlabel metal2 1055 -2688 1055 -2688 0 net=12680
rlabel metal2 1059 -2690 1059 -2690 0 net=3177
rlabel metal2 1269 -2690 1269 -2690 0 net=12955
rlabel metal2 1234 -2692 1234 -2692 0 net=9837
rlabel metal2 1227 -2694 1227 -2694 0 net=9723
rlabel metal2 1227 -2696 1227 -2696 0 net=10141
rlabel metal2 1255 -2698 1255 -2698 0 net=9893
rlabel metal2 1255 -2700 1255 -2700 0 net=11243
rlabel metal2 1423 -2702 1423 -2702 0 net=11093
rlabel metal2 1423 -2704 1423 -2704 0 net=11193
rlabel metal2 1192 -2706 1192 -2706 0 net=11347
rlabel metal2 30 -2717 30 -2717 0 net=4950
rlabel metal2 737 -2717 737 -2717 0 net=4811
rlabel metal2 842 -2717 842 -2717 0 net=11630
rlabel metal2 1769 -2717 1769 -2717 0 net=12952
rlabel metal2 44 -2719 44 -2719 0 net=5824
rlabel metal2 72 -2719 72 -2719 0 net=5048
rlabel metal2 646 -2719 646 -2719 0 net=4687
rlabel metal2 646 -2719 646 -2719 0 net=4687
rlabel metal2 712 -2719 712 -2719 0 net=314
rlabel metal2 1290 -2719 1290 -2719 0 net=11055
rlabel metal2 1433 -2719 1433 -2719 0 net=11094
rlabel metal2 1493 -2719 1493 -2719 0 net=11807
rlabel metal2 1780 -2719 1780 -2719 0 net=7508
rlabel metal2 58 -2721 58 -2721 0 net=4165
rlabel metal2 96 -2721 96 -2721 0 net=7980
rlabel metal2 184 -2721 184 -2721 0 net=1621
rlabel metal2 184 -2721 184 -2721 0 net=1621
rlabel metal2 198 -2721 198 -2721 0 net=1013
rlabel metal2 1783 -2721 1783 -2721 0 net=12614
rlabel metal2 58 -2723 58 -2723 0 net=5797
rlabel metal2 621 -2723 621 -2723 0 net=5451
rlabel metal2 775 -2723 775 -2723 0 net=11485
rlabel metal2 65 -2725 65 -2725 0 net=5693
rlabel metal2 1129 -2725 1129 -2725 0 net=3178
rlabel metal2 1297 -2725 1297 -2725 0 net=10575
rlabel metal2 100 -2727 100 -2727 0 net=2753
rlabel metal2 107 -2727 107 -2727 0 net=2076
rlabel metal2 534 -2727 534 -2727 0 net=6258
rlabel metal2 891 -2727 891 -2727 0 net=6156
rlabel metal2 1003 -2727 1003 -2727 0 net=6952
rlabel metal2 1328 -2727 1328 -2727 0 net=13428
rlabel metal2 100 -2729 100 -2729 0 net=1559
rlabel metal2 198 -2729 198 -2729 0 net=4097
rlabel metal2 275 -2729 275 -2729 0 net=1637
rlabel metal2 275 -2729 275 -2729 0 net=1637
rlabel metal2 289 -2729 289 -2729 0 net=2421
rlabel metal2 401 -2729 401 -2729 0 net=2508
rlabel metal2 425 -2729 425 -2729 0 net=8563
rlabel metal2 660 -2729 660 -2729 0 net=6943
rlabel metal2 919 -2729 919 -2729 0 net=9724
rlabel metal2 1297 -2729 1297 -2729 0 net=10703
rlabel metal2 1346 -2729 1346 -2729 0 net=10873
rlabel metal2 1675 -2729 1675 -2729 0 net=13415
rlabel metal2 107 -2731 107 -2731 0 net=3017
rlabel metal2 464 -2731 464 -2731 0 net=6274
rlabel metal2 1318 -2731 1318 -2731 0 net=12764
rlabel metal2 114 -2733 114 -2733 0 net=3719
rlabel metal2 114 -2733 114 -2733 0 net=3719
rlabel metal2 142 -2733 142 -2733 0 net=4897
rlabel metal2 842 -2733 842 -2733 0 net=6521
rlabel metal2 863 -2733 863 -2733 0 net=8054
rlabel metal2 1318 -2733 1318 -2733 0 net=11349
rlabel metal2 1605 -2733 1605 -2733 0 net=12801
rlabel metal2 149 -2735 149 -2735 0 net=2191
rlabel metal2 201 -2735 201 -2735 0 net=5992
rlabel metal2 292 -2735 292 -2735 0 net=3344
rlabel metal2 534 -2735 534 -2735 0 net=5333
rlabel metal2 849 -2735 849 -2735 0 net=9894
rlabel metal2 1325 -2735 1325 -2735 0 net=11195
rlabel metal2 1437 -2735 1437 -2735 0 net=12077
rlabel metal2 1626 -2735 1626 -2735 0 net=13003
rlabel metal2 205 -2737 205 -2737 0 net=1529
rlabel metal2 226 -2737 226 -2737 0 net=3431
rlabel metal2 436 -2737 436 -2737 0 net=5528
rlabel metal2 660 -2737 660 -2737 0 net=515
rlabel metal2 667 -2737 667 -2737 0 net=6747
rlabel metal2 1003 -2737 1003 -2737 0 net=8319
rlabel metal2 1080 -2737 1080 -2737 0 net=7342
rlabel metal2 1332 -2737 1332 -2737 0 net=8760
rlabel metal2 128 -2739 128 -2739 0 net=3189
rlabel metal2 226 -2739 226 -2739 0 net=4525
rlabel metal2 632 -2739 632 -2739 0 net=4751
rlabel metal2 705 -2739 705 -2739 0 net=10959
rlabel metal2 1346 -2739 1346 -2739 0 net=11013
rlabel metal2 1549 -2739 1549 -2739 0 net=12393
rlabel metal2 1647 -2739 1647 -2739 0 net=13243
rlabel metal2 1773 -2739 1773 -2739 0 net=11957
rlabel metal2 79 -2741 79 -2741 0 net=8597
rlabel metal2 170 -2741 170 -2741 0 net=7737
rlabel metal2 716 -2741 716 -2741 0 net=2712
rlabel metal2 863 -2741 863 -2741 0 net=9603
rlabel metal2 1241 -2741 1241 -2741 0 net=11137
rlabel metal2 1584 -2741 1584 -2741 0 net=12715
rlabel metal2 1682 -2741 1682 -2741 0 net=13479
rlabel metal2 61 -2743 61 -2743 0 net=11081
rlabel metal2 1237 -2743 1237 -2743 0 net=12831
rlabel metal2 79 -2745 79 -2745 0 net=4035
rlabel metal2 170 -2745 170 -2745 0 net=4437
rlabel metal2 436 -2745 436 -2745 0 net=6233
rlabel metal2 716 -2745 716 -2745 0 net=5619
rlabel metal2 852 -2745 852 -2745 0 net=5888
rlabel metal2 884 -2745 884 -2745 0 net=7298
rlabel metal2 1283 -2745 1283 -2745 0 net=636
rlabel metal2 37 -2747 37 -2747 0 net=6403
rlabel metal2 443 -2747 443 -2747 0 net=3923
rlabel metal2 562 -2747 562 -2747 0 net=3711
rlabel metal2 695 -2747 695 -2747 0 net=6815
rlabel metal2 877 -2747 877 -2747 0 net=5721
rlabel metal2 1388 -2747 1388 -2747 0 net=11213
rlabel metal2 37 -2749 37 -2749 0 net=8385
rlabel metal2 261 -2749 261 -2749 0 net=3167
rlabel metal2 9 -2751 9 -2751 0 net=4889
rlabel metal2 303 -2751 303 -2751 0 net=1908
rlabel metal2 884 -2751 884 -2751 0 net=6607
rlabel metal2 1080 -2751 1080 -2751 0 net=9153
rlabel metal2 1101 -2751 1101 -2751 0 net=9217
rlabel metal2 1101 -2751 1101 -2751 0 net=9217
rlabel metal2 1108 -2751 1108 -2751 0 net=9313
rlabel metal2 1108 -2751 1108 -2751 0 net=9313
rlabel metal2 1118 -2751 1118 -2751 0 net=12962
rlabel metal2 44 -2753 44 -2753 0 net=9933
rlabel metal2 303 -2753 303 -2753 0 net=3143
rlabel metal2 464 -2753 464 -2753 0 net=8963
rlabel metal2 919 -2753 919 -2753 0 net=7303
rlabel metal2 1010 -2753 1010 -2753 0 net=6956
rlabel metal2 1087 -2753 1087 -2753 0 net=5450
rlabel metal2 1661 -2753 1661 -2753 0 net=13693
rlabel metal2 268 -2755 268 -2755 0 net=2639
rlabel metal2 478 -2755 478 -2755 0 net=4058
rlabel metal2 513 -2755 513 -2755 0 net=3987
rlabel metal2 541 -2755 541 -2755 0 net=4451
rlabel metal2 611 -2755 611 -2755 0 net=5273
rlabel metal2 744 -2755 744 -2755 0 net=5671
rlabel metal2 940 -2755 940 -2755 0 net=10921
rlabel metal2 1720 -2755 1720 -2755 0 net=8007
rlabel metal2 135 -2757 135 -2757 0 net=1603
rlabel metal2 331 -2757 331 -2757 0 net=2084
rlabel metal2 569 -2757 569 -2757 0 net=4448
rlabel metal2 940 -2757 940 -2757 0 net=5837
rlabel metal2 1164 -2757 1164 -2757 0 net=9461
rlabel metal2 135 -2759 135 -2759 0 net=10279
rlabel metal2 310 -2759 310 -2759 0 net=6027
rlabel metal2 338 -2759 338 -2759 0 net=2767
rlabel metal2 527 -2759 527 -2759 0 net=4275
rlabel metal2 954 -2759 954 -2759 0 net=7107
rlabel metal2 982 -2759 982 -2759 0 net=9045
rlabel metal2 1013 -2759 1013 -2759 0 net=11679
rlabel metal2 51 -2761 51 -2761 0 net=7751
rlabel metal2 310 -2761 310 -2761 0 net=4147
rlabel metal2 1017 -2761 1017 -2761 0 net=13774
rlabel metal2 51 -2763 51 -2763 0 net=5437
rlabel metal2 562 -2763 562 -2763 0 net=5856
rlabel metal2 786 -2763 786 -2763 0 net=10625
rlabel metal2 1052 -2763 1052 -2763 0 net=8255
rlabel metal2 1094 -2763 1094 -2763 0 net=12181
rlabel metal2 1745 -2763 1745 -2763 0 net=13301
rlabel metal2 324 -2765 324 -2765 0 net=3672
rlabel metal2 866 -2765 866 -2765 0 net=12601
rlabel metal2 324 -2767 324 -2767 0 net=1747
rlabel metal2 355 -2767 355 -2767 0 net=1974
rlabel metal2 961 -2767 961 -2767 0 net=8545
rlabel metal2 1150 -2767 1150 -2767 0 net=13724
rlabel metal2 338 -2769 338 -2769 0 net=3203
rlabel metal2 569 -2769 569 -2769 0 net=4239
rlabel metal2 695 -2769 695 -2769 0 net=5569
rlabel metal2 821 -2769 821 -2769 0 net=5741
rlabel metal2 982 -2769 982 -2769 0 net=9321
rlabel metal2 1199 -2769 1199 -2769 0 net=11128
rlabel metal2 1633 -2769 1633 -2769 0 net=13531
rlabel metal2 345 -2771 345 -2771 0 net=2159
rlabel metal2 457 -2771 457 -2771 0 net=2651
rlabel metal2 1031 -2771 1031 -2771 0 net=8125
rlabel metal2 1073 -2771 1073 -2771 0 net=10475
rlabel metal2 1430 -2771 1430 -2771 0 net=11465
rlabel metal2 345 -2773 345 -2773 0 net=4919
rlabel metal2 1143 -2773 1143 -2773 0 net=9799
rlabel metal2 1276 -2773 1276 -2773 0 net=10913
rlabel metal2 1514 -2773 1514 -2773 0 net=12063
rlabel metal2 1633 -2773 1633 -2773 0 net=13031
rlabel metal2 380 -2775 380 -2775 0 net=2473
rlabel metal2 499 -2775 499 -2775 0 net=5407
rlabel metal2 751 -2775 751 -2775 0 net=10245
rlabel metal2 1311 -2775 1311 -2775 0 net=11707
rlabel metal2 1542 -2775 1542 -2775 0 net=12141
rlabel metal2 380 -2777 380 -2777 0 net=2673
rlabel metal2 478 -2777 478 -2777 0 net=3869
rlabel metal2 583 -2777 583 -2777 0 net=6600
rlabel metal2 1458 -2777 1458 -2777 0 net=11723
rlabel metal2 1556 -2777 1556 -2777 0 net=13269
rlabel metal2 408 -2779 408 -2779 0 net=3297
rlabel metal2 583 -2779 583 -2779 0 net=8325
rlabel metal2 807 -2779 807 -2779 0 net=6035
rlabel metal2 996 -2779 996 -2779 0 net=7777
rlabel metal2 1129 -2779 1129 -2779 0 net=13547
rlabel metal2 1696 -2779 1696 -2779 0 net=13545
rlabel metal2 415 -2781 415 -2781 0 net=2695
rlabel metal2 520 -2781 520 -2781 0 net=6779
rlabel metal2 1031 -2781 1031 -2781 0 net=11869
rlabel metal2 1500 -2781 1500 -2781 0 net=7865
rlabel metal2 415 -2783 415 -2783 0 net=3061
rlabel metal2 520 -2783 520 -2783 0 net=3797
rlabel metal2 590 -2783 590 -2783 0 net=4329
rlabel metal2 247 -2785 247 -2785 0 net=6225
rlabel metal2 597 -2785 597 -2785 0 net=5113
rlabel metal2 1150 -2785 1150 -2785 0 net=10367
rlabel metal2 1178 -2785 1178 -2785 0 net=12016
rlabel metal2 247 -2787 247 -2787 0 net=4665
rlabel metal2 548 -2787 548 -2787 0 net=3668
rlabel metal2 1171 -2787 1171 -2787 0 net=10143
rlabel metal2 1374 -2787 1374 -2787 0 net=11073
rlabel metal2 177 -2789 177 -2789 0 net=5487
rlabel metal2 607 -2789 607 -2789 0 net=5895
rlabel metal2 947 -2789 947 -2789 0 net=6603
rlabel metal2 1402 -2789 1402 -2789 0 net=11185
rlabel metal2 121 -2791 121 -2791 0 net=3473
rlabel metal2 296 -2791 296 -2791 0 net=5397
rlabel metal2 1402 -2791 1402 -2791 0 net=12447
rlabel metal2 121 -2793 121 -2793 0 net=2147
rlabel metal2 296 -2793 296 -2793 0 net=1859
rlabel metal2 1465 -2793 1465 -2793 0 net=11501
rlabel metal2 1591 -2793 1591 -2793 0 net=12733
rlabel metal2 212 -2795 212 -2795 0 net=4369
rlabel metal2 317 -2795 317 -2795 0 net=1993
rlabel metal2 471 -2795 471 -2795 0 net=3613
rlabel metal2 618 -2795 618 -2795 0 net=5134
rlabel metal2 1465 -2795 1465 -2795 0 net=11885
rlabel metal2 1619 -2795 1619 -2795 0 net=13329
rlabel metal2 212 -2797 212 -2797 0 net=1795
rlabel metal2 317 -2797 317 -2797 0 net=6861
rlabel metal2 1472 -2797 1472 -2797 0 net=11965
rlabel metal2 1703 -2797 1703 -2797 0 net=13643
rlabel metal2 254 -2799 254 -2799 0 net=2395
rlabel metal2 485 -2799 485 -2799 0 net=3387
rlabel metal2 618 -2799 618 -2799 0 net=6595
rlabel metal2 912 -2799 912 -2799 0 net=12241
rlabel metal2 163 -2801 163 -2801 0 net=3278
rlabel metal2 635 -2801 635 -2801 0 net=8043
rlabel metal2 975 -2801 975 -2801 0 net=12411
rlabel metal2 163 -2803 163 -2803 0 net=2277
rlabel metal2 254 -2803 254 -2803 0 net=6105
rlabel metal2 912 -2803 912 -2803 0 net=6451
rlabel metal2 975 -2803 975 -2803 0 net=7617
rlabel metal2 1185 -2803 1185 -2803 0 net=9817
rlabel metal2 1381 -2803 1381 -2803 0 net=10977
rlabel metal2 191 -2805 191 -2805 0 net=2609
rlabel metal2 681 -2805 681 -2805 0 net=7837
rlabel metal2 926 -2805 926 -2805 0 net=6905
rlabel metal2 1038 -2805 1038 -2805 0 net=8069
rlabel metal2 1255 -2805 1255 -2805 0 net=11245
rlabel metal2 1381 -2805 1381 -2805 0 net=11451
rlabel metal2 1479 -2805 1479 -2805 0 net=11987
rlabel metal2 450 -2807 450 -2807 0 net=3097
rlabel metal2 709 -2807 709 -2807 0 net=5925
rlabel metal2 968 -2807 968 -2807 0 net=8979
rlabel metal2 1087 -2807 1087 -2807 0 net=9073
rlabel metal2 1255 -2807 1255 -2807 0 net=10675
rlabel metal2 1444 -2807 1444 -2807 0 net=12957
rlabel metal2 394 -2809 394 -2809 0 net=3213
rlabel metal2 709 -2809 709 -2809 0 net=946
rlabel metal2 1024 -2809 1024 -2809 0 net=8021
rlabel metal2 1304 -2809 1304 -2809 0 net=11643
rlabel metal2 1528 -2809 1528 -2809 0 net=12277
rlabel metal2 1640 -2809 1640 -2809 0 net=13223
rlabel metal2 394 -2811 394 -2811 0 net=5057
rlabel metal2 1066 -2811 1066 -2811 0 net=10560
rlabel metal2 1367 -2811 1367 -2811 0 net=11161
rlabel metal2 1577 -2811 1577 -2811 0 net=12693
rlabel metal2 1668 -2811 1668 -2811 0 net=13403
rlabel metal2 674 -2813 674 -2813 0 net=4969
rlabel metal2 1020 -2813 1020 -2813 0 net=11549
rlabel metal2 1500 -2813 1500 -2813 0 net=9175
rlabel metal2 758 -2815 758 -2815 0 net=5251
rlabel metal2 1020 -2815 1020 -2815 0 net=687
rlabel metal2 1220 -2815 1220 -2815 0 net=9839
rlabel metal2 1535 -2815 1535 -2815 0 net=12045
rlabel metal2 800 -2817 800 -2817 0 net=6623
rlabel metal2 1136 -2817 1136 -2817 0 net=8919
rlabel metal2 1409 -2817 1409 -2817 0 net=12309
rlabel metal2 814 -2819 814 -2819 0 net=9347
rlabel metal2 1136 -2819 1136 -2819 0 net=10057
rlabel metal2 1409 -2819 1409 -2819 0 net=11601
rlabel metal2 814 -2821 814 -2821 0 net=3479
rlabel metal2 905 -2823 905 -2823 0 net=10745
rlabel metal2 898 -2825 898 -2825 0 net=6727
rlabel metal2 1157 -2825 1157 -2825 0 net=9631
rlabel metal2 733 -2827 733 -2827 0 net=7313
rlabel metal2 1122 -2827 1122 -2827 0 net=9265
rlabel metal2 23 -2838 23 -2838 0 net=2423
rlabel metal2 331 -2838 331 -2838 0 net=6028
rlabel metal2 621 -2838 621 -2838 0 net=11870
rlabel metal2 1097 -2838 1097 -2838 0 net=13404
rlabel metal2 1713 -2838 1713 -2838 0 net=13302
rlabel metal2 44 -2840 44 -2840 0 net=9934
rlabel metal2 656 -2840 656 -2840 0 net=10746
rlabel metal2 1433 -2840 1433 -2840 0 net=13532
rlabel metal2 1717 -2840 1717 -2840 0 net=11958
rlabel metal2 79 -2842 79 -2842 0 net=4037
rlabel metal2 660 -2842 660 -2842 0 net=10246
rlabel metal2 1283 -2842 1283 -2842 0 net=13416
rlabel metal2 1720 -2842 1720 -2842 0 net=11186
rlabel metal2 93 -2844 93 -2844 0 net=9697
rlabel metal2 1339 -2844 1339 -2844 0 net=12833
rlabel metal2 1654 -2844 1654 -2844 0 net=13549
rlabel metal2 1727 -2844 1727 -2844 0 net=8008
rlabel metal2 93 -2846 93 -2846 0 net=2149
rlabel metal2 128 -2846 128 -2846 0 net=8598
rlabel metal2 859 -2846 859 -2846 0 net=13546
rlabel metal2 96 -2848 96 -2848 0 net=202
rlabel metal2 712 -2848 712 -2848 0 net=10626
rlabel metal2 824 -2848 824 -2848 0 net=11486
rlabel metal2 1549 -2848 1549 -2848 0 net=12395
rlabel metal2 1549 -2848 1549 -2848 0 net=12395
rlabel metal2 1598 -2848 1598 -2848 0 net=12047
rlabel metal2 100 -2850 100 -2850 0 net=1560
rlabel metal2 681 -2850 681 -2850 0 net=7839
rlabel metal2 1013 -2850 1013 -2850 0 net=11214
rlabel metal2 1465 -2850 1465 -2850 0 net=11887
rlabel metal2 1591 -2850 1591 -2850 0 net=12735
rlabel metal2 1647 -2850 1647 -2850 0 net=13245
rlabel metal2 37 -2852 37 -2852 0 net=8387
rlabel metal2 730 -2852 730 -2852 0 net=5723
rlabel metal2 915 -2852 915 -2852 0 net=10960
rlabel metal2 1342 -2852 1342 -2852 0 net=11502
rlabel metal2 1640 -2852 1640 -2852 0 net=13225
rlabel metal2 51 -2854 51 -2854 0 net=5439
rlabel metal2 107 -2854 107 -2854 0 net=3018
rlabel metal2 870 -2854 870 -2854 0 net=6728
rlabel metal2 947 -2854 947 -2854 0 net=8045
rlabel metal2 1024 -2854 1024 -2854 0 net=8022
rlabel metal2 1150 -2854 1150 -2854 0 net=10369
rlabel metal2 1353 -2854 1353 -2854 0 net=13480
rlabel metal2 51 -2856 51 -2856 0 net=4167
rlabel metal2 107 -2856 107 -2856 0 net=9266
rlabel metal2 1178 -2856 1178 -2856 0 net=13644
rlabel metal2 72 -2858 72 -2858 0 net=1749
rlabel metal2 359 -2858 359 -2858 0 net=6405
rlabel metal2 765 -2858 765 -2858 0 net=5927
rlabel metal2 877 -2858 877 -2858 0 net=6675
rlabel metal2 1024 -2858 1024 -2858 0 net=12064
rlabel metal2 1661 -2858 1661 -2858 0 net=13695
rlabel metal2 1703 -2858 1703 -2858 0 net=1124
rlabel metal2 121 -2860 121 -2860 0 net=2611
rlabel metal2 226 -2860 226 -2860 0 net=4527
rlabel metal2 366 -2860 366 -2860 0 net=2640
rlabel metal2 499 -2860 499 -2860 0 net=3871
rlabel metal2 499 -2860 499 -2860 0 net=3871
rlabel metal2 520 -2860 520 -2860 0 net=3798
rlabel metal2 1101 -2860 1101 -2860 0 net=9219
rlabel metal2 1199 -2860 1199 -2860 0 net=10914
rlabel metal2 1353 -2860 1353 -2860 0 net=11075
rlabel metal2 1381 -2860 1381 -2860 0 net=11453
rlabel metal2 1444 -2860 1444 -2860 0 net=12959
rlabel metal2 1640 -2860 1640 -2860 0 net=13345
rlabel metal2 65 -2862 65 -2862 0 net=5695
rlabel metal2 555 -2862 555 -2862 0 net=8126
rlabel metal2 1066 -2862 1066 -2862 0 net=8351
rlabel metal2 1115 -2862 1115 -2862 0 net=9462
rlabel metal2 1202 -2862 1202 -2862 0 net=10874
rlabel metal2 1514 -2862 1514 -2862 0 net=12279
rlabel metal2 65 -2864 65 -2864 0 net=3169
rlabel metal2 275 -2864 275 -2864 0 net=1638
rlabel metal2 366 -2864 366 -2864 0 net=2675
rlabel metal2 429 -2864 429 -2864 0 net=1995
rlabel metal2 464 -2864 464 -2864 0 net=8965
rlabel metal2 1227 -2864 1227 -2864 0 net=6605
rlabel metal2 128 -2866 128 -2866 0 net=2175
rlabel metal2 247 -2866 247 -2866 0 net=4666
rlabel metal2 1066 -2866 1066 -2866 0 net=8437
rlabel metal2 1237 -2866 1237 -2866 0 net=9176
rlabel metal2 135 -2868 135 -2868 0 net=10280
rlabel metal2 429 -2868 429 -2868 0 net=4453
rlabel metal2 555 -2868 555 -2868 0 net=4689
rlabel metal2 674 -2868 674 -2868 0 net=4971
rlabel metal2 1125 -2868 1125 -2868 0 net=12142
rlabel metal2 142 -2870 142 -2870 0 net=4899
rlabel metal2 737 -2870 737 -2870 0 net=5453
rlabel metal2 779 -2870 779 -2870 0 net=6817
rlabel metal2 954 -2870 954 -2870 0 net=7109
rlabel metal2 954 -2870 954 -2870 0 net=7109
rlabel metal2 968 -2870 968 -2870 0 net=8981
rlabel metal2 1136 -2870 1136 -2870 0 net=10059
rlabel metal2 1311 -2870 1311 -2870 0 net=11709
rlabel metal2 1500 -2870 1500 -2870 0 net=12243
rlabel metal2 1535 -2870 1535 -2870 0 net=12311
rlabel metal2 86 -2872 86 -2872 0 net=4890
rlabel metal2 145 -2872 145 -2872 0 net=11483
rlabel metal2 86 -2874 86 -2874 0 net=3721
rlabel metal2 170 -2874 170 -2874 0 net=4438
rlabel metal2 604 -2874 604 -2874 0 net=8565
rlabel metal2 1164 -2874 1164 -2874 0 net=10145
rlabel metal2 1227 -2874 1227 -2874 0 net=7867
rlabel metal2 58 -2876 58 -2876 0 net=5799
rlabel metal2 156 -2876 156 -2876 0 net=2193
rlabel metal2 226 -2876 226 -2876 0 net=138
rlabel metal2 471 -2876 471 -2876 0 net=3615
rlabel metal2 471 -2876 471 -2876 0 net=3615
rlabel metal2 562 -2876 562 -2876 0 net=12647
rlabel metal2 58 -2878 58 -2878 0 net=4039
rlabel metal2 786 -2878 786 -2878 0 net=5579
rlabel metal2 1171 -2878 1171 -2878 0 net=11551
rlabel metal2 1437 -2878 1437 -2878 0 net=12079
rlabel metal2 156 -2880 156 -2880 0 net=1623
rlabel metal2 240 -2880 240 -2880 0 net=4371
rlabel metal2 254 -2880 254 -2880 0 net=6106
rlabel metal2 971 -2880 971 -2880 0 net=10704
rlabel metal2 1311 -2880 1311 -2880 0 net=10845
rlabel metal2 149 -2882 149 -2882 0 net=2755
rlabel metal2 261 -2882 261 -2882 0 net=3433
rlabel metal2 380 -2882 380 -2882 0 net=3119
rlabel metal2 576 -2882 576 -2882 0 net=6227
rlabel metal2 646 -2882 646 -2882 0 net=6781
rlabel metal2 821 -2882 821 -2882 0 net=6037
rlabel metal2 982 -2882 982 -2882 0 net=9323
rlabel metal2 1234 -2882 1234 -2882 0 net=11645
rlabel metal2 1318 -2882 1318 -2882 0 net=11351
rlabel metal2 1423 -2882 1423 -2882 0 net=11681
rlabel metal2 1444 -2882 1444 -2882 0 net=12695
rlabel metal2 149 -2884 149 -2884 0 net=3205
rlabel metal2 373 -2884 373 -2884 0 net=2475
rlabel metal2 394 -2884 394 -2884 0 net=5058
rlabel metal2 562 -2884 562 -2884 0 net=4241
rlabel metal2 576 -2884 576 -2884 0 net=1773
rlabel metal2 898 -2884 898 -2884 0 net=7315
rlabel metal2 989 -2884 989 -2884 0 net=9047
rlabel metal2 1255 -2884 1255 -2884 0 net=10677
rlabel metal2 1318 -2884 1318 -2884 0 net=10979
rlabel metal2 184 -2886 184 -2886 0 net=5409
rlabel metal2 667 -2886 667 -2886 0 net=6749
rlabel metal2 933 -2886 933 -2886 0 net=9349
rlabel metal2 1479 -2886 1479 -2886 0 net=11989
rlabel metal2 1570 -2886 1570 -2886 0 net=12603
rlabel metal2 233 -2888 233 -2888 0 net=7753
rlabel metal2 394 -2888 394 -2888 0 net=2161
rlabel metal2 590 -2888 590 -2888 0 net=4331
rlabel metal2 625 -2888 625 -2888 0 net=5319
rlabel metal2 1143 -2888 1143 -2888 0 net=9801
rlabel metal2 1262 -2888 1262 -2888 0 net=11247
rlabel metal2 1458 -2888 1458 -2888 0 net=11725
rlabel metal2 1486 -2888 1486 -2888 0 net=12413
rlabel metal2 1570 -2888 1570 -2888 0 net=12717
rlabel metal2 233 -2890 233 -2890 0 net=1843
rlabel metal2 1185 -2890 1185 -2890 0 net=9819
rlabel metal2 1269 -2890 1269 -2890 0 net=8921
rlabel metal2 1325 -2890 1325 -2890 0 net=11197
rlabel metal2 1409 -2890 1409 -2890 0 net=11603
rlabel metal2 240 -2892 240 -2892 0 net=1605
rlabel metal2 275 -2892 275 -2892 0 net=3481
rlabel metal2 828 -2892 828 -2892 0 net=5743
rlabel metal2 849 -2892 849 -2892 0 net=10576
rlabel metal2 1367 -2892 1367 -2892 0 net=11163
rlabel metal2 1472 -2892 1472 -2892 0 net=11967
rlabel metal2 268 -2894 268 -2894 0 net=3713
rlabel metal2 653 -2894 653 -2894 0 net=7739
rlabel metal2 1185 -2894 1185 -2894 0 net=9633
rlabel metal2 1213 -2894 1213 -2894 0 net=11083
rlabel metal2 1472 -2894 1472 -2894 0 net=11809
rlabel metal2 282 -2896 282 -2896 0 net=2397
rlabel metal2 415 -2896 415 -2896 0 net=3063
rlabel metal2 439 -2896 439 -2896 0 net=8959
rlabel metal2 198 -2898 198 -2898 0 net=4099
rlabel metal2 527 -2898 527 -2898 0 net=4277
rlabel metal2 590 -2898 590 -2898 0 net=5621
rlabel metal2 737 -2898 737 -2898 0 net=5839
rlabel metal2 1059 -2898 1059 -2898 0 net=7779
rlabel metal2 1220 -2898 1220 -2898 0 net=9841
rlabel metal2 1325 -2898 1325 -2898 0 net=11015
rlabel metal2 1356 -2898 1356 -2898 0 net=13330
rlabel metal2 110 -2900 110 -2900 0 net=9429
rlabel metal2 751 -2900 751 -2900 0 net=6597
rlabel metal2 1052 -2900 1052 -2900 0 net=8257
rlabel metal2 1069 -2900 1069 -2900 0 net=11751
rlabel metal2 198 -2902 198 -2902 0 net=1531
rlabel metal2 212 -2902 212 -2902 0 net=1797
rlabel metal2 289 -2902 289 -2902 0 net=4149
rlabel metal2 317 -2902 317 -2902 0 net=6863
rlabel metal2 1052 -2902 1052 -2902 0 net=13270
rlabel metal2 163 -2904 163 -2904 0 net=2278
rlabel metal2 212 -2904 212 -2904 0 net=2131
rlabel metal2 1290 -2904 1290 -2904 0 net=11057
rlabel metal2 1402 -2904 1402 -2904 0 net=12449
rlabel metal2 163 -2906 163 -2906 0 net=8637
rlabel metal2 1206 -2906 1206 -2906 0 net=10923
rlabel metal2 303 -2908 303 -2908 0 net=3145
rlabel metal2 324 -2908 324 -2908 0 net=2769
rlabel metal2 506 -2908 506 -2908 0 net=2697
rlabel metal2 653 -2908 653 -2908 0 net=13379
rlabel metal2 208 -2910 208 -2910 0 net=4005
rlabel metal2 310 -2910 310 -2910 0 net=2653
rlabel metal2 506 -2910 506 -2910 0 net=5115
rlabel metal2 663 -2910 663 -2910 0 net=5121
rlabel metal2 835 -2910 835 -2910 0 net=9075
rlabel metal2 1094 -2910 1094 -2910 0 net=12183
rlabel metal2 219 -2912 219 -2912 0 net=3191
rlabel metal2 667 -2912 667 -2912 0 net=3585
rlabel metal2 1073 -2912 1073 -2912 0 net=10477
rlabel metal2 1402 -2912 1402 -2912 0 net=11467
rlabel metal2 219 -2914 219 -2914 0 net=238
rlabel metal2 1038 -2914 1038 -2914 0 net=8071
rlabel metal2 1080 -2914 1080 -2914 0 net=9155
rlabel metal2 1241 -2914 1241 -2914 0 net=11139
rlabel metal2 338 -2916 338 -2916 0 net=3299
rlabel metal2 436 -2916 436 -2916 0 net=6235
rlabel metal2 674 -2916 674 -2916 0 net=4607
rlabel metal2 891 -2916 891 -2916 0 net=6945
rlabel metal2 191 -2918 191 -2918 0 net=1673
rlabel metal2 688 -2918 688 -2918 0 net=5399
rlabel metal2 800 -2918 800 -2918 0 net=6625
rlabel metal2 961 -2918 961 -2918 0 net=8547
rlabel metal2 331 -2920 331 -2920 0 net=3123
rlabel metal2 926 -2920 926 -2920 0 net=6907
rlabel metal2 975 -2920 975 -2920 0 net=7619
rlabel metal2 1108 -2920 1108 -2920 0 net=9315
rlabel metal2 345 -2922 345 -2922 0 net=4921
rlabel metal2 688 -2922 688 -2922 0 net=5007
rlabel metal2 1108 -2922 1108 -2922 0 net=8355
rlabel metal2 177 -2924 177 -2924 0 net=3475
rlabel metal2 401 -2924 401 -2924 0 net=3215
rlabel metal2 695 -2924 695 -2924 0 net=5571
rlabel metal2 807 -2924 807 -2924 0 net=6609
rlabel metal2 919 -2924 919 -2924 0 net=7305
rlabel metal2 1003 -2924 1003 -2924 0 net=8321
rlabel metal2 1430 -2924 1430 -2924 0 net=12803
rlabel metal2 177 -2926 177 -2926 0 net=3389
rlabel metal2 534 -2926 534 -2926 0 net=5335
rlabel metal2 723 -2926 723 -2926 0 net=8327
rlabel metal2 1605 -2926 1605 -2926 0 net=13005
rlabel metal2 443 -2928 443 -2928 0 net=3925
rlabel metal2 485 -2928 485 -2928 0 net=11769
rlabel metal2 723 -2928 723 -2928 0 net=5253
rlabel metal2 793 -2928 793 -2928 0 net=5897
rlabel metal2 926 -2928 926 -2928 0 net=5631
rlabel metal2 1626 -2928 1626 -2928 0 net=13033
rlabel metal2 443 -2930 443 -2930 0 net=3989
rlabel metal2 733 -2930 733 -2930 0 net=13107
rlabel metal2 478 -2932 478 -2932 0 net=1981
rlabel metal2 744 -2932 744 -2932 0 net=5673
rlabel metal2 842 -2932 842 -2932 0 net=6523
rlabel metal2 478 -2934 478 -2934 0 net=3809
rlabel metal2 492 -2936 492 -2936 0 net=3098
rlabel metal2 611 -2936 611 -2936 0 net=5275
rlabel metal2 758 -2936 758 -2936 0 net=4813
rlabel metal2 863 -2936 863 -2936 0 net=9605
rlabel metal2 492 -2938 492 -2938 0 net=4207
rlabel metal2 663 -2938 663 -2938 0 net=4565
rlabel metal2 863 -2938 863 -2938 0 net=9679
rlabel metal2 548 -2940 548 -2940 0 net=5489
rlabel metal2 884 -2940 884 -2940 0 net=6453
rlabel metal2 82 -2942 82 -2942 0 net=3289
rlabel metal2 611 -2942 611 -2942 0 net=4753
rlabel metal2 912 -2942 912 -2942 0 net=11863
rlabel metal2 296 -2944 296 -2944 0 net=1861
rlabel metal2 166 -2946 166 -2946 0 net=7517
rlabel metal2 30 -2957 30 -2957 0 net=2151
rlabel metal2 100 -2957 100 -2957 0 net=5441
rlabel metal2 439 -2957 439 -2957 0 net=5122
rlabel metal2 821 -2957 821 -2957 0 net=5929
rlabel metal2 863 -2957 863 -2957 0 net=11604
rlabel metal2 1640 -2957 1640 -2957 0 net=12048
rlabel metal2 37 -2959 37 -2959 0 net=4151
rlabel metal2 303 -2959 303 -2959 0 net=4007
rlabel metal2 369 -2959 369 -2959 0 net=1225
rlabel metal2 541 -2959 541 -2959 0 net=1996
rlabel metal2 663 -2959 663 -2959 0 net=6946
rlabel metal2 1332 -2959 1332 -2959 0 net=11888
rlabel metal2 1577 -2959 1577 -2959 0 net=12604
rlabel metal2 44 -2961 44 -2961 0 net=2163
rlabel metal2 450 -2961 450 -2961 0 net=3927
rlabel metal2 548 -2961 548 -2961 0 net=3291
rlabel metal2 842 -2961 842 -2961 0 net=4566
rlabel metal2 1027 -2961 1027 -2961 0 net=6606
rlabel metal2 23 -2963 23 -2963 0 net=2424
rlabel metal2 499 -2963 499 -2963 0 net=3873
rlabel metal2 611 -2963 611 -2963 0 net=4755
rlabel metal2 674 -2963 674 -2963 0 net=4608
rlabel metal2 1020 -2963 1020 -2963 0 net=9316
rlabel metal2 1332 -2963 1332 -2963 0 net=11199
rlabel metal2 1458 -2963 1458 -2963 0 net=11753
rlabel metal2 72 -2965 72 -2965 0 net=1750
rlabel metal2 499 -2965 499 -2965 0 net=5009
rlabel metal2 740 -2965 740 -2965 0 net=7740
rlabel metal2 1171 -2965 1171 -2965 0 net=11553
rlabel metal2 1458 -2965 1458 -2965 0 net=11865
rlabel metal2 1577 -2965 1577 -2965 0 net=13007
rlabel metal2 51 -2967 51 -2967 0 net=4169
rlabel metal2 79 -2967 79 -2967 0 net=3192
rlabel metal2 569 -2967 569 -2967 0 net=4279
rlabel metal2 618 -2967 618 -2967 0 net=6229
rlabel metal2 849 -2967 849 -2967 0 net=4972
rlabel metal2 1150 -2967 1150 -2967 0 net=9221
rlabel metal2 1199 -2967 1199 -2967 0 net=12080
rlabel metal2 1605 -2967 1605 -2967 0 net=13227
rlabel metal2 51 -2969 51 -2969 0 net=2133
rlabel metal2 219 -2969 219 -2969 0 net=7840
rlabel metal2 1010 -2969 1010 -2969 0 net=9049
rlabel metal2 1199 -2969 1199 -2969 0 net=9681
rlabel metal2 1339 -2969 1339 -2969 0 net=12835
rlabel metal2 1647 -2969 1647 -2969 0 net=13697
rlabel metal2 65 -2971 65 -2971 0 net=3171
rlabel metal2 261 -2971 261 -2971 0 net=3434
rlabel metal2 408 -2971 408 -2971 0 net=4463
rlabel metal2 492 -2971 492 -2971 0 net=4209
rlabel metal2 604 -2971 604 -2971 0 net=4332
rlabel metal2 674 -2971 674 -2971 0 net=5675
rlabel metal2 835 -2971 835 -2971 0 net=9077
rlabel metal2 1164 -2971 1164 -2971 0 net=10147
rlabel metal2 1339 -2971 1339 -2971 0 net=11249
rlabel metal2 1465 -2971 1465 -2971 0 net=11969
rlabel metal2 65 -2973 65 -2973 0 net=5889
rlabel metal2 261 -2973 261 -2973 0 net=1983
rlabel metal2 604 -2973 604 -2973 0 net=4815
rlabel metal2 782 -2973 782 -2973 0 net=12414
rlabel metal2 82 -2975 82 -2975 0 net=8966
rlabel metal2 1213 -2975 1213 -2975 0 net=9803
rlabel metal2 1297 -2975 1297 -2975 0 net=10679
rlabel metal2 1486 -2975 1486 -2975 0 net=12185
rlabel metal2 1535 -2975 1535 -2975 0 net=12649
rlabel metal2 93 -2977 93 -2977 0 net=4243
rlabel metal2 793 -2977 793 -2977 0 net=5633
rlabel metal2 943 -2977 943 -2977 0 net=11454
rlabel metal2 1430 -2977 1430 -2977 0 net=12805
rlabel metal2 79 -2979 79 -2979 0 net=11759
rlabel metal2 1430 -2979 1430 -2979 0 net=13381
rlabel metal2 100 -2981 100 -2981 0 net=5891
rlabel metal2 835 -2981 835 -2981 0 net=6864
rlabel metal2 996 -2981 996 -2981 0 net=7621
rlabel metal2 1052 -2981 1052 -2981 0 net=8259
rlabel metal2 1094 -2981 1094 -2981 0 net=10981
rlabel metal2 1493 -2981 1493 -2981 0 net=12281
rlabel metal2 107 -2983 107 -2983 0 net=7929
rlabel metal2 1031 -2983 1031 -2983 0 net=12960
rlabel metal2 107 -2985 107 -2985 0 net=3991
rlabel metal2 562 -2985 562 -2985 0 net=3511
rlabel metal2 891 -2985 891 -2985 0 net=6525
rlabel metal2 891 -2985 891 -2985 0 net=6525
rlabel metal2 901 -2985 901 -2985 0 net=9350
rlabel metal2 1514 -2985 1514 -2985 0 net=12397
rlabel metal2 1591 -2985 1591 -2985 0 net=13109
rlabel metal2 110 -2987 110 -2987 0 net=2756
rlabel metal2 268 -2987 268 -2987 0 net=3714
rlabel metal2 1115 -2987 1115 -2987 0 net=8567
rlabel metal2 1136 -2987 1136 -2987 0 net=9325
rlabel metal2 1202 -2987 1202 -2987 0 net=11757
rlabel metal2 121 -2989 121 -2989 0 net=2612
rlabel metal2 660 -2989 660 -2989 0 net=5725
rlabel metal2 849 -2989 849 -2989 0 net=6455
rlabel metal2 905 -2989 905 -2989 0 net=6627
rlabel metal2 905 -2989 905 -2989 0 net=6627
rlabel metal2 926 -2989 926 -2989 0 net=6819
rlabel metal2 982 -2989 982 -2989 0 net=7317
rlabel metal2 1045 -2989 1045 -2989 0 net=8983
rlabel metal2 1136 -2989 1136 -2989 0 net=11085
rlabel metal2 1423 -2989 1423 -2989 0 net=13551
rlabel metal2 82 -2991 82 -2991 0 net=8219
rlabel metal2 1055 -2991 1055 -2991 0 net=11990
rlabel metal2 1549 -2991 1549 -2991 0 net=12719
rlabel metal2 121 -2993 121 -2993 0 net=2399
rlabel metal2 408 -2993 408 -2993 0 net=4101
rlabel metal2 443 -2993 443 -2993 0 net=3587
rlabel metal2 852 -2993 852 -2993 0 net=5898
rlabel metal2 947 -2993 947 -2993 0 net=7110
rlabel metal2 989 -2993 989 -2993 0 net=8073
rlabel metal2 1122 -2993 1122 -2993 0 net=9157
rlabel metal2 1220 -2993 1220 -2993 0 net=9821
rlabel metal2 1297 -2993 1297 -2993 0 net=11077
rlabel metal2 1521 -2993 1521 -2993 0 net=12451
rlabel metal2 1570 -2993 1570 -2993 0 net=12737
rlabel metal2 89 -2995 89 -2995 0 net=8741
rlabel metal2 1255 -2995 1255 -2995 0 net=10479
rlabel metal2 1318 -2995 1318 -2995 0 net=11141
rlabel metal2 1598 -2995 1598 -2995 0 net=13035
rlabel metal2 142 -2997 142 -2997 0 net=7519
rlabel metal2 1010 -2997 1010 -2997 0 net=7869
rlabel metal2 1262 -2997 1262 -2997 0 net=10847
rlabel metal2 1367 -2997 1367 -2997 0 net=11353
rlabel metal2 1626 -2997 1626 -2997 0 net=13347
rlabel metal2 145 -2999 145 -2999 0 net=4038
rlabel metal2 632 -2999 632 -2999 0 net=1863
rlabel metal2 856 -2999 856 -2999 0 net=6039
rlabel metal2 877 -2999 877 -2999 0 net=6677
rlabel metal2 954 -2999 954 -2999 0 net=6909
rlabel metal2 968 -2999 968 -2999 0 net=8509
rlabel metal2 1227 -2999 1227 -2999 0 net=11059
rlabel metal2 156 -3001 156 -3001 0 net=1625
rlabel metal2 268 -3001 268 -3001 0 net=3121
rlabel metal2 415 -3001 415 -3001 0 net=3065
rlabel metal2 506 -3001 506 -3001 0 net=5117
rlabel metal2 156 -3003 156 -3003 0 net=5581
rlabel metal2 880 -3003 880 -3003 0 net=6753
rlabel metal2 163 -3005 163 -3005 0 net=6598
rlabel metal2 961 -3005 961 -3005 0 net=7199
rlabel metal2 1346 -3005 1346 -3005 0 net=11263
rlabel metal2 86 -3007 86 -3007 0 net=3723
rlabel metal2 170 -3007 170 -3007 0 net=2194
rlabel metal2 282 -3007 282 -3007 0 net=1799
rlabel metal2 401 -3007 401 -3007 0 net=3217
rlabel metal2 583 -3007 583 -3007 0 net=4075
rlabel metal2 968 -3007 968 -3007 0 net=7307
rlabel metal2 1017 -3007 1017 -3007 0 net=8047
rlabel metal2 1034 -3007 1034 -3007 0 net=11484
rlabel metal2 86 -3009 86 -3009 0 net=10924
rlabel metal2 128 -3011 128 -3011 0 net=2177
rlabel metal2 275 -3011 275 -3011 0 net=3483
rlabel metal2 289 -3011 289 -3011 0 net=1775
rlabel metal2 632 -3011 632 -3011 0 net=6177
rlabel metal2 884 -3011 884 -3011 0 net=8357
rlabel metal2 1234 -3011 1234 -3011 0 net=11647
rlabel metal2 1612 -3011 1612 -3011 0 net=13247
rlabel metal2 58 -3013 58 -3013 0 net=4041
rlabel metal2 639 -3013 639 -3013 0 net=4923
rlabel metal2 702 -3013 702 -3013 0 net=4900
rlabel metal2 898 -3013 898 -3013 0 net=6751
rlabel metal2 1059 -3013 1059 -3013 0 net=8329
rlabel metal2 1108 -3013 1108 -3013 0 net=8549
rlabel metal2 1234 -3013 1234 -3013 0 net=10061
rlabel metal2 58 -3015 58 -3015 0 net=1352
rlabel metal2 138 -3015 138 -3015 0 net=1649
rlabel metal2 303 -3015 303 -3015 0 net=3811
rlabel metal2 513 -3015 513 -3015 0 net=3853
rlabel metal2 1192 -3015 1192 -3015 0 net=7781
rlabel metal2 128 -3017 128 -3017 0 net=5337
rlabel metal2 702 -3017 702 -3017 0 net=5255
rlabel metal2 789 -3017 789 -3017 0 net=11283
rlabel metal2 1185 -3017 1185 -3017 0 net=9635
rlabel metal2 1206 -3017 1206 -3017 0 net=9699
rlabel metal2 170 -3019 170 -3019 0 net=1675
rlabel metal2 205 -3019 205 -3019 0 net=7518
rlabel metal2 317 -3019 317 -3019 0 net=3147
rlabel metal2 478 -3019 478 -3019 0 net=4691
rlabel metal2 639 -3019 639 -3019 0 net=6783
rlabel metal2 656 -3019 656 -3019 0 net=11023
rlabel metal2 61 -3021 61 -3021 0 net=3039
rlabel metal2 646 -3021 646 -3021 0 net=8353
rlabel metal2 1248 -3021 1248 -3021 0 net=10371
rlabel metal2 177 -3023 177 -3023 0 net=3390
rlabel metal2 709 -3023 709 -3023 0 net=6407
rlabel metal2 898 -3023 898 -3023 0 net=8438
rlabel metal2 1283 -3023 1283 -3023 0 net=11017
rlabel metal2 177 -3025 177 -3025 0 net=2477
rlabel metal2 401 -3025 401 -3025 0 net=4455
rlabel metal2 681 -3025 681 -3025 0 net=8389
rlabel metal2 1325 -3025 1325 -3025 0 net=11165
rlabel metal2 114 -3027 114 -3027 0 net=5801
rlabel metal2 464 -3027 464 -3027 0 net=5223
rlabel metal2 688 -3027 688 -3027 0 net=8507
rlabel metal2 1374 -3027 1374 -3027 0 net=11469
rlabel metal2 149 -3029 149 -3029 0 net=3207
rlabel metal2 709 -3029 709 -3029 0 net=5401
rlabel metal2 912 -3029 912 -3029 0 net=12725
rlabel metal2 149 -3031 149 -3031 0 net=8638
rlabel metal2 1304 -3031 1304 -3031 0 net=8923
rlabel metal2 187 -3033 187 -3033 0 net=12487
rlabel metal2 191 -3035 191 -3035 0 net=1533
rlabel metal2 205 -3035 205 -3035 0 net=7754
rlabel metal2 716 -3035 716 -3035 0 net=9431
rlabel metal2 1269 -3035 1269 -3035 0 net=9843
rlabel metal2 310 -3037 310 -3037 0 net=2655
rlabel metal2 338 -3037 338 -3037 0 net=3301
rlabel metal2 387 -3037 387 -3037 0 net=2699
rlabel metal2 716 -3037 716 -3037 0 net=5277
rlabel metal2 751 -3037 751 -3037 0 net=5491
rlabel metal2 1003 -3037 1003 -3037 0 net=9607
rlabel metal2 1269 -3037 1269 -3037 0 net=11683
rlabel metal2 184 -3039 184 -3039 0 net=5411
rlabel metal2 1066 -3039 1066 -3039 0 net=8323
rlabel metal2 184 -3041 184 -3041 0 net=5572
rlabel metal2 1080 -3041 1080 -3041 0 net=8960
rlabel metal2 310 -3043 310 -3043 0 net=5321
rlabel metal2 723 -3043 723 -3043 0 net=7235
rlabel metal2 800 -3043 800 -3043 0 net=13275
rlabel metal2 324 -3045 324 -3045 0 net=2771
rlabel metal2 345 -3045 345 -3045 0 net=3477
rlabel metal2 1409 -3045 1409 -3045 0 net=11711
rlabel metal2 324 -3047 324 -3047 0 net=3125
rlabel metal2 345 -3047 345 -3047 0 net=11455
rlabel metal2 786 -3047 786 -3047 0 net=11889
rlabel metal2 331 -3049 331 -3049 0 net=2677
rlabel metal2 485 -3049 485 -3049 0 net=11771
rlabel metal2 114 -3051 114 -3051 0 net=2583
rlabel metal2 485 -3051 485 -3051 0 net=5623
rlabel metal2 352 -3053 352 -3053 0 net=4529
rlabel metal2 520 -3053 520 -3053 0 net=5697
rlabel metal2 152 -3055 152 -3055 0 net=2841
rlabel metal2 359 -3055 359 -3055 0 net=3225
rlabel metal2 590 -3055 590 -3055 0 net=2997
rlabel metal2 471 -3057 471 -3057 0 net=3617
rlabel metal2 527 -3057 527 -3057 0 net=5455
rlabel metal2 915 -3057 915 -3057 0 net=11726
rlabel metal2 471 -3059 471 -3059 0 net=5841
rlabel metal2 765 -3059 765 -3059 0 net=6611
rlabel metal2 1479 -3059 1479 -3059 0 net=12245
rlabel metal2 534 -3061 534 -3061 0 net=7697
rlabel metal2 1500 -3061 1500 -3061 0 net=12313
rlabel metal2 233 -3063 233 -3063 0 net=1845
rlabel metal2 737 -3063 737 -3063 0 net=11587
rlabel metal2 1444 -3063 1444 -3063 0 net=12697
rlabel metal2 233 -3065 233 -3065 0 net=1607
rlabel metal2 807 -3065 807 -3065 0 net=5745
rlabel metal2 1444 -3065 1444 -3065 0 net=11811
rlabel metal2 240 -3067 240 -3067 0 net=4373
rlabel metal2 828 -3067 828 -3067 0 net=12439
rlabel metal2 247 -3069 247 -3069 0 net=1505
rlabel metal2 831 -3069 831 -3069 0 net=12099
rlabel metal2 597 -3071 597 -3071 0 net=6237
rlabel metal2 597 -3073 597 -3073 0 net=5283
rlabel metal2 30 -3084 30 -3084 0 net=2152
rlabel metal2 478 -3084 478 -3084 0 net=4692
rlabel metal2 646 -3084 646 -3084 0 net=8354
rlabel metal2 999 -3084 999 -3084 0 net=11758
rlabel metal2 37 -3086 37 -3086 0 net=4152
rlabel metal2 114 -3086 114 -3086 0 net=2585
rlabel metal2 215 -3086 215 -3086 0 net=1626
rlabel metal2 275 -3086 275 -3086 0 net=1650
rlabel metal2 814 -3086 814 -3086 0 net=3292
rlabel metal2 1090 -3086 1090 -3086 0 net=10680
rlabel metal2 1475 -3086 1475 -3086 0 net=12738
rlabel metal2 61 -3088 61 -3088 0 net=3478
rlabel metal2 656 -3088 656 -3088 0 net=6238
rlabel metal2 789 -3088 789 -3088 0 net=6230
rlabel metal2 877 -3088 877 -3088 0 net=9222
rlabel metal2 1388 -3088 1388 -3088 0 net=12807
rlabel metal2 65 -3090 65 -3090 0 net=5890
rlabel metal2 82 -3090 82 -3090 0 net=5442
rlabel metal2 471 -3090 471 -3090 0 net=5842
rlabel metal2 842 -3090 842 -3090 0 net=7521
rlabel metal2 1020 -3090 1020 -3090 0 net=11866
rlabel metal2 79 -3092 79 -3092 0 net=11457
rlabel metal2 716 -3092 716 -3092 0 net=5278
rlabel metal2 933 -3092 933 -3092 0 net=6752
rlabel metal2 1171 -3092 1171 -3092 0 net=11251
rlabel metal2 1444 -3092 1444 -3092 0 net=11813
rlabel metal2 86 -3094 86 -3094 0 net=2479
rlabel metal2 184 -3094 184 -3094 0 net=874
rlabel metal2 975 -3094 975 -3094 0 net=8049
rlabel metal2 1062 -3094 1062 -3094 0 net=12836
rlabel metal2 117 -3096 117 -3096 0 net=8390
rlabel metal2 1339 -3096 1339 -3096 0 net=12489
rlabel metal2 131 -3098 131 -3098 0 net=3837
rlabel metal2 219 -3098 219 -3098 0 net=3173
rlabel metal2 254 -3098 254 -3098 0 net=6821
rlabel metal2 933 -3098 933 -3098 0 net=9683
rlabel metal2 1276 -3098 1276 -3098 0 net=13383
rlabel metal2 135 -3100 135 -3100 0 net=3724
rlabel metal2 177 -3100 177 -3100 0 net=4375
rlabel metal2 282 -3100 282 -3100 0 net=3484
rlabel metal2 404 -3100 404 -3100 0 net=3817
rlabel metal2 453 -3100 453 -3100 0 net=11981
rlabel metal2 940 -3100 940 -3100 0 net=11285
rlabel metal2 1423 -3100 1423 -3100 0 net=13553
rlabel metal2 51 -3102 51 -3102 0 net=2135
rlabel metal2 303 -3102 303 -3102 0 net=3812
rlabel metal2 527 -3102 527 -3102 0 net=5457
rlabel metal2 674 -3102 674 -3102 0 net=5676
rlabel metal2 779 -3102 779 -3102 0 net=7318
rlabel metal2 1083 -3102 1083 -3102 0 net=11354
rlabel metal2 1423 -3102 1423 -3102 0 net=13229
rlabel metal2 93 -3104 93 -3104 0 net=4245
rlabel metal2 317 -3104 317 -3104 0 net=2657
rlabel metal2 317 -3104 317 -3104 0 net=2657
rlabel metal2 324 -3104 324 -3104 0 net=3127
rlabel metal2 324 -3104 324 -3104 0 net=3127
rlabel metal2 345 -3104 345 -3104 0 net=2843
rlabel metal2 366 -3104 366 -3104 0 net=4076
rlabel metal2 593 -3104 593 -3104 0 net=5726
rlabel metal2 674 -3104 674 -3104 0 net=5413
rlabel metal2 758 -3104 758 -3104 0 net=6679
rlabel metal2 940 -3104 940 -3104 0 net=8331
rlabel metal2 1367 -3104 1367 -3104 0 net=12699
rlabel metal2 1605 -3104 1605 -3104 0 net=13699
rlabel metal2 93 -3106 93 -3106 0 net=7001
rlabel metal2 744 -3106 744 -3106 0 net=6527
rlabel metal2 919 -3106 919 -3106 0 net=8261
rlabel metal2 1430 -3106 1430 -3106 0 net=13249
rlabel metal2 135 -3108 135 -3108 0 net=5225
rlabel metal2 684 -3108 684 -3108 0 net=5118
rlabel metal2 142 -3110 142 -3110 0 net=12186
rlabel metal2 142 -3112 142 -3112 0 net=5699
rlabel metal2 793 -3112 793 -3112 0 net=5634
rlabel metal2 800 -3112 800 -3112 0 net=6889
rlabel metal2 877 -3112 877 -3112 0 net=7931
rlabel metal2 1031 -3112 1031 -3112 0 net=8317
rlabel metal2 1360 -3112 1360 -3112 0 net=12651
rlabel metal2 145 -3114 145 -3114 0 net=1676
rlabel metal2 184 -3114 184 -3114 0 net=3855
rlabel metal2 534 -3114 534 -3114 0 net=1846
rlabel metal2 838 -3114 838 -3114 0 net=8324
rlabel metal2 1486 -3114 1486 -3114 0 net=13349
rlabel metal2 121 -3116 121 -3116 0 net=2400
rlabel metal2 562 -3116 562 -3116 0 net=3513
rlabel metal2 660 -3116 660 -3116 0 net=5711
rlabel metal2 793 -3116 793 -3116 0 net=11754
rlabel metal2 100 -3118 100 -3118 0 net=5893
rlabel metal2 149 -3118 149 -3118 0 net=11588
rlabel metal2 89 -3120 89 -3120 0 net=11037
rlabel metal2 152 -3120 152 -3120 0 net=3122
rlabel metal2 348 -3120 348 -3120 0 net=1800
rlabel metal2 394 -3120 394 -3120 0 net=3219
rlabel metal2 562 -3120 562 -3120 0 net=5931
rlabel metal2 828 -3120 828 -3120 0 net=7309
rlabel metal2 982 -3120 982 -3120 0 net=8985
rlabel metal2 44 -3122 44 -3122 0 net=2165
rlabel metal2 352 -3122 352 -3122 0 net=2999
rlabel metal2 618 -3122 618 -3122 0 net=5257
rlabel metal2 716 -3122 716 -3122 0 net=13469
rlabel metal2 947 -3122 947 -3122 0 net=9158
rlabel metal2 152 -3124 152 -3124 0 net=10
rlabel metal2 821 -3124 821 -3124 0 net=8508
rlabel metal2 1129 -3124 1129 -3124 0 net=11019
rlabel metal2 156 -3126 156 -3126 0 net=5583
rlabel metal2 576 -3126 576 -3126 0 net=4042
rlabel metal2 1066 -3126 1066 -3126 0 net=10063
rlabel metal2 1283 -3126 1283 -3126 0 net=11971
rlabel metal2 156 -3128 156 -3128 0 net=4757
rlabel metal2 688 -3128 688 -3128 0 net=7236
rlabel metal2 730 -3128 730 -3128 0 net=1865
rlabel metal2 835 -3128 835 -3128 0 net=6754
rlabel metal2 163 -3130 163 -3130 0 net=6737
rlabel metal2 772 -3130 772 -3130 0 net=8511
rlabel metal2 1164 -3130 1164 -3130 0 net=11685
rlabel metal2 170 -3132 170 -3132 0 net=4457
rlabel metal2 429 -3132 429 -3132 0 net=5803
rlabel metal2 653 -3132 653 -3132 0 net=5921
rlabel metal2 691 -3132 691 -3132 0 net=13036
rlabel metal2 191 -3134 191 -3134 0 net=1534
rlabel metal2 219 -3134 219 -3134 0 net=3589
rlabel metal2 457 -3134 457 -3134 0 net=4465
rlabel metal2 579 -3134 579 -3134 0 net=10851
rlabel metal2 1234 -3134 1234 -3134 0 net=11713
rlabel metal2 128 -3136 128 -3136 0 net=5339
rlabel metal2 478 -3136 478 -3136 0 net=5493
rlabel metal2 786 -3136 786 -3136 0 net=7377
rlabel metal2 947 -3136 947 -3136 0 net=8924
rlabel metal2 1409 -3136 1409 -3136 0 net=12398
rlabel metal2 72 -3138 72 -3138 0 net=4170
rlabel metal2 191 -3138 191 -3138 0 net=1507
rlabel metal2 261 -3138 261 -3138 0 net=1985
rlabel metal2 492 -3138 492 -3138 0 net=4531
rlabel metal2 681 -3138 681 -3138 0 net=9543
rlabel metal2 730 -3138 730 -3138 0 net=6457
rlabel metal2 898 -3138 898 -3138 0 net=8075
rlabel metal2 1003 -3138 1003 -3138 0 net=7699
rlabel metal2 1269 -3138 1269 -3138 0 net=12453
rlabel metal2 72 -3140 72 -3140 0 net=2179
rlabel metal2 233 -3140 233 -3140 0 net=1609
rlabel metal2 261 -3140 261 -3140 0 net=1777
rlabel metal2 366 -3140 366 -3140 0 net=3067
rlabel metal2 432 -3140 432 -3140 0 net=3208
rlabel metal2 492 -3140 492 -3140 0 net=3874
rlabel metal2 695 -3140 695 -3140 0 net=5135
rlabel metal2 849 -3140 849 -3140 0 net=6911
rlabel metal2 968 -3140 968 -3140 0 net=11061
rlabel metal2 1297 -3140 1297 -3140 0 net=11079
rlabel metal2 198 -3142 198 -3142 0 net=1016
rlabel metal2 1178 -3142 1178 -3142 0 net=9326
rlabel metal2 1325 -3142 1325 -3142 0 net=11167
rlabel metal2 149 -3144 149 -3144 0 net=10831
rlabel metal2 1178 -3144 1178 -3144 0 net=11649
rlabel metal2 1325 -3144 1325 -3144 0 net=12315
rlabel metal2 198 -3146 198 -3146 0 net=6409
rlabel metal2 954 -3146 954 -3146 0 net=9079
rlabel metal2 1227 -3146 1227 -3146 0 net=11761
rlabel metal2 369 -3148 369 -3148 0 net=4102
rlabel metal2 537 -3148 537 -3148 0 net=13115
rlabel metal2 226 -3150 226 -3150 0 net=4817
rlabel metal2 702 -3150 702 -3150 0 net=6041
rlabel metal2 870 -3150 870 -3150 0 net=6399
rlabel metal2 233 -3152 233 -3152 0 net=4281
rlabel metal2 737 -3152 737 -3152 0 net=6613
rlabel metal2 856 -3152 856 -3152 0 net=8359
rlabel metal2 989 -3152 989 -3152 0 net=11773
rlabel metal2 373 -3154 373 -3154 0 net=3303
rlabel metal2 548 -3154 548 -3154 0 net=4925
rlabel metal2 751 -3154 751 -3154 0 net=6629
rlabel metal2 1003 -3154 1003 -3154 0 net=9433
rlabel metal2 1311 -3154 1311 -3154 0 net=12247
rlabel metal2 107 -3156 107 -3156 0 net=3993
rlabel metal2 380 -3156 380 -3156 0 net=3929
rlabel metal2 597 -3156 597 -3156 0 net=5285
rlabel metal2 611 -3156 611 -3156 0 net=5403
rlabel metal2 765 -3156 765 -3156 0 net=6803
rlabel metal2 1024 -3156 1024 -3156 0 net=8569
rlabel metal2 1122 -3156 1122 -3156 0 net=8743
rlabel metal2 107 -3158 107 -3158 0 net=6785
rlabel metal2 667 -3158 667 -3158 0 net=6179
rlabel metal2 884 -3158 884 -3158 0 net=7871
rlabel metal2 1038 -3158 1038 -3158 0 net=10373
rlabel metal2 1402 -3158 1402 -3158 0 net=13111
rlabel metal2 387 -3160 387 -3160 0 net=2701
rlabel metal2 471 -3160 471 -3160 0 net=10111
rlabel metal2 905 -3160 905 -3160 0 net=8101
rlabel metal2 1052 -3160 1052 -3160 0 net=9823
rlabel metal2 1248 -3160 1248 -3160 0 net=12441
rlabel metal2 387 -3162 387 -3162 0 net=9051
rlabel metal2 1150 -3162 1150 -3162 0 net=9805
rlabel metal2 1220 -3162 1220 -3162 0 net=11555
rlabel metal2 1437 -3162 1437 -3162 0 net=13277
rlabel metal2 401 -3164 401 -3164 0 net=3618
rlabel metal2 590 -3164 590 -3164 0 net=4575
rlabel metal2 632 -3164 632 -3164 0 net=11511
rlabel metal2 1304 -3164 1304 -3164 0 net=9845
rlabel metal2 114 -3166 114 -3166 0 net=8267
rlabel metal2 632 -3166 632 -3166 0 net=7201
rlabel metal2 978 -3166 978 -3166 0 net=12127
rlabel metal2 1381 -3166 1381 -3166 0 net=12727
rlabel metal2 408 -3168 408 -3168 0 net=4211
rlabel metal2 639 -3168 639 -3168 0 net=9701
rlabel metal2 429 -3170 429 -3170 0 net=5209
rlabel metal2 709 -3170 709 -3170 0 net=5747
rlabel metal2 912 -3170 912 -3170 0 net=8221
rlabel metal2 1094 -3170 1094 -3170 0 net=10983
rlabel metal2 1122 -3170 1122 -3170 0 net=11143
rlabel metal2 576 -3172 576 -3172 0 net=7543
rlabel metal2 961 -3172 961 -3172 0 net=8551
rlabel metal2 1136 -3172 1136 -3172 0 net=11087
rlabel metal2 1185 -3172 1185 -3172 0 net=9609
rlabel metal2 1045 -3174 1045 -3174 0 net=9637
rlabel metal2 1206 -3174 1206 -3174 0 net=11471
rlabel metal2 1094 -3176 1094 -3176 0 net=10849
rlabel metal2 1318 -3176 1318 -3176 0 net=12283
rlabel metal2 996 -3178 996 -3178 0 net=7623
rlabel metal2 996 -3180 996 -3180 0 net=12879
rlabel metal2 1017 -3182 1017 -3182 0 net=11913
rlabel metal2 1374 -3182 1374 -3182 0 net=12721
rlabel metal2 1017 -3184 1017 -3184 0 net=11025
rlabel metal2 1108 -3186 1108 -3186 0 net=7783
rlabel metal2 1136 -3188 1136 -3188 0 net=10481
rlabel metal2 1290 -3188 1290 -3188 0 net=12101
rlabel metal2 1143 -3190 1143 -3190 0 net=10149
rlabel metal2 1255 -3190 1255 -3190 0 net=11891
rlabel metal2 450 -3192 450 -3192 0 net=13579
rlabel metal2 310 -3194 310 -3194 0 net=5323
rlabel metal2 1185 -3194 1185 -3194 0 net=11201
rlabel metal2 310 -3196 310 -3196 0 net=2679
rlabel metal2 621 -3196 621 -3196 0 net=12473
rlabel metal2 331 -3198 331 -3198 0 net=3149
rlabel metal2 1192 -3198 1192 -3198 0 net=11265
rlabel metal2 422 -3200 422 -3200 0 net=5625
rlabel metal2 1241 -3200 1241 -3200 0 net=13009
rlabel metal2 296 -3202 296 -3202 0 net=3041
rlabel metal2 1346 -3202 1346 -3202 0 net=6761
rlabel metal2 296 -3204 296 -3204 0 net=2773
rlabel metal2 338 -3206 338 -3206 0 net=3227
rlabel metal2 359 -3208 359 -3208 0 net=4009
rlabel metal2 499 -3210 499 -3210 0 net=5011
rlabel metal2 275 -3212 275 -3212 0 net=3231
rlabel metal2 65 -3223 65 -3223 0 net=462
rlabel metal2 121 -3223 121 -3223 0 net=5894
rlabel metal2 502 -3223 502 -3223 0 net=13470
rlabel metal2 779 -3223 779 -3223 0 net=6400
rlabel metal2 880 -3223 880 -3223 0 net=8318
rlabel metal2 1059 -3223 1059 -3223 0 net=12475
rlabel metal2 1346 -3223 1346 -3223 0 net=9610
rlabel metal2 1584 -3223 1584 -3223 0 net=13701
rlabel metal2 72 -3225 72 -3225 0 net=2180
rlabel metal2 485 -3225 485 -3225 0 net=3042
rlabel metal2 593 -3225 593 -3225 0 net=5414
rlabel metal2 684 -3225 684 -3225 0 net=7378
rlabel metal2 800 -3225 800 -3225 0 net=6890
rlabel metal2 1409 -3225 1409 -3225 0 net=11168
rlabel metal2 86 -3227 86 -3227 0 net=2480
rlabel metal2 404 -3227 404 -3227 0 net=4532
rlabel metal2 544 -3227 544 -3227 0 net=5012
rlabel metal2 576 -3227 576 -3227 0 net=5404
rlabel metal2 625 -3227 625 -3227 0 net=5458
rlabel metal2 800 -3227 800 -3227 0 net=6913
rlabel metal2 894 -3227 894 -3227 0 net=11088
rlabel metal2 1185 -3227 1185 -3227 0 net=11202
rlabel metal2 1297 -3227 1297 -3227 0 net=7625
rlabel metal2 142 -3229 142 -3229 0 net=5701
rlabel metal2 597 -3229 597 -3229 0 net=4577
rlabel metal2 597 -3229 597 -3229 0 net=4577
rlabel metal2 611 -3229 611 -3229 0 net=6615
rlabel metal2 849 -3229 849 -3229 0 net=9081
rlabel metal2 999 -3229 999 -3229 0 net=9434
rlabel metal2 1010 -3229 1010 -3229 0 net=12454
rlabel metal2 1300 -3229 1300 -3229 0 net=6762
rlabel metal2 149 -3231 149 -3231 0 net=1508
rlabel metal2 212 -3231 212 -3231 0 net=2587
rlabel metal2 243 -3231 243 -3231 0 net=2658
rlabel metal2 324 -3231 324 -3231 0 net=3128
rlabel metal2 1020 -3231 1020 -3231 0 net=10482
rlabel metal2 1269 -3231 1269 -3231 0 net=12729
rlabel metal2 1458 -3231 1458 -3231 0 net=11814
rlabel metal2 107 -3233 107 -3233 0 net=6787
rlabel metal2 226 -3233 226 -3233 0 net=4819
rlabel metal2 492 -3233 492 -3233 0 net=8512
rlabel metal2 905 -3233 905 -3233 0 net=8102
rlabel metal2 1010 -3233 1010 -3233 0 net=11473
rlabel metal2 1325 -3233 1325 -3233 0 net=12317
rlabel metal2 1332 -3233 1332 -3233 0 net=12809
rlabel metal2 152 -3235 152 -3235 0 net=4010
rlabel metal2 387 -3235 387 -3235 0 net=9053
rlabel metal2 415 -3235 415 -3235 0 net=3304
rlabel metal2 544 -3235 544 -3235 0 net=641
rlabel metal2 905 -3235 905 -3235 0 net=12442
rlabel metal2 1325 -3235 1325 -3235 0 net=12653
rlabel metal2 1381 -3235 1381 -3235 0 net=9847
rlabel metal2 156 -3237 156 -3237 0 net=4758
rlabel metal2 541 -3237 541 -3237 0 net=1009
rlabel metal2 954 -3237 954 -3237 0 net=11287
rlabel metal2 1346 -3237 1346 -3237 0 net=13231
rlabel metal2 170 -3239 170 -3239 0 net=4458
rlabel metal2 499 -3239 499 -3239 0 net=4927
rlabel metal2 555 -3239 555 -3239 0 net=5287
rlabel metal2 625 -3239 625 -3239 0 net=7545
rlabel metal2 940 -3239 940 -3239 0 net=8332
rlabel metal2 1031 -3239 1031 -3239 0 net=11557
rlabel metal2 1349 -3239 1349 -3239 0 net=11080
rlabel metal2 93 -3241 93 -3241 0 net=7003
rlabel metal2 177 -3241 177 -3241 0 net=4376
rlabel metal2 359 -3241 359 -3241 0 net=3221
rlabel metal2 429 -3241 429 -3241 0 net=5324
rlabel metal2 457 -3241 457 -3241 0 net=5341
rlabel metal2 604 -3241 604 -3241 0 net=6181
rlabel metal2 705 -3241 705 -3241 0 net=11026
rlabel metal2 1087 -3241 1087 -3241 0 net=12285
rlabel metal2 1353 -3241 1353 -3241 0 net=13350
rlabel metal2 191 -3243 191 -3243 0 net=3839
rlabel metal2 226 -3243 226 -3243 0 net=4487
rlabel metal2 940 -3243 940 -3243 0 net=8987
rlabel metal2 996 -3243 996 -3243 0 net=11253
rlabel metal2 1199 -3243 1199 -3243 0 net=13011
rlabel metal2 1283 -3243 1283 -3243 0 net=11973
rlabel metal2 1388 -3243 1388 -3243 0 net=12881
rlabel metal2 205 -3245 205 -3245 0 net=7203
rlabel metal2 653 -3245 653 -3245 0 net=6043
rlabel metal2 709 -3245 709 -3245 0 net=5748
rlabel metal2 919 -3245 919 -3245 0 net=8263
rlabel metal2 233 -3247 233 -3247 0 net=4283
rlabel metal2 233 -3247 233 -3247 0 net=4283
rlabel metal2 247 -3247 247 -3247 0 net=1610
rlabel metal2 520 -3247 520 -3247 0 net=8269
rlabel metal2 919 -3247 919 -3247 0 net=10833
rlabel metal2 1090 -3247 1090 -3247 0 net=11650
rlabel metal2 1220 -3247 1220 -3247 0 net=13279
rlabel metal2 135 -3249 135 -3249 0 net=5227
rlabel metal2 254 -3249 254 -3249 0 net=6822
rlabel metal2 709 -3249 709 -3249 0 net=8615
rlabel metal2 947 -3249 947 -3249 0 net=10985
rlabel metal2 1129 -3249 1129 -3249 0 net=11020
rlabel metal2 1234 -3249 1234 -3249 0 net=11715
rlabel metal2 128 -3251 128 -3251 0 net=10115
rlabel metal2 254 -3251 254 -3251 0 net=3453
rlabel metal2 716 -3251 716 -3251 0 net=7311
rlabel metal2 891 -3251 891 -3251 0 net=561
rlabel metal2 1234 -3251 1234 -3251 0 net=12129
rlabel metal2 261 -3253 261 -3253 0 net=1779
rlabel metal2 429 -3253 429 -3253 0 net=4131
rlabel metal2 828 -3253 828 -3253 0 net=8745
rlabel metal2 261 -3255 261 -3255 0 net=3151
rlabel metal2 338 -3255 338 -3255 0 net=3228
rlabel metal2 450 -3255 450 -3255 0 net=5495
rlabel metal2 520 -3255 520 -3255 0 net=5211
rlabel metal2 632 -3255 632 -3255 0 net=6459
rlabel metal2 737 -3255 737 -3255 0 net=7701
rlabel metal2 1080 -3255 1080 -3255 0 net=11915
rlabel metal2 1304 -3255 1304 -3255 0 net=1707
rlabel metal2 198 -3257 198 -3257 0 net=6411
rlabel metal2 751 -3257 751 -3257 0 net=6631
rlabel metal2 1171 -3257 1171 -3257 0 net=13385
rlabel metal2 79 -3259 79 -3259 0 net=11459
rlabel metal2 268 -3259 268 -3259 0 net=2167
rlabel metal2 268 -3259 268 -3259 0 net=2167
rlabel metal2 275 -3259 275 -3259 0 net=3233
rlabel metal2 352 -3259 352 -3259 0 net=3001
rlabel metal2 548 -3259 548 -3259 0 net=5713
rlabel metal2 667 -3259 667 -3259 0 net=6529
rlabel metal2 751 -3259 751 -3259 0 net=11763
rlabel metal2 1276 -3259 1276 -3259 0 net=12723
rlabel metal2 184 -3261 184 -3261 0 net=3857
rlabel metal2 282 -3261 282 -3261 0 net=2137
rlabel metal2 352 -3261 352 -3261 0 net=4213
rlabel metal2 422 -3261 422 -3261 0 net=5627
rlabel metal2 660 -3261 660 -3261 0 net=10281
rlabel metal2 723 -3261 723 -3261 0 net=9545
rlabel metal2 891 -3261 891 -3261 0 net=10529
rlabel metal2 163 -3263 163 -3263 0 net=6739
rlabel metal2 422 -3263 422 -3263 0 net=5259
rlabel metal2 681 -3263 681 -3263 0 net=5137
rlabel metal2 723 -3263 723 -3263 0 net=7523
rlabel metal2 968 -3263 968 -3263 0 net=11063
rlabel metal2 1052 -3263 1052 -3263 0 net=9825
rlabel metal2 100 -3265 100 -3265 0 net=11039
rlabel metal2 184 -3265 184 -3265 0 net=9487
rlabel metal2 618 -3265 618 -3265 0 net=11774
rlabel metal2 1045 -3265 1045 -3265 0 net=9639
rlabel metal2 1073 -3265 1073 -3265 0 net=10151
rlabel metal2 1213 -3265 1213 -3265 0 net=11513
rlabel metal2 282 -3267 282 -3267 0 net=6507
rlabel metal2 968 -3267 968 -3267 0 net=10375
rlabel metal2 1045 -3267 1045 -3267 0 net=11893
rlabel metal2 296 -3269 296 -3269 0 net=2775
rlabel metal2 373 -3269 373 -3269 0 net=3995
rlabel metal2 457 -3269 457 -3269 0 net=3027
rlabel metal2 814 -3269 814 -3269 0 net=1867
rlabel metal2 1094 -3269 1094 -3269 0 net=10850
rlabel metal2 296 -3271 296 -3271 0 net=3931
rlabel metal2 387 -3271 387 -3271 0 net=1987
rlabel metal2 471 -3271 471 -3271 0 net=5083
rlabel metal2 534 -3271 534 -3271 0 net=2965
rlabel metal2 1094 -3271 1094 -3271 0 net=12103
rlabel metal2 303 -3273 303 -3273 0 net=4247
rlabel metal2 380 -3273 380 -3273 0 net=4467
rlabel metal2 695 -3273 695 -3273 0 net=7933
rlabel metal2 1101 -3273 1101 -3273 0 net=10853
rlabel metal2 1290 -3273 1290 -3273 0 net=13555
rlabel metal2 303 -3275 303 -3275 0 net=2681
rlabel metal2 317 -3275 317 -3275 0 net=2845
rlabel metal2 443 -3275 443 -3275 0 net=3514
rlabel metal2 744 -3275 744 -3275 0 net=9413
rlabel metal2 842 -3275 842 -3275 0 net=12491
rlabel metal2 177 -3277 177 -3277 0 net=9641
rlabel metal2 513 -3277 513 -3277 0 net=5805
rlabel metal2 758 -3277 758 -3277 0 net=6680
rlabel metal2 1101 -3277 1101 -3277 0 net=13117
rlabel metal2 289 -3279 289 -3279 0 net=3175
rlabel metal2 464 -3279 464 -3279 0 net=2703
rlabel metal2 758 -3279 758 -3279 0 net=7873
rlabel metal2 1115 -3279 1115 -3279 0 net=13251
rlabel metal2 289 -3281 289 -3281 0 net=3819
rlabel metal2 464 -3281 464 -3281 0 net=5923
rlabel metal2 772 -3281 772 -3281 0 net=11745
rlabel metal2 1311 -3281 1311 -3281 0 net=12249
rlabel metal2 366 -3283 366 -3283 0 net=3068
rlabel metal2 793 -3283 793 -3283 0 net=8553
rlabel metal2 1129 -3283 1129 -3283 0 net=11686
rlabel metal2 1311 -3283 1311 -3283 0 net=12701
rlabel metal2 219 -3285 219 -3285 0 net=3591
rlabel metal2 814 -3285 814 -3285 0 net=8571
rlabel metal2 1143 -3285 1143 -3285 0 net=9807
rlabel metal2 1164 -3285 1164 -3285 0 net=11267
rlabel metal2 1328 -3285 1328 -3285 0 net=1
rlabel metal2 219 -3287 219 -3287 0 net=5933
rlabel metal2 821 -3287 821 -3287 0 net=9685
rlabel metal2 1150 -3287 1150 -3287 0 net=5179
rlabel metal2 506 -3289 506 -3289 0 net=5585
rlabel metal2 856 -3289 856 -3289 0 net=8361
rlabel metal2 915 -3289 915 -3289 0 net=7111
rlabel metal2 1192 -3289 1192 -3289 0 net=13113
rlabel metal2 506 -3291 506 -3291 0 net=6805
rlabel metal2 856 -3291 856 -3291 0 net=8077
rlabel metal2 926 -3291 926 -3291 0 net=11983
rlabel metal2 765 -3293 765 -3293 0 net=8223
rlabel metal2 926 -3293 926 -3293 0 net=10065
rlabel metal2 863 -3295 863 -3295 0 net=10113
rlabel metal2 1066 -3295 1066 -3295 0 net=4081
rlabel metal2 639 -3297 639 -3297 0 net=9703
rlabel metal2 912 -3297 912 -3297 0 net=8050
rlabel metal2 639 -3299 639 -3299 0 net=12511
rlabel metal2 933 -3299 933 -3299 0 net=7785
rlabel metal2 835 -3301 835 -3301 0 net=4153
rlabel metal2 975 -3303 975 -3303 0 net=11145
rlabel metal2 1122 -3305 1122 -3305 0 net=13581
rlabel metal2 131 -3316 131 -3316 0 net=10116
rlabel metal2 163 -3316 163 -3316 0 net=11040
rlabel metal2 590 -3316 590 -3316 0 net=5342
rlabel metal2 691 -3316 691 -3316 0 net=10854
rlabel metal2 1178 -3316 1178 -3316 0 net=1096
rlabel metal2 1577 -3316 1577 -3316 0 net=13703
rlabel metal2 205 -3318 205 -3318 0 net=7205
rlabel metal2 590 -3318 590 -3318 0 net=12493
rlabel metal2 870 -3318 870 -3318 0 net=13114
rlabel metal2 1209 -3318 1209 -3318 0 net=12724
rlabel metal2 1360 -3318 1360 -3318 0 net=12319
rlabel metal2 1388 -3318 1388 -3318 0 net=12883
rlabel metal2 1388 -3318 1388 -3318 0 net=12883
rlabel metal2 233 -3320 233 -3320 0 net=4285
rlabel metal2 506 -3320 506 -3320 0 net=6806
rlabel metal2 870 -3320 870 -3320 0 net=13131
rlabel metal2 1003 -3320 1003 -3320 0 net=11064
rlabel metal2 1111 -3320 1111 -3320 0 net=13556
rlabel metal2 212 -3322 212 -3322 0 net=6789
rlabel metal2 513 -3322 513 -3322 0 net=5806
rlabel metal2 614 -3322 614 -3322 0 net=5180
rlabel metal2 1153 -3322 1153 -3322 0 net=12130
rlabel metal2 1248 -3322 1248 -3322 0 net=12654
rlabel metal2 247 -3324 247 -3324 0 net=5228
rlabel metal2 464 -3324 464 -3324 0 net=5924
rlabel metal2 705 -3324 705 -3324 0 net=1478
rlabel metal2 880 -3324 880 -3324 0 net=6632
rlabel metal2 1192 -3324 1192 -3324 0 net=8265
rlabel metal2 198 -3326 198 -3326 0 net=11461
rlabel metal2 268 -3326 268 -3326 0 net=2168
rlabel metal2 621 -3326 621 -3326 0 net=7
rlabel metal2 915 -3326 915 -3326 0 net=9808
rlabel metal2 1199 -3326 1199 -3326 0 net=13013
rlabel metal2 1262 -3326 1262 -3326 0 net=12702
rlabel metal2 240 -3328 240 -3328 0 net=2589
rlabel metal2 310 -3328 310 -3328 0 net=3176
rlabel metal2 429 -3328 429 -3328 0 net=4133
rlabel metal2 429 -3328 429 -3328 0 net=4133
rlabel metal2 436 -3328 436 -3328 0 net=5085
rlabel metal2 485 -3328 485 -3328 0 net=4820
rlabel metal2 961 -3328 961 -3328 0 net=7112
rlabel metal2 1171 -3328 1171 -3328 0 net=13387
rlabel metal2 1213 -3328 1213 -3328 0 net=11716
rlabel metal2 1311 -3328 1311 -3328 0 net=12811
rlabel metal2 177 -3330 177 -3330 0 net=9643
rlabel metal2 359 -3330 359 -3330 0 net=3223
rlabel metal2 523 -3330 523 -3330 0 net=13591
rlabel metal2 716 -3330 716 -3330 0 net=7312
rlabel metal2 894 -3330 894 -3330 0 net=832
rlabel metal2 1234 -3330 1234 -3330 0 net=9827
rlabel metal2 1332 -3330 1332 -3330 0 net=9849
rlabel metal2 359 -3332 359 -3332 0 net=3593
rlabel metal2 380 -3332 380 -3332 0 net=4469
rlabel metal2 471 -3332 471 -3332 0 net=4929
rlabel metal2 618 -3332 618 -3332 0 net=8617
rlabel metal2 716 -3332 716 -3332 0 net=8271
rlabel metal2 789 -3332 789 -3332 0 net=6914
rlabel metal2 901 -3332 901 -3332 0 net=8988
rlabel metal2 947 -3332 947 -3332 0 net=10987
rlabel metal2 1171 -3332 1171 -3332 0 net=7627
rlabel metal2 1353 -3332 1353 -3332 0 net=11975
rlabel metal2 170 -3334 170 -3334 0 net=7004
rlabel metal2 632 -3334 632 -3334 0 net=6460
rlabel metal2 947 -3334 947 -3334 0 net=10376
rlabel metal2 982 -3334 982 -3334 0 net=11268
rlabel metal2 1213 -3334 1213 -3334 0 net=11443
rlabel metal2 275 -3336 275 -3336 0 net=3859
rlabel metal2 380 -3336 380 -3336 0 net=3045
rlabel metal2 478 -3336 478 -3336 0 net=3003
rlabel metal2 632 -3336 632 -3336 0 net=7525
rlabel metal2 730 -3336 730 -3336 0 net=6412
rlabel metal2 898 -3336 898 -3336 0 net=10067
rlabel metal2 961 -3336 961 -3336 0 net=13119
rlabel metal2 1164 -3336 1164 -3336 0 net=12730
rlabel metal2 394 -3338 394 -3338 0 net=1781
rlabel metal2 478 -3338 478 -3338 0 net=5213
rlabel metal2 639 -3338 639 -3338 0 net=12513
rlabel metal2 891 -3338 891 -3338 0 net=10531
rlabel metal2 982 -3338 982 -3338 0 net=13583
rlabel metal2 1241 -3338 1241 -3338 0 net=12251
rlabel metal2 345 -3340 345 -3340 0 net=2985
rlabel metal2 401 -3340 401 -3340 0 net=3997
rlabel metal2 576 -3340 576 -3340 0 net=5703
rlabel metal2 667 -3340 667 -3340 0 net=6531
rlabel metal2 996 -3340 996 -3340 0 net=11255
rlabel metal2 282 -3342 282 -3342 0 net=6509
rlabel metal2 548 -3342 548 -3342 0 net=5714
rlabel metal2 667 -3342 667 -3342 0 net=9415
rlabel metal2 758 -3342 758 -3342 0 net=7875
rlabel metal2 1003 -3342 1003 -3342 0 net=12287
rlabel metal2 1094 -3342 1094 -3342 0 net=12105
rlabel metal2 184 -3344 184 -3344 0 net=9489
rlabel metal2 317 -3344 317 -3344 0 net=2847
rlabel metal2 530 -3344 530 -3344 0 net=3643
rlabel metal2 226 -3346 226 -3346 0 net=4489
rlabel metal2 583 -3346 583 -3346 0 net=2705
rlabel metal2 863 -3346 863 -3346 0 net=9705
rlabel metal2 1013 -3346 1013 -3346 0 net=13280
rlabel metal2 219 -3348 219 -3348 0 net=5935
rlabel metal2 674 -3348 674 -3348 0 net=8747
rlabel metal2 1024 -3348 1024 -3348 0 net=11984
rlabel metal2 317 -3350 317 -3350 0 net=3235
rlabel metal2 408 -3350 408 -3350 0 net=6741
rlabel metal2 1024 -3350 1024 -3350 0 net=11514
rlabel metal2 296 -3352 296 -3352 0 net=3933
rlabel metal2 373 -3352 373 -3352 0 net=4249
rlabel metal2 709 -3352 709 -3352 0 net=11747
rlabel metal2 828 -3352 828 -3352 0 net=8363
rlabel metal2 1031 -3352 1031 -3352 0 net=11559
rlabel metal2 1038 -3352 1038 -3352 0 net=1868
rlabel metal2 191 -3354 191 -3354 0 net=3840
rlabel metal2 660 -3354 660 -3354 0 net=10283
rlabel metal2 814 -3354 814 -3354 0 net=8573
rlabel metal2 989 -3354 989 -3354 0 net=10114
rlabel metal2 1045 -3354 1045 -3354 0 net=11895
rlabel metal2 1185 -3354 1185 -3354 0 net=3345
rlabel metal2 261 -3356 261 -3356 0 net=3152
rlabel metal2 660 -3356 660 -3356 0 net=8225
rlabel metal2 849 -3356 849 -3356 0 net=9083
rlabel metal2 1031 -3356 1031 -3356 0 net=13253
rlabel metal2 1206 -3356 1206 -3356 0 net=12615
rlabel metal2 681 -3358 681 -3358 0 net=5139
rlabel metal2 681 -3360 681 -3360 0 net=10433
rlabel metal2 1066 -3360 1066 -3360 0 net=4083
rlabel metal2 702 -3362 702 -3362 0 net=7823
rlabel metal2 786 -3362 786 -3362 0 net=5641
rlabel metal2 1045 -3362 1045 -3362 0 net=10153
rlabel metal2 1080 -3362 1080 -3362 0 net=11917
rlabel metal2 646 -3364 646 -3364 0 net=9055
rlabel metal2 723 -3364 723 -3364 0 net=8555
rlabel metal2 856 -3364 856 -3364 0 net=8079
rlabel metal2 611 -3366 611 -3366 0 net=6617
rlabel metal2 856 -3366 856 -3366 0 net=12089
rlabel metal2 254 -3368 254 -3368 0 net=3454
rlabel metal2 646 -3368 646 -3368 0 net=11765
rlabel metal2 786 -3368 786 -3368 0 net=5119
rlabel metal2 933 -3368 933 -3368 0 net=7787
rlabel metal2 737 -3370 737 -3370 0 net=7703
rlabel metal2 1052 -3370 1052 -3370 0 net=9640
rlabel metal2 737 -3372 737 -3372 0 net=9547
rlabel metal2 933 -3372 933 -3372 0 net=12083
rlabel metal2 1066 -3372 1066 -3372 0 net=2549
rlabel metal2 387 -3374 387 -3374 0 net=1988
rlabel metal2 1265 -3374 1265 -3374 0 net=13232
rlabel metal2 387 -3376 387 -3376 0 net=3029
rlabel metal2 597 -3376 597 -3376 0 net=4579
rlabel metal2 450 -3378 450 -3378 0 net=5497
rlabel metal2 597 -3378 597 -3378 0 net=7935
rlabel metal2 744 -3378 744 -3378 0 net=9687
rlabel metal2 450 -3380 450 -3380 0 net=6231
rlabel metal2 695 -3380 695 -3380 0 net=4155
rlabel metal2 527 -3382 527 -3382 0 net=2967
rlabel metal2 562 -3382 562 -3382 0 net=5587
rlabel metal2 534 -3384 534 -3384 0 net=5289
rlabel metal2 562 -3384 562 -3384 0 net=5629
rlabel metal2 751 -3384 751 -3384 0 net=8993
rlabel metal2 555 -3386 555 -3386 0 net=7547
rlabel metal2 821 -3386 821 -3386 0 net=10835
rlabel metal2 569 -3388 569 -3388 0 net=6183
rlabel metal2 625 -3388 625 -3388 0 net=6045
rlabel metal2 912 -3388 912 -3388 0 net=11289
rlabel metal2 422 -3390 422 -3390 0 net=5261
rlabel metal2 919 -3390 919 -3390 0 net=11147
rlabel metal2 338 -3392 338 -3392 0 net=2139
rlabel metal2 604 -3392 604 -3392 0 net=6681
rlabel metal2 954 -3392 954 -3392 0 net=12627
rlabel metal2 338 -3394 338 -3394 0 net=4215
rlabel metal2 905 -3394 905 -3394 0 net=11475
rlabel metal2 324 -3396 324 -3396 0 net=2777
rlabel metal2 975 -3396 975 -3396 0 net=12477
rlabel metal2 303 -3398 303 -3398 0 net=2683
rlabel metal2 1059 -3398 1059 -3398 0 net=1708
rlabel metal2 289 -3400 289 -3400 0 net=3821
rlabel metal2 289 -3402 289 -3402 0 net=3687
rlabel metal2 240 -3413 240 -3413 0 net=9645
rlabel metal2 268 -3413 268 -3413 0 net=2590
rlabel metal2 338 -3413 338 -3413 0 net=4216
rlabel metal2 376 -3413 376 -3413 0 net=6232
rlabel metal2 457 -3413 457 -3413 0 net=5498
rlabel metal2 485 -3413 485 -3413 0 net=3005
rlabel metal2 632 -3413 632 -3413 0 net=7527
rlabel metal2 632 -3413 632 -3413 0 net=7527
rlabel metal2 639 -3413 639 -3413 0 net=5705
rlabel metal2 639 -3413 639 -3413 0 net=5705
rlabel metal2 663 -3413 663 -3413 0 net=716
rlabel metal2 1041 -3413 1041 -3413 0 net=10154
rlabel metal2 1052 -3413 1052 -3413 0 net=7789
rlabel metal2 1111 -3413 1111 -3413 0 net=8266
rlabel metal2 1199 -3413 1199 -3413 0 net=13388
rlabel metal2 1248 -3413 1248 -3413 0 net=13015
rlabel metal2 1304 -3413 1304 -3413 0 net=12813
rlabel metal2 1318 -3413 1318 -3413 0 net=11445
rlabel metal2 1374 -3413 1374 -3413 0 net=12321
rlabel metal2 1577 -3413 1577 -3413 0 net=13705
rlabel metal2 1577 -3413 1577 -3413 0 net=13705
rlabel metal2 247 -3415 247 -3415 0 net=11462
rlabel metal2 317 -3415 317 -3415 0 net=3237
rlabel metal2 499 -3415 499 -3415 0 net=6682
rlabel metal2 688 -3415 688 -3415 0 net=13593
rlabel metal2 688 -3415 688 -3415 0 net=13593
rlabel metal2 702 -3415 702 -3415 0 net=9056
rlabel metal2 824 -3415 824 -3415 0 net=13584
rlabel metal2 989 -3415 989 -3415 0 net=9084
rlabel metal2 1073 -3415 1073 -3415 0 net=11257
rlabel metal2 1122 -3415 1122 -3415 0 net=12107
rlabel metal2 1129 -3415 1129 -3415 0 net=11918
rlabel metal2 1185 -3415 1185 -3415 0 net=3347
rlabel metal2 1318 -3415 1318 -3415 0 net=9851
rlabel metal2 1381 -3415 1381 -3415 0 net=11977
rlabel metal2 282 -3417 282 -3417 0 net=9491
rlabel metal2 324 -3417 324 -3417 0 net=2685
rlabel metal2 352 -3417 352 -3417 0 net=2779
rlabel metal2 394 -3417 394 -3417 0 net=2987
rlabel metal2 513 -3417 513 -3417 0 net=3224
rlabel metal2 702 -3417 702 -3417 0 net=9549
rlabel metal2 793 -3417 793 -3417 0 net=6618
rlabel metal2 863 -3417 863 -3417 0 net=6742
rlabel metal2 1381 -3417 1381 -3417 0 net=12885
rlabel metal2 366 -3419 366 -3419 0 net=3861
rlabel metal2 415 -3419 415 -3419 0 net=2849
rlabel metal2 520 -3419 520 -3419 0 net=2968
rlabel metal2 562 -3419 562 -3419 0 net=5630
rlabel metal2 733 -3419 733 -3419 0 net=5120
rlabel metal2 800 -3419 800 -3419 0 net=5141
rlabel metal2 842 -3419 842 -3419 0 net=6533
rlabel metal2 884 -3419 884 -3419 0 net=8574
rlabel metal2 898 -3419 898 -3419 0 net=10068
rlabel metal2 1017 -3419 1017 -3419 0 net=13254
rlabel metal2 1080 -3419 1080 -3419 0 net=8081
rlabel metal2 359 -3421 359 -3421 0 net=3595
rlabel metal2 562 -3421 562 -3421 0 net=12495
rlabel metal2 625 -3421 625 -3421 0 net=6047
rlabel metal2 751 -3421 751 -3421 0 net=8995
rlabel metal2 898 -3421 898 -3421 0 net=11477
rlabel metal2 919 -3421 919 -3421 0 net=11149
rlabel metal2 996 -3421 996 -3421 0 net=9706
rlabel metal2 1024 -3421 1024 -3421 0 net=7628
rlabel metal2 359 -3423 359 -3423 0 net=6553
rlabel metal2 569 -3423 569 -3423 0 net=6185
rlabel metal2 569 -3423 569 -3423 0 net=6185
rlabel metal2 576 -3423 576 -3423 0 net=7937
rlabel metal2 625 -3423 625 -3423 0 net=11767
rlabel metal2 681 -3423 681 -3423 0 net=10435
rlabel metal2 758 -3423 758 -3423 0 net=2707
rlabel metal2 807 -3423 807 -3423 0 net=4581
rlabel metal2 849 -3423 849 -3423 0 net=5643
rlabel metal2 919 -3423 919 -3423 0 net=13121
rlabel metal2 968 -3423 968 -3423 0 net=7876
rlabel metal2 366 -3425 366 -3425 0 net=3031
rlabel metal2 415 -3425 415 -3425 0 net=5087
rlabel metal2 443 -3425 443 -3425 0 net=4470
rlabel metal2 597 -3425 597 -3425 0 net=4157
rlabel metal2 751 -3425 751 -3425 0 net=11821
rlabel metal2 877 -3425 877 -3425 0 net=5649
rlabel metal2 1031 -3425 1031 -3425 0 net=12201
rlabel metal2 1153 -3425 1153 -3425 0 net=12616
rlabel metal2 303 -3427 303 -3427 0 net=3823
rlabel metal2 450 -3427 450 -3427 0 net=5215
rlabel metal2 492 -3427 492 -3427 0 net=4286
rlabel metal2 618 -3427 618 -3427 0 net=8619
rlabel metal2 758 -3427 758 -3427 0 net=10837
rlabel metal2 877 -3427 877 -3427 0 net=7051
rlabel metal2 940 -3427 940 -3427 0 net=7705
rlabel metal2 1087 -3427 1087 -3427 0 net=3645
rlabel metal2 380 -3429 380 -3429 0 net=3047
rlabel metal2 408 -3429 408 -3429 0 net=4251
rlabel metal2 464 -3429 464 -3429 0 net=1783
rlabel metal2 548 -3429 548 -3429 0 net=4490
rlabel metal2 814 -3429 814 -3429 0 net=8365
rlabel metal2 912 -3429 912 -3429 0 net=11291
rlabel metal2 954 -3429 954 -3429 0 net=12629
rlabel metal2 1003 -3429 1003 -3429 0 net=12289
rlabel metal2 1101 -3429 1101 -3429 0 net=11561
rlabel metal2 1122 -3429 1122 -3429 0 net=10989
rlabel metal2 1157 -3429 1157 -3429 0 net=9828
rlabel metal2 331 -3431 331 -3431 0 net=3935
rlabel metal2 401 -3431 401 -3431 0 net=3999
rlabel metal2 471 -3431 471 -3431 0 net=4931
rlabel metal2 492 -3431 492 -3431 0 net=5291
rlabel metal2 548 -3431 548 -3431 0 net=7549
rlabel metal2 579 -3431 579 -3431 0 net=10391
rlabel metal2 1094 -3431 1094 -3431 0 net=4085
rlabel metal2 1129 -3431 1129 -3431 0 net=10499
rlabel metal2 299 -3433 299 -3433 0 net=2731
rlabel metal2 422 -3433 422 -3433 0 net=2140
rlabel metal2 534 -3433 534 -3433 0 net=7207
rlabel metal2 646 -3433 646 -3433 0 net=8227
rlabel metal2 681 -3433 681 -3433 0 net=11749
rlabel metal2 772 -3433 772 -3433 0 net=10285
rlabel metal2 912 -3433 912 -3433 0 net=10533
rlabel metal2 933 -3433 933 -3433 0 net=12085
rlabel metal2 961 -3433 961 -3433 0 net=12479
rlabel metal2 1003 -3433 1003 -3433 0 net=2551
rlabel metal2 1136 -3433 1136 -3433 0 net=11897
rlabel metal2 1206 -3433 1206 -3433 0 net=12253
rlabel metal2 345 -3435 345 -3435 0 net=6511
rlabel metal2 429 -3435 429 -3435 0 net=4135
rlabel metal2 429 -3435 429 -3435 0 net=4135
rlabel metal2 471 -3435 471 -3435 0 net=8531
rlabel metal2 709 -3435 709 -3435 0 net=9689
rlabel metal2 765 -3435 765 -3435 0 net=7825
rlabel metal2 1384 -3435 1384 -3435 0 net=1
rlabel metal2 310 -3437 310 -3437 0 net=3689
rlabel metal2 485 -3437 485 -3437 0 net=3753
rlabel metal2 716 -3437 716 -3437 0 net=8273
rlabel metal2 779 -3437 779 -3437 0 net=12515
rlabel metal2 821 -3437 821 -3437 0 net=752
rlabel metal2 310 -3439 310 -3439 0 net=1769
rlabel metal2 506 -3439 506 -3439 0 net=6791
rlabel metal2 653 -3439 653 -3439 0 net=5263
rlabel metal2 828 -3439 828 -3439 0 net=5589
rlabel metal2 933 -3439 933 -3439 0 net=2713
rlabel metal2 506 -3441 506 -3441 0 net=1496
rlabel metal2 674 -3441 674 -3441 0 net=8748
rlabel metal2 723 -3441 723 -3441 0 net=8557
rlabel metal2 835 -3441 835 -3441 0 net=8115
rlabel metal2 667 -3443 667 -3443 0 net=9417
rlabel metal2 723 -3443 723 -3443 0 net=7719
rlabel metal2 870 -3443 870 -3443 0 net=13133
rlabel metal2 614 -3445 614 -3445 0 net=3459
rlabel metal2 744 -3445 744 -3445 0 net=12091
rlabel metal2 870 -3445 870 -3445 0 net=1691
rlabel metal2 583 -3447 583 -3447 0 net=5937
rlabel metal2 583 -3449 583 -3449 0 net=6301
rlabel metal2 261 -3460 261 -3460 0 net=9647
rlabel metal2 296 -3460 296 -3460 0 net=1771
rlabel metal2 317 -3460 317 -3460 0 net=9492
rlabel metal2 359 -3460 359 -3460 0 net=6554
rlabel metal2 439 -3460 439 -3460 0 net=417
rlabel metal2 660 -3460 660 -3460 0 net=1232
rlabel metal2 737 -3460 737 -3460 0 net=10437
rlabel metal2 737 -3460 737 -3460 0 net=10437
rlabel metal2 793 -3460 793 -3460 0 net=12517
rlabel metal2 793 -3460 793 -3460 0 net=12517
rlabel metal2 800 -3460 800 -3460 0 net=5142
rlabel metal2 821 -3460 821 -3460 0 net=5590
rlabel metal2 842 -3460 842 -3460 0 net=4582
rlabel metal2 933 -3460 933 -3460 0 net=2715
rlabel metal2 933 -3460 933 -3460 0 net=2715
rlabel metal2 940 -3460 940 -3460 0 net=11293
rlabel metal2 947 -3460 947 -3460 0 net=13134
rlabel metal2 1010 -3460 1010 -3460 0 net=5651
rlabel metal2 1066 -3460 1066 -3460 0 net=11259
rlabel metal2 1087 -3460 1087 -3460 0 net=11562
rlabel metal2 1115 -3460 1115 -3460 0 net=4087
rlabel metal2 1136 -3460 1136 -3460 0 net=11899
rlabel metal2 1136 -3460 1136 -3460 0 net=11899
rlabel metal2 1143 -3460 1143 -3460 0 net=12109
rlabel metal2 1181 -3460 1181 -3460 0 net=9057
rlabel metal2 1577 -3460 1577 -3460 0 net=13707
rlabel metal2 1577 -3460 1577 -3460 0 net=13707
rlabel metal2 373 -3462 373 -3462 0 net=2780
rlabel metal2 401 -3462 401 -3462 0 net=2732
rlabel metal2 604 -3462 604 -3462 0 net=12523
rlabel metal2 604 -3462 604 -3462 0 net=12523
rlabel metal2 611 -3462 611 -3462 0 net=3006
rlabel metal2 786 -3462 786 -3462 0 net=2709
rlabel metal2 807 -3462 807 -3462 0 net=8367
rlabel metal2 828 -3462 828 -3462 0 net=1693
rlabel metal2 877 -3462 877 -3462 0 net=7053
rlabel metal2 877 -3462 877 -3462 0 net=7053
rlabel metal2 940 -3462 940 -3462 0 net=12481
rlabel metal2 968 -3462 968 -3462 0 net=12630
rlabel metal2 989 -3462 989 -3462 0 net=11151
rlabel metal2 1017 -3462 1017 -3462 0 net=7707
rlabel metal2 1052 -3462 1052 -3462 0 net=7791
rlabel metal2 1052 -3462 1052 -3462 0 net=7791
rlabel metal2 1073 -3462 1073 -3462 0 net=10501
rlabel metal2 1185 -3462 1185 -3462 0 net=12255
rlabel metal2 1213 -3462 1213 -3462 0 net=3647
rlabel metal2 1269 -3462 1269 -3462 0 net=13017
rlabel metal2 1297 -3462 1297 -3462 0 net=9852
rlabel metal2 1374 -3462 1374 -3462 0 net=12887
rlabel metal2 1388 -3462 1388 -3462 0 net=11979
rlabel metal2 1388 -3462 1388 -3462 0 net=11979
rlabel metal2 1395 -3462 1395 -3462 0 net=12323
rlabel metal2 1395 -3462 1395 -3462 0 net=12323
rlabel metal2 345 -3464 345 -3464 0 net=3691
rlabel metal2 380 -3464 380 -3464 0 net=3937
rlabel metal2 485 -3464 485 -3464 0 net=3755
rlabel metal2 485 -3464 485 -3464 0 net=3755
rlabel metal2 520 -3464 520 -3464 0 net=3596
rlabel metal2 618 -3464 618 -3464 0 net=11768
rlabel metal2 632 -3464 632 -3464 0 net=7528
rlabel metal2 667 -3464 667 -3464 0 net=3460
rlabel metal2 765 -3464 765 -3464 0 net=8275
rlabel metal2 852 -3464 852 -3464 0 net=13122
rlabel metal2 975 -3464 975 -3464 0 net=7827
rlabel metal2 1080 -3464 1080 -3464 0 net=10393
rlabel metal2 1300 -3464 1300 -3464 0 net=12814
rlabel metal2 1346 -3464 1346 -3464 0 net=11446
rlabel metal2 366 -3466 366 -3466 0 net=3033
rlabel metal2 387 -3466 387 -3466 0 net=3048
rlabel metal2 506 -3466 506 -3466 0 net=12673
rlabel metal2 618 -3466 618 -3466 0 net=7721
rlabel metal2 758 -3466 758 -3466 0 net=10839
rlabel metal2 772 -3466 772 -3466 0 net=8559
rlabel metal2 856 -3466 856 -3466 0 net=5939
rlabel metal2 975 -3466 975 -3466 0 net=2553
rlabel metal2 1024 -3466 1024 -3466 0 net=12291
rlabel metal2 1024 -3466 1024 -3466 0 net=12291
rlabel metal2 1115 -3466 1115 -3466 0 net=10991
rlabel metal2 1192 -3466 1192 -3466 0 net=3349
rlabel metal2 1192 -3466 1192 -3466 0 net=3349
rlabel metal2 1199 -3466 1199 -3466 0 net=8083
rlabel metal2 338 -3468 338 -3468 0 net=2687
rlabel metal2 450 -3468 450 -3468 0 net=5217
rlabel metal2 527 -3468 527 -3468 0 net=1784
rlabel metal2 639 -3468 639 -3468 0 net=5707
rlabel metal2 639 -3468 639 -3468 0 net=5707
rlabel metal2 653 -3468 653 -3468 0 net=11750
rlabel metal2 695 -3468 695 -3468 0 net=8621
rlabel metal2 891 -3468 891 -3468 0 net=5645
rlabel metal2 926 -3468 926 -3468 0 net=6303
rlabel metal2 1118 -3468 1118 -3468 0 net=1
rlabel metal2 429 -3470 429 -3470 0 net=4137
rlabel metal2 499 -3470 499 -3470 0 net=2989
rlabel metal2 534 -3470 534 -3470 0 net=7209
rlabel metal2 653 -3470 653 -3470 0 net=30
rlabel metal2 394 -3472 394 -3472 0 net=3863
rlabel metal2 457 -3472 457 -3472 0 net=3239
rlabel metal2 534 -3472 534 -3472 0 net=2813
rlabel metal2 695 -3472 695 -3472 0 net=12093
rlabel metal2 884 -3472 884 -3472 0 net=8997
rlabel metal2 905 -3472 905 -3472 0 net=10287
rlabel metal2 1003 -3472 1003 -3472 0 net=1362
rlabel metal2 436 -3474 436 -3474 0 net=4253
rlabel metal2 541 -3474 541 -3474 0 net=8532
rlabel metal2 702 -3474 702 -3474 0 net=9551
rlabel metal2 723 -3474 723 -3474 0 net=11822
rlabel metal2 863 -3474 863 -3474 0 net=6535
rlabel metal2 898 -3474 898 -3474 0 net=11479
rlabel metal2 478 -3476 478 -3476 0 net=4933
rlabel metal2 548 -3476 548 -3476 0 net=7550
rlabel metal2 688 -3476 688 -3476 0 net=13595
rlabel metal2 709 -3476 709 -3476 0 net=9691
rlabel metal2 898 -3476 898 -3476 0 net=10535
rlabel metal2 464 -3478 464 -3478 0 net=4001
rlabel metal2 548 -3478 548 -3478 0 net=7939
rlabel metal2 646 -3478 646 -3478 0 net=8229
rlabel metal2 730 -3478 730 -3478 0 net=6049
rlabel metal2 779 -3478 779 -3478 0 net=5264
rlabel metal2 555 -3480 555 -3480 0 net=6793
rlabel metal2 674 -3480 674 -3480 0 net=9419
rlabel metal2 730 -3480 730 -3480 0 net=8116
rlabel metal2 492 -3482 492 -3482 0 net=5293
rlabel metal2 562 -3482 562 -3482 0 net=12497
rlabel metal2 744 -3482 744 -3482 0 net=13493
rlabel metal2 443 -3484 443 -3484 0 net=3825
rlabel metal2 513 -3484 513 -3484 0 net=2851
rlabel metal2 569 -3484 569 -3484 0 net=6187
rlabel metal2 996 -3484 996 -3484 0 net=12203
rlabel metal2 415 -3486 415 -3486 0 net=5089
rlabel metal2 569 -3486 569 -3486 0 net=4159
rlabel metal2 422 -3488 422 -3488 0 net=6513
rlabel metal2 422 -3490 422 -3490 0 net=10007
rlabel metal2 268 -3501 268 -3501 0 net=9648
rlabel metal2 285 -3501 285 -3501 0 net=1772
rlabel metal2 366 -3501 366 -3501 0 net=2689
rlabel metal2 390 -3501 390 -3501 0 net=7259
rlabel metal2 408 -3501 408 -3501 0 net=3938
rlabel metal2 450 -3501 450 -3501 0 net=4138
rlabel metal2 506 -3501 506 -3501 0 net=5218
rlabel metal2 583 -3501 583 -3501 0 net=6795
rlabel metal2 604 -3501 604 -3501 0 net=12525
rlabel metal2 604 -3501 604 -3501 0 net=12525
rlabel metal2 632 -3501 632 -3501 0 net=7210
rlabel metal2 733 -3501 733 -3501 0 net=520
rlabel metal2 1192 -3501 1192 -3501 0 net=3351
rlabel metal2 1192 -3501 1192 -3501 0 net=3351
rlabel metal2 1234 -3501 1234 -3501 0 net=8084
rlabel metal2 1374 -3501 1374 -3501 0 net=12889
rlabel metal2 1384 -3501 1384 -3501 0 net=11980
rlabel metal2 1395 -3501 1395 -3501 0 net=12325
rlabel metal2 1395 -3501 1395 -3501 0 net=12325
rlabel metal2 1416 -3501 1416 -3501 0 net=9059
rlabel metal2 1577 -3501 1577 -3501 0 net=13708
rlabel metal2 1577 -3501 1577 -3501 0 net=13708
rlabel metal2 373 -3503 373 -3503 0 net=3693
rlabel metal2 443 -3503 443 -3503 0 net=5091
rlabel metal2 457 -3503 457 -3503 0 net=4255
rlabel metal2 492 -3503 492 -3503 0 net=3827
rlabel metal2 520 -3503 520 -3503 0 net=7940
rlabel metal2 562 -3503 562 -3503 0 net=2853
rlabel metal2 590 -3503 590 -3503 0 net=12674
rlabel metal2 674 -3503 674 -3503 0 net=12095
rlabel metal2 702 -3503 702 -3503 0 net=13597
rlabel metal2 702 -3503 702 -3503 0 net=13597
rlabel metal2 737 -3503 737 -3503 0 net=10438
rlabel metal2 758 -3503 758 -3503 0 net=8623
rlabel metal2 786 -3503 786 -3503 0 net=8277
rlabel metal2 821 -3503 821 -3503 0 net=9693
rlabel metal2 905 -3503 905 -3503 0 net=11480
rlabel metal2 940 -3503 940 -3503 0 net=12483
rlabel metal2 940 -3503 940 -3503 0 net=12483
rlabel metal2 947 -3503 947 -3503 0 net=5940
rlabel metal2 1045 -3503 1045 -3503 0 net=7709
rlabel metal2 1059 -3503 1059 -3503 0 net=5652
rlabel metal2 1115 -3503 1115 -3503 0 net=10993
rlabel metal2 1115 -3503 1115 -3503 0 net=10993
rlabel metal2 1122 -3503 1122 -3503 0 net=4089
rlabel metal2 1136 -3503 1136 -3503 0 net=11901
rlabel metal2 1136 -3503 1136 -3503 0 net=11901
rlabel metal2 1157 -3503 1157 -3503 0 net=12111
rlabel metal2 1178 -3503 1178 -3503 0 net=12257
rlabel metal2 1248 -3503 1248 -3503 0 net=3649
rlabel metal2 1269 -3503 1269 -3503 0 net=10395
rlabel metal2 380 -3505 380 -3505 0 net=3035
rlabel metal2 380 -3505 380 -3505 0 net=3035
rlabel metal2 429 -3505 429 -3505 0 net=3865
rlabel metal2 478 -3505 478 -3505 0 net=4003
rlabel metal2 527 -3505 527 -3505 0 net=2990
rlabel metal2 576 -3505 576 -3505 0 net=12499
rlabel metal2 646 -3505 646 -3505 0 net=6188
rlabel metal2 758 -3505 758 -3505 0 net=6051
rlabel metal2 786 -3505 786 -3505 0 net=12519
rlabel metal2 800 -3505 800 -3505 0 net=2710
rlabel metal2 842 -3505 842 -3505 0 net=6555
rlabel metal2 1020 -3505 1020 -3505 0 net=10502
rlabel metal2 1080 -3505 1080 -3505 0 net=6305
rlabel metal2 1276 -3505 1276 -3505 0 net=13018
rlabel metal2 1276 -3505 1276 -3505 0 net=13018
rlabel metal2 429 -3507 429 -3507 0 net=12337
rlabel metal2 499 -3507 499 -3507 0 net=3241
rlabel metal2 541 -3507 541 -3507 0 net=4935
rlabel metal2 576 -3507 576 -3507 0 net=7723
rlabel metal2 639 -3507 639 -3507 0 net=5709
rlabel metal2 653 -3507 653 -3507 0 net=13495
rlabel metal2 765 -3507 765 -3507 0 net=10841
rlabel metal2 800 -3507 800 -3507 0 net=8369
rlabel metal2 884 -3507 884 -3507 0 net=6537
rlabel metal2 957 -3507 957 -3507 0 net=12204
rlabel metal2 1003 -3507 1003 -3507 0 net=1215
rlabel metal2 1003 -3507 1003 -3507 0 net=1215
rlabel metal2 1010 -3507 1010 -3507 0 net=11152
rlabel metal2 1045 -3507 1045 -3507 0 net=7793
rlabel metal2 1062 -3507 1062 -3507 0 net=11260
rlabel metal2 485 -3509 485 -3509 0 net=3757
rlabel metal2 513 -3509 513 -3509 0 net=6515
rlabel metal2 688 -3509 688 -3509 0 net=9421
rlabel metal2 709 -3509 709 -3509 0 net=8231
rlabel metal2 807 -3509 807 -3509 0 net=8561
rlabel metal2 877 -3509 877 -3509 0 net=7055
rlabel metal2 961 -3509 961 -3509 0 net=12088
rlabel metal2 968 -3509 968 -3509 0 net=2555
rlabel metal2 1024 -3509 1024 -3509 0 net=12292
rlabel metal2 1038 -3509 1038 -3509 0 net=7829
rlabel metal2 471 -3511 471 -3511 0 net=10009
rlabel metal2 513 -3511 513 -3511 0 net=2815
rlabel metal2 709 -3511 709 -3511 0 net=9553
rlabel metal2 765 -3511 765 -3511 0 net=13171
rlabel metal2 1048 -3511 1048 -3511 0 net=1
rlabel metal2 534 -3513 534 -3513 0 net=4161
rlabel metal2 814 -3513 814 -3513 0 net=1695
rlabel metal2 877 -3513 877 -3513 0 net=10537
rlabel metal2 954 -3513 954 -3513 0 net=11294
rlabel metal2 555 -3515 555 -3515 0 net=5295
rlabel metal2 891 -3515 891 -3515 0 net=8999
rlabel metal2 926 -3515 926 -3515 0 net=10288
rlabel metal2 926 -3517 926 -3517 0 net=2717
rlabel metal2 919 -3519 919 -3519 0 net=5647
rlabel metal2 919 -3521 919 -3521 0 net=5075
rlabel metal2 380 -3532 380 -3532 0 net=3037
rlabel metal2 380 -3532 380 -3532 0 net=3037
rlabel metal2 387 -3532 387 -3532 0 net=2691
rlabel metal2 408 -3532 408 -3532 0 net=12339
rlabel metal2 450 -3532 450 -3532 0 net=5093
rlabel metal2 464 -3532 464 -3532 0 net=4256
rlabel metal2 478 -3532 478 -3532 0 net=10605
rlabel metal2 478 -3532 478 -3532 0 net=10605
rlabel metal2 506 -3532 506 -3532 0 net=3828
rlabel metal2 527 -3532 527 -3532 0 net=3242
rlabel metal2 527 -3532 527 -3532 0 net=3242
rlabel metal2 548 -3532 548 -3532 0 net=4937
rlabel metal2 548 -3532 548 -3532 0 net=4937
rlabel metal2 558 -3532 558 -3532 0 net=868
rlabel metal2 1115 -3532 1115 -3532 0 net=10995
rlabel metal2 1115 -3532 1115 -3532 0 net=10995
rlabel metal2 1129 -3532 1129 -3532 0 net=4091
rlabel metal2 1129 -3532 1129 -3532 0 net=4091
rlabel metal2 1136 -3532 1136 -3532 0 net=11903
rlabel metal2 1136 -3532 1136 -3532 0 net=11903
rlabel metal2 1157 -3532 1157 -3532 0 net=12112
rlabel metal2 1178 -3532 1178 -3532 0 net=12259
rlabel metal2 1178 -3532 1178 -3532 0 net=12259
rlabel metal2 1192 -3532 1192 -3532 0 net=3353
rlabel metal2 1192 -3532 1192 -3532 0 net=3353
rlabel metal2 1262 -3532 1262 -3532 0 net=3650
rlabel metal2 1339 -3532 1339 -3532 0 net=10397
rlabel metal2 1381 -3532 1381 -3532 0 net=12891
rlabel metal2 1395 -3532 1395 -3532 0 net=12327
rlabel metal2 1395 -3532 1395 -3532 0 net=12327
rlabel metal2 1500 -3532 1500 -3532 0 net=9060
rlabel metal2 387 -3534 387 -3534 0 net=3695
rlabel metal2 443 -3534 443 -3534 0 net=3867
rlabel metal2 506 -3534 506 -3534 0 net=2817
rlabel metal2 565 -3534 565 -3534 0 net=13496
rlabel metal2 660 -3534 660 -3534 0 net=12096
rlabel metal2 695 -3534 695 -3534 0 net=9422
rlabel metal2 730 -3534 730 -3534 0 net=8233
rlabel metal2 758 -3534 758 -3534 0 net=6053
rlabel metal2 758 -3534 758 -3534 0 net=6053
rlabel metal2 786 -3534 786 -3534 0 net=12521
rlabel metal2 786 -3534 786 -3534 0 net=12521
rlabel metal2 796 -3534 796 -3534 0 net=8370
rlabel metal2 807 -3534 807 -3534 0 net=8562
rlabel metal2 884 -3534 884 -3534 0 net=7056
rlabel metal2 898 -3534 898 -3534 0 net=9001
rlabel metal2 898 -3534 898 -3534 0 net=9001
rlabel metal2 905 -3534 905 -3534 0 net=6539
rlabel metal2 905 -3534 905 -3534 0 net=6539
rlabel metal2 926 -3534 926 -3534 0 net=2718
rlabel metal2 957 -3534 957 -3534 0 net=2556
rlabel metal2 1038 -3534 1038 -3534 0 net=7794
rlabel metal2 1052 -3534 1052 -3534 0 net=7710
rlabel metal2 1073 -3534 1073 -3534 0 net=7830
rlabel metal2 1143 -3534 1143 -3534 0 net=6307
rlabel metal2 394 -3536 394 -3536 0 net=7261
rlabel metal2 499 -3536 499 -3536 0 net=3759
rlabel metal2 565 -3536 565 -3536 0 net=7724
rlabel metal2 604 -3536 604 -3536 0 net=12526
rlabel metal2 646 -3536 646 -3536 0 net=5710
rlabel metal2 667 -3536 667 -3536 0 net=13173
rlabel metal2 779 -3536 779 -3536 0 net=8625
rlabel metal2 814 -3536 814 -3536 0 net=1697
rlabel metal2 814 -3536 814 -3536 0 net=1697
rlabel metal2 877 -3536 877 -3536 0 net=10539
rlabel metal2 919 -3536 919 -3536 0 net=5077
rlabel metal2 933 -3536 933 -3536 0 net=5648
rlabel metal2 940 -3536 940 -3536 0 net=12485
rlabel metal2 940 -3536 940 -3536 0 net=12485
rlabel metal2 492 -3538 492 -3538 0 net=4004
rlabel metal2 569 -3538 569 -3538 0 net=5297
rlabel metal2 569 -3538 569 -3538 0 net=5297
rlabel metal2 576 -3538 576 -3538 0 net=12500
rlabel metal2 702 -3538 702 -3538 0 net=9554
rlabel metal2 772 -3538 772 -3538 0 net=10843
rlabel metal2 793 -3538 793 -3538 0 net=8279
rlabel metal2 863 -3538 863 -3538 0 net=9695
rlabel metal2 485 -3540 485 -3540 0 net=10011
rlabel metal2 590 -3540 590 -3540 0 net=6797
rlabel metal2 772 -3540 772 -3540 0 net=6557
rlabel metal2 583 -3542 583 -3542 0 net=2855
rlabel metal2 555 -3544 555 -3544 0 net=2733
rlabel metal2 541 -3546 541 -3546 0 net=6517
rlabel metal2 534 -3548 534 -3548 0 net=4163
rlabel metal2 534 -3550 534 -3550 0 net=6469
rlabel metal2 387 -3561 387 -3561 0 net=3697
rlabel metal2 387 -3561 387 -3561 0 net=3697
rlabel metal2 394 -3561 394 -3561 0 net=2692
rlabel metal2 394 -3561 394 -3561 0 net=2692
rlabel metal2 401 -3561 401 -3561 0 net=7262
rlabel metal2 408 -3561 408 -3561 0 net=12341
rlabel metal2 408 -3561 408 -3561 0 net=12341
rlabel metal2 457 -3561 457 -3561 0 net=5095
rlabel metal2 474 -3561 474 -3561 0 net=10606
rlabel metal2 492 -3561 492 -3561 0 net=10013
rlabel metal2 492 -3561 492 -3561 0 net=10013
rlabel metal2 499 -3561 499 -3561 0 net=3760
rlabel metal2 527 -3561 527 -3561 0 net=4164
rlabel metal2 555 -3561 555 -3561 0 net=6518
rlabel metal2 569 -3561 569 -3561 0 net=5298
rlabel metal2 579 -3561 579 -3561 0 net=2856
rlabel metal2 632 -3561 632 -3561 0 net=13175
rlabel metal2 702 -3561 702 -3561 0 net=13600
rlabel metal2 737 -3561 737 -3561 0 net=8234
rlabel metal2 758 -3561 758 -3561 0 net=6054
rlabel metal2 768 -3561 768 -3561 0 net=10844
rlabel metal2 786 -3561 786 -3561 0 net=12522
rlabel metal2 800 -3561 800 -3561 0 net=8627
rlabel metal2 800 -3561 800 -3561 0 net=8627
rlabel metal2 877 -3561 877 -3561 0 net=9696
rlabel metal2 901 -3561 901 -3561 0 net=6540
rlabel metal2 926 -3561 926 -3561 0 net=5078
rlabel metal2 1111 -3561 1111 -3561 0 net=10996
rlabel metal2 1132 -3561 1132 -3561 0 net=11904
rlabel metal2 1164 -3561 1164 -3561 0 net=6309
rlabel metal2 1178 -3561 1178 -3561 0 net=12261
rlabel metal2 1192 -3561 1192 -3561 0 net=3355
rlabel metal2 1391 -3561 1391 -3561 0 net=12328
rlabel metal2 380 -3563 380 -3563 0 net=3038
rlabel metal2 450 -3563 450 -3563 0 net=3868
rlabel metal2 502 -3563 502 -3563 0 net=2818
rlabel metal2 530 -3563 530 -3563 0 net=6470
rlabel metal2 548 -3563 548 -3563 0 net=4939
rlabel metal2 576 -3563 576 -3563 0 net=2734
rlabel metal2 590 -3563 590 -3563 0 net=6799
rlabel metal2 590 -3563 590 -3563 0 net=6799
rlabel metal2 758 -3563 758 -3563 0 net=6559
rlabel metal2 793 -3563 793 -3563 0 net=8280
rlabel metal2 884 -3563 884 -3563 0 net=10541
rlabel metal2 884 -3563 884 -3563 0 net=10541
rlabel metal2 891 -3563 891 -3563 0 net=9002
rlabel metal2 933 -3563 933 -3563 0 net=12486
rlabel metal2 1129 -3563 1129 -3563 0 net=4093
rlabel metal2 1388 -3563 1388 -3563 0 net=12893
rlabel metal2 807 -3565 807 -3565 0 net=1698
rlabel metal2 1360 -3565 1360 -3565 0 net=10398
rlabel metal2 387 -3576 387 -3576 0 net=3698
rlabel metal2 457 -3576 457 -3576 0 net=5096
rlabel metal2 492 -3576 492 -3576 0 net=10014
rlabel metal2 562 -3576 562 -3576 0 net=4940
rlabel metal2 590 -3576 590 -3576 0 net=6800
rlabel metal2 600 -3576 600 -3576 0 net=13176
rlabel metal2 747 -3576 747 -3576 0 net=6560
rlabel metal2 800 -3576 800 -3576 0 net=8628
rlabel metal2 884 -3576 884 -3576 0 net=10542
rlabel metal2 1129 -3576 1129 -3576 0 net=4094
rlabel metal2 1171 -3576 1171 -3576 0 net=6310
rlabel metal2 1195 -3576 1195 -3576 0 net=3356
rlabel metal2 1388 -3576 1388 -3576 0 net=12894
rlabel metal2 397 -3578 397 -3578 0 net=12342
rlabel metal2 1178 -3578 1178 -3578 0 net=12262
<< end >>
