magic
tech scmos
timestamp 1555017904 
<< pdiffusion >>
rect 1 -10 7 -4
rect 8 -10 14 -4
rect 15 -10 21 -4
rect 22 -10 28 -4
rect 29 -10 35 -4
rect 36 -10 42 -4
rect 85 -10 91 -4
rect 92 -10 95 -4
rect 99 -10 105 -4
rect 106 -10 112 -4
rect 113 -10 119 -4
rect 120 -10 123 -4
rect 127 -10 130 -4
rect 141 -10 147 -4
rect 204 -10 207 -4
rect 211 -10 217 -4
rect 218 -10 224 -4
rect 225 -10 228 -4
rect 232 -10 238 -4
rect 239 -10 242 -4
rect 246 -10 252 -4
rect 253 -10 259 -4
rect 260 -10 266 -4
rect 267 -10 270 -4
rect 281 -10 287 -4
rect 323 -10 326 -4
rect 330 -10 336 -4
rect 337 -10 343 -4
rect 428 -10 431 -4
rect 449 -10 455 -4
rect 463 -10 466 -4
rect 484 -10 490 -4
rect 505 -10 511 -4
rect 526 -10 532 -4
rect 533 -10 536 -4
rect 547 -10 553 -4
rect 582 -10 588 -4
rect 589 -10 595 -4
rect 596 -10 599 -4
rect 603 -10 609 -4
rect 659 -10 665 -4
rect 666 -10 669 -4
rect 1 -29 7 -23
rect 8 -29 14 -23
rect 15 -29 21 -23
rect 22 -29 28 -23
rect 29 -29 35 -23
rect 99 -29 105 -23
rect 113 -29 119 -23
rect 134 -29 137 -23
rect 169 -29 175 -23
rect 176 -29 179 -23
rect 183 -29 186 -23
rect 190 -29 196 -23
rect 197 -29 200 -23
rect 204 -29 210 -23
rect 211 -29 217 -23
rect 218 -29 221 -23
rect 225 -29 228 -23
rect 232 -29 238 -23
rect 239 -29 245 -23
rect 246 -29 249 -23
rect 253 -29 256 -23
rect 260 -29 263 -23
rect 267 -29 270 -23
rect 274 -29 277 -23
rect 281 -29 284 -23
rect 288 -29 291 -23
rect 295 -29 301 -23
rect 302 -29 308 -23
rect 309 -29 312 -23
rect 316 -29 319 -23
rect 323 -29 326 -23
rect 330 -29 336 -23
rect 337 -29 343 -23
rect 344 -29 350 -23
rect 358 -29 361 -23
rect 372 -29 375 -23
rect 379 -29 385 -23
rect 414 -29 417 -23
rect 421 -29 427 -23
rect 428 -29 431 -23
rect 435 -29 441 -23
rect 442 -29 448 -23
rect 449 -29 455 -23
rect 463 -29 469 -23
rect 470 -29 473 -23
rect 491 -29 494 -23
rect 505 -29 508 -23
rect 512 -29 518 -23
rect 519 -29 525 -23
rect 526 -29 529 -23
rect 540 -29 543 -23
rect 554 -29 560 -23
rect 561 -29 567 -23
rect 568 -29 571 -23
rect 575 -29 578 -23
rect 603 -29 606 -23
rect 610 -29 613 -23
rect 617 -29 620 -23
rect 673 -29 676 -23
rect 1 -60 7 -54
rect 8 -60 14 -54
rect 15 -60 21 -54
rect 22 -60 28 -54
rect 85 -60 88 -54
rect 92 -60 95 -54
rect 113 -60 116 -54
rect 120 -60 123 -54
rect 127 -60 130 -54
rect 134 -60 137 -54
rect 141 -60 147 -54
rect 148 -60 154 -54
rect 155 -60 158 -54
rect 162 -60 165 -54
rect 169 -60 175 -54
rect 176 -60 182 -54
rect 183 -60 189 -54
rect 190 -60 193 -54
rect 197 -60 203 -54
rect 204 -60 207 -54
rect 211 -60 214 -54
rect 218 -60 221 -54
rect 225 -60 228 -54
rect 232 -60 238 -54
rect 239 -60 245 -54
rect 246 -60 252 -54
rect 253 -60 256 -54
rect 260 -60 263 -54
rect 267 -60 270 -54
rect 274 -60 280 -54
rect 281 -60 284 -54
rect 288 -60 291 -54
rect 295 -60 301 -54
rect 302 -60 305 -54
rect 309 -60 315 -54
rect 316 -60 319 -54
rect 323 -60 326 -54
rect 330 -60 333 -54
rect 337 -60 343 -54
rect 344 -60 347 -54
rect 351 -60 354 -54
rect 358 -60 364 -54
rect 365 -60 368 -54
rect 372 -60 378 -54
rect 379 -60 385 -54
rect 386 -60 389 -54
rect 393 -60 396 -54
rect 400 -60 403 -54
rect 407 -60 410 -54
rect 414 -60 420 -54
rect 421 -60 424 -54
rect 428 -60 431 -54
rect 435 -60 438 -54
rect 442 -60 445 -54
rect 463 -60 469 -54
rect 470 -60 473 -54
rect 477 -60 480 -54
rect 484 -60 487 -54
rect 491 -60 497 -54
rect 498 -60 501 -54
rect 505 -60 508 -54
rect 519 -60 522 -54
rect 526 -60 532 -54
rect 533 -60 536 -54
rect 540 -60 543 -54
rect 547 -60 553 -54
rect 554 -60 560 -54
rect 561 -60 564 -54
rect 568 -60 571 -54
rect 575 -60 578 -54
rect 582 -60 588 -54
rect 589 -60 592 -54
rect 596 -60 599 -54
rect 603 -60 606 -54
rect 610 -60 613 -54
rect 624 -60 627 -54
rect 631 -60 634 -54
rect 638 -60 641 -54
rect 645 -60 648 -54
rect 652 -60 655 -54
rect 659 -60 665 -54
rect 666 -60 669 -54
rect 673 -60 679 -54
rect 680 -60 683 -54
rect 701 -60 704 -54
rect 764 -60 770 -54
rect 771 -60 774 -54
rect 841 -60 844 -54
rect 1 -129 7 -123
rect 8 -129 14 -123
rect 15 -129 21 -123
rect 22 -129 28 -123
rect 29 -129 32 -123
rect 36 -129 39 -123
rect 43 -129 49 -123
rect 50 -129 56 -123
rect 57 -129 63 -123
rect 64 -129 67 -123
rect 71 -129 74 -123
rect 78 -129 84 -123
rect 85 -129 88 -123
rect 92 -129 95 -123
rect 99 -129 105 -123
rect 106 -129 109 -123
rect 113 -129 119 -123
rect 120 -129 123 -123
rect 127 -129 133 -123
rect 134 -129 140 -123
rect 141 -129 144 -123
rect 148 -129 154 -123
rect 155 -129 161 -123
rect 162 -129 165 -123
rect 169 -129 175 -123
rect 176 -129 179 -123
rect 183 -129 186 -123
rect 190 -129 193 -123
rect 197 -129 200 -123
rect 204 -129 207 -123
rect 211 -129 214 -123
rect 218 -129 221 -123
rect 225 -129 231 -123
rect 232 -129 235 -123
rect 239 -129 242 -123
rect 246 -129 252 -123
rect 253 -129 256 -123
rect 260 -129 263 -123
rect 267 -129 270 -123
rect 274 -129 280 -123
rect 281 -129 284 -123
rect 288 -129 291 -123
rect 295 -129 298 -123
rect 302 -129 305 -123
rect 309 -129 312 -123
rect 316 -129 322 -123
rect 323 -129 326 -123
rect 330 -129 333 -123
rect 337 -129 340 -123
rect 344 -129 350 -123
rect 351 -129 357 -123
rect 358 -129 361 -123
rect 365 -129 368 -123
rect 372 -129 378 -123
rect 379 -129 382 -123
rect 386 -129 392 -123
rect 393 -129 399 -123
rect 400 -129 403 -123
rect 407 -129 410 -123
rect 414 -129 420 -123
rect 421 -129 424 -123
rect 428 -129 431 -123
rect 435 -129 438 -123
rect 442 -129 445 -123
rect 449 -129 452 -123
rect 456 -129 459 -123
rect 463 -129 466 -123
rect 470 -129 473 -123
rect 477 -129 480 -123
rect 484 -129 487 -123
rect 491 -129 494 -123
rect 498 -129 504 -123
rect 505 -129 511 -123
rect 512 -129 515 -123
rect 519 -129 522 -123
rect 526 -129 529 -123
rect 533 -129 536 -123
rect 540 -129 543 -123
rect 547 -129 550 -123
rect 554 -129 557 -123
rect 561 -129 564 -123
rect 568 -129 571 -123
rect 575 -129 578 -123
rect 582 -129 588 -123
rect 589 -129 592 -123
rect 596 -129 599 -123
rect 603 -129 606 -123
rect 610 -129 613 -123
rect 617 -129 620 -123
rect 624 -129 627 -123
rect 631 -129 634 -123
rect 638 -129 641 -123
rect 645 -129 648 -123
rect 652 -129 655 -123
rect 659 -129 665 -123
rect 666 -129 669 -123
rect 673 -129 676 -123
rect 680 -129 683 -123
rect 687 -129 690 -123
rect 694 -129 697 -123
rect 701 -129 704 -123
rect 708 -129 711 -123
rect 715 -129 718 -123
rect 722 -129 725 -123
rect 729 -129 732 -123
rect 736 -129 739 -123
rect 743 -129 746 -123
rect 750 -129 753 -123
rect 757 -129 760 -123
rect 764 -129 767 -123
rect 771 -129 774 -123
rect 778 -129 781 -123
rect 785 -129 788 -123
rect 792 -129 795 -123
rect 799 -129 802 -123
rect 806 -129 809 -123
rect 813 -129 816 -123
rect 820 -129 823 -123
rect 827 -129 830 -123
rect 834 -129 837 -123
rect 841 -129 847 -123
rect 869 -129 872 -123
rect 876 -129 879 -123
rect 1107 -129 1113 -123
rect 1 -218 7 -212
rect 8 -218 14 -212
rect 15 -218 21 -212
rect 22 -218 25 -212
rect 29 -218 32 -212
rect 36 -218 39 -212
rect 43 -218 46 -212
rect 50 -218 53 -212
rect 57 -218 60 -212
rect 64 -218 67 -212
rect 71 -218 77 -212
rect 78 -218 81 -212
rect 85 -218 91 -212
rect 92 -218 95 -212
rect 99 -218 102 -212
rect 106 -218 112 -212
rect 113 -218 116 -212
rect 120 -218 126 -212
rect 127 -218 130 -212
rect 134 -218 137 -212
rect 141 -218 147 -212
rect 148 -218 154 -212
rect 155 -218 158 -212
rect 162 -218 165 -212
rect 169 -218 172 -212
rect 176 -218 182 -212
rect 183 -218 186 -212
rect 190 -218 193 -212
rect 197 -218 200 -212
rect 204 -218 210 -212
rect 211 -218 217 -212
rect 218 -218 224 -212
rect 225 -218 231 -212
rect 232 -218 238 -212
rect 239 -218 242 -212
rect 246 -218 252 -212
rect 253 -218 256 -212
rect 260 -218 263 -212
rect 267 -218 270 -212
rect 274 -218 277 -212
rect 281 -218 284 -212
rect 288 -218 291 -212
rect 295 -218 301 -212
rect 302 -218 305 -212
rect 309 -218 312 -212
rect 316 -218 319 -212
rect 323 -218 329 -212
rect 330 -218 336 -212
rect 337 -218 340 -212
rect 344 -218 350 -212
rect 351 -218 354 -212
rect 358 -218 364 -212
rect 365 -218 368 -212
rect 372 -218 375 -212
rect 379 -218 382 -212
rect 386 -218 392 -212
rect 393 -218 399 -212
rect 400 -218 406 -212
rect 407 -218 410 -212
rect 414 -218 417 -212
rect 421 -218 424 -212
rect 428 -218 431 -212
rect 435 -218 438 -212
rect 442 -218 445 -212
rect 449 -218 452 -212
rect 456 -218 462 -212
rect 463 -218 466 -212
rect 470 -218 473 -212
rect 477 -218 480 -212
rect 484 -218 487 -212
rect 491 -218 497 -212
rect 498 -218 501 -212
rect 505 -218 508 -212
rect 512 -218 515 -212
rect 519 -218 525 -212
rect 526 -218 529 -212
rect 533 -218 536 -212
rect 540 -218 543 -212
rect 547 -218 550 -212
rect 554 -218 557 -212
rect 561 -218 564 -212
rect 568 -218 571 -212
rect 575 -218 581 -212
rect 582 -218 585 -212
rect 589 -218 592 -212
rect 596 -218 599 -212
rect 603 -218 606 -212
rect 610 -218 613 -212
rect 617 -218 623 -212
rect 624 -218 630 -212
rect 631 -218 634 -212
rect 638 -218 641 -212
rect 645 -218 648 -212
rect 652 -218 658 -212
rect 659 -218 662 -212
rect 666 -218 669 -212
rect 673 -218 676 -212
rect 680 -218 683 -212
rect 687 -218 690 -212
rect 694 -218 697 -212
rect 701 -218 704 -212
rect 708 -218 711 -212
rect 715 -218 718 -212
rect 722 -218 725 -212
rect 729 -218 732 -212
rect 736 -218 742 -212
rect 743 -218 746 -212
rect 750 -218 753 -212
rect 757 -218 760 -212
rect 764 -218 767 -212
rect 771 -218 774 -212
rect 778 -218 781 -212
rect 785 -218 788 -212
rect 792 -218 795 -212
rect 799 -218 802 -212
rect 806 -218 809 -212
rect 813 -218 816 -212
rect 820 -218 823 -212
rect 827 -218 830 -212
rect 834 -218 837 -212
rect 841 -218 844 -212
rect 848 -218 851 -212
rect 855 -218 858 -212
rect 862 -218 865 -212
rect 869 -218 872 -212
rect 876 -218 879 -212
rect 883 -218 886 -212
rect 890 -218 893 -212
rect 897 -218 900 -212
rect 904 -218 907 -212
rect 911 -218 914 -212
rect 918 -218 921 -212
rect 925 -218 928 -212
rect 932 -218 935 -212
rect 939 -218 942 -212
rect 946 -218 949 -212
rect 953 -218 956 -212
rect 1107 -218 1110 -212
rect 1 -301 7 -295
rect 8 -301 14 -295
rect 15 -301 18 -295
rect 22 -301 25 -295
rect 29 -301 32 -295
rect 36 -301 39 -295
rect 43 -301 49 -295
rect 50 -301 53 -295
rect 57 -301 60 -295
rect 64 -301 70 -295
rect 71 -301 74 -295
rect 78 -301 81 -295
rect 85 -301 88 -295
rect 92 -301 95 -295
rect 99 -301 105 -295
rect 106 -301 109 -295
rect 113 -301 119 -295
rect 120 -301 126 -295
rect 127 -301 133 -295
rect 134 -301 140 -295
rect 141 -301 144 -295
rect 148 -301 151 -295
rect 155 -301 158 -295
rect 162 -301 168 -295
rect 169 -301 175 -295
rect 176 -301 179 -295
rect 183 -301 189 -295
rect 190 -301 196 -295
rect 197 -301 200 -295
rect 204 -301 210 -295
rect 211 -301 214 -295
rect 218 -301 221 -295
rect 225 -301 228 -295
rect 232 -301 235 -295
rect 239 -301 242 -295
rect 246 -301 249 -295
rect 253 -301 259 -295
rect 260 -301 263 -295
rect 267 -301 270 -295
rect 274 -301 277 -295
rect 281 -301 284 -295
rect 288 -301 291 -295
rect 295 -301 301 -295
rect 302 -301 305 -295
rect 309 -301 312 -295
rect 316 -301 322 -295
rect 323 -301 326 -295
rect 330 -301 333 -295
rect 337 -301 340 -295
rect 344 -301 347 -295
rect 351 -301 357 -295
rect 358 -301 364 -295
rect 365 -301 368 -295
rect 372 -301 378 -295
rect 379 -301 382 -295
rect 386 -301 389 -295
rect 393 -301 399 -295
rect 400 -301 406 -295
rect 407 -301 410 -295
rect 414 -301 417 -295
rect 421 -301 424 -295
rect 428 -301 431 -295
rect 435 -301 441 -295
rect 442 -301 445 -295
rect 449 -301 452 -295
rect 456 -301 459 -295
rect 463 -301 469 -295
rect 470 -301 473 -295
rect 477 -301 480 -295
rect 484 -301 490 -295
rect 491 -301 494 -295
rect 498 -301 504 -295
rect 505 -301 508 -295
rect 512 -301 515 -295
rect 519 -301 525 -295
rect 526 -301 529 -295
rect 533 -301 536 -295
rect 540 -301 543 -295
rect 547 -301 550 -295
rect 554 -301 557 -295
rect 561 -301 564 -295
rect 568 -301 571 -295
rect 575 -301 578 -295
rect 582 -301 585 -295
rect 589 -301 592 -295
rect 596 -301 599 -295
rect 603 -301 606 -295
rect 610 -301 613 -295
rect 617 -301 620 -295
rect 624 -301 627 -295
rect 631 -301 634 -295
rect 638 -301 641 -295
rect 645 -301 648 -295
rect 652 -301 655 -295
rect 659 -301 665 -295
rect 666 -301 669 -295
rect 673 -301 676 -295
rect 680 -301 683 -295
rect 687 -301 690 -295
rect 694 -301 697 -295
rect 701 -301 704 -295
rect 708 -301 711 -295
rect 715 -301 718 -295
rect 722 -301 725 -295
rect 729 -301 732 -295
rect 736 -301 739 -295
rect 743 -301 746 -295
rect 750 -301 753 -295
rect 757 -301 760 -295
rect 764 -301 767 -295
rect 771 -301 774 -295
rect 778 -301 781 -295
rect 785 -301 788 -295
rect 792 -301 795 -295
rect 799 -301 802 -295
rect 806 -301 809 -295
rect 813 -301 816 -295
rect 820 -301 823 -295
rect 827 -301 830 -295
rect 834 -301 837 -295
rect 841 -301 844 -295
rect 848 -301 851 -295
rect 855 -301 858 -295
rect 862 -301 865 -295
rect 869 -301 872 -295
rect 876 -301 879 -295
rect 883 -301 889 -295
rect 890 -301 896 -295
rect 897 -301 903 -295
rect 904 -301 910 -295
rect 911 -301 914 -295
rect 918 -301 921 -295
rect 1107 -301 1110 -295
rect 1 -396 7 -390
rect 8 -396 11 -390
rect 15 -396 21 -390
rect 22 -396 25 -390
rect 29 -396 35 -390
rect 36 -396 39 -390
rect 43 -396 46 -390
rect 50 -396 53 -390
rect 57 -396 60 -390
rect 64 -396 70 -390
rect 71 -396 74 -390
rect 78 -396 84 -390
rect 85 -396 88 -390
rect 92 -396 98 -390
rect 99 -396 102 -390
rect 106 -396 112 -390
rect 113 -396 119 -390
rect 120 -396 126 -390
rect 127 -396 130 -390
rect 134 -396 140 -390
rect 141 -396 144 -390
rect 148 -396 151 -390
rect 155 -396 161 -390
rect 162 -396 165 -390
rect 169 -396 175 -390
rect 176 -396 179 -390
rect 183 -396 189 -390
rect 190 -396 193 -390
rect 197 -396 200 -390
rect 204 -396 207 -390
rect 211 -396 217 -390
rect 218 -396 221 -390
rect 225 -396 228 -390
rect 232 -396 235 -390
rect 239 -396 242 -390
rect 246 -396 252 -390
rect 253 -396 259 -390
rect 260 -396 266 -390
rect 267 -396 270 -390
rect 274 -396 277 -390
rect 281 -396 284 -390
rect 288 -396 291 -390
rect 295 -396 298 -390
rect 302 -396 308 -390
rect 309 -396 312 -390
rect 316 -396 322 -390
rect 323 -396 329 -390
rect 330 -396 333 -390
rect 337 -396 343 -390
rect 344 -396 347 -390
rect 351 -396 354 -390
rect 358 -396 361 -390
rect 365 -396 368 -390
rect 372 -396 378 -390
rect 379 -396 385 -390
rect 386 -396 389 -390
rect 393 -396 399 -390
rect 400 -396 403 -390
rect 407 -396 410 -390
rect 414 -396 417 -390
rect 421 -396 424 -390
rect 428 -396 431 -390
rect 435 -396 438 -390
rect 442 -396 445 -390
rect 449 -396 452 -390
rect 456 -396 459 -390
rect 463 -396 466 -390
rect 470 -396 476 -390
rect 477 -396 480 -390
rect 484 -396 487 -390
rect 491 -396 497 -390
rect 498 -396 501 -390
rect 505 -396 508 -390
rect 512 -396 518 -390
rect 519 -396 522 -390
rect 526 -396 529 -390
rect 533 -396 536 -390
rect 540 -396 546 -390
rect 547 -396 550 -390
rect 554 -396 557 -390
rect 561 -396 564 -390
rect 568 -396 571 -390
rect 575 -396 578 -390
rect 582 -396 585 -390
rect 589 -396 592 -390
rect 596 -396 599 -390
rect 603 -396 606 -390
rect 610 -396 613 -390
rect 617 -396 620 -390
rect 624 -396 630 -390
rect 631 -396 634 -390
rect 638 -396 641 -390
rect 645 -396 648 -390
rect 652 -396 655 -390
rect 659 -396 662 -390
rect 666 -396 672 -390
rect 673 -396 676 -390
rect 680 -396 683 -390
rect 687 -396 690 -390
rect 694 -396 697 -390
rect 701 -396 704 -390
rect 708 -396 711 -390
rect 715 -396 718 -390
rect 722 -396 725 -390
rect 729 -396 732 -390
rect 736 -396 739 -390
rect 743 -396 746 -390
rect 750 -396 753 -390
rect 757 -396 760 -390
rect 764 -396 767 -390
rect 771 -396 774 -390
rect 778 -396 781 -390
rect 785 -396 788 -390
rect 792 -396 795 -390
rect 799 -396 802 -390
rect 806 -396 809 -390
rect 813 -396 816 -390
rect 820 -396 823 -390
rect 827 -396 830 -390
rect 834 -396 837 -390
rect 841 -396 844 -390
rect 848 -396 851 -390
rect 855 -396 858 -390
rect 862 -396 865 -390
rect 869 -396 872 -390
rect 876 -396 882 -390
rect 883 -396 889 -390
rect 890 -396 893 -390
rect 897 -396 900 -390
rect 904 -396 907 -390
rect 932 -396 935 -390
rect 1107 -396 1110 -390
rect 1 -485 4 -479
rect 8 -485 14 -479
rect 15 -485 18 -479
rect 22 -485 25 -479
rect 29 -485 32 -479
rect 36 -485 39 -479
rect 43 -485 46 -479
rect 50 -485 53 -479
rect 57 -485 63 -479
rect 64 -485 70 -479
rect 71 -485 74 -479
rect 78 -485 81 -479
rect 85 -485 88 -479
rect 92 -485 95 -479
rect 99 -485 102 -479
rect 106 -485 109 -479
rect 113 -485 116 -479
rect 120 -485 126 -479
rect 127 -485 133 -479
rect 134 -485 137 -479
rect 141 -485 147 -479
rect 148 -485 151 -479
rect 155 -485 158 -479
rect 162 -485 165 -479
rect 169 -485 172 -479
rect 176 -485 182 -479
rect 183 -485 186 -479
rect 190 -485 193 -479
rect 197 -485 203 -479
rect 204 -485 210 -479
rect 211 -485 214 -479
rect 218 -485 221 -479
rect 225 -485 228 -479
rect 232 -485 235 -479
rect 239 -485 242 -479
rect 246 -485 249 -479
rect 253 -485 256 -479
rect 260 -485 263 -479
rect 267 -485 270 -479
rect 274 -485 277 -479
rect 281 -485 287 -479
rect 288 -485 291 -479
rect 295 -485 298 -479
rect 302 -485 305 -479
rect 309 -485 312 -479
rect 316 -485 319 -479
rect 323 -485 329 -479
rect 330 -485 333 -479
rect 337 -485 340 -479
rect 344 -485 350 -479
rect 351 -485 357 -479
rect 358 -485 361 -479
rect 365 -485 368 -479
rect 372 -485 375 -479
rect 379 -485 385 -479
rect 386 -485 389 -479
rect 393 -485 399 -479
rect 400 -485 403 -479
rect 407 -485 410 -479
rect 414 -485 420 -479
rect 421 -485 427 -479
rect 428 -485 431 -479
rect 435 -485 438 -479
rect 442 -485 445 -479
rect 449 -485 452 -479
rect 456 -485 462 -479
rect 463 -485 466 -479
rect 470 -485 476 -479
rect 477 -485 483 -479
rect 484 -485 487 -479
rect 491 -485 494 -479
rect 498 -485 504 -479
rect 505 -485 508 -479
rect 512 -485 515 -479
rect 519 -485 522 -479
rect 526 -485 529 -479
rect 533 -485 539 -479
rect 540 -485 543 -479
rect 547 -485 550 -479
rect 554 -485 560 -479
rect 561 -485 567 -479
rect 568 -485 574 -479
rect 575 -485 581 -479
rect 582 -485 585 -479
rect 589 -485 592 -479
rect 596 -485 599 -479
rect 603 -485 606 -479
rect 610 -485 613 -479
rect 617 -485 620 -479
rect 624 -485 627 -479
rect 631 -485 637 -479
rect 638 -485 644 -479
rect 645 -485 648 -479
rect 652 -485 655 -479
rect 659 -485 662 -479
rect 666 -485 669 -479
rect 673 -485 676 -479
rect 680 -485 683 -479
rect 687 -485 693 -479
rect 694 -485 697 -479
rect 701 -485 704 -479
rect 708 -485 711 -479
rect 715 -485 718 -479
rect 722 -485 725 -479
rect 729 -485 732 -479
rect 736 -485 739 -479
rect 743 -485 746 -479
rect 750 -485 753 -479
rect 757 -485 760 -479
rect 764 -485 767 -479
rect 771 -485 774 -479
rect 778 -485 781 -479
rect 785 -485 788 -479
rect 792 -485 795 -479
rect 799 -485 802 -479
rect 806 -485 809 -479
rect 813 -485 819 -479
rect 820 -485 823 -479
rect 827 -485 830 -479
rect 834 -485 837 -479
rect 841 -485 844 -479
rect 848 -485 851 -479
rect 855 -485 858 -479
rect 862 -485 865 -479
rect 869 -485 872 -479
rect 876 -485 879 -479
rect 883 -485 886 -479
rect 890 -485 893 -479
rect 897 -485 900 -479
rect 904 -485 907 -479
rect 911 -485 914 -479
rect 918 -485 921 -479
rect 925 -485 928 -479
rect 932 -485 935 -479
rect 939 -485 942 -479
rect 946 -485 949 -479
rect 953 -485 956 -479
rect 960 -485 963 -479
rect 967 -485 970 -479
rect 974 -485 977 -479
rect 981 -485 984 -479
rect 988 -485 991 -479
rect 995 -485 998 -479
rect 1002 -485 1005 -479
rect 1009 -485 1012 -479
rect 1016 -485 1019 -479
rect 1023 -485 1026 -479
rect 1030 -485 1036 -479
rect 1037 -485 1043 -479
rect 1044 -485 1047 -479
rect 1114 -485 1117 -479
rect 1 -602 7 -596
rect 8 -602 11 -596
rect 15 -602 18 -596
rect 22 -602 28 -596
rect 29 -602 32 -596
rect 36 -602 42 -596
rect 43 -602 46 -596
rect 50 -602 53 -596
rect 57 -602 60 -596
rect 64 -602 67 -596
rect 71 -602 74 -596
rect 78 -602 81 -596
rect 85 -602 88 -596
rect 92 -602 98 -596
rect 99 -602 105 -596
rect 106 -602 112 -596
rect 113 -602 116 -596
rect 120 -602 123 -596
rect 127 -602 130 -596
rect 134 -602 140 -596
rect 141 -602 144 -596
rect 148 -602 151 -596
rect 155 -602 158 -596
rect 162 -602 168 -596
rect 169 -602 172 -596
rect 176 -602 182 -596
rect 183 -602 186 -596
rect 190 -602 193 -596
rect 197 -602 200 -596
rect 204 -602 210 -596
rect 211 -602 217 -596
rect 218 -602 224 -596
rect 225 -602 228 -596
rect 232 -602 235 -596
rect 239 -602 242 -596
rect 246 -602 249 -596
rect 253 -602 256 -596
rect 260 -602 263 -596
rect 267 -602 273 -596
rect 274 -602 277 -596
rect 281 -602 284 -596
rect 288 -602 291 -596
rect 295 -602 298 -596
rect 302 -602 305 -596
rect 309 -602 312 -596
rect 316 -602 319 -596
rect 323 -602 326 -596
rect 330 -602 333 -596
rect 337 -602 343 -596
rect 344 -602 350 -596
rect 351 -602 354 -596
rect 358 -602 361 -596
rect 365 -602 368 -596
rect 372 -602 375 -596
rect 379 -602 382 -596
rect 386 -602 389 -596
rect 393 -602 396 -596
rect 400 -602 403 -596
rect 407 -602 410 -596
rect 414 -602 417 -596
rect 421 -602 424 -596
rect 428 -602 431 -596
rect 435 -602 441 -596
rect 442 -602 445 -596
rect 449 -602 452 -596
rect 456 -602 459 -596
rect 463 -602 469 -596
rect 470 -602 476 -596
rect 477 -602 480 -596
rect 484 -602 487 -596
rect 491 -602 494 -596
rect 498 -602 501 -596
rect 505 -602 508 -596
rect 512 -602 515 -596
rect 519 -602 525 -596
rect 526 -602 532 -596
rect 533 -602 539 -596
rect 540 -602 543 -596
rect 547 -602 553 -596
rect 554 -602 557 -596
rect 561 -602 567 -596
rect 568 -602 574 -596
rect 575 -602 581 -596
rect 582 -602 585 -596
rect 589 -602 592 -596
rect 596 -602 602 -596
rect 603 -602 606 -596
rect 610 -602 613 -596
rect 617 -602 620 -596
rect 624 -602 627 -596
rect 631 -602 637 -596
rect 638 -602 641 -596
rect 645 -602 648 -596
rect 652 -602 655 -596
rect 659 -602 662 -596
rect 666 -602 669 -596
rect 673 -602 676 -596
rect 680 -602 686 -596
rect 687 -602 690 -596
rect 694 -602 697 -596
rect 701 -602 704 -596
rect 708 -602 714 -596
rect 715 -602 718 -596
rect 722 -602 725 -596
rect 729 -602 735 -596
rect 736 -602 739 -596
rect 743 -602 746 -596
rect 750 -602 753 -596
rect 757 -602 760 -596
rect 764 -602 767 -596
rect 771 -602 774 -596
rect 778 -602 781 -596
rect 785 -602 788 -596
rect 792 -602 795 -596
rect 799 -602 802 -596
rect 806 -602 809 -596
rect 813 -602 816 -596
rect 820 -602 823 -596
rect 827 -602 830 -596
rect 834 -602 837 -596
rect 841 -602 844 -596
rect 848 -602 851 -596
rect 855 -602 858 -596
rect 862 -602 865 -596
rect 869 -602 872 -596
rect 876 -602 879 -596
rect 883 -602 886 -596
rect 890 -602 893 -596
rect 897 -602 900 -596
rect 904 -602 907 -596
rect 911 -602 914 -596
rect 918 -602 921 -596
rect 925 -602 928 -596
rect 932 -602 935 -596
rect 939 -602 942 -596
rect 946 -602 949 -596
rect 953 -602 956 -596
rect 960 -602 963 -596
rect 967 -602 970 -596
rect 974 -602 977 -596
rect 981 -602 984 -596
rect 988 -602 991 -596
rect 995 -602 998 -596
rect 1002 -602 1005 -596
rect 1009 -602 1012 -596
rect 1016 -602 1019 -596
rect 1023 -602 1026 -596
rect 1030 -602 1033 -596
rect 1037 -602 1040 -596
rect 1044 -602 1047 -596
rect 1051 -602 1054 -596
rect 1058 -602 1061 -596
rect 1065 -602 1068 -596
rect 1072 -602 1075 -596
rect 1079 -602 1082 -596
rect 1086 -602 1089 -596
rect 1093 -602 1096 -596
rect 1100 -602 1106 -596
rect 1107 -602 1113 -596
rect 1114 -602 1117 -596
rect 1121 -602 1124 -596
rect 1128 -602 1131 -596
rect 1 -703 4 -697
rect 8 -703 14 -697
rect 15 -703 18 -697
rect 22 -703 25 -697
rect 29 -703 32 -697
rect 36 -703 39 -697
rect 43 -703 49 -697
rect 50 -703 53 -697
rect 57 -703 60 -697
rect 64 -703 67 -697
rect 71 -703 74 -697
rect 78 -703 84 -697
rect 85 -703 88 -697
rect 92 -703 95 -697
rect 99 -703 102 -697
rect 106 -703 109 -697
rect 113 -703 119 -697
rect 120 -703 126 -697
rect 127 -703 133 -697
rect 134 -703 137 -697
rect 141 -703 144 -697
rect 148 -703 151 -697
rect 155 -703 158 -697
rect 162 -703 165 -697
rect 169 -703 175 -697
rect 176 -703 179 -697
rect 183 -703 186 -697
rect 190 -703 196 -697
rect 197 -703 203 -697
rect 204 -703 210 -697
rect 211 -703 214 -697
rect 218 -703 221 -697
rect 225 -703 231 -697
rect 232 -703 235 -697
rect 239 -703 242 -697
rect 246 -703 249 -697
rect 253 -703 256 -697
rect 260 -703 263 -697
rect 267 -703 270 -697
rect 274 -703 277 -697
rect 281 -703 284 -697
rect 288 -703 294 -697
rect 295 -703 298 -697
rect 302 -703 305 -697
rect 309 -703 315 -697
rect 316 -703 319 -697
rect 323 -703 326 -697
rect 330 -703 333 -697
rect 337 -703 340 -697
rect 344 -703 347 -697
rect 351 -703 354 -697
rect 358 -703 364 -697
rect 365 -703 368 -697
rect 372 -703 375 -697
rect 379 -703 382 -697
rect 386 -703 389 -697
rect 393 -703 396 -697
rect 400 -703 403 -697
rect 407 -703 410 -697
rect 414 -703 417 -697
rect 421 -703 424 -697
rect 428 -703 431 -697
rect 435 -703 438 -697
rect 442 -703 448 -697
rect 449 -703 455 -697
rect 456 -703 462 -697
rect 463 -703 469 -697
rect 470 -703 473 -697
rect 477 -703 483 -697
rect 484 -703 487 -697
rect 491 -703 497 -697
rect 498 -703 501 -697
rect 505 -703 508 -697
rect 512 -703 518 -697
rect 519 -703 522 -697
rect 526 -703 529 -697
rect 533 -703 536 -697
rect 540 -703 546 -697
rect 547 -703 550 -697
rect 554 -703 557 -697
rect 561 -703 567 -697
rect 568 -703 571 -697
rect 575 -703 578 -697
rect 582 -703 585 -697
rect 589 -703 592 -697
rect 596 -703 599 -697
rect 603 -703 609 -697
rect 610 -703 613 -697
rect 617 -703 620 -697
rect 624 -703 627 -697
rect 631 -703 634 -697
rect 638 -703 641 -697
rect 645 -703 648 -697
rect 652 -703 655 -697
rect 659 -703 662 -697
rect 666 -703 672 -697
rect 673 -703 676 -697
rect 680 -703 683 -697
rect 687 -703 690 -697
rect 694 -703 697 -697
rect 701 -703 704 -697
rect 708 -703 711 -697
rect 715 -703 718 -697
rect 722 -703 728 -697
rect 729 -703 732 -697
rect 736 -703 739 -697
rect 743 -703 749 -697
rect 750 -703 753 -697
rect 757 -703 760 -697
rect 764 -703 767 -697
rect 771 -703 777 -697
rect 778 -703 781 -697
rect 785 -703 791 -697
rect 792 -703 795 -697
rect 799 -703 802 -697
rect 806 -703 809 -697
rect 813 -703 816 -697
rect 820 -703 823 -697
rect 827 -703 830 -697
rect 834 -703 837 -697
rect 841 -703 844 -697
rect 848 -703 851 -697
rect 855 -703 858 -697
rect 862 -703 865 -697
rect 869 -703 872 -697
rect 876 -703 879 -697
rect 883 -703 886 -697
rect 890 -703 893 -697
rect 897 -703 900 -697
rect 904 -703 907 -697
rect 911 -703 914 -697
rect 918 -703 921 -697
rect 925 -703 928 -697
rect 932 -703 935 -697
rect 939 -703 942 -697
rect 946 -703 949 -697
rect 953 -703 956 -697
rect 960 -703 963 -697
rect 967 -703 970 -697
rect 974 -703 977 -697
rect 981 -703 984 -697
rect 988 -703 991 -697
rect 995 -703 998 -697
rect 1002 -703 1005 -697
rect 1009 -703 1012 -697
rect 1016 -703 1019 -697
rect 1023 -703 1026 -697
rect 1030 -703 1033 -697
rect 1037 -703 1040 -697
rect 1044 -703 1047 -697
rect 1051 -703 1054 -697
rect 1058 -703 1061 -697
rect 1065 -703 1068 -697
rect 1072 -703 1075 -697
rect 1079 -703 1085 -697
rect 1086 -703 1089 -697
rect 1093 -703 1096 -697
rect 1100 -703 1103 -697
rect 1107 -703 1113 -697
rect 1114 -703 1117 -697
rect 1121 -703 1124 -697
rect 1128 -703 1131 -697
rect 1135 -703 1141 -697
rect 1142 -703 1145 -697
rect 1149 -703 1152 -697
rect 1156 -703 1159 -697
rect 22 -780 25 -774
rect 29 -780 35 -774
rect 36 -780 39 -774
rect 43 -780 46 -774
rect 50 -780 53 -774
rect 57 -780 60 -774
rect 64 -780 67 -774
rect 71 -780 74 -774
rect 78 -780 81 -774
rect 85 -780 91 -774
rect 92 -780 95 -774
rect 99 -780 105 -774
rect 106 -780 109 -774
rect 113 -780 116 -774
rect 120 -780 123 -774
rect 127 -780 130 -774
rect 134 -780 140 -774
rect 141 -780 144 -774
rect 148 -780 154 -774
rect 155 -780 161 -774
rect 162 -780 165 -774
rect 169 -780 175 -774
rect 176 -780 179 -774
rect 183 -780 186 -774
rect 190 -780 193 -774
rect 197 -780 200 -774
rect 204 -780 210 -774
rect 211 -780 214 -774
rect 218 -780 221 -774
rect 225 -780 228 -774
rect 232 -780 235 -774
rect 239 -780 242 -774
rect 246 -780 249 -774
rect 253 -780 256 -774
rect 260 -780 263 -774
rect 267 -780 270 -774
rect 274 -780 277 -774
rect 281 -780 284 -774
rect 288 -780 294 -774
rect 295 -780 298 -774
rect 302 -780 305 -774
rect 309 -780 315 -774
rect 316 -780 319 -774
rect 323 -780 329 -774
rect 330 -780 333 -774
rect 337 -780 340 -774
rect 344 -780 347 -774
rect 351 -780 354 -774
rect 358 -780 361 -774
rect 365 -780 371 -774
rect 372 -780 375 -774
rect 379 -780 382 -774
rect 386 -780 389 -774
rect 393 -780 396 -774
rect 400 -780 403 -774
rect 407 -780 410 -774
rect 414 -780 417 -774
rect 421 -780 424 -774
rect 428 -780 431 -774
rect 435 -780 438 -774
rect 442 -780 448 -774
rect 449 -780 452 -774
rect 456 -780 462 -774
rect 463 -780 469 -774
rect 470 -780 473 -774
rect 477 -780 480 -774
rect 484 -780 487 -774
rect 491 -780 497 -774
rect 498 -780 501 -774
rect 505 -780 508 -774
rect 512 -780 515 -774
rect 519 -780 522 -774
rect 526 -780 532 -774
rect 533 -780 539 -774
rect 540 -780 543 -774
rect 547 -780 550 -774
rect 554 -780 557 -774
rect 561 -780 564 -774
rect 568 -780 571 -774
rect 575 -780 578 -774
rect 582 -780 585 -774
rect 589 -780 592 -774
rect 596 -780 599 -774
rect 603 -780 606 -774
rect 610 -780 613 -774
rect 617 -780 623 -774
rect 624 -780 627 -774
rect 631 -780 634 -774
rect 638 -780 641 -774
rect 645 -780 648 -774
rect 652 -780 658 -774
rect 659 -780 665 -774
rect 666 -780 669 -774
rect 673 -780 676 -774
rect 680 -780 683 -774
rect 687 -780 690 -774
rect 694 -780 697 -774
rect 701 -780 707 -774
rect 708 -780 711 -774
rect 715 -780 721 -774
rect 722 -780 725 -774
rect 729 -780 732 -774
rect 736 -780 739 -774
rect 743 -780 746 -774
rect 750 -780 753 -774
rect 757 -780 763 -774
rect 764 -780 767 -774
rect 771 -780 777 -774
rect 778 -780 781 -774
rect 785 -780 788 -774
rect 792 -780 798 -774
rect 799 -780 802 -774
rect 806 -780 809 -774
rect 813 -780 816 -774
rect 820 -780 823 -774
rect 827 -780 830 -774
rect 834 -780 837 -774
rect 841 -780 844 -774
rect 848 -780 851 -774
rect 855 -780 858 -774
rect 862 -780 865 -774
rect 869 -780 872 -774
rect 876 -780 882 -774
rect 883 -780 886 -774
rect 890 -780 893 -774
rect 897 -780 900 -774
rect 904 -780 907 -774
rect 911 -780 914 -774
rect 918 -780 921 -774
rect 925 -780 928 -774
rect 932 -780 938 -774
rect 939 -780 945 -774
rect 946 -780 952 -774
rect 953 -780 959 -774
rect 960 -780 963 -774
rect 967 -780 970 -774
rect 974 -780 977 -774
rect 981 -780 984 -774
rect 988 -780 991 -774
rect 995 -780 998 -774
rect 1002 -780 1005 -774
rect 1009 -780 1015 -774
rect 1030 -780 1033 -774
rect 1121 -780 1124 -774
rect 1 -867 4 -861
rect 8 -867 14 -861
rect 15 -867 18 -861
rect 22 -867 25 -861
rect 29 -867 32 -861
rect 36 -867 42 -861
rect 43 -867 46 -861
rect 50 -867 53 -861
rect 57 -867 60 -861
rect 64 -867 67 -861
rect 71 -867 77 -861
rect 78 -867 84 -861
rect 85 -867 88 -861
rect 92 -867 95 -861
rect 99 -867 102 -861
rect 106 -867 109 -861
rect 113 -867 116 -861
rect 120 -867 123 -861
rect 127 -867 130 -861
rect 134 -867 137 -861
rect 141 -867 144 -861
rect 148 -867 151 -861
rect 155 -867 158 -861
rect 162 -867 165 -861
rect 169 -867 172 -861
rect 176 -867 179 -861
rect 183 -867 186 -861
rect 190 -867 196 -861
rect 197 -867 200 -861
rect 204 -867 207 -861
rect 211 -867 214 -861
rect 218 -867 224 -861
rect 225 -867 231 -861
rect 232 -867 235 -861
rect 239 -867 242 -861
rect 246 -867 249 -861
rect 253 -867 256 -861
rect 260 -867 266 -861
rect 267 -867 270 -861
rect 274 -867 277 -861
rect 281 -867 284 -861
rect 288 -867 291 -861
rect 295 -867 298 -861
rect 302 -867 305 -861
rect 309 -867 312 -861
rect 316 -867 319 -861
rect 323 -867 329 -861
rect 330 -867 333 -861
rect 337 -867 343 -861
rect 344 -867 347 -861
rect 351 -867 357 -861
rect 358 -867 361 -861
rect 365 -867 368 -861
rect 372 -867 375 -861
rect 379 -867 385 -861
rect 386 -867 389 -861
rect 393 -867 399 -861
rect 400 -867 403 -861
rect 407 -867 410 -861
rect 414 -867 417 -861
rect 421 -867 424 -861
rect 428 -867 434 -861
rect 435 -867 438 -861
rect 442 -867 445 -861
rect 449 -867 455 -861
rect 456 -867 459 -861
rect 463 -867 466 -861
rect 470 -867 473 -861
rect 477 -867 483 -861
rect 484 -867 487 -861
rect 491 -867 494 -861
rect 498 -867 504 -861
rect 505 -867 508 -861
rect 512 -867 515 -861
rect 519 -867 522 -861
rect 526 -867 529 -861
rect 533 -867 536 -861
rect 540 -867 546 -861
rect 547 -867 550 -861
rect 554 -867 560 -861
rect 561 -867 567 -861
rect 568 -867 571 -861
rect 575 -867 581 -861
rect 582 -867 585 -861
rect 589 -867 595 -861
rect 596 -867 599 -861
rect 603 -867 609 -861
rect 610 -867 616 -861
rect 617 -867 620 -861
rect 624 -867 627 -861
rect 631 -867 637 -861
rect 638 -867 641 -861
rect 645 -867 648 -861
rect 652 -867 658 -861
rect 659 -867 662 -861
rect 666 -867 669 -861
rect 673 -867 676 -861
rect 680 -867 683 -861
rect 687 -867 690 -861
rect 694 -867 697 -861
rect 701 -867 704 -861
rect 708 -867 711 -861
rect 715 -867 718 -861
rect 722 -867 725 -861
rect 729 -867 732 -861
rect 736 -867 739 -861
rect 743 -867 746 -861
rect 750 -867 753 -861
rect 757 -867 760 -861
rect 764 -867 770 -861
rect 771 -867 774 -861
rect 778 -867 781 -861
rect 785 -867 788 -861
rect 792 -867 795 -861
rect 799 -867 802 -861
rect 806 -867 809 -861
rect 813 -867 816 -861
rect 820 -867 823 -861
rect 827 -867 830 -861
rect 834 -867 837 -861
rect 841 -867 844 -861
rect 848 -867 851 -861
rect 855 -867 858 -861
rect 862 -867 868 -861
rect 869 -867 872 -861
rect 876 -867 879 -861
rect 883 -867 886 -861
rect 890 -867 893 -861
rect 897 -867 900 -861
rect 904 -867 907 -861
rect 911 -867 914 -861
rect 918 -867 921 -861
rect 925 -867 928 -861
rect 932 -867 935 -861
rect 939 -867 942 -861
rect 946 -867 949 -861
rect 953 -867 956 -861
rect 960 -867 963 -861
rect 967 -867 970 -861
rect 974 -867 977 -861
rect 981 -867 984 -861
rect 988 -867 991 -861
rect 995 -867 998 -861
rect 1002 -867 1005 -861
rect 1009 -867 1012 -861
rect 1016 -867 1019 -861
rect 1023 -867 1026 -861
rect 1030 -867 1033 -861
rect 1037 -867 1040 -861
rect 1044 -867 1047 -861
rect 1051 -867 1054 -861
rect 1058 -867 1061 -861
rect 1065 -867 1068 -861
rect 1072 -867 1075 -861
rect 1079 -867 1082 -861
rect 1086 -867 1089 -861
rect 1093 -867 1099 -861
rect 1100 -867 1103 -861
rect 1107 -867 1110 -861
rect 1114 -867 1117 -861
rect 1121 -867 1124 -861
rect 1128 -867 1134 -861
rect 1135 -867 1141 -861
rect 1142 -867 1145 -861
rect 1149 -867 1155 -861
rect 1 -968 7 -962
rect 8 -968 11 -962
rect 15 -968 21 -962
rect 22 -968 25 -962
rect 29 -968 35 -962
rect 36 -968 42 -962
rect 43 -968 46 -962
rect 50 -968 53 -962
rect 57 -968 60 -962
rect 64 -968 70 -962
rect 71 -968 77 -962
rect 78 -968 84 -962
rect 85 -968 88 -962
rect 92 -968 95 -962
rect 99 -968 102 -962
rect 106 -968 109 -962
rect 113 -968 116 -962
rect 120 -968 123 -962
rect 127 -968 130 -962
rect 134 -968 137 -962
rect 141 -968 144 -962
rect 148 -968 154 -962
rect 155 -968 158 -962
rect 162 -968 165 -962
rect 169 -968 172 -962
rect 176 -968 179 -962
rect 183 -968 186 -962
rect 190 -968 193 -962
rect 197 -968 200 -962
rect 204 -968 207 -962
rect 211 -968 214 -962
rect 218 -968 221 -962
rect 225 -968 228 -962
rect 232 -968 235 -962
rect 239 -968 242 -962
rect 246 -968 249 -962
rect 253 -968 256 -962
rect 260 -968 263 -962
rect 267 -968 270 -962
rect 274 -968 277 -962
rect 281 -968 287 -962
rect 288 -968 291 -962
rect 295 -968 301 -962
rect 302 -968 308 -962
rect 309 -968 312 -962
rect 316 -968 319 -962
rect 323 -968 326 -962
rect 330 -968 333 -962
rect 337 -968 340 -962
rect 344 -968 347 -962
rect 351 -968 354 -962
rect 358 -968 364 -962
rect 365 -968 368 -962
rect 372 -968 375 -962
rect 379 -968 382 -962
rect 386 -968 389 -962
rect 393 -968 396 -962
rect 400 -968 403 -962
rect 407 -968 410 -962
rect 414 -968 420 -962
rect 421 -968 424 -962
rect 428 -968 431 -962
rect 435 -968 441 -962
rect 442 -968 448 -962
rect 449 -968 452 -962
rect 456 -968 459 -962
rect 463 -968 469 -962
rect 470 -968 476 -962
rect 477 -968 483 -962
rect 484 -968 487 -962
rect 491 -968 494 -962
rect 498 -968 504 -962
rect 505 -968 511 -962
rect 512 -968 515 -962
rect 519 -968 522 -962
rect 526 -968 529 -962
rect 533 -968 539 -962
rect 540 -968 546 -962
rect 547 -968 550 -962
rect 554 -968 557 -962
rect 561 -968 564 -962
rect 568 -968 574 -962
rect 575 -968 581 -962
rect 582 -968 585 -962
rect 589 -968 595 -962
rect 596 -968 599 -962
rect 603 -968 606 -962
rect 610 -968 616 -962
rect 617 -968 623 -962
rect 624 -968 630 -962
rect 631 -968 637 -962
rect 638 -968 641 -962
rect 645 -968 648 -962
rect 652 -968 655 -962
rect 659 -968 662 -962
rect 666 -968 669 -962
rect 673 -968 676 -962
rect 680 -968 683 -962
rect 687 -968 693 -962
rect 694 -968 700 -962
rect 701 -968 704 -962
rect 708 -968 711 -962
rect 715 -968 718 -962
rect 722 -968 725 -962
rect 729 -968 732 -962
rect 736 -968 739 -962
rect 743 -968 746 -962
rect 750 -968 753 -962
rect 757 -968 760 -962
rect 764 -968 767 -962
rect 771 -968 774 -962
rect 778 -968 781 -962
rect 785 -968 788 -962
rect 792 -968 795 -962
rect 799 -968 802 -962
rect 806 -968 809 -962
rect 813 -968 816 -962
rect 820 -968 823 -962
rect 827 -968 830 -962
rect 834 -968 837 -962
rect 841 -968 844 -962
rect 848 -968 851 -962
rect 855 -968 861 -962
rect 862 -968 865 -962
rect 869 -968 872 -962
rect 876 -968 879 -962
rect 883 -968 886 -962
rect 890 -968 893 -962
rect 897 -968 900 -962
rect 904 -968 907 -962
rect 911 -968 914 -962
rect 918 -968 921 -962
rect 925 -968 928 -962
rect 932 -968 935 -962
rect 939 -968 942 -962
rect 946 -968 949 -962
rect 953 -968 956 -962
rect 960 -968 963 -962
rect 967 -968 970 -962
rect 974 -968 977 -962
rect 981 -968 984 -962
rect 988 -968 991 -962
rect 995 -968 998 -962
rect 1002 -968 1005 -962
rect 1009 -968 1012 -962
rect 1016 -968 1019 -962
rect 1023 -968 1026 -962
rect 1030 -968 1033 -962
rect 1037 -968 1040 -962
rect 1044 -968 1047 -962
rect 1051 -968 1054 -962
rect 1058 -968 1061 -962
rect 1065 -968 1068 -962
rect 1072 -968 1075 -962
rect 1079 -968 1082 -962
rect 1086 -968 1089 -962
rect 1093 -968 1096 -962
rect 1100 -968 1103 -962
rect 1107 -968 1110 -962
rect 1114 -968 1117 -962
rect 1121 -968 1124 -962
rect 1128 -968 1131 -962
rect 1135 -968 1138 -962
rect 1142 -968 1145 -962
rect 1149 -968 1152 -962
rect 1156 -968 1159 -962
rect 1 -1083 7 -1077
rect 8 -1083 11 -1077
rect 15 -1083 18 -1077
rect 22 -1083 25 -1077
rect 29 -1083 32 -1077
rect 36 -1083 39 -1077
rect 43 -1083 46 -1077
rect 50 -1083 56 -1077
rect 57 -1083 60 -1077
rect 64 -1083 70 -1077
rect 71 -1083 74 -1077
rect 78 -1083 84 -1077
rect 85 -1083 88 -1077
rect 92 -1083 95 -1077
rect 99 -1083 105 -1077
rect 106 -1083 112 -1077
rect 113 -1083 116 -1077
rect 120 -1083 123 -1077
rect 127 -1083 130 -1077
rect 134 -1083 137 -1077
rect 141 -1083 144 -1077
rect 148 -1083 151 -1077
rect 155 -1083 158 -1077
rect 162 -1083 168 -1077
rect 169 -1083 172 -1077
rect 176 -1083 179 -1077
rect 183 -1083 186 -1077
rect 190 -1083 196 -1077
rect 197 -1083 203 -1077
rect 204 -1083 207 -1077
rect 211 -1083 217 -1077
rect 218 -1083 221 -1077
rect 225 -1083 231 -1077
rect 232 -1083 235 -1077
rect 239 -1083 242 -1077
rect 246 -1083 249 -1077
rect 253 -1083 256 -1077
rect 260 -1083 263 -1077
rect 267 -1083 273 -1077
rect 274 -1083 277 -1077
rect 281 -1083 287 -1077
rect 288 -1083 291 -1077
rect 295 -1083 298 -1077
rect 302 -1083 305 -1077
rect 309 -1083 312 -1077
rect 316 -1083 319 -1077
rect 323 -1083 329 -1077
rect 330 -1083 333 -1077
rect 337 -1083 340 -1077
rect 344 -1083 347 -1077
rect 351 -1083 354 -1077
rect 358 -1083 361 -1077
rect 365 -1083 368 -1077
rect 372 -1083 375 -1077
rect 379 -1083 382 -1077
rect 386 -1083 392 -1077
rect 393 -1083 399 -1077
rect 400 -1083 403 -1077
rect 407 -1083 410 -1077
rect 414 -1083 417 -1077
rect 421 -1083 424 -1077
rect 428 -1083 431 -1077
rect 435 -1083 438 -1077
rect 442 -1083 445 -1077
rect 449 -1083 452 -1077
rect 456 -1083 459 -1077
rect 463 -1083 466 -1077
rect 470 -1083 473 -1077
rect 477 -1083 480 -1077
rect 484 -1083 490 -1077
rect 491 -1083 497 -1077
rect 498 -1083 504 -1077
rect 505 -1083 508 -1077
rect 512 -1083 515 -1077
rect 519 -1083 522 -1077
rect 526 -1083 529 -1077
rect 533 -1083 536 -1077
rect 540 -1083 546 -1077
rect 547 -1083 550 -1077
rect 554 -1083 560 -1077
rect 561 -1083 564 -1077
rect 568 -1083 574 -1077
rect 575 -1083 578 -1077
rect 582 -1083 588 -1077
rect 589 -1083 592 -1077
rect 596 -1083 602 -1077
rect 603 -1083 609 -1077
rect 610 -1083 613 -1077
rect 617 -1083 620 -1077
rect 624 -1083 627 -1077
rect 631 -1083 637 -1077
rect 638 -1083 641 -1077
rect 645 -1083 648 -1077
rect 652 -1083 655 -1077
rect 659 -1083 662 -1077
rect 666 -1083 669 -1077
rect 673 -1083 676 -1077
rect 680 -1083 686 -1077
rect 687 -1083 690 -1077
rect 694 -1083 697 -1077
rect 701 -1083 704 -1077
rect 708 -1083 711 -1077
rect 715 -1083 718 -1077
rect 722 -1083 728 -1077
rect 729 -1083 732 -1077
rect 736 -1083 742 -1077
rect 743 -1083 746 -1077
rect 750 -1083 753 -1077
rect 757 -1083 760 -1077
rect 764 -1083 767 -1077
rect 771 -1083 774 -1077
rect 778 -1083 781 -1077
rect 785 -1083 788 -1077
rect 792 -1083 795 -1077
rect 799 -1083 802 -1077
rect 806 -1083 809 -1077
rect 813 -1083 819 -1077
rect 820 -1083 823 -1077
rect 827 -1083 830 -1077
rect 834 -1083 837 -1077
rect 841 -1083 844 -1077
rect 848 -1083 851 -1077
rect 855 -1083 858 -1077
rect 862 -1083 865 -1077
rect 869 -1083 872 -1077
rect 876 -1083 879 -1077
rect 883 -1083 886 -1077
rect 890 -1083 893 -1077
rect 897 -1083 900 -1077
rect 904 -1083 907 -1077
rect 911 -1083 914 -1077
rect 918 -1083 921 -1077
rect 925 -1083 928 -1077
rect 932 -1083 935 -1077
rect 939 -1083 942 -1077
rect 946 -1083 949 -1077
rect 953 -1083 956 -1077
rect 960 -1083 963 -1077
rect 967 -1083 970 -1077
rect 974 -1083 977 -1077
rect 981 -1083 984 -1077
rect 988 -1083 991 -1077
rect 995 -1083 998 -1077
rect 1002 -1083 1005 -1077
rect 1009 -1083 1012 -1077
rect 1016 -1083 1019 -1077
rect 1023 -1083 1026 -1077
rect 1030 -1083 1033 -1077
rect 1037 -1083 1043 -1077
rect 1044 -1083 1047 -1077
rect 1051 -1083 1054 -1077
rect 1058 -1083 1064 -1077
rect 1065 -1083 1068 -1077
rect 1072 -1083 1075 -1077
rect 1079 -1083 1082 -1077
rect 1128 -1083 1131 -1077
rect 1142 -1083 1145 -1077
rect 1 -1172 7 -1166
rect 8 -1172 11 -1166
rect 15 -1172 21 -1166
rect 22 -1172 25 -1166
rect 29 -1172 32 -1166
rect 36 -1172 42 -1166
rect 43 -1172 46 -1166
rect 50 -1172 53 -1166
rect 57 -1172 63 -1166
rect 64 -1172 67 -1166
rect 71 -1172 74 -1166
rect 78 -1172 81 -1166
rect 85 -1172 88 -1166
rect 92 -1172 95 -1166
rect 99 -1172 105 -1166
rect 106 -1172 109 -1166
rect 113 -1172 116 -1166
rect 120 -1172 123 -1166
rect 127 -1172 130 -1166
rect 134 -1172 137 -1166
rect 141 -1172 147 -1166
rect 148 -1172 154 -1166
rect 155 -1172 158 -1166
rect 162 -1172 168 -1166
rect 169 -1172 175 -1166
rect 176 -1172 179 -1166
rect 183 -1172 186 -1166
rect 190 -1172 193 -1166
rect 197 -1172 200 -1166
rect 204 -1172 207 -1166
rect 211 -1172 214 -1166
rect 218 -1172 224 -1166
rect 225 -1172 228 -1166
rect 232 -1172 235 -1166
rect 239 -1172 242 -1166
rect 246 -1172 249 -1166
rect 253 -1172 256 -1166
rect 260 -1172 263 -1166
rect 267 -1172 270 -1166
rect 274 -1172 277 -1166
rect 281 -1172 287 -1166
rect 288 -1172 291 -1166
rect 295 -1172 298 -1166
rect 302 -1172 305 -1166
rect 309 -1172 315 -1166
rect 316 -1172 319 -1166
rect 323 -1172 326 -1166
rect 330 -1172 333 -1166
rect 337 -1172 340 -1166
rect 344 -1172 350 -1166
rect 351 -1172 357 -1166
rect 358 -1172 364 -1166
rect 365 -1172 368 -1166
rect 372 -1172 375 -1166
rect 379 -1172 385 -1166
rect 386 -1172 389 -1166
rect 393 -1172 396 -1166
rect 400 -1172 403 -1166
rect 407 -1172 413 -1166
rect 414 -1172 420 -1166
rect 421 -1172 424 -1166
rect 428 -1172 431 -1166
rect 435 -1172 438 -1166
rect 442 -1172 445 -1166
rect 449 -1172 452 -1166
rect 456 -1172 459 -1166
rect 463 -1172 469 -1166
rect 470 -1172 473 -1166
rect 477 -1172 483 -1166
rect 484 -1172 487 -1166
rect 491 -1172 494 -1166
rect 498 -1172 504 -1166
rect 505 -1172 508 -1166
rect 512 -1172 515 -1166
rect 519 -1172 525 -1166
rect 526 -1172 529 -1166
rect 533 -1172 536 -1166
rect 540 -1172 543 -1166
rect 547 -1172 550 -1166
rect 554 -1172 560 -1166
rect 561 -1172 567 -1166
rect 568 -1172 571 -1166
rect 575 -1172 578 -1166
rect 582 -1172 585 -1166
rect 589 -1172 592 -1166
rect 596 -1172 602 -1166
rect 603 -1172 606 -1166
rect 610 -1172 613 -1166
rect 617 -1172 620 -1166
rect 624 -1172 627 -1166
rect 631 -1172 634 -1166
rect 638 -1172 641 -1166
rect 645 -1172 648 -1166
rect 652 -1172 655 -1166
rect 659 -1172 662 -1166
rect 666 -1172 669 -1166
rect 673 -1172 676 -1166
rect 680 -1172 683 -1166
rect 687 -1172 693 -1166
rect 694 -1172 697 -1166
rect 701 -1172 704 -1166
rect 708 -1172 711 -1166
rect 715 -1172 718 -1166
rect 722 -1172 725 -1166
rect 729 -1172 735 -1166
rect 736 -1172 742 -1166
rect 743 -1172 746 -1166
rect 750 -1172 753 -1166
rect 757 -1172 760 -1166
rect 764 -1172 767 -1166
rect 771 -1172 774 -1166
rect 778 -1172 781 -1166
rect 785 -1172 791 -1166
rect 792 -1172 795 -1166
rect 799 -1172 802 -1166
rect 806 -1172 809 -1166
rect 813 -1172 816 -1166
rect 820 -1172 823 -1166
rect 827 -1172 830 -1166
rect 834 -1172 837 -1166
rect 841 -1172 844 -1166
rect 848 -1172 851 -1166
rect 855 -1172 861 -1166
rect 862 -1172 865 -1166
rect 869 -1172 872 -1166
rect 876 -1172 879 -1166
rect 883 -1172 886 -1166
rect 890 -1172 893 -1166
rect 897 -1172 900 -1166
rect 904 -1172 907 -1166
rect 911 -1172 914 -1166
rect 918 -1172 921 -1166
rect 925 -1172 928 -1166
rect 932 -1172 935 -1166
rect 939 -1172 942 -1166
rect 946 -1172 949 -1166
rect 953 -1172 956 -1166
rect 960 -1172 963 -1166
rect 967 -1172 970 -1166
rect 974 -1172 977 -1166
rect 981 -1172 984 -1166
rect 988 -1172 991 -1166
rect 995 -1172 998 -1166
rect 1002 -1172 1005 -1166
rect 1009 -1172 1012 -1166
rect 1016 -1172 1019 -1166
rect 1023 -1172 1026 -1166
rect 1030 -1172 1033 -1166
rect 1037 -1172 1043 -1166
rect 1044 -1172 1047 -1166
rect 1051 -1172 1054 -1166
rect 1058 -1172 1061 -1166
rect 1065 -1172 1068 -1166
rect 1072 -1172 1078 -1166
rect 1121 -1172 1124 -1166
rect 1149 -1172 1152 -1166
rect 1 -1255 4 -1249
rect 8 -1255 11 -1249
rect 15 -1255 18 -1249
rect 22 -1255 28 -1249
rect 29 -1255 32 -1249
rect 36 -1255 39 -1249
rect 43 -1255 49 -1249
rect 50 -1255 53 -1249
rect 57 -1255 60 -1249
rect 64 -1255 67 -1249
rect 71 -1255 77 -1249
rect 78 -1255 81 -1249
rect 85 -1255 88 -1249
rect 92 -1255 98 -1249
rect 99 -1255 102 -1249
rect 106 -1255 109 -1249
rect 113 -1255 116 -1249
rect 120 -1255 123 -1249
rect 127 -1255 130 -1249
rect 134 -1255 137 -1249
rect 141 -1255 144 -1249
rect 148 -1255 151 -1249
rect 155 -1255 161 -1249
rect 162 -1255 165 -1249
rect 169 -1255 172 -1249
rect 176 -1255 179 -1249
rect 183 -1255 189 -1249
rect 190 -1255 196 -1249
rect 197 -1255 203 -1249
rect 204 -1255 207 -1249
rect 211 -1255 214 -1249
rect 218 -1255 221 -1249
rect 225 -1255 228 -1249
rect 232 -1255 235 -1249
rect 239 -1255 242 -1249
rect 246 -1255 249 -1249
rect 253 -1255 256 -1249
rect 260 -1255 263 -1249
rect 267 -1255 273 -1249
rect 274 -1255 277 -1249
rect 281 -1255 284 -1249
rect 288 -1255 294 -1249
rect 295 -1255 298 -1249
rect 302 -1255 308 -1249
rect 309 -1255 312 -1249
rect 316 -1255 319 -1249
rect 323 -1255 326 -1249
rect 330 -1255 333 -1249
rect 337 -1255 340 -1249
rect 344 -1255 347 -1249
rect 351 -1255 354 -1249
rect 358 -1255 364 -1249
rect 365 -1255 371 -1249
rect 372 -1255 378 -1249
rect 379 -1255 382 -1249
rect 386 -1255 389 -1249
rect 393 -1255 396 -1249
rect 400 -1255 403 -1249
rect 407 -1255 410 -1249
rect 414 -1255 417 -1249
rect 421 -1255 424 -1249
rect 428 -1255 431 -1249
rect 435 -1255 441 -1249
rect 442 -1255 445 -1249
rect 449 -1255 452 -1249
rect 456 -1255 462 -1249
rect 463 -1255 466 -1249
rect 470 -1255 473 -1249
rect 477 -1255 480 -1249
rect 484 -1255 487 -1249
rect 491 -1255 497 -1249
rect 498 -1255 501 -1249
rect 505 -1255 511 -1249
rect 512 -1255 515 -1249
rect 519 -1255 522 -1249
rect 526 -1255 529 -1249
rect 533 -1255 539 -1249
rect 540 -1255 543 -1249
rect 547 -1255 550 -1249
rect 554 -1255 557 -1249
rect 561 -1255 564 -1249
rect 568 -1255 571 -1249
rect 575 -1255 578 -1249
rect 582 -1255 585 -1249
rect 589 -1255 592 -1249
rect 596 -1255 602 -1249
rect 603 -1255 606 -1249
rect 610 -1255 613 -1249
rect 617 -1255 620 -1249
rect 624 -1255 627 -1249
rect 631 -1255 637 -1249
rect 638 -1255 644 -1249
rect 645 -1255 648 -1249
rect 652 -1255 658 -1249
rect 659 -1255 662 -1249
rect 666 -1255 672 -1249
rect 673 -1255 676 -1249
rect 680 -1255 686 -1249
rect 687 -1255 690 -1249
rect 694 -1255 697 -1249
rect 701 -1255 707 -1249
rect 708 -1255 711 -1249
rect 715 -1255 721 -1249
rect 722 -1255 725 -1249
rect 729 -1255 732 -1249
rect 736 -1255 739 -1249
rect 743 -1255 746 -1249
rect 750 -1255 753 -1249
rect 757 -1255 760 -1249
rect 764 -1255 767 -1249
rect 771 -1255 774 -1249
rect 778 -1255 781 -1249
rect 785 -1255 791 -1249
rect 792 -1255 795 -1249
rect 799 -1255 802 -1249
rect 806 -1255 809 -1249
rect 813 -1255 816 -1249
rect 820 -1255 823 -1249
rect 827 -1255 833 -1249
rect 834 -1255 837 -1249
rect 841 -1255 844 -1249
rect 848 -1255 851 -1249
rect 855 -1255 858 -1249
rect 862 -1255 865 -1249
rect 869 -1255 872 -1249
rect 876 -1255 879 -1249
rect 883 -1255 886 -1249
rect 890 -1255 893 -1249
rect 897 -1255 900 -1249
rect 904 -1255 907 -1249
rect 911 -1255 914 -1249
rect 918 -1255 921 -1249
rect 925 -1255 928 -1249
rect 932 -1255 935 -1249
rect 939 -1255 942 -1249
rect 946 -1255 949 -1249
rect 953 -1255 956 -1249
rect 960 -1255 963 -1249
rect 967 -1255 973 -1249
rect 974 -1255 977 -1249
rect 981 -1255 984 -1249
rect 988 -1255 991 -1249
rect 995 -1255 998 -1249
rect 1002 -1255 1005 -1249
rect 1009 -1255 1012 -1249
rect 1016 -1255 1019 -1249
rect 1023 -1255 1026 -1249
rect 1030 -1255 1033 -1249
rect 1037 -1255 1040 -1249
rect 1044 -1255 1047 -1249
rect 1051 -1255 1054 -1249
rect 1058 -1255 1061 -1249
rect 1065 -1255 1068 -1249
rect 1072 -1255 1075 -1249
rect 1079 -1255 1082 -1249
rect 1086 -1255 1089 -1249
rect 1093 -1255 1096 -1249
rect 1100 -1255 1103 -1249
rect 1107 -1255 1110 -1249
rect 1114 -1255 1120 -1249
rect 1121 -1255 1124 -1249
rect 1128 -1255 1134 -1249
rect 1135 -1255 1138 -1249
rect 1142 -1255 1145 -1249
rect 1149 -1255 1152 -1249
rect 1156 -1255 1159 -1249
rect 1163 -1255 1166 -1249
rect 1 -1348 4 -1342
rect 8 -1348 11 -1342
rect 15 -1348 18 -1342
rect 22 -1348 28 -1342
rect 29 -1348 35 -1342
rect 36 -1348 39 -1342
rect 43 -1348 46 -1342
rect 50 -1348 53 -1342
rect 57 -1348 60 -1342
rect 64 -1348 70 -1342
rect 71 -1348 74 -1342
rect 78 -1348 81 -1342
rect 85 -1348 88 -1342
rect 92 -1348 98 -1342
rect 99 -1348 105 -1342
rect 106 -1348 109 -1342
rect 113 -1348 116 -1342
rect 120 -1348 123 -1342
rect 127 -1348 130 -1342
rect 134 -1348 137 -1342
rect 141 -1348 144 -1342
rect 148 -1348 151 -1342
rect 155 -1348 158 -1342
rect 162 -1348 168 -1342
rect 169 -1348 172 -1342
rect 176 -1348 182 -1342
rect 183 -1348 186 -1342
rect 190 -1348 193 -1342
rect 197 -1348 200 -1342
rect 204 -1348 207 -1342
rect 211 -1348 217 -1342
rect 218 -1348 221 -1342
rect 225 -1348 228 -1342
rect 232 -1348 235 -1342
rect 239 -1348 242 -1342
rect 246 -1348 249 -1342
rect 253 -1348 256 -1342
rect 260 -1348 263 -1342
rect 267 -1348 270 -1342
rect 274 -1348 277 -1342
rect 281 -1348 284 -1342
rect 288 -1348 294 -1342
rect 295 -1348 298 -1342
rect 302 -1348 305 -1342
rect 309 -1348 312 -1342
rect 316 -1348 319 -1342
rect 323 -1348 326 -1342
rect 330 -1348 333 -1342
rect 337 -1348 340 -1342
rect 344 -1348 350 -1342
rect 351 -1348 354 -1342
rect 358 -1348 361 -1342
rect 365 -1348 368 -1342
rect 372 -1348 375 -1342
rect 379 -1348 382 -1342
rect 386 -1348 389 -1342
rect 393 -1348 396 -1342
rect 400 -1348 406 -1342
rect 407 -1348 413 -1342
rect 414 -1348 417 -1342
rect 421 -1348 424 -1342
rect 428 -1348 431 -1342
rect 435 -1348 441 -1342
rect 442 -1348 445 -1342
rect 449 -1348 452 -1342
rect 456 -1348 462 -1342
rect 463 -1348 466 -1342
rect 470 -1348 473 -1342
rect 477 -1348 480 -1342
rect 484 -1348 487 -1342
rect 491 -1348 497 -1342
rect 498 -1348 501 -1342
rect 505 -1348 508 -1342
rect 512 -1348 515 -1342
rect 519 -1348 525 -1342
rect 526 -1348 529 -1342
rect 533 -1348 539 -1342
rect 540 -1348 546 -1342
rect 547 -1348 550 -1342
rect 554 -1348 557 -1342
rect 561 -1348 564 -1342
rect 568 -1348 574 -1342
rect 575 -1348 578 -1342
rect 582 -1348 585 -1342
rect 589 -1348 592 -1342
rect 596 -1348 599 -1342
rect 603 -1348 609 -1342
rect 610 -1348 616 -1342
rect 617 -1348 623 -1342
rect 624 -1348 630 -1342
rect 631 -1348 634 -1342
rect 638 -1348 641 -1342
rect 645 -1348 648 -1342
rect 652 -1348 655 -1342
rect 659 -1348 662 -1342
rect 666 -1348 669 -1342
rect 673 -1348 676 -1342
rect 680 -1348 686 -1342
rect 687 -1348 690 -1342
rect 694 -1348 697 -1342
rect 701 -1348 704 -1342
rect 708 -1348 711 -1342
rect 715 -1348 718 -1342
rect 722 -1348 725 -1342
rect 729 -1348 735 -1342
rect 736 -1348 739 -1342
rect 743 -1348 746 -1342
rect 750 -1348 753 -1342
rect 757 -1348 760 -1342
rect 764 -1348 767 -1342
rect 771 -1348 777 -1342
rect 778 -1348 781 -1342
rect 785 -1348 788 -1342
rect 792 -1348 798 -1342
rect 799 -1348 802 -1342
rect 806 -1348 809 -1342
rect 813 -1348 816 -1342
rect 820 -1348 823 -1342
rect 827 -1348 833 -1342
rect 834 -1348 837 -1342
rect 841 -1348 844 -1342
rect 848 -1348 851 -1342
rect 855 -1348 858 -1342
rect 862 -1348 865 -1342
rect 869 -1348 872 -1342
rect 876 -1348 879 -1342
rect 883 -1348 886 -1342
rect 890 -1348 893 -1342
rect 897 -1348 900 -1342
rect 904 -1348 907 -1342
rect 911 -1348 914 -1342
rect 918 -1348 921 -1342
rect 925 -1348 928 -1342
rect 932 -1348 935 -1342
rect 939 -1348 942 -1342
rect 946 -1348 952 -1342
rect 953 -1348 956 -1342
rect 960 -1348 963 -1342
rect 967 -1348 970 -1342
rect 974 -1348 977 -1342
rect 981 -1348 984 -1342
rect 988 -1348 991 -1342
rect 995 -1348 1001 -1342
rect 1002 -1348 1005 -1342
rect 1009 -1348 1012 -1342
rect 1016 -1348 1019 -1342
rect 1023 -1348 1026 -1342
rect 1030 -1348 1033 -1342
rect 1037 -1348 1040 -1342
rect 1044 -1348 1047 -1342
rect 1051 -1348 1054 -1342
rect 1058 -1348 1061 -1342
rect 1065 -1348 1068 -1342
rect 1072 -1348 1075 -1342
rect 1079 -1348 1082 -1342
rect 1086 -1348 1089 -1342
rect 1093 -1348 1096 -1342
rect 1100 -1348 1103 -1342
rect 1107 -1348 1110 -1342
rect 1114 -1348 1117 -1342
rect 1121 -1348 1124 -1342
rect 1128 -1348 1131 -1342
rect 1135 -1348 1141 -1342
rect 1142 -1348 1145 -1342
rect 1149 -1348 1155 -1342
rect 1156 -1348 1159 -1342
rect 1163 -1348 1166 -1342
rect 1170 -1348 1173 -1342
rect 1 -1455 4 -1449
rect 8 -1455 14 -1449
rect 15 -1455 18 -1449
rect 22 -1455 25 -1449
rect 29 -1455 32 -1449
rect 36 -1455 39 -1449
rect 43 -1455 46 -1449
rect 50 -1455 53 -1449
rect 57 -1455 60 -1449
rect 64 -1455 67 -1449
rect 71 -1455 74 -1449
rect 78 -1455 81 -1449
rect 85 -1455 88 -1449
rect 92 -1455 95 -1449
rect 99 -1455 105 -1449
rect 106 -1455 112 -1449
rect 113 -1455 119 -1449
rect 120 -1455 126 -1449
rect 127 -1455 130 -1449
rect 134 -1455 137 -1449
rect 141 -1455 144 -1449
rect 148 -1455 151 -1449
rect 155 -1455 158 -1449
rect 162 -1455 165 -1449
rect 169 -1455 172 -1449
rect 176 -1455 182 -1449
rect 183 -1455 189 -1449
rect 190 -1455 196 -1449
rect 197 -1455 200 -1449
rect 204 -1455 207 -1449
rect 211 -1455 217 -1449
rect 218 -1455 221 -1449
rect 225 -1455 228 -1449
rect 232 -1455 235 -1449
rect 239 -1455 242 -1449
rect 246 -1455 249 -1449
rect 253 -1455 259 -1449
rect 260 -1455 263 -1449
rect 267 -1455 270 -1449
rect 274 -1455 277 -1449
rect 281 -1455 284 -1449
rect 288 -1455 291 -1449
rect 295 -1455 298 -1449
rect 302 -1455 305 -1449
rect 309 -1455 312 -1449
rect 316 -1455 319 -1449
rect 323 -1455 326 -1449
rect 330 -1455 336 -1449
rect 337 -1455 340 -1449
rect 344 -1455 347 -1449
rect 351 -1455 354 -1449
rect 358 -1455 361 -1449
rect 365 -1455 368 -1449
rect 372 -1455 375 -1449
rect 379 -1455 382 -1449
rect 386 -1455 389 -1449
rect 393 -1455 396 -1449
rect 400 -1455 406 -1449
rect 407 -1455 413 -1449
rect 414 -1455 417 -1449
rect 421 -1455 424 -1449
rect 428 -1455 434 -1449
rect 435 -1455 441 -1449
rect 442 -1455 448 -1449
rect 449 -1455 452 -1449
rect 456 -1455 459 -1449
rect 463 -1455 466 -1449
rect 470 -1455 473 -1449
rect 477 -1455 483 -1449
rect 484 -1455 490 -1449
rect 491 -1455 497 -1449
rect 498 -1455 504 -1449
rect 505 -1455 511 -1449
rect 512 -1455 515 -1449
rect 519 -1455 522 -1449
rect 526 -1455 529 -1449
rect 533 -1455 536 -1449
rect 540 -1455 543 -1449
rect 547 -1455 553 -1449
rect 554 -1455 557 -1449
rect 561 -1455 564 -1449
rect 568 -1455 574 -1449
rect 575 -1455 581 -1449
rect 582 -1455 585 -1449
rect 589 -1455 592 -1449
rect 596 -1455 602 -1449
rect 603 -1455 606 -1449
rect 610 -1455 616 -1449
rect 617 -1455 620 -1449
rect 624 -1455 627 -1449
rect 631 -1455 634 -1449
rect 638 -1455 641 -1449
rect 645 -1455 648 -1449
rect 652 -1455 655 -1449
rect 659 -1455 662 -1449
rect 666 -1455 669 -1449
rect 673 -1455 676 -1449
rect 680 -1455 683 -1449
rect 687 -1455 693 -1449
rect 694 -1455 697 -1449
rect 701 -1455 707 -1449
rect 708 -1455 711 -1449
rect 715 -1455 718 -1449
rect 722 -1455 725 -1449
rect 729 -1455 732 -1449
rect 736 -1455 739 -1449
rect 743 -1455 749 -1449
rect 750 -1455 753 -1449
rect 757 -1455 760 -1449
rect 764 -1455 767 -1449
rect 771 -1455 774 -1449
rect 778 -1455 781 -1449
rect 785 -1455 788 -1449
rect 792 -1455 795 -1449
rect 799 -1455 802 -1449
rect 806 -1455 809 -1449
rect 813 -1455 816 -1449
rect 820 -1455 823 -1449
rect 827 -1455 830 -1449
rect 834 -1455 837 -1449
rect 841 -1455 844 -1449
rect 848 -1455 851 -1449
rect 855 -1455 861 -1449
rect 862 -1455 865 -1449
rect 869 -1455 872 -1449
rect 876 -1455 879 -1449
rect 883 -1455 886 -1449
rect 890 -1455 893 -1449
rect 897 -1455 900 -1449
rect 904 -1455 907 -1449
rect 911 -1455 914 -1449
rect 918 -1455 921 -1449
rect 925 -1455 928 -1449
rect 932 -1455 935 -1449
rect 939 -1455 942 -1449
rect 946 -1455 949 -1449
rect 953 -1455 956 -1449
rect 960 -1455 963 -1449
rect 967 -1455 970 -1449
rect 974 -1455 977 -1449
rect 981 -1455 984 -1449
rect 988 -1455 991 -1449
rect 995 -1455 998 -1449
rect 1002 -1455 1005 -1449
rect 1009 -1455 1012 -1449
rect 1016 -1455 1019 -1449
rect 1023 -1455 1026 -1449
rect 1030 -1455 1033 -1449
rect 1037 -1455 1040 -1449
rect 1044 -1455 1047 -1449
rect 1051 -1455 1054 -1449
rect 1058 -1455 1064 -1449
rect 1065 -1455 1068 -1449
rect 1072 -1455 1075 -1449
rect 1079 -1455 1082 -1449
rect 1086 -1455 1092 -1449
rect 1093 -1455 1096 -1449
rect 1107 -1455 1110 -1449
rect 1 -1546 4 -1540
rect 8 -1546 11 -1540
rect 15 -1546 18 -1540
rect 22 -1546 25 -1540
rect 29 -1546 35 -1540
rect 36 -1546 42 -1540
rect 43 -1546 46 -1540
rect 50 -1546 53 -1540
rect 57 -1546 60 -1540
rect 64 -1546 67 -1540
rect 71 -1546 74 -1540
rect 78 -1546 81 -1540
rect 85 -1546 88 -1540
rect 92 -1546 98 -1540
rect 99 -1546 102 -1540
rect 106 -1546 109 -1540
rect 113 -1546 116 -1540
rect 120 -1546 123 -1540
rect 127 -1546 130 -1540
rect 134 -1546 137 -1540
rect 141 -1546 147 -1540
rect 148 -1546 151 -1540
rect 155 -1546 161 -1540
rect 162 -1546 168 -1540
rect 169 -1546 172 -1540
rect 176 -1546 182 -1540
rect 183 -1546 186 -1540
rect 190 -1546 193 -1540
rect 197 -1546 200 -1540
rect 204 -1546 210 -1540
rect 211 -1546 217 -1540
rect 218 -1546 224 -1540
rect 225 -1546 228 -1540
rect 232 -1546 235 -1540
rect 239 -1546 242 -1540
rect 246 -1546 252 -1540
rect 253 -1546 256 -1540
rect 260 -1546 263 -1540
rect 267 -1546 270 -1540
rect 274 -1546 280 -1540
rect 281 -1546 284 -1540
rect 288 -1546 294 -1540
rect 295 -1546 298 -1540
rect 302 -1546 305 -1540
rect 309 -1546 312 -1540
rect 316 -1546 319 -1540
rect 323 -1546 329 -1540
rect 330 -1546 333 -1540
rect 337 -1546 340 -1540
rect 344 -1546 347 -1540
rect 351 -1546 354 -1540
rect 358 -1546 364 -1540
rect 365 -1546 368 -1540
rect 372 -1546 375 -1540
rect 379 -1546 382 -1540
rect 386 -1546 389 -1540
rect 393 -1546 396 -1540
rect 400 -1546 403 -1540
rect 407 -1546 410 -1540
rect 414 -1546 417 -1540
rect 421 -1546 424 -1540
rect 428 -1546 431 -1540
rect 435 -1546 438 -1540
rect 442 -1546 445 -1540
rect 449 -1546 452 -1540
rect 456 -1546 462 -1540
rect 463 -1546 469 -1540
rect 470 -1546 476 -1540
rect 477 -1546 483 -1540
rect 484 -1546 490 -1540
rect 491 -1546 494 -1540
rect 498 -1546 501 -1540
rect 505 -1546 508 -1540
rect 512 -1546 518 -1540
rect 519 -1546 525 -1540
rect 526 -1546 529 -1540
rect 533 -1546 539 -1540
rect 540 -1546 543 -1540
rect 547 -1546 550 -1540
rect 554 -1546 557 -1540
rect 561 -1546 567 -1540
rect 568 -1546 571 -1540
rect 575 -1546 578 -1540
rect 582 -1546 585 -1540
rect 589 -1546 595 -1540
rect 596 -1546 599 -1540
rect 603 -1546 606 -1540
rect 610 -1546 613 -1540
rect 617 -1546 620 -1540
rect 624 -1546 627 -1540
rect 631 -1546 634 -1540
rect 638 -1546 641 -1540
rect 645 -1546 648 -1540
rect 652 -1546 655 -1540
rect 659 -1546 665 -1540
rect 666 -1546 672 -1540
rect 673 -1546 679 -1540
rect 680 -1546 683 -1540
rect 687 -1546 693 -1540
rect 694 -1546 697 -1540
rect 701 -1546 704 -1540
rect 708 -1546 711 -1540
rect 715 -1546 718 -1540
rect 722 -1546 725 -1540
rect 729 -1546 732 -1540
rect 736 -1546 739 -1540
rect 743 -1546 746 -1540
rect 750 -1546 753 -1540
rect 757 -1546 760 -1540
rect 764 -1546 767 -1540
rect 771 -1546 777 -1540
rect 778 -1546 781 -1540
rect 785 -1546 788 -1540
rect 792 -1546 795 -1540
rect 799 -1546 802 -1540
rect 806 -1546 809 -1540
rect 813 -1546 816 -1540
rect 820 -1546 823 -1540
rect 827 -1546 830 -1540
rect 834 -1546 837 -1540
rect 841 -1546 844 -1540
rect 848 -1546 851 -1540
rect 855 -1546 858 -1540
rect 862 -1546 865 -1540
rect 869 -1546 872 -1540
rect 876 -1546 879 -1540
rect 883 -1546 886 -1540
rect 890 -1546 893 -1540
rect 897 -1546 900 -1540
rect 904 -1546 907 -1540
rect 911 -1546 914 -1540
rect 918 -1546 921 -1540
rect 925 -1546 928 -1540
rect 932 -1546 935 -1540
rect 939 -1546 942 -1540
rect 946 -1546 949 -1540
rect 953 -1546 956 -1540
rect 960 -1546 963 -1540
rect 967 -1546 970 -1540
rect 974 -1546 977 -1540
rect 981 -1546 984 -1540
rect 988 -1546 991 -1540
rect 995 -1546 998 -1540
rect 1002 -1546 1005 -1540
rect 1009 -1546 1015 -1540
rect 1016 -1546 1019 -1540
rect 1023 -1546 1026 -1540
rect 1030 -1546 1036 -1540
rect 1037 -1546 1040 -1540
rect 1044 -1546 1047 -1540
rect 1058 -1546 1061 -1540
rect 1072 -1546 1075 -1540
rect 1093 -1546 1096 -1540
rect 1 -1635 7 -1629
rect 8 -1635 11 -1629
rect 15 -1635 18 -1629
rect 22 -1635 25 -1629
rect 29 -1635 32 -1629
rect 36 -1635 39 -1629
rect 43 -1635 46 -1629
rect 50 -1635 53 -1629
rect 57 -1635 63 -1629
rect 64 -1635 67 -1629
rect 71 -1635 74 -1629
rect 78 -1635 84 -1629
rect 85 -1635 88 -1629
rect 92 -1635 98 -1629
rect 99 -1635 102 -1629
rect 106 -1635 109 -1629
rect 113 -1635 116 -1629
rect 120 -1635 123 -1629
rect 127 -1635 130 -1629
rect 134 -1635 140 -1629
rect 141 -1635 147 -1629
rect 148 -1635 151 -1629
rect 155 -1635 158 -1629
rect 162 -1635 165 -1629
rect 169 -1635 172 -1629
rect 176 -1635 179 -1629
rect 183 -1635 189 -1629
rect 190 -1635 196 -1629
rect 197 -1635 203 -1629
rect 204 -1635 207 -1629
rect 211 -1635 214 -1629
rect 218 -1635 224 -1629
rect 225 -1635 231 -1629
rect 232 -1635 235 -1629
rect 239 -1635 242 -1629
rect 246 -1635 252 -1629
rect 253 -1635 256 -1629
rect 260 -1635 263 -1629
rect 267 -1635 270 -1629
rect 274 -1635 277 -1629
rect 281 -1635 284 -1629
rect 288 -1635 291 -1629
rect 295 -1635 298 -1629
rect 302 -1635 308 -1629
rect 309 -1635 312 -1629
rect 316 -1635 319 -1629
rect 323 -1635 329 -1629
rect 330 -1635 333 -1629
rect 337 -1635 340 -1629
rect 344 -1635 347 -1629
rect 351 -1635 357 -1629
rect 358 -1635 361 -1629
rect 365 -1635 368 -1629
rect 372 -1635 378 -1629
rect 379 -1635 382 -1629
rect 386 -1635 389 -1629
rect 393 -1635 396 -1629
rect 400 -1635 403 -1629
rect 407 -1635 410 -1629
rect 414 -1635 417 -1629
rect 421 -1635 427 -1629
rect 428 -1635 431 -1629
rect 435 -1635 438 -1629
rect 442 -1635 448 -1629
rect 449 -1635 452 -1629
rect 456 -1635 462 -1629
rect 463 -1635 469 -1629
rect 470 -1635 473 -1629
rect 477 -1635 480 -1629
rect 484 -1635 487 -1629
rect 491 -1635 494 -1629
rect 498 -1635 501 -1629
rect 505 -1635 508 -1629
rect 512 -1635 515 -1629
rect 519 -1635 522 -1629
rect 526 -1635 529 -1629
rect 533 -1635 539 -1629
rect 540 -1635 543 -1629
rect 547 -1635 550 -1629
rect 554 -1635 557 -1629
rect 561 -1635 564 -1629
rect 568 -1635 574 -1629
rect 575 -1635 578 -1629
rect 582 -1635 588 -1629
rect 589 -1635 592 -1629
rect 596 -1635 599 -1629
rect 603 -1635 606 -1629
rect 610 -1635 616 -1629
rect 617 -1635 620 -1629
rect 624 -1635 630 -1629
rect 631 -1635 637 -1629
rect 638 -1635 641 -1629
rect 645 -1635 648 -1629
rect 652 -1635 655 -1629
rect 659 -1635 662 -1629
rect 666 -1635 669 -1629
rect 673 -1635 679 -1629
rect 680 -1635 686 -1629
rect 687 -1635 690 -1629
rect 694 -1635 697 -1629
rect 701 -1635 704 -1629
rect 708 -1635 711 -1629
rect 715 -1635 718 -1629
rect 722 -1635 725 -1629
rect 729 -1635 732 -1629
rect 736 -1635 739 -1629
rect 743 -1635 746 -1629
rect 750 -1635 753 -1629
rect 757 -1635 760 -1629
rect 764 -1635 767 -1629
rect 771 -1635 774 -1629
rect 778 -1635 784 -1629
rect 785 -1635 788 -1629
rect 792 -1635 795 -1629
rect 799 -1635 802 -1629
rect 806 -1635 809 -1629
rect 813 -1635 816 -1629
rect 820 -1635 823 -1629
rect 827 -1635 830 -1629
rect 834 -1635 837 -1629
rect 841 -1635 844 -1629
rect 848 -1635 851 -1629
rect 855 -1635 861 -1629
rect 862 -1635 865 -1629
rect 869 -1635 872 -1629
rect 876 -1635 879 -1629
rect 883 -1635 886 -1629
rect 890 -1635 893 -1629
rect 897 -1635 900 -1629
rect 904 -1635 907 -1629
rect 911 -1635 914 -1629
rect 918 -1635 921 -1629
rect 925 -1635 928 -1629
rect 932 -1635 935 -1629
rect 939 -1635 942 -1629
rect 946 -1635 949 -1629
rect 953 -1635 956 -1629
rect 960 -1635 963 -1629
rect 967 -1635 970 -1629
rect 974 -1635 977 -1629
rect 981 -1635 984 -1629
rect 988 -1635 991 -1629
rect 995 -1635 998 -1629
rect 1002 -1635 1005 -1629
rect 1009 -1635 1012 -1629
rect 1016 -1635 1019 -1629
rect 1023 -1635 1026 -1629
rect 1030 -1635 1033 -1629
rect 1037 -1635 1040 -1629
rect 1044 -1635 1047 -1629
rect 1051 -1635 1054 -1629
rect 1058 -1635 1064 -1629
rect 1065 -1635 1071 -1629
rect 1072 -1635 1075 -1629
rect 1079 -1635 1082 -1629
rect 1086 -1635 1089 -1629
rect 1093 -1635 1096 -1629
rect 1100 -1635 1103 -1629
rect 1107 -1635 1110 -1629
rect 1114 -1635 1117 -1629
rect 22 -1720 25 -1714
rect 29 -1720 32 -1714
rect 36 -1720 39 -1714
rect 43 -1720 46 -1714
rect 50 -1720 56 -1714
rect 57 -1720 60 -1714
rect 64 -1720 70 -1714
rect 71 -1720 74 -1714
rect 78 -1720 81 -1714
rect 85 -1720 88 -1714
rect 92 -1720 95 -1714
rect 99 -1720 102 -1714
rect 106 -1720 109 -1714
rect 113 -1720 116 -1714
rect 120 -1720 123 -1714
rect 127 -1720 130 -1714
rect 134 -1720 137 -1714
rect 141 -1720 144 -1714
rect 148 -1720 151 -1714
rect 155 -1720 161 -1714
rect 162 -1720 165 -1714
rect 169 -1720 172 -1714
rect 176 -1720 179 -1714
rect 183 -1720 186 -1714
rect 190 -1720 193 -1714
rect 197 -1720 200 -1714
rect 204 -1720 207 -1714
rect 211 -1720 214 -1714
rect 218 -1720 224 -1714
rect 225 -1720 228 -1714
rect 232 -1720 235 -1714
rect 239 -1720 242 -1714
rect 246 -1720 249 -1714
rect 253 -1720 256 -1714
rect 260 -1720 263 -1714
rect 267 -1720 270 -1714
rect 274 -1720 277 -1714
rect 281 -1720 284 -1714
rect 288 -1720 291 -1714
rect 295 -1720 298 -1714
rect 302 -1720 308 -1714
rect 309 -1720 315 -1714
rect 316 -1720 319 -1714
rect 323 -1720 329 -1714
rect 330 -1720 333 -1714
rect 337 -1720 343 -1714
rect 344 -1720 347 -1714
rect 351 -1720 357 -1714
rect 358 -1720 364 -1714
rect 365 -1720 368 -1714
rect 372 -1720 378 -1714
rect 379 -1720 385 -1714
rect 386 -1720 389 -1714
rect 393 -1720 396 -1714
rect 400 -1720 403 -1714
rect 407 -1720 410 -1714
rect 414 -1720 417 -1714
rect 421 -1720 427 -1714
rect 428 -1720 434 -1714
rect 435 -1720 438 -1714
rect 442 -1720 445 -1714
rect 449 -1720 452 -1714
rect 456 -1720 459 -1714
rect 463 -1720 466 -1714
rect 470 -1720 473 -1714
rect 477 -1720 483 -1714
rect 484 -1720 490 -1714
rect 491 -1720 497 -1714
rect 498 -1720 501 -1714
rect 505 -1720 508 -1714
rect 512 -1720 515 -1714
rect 519 -1720 525 -1714
rect 526 -1720 532 -1714
rect 533 -1720 536 -1714
rect 540 -1720 543 -1714
rect 547 -1720 550 -1714
rect 554 -1720 557 -1714
rect 561 -1720 564 -1714
rect 568 -1720 571 -1714
rect 575 -1720 581 -1714
rect 582 -1720 588 -1714
rect 589 -1720 592 -1714
rect 596 -1720 599 -1714
rect 603 -1720 609 -1714
rect 610 -1720 613 -1714
rect 617 -1720 620 -1714
rect 624 -1720 627 -1714
rect 631 -1720 634 -1714
rect 638 -1720 641 -1714
rect 645 -1720 648 -1714
rect 652 -1720 658 -1714
rect 659 -1720 665 -1714
rect 666 -1720 669 -1714
rect 673 -1720 679 -1714
rect 680 -1720 683 -1714
rect 687 -1720 693 -1714
rect 694 -1720 697 -1714
rect 701 -1720 704 -1714
rect 708 -1720 711 -1714
rect 715 -1720 718 -1714
rect 722 -1720 725 -1714
rect 729 -1720 732 -1714
rect 736 -1720 739 -1714
rect 743 -1720 746 -1714
rect 750 -1720 756 -1714
rect 757 -1720 763 -1714
rect 764 -1720 767 -1714
rect 771 -1720 774 -1714
rect 778 -1720 781 -1714
rect 785 -1720 788 -1714
rect 792 -1720 795 -1714
rect 799 -1720 802 -1714
rect 806 -1720 809 -1714
rect 813 -1720 819 -1714
rect 820 -1720 823 -1714
rect 827 -1720 830 -1714
rect 834 -1720 837 -1714
rect 841 -1720 844 -1714
rect 848 -1720 851 -1714
rect 855 -1720 858 -1714
rect 862 -1720 865 -1714
rect 869 -1720 872 -1714
rect 876 -1720 879 -1714
rect 883 -1720 886 -1714
rect 890 -1720 893 -1714
rect 897 -1720 900 -1714
rect 904 -1720 910 -1714
rect 911 -1720 914 -1714
rect 918 -1720 921 -1714
rect 925 -1720 931 -1714
rect 932 -1720 935 -1714
rect 939 -1720 942 -1714
rect 946 -1720 949 -1714
rect 953 -1720 956 -1714
rect 960 -1720 963 -1714
rect 967 -1720 970 -1714
rect 1065 -1720 1071 -1714
rect 1093 -1720 1096 -1714
rect 1 -1811 4 -1805
rect 8 -1811 14 -1805
rect 15 -1811 18 -1805
rect 22 -1811 25 -1805
rect 29 -1811 32 -1805
rect 36 -1811 39 -1805
rect 43 -1811 46 -1805
rect 50 -1811 53 -1805
rect 57 -1811 60 -1805
rect 64 -1811 67 -1805
rect 71 -1811 74 -1805
rect 78 -1811 81 -1805
rect 85 -1811 88 -1805
rect 92 -1811 98 -1805
rect 99 -1811 105 -1805
rect 106 -1811 112 -1805
rect 113 -1811 119 -1805
rect 120 -1811 123 -1805
rect 127 -1811 130 -1805
rect 134 -1811 140 -1805
rect 141 -1811 144 -1805
rect 148 -1811 154 -1805
rect 155 -1811 158 -1805
rect 162 -1811 165 -1805
rect 169 -1811 172 -1805
rect 176 -1811 179 -1805
rect 183 -1811 189 -1805
rect 190 -1811 193 -1805
rect 197 -1811 203 -1805
rect 204 -1811 210 -1805
rect 211 -1811 214 -1805
rect 218 -1811 224 -1805
rect 225 -1811 228 -1805
rect 232 -1811 235 -1805
rect 239 -1811 242 -1805
rect 246 -1811 252 -1805
rect 253 -1811 256 -1805
rect 260 -1811 263 -1805
rect 267 -1811 270 -1805
rect 274 -1811 277 -1805
rect 281 -1811 284 -1805
rect 288 -1811 291 -1805
rect 295 -1811 298 -1805
rect 302 -1811 308 -1805
rect 309 -1811 312 -1805
rect 316 -1811 319 -1805
rect 323 -1811 326 -1805
rect 330 -1811 333 -1805
rect 337 -1811 340 -1805
rect 344 -1811 350 -1805
rect 351 -1811 357 -1805
rect 358 -1811 361 -1805
rect 365 -1811 368 -1805
rect 372 -1811 375 -1805
rect 379 -1811 382 -1805
rect 386 -1811 389 -1805
rect 393 -1811 396 -1805
rect 400 -1811 403 -1805
rect 407 -1811 410 -1805
rect 414 -1811 420 -1805
rect 421 -1811 427 -1805
rect 428 -1811 434 -1805
rect 435 -1811 438 -1805
rect 442 -1811 445 -1805
rect 449 -1811 452 -1805
rect 456 -1811 459 -1805
rect 463 -1811 466 -1805
rect 470 -1811 473 -1805
rect 477 -1811 480 -1805
rect 484 -1811 487 -1805
rect 491 -1811 494 -1805
rect 498 -1811 504 -1805
rect 505 -1811 508 -1805
rect 512 -1811 515 -1805
rect 519 -1811 525 -1805
rect 526 -1811 532 -1805
rect 533 -1811 536 -1805
rect 540 -1811 543 -1805
rect 547 -1811 553 -1805
rect 554 -1811 557 -1805
rect 561 -1811 564 -1805
rect 568 -1811 571 -1805
rect 575 -1811 578 -1805
rect 582 -1811 585 -1805
rect 589 -1811 592 -1805
rect 596 -1811 602 -1805
rect 603 -1811 609 -1805
rect 610 -1811 616 -1805
rect 617 -1811 620 -1805
rect 624 -1811 630 -1805
rect 631 -1811 634 -1805
rect 638 -1811 641 -1805
rect 645 -1811 648 -1805
rect 652 -1811 655 -1805
rect 659 -1811 662 -1805
rect 666 -1811 672 -1805
rect 673 -1811 676 -1805
rect 680 -1811 683 -1805
rect 687 -1811 693 -1805
rect 694 -1811 697 -1805
rect 701 -1811 704 -1805
rect 708 -1811 714 -1805
rect 715 -1811 718 -1805
rect 722 -1811 725 -1805
rect 729 -1811 732 -1805
rect 736 -1811 739 -1805
rect 743 -1811 746 -1805
rect 750 -1811 753 -1805
rect 757 -1811 760 -1805
rect 764 -1811 770 -1805
rect 771 -1811 774 -1805
rect 778 -1811 781 -1805
rect 785 -1811 788 -1805
rect 792 -1811 795 -1805
rect 799 -1811 802 -1805
rect 806 -1811 809 -1805
rect 813 -1811 816 -1805
rect 820 -1811 823 -1805
rect 827 -1811 830 -1805
rect 834 -1811 837 -1805
rect 841 -1811 844 -1805
rect 848 -1811 851 -1805
rect 855 -1811 858 -1805
rect 862 -1811 865 -1805
rect 869 -1811 872 -1805
rect 876 -1811 879 -1805
rect 883 -1811 886 -1805
rect 890 -1811 893 -1805
rect 897 -1811 900 -1805
rect 904 -1811 907 -1805
rect 911 -1811 914 -1805
rect 918 -1811 921 -1805
rect 925 -1811 928 -1805
rect 932 -1811 938 -1805
rect 939 -1811 942 -1805
rect 946 -1811 949 -1805
rect 953 -1811 956 -1805
rect 960 -1811 963 -1805
rect 967 -1811 970 -1805
rect 974 -1811 977 -1805
rect 981 -1811 984 -1805
rect 988 -1811 991 -1805
rect 995 -1811 998 -1805
rect 1002 -1811 1005 -1805
rect 1009 -1811 1012 -1805
rect 1016 -1811 1019 -1805
rect 1023 -1811 1026 -1805
rect 1030 -1811 1033 -1805
rect 1037 -1811 1040 -1805
rect 1044 -1811 1047 -1805
rect 1051 -1811 1057 -1805
rect 1058 -1811 1061 -1805
rect 1086 -1811 1089 -1805
rect 1093 -1811 1096 -1805
rect 1 -1902 7 -1896
rect 8 -1902 11 -1896
rect 15 -1902 21 -1896
rect 22 -1902 28 -1896
rect 29 -1902 32 -1896
rect 36 -1902 42 -1896
rect 43 -1902 49 -1896
rect 50 -1902 56 -1896
rect 57 -1902 60 -1896
rect 64 -1902 70 -1896
rect 71 -1902 74 -1896
rect 78 -1902 84 -1896
rect 85 -1902 88 -1896
rect 92 -1902 95 -1896
rect 99 -1902 102 -1896
rect 106 -1902 109 -1896
rect 113 -1902 119 -1896
rect 120 -1902 126 -1896
rect 127 -1902 130 -1896
rect 134 -1902 137 -1896
rect 141 -1902 144 -1896
rect 148 -1902 154 -1896
rect 155 -1902 161 -1896
rect 162 -1902 165 -1896
rect 169 -1902 172 -1896
rect 176 -1902 179 -1896
rect 183 -1902 186 -1896
rect 190 -1902 196 -1896
rect 197 -1902 200 -1896
rect 204 -1902 207 -1896
rect 211 -1902 214 -1896
rect 218 -1902 224 -1896
rect 225 -1902 228 -1896
rect 232 -1902 235 -1896
rect 239 -1902 242 -1896
rect 246 -1902 249 -1896
rect 253 -1902 256 -1896
rect 260 -1902 263 -1896
rect 267 -1902 270 -1896
rect 274 -1902 277 -1896
rect 281 -1902 284 -1896
rect 288 -1902 291 -1896
rect 295 -1902 298 -1896
rect 302 -1902 305 -1896
rect 309 -1902 312 -1896
rect 316 -1902 319 -1896
rect 323 -1902 326 -1896
rect 330 -1902 333 -1896
rect 337 -1902 340 -1896
rect 344 -1902 347 -1896
rect 351 -1902 354 -1896
rect 358 -1902 364 -1896
rect 365 -1902 371 -1896
rect 372 -1902 375 -1896
rect 379 -1902 382 -1896
rect 386 -1902 392 -1896
rect 393 -1902 396 -1896
rect 400 -1902 403 -1896
rect 407 -1902 410 -1896
rect 414 -1902 420 -1896
rect 421 -1902 424 -1896
rect 428 -1902 431 -1896
rect 435 -1902 438 -1896
rect 442 -1902 448 -1896
rect 449 -1902 455 -1896
rect 456 -1902 459 -1896
rect 463 -1902 466 -1896
rect 470 -1902 473 -1896
rect 477 -1902 483 -1896
rect 484 -1902 490 -1896
rect 491 -1902 494 -1896
rect 498 -1902 504 -1896
rect 505 -1902 508 -1896
rect 512 -1902 515 -1896
rect 519 -1902 522 -1896
rect 526 -1902 532 -1896
rect 533 -1902 536 -1896
rect 540 -1902 543 -1896
rect 547 -1902 553 -1896
rect 554 -1902 560 -1896
rect 561 -1902 564 -1896
rect 568 -1902 571 -1896
rect 575 -1902 578 -1896
rect 582 -1902 585 -1896
rect 589 -1902 592 -1896
rect 596 -1902 599 -1896
rect 603 -1902 606 -1896
rect 610 -1902 613 -1896
rect 617 -1902 623 -1896
rect 624 -1902 627 -1896
rect 631 -1902 637 -1896
rect 638 -1902 641 -1896
rect 645 -1902 648 -1896
rect 652 -1902 655 -1896
rect 659 -1902 662 -1896
rect 666 -1902 672 -1896
rect 673 -1902 676 -1896
rect 680 -1902 683 -1896
rect 687 -1902 693 -1896
rect 694 -1902 697 -1896
rect 701 -1902 704 -1896
rect 708 -1902 711 -1896
rect 715 -1902 718 -1896
rect 722 -1902 725 -1896
rect 729 -1902 735 -1896
rect 736 -1902 739 -1896
rect 743 -1902 746 -1896
rect 750 -1902 753 -1896
rect 757 -1902 760 -1896
rect 764 -1902 767 -1896
rect 771 -1902 774 -1896
rect 778 -1902 781 -1896
rect 785 -1902 788 -1896
rect 792 -1902 795 -1896
rect 799 -1902 802 -1896
rect 806 -1902 809 -1896
rect 813 -1902 816 -1896
rect 820 -1902 823 -1896
rect 827 -1902 830 -1896
rect 834 -1902 837 -1896
rect 841 -1902 844 -1896
rect 848 -1902 851 -1896
rect 855 -1902 858 -1896
rect 862 -1902 865 -1896
rect 869 -1902 872 -1896
rect 876 -1902 879 -1896
rect 883 -1902 886 -1896
rect 890 -1902 893 -1896
rect 897 -1902 900 -1896
rect 904 -1902 907 -1896
rect 911 -1902 914 -1896
rect 918 -1902 921 -1896
rect 925 -1902 928 -1896
rect 932 -1902 935 -1896
rect 939 -1902 942 -1896
rect 946 -1902 949 -1896
rect 953 -1902 956 -1896
rect 960 -1902 963 -1896
rect 967 -1902 970 -1896
rect 974 -1902 977 -1896
rect 981 -1902 984 -1896
rect 988 -1902 991 -1896
rect 995 -1902 998 -1896
rect 1002 -1902 1005 -1896
rect 1009 -1902 1012 -1896
rect 1016 -1902 1019 -1896
rect 1023 -1902 1026 -1896
rect 1030 -1902 1033 -1896
rect 1037 -1902 1040 -1896
rect 1044 -1902 1047 -1896
rect 1051 -1902 1054 -1896
rect 1058 -1902 1061 -1896
rect 1065 -1902 1071 -1896
rect 1072 -1902 1075 -1896
rect 1086 -1902 1089 -1896
rect 1100 -1902 1103 -1896
rect 1 -2007 7 -2001
rect 8 -2007 11 -2001
rect 15 -2007 18 -2001
rect 22 -2007 28 -2001
rect 29 -2007 35 -2001
rect 36 -2007 39 -2001
rect 43 -2007 46 -2001
rect 50 -2007 56 -2001
rect 57 -2007 63 -2001
rect 64 -2007 67 -2001
rect 71 -2007 77 -2001
rect 78 -2007 84 -2001
rect 85 -2007 91 -2001
rect 92 -2007 95 -2001
rect 99 -2007 102 -2001
rect 106 -2007 112 -2001
rect 113 -2007 116 -2001
rect 120 -2007 123 -2001
rect 127 -2007 130 -2001
rect 134 -2007 140 -2001
rect 141 -2007 144 -2001
rect 148 -2007 154 -2001
rect 155 -2007 158 -2001
rect 162 -2007 165 -2001
rect 169 -2007 172 -2001
rect 176 -2007 182 -2001
rect 183 -2007 186 -2001
rect 190 -2007 193 -2001
rect 197 -2007 200 -2001
rect 204 -2007 210 -2001
rect 211 -2007 214 -2001
rect 218 -2007 224 -2001
rect 225 -2007 231 -2001
rect 232 -2007 235 -2001
rect 239 -2007 242 -2001
rect 246 -2007 249 -2001
rect 253 -2007 256 -2001
rect 260 -2007 263 -2001
rect 267 -2007 270 -2001
rect 274 -2007 277 -2001
rect 281 -2007 284 -2001
rect 288 -2007 291 -2001
rect 295 -2007 298 -2001
rect 302 -2007 305 -2001
rect 309 -2007 312 -2001
rect 316 -2007 319 -2001
rect 323 -2007 326 -2001
rect 330 -2007 333 -2001
rect 337 -2007 340 -2001
rect 344 -2007 350 -2001
rect 351 -2007 354 -2001
rect 358 -2007 361 -2001
rect 365 -2007 371 -2001
rect 372 -2007 378 -2001
rect 379 -2007 382 -2001
rect 386 -2007 389 -2001
rect 393 -2007 396 -2001
rect 400 -2007 403 -2001
rect 407 -2007 413 -2001
rect 414 -2007 417 -2001
rect 421 -2007 424 -2001
rect 428 -2007 431 -2001
rect 435 -2007 441 -2001
rect 442 -2007 445 -2001
rect 449 -2007 452 -2001
rect 456 -2007 459 -2001
rect 463 -2007 466 -2001
rect 470 -2007 473 -2001
rect 477 -2007 480 -2001
rect 484 -2007 487 -2001
rect 491 -2007 494 -2001
rect 498 -2007 501 -2001
rect 505 -2007 508 -2001
rect 512 -2007 518 -2001
rect 519 -2007 522 -2001
rect 526 -2007 532 -2001
rect 533 -2007 536 -2001
rect 540 -2007 543 -2001
rect 547 -2007 550 -2001
rect 554 -2007 557 -2001
rect 561 -2007 564 -2001
rect 568 -2007 571 -2001
rect 575 -2007 578 -2001
rect 582 -2007 585 -2001
rect 589 -2007 595 -2001
rect 596 -2007 599 -2001
rect 603 -2007 606 -2001
rect 610 -2007 613 -2001
rect 617 -2007 623 -2001
rect 624 -2007 627 -2001
rect 631 -2007 637 -2001
rect 638 -2007 641 -2001
rect 645 -2007 651 -2001
rect 652 -2007 655 -2001
rect 659 -2007 662 -2001
rect 666 -2007 669 -2001
rect 673 -2007 676 -2001
rect 680 -2007 683 -2001
rect 687 -2007 690 -2001
rect 694 -2007 697 -2001
rect 701 -2007 704 -2001
rect 708 -2007 711 -2001
rect 715 -2007 718 -2001
rect 722 -2007 725 -2001
rect 729 -2007 732 -2001
rect 736 -2007 739 -2001
rect 743 -2007 749 -2001
rect 750 -2007 753 -2001
rect 757 -2007 760 -2001
rect 764 -2007 770 -2001
rect 771 -2007 774 -2001
rect 778 -2007 784 -2001
rect 785 -2007 788 -2001
rect 792 -2007 795 -2001
rect 799 -2007 802 -2001
rect 806 -2007 809 -2001
rect 813 -2007 816 -2001
rect 820 -2007 823 -2001
rect 827 -2007 830 -2001
rect 834 -2007 837 -2001
rect 841 -2007 844 -2001
rect 848 -2007 851 -2001
rect 855 -2007 858 -2001
rect 862 -2007 865 -2001
rect 869 -2007 872 -2001
rect 876 -2007 879 -2001
rect 883 -2007 886 -2001
rect 890 -2007 893 -2001
rect 897 -2007 900 -2001
rect 904 -2007 907 -2001
rect 911 -2007 914 -2001
rect 918 -2007 921 -2001
rect 925 -2007 931 -2001
rect 932 -2007 935 -2001
rect 939 -2007 942 -2001
rect 946 -2007 949 -2001
rect 953 -2007 956 -2001
rect 960 -2007 963 -2001
rect 967 -2007 970 -2001
rect 974 -2007 977 -2001
rect 981 -2007 984 -2001
rect 988 -2007 991 -2001
rect 995 -2007 998 -2001
rect 1002 -2007 1005 -2001
rect 1009 -2007 1012 -2001
rect 1016 -2007 1019 -2001
rect 1023 -2007 1026 -2001
rect 1030 -2007 1033 -2001
rect 1037 -2007 1040 -2001
rect 1044 -2007 1047 -2001
rect 1051 -2007 1054 -2001
rect 1058 -2007 1061 -2001
rect 1065 -2007 1068 -2001
rect 1072 -2007 1075 -2001
rect 1079 -2007 1082 -2001
rect 1086 -2007 1089 -2001
rect 1093 -2007 1099 -2001
rect 1100 -2007 1106 -2001
rect 1107 -2007 1110 -2001
rect 1114 -2007 1117 -2001
rect 1 -2120 4 -2114
rect 8 -2120 11 -2114
rect 15 -2120 18 -2114
rect 22 -2120 25 -2114
rect 29 -2120 32 -2114
rect 36 -2120 39 -2114
rect 43 -2120 46 -2114
rect 50 -2120 53 -2114
rect 57 -2120 63 -2114
rect 64 -2120 67 -2114
rect 71 -2120 77 -2114
rect 78 -2120 84 -2114
rect 85 -2120 91 -2114
rect 92 -2120 98 -2114
rect 99 -2120 102 -2114
rect 106 -2120 112 -2114
rect 113 -2120 119 -2114
rect 120 -2120 126 -2114
rect 127 -2120 130 -2114
rect 134 -2120 140 -2114
rect 141 -2120 144 -2114
rect 148 -2120 154 -2114
rect 155 -2120 158 -2114
rect 162 -2120 165 -2114
rect 169 -2120 172 -2114
rect 176 -2120 179 -2114
rect 183 -2120 186 -2114
rect 190 -2120 193 -2114
rect 197 -2120 200 -2114
rect 204 -2120 207 -2114
rect 211 -2120 214 -2114
rect 218 -2120 224 -2114
rect 225 -2120 228 -2114
rect 232 -2120 235 -2114
rect 239 -2120 242 -2114
rect 246 -2120 249 -2114
rect 253 -2120 256 -2114
rect 260 -2120 263 -2114
rect 267 -2120 270 -2114
rect 274 -2120 277 -2114
rect 281 -2120 284 -2114
rect 288 -2120 294 -2114
rect 295 -2120 298 -2114
rect 302 -2120 305 -2114
rect 309 -2120 312 -2114
rect 316 -2120 319 -2114
rect 323 -2120 326 -2114
rect 330 -2120 333 -2114
rect 337 -2120 343 -2114
rect 344 -2120 347 -2114
rect 351 -2120 357 -2114
rect 358 -2120 361 -2114
rect 365 -2120 368 -2114
rect 372 -2120 375 -2114
rect 379 -2120 382 -2114
rect 386 -2120 389 -2114
rect 393 -2120 396 -2114
rect 400 -2120 403 -2114
rect 407 -2120 413 -2114
rect 414 -2120 420 -2114
rect 421 -2120 424 -2114
rect 428 -2120 431 -2114
rect 435 -2120 438 -2114
rect 442 -2120 445 -2114
rect 449 -2120 455 -2114
rect 456 -2120 462 -2114
rect 463 -2120 466 -2114
rect 470 -2120 473 -2114
rect 477 -2120 480 -2114
rect 484 -2120 487 -2114
rect 491 -2120 494 -2114
rect 498 -2120 504 -2114
rect 505 -2120 508 -2114
rect 512 -2120 515 -2114
rect 519 -2120 522 -2114
rect 526 -2120 532 -2114
rect 533 -2120 536 -2114
rect 540 -2120 543 -2114
rect 547 -2120 553 -2114
rect 554 -2120 557 -2114
rect 561 -2120 564 -2114
rect 568 -2120 574 -2114
rect 575 -2120 581 -2114
rect 582 -2120 585 -2114
rect 589 -2120 592 -2114
rect 596 -2120 599 -2114
rect 603 -2120 606 -2114
rect 610 -2120 616 -2114
rect 617 -2120 620 -2114
rect 624 -2120 630 -2114
rect 631 -2120 634 -2114
rect 638 -2120 644 -2114
rect 645 -2120 648 -2114
rect 652 -2120 658 -2114
rect 659 -2120 662 -2114
rect 666 -2120 669 -2114
rect 673 -2120 676 -2114
rect 680 -2120 683 -2114
rect 687 -2120 693 -2114
rect 694 -2120 697 -2114
rect 701 -2120 704 -2114
rect 708 -2120 711 -2114
rect 715 -2120 718 -2114
rect 722 -2120 725 -2114
rect 729 -2120 732 -2114
rect 736 -2120 742 -2114
rect 743 -2120 746 -2114
rect 750 -2120 753 -2114
rect 757 -2120 763 -2114
rect 764 -2120 767 -2114
rect 771 -2120 774 -2114
rect 778 -2120 781 -2114
rect 785 -2120 788 -2114
rect 792 -2120 795 -2114
rect 799 -2120 802 -2114
rect 806 -2120 809 -2114
rect 813 -2120 816 -2114
rect 820 -2120 823 -2114
rect 827 -2120 830 -2114
rect 834 -2120 837 -2114
rect 841 -2120 844 -2114
rect 848 -2120 851 -2114
rect 855 -2120 858 -2114
rect 862 -2120 865 -2114
rect 869 -2120 872 -2114
rect 876 -2120 879 -2114
rect 883 -2120 886 -2114
rect 890 -2120 893 -2114
rect 897 -2120 900 -2114
rect 904 -2120 907 -2114
rect 911 -2120 914 -2114
rect 918 -2120 921 -2114
rect 925 -2120 928 -2114
rect 932 -2120 935 -2114
rect 939 -2120 945 -2114
rect 946 -2120 949 -2114
rect 953 -2120 956 -2114
rect 960 -2120 963 -2114
rect 967 -2120 970 -2114
rect 974 -2120 977 -2114
rect 981 -2120 984 -2114
rect 988 -2120 991 -2114
rect 995 -2120 998 -2114
rect 1002 -2120 1005 -2114
rect 1009 -2120 1012 -2114
rect 1016 -2120 1019 -2114
rect 1023 -2120 1026 -2114
rect 1030 -2120 1033 -2114
rect 1037 -2120 1040 -2114
rect 1044 -2120 1047 -2114
rect 1051 -2120 1054 -2114
rect 1058 -2120 1061 -2114
rect 1065 -2120 1068 -2114
rect 1072 -2120 1075 -2114
rect 1079 -2120 1082 -2114
rect 1086 -2120 1089 -2114
rect 1093 -2120 1096 -2114
rect 1100 -2120 1106 -2114
rect 1107 -2120 1110 -2114
rect 1114 -2120 1117 -2114
rect 1121 -2120 1124 -2114
rect 1 -2215 4 -2209
rect 8 -2215 11 -2209
rect 15 -2215 18 -2209
rect 22 -2215 25 -2209
rect 29 -2215 35 -2209
rect 36 -2215 42 -2209
rect 43 -2215 46 -2209
rect 50 -2215 53 -2209
rect 57 -2215 60 -2209
rect 64 -2215 67 -2209
rect 71 -2215 77 -2209
rect 78 -2215 81 -2209
rect 85 -2215 88 -2209
rect 92 -2215 95 -2209
rect 99 -2215 102 -2209
rect 106 -2215 109 -2209
rect 113 -2215 116 -2209
rect 120 -2215 126 -2209
rect 127 -2215 130 -2209
rect 134 -2215 137 -2209
rect 141 -2215 144 -2209
rect 148 -2215 151 -2209
rect 155 -2215 158 -2209
rect 162 -2215 168 -2209
rect 169 -2215 175 -2209
rect 176 -2215 182 -2209
rect 183 -2215 189 -2209
rect 190 -2215 196 -2209
rect 197 -2215 200 -2209
rect 204 -2215 210 -2209
rect 211 -2215 214 -2209
rect 218 -2215 221 -2209
rect 225 -2215 228 -2209
rect 232 -2215 235 -2209
rect 239 -2215 242 -2209
rect 246 -2215 249 -2209
rect 253 -2215 256 -2209
rect 260 -2215 263 -2209
rect 267 -2215 270 -2209
rect 274 -2215 277 -2209
rect 281 -2215 284 -2209
rect 288 -2215 291 -2209
rect 295 -2215 298 -2209
rect 302 -2215 305 -2209
rect 309 -2215 312 -2209
rect 316 -2215 322 -2209
rect 323 -2215 326 -2209
rect 330 -2215 333 -2209
rect 337 -2215 343 -2209
rect 344 -2215 347 -2209
rect 351 -2215 357 -2209
rect 358 -2215 361 -2209
rect 365 -2215 368 -2209
rect 372 -2215 378 -2209
rect 379 -2215 382 -2209
rect 386 -2215 389 -2209
rect 393 -2215 399 -2209
rect 400 -2215 403 -2209
rect 407 -2215 410 -2209
rect 414 -2215 417 -2209
rect 421 -2215 424 -2209
rect 428 -2215 434 -2209
rect 435 -2215 441 -2209
rect 442 -2215 445 -2209
rect 449 -2215 452 -2209
rect 456 -2215 459 -2209
rect 463 -2215 466 -2209
rect 470 -2215 473 -2209
rect 477 -2215 480 -2209
rect 484 -2215 487 -2209
rect 491 -2215 494 -2209
rect 498 -2215 504 -2209
rect 505 -2215 511 -2209
rect 512 -2215 515 -2209
rect 519 -2215 525 -2209
rect 526 -2215 529 -2209
rect 533 -2215 536 -2209
rect 540 -2215 543 -2209
rect 547 -2215 550 -2209
rect 554 -2215 557 -2209
rect 561 -2215 567 -2209
rect 568 -2215 574 -2209
rect 575 -2215 578 -2209
rect 582 -2215 585 -2209
rect 589 -2215 595 -2209
rect 596 -2215 602 -2209
rect 603 -2215 609 -2209
rect 610 -2215 613 -2209
rect 617 -2215 620 -2209
rect 624 -2215 627 -2209
rect 631 -2215 634 -2209
rect 638 -2215 641 -2209
rect 645 -2215 648 -2209
rect 652 -2215 655 -2209
rect 659 -2215 662 -2209
rect 666 -2215 672 -2209
rect 673 -2215 676 -2209
rect 680 -2215 686 -2209
rect 687 -2215 693 -2209
rect 694 -2215 700 -2209
rect 701 -2215 704 -2209
rect 708 -2215 711 -2209
rect 715 -2215 718 -2209
rect 722 -2215 728 -2209
rect 729 -2215 732 -2209
rect 736 -2215 739 -2209
rect 743 -2215 746 -2209
rect 750 -2215 753 -2209
rect 757 -2215 760 -2209
rect 764 -2215 767 -2209
rect 771 -2215 774 -2209
rect 778 -2215 781 -2209
rect 785 -2215 788 -2209
rect 792 -2215 795 -2209
rect 799 -2215 802 -2209
rect 806 -2215 809 -2209
rect 813 -2215 816 -2209
rect 820 -2215 823 -2209
rect 827 -2215 830 -2209
rect 834 -2215 837 -2209
rect 841 -2215 844 -2209
rect 848 -2215 851 -2209
rect 855 -2215 858 -2209
rect 862 -2215 865 -2209
rect 869 -2215 875 -2209
rect 876 -2215 879 -2209
rect 883 -2215 886 -2209
rect 890 -2215 893 -2209
rect 897 -2215 900 -2209
rect 904 -2215 907 -2209
rect 911 -2215 914 -2209
rect 918 -2215 921 -2209
rect 925 -2215 928 -2209
rect 932 -2215 935 -2209
rect 939 -2215 942 -2209
rect 946 -2215 949 -2209
rect 953 -2215 956 -2209
rect 960 -2215 963 -2209
rect 967 -2215 970 -2209
rect 974 -2215 977 -2209
rect 981 -2215 984 -2209
rect 988 -2215 991 -2209
rect 995 -2215 998 -2209
rect 1002 -2215 1005 -2209
rect 1009 -2215 1012 -2209
rect 1016 -2215 1019 -2209
rect 1023 -2215 1026 -2209
rect 1030 -2215 1033 -2209
rect 1037 -2215 1040 -2209
rect 1044 -2215 1047 -2209
rect 1051 -2215 1057 -2209
rect 1 -2284 4 -2278
rect 8 -2284 11 -2278
rect 15 -2284 18 -2278
rect 22 -2284 25 -2278
rect 29 -2284 32 -2278
rect 36 -2284 39 -2278
rect 43 -2284 46 -2278
rect 50 -2284 56 -2278
rect 57 -2284 63 -2278
rect 64 -2284 67 -2278
rect 71 -2284 74 -2278
rect 78 -2284 84 -2278
rect 85 -2284 88 -2278
rect 92 -2284 95 -2278
rect 99 -2284 105 -2278
rect 106 -2284 112 -2278
rect 113 -2284 116 -2278
rect 120 -2284 123 -2278
rect 127 -2284 133 -2278
rect 134 -2284 137 -2278
rect 141 -2284 144 -2278
rect 148 -2284 151 -2278
rect 155 -2284 158 -2278
rect 162 -2284 165 -2278
rect 169 -2284 172 -2278
rect 176 -2284 182 -2278
rect 183 -2284 186 -2278
rect 190 -2284 193 -2278
rect 197 -2284 203 -2278
rect 204 -2284 207 -2278
rect 211 -2284 217 -2278
rect 218 -2284 224 -2278
rect 225 -2284 228 -2278
rect 232 -2284 235 -2278
rect 239 -2284 242 -2278
rect 246 -2284 249 -2278
rect 253 -2284 256 -2278
rect 260 -2284 263 -2278
rect 267 -2284 270 -2278
rect 274 -2284 277 -2278
rect 281 -2284 284 -2278
rect 288 -2284 294 -2278
rect 295 -2284 298 -2278
rect 302 -2284 305 -2278
rect 309 -2284 312 -2278
rect 316 -2284 319 -2278
rect 323 -2284 329 -2278
rect 330 -2284 333 -2278
rect 337 -2284 340 -2278
rect 344 -2284 350 -2278
rect 351 -2284 357 -2278
rect 358 -2284 361 -2278
rect 365 -2284 371 -2278
rect 372 -2284 375 -2278
rect 379 -2284 385 -2278
rect 386 -2284 389 -2278
rect 393 -2284 396 -2278
rect 400 -2284 403 -2278
rect 407 -2284 410 -2278
rect 414 -2284 417 -2278
rect 421 -2284 424 -2278
rect 428 -2284 431 -2278
rect 435 -2284 438 -2278
rect 442 -2284 445 -2278
rect 449 -2284 452 -2278
rect 456 -2284 459 -2278
rect 463 -2284 469 -2278
rect 470 -2284 473 -2278
rect 477 -2284 483 -2278
rect 484 -2284 490 -2278
rect 491 -2284 494 -2278
rect 498 -2284 504 -2278
rect 505 -2284 508 -2278
rect 512 -2284 515 -2278
rect 519 -2284 522 -2278
rect 526 -2284 529 -2278
rect 533 -2284 536 -2278
rect 540 -2284 546 -2278
rect 547 -2284 550 -2278
rect 554 -2284 557 -2278
rect 561 -2284 564 -2278
rect 568 -2284 571 -2278
rect 575 -2284 581 -2278
rect 582 -2284 588 -2278
rect 589 -2284 592 -2278
rect 596 -2284 599 -2278
rect 603 -2284 606 -2278
rect 610 -2284 613 -2278
rect 617 -2284 620 -2278
rect 624 -2284 627 -2278
rect 631 -2284 634 -2278
rect 638 -2284 641 -2278
rect 645 -2284 648 -2278
rect 652 -2284 655 -2278
rect 659 -2284 662 -2278
rect 666 -2284 669 -2278
rect 673 -2284 676 -2278
rect 680 -2284 686 -2278
rect 687 -2284 690 -2278
rect 694 -2284 697 -2278
rect 701 -2284 704 -2278
rect 708 -2284 711 -2278
rect 715 -2284 721 -2278
rect 722 -2284 725 -2278
rect 729 -2284 732 -2278
rect 736 -2284 739 -2278
rect 743 -2284 746 -2278
rect 750 -2284 753 -2278
rect 757 -2284 760 -2278
rect 764 -2284 770 -2278
rect 771 -2284 774 -2278
rect 778 -2284 781 -2278
rect 785 -2284 788 -2278
rect 792 -2284 795 -2278
rect 799 -2284 802 -2278
rect 806 -2284 809 -2278
rect 813 -2284 816 -2278
rect 820 -2284 823 -2278
rect 827 -2284 830 -2278
rect 834 -2284 837 -2278
rect 841 -2284 844 -2278
rect 848 -2284 851 -2278
rect 855 -2284 858 -2278
rect 862 -2284 865 -2278
rect 869 -2284 872 -2278
rect 876 -2284 879 -2278
rect 883 -2284 886 -2278
rect 890 -2284 893 -2278
rect 897 -2284 903 -2278
rect 904 -2284 910 -2278
rect 911 -2284 917 -2278
rect 918 -2284 924 -2278
rect 925 -2284 931 -2278
rect 932 -2284 935 -2278
rect 939 -2284 942 -2278
rect 946 -2284 949 -2278
rect 953 -2284 956 -2278
rect 960 -2284 963 -2278
rect 967 -2284 973 -2278
rect 974 -2284 977 -2278
rect 1 -2371 4 -2365
rect 8 -2371 14 -2365
rect 15 -2371 18 -2365
rect 22 -2371 25 -2365
rect 29 -2371 32 -2365
rect 36 -2371 39 -2365
rect 43 -2371 49 -2365
rect 50 -2371 56 -2365
rect 57 -2371 60 -2365
rect 64 -2371 67 -2365
rect 71 -2371 74 -2365
rect 78 -2371 81 -2365
rect 85 -2371 88 -2365
rect 92 -2371 98 -2365
rect 99 -2371 102 -2365
rect 106 -2371 112 -2365
rect 113 -2371 116 -2365
rect 120 -2371 123 -2365
rect 127 -2371 130 -2365
rect 134 -2371 137 -2365
rect 141 -2371 144 -2365
rect 148 -2371 151 -2365
rect 155 -2371 161 -2365
rect 162 -2371 165 -2365
rect 169 -2371 172 -2365
rect 176 -2371 179 -2365
rect 183 -2371 186 -2365
rect 190 -2371 193 -2365
rect 197 -2371 200 -2365
rect 204 -2371 207 -2365
rect 211 -2371 214 -2365
rect 218 -2371 224 -2365
rect 225 -2371 231 -2365
rect 232 -2371 235 -2365
rect 239 -2371 242 -2365
rect 246 -2371 249 -2365
rect 253 -2371 256 -2365
rect 260 -2371 263 -2365
rect 267 -2371 273 -2365
rect 274 -2371 277 -2365
rect 281 -2371 284 -2365
rect 288 -2371 291 -2365
rect 295 -2371 298 -2365
rect 302 -2371 305 -2365
rect 309 -2371 315 -2365
rect 316 -2371 319 -2365
rect 323 -2371 326 -2365
rect 330 -2371 336 -2365
rect 337 -2371 343 -2365
rect 344 -2371 347 -2365
rect 351 -2371 357 -2365
rect 358 -2371 364 -2365
rect 365 -2371 368 -2365
rect 372 -2371 378 -2365
rect 379 -2371 382 -2365
rect 386 -2371 389 -2365
rect 393 -2371 399 -2365
rect 400 -2371 406 -2365
rect 407 -2371 410 -2365
rect 414 -2371 420 -2365
rect 421 -2371 424 -2365
rect 428 -2371 431 -2365
rect 435 -2371 438 -2365
rect 442 -2371 445 -2365
rect 449 -2371 452 -2365
rect 456 -2371 462 -2365
rect 463 -2371 469 -2365
rect 470 -2371 473 -2365
rect 477 -2371 483 -2365
rect 484 -2371 487 -2365
rect 491 -2371 494 -2365
rect 498 -2371 501 -2365
rect 505 -2371 508 -2365
rect 512 -2371 515 -2365
rect 519 -2371 525 -2365
rect 526 -2371 529 -2365
rect 533 -2371 539 -2365
rect 540 -2371 543 -2365
rect 547 -2371 550 -2365
rect 554 -2371 560 -2365
rect 561 -2371 567 -2365
rect 568 -2371 571 -2365
rect 575 -2371 578 -2365
rect 582 -2371 588 -2365
rect 589 -2371 592 -2365
rect 596 -2371 599 -2365
rect 603 -2371 606 -2365
rect 610 -2371 613 -2365
rect 617 -2371 620 -2365
rect 624 -2371 627 -2365
rect 631 -2371 634 -2365
rect 638 -2371 644 -2365
rect 645 -2371 648 -2365
rect 652 -2371 655 -2365
rect 659 -2371 662 -2365
rect 666 -2371 669 -2365
rect 673 -2371 676 -2365
rect 680 -2371 683 -2365
rect 687 -2371 690 -2365
rect 694 -2371 697 -2365
rect 701 -2371 707 -2365
rect 708 -2371 711 -2365
rect 715 -2371 718 -2365
rect 722 -2371 725 -2365
rect 729 -2371 732 -2365
rect 736 -2371 739 -2365
rect 743 -2371 746 -2365
rect 750 -2371 753 -2365
rect 757 -2371 760 -2365
rect 764 -2371 767 -2365
rect 771 -2371 777 -2365
rect 778 -2371 781 -2365
rect 785 -2371 788 -2365
rect 792 -2371 795 -2365
rect 799 -2371 805 -2365
rect 806 -2371 809 -2365
rect 813 -2371 816 -2365
rect 820 -2371 823 -2365
rect 827 -2371 830 -2365
rect 834 -2371 837 -2365
rect 841 -2371 844 -2365
rect 848 -2371 851 -2365
rect 855 -2371 858 -2365
rect 862 -2371 865 -2365
rect 869 -2371 875 -2365
rect 876 -2371 879 -2365
rect 883 -2371 886 -2365
rect 890 -2371 893 -2365
rect 925 -2371 931 -2365
rect 946 -2371 949 -2365
rect 29 -2436 35 -2430
rect 57 -2436 63 -2430
rect 64 -2436 67 -2430
rect 71 -2436 77 -2430
rect 78 -2436 81 -2430
rect 85 -2436 88 -2430
rect 92 -2436 95 -2430
rect 99 -2436 102 -2430
rect 106 -2436 109 -2430
rect 113 -2436 116 -2430
rect 120 -2436 123 -2430
rect 127 -2436 130 -2430
rect 134 -2436 140 -2430
rect 141 -2436 144 -2430
rect 148 -2436 154 -2430
rect 155 -2436 161 -2430
rect 162 -2436 165 -2430
rect 169 -2436 172 -2430
rect 176 -2436 179 -2430
rect 183 -2436 189 -2430
rect 190 -2436 193 -2430
rect 197 -2436 200 -2430
rect 204 -2436 210 -2430
rect 211 -2436 217 -2430
rect 218 -2436 224 -2430
rect 225 -2436 228 -2430
rect 232 -2436 235 -2430
rect 239 -2436 242 -2430
rect 246 -2436 249 -2430
rect 253 -2436 256 -2430
rect 260 -2436 263 -2430
rect 267 -2436 270 -2430
rect 274 -2436 277 -2430
rect 281 -2436 284 -2430
rect 288 -2436 291 -2430
rect 295 -2436 301 -2430
rect 302 -2436 305 -2430
rect 309 -2436 312 -2430
rect 316 -2436 319 -2430
rect 323 -2436 326 -2430
rect 330 -2436 336 -2430
rect 337 -2436 340 -2430
rect 344 -2436 347 -2430
rect 351 -2436 354 -2430
rect 358 -2436 361 -2430
rect 365 -2436 368 -2430
rect 372 -2436 378 -2430
rect 379 -2436 382 -2430
rect 386 -2436 389 -2430
rect 393 -2436 399 -2430
rect 400 -2436 403 -2430
rect 407 -2436 413 -2430
rect 414 -2436 417 -2430
rect 421 -2436 424 -2430
rect 428 -2436 434 -2430
rect 435 -2436 438 -2430
rect 442 -2436 445 -2430
rect 449 -2436 452 -2430
rect 456 -2436 462 -2430
rect 463 -2436 469 -2430
rect 470 -2436 476 -2430
rect 477 -2436 483 -2430
rect 484 -2436 490 -2430
rect 491 -2436 494 -2430
rect 498 -2436 501 -2430
rect 505 -2436 508 -2430
rect 512 -2436 515 -2430
rect 519 -2436 522 -2430
rect 526 -2436 529 -2430
rect 533 -2436 536 -2430
rect 540 -2436 546 -2430
rect 547 -2436 553 -2430
rect 554 -2436 557 -2430
rect 561 -2436 564 -2430
rect 568 -2436 571 -2430
rect 575 -2436 581 -2430
rect 582 -2436 585 -2430
rect 589 -2436 592 -2430
rect 596 -2436 599 -2430
rect 603 -2436 606 -2430
rect 610 -2436 613 -2430
rect 617 -2436 620 -2430
rect 624 -2436 630 -2430
rect 631 -2436 634 -2430
rect 638 -2436 641 -2430
rect 645 -2436 648 -2430
rect 652 -2436 655 -2430
rect 659 -2436 662 -2430
rect 666 -2436 669 -2430
rect 673 -2436 676 -2430
rect 680 -2436 683 -2430
rect 701 -2436 704 -2430
rect 708 -2436 711 -2430
rect 715 -2436 718 -2430
rect 722 -2436 728 -2430
rect 729 -2436 735 -2430
rect 736 -2436 739 -2430
rect 743 -2436 746 -2430
rect 750 -2436 756 -2430
rect 757 -2436 763 -2430
rect 764 -2436 767 -2430
rect 771 -2436 774 -2430
rect 778 -2436 784 -2430
rect 806 -2436 809 -2430
rect 827 -2436 830 -2430
rect 883 -2436 886 -2430
rect 890 -2436 893 -2430
rect 925 -2436 928 -2430
rect 939 -2436 942 -2430
rect 1 -2477 7 -2471
rect 64 -2477 70 -2471
rect 71 -2477 74 -2471
rect 99 -2477 102 -2471
rect 106 -2477 109 -2471
rect 113 -2477 119 -2471
rect 120 -2477 123 -2471
rect 127 -2477 133 -2471
rect 134 -2477 137 -2471
rect 162 -2477 165 -2471
rect 169 -2477 172 -2471
rect 176 -2477 179 -2471
rect 183 -2477 189 -2471
rect 190 -2477 193 -2471
rect 197 -2477 200 -2471
rect 204 -2477 207 -2471
rect 218 -2477 221 -2471
rect 225 -2477 228 -2471
rect 232 -2477 238 -2471
rect 239 -2477 245 -2471
rect 246 -2477 249 -2471
rect 253 -2477 259 -2471
rect 260 -2477 266 -2471
rect 267 -2477 270 -2471
rect 274 -2477 277 -2471
rect 281 -2477 284 -2471
rect 288 -2477 291 -2471
rect 295 -2477 301 -2471
rect 302 -2477 305 -2471
rect 309 -2477 312 -2471
rect 316 -2477 319 -2471
rect 323 -2477 329 -2471
rect 330 -2477 333 -2471
rect 337 -2477 340 -2471
rect 344 -2477 350 -2471
rect 351 -2477 354 -2471
rect 358 -2477 361 -2471
rect 365 -2477 371 -2471
rect 372 -2477 378 -2471
rect 379 -2477 382 -2471
rect 386 -2477 392 -2471
rect 393 -2477 396 -2471
rect 400 -2477 403 -2471
rect 407 -2477 410 -2471
rect 414 -2477 417 -2471
rect 421 -2477 424 -2471
rect 428 -2477 434 -2471
rect 435 -2477 438 -2471
rect 442 -2477 445 -2471
rect 449 -2477 455 -2471
rect 456 -2477 459 -2471
rect 463 -2477 469 -2471
rect 470 -2477 473 -2471
rect 477 -2477 480 -2471
rect 498 -2477 504 -2471
rect 505 -2477 508 -2471
rect 512 -2477 515 -2471
rect 519 -2477 525 -2471
rect 526 -2477 532 -2471
rect 533 -2477 539 -2471
rect 540 -2477 543 -2471
rect 547 -2477 550 -2471
rect 568 -2477 571 -2471
rect 575 -2477 578 -2471
rect 582 -2477 588 -2471
rect 589 -2477 595 -2471
rect 596 -2477 602 -2471
rect 603 -2477 606 -2471
rect 610 -2477 613 -2471
rect 624 -2477 627 -2471
rect 638 -2477 644 -2471
rect 659 -2477 662 -2471
rect 673 -2477 676 -2471
rect 680 -2477 683 -2471
rect 687 -2477 690 -2471
rect 694 -2477 700 -2471
rect 708 -2477 711 -2471
rect 715 -2477 718 -2471
rect 722 -2477 725 -2471
rect 729 -2477 732 -2471
rect 736 -2477 739 -2471
rect 757 -2477 763 -2471
rect 764 -2477 767 -2471
rect 883 -2477 886 -2471
rect 890 -2477 893 -2471
rect 932 -2477 938 -2471
rect 939 -2477 942 -2471
rect 1 -2504 7 -2498
rect 85 -2504 88 -2498
rect 92 -2504 98 -2498
rect 99 -2504 105 -2498
rect 106 -2504 112 -2498
rect 113 -2504 119 -2498
rect 120 -2504 123 -2498
rect 134 -2504 140 -2498
rect 141 -2504 144 -2498
rect 148 -2504 151 -2498
rect 155 -2504 161 -2498
rect 162 -2504 168 -2498
rect 169 -2504 172 -2498
rect 176 -2504 179 -2498
rect 183 -2504 189 -2498
rect 190 -2504 196 -2498
rect 197 -2504 203 -2498
rect 204 -2504 207 -2498
rect 211 -2504 214 -2498
rect 218 -2504 224 -2498
rect 225 -2504 228 -2498
rect 232 -2504 235 -2498
rect 239 -2504 242 -2498
rect 246 -2504 249 -2498
rect 253 -2504 256 -2498
rect 260 -2504 263 -2498
rect 267 -2504 273 -2498
rect 274 -2504 277 -2498
rect 281 -2504 287 -2498
rect 288 -2504 291 -2498
rect 295 -2504 301 -2498
rect 302 -2504 308 -2498
rect 309 -2504 312 -2498
rect 316 -2504 319 -2498
rect 323 -2504 326 -2498
rect 330 -2504 333 -2498
rect 351 -2504 354 -2498
rect 358 -2504 364 -2498
rect 379 -2504 382 -2498
rect 386 -2504 392 -2498
rect 393 -2504 396 -2498
rect 400 -2504 406 -2498
rect 407 -2504 410 -2498
rect 414 -2504 420 -2498
rect 421 -2504 427 -2498
rect 442 -2504 445 -2498
rect 449 -2504 452 -2498
rect 519 -2504 525 -2498
rect 526 -2504 529 -2498
rect 603 -2504 606 -2498
rect 610 -2504 613 -2498
rect 659 -2504 662 -2498
rect 666 -2504 669 -2498
rect 680 -2504 683 -2498
rect 687 -2504 690 -2498
rect 694 -2504 697 -2498
rect 701 -2504 707 -2498
rect 708 -2504 711 -2498
rect 715 -2504 718 -2498
rect 722 -2504 725 -2498
rect 729 -2504 735 -2498
rect 736 -2504 742 -2498
rect 743 -2504 749 -2498
rect 750 -2504 753 -2498
rect 757 -2504 760 -2498
rect 883 -2504 889 -2498
rect 890 -2504 893 -2498
rect 932 -2504 935 -2498
rect 939 -2504 945 -2498
rect 946 -2504 949 -2498
rect 1 -2523 7 -2517
rect 8 -2523 11 -2517
rect 99 -2523 105 -2517
rect 106 -2523 109 -2517
rect 113 -2523 116 -2517
rect 120 -2523 126 -2517
rect 127 -2523 133 -2517
rect 155 -2523 161 -2517
rect 162 -2523 165 -2517
rect 169 -2523 175 -2517
rect 176 -2523 182 -2517
rect 183 -2523 186 -2517
rect 190 -2523 193 -2517
rect 197 -2523 203 -2517
rect 225 -2523 231 -2517
rect 267 -2523 273 -2517
rect 274 -2523 280 -2517
rect 281 -2523 287 -2517
rect 288 -2523 294 -2517
rect 295 -2523 298 -2517
rect 302 -2523 308 -2517
rect 309 -2523 312 -2517
rect 337 -2523 343 -2517
rect 344 -2523 347 -2517
rect 358 -2523 364 -2517
rect 379 -2523 385 -2517
rect 393 -2523 399 -2517
rect 400 -2523 406 -2517
rect 449 -2523 452 -2517
rect 456 -2523 462 -2517
rect 519 -2523 525 -2517
rect 596 -2523 602 -2517
rect 603 -2523 606 -2517
rect 659 -2523 665 -2517
rect 666 -2523 669 -2517
rect 687 -2523 693 -2517
rect 708 -2523 714 -2517
rect 715 -2523 718 -2517
rect 722 -2523 728 -2517
rect 729 -2523 732 -2517
rect 736 -2523 742 -2517
<< polysilicon >>
rect 86 -11 87 -9
rect 89 -11 90 -9
rect 93 -5 94 -3
rect 93 -11 94 -9
rect 100 -5 101 -3
rect 100 -11 101 -9
rect 107 -5 108 -3
rect 107 -11 108 -9
rect 117 -5 118 -3
rect 121 -5 122 -3
rect 121 -11 122 -9
rect 128 -5 129 -3
rect 128 -11 129 -9
rect 145 -11 146 -9
rect 205 -5 206 -3
rect 205 -11 206 -9
rect 212 -5 213 -3
rect 215 -5 216 -3
rect 219 -11 220 -9
rect 222 -11 223 -9
rect 226 -5 227 -3
rect 226 -11 227 -9
rect 233 -5 234 -3
rect 236 -5 237 -3
rect 240 -5 241 -3
rect 240 -11 241 -9
rect 247 -5 248 -3
rect 250 -11 251 -9
rect 257 -11 258 -9
rect 261 -5 262 -3
rect 268 -5 269 -3
rect 268 -11 269 -9
rect 282 -11 283 -9
rect 324 -5 325 -3
rect 324 -11 325 -9
rect 334 -5 335 -3
rect 341 -11 342 -9
rect 429 -5 430 -3
rect 429 -11 430 -9
rect 450 -5 451 -3
rect 450 -11 451 -9
rect 464 -5 465 -3
rect 464 -11 465 -9
rect 488 -5 489 -3
rect 485 -11 486 -9
rect 509 -11 510 -9
rect 530 -5 531 -3
rect 534 -5 535 -3
rect 534 -11 535 -9
rect 548 -11 549 -9
rect 583 -5 584 -3
rect 590 -11 591 -9
rect 597 -5 598 -3
rect 597 -11 598 -9
rect 607 -11 608 -9
rect 660 -5 661 -3
rect 667 -5 668 -3
rect 667 -11 668 -9
rect 100 -24 101 -22
rect 103 -24 104 -22
rect 100 -30 101 -28
rect 103 -30 104 -28
rect 117 -24 118 -22
rect 135 -24 136 -22
rect 135 -30 136 -28
rect 173 -24 174 -22
rect 177 -24 178 -22
rect 177 -30 178 -28
rect 184 -24 185 -22
rect 184 -30 185 -28
rect 194 -30 195 -28
rect 198 -24 199 -22
rect 198 -30 199 -28
rect 205 -24 206 -22
rect 212 -24 213 -22
rect 215 -24 216 -22
rect 212 -30 213 -28
rect 219 -24 220 -22
rect 219 -30 220 -28
rect 226 -24 227 -22
rect 226 -30 227 -28
rect 233 -24 234 -22
rect 236 -24 237 -22
rect 240 -24 241 -22
rect 247 -24 248 -22
rect 247 -30 248 -28
rect 254 -24 255 -22
rect 254 -30 255 -28
rect 261 -24 262 -22
rect 261 -30 262 -28
rect 268 -24 269 -22
rect 268 -30 269 -28
rect 275 -24 276 -22
rect 275 -30 276 -28
rect 282 -24 283 -22
rect 282 -30 283 -28
rect 289 -24 290 -22
rect 289 -30 290 -28
rect 296 -30 297 -28
rect 303 -24 304 -22
rect 306 -24 307 -22
rect 310 -24 311 -22
rect 310 -30 311 -28
rect 317 -24 318 -22
rect 317 -30 318 -28
rect 324 -24 325 -22
rect 324 -30 325 -28
rect 331 -24 332 -22
rect 338 -30 339 -28
rect 348 -24 349 -22
rect 348 -30 349 -28
rect 359 -24 360 -22
rect 359 -30 360 -28
rect 373 -24 374 -22
rect 373 -30 374 -28
rect 383 -30 384 -28
rect 415 -24 416 -22
rect 415 -30 416 -28
rect 422 -30 423 -28
rect 429 -24 430 -22
rect 429 -30 430 -28
rect 439 -24 440 -22
rect 446 -24 447 -22
rect 446 -30 447 -28
rect 453 -24 454 -22
rect 464 -30 465 -28
rect 467 -30 468 -28
rect 471 -24 472 -22
rect 471 -30 472 -28
rect 492 -24 493 -22
rect 492 -30 493 -28
rect 506 -24 507 -22
rect 506 -30 507 -28
rect 513 -24 514 -22
rect 513 -30 514 -28
rect 520 -30 521 -28
rect 527 -24 528 -22
rect 527 -30 528 -28
rect 541 -24 542 -22
rect 541 -30 542 -28
rect 555 -30 556 -28
rect 562 -24 563 -22
rect 569 -24 570 -22
rect 569 -30 570 -28
rect 576 -24 577 -22
rect 576 -30 577 -28
rect 604 -24 605 -22
rect 604 -30 605 -28
rect 611 -24 612 -22
rect 611 -30 612 -28
rect 618 -24 619 -22
rect 618 -30 619 -28
rect 674 -24 675 -22
rect 674 -30 675 -28
rect 86 -55 87 -53
rect 86 -61 87 -59
rect 93 -55 94 -53
rect 93 -61 94 -59
rect 114 -55 115 -53
rect 114 -61 115 -59
rect 121 -55 122 -53
rect 121 -61 122 -59
rect 128 -55 129 -53
rect 128 -61 129 -59
rect 135 -55 136 -53
rect 135 -61 136 -59
rect 145 -55 146 -53
rect 149 -61 150 -59
rect 156 -55 157 -53
rect 156 -61 157 -59
rect 163 -55 164 -53
rect 163 -61 164 -59
rect 173 -55 174 -53
rect 170 -61 171 -59
rect 173 -61 174 -59
rect 177 -55 178 -53
rect 177 -61 178 -59
rect 187 -55 188 -53
rect 184 -61 185 -59
rect 191 -55 192 -53
rect 191 -61 192 -59
rect 198 -55 199 -53
rect 201 -55 202 -53
rect 205 -55 206 -53
rect 205 -61 206 -59
rect 212 -55 213 -53
rect 212 -61 213 -59
rect 219 -55 220 -53
rect 219 -61 220 -59
rect 226 -55 227 -53
rect 226 -61 227 -59
rect 236 -55 237 -53
rect 233 -61 234 -59
rect 240 -61 241 -59
rect 243 -61 244 -59
rect 247 -55 248 -53
rect 250 -55 251 -53
rect 250 -61 251 -59
rect 254 -55 255 -53
rect 254 -61 255 -59
rect 261 -55 262 -53
rect 261 -61 262 -59
rect 268 -55 269 -53
rect 268 -61 269 -59
rect 275 -55 276 -53
rect 275 -61 276 -59
rect 282 -55 283 -53
rect 282 -61 283 -59
rect 289 -55 290 -53
rect 289 -61 290 -59
rect 299 -55 300 -53
rect 296 -61 297 -59
rect 303 -55 304 -53
rect 303 -61 304 -59
rect 313 -55 314 -53
rect 310 -61 311 -59
rect 317 -55 318 -53
rect 317 -61 318 -59
rect 324 -55 325 -53
rect 324 -61 325 -59
rect 331 -55 332 -53
rect 331 -61 332 -59
rect 338 -55 339 -53
rect 341 -55 342 -53
rect 341 -61 342 -59
rect 345 -55 346 -53
rect 345 -61 346 -59
rect 352 -55 353 -53
rect 352 -61 353 -59
rect 359 -61 360 -59
rect 366 -55 367 -53
rect 366 -61 367 -59
rect 373 -55 374 -53
rect 373 -61 374 -59
rect 383 -55 384 -53
rect 380 -61 381 -59
rect 387 -55 388 -53
rect 387 -61 388 -59
rect 394 -55 395 -53
rect 394 -61 395 -59
rect 401 -55 402 -53
rect 401 -61 402 -59
rect 408 -55 409 -53
rect 408 -61 409 -59
rect 418 -61 419 -59
rect 422 -55 423 -53
rect 422 -61 423 -59
rect 429 -55 430 -53
rect 429 -61 430 -59
rect 436 -55 437 -53
rect 436 -61 437 -59
rect 443 -55 444 -53
rect 443 -61 444 -59
rect 464 -55 465 -53
rect 467 -61 468 -59
rect 471 -55 472 -53
rect 471 -61 472 -59
rect 478 -55 479 -53
rect 478 -61 479 -59
rect 485 -55 486 -53
rect 485 -61 486 -59
rect 492 -61 493 -59
rect 495 -61 496 -59
rect 499 -55 500 -53
rect 499 -61 500 -59
rect 506 -55 507 -53
rect 506 -61 507 -59
rect 520 -55 521 -53
rect 520 -61 521 -59
rect 527 -55 528 -53
rect 530 -61 531 -59
rect 534 -55 535 -53
rect 534 -61 535 -59
rect 541 -55 542 -53
rect 541 -61 542 -59
rect 551 -55 552 -53
rect 548 -61 549 -59
rect 555 -55 556 -53
rect 555 -61 556 -59
rect 562 -55 563 -53
rect 562 -61 563 -59
rect 569 -55 570 -53
rect 569 -61 570 -59
rect 576 -55 577 -53
rect 576 -61 577 -59
rect 586 -55 587 -53
rect 583 -61 584 -59
rect 586 -61 587 -59
rect 590 -55 591 -53
rect 590 -61 591 -59
rect 597 -55 598 -53
rect 597 -61 598 -59
rect 604 -55 605 -53
rect 604 -61 605 -59
rect 611 -55 612 -53
rect 611 -61 612 -59
rect 625 -55 626 -53
rect 625 -61 626 -59
rect 632 -55 633 -53
rect 632 -61 633 -59
rect 639 -55 640 -53
rect 639 -61 640 -59
rect 646 -55 647 -53
rect 646 -61 647 -59
rect 653 -55 654 -53
rect 653 -61 654 -59
rect 663 -55 664 -53
rect 660 -61 661 -59
rect 667 -55 668 -53
rect 667 -61 668 -59
rect 677 -55 678 -53
rect 681 -55 682 -53
rect 681 -61 682 -59
rect 702 -55 703 -53
rect 702 -61 703 -59
rect 765 -55 766 -53
rect 765 -61 766 -59
rect 772 -55 773 -53
rect 772 -61 773 -59
rect 842 -55 843 -53
rect 842 -61 843 -59
rect 30 -124 31 -122
rect 30 -130 31 -128
rect 37 -124 38 -122
rect 37 -130 38 -128
rect 47 -124 48 -122
rect 51 -124 52 -122
rect 51 -130 52 -128
rect 58 -124 59 -122
rect 61 -124 62 -122
rect 58 -130 59 -128
rect 65 -124 66 -122
rect 65 -130 66 -128
rect 72 -124 73 -122
rect 72 -130 73 -128
rect 79 -124 80 -122
rect 79 -130 80 -128
rect 86 -124 87 -122
rect 86 -130 87 -128
rect 93 -124 94 -122
rect 93 -130 94 -128
rect 100 -124 101 -122
rect 103 -124 104 -122
rect 107 -124 108 -122
rect 107 -130 108 -128
rect 117 -124 118 -122
rect 114 -130 115 -128
rect 117 -130 118 -128
rect 121 -124 122 -122
rect 121 -130 122 -128
rect 128 -124 129 -122
rect 128 -130 129 -128
rect 135 -124 136 -122
rect 135 -130 136 -128
rect 142 -124 143 -122
rect 142 -130 143 -128
rect 152 -124 153 -122
rect 149 -130 150 -128
rect 152 -130 153 -128
rect 156 -124 157 -122
rect 159 -124 160 -122
rect 156 -130 157 -128
rect 159 -130 160 -128
rect 163 -124 164 -122
rect 163 -130 164 -128
rect 173 -124 174 -122
rect 170 -130 171 -128
rect 173 -130 174 -128
rect 177 -124 178 -122
rect 177 -130 178 -128
rect 184 -124 185 -122
rect 184 -130 185 -128
rect 191 -124 192 -122
rect 191 -130 192 -128
rect 198 -124 199 -122
rect 198 -130 199 -128
rect 205 -124 206 -122
rect 205 -130 206 -128
rect 212 -124 213 -122
rect 212 -130 213 -128
rect 219 -124 220 -122
rect 219 -130 220 -128
rect 226 -124 227 -122
rect 229 -124 230 -122
rect 226 -130 227 -128
rect 229 -130 230 -128
rect 233 -124 234 -122
rect 233 -130 234 -128
rect 240 -124 241 -122
rect 240 -130 241 -128
rect 247 -124 248 -122
rect 254 -124 255 -122
rect 254 -130 255 -128
rect 261 -124 262 -122
rect 261 -130 262 -128
rect 268 -124 269 -122
rect 268 -130 269 -128
rect 275 -124 276 -122
rect 278 -124 279 -122
rect 275 -130 276 -128
rect 282 -124 283 -122
rect 282 -130 283 -128
rect 289 -124 290 -122
rect 289 -130 290 -128
rect 296 -124 297 -122
rect 296 -130 297 -128
rect 303 -124 304 -122
rect 303 -130 304 -128
rect 310 -124 311 -122
rect 310 -130 311 -128
rect 317 -124 318 -122
rect 320 -124 321 -122
rect 317 -130 318 -128
rect 320 -130 321 -128
rect 324 -124 325 -122
rect 324 -130 325 -128
rect 331 -124 332 -122
rect 331 -130 332 -128
rect 338 -124 339 -122
rect 338 -130 339 -128
rect 345 -130 346 -128
rect 348 -130 349 -128
rect 355 -124 356 -122
rect 352 -130 353 -128
rect 355 -130 356 -128
rect 359 -124 360 -122
rect 359 -130 360 -128
rect 366 -124 367 -122
rect 366 -130 367 -128
rect 376 -124 377 -122
rect 376 -130 377 -128
rect 380 -124 381 -122
rect 380 -130 381 -128
rect 387 -124 388 -122
rect 390 -124 391 -122
rect 397 -124 398 -122
rect 394 -130 395 -128
rect 397 -130 398 -128
rect 401 -124 402 -122
rect 401 -130 402 -128
rect 408 -124 409 -122
rect 408 -130 409 -128
rect 415 -124 416 -122
rect 418 -130 419 -128
rect 422 -124 423 -122
rect 422 -130 423 -128
rect 429 -124 430 -122
rect 429 -130 430 -128
rect 436 -124 437 -122
rect 436 -130 437 -128
rect 443 -124 444 -122
rect 443 -130 444 -128
rect 450 -124 451 -122
rect 450 -130 451 -128
rect 457 -124 458 -122
rect 457 -130 458 -128
rect 464 -124 465 -122
rect 464 -130 465 -128
rect 471 -124 472 -122
rect 471 -130 472 -128
rect 478 -124 479 -122
rect 478 -130 479 -128
rect 485 -124 486 -122
rect 485 -130 486 -128
rect 492 -124 493 -122
rect 492 -130 493 -128
rect 499 -124 500 -122
rect 502 -124 503 -122
rect 499 -130 500 -128
rect 509 -124 510 -122
rect 506 -130 507 -128
rect 509 -130 510 -128
rect 513 -124 514 -122
rect 513 -130 514 -128
rect 520 -124 521 -122
rect 520 -130 521 -128
rect 527 -124 528 -122
rect 527 -130 528 -128
rect 534 -124 535 -122
rect 534 -130 535 -128
rect 541 -124 542 -122
rect 541 -130 542 -128
rect 548 -124 549 -122
rect 548 -130 549 -128
rect 555 -124 556 -122
rect 555 -130 556 -128
rect 562 -124 563 -122
rect 562 -130 563 -128
rect 569 -124 570 -122
rect 569 -130 570 -128
rect 576 -124 577 -122
rect 576 -130 577 -128
rect 586 -124 587 -122
rect 583 -130 584 -128
rect 590 -124 591 -122
rect 590 -130 591 -128
rect 597 -124 598 -122
rect 597 -130 598 -128
rect 604 -124 605 -122
rect 604 -130 605 -128
rect 611 -124 612 -122
rect 611 -130 612 -128
rect 618 -124 619 -122
rect 618 -130 619 -128
rect 625 -124 626 -122
rect 625 -130 626 -128
rect 632 -124 633 -122
rect 632 -130 633 -128
rect 639 -124 640 -122
rect 639 -130 640 -128
rect 646 -124 647 -122
rect 646 -130 647 -128
rect 653 -124 654 -122
rect 653 -130 654 -128
rect 660 -130 661 -128
rect 667 -124 668 -122
rect 667 -130 668 -128
rect 674 -124 675 -122
rect 674 -130 675 -128
rect 681 -124 682 -122
rect 681 -130 682 -128
rect 688 -124 689 -122
rect 688 -130 689 -128
rect 695 -124 696 -122
rect 695 -130 696 -128
rect 702 -124 703 -122
rect 702 -130 703 -128
rect 709 -124 710 -122
rect 709 -130 710 -128
rect 716 -124 717 -122
rect 716 -130 717 -128
rect 723 -124 724 -122
rect 723 -130 724 -128
rect 730 -124 731 -122
rect 730 -130 731 -128
rect 737 -124 738 -122
rect 737 -130 738 -128
rect 744 -124 745 -122
rect 744 -130 745 -128
rect 751 -124 752 -122
rect 751 -130 752 -128
rect 758 -124 759 -122
rect 758 -130 759 -128
rect 765 -124 766 -122
rect 765 -130 766 -128
rect 772 -124 773 -122
rect 772 -130 773 -128
rect 779 -124 780 -122
rect 779 -130 780 -128
rect 786 -124 787 -122
rect 786 -130 787 -128
rect 793 -124 794 -122
rect 793 -130 794 -128
rect 800 -124 801 -122
rect 800 -130 801 -128
rect 807 -124 808 -122
rect 807 -130 808 -128
rect 814 -124 815 -122
rect 814 -130 815 -128
rect 821 -124 822 -122
rect 821 -130 822 -128
rect 828 -124 829 -122
rect 828 -130 829 -128
rect 835 -124 836 -122
rect 835 -130 836 -128
rect 842 -124 843 -122
rect 842 -130 843 -128
rect 870 -124 871 -122
rect 870 -130 871 -128
rect 877 -124 878 -122
rect 877 -130 878 -128
rect 1108 -130 1109 -128
rect 23 -213 24 -211
rect 23 -219 24 -217
rect 30 -213 31 -211
rect 30 -219 31 -217
rect 37 -213 38 -211
rect 37 -219 38 -217
rect 44 -213 45 -211
rect 44 -219 45 -217
rect 51 -213 52 -211
rect 51 -219 52 -217
rect 58 -213 59 -211
rect 58 -219 59 -217
rect 65 -213 66 -211
rect 65 -219 66 -217
rect 72 -213 73 -211
rect 72 -219 73 -217
rect 79 -213 80 -211
rect 79 -219 80 -217
rect 89 -213 90 -211
rect 93 -213 94 -211
rect 93 -219 94 -217
rect 100 -213 101 -211
rect 100 -219 101 -217
rect 110 -213 111 -211
rect 114 -213 115 -211
rect 114 -219 115 -217
rect 124 -213 125 -211
rect 121 -219 122 -217
rect 128 -213 129 -211
rect 128 -219 129 -217
rect 135 -213 136 -211
rect 135 -219 136 -217
rect 142 -213 143 -211
rect 145 -213 146 -211
rect 142 -219 143 -217
rect 152 -213 153 -211
rect 149 -219 150 -217
rect 152 -219 153 -217
rect 156 -213 157 -211
rect 156 -219 157 -217
rect 163 -213 164 -211
rect 163 -219 164 -217
rect 170 -213 171 -211
rect 170 -219 171 -217
rect 180 -213 181 -211
rect 177 -219 178 -217
rect 184 -213 185 -211
rect 184 -219 185 -217
rect 191 -213 192 -211
rect 191 -219 192 -217
rect 198 -213 199 -211
rect 198 -219 199 -217
rect 205 -213 206 -211
rect 208 -213 209 -211
rect 205 -219 206 -217
rect 208 -219 209 -217
rect 212 -213 213 -211
rect 215 -213 216 -211
rect 212 -219 213 -217
rect 219 -213 220 -211
rect 219 -219 220 -217
rect 222 -219 223 -217
rect 229 -219 230 -217
rect 233 -213 234 -211
rect 240 -213 241 -211
rect 240 -219 241 -217
rect 250 -213 251 -211
rect 247 -219 248 -217
rect 254 -213 255 -211
rect 254 -219 255 -217
rect 261 -213 262 -211
rect 261 -219 262 -217
rect 268 -213 269 -211
rect 268 -219 269 -217
rect 275 -213 276 -211
rect 275 -219 276 -217
rect 282 -213 283 -211
rect 282 -219 283 -217
rect 289 -213 290 -211
rect 289 -219 290 -217
rect 296 -213 297 -211
rect 299 -213 300 -211
rect 299 -219 300 -217
rect 303 -213 304 -211
rect 303 -219 304 -217
rect 310 -213 311 -211
rect 310 -219 311 -217
rect 317 -213 318 -211
rect 317 -219 318 -217
rect 324 -213 325 -211
rect 327 -213 328 -211
rect 324 -219 325 -217
rect 334 -213 335 -211
rect 331 -219 332 -217
rect 334 -219 335 -217
rect 338 -213 339 -211
rect 338 -219 339 -217
rect 345 -213 346 -211
rect 348 -213 349 -211
rect 352 -213 353 -211
rect 352 -219 353 -217
rect 359 -213 360 -211
rect 362 -213 363 -211
rect 359 -219 360 -217
rect 362 -219 363 -217
rect 366 -213 367 -211
rect 366 -219 367 -217
rect 373 -213 374 -211
rect 373 -219 374 -217
rect 380 -213 381 -211
rect 380 -219 381 -217
rect 387 -213 388 -211
rect 387 -219 388 -217
rect 394 -213 395 -211
rect 397 -219 398 -217
rect 401 -213 402 -211
rect 401 -219 402 -217
rect 404 -219 405 -217
rect 408 -213 409 -211
rect 408 -219 409 -217
rect 415 -213 416 -211
rect 415 -219 416 -217
rect 422 -213 423 -211
rect 422 -219 423 -217
rect 429 -213 430 -211
rect 429 -219 430 -217
rect 436 -213 437 -211
rect 436 -219 437 -217
rect 443 -213 444 -211
rect 443 -219 444 -217
rect 450 -213 451 -211
rect 450 -219 451 -217
rect 457 -219 458 -217
rect 464 -213 465 -211
rect 464 -219 465 -217
rect 471 -213 472 -211
rect 471 -219 472 -217
rect 478 -213 479 -211
rect 478 -219 479 -217
rect 485 -213 486 -211
rect 485 -219 486 -217
rect 492 -213 493 -211
rect 495 -213 496 -211
rect 495 -219 496 -217
rect 499 -213 500 -211
rect 499 -219 500 -217
rect 506 -213 507 -211
rect 506 -219 507 -217
rect 513 -213 514 -211
rect 513 -219 514 -217
rect 520 -213 521 -211
rect 523 -213 524 -211
rect 520 -219 521 -217
rect 527 -213 528 -211
rect 527 -219 528 -217
rect 534 -213 535 -211
rect 534 -219 535 -217
rect 541 -213 542 -211
rect 541 -219 542 -217
rect 548 -213 549 -211
rect 548 -219 549 -217
rect 555 -213 556 -211
rect 555 -219 556 -217
rect 562 -213 563 -211
rect 562 -219 563 -217
rect 569 -213 570 -211
rect 569 -219 570 -217
rect 576 -213 577 -211
rect 579 -213 580 -211
rect 576 -219 577 -217
rect 579 -219 580 -217
rect 583 -213 584 -211
rect 583 -219 584 -217
rect 590 -213 591 -211
rect 590 -219 591 -217
rect 597 -213 598 -211
rect 597 -219 598 -217
rect 604 -213 605 -211
rect 604 -219 605 -217
rect 611 -213 612 -211
rect 611 -219 612 -217
rect 618 -213 619 -211
rect 618 -219 619 -217
rect 621 -219 622 -217
rect 625 -213 626 -211
rect 628 -219 629 -217
rect 632 -213 633 -211
rect 632 -219 633 -217
rect 639 -213 640 -211
rect 639 -219 640 -217
rect 646 -213 647 -211
rect 646 -219 647 -217
rect 653 -213 654 -211
rect 656 -213 657 -211
rect 653 -219 654 -217
rect 660 -213 661 -211
rect 660 -219 661 -217
rect 667 -213 668 -211
rect 667 -219 668 -217
rect 674 -213 675 -211
rect 674 -219 675 -217
rect 681 -213 682 -211
rect 681 -219 682 -217
rect 688 -213 689 -211
rect 688 -219 689 -217
rect 695 -213 696 -211
rect 695 -219 696 -217
rect 702 -213 703 -211
rect 702 -219 703 -217
rect 709 -213 710 -211
rect 709 -219 710 -217
rect 716 -213 717 -211
rect 716 -219 717 -217
rect 723 -213 724 -211
rect 723 -219 724 -217
rect 730 -213 731 -211
rect 730 -219 731 -217
rect 737 -213 738 -211
rect 740 -219 741 -217
rect 744 -213 745 -211
rect 744 -219 745 -217
rect 751 -213 752 -211
rect 751 -219 752 -217
rect 758 -213 759 -211
rect 758 -219 759 -217
rect 765 -213 766 -211
rect 765 -219 766 -217
rect 772 -213 773 -211
rect 772 -219 773 -217
rect 779 -213 780 -211
rect 779 -219 780 -217
rect 786 -213 787 -211
rect 786 -219 787 -217
rect 793 -213 794 -211
rect 793 -219 794 -217
rect 800 -213 801 -211
rect 800 -219 801 -217
rect 807 -213 808 -211
rect 807 -219 808 -217
rect 814 -213 815 -211
rect 814 -219 815 -217
rect 821 -213 822 -211
rect 821 -219 822 -217
rect 828 -213 829 -211
rect 828 -219 829 -217
rect 835 -213 836 -211
rect 835 -219 836 -217
rect 842 -213 843 -211
rect 842 -219 843 -217
rect 849 -213 850 -211
rect 849 -219 850 -217
rect 856 -213 857 -211
rect 856 -219 857 -217
rect 863 -213 864 -211
rect 863 -219 864 -217
rect 870 -213 871 -211
rect 870 -219 871 -217
rect 877 -213 878 -211
rect 877 -219 878 -217
rect 884 -213 885 -211
rect 884 -219 885 -217
rect 891 -213 892 -211
rect 891 -219 892 -217
rect 898 -213 899 -211
rect 898 -219 899 -217
rect 905 -213 906 -211
rect 905 -219 906 -217
rect 912 -213 913 -211
rect 912 -219 913 -217
rect 919 -213 920 -211
rect 919 -219 920 -217
rect 926 -213 927 -211
rect 926 -219 927 -217
rect 933 -213 934 -211
rect 933 -219 934 -217
rect 940 -213 941 -211
rect 940 -219 941 -217
rect 947 -213 948 -211
rect 947 -219 948 -217
rect 954 -213 955 -211
rect 954 -219 955 -217
rect 1108 -213 1109 -211
rect 1108 -219 1109 -217
rect 16 -296 17 -294
rect 16 -302 17 -300
rect 23 -296 24 -294
rect 23 -302 24 -300
rect 30 -296 31 -294
rect 30 -302 31 -300
rect 37 -296 38 -294
rect 37 -302 38 -300
rect 47 -296 48 -294
rect 47 -302 48 -300
rect 51 -296 52 -294
rect 51 -302 52 -300
rect 58 -296 59 -294
rect 58 -302 59 -300
rect 65 -296 66 -294
rect 68 -296 69 -294
rect 65 -302 66 -300
rect 68 -302 69 -300
rect 72 -296 73 -294
rect 72 -302 73 -300
rect 79 -296 80 -294
rect 79 -302 80 -300
rect 86 -296 87 -294
rect 86 -302 87 -300
rect 93 -296 94 -294
rect 93 -302 94 -300
rect 100 -296 101 -294
rect 100 -302 101 -300
rect 103 -302 104 -300
rect 107 -296 108 -294
rect 107 -302 108 -300
rect 114 -296 115 -294
rect 117 -296 118 -294
rect 117 -302 118 -300
rect 121 -296 122 -294
rect 121 -302 122 -300
rect 128 -302 129 -300
rect 131 -302 132 -300
rect 135 -296 136 -294
rect 138 -296 139 -294
rect 135 -302 136 -300
rect 142 -296 143 -294
rect 142 -302 143 -300
rect 149 -296 150 -294
rect 149 -302 150 -300
rect 156 -296 157 -294
rect 156 -302 157 -300
rect 166 -296 167 -294
rect 163 -302 164 -300
rect 166 -302 167 -300
rect 170 -296 171 -294
rect 173 -296 174 -294
rect 170 -302 171 -300
rect 173 -302 174 -300
rect 177 -296 178 -294
rect 177 -302 178 -300
rect 184 -296 185 -294
rect 184 -302 185 -300
rect 191 -296 192 -294
rect 194 -296 195 -294
rect 191 -302 192 -300
rect 194 -302 195 -300
rect 198 -296 199 -294
rect 198 -302 199 -300
rect 205 -296 206 -294
rect 205 -302 206 -300
rect 208 -302 209 -300
rect 212 -296 213 -294
rect 212 -302 213 -300
rect 219 -296 220 -294
rect 219 -302 220 -300
rect 226 -296 227 -294
rect 226 -302 227 -300
rect 233 -296 234 -294
rect 233 -302 234 -300
rect 240 -296 241 -294
rect 240 -302 241 -300
rect 247 -296 248 -294
rect 247 -302 248 -300
rect 254 -296 255 -294
rect 257 -296 258 -294
rect 261 -296 262 -294
rect 261 -302 262 -300
rect 268 -296 269 -294
rect 268 -302 269 -300
rect 275 -296 276 -294
rect 275 -302 276 -300
rect 282 -296 283 -294
rect 282 -302 283 -300
rect 289 -296 290 -294
rect 289 -302 290 -300
rect 296 -296 297 -294
rect 299 -296 300 -294
rect 296 -302 297 -300
rect 299 -302 300 -300
rect 303 -296 304 -294
rect 303 -302 304 -300
rect 310 -296 311 -294
rect 310 -302 311 -300
rect 317 -296 318 -294
rect 320 -302 321 -300
rect 324 -296 325 -294
rect 324 -302 325 -300
rect 331 -296 332 -294
rect 331 -302 332 -300
rect 338 -296 339 -294
rect 338 -302 339 -300
rect 345 -296 346 -294
rect 345 -302 346 -300
rect 355 -296 356 -294
rect 352 -302 353 -300
rect 355 -302 356 -300
rect 362 -296 363 -294
rect 359 -302 360 -300
rect 366 -296 367 -294
rect 366 -302 367 -300
rect 373 -296 374 -294
rect 373 -302 374 -300
rect 380 -296 381 -294
rect 380 -302 381 -300
rect 387 -296 388 -294
rect 387 -302 388 -300
rect 394 -296 395 -294
rect 397 -302 398 -300
rect 401 -296 402 -294
rect 401 -302 402 -300
rect 404 -302 405 -300
rect 408 -296 409 -294
rect 408 -302 409 -300
rect 415 -296 416 -294
rect 415 -302 416 -300
rect 422 -296 423 -294
rect 422 -302 423 -300
rect 429 -296 430 -294
rect 429 -302 430 -300
rect 436 -296 437 -294
rect 436 -302 437 -300
rect 439 -302 440 -300
rect 443 -296 444 -294
rect 443 -302 444 -300
rect 450 -296 451 -294
rect 450 -302 451 -300
rect 457 -296 458 -294
rect 457 -302 458 -300
rect 467 -296 468 -294
rect 464 -302 465 -300
rect 467 -302 468 -300
rect 471 -296 472 -294
rect 471 -302 472 -300
rect 478 -296 479 -294
rect 478 -302 479 -300
rect 485 -296 486 -294
rect 488 -296 489 -294
rect 485 -302 486 -300
rect 488 -302 489 -300
rect 492 -296 493 -294
rect 492 -302 493 -300
rect 499 -296 500 -294
rect 502 -296 503 -294
rect 506 -296 507 -294
rect 506 -302 507 -300
rect 513 -296 514 -294
rect 513 -302 514 -300
rect 520 -296 521 -294
rect 523 -302 524 -300
rect 527 -296 528 -294
rect 527 -302 528 -300
rect 534 -296 535 -294
rect 534 -302 535 -300
rect 541 -296 542 -294
rect 541 -302 542 -300
rect 548 -296 549 -294
rect 548 -302 549 -300
rect 555 -296 556 -294
rect 555 -302 556 -300
rect 562 -296 563 -294
rect 562 -302 563 -300
rect 569 -296 570 -294
rect 569 -302 570 -300
rect 576 -296 577 -294
rect 576 -302 577 -300
rect 583 -296 584 -294
rect 583 -302 584 -300
rect 590 -296 591 -294
rect 590 -302 591 -300
rect 597 -296 598 -294
rect 597 -302 598 -300
rect 604 -296 605 -294
rect 604 -302 605 -300
rect 611 -296 612 -294
rect 611 -302 612 -300
rect 618 -296 619 -294
rect 618 -302 619 -300
rect 625 -296 626 -294
rect 625 -302 626 -300
rect 632 -296 633 -294
rect 632 -302 633 -300
rect 639 -296 640 -294
rect 639 -302 640 -300
rect 646 -296 647 -294
rect 646 -302 647 -300
rect 653 -296 654 -294
rect 653 -302 654 -300
rect 663 -296 664 -294
rect 667 -296 668 -294
rect 667 -302 668 -300
rect 674 -296 675 -294
rect 674 -302 675 -300
rect 681 -296 682 -294
rect 681 -302 682 -300
rect 688 -296 689 -294
rect 688 -302 689 -300
rect 695 -296 696 -294
rect 695 -302 696 -300
rect 702 -296 703 -294
rect 702 -302 703 -300
rect 709 -296 710 -294
rect 709 -302 710 -300
rect 716 -296 717 -294
rect 716 -302 717 -300
rect 723 -296 724 -294
rect 723 -302 724 -300
rect 730 -296 731 -294
rect 730 -302 731 -300
rect 737 -296 738 -294
rect 737 -302 738 -300
rect 744 -296 745 -294
rect 744 -302 745 -300
rect 751 -296 752 -294
rect 751 -302 752 -300
rect 758 -296 759 -294
rect 758 -302 759 -300
rect 765 -296 766 -294
rect 765 -302 766 -300
rect 772 -296 773 -294
rect 772 -302 773 -300
rect 779 -296 780 -294
rect 779 -302 780 -300
rect 786 -296 787 -294
rect 786 -302 787 -300
rect 793 -296 794 -294
rect 793 -302 794 -300
rect 800 -296 801 -294
rect 800 -302 801 -300
rect 807 -296 808 -294
rect 807 -302 808 -300
rect 814 -296 815 -294
rect 814 -302 815 -300
rect 821 -296 822 -294
rect 821 -302 822 -300
rect 828 -296 829 -294
rect 828 -302 829 -300
rect 835 -296 836 -294
rect 835 -302 836 -300
rect 842 -296 843 -294
rect 842 -302 843 -300
rect 849 -296 850 -294
rect 849 -302 850 -300
rect 856 -296 857 -294
rect 856 -302 857 -300
rect 863 -296 864 -294
rect 863 -302 864 -300
rect 870 -296 871 -294
rect 870 -302 871 -300
rect 877 -296 878 -294
rect 877 -302 878 -300
rect 887 -296 888 -294
rect 884 -302 885 -300
rect 894 -302 895 -300
rect 898 -296 899 -294
rect 905 -296 906 -294
rect 908 -296 909 -294
rect 912 -296 913 -294
rect 912 -302 913 -300
rect 919 -296 920 -294
rect 919 -302 920 -300
rect 1108 -296 1109 -294
rect 1108 -302 1109 -300
rect 9 -391 10 -389
rect 9 -397 10 -395
rect 16 -391 17 -389
rect 23 -391 24 -389
rect 23 -397 24 -395
rect 30 -397 31 -395
rect 37 -391 38 -389
rect 37 -397 38 -395
rect 44 -391 45 -389
rect 44 -397 45 -395
rect 51 -391 52 -389
rect 51 -397 52 -395
rect 58 -391 59 -389
rect 58 -397 59 -395
rect 65 -391 66 -389
rect 68 -391 69 -389
rect 72 -391 73 -389
rect 72 -397 73 -395
rect 79 -391 80 -389
rect 82 -391 83 -389
rect 79 -397 80 -395
rect 82 -397 83 -395
rect 86 -391 87 -389
rect 86 -397 87 -395
rect 96 -391 97 -389
rect 93 -397 94 -395
rect 96 -397 97 -395
rect 100 -391 101 -389
rect 100 -397 101 -395
rect 107 -391 108 -389
rect 110 -391 111 -389
rect 110 -397 111 -395
rect 114 -391 115 -389
rect 117 -397 118 -395
rect 121 -391 122 -389
rect 124 -391 125 -389
rect 121 -397 122 -395
rect 128 -391 129 -389
rect 128 -397 129 -395
rect 135 -391 136 -389
rect 138 -397 139 -395
rect 142 -391 143 -389
rect 142 -397 143 -395
rect 149 -391 150 -389
rect 149 -397 150 -395
rect 159 -391 160 -389
rect 156 -397 157 -395
rect 163 -391 164 -389
rect 163 -397 164 -395
rect 170 -391 171 -389
rect 173 -391 174 -389
rect 170 -397 171 -395
rect 173 -397 174 -395
rect 177 -391 178 -389
rect 177 -397 178 -395
rect 187 -391 188 -389
rect 184 -397 185 -395
rect 187 -397 188 -395
rect 191 -391 192 -389
rect 191 -397 192 -395
rect 198 -391 199 -389
rect 198 -397 199 -395
rect 205 -391 206 -389
rect 205 -397 206 -395
rect 215 -391 216 -389
rect 219 -391 220 -389
rect 219 -397 220 -395
rect 226 -391 227 -389
rect 226 -397 227 -395
rect 233 -391 234 -389
rect 233 -397 234 -395
rect 240 -391 241 -389
rect 240 -397 241 -395
rect 247 -391 248 -389
rect 250 -391 251 -389
rect 247 -397 248 -395
rect 250 -397 251 -395
rect 254 -391 255 -389
rect 257 -391 258 -389
rect 254 -397 255 -395
rect 261 -391 262 -389
rect 264 -391 265 -389
rect 261 -397 262 -395
rect 264 -397 265 -395
rect 268 -391 269 -389
rect 268 -397 269 -395
rect 275 -391 276 -389
rect 275 -397 276 -395
rect 282 -391 283 -389
rect 282 -397 283 -395
rect 289 -391 290 -389
rect 289 -397 290 -395
rect 296 -391 297 -389
rect 296 -397 297 -395
rect 303 -391 304 -389
rect 306 -391 307 -389
rect 306 -397 307 -395
rect 310 -391 311 -389
rect 310 -397 311 -395
rect 317 -391 318 -389
rect 320 -391 321 -389
rect 317 -397 318 -395
rect 320 -397 321 -395
rect 324 -391 325 -389
rect 324 -397 325 -395
rect 327 -397 328 -395
rect 331 -391 332 -389
rect 331 -397 332 -395
rect 341 -391 342 -389
rect 341 -397 342 -395
rect 345 -391 346 -389
rect 345 -397 346 -395
rect 352 -391 353 -389
rect 352 -397 353 -395
rect 359 -391 360 -389
rect 359 -397 360 -395
rect 366 -391 367 -389
rect 366 -397 367 -395
rect 373 -391 374 -389
rect 373 -397 374 -395
rect 380 -397 381 -395
rect 383 -397 384 -395
rect 387 -391 388 -389
rect 387 -397 388 -395
rect 394 -391 395 -389
rect 397 -391 398 -389
rect 394 -397 395 -395
rect 401 -391 402 -389
rect 401 -397 402 -395
rect 408 -391 409 -389
rect 408 -397 409 -395
rect 415 -391 416 -389
rect 415 -397 416 -395
rect 422 -391 423 -389
rect 422 -397 423 -395
rect 429 -391 430 -389
rect 429 -397 430 -395
rect 436 -391 437 -389
rect 436 -397 437 -395
rect 443 -391 444 -389
rect 443 -397 444 -395
rect 450 -391 451 -389
rect 450 -397 451 -395
rect 457 -391 458 -389
rect 457 -397 458 -395
rect 464 -391 465 -389
rect 464 -397 465 -395
rect 474 -391 475 -389
rect 471 -397 472 -395
rect 474 -397 475 -395
rect 478 -391 479 -389
rect 478 -397 479 -395
rect 485 -391 486 -389
rect 485 -397 486 -395
rect 492 -397 493 -395
rect 495 -397 496 -395
rect 499 -391 500 -389
rect 499 -397 500 -395
rect 506 -391 507 -389
rect 506 -397 507 -395
rect 513 -391 514 -389
rect 516 -391 517 -389
rect 516 -397 517 -395
rect 520 -391 521 -389
rect 520 -397 521 -395
rect 527 -391 528 -389
rect 527 -397 528 -395
rect 534 -391 535 -389
rect 534 -397 535 -395
rect 541 -391 542 -389
rect 544 -391 545 -389
rect 541 -397 542 -395
rect 544 -397 545 -395
rect 548 -391 549 -389
rect 548 -397 549 -395
rect 555 -391 556 -389
rect 555 -397 556 -395
rect 562 -391 563 -389
rect 562 -397 563 -395
rect 569 -391 570 -389
rect 569 -397 570 -395
rect 576 -391 577 -389
rect 576 -397 577 -395
rect 583 -391 584 -389
rect 583 -397 584 -395
rect 590 -391 591 -389
rect 590 -397 591 -395
rect 597 -391 598 -389
rect 597 -397 598 -395
rect 604 -391 605 -389
rect 604 -397 605 -395
rect 611 -391 612 -389
rect 611 -397 612 -395
rect 618 -391 619 -389
rect 618 -397 619 -395
rect 628 -391 629 -389
rect 625 -397 626 -395
rect 628 -397 629 -395
rect 632 -391 633 -389
rect 632 -397 633 -395
rect 639 -391 640 -389
rect 639 -397 640 -395
rect 646 -391 647 -389
rect 646 -397 647 -395
rect 653 -391 654 -389
rect 653 -397 654 -395
rect 660 -391 661 -389
rect 660 -397 661 -395
rect 670 -391 671 -389
rect 667 -397 668 -395
rect 674 -391 675 -389
rect 674 -397 675 -395
rect 681 -391 682 -389
rect 681 -397 682 -395
rect 688 -391 689 -389
rect 688 -397 689 -395
rect 695 -391 696 -389
rect 695 -397 696 -395
rect 702 -391 703 -389
rect 702 -397 703 -395
rect 709 -391 710 -389
rect 709 -397 710 -395
rect 716 -391 717 -389
rect 716 -397 717 -395
rect 723 -391 724 -389
rect 723 -397 724 -395
rect 730 -391 731 -389
rect 730 -397 731 -395
rect 737 -391 738 -389
rect 737 -397 738 -395
rect 744 -391 745 -389
rect 744 -397 745 -395
rect 751 -391 752 -389
rect 751 -397 752 -395
rect 758 -391 759 -389
rect 758 -397 759 -395
rect 765 -391 766 -389
rect 765 -397 766 -395
rect 772 -391 773 -389
rect 772 -397 773 -395
rect 779 -391 780 -389
rect 779 -397 780 -395
rect 786 -391 787 -389
rect 786 -397 787 -395
rect 793 -391 794 -389
rect 793 -397 794 -395
rect 800 -391 801 -389
rect 800 -397 801 -395
rect 807 -391 808 -389
rect 807 -397 808 -395
rect 814 -391 815 -389
rect 814 -397 815 -395
rect 821 -391 822 -389
rect 821 -397 822 -395
rect 828 -391 829 -389
rect 828 -397 829 -395
rect 835 -391 836 -389
rect 835 -397 836 -395
rect 842 -391 843 -389
rect 842 -397 843 -395
rect 849 -391 850 -389
rect 849 -397 850 -395
rect 856 -391 857 -389
rect 856 -397 857 -395
rect 863 -391 864 -389
rect 863 -397 864 -395
rect 870 -391 871 -389
rect 870 -397 871 -395
rect 877 -391 878 -389
rect 880 -391 881 -389
rect 877 -397 878 -395
rect 884 -391 885 -389
rect 887 -391 888 -389
rect 884 -397 885 -395
rect 891 -391 892 -389
rect 891 -397 892 -395
rect 898 -391 899 -389
rect 898 -397 899 -395
rect 905 -391 906 -389
rect 905 -397 906 -395
rect 933 -391 934 -389
rect 933 -397 934 -395
rect 1108 -391 1109 -389
rect 1108 -397 1109 -395
rect 2 -480 3 -478
rect 2 -486 3 -484
rect 12 -480 13 -478
rect 16 -480 17 -478
rect 16 -486 17 -484
rect 23 -480 24 -478
rect 23 -486 24 -484
rect 30 -480 31 -478
rect 30 -486 31 -484
rect 37 -480 38 -478
rect 37 -486 38 -484
rect 44 -480 45 -478
rect 44 -486 45 -484
rect 51 -480 52 -478
rect 51 -486 52 -484
rect 61 -480 62 -478
rect 61 -486 62 -484
rect 65 -480 66 -478
rect 68 -480 69 -478
rect 72 -480 73 -478
rect 72 -486 73 -484
rect 79 -480 80 -478
rect 79 -486 80 -484
rect 86 -480 87 -478
rect 86 -486 87 -484
rect 93 -480 94 -478
rect 93 -486 94 -484
rect 100 -480 101 -478
rect 100 -486 101 -484
rect 107 -480 108 -478
rect 107 -486 108 -484
rect 114 -480 115 -478
rect 114 -486 115 -484
rect 121 -480 122 -478
rect 124 -480 125 -478
rect 131 -480 132 -478
rect 128 -486 129 -484
rect 135 -480 136 -478
rect 135 -486 136 -484
rect 142 -480 143 -478
rect 145 -480 146 -478
rect 142 -486 143 -484
rect 145 -486 146 -484
rect 149 -480 150 -478
rect 149 -486 150 -484
rect 156 -480 157 -478
rect 156 -486 157 -484
rect 163 -480 164 -478
rect 163 -486 164 -484
rect 170 -480 171 -478
rect 170 -486 171 -484
rect 177 -480 178 -478
rect 180 -480 181 -478
rect 184 -480 185 -478
rect 184 -486 185 -484
rect 191 -480 192 -478
rect 191 -486 192 -484
rect 198 -480 199 -478
rect 198 -486 199 -484
rect 205 -480 206 -478
rect 208 -486 209 -484
rect 212 -480 213 -478
rect 212 -486 213 -484
rect 219 -480 220 -478
rect 219 -486 220 -484
rect 226 -480 227 -478
rect 226 -486 227 -484
rect 233 -480 234 -478
rect 233 -486 234 -484
rect 240 -480 241 -478
rect 240 -486 241 -484
rect 247 -480 248 -478
rect 247 -486 248 -484
rect 254 -480 255 -478
rect 254 -486 255 -484
rect 261 -480 262 -478
rect 261 -486 262 -484
rect 268 -480 269 -478
rect 268 -486 269 -484
rect 275 -480 276 -478
rect 275 -486 276 -484
rect 282 -486 283 -484
rect 285 -486 286 -484
rect 289 -480 290 -478
rect 289 -486 290 -484
rect 296 -480 297 -478
rect 296 -486 297 -484
rect 303 -480 304 -478
rect 303 -486 304 -484
rect 310 -480 311 -478
rect 310 -486 311 -484
rect 317 -480 318 -478
rect 317 -486 318 -484
rect 324 -480 325 -478
rect 327 -480 328 -478
rect 324 -486 325 -484
rect 327 -486 328 -484
rect 331 -480 332 -478
rect 331 -486 332 -484
rect 338 -480 339 -478
rect 338 -486 339 -484
rect 345 -480 346 -478
rect 348 -486 349 -484
rect 352 -480 353 -478
rect 352 -486 353 -484
rect 355 -486 356 -484
rect 359 -480 360 -478
rect 359 -486 360 -484
rect 366 -480 367 -478
rect 366 -486 367 -484
rect 373 -480 374 -478
rect 373 -486 374 -484
rect 380 -480 381 -478
rect 383 -480 384 -478
rect 383 -486 384 -484
rect 387 -480 388 -478
rect 387 -486 388 -484
rect 397 -480 398 -478
rect 397 -486 398 -484
rect 401 -480 402 -478
rect 401 -486 402 -484
rect 408 -480 409 -478
rect 408 -486 409 -484
rect 415 -486 416 -484
rect 418 -486 419 -484
rect 422 -480 423 -478
rect 425 -480 426 -478
rect 422 -486 423 -484
rect 425 -486 426 -484
rect 429 -480 430 -478
rect 429 -486 430 -484
rect 436 -480 437 -478
rect 436 -486 437 -484
rect 443 -480 444 -478
rect 443 -486 444 -484
rect 450 -480 451 -478
rect 450 -486 451 -484
rect 457 -480 458 -478
rect 460 -480 461 -478
rect 457 -486 458 -484
rect 460 -486 461 -484
rect 464 -480 465 -478
rect 464 -486 465 -484
rect 474 -480 475 -478
rect 471 -486 472 -484
rect 481 -480 482 -478
rect 481 -486 482 -484
rect 485 -480 486 -478
rect 485 -486 486 -484
rect 492 -480 493 -478
rect 492 -486 493 -484
rect 499 -480 500 -478
rect 502 -480 503 -478
rect 502 -486 503 -484
rect 506 -480 507 -478
rect 506 -486 507 -484
rect 513 -480 514 -478
rect 513 -486 514 -484
rect 520 -480 521 -478
rect 520 -486 521 -484
rect 527 -480 528 -478
rect 527 -486 528 -484
rect 534 -480 535 -478
rect 534 -486 535 -484
rect 537 -486 538 -484
rect 541 -480 542 -478
rect 541 -486 542 -484
rect 548 -480 549 -478
rect 548 -486 549 -484
rect 555 -480 556 -478
rect 558 -480 559 -478
rect 555 -486 556 -484
rect 562 -486 563 -484
rect 565 -486 566 -484
rect 569 -480 570 -478
rect 572 -480 573 -478
rect 569 -486 570 -484
rect 572 -486 573 -484
rect 576 -480 577 -478
rect 579 -480 580 -478
rect 583 -480 584 -478
rect 583 -486 584 -484
rect 590 -480 591 -478
rect 590 -486 591 -484
rect 597 -480 598 -478
rect 597 -486 598 -484
rect 604 -480 605 -478
rect 604 -486 605 -484
rect 611 -480 612 -478
rect 611 -486 612 -484
rect 618 -480 619 -478
rect 618 -486 619 -484
rect 625 -480 626 -478
rect 625 -486 626 -484
rect 635 -480 636 -478
rect 632 -486 633 -484
rect 635 -486 636 -484
rect 642 -486 643 -484
rect 646 -480 647 -478
rect 646 -486 647 -484
rect 653 -480 654 -478
rect 653 -486 654 -484
rect 660 -480 661 -478
rect 660 -486 661 -484
rect 667 -480 668 -478
rect 667 -486 668 -484
rect 674 -480 675 -478
rect 674 -486 675 -484
rect 681 -480 682 -478
rect 681 -486 682 -484
rect 688 -480 689 -478
rect 688 -486 689 -484
rect 695 -480 696 -478
rect 695 -486 696 -484
rect 702 -480 703 -478
rect 702 -486 703 -484
rect 709 -480 710 -478
rect 709 -486 710 -484
rect 716 -480 717 -478
rect 716 -486 717 -484
rect 723 -480 724 -478
rect 723 -486 724 -484
rect 730 -480 731 -478
rect 730 -486 731 -484
rect 737 -480 738 -478
rect 737 -486 738 -484
rect 744 -480 745 -478
rect 744 -486 745 -484
rect 751 -480 752 -478
rect 751 -486 752 -484
rect 758 -480 759 -478
rect 758 -486 759 -484
rect 765 -480 766 -478
rect 765 -486 766 -484
rect 772 -480 773 -478
rect 772 -486 773 -484
rect 779 -480 780 -478
rect 779 -486 780 -484
rect 786 -480 787 -478
rect 786 -486 787 -484
rect 793 -480 794 -478
rect 793 -486 794 -484
rect 800 -480 801 -478
rect 800 -486 801 -484
rect 807 -480 808 -478
rect 807 -486 808 -484
rect 814 -486 815 -484
rect 817 -486 818 -484
rect 821 -480 822 -478
rect 821 -486 822 -484
rect 828 -480 829 -478
rect 828 -486 829 -484
rect 835 -480 836 -478
rect 835 -486 836 -484
rect 842 -480 843 -478
rect 842 -486 843 -484
rect 849 -480 850 -478
rect 849 -486 850 -484
rect 856 -480 857 -478
rect 856 -486 857 -484
rect 863 -480 864 -478
rect 863 -486 864 -484
rect 870 -480 871 -478
rect 870 -486 871 -484
rect 877 -480 878 -478
rect 877 -486 878 -484
rect 884 -480 885 -478
rect 884 -486 885 -484
rect 891 -480 892 -478
rect 891 -486 892 -484
rect 898 -480 899 -478
rect 898 -486 899 -484
rect 905 -480 906 -478
rect 905 -486 906 -484
rect 912 -480 913 -478
rect 912 -486 913 -484
rect 919 -480 920 -478
rect 919 -486 920 -484
rect 926 -480 927 -478
rect 926 -486 927 -484
rect 933 -480 934 -478
rect 933 -486 934 -484
rect 940 -480 941 -478
rect 940 -486 941 -484
rect 947 -480 948 -478
rect 947 -486 948 -484
rect 954 -480 955 -478
rect 954 -486 955 -484
rect 961 -480 962 -478
rect 961 -486 962 -484
rect 968 -480 969 -478
rect 968 -486 969 -484
rect 975 -480 976 -478
rect 975 -486 976 -484
rect 982 -480 983 -478
rect 982 -486 983 -484
rect 989 -480 990 -478
rect 989 -486 990 -484
rect 996 -480 997 -478
rect 996 -486 997 -484
rect 1003 -480 1004 -478
rect 1003 -486 1004 -484
rect 1010 -480 1011 -478
rect 1010 -486 1011 -484
rect 1017 -480 1018 -478
rect 1017 -486 1018 -484
rect 1024 -480 1025 -478
rect 1024 -486 1025 -484
rect 1031 -480 1032 -478
rect 1034 -480 1035 -478
rect 1038 -480 1039 -478
rect 1045 -480 1046 -478
rect 1045 -486 1046 -484
rect 1115 -480 1116 -478
rect 1115 -486 1116 -484
rect 2 -603 3 -601
rect 5 -603 6 -601
rect 9 -597 10 -595
rect 9 -603 10 -601
rect 16 -597 17 -595
rect 16 -603 17 -601
rect 26 -597 27 -595
rect 26 -603 27 -601
rect 30 -597 31 -595
rect 30 -603 31 -601
rect 37 -603 38 -601
rect 40 -603 41 -601
rect 44 -597 45 -595
rect 44 -603 45 -601
rect 51 -597 52 -595
rect 51 -603 52 -601
rect 58 -597 59 -595
rect 58 -603 59 -601
rect 65 -597 66 -595
rect 65 -603 66 -601
rect 72 -597 73 -595
rect 72 -603 73 -601
rect 79 -597 80 -595
rect 79 -603 80 -601
rect 86 -597 87 -595
rect 86 -603 87 -601
rect 93 -597 94 -595
rect 96 -597 97 -595
rect 93 -603 94 -601
rect 100 -597 101 -595
rect 100 -603 101 -601
rect 103 -603 104 -601
rect 107 -597 108 -595
rect 107 -603 108 -601
rect 114 -597 115 -595
rect 114 -603 115 -601
rect 121 -597 122 -595
rect 121 -603 122 -601
rect 128 -597 129 -595
rect 128 -603 129 -601
rect 135 -597 136 -595
rect 138 -597 139 -595
rect 135 -603 136 -601
rect 138 -603 139 -601
rect 142 -597 143 -595
rect 142 -603 143 -601
rect 149 -597 150 -595
rect 149 -603 150 -601
rect 156 -597 157 -595
rect 156 -603 157 -601
rect 163 -597 164 -595
rect 166 -597 167 -595
rect 163 -603 164 -601
rect 170 -597 171 -595
rect 170 -603 171 -601
rect 180 -597 181 -595
rect 177 -603 178 -601
rect 184 -597 185 -595
rect 184 -603 185 -601
rect 191 -597 192 -595
rect 191 -603 192 -601
rect 198 -597 199 -595
rect 198 -603 199 -601
rect 205 -597 206 -595
rect 208 -597 209 -595
rect 205 -603 206 -601
rect 212 -597 213 -595
rect 215 -597 216 -595
rect 212 -603 213 -601
rect 215 -603 216 -601
rect 219 -597 220 -595
rect 219 -603 220 -601
rect 222 -603 223 -601
rect 226 -597 227 -595
rect 226 -603 227 -601
rect 233 -597 234 -595
rect 233 -603 234 -601
rect 240 -597 241 -595
rect 240 -603 241 -601
rect 247 -597 248 -595
rect 247 -603 248 -601
rect 254 -597 255 -595
rect 254 -603 255 -601
rect 261 -597 262 -595
rect 261 -603 262 -601
rect 268 -597 269 -595
rect 271 -597 272 -595
rect 268 -603 269 -601
rect 275 -597 276 -595
rect 275 -603 276 -601
rect 282 -597 283 -595
rect 282 -603 283 -601
rect 289 -597 290 -595
rect 289 -603 290 -601
rect 296 -597 297 -595
rect 296 -603 297 -601
rect 303 -597 304 -595
rect 303 -603 304 -601
rect 310 -597 311 -595
rect 310 -603 311 -601
rect 317 -597 318 -595
rect 317 -603 318 -601
rect 324 -597 325 -595
rect 324 -603 325 -601
rect 331 -597 332 -595
rect 331 -603 332 -601
rect 341 -597 342 -595
rect 338 -603 339 -601
rect 341 -603 342 -601
rect 345 -597 346 -595
rect 348 -597 349 -595
rect 345 -603 346 -601
rect 348 -603 349 -601
rect 352 -597 353 -595
rect 352 -603 353 -601
rect 359 -597 360 -595
rect 359 -603 360 -601
rect 366 -597 367 -595
rect 366 -603 367 -601
rect 373 -597 374 -595
rect 373 -603 374 -601
rect 380 -597 381 -595
rect 380 -603 381 -601
rect 387 -597 388 -595
rect 387 -603 388 -601
rect 394 -597 395 -595
rect 394 -603 395 -601
rect 401 -597 402 -595
rect 401 -603 402 -601
rect 408 -597 409 -595
rect 408 -603 409 -601
rect 415 -597 416 -595
rect 415 -603 416 -601
rect 422 -597 423 -595
rect 422 -603 423 -601
rect 429 -597 430 -595
rect 429 -603 430 -601
rect 436 -597 437 -595
rect 439 -603 440 -601
rect 443 -597 444 -595
rect 443 -603 444 -601
rect 450 -597 451 -595
rect 450 -603 451 -601
rect 457 -597 458 -595
rect 457 -603 458 -601
rect 464 -597 465 -595
rect 467 -603 468 -601
rect 471 -597 472 -595
rect 474 -597 475 -595
rect 471 -603 472 -601
rect 474 -603 475 -601
rect 478 -597 479 -595
rect 478 -603 479 -601
rect 485 -597 486 -595
rect 485 -603 486 -601
rect 492 -597 493 -595
rect 492 -603 493 -601
rect 499 -597 500 -595
rect 499 -603 500 -601
rect 506 -597 507 -595
rect 506 -603 507 -601
rect 513 -597 514 -595
rect 513 -603 514 -601
rect 523 -597 524 -595
rect 520 -603 521 -601
rect 523 -603 524 -601
rect 527 -597 528 -595
rect 530 -597 531 -595
rect 534 -597 535 -595
rect 537 -597 538 -595
rect 534 -603 535 -601
rect 541 -597 542 -595
rect 541 -603 542 -601
rect 548 -597 549 -595
rect 551 -597 552 -595
rect 548 -603 549 -601
rect 551 -603 552 -601
rect 555 -597 556 -595
rect 555 -603 556 -601
rect 562 -597 563 -595
rect 565 -597 566 -595
rect 562 -603 563 -601
rect 572 -597 573 -595
rect 569 -603 570 -601
rect 572 -603 573 -601
rect 576 -597 577 -595
rect 579 -597 580 -595
rect 576 -603 577 -601
rect 579 -603 580 -601
rect 583 -597 584 -595
rect 583 -603 584 -601
rect 590 -597 591 -595
rect 590 -603 591 -601
rect 597 -597 598 -595
rect 600 -597 601 -595
rect 597 -603 598 -601
rect 604 -597 605 -595
rect 604 -603 605 -601
rect 611 -597 612 -595
rect 611 -603 612 -601
rect 618 -597 619 -595
rect 618 -603 619 -601
rect 625 -597 626 -595
rect 625 -603 626 -601
rect 632 -597 633 -595
rect 632 -603 633 -601
rect 639 -597 640 -595
rect 639 -603 640 -601
rect 646 -597 647 -595
rect 646 -603 647 -601
rect 653 -597 654 -595
rect 653 -603 654 -601
rect 660 -597 661 -595
rect 660 -603 661 -601
rect 667 -597 668 -595
rect 667 -603 668 -601
rect 674 -597 675 -595
rect 674 -603 675 -601
rect 681 -597 682 -595
rect 684 -597 685 -595
rect 684 -603 685 -601
rect 688 -597 689 -595
rect 688 -603 689 -601
rect 695 -597 696 -595
rect 695 -603 696 -601
rect 702 -597 703 -595
rect 702 -603 703 -601
rect 709 -597 710 -595
rect 712 -597 713 -595
rect 712 -603 713 -601
rect 716 -597 717 -595
rect 716 -603 717 -601
rect 723 -597 724 -595
rect 723 -603 724 -601
rect 733 -603 734 -601
rect 737 -597 738 -595
rect 737 -603 738 -601
rect 744 -597 745 -595
rect 744 -603 745 -601
rect 751 -597 752 -595
rect 751 -603 752 -601
rect 758 -597 759 -595
rect 758 -603 759 -601
rect 765 -597 766 -595
rect 765 -603 766 -601
rect 772 -597 773 -595
rect 772 -603 773 -601
rect 779 -597 780 -595
rect 779 -603 780 -601
rect 786 -597 787 -595
rect 786 -603 787 -601
rect 793 -597 794 -595
rect 793 -603 794 -601
rect 800 -597 801 -595
rect 800 -603 801 -601
rect 807 -597 808 -595
rect 807 -603 808 -601
rect 814 -597 815 -595
rect 814 -603 815 -601
rect 821 -597 822 -595
rect 821 -603 822 -601
rect 828 -597 829 -595
rect 828 -603 829 -601
rect 835 -597 836 -595
rect 835 -603 836 -601
rect 842 -597 843 -595
rect 842 -603 843 -601
rect 849 -597 850 -595
rect 849 -603 850 -601
rect 856 -597 857 -595
rect 856 -603 857 -601
rect 863 -597 864 -595
rect 863 -603 864 -601
rect 870 -597 871 -595
rect 870 -603 871 -601
rect 877 -597 878 -595
rect 877 -603 878 -601
rect 884 -597 885 -595
rect 884 -603 885 -601
rect 891 -597 892 -595
rect 891 -603 892 -601
rect 898 -597 899 -595
rect 898 -603 899 -601
rect 905 -597 906 -595
rect 905 -603 906 -601
rect 912 -597 913 -595
rect 912 -603 913 -601
rect 919 -597 920 -595
rect 919 -603 920 -601
rect 926 -597 927 -595
rect 926 -603 927 -601
rect 933 -597 934 -595
rect 933 -603 934 -601
rect 940 -597 941 -595
rect 940 -603 941 -601
rect 947 -597 948 -595
rect 947 -603 948 -601
rect 954 -597 955 -595
rect 954 -603 955 -601
rect 961 -597 962 -595
rect 961 -603 962 -601
rect 968 -597 969 -595
rect 968 -603 969 -601
rect 975 -597 976 -595
rect 975 -603 976 -601
rect 982 -597 983 -595
rect 982 -603 983 -601
rect 989 -597 990 -595
rect 989 -603 990 -601
rect 996 -597 997 -595
rect 996 -603 997 -601
rect 1003 -597 1004 -595
rect 1003 -603 1004 -601
rect 1010 -597 1011 -595
rect 1010 -603 1011 -601
rect 1017 -597 1018 -595
rect 1017 -603 1018 -601
rect 1024 -597 1025 -595
rect 1024 -603 1025 -601
rect 1031 -597 1032 -595
rect 1031 -603 1032 -601
rect 1038 -597 1039 -595
rect 1038 -603 1039 -601
rect 1045 -597 1046 -595
rect 1045 -603 1046 -601
rect 1052 -597 1053 -595
rect 1052 -603 1053 -601
rect 1059 -597 1060 -595
rect 1059 -603 1060 -601
rect 1066 -597 1067 -595
rect 1066 -603 1067 -601
rect 1073 -597 1074 -595
rect 1073 -603 1074 -601
rect 1080 -597 1081 -595
rect 1080 -603 1081 -601
rect 1087 -597 1088 -595
rect 1087 -603 1088 -601
rect 1094 -597 1095 -595
rect 1094 -603 1095 -601
rect 1101 -603 1102 -601
rect 1111 -597 1112 -595
rect 1108 -603 1109 -601
rect 1115 -597 1116 -595
rect 1115 -603 1116 -601
rect 1122 -597 1123 -595
rect 1122 -603 1123 -601
rect 1129 -597 1130 -595
rect 1129 -603 1130 -601
rect 2 -698 3 -696
rect 2 -704 3 -702
rect 9 -704 10 -702
rect 16 -698 17 -696
rect 16 -704 17 -702
rect 23 -698 24 -696
rect 23 -704 24 -702
rect 30 -698 31 -696
rect 30 -704 31 -702
rect 37 -698 38 -696
rect 37 -704 38 -702
rect 44 -698 45 -696
rect 47 -698 48 -696
rect 51 -698 52 -696
rect 51 -704 52 -702
rect 58 -698 59 -696
rect 58 -704 59 -702
rect 65 -698 66 -696
rect 65 -704 66 -702
rect 72 -698 73 -696
rect 72 -704 73 -702
rect 82 -698 83 -696
rect 79 -704 80 -702
rect 82 -704 83 -702
rect 86 -698 87 -696
rect 86 -704 87 -702
rect 93 -698 94 -696
rect 93 -704 94 -702
rect 100 -698 101 -696
rect 100 -704 101 -702
rect 107 -698 108 -696
rect 107 -704 108 -702
rect 117 -698 118 -696
rect 114 -704 115 -702
rect 124 -698 125 -696
rect 121 -704 122 -702
rect 124 -704 125 -702
rect 128 -698 129 -696
rect 131 -698 132 -696
rect 131 -704 132 -702
rect 135 -698 136 -696
rect 135 -704 136 -702
rect 142 -698 143 -696
rect 142 -704 143 -702
rect 149 -698 150 -696
rect 149 -704 150 -702
rect 156 -698 157 -696
rect 156 -704 157 -702
rect 163 -698 164 -696
rect 163 -704 164 -702
rect 173 -698 174 -696
rect 170 -704 171 -702
rect 177 -698 178 -696
rect 177 -704 178 -702
rect 184 -698 185 -696
rect 184 -704 185 -702
rect 191 -698 192 -696
rect 191 -704 192 -702
rect 201 -698 202 -696
rect 198 -704 199 -702
rect 205 -698 206 -696
rect 205 -704 206 -702
rect 208 -704 209 -702
rect 212 -698 213 -696
rect 212 -704 213 -702
rect 219 -698 220 -696
rect 219 -704 220 -702
rect 226 -704 227 -702
rect 233 -698 234 -696
rect 233 -704 234 -702
rect 240 -698 241 -696
rect 240 -704 241 -702
rect 247 -698 248 -696
rect 247 -704 248 -702
rect 254 -698 255 -696
rect 254 -704 255 -702
rect 261 -698 262 -696
rect 261 -704 262 -702
rect 268 -698 269 -696
rect 268 -704 269 -702
rect 275 -698 276 -696
rect 275 -704 276 -702
rect 282 -698 283 -696
rect 282 -704 283 -702
rect 292 -698 293 -696
rect 289 -704 290 -702
rect 292 -704 293 -702
rect 296 -698 297 -696
rect 296 -704 297 -702
rect 303 -698 304 -696
rect 303 -704 304 -702
rect 313 -698 314 -696
rect 310 -704 311 -702
rect 317 -698 318 -696
rect 317 -704 318 -702
rect 324 -698 325 -696
rect 324 -704 325 -702
rect 331 -698 332 -696
rect 331 -704 332 -702
rect 338 -698 339 -696
rect 338 -704 339 -702
rect 345 -698 346 -696
rect 345 -704 346 -702
rect 352 -698 353 -696
rect 352 -704 353 -702
rect 359 -698 360 -696
rect 362 -698 363 -696
rect 359 -704 360 -702
rect 362 -704 363 -702
rect 366 -698 367 -696
rect 366 -704 367 -702
rect 373 -698 374 -696
rect 373 -704 374 -702
rect 380 -698 381 -696
rect 380 -704 381 -702
rect 387 -698 388 -696
rect 387 -704 388 -702
rect 394 -698 395 -696
rect 394 -704 395 -702
rect 401 -698 402 -696
rect 401 -704 402 -702
rect 408 -698 409 -696
rect 408 -704 409 -702
rect 415 -698 416 -696
rect 415 -704 416 -702
rect 422 -698 423 -696
rect 422 -704 423 -702
rect 429 -698 430 -696
rect 429 -704 430 -702
rect 436 -698 437 -696
rect 436 -704 437 -702
rect 443 -698 444 -696
rect 443 -704 444 -702
rect 446 -704 447 -702
rect 450 -698 451 -696
rect 453 -698 454 -696
rect 453 -704 454 -702
rect 457 -698 458 -696
rect 460 -698 461 -696
rect 457 -704 458 -702
rect 460 -704 461 -702
rect 467 -698 468 -696
rect 464 -704 465 -702
rect 467 -704 468 -702
rect 471 -698 472 -696
rect 471 -704 472 -702
rect 478 -698 479 -696
rect 481 -698 482 -696
rect 478 -704 479 -702
rect 485 -698 486 -696
rect 485 -704 486 -702
rect 492 -698 493 -696
rect 495 -698 496 -696
rect 495 -704 496 -702
rect 499 -698 500 -696
rect 499 -704 500 -702
rect 506 -698 507 -696
rect 506 -704 507 -702
rect 513 -698 514 -696
rect 516 -698 517 -696
rect 513 -704 514 -702
rect 516 -704 517 -702
rect 520 -698 521 -696
rect 520 -704 521 -702
rect 527 -698 528 -696
rect 527 -704 528 -702
rect 534 -698 535 -696
rect 534 -704 535 -702
rect 541 -698 542 -696
rect 544 -698 545 -696
rect 544 -704 545 -702
rect 548 -698 549 -696
rect 548 -704 549 -702
rect 555 -698 556 -696
rect 555 -704 556 -702
rect 562 -698 563 -696
rect 565 -698 566 -696
rect 562 -704 563 -702
rect 569 -698 570 -696
rect 569 -704 570 -702
rect 576 -698 577 -696
rect 576 -704 577 -702
rect 583 -698 584 -696
rect 583 -704 584 -702
rect 590 -698 591 -696
rect 590 -704 591 -702
rect 597 -698 598 -696
rect 597 -704 598 -702
rect 604 -698 605 -696
rect 607 -698 608 -696
rect 611 -698 612 -696
rect 611 -704 612 -702
rect 618 -698 619 -696
rect 618 -704 619 -702
rect 625 -698 626 -696
rect 625 -704 626 -702
rect 632 -698 633 -696
rect 632 -704 633 -702
rect 639 -698 640 -696
rect 639 -704 640 -702
rect 646 -698 647 -696
rect 646 -704 647 -702
rect 653 -698 654 -696
rect 653 -704 654 -702
rect 660 -698 661 -696
rect 660 -704 661 -702
rect 667 -698 668 -696
rect 674 -698 675 -696
rect 674 -704 675 -702
rect 681 -698 682 -696
rect 681 -704 682 -702
rect 688 -698 689 -696
rect 688 -704 689 -702
rect 695 -698 696 -696
rect 695 -704 696 -702
rect 702 -698 703 -696
rect 702 -704 703 -702
rect 709 -698 710 -696
rect 709 -704 710 -702
rect 716 -698 717 -696
rect 716 -704 717 -702
rect 723 -698 724 -696
rect 726 -698 727 -696
rect 723 -704 724 -702
rect 726 -704 727 -702
rect 730 -698 731 -696
rect 730 -704 731 -702
rect 737 -698 738 -696
rect 737 -704 738 -702
rect 747 -704 748 -702
rect 751 -698 752 -696
rect 751 -704 752 -702
rect 758 -698 759 -696
rect 758 -704 759 -702
rect 765 -698 766 -696
rect 765 -704 766 -702
rect 775 -698 776 -696
rect 772 -704 773 -702
rect 775 -704 776 -702
rect 779 -698 780 -696
rect 779 -704 780 -702
rect 786 -698 787 -696
rect 789 -698 790 -696
rect 786 -704 787 -702
rect 793 -698 794 -696
rect 793 -704 794 -702
rect 800 -698 801 -696
rect 800 -704 801 -702
rect 807 -698 808 -696
rect 807 -704 808 -702
rect 814 -698 815 -696
rect 814 -704 815 -702
rect 821 -698 822 -696
rect 821 -704 822 -702
rect 828 -698 829 -696
rect 828 -704 829 -702
rect 835 -698 836 -696
rect 835 -704 836 -702
rect 842 -698 843 -696
rect 842 -704 843 -702
rect 849 -698 850 -696
rect 849 -704 850 -702
rect 856 -698 857 -696
rect 856 -704 857 -702
rect 863 -698 864 -696
rect 863 -704 864 -702
rect 870 -698 871 -696
rect 870 -704 871 -702
rect 877 -698 878 -696
rect 877 -704 878 -702
rect 884 -698 885 -696
rect 884 -704 885 -702
rect 891 -698 892 -696
rect 891 -704 892 -702
rect 898 -698 899 -696
rect 898 -704 899 -702
rect 905 -698 906 -696
rect 905 -704 906 -702
rect 912 -698 913 -696
rect 912 -704 913 -702
rect 919 -698 920 -696
rect 919 -704 920 -702
rect 926 -698 927 -696
rect 926 -704 927 -702
rect 933 -698 934 -696
rect 933 -704 934 -702
rect 940 -698 941 -696
rect 940 -704 941 -702
rect 947 -698 948 -696
rect 947 -704 948 -702
rect 954 -698 955 -696
rect 954 -704 955 -702
rect 961 -698 962 -696
rect 961 -704 962 -702
rect 968 -698 969 -696
rect 968 -704 969 -702
rect 975 -698 976 -696
rect 975 -704 976 -702
rect 982 -698 983 -696
rect 982 -704 983 -702
rect 989 -698 990 -696
rect 989 -704 990 -702
rect 996 -698 997 -696
rect 996 -704 997 -702
rect 1003 -698 1004 -696
rect 1003 -704 1004 -702
rect 1010 -698 1011 -696
rect 1010 -704 1011 -702
rect 1017 -698 1018 -696
rect 1017 -704 1018 -702
rect 1024 -698 1025 -696
rect 1024 -704 1025 -702
rect 1031 -698 1032 -696
rect 1031 -704 1032 -702
rect 1038 -698 1039 -696
rect 1038 -704 1039 -702
rect 1045 -698 1046 -696
rect 1045 -704 1046 -702
rect 1052 -698 1053 -696
rect 1052 -704 1053 -702
rect 1059 -698 1060 -696
rect 1059 -704 1060 -702
rect 1066 -698 1067 -696
rect 1066 -704 1067 -702
rect 1073 -698 1074 -696
rect 1073 -704 1074 -702
rect 1080 -698 1081 -696
rect 1080 -704 1081 -702
rect 1083 -704 1084 -702
rect 1087 -698 1088 -696
rect 1087 -704 1088 -702
rect 1094 -698 1095 -696
rect 1094 -704 1095 -702
rect 1101 -698 1102 -696
rect 1101 -704 1102 -702
rect 1111 -698 1112 -696
rect 1111 -704 1112 -702
rect 1115 -698 1116 -696
rect 1115 -704 1116 -702
rect 1122 -698 1123 -696
rect 1122 -704 1123 -702
rect 1129 -698 1130 -696
rect 1129 -704 1130 -702
rect 1139 -698 1140 -696
rect 1143 -698 1144 -696
rect 1143 -704 1144 -702
rect 1150 -698 1151 -696
rect 1150 -704 1151 -702
rect 1157 -698 1158 -696
rect 1157 -704 1158 -702
rect 23 -775 24 -773
rect 23 -781 24 -779
rect 30 -775 31 -773
rect 37 -775 38 -773
rect 37 -781 38 -779
rect 44 -775 45 -773
rect 44 -781 45 -779
rect 51 -775 52 -773
rect 51 -781 52 -779
rect 58 -775 59 -773
rect 58 -781 59 -779
rect 65 -775 66 -773
rect 65 -781 66 -779
rect 72 -775 73 -773
rect 72 -781 73 -779
rect 79 -775 80 -773
rect 79 -781 80 -779
rect 86 -775 87 -773
rect 89 -775 90 -773
rect 86 -781 87 -779
rect 93 -775 94 -773
rect 93 -781 94 -779
rect 100 -775 101 -773
rect 103 -775 104 -773
rect 103 -781 104 -779
rect 107 -775 108 -773
rect 107 -781 108 -779
rect 114 -775 115 -773
rect 114 -781 115 -779
rect 121 -775 122 -773
rect 121 -781 122 -779
rect 128 -775 129 -773
rect 128 -781 129 -779
rect 135 -775 136 -773
rect 135 -781 136 -779
rect 138 -781 139 -779
rect 142 -775 143 -773
rect 142 -781 143 -779
rect 149 -775 150 -773
rect 152 -775 153 -773
rect 152 -781 153 -779
rect 156 -775 157 -773
rect 159 -775 160 -773
rect 156 -781 157 -779
rect 163 -775 164 -773
rect 163 -781 164 -779
rect 170 -775 171 -773
rect 173 -775 174 -773
rect 173 -781 174 -779
rect 177 -775 178 -773
rect 177 -781 178 -779
rect 184 -775 185 -773
rect 184 -781 185 -779
rect 191 -775 192 -773
rect 191 -781 192 -779
rect 198 -775 199 -773
rect 198 -781 199 -779
rect 208 -775 209 -773
rect 208 -781 209 -779
rect 212 -775 213 -773
rect 212 -781 213 -779
rect 219 -775 220 -773
rect 219 -781 220 -779
rect 226 -775 227 -773
rect 226 -781 227 -779
rect 233 -775 234 -773
rect 233 -781 234 -779
rect 240 -775 241 -773
rect 240 -781 241 -779
rect 247 -775 248 -773
rect 247 -781 248 -779
rect 254 -775 255 -773
rect 254 -781 255 -779
rect 261 -775 262 -773
rect 261 -781 262 -779
rect 268 -775 269 -773
rect 268 -781 269 -779
rect 275 -775 276 -773
rect 275 -781 276 -779
rect 282 -775 283 -773
rect 282 -781 283 -779
rect 289 -775 290 -773
rect 292 -775 293 -773
rect 292 -781 293 -779
rect 296 -775 297 -773
rect 296 -781 297 -779
rect 303 -775 304 -773
rect 303 -781 304 -779
rect 310 -775 311 -773
rect 313 -781 314 -779
rect 317 -775 318 -773
rect 317 -781 318 -779
rect 324 -775 325 -773
rect 327 -775 328 -773
rect 324 -781 325 -779
rect 331 -775 332 -773
rect 331 -781 332 -779
rect 338 -775 339 -773
rect 338 -781 339 -779
rect 345 -775 346 -773
rect 345 -781 346 -779
rect 352 -775 353 -773
rect 352 -781 353 -779
rect 359 -775 360 -773
rect 359 -781 360 -779
rect 369 -775 370 -773
rect 366 -781 367 -779
rect 369 -781 370 -779
rect 373 -775 374 -773
rect 373 -781 374 -779
rect 380 -775 381 -773
rect 380 -781 381 -779
rect 387 -775 388 -773
rect 387 -781 388 -779
rect 394 -775 395 -773
rect 394 -781 395 -779
rect 401 -775 402 -773
rect 401 -781 402 -779
rect 408 -775 409 -773
rect 408 -781 409 -779
rect 415 -775 416 -773
rect 415 -781 416 -779
rect 422 -775 423 -773
rect 422 -781 423 -779
rect 429 -775 430 -773
rect 429 -781 430 -779
rect 436 -775 437 -773
rect 436 -781 437 -779
rect 443 -775 444 -773
rect 446 -775 447 -773
rect 443 -781 444 -779
rect 446 -781 447 -779
rect 450 -775 451 -773
rect 450 -781 451 -779
rect 457 -775 458 -773
rect 460 -775 461 -773
rect 457 -781 458 -779
rect 460 -781 461 -779
rect 464 -781 465 -779
rect 467 -781 468 -779
rect 471 -775 472 -773
rect 471 -781 472 -779
rect 478 -775 479 -773
rect 478 -781 479 -779
rect 485 -775 486 -773
rect 485 -781 486 -779
rect 492 -775 493 -773
rect 492 -781 493 -779
rect 495 -781 496 -779
rect 499 -775 500 -773
rect 499 -781 500 -779
rect 506 -775 507 -773
rect 506 -781 507 -779
rect 513 -775 514 -773
rect 513 -781 514 -779
rect 520 -775 521 -773
rect 520 -781 521 -779
rect 527 -775 528 -773
rect 527 -781 528 -779
rect 530 -781 531 -779
rect 534 -775 535 -773
rect 537 -775 538 -773
rect 534 -781 535 -779
rect 537 -781 538 -779
rect 541 -775 542 -773
rect 541 -781 542 -779
rect 548 -775 549 -773
rect 548 -781 549 -779
rect 555 -775 556 -773
rect 555 -781 556 -779
rect 562 -775 563 -773
rect 562 -781 563 -779
rect 569 -775 570 -773
rect 569 -781 570 -779
rect 576 -775 577 -773
rect 576 -781 577 -779
rect 583 -775 584 -773
rect 583 -781 584 -779
rect 590 -775 591 -773
rect 590 -781 591 -779
rect 597 -775 598 -773
rect 597 -781 598 -779
rect 604 -775 605 -773
rect 604 -781 605 -779
rect 611 -775 612 -773
rect 611 -781 612 -779
rect 618 -775 619 -773
rect 618 -781 619 -779
rect 621 -781 622 -779
rect 625 -775 626 -773
rect 625 -781 626 -779
rect 632 -775 633 -773
rect 632 -781 633 -779
rect 639 -775 640 -773
rect 639 -781 640 -779
rect 646 -775 647 -773
rect 646 -781 647 -779
rect 653 -775 654 -773
rect 656 -775 657 -773
rect 653 -781 654 -779
rect 656 -781 657 -779
rect 660 -775 661 -773
rect 663 -775 664 -773
rect 660 -781 661 -779
rect 663 -781 664 -779
rect 667 -775 668 -773
rect 667 -781 668 -779
rect 674 -775 675 -773
rect 674 -781 675 -779
rect 681 -775 682 -773
rect 681 -781 682 -779
rect 688 -775 689 -773
rect 688 -781 689 -779
rect 695 -775 696 -773
rect 695 -781 696 -779
rect 702 -775 703 -773
rect 705 -775 706 -773
rect 702 -781 703 -779
rect 705 -781 706 -779
rect 709 -775 710 -773
rect 709 -781 710 -779
rect 716 -775 717 -773
rect 719 -775 720 -773
rect 719 -781 720 -779
rect 723 -775 724 -773
rect 723 -781 724 -779
rect 730 -775 731 -773
rect 730 -781 731 -779
rect 737 -775 738 -773
rect 737 -781 738 -779
rect 744 -775 745 -773
rect 744 -781 745 -779
rect 751 -775 752 -773
rect 751 -781 752 -779
rect 758 -775 759 -773
rect 761 -775 762 -773
rect 765 -775 766 -773
rect 765 -781 766 -779
rect 772 -775 773 -773
rect 775 -775 776 -773
rect 772 -781 773 -779
rect 775 -781 776 -779
rect 779 -775 780 -773
rect 779 -781 780 -779
rect 786 -775 787 -773
rect 786 -781 787 -779
rect 793 -781 794 -779
rect 796 -781 797 -779
rect 800 -775 801 -773
rect 800 -781 801 -779
rect 807 -775 808 -773
rect 807 -781 808 -779
rect 814 -775 815 -773
rect 814 -781 815 -779
rect 821 -775 822 -773
rect 821 -781 822 -779
rect 828 -775 829 -773
rect 828 -781 829 -779
rect 835 -775 836 -773
rect 835 -781 836 -779
rect 842 -775 843 -773
rect 842 -781 843 -779
rect 849 -775 850 -773
rect 849 -781 850 -779
rect 856 -775 857 -773
rect 856 -781 857 -779
rect 863 -775 864 -773
rect 863 -781 864 -779
rect 870 -775 871 -773
rect 870 -781 871 -779
rect 880 -775 881 -773
rect 877 -781 878 -779
rect 884 -775 885 -773
rect 884 -781 885 -779
rect 891 -775 892 -773
rect 891 -781 892 -779
rect 898 -775 899 -773
rect 898 -781 899 -779
rect 905 -775 906 -773
rect 905 -781 906 -779
rect 912 -775 913 -773
rect 912 -781 913 -779
rect 919 -775 920 -773
rect 919 -781 920 -779
rect 926 -775 927 -773
rect 926 -781 927 -779
rect 933 -775 934 -773
rect 936 -775 937 -773
rect 936 -781 937 -779
rect 940 -775 941 -773
rect 940 -781 941 -779
rect 950 -775 951 -773
rect 947 -781 948 -779
rect 954 -775 955 -773
rect 957 -781 958 -779
rect 961 -775 962 -773
rect 961 -781 962 -779
rect 968 -775 969 -773
rect 968 -781 969 -779
rect 975 -775 976 -773
rect 975 -781 976 -779
rect 982 -775 983 -773
rect 982 -781 983 -779
rect 989 -775 990 -773
rect 989 -781 990 -779
rect 996 -775 997 -773
rect 996 -781 997 -779
rect 1003 -775 1004 -773
rect 1003 -781 1004 -779
rect 1010 -781 1011 -779
rect 1031 -775 1032 -773
rect 1031 -781 1032 -779
rect 1122 -775 1123 -773
rect 1122 -781 1123 -779
rect 2 -862 3 -860
rect 2 -868 3 -866
rect 12 -868 13 -866
rect 16 -862 17 -860
rect 16 -868 17 -866
rect 23 -862 24 -860
rect 23 -868 24 -866
rect 30 -862 31 -860
rect 30 -868 31 -866
rect 37 -862 38 -860
rect 40 -862 41 -860
rect 44 -862 45 -860
rect 44 -868 45 -866
rect 51 -862 52 -860
rect 51 -868 52 -866
rect 58 -862 59 -860
rect 58 -868 59 -866
rect 65 -862 66 -860
rect 65 -868 66 -866
rect 75 -862 76 -860
rect 72 -868 73 -866
rect 75 -868 76 -866
rect 82 -862 83 -860
rect 79 -868 80 -866
rect 82 -868 83 -866
rect 86 -862 87 -860
rect 86 -868 87 -866
rect 93 -862 94 -860
rect 93 -868 94 -866
rect 100 -862 101 -860
rect 100 -868 101 -866
rect 107 -862 108 -860
rect 107 -868 108 -866
rect 114 -862 115 -860
rect 114 -868 115 -866
rect 121 -862 122 -860
rect 121 -868 122 -866
rect 128 -862 129 -860
rect 128 -868 129 -866
rect 135 -862 136 -860
rect 135 -868 136 -866
rect 142 -862 143 -860
rect 142 -868 143 -866
rect 149 -862 150 -860
rect 149 -868 150 -866
rect 156 -862 157 -860
rect 156 -868 157 -866
rect 163 -862 164 -860
rect 163 -868 164 -866
rect 170 -862 171 -860
rect 170 -868 171 -866
rect 177 -862 178 -860
rect 177 -868 178 -866
rect 184 -862 185 -860
rect 184 -868 185 -866
rect 194 -862 195 -860
rect 191 -868 192 -866
rect 194 -868 195 -866
rect 198 -862 199 -860
rect 198 -868 199 -866
rect 205 -862 206 -860
rect 205 -868 206 -866
rect 212 -862 213 -860
rect 212 -868 213 -866
rect 219 -862 220 -860
rect 222 -862 223 -860
rect 222 -868 223 -866
rect 226 -862 227 -860
rect 226 -868 227 -866
rect 229 -868 230 -866
rect 233 -862 234 -860
rect 233 -868 234 -866
rect 240 -862 241 -860
rect 240 -868 241 -866
rect 247 -862 248 -860
rect 247 -868 248 -866
rect 254 -862 255 -860
rect 254 -868 255 -866
rect 261 -862 262 -860
rect 268 -862 269 -860
rect 268 -868 269 -866
rect 275 -862 276 -860
rect 275 -868 276 -866
rect 282 -862 283 -860
rect 282 -868 283 -866
rect 289 -862 290 -860
rect 289 -868 290 -866
rect 296 -862 297 -860
rect 296 -868 297 -866
rect 303 -862 304 -860
rect 303 -868 304 -866
rect 310 -862 311 -860
rect 310 -868 311 -866
rect 317 -862 318 -860
rect 317 -868 318 -866
rect 324 -862 325 -860
rect 327 -862 328 -860
rect 324 -868 325 -866
rect 331 -862 332 -860
rect 331 -868 332 -866
rect 338 -862 339 -860
rect 341 -862 342 -860
rect 338 -868 339 -866
rect 341 -868 342 -866
rect 345 -862 346 -860
rect 345 -868 346 -866
rect 352 -862 353 -860
rect 355 -862 356 -860
rect 352 -868 353 -866
rect 355 -868 356 -866
rect 359 -862 360 -860
rect 359 -868 360 -866
rect 366 -862 367 -860
rect 366 -868 367 -866
rect 373 -862 374 -860
rect 373 -868 374 -866
rect 383 -862 384 -860
rect 380 -868 381 -866
rect 383 -868 384 -866
rect 387 -862 388 -860
rect 387 -868 388 -866
rect 394 -862 395 -860
rect 394 -868 395 -866
rect 397 -868 398 -866
rect 401 -862 402 -860
rect 401 -868 402 -866
rect 408 -862 409 -860
rect 408 -868 409 -866
rect 415 -862 416 -860
rect 415 -868 416 -866
rect 422 -862 423 -860
rect 422 -868 423 -866
rect 429 -868 430 -866
rect 432 -868 433 -866
rect 436 -862 437 -860
rect 436 -868 437 -866
rect 443 -862 444 -860
rect 443 -868 444 -866
rect 450 -862 451 -860
rect 453 -862 454 -860
rect 450 -868 451 -866
rect 453 -868 454 -866
rect 457 -862 458 -860
rect 457 -868 458 -866
rect 464 -862 465 -860
rect 464 -868 465 -866
rect 471 -862 472 -860
rect 471 -868 472 -866
rect 478 -862 479 -860
rect 481 -862 482 -860
rect 481 -868 482 -866
rect 485 -862 486 -860
rect 485 -868 486 -866
rect 492 -862 493 -860
rect 492 -868 493 -866
rect 499 -862 500 -860
rect 502 -862 503 -860
rect 499 -868 500 -866
rect 506 -862 507 -860
rect 506 -868 507 -866
rect 513 -862 514 -860
rect 513 -868 514 -866
rect 520 -862 521 -860
rect 520 -868 521 -866
rect 527 -862 528 -860
rect 527 -868 528 -866
rect 534 -862 535 -860
rect 534 -868 535 -866
rect 541 -862 542 -860
rect 541 -868 542 -866
rect 544 -868 545 -866
rect 548 -862 549 -860
rect 548 -868 549 -866
rect 555 -862 556 -860
rect 555 -868 556 -866
rect 558 -868 559 -866
rect 565 -862 566 -860
rect 562 -868 563 -866
rect 565 -868 566 -866
rect 569 -862 570 -860
rect 569 -868 570 -866
rect 576 -862 577 -860
rect 579 -862 580 -860
rect 576 -868 577 -866
rect 579 -868 580 -866
rect 583 -862 584 -860
rect 583 -868 584 -866
rect 593 -862 594 -860
rect 590 -868 591 -866
rect 593 -868 594 -866
rect 597 -862 598 -860
rect 597 -868 598 -866
rect 604 -862 605 -860
rect 607 -862 608 -860
rect 604 -868 605 -866
rect 611 -862 612 -860
rect 614 -862 615 -860
rect 611 -868 612 -866
rect 614 -868 615 -866
rect 618 -862 619 -860
rect 618 -868 619 -866
rect 625 -862 626 -860
rect 625 -868 626 -866
rect 632 -862 633 -860
rect 635 -862 636 -860
rect 632 -868 633 -866
rect 635 -868 636 -866
rect 639 -862 640 -860
rect 639 -868 640 -866
rect 646 -862 647 -860
rect 646 -868 647 -866
rect 653 -862 654 -860
rect 656 -862 657 -860
rect 660 -862 661 -860
rect 660 -868 661 -866
rect 667 -862 668 -860
rect 667 -868 668 -866
rect 674 -862 675 -860
rect 674 -868 675 -866
rect 681 -862 682 -860
rect 681 -868 682 -866
rect 688 -862 689 -860
rect 688 -868 689 -866
rect 695 -862 696 -860
rect 695 -868 696 -866
rect 702 -862 703 -860
rect 702 -868 703 -866
rect 709 -862 710 -860
rect 709 -868 710 -866
rect 716 -862 717 -860
rect 716 -868 717 -866
rect 723 -862 724 -860
rect 723 -868 724 -866
rect 730 -862 731 -860
rect 730 -868 731 -866
rect 737 -862 738 -860
rect 737 -868 738 -866
rect 744 -862 745 -860
rect 744 -868 745 -866
rect 751 -862 752 -860
rect 751 -868 752 -866
rect 758 -862 759 -860
rect 758 -868 759 -866
rect 765 -862 766 -860
rect 768 -862 769 -860
rect 768 -868 769 -866
rect 772 -862 773 -860
rect 772 -868 773 -866
rect 779 -862 780 -860
rect 779 -868 780 -866
rect 786 -862 787 -860
rect 786 -868 787 -866
rect 793 -862 794 -860
rect 793 -868 794 -866
rect 800 -862 801 -860
rect 800 -868 801 -866
rect 807 -862 808 -860
rect 807 -868 808 -866
rect 814 -862 815 -860
rect 814 -868 815 -866
rect 821 -862 822 -860
rect 821 -868 822 -866
rect 828 -862 829 -860
rect 828 -868 829 -866
rect 835 -862 836 -860
rect 835 -868 836 -866
rect 842 -862 843 -860
rect 842 -868 843 -866
rect 849 -862 850 -860
rect 849 -868 850 -866
rect 856 -862 857 -860
rect 856 -868 857 -866
rect 863 -862 864 -860
rect 866 -862 867 -860
rect 870 -862 871 -860
rect 870 -868 871 -866
rect 877 -862 878 -860
rect 877 -868 878 -866
rect 884 -862 885 -860
rect 884 -868 885 -866
rect 891 -862 892 -860
rect 891 -868 892 -866
rect 898 -862 899 -860
rect 898 -868 899 -866
rect 905 -862 906 -860
rect 905 -868 906 -866
rect 912 -862 913 -860
rect 912 -868 913 -866
rect 919 -862 920 -860
rect 919 -868 920 -866
rect 926 -862 927 -860
rect 926 -868 927 -866
rect 933 -862 934 -860
rect 933 -868 934 -866
rect 940 -862 941 -860
rect 940 -868 941 -866
rect 947 -862 948 -860
rect 947 -868 948 -866
rect 954 -862 955 -860
rect 954 -868 955 -866
rect 961 -862 962 -860
rect 961 -868 962 -866
rect 968 -862 969 -860
rect 968 -868 969 -866
rect 975 -862 976 -860
rect 975 -868 976 -866
rect 982 -862 983 -860
rect 982 -868 983 -866
rect 989 -862 990 -860
rect 989 -868 990 -866
rect 996 -862 997 -860
rect 996 -868 997 -866
rect 1003 -862 1004 -860
rect 1003 -868 1004 -866
rect 1010 -862 1011 -860
rect 1010 -868 1011 -866
rect 1017 -862 1018 -860
rect 1017 -868 1018 -866
rect 1024 -862 1025 -860
rect 1024 -868 1025 -866
rect 1031 -862 1032 -860
rect 1031 -868 1032 -866
rect 1038 -862 1039 -860
rect 1038 -868 1039 -866
rect 1045 -862 1046 -860
rect 1045 -868 1046 -866
rect 1052 -862 1053 -860
rect 1052 -868 1053 -866
rect 1059 -862 1060 -860
rect 1059 -868 1060 -866
rect 1066 -862 1067 -860
rect 1066 -868 1067 -866
rect 1073 -862 1074 -860
rect 1073 -868 1074 -866
rect 1080 -862 1081 -860
rect 1080 -868 1081 -866
rect 1087 -862 1088 -860
rect 1087 -868 1088 -866
rect 1094 -862 1095 -860
rect 1097 -868 1098 -866
rect 1101 -862 1102 -860
rect 1101 -868 1102 -866
rect 1108 -862 1109 -860
rect 1108 -868 1109 -866
rect 1115 -862 1116 -860
rect 1115 -868 1116 -866
rect 1122 -862 1123 -860
rect 1122 -868 1123 -866
rect 1129 -868 1130 -866
rect 1139 -862 1140 -860
rect 1136 -868 1137 -866
rect 1143 -862 1144 -860
rect 1143 -868 1144 -866
rect 1150 -862 1151 -860
rect 1153 -862 1154 -860
rect 2 -969 3 -967
rect 9 -963 10 -961
rect 9 -969 10 -967
rect 16 -963 17 -961
rect 16 -969 17 -967
rect 23 -963 24 -961
rect 23 -969 24 -967
rect 30 -963 31 -961
rect 30 -969 31 -967
rect 37 -963 38 -961
rect 37 -969 38 -967
rect 44 -963 45 -961
rect 44 -969 45 -967
rect 51 -963 52 -961
rect 51 -969 52 -967
rect 58 -963 59 -961
rect 58 -969 59 -967
rect 65 -963 66 -961
rect 65 -969 66 -967
rect 68 -969 69 -967
rect 72 -963 73 -961
rect 75 -963 76 -961
rect 72 -969 73 -967
rect 75 -969 76 -967
rect 79 -963 80 -961
rect 82 -963 83 -961
rect 82 -969 83 -967
rect 86 -963 87 -961
rect 86 -969 87 -967
rect 93 -963 94 -961
rect 93 -969 94 -967
rect 100 -963 101 -961
rect 100 -969 101 -967
rect 107 -963 108 -961
rect 107 -969 108 -967
rect 114 -963 115 -961
rect 114 -969 115 -967
rect 121 -963 122 -961
rect 121 -969 122 -967
rect 128 -963 129 -961
rect 128 -969 129 -967
rect 135 -963 136 -961
rect 135 -969 136 -967
rect 142 -963 143 -961
rect 142 -969 143 -967
rect 149 -963 150 -961
rect 152 -963 153 -961
rect 156 -963 157 -961
rect 156 -969 157 -967
rect 163 -963 164 -961
rect 163 -969 164 -967
rect 170 -963 171 -961
rect 170 -969 171 -967
rect 177 -963 178 -961
rect 177 -969 178 -967
rect 184 -963 185 -961
rect 184 -969 185 -967
rect 191 -963 192 -961
rect 191 -969 192 -967
rect 198 -963 199 -961
rect 198 -969 199 -967
rect 205 -963 206 -961
rect 205 -969 206 -967
rect 212 -963 213 -961
rect 212 -969 213 -967
rect 219 -963 220 -961
rect 219 -969 220 -967
rect 226 -963 227 -961
rect 226 -969 227 -967
rect 233 -963 234 -961
rect 233 -969 234 -967
rect 240 -963 241 -961
rect 240 -969 241 -967
rect 247 -963 248 -961
rect 247 -969 248 -967
rect 254 -963 255 -961
rect 254 -969 255 -967
rect 261 -963 262 -961
rect 261 -969 262 -967
rect 268 -963 269 -961
rect 268 -969 269 -967
rect 275 -963 276 -961
rect 275 -969 276 -967
rect 282 -969 283 -967
rect 285 -969 286 -967
rect 289 -963 290 -961
rect 289 -969 290 -967
rect 299 -963 300 -961
rect 303 -963 304 -961
rect 303 -969 304 -967
rect 306 -969 307 -967
rect 310 -963 311 -961
rect 310 -969 311 -967
rect 317 -963 318 -961
rect 317 -969 318 -967
rect 324 -963 325 -961
rect 324 -969 325 -967
rect 331 -963 332 -961
rect 331 -969 332 -967
rect 338 -963 339 -961
rect 338 -969 339 -967
rect 345 -963 346 -961
rect 345 -969 346 -967
rect 352 -963 353 -961
rect 352 -969 353 -967
rect 359 -963 360 -961
rect 362 -963 363 -961
rect 362 -969 363 -967
rect 366 -963 367 -961
rect 366 -969 367 -967
rect 373 -963 374 -961
rect 373 -969 374 -967
rect 380 -963 381 -961
rect 380 -969 381 -967
rect 387 -963 388 -961
rect 387 -969 388 -967
rect 394 -963 395 -961
rect 394 -969 395 -967
rect 401 -963 402 -961
rect 401 -969 402 -967
rect 408 -963 409 -961
rect 408 -969 409 -967
rect 415 -963 416 -961
rect 418 -963 419 -961
rect 415 -969 416 -967
rect 418 -969 419 -967
rect 422 -963 423 -961
rect 422 -969 423 -967
rect 429 -963 430 -961
rect 429 -969 430 -967
rect 439 -963 440 -961
rect 436 -969 437 -967
rect 439 -969 440 -967
rect 443 -963 444 -961
rect 446 -963 447 -961
rect 446 -969 447 -967
rect 450 -963 451 -961
rect 450 -969 451 -967
rect 457 -963 458 -961
rect 457 -969 458 -967
rect 464 -963 465 -961
rect 467 -969 468 -967
rect 471 -963 472 -961
rect 471 -969 472 -967
rect 474 -969 475 -967
rect 478 -963 479 -961
rect 481 -963 482 -961
rect 478 -969 479 -967
rect 481 -969 482 -967
rect 485 -963 486 -961
rect 485 -969 486 -967
rect 492 -963 493 -961
rect 492 -969 493 -967
rect 502 -963 503 -961
rect 499 -969 500 -967
rect 502 -969 503 -967
rect 506 -963 507 -961
rect 506 -969 507 -967
rect 513 -963 514 -961
rect 513 -969 514 -967
rect 520 -963 521 -961
rect 520 -969 521 -967
rect 527 -963 528 -961
rect 527 -969 528 -967
rect 537 -963 538 -961
rect 534 -969 535 -967
rect 541 -963 542 -961
rect 544 -963 545 -961
rect 544 -969 545 -967
rect 548 -963 549 -961
rect 548 -969 549 -967
rect 555 -963 556 -961
rect 555 -969 556 -967
rect 562 -963 563 -961
rect 562 -969 563 -967
rect 569 -963 570 -961
rect 572 -963 573 -961
rect 569 -969 570 -967
rect 572 -969 573 -967
rect 576 -963 577 -961
rect 579 -963 580 -961
rect 579 -969 580 -967
rect 583 -963 584 -961
rect 583 -969 584 -967
rect 593 -963 594 -961
rect 590 -969 591 -967
rect 593 -969 594 -967
rect 597 -963 598 -961
rect 597 -969 598 -967
rect 604 -963 605 -961
rect 604 -969 605 -967
rect 614 -963 615 -961
rect 611 -969 612 -967
rect 614 -969 615 -967
rect 618 -963 619 -961
rect 621 -963 622 -961
rect 618 -969 619 -967
rect 621 -969 622 -967
rect 625 -963 626 -961
rect 625 -969 626 -967
rect 628 -969 629 -967
rect 632 -963 633 -961
rect 635 -969 636 -967
rect 639 -963 640 -961
rect 639 -969 640 -967
rect 646 -963 647 -961
rect 646 -969 647 -967
rect 653 -963 654 -961
rect 653 -969 654 -967
rect 660 -963 661 -961
rect 660 -969 661 -967
rect 667 -963 668 -961
rect 667 -969 668 -967
rect 674 -963 675 -961
rect 674 -969 675 -967
rect 681 -963 682 -961
rect 681 -969 682 -967
rect 688 -963 689 -961
rect 691 -963 692 -961
rect 691 -969 692 -967
rect 698 -963 699 -961
rect 698 -969 699 -967
rect 702 -963 703 -961
rect 702 -969 703 -967
rect 709 -963 710 -961
rect 709 -969 710 -967
rect 716 -963 717 -961
rect 716 -969 717 -967
rect 723 -963 724 -961
rect 723 -969 724 -967
rect 730 -963 731 -961
rect 730 -969 731 -967
rect 737 -963 738 -961
rect 737 -969 738 -967
rect 744 -963 745 -961
rect 744 -969 745 -967
rect 751 -963 752 -961
rect 751 -969 752 -967
rect 758 -963 759 -961
rect 758 -969 759 -967
rect 765 -963 766 -961
rect 765 -969 766 -967
rect 772 -963 773 -961
rect 772 -969 773 -967
rect 779 -963 780 -961
rect 779 -969 780 -967
rect 786 -963 787 -961
rect 786 -969 787 -967
rect 793 -963 794 -961
rect 793 -969 794 -967
rect 800 -963 801 -961
rect 800 -969 801 -967
rect 807 -963 808 -961
rect 807 -969 808 -967
rect 814 -963 815 -961
rect 814 -969 815 -967
rect 821 -963 822 -961
rect 821 -969 822 -967
rect 828 -963 829 -961
rect 828 -969 829 -967
rect 835 -963 836 -961
rect 835 -969 836 -967
rect 842 -963 843 -961
rect 842 -969 843 -967
rect 849 -963 850 -961
rect 849 -969 850 -967
rect 856 -969 857 -967
rect 859 -969 860 -967
rect 863 -963 864 -961
rect 863 -969 864 -967
rect 870 -963 871 -961
rect 870 -969 871 -967
rect 877 -963 878 -961
rect 877 -969 878 -967
rect 884 -963 885 -961
rect 884 -969 885 -967
rect 891 -963 892 -961
rect 891 -969 892 -967
rect 898 -963 899 -961
rect 898 -969 899 -967
rect 905 -963 906 -961
rect 905 -969 906 -967
rect 912 -963 913 -961
rect 912 -969 913 -967
rect 919 -963 920 -961
rect 919 -969 920 -967
rect 926 -963 927 -961
rect 926 -969 927 -967
rect 933 -963 934 -961
rect 933 -969 934 -967
rect 940 -963 941 -961
rect 940 -969 941 -967
rect 947 -963 948 -961
rect 947 -969 948 -967
rect 954 -963 955 -961
rect 954 -969 955 -967
rect 961 -963 962 -961
rect 961 -969 962 -967
rect 968 -963 969 -961
rect 968 -969 969 -967
rect 975 -963 976 -961
rect 975 -969 976 -967
rect 982 -963 983 -961
rect 982 -969 983 -967
rect 989 -963 990 -961
rect 989 -969 990 -967
rect 996 -963 997 -961
rect 996 -969 997 -967
rect 1003 -963 1004 -961
rect 1003 -969 1004 -967
rect 1010 -963 1011 -961
rect 1010 -969 1011 -967
rect 1017 -963 1018 -961
rect 1017 -969 1018 -967
rect 1024 -963 1025 -961
rect 1024 -969 1025 -967
rect 1031 -963 1032 -961
rect 1031 -969 1032 -967
rect 1038 -963 1039 -961
rect 1038 -969 1039 -967
rect 1045 -963 1046 -961
rect 1045 -969 1046 -967
rect 1052 -963 1053 -961
rect 1052 -969 1053 -967
rect 1059 -963 1060 -961
rect 1059 -969 1060 -967
rect 1066 -963 1067 -961
rect 1066 -969 1067 -967
rect 1073 -963 1074 -961
rect 1073 -969 1074 -967
rect 1080 -963 1081 -961
rect 1080 -969 1081 -967
rect 1087 -963 1088 -961
rect 1087 -969 1088 -967
rect 1094 -963 1095 -961
rect 1094 -969 1095 -967
rect 1101 -963 1102 -961
rect 1101 -969 1102 -967
rect 1108 -963 1109 -961
rect 1108 -969 1109 -967
rect 1115 -963 1116 -961
rect 1115 -969 1116 -967
rect 1122 -963 1123 -961
rect 1122 -969 1123 -967
rect 1129 -963 1130 -961
rect 1129 -969 1130 -967
rect 1136 -963 1137 -961
rect 1136 -969 1137 -967
rect 1143 -963 1144 -961
rect 1143 -969 1144 -967
rect 1150 -963 1151 -961
rect 1150 -969 1151 -967
rect 1157 -963 1158 -961
rect 1157 -969 1158 -967
rect 2 -1078 3 -1076
rect 9 -1078 10 -1076
rect 9 -1084 10 -1082
rect 16 -1078 17 -1076
rect 16 -1084 17 -1082
rect 23 -1078 24 -1076
rect 23 -1084 24 -1082
rect 30 -1078 31 -1076
rect 30 -1084 31 -1082
rect 37 -1078 38 -1076
rect 37 -1084 38 -1082
rect 44 -1078 45 -1076
rect 44 -1084 45 -1082
rect 51 -1078 52 -1076
rect 51 -1084 52 -1082
rect 54 -1084 55 -1082
rect 58 -1078 59 -1076
rect 58 -1084 59 -1082
rect 68 -1078 69 -1076
rect 65 -1084 66 -1082
rect 68 -1084 69 -1082
rect 72 -1078 73 -1076
rect 72 -1084 73 -1082
rect 82 -1078 83 -1076
rect 79 -1084 80 -1082
rect 86 -1078 87 -1076
rect 86 -1084 87 -1082
rect 93 -1078 94 -1076
rect 93 -1084 94 -1082
rect 100 -1084 101 -1082
rect 103 -1084 104 -1082
rect 107 -1078 108 -1076
rect 110 -1084 111 -1082
rect 114 -1078 115 -1076
rect 114 -1084 115 -1082
rect 121 -1078 122 -1076
rect 121 -1084 122 -1082
rect 128 -1078 129 -1076
rect 128 -1084 129 -1082
rect 135 -1078 136 -1076
rect 135 -1084 136 -1082
rect 142 -1078 143 -1076
rect 142 -1084 143 -1082
rect 149 -1078 150 -1076
rect 149 -1084 150 -1082
rect 156 -1078 157 -1076
rect 156 -1084 157 -1082
rect 163 -1078 164 -1076
rect 166 -1078 167 -1076
rect 166 -1084 167 -1082
rect 170 -1078 171 -1076
rect 170 -1084 171 -1082
rect 177 -1078 178 -1076
rect 177 -1084 178 -1082
rect 184 -1078 185 -1076
rect 184 -1084 185 -1082
rect 191 -1078 192 -1076
rect 194 -1078 195 -1076
rect 191 -1084 192 -1082
rect 198 -1078 199 -1076
rect 198 -1084 199 -1082
rect 205 -1078 206 -1076
rect 205 -1084 206 -1082
rect 212 -1084 213 -1082
rect 215 -1084 216 -1082
rect 219 -1078 220 -1076
rect 219 -1084 220 -1082
rect 229 -1078 230 -1076
rect 226 -1084 227 -1082
rect 233 -1078 234 -1076
rect 233 -1084 234 -1082
rect 240 -1078 241 -1076
rect 240 -1084 241 -1082
rect 247 -1078 248 -1076
rect 247 -1084 248 -1082
rect 254 -1078 255 -1076
rect 254 -1084 255 -1082
rect 261 -1078 262 -1076
rect 261 -1084 262 -1082
rect 268 -1078 269 -1076
rect 271 -1078 272 -1076
rect 275 -1078 276 -1076
rect 275 -1084 276 -1082
rect 282 -1078 283 -1076
rect 285 -1084 286 -1082
rect 289 -1078 290 -1076
rect 289 -1084 290 -1082
rect 296 -1078 297 -1076
rect 296 -1084 297 -1082
rect 303 -1078 304 -1076
rect 303 -1084 304 -1082
rect 310 -1078 311 -1076
rect 310 -1084 311 -1082
rect 317 -1078 318 -1076
rect 317 -1084 318 -1082
rect 324 -1078 325 -1076
rect 324 -1084 325 -1082
rect 331 -1078 332 -1076
rect 331 -1084 332 -1082
rect 338 -1078 339 -1076
rect 338 -1084 339 -1082
rect 345 -1078 346 -1076
rect 345 -1084 346 -1082
rect 352 -1078 353 -1076
rect 352 -1084 353 -1082
rect 359 -1078 360 -1076
rect 359 -1084 360 -1082
rect 366 -1078 367 -1076
rect 366 -1084 367 -1082
rect 373 -1078 374 -1076
rect 373 -1084 374 -1082
rect 380 -1078 381 -1076
rect 380 -1084 381 -1082
rect 387 -1078 388 -1076
rect 390 -1078 391 -1076
rect 387 -1084 388 -1082
rect 390 -1084 391 -1082
rect 394 -1078 395 -1076
rect 397 -1078 398 -1076
rect 394 -1084 395 -1082
rect 397 -1084 398 -1082
rect 401 -1078 402 -1076
rect 401 -1084 402 -1082
rect 408 -1078 409 -1076
rect 408 -1084 409 -1082
rect 415 -1078 416 -1076
rect 415 -1084 416 -1082
rect 422 -1078 423 -1076
rect 422 -1084 423 -1082
rect 429 -1078 430 -1076
rect 429 -1084 430 -1082
rect 436 -1078 437 -1076
rect 436 -1084 437 -1082
rect 443 -1078 444 -1076
rect 443 -1084 444 -1082
rect 450 -1078 451 -1076
rect 450 -1084 451 -1082
rect 457 -1078 458 -1076
rect 457 -1084 458 -1082
rect 464 -1078 465 -1076
rect 464 -1084 465 -1082
rect 471 -1078 472 -1076
rect 471 -1084 472 -1082
rect 478 -1078 479 -1076
rect 478 -1084 479 -1082
rect 488 -1078 489 -1076
rect 485 -1084 486 -1082
rect 488 -1084 489 -1082
rect 492 -1078 493 -1076
rect 495 -1078 496 -1076
rect 495 -1084 496 -1082
rect 502 -1078 503 -1076
rect 499 -1084 500 -1082
rect 502 -1084 503 -1082
rect 506 -1078 507 -1076
rect 506 -1084 507 -1082
rect 513 -1078 514 -1076
rect 513 -1084 514 -1082
rect 520 -1078 521 -1076
rect 520 -1084 521 -1082
rect 527 -1078 528 -1076
rect 527 -1084 528 -1082
rect 534 -1078 535 -1076
rect 534 -1084 535 -1082
rect 541 -1078 542 -1076
rect 541 -1084 542 -1082
rect 544 -1084 545 -1082
rect 548 -1078 549 -1076
rect 548 -1084 549 -1082
rect 555 -1078 556 -1076
rect 558 -1078 559 -1076
rect 555 -1084 556 -1082
rect 558 -1084 559 -1082
rect 562 -1078 563 -1076
rect 562 -1084 563 -1082
rect 569 -1078 570 -1076
rect 572 -1078 573 -1076
rect 572 -1084 573 -1082
rect 576 -1078 577 -1076
rect 576 -1084 577 -1082
rect 583 -1078 584 -1076
rect 583 -1084 584 -1082
rect 586 -1084 587 -1082
rect 590 -1078 591 -1076
rect 590 -1084 591 -1082
rect 600 -1078 601 -1076
rect 597 -1084 598 -1082
rect 604 -1078 605 -1076
rect 607 -1078 608 -1076
rect 604 -1084 605 -1082
rect 607 -1084 608 -1082
rect 611 -1078 612 -1076
rect 611 -1084 612 -1082
rect 618 -1078 619 -1076
rect 618 -1084 619 -1082
rect 625 -1078 626 -1076
rect 625 -1084 626 -1082
rect 632 -1078 633 -1076
rect 635 -1078 636 -1076
rect 632 -1084 633 -1082
rect 635 -1084 636 -1082
rect 639 -1078 640 -1076
rect 639 -1084 640 -1082
rect 646 -1078 647 -1076
rect 646 -1084 647 -1082
rect 653 -1078 654 -1076
rect 653 -1084 654 -1082
rect 660 -1078 661 -1076
rect 660 -1084 661 -1082
rect 667 -1078 668 -1076
rect 667 -1084 668 -1082
rect 674 -1078 675 -1076
rect 674 -1084 675 -1082
rect 681 -1078 682 -1076
rect 681 -1084 682 -1082
rect 684 -1084 685 -1082
rect 688 -1078 689 -1076
rect 688 -1084 689 -1082
rect 695 -1078 696 -1076
rect 695 -1084 696 -1082
rect 702 -1078 703 -1076
rect 702 -1084 703 -1082
rect 709 -1078 710 -1076
rect 709 -1084 710 -1082
rect 716 -1078 717 -1076
rect 716 -1084 717 -1082
rect 723 -1078 724 -1076
rect 726 -1078 727 -1076
rect 730 -1078 731 -1076
rect 730 -1084 731 -1082
rect 737 -1078 738 -1076
rect 740 -1078 741 -1076
rect 737 -1084 738 -1082
rect 744 -1078 745 -1076
rect 744 -1084 745 -1082
rect 751 -1078 752 -1076
rect 751 -1084 752 -1082
rect 758 -1078 759 -1076
rect 758 -1084 759 -1082
rect 765 -1078 766 -1076
rect 765 -1084 766 -1082
rect 772 -1078 773 -1076
rect 772 -1084 773 -1082
rect 779 -1078 780 -1076
rect 779 -1084 780 -1082
rect 786 -1078 787 -1076
rect 786 -1084 787 -1082
rect 793 -1078 794 -1076
rect 793 -1084 794 -1082
rect 800 -1078 801 -1076
rect 800 -1084 801 -1082
rect 807 -1078 808 -1076
rect 807 -1084 808 -1082
rect 814 -1084 815 -1082
rect 817 -1084 818 -1082
rect 821 -1078 822 -1076
rect 821 -1084 822 -1082
rect 828 -1078 829 -1076
rect 828 -1084 829 -1082
rect 835 -1078 836 -1076
rect 835 -1084 836 -1082
rect 842 -1078 843 -1076
rect 842 -1084 843 -1082
rect 849 -1078 850 -1076
rect 849 -1084 850 -1082
rect 856 -1078 857 -1076
rect 856 -1084 857 -1082
rect 863 -1078 864 -1076
rect 863 -1084 864 -1082
rect 870 -1078 871 -1076
rect 870 -1084 871 -1082
rect 877 -1078 878 -1076
rect 877 -1084 878 -1082
rect 884 -1078 885 -1076
rect 884 -1084 885 -1082
rect 891 -1078 892 -1076
rect 891 -1084 892 -1082
rect 898 -1078 899 -1076
rect 898 -1084 899 -1082
rect 905 -1078 906 -1076
rect 905 -1084 906 -1082
rect 912 -1078 913 -1076
rect 912 -1084 913 -1082
rect 919 -1078 920 -1076
rect 919 -1084 920 -1082
rect 926 -1078 927 -1076
rect 926 -1084 927 -1082
rect 933 -1078 934 -1076
rect 933 -1084 934 -1082
rect 940 -1078 941 -1076
rect 940 -1084 941 -1082
rect 947 -1078 948 -1076
rect 947 -1084 948 -1082
rect 954 -1078 955 -1076
rect 954 -1084 955 -1082
rect 961 -1078 962 -1076
rect 961 -1084 962 -1082
rect 968 -1078 969 -1076
rect 968 -1084 969 -1082
rect 975 -1078 976 -1076
rect 975 -1084 976 -1082
rect 982 -1078 983 -1076
rect 982 -1084 983 -1082
rect 989 -1078 990 -1076
rect 989 -1084 990 -1082
rect 996 -1078 997 -1076
rect 996 -1084 997 -1082
rect 1003 -1078 1004 -1076
rect 1003 -1084 1004 -1082
rect 1010 -1078 1011 -1076
rect 1010 -1084 1011 -1082
rect 1017 -1078 1018 -1076
rect 1017 -1084 1018 -1082
rect 1024 -1078 1025 -1076
rect 1024 -1084 1025 -1082
rect 1031 -1078 1032 -1076
rect 1031 -1084 1032 -1082
rect 1041 -1078 1042 -1076
rect 1038 -1084 1039 -1082
rect 1041 -1084 1042 -1082
rect 1045 -1078 1046 -1076
rect 1045 -1084 1046 -1082
rect 1052 -1078 1053 -1076
rect 1052 -1084 1053 -1082
rect 1059 -1084 1060 -1082
rect 1066 -1078 1067 -1076
rect 1066 -1084 1067 -1082
rect 1073 -1078 1074 -1076
rect 1073 -1084 1074 -1082
rect 1080 -1078 1081 -1076
rect 1080 -1084 1081 -1082
rect 1129 -1078 1130 -1076
rect 1129 -1084 1130 -1082
rect 1143 -1078 1144 -1076
rect 1143 -1084 1144 -1082
rect 5 -1167 6 -1165
rect 9 -1167 10 -1165
rect 9 -1173 10 -1171
rect 16 -1173 17 -1171
rect 19 -1173 20 -1171
rect 23 -1167 24 -1165
rect 23 -1173 24 -1171
rect 30 -1167 31 -1165
rect 30 -1173 31 -1171
rect 37 -1167 38 -1165
rect 40 -1167 41 -1165
rect 37 -1173 38 -1171
rect 44 -1167 45 -1165
rect 44 -1173 45 -1171
rect 51 -1167 52 -1165
rect 51 -1173 52 -1171
rect 61 -1167 62 -1165
rect 58 -1173 59 -1171
rect 61 -1173 62 -1171
rect 65 -1167 66 -1165
rect 65 -1173 66 -1171
rect 72 -1167 73 -1165
rect 72 -1173 73 -1171
rect 79 -1167 80 -1165
rect 79 -1173 80 -1171
rect 86 -1167 87 -1165
rect 86 -1173 87 -1171
rect 93 -1167 94 -1165
rect 93 -1173 94 -1171
rect 100 -1167 101 -1165
rect 100 -1173 101 -1171
rect 107 -1167 108 -1165
rect 107 -1173 108 -1171
rect 114 -1167 115 -1165
rect 114 -1173 115 -1171
rect 121 -1167 122 -1165
rect 121 -1173 122 -1171
rect 128 -1167 129 -1165
rect 128 -1173 129 -1171
rect 135 -1167 136 -1165
rect 135 -1173 136 -1171
rect 142 -1173 143 -1171
rect 145 -1173 146 -1171
rect 152 -1167 153 -1165
rect 152 -1173 153 -1171
rect 156 -1167 157 -1165
rect 156 -1173 157 -1171
rect 163 -1167 164 -1165
rect 163 -1173 164 -1171
rect 170 -1167 171 -1165
rect 170 -1173 171 -1171
rect 177 -1167 178 -1165
rect 177 -1173 178 -1171
rect 184 -1167 185 -1165
rect 184 -1173 185 -1171
rect 191 -1167 192 -1165
rect 191 -1173 192 -1171
rect 198 -1167 199 -1165
rect 198 -1173 199 -1171
rect 205 -1167 206 -1165
rect 205 -1173 206 -1171
rect 212 -1167 213 -1165
rect 212 -1173 213 -1171
rect 219 -1167 220 -1165
rect 222 -1173 223 -1171
rect 226 -1167 227 -1165
rect 226 -1173 227 -1171
rect 233 -1167 234 -1165
rect 233 -1173 234 -1171
rect 240 -1167 241 -1165
rect 240 -1173 241 -1171
rect 247 -1167 248 -1165
rect 247 -1173 248 -1171
rect 254 -1167 255 -1165
rect 254 -1173 255 -1171
rect 261 -1167 262 -1165
rect 261 -1173 262 -1171
rect 268 -1167 269 -1165
rect 268 -1173 269 -1171
rect 275 -1167 276 -1165
rect 275 -1173 276 -1171
rect 282 -1167 283 -1165
rect 282 -1173 283 -1171
rect 285 -1173 286 -1171
rect 289 -1167 290 -1165
rect 289 -1173 290 -1171
rect 296 -1167 297 -1165
rect 296 -1173 297 -1171
rect 303 -1167 304 -1165
rect 303 -1173 304 -1171
rect 313 -1167 314 -1165
rect 310 -1173 311 -1171
rect 313 -1173 314 -1171
rect 317 -1167 318 -1165
rect 317 -1173 318 -1171
rect 324 -1167 325 -1165
rect 324 -1173 325 -1171
rect 331 -1167 332 -1165
rect 331 -1173 332 -1171
rect 338 -1167 339 -1165
rect 338 -1173 339 -1171
rect 345 -1167 346 -1165
rect 348 -1167 349 -1165
rect 345 -1173 346 -1171
rect 348 -1173 349 -1171
rect 352 -1167 353 -1165
rect 355 -1167 356 -1165
rect 352 -1173 353 -1171
rect 355 -1173 356 -1171
rect 359 -1173 360 -1171
rect 362 -1173 363 -1171
rect 366 -1167 367 -1165
rect 366 -1173 367 -1171
rect 373 -1167 374 -1165
rect 373 -1173 374 -1171
rect 380 -1167 381 -1165
rect 383 -1167 384 -1165
rect 380 -1173 381 -1171
rect 383 -1173 384 -1171
rect 387 -1167 388 -1165
rect 387 -1173 388 -1171
rect 394 -1167 395 -1165
rect 394 -1173 395 -1171
rect 401 -1167 402 -1165
rect 401 -1173 402 -1171
rect 408 -1167 409 -1165
rect 411 -1167 412 -1165
rect 415 -1167 416 -1165
rect 418 -1167 419 -1165
rect 415 -1173 416 -1171
rect 418 -1173 419 -1171
rect 422 -1167 423 -1165
rect 422 -1173 423 -1171
rect 429 -1167 430 -1165
rect 429 -1173 430 -1171
rect 436 -1167 437 -1165
rect 436 -1173 437 -1171
rect 443 -1167 444 -1165
rect 443 -1173 444 -1171
rect 450 -1167 451 -1165
rect 450 -1173 451 -1171
rect 457 -1167 458 -1165
rect 457 -1173 458 -1171
rect 464 -1167 465 -1165
rect 467 -1167 468 -1165
rect 464 -1173 465 -1171
rect 467 -1173 468 -1171
rect 471 -1167 472 -1165
rect 471 -1173 472 -1171
rect 481 -1167 482 -1165
rect 478 -1173 479 -1171
rect 481 -1173 482 -1171
rect 485 -1167 486 -1165
rect 485 -1173 486 -1171
rect 492 -1167 493 -1165
rect 492 -1173 493 -1171
rect 499 -1167 500 -1165
rect 502 -1167 503 -1165
rect 499 -1173 500 -1171
rect 502 -1173 503 -1171
rect 506 -1167 507 -1165
rect 506 -1173 507 -1171
rect 513 -1167 514 -1165
rect 513 -1173 514 -1171
rect 520 -1167 521 -1165
rect 523 -1167 524 -1165
rect 523 -1173 524 -1171
rect 527 -1167 528 -1165
rect 527 -1173 528 -1171
rect 534 -1167 535 -1165
rect 534 -1173 535 -1171
rect 541 -1167 542 -1165
rect 541 -1173 542 -1171
rect 548 -1167 549 -1165
rect 548 -1173 549 -1171
rect 555 -1167 556 -1165
rect 558 -1167 559 -1165
rect 555 -1173 556 -1171
rect 558 -1173 559 -1171
rect 565 -1167 566 -1165
rect 562 -1173 563 -1171
rect 569 -1167 570 -1165
rect 569 -1173 570 -1171
rect 576 -1167 577 -1165
rect 576 -1173 577 -1171
rect 583 -1167 584 -1165
rect 583 -1173 584 -1171
rect 590 -1167 591 -1165
rect 590 -1173 591 -1171
rect 597 -1173 598 -1171
rect 600 -1173 601 -1171
rect 604 -1167 605 -1165
rect 604 -1173 605 -1171
rect 611 -1167 612 -1165
rect 611 -1173 612 -1171
rect 618 -1167 619 -1165
rect 618 -1173 619 -1171
rect 625 -1167 626 -1165
rect 625 -1173 626 -1171
rect 632 -1167 633 -1165
rect 632 -1173 633 -1171
rect 639 -1167 640 -1165
rect 639 -1173 640 -1171
rect 646 -1167 647 -1165
rect 646 -1173 647 -1171
rect 653 -1167 654 -1165
rect 653 -1173 654 -1171
rect 660 -1167 661 -1165
rect 660 -1173 661 -1171
rect 667 -1167 668 -1165
rect 667 -1173 668 -1171
rect 674 -1167 675 -1165
rect 674 -1173 675 -1171
rect 681 -1167 682 -1165
rect 681 -1173 682 -1171
rect 691 -1167 692 -1165
rect 688 -1173 689 -1171
rect 695 -1167 696 -1165
rect 695 -1173 696 -1171
rect 702 -1167 703 -1165
rect 702 -1173 703 -1171
rect 709 -1167 710 -1165
rect 709 -1173 710 -1171
rect 716 -1167 717 -1165
rect 716 -1173 717 -1171
rect 723 -1167 724 -1165
rect 723 -1173 724 -1171
rect 730 -1167 731 -1165
rect 733 -1167 734 -1165
rect 730 -1173 731 -1171
rect 733 -1173 734 -1171
rect 740 -1167 741 -1165
rect 737 -1173 738 -1171
rect 744 -1167 745 -1165
rect 744 -1173 745 -1171
rect 751 -1167 752 -1165
rect 751 -1173 752 -1171
rect 758 -1167 759 -1165
rect 758 -1173 759 -1171
rect 765 -1167 766 -1165
rect 765 -1173 766 -1171
rect 772 -1167 773 -1165
rect 772 -1173 773 -1171
rect 779 -1167 780 -1165
rect 779 -1173 780 -1171
rect 786 -1167 787 -1165
rect 789 -1167 790 -1165
rect 786 -1173 787 -1171
rect 789 -1173 790 -1171
rect 793 -1167 794 -1165
rect 793 -1173 794 -1171
rect 800 -1167 801 -1165
rect 800 -1173 801 -1171
rect 807 -1167 808 -1165
rect 807 -1173 808 -1171
rect 814 -1167 815 -1165
rect 814 -1173 815 -1171
rect 821 -1167 822 -1165
rect 821 -1173 822 -1171
rect 828 -1167 829 -1165
rect 828 -1173 829 -1171
rect 835 -1167 836 -1165
rect 835 -1173 836 -1171
rect 842 -1167 843 -1165
rect 842 -1173 843 -1171
rect 849 -1167 850 -1165
rect 849 -1173 850 -1171
rect 856 -1167 857 -1165
rect 859 -1173 860 -1171
rect 863 -1167 864 -1165
rect 863 -1173 864 -1171
rect 870 -1167 871 -1165
rect 870 -1173 871 -1171
rect 877 -1167 878 -1165
rect 877 -1173 878 -1171
rect 884 -1167 885 -1165
rect 884 -1173 885 -1171
rect 891 -1167 892 -1165
rect 891 -1173 892 -1171
rect 898 -1167 899 -1165
rect 898 -1173 899 -1171
rect 905 -1167 906 -1165
rect 905 -1173 906 -1171
rect 912 -1167 913 -1165
rect 912 -1173 913 -1171
rect 919 -1167 920 -1165
rect 919 -1173 920 -1171
rect 926 -1167 927 -1165
rect 926 -1173 927 -1171
rect 933 -1167 934 -1165
rect 933 -1173 934 -1171
rect 940 -1167 941 -1165
rect 940 -1173 941 -1171
rect 947 -1167 948 -1165
rect 947 -1173 948 -1171
rect 954 -1167 955 -1165
rect 954 -1173 955 -1171
rect 961 -1167 962 -1165
rect 961 -1173 962 -1171
rect 968 -1167 969 -1165
rect 968 -1173 969 -1171
rect 975 -1167 976 -1165
rect 975 -1173 976 -1171
rect 982 -1167 983 -1165
rect 982 -1173 983 -1171
rect 989 -1167 990 -1165
rect 989 -1173 990 -1171
rect 996 -1167 997 -1165
rect 996 -1173 997 -1171
rect 1003 -1167 1004 -1165
rect 1003 -1173 1004 -1171
rect 1010 -1167 1011 -1165
rect 1010 -1173 1011 -1171
rect 1017 -1167 1018 -1165
rect 1017 -1173 1018 -1171
rect 1024 -1167 1025 -1165
rect 1024 -1173 1025 -1171
rect 1031 -1167 1032 -1165
rect 1031 -1173 1032 -1171
rect 1038 -1167 1039 -1165
rect 1041 -1167 1042 -1165
rect 1038 -1173 1039 -1171
rect 1041 -1173 1042 -1171
rect 1045 -1167 1046 -1165
rect 1045 -1173 1046 -1171
rect 1052 -1167 1053 -1165
rect 1052 -1173 1053 -1171
rect 1059 -1167 1060 -1165
rect 1059 -1173 1060 -1171
rect 1066 -1167 1067 -1165
rect 1066 -1173 1067 -1171
rect 1073 -1167 1074 -1165
rect 1076 -1167 1077 -1165
rect 1122 -1167 1123 -1165
rect 1122 -1173 1123 -1171
rect 1150 -1167 1151 -1165
rect 1150 -1173 1151 -1171
rect 2 -1250 3 -1248
rect 2 -1256 3 -1254
rect 9 -1250 10 -1248
rect 9 -1256 10 -1254
rect 16 -1250 17 -1248
rect 16 -1256 17 -1254
rect 23 -1250 24 -1248
rect 30 -1250 31 -1248
rect 30 -1256 31 -1254
rect 37 -1250 38 -1248
rect 37 -1256 38 -1254
rect 44 -1250 45 -1248
rect 44 -1256 45 -1254
rect 47 -1256 48 -1254
rect 51 -1250 52 -1248
rect 51 -1256 52 -1254
rect 58 -1250 59 -1248
rect 58 -1256 59 -1254
rect 65 -1250 66 -1248
rect 65 -1256 66 -1254
rect 72 -1256 73 -1254
rect 79 -1250 80 -1248
rect 79 -1256 80 -1254
rect 86 -1250 87 -1248
rect 86 -1256 87 -1254
rect 93 -1250 94 -1248
rect 96 -1250 97 -1248
rect 100 -1250 101 -1248
rect 100 -1256 101 -1254
rect 107 -1250 108 -1248
rect 107 -1256 108 -1254
rect 114 -1250 115 -1248
rect 114 -1256 115 -1254
rect 121 -1250 122 -1248
rect 121 -1256 122 -1254
rect 128 -1250 129 -1248
rect 128 -1256 129 -1254
rect 135 -1250 136 -1248
rect 135 -1256 136 -1254
rect 142 -1250 143 -1248
rect 142 -1256 143 -1254
rect 149 -1250 150 -1248
rect 149 -1256 150 -1254
rect 159 -1250 160 -1248
rect 156 -1256 157 -1254
rect 159 -1256 160 -1254
rect 163 -1250 164 -1248
rect 163 -1256 164 -1254
rect 170 -1250 171 -1248
rect 170 -1256 171 -1254
rect 177 -1250 178 -1248
rect 177 -1256 178 -1254
rect 184 -1250 185 -1248
rect 184 -1256 185 -1254
rect 187 -1256 188 -1254
rect 194 -1250 195 -1248
rect 191 -1256 192 -1254
rect 194 -1256 195 -1254
rect 201 -1250 202 -1248
rect 198 -1256 199 -1254
rect 205 -1250 206 -1248
rect 205 -1256 206 -1254
rect 212 -1250 213 -1248
rect 212 -1256 213 -1254
rect 219 -1250 220 -1248
rect 219 -1256 220 -1254
rect 226 -1250 227 -1248
rect 226 -1256 227 -1254
rect 233 -1250 234 -1248
rect 233 -1256 234 -1254
rect 240 -1250 241 -1248
rect 240 -1256 241 -1254
rect 247 -1250 248 -1248
rect 247 -1256 248 -1254
rect 254 -1250 255 -1248
rect 254 -1256 255 -1254
rect 261 -1250 262 -1248
rect 261 -1256 262 -1254
rect 268 -1250 269 -1248
rect 271 -1250 272 -1248
rect 268 -1256 269 -1254
rect 271 -1256 272 -1254
rect 275 -1250 276 -1248
rect 275 -1256 276 -1254
rect 282 -1250 283 -1248
rect 282 -1256 283 -1254
rect 289 -1250 290 -1248
rect 289 -1256 290 -1254
rect 292 -1256 293 -1254
rect 296 -1250 297 -1248
rect 296 -1256 297 -1254
rect 303 -1250 304 -1248
rect 303 -1256 304 -1254
rect 310 -1250 311 -1248
rect 310 -1256 311 -1254
rect 317 -1250 318 -1248
rect 317 -1256 318 -1254
rect 324 -1250 325 -1248
rect 324 -1256 325 -1254
rect 331 -1250 332 -1248
rect 331 -1256 332 -1254
rect 338 -1250 339 -1248
rect 338 -1256 339 -1254
rect 345 -1250 346 -1248
rect 345 -1256 346 -1254
rect 352 -1250 353 -1248
rect 352 -1256 353 -1254
rect 359 -1250 360 -1248
rect 359 -1256 360 -1254
rect 366 -1250 367 -1248
rect 369 -1250 370 -1248
rect 366 -1256 367 -1254
rect 369 -1256 370 -1254
rect 373 -1250 374 -1248
rect 376 -1250 377 -1248
rect 380 -1250 381 -1248
rect 380 -1256 381 -1254
rect 387 -1250 388 -1248
rect 387 -1256 388 -1254
rect 394 -1250 395 -1248
rect 394 -1256 395 -1254
rect 401 -1250 402 -1248
rect 401 -1256 402 -1254
rect 408 -1250 409 -1248
rect 408 -1256 409 -1254
rect 415 -1250 416 -1248
rect 415 -1256 416 -1254
rect 422 -1250 423 -1248
rect 422 -1256 423 -1254
rect 429 -1250 430 -1248
rect 429 -1256 430 -1254
rect 436 -1250 437 -1248
rect 436 -1256 437 -1254
rect 443 -1250 444 -1248
rect 443 -1256 444 -1254
rect 450 -1250 451 -1248
rect 457 -1250 458 -1248
rect 460 -1250 461 -1248
rect 457 -1256 458 -1254
rect 460 -1256 461 -1254
rect 464 -1250 465 -1248
rect 464 -1256 465 -1254
rect 471 -1250 472 -1248
rect 471 -1256 472 -1254
rect 478 -1250 479 -1248
rect 478 -1256 479 -1254
rect 485 -1250 486 -1248
rect 485 -1256 486 -1254
rect 492 -1250 493 -1248
rect 492 -1256 493 -1254
rect 495 -1256 496 -1254
rect 499 -1250 500 -1248
rect 499 -1256 500 -1254
rect 506 -1250 507 -1248
rect 509 -1250 510 -1248
rect 506 -1256 507 -1254
rect 509 -1256 510 -1254
rect 513 -1250 514 -1248
rect 513 -1256 514 -1254
rect 520 -1250 521 -1248
rect 520 -1256 521 -1254
rect 527 -1250 528 -1248
rect 527 -1256 528 -1254
rect 537 -1250 538 -1248
rect 534 -1256 535 -1254
rect 541 -1250 542 -1248
rect 541 -1256 542 -1254
rect 548 -1250 549 -1248
rect 548 -1256 549 -1254
rect 555 -1250 556 -1248
rect 555 -1256 556 -1254
rect 562 -1250 563 -1248
rect 562 -1256 563 -1254
rect 569 -1250 570 -1248
rect 569 -1256 570 -1254
rect 576 -1250 577 -1248
rect 576 -1256 577 -1254
rect 583 -1250 584 -1248
rect 583 -1256 584 -1254
rect 590 -1250 591 -1248
rect 590 -1256 591 -1254
rect 600 -1250 601 -1248
rect 597 -1256 598 -1254
rect 600 -1256 601 -1254
rect 604 -1250 605 -1248
rect 604 -1256 605 -1254
rect 611 -1250 612 -1248
rect 611 -1256 612 -1254
rect 618 -1250 619 -1248
rect 618 -1256 619 -1254
rect 625 -1250 626 -1248
rect 625 -1256 626 -1254
rect 632 -1256 633 -1254
rect 635 -1256 636 -1254
rect 642 -1250 643 -1248
rect 639 -1256 640 -1254
rect 642 -1256 643 -1254
rect 646 -1250 647 -1248
rect 646 -1256 647 -1254
rect 656 -1250 657 -1248
rect 653 -1256 654 -1254
rect 656 -1256 657 -1254
rect 660 -1250 661 -1248
rect 660 -1256 661 -1254
rect 667 -1250 668 -1248
rect 670 -1250 671 -1248
rect 667 -1256 668 -1254
rect 670 -1256 671 -1254
rect 674 -1250 675 -1248
rect 674 -1256 675 -1254
rect 681 -1250 682 -1248
rect 684 -1250 685 -1248
rect 688 -1250 689 -1248
rect 688 -1256 689 -1254
rect 695 -1250 696 -1248
rect 695 -1256 696 -1254
rect 702 -1250 703 -1248
rect 705 -1250 706 -1248
rect 705 -1256 706 -1254
rect 709 -1250 710 -1248
rect 709 -1256 710 -1254
rect 716 -1250 717 -1248
rect 719 -1250 720 -1248
rect 723 -1250 724 -1248
rect 723 -1256 724 -1254
rect 730 -1250 731 -1248
rect 730 -1256 731 -1254
rect 737 -1250 738 -1248
rect 737 -1256 738 -1254
rect 744 -1250 745 -1248
rect 744 -1256 745 -1254
rect 751 -1250 752 -1248
rect 751 -1256 752 -1254
rect 758 -1250 759 -1248
rect 758 -1256 759 -1254
rect 765 -1250 766 -1248
rect 765 -1256 766 -1254
rect 772 -1250 773 -1248
rect 772 -1256 773 -1254
rect 779 -1250 780 -1248
rect 779 -1256 780 -1254
rect 786 -1250 787 -1248
rect 789 -1256 790 -1254
rect 793 -1250 794 -1248
rect 793 -1256 794 -1254
rect 800 -1250 801 -1248
rect 800 -1256 801 -1254
rect 807 -1250 808 -1248
rect 807 -1256 808 -1254
rect 814 -1250 815 -1248
rect 814 -1256 815 -1254
rect 821 -1250 822 -1248
rect 821 -1256 822 -1254
rect 828 -1256 829 -1254
rect 831 -1256 832 -1254
rect 835 -1250 836 -1248
rect 835 -1256 836 -1254
rect 842 -1250 843 -1248
rect 842 -1256 843 -1254
rect 849 -1250 850 -1248
rect 849 -1256 850 -1254
rect 856 -1250 857 -1248
rect 856 -1256 857 -1254
rect 863 -1250 864 -1248
rect 863 -1256 864 -1254
rect 870 -1250 871 -1248
rect 870 -1256 871 -1254
rect 877 -1250 878 -1248
rect 877 -1256 878 -1254
rect 884 -1250 885 -1248
rect 884 -1256 885 -1254
rect 891 -1250 892 -1248
rect 891 -1256 892 -1254
rect 898 -1250 899 -1248
rect 898 -1256 899 -1254
rect 905 -1250 906 -1248
rect 905 -1256 906 -1254
rect 912 -1250 913 -1248
rect 912 -1256 913 -1254
rect 919 -1250 920 -1248
rect 919 -1256 920 -1254
rect 926 -1250 927 -1248
rect 926 -1256 927 -1254
rect 933 -1250 934 -1248
rect 933 -1256 934 -1254
rect 940 -1250 941 -1248
rect 940 -1256 941 -1254
rect 947 -1250 948 -1248
rect 947 -1256 948 -1254
rect 954 -1250 955 -1248
rect 954 -1256 955 -1254
rect 961 -1250 962 -1248
rect 961 -1256 962 -1254
rect 968 -1250 969 -1248
rect 968 -1256 969 -1254
rect 975 -1250 976 -1248
rect 975 -1256 976 -1254
rect 982 -1250 983 -1248
rect 982 -1256 983 -1254
rect 989 -1250 990 -1248
rect 989 -1256 990 -1254
rect 996 -1250 997 -1248
rect 996 -1256 997 -1254
rect 1003 -1250 1004 -1248
rect 1003 -1256 1004 -1254
rect 1010 -1250 1011 -1248
rect 1010 -1256 1011 -1254
rect 1017 -1250 1018 -1248
rect 1017 -1256 1018 -1254
rect 1024 -1250 1025 -1248
rect 1024 -1256 1025 -1254
rect 1027 -1256 1028 -1254
rect 1031 -1250 1032 -1248
rect 1031 -1256 1032 -1254
rect 1038 -1250 1039 -1248
rect 1038 -1256 1039 -1254
rect 1045 -1250 1046 -1248
rect 1045 -1256 1046 -1254
rect 1052 -1250 1053 -1248
rect 1052 -1256 1053 -1254
rect 1059 -1250 1060 -1248
rect 1059 -1256 1060 -1254
rect 1066 -1250 1067 -1248
rect 1066 -1256 1067 -1254
rect 1073 -1250 1074 -1248
rect 1073 -1256 1074 -1254
rect 1080 -1250 1081 -1248
rect 1080 -1256 1081 -1254
rect 1087 -1250 1088 -1248
rect 1087 -1256 1088 -1254
rect 1094 -1250 1095 -1248
rect 1094 -1256 1095 -1254
rect 1101 -1250 1102 -1248
rect 1101 -1256 1102 -1254
rect 1108 -1250 1109 -1248
rect 1108 -1256 1109 -1254
rect 1115 -1250 1116 -1248
rect 1118 -1250 1119 -1248
rect 1115 -1256 1116 -1254
rect 1122 -1250 1123 -1248
rect 1122 -1256 1123 -1254
rect 1129 -1250 1130 -1248
rect 1132 -1256 1133 -1254
rect 1136 -1250 1137 -1248
rect 1136 -1256 1137 -1254
rect 1143 -1250 1144 -1248
rect 1143 -1256 1144 -1254
rect 1150 -1250 1151 -1248
rect 1150 -1256 1151 -1254
rect 1157 -1250 1158 -1248
rect 1157 -1256 1158 -1254
rect 1164 -1250 1165 -1248
rect 1164 -1256 1165 -1254
rect 2 -1343 3 -1341
rect 2 -1349 3 -1347
rect 9 -1343 10 -1341
rect 9 -1349 10 -1347
rect 16 -1343 17 -1341
rect 16 -1349 17 -1347
rect 23 -1343 24 -1341
rect 26 -1343 27 -1341
rect 26 -1349 27 -1347
rect 33 -1343 34 -1341
rect 30 -1349 31 -1347
rect 33 -1349 34 -1347
rect 37 -1343 38 -1341
rect 37 -1349 38 -1347
rect 44 -1343 45 -1341
rect 44 -1349 45 -1347
rect 51 -1343 52 -1341
rect 51 -1349 52 -1347
rect 58 -1343 59 -1341
rect 58 -1349 59 -1347
rect 65 -1349 66 -1347
rect 68 -1349 69 -1347
rect 72 -1343 73 -1341
rect 72 -1349 73 -1347
rect 79 -1343 80 -1341
rect 79 -1349 80 -1347
rect 86 -1343 87 -1341
rect 86 -1349 87 -1347
rect 96 -1343 97 -1341
rect 93 -1349 94 -1347
rect 96 -1349 97 -1347
rect 100 -1343 101 -1341
rect 103 -1343 104 -1341
rect 100 -1349 101 -1347
rect 103 -1349 104 -1347
rect 107 -1343 108 -1341
rect 107 -1349 108 -1347
rect 114 -1343 115 -1341
rect 114 -1349 115 -1347
rect 121 -1343 122 -1341
rect 121 -1349 122 -1347
rect 128 -1343 129 -1341
rect 128 -1349 129 -1347
rect 135 -1343 136 -1341
rect 135 -1349 136 -1347
rect 142 -1343 143 -1341
rect 142 -1349 143 -1347
rect 149 -1343 150 -1341
rect 149 -1349 150 -1347
rect 156 -1343 157 -1341
rect 156 -1349 157 -1347
rect 163 -1349 164 -1347
rect 170 -1343 171 -1341
rect 170 -1349 171 -1347
rect 180 -1343 181 -1341
rect 177 -1349 178 -1347
rect 184 -1343 185 -1341
rect 184 -1349 185 -1347
rect 191 -1343 192 -1341
rect 191 -1349 192 -1347
rect 198 -1343 199 -1341
rect 198 -1349 199 -1347
rect 205 -1343 206 -1341
rect 205 -1349 206 -1347
rect 212 -1343 213 -1341
rect 215 -1343 216 -1341
rect 212 -1349 213 -1347
rect 215 -1349 216 -1347
rect 219 -1343 220 -1341
rect 219 -1349 220 -1347
rect 226 -1343 227 -1341
rect 226 -1349 227 -1347
rect 233 -1343 234 -1341
rect 233 -1349 234 -1347
rect 240 -1343 241 -1341
rect 240 -1349 241 -1347
rect 247 -1343 248 -1341
rect 247 -1349 248 -1347
rect 254 -1343 255 -1341
rect 254 -1349 255 -1347
rect 261 -1343 262 -1341
rect 261 -1349 262 -1347
rect 268 -1343 269 -1341
rect 268 -1349 269 -1347
rect 275 -1343 276 -1341
rect 275 -1349 276 -1347
rect 282 -1343 283 -1341
rect 282 -1349 283 -1347
rect 289 -1343 290 -1341
rect 292 -1349 293 -1347
rect 296 -1343 297 -1341
rect 296 -1349 297 -1347
rect 303 -1343 304 -1341
rect 303 -1349 304 -1347
rect 310 -1343 311 -1341
rect 310 -1349 311 -1347
rect 317 -1343 318 -1341
rect 317 -1349 318 -1347
rect 324 -1343 325 -1341
rect 324 -1349 325 -1347
rect 331 -1343 332 -1341
rect 331 -1349 332 -1347
rect 338 -1343 339 -1341
rect 338 -1349 339 -1347
rect 345 -1343 346 -1341
rect 348 -1343 349 -1341
rect 345 -1349 346 -1347
rect 348 -1349 349 -1347
rect 352 -1343 353 -1341
rect 352 -1349 353 -1347
rect 359 -1343 360 -1341
rect 359 -1349 360 -1347
rect 366 -1343 367 -1341
rect 366 -1349 367 -1347
rect 373 -1343 374 -1341
rect 373 -1349 374 -1347
rect 380 -1343 381 -1341
rect 380 -1349 381 -1347
rect 387 -1343 388 -1341
rect 387 -1349 388 -1347
rect 394 -1343 395 -1341
rect 394 -1349 395 -1347
rect 401 -1343 402 -1341
rect 404 -1343 405 -1341
rect 401 -1349 402 -1347
rect 408 -1343 409 -1341
rect 411 -1343 412 -1341
rect 408 -1349 409 -1347
rect 411 -1349 412 -1347
rect 415 -1343 416 -1341
rect 415 -1349 416 -1347
rect 422 -1343 423 -1341
rect 422 -1349 423 -1347
rect 429 -1343 430 -1341
rect 429 -1349 430 -1347
rect 436 -1343 437 -1341
rect 439 -1343 440 -1341
rect 439 -1349 440 -1347
rect 443 -1343 444 -1341
rect 443 -1349 444 -1347
rect 450 -1349 451 -1347
rect 457 -1343 458 -1341
rect 460 -1343 461 -1341
rect 457 -1349 458 -1347
rect 460 -1349 461 -1347
rect 464 -1343 465 -1341
rect 464 -1349 465 -1347
rect 471 -1343 472 -1341
rect 471 -1349 472 -1347
rect 478 -1343 479 -1341
rect 478 -1349 479 -1347
rect 485 -1343 486 -1341
rect 485 -1349 486 -1347
rect 492 -1343 493 -1341
rect 495 -1349 496 -1347
rect 499 -1343 500 -1341
rect 499 -1349 500 -1347
rect 506 -1343 507 -1341
rect 506 -1349 507 -1347
rect 513 -1343 514 -1341
rect 513 -1349 514 -1347
rect 520 -1343 521 -1341
rect 523 -1343 524 -1341
rect 523 -1349 524 -1347
rect 527 -1343 528 -1341
rect 527 -1349 528 -1347
rect 534 -1343 535 -1341
rect 537 -1343 538 -1341
rect 534 -1349 535 -1347
rect 537 -1349 538 -1347
rect 541 -1343 542 -1341
rect 544 -1343 545 -1341
rect 544 -1349 545 -1347
rect 548 -1343 549 -1341
rect 548 -1349 549 -1347
rect 555 -1343 556 -1341
rect 555 -1349 556 -1347
rect 562 -1343 563 -1341
rect 562 -1349 563 -1347
rect 569 -1343 570 -1341
rect 572 -1343 573 -1341
rect 569 -1349 570 -1347
rect 576 -1343 577 -1341
rect 576 -1349 577 -1347
rect 583 -1343 584 -1341
rect 583 -1349 584 -1347
rect 590 -1343 591 -1341
rect 590 -1349 591 -1347
rect 597 -1343 598 -1341
rect 597 -1349 598 -1347
rect 604 -1343 605 -1341
rect 607 -1343 608 -1341
rect 604 -1349 605 -1347
rect 611 -1343 612 -1341
rect 611 -1349 612 -1347
rect 614 -1349 615 -1347
rect 618 -1343 619 -1341
rect 621 -1343 622 -1341
rect 618 -1349 619 -1347
rect 628 -1343 629 -1341
rect 625 -1349 626 -1347
rect 632 -1343 633 -1341
rect 632 -1349 633 -1347
rect 639 -1343 640 -1341
rect 639 -1349 640 -1347
rect 646 -1343 647 -1341
rect 646 -1349 647 -1347
rect 653 -1343 654 -1341
rect 653 -1349 654 -1347
rect 660 -1343 661 -1341
rect 660 -1349 661 -1347
rect 667 -1343 668 -1341
rect 667 -1349 668 -1347
rect 674 -1343 675 -1341
rect 674 -1349 675 -1347
rect 681 -1343 682 -1341
rect 684 -1343 685 -1341
rect 681 -1349 682 -1347
rect 688 -1343 689 -1341
rect 688 -1349 689 -1347
rect 695 -1343 696 -1341
rect 695 -1349 696 -1347
rect 702 -1343 703 -1341
rect 702 -1349 703 -1347
rect 709 -1343 710 -1341
rect 709 -1349 710 -1347
rect 716 -1343 717 -1341
rect 716 -1349 717 -1347
rect 723 -1343 724 -1341
rect 723 -1349 724 -1347
rect 733 -1343 734 -1341
rect 733 -1349 734 -1347
rect 737 -1343 738 -1341
rect 737 -1349 738 -1347
rect 744 -1343 745 -1341
rect 744 -1349 745 -1347
rect 751 -1343 752 -1341
rect 751 -1349 752 -1347
rect 758 -1343 759 -1341
rect 758 -1349 759 -1347
rect 765 -1343 766 -1341
rect 765 -1349 766 -1347
rect 772 -1343 773 -1341
rect 772 -1349 773 -1347
rect 775 -1349 776 -1347
rect 779 -1343 780 -1341
rect 779 -1349 780 -1347
rect 786 -1343 787 -1341
rect 786 -1349 787 -1347
rect 793 -1343 794 -1341
rect 796 -1343 797 -1341
rect 793 -1349 794 -1347
rect 800 -1343 801 -1341
rect 800 -1349 801 -1347
rect 807 -1343 808 -1341
rect 807 -1349 808 -1347
rect 814 -1343 815 -1341
rect 814 -1349 815 -1347
rect 821 -1343 822 -1341
rect 821 -1349 822 -1347
rect 828 -1343 829 -1341
rect 831 -1343 832 -1341
rect 828 -1349 829 -1347
rect 835 -1343 836 -1341
rect 835 -1349 836 -1347
rect 842 -1343 843 -1341
rect 842 -1349 843 -1347
rect 849 -1343 850 -1341
rect 849 -1349 850 -1347
rect 856 -1343 857 -1341
rect 856 -1349 857 -1347
rect 863 -1343 864 -1341
rect 863 -1349 864 -1347
rect 870 -1343 871 -1341
rect 870 -1349 871 -1347
rect 877 -1343 878 -1341
rect 877 -1349 878 -1347
rect 884 -1343 885 -1341
rect 884 -1349 885 -1347
rect 891 -1343 892 -1341
rect 891 -1349 892 -1347
rect 898 -1343 899 -1341
rect 898 -1349 899 -1347
rect 905 -1343 906 -1341
rect 905 -1349 906 -1347
rect 912 -1343 913 -1341
rect 912 -1349 913 -1347
rect 919 -1343 920 -1341
rect 919 -1349 920 -1347
rect 926 -1343 927 -1341
rect 926 -1349 927 -1347
rect 933 -1343 934 -1341
rect 933 -1349 934 -1347
rect 940 -1343 941 -1341
rect 940 -1349 941 -1347
rect 947 -1343 948 -1341
rect 950 -1349 951 -1347
rect 954 -1343 955 -1341
rect 954 -1349 955 -1347
rect 961 -1343 962 -1341
rect 961 -1349 962 -1347
rect 968 -1343 969 -1341
rect 968 -1349 969 -1347
rect 975 -1343 976 -1341
rect 975 -1349 976 -1347
rect 982 -1343 983 -1341
rect 982 -1349 983 -1347
rect 989 -1343 990 -1341
rect 989 -1349 990 -1347
rect 996 -1343 997 -1341
rect 1003 -1343 1004 -1341
rect 1003 -1349 1004 -1347
rect 1010 -1343 1011 -1341
rect 1010 -1349 1011 -1347
rect 1017 -1343 1018 -1341
rect 1017 -1349 1018 -1347
rect 1024 -1343 1025 -1341
rect 1027 -1343 1028 -1341
rect 1024 -1349 1025 -1347
rect 1031 -1343 1032 -1341
rect 1031 -1349 1032 -1347
rect 1038 -1343 1039 -1341
rect 1038 -1349 1039 -1347
rect 1045 -1343 1046 -1341
rect 1045 -1349 1046 -1347
rect 1052 -1343 1053 -1341
rect 1052 -1349 1053 -1347
rect 1059 -1343 1060 -1341
rect 1059 -1349 1060 -1347
rect 1066 -1343 1067 -1341
rect 1066 -1349 1067 -1347
rect 1073 -1343 1074 -1341
rect 1073 -1349 1074 -1347
rect 1080 -1343 1081 -1341
rect 1080 -1349 1081 -1347
rect 1087 -1343 1088 -1341
rect 1087 -1349 1088 -1347
rect 1094 -1343 1095 -1341
rect 1094 -1349 1095 -1347
rect 1101 -1343 1102 -1341
rect 1101 -1349 1102 -1347
rect 1108 -1343 1109 -1341
rect 1108 -1349 1109 -1347
rect 1115 -1343 1116 -1341
rect 1115 -1349 1116 -1347
rect 1122 -1343 1123 -1341
rect 1122 -1349 1123 -1347
rect 1129 -1343 1130 -1341
rect 1129 -1349 1130 -1347
rect 1136 -1343 1137 -1341
rect 1136 -1349 1137 -1347
rect 1143 -1343 1144 -1341
rect 1143 -1349 1144 -1347
rect 1150 -1349 1151 -1347
rect 1153 -1349 1154 -1347
rect 1157 -1343 1158 -1341
rect 1157 -1349 1158 -1347
rect 1164 -1343 1165 -1341
rect 1164 -1349 1165 -1347
rect 1171 -1343 1172 -1341
rect 1171 -1349 1172 -1347
rect 2 -1450 3 -1448
rect 2 -1456 3 -1454
rect 9 -1456 10 -1454
rect 16 -1450 17 -1448
rect 16 -1456 17 -1454
rect 23 -1450 24 -1448
rect 23 -1456 24 -1454
rect 30 -1450 31 -1448
rect 30 -1456 31 -1454
rect 37 -1450 38 -1448
rect 37 -1456 38 -1454
rect 44 -1450 45 -1448
rect 44 -1456 45 -1454
rect 51 -1450 52 -1448
rect 51 -1456 52 -1454
rect 58 -1450 59 -1448
rect 58 -1456 59 -1454
rect 65 -1450 66 -1448
rect 65 -1456 66 -1454
rect 72 -1450 73 -1448
rect 72 -1456 73 -1454
rect 79 -1450 80 -1448
rect 79 -1456 80 -1454
rect 86 -1450 87 -1448
rect 86 -1456 87 -1454
rect 93 -1450 94 -1448
rect 93 -1456 94 -1454
rect 100 -1450 101 -1448
rect 103 -1450 104 -1448
rect 103 -1456 104 -1454
rect 110 -1450 111 -1448
rect 107 -1456 108 -1454
rect 110 -1456 111 -1454
rect 114 -1456 115 -1454
rect 121 -1450 122 -1448
rect 124 -1456 125 -1454
rect 128 -1450 129 -1448
rect 128 -1456 129 -1454
rect 135 -1450 136 -1448
rect 135 -1456 136 -1454
rect 142 -1450 143 -1448
rect 142 -1456 143 -1454
rect 149 -1450 150 -1448
rect 149 -1456 150 -1454
rect 156 -1450 157 -1448
rect 156 -1456 157 -1454
rect 163 -1450 164 -1448
rect 163 -1456 164 -1454
rect 170 -1450 171 -1448
rect 170 -1456 171 -1454
rect 177 -1450 178 -1448
rect 177 -1456 178 -1454
rect 180 -1456 181 -1454
rect 187 -1450 188 -1448
rect 184 -1456 185 -1454
rect 187 -1456 188 -1454
rect 194 -1450 195 -1448
rect 191 -1456 192 -1454
rect 194 -1456 195 -1454
rect 198 -1450 199 -1448
rect 198 -1456 199 -1454
rect 205 -1450 206 -1448
rect 205 -1456 206 -1454
rect 212 -1456 213 -1454
rect 215 -1456 216 -1454
rect 219 -1450 220 -1448
rect 219 -1456 220 -1454
rect 226 -1450 227 -1448
rect 226 -1456 227 -1454
rect 233 -1450 234 -1448
rect 233 -1456 234 -1454
rect 240 -1450 241 -1448
rect 240 -1456 241 -1454
rect 247 -1450 248 -1448
rect 247 -1456 248 -1454
rect 254 -1450 255 -1448
rect 254 -1456 255 -1454
rect 257 -1456 258 -1454
rect 261 -1450 262 -1448
rect 261 -1456 262 -1454
rect 268 -1450 269 -1448
rect 268 -1456 269 -1454
rect 275 -1450 276 -1448
rect 275 -1456 276 -1454
rect 282 -1450 283 -1448
rect 282 -1456 283 -1454
rect 289 -1450 290 -1448
rect 289 -1456 290 -1454
rect 296 -1450 297 -1448
rect 296 -1456 297 -1454
rect 303 -1450 304 -1448
rect 303 -1456 304 -1454
rect 310 -1450 311 -1448
rect 310 -1456 311 -1454
rect 317 -1450 318 -1448
rect 317 -1456 318 -1454
rect 324 -1450 325 -1448
rect 324 -1456 325 -1454
rect 331 -1450 332 -1448
rect 334 -1450 335 -1448
rect 331 -1456 332 -1454
rect 334 -1456 335 -1454
rect 338 -1450 339 -1448
rect 338 -1456 339 -1454
rect 345 -1450 346 -1448
rect 345 -1456 346 -1454
rect 352 -1450 353 -1448
rect 352 -1456 353 -1454
rect 359 -1450 360 -1448
rect 359 -1456 360 -1454
rect 366 -1450 367 -1448
rect 366 -1456 367 -1454
rect 373 -1450 374 -1448
rect 373 -1456 374 -1454
rect 380 -1450 381 -1448
rect 380 -1456 381 -1454
rect 387 -1450 388 -1448
rect 387 -1456 388 -1454
rect 394 -1450 395 -1448
rect 394 -1456 395 -1454
rect 401 -1450 402 -1448
rect 404 -1450 405 -1448
rect 404 -1456 405 -1454
rect 408 -1450 409 -1448
rect 408 -1456 409 -1454
rect 411 -1456 412 -1454
rect 415 -1450 416 -1448
rect 415 -1456 416 -1454
rect 422 -1450 423 -1448
rect 422 -1456 423 -1454
rect 432 -1450 433 -1448
rect 432 -1456 433 -1454
rect 436 -1450 437 -1448
rect 439 -1450 440 -1448
rect 439 -1456 440 -1454
rect 446 -1450 447 -1448
rect 443 -1456 444 -1454
rect 450 -1450 451 -1448
rect 450 -1456 451 -1454
rect 457 -1450 458 -1448
rect 457 -1456 458 -1454
rect 464 -1450 465 -1448
rect 464 -1456 465 -1454
rect 471 -1450 472 -1448
rect 471 -1456 472 -1454
rect 478 -1450 479 -1448
rect 485 -1450 486 -1448
rect 488 -1450 489 -1448
rect 485 -1456 486 -1454
rect 492 -1450 493 -1448
rect 495 -1450 496 -1448
rect 495 -1456 496 -1454
rect 499 -1450 500 -1448
rect 502 -1450 503 -1448
rect 499 -1456 500 -1454
rect 502 -1456 503 -1454
rect 506 -1450 507 -1448
rect 509 -1450 510 -1448
rect 506 -1456 507 -1454
rect 509 -1456 510 -1454
rect 513 -1450 514 -1448
rect 513 -1456 514 -1454
rect 520 -1450 521 -1448
rect 520 -1456 521 -1454
rect 527 -1450 528 -1448
rect 527 -1456 528 -1454
rect 534 -1450 535 -1448
rect 534 -1456 535 -1454
rect 541 -1450 542 -1448
rect 541 -1456 542 -1454
rect 548 -1450 549 -1448
rect 548 -1456 549 -1454
rect 551 -1456 552 -1454
rect 555 -1450 556 -1448
rect 555 -1456 556 -1454
rect 562 -1450 563 -1448
rect 562 -1456 563 -1454
rect 569 -1450 570 -1448
rect 569 -1456 570 -1454
rect 576 -1450 577 -1448
rect 579 -1450 580 -1448
rect 576 -1456 577 -1454
rect 579 -1456 580 -1454
rect 583 -1450 584 -1448
rect 583 -1456 584 -1454
rect 590 -1450 591 -1448
rect 590 -1456 591 -1454
rect 600 -1450 601 -1448
rect 600 -1456 601 -1454
rect 604 -1450 605 -1448
rect 604 -1456 605 -1454
rect 611 -1450 612 -1448
rect 611 -1456 612 -1454
rect 614 -1456 615 -1454
rect 618 -1450 619 -1448
rect 618 -1456 619 -1454
rect 625 -1450 626 -1448
rect 625 -1456 626 -1454
rect 632 -1450 633 -1448
rect 632 -1456 633 -1454
rect 639 -1450 640 -1448
rect 639 -1456 640 -1454
rect 646 -1450 647 -1448
rect 646 -1456 647 -1454
rect 653 -1450 654 -1448
rect 653 -1456 654 -1454
rect 660 -1450 661 -1448
rect 660 -1456 661 -1454
rect 667 -1450 668 -1448
rect 667 -1456 668 -1454
rect 674 -1450 675 -1448
rect 674 -1456 675 -1454
rect 681 -1450 682 -1448
rect 681 -1456 682 -1454
rect 688 -1450 689 -1448
rect 691 -1450 692 -1448
rect 691 -1456 692 -1454
rect 695 -1450 696 -1448
rect 695 -1456 696 -1454
rect 702 -1450 703 -1448
rect 705 -1456 706 -1454
rect 709 -1450 710 -1448
rect 709 -1456 710 -1454
rect 716 -1450 717 -1448
rect 716 -1456 717 -1454
rect 723 -1450 724 -1448
rect 723 -1456 724 -1454
rect 730 -1450 731 -1448
rect 730 -1456 731 -1454
rect 737 -1450 738 -1448
rect 737 -1456 738 -1454
rect 744 -1450 745 -1448
rect 744 -1456 745 -1454
rect 747 -1456 748 -1454
rect 751 -1450 752 -1448
rect 751 -1456 752 -1454
rect 758 -1450 759 -1448
rect 758 -1456 759 -1454
rect 765 -1450 766 -1448
rect 765 -1456 766 -1454
rect 772 -1450 773 -1448
rect 772 -1456 773 -1454
rect 779 -1450 780 -1448
rect 779 -1456 780 -1454
rect 786 -1450 787 -1448
rect 786 -1456 787 -1454
rect 793 -1450 794 -1448
rect 793 -1456 794 -1454
rect 800 -1450 801 -1448
rect 800 -1456 801 -1454
rect 807 -1450 808 -1448
rect 807 -1456 808 -1454
rect 814 -1450 815 -1448
rect 814 -1456 815 -1454
rect 821 -1450 822 -1448
rect 821 -1456 822 -1454
rect 828 -1450 829 -1448
rect 828 -1456 829 -1454
rect 835 -1450 836 -1448
rect 835 -1456 836 -1454
rect 842 -1450 843 -1448
rect 842 -1456 843 -1454
rect 849 -1450 850 -1448
rect 849 -1456 850 -1454
rect 856 -1450 857 -1448
rect 856 -1456 857 -1454
rect 859 -1456 860 -1454
rect 863 -1450 864 -1448
rect 863 -1456 864 -1454
rect 870 -1450 871 -1448
rect 870 -1456 871 -1454
rect 877 -1450 878 -1448
rect 877 -1456 878 -1454
rect 884 -1450 885 -1448
rect 884 -1456 885 -1454
rect 891 -1450 892 -1448
rect 891 -1456 892 -1454
rect 898 -1450 899 -1448
rect 898 -1456 899 -1454
rect 905 -1450 906 -1448
rect 905 -1456 906 -1454
rect 912 -1450 913 -1448
rect 912 -1456 913 -1454
rect 919 -1450 920 -1448
rect 919 -1456 920 -1454
rect 926 -1450 927 -1448
rect 926 -1456 927 -1454
rect 933 -1450 934 -1448
rect 933 -1456 934 -1454
rect 940 -1450 941 -1448
rect 940 -1456 941 -1454
rect 947 -1450 948 -1448
rect 947 -1456 948 -1454
rect 954 -1450 955 -1448
rect 954 -1456 955 -1454
rect 961 -1450 962 -1448
rect 961 -1456 962 -1454
rect 968 -1450 969 -1448
rect 968 -1456 969 -1454
rect 975 -1450 976 -1448
rect 975 -1456 976 -1454
rect 982 -1450 983 -1448
rect 982 -1456 983 -1454
rect 989 -1450 990 -1448
rect 989 -1456 990 -1454
rect 996 -1450 997 -1448
rect 996 -1456 997 -1454
rect 1003 -1450 1004 -1448
rect 1003 -1456 1004 -1454
rect 1010 -1450 1011 -1448
rect 1010 -1456 1011 -1454
rect 1017 -1450 1018 -1448
rect 1017 -1456 1018 -1454
rect 1024 -1450 1025 -1448
rect 1024 -1456 1025 -1454
rect 1031 -1450 1032 -1448
rect 1031 -1456 1032 -1454
rect 1038 -1450 1039 -1448
rect 1038 -1456 1039 -1454
rect 1045 -1450 1046 -1448
rect 1045 -1456 1046 -1454
rect 1052 -1450 1053 -1448
rect 1052 -1456 1053 -1454
rect 1062 -1450 1063 -1448
rect 1062 -1456 1063 -1454
rect 1066 -1450 1067 -1448
rect 1066 -1456 1067 -1454
rect 1073 -1450 1074 -1448
rect 1073 -1456 1074 -1454
rect 1080 -1450 1081 -1448
rect 1080 -1456 1081 -1454
rect 1087 -1450 1088 -1448
rect 1094 -1450 1095 -1448
rect 1094 -1456 1095 -1454
rect 1108 -1450 1109 -1448
rect 1108 -1456 1109 -1454
rect 2 -1541 3 -1539
rect 2 -1547 3 -1545
rect 9 -1541 10 -1539
rect 9 -1547 10 -1545
rect 16 -1541 17 -1539
rect 16 -1547 17 -1545
rect 23 -1541 24 -1539
rect 23 -1547 24 -1545
rect 30 -1541 31 -1539
rect 33 -1541 34 -1539
rect 33 -1547 34 -1545
rect 37 -1541 38 -1539
rect 37 -1547 38 -1545
rect 40 -1547 41 -1545
rect 44 -1541 45 -1539
rect 44 -1547 45 -1545
rect 51 -1541 52 -1539
rect 51 -1547 52 -1545
rect 58 -1541 59 -1539
rect 58 -1547 59 -1545
rect 65 -1541 66 -1539
rect 65 -1547 66 -1545
rect 72 -1541 73 -1539
rect 72 -1547 73 -1545
rect 79 -1541 80 -1539
rect 79 -1547 80 -1545
rect 86 -1541 87 -1539
rect 86 -1547 87 -1545
rect 93 -1541 94 -1539
rect 96 -1541 97 -1539
rect 100 -1541 101 -1539
rect 100 -1547 101 -1545
rect 107 -1541 108 -1539
rect 107 -1547 108 -1545
rect 114 -1541 115 -1539
rect 114 -1547 115 -1545
rect 121 -1541 122 -1539
rect 121 -1547 122 -1545
rect 128 -1541 129 -1539
rect 128 -1547 129 -1545
rect 135 -1541 136 -1539
rect 135 -1547 136 -1545
rect 145 -1541 146 -1539
rect 145 -1547 146 -1545
rect 149 -1541 150 -1539
rect 149 -1547 150 -1545
rect 156 -1541 157 -1539
rect 156 -1547 157 -1545
rect 163 -1541 164 -1539
rect 166 -1541 167 -1539
rect 163 -1547 164 -1545
rect 166 -1547 167 -1545
rect 170 -1541 171 -1539
rect 170 -1547 171 -1545
rect 177 -1541 178 -1539
rect 180 -1547 181 -1545
rect 184 -1541 185 -1539
rect 184 -1547 185 -1545
rect 191 -1541 192 -1539
rect 191 -1547 192 -1545
rect 198 -1541 199 -1539
rect 198 -1547 199 -1545
rect 205 -1541 206 -1539
rect 208 -1547 209 -1545
rect 212 -1541 213 -1539
rect 215 -1541 216 -1539
rect 212 -1547 213 -1545
rect 219 -1541 220 -1539
rect 219 -1547 220 -1545
rect 226 -1541 227 -1539
rect 226 -1547 227 -1545
rect 233 -1541 234 -1539
rect 233 -1547 234 -1545
rect 240 -1541 241 -1539
rect 240 -1547 241 -1545
rect 247 -1541 248 -1539
rect 250 -1547 251 -1545
rect 254 -1541 255 -1539
rect 254 -1547 255 -1545
rect 261 -1541 262 -1539
rect 261 -1547 262 -1545
rect 268 -1541 269 -1539
rect 268 -1547 269 -1545
rect 278 -1547 279 -1545
rect 282 -1541 283 -1539
rect 282 -1547 283 -1545
rect 289 -1541 290 -1539
rect 292 -1541 293 -1539
rect 292 -1547 293 -1545
rect 296 -1541 297 -1539
rect 296 -1547 297 -1545
rect 303 -1541 304 -1539
rect 303 -1547 304 -1545
rect 310 -1541 311 -1539
rect 310 -1547 311 -1545
rect 317 -1541 318 -1539
rect 317 -1547 318 -1545
rect 324 -1541 325 -1539
rect 327 -1541 328 -1539
rect 324 -1547 325 -1545
rect 331 -1541 332 -1539
rect 331 -1547 332 -1545
rect 338 -1541 339 -1539
rect 338 -1547 339 -1545
rect 345 -1541 346 -1539
rect 345 -1547 346 -1545
rect 352 -1541 353 -1539
rect 352 -1547 353 -1545
rect 359 -1541 360 -1539
rect 359 -1547 360 -1545
rect 366 -1541 367 -1539
rect 366 -1547 367 -1545
rect 373 -1541 374 -1539
rect 373 -1547 374 -1545
rect 380 -1541 381 -1539
rect 380 -1547 381 -1545
rect 387 -1541 388 -1539
rect 387 -1547 388 -1545
rect 394 -1541 395 -1539
rect 394 -1547 395 -1545
rect 401 -1541 402 -1539
rect 401 -1547 402 -1545
rect 408 -1541 409 -1539
rect 408 -1547 409 -1545
rect 415 -1541 416 -1539
rect 415 -1547 416 -1545
rect 422 -1541 423 -1539
rect 422 -1547 423 -1545
rect 429 -1541 430 -1539
rect 429 -1547 430 -1545
rect 436 -1541 437 -1539
rect 436 -1547 437 -1545
rect 443 -1541 444 -1539
rect 443 -1547 444 -1545
rect 450 -1541 451 -1539
rect 450 -1547 451 -1545
rect 457 -1541 458 -1539
rect 457 -1547 458 -1545
rect 460 -1547 461 -1545
rect 467 -1541 468 -1539
rect 464 -1547 465 -1545
rect 467 -1547 468 -1545
rect 471 -1547 472 -1545
rect 478 -1541 479 -1539
rect 481 -1541 482 -1539
rect 478 -1547 479 -1545
rect 485 -1541 486 -1539
rect 485 -1547 486 -1545
rect 492 -1541 493 -1539
rect 492 -1547 493 -1545
rect 499 -1541 500 -1539
rect 499 -1547 500 -1545
rect 506 -1541 507 -1539
rect 506 -1547 507 -1545
rect 513 -1541 514 -1539
rect 516 -1541 517 -1539
rect 516 -1547 517 -1545
rect 523 -1541 524 -1539
rect 520 -1547 521 -1545
rect 523 -1547 524 -1545
rect 527 -1541 528 -1539
rect 527 -1547 528 -1545
rect 534 -1541 535 -1539
rect 537 -1541 538 -1539
rect 534 -1547 535 -1545
rect 537 -1547 538 -1545
rect 541 -1541 542 -1539
rect 541 -1547 542 -1545
rect 548 -1541 549 -1539
rect 548 -1547 549 -1545
rect 555 -1541 556 -1539
rect 555 -1547 556 -1545
rect 562 -1541 563 -1539
rect 562 -1547 563 -1545
rect 565 -1547 566 -1545
rect 569 -1541 570 -1539
rect 569 -1547 570 -1545
rect 576 -1541 577 -1539
rect 576 -1547 577 -1545
rect 583 -1541 584 -1539
rect 583 -1547 584 -1545
rect 590 -1541 591 -1539
rect 590 -1547 591 -1545
rect 593 -1547 594 -1545
rect 597 -1541 598 -1539
rect 597 -1547 598 -1545
rect 604 -1541 605 -1539
rect 604 -1547 605 -1545
rect 611 -1541 612 -1539
rect 611 -1547 612 -1545
rect 618 -1541 619 -1539
rect 618 -1547 619 -1545
rect 625 -1541 626 -1539
rect 625 -1547 626 -1545
rect 632 -1541 633 -1539
rect 632 -1547 633 -1545
rect 639 -1541 640 -1539
rect 639 -1547 640 -1545
rect 646 -1541 647 -1539
rect 646 -1547 647 -1545
rect 653 -1541 654 -1539
rect 653 -1547 654 -1545
rect 663 -1541 664 -1539
rect 663 -1547 664 -1545
rect 670 -1541 671 -1539
rect 667 -1547 668 -1545
rect 670 -1547 671 -1545
rect 674 -1541 675 -1539
rect 677 -1541 678 -1539
rect 674 -1547 675 -1545
rect 677 -1547 678 -1545
rect 681 -1541 682 -1539
rect 681 -1547 682 -1545
rect 688 -1541 689 -1539
rect 691 -1541 692 -1539
rect 695 -1541 696 -1539
rect 695 -1547 696 -1545
rect 702 -1541 703 -1539
rect 702 -1547 703 -1545
rect 709 -1541 710 -1539
rect 709 -1547 710 -1545
rect 716 -1541 717 -1539
rect 716 -1547 717 -1545
rect 723 -1541 724 -1539
rect 723 -1547 724 -1545
rect 730 -1541 731 -1539
rect 730 -1547 731 -1545
rect 737 -1541 738 -1539
rect 737 -1547 738 -1545
rect 744 -1541 745 -1539
rect 744 -1547 745 -1545
rect 751 -1541 752 -1539
rect 751 -1547 752 -1545
rect 758 -1541 759 -1539
rect 758 -1547 759 -1545
rect 765 -1541 766 -1539
rect 765 -1547 766 -1545
rect 772 -1547 773 -1545
rect 775 -1547 776 -1545
rect 779 -1541 780 -1539
rect 779 -1547 780 -1545
rect 786 -1541 787 -1539
rect 786 -1547 787 -1545
rect 793 -1541 794 -1539
rect 793 -1547 794 -1545
rect 800 -1541 801 -1539
rect 800 -1547 801 -1545
rect 807 -1541 808 -1539
rect 807 -1547 808 -1545
rect 814 -1541 815 -1539
rect 814 -1547 815 -1545
rect 821 -1541 822 -1539
rect 821 -1547 822 -1545
rect 828 -1541 829 -1539
rect 828 -1547 829 -1545
rect 835 -1541 836 -1539
rect 835 -1547 836 -1545
rect 842 -1541 843 -1539
rect 842 -1547 843 -1545
rect 849 -1541 850 -1539
rect 849 -1547 850 -1545
rect 856 -1541 857 -1539
rect 856 -1547 857 -1545
rect 863 -1541 864 -1539
rect 863 -1547 864 -1545
rect 870 -1541 871 -1539
rect 870 -1547 871 -1545
rect 877 -1541 878 -1539
rect 877 -1547 878 -1545
rect 884 -1541 885 -1539
rect 884 -1547 885 -1545
rect 891 -1541 892 -1539
rect 891 -1547 892 -1545
rect 898 -1541 899 -1539
rect 898 -1547 899 -1545
rect 905 -1541 906 -1539
rect 905 -1547 906 -1545
rect 912 -1541 913 -1539
rect 912 -1547 913 -1545
rect 919 -1541 920 -1539
rect 919 -1547 920 -1545
rect 926 -1541 927 -1539
rect 926 -1547 927 -1545
rect 933 -1541 934 -1539
rect 933 -1547 934 -1545
rect 940 -1541 941 -1539
rect 940 -1547 941 -1545
rect 947 -1541 948 -1539
rect 947 -1547 948 -1545
rect 954 -1541 955 -1539
rect 954 -1547 955 -1545
rect 961 -1541 962 -1539
rect 961 -1547 962 -1545
rect 968 -1541 969 -1539
rect 968 -1547 969 -1545
rect 975 -1541 976 -1539
rect 975 -1547 976 -1545
rect 982 -1541 983 -1539
rect 982 -1547 983 -1545
rect 989 -1541 990 -1539
rect 989 -1547 990 -1545
rect 996 -1541 997 -1539
rect 996 -1547 997 -1545
rect 1003 -1541 1004 -1539
rect 1003 -1547 1004 -1545
rect 1010 -1541 1011 -1539
rect 1017 -1541 1018 -1539
rect 1017 -1547 1018 -1545
rect 1024 -1541 1025 -1539
rect 1024 -1547 1025 -1545
rect 1031 -1541 1032 -1539
rect 1031 -1547 1032 -1545
rect 1034 -1547 1035 -1545
rect 1038 -1541 1039 -1539
rect 1038 -1547 1039 -1545
rect 1045 -1541 1046 -1539
rect 1045 -1547 1046 -1545
rect 1059 -1541 1060 -1539
rect 1059 -1547 1060 -1545
rect 1073 -1541 1074 -1539
rect 1073 -1547 1074 -1545
rect 1094 -1541 1095 -1539
rect 1094 -1547 1095 -1545
rect 5 -1630 6 -1628
rect 9 -1630 10 -1628
rect 9 -1636 10 -1634
rect 16 -1630 17 -1628
rect 16 -1636 17 -1634
rect 23 -1630 24 -1628
rect 23 -1636 24 -1634
rect 30 -1630 31 -1628
rect 30 -1636 31 -1634
rect 37 -1630 38 -1628
rect 37 -1636 38 -1634
rect 44 -1630 45 -1628
rect 44 -1636 45 -1634
rect 51 -1630 52 -1628
rect 51 -1636 52 -1634
rect 58 -1630 59 -1628
rect 58 -1636 59 -1634
rect 61 -1636 62 -1634
rect 65 -1630 66 -1628
rect 65 -1636 66 -1634
rect 72 -1630 73 -1628
rect 72 -1636 73 -1634
rect 79 -1630 80 -1628
rect 82 -1630 83 -1628
rect 82 -1636 83 -1634
rect 86 -1630 87 -1628
rect 86 -1636 87 -1634
rect 93 -1630 94 -1628
rect 96 -1630 97 -1628
rect 96 -1636 97 -1634
rect 100 -1630 101 -1628
rect 100 -1636 101 -1634
rect 107 -1630 108 -1628
rect 107 -1636 108 -1634
rect 114 -1630 115 -1628
rect 114 -1636 115 -1634
rect 121 -1630 122 -1628
rect 121 -1636 122 -1634
rect 128 -1630 129 -1628
rect 128 -1636 129 -1634
rect 135 -1636 136 -1634
rect 138 -1636 139 -1634
rect 145 -1630 146 -1628
rect 142 -1636 143 -1634
rect 149 -1630 150 -1628
rect 149 -1636 150 -1634
rect 156 -1630 157 -1628
rect 156 -1636 157 -1634
rect 163 -1630 164 -1628
rect 163 -1636 164 -1634
rect 170 -1630 171 -1628
rect 170 -1636 171 -1634
rect 177 -1630 178 -1628
rect 177 -1636 178 -1634
rect 184 -1636 185 -1634
rect 187 -1636 188 -1634
rect 191 -1630 192 -1628
rect 191 -1636 192 -1634
rect 201 -1630 202 -1628
rect 198 -1636 199 -1634
rect 201 -1636 202 -1634
rect 205 -1630 206 -1628
rect 205 -1636 206 -1634
rect 212 -1630 213 -1628
rect 212 -1636 213 -1634
rect 222 -1630 223 -1628
rect 222 -1636 223 -1634
rect 226 -1630 227 -1628
rect 229 -1630 230 -1628
rect 226 -1636 227 -1634
rect 233 -1630 234 -1628
rect 233 -1636 234 -1634
rect 240 -1630 241 -1628
rect 240 -1636 241 -1634
rect 247 -1630 248 -1628
rect 254 -1630 255 -1628
rect 254 -1636 255 -1634
rect 261 -1630 262 -1628
rect 261 -1636 262 -1634
rect 268 -1630 269 -1628
rect 268 -1636 269 -1634
rect 275 -1630 276 -1628
rect 275 -1636 276 -1634
rect 282 -1630 283 -1628
rect 282 -1636 283 -1634
rect 289 -1630 290 -1628
rect 289 -1636 290 -1634
rect 296 -1630 297 -1628
rect 296 -1636 297 -1634
rect 303 -1636 304 -1634
rect 306 -1636 307 -1634
rect 310 -1630 311 -1628
rect 310 -1636 311 -1634
rect 317 -1630 318 -1628
rect 317 -1636 318 -1634
rect 327 -1630 328 -1628
rect 324 -1636 325 -1634
rect 327 -1636 328 -1634
rect 331 -1630 332 -1628
rect 331 -1636 332 -1634
rect 338 -1630 339 -1628
rect 338 -1636 339 -1634
rect 345 -1630 346 -1628
rect 345 -1636 346 -1634
rect 352 -1630 353 -1628
rect 355 -1630 356 -1628
rect 355 -1636 356 -1634
rect 359 -1630 360 -1628
rect 359 -1636 360 -1634
rect 366 -1630 367 -1628
rect 366 -1636 367 -1634
rect 373 -1630 374 -1628
rect 376 -1630 377 -1628
rect 373 -1636 374 -1634
rect 376 -1636 377 -1634
rect 380 -1630 381 -1628
rect 380 -1636 381 -1634
rect 387 -1630 388 -1628
rect 387 -1636 388 -1634
rect 394 -1630 395 -1628
rect 394 -1636 395 -1634
rect 401 -1630 402 -1628
rect 401 -1636 402 -1634
rect 408 -1630 409 -1628
rect 408 -1636 409 -1634
rect 415 -1630 416 -1628
rect 415 -1636 416 -1634
rect 425 -1630 426 -1628
rect 422 -1636 423 -1634
rect 425 -1636 426 -1634
rect 429 -1630 430 -1628
rect 429 -1636 430 -1634
rect 436 -1630 437 -1628
rect 436 -1636 437 -1634
rect 443 -1630 444 -1628
rect 446 -1636 447 -1634
rect 450 -1630 451 -1628
rect 450 -1636 451 -1634
rect 457 -1630 458 -1628
rect 457 -1636 458 -1634
rect 460 -1636 461 -1634
rect 464 -1630 465 -1628
rect 464 -1636 465 -1634
rect 471 -1630 472 -1628
rect 471 -1636 472 -1634
rect 478 -1630 479 -1628
rect 478 -1636 479 -1634
rect 485 -1630 486 -1628
rect 485 -1636 486 -1634
rect 492 -1630 493 -1628
rect 492 -1636 493 -1634
rect 499 -1630 500 -1628
rect 499 -1636 500 -1634
rect 506 -1630 507 -1628
rect 506 -1636 507 -1634
rect 513 -1630 514 -1628
rect 513 -1636 514 -1634
rect 520 -1630 521 -1628
rect 520 -1636 521 -1634
rect 527 -1630 528 -1628
rect 527 -1636 528 -1634
rect 534 -1630 535 -1628
rect 537 -1636 538 -1634
rect 541 -1630 542 -1628
rect 541 -1636 542 -1634
rect 548 -1630 549 -1628
rect 548 -1636 549 -1634
rect 555 -1630 556 -1628
rect 555 -1636 556 -1634
rect 562 -1630 563 -1628
rect 562 -1636 563 -1634
rect 569 -1630 570 -1628
rect 569 -1636 570 -1634
rect 572 -1636 573 -1634
rect 576 -1630 577 -1628
rect 576 -1636 577 -1634
rect 586 -1630 587 -1628
rect 583 -1636 584 -1634
rect 590 -1630 591 -1628
rect 590 -1636 591 -1634
rect 597 -1630 598 -1628
rect 597 -1636 598 -1634
rect 604 -1630 605 -1628
rect 604 -1636 605 -1634
rect 611 -1630 612 -1628
rect 614 -1630 615 -1628
rect 614 -1636 615 -1634
rect 618 -1630 619 -1628
rect 618 -1636 619 -1634
rect 625 -1630 626 -1628
rect 625 -1636 626 -1634
rect 632 -1630 633 -1628
rect 635 -1630 636 -1628
rect 632 -1636 633 -1634
rect 639 -1630 640 -1628
rect 639 -1636 640 -1634
rect 646 -1630 647 -1628
rect 646 -1636 647 -1634
rect 653 -1630 654 -1628
rect 653 -1636 654 -1634
rect 660 -1630 661 -1628
rect 660 -1636 661 -1634
rect 667 -1630 668 -1628
rect 667 -1636 668 -1634
rect 674 -1630 675 -1628
rect 677 -1630 678 -1628
rect 674 -1636 675 -1634
rect 677 -1636 678 -1634
rect 684 -1630 685 -1628
rect 681 -1636 682 -1634
rect 684 -1636 685 -1634
rect 688 -1630 689 -1628
rect 688 -1636 689 -1634
rect 695 -1630 696 -1628
rect 695 -1636 696 -1634
rect 702 -1630 703 -1628
rect 702 -1636 703 -1634
rect 709 -1630 710 -1628
rect 709 -1636 710 -1634
rect 716 -1630 717 -1628
rect 716 -1636 717 -1634
rect 723 -1630 724 -1628
rect 723 -1636 724 -1634
rect 730 -1630 731 -1628
rect 730 -1636 731 -1634
rect 737 -1630 738 -1628
rect 737 -1636 738 -1634
rect 744 -1630 745 -1628
rect 744 -1636 745 -1634
rect 751 -1630 752 -1628
rect 751 -1636 752 -1634
rect 758 -1630 759 -1628
rect 758 -1636 759 -1634
rect 765 -1630 766 -1628
rect 765 -1636 766 -1634
rect 772 -1630 773 -1628
rect 772 -1636 773 -1634
rect 779 -1630 780 -1628
rect 779 -1636 780 -1634
rect 786 -1630 787 -1628
rect 786 -1636 787 -1634
rect 793 -1630 794 -1628
rect 793 -1636 794 -1634
rect 800 -1630 801 -1628
rect 800 -1636 801 -1634
rect 807 -1630 808 -1628
rect 807 -1636 808 -1634
rect 814 -1630 815 -1628
rect 814 -1636 815 -1634
rect 821 -1630 822 -1628
rect 821 -1636 822 -1634
rect 828 -1630 829 -1628
rect 828 -1636 829 -1634
rect 835 -1630 836 -1628
rect 835 -1636 836 -1634
rect 842 -1630 843 -1628
rect 842 -1636 843 -1634
rect 849 -1630 850 -1628
rect 849 -1636 850 -1634
rect 856 -1630 857 -1628
rect 859 -1630 860 -1628
rect 856 -1636 857 -1634
rect 863 -1630 864 -1628
rect 863 -1636 864 -1634
rect 870 -1630 871 -1628
rect 870 -1636 871 -1634
rect 877 -1630 878 -1628
rect 877 -1636 878 -1634
rect 884 -1630 885 -1628
rect 884 -1636 885 -1634
rect 891 -1630 892 -1628
rect 891 -1636 892 -1634
rect 898 -1630 899 -1628
rect 898 -1636 899 -1634
rect 905 -1630 906 -1628
rect 905 -1636 906 -1634
rect 912 -1630 913 -1628
rect 912 -1636 913 -1634
rect 919 -1630 920 -1628
rect 919 -1636 920 -1634
rect 926 -1630 927 -1628
rect 926 -1636 927 -1634
rect 933 -1630 934 -1628
rect 933 -1636 934 -1634
rect 940 -1630 941 -1628
rect 940 -1636 941 -1634
rect 947 -1630 948 -1628
rect 947 -1636 948 -1634
rect 954 -1630 955 -1628
rect 954 -1636 955 -1634
rect 961 -1630 962 -1628
rect 961 -1636 962 -1634
rect 968 -1630 969 -1628
rect 968 -1636 969 -1634
rect 975 -1630 976 -1628
rect 975 -1636 976 -1634
rect 982 -1630 983 -1628
rect 982 -1636 983 -1634
rect 989 -1630 990 -1628
rect 989 -1636 990 -1634
rect 996 -1630 997 -1628
rect 996 -1636 997 -1634
rect 1003 -1630 1004 -1628
rect 1003 -1636 1004 -1634
rect 1010 -1630 1011 -1628
rect 1010 -1636 1011 -1634
rect 1017 -1630 1018 -1628
rect 1017 -1636 1018 -1634
rect 1024 -1630 1025 -1628
rect 1024 -1636 1025 -1634
rect 1031 -1630 1032 -1628
rect 1031 -1636 1032 -1634
rect 1038 -1630 1039 -1628
rect 1038 -1636 1039 -1634
rect 1045 -1630 1046 -1628
rect 1045 -1636 1046 -1634
rect 1052 -1630 1053 -1628
rect 1052 -1636 1053 -1634
rect 1062 -1630 1063 -1628
rect 1059 -1636 1060 -1634
rect 1062 -1636 1063 -1634
rect 1069 -1630 1070 -1628
rect 1069 -1636 1070 -1634
rect 1073 -1630 1074 -1628
rect 1073 -1636 1074 -1634
rect 1080 -1630 1081 -1628
rect 1080 -1636 1081 -1634
rect 1087 -1630 1088 -1628
rect 1087 -1636 1088 -1634
rect 1094 -1630 1095 -1628
rect 1094 -1636 1095 -1634
rect 1101 -1630 1102 -1628
rect 1101 -1636 1102 -1634
rect 1108 -1630 1109 -1628
rect 1108 -1636 1109 -1634
rect 1115 -1630 1116 -1628
rect 1115 -1636 1116 -1634
rect 23 -1715 24 -1713
rect 23 -1721 24 -1719
rect 30 -1715 31 -1713
rect 30 -1721 31 -1719
rect 37 -1715 38 -1713
rect 37 -1721 38 -1719
rect 44 -1715 45 -1713
rect 44 -1721 45 -1719
rect 51 -1715 52 -1713
rect 54 -1715 55 -1713
rect 58 -1715 59 -1713
rect 58 -1721 59 -1719
rect 65 -1715 66 -1713
rect 68 -1715 69 -1713
rect 65 -1721 66 -1719
rect 72 -1715 73 -1713
rect 72 -1721 73 -1719
rect 79 -1715 80 -1713
rect 79 -1721 80 -1719
rect 86 -1715 87 -1713
rect 86 -1721 87 -1719
rect 93 -1715 94 -1713
rect 93 -1721 94 -1719
rect 100 -1715 101 -1713
rect 100 -1721 101 -1719
rect 107 -1715 108 -1713
rect 107 -1721 108 -1719
rect 114 -1715 115 -1713
rect 114 -1721 115 -1719
rect 121 -1715 122 -1713
rect 121 -1721 122 -1719
rect 128 -1715 129 -1713
rect 128 -1721 129 -1719
rect 135 -1715 136 -1713
rect 135 -1721 136 -1719
rect 142 -1715 143 -1713
rect 142 -1721 143 -1719
rect 149 -1715 150 -1713
rect 149 -1721 150 -1719
rect 159 -1715 160 -1713
rect 156 -1721 157 -1719
rect 159 -1721 160 -1719
rect 163 -1715 164 -1713
rect 163 -1721 164 -1719
rect 170 -1715 171 -1713
rect 170 -1721 171 -1719
rect 177 -1715 178 -1713
rect 177 -1721 178 -1719
rect 184 -1715 185 -1713
rect 184 -1721 185 -1719
rect 191 -1715 192 -1713
rect 191 -1721 192 -1719
rect 198 -1715 199 -1713
rect 198 -1721 199 -1719
rect 205 -1715 206 -1713
rect 205 -1721 206 -1719
rect 212 -1715 213 -1713
rect 212 -1721 213 -1719
rect 222 -1721 223 -1719
rect 226 -1715 227 -1713
rect 226 -1721 227 -1719
rect 233 -1715 234 -1713
rect 233 -1721 234 -1719
rect 240 -1715 241 -1713
rect 240 -1721 241 -1719
rect 247 -1715 248 -1713
rect 247 -1721 248 -1719
rect 254 -1715 255 -1713
rect 254 -1721 255 -1719
rect 261 -1715 262 -1713
rect 261 -1721 262 -1719
rect 268 -1715 269 -1713
rect 268 -1721 269 -1719
rect 275 -1715 276 -1713
rect 275 -1721 276 -1719
rect 282 -1715 283 -1713
rect 282 -1721 283 -1719
rect 289 -1715 290 -1713
rect 289 -1721 290 -1719
rect 296 -1715 297 -1713
rect 296 -1721 297 -1719
rect 303 -1715 304 -1713
rect 303 -1721 304 -1719
rect 310 -1715 311 -1713
rect 313 -1715 314 -1713
rect 310 -1721 311 -1719
rect 317 -1715 318 -1713
rect 317 -1721 318 -1719
rect 327 -1715 328 -1713
rect 324 -1721 325 -1719
rect 331 -1715 332 -1713
rect 331 -1721 332 -1719
rect 341 -1715 342 -1713
rect 341 -1721 342 -1719
rect 345 -1715 346 -1713
rect 345 -1721 346 -1719
rect 355 -1715 356 -1713
rect 352 -1721 353 -1719
rect 355 -1721 356 -1719
rect 359 -1715 360 -1713
rect 362 -1715 363 -1713
rect 362 -1721 363 -1719
rect 366 -1715 367 -1713
rect 366 -1721 367 -1719
rect 373 -1715 374 -1713
rect 376 -1715 377 -1713
rect 373 -1721 374 -1719
rect 376 -1721 377 -1719
rect 380 -1715 381 -1713
rect 383 -1715 384 -1713
rect 380 -1721 381 -1719
rect 383 -1721 384 -1719
rect 387 -1715 388 -1713
rect 387 -1721 388 -1719
rect 394 -1715 395 -1713
rect 394 -1721 395 -1719
rect 401 -1715 402 -1713
rect 401 -1721 402 -1719
rect 408 -1715 409 -1713
rect 408 -1721 409 -1719
rect 415 -1715 416 -1713
rect 415 -1721 416 -1719
rect 422 -1715 423 -1713
rect 425 -1721 426 -1719
rect 429 -1715 430 -1713
rect 429 -1721 430 -1719
rect 436 -1715 437 -1713
rect 436 -1721 437 -1719
rect 443 -1715 444 -1713
rect 443 -1721 444 -1719
rect 450 -1715 451 -1713
rect 450 -1721 451 -1719
rect 457 -1715 458 -1713
rect 457 -1721 458 -1719
rect 464 -1715 465 -1713
rect 464 -1721 465 -1719
rect 471 -1715 472 -1713
rect 471 -1721 472 -1719
rect 478 -1715 479 -1713
rect 481 -1715 482 -1713
rect 485 -1715 486 -1713
rect 488 -1715 489 -1713
rect 485 -1721 486 -1719
rect 488 -1721 489 -1719
rect 492 -1721 493 -1719
rect 495 -1721 496 -1719
rect 499 -1715 500 -1713
rect 499 -1721 500 -1719
rect 506 -1715 507 -1713
rect 506 -1721 507 -1719
rect 513 -1715 514 -1713
rect 513 -1721 514 -1719
rect 523 -1715 524 -1713
rect 520 -1721 521 -1719
rect 523 -1721 524 -1719
rect 527 -1715 528 -1713
rect 527 -1721 528 -1719
rect 530 -1721 531 -1719
rect 534 -1715 535 -1713
rect 534 -1721 535 -1719
rect 541 -1715 542 -1713
rect 541 -1721 542 -1719
rect 548 -1715 549 -1713
rect 548 -1721 549 -1719
rect 555 -1715 556 -1713
rect 555 -1721 556 -1719
rect 562 -1715 563 -1713
rect 562 -1721 563 -1719
rect 569 -1715 570 -1713
rect 569 -1721 570 -1719
rect 579 -1715 580 -1713
rect 576 -1721 577 -1719
rect 579 -1721 580 -1719
rect 586 -1715 587 -1713
rect 586 -1721 587 -1719
rect 590 -1715 591 -1713
rect 590 -1721 591 -1719
rect 597 -1715 598 -1713
rect 597 -1721 598 -1719
rect 607 -1715 608 -1713
rect 604 -1721 605 -1719
rect 607 -1721 608 -1719
rect 611 -1715 612 -1713
rect 611 -1721 612 -1719
rect 618 -1715 619 -1713
rect 618 -1721 619 -1719
rect 625 -1715 626 -1713
rect 625 -1721 626 -1719
rect 632 -1715 633 -1713
rect 632 -1721 633 -1719
rect 639 -1715 640 -1713
rect 639 -1721 640 -1719
rect 646 -1715 647 -1713
rect 646 -1721 647 -1719
rect 653 -1715 654 -1713
rect 656 -1715 657 -1713
rect 653 -1721 654 -1719
rect 660 -1715 661 -1713
rect 663 -1715 664 -1713
rect 660 -1721 661 -1719
rect 667 -1715 668 -1713
rect 667 -1721 668 -1719
rect 674 -1715 675 -1713
rect 674 -1721 675 -1719
rect 677 -1721 678 -1719
rect 681 -1715 682 -1713
rect 681 -1721 682 -1719
rect 691 -1715 692 -1713
rect 688 -1721 689 -1719
rect 695 -1715 696 -1713
rect 695 -1721 696 -1719
rect 702 -1715 703 -1713
rect 702 -1721 703 -1719
rect 709 -1715 710 -1713
rect 709 -1721 710 -1719
rect 716 -1715 717 -1713
rect 716 -1721 717 -1719
rect 723 -1715 724 -1713
rect 723 -1721 724 -1719
rect 730 -1715 731 -1713
rect 730 -1721 731 -1719
rect 737 -1715 738 -1713
rect 737 -1721 738 -1719
rect 744 -1715 745 -1713
rect 744 -1721 745 -1719
rect 751 -1715 752 -1713
rect 751 -1721 752 -1719
rect 758 -1715 759 -1713
rect 761 -1715 762 -1713
rect 761 -1721 762 -1719
rect 765 -1715 766 -1713
rect 765 -1721 766 -1719
rect 772 -1715 773 -1713
rect 772 -1721 773 -1719
rect 779 -1715 780 -1713
rect 779 -1721 780 -1719
rect 786 -1715 787 -1713
rect 786 -1721 787 -1719
rect 793 -1715 794 -1713
rect 793 -1721 794 -1719
rect 800 -1715 801 -1713
rect 800 -1721 801 -1719
rect 807 -1715 808 -1713
rect 807 -1721 808 -1719
rect 817 -1721 818 -1719
rect 821 -1715 822 -1713
rect 821 -1721 822 -1719
rect 828 -1715 829 -1713
rect 828 -1721 829 -1719
rect 835 -1715 836 -1713
rect 835 -1721 836 -1719
rect 842 -1715 843 -1713
rect 842 -1721 843 -1719
rect 849 -1715 850 -1713
rect 849 -1721 850 -1719
rect 856 -1715 857 -1713
rect 856 -1721 857 -1719
rect 863 -1715 864 -1713
rect 863 -1721 864 -1719
rect 870 -1715 871 -1713
rect 870 -1721 871 -1719
rect 877 -1715 878 -1713
rect 877 -1721 878 -1719
rect 884 -1715 885 -1713
rect 884 -1721 885 -1719
rect 891 -1715 892 -1713
rect 891 -1721 892 -1719
rect 898 -1715 899 -1713
rect 898 -1721 899 -1719
rect 905 -1715 906 -1713
rect 905 -1721 906 -1719
rect 908 -1721 909 -1719
rect 912 -1715 913 -1713
rect 912 -1721 913 -1719
rect 919 -1715 920 -1713
rect 919 -1721 920 -1719
rect 926 -1721 927 -1719
rect 929 -1721 930 -1719
rect 933 -1715 934 -1713
rect 933 -1721 934 -1719
rect 940 -1715 941 -1713
rect 940 -1721 941 -1719
rect 947 -1715 948 -1713
rect 947 -1721 948 -1719
rect 954 -1715 955 -1713
rect 954 -1721 955 -1719
rect 961 -1715 962 -1713
rect 961 -1721 962 -1719
rect 968 -1715 969 -1713
rect 968 -1721 969 -1719
rect 1066 -1715 1067 -1713
rect 1069 -1721 1070 -1719
rect 1094 -1715 1095 -1713
rect 1094 -1721 1095 -1719
rect 2 -1806 3 -1804
rect 2 -1812 3 -1810
rect 9 -1812 10 -1810
rect 16 -1806 17 -1804
rect 16 -1812 17 -1810
rect 23 -1806 24 -1804
rect 23 -1812 24 -1810
rect 30 -1806 31 -1804
rect 30 -1812 31 -1810
rect 37 -1806 38 -1804
rect 37 -1812 38 -1810
rect 44 -1806 45 -1804
rect 44 -1812 45 -1810
rect 51 -1806 52 -1804
rect 51 -1812 52 -1810
rect 58 -1806 59 -1804
rect 58 -1812 59 -1810
rect 65 -1806 66 -1804
rect 65 -1812 66 -1810
rect 72 -1806 73 -1804
rect 72 -1812 73 -1810
rect 79 -1806 80 -1804
rect 79 -1812 80 -1810
rect 86 -1806 87 -1804
rect 86 -1812 87 -1810
rect 93 -1812 94 -1810
rect 96 -1812 97 -1810
rect 100 -1806 101 -1804
rect 100 -1812 101 -1810
rect 103 -1812 104 -1810
rect 107 -1806 108 -1804
rect 107 -1812 108 -1810
rect 117 -1806 118 -1804
rect 114 -1812 115 -1810
rect 117 -1812 118 -1810
rect 121 -1806 122 -1804
rect 121 -1812 122 -1810
rect 128 -1806 129 -1804
rect 128 -1812 129 -1810
rect 135 -1806 136 -1804
rect 138 -1806 139 -1804
rect 135 -1812 136 -1810
rect 142 -1806 143 -1804
rect 142 -1812 143 -1810
rect 149 -1806 150 -1804
rect 149 -1812 150 -1810
rect 156 -1806 157 -1804
rect 156 -1812 157 -1810
rect 163 -1806 164 -1804
rect 163 -1812 164 -1810
rect 170 -1806 171 -1804
rect 170 -1812 171 -1810
rect 177 -1806 178 -1804
rect 177 -1812 178 -1810
rect 184 -1806 185 -1804
rect 191 -1806 192 -1804
rect 191 -1812 192 -1810
rect 198 -1806 199 -1804
rect 198 -1812 199 -1810
rect 201 -1812 202 -1810
rect 205 -1812 206 -1810
rect 208 -1812 209 -1810
rect 212 -1806 213 -1804
rect 212 -1812 213 -1810
rect 219 -1806 220 -1804
rect 222 -1806 223 -1804
rect 219 -1812 220 -1810
rect 226 -1806 227 -1804
rect 226 -1812 227 -1810
rect 233 -1806 234 -1804
rect 233 -1812 234 -1810
rect 240 -1806 241 -1804
rect 240 -1812 241 -1810
rect 247 -1806 248 -1804
rect 247 -1812 248 -1810
rect 250 -1812 251 -1810
rect 254 -1806 255 -1804
rect 254 -1812 255 -1810
rect 261 -1806 262 -1804
rect 261 -1812 262 -1810
rect 268 -1806 269 -1804
rect 268 -1812 269 -1810
rect 275 -1806 276 -1804
rect 275 -1812 276 -1810
rect 282 -1806 283 -1804
rect 282 -1812 283 -1810
rect 289 -1806 290 -1804
rect 289 -1812 290 -1810
rect 296 -1806 297 -1804
rect 296 -1812 297 -1810
rect 303 -1806 304 -1804
rect 306 -1806 307 -1804
rect 306 -1812 307 -1810
rect 310 -1806 311 -1804
rect 310 -1812 311 -1810
rect 317 -1806 318 -1804
rect 317 -1812 318 -1810
rect 324 -1806 325 -1804
rect 324 -1812 325 -1810
rect 331 -1806 332 -1804
rect 331 -1812 332 -1810
rect 338 -1806 339 -1804
rect 338 -1812 339 -1810
rect 348 -1806 349 -1804
rect 348 -1812 349 -1810
rect 352 -1806 353 -1804
rect 352 -1812 353 -1810
rect 355 -1812 356 -1810
rect 359 -1806 360 -1804
rect 359 -1812 360 -1810
rect 366 -1806 367 -1804
rect 366 -1812 367 -1810
rect 373 -1806 374 -1804
rect 373 -1812 374 -1810
rect 380 -1806 381 -1804
rect 380 -1812 381 -1810
rect 387 -1806 388 -1804
rect 387 -1812 388 -1810
rect 394 -1806 395 -1804
rect 394 -1812 395 -1810
rect 401 -1806 402 -1804
rect 401 -1812 402 -1810
rect 408 -1806 409 -1804
rect 408 -1812 409 -1810
rect 415 -1806 416 -1804
rect 418 -1806 419 -1804
rect 415 -1812 416 -1810
rect 418 -1812 419 -1810
rect 425 -1806 426 -1804
rect 422 -1812 423 -1810
rect 425 -1812 426 -1810
rect 429 -1806 430 -1804
rect 432 -1806 433 -1804
rect 429 -1812 430 -1810
rect 432 -1812 433 -1810
rect 436 -1806 437 -1804
rect 436 -1812 437 -1810
rect 443 -1806 444 -1804
rect 443 -1812 444 -1810
rect 450 -1806 451 -1804
rect 450 -1812 451 -1810
rect 457 -1806 458 -1804
rect 457 -1812 458 -1810
rect 464 -1806 465 -1804
rect 464 -1812 465 -1810
rect 471 -1806 472 -1804
rect 471 -1812 472 -1810
rect 478 -1806 479 -1804
rect 478 -1812 479 -1810
rect 485 -1806 486 -1804
rect 485 -1812 486 -1810
rect 492 -1806 493 -1804
rect 492 -1812 493 -1810
rect 499 -1806 500 -1804
rect 502 -1806 503 -1804
rect 499 -1812 500 -1810
rect 506 -1806 507 -1804
rect 506 -1812 507 -1810
rect 513 -1806 514 -1804
rect 513 -1812 514 -1810
rect 520 -1806 521 -1804
rect 520 -1812 521 -1810
rect 523 -1812 524 -1810
rect 527 -1806 528 -1804
rect 530 -1806 531 -1804
rect 527 -1812 528 -1810
rect 534 -1806 535 -1804
rect 534 -1812 535 -1810
rect 541 -1806 542 -1804
rect 541 -1812 542 -1810
rect 548 -1806 549 -1804
rect 551 -1812 552 -1810
rect 555 -1806 556 -1804
rect 555 -1812 556 -1810
rect 562 -1806 563 -1804
rect 562 -1812 563 -1810
rect 569 -1806 570 -1804
rect 569 -1812 570 -1810
rect 576 -1806 577 -1804
rect 576 -1812 577 -1810
rect 583 -1806 584 -1804
rect 583 -1812 584 -1810
rect 590 -1806 591 -1804
rect 590 -1812 591 -1810
rect 597 -1806 598 -1804
rect 600 -1806 601 -1804
rect 604 -1806 605 -1804
rect 604 -1812 605 -1810
rect 611 -1806 612 -1804
rect 611 -1812 612 -1810
rect 614 -1812 615 -1810
rect 618 -1806 619 -1804
rect 618 -1812 619 -1810
rect 625 -1806 626 -1804
rect 625 -1812 626 -1810
rect 628 -1812 629 -1810
rect 632 -1806 633 -1804
rect 632 -1812 633 -1810
rect 639 -1806 640 -1804
rect 639 -1812 640 -1810
rect 646 -1806 647 -1804
rect 646 -1812 647 -1810
rect 653 -1806 654 -1804
rect 653 -1812 654 -1810
rect 660 -1806 661 -1804
rect 660 -1812 661 -1810
rect 667 -1806 668 -1804
rect 670 -1806 671 -1804
rect 670 -1812 671 -1810
rect 674 -1806 675 -1804
rect 674 -1812 675 -1810
rect 681 -1806 682 -1804
rect 681 -1812 682 -1810
rect 688 -1806 689 -1804
rect 691 -1806 692 -1804
rect 691 -1812 692 -1810
rect 695 -1806 696 -1804
rect 695 -1812 696 -1810
rect 702 -1806 703 -1804
rect 702 -1812 703 -1810
rect 712 -1806 713 -1804
rect 709 -1812 710 -1810
rect 712 -1812 713 -1810
rect 716 -1806 717 -1804
rect 716 -1812 717 -1810
rect 723 -1806 724 -1804
rect 723 -1812 724 -1810
rect 730 -1806 731 -1804
rect 730 -1812 731 -1810
rect 737 -1806 738 -1804
rect 737 -1812 738 -1810
rect 744 -1806 745 -1804
rect 744 -1812 745 -1810
rect 751 -1806 752 -1804
rect 751 -1812 752 -1810
rect 758 -1806 759 -1804
rect 758 -1812 759 -1810
rect 765 -1806 766 -1804
rect 765 -1812 766 -1810
rect 772 -1806 773 -1804
rect 772 -1812 773 -1810
rect 779 -1806 780 -1804
rect 779 -1812 780 -1810
rect 786 -1806 787 -1804
rect 786 -1812 787 -1810
rect 793 -1806 794 -1804
rect 793 -1812 794 -1810
rect 800 -1806 801 -1804
rect 800 -1812 801 -1810
rect 807 -1806 808 -1804
rect 807 -1812 808 -1810
rect 814 -1806 815 -1804
rect 814 -1812 815 -1810
rect 821 -1806 822 -1804
rect 821 -1812 822 -1810
rect 828 -1806 829 -1804
rect 828 -1812 829 -1810
rect 835 -1806 836 -1804
rect 835 -1812 836 -1810
rect 842 -1806 843 -1804
rect 842 -1812 843 -1810
rect 849 -1806 850 -1804
rect 849 -1812 850 -1810
rect 856 -1806 857 -1804
rect 856 -1812 857 -1810
rect 863 -1806 864 -1804
rect 863 -1812 864 -1810
rect 870 -1806 871 -1804
rect 870 -1812 871 -1810
rect 877 -1806 878 -1804
rect 877 -1812 878 -1810
rect 884 -1806 885 -1804
rect 884 -1812 885 -1810
rect 891 -1806 892 -1804
rect 891 -1812 892 -1810
rect 898 -1806 899 -1804
rect 898 -1812 899 -1810
rect 905 -1806 906 -1804
rect 905 -1812 906 -1810
rect 912 -1806 913 -1804
rect 912 -1812 913 -1810
rect 919 -1806 920 -1804
rect 919 -1812 920 -1810
rect 926 -1806 927 -1804
rect 926 -1812 927 -1810
rect 933 -1812 934 -1810
rect 940 -1806 941 -1804
rect 940 -1812 941 -1810
rect 947 -1806 948 -1804
rect 947 -1812 948 -1810
rect 954 -1806 955 -1804
rect 954 -1812 955 -1810
rect 961 -1806 962 -1804
rect 961 -1812 962 -1810
rect 968 -1806 969 -1804
rect 968 -1812 969 -1810
rect 975 -1806 976 -1804
rect 975 -1812 976 -1810
rect 982 -1806 983 -1804
rect 982 -1812 983 -1810
rect 989 -1806 990 -1804
rect 989 -1812 990 -1810
rect 996 -1806 997 -1804
rect 996 -1812 997 -1810
rect 1003 -1806 1004 -1804
rect 1003 -1812 1004 -1810
rect 1010 -1806 1011 -1804
rect 1010 -1812 1011 -1810
rect 1017 -1806 1018 -1804
rect 1017 -1812 1018 -1810
rect 1024 -1806 1025 -1804
rect 1024 -1812 1025 -1810
rect 1031 -1806 1032 -1804
rect 1031 -1812 1032 -1810
rect 1038 -1806 1039 -1804
rect 1038 -1812 1039 -1810
rect 1045 -1806 1046 -1804
rect 1045 -1812 1046 -1810
rect 1052 -1806 1053 -1804
rect 1055 -1806 1056 -1804
rect 1055 -1812 1056 -1810
rect 1059 -1806 1060 -1804
rect 1059 -1812 1060 -1810
rect 1087 -1806 1088 -1804
rect 1087 -1812 1088 -1810
rect 1094 -1806 1095 -1804
rect 1094 -1812 1095 -1810
rect 5 -1897 6 -1895
rect 9 -1897 10 -1895
rect 9 -1903 10 -1901
rect 16 -1897 17 -1895
rect 19 -1903 20 -1901
rect 23 -1897 24 -1895
rect 23 -1903 24 -1901
rect 30 -1897 31 -1895
rect 30 -1903 31 -1901
rect 40 -1897 41 -1895
rect 40 -1903 41 -1901
rect 44 -1897 45 -1895
rect 47 -1897 48 -1895
rect 44 -1903 45 -1901
rect 47 -1903 48 -1901
rect 51 -1897 52 -1895
rect 54 -1897 55 -1895
rect 51 -1903 52 -1901
rect 54 -1903 55 -1901
rect 58 -1897 59 -1895
rect 58 -1903 59 -1901
rect 65 -1897 66 -1895
rect 68 -1897 69 -1895
rect 72 -1897 73 -1895
rect 72 -1903 73 -1901
rect 79 -1897 80 -1895
rect 82 -1897 83 -1895
rect 82 -1903 83 -1901
rect 86 -1897 87 -1895
rect 86 -1903 87 -1901
rect 93 -1897 94 -1895
rect 93 -1903 94 -1901
rect 100 -1897 101 -1895
rect 100 -1903 101 -1901
rect 107 -1897 108 -1895
rect 107 -1903 108 -1901
rect 114 -1897 115 -1895
rect 117 -1897 118 -1895
rect 117 -1903 118 -1901
rect 121 -1897 122 -1895
rect 124 -1897 125 -1895
rect 121 -1903 122 -1901
rect 124 -1903 125 -1901
rect 128 -1897 129 -1895
rect 128 -1903 129 -1901
rect 135 -1897 136 -1895
rect 135 -1903 136 -1901
rect 142 -1897 143 -1895
rect 142 -1903 143 -1901
rect 149 -1903 150 -1901
rect 152 -1903 153 -1901
rect 156 -1897 157 -1895
rect 156 -1903 157 -1901
rect 159 -1903 160 -1901
rect 163 -1897 164 -1895
rect 163 -1903 164 -1901
rect 170 -1897 171 -1895
rect 170 -1903 171 -1901
rect 177 -1897 178 -1895
rect 177 -1903 178 -1901
rect 184 -1897 185 -1895
rect 184 -1903 185 -1901
rect 194 -1897 195 -1895
rect 194 -1903 195 -1901
rect 198 -1897 199 -1895
rect 198 -1903 199 -1901
rect 205 -1897 206 -1895
rect 205 -1903 206 -1901
rect 212 -1897 213 -1895
rect 212 -1903 213 -1901
rect 222 -1903 223 -1901
rect 226 -1897 227 -1895
rect 226 -1903 227 -1901
rect 233 -1897 234 -1895
rect 233 -1903 234 -1901
rect 240 -1897 241 -1895
rect 240 -1903 241 -1901
rect 247 -1897 248 -1895
rect 247 -1903 248 -1901
rect 254 -1897 255 -1895
rect 254 -1903 255 -1901
rect 261 -1897 262 -1895
rect 261 -1903 262 -1901
rect 268 -1897 269 -1895
rect 268 -1903 269 -1901
rect 275 -1897 276 -1895
rect 275 -1903 276 -1901
rect 282 -1897 283 -1895
rect 282 -1903 283 -1901
rect 289 -1897 290 -1895
rect 289 -1903 290 -1901
rect 296 -1897 297 -1895
rect 296 -1903 297 -1901
rect 303 -1897 304 -1895
rect 303 -1903 304 -1901
rect 310 -1897 311 -1895
rect 310 -1903 311 -1901
rect 317 -1897 318 -1895
rect 317 -1903 318 -1901
rect 324 -1897 325 -1895
rect 324 -1903 325 -1901
rect 331 -1897 332 -1895
rect 331 -1903 332 -1901
rect 338 -1897 339 -1895
rect 338 -1903 339 -1901
rect 345 -1897 346 -1895
rect 345 -1903 346 -1901
rect 352 -1897 353 -1895
rect 352 -1903 353 -1901
rect 359 -1897 360 -1895
rect 362 -1897 363 -1895
rect 359 -1903 360 -1901
rect 366 -1897 367 -1895
rect 369 -1897 370 -1895
rect 366 -1903 367 -1901
rect 369 -1903 370 -1901
rect 373 -1897 374 -1895
rect 373 -1903 374 -1901
rect 380 -1897 381 -1895
rect 380 -1903 381 -1901
rect 387 -1897 388 -1895
rect 390 -1897 391 -1895
rect 390 -1903 391 -1901
rect 394 -1897 395 -1895
rect 394 -1903 395 -1901
rect 401 -1897 402 -1895
rect 401 -1903 402 -1901
rect 408 -1897 409 -1895
rect 408 -1903 409 -1901
rect 418 -1897 419 -1895
rect 415 -1903 416 -1901
rect 422 -1897 423 -1895
rect 422 -1903 423 -1901
rect 429 -1897 430 -1895
rect 429 -1903 430 -1901
rect 436 -1897 437 -1895
rect 436 -1903 437 -1901
rect 443 -1897 444 -1895
rect 446 -1897 447 -1895
rect 450 -1897 451 -1895
rect 453 -1903 454 -1901
rect 457 -1897 458 -1895
rect 457 -1903 458 -1901
rect 464 -1897 465 -1895
rect 464 -1903 465 -1901
rect 471 -1897 472 -1895
rect 471 -1903 472 -1901
rect 478 -1897 479 -1895
rect 481 -1897 482 -1895
rect 478 -1903 479 -1901
rect 481 -1903 482 -1901
rect 485 -1897 486 -1895
rect 488 -1897 489 -1895
rect 485 -1903 486 -1901
rect 492 -1897 493 -1895
rect 492 -1903 493 -1901
rect 502 -1897 503 -1895
rect 499 -1903 500 -1901
rect 502 -1903 503 -1901
rect 506 -1897 507 -1895
rect 506 -1903 507 -1901
rect 513 -1897 514 -1895
rect 513 -1903 514 -1901
rect 520 -1897 521 -1895
rect 520 -1903 521 -1901
rect 527 -1903 528 -1901
rect 530 -1903 531 -1901
rect 534 -1897 535 -1895
rect 534 -1903 535 -1901
rect 541 -1897 542 -1895
rect 541 -1903 542 -1901
rect 548 -1897 549 -1895
rect 551 -1897 552 -1895
rect 548 -1903 549 -1901
rect 551 -1903 552 -1901
rect 555 -1897 556 -1895
rect 558 -1897 559 -1895
rect 558 -1903 559 -1901
rect 562 -1897 563 -1895
rect 562 -1903 563 -1901
rect 569 -1897 570 -1895
rect 569 -1903 570 -1901
rect 576 -1897 577 -1895
rect 576 -1903 577 -1901
rect 583 -1897 584 -1895
rect 583 -1903 584 -1901
rect 590 -1897 591 -1895
rect 590 -1903 591 -1901
rect 597 -1897 598 -1895
rect 597 -1903 598 -1901
rect 604 -1897 605 -1895
rect 604 -1903 605 -1901
rect 611 -1897 612 -1895
rect 611 -1903 612 -1901
rect 621 -1897 622 -1895
rect 618 -1903 619 -1901
rect 621 -1903 622 -1901
rect 625 -1897 626 -1895
rect 625 -1903 626 -1901
rect 632 -1897 633 -1895
rect 635 -1897 636 -1895
rect 632 -1903 633 -1901
rect 635 -1903 636 -1901
rect 639 -1897 640 -1895
rect 639 -1903 640 -1901
rect 646 -1897 647 -1895
rect 646 -1903 647 -1901
rect 653 -1897 654 -1895
rect 653 -1903 654 -1901
rect 660 -1897 661 -1895
rect 660 -1903 661 -1901
rect 667 -1897 668 -1895
rect 670 -1897 671 -1895
rect 667 -1903 668 -1901
rect 670 -1903 671 -1901
rect 674 -1897 675 -1895
rect 674 -1903 675 -1901
rect 681 -1897 682 -1895
rect 681 -1903 682 -1901
rect 688 -1897 689 -1895
rect 688 -1903 689 -1901
rect 695 -1897 696 -1895
rect 695 -1903 696 -1901
rect 702 -1897 703 -1895
rect 702 -1903 703 -1901
rect 709 -1897 710 -1895
rect 709 -1903 710 -1901
rect 716 -1897 717 -1895
rect 716 -1903 717 -1901
rect 723 -1897 724 -1895
rect 723 -1903 724 -1901
rect 730 -1897 731 -1895
rect 733 -1897 734 -1895
rect 730 -1903 731 -1901
rect 737 -1897 738 -1895
rect 737 -1903 738 -1901
rect 744 -1897 745 -1895
rect 744 -1903 745 -1901
rect 751 -1897 752 -1895
rect 751 -1903 752 -1901
rect 758 -1897 759 -1895
rect 758 -1903 759 -1901
rect 765 -1897 766 -1895
rect 765 -1903 766 -1901
rect 772 -1897 773 -1895
rect 772 -1903 773 -1901
rect 779 -1897 780 -1895
rect 779 -1903 780 -1901
rect 786 -1897 787 -1895
rect 786 -1903 787 -1901
rect 793 -1897 794 -1895
rect 793 -1903 794 -1901
rect 800 -1897 801 -1895
rect 800 -1903 801 -1901
rect 807 -1897 808 -1895
rect 807 -1903 808 -1901
rect 814 -1897 815 -1895
rect 814 -1903 815 -1901
rect 821 -1897 822 -1895
rect 821 -1903 822 -1901
rect 828 -1897 829 -1895
rect 828 -1903 829 -1901
rect 835 -1897 836 -1895
rect 835 -1903 836 -1901
rect 842 -1897 843 -1895
rect 842 -1903 843 -1901
rect 849 -1897 850 -1895
rect 849 -1903 850 -1901
rect 856 -1897 857 -1895
rect 856 -1903 857 -1901
rect 863 -1897 864 -1895
rect 863 -1903 864 -1901
rect 870 -1897 871 -1895
rect 870 -1903 871 -1901
rect 877 -1897 878 -1895
rect 877 -1903 878 -1901
rect 884 -1897 885 -1895
rect 884 -1903 885 -1901
rect 891 -1897 892 -1895
rect 891 -1903 892 -1901
rect 898 -1897 899 -1895
rect 898 -1903 899 -1901
rect 905 -1897 906 -1895
rect 905 -1903 906 -1901
rect 912 -1897 913 -1895
rect 912 -1903 913 -1901
rect 919 -1897 920 -1895
rect 919 -1903 920 -1901
rect 926 -1897 927 -1895
rect 926 -1903 927 -1901
rect 933 -1897 934 -1895
rect 933 -1903 934 -1901
rect 940 -1897 941 -1895
rect 940 -1903 941 -1901
rect 947 -1897 948 -1895
rect 947 -1903 948 -1901
rect 954 -1897 955 -1895
rect 954 -1903 955 -1901
rect 961 -1897 962 -1895
rect 961 -1903 962 -1901
rect 968 -1897 969 -1895
rect 968 -1903 969 -1901
rect 975 -1897 976 -1895
rect 975 -1903 976 -1901
rect 982 -1897 983 -1895
rect 982 -1903 983 -1901
rect 989 -1897 990 -1895
rect 989 -1903 990 -1901
rect 996 -1897 997 -1895
rect 996 -1903 997 -1901
rect 1003 -1897 1004 -1895
rect 1003 -1903 1004 -1901
rect 1010 -1897 1011 -1895
rect 1010 -1903 1011 -1901
rect 1017 -1897 1018 -1895
rect 1017 -1903 1018 -1901
rect 1024 -1897 1025 -1895
rect 1024 -1903 1025 -1901
rect 1031 -1897 1032 -1895
rect 1031 -1903 1032 -1901
rect 1038 -1897 1039 -1895
rect 1038 -1903 1039 -1901
rect 1045 -1897 1046 -1895
rect 1045 -1903 1046 -1901
rect 1052 -1897 1053 -1895
rect 1052 -1903 1053 -1901
rect 1059 -1897 1060 -1895
rect 1059 -1903 1060 -1901
rect 1069 -1897 1070 -1895
rect 1066 -1903 1067 -1901
rect 1069 -1903 1070 -1901
rect 1073 -1897 1074 -1895
rect 1073 -1903 1074 -1901
rect 1087 -1897 1088 -1895
rect 1087 -1903 1088 -1901
rect 1101 -1897 1102 -1895
rect 1101 -1903 1102 -1901
rect 2 -2002 3 -2000
rect 9 -2002 10 -2000
rect 9 -2008 10 -2006
rect 16 -2002 17 -2000
rect 16 -2008 17 -2006
rect 23 -2002 24 -2000
rect 26 -2008 27 -2006
rect 30 -2002 31 -2000
rect 33 -2002 34 -2000
rect 30 -2008 31 -2006
rect 33 -2008 34 -2006
rect 37 -2002 38 -2000
rect 37 -2008 38 -2006
rect 44 -2002 45 -2000
rect 44 -2008 45 -2006
rect 54 -2002 55 -2000
rect 51 -2008 52 -2006
rect 54 -2008 55 -2006
rect 58 -2002 59 -2000
rect 61 -2002 62 -2000
rect 58 -2008 59 -2006
rect 65 -2002 66 -2000
rect 65 -2008 66 -2006
rect 75 -2002 76 -2000
rect 75 -2008 76 -2006
rect 79 -2008 80 -2006
rect 86 -2008 87 -2006
rect 89 -2008 90 -2006
rect 93 -2002 94 -2000
rect 93 -2008 94 -2006
rect 100 -2002 101 -2000
rect 100 -2008 101 -2006
rect 107 -2002 108 -2000
rect 107 -2008 108 -2006
rect 110 -2008 111 -2006
rect 114 -2002 115 -2000
rect 114 -2008 115 -2006
rect 121 -2002 122 -2000
rect 121 -2008 122 -2006
rect 128 -2002 129 -2000
rect 128 -2008 129 -2006
rect 135 -2008 136 -2006
rect 138 -2008 139 -2006
rect 142 -2002 143 -2000
rect 142 -2008 143 -2006
rect 149 -2002 150 -2000
rect 152 -2002 153 -2000
rect 149 -2008 150 -2006
rect 152 -2008 153 -2006
rect 156 -2002 157 -2000
rect 156 -2008 157 -2006
rect 163 -2002 164 -2000
rect 163 -2008 164 -2006
rect 170 -2002 171 -2000
rect 170 -2008 171 -2006
rect 180 -2002 181 -2000
rect 177 -2008 178 -2006
rect 180 -2008 181 -2006
rect 184 -2002 185 -2000
rect 184 -2008 185 -2006
rect 191 -2002 192 -2000
rect 191 -2008 192 -2006
rect 198 -2002 199 -2000
rect 198 -2008 199 -2006
rect 205 -2002 206 -2000
rect 208 -2002 209 -2000
rect 212 -2002 213 -2000
rect 212 -2008 213 -2006
rect 219 -2002 220 -2000
rect 222 -2002 223 -2000
rect 222 -2008 223 -2006
rect 229 -2002 230 -2000
rect 226 -2008 227 -2006
rect 229 -2008 230 -2006
rect 233 -2002 234 -2000
rect 233 -2008 234 -2006
rect 240 -2002 241 -2000
rect 240 -2008 241 -2006
rect 247 -2002 248 -2000
rect 247 -2008 248 -2006
rect 254 -2002 255 -2000
rect 254 -2008 255 -2006
rect 261 -2002 262 -2000
rect 261 -2008 262 -2006
rect 268 -2002 269 -2000
rect 268 -2008 269 -2006
rect 275 -2002 276 -2000
rect 275 -2008 276 -2006
rect 282 -2002 283 -2000
rect 282 -2008 283 -2006
rect 289 -2002 290 -2000
rect 289 -2008 290 -2006
rect 296 -2002 297 -2000
rect 296 -2008 297 -2006
rect 303 -2002 304 -2000
rect 303 -2008 304 -2006
rect 310 -2002 311 -2000
rect 310 -2008 311 -2006
rect 317 -2002 318 -2000
rect 317 -2008 318 -2006
rect 324 -2002 325 -2000
rect 324 -2008 325 -2006
rect 331 -2002 332 -2000
rect 331 -2008 332 -2006
rect 338 -2002 339 -2000
rect 338 -2008 339 -2006
rect 345 -2002 346 -2000
rect 348 -2002 349 -2000
rect 345 -2008 346 -2006
rect 348 -2008 349 -2006
rect 352 -2002 353 -2000
rect 352 -2008 353 -2006
rect 359 -2002 360 -2000
rect 359 -2008 360 -2006
rect 366 -2002 367 -2000
rect 369 -2002 370 -2000
rect 366 -2008 367 -2006
rect 369 -2008 370 -2006
rect 373 -2002 374 -2000
rect 376 -2002 377 -2000
rect 373 -2008 374 -2006
rect 376 -2008 377 -2006
rect 380 -2002 381 -2000
rect 380 -2008 381 -2006
rect 387 -2002 388 -2000
rect 387 -2008 388 -2006
rect 394 -2002 395 -2000
rect 394 -2008 395 -2006
rect 401 -2002 402 -2000
rect 401 -2008 402 -2006
rect 408 -2002 409 -2000
rect 408 -2008 409 -2006
rect 411 -2008 412 -2006
rect 415 -2002 416 -2000
rect 415 -2008 416 -2006
rect 422 -2002 423 -2000
rect 422 -2008 423 -2006
rect 429 -2002 430 -2000
rect 429 -2008 430 -2006
rect 436 -2002 437 -2000
rect 439 -2008 440 -2006
rect 443 -2002 444 -2000
rect 443 -2008 444 -2006
rect 450 -2002 451 -2000
rect 450 -2008 451 -2006
rect 457 -2002 458 -2000
rect 457 -2008 458 -2006
rect 464 -2002 465 -2000
rect 464 -2008 465 -2006
rect 471 -2002 472 -2000
rect 471 -2008 472 -2006
rect 478 -2002 479 -2000
rect 478 -2008 479 -2006
rect 485 -2002 486 -2000
rect 485 -2008 486 -2006
rect 492 -2002 493 -2000
rect 492 -2008 493 -2006
rect 499 -2002 500 -2000
rect 499 -2008 500 -2006
rect 506 -2002 507 -2000
rect 506 -2008 507 -2006
rect 516 -2002 517 -2000
rect 516 -2008 517 -2006
rect 520 -2002 521 -2000
rect 520 -2008 521 -2006
rect 527 -2002 528 -2000
rect 530 -2002 531 -2000
rect 527 -2008 528 -2006
rect 530 -2008 531 -2006
rect 534 -2002 535 -2000
rect 534 -2008 535 -2006
rect 541 -2002 542 -2000
rect 541 -2008 542 -2006
rect 548 -2002 549 -2000
rect 548 -2008 549 -2006
rect 555 -2002 556 -2000
rect 555 -2008 556 -2006
rect 562 -2002 563 -2000
rect 562 -2008 563 -2006
rect 569 -2002 570 -2000
rect 569 -2008 570 -2006
rect 576 -2002 577 -2000
rect 576 -2008 577 -2006
rect 583 -2002 584 -2000
rect 583 -2008 584 -2006
rect 590 -2008 591 -2006
rect 593 -2008 594 -2006
rect 597 -2002 598 -2000
rect 597 -2008 598 -2006
rect 604 -2002 605 -2000
rect 604 -2008 605 -2006
rect 611 -2002 612 -2000
rect 611 -2008 612 -2006
rect 618 -2002 619 -2000
rect 621 -2002 622 -2000
rect 618 -2008 619 -2006
rect 625 -2002 626 -2000
rect 625 -2008 626 -2006
rect 635 -2002 636 -2000
rect 635 -2008 636 -2006
rect 639 -2002 640 -2000
rect 639 -2008 640 -2006
rect 646 -2002 647 -2000
rect 649 -2002 650 -2000
rect 646 -2008 647 -2006
rect 649 -2008 650 -2006
rect 653 -2002 654 -2000
rect 653 -2008 654 -2006
rect 660 -2002 661 -2000
rect 660 -2008 661 -2006
rect 667 -2002 668 -2000
rect 667 -2008 668 -2006
rect 674 -2002 675 -2000
rect 674 -2008 675 -2006
rect 681 -2002 682 -2000
rect 681 -2008 682 -2006
rect 688 -2002 689 -2000
rect 688 -2008 689 -2006
rect 695 -2002 696 -2000
rect 695 -2008 696 -2006
rect 702 -2002 703 -2000
rect 702 -2008 703 -2006
rect 709 -2002 710 -2000
rect 709 -2008 710 -2006
rect 716 -2002 717 -2000
rect 716 -2008 717 -2006
rect 723 -2002 724 -2000
rect 723 -2008 724 -2006
rect 730 -2002 731 -2000
rect 730 -2008 731 -2006
rect 737 -2002 738 -2000
rect 737 -2008 738 -2006
rect 744 -2008 745 -2006
rect 751 -2002 752 -2000
rect 751 -2008 752 -2006
rect 758 -2002 759 -2000
rect 758 -2008 759 -2006
rect 765 -2002 766 -2000
rect 768 -2002 769 -2000
rect 765 -2008 766 -2006
rect 768 -2008 769 -2006
rect 772 -2002 773 -2000
rect 772 -2008 773 -2006
rect 779 -2008 780 -2006
rect 782 -2008 783 -2006
rect 786 -2002 787 -2000
rect 786 -2008 787 -2006
rect 793 -2002 794 -2000
rect 793 -2008 794 -2006
rect 800 -2002 801 -2000
rect 800 -2008 801 -2006
rect 807 -2002 808 -2000
rect 807 -2008 808 -2006
rect 814 -2002 815 -2000
rect 814 -2008 815 -2006
rect 821 -2002 822 -2000
rect 821 -2008 822 -2006
rect 828 -2002 829 -2000
rect 828 -2008 829 -2006
rect 835 -2002 836 -2000
rect 835 -2008 836 -2006
rect 842 -2002 843 -2000
rect 842 -2008 843 -2006
rect 849 -2002 850 -2000
rect 849 -2008 850 -2006
rect 856 -2002 857 -2000
rect 856 -2008 857 -2006
rect 863 -2002 864 -2000
rect 863 -2008 864 -2006
rect 870 -2002 871 -2000
rect 870 -2008 871 -2006
rect 877 -2002 878 -2000
rect 877 -2008 878 -2006
rect 884 -2002 885 -2000
rect 884 -2008 885 -2006
rect 891 -2002 892 -2000
rect 891 -2008 892 -2006
rect 898 -2002 899 -2000
rect 898 -2008 899 -2006
rect 905 -2002 906 -2000
rect 905 -2008 906 -2006
rect 912 -2002 913 -2000
rect 912 -2008 913 -2006
rect 919 -2002 920 -2000
rect 919 -2008 920 -2006
rect 929 -2008 930 -2006
rect 933 -2002 934 -2000
rect 933 -2008 934 -2006
rect 940 -2002 941 -2000
rect 940 -2008 941 -2006
rect 947 -2002 948 -2000
rect 947 -2008 948 -2006
rect 954 -2002 955 -2000
rect 954 -2008 955 -2006
rect 961 -2002 962 -2000
rect 961 -2008 962 -2006
rect 968 -2002 969 -2000
rect 968 -2008 969 -2006
rect 975 -2002 976 -2000
rect 975 -2008 976 -2006
rect 982 -2002 983 -2000
rect 982 -2008 983 -2006
rect 989 -2002 990 -2000
rect 989 -2008 990 -2006
rect 996 -2002 997 -2000
rect 996 -2008 997 -2006
rect 1003 -2002 1004 -2000
rect 1003 -2008 1004 -2006
rect 1010 -2002 1011 -2000
rect 1010 -2008 1011 -2006
rect 1017 -2002 1018 -2000
rect 1017 -2008 1018 -2006
rect 1024 -2002 1025 -2000
rect 1024 -2008 1025 -2006
rect 1031 -2002 1032 -2000
rect 1031 -2008 1032 -2006
rect 1038 -2002 1039 -2000
rect 1038 -2008 1039 -2006
rect 1045 -2002 1046 -2000
rect 1045 -2008 1046 -2006
rect 1052 -2002 1053 -2000
rect 1052 -2008 1053 -2006
rect 1059 -2002 1060 -2000
rect 1059 -2008 1060 -2006
rect 1066 -2002 1067 -2000
rect 1066 -2008 1067 -2006
rect 1073 -2002 1074 -2000
rect 1073 -2008 1074 -2006
rect 1080 -2002 1081 -2000
rect 1080 -2008 1081 -2006
rect 1087 -2002 1088 -2000
rect 1087 -2008 1088 -2006
rect 1097 -2002 1098 -2000
rect 1094 -2008 1095 -2006
rect 1104 -2002 1105 -2000
rect 1101 -2008 1102 -2006
rect 1104 -2008 1105 -2006
rect 1108 -2002 1109 -2000
rect 1108 -2008 1109 -2006
rect 1115 -2002 1116 -2000
rect 1115 -2008 1116 -2006
rect 2 -2115 3 -2113
rect 2 -2121 3 -2119
rect 9 -2115 10 -2113
rect 9 -2121 10 -2119
rect 16 -2115 17 -2113
rect 16 -2121 17 -2119
rect 23 -2115 24 -2113
rect 23 -2121 24 -2119
rect 30 -2115 31 -2113
rect 30 -2121 31 -2119
rect 37 -2115 38 -2113
rect 37 -2121 38 -2119
rect 44 -2115 45 -2113
rect 44 -2121 45 -2119
rect 51 -2115 52 -2113
rect 51 -2121 52 -2119
rect 58 -2115 59 -2113
rect 58 -2121 59 -2119
rect 61 -2121 62 -2119
rect 65 -2115 66 -2113
rect 65 -2121 66 -2119
rect 72 -2115 73 -2113
rect 75 -2115 76 -2113
rect 72 -2121 73 -2119
rect 75 -2121 76 -2119
rect 79 -2115 80 -2113
rect 82 -2115 83 -2113
rect 79 -2121 80 -2119
rect 82 -2121 83 -2119
rect 86 -2115 87 -2113
rect 89 -2115 90 -2113
rect 86 -2121 87 -2119
rect 89 -2121 90 -2119
rect 93 -2115 94 -2113
rect 96 -2115 97 -2113
rect 93 -2121 94 -2119
rect 96 -2121 97 -2119
rect 100 -2115 101 -2113
rect 100 -2121 101 -2119
rect 107 -2115 108 -2113
rect 110 -2115 111 -2113
rect 107 -2121 108 -2119
rect 110 -2121 111 -2119
rect 114 -2115 115 -2113
rect 117 -2115 118 -2113
rect 117 -2121 118 -2119
rect 121 -2115 122 -2113
rect 121 -2121 122 -2119
rect 124 -2121 125 -2119
rect 128 -2115 129 -2113
rect 128 -2121 129 -2119
rect 135 -2115 136 -2113
rect 138 -2115 139 -2113
rect 138 -2121 139 -2119
rect 142 -2115 143 -2113
rect 142 -2121 143 -2119
rect 149 -2115 150 -2113
rect 152 -2115 153 -2113
rect 149 -2121 150 -2119
rect 152 -2121 153 -2119
rect 156 -2115 157 -2113
rect 156 -2121 157 -2119
rect 163 -2115 164 -2113
rect 163 -2121 164 -2119
rect 170 -2115 171 -2113
rect 170 -2121 171 -2119
rect 177 -2115 178 -2113
rect 177 -2121 178 -2119
rect 184 -2115 185 -2113
rect 184 -2121 185 -2119
rect 191 -2115 192 -2113
rect 191 -2121 192 -2119
rect 198 -2115 199 -2113
rect 198 -2121 199 -2119
rect 205 -2115 206 -2113
rect 205 -2121 206 -2119
rect 212 -2115 213 -2113
rect 212 -2121 213 -2119
rect 222 -2115 223 -2113
rect 226 -2115 227 -2113
rect 226 -2121 227 -2119
rect 233 -2115 234 -2113
rect 233 -2121 234 -2119
rect 240 -2115 241 -2113
rect 240 -2121 241 -2119
rect 247 -2115 248 -2113
rect 247 -2121 248 -2119
rect 254 -2115 255 -2113
rect 254 -2121 255 -2119
rect 261 -2115 262 -2113
rect 261 -2121 262 -2119
rect 268 -2115 269 -2113
rect 268 -2121 269 -2119
rect 275 -2115 276 -2113
rect 275 -2121 276 -2119
rect 282 -2115 283 -2113
rect 282 -2121 283 -2119
rect 289 -2115 290 -2113
rect 289 -2121 290 -2119
rect 292 -2121 293 -2119
rect 296 -2115 297 -2113
rect 296 -2121 297 -2119
rect 303 -2115 304 -2113
rect 303 -2121 304 -2119
rect 310 -2115 311 -2113
rect 310 -2121 311 -2119
rect 317 -2115 318 -2113
rect 317 -2121 318 -2119
rect 324 -2115 325 -2113
rect 324 -2121 325 -2119
rect 331 -2115 332 -2113
rect 331 -2121 332 -2119
rect 338 -2115 339 -2113
rect 341 -2115 342 -2113
rect 338 -2121 339 -2119
rect 341 -2121 342 -2119
rect 345 -2115 346 -2113
rect 345 -2121 346 -2119
rect 352 -2115 353 -2113
rect 355 -2115 356 -2113
rect 359 -2115 360 -2113
rect 359 -2121 360 -2119
rect 366 -2115 367 -2113
rect 366 -2121 367 -2119
rect 373 -2115 374 -2113
rect 373 -2121 374 -2119
rect 380 -2115 381 -2113
rect 380 -2121 381 -2119
rect 387 -2115 388 -2113
rect 387 -2121 388 -2119
rect 394 -2115 395 -2113
rect 394 -2121 395 -2119
rect 401 -2115 402 -2113
rect 401 -2121 402 -2119
rect 411 -2115 412 -2113
rect 408 -2121 409 -2119
rect 415 -2115 416 -2113
rect 418 -2115 419 -2113
rect 415 -2121 416 -2119
rect 418 -2121 419 -2119
rect 422 -2115 423 -2113
rect 422 -2121 423 -2119
rect 429 -2115 430 -2113
rect 429 -2121 430 -2119
rect 436 -2115 437 -2113
rect 436 -2121 437 -2119
rect 443 -2115 444 -2113
rect 443 -2121 444 -2119
rect 450 -2115 451 -2113
rect 453 -2115 454 -2113
rect 453 -2121 454 -2119
rect 460 -2115 461 -2113
rect 464 -2115 465 -2113
rect 464 -2121 465 -2119
rect 471 -2115 472 -2113
rect 471 -2121 472 -2119
rect 478 -2115 479 -2113
rect 478 -2121 479 -2119
rect 485 -2115 486 -2113
rect 485 -2121 486 -2119
rect 492 -2115 493 -2113
rect 492 -2121 493 -2119
rect 499 -2115 500 -2113
rect 502 -2115 503 -2113
rect 506 -2115 507 -2113
rect 506 -2121 507 -2119
rect 513 -2115 514 -2113
rect 513 -2121 514 -2119
rect 520 -2115 521 -2113
rect 520 -2121 521 -2119
rect 527 -2115 528 -2113
rect 527 -2121 528 -2119
rect 530 -2121 531 -2119
rect 534 -2115 535 -2113
rect 534 -2121 535 -2119
rect 541 -2115 542 -2113
rect 541 -2121 542 -2119
rect 548 -2115 549 -2113
rect 548 -2121 549 -2119
rect 551 -2121 552 -2119
rect 555 -2115 556 -2113
rect 555 -2121 556 -2119
rect 562 -2115 563 -2113
rect 562 -2121 563 -2119
rect 572 -2115 573 -2113
rect 569 -2121 570 -2119
rect 579 -2115 580 -2113
rect 576 -2121 577 -2119
rect 579 -2121 580 -2119
rect 583 -2115 584 -2113
rect 583 -2121 584 -2119
rect 590 -2115 591 -2113
rect 590 -2121 591 -2119
rect 597 -2115 598 -2113
rect 597 -2121 598 -2119
rect 604 -2115 605 -2113
rect 604 -2121 605 -2119
rect 614 -2115 615 -2113
rect 611 -2121 612 -2119
rect 618 -2115 619 -2113
rect 618 -2121 619 -2119
rect 625 -2121 626 -2119
rect 628 -2121 629 -2119
rect 632 -2115 633 -2113
rect 632 -2121 633 -2119
rect 639 -2115 640 -2113
rect 642 -2115 643 -2113
rect 639 -2121 640 -2119
rect 642 -2121 643 -2119
rect 646 -2115 647 -2113
rect 646 -2121 647 -2119
rect 653 -2115 654 -2113
rect 656 -2121 657 -2119
rect 660 -2115 661 -2113
rect 660 -2121 661 -2119
rect 667 -2115 668 -2113
rect 667 -2121 668 -2119
rect 674 -2115 675 -2113
rect 674 -2121 675 -2119
rect 681 -2115 682 -2113
rect 681 -2121 682 -2119
rect 688 -2115 689 -2113
rect 691 -2115 692 -2113
rect 691 -2121 692 -2119
rect 695 -2115 696 -2113
rect 695 -2121 696 -2119
rect 702 -2115 703 -2113
rect 702 -2121 703 -2119
rect 709 -2115 710 -2113
rect 709 -2121 710 -2119
rect 716 -2115 717 -2113
rect 716 -2121 717 -2119
rect 723 -2115 724 -2113
rect 723 -2121 724 -2119
rect 730 -2115 731 -2113
rect 730 -2121 731 -2119
rect 737 -2115 738 -2113
rect 737 -2121 738 -2119
rect 740 -2121 741 -2119
rect 744 -2115 745 -2113
rect 744 -2121 745 -2119
rect 751 -2115 752 -2113
rect 751 -2121 752 -2119
rect 758 -2115 759 -2113
rect 761 -2115 762 -2113
rect 758 -2121 759 -2119
rect 761 -2121 762 -2119
rect 765 -2115 766 -2113
rect 765 -2121 766 -2119
rect 772 -2115 773 -2113
rect 772 -2121 773 -2119
rect 779 -2115 780 -2113
rect 779 -2121 780 -2119
rect 786 -2115 787 -2113
rect 786 -2121 787 -2119
rect 793 -2115 794 -2113
rect 793 -2121 794 -2119
rect 800 -2115 801 -2113
rect 800 -2121 801 -2119
rect 807 -2115 808 -2113
rect 807 -2121 808 -2119
rect 814 -2115 815 -2113
rect 814 -2121 815 -2119
rect 821 -2115 822 -2113
rect 821 -2121 822 -2119
rect 828 -2115 829 -2113
rect 828 -2121 829 -2119
rect 835 -2115 836 -2113
rect 835 -2121 836 -2119
rect 842 -2115 843 -2113
rect 842 -2121 843 -2119
rect 849 -2115 850 -2113
rect 849 -2121 850 -2119
rect 856 -2115 857 -2113
rect 856 -2121 857 -2119
rect 863 -2115 864 -2113
rect 863 -2121 864 -2119
rect 870 -2115 871 -2113
rect 870 -2121 871 -2119
rect 877 -2115 878 -2113
rect 877 -2121 878 -2119
rect 884 -2115 885 -2113
rect 884 -2121 885 -2119
rect 891 -2115 892 -2113
rect 891 -2121 892 -2119
rect 898 -2115 899 -2113
rect 898 -2121 899 -2119
rect 905 -2115 906 -2113
rect 905 -2121 906 -2119
rect 912 -2115 913 -2113
rect 912 -2121 913 -2119
rect 919 -2115 920 -2113
rect 919 -2121 920 -2119
rect 926 -2115 927 -2113
rect 926 -2121 927 -2119
rect 933 -2115 934 -2113
rect 933 -2121 934 -2119
rect 943 -2115 944 -2113
rect 947 -2115 948 -2113
rect 947 -2121 948 -2119
rect 954 -2115 955 -2113
rect 954 -2121 955 -2119
rect 961 -2115 962 -2113
rect 961 -2121 962 -2119
rect 968 -2115 969 -2113
rect 968 -2121 969 -2119
rect 975 -2115 976 -2113
rect 975 -2121 976 -2119
rect 982 -2115 983 -2113
rect 982 -2121 983 -2119
rect 989 -2115 990 -2113
rect 989 -2121 990 -2119
rect 996 -2115 997 -2113
rect 996 -2121 997 -2119
rect 1003 -2115 1004 -2113
rect 1003 -2121 1004 -2119
rect 1010 -2115 1011 -2113
rect 1010 -2121 1011 -2119
rect 1017 -2115 1018 -2113
rect 1017 -2121 1018 -2119
rect 1024 -2115 1025 -2113
rect 1024 -2121 1025 -2119
rect 1031 -2115 1032 -2113
rect 1031 -2121 1032 -2119
rect 1038 -2115 1039 -2113
rect 1038 -2121 1039 -2119
rect 1045 -2115 1046 -2113
rect 1045 -2121 1046 -2119
rect 1052 -2115 1053 -2113
rect 1052 -2121 1053 -2119
rect 1059 -2115 1060 -2113
rect 1059 -2121 1060 -2119
rect 1066 -2115 1067 -2113
rect 1066 -2121 1067 -2119
rect 1073 -2115 1074 -2113
rect 1073 -2121 1074 -2119
rect 1080 -2115 1081 -2113
rect 1080 -2121 1081 -2119
rect 1087 -2115 1088 -2113
rect 1087 -2121 1088 -2119
rect 1094 -2115 1095 -2113
rect 1094 -2121 1095 -2119
rect 1101 -2115 1102 -2113
rect 1101 -2121 1102 -2119
rect 1108 -2115 1109 -2113
rect 1108 -2121 1109 -2119
rect 1115 -2115 1116 -2113
rect 1115 -2121 1116 -2119
rect 1122 -2115 1123 -2113
rect 1122 -2121 1123 -2119
rect 2 -2210 3 -2208
rect 2 -2216 3 -2214
rect 9 -2210 10 -2208
rect 9 -2216 10 -2214
rect 16 -2210 17 -2208
rect 16 -2216 17 -2214
rect 23 -2210 24 -2208
rect 23 -2216 24 -2214
rect 30 -2216 31 -2214
rect 33 -2216 34 -2214
rect 40 -2210 41 -2208
rect 37 -2216 38 -2214
rect 44 -2210 45 -2208
rect 44 -2216 45 -2214
rect 51 -2210 52 -2208
rect 51 -2216 52 -2214
rect 58 -2210 59 -2208
rect 58 -2216 59 -2214
rect 65 -2210 66 -2208
rect 65 -2216 66 -2214
rect 72 -2210 73 -2208
rect 75 -2210 76 -2208
rect 79 -2210 80 -2208
rect 79 -2216 80 -2214
rect 86 -2210 87 -2208
rect 86 -2216 87 -2214
rect 93 -2210 94 -2208
rect 93 -2216 94 -2214
rect 100 -2210 101 -2208
rect 100 -2216 101 -2214
rect 107 -2210 108 -2208
rect 107 -2216 108 -2214
rect 114 -2210 115 -2208
rect 114 -2216 115 -2214
rect 121 -2210 122 -2208
rect 124 -2210 125 -2208
rect 121 -2216 122 -2214
rect 128 -2210 129 -2208
rect 128 -2216 129 -2214
rect 135 -2210 136 -2208
rect 135 -2216 136 -2214
rect 142 -2210 143 -2208
rect 142 -2216 143 -2214
rect 149 -2210 150 -2208
rect 149 -2216 150 -2214
rect 156 -2210 157 -2208
rect 156 -2216 157 -2214
rect 166 -2210 167 -2208
rect 163 -2216 164 -2214
rect 166 -2216 167 -2214
rect 173 -2210 174 -2208
rect 173 -2216 174 -2214
rect 177 -2210 178 -2208
rect 187 -2216 188 -2214
rect 191 -2210 192 -2208
rect 194 -2216 195 -2214
rect 198 -2210 199 -2208
rect 198 -2216 199 -2214
rect 205 -2210 206 -2208
rect 205 -2216 206 -2214
rect 208 -2216 209 -2214
rect 212 -2210 213 -2208
rect 212 -2216 213 -2214
rect 219 -2210 220 -2208
rect 219 -2216 220 -2214
rect 226 -2210 227 -2208
rect 226 -2216 227 -2214
rect 233 -2210 234 -2208
rect 233 -2216 234 -2214
rect 240 -2210 241 -2208
rect 240 -2216 241 -2214
rect 247 -2210 248 -2208
rect 247 -2216 248 -2214
rect 254 -2210 255 -2208
rect 254 -2216 255 -2214
rect 261 -2210 262 -2208
rect 261 -2216 262 -2214
rect 268 -2210 269 -2208
rect 268 -2216 269 -2214
rect 275 -2210 276 -2208
rect 275 -2216 276 -2214
rect 282 -2210 283 -2208
rect 282 -2216 283 -2214
rect 289 -2210 290 -2208
rect 289 -2216 290 -2214
rect 296 -2210 297 -2208
rect 296 -2216 297 -2214
rect 303 -2210 304 -2208
rect 303 -2216 304 -2214
rect 310 -2210 311 -2208
rect 310 -2216 311 -2214
rect 320 -2210 321 -2208
rect 317 -2216 318 -2214
rect 324 -2210 325 -2208
rect 324 -2216 325 -2214
rect 331 -2210 332 -2208
rect 331 -2216 332 -2214
rect 338 -2210 339 -2208
rect 341 -2210 342 -2208
rect 338 -2216 339 -2214
rect 341 -2216 342 -2214
rect 345 -2210 346 -2208
rect 345 -2216 346 -2214
rect 355 -2210 356 -2208
rect 352 -2216 353 -2214
rect 355 -2216 356 -2214
rect 359 -2210 360 -2208
rect 359 -2216 360 -2214
rect 366 -2210 367 -2208
rect 366 -2216 367 -2214
rect 376 -2210 377 -2208
rect 380 -2210 381 -2208
rect 380 -2216 381 -2214
rect 387 -2210 388 -2208
rect 387 -2216 388 -2214
rect 397 -2210 398 -2208
rect 394 -2216 395 -2214
rect 397 -2216 398 -2214
rect 401 -2210 402 -2208
rect 401 -2216 402 -2214
rect 408 -2210 409 -2208
rect 408 -2216 409 -2214
rect 415 -2210 416 -2208
rect 415 -2216 416 -2214
rect 422 -2210 423 -2208
rect 422 -2216 423 -2214
rect 429 -2210 430 -2208
rect 432 -2210 433 -2208
rect 429 -2216 430 -2214
rect 436 -2210 437 -2208
rect 439 -2210 440 -2208
rect 439 -2216 440 -2214
rect 443 -2210 444 -2208
rect 443 -2216 444 -2214
rect 450 -2210 451 -2208
rect 450 -2216 451 -2214
rect 457 -2210 458 -2208
rect 457 -2216 458 -2214
rect 464 -2210 465 -2208
rect 464 -2216 465 -2214
rect 471 -2210 472 -2208
rect 471 -2216 472 -2214
rect 478 -2210 479 -2208
rect 478 -2216 479 -2214
rect 485 -2210 486 -2208
rect 485 -2216 486 -2214
rect 492 -2210 493 -2208
rect 492 -2216 493 -2214
rect 499 -2210 500 -2208
rect 502 -2210 503 -2208
rect 502 -2216 503 -2214
rect 509 -2210 510 -2208
rect 509 -2216 510 -2214
rect 513 -2210 514 -2208
rect 513 -2216 514 -2214
rect 520 -2210 521 -2208
rect 523 -2210 524 -2208
rect 523 -2216 524 -2214
rect 527 -2210 528 -2208
rect 527 -2216 528 -2214
rect 534 -2210 535 -2208
rect 534 -2216 535 -2214
rect 541 -2210 542 -2208
rect 541 -2216 542 -2214
rect 548 -2210 549 -2208
rect 548 -2216 549 -2214
rect 555 -2210 556 -2208
rect 555 -2216 556 -2214
rect 565 -2210 566 -2208
rect 565 -2216 566 -2214
rect 572 -2210 573 -2208
rect 572 -2216 573 -2214
rect 576 -2210 577 -2208
rect 576 -2216 577 -2214
rect 583 -2210 584 -2208
rect 583 -2216 584 -2214
rect 590 -2210 591 -2208
rect 593 -2210 594 -2208
rect 590 -2216 591 -2214
rect 593 -2216 594 -2214
rect 597 -2210 598 -2208
rect 600 -2210 601 -2208
rect 604 -2210 605 -2208
rect 607 -2210 608 -2208
rect 604 -2216 605 -2214
rect 611 -2210 612 -2208
rect 611 -2216 612 -2214
rect 618 -2210 619 -2208
rect 618 -2216 619 -2214
rect 625 -2210 626 -2208
rect 625 -2216 626 -2214
rect 632 -2210 633 -2208
rect 632 -2216 633 -2214
rect 639 -2210 640 -2208
rect 639 -2216 640 -2214
rect 646 -2210 647 -2208
rect 646 -2216 647 -2214
rect 653 -2210 654 -2208
rect 653 -2216 654 -2214
rect 660 -2210 661 -2208
rect 660 -2216 661 -2214
rect 667 -2210 668 -2208
rect 670 -2210 671 -2208
rect 670 -2216 671 -2214
rect 674 -2210 675 -2208
rect 674 -2216 675 -2214
rect 684 -2210 685 -2208
rect 681 -2216 682 -2214
rect 684 -2216 685 -2214
rect 688 -2210 689 -2208
rect 691 -2216 692 -2214
rect 695 -2210 696 -2208
rect 698 -2210 699 -2208
rect 695 -2216 696 -2214
rect 698 -2216 699 -2214
rect 702 -2210 703 -2208
rect 702 -2216 703 -2214
rect 709 -2210 710 -2208
rect 709 -2216 710 -2214
rect 716 -2210 717 -2208
rect 716 -2216 717 -2214
rect 723 -2210 724 -2208
rect 726 -2210 727 -2208
rect 723 -2216 724 -2214
rect 726 -2216 727 -2214
rect 730 -2210 731 -2208
rect 730 -2216 731 -2214
rect 737 -2210 738 -2208
rect 737 -2216 738 -2214
rect 744 -2210 745 -2208
rect 744 -2216 745 -2214
rect 751 -2210 752 -2208
rect 751 -2216 752 -2214
rect 758 -2210 759 -2208
rect 758 -2216 759 -2214
rect 765 -2210 766 -2208
rect 765 -2216 766 -2214
rect 772 -2210 773 -2208
rect 772 -2216 773 -2214
rect 779 -2210 780 -2208
rect 779 -2216 780 -2214
rect 786 -2210 787 -2208
rect 786 -2216 787 -2214
rect 793 -2210 794 -2208
rect 793 -2216 794 -2214
rect 800 -2210 801 -2208
rect 800 -2216 801 -2214
rect 807 -2210 808 -2208
rect 807 -2216 808 -2214
rect 814 -2210 815 -2208
rect 814 -2216 815 -2214
rect 821 -2210 822 -2208
rect 821 -2216 822 -2214
rect 828 -2210 829 -2208
rect 828 -2216 829 -2214
rect 835 -2210 836 -2208
rect 835 -2216 836 -2214
rect 842 -2210 843 -2208
rect 842 -2216 843 -2214
rect 849 -2210 850 -2208
rect 849 -2216 850 -2214
rect 856 -2210 857 -2208
rect 856 -2216 857 -2214
rect 863 -2210 864 -2208
rect 863 -2216 864 -2214
rect 873 -2210 874 -2208
rect 877 -2210 878 -2208
rect 877 -2216 878 -2214
rect 884 -2210 885 -2208
rect 884 -2216 885 -2214
rect 891 -2210 892 -2208
rect 891 -2216 892 -2214
rect 898 -2210 899 -2208
rect 898 -2216 899 -2214
rect 905 -2210 906 -2208
rect 905 -2216 906 -2214
rect 912 -2210 913 -2208
rect 912 -2216 913 -2214
rect 919 -2210 920 -2208
rect 919 -2216 920 -2214
rect 926 -2210 927 -2208
rect 926 -2216 927 -2214
rect 933 -2210 934 -2208
rect 933 -2216 934 -2214
rect 940 -2210 941 -2208
rect 940 -2216 941 -2214
rect 947 -2210 948 -2208
rect 947 -2216 948 -2214
rect 954 -2210 955 -2208
rect 954 -2216 955 -2214
rect 961 -2210 962 -2208
rect 961 -2216 962 -2214
rect 968 -2210 969 -2208
rect 968 -2216 969 -2214
rect 975 -2210 976 -2208
rect 975 -2216 976 -2214
rect 982 -2210 983 -2208
rect 982 -2216 983 -2214
rect 989 -2210 990 -2208
rect 989 -2216 990 -2214
rect 996 -2210 997 -2208
rect 996 -2216 997 -2214
rect 1003 -2210 1004 -2208
rect 1003 -2216 1004 -2214
rect 1010 -2210 1011 -2208
rect 1010 -2216 1011 -2214
rect 1017 -2210 1018 -2208
rect 1017 -2216 1018 -2214
rect 1024 -2210 1025 -2208
rect 1024 -2216 1025 -2214
rect 1031 -2210 1032 -2208
rect 1031 -2216 1032 -2214
rect 1038 -2210 1039 -2208
rect 1038 -2216 1039 -2214
rect 1045 -2210 1046 -2208
rect 1045 -2216 1046 -2214
rect 1055 -2210 1056 -2208
rect 2 -2279 3 -2277
rect 2 -2285 3 -2283
rect 9 -2279 10 -2277
rect 9 -2285 10 -2283
rect 16 -2279 17 -2277
rect 16 -2285 17 -2283
rect 23 -2279 24 -2277
rect 23 -2285 24 -2283
rect 30 -2279 31 -2277
rect 30 -2285 31 -2283
rect 37 -2279 38 -2277
rect 37 -2285 38 -2283
rect 44 -2279 45 -2277
rect 44 -2285 45 -2283
rect 51 -2279 52 -2277
rect 51 -2285 52 -2283
rect 54 -2285 55 -2283
rect 58 -2279 59 -2277
rect 58 -2285 59 -2283
rect 61 -2285 62 -2283
rect 65 -2279 66 -2277
rect 65 -2285 66 -2283
rect 72 -2279 73 -2277
rect 72 -2285 73 -2283
rect 79 -2285 80 -2283
rect 82 -2285 83 -2283
rect 86 -2279 87 -2277
rect 86 -2285 87 -2283
rect 93 -2279 94 -2277
rect 93 -2285 94 -2283
rect 103 -2279 104 -2277
rect 100 -2285 101 -2283
rect 103 -2285 104 -2283
rect 107 -2279 108 -2277
rect 107 -2285 108 -2283
rect 110 -2285 111 -2283
rect 114 -2279 115 -2277
rect 114 -2285 115 -2283
rect 121 -2279 122 -2277
rect 121 -2285 122 -2283
rect 128 -2285 129 -2283
rect 131 -2285 132 -2283
rect 135 -2279 136 -2277
rect 135 -2285 136 -2283
rect 142 -2279 143 -2277
rect 142 -2285 143 -2283
rect 149 -2279 150 -2277
rect 149 -2285 150 -2283
rect 156 -2279 157 -2277
rect 156 -2285 157 -2283
rect 163 -2279 164 -2277
rect 163 -2285 164 -2283
rect 170 -2279 171 -2277
rect 170 -2285 171 -2283
rect 177 -2279 178 -2277
rect 177 -2285 178 -2283
rect 180 -2285 181 -2283
rect 184 -2279 185 -2277
rect 184 -2285 185 -2283
rect 191 -2279 192 -2277
rect 191 -2285 192 -2283
rect 198 -2279 199 -2277
rect 201 -2279 202 -2277
rect 198 -2285 199 -2283
rect 205 -2279 206 -2277
rect 205 -2285 206 -2283
rect 212 -2279 213 -2277
rect 215 -2279 216 -2277
rect 215 -2285 216 -2283
rect 219 -2279 220 -2277
rect 226 -2279 227 -2277
rect 226 -2285 227 -2283
rect 233 -2279 234 -2277
rect 233 -2285 234 -2283
rect 240 -2279 241 -2277
rect 240 -2285 241 -2283
rect 247 -2279 248 -2277
rect 247 -2285 248 -2283
rect 254 -2279 255 -2277
rect 254 -2285 255 -2283
rect 261 -2279 262 -2277
rect 261 -2285 262 -2283
rect 268 -2279 269 -2277
rect 268 -2285 269 -2283
rect 275 -2279 276 -2277
rect 275 -2285 276 -2283
rect 282 -2279 283 -2277
rect 282 -2285 283 -2283
rect 292 -2279 293 -2277
rect 289 -2285 290 -2283
rect 292 -2285 293 -2283
rect 296 -2279 297 -2277
rect 296 -2285 297 -2283
rect 303 -2279 304 -2277
rect 303 -2285 304 -2283
rect 310 -2279 311 -2277
rect 310 -2285 311 -2283
rect 317 -2279 318 -2277
rect 317 -2285 318 -2283
rect 324 -2279 325 -2277
rect 327 -2279 328 -2277
rect 331 -2279 332 -2277
rect 331 -2285 332 -2283
rect 338 -2279 339 -2277
rect 338 -2285 339 -2283
rect 348 -2279 349 -2277
rect 348 -2285 349 -2283
rect 352 -2279 353 -2277
rect 355 -2279 356 -2277
rect 352 -2285 353 -2283
rect 355 -2285 356 -2283
rect 359 -2279 360 -2277
rect 359 -2285 360 -2283
rect 369 -2279 370 -2277
rect 366 -2285 367 -2283
rect 373 -2279 374 -2277
rect 373 -2285 374 -2283
rect 380 -2279 381 -2277
rect 383 -2279 384 -2277
rect 380 -2285 381 -2283
rect 383 -2285 384 -2283
rect 387 -2279 388 -2277
rect 387 -2285 388 -2283
rect 394 -2279 395 -2277
rect 394 -2285 395 -2283
rect 401 -2279 402 -2277
rect 401 -2285 402 -2283
rect 408 -2279 409 -2277
rect 408 -2285 409 -2283
rect 415 -2279 416 -2277
rect 415 -2285 416 -2283
rect 422 -2279 423 -2277
rect 422 -2285 423 -2283
rect 429 -2279 430 -2277
rect 429 -2285 430 -2283
rect 436 -2279 437 -2277
rect 436 -2285 437 -2283
rect 443 -2279 444 -2277
rect 443 -2285 444 -2283
rect 450 -2279 451 -2277
rect 450 -2285 451 -2283
rect 457 -2279 458 -2277
rect 457 -2285 458 -2283
rect 464 -2279 465 -2277
rect 467 -2279 468 -2277
rect 464 -2285 465 -2283
rect 467 -2285 468 -2283
rect 471 -2279 472 -2277
rect 471 -2285 472 -2283
rect 478 -2279 479 -2277
rect 481 -2279 482 -2277
rect 481 -2285 482 -2283
rect 485 -2279 486 -2277
rect 488 -2279 489 -2277
rect 485 -2285 486 -2283
rect 488 -2285 489 -2283
rect 492 -2279 493 -2277
rect 492 -2285 493 -2283
rect 499 -2279 500 -2277
rect 502 -2279 503 -2277
rect 502 -2285 503 -2283
rect 506 -2279 507 -2277
rect 506 -2285 507 -2283
rect 513 -2279 514 -2277
rect 513 -2285 514 -2283
rect 520 -2279 521 -2277
rect 520 -2285 521 -2283
rect 527 -2279 528 -2277
rect 527 -2285 528 -2283
rect 534 -2279 535 -2277
rect 534 -2285 535 -2283
rect 541 -2279 542 -2277
rect 544 -2279 545 -2277
rect 541 -2285 542 -2283
rect 544 -2285 545 -2283
rect 548 -2279 549 -2277
rect 548 -2285 549 -2283
rect 555 -2279 556 -2277
rect 555 -2285 556 -2283
rect 562 -2279 563 -2277
rect 562 -2285 563 -2283
rect 569 -2279 570 -2277
rect 569 -2285 570 -2283
rect 576 -2279 577 -2277
rect 579 -2279 580 -2277
rect 576 -2285 577 -2283
rect 579 -2285 580 -2283
rect 583 -2279 584 -2277
rect 583 -2285 584 -2283
rect 590 -2279 591 -2277
rect 590 -2285 591 -2283
rect 597 -2279 598 -2277
rect 597 -2285 598 -2283
rect 604 -2279 605 -2277
rect 604 -2285 605 -2283
rect 611 -2279 612 -2277
rect 611 -2285 612 -2283
rect 618 -2279 619 -2277
rect 618 -2285 619 -2283
rect 625 -2279 626 -2277
rect 625 -2285 626 -2283
rect 632 -2279 633 -2277
rect 632 -2285 633 -2283
rect 639 -2279 640 -2277
rect 639 -2285 640 -2283
rect 646 -2279 647 -2277
rect 646 -2285 647 -2283
rect 653 -2279 654 -2277
rect 653 -2285 654 -2283
rect 660 -2279 661 -2277
rect 660 -2285 661 -2283
rect 667 -2279 668 -2277
rect 667 -2285 668 -2283
rect 674 -2279 675 -2277
rect 674 -2285 675 -2283
rect 681 -2279 682 -2277
rect 684 -2279 685 -2277
rect 681 -2285 682 -2283
rect 684 -2285 685 -2283
rect 688 -2279 689 -2277
rect 688 -2285 689 -2283
rect 695 -2279 696 -2277
rect 695 -2285 696 -2283
rect 702 -2279 703 -2277
rect 702 -2285 703 -2283
rect 709 -2279 710 -2277
rect 709 -2285 710 -2283
rect 716 -2279 717 -2277
rect 716 -2285 717 -2283
rect 723 -2279 724 -2277
rect 723 -2285 724 -2283
rect 730 -2279 731 -2277
rect 730 -2285 731 -2283
rect 737 -2279 738 -2277
rect 737 -2285 738 -2283
rect 744 -2279 745 -2277
rect 744 -2285 745 -2283
rect 751 -2279 752 -2277
rect 751 -2285 752 -2283
rect 758 -2279 759 -2277
rect 758 -2285 759 -2283
rect 768 -2279 769 -2277
rect 768 -2285 769 -2283
rect 772 -2279 773 -2277
rect 772 -2285 773 -2283
rect 779 -2279 780 -2277
rect 779 -2285 780 -2283
rect 786 -2279 787 -2277
rect 786 -2285 787 -2283
rect 793 -2279 794 -2277
rect 793 -2285 794 -2283
rect 800 -2279 801 -2277
rect 800 -2285 801 -2283
rect 807 -2279 808 -2277
rect 807 -2285 808 -2283
rect 814 -2279 815 -2277
rect 814 -2285 815 -2283
rect 821 -2279 822 -2277
rect 821 -2285 822 -2283
rect 828 -2279 829 -2277
rect 828 -2285 829 -2283
rect 835 -2279 836 -2277
rect 835 -2285 836 -2283
rect 842 -2279 843 -2277
rect 842 -2285 843 -2283
rect 849 -2279 850 -2277
rect 849 -2285 850 -2283
rect 856 -2279 857 -2277
rect 856 -2285 857 -2283
rect 863 -2279 864 -2277
rect 863 -2285 864 -2283
rect 870 -2279 871 -2277
rect 870 -2285 871 -2283
rect 877 -2279 878 -2277
rect 877 -2285 878 -2283
rect 884 -2279 885 -2277
rect 884 -2285 885 -2283
rect 891 -2279 892 -2277
rect 891 -2285 892 -2283
rect 898 -2279 899 -2277
rect 898 -2285 899 -2283
rect 901 -2285 902 -2283
rect 905 -2285 906 -2283
rect 908 -2285 909 -2283
rect 912 -2279 913 -2277
rect 912 -2285 913 -2283
rect 922 -2279 923 -2277
rect 922 -2285 923 -2283
rect 929 -2279 930 -2277
rect 926 -2285 927 -2283
rect 933 -2279 934 -2277
rect 933 -2285 934 -2283
rect 940 -2279 941 -2277
rect 940 -2285 941 -2283
rect 947 -2279 948 -2277
rect 947 -2285 948 -2283
rect 954 -2279 955 -2277
rect 954 -2285 955 -2283
rect 961 -2279 962 -2277
rect 961 -2285 962 -2283
rect 968 -2279 969 -2277
rect 975 -2279 976 -2277
rect 975 -2285 976 -2283
rect 2 -2366 3 -2364
rect 2 -2372 3 -2370
rect 12 -2366 13 -2364
rect 16 -2366 17 -2364
rect 16 -2372 17 -2370
rect 23 -2366 24 -2364
rect 23 -2372 24 -2370
rect 30 -2366 31 -2364
rect 30 -2372 31 -2370
rect 37 -2366 38 -2364
rect 37 -2372 38 -2370
rect 44 -2366 45 -2364
rect 47 -2366 48 -2364
rect 44 -2372 45 -2370
rect 51 -2366 52 -2364
rect 54 -2366 55 -2364
rect 51 -2372 52 -2370
rect 58 -2366 59 -2364
rect 58 -2372 59 -2370
rect 65 -2366 66 -2364
rect 65 -2372 66 -2370
rect 72 -2366 73 -2364
rect 72 -2372 73 -2370
rect 79 -2366 80 -2364
rect 79 -2372 80 -2370
rect 86 -2366 87 -2364
rect 86 -2372 87 -2370
rect 93 -2366 94 -2364
rect 93 -2372 94 -2370
rect 100 -2366 101 -2364
rect 100 -2372 101 -2370
rect 107 -2366 108 -2364
rect 110 -2366 111 -2364
rect 107 -2372 108 -2370
rect 114 -2366 115 -2364
rect 114 -2372 115 -2370
rect 121 -2366 122 -2364
rect 121 -2372 122 -2370
rect 128 -2366 129 -2364
rect 128 -2372 129 -2370
rect 135 -2366 136 -2364
rect 135 -2372 136 -2370
rect 142 -2366 143 -2364
rect 142 -2372 143 -2370
rect 149 -2366 150 -2364
rect 149 -2372 150 -2370
rect 156 -2366 157 -2364
rect 159 -2366 160 -2364
rect 156 -2372 157 -2370
rect 163 -2366 164 -2364
rect 163 -2372 164 -2370
rect 170 -2366 171 -2364
rect 170 -2372 171 -2370
rect 177 -2366 178 -2364
rect 177 -2372 178 -2370
rect 184 -2366 185 -2364
rect 184 -2372 185 -2370
rect 191 -2366 192 -2364
rect 191 -2372 192 -2370
rect 198 -2366 199 -2364
rect 198 -2372 199 -2370
rect 205 -2366 206 -2364
rect 205 -2372 206 -2370
rect 212 -2366 213 -2364
rect 212 -2372 213 -2370
rect 219 -2372 220 -2370
rect 222 -2372 223 -2370
rect 229 -2366 230 -2364
rect 226 -2372 227 -2370
rect 233 -2366 234 -2364
rect 233 -2372 234 -2370
rect 240 -2366 241 -2364
rect 240 -2372 241 -2370
rect 247 -2366 248 -2364
rect 247 -2372 248 -2370
rect 254 -2366 255 -2364
rect 254 -2372 255 -2370
rect 261 -2366 262 -2364
rect 261 -2372 262 -2370
rect 268 -2366 269 -2364
rect 271 -2372 272 -2370
rect 275 -2366 276 -2364
rect 275 -2372 276 -2370
rect 282 -2366 283 -2364
rect 282 -2372 283 -2370
rect 289 -2366 290 -2364
rect 289 -2372 290 -2370
rect 296 -2366 297 -2364
rect 296 -2372 297 -2370
rect 303 -2366 304 -2364
rect 303 -2372 304 -2370
rect 310 -2366 311 -2364
rect 313 -2366 314 -2364
rect 310 -2372 311 -2370
rect 313 -2372 314 -2370
rect 317 -2366 318 -2364
rect 317 -2372 318 -2370
rect 324 -2366 325 -2364
rect 324 -2372 325 -2370
rect 334 -2366 335 -2364
rect 331 -2372 332 -2370
rect 334 -2372 335 -2370
rect 338 -2366 339 -2364
rect 341 -2366 342 -2364
rect 341 -2372 342 -2370
rect 345 -2366 346 -2364
rect 345 -2372 346 -2370
rect 355 -2366 356 -2364
rect 355 -2372 356 -2370
rect 359 -2366 360 -2364
rect 362 -2366 363 -2364
rect 366 -2366 367 -2364
rect 366 -2372 367 -2370
rect 373 -2366 374 -2364
rect 376 -2366 377 -2364
rect 380 -2366 381 -2364
rect 380 -2372 381 -2370
rect 387 -2366 388 -2364
rect 387 -2372 388 -2370
rect 394 -2366 395 -2364
rect 397 -2366 398 -2364
rect 401 -2366 402 -2364
rect 401 -2372 402 -2370
rect 404 -2372 405 -2370
rect 408 -2366 409 -2364
rect 408 -2372 409 -2370
rect 415 -2366 416 -2364
rect 415 -2372 416 -2370
rect 418 -2372 419 -2370
rect 422 -2366 423 -2364
rect 422 -2372 423 -2370
rect 429 -2366 430 -2364
rect 429 -2372 430 -2370
rect 436 -2366 437 -2364
rect 436 -2372 437 -2370
rect 443 -2366 444 -2364
rect 443 -2372 444 -2370
rect 450 -2366 451 -2364
rect 450 -2372 451 -2370
rect 457 -2372 458 -2370
rect 464 -2366 465 -2364
rect 467 -2366 468 -2364
rect 464 -2372 465 -2370
rect 471 -2366 472 -2364
rect 471 -2372 472 -2370
rect 478 -2366 479 -2364
rect 485 -2366 486 -2364
rect 485 -2372 486 -2370
rect 492 -2366 493 -2364
rect 492 -2372 493 -2370
rect 499 -2366 500 -2364
rect 499 -2372 500 -2370
rect 506 -2366 507 -2364
rect 506 -2372 507 -2370
rect 513 -2366 514 -2364
rect 513 -2372 514 -2370
rect 523 -2366 524 -2364
rect 523 -2372 524 -2370
rect 527 -2366 528 -2364
rect 527 -2372 528 -2370
rect 537 -2366 538 -2364
rect 534 -2372 535 -2370
rect 541 -2366 542 -2364
rect 541 -2372 542 -2370
rect 548 -2366 549 -2364
rect 548 -2372 549 -2370
rect 555 -2366 556 -2364
rect 558 -2372 559 -2370
rect 562 -2366 563 -2364
rect 565 -2366 566 -2364
rect 565 -2372 566 -2370
rect 569 -2366 570 -2364
rect 569 -2372 570 -2370
rect 576 -2366 577 -2364
rect 576 -2372 577 -2370
rect 583 -2366 584 -2364
rect 586 -2366 587 -2364
rect 590 -2366 591 -2364
rect 590 -2372 591 -2370
rect 597 -2366 598 -2364
rect 597 -2372 598 -2370
rect 604 -2366 605 -2364
rect 604 -2372 605 -2370
rect 611 -2366 612 -2364
rect 611 -2372 612 -2370
rect 618 -2366 619 -2364
rect 618 -2372 619 -2370
rect 625 -2366 626 -2364
rect 625 -2372 626 -2370
rect 632 -2366 633 -2364
rect 632 -2372 633 -2370
rect 639 -2366 640 -2364
rect 642 -2366 643 -2364
rect 639 -2372 640 -2370
rect 646 -2366 647 -2364
rect 646 -2372 647 -2370
rect 653 -2366 654 -2364
rect 653 -2372 654 -2370
rect 660 -2366 661 -2364
rect 660 -2372 661 -2370
rect 667 -2366 668 -2364
rect 667 -2372 668 -2370
rect 674 -2366 675 -2364
rect 674 -2372 675 -2370
rect 681 -2366 682 -2364
rect 681 -2372 682 -2370
rect 688 -2366 689 -2364
rect 688 -2372 689 -2370
rect 695 -2366 696 -2364
rect 695 -2372 696 -2370
rect 702 -2366 703 -2364
rect 705 -2366 706 -2364
rect 709 -2366 710 -2364
rect 709 -2372 710 -2370
rect 716 -2366 717 -2364
rect 716 -2372 717 -2370
rect 723 -2366 724 -2364
rect 723 -2372 724 -2370
rect 730 -2366 731 -2364
rect 730 -2372 731 -2370
rect 737 -2366 738 -2364
rect 737 -2372 738 -2370
rect 744 -2366 745 -2364
rect 744 -2372 745 -2370
rect 751 -2366 752 -2364
rect 751 -2372 752 -2370
rect 758 -2366 759 -2364
rect 758 -2372 759 -2370
rect 765 -2366 766 -2364
rect 765 -2372 766 -2370
rect 772 -2366 773 -2364
rect 772 -2372 773 -2370
rect 779 -2366 780 -2364
rect 779 -2372 780 -2370
rect 786 -2366 787 -2364
rect 786 -2372 787 -2370
rect 793 -2366 794 -2364
rect 793 -2372 794 -2370
rect 800 -2366 801 -2364
rect 807 -2366 808 -2364
rect 807 -2372 808 -2370
rect 814 -2366 815 -2364
rect 814 -2372 815 -2370
rect 821 -2366 822 -2364
rect 821 -2372 822 -2370
rect 828 -2366 829 -2364
rect 828 -2372 829 -2370
rect 835 -2366 836 -2364
rect 835 -2372 836 -2370
rect 842 -2366 843 -2364
rect 842 -2372 843 -2370
rect 849 -2366 850 -2364
rect 849 -2372 850 -2370
rect 856 -2366 857 -2364
rect 856 -2372 857 -2370
rect 863 -2366 864 -2364
rect 863 -2372 864 -2370
rect 870 -2366 871 -2364
rect 877 -2366 878 -2364
rect 877 -2372 878 -2370
rect 884 -2366 885 -2364
rect 884 -2372 885 -2370
rect 891 -2366 892 -2364
rect 891 -2372 892 -2370
rect 929 -2366 930 -2364
rect 926 -2372 927 -2370
rect 947 -2366 948 -2364
rect 947 -2372 948 -2370
rect 30 -2431 31 -2429
rect 58 -2431 59 -2429
rect 61 -2431 62 -2429
rect 65 -2431 66 -2429
rect 65 -2437 66 -2435
rect 72 -2431 73 -2429
rect 79 -2431 80 -2429
rect 79 -2437 80 -2435
rect 86 -2431 87 -2429
rect 86 -2437 87 -2435
rect 93 -2431 94 -2429
rect 93 -2437 94 -2435
rect 100 -2431 101 -2429
rect 100 -2437 101 -2435
rect 107 -2431 108 -2429
rect 107 -2437 108 -2435
rect 114 -2431 115 -2429
rect 114 -2437 115 -2435
rect 121 -2431 122 -2429
rect 121 -2437 122 -2435
rect 128 -2431 129 -2429
rect 128 -2437 129 -2435
rect 138 -2431 139 -2429
rect 142 -2431 143 -2429
rect 142 -2437 143 -2435
rect 149 -2431 150 -2429
rect 152 -2431 153 -2429
rect 149 -2437 150 -2435
rect 152 -2437 153 -2435
rect 156 -2431 157 -2429
rect 156 -2437 157 -2435
rect 159 -2437 160 -2435
rect 163 -2431 164 -2429
rect 163 -2437 164 -2435
rect 170 -2431 171 -2429
rect 170 -2437 171 -2435
rect 177 -2431 178 -2429
rect 177 -2437 178 -2435
rect 184 -2431 185 -2429
rect 184 -2437 185 -2435
rect 191 -2431 192 -2429
rect 191 -2437 192 -2435
rect 198 -2431 199 -2429
rect 198 -2437 199 -2435
rect 208 -2431 209 -2429
rect 208 -2437 209 -2435
rect 215 -2431 216 -2429
rect 212 -2437 213 -2435
rect 215 -2437 216 -2435
rect 219 -2431 220 -2429
rect 222 -2431 223 -2429
rect 219 -2437 220 -2435
rect 222 -2437 223 -2435
rect 226 -2431 227 -2429
rect 226 -2437 227 -2435
rect 233 -2431 234 -2429
rect 233 -2437 234 -2435
rect 240 -2431 241 -2429
rect 240 -2437 241 -2435
rect 247 -2431 248 -2429
rect 247 -2437 248 -2435
rect 254 -2431 255 -2429
rect 254 -2437 255 -2435
rect 261 -2431 262 -2429
rect 261 -2437 262 -2435
rect 268 -2431 269 -2429
rect 268 -2437 269 -2435
rect 275 -2431 276 -2429
rect 275 -2437 276 -2435
rect 282 -2431 283 -2429
rect 282 -2437 283 -2435
rect 289 -2431 290 -2429
rect 289 -2437 290 -2435
rect 296 -2431 297 -2429
rect 296 -2437 297 -2435
rect 303 -2431 304 -2429
rect 303 -2437 304 -2435
rect 310 -2431 311 -2429
rect 310 -2437 311 -2435
rect 317 -2431 318 -2429
rect 317 -2437 318 -2435
rect 324 -2431 325 -2429
rect 324 -2437 325 -2435
rect 331 -2431 332 -2429
rect 334 -2431 335 -2429
rect 331 -2437 332 -2435
rect 334 -2437 335 -2435
rect 338 -2431 339 -2429
rect 338 -2437 339 -2435
rect 345 -2431 346 -2429
rect 345 -2437 346 -2435
rect 352 -2431 353 -2429
rect 352 -2437 353 -2435
rect 359 -2431 360 -2429
rect 359 -2437 360 -2435
rect 366 -2431 367 -2429
rect 366 -2437 367 -2435
rect 373 -2431 374 -2429
rect 376 -2431 377 -2429
rect 380 -2431 381 -2429
rect 380 -2437 381 -2435
rect 387 -2431 388 -2429
rect 387 -2437 388 -2435
rect 394 -2431 395 -2429
rect 397 -2431 398 -2429
rect 394 -2437 395 -2435
rect 397 -2437 398 -2435
rect 401 -2431 402 -2429
rect 401 -2437 402 -2435
rect 408 -2431 409 -2429
rect 411 -2431 412 -2429
rect 408 -2437 409 -2435
rect 415 -2431 416 -2429
rect 415 -2437 416 -2435
rect 422 -2431 423 -2429
rect 422 -2437 423 -2435
rect 429 -2431 430 -2429
rect 432 -2437 433 -2435
rect 436 -2431 437 -2429
rect 436 -2437 437 -2435
rect 443 -2431 444 -2429
rect 443 -2437 444 -2435
rect 450 -2431 451 -2429
rect 450 -2437 451 -2435
rect 457 -2431 458 -2429
rect 460 -2431 461 -2429
rect 460 -2437 461 -2435
rect 464 -2431 465 -2429
rect 464 -2437 465 -2435
rect 467 -2437 468 -2435
rect 471 -2431 472 -2429
rect 471 -2437 472 -2435
rect 474 -2437 475 -2435
rect 481 -2431 482 -2429
rect 478 -2437 479 -2435
rect 481 -2437 482 -2435
rect 488 -2431 489 -2429
rect 485 -2437 486 -2435
rect 488 -2437 489 -2435
rect 492 -2431 493 -2429
rect 492 -2437 493 -2435
rect 499 -2431 500 -2429
rect 499 -2437 500 -2435
rect 506 -2431 507 -2429
rect 506 -2437 507 -2435
rect 513 -2431 514 -2429
rect 513 -2437 514 -2435
rect 520 -2431 521 -2429
rect 520 -2437 521 -2435
rect 527 -2431 528 -2429
rect 527 -2437 528 -2435
rect 534 -2431 535 -2429
rect 534 -2437 535 -2435
rect 544 -2431 545 -2429
rect 548 -2431 549 -2429
rect 551 -2431 552 -2429
rect 551 -2437 552 -2435
rect 555 -2431 556 -2429
rect 555 -2437 556 -2435
rect 562 -2431 563 -2429
rect 562 -2437 563 -2435
rect 569 -2431 570 -2429
rect 569 -2437 570 -2435
rect 576 -2437 577 -2435
rect 579 -2437 580 -2435
rect 583 -2431 584 -2429
rect 583 -2437 584 -2435
rect 590 -2431 591 -2429
rect 590 -2437 591 -2435
rect 597 -2431 598 -2429
rect 597 -2437 598 -2435
rect 604 -2431 605 -2429
rect 604 -2437 605 -2435
rect 611 -2431 612 -2429
rect 611 -2437 612 -2435
rect 618 -2431 619 -2429
rect 618 -2437 619 -2435
rect 628 -2431 629 -2429
rect 625 -2437 626 -2435
rect 632 -2431 633 -2429
rect 632 -2437 633 -2435
rect 639 -2431 640 -2429
rect 639 -2437 640 -2435
rect 646 -2431 647 -2429
rect 646 -2437 647 -2435
rect 653 -2431 654 -2429
rect 653 -2437 654 -2435
rect 660 -2431 661 -2429
rect 660 -2437 661 -2435
rect 667 -2431 668 -2429
rect 667 -2437 668 -2435
rect 674 -2431 675 -2429
rect 674 -2437 675 -2435
rect 681 -2431 682 -2429
rect 681 -2437 682 -2435
rect 702 -2431 703 -2429
rect 702 -2437 703 -2435
rect 709 -2431 710 -2429
rect 709 -2437 710 -2435
rect 716 -2431 717 -2429
rect 716 -2437 717 -2435
rect 723 -2431 724 -2429
rect 726 -2431 727 -2429
rect 723 -2437 724 -2435
rect 726 -2437 727 -2435
rect 730 -2437 731 -2435
rect 733 -2437 734 -2435
rect 737 -2431 738 -2429
rect 737 -2437 738 -2435
rect 744 -2431 745 -2429
rect 744 -2437 745 -2435
rect 754 -2431 755 -2429
rect 754 -2437 755 -2435
rect 761 -2431 762 -2429
rect 758 -2437 759 -2435
rect 761 -2437 762 -2435
rect 765 -2431 766 -2429
rect 765 -2437 766 -2435
rect 772 -2431 773 -2429
rect 772 -2437 773 -2435
rect 779 -2437 780 -2435
rect 807 -2431 808 -2429
rect 807 -2437 808 -2435
rect 828 -2431 829 -2429
rect 828 -2437 829 -2435
rect 884 -2431 885 -2429
rect 884 -2437 885 -2435
rect 891 -2431 892 -2429
rect 891 -2437 892 -2435
rect 926 -2431 927 -2429
rect 926 -2437 927 -2435
rect 940 -2431 941 -2429
rect 940 -2437 941 -2435
rect 5 -2478 6 -2476
rect 65 -2478 66 -2476
rect 72 -2472 73 -2470
rect 72 -2478 73 -2476
rect 100 -2472 101 -2470
rect 100 -2478 101 -2476
rect 107 -2472 108 -2470
rect 107 -2478 108 -2476
rect 114 -2472 115 -2470
rect 117 -2472 118 -2470
rect 114 -2478 115 -2476
rect 121 -2472 122 -2470
rect 121 -2478 122 -2476
rect 131 -2472 132 -2470
rect 131 -2478 132 -2476
rect 135 -2472 136 -2470
rect 135 -2478 136 -2476
rect 163 -2472 164 -2470
rect 163 -2478 164 -2476
rect 170 -2472 171 -2470
rect 170 -2478 171 -2476
rect 177 -2472 178 -2470
rect 177 -2478 178 -2476
rect 184 -2472 185 -2470
rect 187 -2478 188 -2476
rect 191 -2472 192 -2470
rect 191 -2478 192 -2476
rect 198 -2472 199 -2470
rect 198 -2478 199 -2476
rect 205 -2472 206 -2470
rect 205 -2478 206 -2476
rect 219 -2472 220 -2470
rect 219 -2478 220 -2476
rect 226 -2472 227 -2470
rect 226 -2478 227 -2476
rect 233 -2472 234 -2470
rect 233 -2478 234 -2476
rect 236 -2478 237 -2476
rect 240 -2472 241 -2470
rect 247 -2472 248 -2470
rect 247 -2478 248 -2476
rect 257 -2472 258 -2470
rect 264 -2472 265 -2470
rect 261 -2478 262 -2476
rect 268 -2472 269 -2470
rect 268 -2478 269 -2476
rect 275 -2472 276 -2470
rect 275 -2478 276 -2476
rect 282 -2472 283 -2470
rect 282 -2478 283 -2476
rect 289 -2472 290 -2470
rect 289 -2478 290 -2476
rect 299 -2472 300 -2470
rect 296 -2478 297 -2476
rect 303 -2472 304 -2470
rect 303 -2478 304 -2476
rect 310 -2472 311 -2470
rect 310 -2478 311 -2476
rect 317 -2472 318 -2470
rect 317 -2478 318 -2476
rect 324 -2478 325 -2476
rect 331 -2472 332 -2470
rect 331 -2478 332 -2476
rect 338 -2472 339 -2470
rect 338 -2478 339 -2476
rect 345 -2472 346 -2470
rect 348 -2472 349 -2470
rect 352 -2472 353 -2470
rect 352 -2478 353 -2476
rect 359 -2472 360 -2470
rect 359 -2478 360 -2476
rect 369 -2472 370 -2470
rect 366 -2478 367 -2476
rect 373 -2472 374 -2470
rect 373 -2478 374 -2476
rect 376 -2478 377 -2476
rect 380 -2472 381 -2470
rect 380 -2478 381 -2476
rect 387 -2472 388 -2470
rect 390 -2472 391 -2470
rect 394 -2472 395 -2470
rect 394 -2478 395 -2476
rect 401 -2472 402 -2470
rect 401 -2478 402 -2476
rect 408 -2472 409 -2470
rect 408 -2478 409 -2476
rect 415 -2472 416 -2470
rect 415 -2478 416 -2476
rect 422 -2472 423 -2470
rect 422 -2478 423 -2476
rect 432 -2472 433 -2470
rect 432 -2478 433 -2476
rect 436 -2472 437 -2470
rect 436 -2478 437 -2476
rect 443 -2472 444 -2470
rect 443 -2478 444 -2476
rect 450 -2472 451 -2470
rect 450 -2478 451 -2476
rect 457 -2472 458 -2470
rect 457 -2478 458 -2476
rect 467 -2478 468 -2476
rect 471 -2472 472 -2470
rect 471 -2478 472 -2476
rect 478 -2472 479 -2470
rect 478 -2478 479 -2476
rect 502 -2472 503 -2470
rect 502 -2478 503 -2476
rect 506 -2472 507 -2470
rect 506 -2478 507 -2476
rect 513 -2472 514 -2470
rect 513 -2478 514 -2476
rect 520 -2478 521 -2476
rect 523 -2478 524 -2476
rect 527 -2478 528 -2476
rect 534 -2472 535 -2470
rect 537 -2478 538 -2476
rect 541 -2472 542 -2470
rect 541 -2478 542 -2476
rect 548 -2472 549 -2470
rect 548 -2478 549 -2476
rect 569 -2472 570 -2470
rect 569 -2478 570 -2476
rect 576 -2472 577 -2470
rect 576 -2478 577 -2476
rect 586 -2478 587 -2476
rect 593 -2472 594 -2470
rect 590 -2478 591 -2476
rect 600 -2472 601 -2470
rect 597 -2478 598 -2476
rect 604 -2472 605 -2470
rect 604 -2478 605 -2476
rect 611 -2472 612 -2470
rect 611 -2478 612 -2476
rect 625 -2472 626 -2470
rect 625 -2478 626 -2476
rect 639 -2472 640 -2470
rect 642 -2472 643 -2470
rect 660 -2472 661 -2470
rect 660 -2478 661 -2476
rect 674 -2472 675 -2470
rect 674 -2478 675 -2476
rect 681 -2472 682 -2470
rect 681 -2478 682 -2476
rect 688 -2472 689 -2470
rect 688 -2478 689 -2476
rect 695 -2472 696 -2470
rect 695 -2478 696 -2476
rect 709 -2472 710 -2470
rect 709 -2478 710 -2476
rect 716 -2472 717 -2470
rect 716 -2478 717 -2476
rect 723 -2472 724 -2470
rect 723 -2478 724 -2476
rect 730 -2472 731 -2470
rect 730 -2478 731 -2476
rect 737 -2472 738 -2470
rect 737 -2478 738 -2476
rect 758 -2472 759 -2470
rect 761 -2472 762 -2470
rect 758 -2478 759 -2476
rect 761 -2478 762 -2476
rect 765 -2472 766 -2470
rect 765 -2478 766 -2476
rect 884 -2472 885 -2470
rect 884 -2478 885 -2476
rect 891 -2472 892 -2470
rect 891 -2478 892 -2476
rect 933 -2472 934 -2470
rect 936 -2478 937 -2476
rect 940 -2472 941 -2470
rect 940 -2478 941 -2476
rect 5 -2499 6 -2497
rect 5 -2505 6 -2503
rect 86 -2499 87 -2497
rect 86 -2505 87 -2503
rect 96 -2499 97 -2497
rect 100 -2499 101 -2497
rect 100 -2505 101 -2503
rect 103 -2505 104 -2503
rect 110 -2499 111 -2497
rect 107 -2505 108 -2503
rect 114 -2499 115 -2497
rect 117 -2505 118 -2503
rect 121 -2499 122 -2497
rect 121 -2505 122 -2503
rect 138 -2499 139 -2497
rect 142 -2499 143 -2497
rect 142 -2505 143 -2503
rect 149 -2499 150 -2497
rect 149 -2505 150 -2503
rect 159 -2499 160 -2497
rect 156 -2505 157 -2503
rect 163 -2505 164 -2503
rect 166 -2505 167 -2503
rect 170 -2499 171 -2497
rect 170 -2505 171 -2503
rect 177 -2499 178 -2497
rect 177 -2505 178 -2503
rect 187 -2505 188 -2503
rect 191 -2505 192 -2503
rect 194 -2505 195 -2503
rect 201 -2499 202 -2497
rect 201 -2505 202 -2503
rect 205 -2499 206 -2497
rect 205 -2505 206 -2503
rect 212 -2499 213 -2497
rect 212 -2505 213 -2503
rect 219 -2499 220 -2497
rect 219 -2505 220 -2503
rect 226 -2499 227 -2497
rect 226 -2505 227 -2503
rect 233 -2499 234 -2497
rect 233 -2505 234 -2503
rect 240 -2499 241 -2497
rect 240 -2505 241 -2503
rect 247 -2499 248 -2497
rect 247 -2505 248 -2503
rect 254 -2499 255 -2497
rect 254 -2505 255 -2503
rect 261 -2499 262 -2497
rect 261 -2505 262 -2503
rect 271 -2499 272 -2497
rect 268 -2505 269 -2503
rect 275 -2499 276 -2497
rect 275 -2505 276 -2503
rect 282 -2505 283 -2503
rect 289 -2499 290 -2497
rect 289 -2505 290 -2503
rect 296 -2499 297 -2497
rect 299 -2505 300 -2503
rect 303 -2499 304 -2497
rect 303 -2505 304 -2503
rect 310 -2499 311 -2497
rect 310 -2505 311 -2503
rect 317 -2499 318 -2497
rect 317 -2505 318 -2503
rect 324 -2499 325 -2497
rect 324 -2505 325 -2503
rect 331 -2499 332 -2497
rect 331 -2505 332 -2503
rect 352 -2499 353 -2497
rect 352 -2505 353 -2503
rect 359 -2499 360 -2497
rect 362 -2499 363 -2497
rect 380 -2499 381 -2497
rect 380 -2505 381 -2503
rect 387 -2505 388 -2503
rect 394 -2499 395 -2497
rect 394 -2505 395 -2503
rect 401 -2499 402 -2497
rect 404 -2499 405 -2497
rect 401 -2505 402 -2503
rect 404 -2505 405 -2503
rect 408 -2499 409 -2497
rect 408 -2505 409 -2503
rect 418 -2505 419 -2503
rect 422 -2499 423 -2497
rect 443 -2499 444 -2497
rect 443 -2505 444 -2503
rect 450 -2499 451 -2497
rect 450 -2505 451 -2503
rect 520 -2499 521 -2497
rect 523 -2499 524 -2497
rect 527 -2499 528 -2497
rect 527 -2505 528 -2503
rect 604 -2499 605 -2497
rect 604 -2505 605 -2503
rect 611 -2499 612 -2497
rect 611 -2505 612 -2503
rect 660 -2499 661 -2497
rect 660 -2505 661 -2503
rect 667 -2499 668 -2497
rect 667 -2505 668 -2503
rect 681 -2499 682 -2497
rect 681 -2505 682 -2503
rect 688 -2499 689 -2497
rect 688 -2505 689 -2503
rect 695 -2499 696 -2497
rect 695 -2505 696 -2503
rect 702 -2505 703 -2503
rect 705 -2505 706 -2503
rect 709 -2499 710 -2497
rect 709 -2505 710 -2503
rect 716 -2499 717 -2497
rect 716 -2505 717 -2503
rect 723 -2499 724 -2497
rect 723 -2505 724 -2503
rect 730 -2499 731 -2497
rect 740 -2505 741 -2503
rect 744 -2499 745 -2497
rect 744 -2505 745 -2503
rect 751 -2499 752 -2497
rect 751 -2505 752 -2503
rect 758 -2499 759 -2497
rect 758 -2505 759 -2503
rect 884 -2499 885 -2497
rect 887 -2505 888 -2503
rect 891 -2499 892 -2497
rect 891 -2505 892 -2503
rect 933 -2499 934 -2497
rect 933 -2505 934 -2503
rect 940 -2505 941 -2503
rect 943 -2505 944 -2503
rect 947 -2499 948 -2497
rect 947 -2505 948 -2503
rect 5 -2524 6 -2522
rect 9 -2518 10 -2516
rect 9 -2524 10 -2522
rect 100 -2524 101 -2522
rect 107 -2518 108 -2516
rect 107 -2524 108 -2522
rect 114 -2518 115 -2516
rect 114 -2524 115 -2522
rect 121 -2524 122 -2522
rect 124 -2524 125 -2522
rect 131 -2524 132 -2522
rect 159 -2518 160 -2516
rect 163 -2518 164 -2516
rect 163 -2524 164 -2522
rect 170 -2524 171 -2522
rect 180 -2518 181 -2516
rect 180 -2524 181 -2522
rect 184 -2518 185 -2516
rect 184 -2524 185 -2522
rect 191 -2518 192 -2516
rect 191 -2524 192 -2522
rect 198 -2524 199 -2522
rect 226 -2518 227 -2516
rect 229 -2518 230 -2516
rect 271 -2518 272 -2516
rect 278 -2518 279 -2516
rect 285 -2518 286 -2516
rect 292 -2524 293 -2522
rect 296 -2518 297 -2516
rect 296 -2524 297 -2522
rect 303 -2524 304 -2522
rect 310 -2518 311 -2516
rect 310 -2524 311 -2522
rect 341 -2518 342 -2516
rect 341 -2524 342 -2522
rect 345 -2518 346 -2516
rect 345 -2524 346 -2522
rect 362 -2518 363 -2516
rect 383 -2518 384 -2516
rect 397 -2518 398 -2516
rect 404 -2518 405 -2516
rect 450 -2518 451 -2516
rect 450 -2524 451 -2522
rect 457 -2518 458 -2516
rect 457 -2524 458 -2522
rect 523 -2518 524 -2516
rect 597 -2518 598 -2516
rect 597 -2524 598 -2522
rect 604 -2518 605 -2516
rect 604 -2524 605 -2522
rect 663 -2518 664 -2516
rect 663 -2524 664 -2522
rect 667 -2518 668 -2516
rect 667 -2524 668 -2522
rect 688 -2518 689 -2516
rect 712 -2518 713 -2516
rect 716 -2518 717 -2516
rect 716 -2524 717 -2522
rect 723 -2524 724 -2522
rect 730 -2518 731 -2516
rect 730 -2524 731 -2522
rect 740 -2524 741 -2522
<< metal1 >>
rect 93 0 101 1
rect 107 0 129 1
rect 205 0 213 1
rect 215 0 237 1
rect 240 0 248 1
rect 261 0 269 1
rect 324 0 335 1
rect 429 0 451 1
rect 464 0 489 1
rect 530 0 535 1
rect 583 0 598 1
rect 660 0 668 1
rect 117 -2 122 -1
rect 226 -2 234 -1
rect 86 -13 104 -12
rect 117 -13 129 -12
rect 135 -13 146 -12
rect 173 -13 199 -12
rect 205 -13 216 -12
rect 226 -13 251 -12
rect 254 -13 269 -12
rect 289 -13 307 -12
rect 310 -13 325 -12
rect 348 -13 360 -12
rect 373 -13 447 -12
rect 450 -13 465 -12
rect 485 -13 528 -12
rect 534 -13 542 -12
rect 548 -13 570 -12
rect 590 -13 605 -12
rect 607 -13 619 -12
rect 667 -13 675 -12
rect 89 -15 101 -14
rect 177 -15 213 -14
rect 219 -15 227 -14
rect 233 -15 248 -14
rect 257 -15 276 -14
rect 317 -15 332 -14
rect 415 -15 430 -14
rect 453 -15 472 -14
rect 492 -15 514 -14
rect 562 -15 577 -14
rect 597 -15 612 -14
rect 93 -17 108 -16
rect 184 -17 206 -16
rect 219 -17 223 -16
rect 261 -17 283 -16
rect 324 -17 342 -16
rect 429 -17 440 -16
rect 506 -17 510 -16
rect 100 -19 122 -18
rect 236 -19 283 -18
rect 268 -21 304 -20
rect 86 -32 104 -31
rect 114 -32 188 -31
rect 191 -32 220 -31
rect 226 -32 230 -31
rect 247 -32 353 -31
rect 359 -32 409 -31
rect 415 -32 423 -31
rect 429 -32 437 -31
rect 446 -32 500 -31
rect 520 -32 535 -31
rect 551 -32 563 -31
rect 569 -32 598 -31
rect 604 -32 640 -31
rect 663 -32 668 -31
rect 674 -32 703 -31
rect 765 -32 843 -31
rect 93 -34 101 -33
rect 121 -34 136 -33
rect 163 -34 237 -33
rect 247 -34 255 -33
rect 275 -34 346 -33
rect 366 -34 374 -33
rect 383 -34 395 -33
rect 471 -34 521 -33
rect 527 -34 591 -33
rect 611 -34 654 -33
rect 677 -34 682 -33
rect 128 -36 146 -35
rect 177 -36 195 -35
rect 198 -36 206 -35
rect 212 -36 276 -35
rect 282 -36 304 -35
rect 313 -36 318 -35
rect 341 -36 423 -35
rect 464 -36 612 -35
rect 618 -36 647 -35
rect 135 -38 269 -37
rect 282 -38 349 -37
rect 373 -38 444 -37
rect 464 -38 626 -37
rect 156 -40 178 -39
rect 184 -40 220 -39
rect 226 -40 262 -39
rect 268 -40 290 -39
rect 296 -40 430 -39
rect 471 -40 587 -39
rect 198 -42 332 -41
rect 383 -42 486 -41
rect 527 -42 633 -41
rect 201 -44 255 -43
rect 289 -44 325 -43
rect 387 -44 468 -43
rect 478 -44 493 -43
rect 541 -44 570 -43
rect 173 -46 325 -45
rect 513 -46 542 -45
rect 555 -46 605 -45
rect 212 -48 300 -47
rect 310 -48 318 -47
rect 555 -48 773 -47
rect 229 -50 262 -49
rect 250 -52 402 -51
rect 30 -63 153 -62
rect 159 -63 251 -62
rect 317 -63 339 -62
rect 429 -63 822 -62
rect 842 -63 878 -62
rect 58 -65 108 -64
rect 114 -65 174 -64
rect 198 -65 206 -64
rect 219 -65 230 -64
rect 233 -65 346 -64
rect 394 -65 430 -64
rect 450 -65 468 -64
rect 471 -65 475 -64
rect 485 -65 514 -64
rect 530 -65 689 -64
rect 702 -65 780 -64
rect 37 -67 174 -66
rect 219 -67 279 -66
rect 317 -67 717 -66
rect 772 -67 871 -66
rect 61 -69 321 -68
rect 324 -69 381 -68
rect 457 -69 556 -68
rect 583 -69 794 -68
rect 65 -71 94 -70
rect 100 -71 206 -70
rect 233 -71 388 -70
rect 464 -71 479 -70
rect 485 -71 500 -70
rect 502 -71 808 -70
rect 72 -73 129 -72
rect 142 -73 244 -72
rect 254 -73 556 -72
rect 590 -73 773 -72
rect 79 -75 87 -74
rect 93 -75 304 -74
rect 331 -75 696 -74
rect 702 -75 766 -74
rect 86 -77 283 -76
rect 289 -77 325 -76
rect 331 -77 353 -76
rect 376 -77 479 -76
rect 495 -77 829 -76
rect 103 -79 283 -78
rect 380 -79 409 -78
rect 471 -79 493 -78
rect 506 -79 510 -78
rect 548 -79 619 -78
rect 625 -79 815 -78
rect 117 -81 171 -80
rect 240 -81 409 -80
rect 474 -81 493 -80
rect 569 -81 626 -80
rect 632 -81 787 -80
rect 51 -83 241 -82
rect 261 -83 304 -82
rect 355 -83 633 -82
rect 639 -83 745 -82
rect 121 -85 255 -84
rect 268 -85 290 -84
rect 387 -85 836 -84
rect 121 -87 164 -86
rect 247 -87 262 -86
rect 268 -87 374 -86
rect 397 -87 549 -86
rect 586 -87 591 -86
rect 604 -87 738 -86
rect 128 -89 675 -88
rect 681 -89 731 -88
rect 149 -91 157 -90
rect 163 -91 419 -90
rect 527 -91 587 -90
rect 597 -91 682 -90
rect 709 -91 843 -90
rect 401 -93 570 -92
rect 576 -93 598 -92
rect 611 -93 724 -92
rect 366 -95 402 -94
rect 443 -95 612 -94
rect 646 -95 759 -94
rect 359 -97 647 -96
rect 653 -97 752 -96
rect 226 -99 360 -98
rect 436 -99 444 -98
rect 520 -99 654 -98
rect 660 -99 766 -98
rect 177 -101 227 -100
rect 310 -101 521 -100
rect 534 -101 640 -100
rect 667 -101 801 -100
rect 156 -103 668 -102
rect 177 -105 213 -104
rect 310 -105 342 -104
rect 415 -105 437 -104
rect 499 -105 535 -104
rect 541 -105 605 -104
rect 191 -107 213 -106
rect 422 -107 542 -106
rect 562 -107 577 -106
rect 47 -109 423 -108
rect 191 -111 391 -110
rect 296 -113 563 -112
rect 275 -115 297 -114
rect 184 -117 276 -116
rect 135 -119 185 -118
rect 135 -121 367 -120
rect 23 -132 122 -131
rect 128 -132 209 -131
rect 226 -132 689 -131
rect 723 -132 864 -131
rect 870 -132 955 -131
rect 30 -134 136 -133
rect 145 -134 416 -133
rect 499 -134 640 -133
rect 751 -134 871 -133
rect 877 -134 913 -133
rect 30 -136 164 -135
rect 170 -136 829 -135
rect 37 -138 101 -137
rect 149 -138 178 -137
rect 250 -138 836 -137
rect 37 -140 206 -139
rect 275 -140 311 -139
rect 317 -140 493 -139
rect 509 -140 738 -139
rect 765 -140 892 -139
rect 44 -142 143 -141
rect 156 -142 822 -141
rect 51 -144 276 -143
rect 299 -144 353 -143
rect 362 -144 920 -143
rect 51 -146 125 -145
rect 142 -146 374 -145
rect 376 -146 570 -145
rect 579 -146 759 -145
rect 772 -146 906 -145
rect 58 -148 647 -147
rect 660 -148 759 -147
rect 779 -148 885 -147
rect 65 -150 115 -149
rect 117 -150 157 -149
rect 159 -150 349 -149
rect 352 -150 542 -149
rect 548 -150 850 -149
rect 79 -152 675 -151
rect 681 -152 780 -151
rect 786 -152 927 -151
rect 79 -154 153 -153
rect 163 -154 199 -153
rect 310 -154 472 -153
rect 495 -154 661 -153
rect 667 -154 766 -153
rect 793 -154 934 -153
rect 86 -156 398 -155
rect 418 -156 640 -155
rect 695 -156 822 -155
rect 89 -158 129 -157
rect 152 -158 857 -157
rect 114 -160 181 -159
rect 198 -160 213 -159
rect 317 -160 409 -159
rect 422 -160 500 -159
rect 513 -160 542 -159
rect 583 -160 899 -159
rect 170 -162 216 -161
rect 320 -162 402 -161
rect 429 -162 514 -161
rect 520 -162 549 -161
rect 583 -162 731 -161
rect 737 -162 878 -161
rect 173 -164 458 -163
rect 464 -164 472 -163
rect 492 -164 696 -163
rect 702 -164 773 -163
rect 800 -164 941 -163
rect 212 -166 304 -165
rect 324 -166 356 -165
rect 359 -166 409 -165
rect 443 -166 787 -165
rect 814 -166 948 -165
rect 65 -168 360 -167
rect 380 -168 465 -167
rect 506 -168 801 -167
rect 93 -170 381 -169
rect 387 -170 430 -169
rect 520 -170 836 -169
rect 93 -172 185 -171
rect 219 -172 304 -171
rect 324 -172 689 -171
rect 709 -172 752 -171
rect 135 -174 220 -173
rect 261 -174 507 -173
rect 523 -174 724 -173
rect 107 -176 262 -175
rect 327 -176 339 -175
rect 345 -176 423 -175
rect 534 -176 570 -175
rect 590 -176 647 -175
rect 716 -176 829 -175
rect 184 -178 192 -177
rect 268 -178 339 -177
rect 348 -178 528 -177
rect 597 -178 731 -177
rect 72 -180 598 -179
rect 611 -180 668 -179
rect 72 -182 703 -181
rect 191 -184 230 -183
rect 268 -184 290 -183
rect 331 -184 444 -183
rect 450 -184 535 -183
rect 555 -184 612 -183
rect 618 -184 710 -183
rect 205 -186 290 -185
rect 334 -186 843 -185
rect 366 -188 451 -187
rect 478 -188 556 -187
rect 618 -188 843 -187
rect 296 -190 367 -189
rect 394 -190 682 -189
rect 282 -192 395 -191
rect 401 -192 675 -191
rect 240 -194 283 -193
rect 296 -194 591 -193
rect 625 -194 794 -193
rect 240 -196 255 -195
rect 478 -196 563 -195
rect 625 -196 815 -195
rect 233 -198 255 -197
rect 345 -198 563 -197
rect 632 -198 717 -197
rect 58 -200 234 -199
rect 485 -200 528 -199
rect 604 -200 633 -199
rect 110 -202 486 -201
rect 576 -202 605 -201
rect 576 -204 745 -203
rect 653 -206 745 -205
rect 653 -208 808 -207
rect 656 -210 808 -209
rect 16 -221 703 -220
rect 723 -221 909 -220
rect 23 -223 209 -222
rect 261 -223 346 -222
rect 352 -223 388 -222
rect 401 -223 829 -222
rect 887 -223 913 -222
rect 23 -225 80 -224
rect 114 -225 234 -224
rect 254 -225 388 -224
rect 471 -225 493 -224
rect 495 -225 906 -224
rect 30 -227 363 -226
rect 366 -227 405 -226
rect 502 -227 556 -226
rect 579 -227 927 -226
rect 30 -229 157 -228
rect 163 -229 223 -228
rect 296 -229 395 -228
rect 555 -229 612 -228
rect 618 -229 864 -228
rect 44 -231 139 -230
rect 142 -231 535 -230
rect 611 -231 668 -230
rect 674 -231 906 -230
rect 51 -233 255 -232
rect 299 -233 402 -232
rect 621 -233 899 -232
rect 51 -235 59 -234
rect 65 -235 262 -234
rect 299 -235 409 -234
rect 618 -235 899 -234
rect 58 -237 468 -236
rect 625 -237 661 -236
rect 663 -237 668 -236
rect 674 -237 689 -236
rect 702 -237 780 -236
rect 807 -237 864 -236
rect 65 -239 108 -238
rect 121 -239 563 -238
rect 628 -239 934 -238
rect 68 -241 367 -240
rect 408 -241 437 -240
rect 541 -241 563 -240
rect 639 -241 913 -240
rect 72 -243 304 -242
rect 317 -243 472 -242
rect 541 -243 549 -242
rect 597 -243 640 -242
rect 653 -243 948 -242
rect 72 -245 339 -244
rect 359 -245 479 -244
rect 527 -245 549 -244
rect 597 -245 710 -244
rect 723 -245 731 -244
rect 737 -245 745 -244
rect 800 -245 808 -244
rect 828 -245 885 -244
rect 79 -247 115 -246
rect 121 -247 171 -246
rect 177 -247 276 -246
rect 289 -247 304 -246
rect 317 -247 535 -246
rect 653 -247 717 -246
rect 730 -247 773 -246
rect 93 -249 276 -248
rect 324 -249 850 -248
rect 100 -251 157 -250
rect 170 -251 857 -250
rect 100 -253 150 -252
rect 173 -253 290 -252
rect 324 -253 521 -252
rect 688 -253 752 -252
rect 814 -253 850 -252
rect 856 -253 920 -252
rect 117 -255 150 -254
rect 177 -255 185 -254
rect 194 -255 507 -254
rect 695 -255 801 -254
rect 814 -255 836 -254
rect 919 -255 955 -254
rect 93 -257 185 -256
rect 198 -257 227 -256
rect 240 -257 696 -256
rect 709 -257 759 -256
rect 37 -259 241 -258
rect 331 -259 465 -258
rect 485 -259 773 -258
rect 37 -261 248 -260
rect 331 -261 570 -260
rect 740 -261 780 -260
rect 47 -263 199 -262
rect 219 -263 479 -262
rect 485 -263 941 -262
rect 135 -265 167 -264
rect 219 -265 230 -264
rect 247 -265 269 -264
rect 338 -265 381 -264
rect 397 -265 836 -264
rect 86 -267 136 -266
rect 142 -267 213 -266
rect 282 -267 381 -266
rect 436 -267 787 -266
rect 128 -269 269 -268
rect 282 -269 356 -268
rect 362 -269 591 -268
rect 744 -269 766 -268
rect 191 -271 213 -270
rect 450 -271 528 -270
rect 583 -271 787 -270
rect 191 -273 430 -272
rect 443 -273 584 -272
rect 590 -273 633 -272
rect 751 -273 822 -272
rect 334 -275 430 -274
rect 488 -275 717 -274
rect 758 -275 794 -274
rect 821 -275 843 -274
rect 415 -277 444 -276
rect 506 -277 514 -276
rect 632 -277 682 -276
rect 793 -277 871 -276
rect 152 -279 514 -278
rect 842 -279 878 -278
rect 257 -281 682 -280
rect 870 -281 892 -280
rect 310 -283 416 -282
rect 422 -283 451 -282
rect 576 -283 878 -282
rect 310 -285 521 -284
rect 373 -287 423 -286
rect 457 -287 577 -286
rect 373 -289 766 -288
rect 457 -291 500 -290
rect 499 -293 570 -292
rect 16 -304 185 -303
rect 240 -304 475 -303
rect 492 -304 521 -303
rect 523 -304 857 -303
rect 863 -304 906 -303
rect 23 -306 101 -305
rect 110 -306 122 -305
rect 124 -306 132 -305
rect 159 -306 251 -305
rect 254 -306 388 -305
rect 394 -306 885 -305
rect 898 -306 913 -305
rect 23 -308 209 -307
rect 233 -308 241 -307
rect 247 -308 321 -307
rect 352 -308 468 -307
rect 544 -308 654 -307
rect 660 -308 745 -307
rect 800 -308 881 -307
rect 30 -310 353 -309
rect 355 -310 507 -309
rect 516 -310 745 -309
rect 835 -310 888 -309
rect 37 -312 97 -311
rect 100 -312 199 -311
rect 233 -312 629 -311
rect 681 -312 934 -311
rect 37 -314 300 -313
rect 306 -314 801 -313
rect 807 -314 836 -313
rect 863 -314 871 -313
rect 877 -314 892 -313
rect 44 -316 104 -315
rect 117 -316 157 -315
rect 170 -316 542 -315
rect 625 -316 654 -315
rect 786 -316 871 -315
rect 877 -316 920 -315
rect 47 -318 556 -317
rect 646 -318 682 -317
rect 716 -318 787 -317
rect 793 -318 808 -317
rect 58 -320 402 -319
rect 422 -320 489 -319
rect 541 -320 724 -319
rect 730 -320 794 -319
rect 58 -322 87 -321
rect 128 -322 136 -321
rect 149 -322 199 -321
rect 268 -322 500 -321
rect 576 -322 717 -321
rect 65 -324 374 -323
rect 439 -324 738 -323
rect 9 -326 66 -325
rect 68 -326 752 -325
rect 68 -328 87 -327
rect 128 -328 164 -327
rect 173 -328 640 -327
rect 702 -328 752 -327
rect 79 -330 115 -329
rect 135 -330 724 -329
rect 79 -332 850 -331
rect 82 -334 507 -333
rect 527 -334 577 -333
rect 597 -334 731 -333
rect 842 -334 850 -333
rect 149 -336 220 -335
rect 268 -336 276 -335
rect 296 -336 444 -335
rect 464 -336 773 -335
rect 16 -338 220 -337
rect 275 -338 486 -337
rect 513 -338 528 -337
rect 583 -338 598 -337
rect 618 -338 640 -337
rect 674 -338 703 -337
rect 709 -338 738 -337
rect 772 -338 780 -337
rect 163 -340 188 -339
rect 191 -340 402 -339
rect 404 -340 619 -339
rect 667 -340 675 -339
rect 688 -340 843 -339
rect 170 -342 192 -341
rect 205 -342 584 -341
rect 709 -342 895 -341
rect 173 -344 332 -343
rect 345 -344 689 -343
rect 779 -344 829 -343
rect 72 -346 346 -345
rect 359 -346 671 -345
rect 814 -346 829 -345
rect 72 -348 122 -347
rect 205 -348 216 -347
rect 289 -348 297 -347
rect 310 -348 388 -347
rect 408 -348 486 -347
rect 513 -348 591 -347
rect 814 -348 822 -347
rect 194 -350 822 -349
rect 226 -352 290 -351
rect 310 -352 416 -351
rect 443 -352 696 -351
rect 212 -354 227 -353
rect 247 -354 416 -353
rect 450 -354 465 -353
rect 471 -354 647 -353
rect 257 -356 409 -355
rect 562 -356 591 -355
rect 632 -356 696 -355
rect 264 -358 563 -357
rect 604 -358 633 -357
rect 282 -360 451 -359
rect 142 -362 283 -361
rect 317 -362 612 -361
rect 107 -364 143 -363
rect 320 -364 423 -363
rect 429 -364 605 -363
rect 107 -366 857 -365
rect 324 -368 430 -367
rect 534 -368 612 -367
rect 324 -370 766 -369
rect 331 -372 885 -371
rect 341 -374 360 -373
rect 366 -374 556 -373
rect 758 -374 766 -373
rect 303 -376 367 -375
rect 373 -376 458 -375
rect 534 -376 570 -375
rect 51 -378 304 -377
rect 338 -378 458 -377
rect 548 -378 570 -377
rect 51 -380 94 -379
rect 380 -380 549 -379
rect 436 -382 759 -381
rect 397 -384 437 -383
rect 397 -386 479 -385
rect 166 -388 479 -387
rect 2 -399 580 -398
rect 611 -399 997 -398
rect 1108 -399 1116 -398
rect 9 -401 31 -400
rect 44 -401 139 -400
rect 145 -401 444 -400
rect 474 -401 843 -400
rect 849 -401 976 -400
rect 982 -401 1032 -400
rect 16 -403 101 -402
rect 107 -403 332 -402
rect 338 -403 367 -402
rect 380 -403 514 -402
rect 569 -403 612 -402
rect 628 -403 871 -402
rect 884 -403 899 -402
rect 933 -403 1046 -402
rect 23 -405 157 -404
rect 170 -405 801 -404
rect 807 -405 955 -404
rect 989 -405 1039 -404
rect 23 -407 52 -406
rect 58 -407 367 -406
rect 380 -407 507 -406
rect 569 -407 822 -406
rect 828 -407 927 -406
rect 37 -409 332 -408
rect 341 -409 402 -408
rect 422 -409 444 -408
rect 474 -409 1025 -408
rect 44 -411 276 -410
rect 296 -411 304 -410
rect 306 -411 808 -410
rect 863 -411 1011 -410
rect 51 -413 311 -412
rect 327 -413 689 -412
rect 702 -413 829 -412
rect 835 -413 864 -412
rect 891 -413 1018 -412
rect 65 -415 584 -414
rect 625 -415 934 -414
rect 79 -417 353 -416
rect 383 -417 549 -416
rect 572 -417 962 -416
rect 79 -419 129 -418
rect 135 -419 521 -418
rect 576 -419 626 -418
rect 635 -419 794 -418
rect 814 -419 892 -418
rect 82 -421 703 -420
rect 709 -421 801 -420
rect 96 -423 822 -422
rect 100 -425 423 -424
rect 478 -425 584 -424
rect 632 -425 710 -424
rect 723 -425 843 -424
rect 114 -427 472 -426
rect 485 -427 549 -426
rect 576 -427 850 -426
rect 117 -429 857 -428
rect 121 -431 388 -430
rect 397 -431 647 -430
rect 667 -431 857 -430
rect 86 -433 388 -432
rect 401 -433 500 -432
rect 506 -433 559 -432
rect 590 -433 647 -432
rect 667 -433 752 -432
rect 765 -433 899 -432
rect 72 -435 87 -434
rect 121 -435 164 -434
rect 170 -435 262 -434
rect 264 -435 563 -434
rect 590 -435 605 -434
rect 681 -435 766 -434
rect 772 -435 913 -434
rect 72 -437 132 -436
rect 149 -437 164 -436
rect 184 -437 619 -436
rect 639 -437 773 -436
rect 786 -437 948 -436
rect 61 -439 619 -438
rect 653 -439 787 -438
rect 149 -441 374 -440
rect 408 -441 521 -440
rect 534 -441 605 -440
rect 688 -441 871 -440
rect 12 -443 409 -442
rect 429 -443 486 -442
rect 492 -443 920 -442
rect 156 -445 178 -444
rect 184 -445 192 -444
rect 198 -445 262 -444
rect 268 -445 321 -444
rect 327 -445 458 -444
rect 460 -445 752 -444
rect 177 -447 213 -446
rect 219 -447 297 -446
rect 352 -447 1004 -446
rect 180 -449 220 -448
rect 233 -449 311 -448
rect 373 -449 528 -448
rect 534 -449 661 -448
rect 716 -449 724 -448
rect 730 -449 885 -448
rect 187 -451 416 -450
rect 425 -451 661 -450
rect 695 -451 731 -450
rect 737 -451 969 -450
rect 191 -453 878 -452
rect 198 -455 227 -454
rect 233 -455 395 -454
rect 429 -455 437 -454
rect 450 -455 528 -454
rect 597 -455 717 -454
rect 744 -455 836 -454
rect 205 -457 227 -456
rect 247 -457 269 -456
rect 275 -457 503 -456
rect 516 -457 738 -456
rect 758 -457 878 -456
rect 93 -459 206 -458
rect 240 -459 248 -458
rect 250 -459 290 -458
rect 317 -459 437 -458
rect 457 -459 941 -458
rect 93 -461 125 -460
rect 142 -461 241 -460
rect 254 -461 1035 -460
rect 68 -463 255 -462
rect 282 -463 384 -462
rect 481 -463 654 -462
rect 674 -463 745 -462
rect 110 -465 318 -464
rect 359 -465 451 -464
rect 495 -465 794 -464
rect 142 -467 682 -466
rect 695 -467 780 -466
rect 173 -469 290 -468
rect 345 -469 360 -468
rect 499 -469 598 -468
rect 30 -471 346 -470
rect 541 -471 675 -470
rect 324 -473 542 -472
rect 544 -473 759 -472
rect 37 -475 325 -474
rect 555 -475 780 -474
rect 492 -477 556 -476
rect 9 -488 633 -487
rect 814 -488 1032 -487
rect 1111 -488 1123 -487
rect 30 -490 34 -489
rect 44 -490 283 -489
rect 285 -490 619 -489
rect 765 -490 815 -489
rect 817 -490 836 -489
rect 954 -490 1039 -489
rect 1115 -490 1130 -489
rect 23 -492 619 -491
rect 772 -492 836 -491
rect 975 -492 1053 -491
rect 30 -494 213 -493
rect 296 -494 356 -493
rect 373 -494 531 -493
rect 555 -494 913 -493
rect 1010 -494 1060 -493
rect 33 -496 213 -495
rect 296 -496 311 -495
rect 317 -496 1074 -495
rect 37 -498 283 -497
rect 310 -498 493 -497
rect 499 -498 552 -497
rect 565 -498 969 -497
rect 1017 -498 1067 -497
rect 44 -500 402 -499
rect 415 -500 766 -499
rect 842 -500 1018 -499
rect 1024 -500 1095 -499
rect 16 -502 416 -501
rect 422 -502 605 -501
rect 709 -502 773 -501
rect 863 -502 976 -501
rect 1045 -502 1116 -501
rect 16 -504 353 -503
rect 359 -504 374 -503
rect 397 -504 808 -503
rect 926 -504 969 -503
rect 982 -504 1046 -503
rect 58 -506 73 -505
rect 79 -506 143 -505
rect 149 -506 395 -505
rect 401 -506 419 -505
rect 425 -506 997 -505
rect 61 -508 640 -507
rect 695 -508 927 -507
rect 940 -508 1011 -507
rect 26 -510 941 -509
rect 65 -512 304 -511
rect 327 -512 423 -511
rect 443 -512 479 -511
rect 481 -512 780 -511
rect 800 -512 864 -511
rect 891 -512 983 -511
rect 72 -514 584 -513
rect 597 -514 843 -513
rect 856 -514 892 -513
rect 919 -514 997 -513
rect 79 -516 94 -515
rect 96 -516 241 -515
rect 261 -516 318 -515
rect 338 -516 461 -515
rect 464 -516 472 -515
rect 474 -516 591 -515
rect 597 -516 829 -515
rect 877 -516 920 -515
rect 51 -518 472 -517
rect 485 -518 493 -517
rect 502 -518 731 -517
rect 758 -518 808 -517
rect 51 -520 332 -519
rect 341 -520 633 -519
rect 712 -520 829 -519
rect 100 -522 360 -521
rect 383 -522 857 -521
rect 2 -524 101 -523
rect 114 -524 381 -523
rect 436 -524 486 -523
rect 506 -524 591 -523
rect 600 -524 955 -523
rect 114 -526 209 -525
rect 261 -526 269 -525
rect 271 -526 780 -525
rect 121 -528 563 -527
rect 569 -528 605 -527
rect 716 -528 801 -527
rect 128 -530 388 -529
rect 457 -530 885 -529
rect 107 -532 388 -531
rect 429 -532 458 -531
rect 506 -532 661 -531
rect 758 -532 850 -531
rect 107 -534 822 -533
rect 128 -536 206 -535
rect 303 -536 437 -535
rect 523 -536 899 -535
rect 135 -538 430 -537
rect 534 -538 710 -537
rect 723 -538 899 -537
rect 135 -540 255 -539
rect 324 -540 885 -539
rect 142 -542 276 -541
rect 324 -542 451 -541
rect 534 -542 696 -541
rect 723 -542 787 -541
rect 145 -544 241 -543
rect 247 -544 255 -543
rect 275 -544 290 -543
rect 331 -544 685 -543
rect 688 -544 787 -543
rect 138 -546 290 -545
rect 345 -546 682 -545
rect 744 -546 822 -545
rect 149 -548 234 -547
rect 247 -548 269 -547
rect 348 -548 675 -547
rect 681 -548 934 -547
rect 86 -550 234 -549
rect 348 -550 444 -549
rect 450 -550 465 -549
rect 527 -550 675 -549
rect 702 -550 745 -549
rect 751 -550 850 -549
rect 86 -552 171 -551
rect 180 -552 227 -551
rect 366 -552 661 -551
rect 93 -554 934 -553
rect 156 -556 353 -555
rect 527 -556 584 -555
rect 611 -556 703 -555
rect 156 -558 216 -557
rect 537 -558 878 -557
rect 163 -560 171 -559
rect 191 -560 227 -559
rect 537 -560 668 -559
rect 163 -562 367 -561
rect 541 -562 752 -561
rect 166 -564 1025 -563
rect 184 -566 192 -565
rect 198 -566 1081 -565
rect 184 -568 220 -567
rect 513 -568 542 -567
rect 555 -568 566 -567
rect 572 -568 794 -567
rect 198 -570 209 -569
rect 219 -570 612 -569
rect 625 -570 717 -569
rect 737 -570 794 -569
rect 408 -572 738 -571
rect 408 -574 577 -573
rect 579 -574 913 -573
rect 513 -576 521 -575
rect 562 -576 1088 -575
rect 625 -578 654 -577
rect 548 -580 654 -579
rect 548 -582 1004 -581
rect 635 -584 668 -583
rect 989 -584 1004 -583
rect 642 -586 689 -585
rect 961 -586 990 -585
rect 905 -588 962 -587
rect 905 -590 948 -589
rect 870 -592 948 -591
rect 572 -594 871 -593
rect 2 -605 234 -604
rect 254 -605 269 -604
rect 289 -605 535 -604
rect 544 -605 1011 -604
rect 1111 -605 1144 -604
rect 2 -607 108 -606
rect 121 -607 269 -606
rect 310 -607 524 -606
rect 534 -607 647 -606
rect 684 -607 1053 -606
rect 1115 -607 1151 -606
rect 5 -609 528 -608
rect 548 -609 899 -608
rect 989 -609 1053 -608
rect 1101 -609 1116 -608
rect 1129 -609 1158 -608
rect 9 -611 213 -610
rect 338 -611 752 -610
rect 898 -611 1046 -610
rect 1094 -611 1102 -610
rect 1129 -611 1140 -610
rect 16 -613 349 -612
rect 362 -613 577 -612
rect 579 -613 1039 -612
rect 1066 -613 1095 -612
rect 16 -615 66 -614
rect 72 -615 517 -614
rect 541 -615 577 -614
rect 604 -615 1109 -614
rect 23 -617 129 -616
rect 135 -617 213 -616
rect 338 -617 458 -616
rect 460 -617 843 -616
rect 926 -617 1067 -616
rect 26 -619 59 -618
rect 65 -619 297 -618
rect 341 -619 612 -618
rect 709 -619 787 -618
rect 926 -619 934 -618
rect 961 -619 990 -618
rect 1024 -619 1046 -618
rect 37 -621 619 -620
rect 712 -621 1088 -620
rect 47 -623 346 -622
rect 366 -623 566 -622
rect 569 -623 738 -622
rect 786 -623 976 -622
rect 1031 -623 1088 -622
rect 51 -625 234 -624
rect 292 -625 612 -624
rect 618 -625 745 -624
rect 905 -625 976 -624
rect 982 -625 1032 -624
rect 44 -627 52 -626
rect 58 -627 171 -626
rect 173 -627 661 -626
rect 730 -627 808 -626
rect 870 -627 906 -626
rect 912 -627 962 -626
rect 968 -627 983 -626
rect 40 -629 661 -628
rect 726 -629 969 -628
rect 44 -631 766 -630
rect 933 -631 941 -630
rect 72 -633 80 -632
rect 86 -633 216 -632
rect 296 -633 598 -632
rect 604 -633 836 -632
rect 940 -633 948 -632
rect 86 -635 143 -634
rect 156 -635 255 -634
rect 317 -635 346 -634
rect 359 -635 367 -634
rect 380 -635 384 -634
rect 394 -635 542 -634
rect 548 -635 556 -634
rect 562 -635 1018 -634
rect 37 -637 360 -636
rect 380 -637 388 -636
rect 394 -637 451 -636
rect 453 -637 486 -636
rect 513 -637 570 -636
rect 572 -637 864 -636
rect 947 -637 955 -636
rect 1003 -637 1018 -636
rect 93 -639 1074 -638
rect 93 -641 220 -640
rect 313 -641 318 -640
rect 387 -641 591 -640
rect 597 -641 689 -640
rect 765 -641 773 -640
rect 828 -641 836 -640
rect 863 -641 920 -640
rect 1059 -641 1074 -640
rect 100 -643 997 -642
rect 100 -645 132 -644
rect 135 -645 223 -644
rect 383 -645 591 -644
rect 625 -645 920 -644
rect 107 -647 185 -646
rect 201 -647 640 -646
rect 688 -647 734 -646
rect 789 -647 997 -646
rect 114 -649 808 -648
rect 117 -651 157 -650
rect 163 -651 283 -650
rect 401 -651 486 -650
rect 495 -651 640 -650
rect 723 -651 829 -650
rect 128 -653 1039 -652
rect 138 -655 801 -654
rect 142 -657 150 -656
rect 163 -657 262 -656
rect 275 -657 283 -656
rect 408 -657 556 -656
rect 562 -657 843 -656
rect 30 -659 150 -658
rect 177 -659 1004 -658
rect 30 -661 83 -660
rect 124 -661 262 -660
rect 275 -661 458 -660
rect 467 -661 654 -660
rect 723 -661 913 -660
rect 177 -663 192 -662
rect 205 -663 353 -662
rect 408 -663 479 -662
rect 513 -663 647 -662
rect 653 -663 703 -662
rect 800 -663 815 -662
rect 184 -665 199 -664
rect 205 -665 325 -664
rect 352 -665 493 -664
rect 520 -665 871 -664
rect 219 -667 248 -666
rect 415 -667 437 -666
rect 439 -667 1011 -666
rect 191 -669 248 -668
rect 415 -669 479 -668
rect 492 -669 675 -668
rect 702 -669 857 -668
rect 226 -671 402 -670
rect 429 -671 626 -670
rect 632 -671 955 -670
rect 422 -673 430 -672
rect 443 -673 521 -672
rect 551 -673 738 -672
rect 775 -673 815 -672
rect 856 -673 892 -672
rect 324 -675 444 -674
rect 450 -675 682 -674
rect 884 -675 892 -674
rect 422 -677 507 -676
rect 583 -677 633 -676
rect 674 -677 696 -676
rect 877 -677 885 -676
rect 103 -679 507 -678
rect 583 -679 608 -678
rect 667 -679 696 -678
rect 849 -679 878 -678
rect 467 -681 1025 -680
rect 471 -683 752 -682
rect 849 -683 1081 -682
rect 471 -685 500 -684
rect 667 -685 759 -684
rect 474 -687 1060 -686
rect 481 -689 500 -688
rect 758 -689 822 -688
rect 716 -691 822 -690
rect 331 -693 717 -692
rect 331 -695 1081 -694
rect 2 -706 115 -705
rect 128 -706 157 -705
rect 208 -706 293 -705
rect 310 -706 486 -705
rect 513 -706 892 -705
rect 936 -706 969 -705
rect 1080 -706 1144 -705
rect 16 -708 370 -707
rect 443 -708 773 -707
rect 775 -708 1032 -707
rect 1083 -708 1151 -707
rect 30 -710 199 -709
rect 268 -710 272 -709
rect 292 -710 402 -709
rect 446 -710 822 -709
rect 880 -710 885 -709
rect 891 -710 1011 -709
rect 1031 -710 1130 -709
rect 44 -712 52 -711
rect 58 -712 290 -711
rect 327 -712 423 -711
rect 436 -712 447 -711
rect 450 -712 591 -711
rect 604 -712 801 -711
rect 821 -712 871 -711
rect 884 -712 948 -711
rect 968 -712 1102 -711
rect 1111 -712 1158 -711
rect 51 -714 157 -713
rect 177 -714 199 -713
rect 268 -714 276 -713
rect 289 -714 472 -713
rect 478 -714 920 -713
rect 58 -716 297 -715
rect 317 -716 423 -715
rect 436 -716 444 -715
rect 453 -716 570 -715
rect 590 -716 941 -715
rect 82 -718 90 -717
rect 114 -718 136 -717
rect 142 -718 160 -717
rect 163 -718 178 -717
rect 233 -718 297 -717
rect 317 -718 395 -717
rect 401 -718 500 -717
rect 516 -718 717 -717
rect 723 -718 955 -717
rect 121 -720 479 -719
rect 485 -720 584 -719
rect 639 -720 664 -719
rect 705 -720 913 -719
rect 919 -720 1004 -719
rect 93 -722 122 -721
rect 131 -722 346 -721
rect 352 -722 461 -721
rect 467 -722 808 -721
rect 870 -722 899 -721
rect 912 -722 997 -721
rect 1003 -722 1046 -721
rect 93 -724 332 -723
rect 338 -724 493 -723
rect 541 -724 647 -723
rect 653 -724 668 -723
rect 688 -724 808 -723
rect 877 -724 899 -723
rect 940 -724 990 -723
rect 996 -724 1018 -723
rect 135 -726 153 -725
rect 163 -726 185 -725
rect 205 -726 332 -725
rect 352 -726 381 -725
rect 457 -726 619 -725
rect 639 -726 675 -725
rect 688 -726 710 -725
rect 716 -726 1053 -725
rect 142 -728 150 -727
rect 173 -728 461 -727
rect 471 -728 507 -727
rect 513 -728 619 -727
rect 646 -728 682 -727
rect 709 -728 731 -727
rect 737 -728 745 -727
rect 747 -728 801 -727
rect 989 -728 1095 -727
rect 65 -730 150 -729
rect 184 -730 388 -729
rect 457 -730 934 -729
rect 37 -732 66 -731
rect 226 -732 339 -731
rect 359 -732 367 -731
rect 380 -732 538 -731
rect 544 -732 1039 -731
rect 30 -734 38 -733
rect 226 -734 727 -733
rect 730 -734 794 -733
rect 863 -734 934 -733
rect 233 -736 255 -735
rect 261 -736 500 -735
rect 506 -736 521 -735
rect 555 -736 570 -735
rect 583 -736 720 -735
rect 723 -736 766 -735
rect 775 -736 976 -735
rect 79 -738 766 -737
rect 786 -738 962 -737
rect 79 -740 87 -739
rect 240 -740 255 -739
rect 261 -740 409 -739
rect 464 -740 521 -739
rect 534 -740 556 -739
rect 562 -740 738 -739
rect 751 -740 951 -739
rect 954 -740 976 -739
rect 23 -742 87 -741
rect 240 -742 304 -741
rect 310 -742 346 -741
rect 362 -742 430 -741
rect 495 -742 675 -741
rect 681 -742 696 -741
rect 702 -742 752 -741
rect 758 -742 773 -741
rect 786 -742 815 -741
rect 856 -742 864 -741
rect 23 -744 125 -743
rect 219 -744 304 -743
rect 324 -744 360 -743
rect 387 -744 416 -743
rect 534 -744 563 -743
rect 597 -744 962 -743
rect 100 -746 430 -745
rect 597 -746 836 -745
rect 856 -746 927 -745
rect 100 -748 192 -747
rect 208 -748 416 -747
rect 653 -748 1067 -747
rect 107 -750 192 -749
rect 212 -750 220 -749
rect 271 -750 276 -749
rect 324 -750 395 -749
rect 408 -750 549 -749
rect 656 -750 696 -749
rect 702 -750 1074 -749
rect 107 -752 248 -751
rect 548 -752 661 -751
rect 758 -752 1060 -751
rect 103 -754 248 -753
rect 660 -754 829 -753
rect 835 -754 983 -753
rect 170 -756 213 -755
rect 814 -756 906 -755
rect 926 -756 1116 -755
rect 9 -758 171 -757
rect 828 -758 843 -757
rect 849 -758 906 -757
rect 982 -758 1088 -757
rect 527 -760 843 -759
rect 849 -760 1025 -759
rect 527 -762 577 -761
rect 576 -764 612 -763
rect 611 -766 626 -765
rect 625 -768 633 -767
rect 632 -770 780 -769
rect 761 -772 780 -771
rect 2 -783 157 -782
rect 173 -783 468 -782
rect 492 -783 1018 -782
rect 1087 -783 1095 -782
rect 1108 -783 1154 -782
rect 16 -785 185 -784
rect 194 -785 395 -784
rect 408 -785 493 -784
rect 499 -785 664 -784
rect 667 -785 717 -784
rect 719 -785 745 -784
rect 779 -785 1046 -784
rect 1122 -785 1144 -784
rect 23 -787 139 -786
rect 149 -787 269 -786
rect 289 -787 346 -786
rect 355 -787 955 -786
rect 957 -787 997 -786
rect 1010 -787 1067 -786
rect 1139 -787 1151 -786
rect 23 -789 87 -788
rect 107 -789 328 -788
rect 341 -789 353 -788
rect 408 -789 482 -788
rect 506 -789 535 -788
rect 537 -789 633 -788
rect 646 -789 1102 -788
rect 30 -791 503 -790
rect 548 -791 668 -790
rect 674 -791 934 -790
rect 947 -791 1004 -790
rect 40 -793 619 -792
rect 621 -793 871 -792
rect 884 -793 1004 -792
rect 51 -795 171 -794
rect 177 -795 185 -794
rect 198 -795 206 -794
rect 208 -795 241 -794
rect 247 -795 507 -794
rect 513 -795 549 -794
rect 562 -795 619 -794
rect 653 -795 843 -794
rect 866 -795 1053 -794
rect 51 -797 461 -796
rect 464 -797 759 -796
rect 768 -797 1011 -796
rect 58 -799 531 -798
rect 541 -799 843 -798
rect 912 -799 997 -798
rect 58 -801 262 -800
rect 268 -801 451 -800
rect 453 -801 906 -800
rect 961 -801 1074 -800
rect 65 -803 101 -802
rect 128 -803 514 -802
rect 593 -803 1060 -802
rect 65 -805 73 -804
rect 75 -805 108 -804
rect 128 -805 227 -804
rect 240 -805 500 -804
rect 604 -805 633 -804
rect 653 -805 1123 -804
rect 86 -807 115 -806
rect 156 -807 325 -806
rect 345 -807 416 -806
rect 422 -807 451 -806
rect 457 -807 927 -806
rect 982 -807 1025 -806
rect 114 -809 297 -808
rect 310 -809 339 -808
rect 359 -809 465 -808
rect 478 -809 675 -808
rect 737 -809 1039 -808
rect 93 -811 297 -810
rect 313 -811 521 -810
rect 527 -811 983 -810
rect 989 -811 1116 -810
rect 93 -813 332 -812
rect 380 -813 528 -812
rect 607 -813 871 -812
rect 877 -813 990 -812
rect 152 -815 360 -814
rect 383 -815 535 -814
rect 614 -815 850 -814
rect 898 -815 906 -814
rect 926 -815 1032 -814
rect 177 -817 293 -816
rect 317 -817 416 -816
rect 422 -817 437 -816
rect 443 -817 591 -816
rect 656 -817 706 -816
rect 744 -817 937 -816
rect 142 -819 444 -818
rect 457 -819 486 -818
rect 495 -819 647 -818
rect 656 -819 948 -818
rect 142 -821 234 -820
rect 254 -821 332 -820
rect 387 -821 542 -820
rect 660 -821 1081 -820
rect 121 -823 255 -822
rect 317 -823 367 -822
rect 387 -823 430 -822
rect 436 -823 703 -822
rect 751 -823 850 -822
rect 863 -823 1032 -822
rect 79 -825 122 -824
rect 198 -825 213 -824
rect 222 -825 248 -824
rect 261 -825 367 -824
rect 401 -825 703 -824
rect 751 -825 941 -824
rect 212 -827 227 -826
rect 233 -827 447 -826
rect 471 -827 486 -826
rect 520 -827 776 -826
rect 779 -827 822 -826
rect 828 -827 878 -826
rect 324 -829 738 -828
rect 765 -829 962 -828
rect 401 -831 636 -830
rect 660 -831 682 -830
rect 723 -831 822 -830
rect 828 -831 976 -830
rect 135 -833 682 -832
rect 772 -833 913 -832
rect 135 -835 164 -834
rect 471 -835 612 -834
rect 688 -835 773 -834
rect 793 -835 920 -834
rect 163 -837 220 -836
rect 478 -837 598 -836
rect 604 -837 976 -836
rect 219 -839 304 -838
rect 555 -839 724 -838
rect 730 -839 794 -838
rect 807 -839 920 -838
rect 282 -841 304 -840
rect 555 -841 801 -840
rect 814 -841 899 -840
rect 191 -843 283 -842
rect 565 -843 766 -842
rect 786 -843 815 -842
rect 835 -843 885 -842
rect 103 -845 836 -844
rect 863 -845 969 -844
rect 82 -847 969 -846
rect 576 -849 598 -848
rect 611 -849 941 -848
rect 352 -851 577 -850
rect 579 -851 808 -850
rect 639 -853 689 -852
rect 695 -853 731 -852
rect 786 -853 857 -852
rect 338 -855 696 -854
rect 709 -855 801 -854
rect 856 -855 892 -854
rect 369 -857 892 -856
rect 394 -859 640 -858
rect 709 -859 797 -858
rect 9 -870 150 -869
rect 198 -870 220 -869
rect 222 -870 283 -869
rect 317 -870 433 -869
rect 481 -870 871 -869
rect 982 -870 1151 -869
rect 12 -872 381 -871
rect 383 -872 545 -871
rect 555 -872 1102 -871
rect 16 -874 153 -873
rect 170 -874 381 -873
rect 394 -874 913 -873
rect 989 -874 1102 -873
rect 30 -876 430 -875
rect 492 -876 580 -875
rect 583 -876 654 -875
rect 768 -876 1032 -875
rect 1052 -876 1158 -875
rect 30 -878 76 -877
rect 79 -878 766 -877
rect 779 -878 871 -877
rect 912 -878 934 -877
rect 1017 -878 1130 -877
rect 58 -880 447 -879
rect 478 -880 493 -879
rect 537 -880 920 -879
rect 933 -880 948 -879
rect 1087 -880 1095 -879
rect 1097 -880 1144 -879
rect 16 -882 59 -881
rect 65 -882 83 -881
rect 93 -882 503 -881
rect 565 -882 703 -881
rect 709 -882 1053 -881
rect 1115 -882 1130 -881
rect 72 -884 1137 -883
rect 75 -886 87 -885
rect 93 -886 157 -885
rect 170 -886 454 -885
rect 572 -886 822 -885
rect 856 -886 983 -885
rect 1108 -886 1116 -885
rect 79 -888 549 -887
rect 576 -888 1088 -887
rect 1108 -888 1123 -887
rect 86 -890 129 -889
rect 135 -890 192 -889
rect 198 -890 206 -889
rect 229 -890 556 -889
rect 562 -890 1123 -889
rect 51 -892 129 -891
rect 135 -892 269 -891
rect 310 -892 318 -891
rect 324 -892 500 -891
rect 548 -892 699 -891
rect 730 -892 822 -891
rect 905 -892 1144 -891
rect 51 -894 416 -893
rect 418 -894 1039 -893
rect 82 -896 192 -895
rect 261 -896 580 -895
rect 590 -896 1074 -895
rect 114 -898 356 -897
rect 359 -898 370 -897
rect 394 -898 423 -897
rect 439 -898 1032 -897
rect 1073 -898 1081 -897
rect 114 -900 241 -899
rect 268 -900 300 -899
rect 310 -900 615 -899
rect 635 -900 1004 -899
rect 1010 -900 1039 -899
rect 142 -902 227 -901
rect 240 -902 346 -901
rect 359 -902 752 -901
rect 758 -902 780 -901
rect 891 -902 906 -901
rect 919 -902 927 -901
rect 947 -902 1025 -901
rect 142 -904 213 -903
rect 226 -904 451 -903
rect 562 -904 598 -903
rect 604 -904 1018 -903
rect 149 -906 584 -905
rect 604 -906 619 -905
rect 639 -906 864 -905
rect 898 -906 927 -905
rect 961 -906 1011 -905
rect 156 -908 402 -907
rect 408 -908 430 -907
rect 443 -908 710 -907
rect 723 -908 731 -907
rect 751 -908 829 -907
rect 961 -908 976 -907
rect 996 -908 1004 -907
rect 163 -910 213 -909
rect 254 -910 598 -909
rect 611 -910 661 -909
rect 674 -910 1081 -909
rect 121 -912 255 -911
rect 324 -912 507 -911
rect 534 -912 619 -911
rect 625 -912 675 -911
rect 695 -912 703 -911
rect 716 -912 724 -911
rect 793 -912 1025 -911
rect 2 -914 794 -913
rect 807 -914 829 -913
rect 884 -914 976 -913
rect 100 -916 122 -915
rect 163 -916 416 -915
rect 443 -916 990 -915
rect 65 -918 101 -917
rect 177 -918 206 -917
rect 331 -918 398 -917
rect 408 -918 458 -917
rect 481 -918 640 -917
rect 646 -918 661 -917
rect 716 -918 801 -917
rect 807 -918 836 -917
rect 877 -918 885 -917
rect 289 -920 332 -919
rect 338 -920 528 -919
rect 541 -920 997 -919
rect 107 -922 339 -921
rect 341 -922 423 -921
rect 450 -922 486 -921
rect 506 -922 1060 -921
rect 107 -924 195 -923
rect 289 -924 437 -923
rect 457 -924 689 -923
rect 814 -924 836 -923
rect 849 -924 878 -923
rect 1059 -924 1067 -923
rect 72 -926 1067 -925
rect 345 -928 465 -927
rect 471 -928 815 -927
rect 352 -930 647 -929
rect 688 -930 787 -929
rect 362 -932 402 -931
rect 464 -932 528 -931
rect 541 -932 1046 -931
rect 366 -934 577 -933
rect 593 -934 801 -933
rect 352 -936 594 -935
rect 614 -936 759 -935
rect 366 -938 374 -937
rect 485 -938 559 -937
rect 569 -938 892 -937
rect 177 -940 570 -939
rect 621 -940 1046 -939
rect 369 -942 472 -941
rect 513 -942 850 -941
rect 373 -944 545 -943
rect 625 -944 843 -943
rect 513 -946 521 -945
rect 632 -946 899 -945
rect 23 -948 521 -947
rect 632 -948 1137 -947
rect 23 -950 388 -949
rect 681 -950 843 -949
rect 247 -952 388 -951
rect 667 -952 682 -951
rect 744 -952 787 -951
rect 233 -954 248 -953
rect 667 -954 773 -953
rect 233 -956 297 -955
rect 691 -956 773 -955
rect 737 -958 745 -957
rect 37 -960 738 -959
rect 9 -971 283 -970
rect 285 -971 311 -970
rect 359 -971 727 -970
rect 859 -971 962 -970
rect 9 -973 486 -972
rect 541 -973 1137 -972
rect 16 -975 598 -974
rect 607 -975 906 -974
rect 16 -977 167 -976
rect 194 -977 381 -976
rect 401 -977 465 -976
rect 467 -977 766 -976
rect 23 -979 437 -978
rect 439 -979 689 -978
rect 691 -979 962 -978
rect 23 -981 391 -980
rect 436 -981 559 -980
rect 569 -981 1116 -980
rect 30 -983 34 -982
rect 37 -983 255 -982
rect 271 -983 325 -982
rect 362 -983 629 -982
rect 632 -983 983 -982
rect 30 -985 654 -984
rect 695 -985 829 -984
rect 982 -985 1046 -984
rect 33 -987 654 -986
rect 698 -987 1053 -986
rect 37 -989 45 -988
rect 65 -989 934 -988
rect 1045 -989 1074 -988
rect 44 -991 528 -990
rect 569 -991 927 -990
rect 933 -991 997 -990
rect 1052 -991 1102 -990
rect 2 -993 927 -992
rect 68 -995 416 -994
rect 422 -995 528 -994
rect 576 -995 675 -994
rect 786 -995 1074 -994
rect 68 -997 339 -996
rect 380 -997 514 -996
rect 579 -997 1025 -996
rect 72 -999 87 -998
rect 114 -999 402 -998
rect 415 -999 521 -998
rect 590 -999 668 -998
rect 674 -999 780 -998
rect 786 -999 913 -998
rect 1024 -999 1123 -998
rect 72 -1001 94 -1000
rect 114 -1001 276 -1000
rect 282 -1001 710 -1000
rect 779 -1001 941 -1000
rect 82 -1003 556 -1002
rect 590 -1003 682 -1002
rect 709 -1003 864 -1002
rect 912 -1003 1032 -1002
rect 82 -1005 794 -1004
rect 842 -1005 941 -1004
rect 1010 -1005 1032 -1004
rect 86 -1007 206 -1006
rect 229 -1007 234 -1006
rect 240 -1007 507 -1006
rect 513 -1007 605 -1006
rect 614 -1007 717 -1006
rect 793 -1007 885 -1006
rect 1010 -1007 1042 -1006
rect 93 -1009 108 -1008
rect 135 -1009 419 -1008
rect 443 -1009 451 -1008
rect 471 -1009 682 -1008
rect 716 -1009 822 -1008
rect 842 -1009 899 -1008
rect 58 -1011 822 -1010
rect 863 -1011 969 -1010
rect 58 -1013 76 -1012
rect 107 -1013 122 -1012
rect 135 -1013 227 -1012
rect 233 -1013 430 -1012
rect 450 -1013 703 -1012
rect 884 -1013 976 -1012
rect 121 -1015 164 -1014
rect 191 -1015 423 -1014
rect 471 -1015 489 -1014
rect 492 -1015 507 -1014
rect 520 -1015 545 -1014
rect 548 -1015 703 -1014
rect 898 -1015 1018 -1014
rect 149 -1017 213 -1016
rect 240 -1017 458 -1016
rect 474 -1017 1018 -1016
rect 163 -1019 206 -1018
rect 254 -1019 741 -1018
rect 947 -1019 969 -1018
rect 975 -1019 1039 -1018
rect 191 -1021 297 -1020
rect 303 -1021 549 -1020
rect 555 -1021 808 -1020
rect 856 -1021 948 -1020
rect 177 -1023 304 -1022
rect 306 -1023 584 -1022
rect 593 -1023 1081 -1022
rect 177 -1025 374 -1024
rect 408 -1025 430 -1024
rect 446 -1025 808 -1024
rect 1080 -1025 1095 -1024
rect 268 -1027 325 -1026
rect 331 -1027 374 -1026
rect 408 -1027 493 -1026
rect 502 -1027 997 -1026
rect 142 -1029 269 -1028
rect 275 -1029 395 -1028
rect 457 -1029 738 -1028
rect 51 -1031 395 -1030
rect 478 -1031 1088 -1030
rect 2 -1033 52 -1032
rect 100 -1033 143 -1032
rect 156 -1033 479 -1032
rect 481 -1033 815 -1032
rect 156 -1035 248 -1034
rect 289 -1035 332 -1034
rect 338 -1035 398 -1034
rect 583 -1035 892 -1034
rect 247 -1037 318 -1036
rect 600 -1037 766 -1036
rect 891 -1037 1004 -1036
rect 289 -1039 346 -1038
rect 618 -1039 829 -1038
rect 1003 -1039 1067 -1038
rect 261 -1041 346 -1040
rect 562 -1041 619 -1040
rect 621 -1041 871 -1040
rect 919 -1041 1067 -1040
rect 261 -1043 353 -1042
rect 499 -1043 920 -1042
rect 310 -1045 388 -1044
rect 562 -1045 573 -1044
rect 635 -1045 752 -1044
rect 870 -1045 990 -1044
rect 317 -1047 535 -1046
rect 572 -1047 906 -1046
rect 989 -1047 1109 -1046
rect 352 -1049 367 -1048
rect 387 -1049 640 -1048
rect 667 -1049 773 -1048
rect 128 -1051 367 -1050
rect 495 -1051 640 -1050
rect 737 -1051 1130 -1050
rect 128 -1053 171 -1052
rect 534 -1053 647 -1052
rect 751 -1053 836 -1052
rect 1129 -1053 1158 -1052
rect 170 -1055 199 -1054
rect 611 -1055 647 -1054
rect 800 -1055 836 -1054
rect 198 -1057 850 -1056
rect 611 -1059 724 -1058
rect 744 -1059 801 -1058
rect 849 -1059 955 -1058
rect 625 -1061 773 -1060
rect 954 -1061 1060 -1060
rect 502 -1063 626 -1062
rect 635 -1063 857 -1062
rect 723 -1065 1144 -1064
rect 730 -1067 745 -1066
rect 1143 -1067 1151 -1066
rect 660 -1069 731 -1068
rect 660 -1071 759 -1070
rect 758 -1073 878 -1072
rect 604 -1075 878 -1074
rect 5 -1086 349 -1085
rect 366 -1086 370 -1085
rect 390 -1086 899 -1085
rect 947 -1086 1039 -1085
rect 1041 -1086 1067 -1085
rect 1076 -1086 1081 -1085
rect 1122 -1086 1130 -1085
rect 1143 -1086 1151 -1085
rect 9 -1088 468 -1087
rect 488 -1088 521 -1087
rect 523 -1088 829 -1087
rect 905 -1088 948 -1087
rect 996 -1088 1060 -1087
rect 9 -1090 31 -1089
rect 40 -1090 899 -1089
rect 982 -1090 997 -1089
rect 1031 -1090 1067 -1089
rect 16 -1092 496 -1091
rect 513 -1092 692 -1091
rect 723 -1092 752 -1091
rect 779 -1092 829 -1091
rect 856 -1092 906 -1091
rect 926 -1092 983 -1091
rect 1017 -1092 1032 -1091
rect 51 -1094 59 -1093
rect 61 -1094 199 -1093
rect 212 -1094 801 -1093
rect 817 -1094 955 -1093
rect 1010 -1094 1018 -1093
rect 51 -1096 276 -1095
rect 324 -1096 409 -1095
rect 418 -1096 990 -1095
rect 1003 -1096 1011 -1095
rect 65 -1098 157 -1097
rect 166 -1098 703 -1097
rect 740 -1098 780 -1097
rect 789 -1098 864 -1097
rect 926 -1098 934 -1097
rect 940 -1098 1004 -1097
rect 65 -1100 73 -1099
rect 79 -1100 206 -1099
rect 212 -1100 220 -1099
rect 268 -1100 332 -1099
rect 366 -1100 395 -1099
rect 397 -1100 444 -1099
rect 450 -1100 514 -1099
rect 527 -1100 636 -1099
rect 639 -1100 703 -1099
rect 751 -1100 815 -1099
rect 835 -1100 857 -1099
rect 870 -1100 941 -1099
rect 975 -1100 990 -1099
rect 68 -1102 503 -1101
rect 541 -1102 955 -1101
rect 79 -1104 94 -1103
rect 100 -1104 108 -1103
rect 114 -1104 199 -1103
rect 205 -1104 262 -1103
rect 324 -1104 1039 -1103
rect 93 -1106 286 -1105
rect 331 -1106 353 -1105
rect 369 -1106 395 -1105
rect 401 -1106 521 -1105
rect 544 -1106 822 -1105
rect 835 -1106 843 -1105
rect 884 -1106 934 -1105
rect 72 -1108 353 -1107
rect 355 -1108 822 -1107
rect 842 -1108 1042 -1107
rect 100 -1110 143 -1109
rect 149 -1110 157 -1109
rect 170 -1110 220 -1109
rect 254 -1110 402 -1109
rect 415 -1110 444 -1109
rect 450 -1110 738 -1109
rect 765 -1110 801 -1109
rect 919 -1110 976 -1109
rect 23 -1112 171 -1111
rect 177 -1112 412 -1111
rect 422 -1112 528 -1111
rect 555 -1112 745 -1111
rect 765 -1112 1074 -1111
rect 23 -1114 38 -1113
rect 103 -1114 689 -1113
rect 744 -1114 759 -1113
rect 772 -1114 885 -1113
rect 891 -1114 920 -1113
rect 114 -1116 129 -1115
rect 152 -1116 314 -1115
rect 383 -1116 1060 -1115
rect 177 -1118 304 -1117
rect 436 -1118 542 -1117
rect 555 -1118 1025 -1117
rect 184 -1120 262 -1119
rect 296 -1120 423 -1119
rect 492 -1120 734 -1119
rect 891 -1120 913 -1119
rect 121 -1122 297 -1121
rect 303 -1122 346 -1121
rect 380 -1122 437 -1121
rect 499 -1122 864 -1121
rect 877 -1122 913 -1121
rect 30 -1124 346 -1123
rect 373 -1124 381 -1123
rect 499 -1124 1074 -1123
rect 44 -1126 374 -1125
rect 502 -1126 787 -1125
rect 44 -1128 573 -1127
rect 576 -1128 598 -1127
rect 607 -1128 619 -1127
rect 632 -1128 759 -1127
rect 110 -1130 878 -1129
rect 121 -1132 290 -1131
rect 387 -1132 633 -1131
rect 639 -1132 710 -1131
rect 163 -1134 290 -1133
rect 481 -1134 787 -1133
rect 184 -1136 409 -1135
rect 565 -1136 815 -1135
rect 191 -1138 276 -1137
rect 569 -1138 612 -1137
rect 618 -1138 647 -1137
rect 653 -1138 773 -1137
rect 86 -1140 192 -1139
rect 215 -1140 486 -1139
rect 558 -1140 647 -1139
rect 684 -1140 962 -1139
rect 86 -1142 318 -1141
rect 415 -1142 612 -1141
rect 709 -1142 717 -1141
rect 849 -1142 962 -1141
rect 54 -1144 717 -1143
rect 807 -1144 850 -1143
rect 128 -1146 559 -1145
rect 583 -1146 682 -1145
rect 226 -1148 388 -1147
rect 471 -1148 682 -1147
rect 135 -1150 227 -1149
rect 240 -1150 577 -1149
rect 586 -1150 871 -1149
rect 135 -1152 535 -1151
rect 562 -1152 584 -1151
rect 604 -1152 654 -1151
rect 240 -1154 339 -1153
rect 457 -1154 472 -1153
rect 478 -1154 486 -1153
rect 534 -1154 696 -1153
rect 247 -1156 255 -1155
rect 310 -1156 339 -1155
rect 359 -1156 458 -1155
rect 548 -1156 605 -1155
rect 625 -1156 808 -1155
rect 233 -1158 248 -1157
rect 317 -1158 465 -1157
rect 548 -1158 661 -1157
rect 674 -1158 696 -1157
rect 37 -1160 234 -1159
rect 282 -1160 675 -1159
rect 464 -1162 626 -1161
rect 660 -1162 731 -1161
rect 730 -1164 1025 -1163
rect 2 -1175 146 -1174
rect 149 -1175 206 -1174
rect 226 -1175 311 -1174
rect 313 -1175 822 -1174
rect 982 -1175 1074 -1174
rect 1115 -1175 1123 -1174
rect 1129 -1175 1158 -1174
rect 16 -1177 276 -1176
rect 303 -1177 409 -1176
rect 460 -1177 472 -1176
rect 485 -1177 489 -1176
rect 506 -1177 521 -1176
rect 558 -1177 696 -1176
rect 730 -1177 934 -1176
rect 989 -1177 1081 -1176
rect 1150 -1177 1165 -1176
rect 16 -1179 381 -1178
rect 383 -1179 479 -1178
rect 485 -1179 605 -1178
rect 653 -1179 731 -1178
rect 751 -1179 857 -1178
rect 863 -1179 934 -1178
rect 996 -1179 1088 -1178
rect 19 -1181 248 -1180
rect 310 -1181 318 -1180
rect 331 -1181 356 -1180
rect 359 -1181 822 -1180
rect 912 -1181 990 -1180
rect 1003 -1181 1095 -1180
rect 23 -1183 38 -1182
rect 58 -1183 941 -1182
rect 947 -1183 1004 -1182
rect 1017 -1183 1109 -1182
rect 23 -1185 363 -1184
rect 380 -1185 402 -1184
rect 443 -1185 472 -1184
rect 478 -1185 538 -1184
rect 562 -1185 808 -1184
rect 877 -1185 941 -1184
rect 1031 -1185 1144 -1184
rect 37 -1187 353 -1186
rect 366 -1187 402 -1186
rect 429 -1187 444 -1186
rect 464 -1187 668 -1186
rect 681 -1187 752 -1186
rect 758 -1187 808 -1186
rect 884 -1187 948 -1186
rect 1041 -1187 1067 -1186
rect 44 -1189 367 -1188
rect 394 -1189 419 -1188
rect 429 -1189 643 -1188
rect 656 -1189 1137 -1188
rect 44 -1191 66 -1190
rect 96 -1191 528 -1190
rect 534 -1191 759 -1190
rect 786 -1191 969 -1190
rect 1045 -1191 1102 -1190
rect 58 -1193 129 -1192
rect 135 -1193 482 -1192
rect 506 -1193 1025 -1192
rect 1052 -1193 1123 -1192
rect 61 -1195 136 -1194
rect 142 -1195 416 -1194
rect 513 -1195 605 -1194
rect 681 -1195 962 -1194
rect 1059 -1195 1151 -1194
rect 65 -1197 195 -1196
rect 198 -1197 286 -1196
rect 289 -1197 353 -1196
rect 394 -1197 556 -1196
rect 562 -1197 577 -1196
rect 597 -1197 661 -1196
rect 688 -1197 1025 -1196
rect 100 -1199 108 -1198
rect 121 -1199 360 -1198
rect 415 -1199 503 -1198
rect 523 -1199 1067 -1198
rect 100 -1201 115 -1200
rect 121 -1201 612 -1200
rect 688 -1201 717 -1200
rect 733 -1201 864 -1200
rect 891 -1201 1018 -1200
rect 79 -1203 115 -1202
rect 128 -1203 178 -1202
rect 184 -1203 206 -1202
rect 222 -1203 276 -1202
rect 296 -1203 332 -1202
rect 345 -1203 773 -1202
rect 786 -1203 1011 -1202
rect 79 -1205 451 -1204
rect 488 -1205 514 -1204
rect 527 -1205 633 -1204
rect 695 -1205 766 -1204
rect 789 -1205 1032 -1204
rect 107 -1207 325 -1206
rect 345 -1207 374 -1206
rect 422 -1207 773 -1206
rect 859 -1207 1053 -1206
rect 72 -1209 325 -1208
rect 373 -1209 815 -1208
rect 905 -1209 962 -1208
rect 975 -1209 1060 -1208
rect 142 -1211 370 -1210
rect 422 -1211 493 -1210
rect 555 -1211 1119 -1210
rect 152 -1213 465 -1212
rect 569 -1213 612 -1212
rect 702 -1213 892 -1212
rect 898 -1213 976 -1212
rect 93 -1215 703 -1214
rect 716 -1215 878 -1214
rect 919 -1215 997 -1214
rect 156 -1217 220 -1216
rect 233 -1217 885 -1216
rect 926 -1217 1011 -1216
rect 86 -1219 234 -1218
rect 240 -1219 297 -1218
rect 436 -1219 451 -1218
rect 467 -1219 570 -1218
rect 576 -1219 591 -1218
rect 670 -1219 920 -1218
rect 954 -1219 1046 -1218
rect 51 -1221 437 -1220
rect 583 -1221 591 -1220
rect 719 -1221 955 -1220
rect 51 -1223 269 -1222
rect 723 -1223 766 -1222
rect 828 -1223 899 -1222
rect 86 -1225 171 -1224
rect 177 -1225 388 -1224
rect 646 -1225 724 -1224
rect 737 -1225 913 -1224
rect 9 -1227 171 -1226
rect 184 -1227 262 -1226
rect 268 -1227 283 -1226
rect 387 -1227 626 -1226
rect 744 -1227 815 -1226
rect 849 -1227 927 -1226
rect 9 -1229 31 -1228
rect 93 -1229 584 -1228
rect 618 -1229 647 -1228
rect 709 -1229 745 -1228
rect 779 -1229 850 -1228
rect 870 -1229 906 -1228
rect 30 -1231 290 -1230
rect 492 -1231 738 -1230
rect 779 -1231 794 -1230
rect 800 -1231 871 -1230
rect 159 -1233 601 -1232
rect 625 -1233 668 -1232
rect 674 -1233 710 -1232
rect 800 -1233 1039 -1232
rect 163 -1235 983 -1234
rect 163 -1237 213 -1236
rect 240 -1237 349 -1236
rect 541 -1237 619 -1236
rect 639 -1237 794 -1236
rect 968 -1237 1039 -1236
rect 191 -1239 227 -1238
rect 247 -1239 304 -1238
rect 509 -1239 542 -1238
rect 548 -1239 675 -1238
rect 201 -1241 318 -1240
rect 499 -1241 549 -1240
rect 600 -1241 843 -1240
rect 212 -1243 272 -1242
rect 282 -1243 339 -1242
rect 457 -1243 500 -1242
rect 705 -1243 843 -1242
rect 254 -1245 262 -1244
rect 338 -1245 685 -1244
rect 254 -1247 377 -1246
rect 457 -1247 661 -1246
rect 2 -1258 73 -1257
rect 159 -1258 388 -1257
rect 404 -1258 528 -1257
rect 534 -1258 619 -1257
rect 632 -1258 815 -1257
rect 821 -1258 1133 -1257
rect 1164 -1258 1172 -1257
rect 2 -1260 52 -1259
rect 72 -1260 269 -1259
rect 282 -1260 304 -1259
rect 317 -1260 440 -1259
rect 443 -1260 447 -1259
rect 485 -1260 703 -1259
rect 705 -1260 1018 -1259
rect 1024 -1260 1028 -1259
rect 1122 -1260 1130 -1259
rect 1157 -1260 1165 -1259
rect 44 -1262 216 -1261
rect 233 -1262 293 -1261
rect 303 -1262 556 -1261
rect 572 -1262 871 -1261
rect 968 -1262 1102 -1261
rect 1122 -1262 1144 -1261
rect 33 -1264 45 -1263
rect 51 -1264 171 -1263
rect 191 -1264 1074 -1263
rect 1143 -1264 1151 -1263
rect 47 -1266 1074 -1265
rect 142 -1268 815 -1267
rect 828 -1268 878 -1267
rect 968 -1268 983 -1267
rect 1024 -1268 1039 -1267
rect 1052 -1268 1102 -1267
rect 142 -1270 213 -1269
rect 233 -1270 297 -1269
rect 317 -1270 412 -1269
rect 443 -1270 465 -1269
rect 471 -1270 486 -1269
rect 492 -1270 605 -1269
rect 618 -1270 675 -1269
rect 684 -1270 962 -1269
rect 9 -1272 213 -1271
rect 240 -1272 370 -1271
rect 408 -1272 507 -1271
rect 523 -1272 899 -1271
rect 905 -1272 962 -1271
rect 9 -1274 255 -1273
rect 261 -1274 272 -1273
rect 282 -1274 661 -1273
rect 667 -1274 990 -1273
rect 16 -1276 605 -1275
rect 632 -1276 752 -1275
rect 786 -1276 808 -1275
rect 828 -1276 1011 -1275
rect 16 -1278 181 -1277
rect 191 -1278 206 -1277
rect 261 -1278 538 -1277
rect 555 -1278 563 -1277
rect 569 -1278 983 -1277
rect 1010 -1278 1081 -1277
rect 114 -1280 241 -1279
rect 268 -1280 339 -1279
rect 359 -1280 388 -1279
rect 436 -1280 808 -1279
rect 831 -1280 1088 -1279
rect 58 -1282 360 -1281
rect 450 -1282 465 -1281
rect 471 -1282 514 -1281
rect 534 -1282 738 -1281
rect 751 -1282 850 -1281
rect 877 -1282 892 -1281
rect 1066 -1282 1088 -1281
rect 58 -1284 195 -1283
rect 205 -1284 248 -1283
rect 289 -1284 374 -1283
rect 457 -1284 1053 -1283
rect 86 -1286 115 -1285
rect 135 -1286 290 -1285
rect 296 -1286 430 -1285
rect 457 -1286 563 -1285
rect 576 -1286 598 -1285
rect 600 -1286 913 -1285
rect 1027 -1286 1039 -1285
rect 1045 -1286 1067 -1285
rect 86 -1288 101 -1287
rect 107 -1288 136 -1287
rect 156 -1288 871 -1287
rect 891 -1288 948 -1287
rect 1003 -1288 1046 -1287
rect 26 -1290 157 -1289
rect 163 -1290 255 -1289
rect 275 -1290 430 -1289
rect 478 -1290 738 -1289
rect 796 -1290 857 -1289
rect 912 -1290 934 -1289
rect 947 -1290 990 -1289
rect 1003 -1290 1032 -1289
rect 37 -1292 276 -1291
rect 324 -1292 570 -1291
rect 590 -1292 675 -1291
rect 688 -1292 822 -1291
rect 835 -1292 906 -1291
rect 933 -1292 955 -1291
rect 1031 -1292 1137 -1291
rect 37 -1294 185 -1293
rect 247 -1294 395 -1293
rect 408 -1294 577 -1293
rect 607 -1294 1081 -1293
rect 1136 -1294 1158 -1293
rect 100 -1296 311 -1295
rect 324 -1296 423 -1295
rect 495 -1296 689 -1295
rect 716 -1296 1116 -1295
rect 107 -1298 129 -1297
rect 170 -1298 636 -1297
rect 639 -1298 1018 -1297
rect 1108 -1298 1116 -1297
rect 30 -1300 129 -1299
rect 184 -1300 188 -1299
rect 310 -1300 416 -1299
rect 499 -1300 528 -1299
rect 541 -1300 591 -1299
rect 621 -1300 832 -1299
rect 849 -1300 976 -1299
rect 1094 -1300 1109 -1299
rect 65 -1302 416 -1301
rect 513 -1302 521 -1301
rect 642 -1302 1060 -1301
rect 121 -1304 640 -1303
rect 646 -1304 668 -1303
rect 670 -1304 766 -1303
rect 779 -1304 836 -1303
rect 842 -1304 1095 -1303
rect 79 -1306 122 -1305
rect 338 -1306 629 -1305
rect 646 -1306 759 -1305
rect 772 -1306 780 -1305
rect 800 -1306 899 -1305
rect 940 -1306 955 -1305
rect 975 -1306 997 -1305
rect 79 -1308 97 -1307
rect 345 -1308 500 -1307
rect 506 -1308 773 -1307
rect 842 -1308 864 -1307
rect 198 -1310 346 -1309
rect 348 -1310 1060 -1309
rect 177 -1312 199 -1311
rect 352 -1312 423 -1311
rect 436 -1312 941 -1311
rect 352 -1314 381 -1313
rect 394 -1314 542 -1313
rect 597 -1314 997 -1313
rect 366 -1316 766 -1315
rect 856 -1316 920 -1315
rect 23 -1318 920 -1317
rect 331 -1320 367 -1319
rect 380 -1320 402 -1319
rect 520 -1320 661 -1319
rect 709 -1320 801 -1319
rect 149 -1322 332 -1321
rect 401 -1322 461 -1321
rect 625 -1322 710 -1321
rect 723 -1322 864 -1321
rect 149 -1324 682 -1323
rect 695 -1324 724 -1323
rect 733 -1324 885 -1323
rect 103 -1326 696 -1325
rect 744 -1326 759 -1325
rect 884 -1326 927 -1325
rect 460 -1328 510 -1327
rect 544 -1328 927 -1327
rect 653 -1330 790 -1329
rect 492 -1332 654 -1331
rect 656 -1332 794 -1331
rect 548 -1334 794 -1333
rect 548 -1336 584 -1335
rect 730 -1336 745 -1335
rect 583 -1338 612 -1337
rect 478 -1340 612 -1339
rect 2 -1351 433 -1350
rect 436 -1351 689 -1350
rect 733 -1351 1046 -1350
rect 1101 -1351 1151 -1350
rect 1153 -1351 1165 -1350
rect 2 -1353 122 -1352
rect 135 -1353 335 -1352
rect 359 -1353 524 -1352
rect 527 -1353 948 -1352
rect 950 -1353 1130 -1352
rect 1136 -1353 1172 -1352
rect 9 -1355 164 -1354
rect 215 -1355 416 -1354
rect 506 -1355 542 -1354
rect 544 -1355 647 -1354
rect 688 -1355 976 -1354
rect 996 -1355 1067 -1354
rect 16 -1357 412 -1356
rect 506 -1357 633 -1356
rect 681 -1357 976 -1356
rect 1031 -1357 1067 -1356
rect 23 -1359 447 -1358
rect 520 -1359 843 -1358
rect 1031 -1359 1095 -1358
rect 26 -1361 241 -1360
rect 275 -1361 528 -1360
rect 537 -1361 899 -1360
rect 1045 -1361 1144 -1360
rect 33 -1363 59 -1362
rect 65 -1363 486 -1362
rect 562 -1363 647 -1362
rect 681 -1363 752 -1362
rect 772 -1363 906 -1362
rect 44 -1365 69 -1364
rect 93 -1365 108 -1364
rect 121 -1365 1081 -1364
rect 44 -1367 87 -1366
rect 100 -1367 206 -1366
rect 212 -1367 1095 -1366
rect 16 -1369 101 -1368
rect 103 -1369 276 -1368
rect 289 -1369 423 -1368
rect 485 -1369 675 -1368
rect 751 -1369 759 -1368
rect 772 -1369 836 -1368
rect 842 -1369 857 -1368
rect 898 -1369 1025 -1368
rect 51 -1371 461 -1370
rect 492 -1371 1081 -1370
rect 51 -1373 353 -1372
rect 359 -1373 381 -1372
rect 387 -1373 906 -1372
rect 58 -1375 248 -1374
rect 268 -1375 381 -1374
rect 387 -1375 500 -1374
rect 600 -1375 1053 -1374
rect 65 -1377 115 -1376
rect 128 -1377 241 -1376
rect 247 -1377 297 -1376
rect 303 -1377 496 -1376
rect 569 -1377 1053 -1376
rect 37 -1379 129 -1378
rect 135 -1379 332 -1378
rect 408 -1379 451 -1378
rect 611 -1379 969 -1378
rect 37 -1381 325 -1380
rect 331 -1381 416 -1380
rect 422 -1381 570 -1380
rect 611 -1381 696 -1380
rect 758 -1381 822 -1380
rect 828 -1381 1109 -1380
rect 72 -1383 87 -1382
rect 103 -1383 178 -1382
rect 187 -1383 409 -1382
rect 443 -1383 451 -1382
rect 509 -1383 969 -1382
rect 1108 -1383 1158 -1382
rect 72 -1385 556 -1384
rect 614 -1385 815 -1384
rect 821 -1385 878 -1384
rect 79 -1387 556 -1386
rect 625 -1387 955 -1386
rect 79 -1389 199 -1388
rect 226 -1389 349 -1388
rect 618 -1389 626 -1388
rect 632 -1389 654 -1388
rect 660 -1389 836 -1388
rect 849 -1389 955 -1388
rect 110 -1391 1025 -1390
rect 149 -1393 405 -1392
rect 653 -1393 808 -1392
rect 814 -1393 1063 -1392
rect 149 -1395 318 -1394
rect 324 -1395 430 -1394
rect 660 -1395 668 -1394
rect 674 -1395 717 -1394
rect 775 -1395 787 -1394
rect 828 -1395 934 -1394
rect 156 -1397 731 -1396
rect 786 -1397 871 -1396
rect 877 -1397 913 -1396
rect 933 -1397 1088 -1396
rect 156 -1399 262 -1398
rect 282 -1399 668 -1398
rect 695 -1399 724 -1398
rect 856 -1399 1060 -1398
rect 163 -1401 185 -1400
rect 191 -1401 206 -1400
rect 219 -1401 283 -1400
rect 292 -1401 496 -1400
rect 716 -1401 766 -1400
rect 870 -1401 885 -1400
rect 912 -1401 1011 -1400
rect 177 -1403 353 -1402
rect 534 -1403 885 -1402
rect 926 -1403 1088 -1402
rect 194 -1405 269 -1404
rect 296 -1405 503 -1404
rect 723 -1405 738 -1404
rect 765 -1405 780 -1404
rect 891 -1405 927 -1404
rect 961 -1405 1011 -1404
rect 198 -1407 605 -1406
rect 737 -1407 745 -1406
rect 779 -1407 801 -1406
rect 961 -1407 983 -1406
rect 30 -1409 801 -1408
rect 982 -1409 990 -1408
rect 30 -1411 143 -1410
rect 219 -1411 234 -1410
rect 254 -1411 262 -1410
rect 310 -1411 440 -1410
rect 471 -1411 535 -1410
rect 604 -1411 710 -1410
rect 793 -1411 892 -1410
rect 989 -1411 1004 -1410
rect 93 -1413 745 -1412
rect 1003 -1413 1074 -1412
rect 142 -1415 171 -1414
rect 226 -1415 458 -1414
rect 464 -1415 472 -1414
rect 639 -1415 710 -1414
rect 1073 -1415 1123 -1414
rect 96 -1417 171 -1416
rect 233 -1417 402 -1416
rect 457 -1417 692 -1416
rect 702 -1417 794 -1416
rect 254 -1419 850 -1418
rect 303 -1421 440 -1420
rect 464 -1421 577 -1420
rect 702 -1421 808 -1420
rect 310 -1423 598 -1422
rect 317 -1425 580 -1424
rect 338 -1427 619 -1426
rect 338 -1429 489 -1428
rect 499 -1429 640 -1428
rect 401 -1431 563 -1430
rect 576 -1431 864 -1430
rect 345 -1433 864 -1432
rect 345 -1435 479 -1434
rect 478 -1437 591 -1436
rect 583 -1439 591 -1438
rect 548 -1441 584 -1440
rect 548 -1443 1018 -1442
rect 1017 -1445 1039 -1444
rect 1038 -1447 1116 -1446
rect 9 -1458 468 -1457
rect 481 -1458 605 -1457
rect 611 -1458 997 -1457
rect 1010 -1458 1060 -1457
rect 16 -1460 496 -1459
rect 499 -1460 948 -1459
rect 996 -1460 1074 -1459
rect 16 -1462 332 -1461
rect 352 -1462 524 -1461
rect 551 -1462 675 -1461
rect 681 -1462 703 -1461
rect 744 -1462 1046 -1461
rect 1062 -1462 1074 -1461
rect 30 -1464 188 -1463
rect 198 -1464 549 -1463
rect 569 -1464 661 -1463
rect 681 -1464 766 -1463
rect 856 -1464 913 -1463
rect 947 -1464 1032 -1463
rect 23 -1466 199 -1465
rect 257 -1466 262 -1465
rect 289 -1466 412 -1465
rect 415 -1466 430 -1465
rect 436 -1466 507 -1465
rect 516 -1466 759 -1465
rect 765 -1466 836 -1465
rect 856 -1466 962 -1465
rect 1017 -1466 1021 -1465
rect 23 -1468 255 -1467
rect 292 -1468 360 -1467
rect 387 -1468 500 -1467
rect 502 -1468 696 -1467
rect 747 -1468 878 -1467
rect 884 -1468 1011 -1467
rect 1017 -1468 1039 -1467
rect 33 -1470 717 -1469
rect 758 -1470 787 -1469
rect 835 -1470 955 -1469
rect 1020 -1470 1039 -1469
rect 44 -1472 111 -1471
rect 114 -1472 269 -1471
rect 310 -1472 510 -1471
rect 541 -1472 549 -1471
rect 569 -1472 664 -1471
rect 695 -1472 920 -1471
rect 933 -1472 962 -1471
rect 30 -1474 45 -1473
rect 51 -1474 216 -1473
rect 254 -1474 297 -1473
rect 310 -1474 328 -1473
rect 331 -1474 374 -1473
rect 387 -1474 479 -1473
rect 485 -1474 668 -1473
rect 730 -1474 920 -1473
rect 954 -1474 1095 -1473
rect 2 -1476 216 -1475
rect 296 -1476 514 -1475
rect 541 -1476 640 -1475
rect 730 -1476 752 -1475
rect 786 -1476 892 -1475
rect 912 -1476 990 -1475
rect 1094 -1476 1109 -1475
rect 2 -1478 97 -1477
rect 103 -1478 675 -1477
rect 688 -1478 990 -1477
rect 51 -1480 325 -1479
rect 345 -1480 416 -1479
rect 422 -1480 507 -1479
rect 576 -1480 822 -1479
rect 859 -1480 934 -1479
rect 37 -1482 325 -1481
rect 373 -1482 381 -1481
rect 394 -1482 405 -1481
rect 408 -1482 745 -1481
rect 821 -1482 906 -1481
rect 9 -1484 38 -1483
rect 65 -1484 192 -1483
rect 233 -1484 752 -1483
rect 863 -1484 1046 -1483
rect 58 -1486 192 -1485
rect 226 -1486 234 -1485
rect 366 -1486 381 -1485
rect 401 -1486 615 -1485
rect 639 -1486 710 -1485
rect 807 -1486 864 -1485
rect 870 -1486 892 -1485
rect 58 -1488 143 -1487
rect 163 -1488 181 -1487
rect 226 -1488 290 -1487
rect 422 -1488 671 -1487
rect 807 -1488 941 -1487
rect 65 -1490 451 -1489
rect 464 -1490 612 -1489
rect 870 -1490 969 -1489
rect 72 -1492 269 -1491
rect 432 -1492 717 -1491
rect 877 -1492 983 -1491
rect 72 -1494 220 -1493
rect 439 -1494 815 -1493
rect 884 -1494 899 -1493
rect 940 -1494 1025 -1493
rect 79 -1496 335 -1495
rect 443 -1496 472 -1495
rect 485 -1496 794 -1495
rect 814 -1496 829 -1495
rect 968 -1496 1004 -1495
rect 1024 -1496 1081 -1495
rect 79 -1498 248 -1497
rect 443 -1498 563 -1497
rect 590 -1498 605 -1497
rect 793 -1498 850 -1497
rect 982 -1498 1053 -1497
rect 86 -1500 146 -1499
rect 163 -1500 521 -1499
rect 534 -1500 591 -1499
rect 597 -1500 647 -1499
rect 779 -1500 850 -1499
rect 1003 -1500 1067 -1499
rect 86 -1502 150 -1501
rect 166 -1502 633 -1501
rect 646 -1502 738 -1501
rect 772 -1502 780 -1501
rect 828 -1502 843 -1501
rect 107 -1504 171 -1503
rect 177 -1504 493 -1503
rect 534 -1504 710 -1503
rect 842 -1504 927 -1503
rect 93 -1506 108 -1505
rect 114 -1506 692 -1505
rect 705 -1506 927 -1505
rect 93 -1508 601 -1507
rect 677 -1508 738 -1507
rect 121 -1510 580 -1509
rect 691 -1510 801 -1509
rect 124 -1512 241 -1511
rect 247 -1512 619 -1511
rect 800 -1512 976 -1511
rect 128 -1514 262 -1513
rect 366 -1514 563 -1513
rect 618 -1514 724 -1513
rect 128 -1516 185 -1515
rect 212 -1516 976 -1515
rect 100 -1518 213 -1517
rect 219 -1518 409 -1517
rect 450 -1518 538 -1517
rect 555 -1518 906 -1517
rect 135 -1520 353 -1519
rect 359 -1520 724 -1519
rect 135 -1522 339 -1521
rect 457 -1522 633 -1521
rect 149 -1524 626 -1523
rect 156 -1526 171 -1525
rect 177 -1526 395 -1525
rect 457 -1526 577 -1525
rect 625 -1526 654 -1525
rect 156 -1528 899 -1527
rect 184 -1530 206 -1529
rect 240 -1530 318 -1529
rect 338 -1530 1032 -1529
rect 194 -1532 654 -1531
rect 205 -1534 346 -1533
rect 527 -1534 556 -1533
rect 275 -1536 318 -1535
rect 527 -1536 584 -1535
rect 513 -1538 584 -1537
rect 2 -1549 248 -1548
rect 254 -1549 290 -1548
rect 352 -1549 360 -1548
rect 376 -1549 437 -1548
rect 457 -1549 920 -1548
rect 940 -1549 1011 -1548
rect 1034 -1549 1039 -1548
rect 1045 -1549 1102 -1548
rect 5 -1551 101 -1550
rect 145 -1551 1053 -1550
rect 1059 -1551 1109 -1550
rect 9 -1553 251 -1552
rect 261 -1553 437 -1552
rect 464 -1553 696 -1552
rect 772 -1553 892 -1552
rect 975 -1553 1046 -1552
rect 1094 -1553 1116 -1552
rect 9 -1555 486 -1554
rect 513 -1555 671 -1554
rect 674 -1555 1018 -1554
rect 1073 -1555 1095 -1554
rect 30 -1557 150 -1556
rect 156 -1557 185 -1556
rect 198 -1557 262 -1556
rect 268 -1557 535 -1556
rect 562 -1557 906 -1556
rect 926 -1557 1018 -1556
rect 33 -1559 41 -1558
rect 51 -1559 461 -1558
rect 471 -1559 752 -1558
rect 821 -1559 892 -1558
rect 989 -1559 1074 -1558
rect 37 -1561 654 -1560
rect 660 -1561 759 -1560
rect 821 -1561 1070 -1560
rect 37 -1563 45 -1562
rect 51 -1563 426 -1562
rect 478 -1563 500 -1562
rect 520 -1563 619 -1562
rect 625 -1563 773 -1562
rect 835 -1563 927 -1562
rect 961 -1563 990 -1562
rect 996 -1563 1081 -1562
rect 65 -1565 500 -1564
rect 534 -1565 899 -1564
rect 16 -1567 66 -1566
rect 72 -1567 521 -1566
rect 565 -1567 1025 -1566
rect 16 -1569 223 -1568
rect 268 -1569 339 -1568
rect 359 -1569 678 -1568
rect 716 -1569 752 -1568
rect 814 -1569 899 -1568
rect 982 -1569 1025 -1568
rect 72 -1571 87 -1570
rect 93 -1571 570 -1570
rect 576 -1571 689 -1570
rect 716 -1571 745 -1570
rect 765 -1571 815 -1570
rect 859 -1571 1004 -1570
rect 79 -1573 150 -1572
rect 163 -1573 472 -1572
rect 478 -1573 675 -1572
rect 684 -1573 745 -1572
rect 765 -1573 864 -1572
rect 870 -1573 920 -1572
rect 933 -1573 1004 -1572
rect 79 -1575 276 -1574
rect 282 -1575 293 -1574
rect 345 -1575 864 -1574
rect 884 -1575 976 -1574
rect 86 -1577 115 -1576
rect 121 -1577 157 -1576
rect 163 -1577 451 -1576
rect 464 -1577 619 -1576
rect 625 -1577 1039 -1576
rect 96 -1579 517 -1578
rect 527 -1579 577 -1578
rect 590 -1579 962 -1578
rect 968 -1579 983 -1578
rect 100 -1581 108 -1580
rect 121 -1581 136 -1580
rect 166 -1581 486 -1580
rect 506 -1581 528 -1580
rect 583 -1581 591 -1580
rect 593 -1581 703 -1580
rect 723 -1581 836 -1580
rect 912 -1581 969 -1580
rect 107 -1583 311 -1582
rect 331 -1583 451 -1582
rect 597 -1583 1088 -1582
rect 128 -1585 146 -1584
rect 177 -1585 402 -1584
rect 597 -1585 605 -1584
rect 611 -1585 678 -1584
rect 723 -1585 731 -1584
rect 793 -1585 871 -1584
rect 114 -1587 612 -1586
rect 614 -1587 941 -1586
rect 128 -1589 353 -1588
rect 366 -1589 402 -1588
rect 429 -1589 605 -1588
rect 632 -1589 906 -1588
rect 180 -1591 423 -1590
rect 457 -1591 794 -1590
rect 800 -1591 934 -1590
rect 201 -1593 682 -1592
rect 730 -1593 850 -1592
rect 205 -1595 209 -1594
rect 212 -1595 230 -1594
rect 233 -1595 507 -1594
rect 635 -1595 703 -1594
rect 800 -1595 1063 -1594
rect 191 -1597 213 -1596
rect 219 -1597 255 -1596
rect 278 -1597 850 -1596
rect 58 -1599 192 -1598
rect 226 -1599 346 -1598
rect 366 -1599 468 -1598
rect 639 -1599 654 -1598
rect 663 -1599 808 -1598
rect 828 -1599 885 -1598
rect 44 -1601 227 -1600
rect 233 -1601 388 -1600
rect 394 -1601 563 -1600
rect 639 -1601 1032 -1600
rect 58 -1603 696 -1602
rect 737 -1603 808 -1602
rect 947 -1603 1032 -1602
rect 240 -1605 332 -1604
rect 355 -1605 395 -1604
rect 408 -1605 430 -1604
rect 646 -1605 913 -1604
rect 947 -1605 955 -1604
rect 240 -1607 318 -1606
rect 324 -1607 633 -1606
rect 667 -1607 780 -1606
rect 877 -1607 955 -1606
rect 282 -1609 587 -1608
rect 709 -1609 878 -1608
rect 303 -1611 318 -1610
rect 373 -1611 388 -1610
rect 408 -1611 416 -1610
rect 492 -1611 647 -1610
rect 737 -1611 787 -1610
rect 23 -1613 493 -1612
rect 523 -1613 710 -1612
rect 758 -1613 780 -1612
rect 786 -1613 857 -1612
rect 23 -1615 297 -1614
rect 310 -1615 328 -1614
rect 338 -1615 374 -1614
rect 415 -1615 570 -1614
rect 775 -1615 829 -1614
rect 856 -1615 997 -1614
rect 296 -1617 381 -1616
rect 537 -1617 668 -1616
rect 380 -1619 444 -1618
rect 443 -1621 542 -1620
rect 541 -1623 556 -1622
rect 548 -1625 556 -1624
rect 82 -1627 549 -1626
rect 9 -1638 342 -1637
rect 355 -1638 605 -1637
rect 607 -1638 927 -1637
rect 1059 -1638 1109 -1637
rect 23 -1640 27 -1639
rect 37 -1640 41 -1639
rect 58 -1640 696 -1639
rect 779 -1640 885 -1639
rect 1066 -1640 1095 -1639
rect 23 -1642 143 -1641
rect 149 -1642 307 -1641
rect 313 -1642 486 -1641
rect 523 -1642 661 -1641
rect 674 -1642 990 -1641
rect 1069 -1642 1116 -1641
rect 37 -1644 199 -1643
rect 222 -1644 521 -1643
rect 534 -1644 577 -1643
rect 583 -1644 948 -1643
rect 1094 -1644 1102 -1643
rect 58 -1646 101 -1645
rect 114 -1646 199 -1645
rect 247 -1646 325 -1645
rect 376 -1646 829 -1645
rect 835 -1646 885 -1645
rect 947 -1646 1074 -1645
rect 51 -1648 115 -1647
rect 135 -1648 444 -1647
rect 450 -1648 486 -1647
rect 572 -1648 913 -1647
rect 16 -1650 136 -1649
rect 138 -1650 332 -1649
rect 383 -1650 762 -1649
rect 786 -1650 829 -1649
rect 912 -1650 997 -1649
rect 61 -1652 664 -1651
rect 684 -1652 892 -1651
rect 65 -1654 101 -1653
rect 142 -1654 178 -1653
rect 187 -1654 507 -1653
rect 586 -1654 1088 -1653
rect 40 -1656 52 -1655
rect 79 -1656 381 -1655
rect 394 -1656 447 -1655
rect 450 -1656 591 -1655
rect 611 -1656 657 -1655
rect 691 -1656 717 -1655
rect 730 -1656 836 -1655
rect 891 -1656 1011 -1655
rect 82 -1658 437 -1657
rect 460 -1658 822 -1657
rect 93 -1660 129 -1659
rect 149 -1660 227 -1659
rect 254 -1660 332 -1659
rect 380 -1660 759 -1659
rect 786 -1660 871 -1659
rect 54 -1662 129 -1661
rect 159 -1662 458 -1661
rect 506 -1662 542 -1661
rect 590 -1662 598 -1661
rect 614 -1662 899 -1661
rect 96 -1664 108 -1663
rect 170 -1664 363 -1663
rect 401 -1664 626 -1663
rect 639 -1664 661 -1663
rect 667 -1664 759 -1663
rect 765 -1664 871 -1663
rect 898 -1664 962 -1663
rect 72 -1666 108 -1665
rect 156 -1666 171 -1665
rect 191 -1666 864 -1665
rect 961 -1666 983 -1665
rect 72 -1668 87 -1667
rect 191 -1668 206 -1667
rect 226 -1668 241 -1667
rect 254 -1668 262 -1667
rect 296 -1668 328 -1667
rect 387 -1668 402 -1667
rect 422 -1668 675 -1667
rect 681 -1668 766 -1667
rect 821 -1668 920 -1667
rect 86 -1670 213 -1669
rect 240 -1670 367 -1669
rect 387 -1670 570 -1669
rect 597 -1670 654 -1669
rect 695 -1670 752 -1669
rect 842 -1670 864 -1669
rect 919 -1670 1032 -1669
rect 65 -1672 654 -1671
rect 702 -1672 780 -1671
rect 842 -1672 955 -1671
rect 163 -1674 262 -1673
rect 296 -1674 311 -1673
rect 317 -1674 356 -1673
rect 366 -1674 493 -1673
rect 618 -1674 1063 -1673
rect 163 -1676 377 -1675
rect 422 -1676 538 -1675
rect 618 -1676 689 -1675
rect 702 -1676 808 -1675
rect 954 -1676 1081 -1675
rect 201 -1678 395 -1677
rect 425 -1678 906 -1677
rect 205 -1680 290 -1679
rect 317 -1680 360 -1679
rect 429 -1680 437 -1679
rect 457 -1680 465 -1679
rect 471 -1680 668 -1679
rect 716 -1680 794 -1679
rect 807 -1680 976 -1679
rect 212 -1682 416 -1681
rect 464 -1682 514 -1681
rect 625 -1682 710 -1681
rect 730 -1682 934 -1681
rect 233 -1684 311 -1683
rect 327 -1684 850 -1683
rect 905 -1684 941 -1683
rect 184 -1686 850 -1685
rect 933 -1686 1046 -1685
rect 44 -1688 185 -1687
rect 233 -1688 339 -1687
rect 359 -1688 570 -1687
rect 632 -1688 682 -1687
rect 709 -1688 738 -1687
rect 744 -1688 794 -1687
rect 940 -1688 1039 -1687
rect 44 -1690 69 -1689
rect 268 -1690 290 -1689
rect 373 -1690 430 -1689
rect 471 -1690 500 -1689
rect 513 -1690 563 -1689
rect 639 -1690 647 -1689
rect 737 -1690 878 -1689
rect 268 -1692 276 -1691
rect 373 -1692 773 -1691
rect 877 -1692 1053 -1691
rect 415 -1694 528 -1693
rect 646 -1694 678 -1693
rect 723 -1694 773 -1693
rect 408 -1696 528 -1695
rect 723 -1696 815 -1695
rect 408 -1698 580 -1697
rect 744 -1698 801 -1697
rect 478 -1700 542 -1699
rect 751 -1700 1025 -1699
rect 30 -1702 479 -1701
rect 481 -1702 563 -1701
rect 800 -1702 969 -1701
rect 30 -1704 122 -1703
rect 488 -1704 633 -1703
rect 968 -1704 1004 -1703
rect 121 -1706 283 -1705
rect 499 -1706 549 -1705
rect 282 -1708 304 -1707
rect 548 -1708 556 -1707
rect 275 -1710 304 -1709
rect 555 -1710 857 -1709
rect 856 -1712 1018 -1711
rect 2 -1723 213 -1722
rect 254 -1723 325 -1722
rect 338 -1723 608 -1722
rect 653 -1723 829 -1722
rect 849 -1723 1018 -1722
rect 1052 -1723 1070 -1722
rect 16 -1725 38 -1724
rect 51 -1725 94 -1724
rect 100 -1725 139 -1724
rect 159 -1725 241 -1724
rect 261 -1725 850 -1724
rect 870 -1725 909 -1724
rect 919 -1725 997 -1724
rect 1055 -1725 1088 -1724
rect 30 -1727 223 -1726
rect 226 -1727 262 -1726
rect 275 -1727 325 -1726
rect 359 -1727 521 -1726
rect 527 -1727 731 -1726
rect 758 -1727 808 -1726
rect 817 -1727 934 -1726
rect 940 -1727 983 -1726
rect 23 -1729 223 -1728
rect 233 -1729 255 -1728
rect 275 -1729 283 -1728
rect 296 -1729 304 -1728
rect 366 -1729 433 -1728
rect 436 -1729 524 -1728
rect 527 -1729 598 -1728
rect 632 -1729 920 -1728
rect 926 -1729 962 -1728
rect 30 -1731 678 -1730
rect 681 -1731 815 -1730
rect 828 -1731 864 -1730
rect 877 -1731 1004 -1730
rect 37 -1733 45 -1732
rect 65 -1733 458 -1732
rect 478 -1733 752 -1732
rect 761 -1733 1046 -1732
rect 44 -1735 122 -1734
rect 212 -1735 318 -1734
rect 366 -1735 381 -1734
rect 408 -1735 654 -1734
rect 660 -1735 990 -1734
rect 65 -1737 206 -1736
rect 219 -1737 318 -1736
rect 380 -1737 465 -1736
rect 495 -1737 500 -1736
rect 534 -1737 661 -1736
rect 674 -1737 857 -1736
rect 863 -1737 913 -1736
rect 926 -1737 948 -1736
rect 954 -1737 1025 -1736
rect 79 -1739 384 -1738
rect 408 -1739 503 -1738
rect 506 -1739 535 -1738
rect 586 -1739 752 -1738
rect 793 -1739 913 -1738
rect 929 -1739 962 -1738
rect 79 -1741 356 -1740
rect 425 -1741 633 -1740
rect 667 -1741 857 -1740
rect 891 -1741 941 -1740
rect 947 -1741 969 -1740
rect 86 -1743 374 -1742
rect 443 -1743 1032 -1742
rect 86 -1745 108 -1744
rect 121 -1745 377 -1744
rect 443 -1745 580 -1744
rect 597 -1745 626 -1744
rect 667 -1745 773 -1744
rect 842 -1745 878 -1744
rect 891 -1745 899 -1744
rect 905 -1745 1039 -1744
rect 100 -1747 290 -1746
rect 296 -1747 419 -1746
rect 450 -1747 584 -1746
rect 670 -1747 899 -1746
rect 107 -1749 143 -1748
rect 156 -1749 675 -1748
rect 681 -1749 710 -1748
rect 716 -1749 1060 -1748
rect 135 -1751 794 -1750
rect 800 -1751 906 -1750
rect 23 -1753 136 -1752
rect 142 -1753 192 -1752
rect 198 -1753 500 -1752
rect 506 -1753 647 -1752
rect 688 -1753 787 -1752
rect 156 -1755 388 -1754
rect 450 -1755 521 -1754
rect 569 -1755 647 -1754
rect 688 -1755 822 -1754
rect 163 -1757 717 -1756
rect 723 -1757 822 -1756
rect 149 -1759 724 -1758
rect 730 -1759 836 -1758
rect 149 -1761 346 -1760
rect 348 -1761 787 -1760
rect 163 -1763 185 -1762
rect 191 -1763 692 -1762
rect 702 -1763 871 -1762
rect 114 -1765 185 -1764
rect 198 -1765 1011 -1764
rect 226 -1767 426 -1766
rect 457 -1767 612 -1766
rect 625 -1767 801 -1766
rect 233 -1769 311 -1768
rect 373 -1769 489 -1768
rect 576 -1769 969 -1768
rect 128 -1771 311 -1770
rect 387 -1771 430 -1770
rect 464 -1771 514 -1770
rect 611 -1771 976 -1770
rect 128 -1773 248 -1772
rect 268 -1773 304 -1772
rect 306 -1773 437 -1772
rect 485 -1773 577 -1772
rect 639 -1773 703 -1772
rect 737 -1773 773 -1772
rect 240 -1775 531 -1774
rect 618 -1775 640 -1774
rect 695 -1775 738 -1774
rect 744 -1775 808 -1774
rect 268 -1777 332 -1776
rect 352 -1777 486 -1776
rect 492 -1777 745 -1776
rect 765 -1777 836 -1776
rect 58 -1779 332 -1778
rect 352 -1779 570 -1778
rect 600 -1779 696 -1778
rect 712 -1779 766 -1778
rect 58 -1781 73 -1780
rect 282 -1781 402 -1780
rect 415 -1781 493 -1780
rect 72 -1783 248 -1782
rect 289 -1783 342 -1782
rect 362 -1783 619 -1782
rect 394 -1785 514 -1784
rect 394 -1787 531 -1786
rect 401 -1789 556 -1788
rect 415 -1791 472 -1790
rect 555 -1791 591 -1790
rect 429 -1793 955 -1792
rect 471 -1795 563 -1794
rect 590 -1795 605 -1794
rect 541 -1797 563 -1796
rect 604 -1797 843 -1796
rect 541 -1799 549 -1798
rect 548 -1801 885 -1800
rect 117 -1803 885 -1802
rect 2 -1814 426 -1813
rect 443 -1814 454 -1813
rect 499 -1814 871 -1813
rect 933 -1814 948 -1813
rect 1010 -1814 1053 -1813
rect 1087 -1814 1102 -1813
rect 5 -1816 528 -1815
rect 604 -1816 703 -1815
rect 709 -1816 997 -1815
rect 1017 -1816 1074 -1815
rect 1087 -1816 1095 -1815
rect 37 -1818 41 -1817
rect 54 -1818 73 -1817
rect 79 -1818 433 -1817
rect 443 -1818 493 -1817
rect 502 -1818 654 -1817
rect 667 -1818 759 -1817
rect 912 -1818 934 -1817
rect 975 -1818 997 -1817
rect 1045 -1818 1056 -1817
rect 47 -1820 73 -1819
rect 93 -1820 850 -1819
rect 891 -1820 913 -1819
rect 926 -1820 1018 -1819
rect 103 -1822 374 -1821
rect 387 -1822 636 -1821
rect 646 -1822 871 -1821
rect 891 -1822 941 -1821
rect 954 -1822 976 -1821
rect 114 -1824 262 -1823
rect 268 -1824 363 -1823
rect 373 -1824 713 -1823
rect 733 -1824 906 -1823
rect 919 -1824 941 -1823
rect 93 -1826 115 -1825
rect 121 -1826 185 -1825
rect 198 -1826 794 -1825
rect 863 -1826 927 -1825
rect 121 -1828 584 -1827
rect 590 -1828 647 -1827
rect 688 -1828 1070 -1827
rect 124 -1830 220 -1829
rect 226 -1830 419 -1829
rect 429 -1830 948 -1829
rect 135 -1832 1011 -1831
rect 135 -1834 192 -1833
rect 194 -1834 591 -1833
rect 614 -1834 822 -1833
rect 877 -1834 906 -1833
rect 163 -1836 353 -1835
rect 366 -1836 878 -1835
rect 884 -1836 920 -1835
rect 163 -1838 552 -1837
rect 569 -1838 710 -1837
rect 737 -1838 850 -1837
rect 898 -1838 955 -1837
rect 198 -1840 360 -1839
rect 394 -1840 605 -1839
rect 628 -1840 682 -1839
rect 695 -1840 703 -1839
rect 723 -1840 738 -1839
rect 751 -1840 759 -1839
rect 765 -1840 899 -1839
rect 201 -1842 269 -1841
rect 282 -1842 388 -1841
rect 415 -1842 752 -1841
rect 772 -1842 864 -1841
rect 208 -1844 234 -1843
rect 250 -1844 619 -1843
rect 695 -1844 717 -1843
rect 723 -1844 801 -1843
rect 814 -1844 822 -1843
rect 842 -1844 885 -1843
rect 226 -1846 559 -1845
rect 576 -1846 794 -1845
rect 800 -1846 808 -1845
rect 814 -1846 1060 -1845
rect 233 -1848 472 -1847
rect 481 -1848 717 -1847
rect 730 -1848 773 -1847
rect 786 -1848 843 -1847
rect 1031 -1848 1060 -1847
rect 254 -1850 360 -1849
rect 366 -1850 577 -1849
rect 583 -1850 626 -1849
rect 691 -1850 808 -1849
rect 989 -1850 1032 -1849
rect 100 -1852 255 -1851
rect 261 -1852 437 -1851
rect 457 -1852 682 -1851
rect 744 -1852 766 -1851
rect 779 -1852 787 -1851
rect 961 -1852 990 -1851
rect 100 -1854 206 -1853
rect 282 -1854 409 -1853
rect 418 -1854 430 -1853
rect 436 -1854 671 -1853
rect 835 -1854 962 -1853
rect 149 -1856 458 -1855
rect 485 -1856 654 -1855
rect 23 -1858 486 -1857
rect 488 -1858 745 -1857
rect 23 -1860 311 -1859
rect 317 -1860 346 -1859
rect 352 -1860 465 -1859
rect 492 -1860 507 -1859
rect 520 -1860 857 -1859
rect 65 -1862 311 -1861
rect 317 -1862 356 -1861
rect 394 -1862 671 -1861
rect 65 -1864 83 -1863
rect 205 -1864 241 -1863
rect 296 -1864 524 -1863
rect 562 -1864 626 -1863
rect 632 -1864 857 -1863
rect 79 -1866 521 -1865
rect 534 -1866 563 -1865
rect 569 -1866 731 -1865
rect 117 -1868 241 -1867
rect 303 -1868 381 -1867
rect 408 -1868 447 -1867
rect 450 -1868 465 -1867
rect 621 -1868 836 -1867
rect 117 -1870 339 -1869
rect 450 -1870 598 -1869
rect 632 -1870 1039 -1869
rect 16 -1872 339 -1871
rect 453 -1872 507 -1871
rect 639 -1872 780 -1871
rect 1003 -1872 1039 -1871
rect 128 -1874 297 -1873
rect 306 -1874 675 -1873
rect 982 -1874 1004 -1873
rect 86 -1876 129 -1875
rect 177 -1876 535 -1875
rect 548 -1876 675 -1875
rect 86 -1878 248 -1877
rect 289 -1878 381 -1877
rect 422 -1878 983 -1877
rect 9 -1880 423 -1879
rect 513 -1880 640 -1879
rect 9 -1882 17 -1881
rect 142 -1882 178 -1881
rect 212 -1882 248 -1881
rect 275 -1882 290 -1881
rect 324 -1882 370 -1881
rect 513 -1882 542 -1881
rect 96 -1884 143 -1883
rect 156 -1884 325 -1883
rect 331 -1884 472 -1883
rect 30 -1886 157 -1885
rect 170 -1886 213 -1885
rect 331 -1886 479 -1885
rect 30 -1888 45 -1887
rect 107 -1888 276 -1887
rect 390 -1888 542 -1887
rect 44 -1890 1046 -1889
rect 51 -1892 108 -1891
rect 170 -1892 349 -1891
rect 478 -1892 661 -1891
rect 51 -1894 69 -1893
rect 551 -1894 661 -1893
rect 2 -1905 528 -1904
rect 530 -1905 1032 -1904
rect 1073 -1905 1109 -1904
rect 9 -1907 41 -1906
rect 44 -1907 129 -1906
rect 142 -1907 192 -1906
rect 194 -1907 493 -1906
rect 502 -1907 535 -1906
rect 551 -1907 850 -1906
rect 1003 -1907 1032 -1906
rect 1045 -1907 1074 -1906
rect 1080 -1907 1088 -1906
rect 1101 -1907 1116 -1906
rect 9 -1909 101 -1908
rect 114 -1909 136 -1908
rect 149 -1909 269 -1908
rect 296 -1909 367 -1908
rect 369 -1909 703 -1908
rect 821 -1909 825 -1908
rect 842 -1909 1067 -1908
rect 16 -1911 482 -1910
rect 485 -1911 696 -1910
rect 702 -1911 1098 -1910
rect 19 -1913 423 -1912
rect 443 -1913 605 -1912
rect 618 -1913 920 -1912
rect 968 -1913 1004 -1912
rect 1024 -1913 1088 -1912
rect 33 -1915 1046 -1914
rect 37 -1917 395 -1916
rect 450 -1917 458 -1916
rect 471 -1917 493 -1916
rect 516 -1917 871 -1916
rect 968 -1917 997 -1916
rect 47 -1919 976 -1918
rect 51 -1921 59 -1920
rect 65 -1921 73 -1920
rect 75 -1921 500 -1920
rect 527 -1921 1039 -1920
rect 58 -1923 395 -1922
rect 453 -1923 1067 -1922
rect 82 -1925 248 -1924
rect 324 -1925 605 -1924
rect 618 -1925 857 -1924
rect 870 -1925 934 -1924
rect 947 -1925 976 -1924
rect 93 -1927 535 -1926
rect 555 -1927 745 -1926
rect 768 -1927 920 -1926
rect 926 -1927 948 -1926
rect 954 -1927 997 -1926
rect 93 -1929 220 -1928
rect 222 -1929 290 -1928
rect 324 -1929 465 -1928
rect 471 -1929 507 -1928
rect 558 -1929 843 -1928
rect 856 -1929 1070 -1928
rect 100 -1931 346 -1930
rect 348 -1931 409 -1930
rect 485 -1931 577 -1930
rect 621 -1931 794 -1930
rect 821 -1931 829 -1930
rect 912 -1931 934 -1930
rect 940 -1931 955 -1930
rect 124 -1933 1060 -1932
rect 128 -1935 377 -1934
rect 387 -1935 402 -1934
rect 506 -1935 738 -1934
rect 824 -1935 829 -1934
rect 835 -1935 941 -1934
rect 1010 -1935 1060 -1934
rect 152 -1937 878 -1936
rect 898 -1937 913 -1936
rect 23 -1939 899 -1938
rect 44 -1941 153 -1940
rect 156 -1941 836 -1940
rect 877 -1941 892 -1940
rect 107 -1943 157 -1942
rect 159 -1943 1025 -1942
rect 107 -1945 143 -1944
rect 184 -1945 269 -1944
rect 338 -1945 458 -1944
rect 576 -1945 612 -1944
rect 621 -1945 1053 -1944
rect 184 -1947 367 -1946
rect 369 -1947 409 -1946
rect 583 -1947 612 -1946
rect 632 -1947 1039 -1946
rect 198 -1949 290 -1948
rect 338 -1949 647 -1948
rect 660 -1949 794 -1948
rect 1017 -1949 1053 -1948
rect 198 -1951 283 -1950
rect 345 -1951 402 -1950
rect 569 -1951 584 -1950
rect 635 -1951 724 -1950
rect 989 -1951 1018 -1950
rect 23 -1953 724 -1952
rect 807 -1953 990 -1952
rect 54 -1955 570 -1954
rect 635 -1955 773 -1954
rect 807 -1955 885 -1954
rect 54 -1957 227 -1956
rect 229 -1957 297 -1956
rect 352 -1957 416 -1956
rect 646 -1957 906 -1956
rect 180 -1959 416 -1958
rect 625 -1959 906 -1958
rect 117 -1961 626 -1960
rect 660 -1961 780 -1960
rect 863 -1961 885 -1960
rect 208 -1963 983 -1962
rect 149 -1965 983 -1964
rect 222 -1967 262 -1966
rect 275 -1967 283 -1966
rect 331 -1967 353 -1966
rect 359 -1967 1011 -1966
rect 163 -1969 276 -1968
rect 331 -1969 374 -1968
rect 390 -1969 892 -1968
rect 163 -1971 531 -1970
rect 670 -1971 850 -1970
rect 240 -1973 423 -1972
rect 681 -1973 738 -1972
rect 751 -1973 864 -1972
rect 240 -1975 255 -1974
rect 359 -1975 381 -1974
rect 667 -1975 682 -1974
rect 688 -1975 962 -1974
rect 86 -1977 381 -1976
rect 520 -1977 668 -1976
rect 674 -1977 962 -1976
rect 61 -1979 521 -1978
rect 597 -1979 689 -1978
rect 695 -1979 710 -1978
rect 751 -1979 815 -1978
rect 233 -1981 598 -1980
rect 649 -1981 815 -1980
rect 212 -1983 234 -1982
rect 247 -1983 731 -1982
rect 758 -1983 773 -1982
rect 121 -1985 213 -1984
rect 254 -1985 304 -1984
rect 373 -1985 465 -1984
rect 653 -1985 675 -1984
rect 709 -1985 717 -1984
rect 730 -1985 801 -1984
rect 121 -1987 206 -1986
rect 303 -1987 311 -1986
rect 548 -1987 717 -1986
rect 758 -1987 766 -1986
rect 170 -1989 801 -1988
rect 170 -1991 178 -1990
rect 205 -1991 500 -1990
rect 548 -1991 1105 -1990
rect 310 -1993 542 -1992
rect 639 -1993 654 -1992
rect 317 -1995 766 -1994
rect 317 -1997 437 -1996
rect 513 -1997 542 -1996
rect 590 -1997 640 -1996
rect 261 -1999 437 -1998
rect 2 -2010 223 -2009
rect 229 -2010 374 -2009
rect 376 -2010 899 -2009
rect 926 -2010 934 -2009
rect 943 -2010 1018 -2009
rect 1080 -2010 1095 -2009
rect 1104 -2010 1109 -2009
rect 1115 -2010 1123 -2009
rect 9 -2012 24 -2011
rect 33 -2012 1025 -2011
rect 1038 -2012 1081 -2011
rect 9 -2014 164 -2013
rect 170 -2014 227 -2013
rect 275 -2014 437 -2013
rect 439 -2014 1067 -2013
rect 1073 -2014 1109 -2013
rect 16 -2016 346 -2015
rect 348 -2016 801 -2015
rect 807 -2016 934 -2015
rect 982 -2016 1018 -2015
rect 1031 -2016 1039 -2015
rect 1045 -2016 1074 -2015
rect 16 -2018 101 -2017
rect 107 -2018 584 -2017
rect 593 -2018 962 -2017
rect 996 -2018 1025 -2017
rect 1059 -2018 1095 -2017
rect 51 -2020 836 -2019
rect 863 -2020 899 -2019
rect 929 -2020 969 -2019
rect 1003 -2020 1046 -2019
rect 54 -2022 346 -2021
rect 380 -2022 461 -2021
rect 464 -2022 647 -2021
rect 688 -2022 780 -2021
rect 782 -2022 822 -2021
rect 835 -2022 913 -2021
rect 940 -2022 962 -2021
rect 975 -2022 1004 -2021
rect 1010 -2022 1067 -2021
rect 37 -2024 381 -2023
rect 394 -2024 647 -2023
rect 691 -2024 1060 -2023
rect 37 -2026 178 -2025
rect 180 -2026 234 -2025
rect 275 -2026 472 -2025
rect 502 -2026 906 -2025
rect 954 -2026 983 -2025
rect 44 -2028 465 -2027
rect 471 -2028 531 -2027
rect 569 -2028 633 -2027
rect 716 -2028 906 -2027
rect 44 -2030 213 -2029
rect 222 -2030 605 -2029
rect 611 -2030 1116 -2029
rect 58 -2032 76 -2031
rect 79 -2032 171 -2031
rect 177 -2032 283 -2031
rect 324 -2032 356 -2031
rect 394 -2032 419 -2031
rect 478 -2032 605 -2031
rect 625 -2032 1032 -2031
rect 58 -2034 850 -2033
rect 870 -2034 976 -2033
rect 65 -2036 367 -2035
rect 408 -2036 535 -2035
rect 579 -2036 780 -2035
rect 821 -2036 829 -2035
rect 842 -2036 864 -2035
rect 877 -2036 997 -2035
rect 65 -2038 129 -2037
rect 135 -2038 493 -2037
rect 513 -2038 724 -2037
rect 744 -2038 773 -2037
rect 842 -2038 892 -2037
rect 51 -2040 136 -2039
rect 149 -2040 528 -2039
rect 534 -2040 563 -2039
rect 667 -2040 871 -2039
rect 884 -2040 1011 -2039
rect 72 -2042 108 -2041
rect 110 -2042 157 -2041
rect 184 -2042 636 -2041
rect 695 -2042 724 -2041
rect 751 -2042 773 -2041
rect 891 -2042 990 -2041
rect 75 -2044 591 -2043
rect 695 -2044 731 -2043
rect 758 -2044 808 -2043
rect 79 -2046 423 -2045
rect 429 -2046 479 -2045
rect 492 -2046 500 -2045
rect 506 -2046 745 -2045
rect 761 -2046 1088 -2045
rect 86 -2048 801 -2047
rect 814 -2048 1088 -2047
rect 86 -2050 752 -2049
rect 765 -2050 1053 -2049
rect 96 -2052 794 -2051
rect 100 -2054 115 -2053
rect 117 -2054 164 -2053
rect 184 -2054 619 -2053
rect 688 -2054 794 -2053
rect 114 -2056 374 -2055
rect 401 -2056 423 -2055
rect 443 -2056 668 -2055
rect 709 -2056 731 -2055
rect 768 -2056 885 -2055
rect 121 -2058 206 -2057
rect 226 -2058 615 -2057
rect 618 -2058 682 -2057
rect 786 -2058 815 -2057
rect 82 -2060 122 -2059
rect 128 -2060 332 -2059
rect 338 -2060 528 -2059
rect 555 -2060 766 -2059
rect 110 -2062 339 -2061
rect 366 -2062 549 -2061
rect 572 -2062 787 -2061
rect 138 -2064 682 -2063
rect 138 -2066 913 -2065
rect 142 -2068 157 -2067
rect 198 -2068 234 -2067
rect 247 -2068 430 -2067
rect 443 -2068 598 -2067
rect 674 -2068 710 -2067
rect 26 -2070 598 -2069
rect 89 -2072 199 -2071
rect 247 -2072 297 -2071
rect 310 -2072 591 -2071
rect 89 -2074 738 -2073
rect 149 -2076 213 -2075
rect 254 -2076 500 -2075
rect 516 -2076 990 -2075
rect 152 -2078 192 -2077
rect 240 -2078 255 -2077
rect 282 -2078 353 -2077
rect 369 -2078 829 -2077
rect 152 -2080 969 -2079
rect 191 -2082 269 -2081
rect 289 -2082 311 -2081
rect 324 -2082 353 -2081
rect 387 -2082 402 -2081
rect 411 -2082 955 -2081
rect 240 -2084 451 -2083
rect 457 -2084 507 -2083
rect 520 -2084 563 -2083
rect 576 -2084 675 -2083
rect 737 -2084 878 -2083
rect 142 -2086 451 -2085
rect 541 -2086 556 -2085
rect 268 -2088 454 -2087
rect 541 -2088 759 -2087
rect 289 -2090 857 -2089
rect 296 -2092 304 -2091
rect 317 -2092 388 -2091
rect 411 -2092 640 -2091
rect 303 -2094 650 -2093
rect 317 -2096 360 -2095
rect 415 -2096 584 -2095
rect 639 -2096 857 -2095
rect 261 -2098 360 -2097
rect 415 -2098 850 -2097
rect 93 -2100 262 -2099
rect 331 -2100 643 -2099
rect 93 -2102 1102 -2101
rect 341 -2104 521 -2103
rect 548 -2104 661 -2103
rect 716 -2104 1102 -2103
rect 485 -2106 661 -2105
rect 485 -2108 703 -2107
rect 653 -2110 703 -2109
rect 653 -2112 1053 -2111
rect 9 -2123 398 -2122
rect 401 -2123 419 -2122
rect 432 -2123 605 -2122
rect 611 -2123 1116 -2122
rect 9 -2125 255 -2124
rect 275 -2125 416 -2124
rect 436 -2125 580 -2124
rect 590 -2125 629 -2124
rect 642 -2125 1011 -2124
rect 1052 -2125 1056 -2124
rect 1101 -2125 1123 -2124
rect 16 -2127 458 -2126
rect 485 -2127 500 -2126
rect 523 -2127 808 -2126
rect 873 -2127 962 -2126
rect 16 -2129 90 -2128
rect 93 -2129 276 -2128
rect 282 -2129 339 -2128
rect 359 -2129 570 -2128
rect 576 -2129 983 -2128
rect 23 -2131 150 -2130
rect 152 -2131 367 -2130
rect 373 -2131 451 -2130
rect 485 -2131 542 -2130
rect 548 -2131 563 -2130
rect 565 -2131 1018 -2130
rect 23 -2133 584 -2132
rect 604 -2133 1046 -2132
rect 30 -2135 41 -2134
rect 58 -2135 171 -2134
rect 173 -2135 346 -2134
rect 366 -2135 381 -2134
rect 394 -2135 584 -2134
rect 611 -2135 710 -2134
rect 730 -2135 734 -2134
rect 737 -2135 997 -2134
rect 1017 -2135 1095 -2134
rect 51 -2137 381 -2136
rect 401 -2137 671 -2136
rect 684 -2137 976 -2136
rect 982 -2137 1088 -2136
rect 51 -2139 339 -2138
rect 376 -2139 409 -2138
rect 415 -2139 699 -2138
rect 723 -2139 738 -2138
rect 807 -2139 878 -2138
rect 940 -2139 955 -2138
rect 961 -2139 1025 -2138
rect 1038 -2139 1046 -2138
rect 58 -2141 388 -2140
rect 408 -2141 493 -2140
rect 530 -2141 990 -2140
rect 61 -2143 542 -2142
rect 548 -2143 552 -2142
rect 555 -2143 573 -2142
rect 593 -2143 1025 -2142
rect 72 -2145 507 -2144
rect 534 -2145 601 -2144
rect 625 -2145 1004 -2144
rect 75 -2147 1011 -2146
rect 75 -2149 661 -2148
rect 691 -2149 815 -2148
rect 891 -2149 955 -2148
rect 989 -2149 1109 -2148
rect 79 -2151 801 -2150
rect 814 -2151 829 -2150
rect 835 -2151 892 -2150
rect 947 -2151 997 -2150
rect 1003 -2151 1081 -2150
rect 79 -2153 192 -2152
rect 219 -2153 342 -2152
rect 443 -2153 510 -2152
rect 534 -2153 668 -2152
rect 695 -2153 878 -2152
rect 947 -2153 969 -2152
rect 86 -2155 472 -2154
rect 527 -2155 969 -2154
rect 72 -2157 87 -2156
rect 93 -2157 192 -2156
rect 226 -2157 577 -2156
rect 625 -2157 703 -2156
rect 730 -2157 843 -2156
rect 96 -2159 598 -2158
rect 653 -2159 696 -2158
rect 702 -2159 773 -2158
rect 786 -2159 801 -2158
rect 828 -2159 864 -2158
rect 107 -2161 290 -2160
rect 317 -2161 388 -2160
rect 443 -2161 465 -2160
rect 471 -2161 762 -2160
rect 765 -2161 773 -2160
rect 779 -2161 787 -2160
rect 835 -2161 871 -2160
rect 37 -2163 780 -2162
rect 863 -2163 906 -2162
rect 44 -2165 290 -2164
rect 320 -2165 976 -2164
rect 44 -2167 213 -2166
rect 226 -2167 304 -2166
rect 324 -2167 360 -2166
rect 453 -2167 1039 -2166
rect 107 -2169 167 -2168
rect 177 -2169 283 -2168
rect 303 -2169 430 -2168
rect 464 -2169 479 -2168
rect 527 -2169 727 -2168
rect 744 -2169 843 -2168
rect 905 -2169 1032 -2168
rect 65 -2171 178 -2170
rect 198 -2171 325 -2170
rect 345 -2171 430 -2170
rect 555 -2171 633 -2170
rect 656 -2171 1074 -2170
rect 65 -2173 269 -2172
rect 422 -2173 479 -2172
rect 597 -2173 934 -2172
rect 110 -2175 591 -2174
rect 632 -2175 647 -2174
rect 660 -2175 682 -2174
rect 733 -2175 745 -2174
rect 751 -2175 766 -2174
rect 114 -2177 122 -2176
rect 128 -2177 136 -2176
rect 138 -2177 857 -2176
rect 82 -2179 129 -2178
rect 142 -2179 503 -2178
rect 513 -2179 752 -2178
rect 117 -2181 794 -2180
rect 142 -2183 241 -2182
rect 261 -2183 342 -2182
rect 422 -2183 741 -2182
rect 149 -2185 157 -2184
rect 163 -2185 255 -2184
rect 261 -2185 297 -2184
rect 436 -2185 934 -2184
rect 121 -2187 297 -2186
rect 513 -2187 724 -2186
rect 124 -2189 157 -2188
rect 184 -2189 241 -2188
rect 268 -2189 332 -2188
rect 639 -2189 794 -2188
rect 2 -2191 640 -2190
rect 646 -2191 675 -2190
rect 688 -2191 857 -2190
rect 2 -2193 759 -2192
rect 124 -2195 1032 -2194
rect 198 -2197 356 -2196
rect 667 -2197 1067 -2196
rect 212 -2199 293 -2198
rect 310 -2199 332 -2198
rect 674 -2199 717 -2198
rect 758 -2199 913 -2198
rect 233 -2201 440 -2200
rect 618 -2201 717 -2200
rect 912 -2201 920 -2200
rect 205 -2203 234 -2202
rect 247 -2203 311 -2202
rect 520 -2203 619 -2202
rect 919 -2203 927 -2202
rect 205 -2205 493 -2204
rect 520 -2205 710 -2204
rect 926 -2205 1060 -2204
rect 247 -2207 608 -2206
rect 9 -2218 206 -2217
rect 208 -2218 640 -2217
rect 653 -2218 671 -2217
rect 691 -2218 864 -2217
rect 870 -2218 969 -2217
rect 9 -2220 339 -2219
rect 341 -2220 486 -2219
rect 488 -2220 780 -2219
rect 856 -2220 930 -2219
rect 16 -2222 104 -2221
rect 121 -2222 255 -2221
rect 282 -2222 318 -2221
rect 348 -2222 367 -2221
rect 373 -2222 472 -2221
rect 485 -2222 689 -2221
rect 695 -2222 983 -2221
rect 30 -2224 346 -2223
rect 355 -2224 388 -2223
rect 394 -2224 1032 -2223
rect 44 -2226 384 -2225
rect 387 -2226 423 -2225
rect 436 -2226 682 -2225
rect 695 -2226 738 -2225
rect 768 -2226 801 -2225
rect 856 -2226 1018 -2225
rect 37 -2228 45 -2227
rect 51 -2228 192 -2227
rect 194 -2228 213 -2227
rect 215 -2228 297 -2227
rect 310 -2228 339 -2227
rect 359 -2228 395 -2227
rect 401 -2228 423 -2227
rect 439 -2228 1011 -2227
rect 30 -2230 52 -2229
rect 93 -2230 174 -2229
rect 177 -2230 304 -2229
rect 317 -2230 325 -2229
rect 331 -2230 356 -2229
rect 359 -2230 580 -2229
rect 590 -2230 836 -2229
rect 863 -2230 1025 -2229
rect 23 -2232 304 -2231
rect 331 -2232 500 -2231
rect 502 -2232 521 -2231
rect 548 -2232 570 -2231
rect 572 -2232 703 -2231
rect 723 -2232 815 -2231
rect 835 -2232 962 -2231
rect 23 -2234 164 -2233
rect 166 -2234 545 -2233
rect 576 -2234 640 -2233
rect 653 -2234 710 -2233
rect 723 -2234 773 -2233
rect 779 -2234 794 -2233
rect 800 -2234 913 -2233
rect 922 -2234 997 -2233
rect 37 -2236 143 -2235
rect 156 -2236 185 -2235
rect 201 -2236 566 -2235
rect 590 -2236 633 -2235
rect 667 -2236 731 -2235
rect 737 -2236 787 -2235
rect 793 -2236 941 -2235
rect 961 -2236 1004 -2235
rect 2 -2238 143 -2237
rect 170 -2238 276 -2237
rect 282 -2238 398 -2237
rect 401 -2238 493 -2237
rect 506 -2238 556 -2237
rect 597 -2238 717 -2237
rect 726 -2238 1046 -2237
rect 2 -2240 115 -2239
rect 121 -2240 584 -2239
rect 604 -2240 619 -2239
rect 681 -2240 731 -2239
rect 758 -2240 787 -2239
rect 814 -2240 829 -2239
rect 940 -2240 990 -2239
rect 79 -2242 164 -2241
rect 198 -2242 276 -2241
rect 296 -2242 328 -2241
rect 408 -2242 510 -2241
rect 513 -2242 633 -2241
rect 698 -2242 906 -2241
rect 93 -2244 108 -2243
rect 114 -2244 129 -2243
rect 135 -2244 293 -2243
rect 380 -2244 409 -2243
rect 429 -2244 514 -2243
rect 527 -2244 556 -2243
rect 583 -2244 843 -2243
rect 100 -2246 108 -2245
rect 135 -2246 150 -2245
rect 156 -2246 199 -2245
rect 205 -2246 220 -2245
rect 226 -2246 381 -2245
rect 429 -2246 542 -2245
rect 548 -2246 577 -2245
rect 604 -2246 647 -2245
rect 709 -2246 766 -2245
rect 772 -2246 850 -2245
rect 65 -2248 150 -2247
rect 212 -2248 269 -2247
rect 450 -2248 563 -2247
rect 618 -2248 626 -2247
rect 646 -2248 685 -2247
rect 716 -2248 892 -2247
rect 33 -2250 269 -2249
rect 450 -2250 745 -2249
rect 758 -2250 822 -2249
rect 828 -2250 934 -2249
rect 65 -2252 188 -2251
rect 226 -2252 290 -2251
rect 352 -2252 745 -2251
rect 821 -2252 976 -2251
rect 72 -2254 220 -2253
rect 240 -2254 325 -2253
rect 352 -2254 465 -2253
rect 467 -2254 528 -2253
rect 541 -2254 878 -2253
rect 891 -2254 1039 -2253
rect 240 -2256 416 -2255
rect 457 -2256 482 -2255
rect 593 -2256 626 -2255
rect 684 -2256 703 -2255
rect 842 -2256 920 -2255
rect 968 -2256 976 -2255
rect 58 -2258 416 -2257
rect 443 -2258 458 -2257
rect 471 -2258 612 -2257
rect 849 -2258 899 -2257
rect 912 -2258 934 -2257
rect 16 -2260 59 -2259
rect 254 -2260 370 -2259
rect 443 -2260 675 -2259
rect 877 -2260 927 -2259
rect 261 -2262 311 -2261
rect 478 -2262 675 -2261
rect 233 -2264 262 -2263
rect 478 -2264 493 -2263
rect 534 -2264 899 -2263
rect 233 -2266 524 -2265
rect 611 -2266 661 -2265
rect 502 -2268 535 -2267
rect 660 -2268 752 -2267
rect 751 -2270 808 -2269
rect 807 -2272 948 -2271
rect 947 -2274 955 -2273
rect 464 -2276 955 -2275
rect 2 -2287 52 -2286
rect 58 -2287 276 -2286
rect 303 -2287 479 -2286
rect 481 -2287 892 -2286
rect 905 -2287 934 -2286
rect 2 -2289 31 -2288
rect 44 -2289 55 -2288
rect 58 -2289 437 -2288
rect 450 -2289 468 -2288
rect 499 -2289 612 -2288
rect 642 -2289 801 -2288
rect 877 -2289 892 -2288
rect 908 -2289 948 -2288
rect 9 -2291 129 -2290
rect 191 -2291 213 -2290
rect 226 -2291 346 -2290
rect 376 -2291 647 -2290
rect 684 -2291 836 -2290
rect 877 -2291 955 -2290
rect 12 -2293 216 -2292
rect 268 -2293 489 -2292
rect 502 -2293 724 -2292
rect 765 -2293 829 -2292
rect 884 -2293 913 -2292
rect 922 -2293 930 -2292
rect 947 -2293 962 -2292
rect 16 -2295 486 -2294
rect 534 -2295 566 -2294
rect 576 -2295 857 -2294
rect 926 -2295 976 -2294
rect 16 -2297 234 -2296
rect 268 -2297 297 -2296
rect 303 -2297 416 -2296
rect 436 -2297 458 -2296
rect 464 -2297 563 -2296
rect 583 -2297 661 -2296
rect 723 -2297 822 -2296
rect 842 -2297 885 -2296
rect 23 -2299 52 -2298
rect 61 -2299 706 -2298
rect 768 -2299 850 -2298
rect 856 -2299 899 -2298
rect 23 -2301 283 -2300
rect 296 -2301 465 -2300
rect 467 -2301 472 -2300
rect 520 -2301 577 -2300
rect 597 -2301 647 -2300
rect 779 -2301 829 -2300
rect 849 -2301 902 -2300
rect 30 -2303 230 -2302
rect 233 -2303 262 -2302
rect 275 -2303 363 -2302
rect 373 -2303 486 -2302
rect 562 -2303 759 -2302
rect 786 -2303 822 -2302
rect 44 -2305 780 -2304
rect 793 -2305 843 -2304
rect 47 -2307 132 -2306
rect 163 -2307 192 -2306
rect 261 -2307 290 -2306
rect 310 -2307 335 -2306
rect 341 -2307 717 -2306
rect 793 -2307 864 -2306
rect 65 -2309 311 -2308
rect 313 -2309 787 -2308
rect 800 -2309 815 -2308
rect 65 -2311 101 -2310
rect 107 -2311 626 -2310
rect 667 -2311 815 -2310
rect 72 -2313 178 -2312
rect 282 -2313 409 -2312
rect 415 -2313 717 -2312
rect 72 -2315 80 -2314
rect 82 -2315 87 -2314
rect 93 -2315 104 -2314
rect 107 -2315 111 -2314
rect 114 -2315 199 -2314
rect 289 -2315 339 -2314
rect 355 -2315 472 -2314
rect 537 -2315 759 -2314
rect 79 -2317 150 -2316
rect 163 -2317 339 -2316
rect 355 -2317 661 -2316
rect 681 -2317 864 -2316
rect 86 -2319 542 -2318
rect 586 -2319 668 -2318
rect 93 -2321 524 -2320
rect 597 -2321 605 -2320
rect 611 -2321 633 -2320
rect 100 -2323 423 -2322
rect 450 -2323 731 -2322
rect 114 -2325 136 -2324
rect 149 -2325 185 -2324
rect 198 -2325 206 -2324
rect 317 -2325 398 -2324
rect 401 -2325 542 -2324
rect 625 -2325 689 -2324
rect 54 -2327 136 -2326
rect 142 -2327 185 -2326
rect 205 -2327 349 -2326
rect 359 -2327 731 -2326
rect 128 -2329 241 -2328
rect 317 -2329 675 -2328
rect 688 -2329 696 -2328
rect 142 -2331 157 -2330
rect 177 -2331 248 -2330
rect 324 -2331 444 -2330
rect 513 -2331 633 -2330
rect 674 -2331 710 -2330
rect 37 -2333 157 -2332
rect 180 -2333 696 -2332
rect 702 -2333 710 -2332
rect 37 -2335 111 -2334
rect 121 -2335 248 -2334
rect 254 -2335 514 -2334
rect 702 -2335 752 -2334
rect 121 -2337 293 -2336
rect 359 -2337 395 -2336
rect 401 -2337 654 -2336
rect 737 -2337 752 -2336
rect 240 -2339 528 -2338
rect 737 -2339 745 -2338
rect 254 -2341 580 -2340
rect 744 -2341 773 -2340
rect 352 -2343 528 -2342
rect 772 -2343 871 -2342
rect 366 -2345 605 -2344
rect 870 -2345 941 -2344
rect 170 -2347 367 -2346
rect 380 -2347 682 -2346
rect 159 -2349 171 -2348
rect 331 -2349 381 -2348
rect 383 -2349 409 -2348
rect 422 -2349 430 -2348
rect 443 -2349 549 -2348
rect 373 -2351 430 -2350
rect 492 -2351 654 -2350
rect 394 -2353 836 -2352
rect 492 -2355 556 -2354
rect 548 -2357 591 -2356
rect 544 -2359 591 -2358
rect 555 -2361 808 -2360
rect 583 -2363 808 -2362
rect 16 -2374 139 -2373
rect 156 -2374 216 -2373
rect 226 -2374 668 -2373
rect 702 -2374 710 -2373
rect 726 -2374 822 -2373
rect 940 -2374 948 -2373
rect 23 -2376 220 -2375
rect 240 -2376 559 -2375
rect 569 -2376 668 -2375
rect 709 -2376 766 -2375
rect 772 -2376 829 -2375
rect 30 -2378 157 -2377
rect 177 -2378 227 -2377
rect 233 -2378 241 -2377
rect 247 -2378 353 -2377
rect 376 -2378 759 -2377
rect 761 -2378 843 -2377
rect 2 -2380 31 -2379
rect 44 -2380 62 -2379
rect 93 -2380 209 -2379
rect 212 -2380 374 -2379
rect 404 -2380 780 -2379
rect 828 -2380 878 -2379
rect 37 -2382 94 -2381
rect 100 -2382 360 -2381
rect 411 -2382 437 -2381
rect 457 -2382 577 -2381
rect 583 -2382 661 -2381
rect 723 -2382 766 -2381
rect 772 -2382 794 -2381
rect 51 -2384 731 -2383
rect 751 -2384 755 -2383
rect 100 -2386 150 -2385
rect 177 -2386 255 -2385
rect 268 -2386 290 -2385
rect 303 -2386 419 -2385
rect 460 -2386 507 -2385
rect 520 -2386 549 -2385
rect 555 -2386 626 -2385
rect 639 -2386 689 -2385
rect 723 -2386 850 -2385
rect 107 -2388 451 -2387
rect 464 -2388 507 -2387
rect 523 -2388 612 -2387
rect 618 -2388 629 -2387
rect 639 -2388 836 -2387
rect 107 -2390 150 -2389
rect 163 -2390 290 -2389
rect 310 -2390 605 -2389
rect 611 -2390 675 -2389
rect 114 -2392 153 -2391
rect 163 -2392 185 -2391
rect 205 -2392 248 -2391
rect 275 -2392 398 -2391
rect 408 -2392 437 -2391
rect 450 -2392 472 -2391
rect 481 -2392 717 -2391
rect 114 -2394 171 -2393
rect 184 -2394 223 -2393
rect 233 -2394 388 -2393
rect 408 -2394 647 -2393
rect 660 -2394 738 -2393
rect 121 -2396 272 -2395
rect 275 -2396 423 -2395
rect 464 -2396 815 -2395
rect 65 -2398 122 -2397
rect 135 -2398 304 -2397
rect 310 -2398 356 -2397
rect 380 -2398 605 -2397
rect 618 -2398 696 -2397
rect 716 -2398 808 -2397
rect 170 -2400 192 -2399
rect 219 -2400 549 -2399
rect 551 -2400 647 -2399
rect 674 -2400 787 -2399
rect 807 -2400 864 -2399
rect 191 -2402 199 -2401
rect 282 -2402 458 -2401
rect 471 -2402 563 -2401
rect 737 -2402 745 -2401
rect 128 -2404 283 -2403
rect 313 -2404 542 -2403
rect 744 -2404 857 -2403
rect 128 -2406 297 -2405
rect 324 -2406 342 -2405
rect 345 -2406 423 -2405
rect 527 -2406 570 -2405
rect 79 -2408 297 -2407
rect 317 -2408 346 -2407
rect 527 -2408 591 -2407
rect 58 -2410 80 -2409
rect 198 -2410 223 -2409
rect 317 -2410 545 -2409
rect 58 -2412 66 -2411
rect 324 -2412 416 -2411
rect 534 -2412 598 -2411
rect 331 -2414 381 -2413
rect 415 -2414 430 -2413
rect 499 -2414 535 -2413
rect 597 -2414 682 -2413
rect 331 -2416 367 -2415
rect 429 -2416 591 -2415
rect 653 -2416 682 -2415
rect 334 -2418 388 -2417
rect 401 -2418 654 -2417
rect 254 -2420 335 -2419
rect 338 -2420 514 -2419
rect 366 -2422 486 -2421
rect 499 -2422 633 -2421
rect 401 -2424 493 -2423
rect 513 -2424 566 -2423
rect 443 -2426 493 -2425
rect 394 -2428 444 -2427
rect 488 -2428 633 -2427
rect 65 -2439 73 -2438
rect 79 -2439 265 -2438
rect 268 -2439 409 -2438
rect 422 -2439 465 -2438
rect 471 -2439 584 -2438
rect 590 -2439 594 -2438
rect 625 -2439 717 -2438
rect 730 -2439 738 -2438
rect 754 -2439 808 -2438
rect 926 -2439 934 -2438
rect 93 -2441 132 -2440
rect 135 -2441 143 -2440
rect 170 -2441 216 -2440
rect 233 -2441 370 -2440
rect 401 -2441 472 -2440
rect 474 -2441 482 -2440
rect 485 -2441 605 -2440
rect 625 -2441 661 -2440
rect 681 -2441 689 -2440
rect 695 -2441 703 -2440
rect 716 -2441 727 -2440
rect 730 -2441 734 -2440
rect 779 -2441 829 -2440
rect 100 -2443 157 -2442
rect 191 -2443 209 -2442
rect 240 -2443 258 -2442
rect 275 -2443 332 -2442
rect 334 -2443 391 -2442
rect 408 -2443 416 -2442
rect 422 -2443 479 -2442
rect 502 -2443 570 -2442
rect 576 -2443 654 -2442
rect 660 -2443 668 -2442
rect 681 -2443 710 -2442
rect 100 -2445 118 -2444
rect 121 -2445 220 -2444
rect 226 -2445 276 -2444
rect 296 -2445 598 -2444
rect 604 -2445 612 -2444
rect 642 -2445 647 -2444
rect 709 -2445 745 -2444
rect 107 -2447 122 -2446
rect 128 -2447 220 -2446
rect 226 -2447 262 -2446
rect 310 -2447 489 -2446
rect 506 -2447 601 -2446
rect 611 -2447 633 -2446
rect 114 -2449 234 -2448
rect 254 -2449 269 -2448
rect 317 -2449 433 -2448
rect 443 -2449 479 -2448
rect 499 -2449 507 -2448
rect 513 -2449 580 -2448
rect 107 -2451 115 -2450
rect 149 -2451 171 -2450
rect 191 -2451 199 -2450
rect 222 -2451 311 -2450
rect 345 -2451 402 -2450
rect 443 -2451 451 -2450
rect 457 -2451 493 -2450
rect 513 -2451 535 -2450
rect 541 -2451 563 -2450
rect 569 -2451 619 -2450
rect 86 -2453 451 -2452
rect 460 -2453 521 -2452
rect 527 -2453 552 -2452
rect 555 -2453 577 -2452
rect 152 -2455 199 -2454
rect 282 -2455 318 -2454
rect 331 -2455 346 -2454
rect 348 -2455 388 -2454
rect 534 -2455 675 -2454
rect 163 -2457 241 -2456
rect 289 -2457 433 -2456
rect 548 -2457 640 -2456
rect 674 -2457 759 -2456
rect 163 -2459 185 -2458
rect 212 -2459 283 -2458
rect 352 -2459 395 -2458
rect 639 -2459 724 -2458
rect 737 -2459 759 -2458
rect 184 -2461 206 -2460
rect 247 -2461 290 -2460
rect 324 -2461 353 -2460
rect 359 -2461 468 -2460
rect 723 -2461 762 -2460
rect 177 -2463 248 -2462
rect 338 -2463 360 -2462
rect 366 -2463 416 -2462
rect 761 -2463 773 -2462
rect 159 -2465 178 -2464
rect 299 -2465 339 -2464
rect 387 -2465 437 -2464
rect 380 -2467 437 -2466
rect 373 -2469 381 -2468
rect 394 -2469 398 -2468
rect 65 -2480 73 -2479
rect 86 -2480 97 -2479
rect 100 -2480 111 -2479
rect 114 -2480 122 -2479
rect 131 -2480 136 -2479
rect 142 -2480 171 -2479
rect 177 -2480 188 -2479
rect 198 -2480 213 -2479
rect 219 -2480 255 -2479
rect 282 -2480 363 -2479
rect 376 -2480 423 -2479
rect 432 -2480 458 -2479
rect 467 -2480 479 -2479
rect 502 -2480 514 -2479
rect 523 -2480 542 -2479
rect 576 -2480 587 -2479
rect 590 -2480 626 -2479
rect 667 -2480 682 -2479
rect 744 -2480 752 -2479
rect 758 -2480 766 -2479
rect 933 -2480 937 -2479
rect 940 -2480 948 -2479
rect 100 -2482 122 -2481
rect 138 -2482 220 -2481
rect 226 -2482 230 -2481
rect 247 -2482 325 -2481
rect 338 -2482 405 -2481
rect 450 -2482 549 -2481
rect 597 -2482 675 -2481
rect 681 -2482 689 -2481
rect 758 -2482 762 -2481
rect 107 -2484 115 -2483
rect 149 -2484 164 -2483
rect 177 -2484 192 -2483
rect 226 -2484 262 -2483
rect 275 -2484 325 -2483
rect 359 -2484 374 -2483
rect 401 -2484 423 -2483
rect 443 -2484 451 -2483
rect 471 -2484 528 -2483
rect 688 -2484 696 -2483
rect 159 -2486 171 -2485
rect 233 -2486 262 -2485
rect 271 -2486 276 -2485
rect 296 -2486 304 -2485
rect 310 -2486 367 -2485
rect 401 -2486 538 -2485
rect 695 -2486 710 -2485
rect 229 -2488 234 -2487
rect 236 -2488 311 -2487
rect 359 -2488 409 -2487
rect 415 -2488 444 -2487
rect 506 -2488 521 -2487
rect 523 -2488 528 -2487
rect 709 -2488 717 -2487
rect 240 -2490 297 -2489
rect 303 -2490 332 -2489
rect 408 -2490 437 -2489
rect 520 -2490 570 -2489
rect 716 -2490 724 -2489
rect 247 -2492 269 -2491
rect 317 -2492 332 -2491
rect 723 -2492 738 -2491
rect 289 -2494 318 -2493
rect 201 -2496 290 -2495
rect 5 -2507 10 -2506
rect 86 -2507 104 -2506
rect 107 -2507 122 -2506
rect 142 -2507 195 -2506
rect 201 -2507 206 -2506
rect 219 -2507 241 -2506
rect 247 -2507 272 -2506
rect 275 -2507 283 -2506
rect 285 -2507 318 -2506
rect 331 -2507 346 -2506
rect 352 -2507 363 -2506
rect 380 -2507 384 -2506
rect 387 -2507 409 -2506
rect 450 -2507 458 -2506
rect 523 -2507 528 -2506
rect 597 -2507 605 -2506
rect 660 -2507 664 -2506
rect 681 -2507 703 -2506
rect 709 -2507 713 -2506
rect 723 -2507 731 -2506
rect 740 -2507 752 -2506
rect 887 -2507 892 -2506
rect 933 -2507 941 -2506
rect 943 -2507 948 -2506
rect 100 -2509 108 -2508
rect 114 -2509 118 -2508
rect 149 -2509 167 -2508
rect 184 -2509 188 -2508
rect 191 -2509 227 -2508
rect 229 -2509 234 -2508
rect 254 -2509 279 -2508
rect 289 -2509 304 -2508
rect 394 -2509 398 -2508
rect 404 -2509 419 -2508
rect 443 -2509 451 -2508
rect 604 -2509 612 -2508
rect 695 -2509 706 -2508
rect 744 -2509 759 -2508
rect 156 -2511 160 -2510
rect 163 -2511 171 -2510
rect 177 -2511 192 -2510
rect 212 -2511 227 -2510
rect 261 -2511 269 -2510
rect 296 -2511 311 -2510
rect 401 -2511 405 -2510
rect 163 -2513 181 -2512
rect 299 -2513 342 -2512
rect 310 -2515 325 -2514
rect 5 -2526 10 -2525
rect 100 -2526 108 -2525
rect 114 -2526 125 -2525
rect 163 -2526 171 -2525
rect 180 -2526 185 -2525
rect 191 -2526 199 -2525
rect 292 -2526 297 -2525
rect 303 -2526 311 -2525
rect 341 -2526 346 -2525
rect 450 -2526 458 -2525
rect 597 -2526 605 -2525
rect 663 -2526 668 -2525
rect 716 -2526 724 -2525
rect 730 -2526 741 -2525
rect 121 -2528 132 -2527
<< m2contact >>
rect 93 0 94 1
rect 100 0 101 1
rect 107 0 108 1
rect 128 0 129 1
rect 205 0 206 1
rect 212 0 213 1
rect 215 0 216 1
rect 236 0 237 1
rect 240 0 241 1
rect 247 0 248 1
rect 261 0 262 1
rect 268 0 269 1
rect 324 0 325 1
rect 334 0 335 1
rect 429 0 430 1
rect 450 0 451 1
rect 464 0 465 1
rect 488 0 489 1
rect 530 0 531 1
rect 534 0 535 1
rect 583 0 584 1
rect 597 0 598 1
rect 660 0 661 1
rect 667 0 668 1
rect 117 -2 118 -1
rect 121 -2 122 -1
rect 226 -2 227 -1
rect 233 -2 234 -1
rect 86 -13 87 -12
rect 103 -13 104 -12
rect 117 -13 118 -12
rect 128 -13 129 -12
rect 135 -13 136 -12
rect 145 -13 146 -12
rect 173 -13 174 -12
rect 198 -13 199 -12
rect 205 -13 206 -12
rect 215 -13 216 -12
rect 226 -13 227 -12
rect 250 -13 251 -12
rect 254 -13 255 -12
rect 268 -13 269 -12
rect 289 -13 290 -12
rect 306 -13 307 -12
rect 310 -13 311 -12
rect 324 -13 325 -12
rect 348 -13 349 -12
rect 359 -13 360 -12
rect 373 -13 374 -12
rect 446 -13 447 -12
rect 450 -13 451 -12
rect 464 -13 465 -12
rect 485 -13 486 -12
rect 527 -13 528 -12
rect 534 -13 535 -12
rect 541 -13 542 -12
rect 548 -13 549 -12
rect 569 -13 570 -12
rect 590 -13 591 -12
rect 604 -13 605 -12
rect 607 -13 608 -12
rect 618 -13 619 -12
rect 667 -13 668 -12
rect 674 -13 675 -12
rect 89 -15 90 -14
rect 100 -15 101 -14
rect 177 -15 178 -14
rect 212 -15 213 -14
rect 219 -15 220 -14
rect 226 -15 227 -14
rect 233 -15 234 -14
rect 247 -15 248 -14
rect 257 -15 258 -14
rect 275 -15 276 -14
rect 317 -15 318 -14
rect 331 -15 332 -14
rect 415 -15 416 -14
rect 429 -15 430 -14
rect 453 -15 454 -14
rect 471 -15 472 -14
rect 492 -15 493 -14
rect 513 -15 514 -14
rect 562 -15 563 -14
rect 576 -15 577 -14
rect 597 -15 598 -14
rect 611 -15 612 -14
rect 93 -17 94 -16
rect 107 -17 108 -16
rect 184 -17 185 -16
rect 205 -17 206 -16
rect 219 -17 220 -16
rect 222 -17 223 -16
rect 261 -17 262 -16
rect 282 -17 283 -16
rect 324 -17 325 -16
rect 341 -17 342 -16
rect 429 -17 430 -16
rect 439 -17 440 -16
rect 506 -17 507 -16
rect 509 -17 510 -16
rect 100 -19 101 -18
rect 121 -19 122 -18
rect 236 -19 237 -18
rect 282 -19 283 -18
rect 268 -21 269 -20
rect 303 -21 304 -20
rect 86 -32 87 -31
rect 103 -32 104 -31
rect 114 -32 115 -31
rect 187 -32 188 -31
rect 191 -32 192 -31
rect 219 -32 220 -31
rect 226 -32 227 -31
rect 229 -32 230 -31
rect 247 -32 248 -31
rect 352 -32 353 -31
rect 359 -32 360 -31
rect 408 -32 409 -31
rect 415 -32 416 -31
rect 422 -32 423 -31
rect 429 -32 430 -31
rect 436 -32 437 -31
rect 446 -32 447 -31
rect 499 -32 500 -31
rect 520 -32 521 -31
rect 534 -32 535 -31
rect 551 -32 552 -31
rect 562 -32 563 -31
rect 569 -32 570 -31
rect 597 -32 598 -31
rect 604 -32 605 -31
rect 639 -32 640 -31
rect 663 -32 664 -31
rect 667 -32 668 -31
rect 674 -32 675 -31
rect 702 -32 703 -31
rect 765 -32 766 -31
rect 842 -32 843 -31
rect 93 -34 94 -33
rect 100 -34 101 -33
rect 121 -34 122 -33
rect 135 -34 136 -33
rect 163 -34 164 -33
rect 236 -34 237 -33
rect 247 -34 248 -33
rect 254 -34 255 -33
rect 275 -34 276 -33
rect 345 -34 346 -33
rect 366 -34 367 -33
rect 373 -34 374 -33
rect 383 -34 384 -33
rect 394 -34 395 -33
rect 471 -34 472 -33
rect 520 -34 521 -33
rect 527 -34 528 -33
rect 590 -34 591 -33
rect 611 -34 612 -33
rect 653 -34 654 -33
rect 677 -34 678 -33
rect 681 -34 682 -33
rect 128 -36 129 -35
rect 145 -36 146 -35
rect 177 -36 178 -35
rect 194 -36 195 -35
rect 198 -36 199 -35
rect 205 -36 206 -35
rect 212 -36 213 -35
rect 275 -36 276 -35
rect 282 -36 283 -35
rect 303 -36 304 -35
rect 313 -36 314 -35
rect 317 -36 318 -35
rect 341 -36 342 -35
rect 422 -36 423 -35
rect 464 -36 465 -35
rect 611 -36 612 -35
rect 618 -36 619 -35
rect 646 -36 647 -35
rect 135 -38 136 -37
rect 268 -38 269 -37
rect 282 -38 283 -37
rect 348 -38 349 -37
rect 373 -38 374 -37
rect 443 -38 444 -37
rect 464 -38 465 -37
rect 625 -38 626 -37
rect 156 -40 157 -39
rect 177 -40 178 -39
rect 184 -40 185 -39
rect 219 -40 220 -39
rect 226 -40 227 -39
rect 261 -40 262 -39
rect 268 -40 269 -39
rect 289 -40 290 -39
rect 296 -40 297 -39
rect 429 -40 430 -39
rect 471 -40 472 -39
rect 586 -40 587 -39
rect 198 -42 199 -41
rect 331 -42 332 -41
rect 383 -42 384 -41
rect 485 -42 486 -41
rect 527 -42 528 -41
rect 632 -42 633 -41
rect 201 -44 202 -43
rect 254 -44 255 -43
rect 289 -44 290 -43
rect 324 -44 325 -43
rect 387 -44 388 -43
rect 467 -44 468 -43
rect 478 -44 479 -43
rect 492 -44 493 -43
rect 541 -44 542 -43
rect 569 -44 570 -43
rect 173 -46 174 -45
rect 324 -46 325 -45
rect 513 -46 514 -45
rect 541 -46 542 -45
rect 555 -46 556 -45
rect 604 -46 605 -45
rect 212 -48 213 -47
rect 299 -48 300 -47
rect 310 -48 311 -47
rect 317 -48 318 -47
rect 555 -48 556 -47
rect 772 -48 773 -47
rect 229 -50 230 -49
rect 261 -50 262 -49
rect 250 -52 251 -51
rect 401 -52 402 -51
rect 30 -63 31 -62
rect 152 -63 153 -62
rect 159 -63 160 -62
rect 250 -63 251 -62
rect 317 -63 318 -62
rect 338 -63 339 -62
rect 429 -63 430 -62
rect 821 -63 822 -62
rect 842 -63 843 -62
rect 877 -63 878 -62
rect 58 -65 59 -64
rect 107 -65 108 -64
rect 114 -65 115 -64
rect 173 -65 174 -64
rect 198 -65 199 -64
rect 205 -65 206 -64
rect 219 -65 220 -64
rect 229 -65 230 -64
rect 233 -65 234 -64
rect 345 -65 346 -64
rect 394 -65 395 -64
rect 429 -65 430 -64
rect 450 -65 451 -64
rect 467 -65 468 -64
rect 471 -65 472 -64
rect 474 -65 475 -64
rect 485 -65 486 -64
rect 513 -65 514 -64
rect 530 -65 531 -64
rect 688 -65 689 -64
rect 702 -65 703 -64
rect 779 -65 780 -64
rect 37 -67 38 -66
rect 173 -67 174 -66
rect 219 -67 220 -66
rect 278 -67 279 -66
rect 317 -67 318 -66
rect 716 -67 717 -66
rect 772 -67 773 -66
rect 870 -67 871 -66
rect 61 -69 62 -68
rect 320 -69 321 -68
rect 324 -69 325 -68
rect 380 -69 381 -68
rect 457 -69 458 -68
rect 555 -69 556 -68
rect 583 -69 584 -68
rect 793 -69 794 -68
rect 65 -71 66 -70
rect 93 -71 94 -70
rect 100 -71 101 -70
rect 205 -71 206 -70
rect 233 -71 234 -70
rect 387 -71 388 -70
rect 464 -71 465 -70
rect 478 -71 479 -70
rect 485 -71 486 -70
rect 499 -71 500 -70
rect 502 -71 503 -70
rect 807 -71 808 -70
rect 72 -73 73 -72
rect 128 -73 129 -72
rect 142 -73 143 -72
rect 243 -73 244 -72
rect 254 -73 255 -72
rect 555 -73 556 -72
rect 590 -73 591 -72
rect 772 -73 773 -72
rect 79 -75 80 -74
rect 86 -75 87 -74
rect 93 -75 94 -74
rect 303 -75 304 -74
rect 331 -75 332 -74
rect 695 -75 696 -74
rect 702 -75 703 -74
rect 765 -75 766 -74
rect 86 -77 87 -76
rect 282 -77 283 -76
rect 289 -77 290 -76
rect 324 -77 325 -76
rect 331 -77 332 -76
rect 352 -77 353 -76
rect 376 -77 377 -76
rect 478 -77 479 -76
rect 495 -77 496 -76
rect 828 -77 829 -76
rect 103 -79 104 -78
rect 282 -79 283 -78
rect 380 -79 381 -78
rect 408 -79 409 -78
rect 471 -79 472 -78
rect 492 -79 493 -78
rect 506 -79 507 -78
rect 509 -79 510 -78
rect 548 -79 549 -78
rect 618 -79 619 -78
rect 625 -79 626 -78
rect 814 -79 815 -78
rect 117 -81 118 -80
rect 170 -81 171 -80
rect 240 -81 241 -80
rect 408 -81 409 -80
rect 474 -81 475 -80
rect 492 -81 493 -80
rect 569 -81 570 -80
rect 625 -81 626 -80
rect 632 -81 633 -80
rect 786 -81 787 -80
rect 51 -83 52 -82
rect 240 -83 241 -82
rect 261 -83 262 -82
rect 303 -83 304 -82
rect 355 -83 356 -82
rect 632 -83 633 -82
rect 639 -83 640 -82
rect 744 -83 745 -82
rect 121 -85 122 -84
rect 254 -85 255 -84
rect 268 -85 269 -84
rect 289 -85 290 -84
rect 387 -85 388 -84
rect 835 -85 836 -84
rect 121 -87 122 -86
rect 163 -87 164 -86
rect 247 -87 248 -86
rect 261 -87 262 -86
rect 268 -87 269 -86
rect 373 -87 374 -86
rect 397 -87 398 -86
rect 548 -87 549 -86
rect 586 -87 587 -86
rect 590 -87 591 -86
rect 604 -87 605 -86
rect 737 -87 738 -86
rect 128 -89 129 -88
rect 674 -89 675 -88
rect 681 -89 682 -88
rect 730 -89 731 -88
rect 149 -91 150 -90
rect 156 -91 157 -90
rect 163 -91 164 -90
rect 418 -91 419 -90
rect 527 -91 528 -90
rect 586 -91 587 -90
rect 597 -91 598 -90
rect 681 -91 682 -90
rect 709 -91 710 -90
rect 842 -91 843 -90
rect 401 -93 402 -92
rect 569 -93 570 -92
rect 576 -93 577 -92
rect 597 -93 598 -92
rect 611 -93 612 -92
rect 723 -93 724 -92
rect 366 -95 367 -94
rect 401 -95 402 -94
rect 443 -95 444 -94
rect 611 -95 612 -94
rect 646 -95 647 -94
rect 758 -95 759 -94
rect 359 -97 360 -96
rect 646 -97 647 -96
rect 653 -97 654 -96
rect 751 -97 752 -96
rect 226 -99 227 -98
rect 359 -99 360 -98
rect 436 -99 437 -98
rect 443 -99 444 -98
rect 520 -99 521 -98
rect 653 -99 654 -98
rect 660 -99 661 -98
rect 765 -99 766 -98
rect 177 -101 178 -100
rect 226 -101 227 -100
rect 310 -101 311 -100
rect 520 -101 521 -100
rect 534 -101 535 -100
rect 639 -101 640 -100
rect 667 -101 668 -100
rect 800 -101 801 -100
rect 156 -103 157 -102
rect 667 -103 668 -102
rect 177 -105 178 -104
rect 212 -105 213 -104
rect 310 -105 311 -104
rect 341 -105 342 -104
rect 415 -105 416 -104
rect 436 -105 437 -104
rect 499 -105 500 -104
rect 534 -105 535 -104
rect 541 -105 542 -104
rect 604 -105 605 -104
rect 191 -107 192 -106
rect 212 -107 213 -106
rect 422 -107 423 -106
rect 541 -107 542 -106
rect 562 -107 563 -106
rect 576 -107 577 -106
rect 47 -109 48 -108
rect 422 -109 423 -108
rect 191 -111 192 -110
rect 390 -111 391 -110
rect 296 -113 297 -112
rect 562 -113 563 -112
rect 275 -115 276 -114
rect 296 -115 297 -114
rect 184 -117 185 -116
rect 275 -117 276 -116
rect 135 -119 136 -118
rect 184 -119 185 -118
rect 135 -121 136 -120
rect 366 -121 367 -120
rect 23 -132 24 -131
rect 121 -132 122 -131
rect 128 -132 129 -131
rect 208 -132 209 -131
rect 226 -132 227 -131
rect 688 -132 689 -131
rect 723 -132 724 -131
rect 863 -132 864 -131
rect 870 -132 871 -131
rect 954 -132 955 -131
rect 30 -134 31 -133
rect 135 -134 136 -133
rect 145 -134 146 -133
rect 415 -134 416 -133
rect 499 -134 500 -133
rect 639 -134 640 -133
rect 751 -134 752 -133
rect 870 -134 871 -133
rect 877 -134 878 -133
rect 912 -134 913 -133
rect 30 -136 31 -135
rect 163 -136 164 -135
rect 170 -136 171 -135
rect 828 -136 829 -135
rect 37 -138 38 -137
rect 100 -138 101 -137
rect 149 -138 150 -137
rect 177 -138 178 -137
rect 250 -138 251 -137
rect 835 -138 836 -137
rect 37 -140 38 -139
rect 205 -140 206 -139
rect 275 -140 276 -139
rect 310 -140 311 -139
rect 317 -140 318 -139
rect 492 -140 493 -139
rect 509 -140 510 -139
rect 737 -140 738 -139
rect 765 -140 766 -139
rect 891 -140 892 -139
rect 44 -142 45 -141
rect 142 -142 143 -141
rect 156 -142 157 -141
rect 821 -142 822 -141
rect 51 -144 52 -143
rect 275 -144 276 -143
rect 299 -144 300 -143
rect 352 -144 353 -143
rect 362 -144 363 -143
rect 919 -144 920 -143
rect 51 -146 52 -145
rect 124 -146 125 -145
rect 142 -146 143 -145
rect 373 -146 374 -145
rect 376 -146 377 -145
rect 569 -146 570 -145
rect 579 -146 580 -145
rect 758 -146 759 -145
rect 772 -146 773 -145
rect 905 -146 906 -145
rect 58 -148 59 -147
rect 646 -148 647 -147
rect 660 -148 661 -147
rect 758 -148 759 -147
rect 779 -148 780 -147
rect 884 -148 885 -147
rect 65 -150 66 -149
rect 114 -150 115 -149
rect 117 -150 118 -149
rect 156 -150 157 -149
rect 159 -150 160 -149
rect 348 -150 349 -149
rect 352 -150 353 -149
rect 541 -150 542 -149
rect 548 -150 549 -149
rect 849 -150 850 -149
rect 79 -152 80 -151
rect 674 -152 675 -151
rect 681 -152 682 -151
rect 779 -152 780 -151
rect 786 -152 787 -151
rect 926 -152 927 -151
rect 79 -154 80 -153
rect 152 -154 153 -153
rect 163 -154 164 -153
rect 198 -154 199 -153
rect 310 -154 311 -153
rect 471 -154 472 -153
rect 495 -154 496 -153
rect 660 -154 661 -153
rect 667 -154 668 -153
rect 765 -154 766 -153
rect 793 -154 794 -153
rect 933 -154 934 -153
rect 86 -156 87 -155
rect 397 -156 398 -155
rect 418 -156 419 -155
rect 639 -156 640 -155
rect 695 -156 696 -155
rect 821 -156 822 -155
rect 89 -158 90 -157
rect 128 -158 129 -157
rect 152 -158 153 -157
rect 856 -158 857 -157
rect 114 -160 115 -159
rect 180 -160 181 -159
rect 198 -160 199 -159
rect 212 -160 213 -159
rect 317 -160 318 -159
rect 408 -160 409 -159
rect 422 -160 423 -159
rect 499 -160 500 -159
rect 513 -160 514 -159
rect 541 -160 542 -159
rect 583 -160 584 -159
rect 898 -160 899 -159
rect 170 -162 171 -161
rect 215 -162 216 -161
rect 320 -162 321 -161
rect 401 -162 402 -161
rect 429 -162 430 -161
rect 513 -162 514 -161
rect 520 -162 521 -161
rect 548 -162 549 -161
rect 583 -162 584 -161
rect 730 -162 731 -161
rect 737 -162 738 -161
rect 877 -162 878 -161
rect 173 -164 174 -163
rect 457 -164 458 -163
rect 464 -164 465 -163
rect 471 -164 472 -163
rect 492 -164 493 -163
rect 695 -164 696 -163
rect 702 -164 703 -163
rect 772 -164 773 -163
rect 800 -164 801 -163
rect 940 -164 941 -163
rect 212 -166 213 -165
rect 303 -166 304 -165
rect 324 -166 325 -165
rect 355 -166 356 -165
rect 359 -166 360 -165
rect 408 -166 409 -165
rect 443 -166 444 -165
rect 786 -166 787 -165
rect 814 -166 815 -165
rect 947 -166 948 -165
rect 65 -168 66 -167
rect 359 -168 360 -167
rect 380 -168 381 -167
rect 464 -168 465 -167
rect 506 -168 507 -167
rect 800 -168 801 -167
rect 93 -170 94 -169
rect 380 -170 381 -169
rect 387 -170 388 -169
rect 429 -170 430 -169
rect 520 -170 521 -169
rect 835 -170 836 -169
rect 93 -172 94 -171
rect 184 -172 185 -171
rect 219 -172 220 -171
rect 303 -172 304 -171
rect 324 -172 325 -171
rect 688 -172 689 -171
rect 709 -172 710 -171
rect 751 -172 752 -171
rect 135 -174 136 -173
rect 219 -174 220 -173
rect 261 -174 262 -173
rect 506 -174 507 -173
rect 523 -174 524 -173
rect 723 -174 724 -173
rect 107 -176 108 -175
rect 261 -176 262 -175
rect 327 -176 328 -175
rect 338 -176 339 -175
rect 345 -176 346 -175
rect 422 -176 423 -175
rect 534 -176 535 -175
rect 569 -176 570 -175
rect 590 -176 591 -175
rect 646 -176 647 -175
rect 716 -176 717 -175
rect 828 -176 829 -175
rect 184 -178 185 -177
rect 191 -178 192 -177
rect 268 -178 269 -177
rect 338 -178 339 -177
rect 348 -178 349 -177
rect 527 -178 528 -177
rect 597 -178 598 -177
rect 730 -178 731 -177
rect 72 -180 73 -179
rect 597 -180 598 -179
rect 611 -180 612 -179
rect 667 -180 668 -179
rect 72 -182 73 -181
rect 702 -182 703 -181
rect 191 -184 192 -183
rect 229 -184 230 -183
rect 268 -184 269 -183
rect 289 -184 290 -183
rect 331 -184 332 -183
rect 443 -184 444 -183
rect 450 -184 451 -183
rect 534 -184 535 -183
rect 555 -184 556 -183
rect 611 -184 612 -183
rect 618 -184 619 -183
rect 709 -184 710 -183
rect 205 -186 206 -185
rect 289 -186 290 -185
rect 334 -186 335 -185
rect 842 -186 843 -185
rect 366 -188 367 -187
rect 450 -188 451 -187
rect 478 -188 479 -187
rect 555 -188 556 -187
rect 618 -188 619 -187
rect 842 -188 843 -187
rect 296 -190 297 -189
rect 366 -190 367 -189
rect 394 -190 395 -189
rect 681 -190 682 -189
rect 282 -192 283 -191
rect 394 -192 395 -191
rect 401 -192 402 -191
rect 674 -192 675 -191
rect 240 -194 241 -193
rect 282 -194 283 -193
rect 296 -194 297 -193
rect 590 -194 591 -193
rect 625 -194 626 -193
rect 793 -194 794 -193
rect 240 -196 241 -195
rect 254 -196 255 -195
rect 478 -196 479 -195
rect 562 -196 563 -195
rect 625 -196 626 -195
rect 814 -196 815 -195
rect 233 -198 234 -197
rect 254 -198 255 -197
rect 345 -198 346 -197
rect 562 -198 563 -197
rect 632 -198 633 -197
rect 716 -198 717 -197
rect 58 -200 59 -199
rect 233 -200 234 -199
rect 485 -200 486 -199
rect 527 -200 528 -199
rect 604 -200 605 -199
rect 632 -200 633 -199
rect 110 -202 111 -201
rect 485 -202 486 -201
rect 576 -202 577 -201
rect 604 -202 605 -201
rect 576 -204 577 -203
rect 744 -204 745 -203
rect 653 -206 654 -205
rect 744 -206 745 -205
rect 653 -208 654 -207
rect 807 -208 808 -207
rect 656 -210 657 -209
rect 807 -210 808 -209
rect 16 -221 17 -220
rect 702 -221 703 -220
rect 723 -221 724 -220
rect 908 -221 909 -220
rect 23 -223 24 -222
rect 208 -223 209 -222
rect 261 -223 262 -222
rect 345 -223 346 -222
rect 352 -223 353 -222
rect 387 -223 388 -222
rect 401 -223 402 -222
rect 828 -223 829 -222
rect 887 -223 888 -222
rect 912 -223 913 -222
rect 23 -225 24 -224
rect 79 -225 80 -224
rect 114 -225 115 -224
rect 233 -225 234 -224
rect 254 -225 255 -224
rect 387 -225 388 -224
rect 471 -225 472 -224
rect 492 -225 493 -224
rect 495 -225 496 -224
rect 905 -225 906 -224
rect 30 -227 31 -226
rect 362 -227 363 -226
rect 366 -227 367 -226
rect 404 -227 405 -226
rect 502 -227 503 -226
rect 555 -227 556 -226
rect 579 -227 580 -226
rect 926 -227 927 -226
rect 30 -229 31 -228
rect 156 -229 157 -228
rect 163 -229 164 -228
rect 222 -229 223 -228
rect 296 -229 297 -228
rect 394 -229 395 -228
rect 555 -229 556 -228
rect 611 -229 612 -228
rect 618 -229 619 -228
rect 863 -229 864 -228
rect 44 -231 45 -230
rect 138 -231 139 -230
rect 142 -231 143 -230
rect 534 -231 535 -230
rect 611 -231 612 -230
rect 667 -231 668 -230
rect 674 -231 675 -230
rect 905 -231 906 -230
rect 51 -233 52 -232
rect 254 -233 255 -232
rect 299 -233 300 -232
rect 401 -233 402 -232
rect 621 -233 622 -232
rect 898 -233 899 -232
rect 51 -235 52 -234
rect 58 -235 59 -234
rect 65 -235 66 -234
rect 261 -235 262 -234
rect 299 -235 300 -234
rect 408 -235 409 -234
rect 618 -235 619 -234
rect 898 -235 899 -234
rect 58 -237 59 -236
rect 467 -237 468 -236
rect 625 -237 626 -236
rect 660 -237 661 -236
rect 663 -237 664 -236
rect 667 -237 668 -236
rect 674 -237 675 -236
rect 688 -237 689 -236
rect 702 -237 703 -236
rect 779 -237 780 -236
rect 807 -237 808 -236
rect 863 -237 864 -236
rect 65 -239 66 -238
rect 107 -239 108 -238
rect 121 -239 122 -238
rect 562 -239 563 -238
rect 628 -239 629 -238
rect 933 -239 934 -238
rect 68 -241 69 -240
rect 366 -241 367 -240
rect 408 -241 409 -240
rect 436 -241 437 -240
rect 541 -241 542 -240
rect 562 -241 563 -240
rect 639 -241 640 -240
rect 912 -241 913 -240
rect 72 -243 73 -242
rect 303 -243 304 -242
rect 317 -243 318 -242
rect 471 -243 472 -242
rect 541 -243 542 -242
rect 548 -243 549 -242
rect 597 -243 598 -242
rect 639 -243 640 -242
rect 653 -243 654 -242
rect 947 -243 948 -242
rect 72 -245 73 -244
rect 338 -245 339 -244
rect 359 -245 360 -244
rect 478 -245 479 -244
rect 527 -245 528 -244
rect 548 -245 549 -244
rect 597 -245 598 -244
rect 709 -245 710 -244
rect 723 -245 724 -244
rect 730 -245 731 -244
rect 737 -245 738 -244
rect 744 -245 745 -244
rect 800 -245 801 -244
rect 807 -245 808 -244
rect 828 -245 829 -244
rect 884 -245 885 -244
rect 79 -247 80 -246
rect 114 -247 115 -246
rect 121 -247 122 -246
rect 170 -247 171 -246
rect 177 -247 178 -246
rect 275 -247 276 -246
rect 289 -247 290 -246
rect 303 -247 304 -246
rect 317 -247 318 -246
rect 534 -247 535 -246
rect 653 -247 654 -246
rect 716 -247 717 -246
rect 730 -247 731 -246
rect 772 -247 773 -246
rect 93 -249 94 -248
rect 275 -249 276 -248
rect 324 -249 325 -248
rect 849 -249 850 -248
rect 100 -251 101 -250
rect 156 -251 157 -250
rect 170 -251 171 -250
rect 856 -251 857 -250
rect 100 -253 101 -252
rect 149 -253 150 -252
rect 173 -253 174 -252
rect 289 -253 290 -252
rect 324 -253 325 -252
rect 520 -253 521 -252
rect 688 -253 689 -252
rect 751 -253 752 -252
rect 814 -253 815 -252
rect 849 -253 850 -252
rect 856 -253 857 -252
rect 919 -253 920 -252
rect 117 -255 118 -254
rect 149 -255 150 -254
rect 177 -255 178 -254
rect 184 -255 185 -254
rect 194 -255 195 -254
rect 506 -255 507 -254
rect 695 -255 696 -254
rect 800 -255 801 -254
rect 814 -255 815 -254
rect 835 -255 836 -254
rect 919 -255 920 -254
rect 954 -255 955 -254
rect 93 -257 94 -256
rect 184 -257 185 -256
rect 198 -257 199 -256
rect 226 -257 227 -256
rect 240 -257 241 -256
rect 695 -257 696 -256
rect 709 -257 710 -256
rect 758 -257 759 -256
rect 37 -259 38 -258
rect 240 -259 241 -258
rect 331 -259 332 -258
rect 464 -259 465 -258
rect 485 -259 486 -258
rect 772 -259 773 -258
rect 37 -261 38 -260
rect 247 -261 248 -260
rect 331 -261 332 -260
rect 569 -261 570 -260
rect 740 -261 741 -260
rect 779 -261 780 -260
rect 47 -263 48 -262
rect 198 -263 199 -262
rect 219 -263 220 -262
rect 478 -263 479 -262
rect 485 -263 486 -262
rect 940 -263 941 -262
rect 135 -265 136 -264
rect 166 -265 167 -264
rect 219 -265 220 -264
rect 229 -265 230 -264
rect 247 -265 248 -264
rect 268 -265 269 -264
rect 338 -265 339 -264
rect 380 -265 381 -264
rect 397 -265 398 -264
rect 835 -265 836 -264
rect 86 -267 87 -266
rect 135 -267 136 -266
rect 142 -267 143 -266
rect 212 -267 213 -266
rect 282 -267 283 -266
rect 380 -267 381 -266
rect 436 -267 437 -266
rect 786 -267 787 -266
rect 128 -269 129 -268
rect 268 -269 269 -268
rect 282 -269 283 -268
rect 355 -269 356 -268
rect 362 -269 363 -268
rect 590 -269 591 -268
rect 744 -269 745 -268
rect 765 -269 766 -268
rect 191 -271 192 -270
rect 212 -271 213 -270
rect 450 -271 451 -270
rect 527 -271 528 -270
rect 583 -271 584 -270
rect 786 -271 787 -270
rect 191 -273 192 -272
rect 429 -273 430 -272
rect 443 -273 444 -272
rect 583 -273 584 -272
rect 590 -273 591 -272
rect 632 -273 633 -272
rect 751 -273 752 -272
rect 821 -273 822 -272
rect 334 -275 335 -274
rect 429 -275 430 -274
rect 488 -275 489 -274
rect 716 -275 717 -274
rect 758 -275 759 -274
rect 793 -275 794 -274
rect 821 -275 822 -274
rect 842 -275 843 -274
rect 415 -277 416 -276
rect 443 -277 444 -276
rect 506 -277 507 -276
rect 513 -277 514 -276
rect 632 -277 633 -276
rect 681 -277 682 -276
rect 793 -277 794 -276
rect 870 -277 871 -276
rect 152 -279 153 -278
rect 513 -279 514 -278
rect 842 -279 843 -278
rect 877 -279 878 -278
rect 257 -281 258 -280
rect 681 -281 682 -280
rect 870 -281 871 -280
rect 891 -281 892 -280
rect 310 -283 311 -282
rect 415 -283 416 -282
rect 422 -283 423 -282
rect 450 -283 451 -282
rect 576 -283 577 -282
rect 877 -283 878 -282
rect 310 -285 311 -284
rect 520 -285 521 -284
rect 373 -287 374 -286
rect 422 -287 423 -286
rect 457 -287 458 -286
rect 576 -287 577 -286
rect 373 -289 374 -288
rect 765 -289 766 -288
rect 457 -291 458 -290
rect 499 -291 500 -290
rect 499 -293 500 -292
rect 569 -293 570 -292
rect 16 -304 17 -303
rect 184 -304 185 -303
rect 240 -304 241 -303
rect 474 -304 475 -303
rect 492 -304 493 -303
rect 520 -304 521 -303
rect 523 -304 524 -303
rect 856 -304 857 -303
rect 863 -304 864 -303
rect 905 -304 906 -303
rect 23 -306 24 -305
rect 100 -306 101 -305
rect 110 -306 111 -305
rect 121 -306 122 -305
rect 124 -306 125 -305
rect 131 -306 132 -305
rect 159 -306 160 -305
rect 250 -306 251 -305
rect 254 -306 255 -305
rect 387 -306 388 -305
rect 394 -306 395 -305
rect 884 -306 885 -305
rect 898 -306 899 -305
rect 912 -306 913 -305
rect 23 -308 24 -307
rect 208 -308 209 -307
rect 233 -308 234 -307
rect 240 -308 241 -307
rect 247 -308 248 -307
rect 320 -308 321 -307
rect 352 -308 353 -307
rect 467 -308 468 -307
rect 544 -308 545 -307
rect 653 -308 654 -307
rect 660 -308 661 -307
rect 744 -308 745 -307
rect 800 -308 801 -307
rect 880 -308 881 -307
rect 30 -310 31 -309
rect 352 -310 353 -309
rect 355 -310 356 -309
rect 506 -310 507 -309
rect 516 -310 517 -309
rect 744 -310 745 -309
rect 835 -310 836 -309
rect 887 -310 888 -309
rect 37 -312 38 -311
rect 96 -312 97 -311
rect 100 -312 101 -311
rect 198 -312 199 -311
rect 233 -312 234 -311
rect 628 -312 629 -311
rect 681 -312 682 -311
rect 933 -312 934 -311
rect 37 -314 38 -313
rect 299 -314 300 -313
rect 306 -314 307 -313
rect 800 -314 801 -313
rect 807 -314 808 -313
rect 835 -314 836 -313
rect 863 -314 864 -313
rect 870 -314 871 -313
rect 877 -314 878 -313
rect 891 -314 892 -313
rect 44 -316 45 -315
rect 103 -316 104 -315
rect 117 -316 118 -315
rect 156 -316 157 -315
rect 170 -316 171 -315
rect 541 -316 542 -315
rect 625 -316 626 -315
rect 653 -316 654 -315
rect 786 -316 787 -315
rect 870 -316 871 -315
rect 877 -316 878 -315
rect 919 -316 920 -315
rect 47 -318 48 -317
rect 555 -318 556 -317
rect 646 -318 647 -317
rect 681 -318 682 -317
rect 716 -318 717 -317
rect 786 -318 787 -317
rect 793 -318 794 -317
rect 807 -318 808 -317
rect 58 -320 59 -319
rect 401 -320 402 -319
rect 422 -320 423 -319
rect 488 -320 489 -319
rect 541 -320 542 -319
rect 723 -320 724 -319
rect 730 -320 731 -319
rect 793 -320 794 -319
rect 58 -322 59 -321
rect 86 -322 87 -321
rect 128 -322 129 -321
rect 135 -322 136 -321
rect 149 -322 150 -321
rect 198 -322 199 -321
rect 268 -322 269 -321
rect 499 -322 500 -321
rect 576 -322 577 -321
rect 716 -322 717 -321
rect 65 -324 66 -323
rect 373 -324 374 -323
rect 439 -324 440 -323
rect 737 -324 738 -323
rect 9 -326 10 -325
rect 65 -326 66 -325
rect 68 -326 69 -325
rect 751 -326 752 -325
rect 68 -328 69 -327
rect 86 -328 87 -327
rect 128 -328 129 -327
rect 163 -328 164 -327
rect 173 -328 174 -327
rect 639 -328 640 -327
rect 702 -328 703 -327
rect 751 -328 752 -327
rect 79 -330 80 -329
rect 114 -330 115 -329
rect 135 -330 136 -329
rect 723 -330 724 -329
rect 79 -332 80 -331
rect 849 -332 850 -331
rect 82 -334 83 -333
rect 506 -334 507 -333
rect 527 -334 528 -333
rect 576 -334 577 -333
rect 597 -334 598 -333
rect 730 -334 731 -333
rect 842 -334 843 -333
rect 849 -334 850 -333
rect 149 -336 150 -335
rect 219 -336 220 -335
rect 268 -336 269 -335
rect 275 -336 276 -335
rect 296 -336 297 -335
rect 443 -336 444 -335
rect 464 -336 465 -335
rect 772 -336 773 -335
rect 16 -338 17 -337
rect 219 -338 220 -337
rect 275 -338 276 -337
rect 485 -338 486 -337
rect 513 -338 514 -337
rect 527 -338 528 -337
rect 583 -338 584 -337
rect 597 -338 598 -337
rect 618 -338 619 -337
rect 639 -338 640 -337
rect 674 -338 675 -337
rect 702 -338 703 -337
rect 709 -338 710 -337
rect 737 -338 738 -337
rect 772 -338 773 -337
rect 779 -338 780 -337
rect 163 -340 164 -339
rect 187 -340 188 -339
rect 191 -340 192 -339
rect 401 -340 402 -339
rect 404 -340 405 -339
rect 618 -340 619 -339
rect 667 -340 668 -339
rect 674 -340 675 -339
rect 688 -340 689 -339
rect 842 -340 843 -339
rect 170 -342 171 -341
rect 191 -342 192 -341
rect 205 -342 206 -341
rect 583 -342 584 -341
rect 709 -342 710 -341
rect 894 -342 895 -341
rect 173 -344 174 -343
rect 331 -344 332 -343
rect 345 -344 346 -343
rect 688 -344 689 -343
rect 779 -344 780 -343
rect 828 -344 829 -343
rect 72 -346 73 -345
rect 345 -346 346 -345
rect 359 -346 360 -345
rect 670 -346 671 -345
rect 814 -346 815 -345
rect 828 -346 829 -345
rect 72 -348 73 -347
rect 121 -348 122 -347
rect 205 -348 206 -347
rect 215 -348 216 -347
rect 289 -348 290 -347
rect 296 -348 297 -347
rect 310 -348 311 -347
rect 387 -348 388 -347
rect 408 -348 409 -347
rect 485 -348 486 -347
rect 513 -348 514 -347
rect 590 -348 591 -347
rect 814 -348 815 -347
rect 821 -348 822 -347
rect 194 -350 195 -349
rect 821 -350 822 -349
rect 226 -352 227 -351
rect 289 -352 290 -351
rect 310 -352 311 -351
rect 415 -352 416 -351
rect 443 -352 444 -351
rect 695 -352 696 -351
rect 212 -354 213 -353
rect 226 -354 227 -353
rect 247 -354 248 -353
rect 415 -354 416 -353
rect 450 -354 451 -353
rect 464 -354 465 -353
rect 471 -354 472 -353
rect 646 -354 647 -353
rect 257 -356 258 -355
rect 408 -356 409 -355
rect 562 -356 563 -355
rect 590 -356 591 -355
rect 632 -356 633 -355
rect 695 -356 696 -355
rect 264 -358 265 -357
rect 562 -358 563 -357
rect 604 -358 605 -357
rect 632 -358 633 -357
rect 282 -360 283 -359
rect 450 -360 451 -359
rect 142 -362 143 -361
rect 282 -362 283 -361
rect 317 -362 318 -361
rect 611 -362 612 -361
rect 107 -364 108 -363
rect 142 -364 143 -363
rect 320 -364 321 -363
rect 422 -364 423 -363
rect 429 -364 430 -363
rect 604 -364 605 -363
rect 107 -366 108 -365
rect 856 -366 857 -365
rect 324 -368 325 -367
rect 429 -368 430 -367
rect 534 -368 535 -367
rect 611 -368 612 -367
rect 324 -370 325 -369
rect 765 -370 766 -369
rect 331 -372 332 -371
rect 884 -372 885 -371
rect 341 -374 342 -373
rect 359 -374 360 -373
rect 366 -374 367 -373
rect 555 -374 556 -373
rect 758 -374 759 -373
rect 765 -374 766 -373
rect 303 -376 304 -375
rect 366 -376 367 -375
rect 373 -376 374 -375
rect 457 -376 458 -375
rect 534 -376 535 -375
rect 569 -376 570 -375
rect 51 -378 52 -377
rect 303 -378 304 -377
rect 338 -378 339 -377
rect 457 -378 458 -377
rect 548 -378 549 -377
rect 569 -378 570 -377
rect 51 -380 52 -379
rect 93 -380 94 -379
rect 380 -380 381 -379
rect 548 -380 549 -379
rect 436 -382 437 -381
rect 758 -382 759 -381
rect 397 -384 398 -383
rect 436 -384 437 -383
rect 397 -386 398 -385
rect 478 -386 479 -385
rect 166 -388 167 -387
rect 478 -388 479 -387
rect 2 -399 3 -398
rect 579 -399 580 -398
rect 611 -399 612 -398
rect 996 -399 997 -398
rect 1108 -399 1109 -398
rect 1115 -399 1116 -398
rect 9 -401 10 -400
rect 30 -401 31 -400
rect 44 -401 45 -400
rect 138 -401 139 -400
rect 145 -401 146 -400
rect 443 -401 444 -400
rect 474 -401 475 -400
rect 842 -401 843 -400
rect 849 -401 850 -400
rect 975 -401 976 -400
rect 982 -401 983 -400
rect 1031 -401 1032 -400
rect 16 -403 17 -402
rect 100 -403 101 -402
rect 107 -403 108 -402
rect 331 -403 332 -402
rect 338 -403 339 -402
rect 366 -403 367 -402
rect 380 -403 381 -402
rect 513 -403 514 -402
rect 569 -403 570 -402
rect 611 -403 612 -402
rect 628 -403 629 -402
rect 870 -403 871 -402
rect 884 -403 885 -402
rect 898 -403 899 -402
rect 933 -403 934 -402
rect 1045 -403 1046 -402
rect 23 -405 24 -404
rect 156 -405 157 -404
rect 170 -405 171 -404
rect 800 -405 801 -404
rect 807 -405 808 -404
rect 954 -405 955 -404
rect 989 -405 990 -404
rect 1038 -405 1039 -404
rect 23 -407 24 -406
rect 51 -407 52 -406
rect 58 -407 59 -406
rect 366 -407 367 -406
rect 380 -407 381 -406
rect 506 -407 507 -406
rect 569 -407 570 -406
rect 821 -407 822 -406
rect 828 -407 829 -406
rect 926 -407 927 -406
rect 37 -409 38 -408
rect 331 -409 332 -408
rect 341 -409 342 -408
rect 401 -409 402 -408
rect 422 -409 423 -408
rect 443 -409 444 -408
rect 474 -409 475 -408
rect 1024 -409 1025 -408
rect 44 -411 45 -410
rect 275 -411 276 -410
rect 296 -411 297 -410
rect 303 -411 304 -410
rect 306 -411 307 -410
rect 807 -411 808 -410
rect 863 -411 864 -410
rect 1010 -411 1011 -410
rect 51 -413 52 -412
rect 310 -413 311 -412
rect 327 -413 328 -412
rect 688 -413 689 -412
rect 702 -413 703 -412
rect 828 -413 829 -412
rect 835 -413 836 -412
rect 863 -413 864 -412
rect 891 -413 892 -412
rect 1017 -413 1018 -412
rect 65 -415 66 -414
rect 583 -415 584 -414
rect 625 -415 626 -414
rect 933 -415 934 -414
rect 79 -417 80 -416
rect 352 -417 353 -416
rect 383 -417 384 -416
rect 548 -417 549 -416
rect 572 -417 573 -416
rect 961 -417 962 -416
rect 79 -419 80 -418
rect 128 -419 129 -418
rect 135 -419 136 -418
rect 520 -419 521 -418
rect 576 -419 577 -418
rect 625 -419 626 -418
rect 635 -419 636 -418
rect 793 -419 794 -418
rect 814 -419 815 -418
rect 891 -419 892 -418
rect 82 -421 83 -420
rect 702 -421 703 -420
rect 709 -421 710 -420
rect 800 -421 801 -420
rect 96 -423 97 -422
rect 821 -423 822 -422
rect 100 -425 101 -424
rect 422 -425 423 -424
rect 478 -425 479 -424
rect 583 -425 584 -424
rect 632 -425 633 -424
rect 709 -425 710 -424
rect 723 -425 724 -424
rect 842 -425 843 -424
rect 114 -427 115 -426
rect 471 -427 472 -426
rect 485 -427 486 -426
rect 548 -427 549 -426
rect 576 -427 577 -426
rect 849 -427 850 -426
rect 117 -429 118 -428
rect 856 -429 857 -428
rect 121 -431 122 -430
rect 387 -431 388 -430
rect 397 -431 398 -430
rect 646 -431 647 -430
rect 667 -431 668 -430
rect 856 -431 857 -430
rect 86 -433 87 -432
rect 387 -433 388 -432
rect 401 -433 402 -432
rect 499 -433 500 -432
rect 506 -433 507 -432
rect 558 -433 559 -432
rect 590 -433 591 -432
rect 646 -433 647 -432
rect 667 -433 668 -432
rect 751 -433 752 -432
rect 765 -433 766 -432
rect 898 -433 899 -432
rect 72 -435 73 -434
rect 86 -435 87 -434
rect 121 -435 122 -434
rect 163 -435 164 -434
rect 170 -435 171 -434
rect 261 -435 262 -434
rect 264 -435 265 -434
rect 562 -435 563 -434
rect 590 -435 591 -434
rect 604 -435 605 -434
rect 681 -435 682 -434
rect 765 -435 766 -434
rect 772 -435 773 -434
rect 912 -435 913 -434
rect 72 -437 73 -436
rect 131 -437 132 -436
rect 149 -437 150 -436
rect 163 -437 164 -436
rect 184 -437 185 -436
rect 618 -437 619 -436
rect 639 -437 640 -436
rect 772 -437 773 -436
rect 786 -437 787 -436
rect 947 -437 948 -436
rect 61 -439 62 -438
rect 618 -439 619 -438
rect 653 -439 654 -438
rect 786 -439 787 -438
rect 149 -441 150 -440
rect 373 -441 374 -440
rect 408 -441 409 -440
rect 520 -441 521 -440
rect 534 -441 535 -440
rect 604 -441 605 -440
rect 688 -441 689 -440
rect 870 -441 871 -440
rect 12 -443 13 -442
rect 408 -443 409 -442
rect 429 -443 430 -442
rect 485 -443 486 -442
rect 492 -443 493 -442
rect 919 -443 920 -442
rect 156 -445 157 -444
rect 177 -445 178 -444
rect 184 -445 185 -444
rect 191 -445 192 -444
rect 198 -445 199 -444
rect 261 -445 262 -444
rect 268 -445 269 -444
rect 320 -445 321 -444
rect 327 -445 328 -444
rect 457 -445 458 -444
rect 460 -445 461 -444
rect 751 -445 752 -444
rect 177 -447 178 -446
rect 212 -447 213 -446
rect 219 -447 220 -446
rect 296 -447 297 -446
rect 352 -447 353 -446
rect 1003 -447 1004 -446
rect 180 -449 181 -448
rect 219 -449 220 -448
rect 233 -449 234 -448
rect 310 -449 311 -448
rect 373 -449 374 -448
rect 527 -449 528 -448
rect 534 -449 535 -448
rect 660 -449 661 -448
rect 716 -449 717 -448
rect 723 -449 724 -448
rect 730 -449 731 -448
rect 884 -449 885 -448
rect 187 -451 188 -450
rect 415 -451 416 -450
rect 425 -451 426 -450
rect 660 -451 661 -450
rect 695 -451 696 -450
rect 730 -451 731 -450
rect 737 -451 738 -450
rect 968 -451 969 -450
rect 191 -453 192 -452
rect 877 -453 878 -452
rect 198 -455 199 -454
rect 226 -455 227 -454
rect 233 -455 234 -454
rect 394 -455 395 -454
rect 429 -455 430 -454
rect 436 -455 437 -454
rect 450 -455 451 -454
rect 527 -455 528 -454
rect 597 -455 598 -454
rect 716 -455 717 -454
rect 744 -455 745 -454
rect 835 -455 836 -454
rect 205 -457 206 -456
rect 226 -457 227 -456
rect 247 -457 248 -456
rect 268 -457 269 -456
rect 275 -457 276 -456
rect 502 -457 503 -456
rect 516 -457 517 -456
rect 737 -457 738 -456
rect 758 -457 759 -456
rect 877 -457 878 -456
rect 93 -459 94 -458
rect 205 -459 206 -458
rect 240 -459 241 -458
rect 247 -459 248 -458
rect 250 -459 251 -458
rect 289 -459 290 -458
rect 317 -459 318 -458
rect 436 -459 437 -458
rect 457 -459 458 -458
rect 940 -459 941 -458
rect 93 -461 94 -460
rect 124 -461 125 -460
rect 142 -461 143 -460
rect 240 -461 241 -460
rect 254 -461 255 -460
rect 1034 -461 1035 -460
rect 68 -463 69 -462
rect 254 -463 255 -462
rect 282 -463 283 -462
rect 383 -463 384 -462
rect 481 -463 482 -462
rect 653 -463 654 -462
rect 674 -463 675 -462
rect 744 -463 745 -462
rect 110 -465 111 -464
rect 317 -465 318 -464
rect 359 -465 360 -464
rect 450 -465 451 -464
rect 495 -465 496 -464
rect 793 -465 794 -464
rect 142 -467 143 -466
rect 681 -467 682 -466
rect 695 -467 696 -466
rect 779 -467 780 -466
rect 173 -469 174 -468
rect 289 -469 290 -468
rect 345 -469 346 -468
rect 359 -469 360 -468
rect 499 -469 500 -468
rect 597 -469 598 -468
rect 30 -471 31 -470
rect 345 -471 346 -470
rect 541 -471 542 -470
rect 674 -471 675 -470
rect 324 -473 325 -472
rect 541 -473 542 -472
rect 544 -473 545 -472
rect 758 -473 759 -472
rect 37 -475 38 -474
rect 324 -475 325 -474
rect 555 -475 556 -474
rect 779 -475 780 -474
rect 492 -477 493 -476
rect 555 -477 556 -476
rect 9 -488 10 -487
rect 632 -488 633 -487
rect 814 -488 815 -487
rect 1031 -488 1032 -487
rect 1111 -488 1112 -487
rect 1122 -488 1123 -487
rect 30 -490 31 -489
rect 33 -490 34 -489
rect 44 -490 45 -489
rect 282 -490 283 -489
rect 285 -490 286 -489
rect 618 -490 619 -489
rect 765 -490 766 -489
rect 814 -490 815 -489
rect 817 -490 818 -489
rect 835 -490 836 -489
rect 954 -490 955 -489
rect 1038 -490 1039 -489
rect 1115 -490 1116 -489
rect 1129 -490 1130 -489
rect 23 -492 24 -491
rect 618 -492 619 -491
rect 772 -492 773 -491
rect 835 -492 836 -491
rect 975 -492 976 -491
rect 1052 -492 1053 -491
rect 30 -494 31 -493
rect 212 -494 213 -493
rect 296 -494 297 -493
rect 355 -494 356 -493
rect 373 -494 374 -493
rect 530 -494 531 -493
rect 555 -494 556 -493
rect 912 -494 913 -493
rect 1010 -494 1011 -493
rect 1059 -494 1060 -493
rect 33 -496 34 -495
rect 212 -496 213 -495
rect 296 -496 297 -495
rect 310 -496 311 -495
rect 317 -496 318 -495
rect 1073 -496 1074 -495
rect 37 -498 38 -497
rect 282 -498 283 -497
rect 310 -498 311 -497
rect 492 -498 493 -497
rect 499 -498 500 -497
rect 551 -498 552 -497
rect 565 -498 566 -497
rect 968 -498 969 -497
rect 1017 -498 1018 -497
rect 1066 -498 1067 -497
rect 44 -500 45 -499
rect 401 -500 402 -499
rect 415 -500 416 -499
rect 765 -500 766 -499
rect 842 -500 843 -499
rect 1017 -500 1018 -499
rect 1024 -500 1025 -499
rect 1094 -500 1095 -499
rect 16 -502 17 -501
rect 415 -502 416 -501
rect 422 -502 423 -501
rect 604 -502 605 -501
rect 709 -502 710 -501
rect 772 -502 773 -501
rect 863 -502 864 -501
rect 975 -502 976 -501
rect 1045 -502 1046 -501
rect 1115 -502 1116 -501
rect 16 -504 17 -503
rect 352 -504 353 -503
rect 359 -504 360 -503
rect 373 -504 374 -503
rect 397 -504 398 -503
rect 807 -504 808 -503
rect 926 -504 927 -503
rect 968 -504 969 -503
rect 982 -504 983 -503
rect 1045 -504 1046 -503
rect 58 -506 59 -505
rect 72 -506 73 -505
rect 79 -506 80 -505
rect 142 -506 143 -505
rect 149 -506 150 -505
rect 394 -506 395 -505
rect 401 -506 402 -505
rect 418 -506 419 -505
rect 425 -506 426 -505
rect 996 -506 997 -505
rect 61 -508 62 -507
rect 639 -508 640 -507
rect 695 -508 696 -507
rect 926 -508 927 -507
rect 940 -508 941 -507
rect 1010 -508 1011 -507
rect 26 -510 27 -509
rect 940 -510 941 -509
rect 65 -512 66 -511
rect 303 -512 304 -511
rect 327 -512 328 -511
rect 422 -512 423 -511
rect 443 -512 444 -511
rect 478 -512 479 -511
rect 481 -512 482 -511
rect 779 -512 780 -511
rect 800 -512 801 -511
rect 863 -512 864 -511
rect 891 -512 892 -511
rect 982 -512 983 -511
rect 72 -514 73 -513
rect 583 -514 584 -513
rect 597 -514 598 -513
rect 842 -514 843 -513
rect 856 -514 857 -513
rect 891 -514 892 -513
rect 919 -514 920 -513
rect 996 -514 997 -513
rect 79 -516 80 -515
rect 93 -516 94 -515
rect 96 -516 97 -515
rect 240 -516 241 -515
rect 261 -516 262 -515
rect 317 -516 318 -515
rect 338 -516 339 -515
rect 460 -516 461 -515
rect 464 -516 465 -515
rect 471 -516 472 -515
rect 474 -516 475 -515
rect 590 -516 591 -515
rect 597 -516 598 -515
rect 828 -516 829 -515
rect 877 -516 878 -515
rect 919 -516 920 -515
rect 51 -518 52 -517
rect 471 -518 472 -517
rect 485 -518 486 -517
rect 492 -518 493 -517
rect 502 -518 503 -517
rect 730 -518 731 -517
rect 758 -518 759 -517
rect 807 -518 808 -517
rect 51 -520 52 -519
rect 331 -520 332 -519
rect 341 -520 342 -519
rect 632 -520 633 -519
rect 712 -520 713 -519
rect 828 -520 829 -519
rect 100 -522 101 -521
rect 359 -522 360 -521
rect 383 -522 384 -521
rect 856 -522 857 -521
rect 2 -524 3 -523
rect 100 -524 101 -523
rect 114 -524 115 -523
rect 380 -524 381 -523
rect 436 -524 437 -523
rect 485 -524 486 -523
rect 506 -524 507 -523
rect 590 -524 591 -523
rect 600 -524 601 -523
rect 954 -524 955 -523
rect 114 -526 115 -525
rect 208 -526 209 -525
rect 261 -526 262 -525
rect 268 -526 269 -525
rect 271 -526 272 -525
rect 779 -526 780 -525
rect 121 -528 122 -527
rect 562 -528 563 -527
rect 569 -528 570 -527
rect 604 -528 605 -527
rect 716 -528 717 -527
rect 800 -528 801 -527
rect 128 -530 129 -529
rect 387 -530 388 -529
rect 457 -530 458 -529
rect 884 -530 885 -529
rect 107 -532 108 -531
rect 387 -532 388 -531
rect 429 -532 430 -531
rect 457 -532 458 -531
rect 506 -532 507 -531
rect 660 -532 661 -531
rect 758 -532 759 -531
rect 849 -532 850 -531
rect 107 -534 108 -533
rect 821 -534 822 -533
rect 128 -536 129 -535
rect 205 -536 206 -535
rect 303 -536 304 -535
rect 436 -536 437 -535
rect 523 -536 524 -535
rect 898 -536 899 -535
rect 135 -538 136 -537
rect 429 -538 430 -537
rect 534 -538 535 -537
rect 709 -538 710 -537
rect 723 -538 724 -537
rect 898 -538 899 -537
rect 135 -540 136 -539
rect 254 -540 255 -539
rect 324 -540 325 -539
rect 884 -540 885 -539
rect 142 -542 143 -541
rect 275 -542 276 -541
rect 324 -542 325 -541
rect 450 -542 451 -541
rect 534 -542 535 -541
rect 695 -542 696 -541
rect 723 -542 724 -541
rect 786 -542 787 -541
rect 145 -544 146 -543
rect 240 -544 241 -543
rect 247 -544 248 -543
rect 254 -544 255 -543
rect 275 -544 276 -543
rect 289 -544 290 -543
rect 331 -544 332 -543
rect 684 -544 685 -543
rect 688 -544 689 -543
rect 786 -544 787 -543
rect 138 -546 139 -545
rect 289 -546 290 -545
rect 345 -546 346 -545
rect 681 -546 682 -545
rect 744 -546 745 -545
rect 821 -546 822 -545
rect 149 -548 150 -547
rect 233 -548 234 -547
rect 247 -548 248 -547
rect 268 -548 269 -547
rect 348 -548 349 -547
rect 674 -548 675 -547
rect 681 -548 682 -547
rect 933 -548 934 -547
rect 86 -550 87 -549
rect 233 -550 234 -549
rect 348 -550 349 -549
rect 443 -550 444 -549
rect 450 -550 451 -549
rect 464 -550 465 -549
rect 527 -550 528 -549
rect 674 -550 675 -549
rect 702 -550 703 -549
rect 744 -550 745 -549
rect 751 -550 752 -549
rect 849 -550 850 -549
rect 86 -552 87 -551
rect 170 -552 171 -551
rect 180 -552 181 -551
rect 226 -552 227 -551
rect 366 -552 367 -551
rect 660 -552 661 -551
rect 93 -554 94 -553
rect 933 -554 934 -553
rect 156 -556 157 -555
rect 352 -556 353 -555
rect 527 -556 528 -555
rect 583 -556 584 -555
rect 611 -556 612 -555
rect 702 -556 703 -555
rect 156 -558 157 -557
rect 215 -558 216 -557
rect 537 -558 538 -557
rect 877 -558 878 -557
rect 163 -560 164 -559
rect 170 -560 171 -559
rect 191 -560 192 -559
rect 226 -560 227 -559
rect 537 -560 538 -559
rect 667 -560 668 -559
rect 163 -562 164 -561
rect 366 -562 367 -561
rect 541 -562 542 -561
rect 751 -562 752 -561
rect 166 -564 167 -563
rect 1024 -564 1025 -563
rect 184 -566 185 -565
rect 191 -566 192 -565
rect 198 -566 199 -565
rect 1080 -566 1081 -565
rect 184 -568 185 -567
rect 219 -568 220 -567
rect 513 -568 514 -567
rect 541 -568 542 -567
rect 555 -568 556 -567
rect 565 -568 566 -567
rect 572 -568 573 -567
rect 793 -568 794 -567
rect 198 -570 199 -569
rect 208 -570 209 -569
rect 219 -570 220 -569
rect 611 -570 612 -569
rect 625 -570 626 -569
rect 716 -570 717 -569
rect 737 -570 738 -569
rect 793 -570 794 -569
rect 408 -572 409 -571
rect 737 -572 738 -571
rect 408 -574 409 -573
rect 576 -574 577 -573
rect 579 -574 580 -573
rect 912 -574 913 -573
rect 513 -576 514 -575
rect 520 -576 521 -575
rect 562 -576 563 -575
rect 1087 -576 1088 -575
rect 625 -578 626 -577
rect 653 -578 654 -577
rect 548 -580 549 -579
rect 653 -580 654 -579
rect 548 -582 549 -581
rect 1003 -582 1004 -581
rect 635 -584 636 -583
rect 667 -584 668 -583
rect 989 -584 990 -583
rect 1003 -584 1004 -583
rect 642 -586 643 -585
rect 688 -586 689 -585
rect 961 -586 962 -585
rect 989 -586 990 -585
rect 905 -588 906 -587
rect 961 -588 962 -587
rect 905 -590 906 -589
rect 947 -590 948 -589
rect 870 -592 871 -591
rect 947 -592 948 -591
rect 572 -594 573 -593
rect 870 -594 871 -593
rect 2 -605 3 -604
rect 233 -605 234 -604
rect 254 -605 255 -604
rect 268 -605 269 -604
rect 289 -605 290 -604
rect 534 -605 535 -604
rect 544 -605 545 -604
rect 1010 -605 1011 -604
rect 1111 -605 1112 -604
rect 1143 -605 1144 -604
rect 2 -607 3 -606
rect 107 -607 108 -606
rect 121 -607 122 -606
rect 268 -607 269 -606
rect 310 -607 311 -606
rect 523 -607 524 -606
rect 534 -607 535 -606
rect 646 -607 647 -606
rect 684 -607 685 -606
rect 1052 -607 1053 -606
rect 1115 -607 1116 -606
rect 1150 -607 1151 -606
rect 5 -609 6 -608
rect 527 -609 528 -608
rect 548 -609 549 -608
rect 898 -609 899 -608
rect 989 -609 990 -608
rect 1052 -609 1053 -608
rect 1101 -609 1102 -608
rect 1115 -609 1116 -608
rect 1129 -609 1130 -608
rect 1157 -609 1158 -608
rect 9 -611 10 -610
rect 212 -611 213 -610
rect 338 -611 339 -610
rect 751 -611 752 -610
rect 898 -611 899 -610
rect 1045 -611 1046 -610
rect 1094 -611 1095 -610
rect 1101 -611 1102 -610
rect 1129 -611 1130 -610
rect 1139 -611 1140 -610
rect 16 -613 17 -612
rect 348 -613 349 -612
rect 362 -613 363 -612
rect 576 -613 577 -612
rect 579 -613 580 -612
rect 1038 -613 1039 -612
rect 1066 -613 1067 -612
rect 1094 -613 1095 -612
rect 16 -615 17 -614
rect 65 -615 66 -614
rect 72 -615 73 -614
rect 516 -615 517 -614
rect 541 -615 542 -614
rect 576 -615 577 -614
rect 604 -615 605 -614
rect 1108 -615 1109 -614
rect 23 -617 24 -616
rect 128 -617 129 -616
rect 135 -617 136 -616
rect 212 -617 213 -616
rect 338 -617 339 -616
rect 457 -617 458 -616
rect 460 -617 461 -616
rect 842 -617 843 -616
rect 926 -617 927 -616
rect 1066 -617 1067 -616
rect 26 -619 27 -618
rect 58 -619 59 -618
rect 65 -619 66 -618
rect 296 -619 297 -618
rect 341 -619 342 -618
rect 611 -619 612 -618
rect 709 -619 710 -618
rect 786 -619 787 -618
rect 926 -619 927 -618
rect 933 -619 934 -618
rect 961 -619 962 -618
rect 989 -619 990 -618
rect 1024 -619 1025 -618
rect 1045 -619 1046 -618
rect 37 -621 38 -620
rect 618 -621 619 -620
rect 712 -621 713 -620
rect 1087 -621 1088 -620
rect 47 -623 48 -622
rect 345 -623 346 -622
rect 366 -623 367 -622
rect 565 -623 566 -622
rect 569 -623 570 -622
rect 737 -623 738 -622
rect 786 -623 787 -622
rect 975 -623 976 -622
rect 1031 -623 1032 -622
rect 1087 -623 1088 -622
rect 51 -625 52 -624
rect 233 -625 234 -624
rect 292 -625 293 -624
rect 611 -625 612 -624
rect 618 -625 619 -624
rect 744 -625 745 -624
rect 905 -625 906 -624
rect 975 -625 976 -624
rect 982 -625 983 -624
rect 1031 -625 1032 -624
rect 44 -627 45 -626
rect 51 -627 52 -626
rect 58 -627 59 -626
rect 170 -627 171 -626
rect 173 -627 174 -626
rect 660 -627 661 -626
rect 730 -627 731 -626
rect 807 -627 808 -626
rect 870 -627 871 -626
rect 905 -627 906 -626
rect 912 -627 913 -626
rect 961 -627 962 -626
rect 968 -627 969 -626
rect 982 -627 983 -626
rect 40 -629 41 -628
rect 660 -629 661 -628
rect 726 -629 727 -628
rect 968 -629 969 -628
rect 44 -631 45 -630
rect 765 -631 766 -630
rect 933 -631 934 -630
rect 940 -631 941 -630
rect 72 -633 73 -632
rect 79 -633 80 -632
rect 86 -633 87 -632
rect 215 -633 216 -632
rect 296 -633 297 -632
rect 597 -633 598 -632
rect 604 -633 605 -632
rect 835 -633 836 -632
rect 940 -633 941 -632
rect 947 -633 948 -632
rect 86 -635 87 -634
rect 142 -635 143 -634
rect 156 -635 157 -634
rect 254 -635 255 -634
rect 317 -635 318 -634
rect 345 -635 346 -634
rect 359 -635 360 -634
rect 366 -635 367 -634
rect 380 -635 381 -634
rect 383 -635 384 -634
rect 394 -635 395 -634
rect 541 -635 542 -634
rect 548 -635 549 -634
rect 555 -635 556 -634
rect 562 -635 563 -634
rect 1017 -635 1018 -634
rect 37 -637 38 -636
rect 359 -637 360 -636
rect 380 -637 381 -636
rect 387 -637 388 -636
rect 394 -637 395 -636
rect 450 -637 451 -636
rect 453 -637 454 -636
rect 485 -637 486 -636
rect 513 -637 514 -636
rect 569 -637 570 -636
rect 572 -637 573 -636
rect 863 -637 864 -636
rect 947 -637 948 -636
rect 954 -637 955 -636
rect 1003 -637 1004 -636
rect 1017 -637 1018 -636
rect 93 -639 94 -638
rect 1073 -639 1074 -638
rect 93 -641 94 -640
rect 219 -641 220 -640
rect 313 -641 314 -640
rect 317 -641 318 -640
rect 387 -641 388 -640
rect 590 -641 591 -640
rect 597 -641 598 -640
rect 688 -641 689 -640
rect 765 -641 766 -640
rect 772 -641 773 -640
rect 828 -641 829 -640
rect 835 -641 836 -640
rect 863 -641 864 -640
rect 919 -641 920 -640
rect 1059 -641 1060 -640
rect 1073 -641 1074 -640
rect 100 -643 101 -642
rect 996 -643 997 -642
rect 100 -645 101 -644
rect 131 -645 132 -644
rect 135 -645 136 -644
rect 222 -645 223 -644
rect 383 -645 384 -644
rect 590 -645 591 -644
rect 625 -645 626 -644
rect 919 -645 920 -644
rect 107 -647 108 -646
rect 184 -647 185 -646
rect 201 -647 202 -646
rect 639 -647 640 -646
rect 688 -647 689 -646
rect 733 -647 734 -646
rect 789 -647 790 -646
rect 996 -647 997 -646
rect 114 -649 115 -648
rect 807 -649 808 -648
rect 117 -651 118 -650
rect 156 -651 157 -650
rect 163 -651 164 -650
rect 282 -651 283 -650
rect 401 -651 402 -650
rect 485 -651 486 -650
rect 495 -651 496 -650
rect 639 -651 640 -650
rect 723 -651 724 -650
rect 828 -651 829 -650
rect 128 -653 129 -652
rect 1038 -653 1039 -652
rect 138 -655 139 -654
rect 800 -655 801 -654
rect 142 -657 143 -656
rect 149 -657 150 -656
rect 163 -657 164 -656
rect 261 -657 262 -656
rect 275 -657 276 -656
rect 282 -657 283 -656
rect 408 -657 409 -656
rect 555 -657 556 -656
rect 562 -657 563 -656
rect 842 -657 843 -656
rect 30 -659 31 -658
rect 149 -659 150 -658
rect 177 -659 178 -658
rect 1003 -659 1004 -658
rect 30 -661 31 -660
rect 82 -661 83 -660
rect 124 -661 125 -660
rect 261 -661 262 -660
rect 275 -661 276 -660
rect 457 -661 458 -660
rect 467 -661 468 -660
rect 653 -661 654 -660
rect 723 -661 724 -660
rect 912 -661 913 -660
rect 177 -663 178 -662
rect 191 -663 192 -662
rect 205 -663 206 -662
rect 352 -663 353 -662
rect 408 -663 409 -662
rect 478 -663 479 -662
rect 513 -663 514 -662
rect 646 -663 647 -662
rect 653 -663 654 -662
rect 702 -663 703 -662
rect 800 -663 801 -662
rect 814 -663 815 -662
rect 184 -665 185 -664
rect 198 -665 199 -664
rect 205 -665 206 -664
rect 324 -665 325 -664
rect 352 -665 353 -664
rect 492 -665 493 -664
rect 520 -665 521 -664
rect 870 -665 871 -664
rect 219 -667 220 -666
rect 247 -667 248 -666
rect 415 -667 416 -666
rect 436 -667 437 -666
rect 439 -667 440 -666
rect 1010 -667 1011 -666
rect 191 -669 192 -668
rect 247 -669 248 -668
rect 415 -669 416 -668
rect 478 -669 479 -668
rect 492 -669 493 -668
rect 674 -669 675 -668
rect 702 -669 703 -668
rect 856 -669 857 -668
rect 226 -671 227 -670
rect 401 -671 402 -670
rect 429 -671 430 -670
rect 625 -671 626 -670
rect 632 -671 633 -670
rect 954 -671 955 -670
rect 422 -673 423 -672
rect 429 -673 430 -672
rect 443 -673 444 -672
rect 520 -673 521 -672
rect 551 -673 552 -672
rect 737 -673 738 -672
rect 775 -673 776 -672
rect 814 -673 815 -672
rect 856 -673 857 -672
rect 891 -673 892 -672
rect 324 -675 325 -674
rect 443 -675 444 -674
rect 450 -675 451 -674
rect 681 -675 682 -674
rect 884 -675 885 -674
rect 891 -675 892 -674
rect 422 -677 423 -676
rect 506 -677 507 -676
rect 583 -677 584 -676
rect 632 -677 633 -676
rect 674 -677 675 -676
rect 695 -677 696 -676
rect 877 -677 878 -676
rect 884 -677 885 -676
rect 103 -679 104 -678
rect 506 -679 507 -678
rect 583 -679 584 -678
rect 607 -679 608 -678
rect 667 -679 668 -678
rect 695 -679 696 -678
rect 849 -679 850 -678
rect 877 -679 878 -678
rect 467 -681 468 -680
rect 1024 -681 1025 -680
rect 471 -683 472 -682
rect 751 -683 752 -682
rect 849 -683 850 -682
rect 1080 -683 1081 -682
rect 471 -685 472 -684
rect 499 -685 500 -684
rect 667 -685 668 -684
rect 758 -685 759 -684
rect 474 -687 475 -686
rect 1059 -687 1060 -686
rect 481 -689 482 -688
rect 499 -689 500 -688
rect 758 -689 759 -688
rect 821 -689 822 -688
rect 716 -691 717 -690
rect 821 -691 822 -690
rect 331 -693 332 -692
rect 716 -693 717 -692
rect 331 -695 332 -694
rect 1080 -695 1081 -694
rect 2 -706 3 -705
rect 114 -706 115 -705
rect 128 -706 129 -705
rect 156 -706 157 -705
rect 208 -706 209 -705
rect 292 -706 293 -705
rect 310 -706 311 -705
rect 485 -706 486 -705
rect 513 -706 514 -705
rect 891 -706 892 -705
rect 936 -706 937 -705
rect 968 -706 969 -705
rect 1080 -706 1081 -705
rect 1143 -706 1144 -705
rect 16 -708 17 -707
rect 369 -708 370 -707
rect 443 -708 444 -707
rect 772 -708 773 -707
rect 775 -708 776 -707
rect 1031 -708 1032 -707
rect 1083 -708 1084 -707
rect 1150 -708 1151 -707
rect 30 -710 31 -709
rect 198 -710 199 -709
rect 268 -710 269 -709
rect 271 -710 272 -709
rect 292 -710 293 -709
rect 401 -710 402 -709
rect 446 -710 447 -709
rect 821 -710 822 -709
rect 880 -710 881 -709
rect 884 -710 885 -709
rect 891 -710 892 -709
rect 1010 -710 1011 -709
rect 1031 -710 1032 -709
rect 1129 -710 1130 -709
rect 44 -712 45 -711
rect 51 -712 52 -711
rect 58 -712 59 -711
rect 289 -712 290 -711
rect 327 -712 328 -711
rect 422 -712 423 -711
rect 436 -712 437 -711
rect 446 -712 447 -711
rect 450 -712 451 -711
rect 590 -712 591 -711
rect 604 -712 605 -711
rect 800 -712 801 -711
rect 821 -712 822 -711
rect 870 -712 871 -711
rect 884 -712 885 -711
rect 947 -712 948 -711
rect 968 -712 969 -711
rect 1101 -712 1102 -711
rect 1111 -712 1112 -711
rect 1157 -712 1158 -711
rect 51 -714 52 -713
rect 156 -714 157 -713
rect 177 -714 178 -713
rect 198 -714 199 -713
rect 268 -714 269 -713
rect 275 -714 276 -713
rect 289 -714 290 -713
rect 471 -714 472 -713
rect 478 -714 479 -713
rect 919 -714 920 -713
rect 58 -716 59 -715
rect 296 -716 297 -715
rect 317 -716 318 -715
rect 422 -716 423 -715
rect 436 -716 437 -715
rect 443 -716 444 -715
rect 453 -716 454 -715
rect 569 -716 570 -715
rect 590 -716 591 -715
rect 940 -716 941 -715
rect 82 -718 83 -717
rect 89 -718 90 -717
rect 114 -718 115 -717
rect 135 -718 136 -717
rect 142 -718 143 -717
rect 159 -718 160 -717
rect 163 -718 164 -717
rect 177 -718 178 -717
rect 233 -718 234 -717
rect 296 -718 297 -717
rect 317 -718 318 -717
rect 394 -718 395 -717
rect 401 -718 402 -717
rect 499 -718 500 -717
rect 516 -718 517 -717
rect 716 -718 717 -717
rect 723 -718 724 -717
rect 954 -718 955 -717
rect 121 -720 122 -719
rect 478 -720 479 -719
rect 485 -720 486 -719
rect 583 -720 584 -719
rect 639 -720 640 -719
rect 663 -720 664 -719
rect 705 -720 706 -719
rect 912 -720 913 -719
rect 919 -720 920 -719
rect 1003 -720 1004 -719
rect 93 -722 94 -721
rect 121 -722 122 -721
rect 131 -722 132 -721
rect 345 -722 346 -721
rect 352 -722 353 -721
rect 460 -722 461 -721
rect 467 -722 468 -721
rect 807 -722 808 -721
rect 870 -722 871 -721
rect 898 -722 899 -721
rect 912 -722 913 -721
rect 996 -722 997 -721
rect 1003 -722 1004 -721
rect 1045 -722 1046 -721
rect 93 -724 94 -723
rect 331 -724 332 -723
rect 338 -724 339 -723
rect 492 -724 493 -723
rect 541 -724 542 -723
rect 646 -724 647 -723
rect 653 -724 654 -723
rect 667 -724 668 -723
rect 688 -724 689 -723
rect 807 -724 808 -723
rect 877 -724 878 -723
rect 898 -724 899 -723
rect 940 -724 941 -723
rect 989 -724 990 -723
rect 996 -724 997 -723
rect 1017 -724 1018 -723
rect 135 -726 136 -725
rect 152 -726 153 -725
rect 163 -726 164 -725
rect 184 -726 185 -725
rect 205 -726 206 -725
rect 331 -726 332 -725
rect 352 -726 353 -725
rect 380 -726 381 -725
rect 457 -726 458 -725
rect 618 -726 619 -725
rect 639 -726 640 -725
rect 674 -726 675 -725
rect 688 -726 689 -725
rect 709 -726 710 -725
rect 716 -726 717 -725
rect 1052 -726 1053 -725
rect 142 -728 143 -727
rect 149 -728 150 -727
rect 173 -728 174 -727
rect 460 -728 461 -727
rect 471 -728 472 -727
rect 506 -728 507 -727
rect 513 -728 514 -727
rect 618 -728 619 -727
rect 646 -728 647 -727
rect 681 -728 682 -727
rect 709 -728 710 -727
rect 730 -728 731 -727
rect 737 -728 738 -727
rect 744 -728 745 -727
rect 747 -728 748 -727
rect 800 -728 801 -727
rect 989 -728 990 -727
rect 1094 -728 1095 -727
rect 65 -730 66 -729
rect 149 -730 150 -729
rect 184 -730 185 -729
rect 387 -730 388 -729
rect 457 -730 458 -729
rect 933 -730 934 -729
rect 37 -732 38 -731
rect 65 -732 66 -731
rect 226 -732 227 -731
rect 338 -732 339 -731
rect 359 -732 360 -731
rect 366 -732 367 -731
rect 380 -732 381 -731
rect 537 -732 538 -731
rect 544 -732 545 -731
rect 1038 -732 1039 -731
rect 30 -734 31 -733
rect 37 -734 38 -733
rect 226 -734 227 -733
rect 726 -734 727 -733
rect 730 -734 731 -733
rect 793 -734 794 -733
rect 863 -734 864 -733
rect 933 -734 934 -733
rect 233 -736 234 -735
rect 254 -736 255 -735
rect 261 -736 262 -735
rect 499 -736 500 -735
rect 506 -736 507 -735
rect 520 -736 521 -735
rect 555 -736 556 -735
rect 569 -736 570 -735
rect 583 -736 584 -735
rect 719 -736 720 -735
rect 723 -736 724 -735
rect 765 -736 766 -735
rect 775 -736 776 -735
rect 975 -736 976 -735
rect 79 -738 80 -737
rect 765 -738 766 -737
rect 786 -738 787 -737
rect 961 -738 962 -737
rect 79 -740 80 -739
rect 86 -740 87 -739
rect 240 -740 241 -739
rect 254 -740 255 -739
rect 261 -740 262 -739
rect 408 -740 409 -739
rect 464 -740 465 -739
rect 520 -740 521 -739
rect 534 -740 535 -739
rect 555 -740 556 -739
rect 562 -740 563 -739
rect 737 -740 738 -739
rect 751 -740 752 -739
rect 950 -740 951 -739
rect 954 -740 955 -739
rect 975 -740 976 -739
rect 23 -742 24 -741
rect 86 -742 87 -741
rect 240 -742 241 -741
rect 303 -742 304 -741
rect 310 -742 311 -741
rect 345 -742 346 -741
rect 362 -742 363 -741
rect 429 -742 430 -741
rect 495 -742 496 -741
rect 674 -742 675 -741
rect 681 -742 682 -741
rect 695 -742 696 -741
rect 702 -742 703 -741
rect 751 -742 752 -741
rect 758 -742 759 -741
rect 772 -742 773 -741
rect 786 -742 787 -741
rect 814 -742 815 -741
rect 856 -742 857 -741
rect 863 -742 864 -741
rect 23 -744 24 -743
rect 124 -744 125 -743
rect 219 -744 220 -743
rect 303 -744 304 -743
rect 324 -744 325 -743
rect 359 -744 360 -743
rect 387 -744 388 -743
rect 415 -744 416 -743
rect 534 -744 535 -743
rect 562 -744 563 -743
rect 597 -744 598 -743
rect 961 -744 962 -743
rect 100 -746 101 -745
rect 429 -746 430 -745
rect 597 -746 598 -745
rect 835 -746 836 -745
rect 856 -746 857 -745
rect 926 -746 927 -745
rect 100 -748 101 -747
rect 191 -748 192 -747
rect 208 -748 209 -747
rect 415 -748 416 -747
rect 653 -748 654 -747
rect 1066 -748 1067 -747
rect 107 -750 108 -749
rect 191 -750 192 -749
rect 212 -750 213 -749
rect 219 -750 220 -749
rect 271 -750 272 -749
rect 275 -750 276 -749
rect 324 -750 325 -749
rect 394 -750 395 -749
rect 408 -750 409 -749
rect 548 -750 549 -749
rect 656 -750 657 -749
rect 695 -750 696 -749
rect 702 -750 703 -749
rect 1073 -750 1074 -749
rect 107 -752 108 -751
rect 247 -752 248 -751
rect 548 -752 549 -751
rect 660 -752 661 -751
rect 758 -752 759 -751
rect 1059 -752 1060 -751
rect 103 -754 104 -753
rect 247 -754 248 -753
rect 660 -754 661 -753
rect 828 -754 829 -753
rect 835 -754 836 -753
rect 982 -754 983 -753
rect 170 -756 171 -755
rect 212 -756 213 -755
rect 814 -756 815 -755
rect 905 -756 906 -755
rect 926 -756 927 -755
rect 1115 -756 1116 -755
rect 9 -758 10 -757
rect 170 -758 171 -757
rect 828 -758 829 -757
rect 842 -758 843 -757
rect 849 -758 850 -757
rect 905 -758 906 -757
rect 982 -758 983 -757
rect 1087 -758 1088 -757
rect 527 -760 528 -759
rect 842 -760 843 -759
rect 849 -760 850 -759
rect 1024 -760 1025 -759
rect 527 -762 528 -761
rect 576 -762 577 -761
rect 576 -764 577 -763
rect 611 -764 612 -763
rect 611 -766 612 -765
rect 625 -766 626 -765
rect 625 -768 626 -767
rect 632 -768 633 -767
rect 632 -770 633 -769
rect 779 -770 780 -769
rect 761 -772 762 -771
rect 779 -772 780 -771
rect 2 -783 3 -782
rect 156 -783 157 -782
rect 173 -783 174 -782
rect 467 -783 468 -782
rect 492 -783 493 -782
rect 1017 -783 1018 -782
rect 1087 -783 1088 -782
rect 1094 -783 1095 -782
rect 1108 -783 1109 -782
rect 1153 -783 1154 -782
rect 16 -785 17 -784
rect 184 -785 185 -784
rect 194 -785 195 -784
rect 394 -785 395 -784
rect 408 -785 409 -784
rect 492 -785 493 -784
rect 499 -785 500 -784
rect 663 -785 664 -784
rect 667 -785 668 -784
rect 716 -785 717 -784
rect 719 -785 720 -784
rect 744 -785 745 -784
rect 779 -785 780 -784
rect 1045 -785 1046 -784
rect 1122 -785 1123 -784
rect 1143 -785 1144 -784
rect 23 -787 24 -786
rect 138 -787 139 -786
rect 149 -787 150 -786
rect 268 -787 269 -786
rect 289 -787 290 -786
rect 345 -787 346 -786
rect 355 -787 356 -786
rect 954 -787 955 -786
rect 957 -787 958 -786
rect 996 -787 997 -786
rect 1010 -787 1011 -786
rect 1066 -787 1067 -786
rect 1139 -787 1140 -786
rect 1150 -787 1151 -786
rect 23 -789 24 -788
rect 86 -789 87 -788
rect 107 -789 108 -788
rect 327 -789 328 -788
rect 341 -789 342 -788
rect 352 -789 353 -788
rect 408 -789 409 -788
rect 481 -789 482 -788
rect 506 -789 507 -788
rect 534 -789 535 -788
rect 537 -789 538 -788
rect 632 -789 633 -788
rect 646 -789 647 -788
rect 1101 -789 1102 -788
rect 30 -791 31 -790
rect 502 -791 503 -790
rect 548 -791 549 -790
rect 667 -791 668 -790
rect 674 -791 675 -790
rect 933 -791 934 -790
rect 947 -791 948 -790
rect 1003 -791 1004 -790
rect 40 -793 41 -792
rect 618 -793 619 -792
rect 621 -793 622 -792
rect 870 -793 871 -792
rect 884 -793 885 -792
rect 1003 -793 1004 -792
rect 51 -795 52 -794
rect 170 -795 171 -794
rect 177 -795 178 -794
rect 184 -795 185 -794
rect 198 -795 199 -794
rect 205 -795 206 -794
rect 208 -795 209 -794
rect 240 -795 241 -794
rect 247 -795 248 -794
rect 506 -795 507 -794
rect 513 -795 514 -794
rect 548 -795 549 -794
rect 562 -795 563 -794
rect 618 -795 619 -794
rect 653 -795 654 -794
rect 842 -795 843 -794
rect 866 -795 867 -794
rect 1052 -795 1053 -794
rect 51 -797 52 -796
rect 460 -797 461 -796
rect 464 -797 465 -796
rect 758 -797 759 -796
rect 768 -797 769 -796
rect 1010 -797 1011 -796
rect 58 -799 59 -798
rect 530 -799 531 -798
rect 541 -799 542 -798
rect 842 -799 843 -798
rect 912 -799 913 -798
rect 996 -799 997 -798
rect 58 -801 59 -800
rect 261 -801 262 -800
rect 268 -801 269 -800
rect 450 -801 451 -800
rect 453 -801 454 -800
rect 905 -801 906 -800
rect 961 -801 962 -800
rect 1073 -801 1074 -800
rect 65 -803 66 -802
rect 100 -803 101 -802
rect 128 -803 129 -802
rect 513 -803 514 -802
rect 593 -803 594 -802
rect 1059 -803 1060 -802
rect 65 -805 66 -804
rect 72 -805 73 -804
rect 75 -805 76 -804
rect 107 -805 108 -804
rect 128 -805 129 -804
rect 226 -805 227 -804
rect 240 -805 241 -804
rect 499 -805 500 -804
rect 604 -805 605 -804
rect 632 -805 633 -804
rect 653 -805 654 -804
rect 1122 -805 1123 -804
rect 86 -807 87 -806
rect 114 -807 115 -806
rect 156 -807 157 -806
rect 324 -807 325 -806
rect 345 -807 346 -806
rect 415 -807 416 -806
rect 422 -807 423 -806
rect 450 -807 451 -806
rect 457 -807 458 -806
rect 926 -807 927 -806
rect 982 -807 983 -806
rect 1024 -807 1025 -806
rect 114 -809 115 -808
rect 296 -809 297 -808
rect 310 -809 311 -808
rect 338 -809 339 -808
rect 359 -809 360 -808
rect 464 -809 465 -808
rect 478 -809 479 -808
rect 674 -809 675 -808
rect 737 -809 738 -808
rect 1038 -809 1039 -808
rect 93 -811 94 -810
rect 296 -811 297 -810
rect 313 -811 314 -810
rect 520 -811 521 -810
rect 527 -811 528 -810
rect 982 -811 983 -810
rect 989 -811 990 -810
rect 1115 -811 1116 -810
rect 93 -813 94 -812
rect 331 -813 332 -812
rect 380 -813 381 -812
rect 527 -813 528 -812
rect 607 -813 608 -812
rect 870 -813 871 -812
rect 877 -813 878 -812
rect 989 -813 990 -812
rect 152 -815 153 -814
rect 359 -815 360 -814
rect 383 -815 384 -814
rect 534 -815 535 -814
rect 614 -815 615 -814
rect 849 -815 850 -814
rect 898 -815 899 -814
rect 905 -815 906 -814
rect 926 -815 927 -814
rect 1031 -815 1032 -814
rect 177 -817 178 -816
rect 292 -817 293 -816
rect 317 -817 318 -816
rect 415 -817 416 -816
rect 422 -817 423 -816
rect 436 -817 437 -816
rect 443 -817 444 -816
rect 590 -817 591 -816
rect 656 -817 657 -816
rect 705 -817 706 -816
rect 744 -817 745 -816
rect 936 -817 937 -816
rect 142 -819 143 -818
rect 443 -819 444 -818
rect 457 -819 458 -818
rect 485 -819 486 -818
rect 495 -819 496 -818
rect 646 -819 647 -818
rect 656 -819 657 -818
rect 947 -819 948 -818
rect 142 -821 143 -820
rect 233 -821 234 -820
rect 254 -821 255 -820
rect 331 -821 332 -820
rect 387 -821 388 -820
rect 541 -821 542 -820
rect 660 -821 661 -820
rect 1080 -821 1081 -820
rect 121 -823 122 -822
rect 254 -823 255 -822
rect 317 -823 318 -822
rect 366 -823 367 -822
rect 387 -823 388 -822
rect 429 -823 430 -822
rect 436 -823 437 -822
rect 702 -823 703 -822
rect 751 -823 752 -822
rect 849 -823 850 -822
rect 863 -823 864 -822
rect 1031 -823 1032 -822
rect 79 -825 80 -824
rect 121 -825 122 -824
rect 198 -825 199 -824
rect 212 -825 213 -824
rect 222 -825 223 -824
rect 247 -825 248 -824
rect 261 -825 262 -824
rect 366 -825 367 -824
rect 401 -825 402 -824
rect 702 -825 703 -824
rect 751 -825 752 -824
rect 940 -825 941 -824
rect 212 -827 213 -826
rect 226 -827 227 -826
rect 233 -827 234 -826
rect 446 -827 447 -826
rect 471 -827 472 -826
rect 485 -827 486 -826
rect 520 -827 521 -826
rect 775 -827 776 -826
rect 779 -827 780 -826
rect 821 -827 822 -826
rect 828 -827 829 -826
rect 877 -827 878 -826
rect 324 -829 325 -828
rect 737 -829 738 -828
rect 765 -829 766 -828
rect 961 -829 962 -828
rect 401 -831 402 -830
rect 635 -831 636 -830
rect 660 -831 661 -830
rect 681 -831 682 -830
rect 723 -831 724 -830
rect 821 -831 822 -830
rect 828 -831 829 -830
rect 975 -831 976 -830
rect 135 -833 136 -832
rect 681 -833 682 -832
rect 772 -833 773 -832
rect 912 -833 913 -832
rect 135 -835 136 -834
rect 163 -835 164 -834
rect 471 -835 472 -834
rect 611 -835 612 -834
rect 688 -835 689 -834
rect 772 -835 773 -834
rect 793 -835 794 -834
rect 919 -835 920 -834
rect 163 -837 164 -836
rect 219 -837 220 -836
rect 478 -837 479 -836
rect 597 -837 598 -836
rect 604 -837 605 -836
rect 975 -837 976 -836
rect 219 -839 220 -838
rect 303 -839 304 -838
rect 555 -839 556 -838
rect 723 -839 724 -838
rect 730 -839 731 -838
rect 793 -839 794 -838
rect 807 -839 808 -838
rect 919 -839 920 -838
rect 282 -841 283 -840
rect 303 -841 304 -840
rect 555 -841 556 -840
rect 800 -841 801 -840
rect 814 -841 815 -840
rect 898 -841 899 -840
rect 191 -843 192 -842
rect 282 -843 283 -842
rect 565 -843 566 -842
rect 765 -843 766 -842
rect 786 -843 787 -842
rect 814 -843 815 -842
rect 835 -843 836 -842
rect 884 -843 885 -842
rect 103 -845 104 -844
rect 835 -845 836 -844
rect 863 -845 864 -844
rect 968 -845 969 -844
rect 82 -847 83 -846
rect 968 -847 969 -846
rect 576 -849 577 -848
rect 597 -849 598 -848
rect 611 -849 612 -848
rect 940 -849 941 -848
rect 352 -851 353 -850
rect 576 -851 577 -850
rect 579 -851 580 -850
rect 807 -851 808 -850
rect 639 -853 640 -852
rect 688 -853 689 -852
rect 695 -853 696 -852
rect 730 -853 731 -852
rect 786 -853 787 -852
rect 856 -853 857 -852
rect 338 -855 339 -854
rect 695 -855 696 -854
rect 709 -855 710 -854
rect 800 -855 801 -854
rect 856 -855 857 -854
rect 891 -855 892 -854
rect 369 -857 370 -856
rect 891 -857 892 -856
rect 394 -859 395 -858
rect 639 -859 640 -858
rect 709 -859 710 -858
rect 796 -859 797 -858
rect 9 -870 10 -869
rect 149 -870 150 -869
rect 198 -870 199 -869
rect 219 -870 220 -869
rect 222 -870 223 -869
rect 282 -870 283 -869
rect 317 -870 318 -869
rect 432 -870 433 -869
rect 481 -870 482 -869
rect 870 -870 871 -869
rect 982 -870 983 -869
rect 1150 -870 1151 -869
rect 12 -872 13 -871
rect 380 -872 381 -871
rect 383 -872 384 -871
rect 544 -872 545 -871
rect 555 -872 556 -871
rect 1101 -872 1102 -871
rect 16 -874 17 -873
rect 152 -874 153 -873
rect 170 -874 171 -873
rect 380 -874 381 -873
rect 394 -874 395 -873
rect 912 -874 913 -873
rect 989 -874 990 -873
rect 1101 -874 1102 -873
rect 30 -876 31 -875
rect 429 -876 430 -875
rect 492 -876 493 -875
rect 579 -876 580 -875
rect 583 -876 584 -875
rect 653 -876 654 -875
rect 768 -876 769 -875
rect 1031 -876 1032 -875
rect 1052 -876 1053 -875
rect 1157 -876 1158 -875
rect 30 -878 31 -877
rect 75 -878 76 -877
rect 79 -878 80 -877
rect 765 -878 766 -877
rect 779 -878 780 -877
rect 870 -878 871 -877
rect 912 -878 913 -877
rect 933 -878 934 -877
rect 1017 -878 1018 -877
rect 1129 -878 1130 -877
rect 58 -880 59 -879
rect 446 -880 447 -879
rect 478 -880 479 -879
rect 492 -880 493 -879
rect 537 -880 538 -879
rect 919 -880 920 -879
rect 933 -880 934 -879
rect 947 -880 948 -879
rect 1087 -880 1088 -879
rect 1094 -880 1095 -879
rect 1097 -880 1098 -879
rect 1143 -880 1144 -879
rect 16 -882 17 -881
rect 58 -882 59 -881
rect 65 -882 66 -881
rect 82 -882 83 -881
rect 93 -882 94 -881
rect 502 -882 503 -881
rect 565 -882 566 -881
rect 702 -882 703 -881
rect 709 -882 710 -881
rect 1052 -882 1053 -881
rect 1115 -882 1116 -881
rect 1129 -882 1130 -881
rect 72 -884 73 -883
rect 1136 -884 1137 -883
rect 75 -886 76 -885
rect 86 -886 87 -885
rect 93 -886 94 -885
rect 156 -886 157 -885
rect 170 -886 171 -885
rect 453 -886 454 -885
rect 572 -886 573 -885
rect 821 -886 822 -885
rect 856 -886 857 -885
rect 982 -886 983 -885
rect 1108 -886 1109 -885
rect 1115 -886 1116 -885
rect 79 -888 80 -887
rect 548 -888 549 -887
rect 576 -888 577 -887
rect 1087 -888 1088 -887
rect 1108 -888 1109 -887
rect 1122 -888 1123 -887
rect 86 -890 87 -889
rect 128 -890 129 -889
rect 135 -890 136 -889
rect 191 -890 192 -889
rect 198 -890 199 -889
rect 205 -890 206 -889
rect 229 -890 230 -889
rect 555 -890 556 -889
rect 562 -890 563 -889
rect 1122 -890 1123 -889
rect 51 -892 52 -891
rect 128 -892 129 -891
rect 135 -892 136 -891
rect 268 -892 269 -891
rect 310 -892 311 -891
rect 317 -892 318 -891
rect 324 -892 325 -891
rect 499 -892 500 -891
rect 548 -892 549 -891
rect 698 -892 699 -891
rect 730 -892 731 -891
rect 821 -892 822 -891
rect 905 -892 906 -891
rect 1143 -892 1144 -891
rect 51 -894 52 -893
rect 415 -894 416 -893
rect 418 -894 419 -893
rect 1038 -894 1039 -893
rect 82 -896 83 -895
rect 191 -896 192 -895
rect 261 -896 262 -895
rect 579 -896 580 -895
rect 590 -896 591 -895
rect 1073 -896 1074 -895
rect 114 -898 115 -897
rect 355 -898 356 -897
rect 359 -898 360 -897
rect 369 -898 370 -897
rect 394 -898 395 -897
rect 422 -898 423 -897
rect 439 -898 440 -897
rect 1031 -898 1032 -897
rect 1073 -898 1074 -897
rect 1080 -898 1081 -897
rect 114 -900 115 -899
rect 240 -900 241 -899
rect 268 -900 269 -899
rect 299 -900 300 -899
rect 310 -900 311 -899
rect 614 -900 615 -899
rect 635 -900 636 -899
rect 1003 -900 1004 -899
rect 1010 -900 1011 -899
rect 1038 -900 1039 -899
rect 142 -902 143 -901
rect 226 -902 227 -901
rect 240 -902 241 -901
rect 345 -902 346 -901
rect 359 -902 360 -901
rect 751 -902 752 -901
rect 758 -902 759 -901
rect 779 -902 780 -901
rect 891 -902 892 -901
rect 905 -902 906 -901
rect 919 -902 920 -901
rect 926 -902 927 -901
rect 947 -902 948 -901
rect 1024 -902 1025 -901
rect 142 -904 143 -903
rect 212 -904 213 -903
rect 226 -904 227 -903
rect 450 -904 451 -903
rect 562 -904 563 -903
rect 597 -904 598 -903
rect 604 -904 605 -903
rect 1017 -904 1018 -903
rect 149 -906 150 -905
rect 583 -906 584 -905
rect 604 -906 605 -905
rect 618 -906 619 -905
rect 639 -906 640 -905
rect 863 -906 864 -905
rect 898 -906 899 -905
rect 926 -906 927 -905
rect 961 -906 962 -905
rect 1010 -906 1011 -905
rect 156 -908 157 -907
rect 401 -908 402 -907
rect 408 -908 409 -907
rect 429 -908 430 -907
rect 443 -908 444 -907
rect 709 -908 710 -907
rect 723 -908 724 -907
rect 730 -908 731 -907
rect 751 -908 752 -907
rect 828 -908 829 -907
rect 961 -908 962 -907
rect 975 -908 976 -907
rect 996 -908 997 -907
rect 1003 -908 1004 -907
rect 163 -910 164 -909
rect 212 -910 213 -909
rect 254 -910 255 -909
rect 597 -910 598 -909
rect 611 -910 612 -909
rect 660 -910 661 -909
rect 674 -910 675 -909
rect 1080 -910 1081 -909
rect 121 -912 122 -911
rect 254 -912 255 -911
rect 324 -912 325 -911
rect 506 -912 507 -911
rect 534 -912 535 -911
rect 618 -912 619 -911
rect 625 -912 626 -911
rect 674 -912 675 -911
rect 695 -912 696 -911
rect 702 -912 703 -911
rect 716 -912 717 -911
rect 723 -912 724 -911
rect 793 -912 794 -911
rect 1024 -912 1025 -911
rect 2 -914 3 -913
rect 793 -914 794 -913
rect 807 -914 808 -913
rect 828 -914 829 -913
rect 884 -914 885 -913
rect 975 -914 976 -913
rect 100 -916 101 -915
rect 121 -916 122 -915
rect 163 -916 164 -915
rect 415 -916 416 -915
rect 443 -916 444 -915
rect 989 -916 990 -915
rect 65 -918 66 -917
rect 100 -918 101 -917
rect 177 -918 178 -917
rect 205 -918 206 -917
rect 331 -918 332 -917
rect 397 -918 398 -917
rect 408 -918 409 -917
rect 457 -918 458 -917
rect 481 -918 482 -917
rect 639 -918 640 -917
rect 646 -918 647 -917
rect 660 -918 661 -917
rect 716 -918 717 -917
rect 800 -918 801 -917
rect 807 -918 808 -917
rect 835 -918 836 -917
rect 877 -918 878 -917
rect 884 -918 885 -917
rect 289 -920 290 -919
rect 331 -920 332 -919
rect 338 -920 339 -919
rect 527 -920 528 -919
rect 541 -920 542 -919
rect 996 -920 997 -919
rect 107 -922 108 -921
rect 338 -922 339 -921
rect 341 -922 342 -921
rect 422 -922 423 -921
rect 450 -922 451 -921
rect 485 -922 486 -921
rect 506 -922 507 -921
rect 1059 -922 1060 -921
rect 107 -924 108 -923
rect 194 -924 195 -923
rect 289 -924 290 -923
rect 436 -924 437 -923
rect 457 -924 458 -923
rect 688 -924 689 -923
rect 814 -924 815 -923
rect 835 -924 836 -923
rect 849 -924 850 -923
rect 877 -924 878 -923
rect 1059 -924 1060 -923
rect 1066 -924 1067 -923
rect 72 -926 73 -925
rect 1066 -926 1067 -925
rect 345 -928 346 -927
rect 464 -928 465 -927
rect 471 -928 472 -927
rect 814 -928 815 -927
rect 352 -930 353 -929
rect 646 -930 647 -929
rect 688 -930 689 -929
rect 786 -930 787 -929
rect 362 -932 363 -931
rect 401 -932 402 -931
rect 464 -932 465 -931
rect 527 -932 528 -931
rect 541 -932 542 -931
rect 1045 -932 1046 -931
rect 366 -934 367 -933
rect 576 -934 577 -933
rect 593 -934 594 -933
rect 800 -934 801 -933
rect 352 -936 353 -935
rect 593 -936 594 -935
rect 614 -936 615 -935
rect 758 -936 759 -935
rect 366 -938 367 -937
rect 373 -938 374 -937
rect 485 -938 486 -937
rect 558 -938 559 -937
rect 569 -938 570 -937
rect 891 -938 892 -937
rect 177 -940 178 -939
rect 569 -940 570 -939
rect 621 -940 622 -939
rect 1045 -940 1046 -939
rect 369 -942 370 -941
rect 471 -942 472 -941
rect 513 -942 514 -941
rect 849 -942 850 -941
rect 373 -944 374 -943
rect 544 -944 545 -943
rect 625 -944 626 -943
rect 842 -944 843 -943
rect 513 -946 514 -945
rect 520 -946 521 -945
rect 632 -946 633 -945
rect 898 -946 899 -945
rect 23 -948 24 -947
rect 520 -948 521 -947
rect 632 -948 633 -947
rect 1136 -948 1137 -947
rect 23 -950 24 -949
rect 387 -950 388 -949
rect 681 -950 682 -949
rect 842 -950 843 -949
rect 247 -952 248 -951
rect 387 -952 388 -951
rect 667 -952 668 -951
rect 681 -952 682 -951
rect 744 -952 745 -951
rect 786 -952 787 -951
rect 233 -954 234 -953
rect 247 -954 248 -953
rect 667 -954 668 -953
rect 772 -954 773 -953
rect 233 -956 234 -955
rect 296 -956 297 -955
rect 691 -956 692 -955
rect 772 -956 773 -955
rect 737 -958 738 -957
rect 744 -958 745 -957
rect 37 -960 38 -959
rect 737 -960 738 -959
rect 9 -971 10 -970
rect 282 -971 283 -970
rect 285 -971 286 -970
rect 310 -971 311 -970
rect 359 -971 360 -970
rect 726 -971 727 -970
rect 859 -971 860 -970
rect 961 -971 962 -970
rect 9 -973 10 -972
rect 485 -973 486 -972
rect 541 -973 542 -972
rect 1136 -973 1137 -972
rect 16 -975 17 -974
rect 597 -975 598 -974
rect 607 -975 608 -974
rect 905 -975 906 -974
rect 16 -977 17 -976
rect 166 -977 167 -976
rect 194 -977 195 -976
rect 380 -977 381 -976
rect 401 -977 402 -976
rect 464 -977 465 -976
rect 467 -977 468 -976
rect 765 -977 766 -976
rect 23 -979 24 -978
rect 436 -979 437 -978
rect 439 -979 440 -978
rect 688 -979 689 -978
rect 691 -979 692 -978
rect 961 -979 962 -978
rect 23 -981 24 -980
rect 390 -981 391 -980
rect 436 -981 437 -980
rect 558 -981 559 -980
rect 569 -981 570 -980
rect 1115 -981 1116 -980
rect 30 -983 31 -982
rect 33 -983 34 -982
rect 37 -983 38 -982
rect 254 -983 255 -982
rect 271 -983 272 -982
rect 324 -983 325 -982
rect 362 -983 363 -982
rect 628 -983 629 -982
rect 632 -983 633 -982
rect 982 -983 983 -982
rect 30 -985 31 -984
rect 653 -985 654 -984
rect 695 -985 696 -984
rect 828 -985 829 -984
rect 982 -985 983 -984
rect 1045 -985 1046 -984
rect 33 -987 34 -986
rect 653 -987 654 -986
rect 698 -987 699 -986
rect 1052 -987 1053 -986
rect 37 -989 38 -988
rect 44 -989 45 -988
rect 65 -989 66 -988
rect 933 -989 934 -988
rect 1045 -989 1046 -988
rect 1073 -989 1074 -988
rect 44 -991 45 -990
rect 527 -991 528 -990
rect 569 -991 570 -990
rect 926 -991 927 -990
rect 933 -991 934 -990
rect 996 -991 997 -990
rect 1052 -991 1053 -990
rect 1101 -991 1102 -990
rect 2 -993 3 -992
rect 926 -993 927 -992
rect 68 -995 69 -994
rect 415 -995 416 -994
rect 422 -995 423 -994
rect 527 -995 528 -994
rect 576 -995 577 -994
rect 674 -995 675 -994
rect 786 -995 787 -994
rect 1073 -995 1074 -994
rect 68 -997 69 -996
rect 338 -997 339 -996
rect 380 -997 381 -996
rect 513 -997 514 -996
rect 579 -997 580 -996
rect 1024 -997 1025 -996
rect 72 -999 73 -998
rect 86 -999 87 -998
rect 114 -999 115 -998
rect 401 -999 402 -998
rect 415 -999 416 -998
rect 520 -999 521 -998
rect 590 -999 591 -998
rect 667 -999 668 -998
rect 674 -999 675 -998
rect 779 -999 780 -998
rect 786 -999 787 -998
rect 912 -999 913 -998
rect 1024 -999 1025 -998
rect 1122 -999 1123 -998
rect 72 -1001 73 -1000
rect 93 -1001 94 -1000
rect 114 -1001 115 -1000
rect 275 -1001 276 -1000
rect 282 -1001 283 -1000
rect 709 -1001 710 -1000
rect 779 -1001 780 -1000
rect 940 -1001 941 -1000
rect 82 -1003 83 -1002
rect 555 -1003 556 -1002
rect 590 -1003 591 -1002
rect 681 -1003 682 -1002
rect 709 -1003 710 -1002
rect 863 -1003 864 -1002
rect 912 -1003 913 -1002
rect 1031 -1003 1032 -1002
rect 82 -1005 83 -1004
rect 793 -1005 794 -1004
rect 842 -1005 843 -1004
rect 940 -1005 941 -1004
rect 1010 -1005 1011 -1004
rect 1031 -1005 1032 -1004
rect 86 -1007 87 -1006
rect 205 -1007 206 -1006
rect 229 -1007 230 -1006
rect 233 -1007 234 -1006
rect 240 -1007 241 -1006
rect 506 -1007 507 -1006
rect 513 -1007 514 -1006
rect 604 -1007 605 -1006
rect 614 -1007 615 -1006
rect 716 -1007 717 -1006
rect 793 -1007 794 -1006
rect 884 -1007 885 -1006
rect 1010 -1007 1011 -1006
rect 1041 -1007 1042 -1006
rect 93 -1009 94 -1008
rect 107 -1009 108 -1008
rect 135 -1009 136 -1008
rect 418 -1009 419 -1008
rect 443 -1009 444 -1008
rect 450 -1009 451 -1008
rect 471 -1009 472 -1008
rect 681 -1009 682 -1008
rect 716 -1009 717 -1008
rect 821 -1009 822 -1008
rect 842 -1009 843 -1008
rect 898 -1009 899 -1008
rect 58 -1011 59 -1010
rect 821 -1011 822 -1010
rect 863 -1011 864 -1010
rect 968 -1011 969 -1010
rect 58 -1013 59 -1012
rect 75 -1013 76 -1012
rect 107 -1013 108 -1012
rect 121 -1013 122 -1012
rect 135 -1013 136 -1012
rect 226 -1013 227 -1012
rect 233 -1013 234 -1012
rect 429 -1013 430 -1012
rect 450 -1013 451 -1012
rect 702 -1013 703 -1012
rect 884 -1013 885 -1012
rect 975 -1013 976 -1012
rect 121 -1015 122 -1014
rect 163 -1015 164 -1014
rect 191 -1015 192 -1014
rect 422 -1015 423 -1014
rect 471 -1015 472 -1014
rect 488 -1015 489 -1014
rect 492 -1015 493 -1014
rect 506 -1015 507 -1014
rect 520 -1015 521 -1014
rect 544 -1015 545 -1014
rect 548 -1015 549 -1014
rect 702 -1015 703 -1014
rect 898 -1015 899 -1014
rect 1017 -1015 1018 -1014
rect 149 -1017 150 -1016
rect 212 -1017 213 -1016
rect 240 -1017 241 -1016
rect 457 -1017 458 -1016
rect 474 -1017 475 -1016
rect 1017 -1017 1018 -1016
rect 163 -1019 164 -1018
rect 205 -1019 206 -1018
rect 254 -1019 255 -1018
rect 740 -1019 741 -1018
rect 947 -1019 948 -1018
rect 968 -1019 969 -1018
rect 975 -1019 976 -1018
rect 1038 -1019 1039 -1018
rect 191 -1021 192 -1020
rect 296 -1021 297 -1020
rect 303 -1021 304 -1020
rect 548 -1021 549 -1020
rect 555 -1021 556 -1020
rect 807 -1021 808 -1020
rect 856 -1021 857 -1020
rect 947 -1021 948 -1020
rect 177 -1023 178 -1022
rect 303 -1023 304 -1022
rect 306 -1023 307 -1022
rect 583 -1023 584 -1022
rect 593 -1023 594 -1022
rect 1080 -1023 1081 -1022
rect 177 -1025 178 -1024
rect 373 -1025 374 -1024
rect 408 -1025 409 -1024
rect 429 -1025 430 -1024
rect 446 -1025 447 -1024
rect 807 -1025 808 -1024
rect 1080 -1025 1081 -1024
rect 1094 -1025 1095 -1024
rect 268 -1027 269 -1026
rect 324 -1027 325 -1026
rect 331 -1027 332 -1026
rect 373 -1027 374 -1026
rect 408 -1027 409 -1026
rect 492 -1027 493 -1026
rect 502 -1027 503 -1026
rect 996 -1027 997 -1026
rect 142 -1029 143 -1028
rect 268 -1029 269 -1028
rect 275 -1029 276 -1028
rect 394 -1029 395 -1028
rect 457 -1029 458 -1028
rect 737 -1029 738 -1028
rect 51 -1031 52 -1030
rect 394 -1031 395 -1030
rect 478 -1031 479 -1030
rect 1087 -1031 1088 -1030
rect 2 -1033 3 -1032
rect 51 -1033 52 -1032
rect 100 -1033 101 -1032
rect 142 -1033 143 -1032
rect 156 -1033 157 -1032
rect 478 -1033 479 -1032
rect 481 -1033 482 -1032
rect 814 -1033 815 -1032
rect 156 -1035 157 -1034
rect 247 -1035 248 -1034
rect 289 -1035 290 -1034
rect 331 -1035 332 -1034
rect 338 -1035 339 -1034
rect 397 -1035 398 -1034
rect 583 -1035 584 -1034
rect 891 -1035 892 -1034
rect 247 -1037 248 -1036
rect 317 -1037 318 -1036
rect 600 -1037 601 -1036
rect 765 -1037 766 -1036
rect 891 -1037 892 -1036
rect 1003 -1037 1004 -1036
rect 289 -1039 290 -1038
rect 345 -1039 346 -1038
rect 618 -1039 619 -1038
rect 828 -1039 829 -1038
rect 1003 -1039 1004 -1038
rect 1066 -1039 1067 -1038
rect 261 -1041 262 -1040
rect 345 -1041 346 -1040
rect 562 -1041 563 -1040
rect 618 -1041 619 -1040
rect 621 -1041 622 -1040
rect 870 -1041 871 -1040
rect 919 -1041 920 -1040
rect 1066 -1041 1067 -1040
rect 261 -1043 262 -1042
rect 352 -1043 353 -1042
rect 499 -1043 500 -1042
rect 919 -1043 920 -1042
rect 310 -1045 311 -1044
rect 387 -1045 388 -1044
rect 562 -1045 563 -1044
rect 572 -1045 573 -1044
rect 635 -1045 636 -1044
rect 751 -1045 752 -1044
rect 870 -1045 871 -1044
rect 989 -1045 990 -1044
rect 317 -1047 318 -1046
rect 534 -1047 535 -1046
rect 572 -1047 573 -1046
rect 905 -1047 906 -1046
rect 989 -1047 990 -1046
rect 1108 -1047 1109 -1046
rect 352 -1049 353 -1048
rect 366 -1049 367 -1048
rect 387 -1049 388 -1048
rect 639 -1049 640 -1048
rect 667 -1049 668 -1048
rect 772 -1049 773 -1048
rect 128 -1051 129 -1050
rect 366 -1051 367 -1050
rect 495 -1051 496 -1050
rect 639 -1051 640 -1050
rect 737 -1051 738 -1050
rect 1129 -1051 1130 -1050
rect 128 -1053 129 -1052
rect 170 -1053 171 -1052
rect 534 -1053 535 -1052
rect 646 -1053 647 -1052
rect 751 -1053 752 -1052
rect 835 -1053 836 -1052
rect 1129 -1053 1130 -1052
rect 1157 -1053 1158 -1052
rect 170 -1055 171 -1054
rect 198 -1055 199 -1054
rect 611 -1055 612 -1054
rect 646 -1055 647 -1054
rect 800 -1055 801 -1054
rect 835 -1055 836 -1054
rect 198 -1057 199 -1056
rect 849 -1057 850 -1056
rect 611 -1059 612 -1058
rect 723 -1059 724 -1058
rect 744 -1059 745 -1058
rect 800 -1059 801 -1058
rect 849 -1059 850 -1058
rect 954 -1059 955 -1058
rect 625 -1061 626 -1060
rect 772 -1061 773 -1060
rect 954 -1061 955 -1060
rect 1059 -1061 1060 -1060
rect 502 -1063 503 -1062
rect 625 -1063 626 -1062
rect 635 -1063 636 -1062
rect 856 -1063 857 -1062
rect 723 -1065 724 -1064
rect 1143 -1065 1144 -1064
rect 730 -1067 731 -1066
rect 744 -1067 745 -1066
rect 1143 -1067 1144 -1066
rect 1150 -1067 1151 -1066
rect 660 -1069 661 -1068
rect 730 -1069 731 -1068
rect 660 -1071 661 -1070
rect 758 -1071 759 -1070
rect 758 -1073 759 -1072
rect 877 -1073 878 -1072
rect 604 -1075 605 -1074
rect 877 -1075 878 -1074
rect 5 -1086 6 -1085
rect 348 -1086 349 -1085
rect 366 -1086 367 -1085
rect 369 -1086 370 -1085
rect 390 -1086 391 -1085
rect 898 -1086 899 -1085
rect 947 -1086 948 -1085
rect 1038 -1086 1039 -1085
rect 1041 -1086 1042 -1085
rect 1066 -1086 1067 -1085
rect 1076 -1086 1077 -1085
rect 1080 -1086 1081 -1085
rect 1122 -1086 1123 -1085
rect 1129 -1086 1130 -1085
rect 1143 -1086 1144 -1085
rect 1150 -1086 1151 -1085
rect 9 -1088 10 -1087
rect 467 -1088 468 -1087
rect 488 -1088 489 -1087
rect 520 -1088 521 -1087
rect 523 -1088 524 -1087
rect 828 -1088 829 -1087
rect 905 -1088 906 -1087
rect 947 -1088 948 -1087
rect 996 -1088 997 -1087
rect 1059 -1088 1060 -1087
rect 9 -1090 10 -1089
rect 30 -1090 31 -1089
rect 40 -1090 41 -1089
rect 898 -1090 899 -1089
rect 982 -1090 983 -1089
rect 996 -1090 997 -1089
rect 1031 -1090 1032 -1089
rect 1066 -1090 1067 -1089
rect 16 -1092 17 -1091
rect 495 -1092 496 -1091
rect 513 -1092 514 -1091
rect 691 -1092 692 -1091
rect 723 -1092 724 -1091
rect 751 -1092 752 -1091
rect 779 -1092 780 -1091
rect 828 -1092 829 -1091
rect 856 -1092 857 -1091
rect 905 -1092 906 -1091
rect 926 -1092 927 -1091
rect 982 -1092 983 -1091
rect 1017 -1092 1018 -1091
rect 1031 -1092 1032 -1091
rect 51 -1094 52 -1093
rect 58 -1094 59 -1093
rect 61 -1094 62 -1093
rect 198 -1094 199 -1093
rect 212 -1094 213 -1093
rect 800 -1094 801 -1093
rect 817 -1094 818 -1093
rect 954 -1094 955 -1093
rect 1010 -1094 1011 -1093
rect 1017 -1094 1018 -1093
rect 51 -1096 52 -1095
rect 275 -1096 276 -1095
rect 324 -1096 325 -1095
rect 408 -1096 409 -1095
rect 418 -1096 419 -1095
rect 989 -1096 990 -1095
rect 1003 -1096 1004 -1095
rect 1010 -1096 1011 -1095
rect 65 -1098 66 -1097
rect 156 -1098 157 -1097
rect 166 -1098 167 -1097
rect 702 -1098 703 -1097
rect 740 -1098 741 -1097
rect 779 -1098 780 -1097
rect 789 -1098 790 -1097
rect 863 -1098 864 -1097
rect 926 -1098 927 -1097
rect 933 -1098 934 -1097
rect 940 -1098 941 -1097
rect 1003 -1098 1004 -1097
rect 65 -1100 66 -1099
rect 72 -1100 73 -1099
rect 79 -1100 80 -1099
rect 205 -1100 206 -1099
rect 212 -1100 213 -1099
rect 219 -1100 220 -1099
rect 268 -1100 269 -1099
rect 331 -1100 332 -1099
rect 366 -1100 367 -1099
rect 394 -1100 395 -1099
rect 397 -1100 398 -1099
rect 443 -1100 444 -1099
rect 450 -1100 451 -1099
rect 513 -1100 514 -1099
rect 527 -1100 528 -1099
rect 635 -1100 636 -1099
rect 639 -1100 640 -1099
rect 702 -1100 703 -1099
rect 751 -1100 752 -1099
rect 814 -1100 815 -1099
rect 835 -1100 836 -1099
rect 856 -1100 857 -1099
rect 870 -1100 871 -1099
rect 940 -1100 941 -1099
rect 975 -1100 976 -1099
rect 989 -1100 990 -1099
rect 68 -1102 69 -1101
rect 502 -1102 503 -1101
rect 541 -1102 542 -1101
rect 954 -1102 955 -1101
rect 79 -1104 80 -1103
rect 93 -1104 94 -1103
rect 100 -1104 101 -1103
rect 107 -1104 108 -1103
rect 114 -1104 115 -1103
rect 198 -1104 199 -1103
rect 205 -1104 206 -1103
rect 261 -1104 262 -1103
rect 324 -1104 325 -1103
rect 1038 -1104 1039 -1103
rect 93 -1106 94 -1105
rect 285 -1106 286 -1105
rect 331 -1106 332 -1105
rect 352 -1106 353 -1105
rect 369 -1106 370 -1105
rect 394 -1106 395 -1105
rect 401 -1106 402 -1105
rect 520 -1106 521 -1105
rect 544 -1106 545 -1105
rect 821 -1106 822 -1105
rect 835 -1106 836 -1105
rect 842 -1106 843 -1105
rect 884 -1106 885 -1105
rect 933 -1106 934 -1105
rect 72 -1108 73 -1107
rect 352 -1108 353 -1107
rect 355 -1108 356 -1107
rect 821 -1108 822 -1107
rect 842 -1108 843 -1107
rect 1041 -1108 1042 -1107
rect 100 -1110 101 -1109
rect 142 -1110 143 -1109
rect 149 -1110 150 -1109
rect 156 -1110 157 -1109
rect 170 -1110 171 -1109
rect 219 -1110 220 -1109
rect 254 -1110 255 -1109
rect 401 -1110 402 -1109
rect 415 -1110 416 -1109
rect 443 -1110 444 -1109
rect 450 -1110 451 -1109
rect 737 -1110 738 -1109
rect 765 -1110 766 -1109
rect 800 -1110 801 -1109
rect 919 -1110 920 -1109
rect 975 -1110 976 -1109
rect 23 -1112 24 -1111
rect 170 -1112 171 -1111
rect 177 -1112 178 -1111
rect 411 -1112 412 -1111
rect 422 -1112 423 -1111
rect 527 -1112 528 -1111
rect 555 -1112 556 -1111
rect 744 -1112 745 -1111
rect 765 -1112 766 -1111
rect 1073 -1112 1074 -1111
rect 23 -1114 24 -1113
rect 37 -1114 38 -1113
rect 103 -1114 104 -1113
rect 688 -1114 689 -1113
rect 744 -1114 745 -1113
rect 758 -1114 759 -1113
rect 772 -1114 773 -1113
rect 884 -1114 885 -1113
rect 891 -1114 892 -1113
rect 919 -1114 920 -1113
rect 114 -1116 115 -1115
rect 128 -1116 129 -1115
rect 152 -1116 153 -1115
rect 313 -1116 314 -1115
rect 383 -1116 384 -1115
rect 1059 -1116 1060 -1115
rect 177 -1118 178 -1117
rect 303 -1118 304 -1117
rect 436 -1118 437 -1117
rect 541 -1118 542 -1117
rect 555 -1118 556 -1117
rect 1024 -1118 1025 -1117
rect 184 -1120 185 -1119
rect 261 -1120 262 -1119
rect 296 -1120 297 -1119
rect 422 -1120 423 -1119
rect 492 -1120 493 -1119
rect 733 -1120 734 -1119
rect 891 -1120 892 -1119
rect 912 -1120 913 -1119
rect 121 -1122 122 -1121
rect 296 -1122 297 -1121
rect 303 -1122 304 -1121
rect 345 -1122 346 -1121
rect 380 -1122 381 -1121
rect 436 -1122 437 -1121
rect 499 -1122 500 -1121
rect 863 -1122 864 -1121
rect 877 -1122 878 -1121
rect 912 -1122 913 -1121
rect 30 -1124 31 -1123
rect 345 -1124 346 -1123
rect 373 -1124 374 -1123
rect 380 -1124 381 -1123
rect 499 -1124 500 -1123
rect 1073 -1124 1074 -1123
rect 44 -1126 45 -1125
rect 373 -1126 374 -1125
rect 502 -1126 503 -1125
rect 786 -1126 787 -1125
rect 44 -1128 45 -1127
rect 572 -1128 573 -1127
rect 576 -1128 577 -1127
rect 597 -1128 598 -1127
rect 607 -1128 608 -1127
rect 618 -1128 619 -1127
rect 632 -1128 633 -1127
rect 758 -1128 759 -1127
rect 110 -1130 111 -1129
rect 877 -1130 878 -1129
rect 121 -1132 122 -1131
rect 289 -1132 290 -1131
rect 387 -1132 388 -1131
rect 632 -1132 633 -1131
rect 639 -1132 640 -1131
rect 709 -1132 710 -1131
rect 163 -1134 164 -1133
rect 289 -1134 290 -1133
rect 481 -1134 482 -1133
rect 786 -1134 787 -1133
rect 184 -1136 185 -1135
rect 408 -1136 409 -1135
rect 565 -1136 566 -1135
rect 814 -1136 815 -1135
rect 191 -1138 192 -1137
rect 275 -1138 276 -1137
rect 569 -1138 570 -1137
rect 611 -1138 612 -1137
rect 618 -1138 619 -1137
rect 646 -1138 647 -1137
rect 653 -1138 654 -1137
rect 772 -1138 773 -1137
rect 86 -1140 87 -1139
rect 191 -1140 192 -1139
rect 215 -1140 216 -1139
rect 485 -1140 486 -1139
rect 558 -1140 559 -1139
rect 646 -1140 647 -1139
rect 684 -1140 685 -1139
rect 961 -1140 962 -1139
rect 86 -1142 87 -1141
rect 317 -1142 318 -1141
rect 415 -1142 416 -1141
rect 611 -1142 612 -1141
rect 709 -1142 710 -1141
rect 716 -1142 717 -1141
rect 849 -1142 850 -1141
rect 961 -1142 962 -1141
rect 54 -1144 55 -1143
rect 716 -1144 717 -1143
rect 807 -1144 808 -1143
rect 849 -1144 850 -1143
rect 128 -1146 129 -1145
rect 558 -1146 559 -1145
rect 583 -1146 584 -1145
rect 681 -1146 682 -1145
rect 226 -1148 227 -1147
rect 387 -1148 388 -1147
rect 471 -1148 472 -1147
rect 681 -1148 682 -1147
rect 135 -1150 136 -1149
rect 226 -1150 227 -1149
rect 240 -1150 241 -1149
rect 576 -1150 577 -1149
rect 586 -1150 587 -1149
rect 870 -1150 871 -1149
rect 135 -1152 136 -1151
rect 534 -1152 535 -1151
rect 562 -1152 563 -1151
rect 583 -1152 584 -1151
rect 604 -1152 605 -1151
rect 653 -1152 654 -1151
rect 240 -1154 241 -1153
rect 338 -1154 339 -1153
rect 457 -1154 458 -1153
rect 471 -1154 472 -1153
rect 478 -1154 479 -1153
rect 485 -1154 486 -1153
rect 534 -1154 535 -1153
rect 695 -1154 696 -1153
rect 247 -1156 248 -1155
rect 254 -1156 255 -1155
rect 310 -1156 311 -1155
rect 338 -1156 339 -1155
rect 359 -1156 360 -1155
rect 457 -1156 458 -1155
rect 548 -1156 549 -1155
rect 604 -1156 605 -1155
rect 625 -1156 626 -1155
rect 807 -1156 808 -1155
rect 233 -1158 234 -1157
rect 247 -1158 248 -1157
rect 317 -1158 318 -1157
rect 464 -1158 465 -1157
rect 548 -1158 549 -1157
rect 660 -1158 661 -1157
rect 674 -1158 675 -1157
rect 695 -1158 696 -1157
rect 37 -1160 38 -1159
rect 233 -1160 234 -1159
rect 282 -1160 283 -1159
rect 674 -1160 675 -1159
rect 464 -1162 465 -1161
rect 625 -1162 626 -1161
rect 660 -1162 661 -1161
rect 730 -1162 731 -1161
rect 730 -1164 731 -1163
rect 1024 -1164 1025 -1163
rect 2 -1175 3 -1174
rect 145 -1175 146 -1174
rect 149 -1175 150 -1174
rect 205 -1175 206 -1174
rect 226 -1175 227 -1174
rect 310 -1175 311 -1174
rect 313 -1175 314 -1174
rect 821 -1175 822 -1174
rect 982 -1175 983 -1174
rect 1073 -1175 1074 -1174
rect 1115 -1175 1116 -1174
rect 1122 -1175 1123 -1174
rect 1129 -1175 1130 -1174
rect 1157 -1175 1158 -1174
rect 16 -1177 17 -1176
rect 275 -1177 276 -1176
rect 303 -1177 304 -1176
rect 408 -1177 409 -1176
rect 460 -1177 461 -1176
rect 471 -1177 472 -1176
rect 485 -1177 486 -1176
rect 488 -1177 489 -1176
rect 506 -1177 507 -1176
rect 520 -1177 521 -1176
rect 558 -1177 559 -1176
rect 695 -1177 696 -1176
rect 730 -1177 731 -1176
rect 933 -1177 934 -1176
rect 989 -1177 990 -1176
rect 1080 -1177 1081 -1176
rect 1150 -1177 1151 -1176
rect 1164 -1177 1165 -1176
rect 16 -1179 17 -1178
rect 380 -1179 381 -1178
rect 383 -1179 384 -1178
rect 478 -1179 479 -1178
rect 485 -1179 486 -1178
rect 604 -1179 605 -1178
rect 653 -1179 654 -1178
rect 730 -1179 731 -1178
rect 751 -1179 752 -1178
rect 856 -1179 857 -1178
rect 863 -1179 864 -1178
rect 933 -1179 934 -1178
rect 996 -1179 997 -1178
rect 1087 -1179 1088 -1178
rect 19 -1181 20 -1180
rect 247 -1181 248 -1180
rect 310 -1181 311 -1180
rect 317 -1181 318 -1180
rect 331 -1181 332 -1180
rect 355 -1181 356 -1180
rect 359 -1181 360 -1180
rect 821 -1181 822 -1180
rect 912 -1181 913 -1180
rect 989 -1181 990 -1180
rect 1003 -1181 1004 -1180
rect 1094 -1181 1095 -1180
rect 23 -1183 24 -1182
rect 37 -1183 38 -1182
rect 58 -1183 59 -1182
rect 940 -1183 941 -1182
rect 947 -1183 948 -1182
rect 1003 -1183 1004 -1182
rect 1017 -1183 1018 -1182
rect 1108 -1183 1109 -1182
rect 23 -1185 24 -1184
rect 362 -1185 363 -1184
rect 380 -1185 381 -1184
rect 401 -1185 402 -1184
rect 443 -1185 444 -1184
rect 471 -1185 472 -1184
rect 478 -1185 479 -1184
rect 537 -1185 538 -1184
rect 562 -1185 563 -1184
rect 807 -1185 808 -1184
rect 877 -1185 878 -1184
rect 940 -1185 941 -1184
rect 1031 -1185 1032 -1184
rect 1143 -1185 1144 -1184
rect 37 -1187 38 -1186
rect 352 -1187 353 -1186
rect 366 -1187 367 -1186
rect 401 -1187 402 -1186
rect 429 -1187 430 -1186
rect 443 -1187 444 -1186
rect 464 -1187 465 -1186
rect 667 -1187 668 -1186
rect 681 -1187 682 -1186
rect 751 -1187 752 -1186
rect 758 -1187 759 -1186
rect 807 -1187 808 -1186
rect 884 -1187 885 -1186
rect 947 -1187 948 -1186
rect 1041 -1187 1042 -1186
rect 1066 -1187 1067 -1186
rect 44 -1189 45 -1188
rect 366 -1189 367 -1188
rect 394 -1189 395 -1188
rect 418 -1189 419 -1188
rect 429 -1189 430 -1188
rect 642 -1189 643 -1188
rect 656 -1189 657 -1188
rect 1136 -1189 1137 -1188
rect 44 -1191 45 -1190
rect 65 -1191 66 -1190
rect 96 -1191 97 -1190
rect 527 -1191 528 -1190
rect 534 -1191 535 -1190
rect 758 -1191 759 -1190
rect 786 -1191 787 -1190
rect 968 -1191 969 -1190
rect 1045 -1191 1046 -1190
rect 1101 -1191 1102 -1190
rect 58 -1193 59 -1192
rect 128 -1193 129 -1192
rect 135 -1193 136 -1192
rect 481 -1193 482 -1192
rect 506 -1193 507 -1192
rect 1024 -1193 1025 -1192
rect 1052 -1193 1053 -1192
rect 1122 -1193 1123 -1192
rect 61 -1195 62 -1194
rect 135 -1195 136 -1194
rect 142 -1195 143 -1194
rect 415 -1195 416 -1194
rect 513 -1195 514 -1194
rect 604 -1195 605 -1194
rect 681 -1195 682 -1194
rect 961 -1195 962 -1194
rect 1059 -1195 1060 -1194
rect 1150 -1195 1151 -1194
rect 65 -1197 66 -1196
rect 194 -1197 195 -1196
rect 198 -1197 199 -1196
rect 285 -1197 286 -1196
rect 289 -1197 290 -1196
rect 352 -1197 353 -1196
rect 394 -1197 395 -1196
rect 555 -1197 556 -1196
rect 562 -1197 563 -1196
rect 576 -1197 577 -1196
rect 597 -1197 598 -1196
rect 660 -1197 661 -1196
rect 688 -1197 689 -1196
rect 1024 -1197 1025 -1196
rect 100 -1199 101 -1198
rect 107 -1199 108 -1198
rect 121 -1199 122 -1198
rect 359 -1199 360 -1198
rect 415 -1199 416 -1198
rect 502 -1199 503 -1198
rect 523 -1199 524 -1198
rect 1066 -1199 1067 -1198
rect 100 -1201 101 -1200
rect 114 -1201 115 -1200
rect 121 -1201 122 -1200
rect 611 -1201 612 -1200
rect 688 -1201 689 -1200
rect 716 -1201 717 -1200
rect 733 -1201 734 -1200
rect 863 -1201 864 -1200
rect 891 -1201 892 -1200
rect 1017 -1201 1018 -1200
rect 79 -1203 80 -1202
rect 114 -1203 115 -1202
rect 128 -1203 129 -1202
rect 177 -1203 178 -1202
rect 184 -1203 185 -1202
rect 205 -1203 206 -1202
rect 222 -1203 223 -1202
rect 275 -1203 276 -1202
rect 296 -1203 297 -1202
rect 331 -1203 332 -1202
rect 345 -1203 346 -1202
rect 772 -1203 773 -1202
rect 786 -1203 787 -1202
rect 1010 -1203 1011 -1202
rect 79 -1205 80 -1204
rect 450 -1205 451 -1204
rect 488 -1205 489 -1204
rect 513 -1205 514 -1204
rect 527 -1205 528 -1204
rect 632 -1205 633 -1204
rect 695 -1205 696 -1204
rect 765 -1205 766 -1204
rect 789 -1205 790 -1204
rect 1031 -1205 1032 -1204
rect 107 -1207 108 -1206
rect 324 -1207 325 -1206
rect 345 -1207 346 -1206
rect 373 -1207 374 -1206
rect 422 -1207 423 -1206
rect 772 -1207 773 -1206
rect 859 -1207 860 -1206
rect 1052 -1207 1053 -1206
rect 72 -1209 73 -1208
rect 324 -1209 325 -1208
rect 373 -1209 374 -1208
rect 814 -1209 815 -1208
rect 905 -1209 906 -1208
rect 961 -1209 962 -1208
rect 975 -1209 976 -1208
rect 1059 -1209 1060 -1208
rect 142 -1211 143 -1210
rect 369 -1211 370 -1210
rect 422 -1211 423 -1210
rect 492 -1211 493 -1210
rect 555 -1211 556 -1210
rect 1118 -1211 1119 -1210
rect 152 -1213 153 -1212
rect 464 -1213 465 -1212
rect 569 -1213 570 -1212
rect 611 -1213 612 -1212
rect 702 -1213 703 -1212
rect 891 -1213 892 -1212
rect 898 -1213 899 -1212
rect 975 -1213 976 -1212
rect 93 -1215 94 -1214
rect 702 -1215 703 -1214
rect 716 -1215 717 -1214
rect 877 -1215 878 -1214
rect 919 -1215 920 -1214
rect 996 -1215 997 -1214
rect 156 -1217 157 -1216
rect 219 -1217 220 -1216
rect 233 -1217 234 -1216
rect 884 -1217 885 -1216
rect 926 -1217 927 -1216
rect 1010 -1217 1011 -1216
rect 86 -1219 87 -1218
rect 233 -1219 234 -1218
rect 240 -1219 241 -1218
rect 296 -1219 297 -1218
rect 436 -1219 437 -1218
rect 450 -1219 451 -1218
rect 467 -1219 468 -1218
rect 569 -1219 570 -1218
rect 576 -1219 577 -1218
rect 590 -1219 591 -1218
rect 670 -1219 671 -1218
rect 919 -1219 920 -1218
rect 954 -1219 955 -1218
rect 1045 -1219 1046 -1218
rect 51 -1221 52 -1220
rect 436 -1221 437 -1220
rect 583 -1221 584 -1220
rect 590 -1221 591 -1220
rect 719 -1221 720 -1220
rect 954 -1221 955 -1220
rect 51 -1223 52 -1222
rect 268 -1223 269 -1222
rect 723 -1223 724 -1222
rect 765 -1223 766 -1222
rect 828 -1223 829 -1222
rect 898 -1223 899 -1222
rect 86 -1225 87 -1224
rect 170 -1225 171 -1224
rect 177 -1225 178 -1224
rect 387 -1225 388 -1224
rect 646 -1225 647 -1224
rect 723 -1225 724 -1224
rect 737 -1225 738 -1224
rect 912 -1225 913 -1224
rect 9 -1227 10 -1226
rect 170 -1227 171 -1226
rect 184 -1227 185 -1226
rect 261 -1227 262 -1226
rect 268 -1227 269 -1226
rect 282 -1227 283 -1226
rect 387 -1227 388 -1226
rect 625 -1227 626 -1226
rect 744 -1227 745 -1226
rect 814 -1227 815 -1226
rect 849 -1227 850 -1226
rect 926 -1227 927 -1226
rect 9 -1229 10 -1228
rect 30 -1229 31 -1228
rect 93 -1229 94 -1228
rect 583 -1229 584 -1228
rect 618 -1229 619 -1228
rect 646 -1229 647 -1228
rect 709 -1229 710 -1228
rect 744 -1229 745 -1228
rect 779 -1229 780 -1228
rect 849 -1229 850 -1228
rect 870 -1229 871 -1228
rect 905 -1229 906 -1228
rect 30 -1231 31 -1230
rect 289 -1231 290 -1230
rect 492 -1231 493 -1230
rect 737 -1231 738 -1230
rect 779 -1231 780 -1230
rect 793 -1231 794 -1230
rect 800 -1231 801 -1230
rect 870 -1231 871 -1230
rect 159 -1233 160 -1232
rect 600 -1233 601 -1232
rect 625 -1233 626 -1232
rect 667 -1233 668 -1232
rect 674 -1233 675 -1232
rect 709 -1233 710 -1232
rect 800 -1233 801 -1232
rect 1038 -1233 1039 -1232
rect 163 -1235 164 -1234
rect 982 -1235 983 -1234
rect 163 -1237 164 -1236
rect 212 -1237 213 -1236
rect 240 -1237 241 -1236
rect 348 -1237 349 -1236
rect 541 -1237 542 -1236
rect 618 -1237 619 -1236
rect 639 -1237 640 -1236
rect 793 -1237 794 -1236
rect 968 -1237 969 -1236
rect 1038 -1237 1039 -1236
rect 191 -1239 192 -1238
rect 226 -1239 227 -1238
rect 247 -1239 248 -1238
rect 303 -1239 304 -1238
rect 509 -1239 510 -1238
rect 541 -1239 542 -1238
rect 548 -1239 549 -1238
rect 674 -1239 675 -1238
rect 201 -1241 202 -1240
rect 317 -1241 318 -1240
rect 499 -1241 500 -1240
rect 548 -1241 549 -1240
rect 600 -1241 601 -1240
rect 842 -1241 843 -1240
rect 212 -1243 213 -1242
rect 271 -1243 272 -1242
rect 282 -1243 283 -1242
rect 338 -1243 339 -1242
rect 457 -1243 458 -1242
rect 499 -1243 500 -1242
rect 705 -1243 706 -1242
rect 842 -1243 843 -1242
rect 254 -1245 255 -1244
rect 261 -1245 262 -1244
rect 338 -1245 339 -1244
rect 684 -1245 685 -1244
rect 254 -1247 255 -1246
rect 376 -1247 377 -1246
rect 457 -1247 458 -1246
rect 660 -1247 661 -1246
rect 2 -1258 3 -1257
rect 72 -1258 73 -1257
rect 159 -1258 160 -1257
rect 387 -1258 388 -1257
rect 404 -1258 405 -1257
rect 527 -1258 528 -1257
rect 534 -1258 535 -1257
rect 618 -1258 619 -1257
rect 632 -1258 633 -1257
rect 814 -1258 815 -1257
rect 821 -1258 822 -1257
rect 1132 -1258 1133 -1257
rect 1164 -1258 1165 -1257
rect 1171 -1258 1172 -1257
rect 2 -1260 3 -1259
rect 51 -1260 52 -1259
rect 72 -1260 73 -1259
rect 268 -1260 269 -1259
rect 282 -1260 283 -1259
rect 303 -1260 304 -1259
rect 317 -1260 318 -1259
rect 439 -1260 440 -1259
rect 443 -1260 444 -1259
rect 446 -1260 447 -1259
rect 485 -1260 486 -1259
rect 702 -1260 703 -1259
rect 705 -1260 706 -1259
rect 1017 -1260 1018 -1259
rect 1024 -1260 1025 -1259
rect 1027 -1260 1028 -1259
rect 1122 -1260 1123 -1259
rect 1129 -1260 1130 -1259
rect 1157 -1260 1158 -1259
rect 1164 -1260 1165 -1259
rect 44 -1262 45 -1261
rect 215 -1262 216 -1261
rect 233 -1262 234 -1261
rect 292 -1262 293 -1261
rect 303 -1262 304 -1261
rect 555 -1262 556 -1261
rect 572 -1262 573 -1261
rect 870 -1262 871 -1261
rect 968 -1262 969 -1261
rect 1101 -1262 1102 -1261
rect 1122 -1262 1123 -1261
rect 1143 -1262 1144 -1261
rect 33 -1264 34 -1263
rect 44 -1264 45 -1263
rect 51 -1264 52 -1263
rect 170 -1264 171 -1263
rect 191 -1264 192 -1263
rect 1073 -1264 1074 -1263
rect 1143 -1264 1144 -1263
rect 1150 -1264 1151 -1263
rect 47 -1266 48 -1265
rect 1073 -1266 1074 -1265
rect 142 -1268 143 -1267
rect 814 -1268 815 -1267
rect 828 -1268 829 -1267
rect 877 -1268 878 -1267
rect 968 -1268 969 -1267
rect 982 -1268 983 -1267
rect 1024 -1268 1025 -1267
rect 1038 -1268 1039 -1267
rect 1052 -1268 1053 -1267
rect 1101 -1268 1102 -1267
rect 142 -1270 143 -1269
rect 212 -1270 213 -1269
rect 233 -1270 234 -1269
rect 296 -1270 297 -1269
rect 317 -1270 318 -1269
rect 411 -1270 412 -1269
rect 443 -1270 444 -1269
rect 464 -1270 465 -1269
rect 471 -1270 472 -1269
rect 485 -1270 486 -1269
rect 492 -1270 493 -1269
rect 604 -1270 605 -1269
rect 618 -1270 619 -1269
rect 674 -1270 675 -1269
rect 684 -1270 685 -1269
rect 961 -1270 962 -1269
rect 9 -1272 10 -1271
rect 212 -1272 213 -1271
rect 240 -1272 241 -1271
rect 369 -1272 370 -1271
rect 408 -1272 409 -1271
rect 506 -1272 507 -1271
rect 523 -1272 524 -1271
rect 898 -1272 899 -1271
rect 905 -1272 906 -1271
rect 961 -1272 962 -1271
rect 9 -1274 10 -1273
rect 254 -1274 255 -1273
rect 261 -1274 262 -1273
rect 271 -1274 272 -1273
rect 282 -1274 283 -1273
rect 660 -1274 661 -1273
rect 667 -1274 668 -1273
rect 989 -1274 990 -1273
rect 16 -1276 17 -1275
rect 604 -1276 605 -1275
rect 632 -1276 633 -1275
rect 751 -1276 752 -1275
rect 786 -1276 787 -1275
rect 807 -1276 808 -1275
rect 828 -1276 829 -1275
rect 1010 -1276 1011 -1275
rect 16 -1278 17 -1277
rect 180 -1278 181 -1277
rect 191 -1278 192 -1277
rect 205 -1278 206 -1277
rect 261 -1278 262 -1277
rect 537 -1278 538 -1277
rect 555 -1278 556 -1277
rect 562 -1278 563 -1277
rect 569 -1278 570 -1277
rect 982 -1278 983 -1277
rect 1010 -1278 1011 -1277
rect 1080 -1278 1081 -1277
rect 114 -1280 115 -1279
rect 240 -1280 241 -1279
rect 268 -1280 269 -1279
rect 338 -1280 339 -1279
rect 359 -1280 360 -1279
rect 387 -1280 388 -1279
rect 436 -1280 437 -1279
rect 807 -1280 808 -1279
rect 831 -1280 832 -1279
rect 1087 -1280 1088 -1279
rect 58 -1282 59 -1281
rect 359 -1282 360 -1281
rect 450 -1282 451 -1281
rect 464 -1282 465 -1281
rect 471 -1282 472 -1281
rect 513 -1282 514 -1281
rect 534 -1282 535 -1281
rect 737 -1282 738 -1281
rect 751 -1282 752 -1281
rect 849 -1282 850 -1281
rect 877 -1282 878 -1281
rect 891 -1282 892 -1281
rect 1066 -1282 1067 -1281
rect 1087 -1282 1088 -1281
rect 58 -1284 59 -1283
rect 194 -1284 195 -1283
rect 205 -1284 206 -1283
rect 247 -1284 248 -1283
rect 289 -1284 290 -1283
rect 373 -1284 374 -1283
rect 457 -1284 458 -1283
rect 1052 -1284 1053 -1283
rect 86 -1286 87 -1285
rect 114 -1286 115 -1285
rect 135 -1286 136 -1285
rect 289 -1286 290 -1285
rect 296 -1286 297 -1285
rect 429 -1286 430 -1285
rect 457 -1286 458 -1285
rect 562 -1286 563 -1285
rect 576 -1286 577 -1285
rect 597 -1286 598 -1285
rect 600 -1286 601 -1285
rect 912 -1286 913 -1285
rect 1027 -1286 1028 -1285
rect 1038 -1286 1039 -1285
rect 1045 -1286 1046 -1285
rect 1066 -1286 1067 -1285
rect 86 -1288 87 -1287
rect 100 -1288 101 -1287
rect 107 -1288 108 -1287
rect 135 -1288 136 -1287
rect 156 -1288 157 -1287
rect 870 -1288 871 -1287
rect 891 -1288 892 -1287
rect 947 -1288 948 -1287
rect 1003 -1288 1004 -1287
rect 1045 -1288 1046 -1287
rect 26 -1290 27 -1289
rect 156 -1290 157 -1289
rect 163 -1290 164 -1289
rect 254 -1290 255 -1289
rect 275 -1290 276 -1289
rect 429 -1290 430 -1289
rect 478 -1290 479 -1289
rect 737 -1290 738 -1289
rect 796 -1290 797 -1289
rect 856 -1290 857 -1289
rect 912 -1290 913 -1289
rect 933 -1290 934 -1289
rect 947 -1290 948 -1289
rect 989 -1290 990 -1289
rect 1003 -1290 1004 -1289
rect 1031 -1290 1032 -1289
rect 37 -1292 38 -1291
rect 275 -1292 276 -1291
rect 324 -1292 325 -1291
rect 569 -1292 570 -1291
rect 590 -1292 591 -1291
rect 674 -1292 675 -1291
rect 688 -1292 689 -1291
rect 821 -1292 822 -1291
rect 835 -1292 836 -1291
rect 905 -1292 906 -1291
rect 933 -1292 934 -1291
rect 954 -1292 955 -1291
rect 1031 -1292 1032 -1291
rect 1136 -1292 1137 -1291
rect 37 -1294 38 -1293
rect 184 -1294 185 -1293
rect 247 -1294 248 -1293
rect 394 -1294 395 -1293
rect 408 -1294 409 -1293
rect 576 -1294 577 -1293
rect 607 -1294 608 -1293
rect 1080 -1294 1081 -1293
rect 1136 -1294 1137 -1293
rect 1157 -1294 1158 -1293
rect 100 -1296 101 -1295
rect 310 -1296 311 -1295
rect 324 -1296 325 -1295
rect 422 -1296 423 -1295
rect 495 -1296 496 -1295
rect 688 -1296 689 -1295
rect 716 -1296 717 -1295
rect 1115 -1296 1116 -1295
rect 107 -1298 108 -1297
rect 128 -1298 129 -1297
rect 170 -1298 171 -1297
rect 635 -1298 636 -1297
rect 639 -1298 640 -1297
rect 1017 -1298 1018 -1297
rect 1108 -1298 1109 -1297
rect 1115 -1298 1116 -1297
rect 30 -1300 31 -1299
rect 128 -1300 129 -1299
rect 184 -1300 185 -1299
rect 187 -1300 188 -1299
rect 310 -1300 311 -1299
rect 415 -1300 416 -1299
rect 499 -1300 500 -1299
rect 527 -1300 528 -1299
rect 541 -1300 542 -1299
rect 590 -1300 591 -1299
rect 621 -1300 622 -1299
rect 831 -1300 832 -1299
rect 849 -1300 850 -1299
rect 975 -1300 976 -1299
rect 1094 -1300 1095 -1299
rect 1108 -1300 1109 -1299
rect 65 -1302 66 -1301
rect 415 -1302 416 -1301
rect 513 -1302 514 -1301
rect 520 -1302 521 -1301
rect 642 -1302 643 -1301
rect 1059 -1302 1060 -1301
rect 121 -1304 122 -1303
rect 639 -1304 640 -1303
rect 646 -1304 647 -1303
rect 667 -1304 668 -1303
rect 670 -1304 671 -1303
rect 765 -1304 766 -1303
rect 779 -1304 780 -1303
rect 835 -1304 836 -1303
rect 842 -1304 843 -1303
rect 1094 -1304 1095 -1303
rect 79 -1306 80 -1305
rect 121 -1306 122 -1305
rect 338 -1306 339 -1305
rect 628 -1306 629 -1305
rect 646 -1306 647 -1305
rect 758 -1306 759 -1305
rect 772 -1306 773 -1305
rect 779 -1306 780 -1305
rect 800 -1306 801 -1305
rect 898 -1306 899 -1305
rect 940 -1306 941 -1305
rect 954 -1306 955 -1305
rect 975 -1306 976 -1305
rect 996 -1306 997 -1305
rect 79 -1308 80 -1307
rect 96 -1308 97 -1307
rect 345 -1308 346 -1307
rect 499 -1308 500 -1307
rect 506 -1308 507 -1307
rect 772 -1308 773 -1307
rect 842 -1308 843 -1307
rect 863 -1308 864 -1307
rect 198 -1310 199 -1309
rect 345 -1310 346 -1309
rect 348 -1310 349 -1309
rect 1059 -1310 1060 -1309
rect 177 -1312 178 -1311
rect 198 -1312 199 -1311
rect 352 -1312 353 -1311
rect 422 -1312 423 -1311
rect 436 -1312 437 -1311
rect 940 -1312 941 -1311
rect 352 -1314 353 -1313
rect 380 -1314 381 -1313
rect 394 -1314 395 -1313
rect 541 -1314 542 -1313
rect 597 -1314 598 -1313
rect 996 -1314 997 -1313
rect 366 -1316 367 -1315
rect 765 -1316 766 -1315
rect 856 -1316 857 -1315
rect 919 -1316 920 -1315
rect 23 -1318 24 -1317
rect 919 -1318 920 -1317
rect 331 -1320 332 -1319
rect 366 -1320 367 -1319
rect 380 -1320 381 -1319
rect 401 -1320 402 -1319
rect 520 -1320 521 -1319
rect 660 -1320 661 -1319
rect 709 -1320 710 -1319
rect 800 -1320 801 -1319
rect 149 -1322 150 -1321
rect 331 -1322 332 -1321
rect 401 -1322 402 -1321
rect 460 -1322 461 -1321
rect 625 -1322 626 -1321
rect 709 -1322 710 -1321
rect 723 -1322 724 -1321
rect 863 -1322 864 -1321
rect 149 -1324 150 -1323
rect 681 -1324 682 -1323
rect 695 -1324 696 -1323
rect 723 -1324 724 -1323
rect 733 -1324 734 -1323
rect 884 -1324 885 -1323
rect 103 -1326 104 -1325
rect 695 -1326 696 -1325
rect 744 -1326 745 -1325
rect 758 -1326 759 -1325
rect 884 -1326 885 -1325
rect 926 -1326 927 -1325
rect 460 -1328 461 -1327
rect 509 -1328 510 -1327
rect 544 -1328 545 -1327
rect 926 -1328 927 -1327
rect 653 -1330 654 -1329
rect 789 -1330 790 -1329
rect 492 -1332 493 -1331
rect 653 -1332 654 -1331
rect 656 -1332 657 -1331
rect 793 -1332 794 -1331
rect 548 -1334 549 -1333
rect 793 -1334 794 -1333
rect 548 -1336 549 -1335
rect 583 -1336 584 -1335
rect 730 -1336 731 -1335
rect 744 -1336 745 -1335
rect 583 -1338 584 -1337
rect 611 -1338 612 -1337
rect 478 -1340 479 -1339
rect 611 -1340 612 -1339
rect 2 -1351 3 -1350
rect 432 -1351 433 -1350
rect 436 -1351 437 -1350
rect 688 -1351 689 -1350
rect 733 -1351 734 -1350
rect 1045 -1351 1046 -1350
rect 1101 -1351 1102 -1350
rect 1150 -1351 1151 -1350
rect 1153 -1351 1154 -1350
rect 1164 -1351 1165 -1350
rect 2 -1353 3 -1352
rect 121 -1353 122 -1352
rect 135 -1353 136 -1352
rect 334 -1353 335 -1352
rect 359 -1353 360 -1352
rect 523 -1353 524 -1352
rect 527 -1353 528 -1352
rect 947 -1353 948 -1352
rect 950 -1353 951 -1352
rect 1129 -1353 1130 -1352
rect 1136 -1353 1137 -1352
rect 1171 -1353 1172 -1352
rect 9 -1355 10 -1354
rect 163 -1355 164 -1354
rect 215 -1355 216 -1354
rect 415 -1355 416 -1354
rect 506 -1355 507 -1354
rect 541 -1355 542 -1354
rect 544 -1355 545 -1354
rect 646 -1355 647 -1354
rect 688 -1355 689 -1354
rect 975 -1355 976 -1354
rect 996 -1355 997 -1354
rect 1066 -1355 1067 -1354
rect 16 -1357 17 -1356
rect 411 -1357 412 -1356
rect 506 -1357 507 -1356
rect 632 -1357 633 -1356
rect 681 -1357 682 -1356
rect 975 -1357 976 -1356
rect 1031 -1357 1032 -1356
rect 1066 -1357 1067 -1356
rect 23 -1359 24 -1358
rect 446 -1359 447 -1358
rect 520 -1359 521 -1358
rect 842 -1359 843 -1358
rect 1031 -1359 1032 -1358
rect 1094 -1359 1095 -1358
rect 26 -1361 27 -1360
rect 240 -1361 241 -1360
rect 275 -1361 276 -1360
rect 527 -1361 528 -1360
rect 537 -1361 538 -1360
rect 898 -1361 899 -1360
rect 1045 -1361 1046 -1360
rect 1143 -1361 1144 -1360
rect 33 -1363 34 -1362
rect 58 -1363 59 -1362
rect 65 -1363 66 -1362
rect 485 -1363 486 -1362
rect 562 -1363 563 -1362
rect 646 -1363 647 -1362
rect 681 -1363 682 -1362
rect 751 -1363 752 -1362
rect 772 -1363 773 -1362
rect 905 -1363 906 -1362
rect 44 -1365 45 -1364
rect 68 -1365 69 -1364
rect 93 -1365 94 -1364
rect 107 -1365 108 -1364
rect 121 -1365 122 -1364
rect 1080 -1365 1081 -1364
rect 44 -1367 45 -1366
rect 86 -1367 87 -1366
rect 100 -1367 101 -1366
rect 205 -1367 206 -1366
rect 212 -1367 213 -1366
rect 1094 -1367 1095 -1366
rect 16 -1369 17 -1368
rect 100 -1369 101 -1368
rect 103 -1369 104 -1368
rect 275 -1369 276 -1368
rect 289 -1369 290 -1368
rect 422 -1369 423 -1368
rect 485 -1369 486 -1368
rect 674 -1369 675 -1368
rect 751 -1369 752 -1368
rect 758 -1369 759 -1368
rect 772 -1369 773 -1368
rect 835 -1369 836 -1368
rect 842 -1369 843 -1368
rect 856 -1369 857 -1368
rect 898 -1369 899 -1368
rect 1024 -1369 1025 -1368
rect 51 -1371 52 -1370
rect 460 -1371 461 -1370
rect 492 -1371 493 -1370
rect 1080 -1371 1081 -1370
rect 51 -1373 52 -1372
rect 352 -1373 353 -1372
rect 359 -1373 360 -1372
rect 380 -1373 381 -1372
rect 387 -1373 388 -1372
rect 905 -1373 906 -1372
rect 58 -1375 59 -1374
rect 247 -1375 248 -1374
rect 268 -1375 269 -1374
rect 380 -1375 381 -1374
rect 387 -1375 388 -1374
rect 499 -1375 500 -1374
rect 600 -1375 601 -1374
rect 1052 -1375 1053 -1374
rect 65 -1377 66 -1376
rect 114 -1377 115 -1376
rect 128 -1377 129 -1376
rect 240 -1377 241 -1376
rect 247 -1377 248 -1376
rect 296 -1377 297 -1376
rect 303 -1377 304 -1376
rect 495 -1377 496 -1376
rect 569 -1377 570 -1376
rect 1052 -1377 1053 -1376
rect 37 -1379 38 -1378
rect 128 -1379 129 -1378
rect 135 -1379 136 -1378
rect 331 -1379 332 -1378
rect 408 -1379 409 -1378
rect 450 -1379 451 -1378
rect 611 -1379 612 -1378
rect 968 -1379 969 -1378
rect 37 -1381 38 -1380
rect 324 -1381 325 -1380
rect 331 -1381 332 -1380
rect 415 -1381 416 -1380
rect 422 -1381 423 -1380
rect 569 -1381 570 -1380
rect 611 -1381 612 -1380
rect 695 -1381 696 -1380
rect 758 -1381 759 -1380
rect 821 -1381 822 -1380
rect 828 -1381 829 -1380
rect 1108 -1381 1109 -1380
rect 72 -1383 73 -1382
rect 86 -1383 87 -1382
rect 103 -1383 104 -1382
rect 177 -1383 178 -1382
rect 187 -1383 188 -1382
rect 408 -1383 409 -1382
rect 443 -1383 444 -1382
rect 450 -1383 451 -1382
rect 509 -1383 510 -1382
rect 968 -1383 969 -1382
rect 1108 -1383 1109 -1382
rect 1157 -1383 1158 -1382
rect 72 -1385 73 -1384
rect 555 -1385 556 -1384
rect 614 -1385 615 -1384
rect 814 -1385 815 -1384
rect 821 -1385 822 -1384
rect 877 -1385 878 -1384
rect 79 -1387 80 -1386
rect 555 -1387 556 -1386
rect 625 -1387 626 -1386
rect 954 -1387 955 -1386
rect 79 -1389 80 -1388
rect 198 -1389 199 -1388
rect 226 -1389 227 -1388
rect 348 -1389 349 -1388
rect 618 -1389 619 -1388
rect 625 -1389 626 -1388
rect 632 -1389 633 -1388
rect 653 -1389 654 -1388
rect 660 -1389 661 -1388
rect 835 -1389 836 -1388
rect 849 -1389 850 -1388
rect 954 -1389 955 -1388
rect 110 -1391 111 -1390
rect 1024 -1391 1025 -1390
rect 149 -1393 150 -1392
rect 404 -1393 405 -1392
rect 653 -1393 654 -1392
rect 807 -1393 808 -1392
rect 814 -1393 815 -1392
rect 1062 -1393 1063 -1392
rect 149 -1395 150 -1394
rect 317 -1395 318 -1394
rect 324 -1395 325 -1394
rect 429 -1395 430 -1394
rect 660 -1395 661 -1394
rect 667 -1395 668 -1394
rect 674 -1395 675 -1394
rect 716 -1395 717 -1394
rect 775 -1395 776 -1394
rect 786 -1395 787 -1394
rect 828 -1395 829 -1394
rect 933 -1395 934 -1394
rect 156 -1397 157 -1396
rect 730 -1397 731 -1396
rect 786 -1397 787 -1396
rect 870 -1397 871 -1396
rect 877 -1397 878 -1396
rect 912 -1397 913 -1396
rect 933 -1397 934 -1396
rect 1087 -1397 1088 -1396
rect 156 -1399 157 -1398
rect 261 -1399 262 -1398
rect 282 -1399 283 -1398
rect 667 -1399 668 -1398
rect 695 -1399 696 -1398
rect 723 -1399 724 -1398
rect 856 -1399 857 -1398
rect 1059 -1399 1060 -1398
rect 163 -1401 164 -1400
rect 184 -1401 185 -1400
rect 191 -1401 192 -1400
rect 205 -1401 206 -1400
rect 219 -1401 220 -1400
rect 282 -1401 283 -1400
rect 292 -1401 293 -1400
rect 495 -1401 496 -1400
rect 716 -1401 717 -1400
rect 765 -1401 766 -1400
rect 870 -1401 871 -1400
rect 884 -1401 885 -1400
rect 912 -1401 913 -1400
rect 1010 -1401 1011 -1400
rect 177 -1403 178 -1402
rect 352 -1403 353 -1402
rect 534 -1403 535 -1402
rect 884 -1403 885 -1402
rect 926 -1403 927 -1402
rect 1087 -1403 1088 -1402
rect 194 -1405 195 -1404
rect 268 -1405 269 -1404
rect 296 -1405 297 -1404
rect 502 -1405 503 -1404
rect 723 -1405 724 -1404
rect 737 -1405 738 -1404
rect 765 -1405 766 -1404
rect 779 -1405 780 -1404
rect 891 -1405 892 -1404
rect 926 -1405 927 -1404
rect 961 -1405 962 -1404
rect 1010 -1405 1011 -1404
rect 198 -1407 199 -1406
rect 604 -1407 605 -1406
rect 737 -1407 738 -1406
rect 744 -1407 745 -1406
rect 779 -1407 780 -1406
rect 800 -1407 801 -1406
rect 961 -1407 962 -1406
rect 982 -1407 983 -1406
rect 30 -1409 31 -1408
rect 800 -1409 801 -1408
rect 982 -1409 983 -1408
rect 989 -1409 990 -1408
rect 30 -1411 31 -1410
rect 142 -1411 143 -1410
rect 219 -1411 220 -1410
rect 233 -1411 234 -1410
rect 254 -1411 255 -1410
rect 261 -1411 262 -1410
rect 310 -1411 311 -1410
rect 439 -1411 440 -1410
rect 471 -1411 472 -1410
rect 534 -1411 535 -1410
rect 604 -1411 605 -1410
rect 709 -1411 710 -1410
rect 793 -1411 794 -1410
rect 891 -1411 892 -1410
rect 989 -1411 990 -1410
rect 1003 -1411 1004 -1410
rect 93 -1413 94 -1412
rect 744 -1413 745 -1412
rect 1003 -1413 1004 -1412
rect 1073 -1413 1074 -1412
rect 142 -1415 143 -1414
rect 170 -1415 171 -1414
rect 226 -1415 227 -1414
rect 457 -1415 458 -1414
rect 464 -1415 465 -1414
rect 471 -1415 472 -1414
rect 639 -1415 640 -1414
rect 709 -1415 710 -1414
rect 1073 -1415 1074 -1414
rect 1122 -1415 1123 -1414
rect 96 -1417 97 -1416
rect 170 -1417 171 -1416
rect 233 -1417 234 -1416
rect 401 -1417 402 -1416
rect 457 -1417 458 -1416
rect 691 -1417 692 -1416
rect 702 -1417 703 -1416
rect 793 -1417 794 -1416
rect 254 -1419 255 -1418
rect 849 -1419 850 -1418
rect 303 -1421 304 -1420
rect 439 -1421 440 -1420
rect 464 -1421 465 -1420
rect 576 -1421 577 -1420
rect 702 -1421 703 -1420
rect 807 -1421 808 -1420
rect 310 -1423 311 -1422
rect 597 -1423 598 -1422
rect 317 -1425 318 -1424
rect 579 -1425 580 -1424
rect 338 -1427 339 -1426
rect 618 -1427 619 -1426
rect 338 -1429 339 -1428
rect 488 -1429 489 -1428
rect 499 -1429 500 -1428
rect 639 -1429 640 -1428
rect 401 -1431 402 -1430
rect 562 -1431 563 -1430
rect 576 -1431 577 -1430
rect 863 -1431 864 -1430
rect 345 -1433 346 -1432
rect 863 -1433 864 -1432
rect 345 -1435 346 -1434
rect 478 -1435 479 -1434
rect 478 -1437 479 -1436
rect 590 -1437 591 -1436
rect 583 -1439 584 -1438
rect 590 -1439 591 -1438
rect 548 -1441 549 -1440
rect 583 -1441 584 -1440
rect 548 -1443 549 -1442
rect 1017 -1443 1018 -1442
rect 1017 -1445 1018 -1444
rect 1038 -1445 1039 -1444
rect 1038 -1447 1039 -1446
rect 1115 -1447 1116 -1446
rect 9 -1458 10 -1457
rect 467 -1458 468 -1457
rect 481 -1458 482 -1457
rect 604 -1458 605 -1457
rect 611 -1458 612 -1457
rect 996 -1458 997 -1457
rect 1010 -1458 1011 -1457
rect 1059 -1458 1060 -1457
rect 16 -1460 17 -1459
rect 495 -1460 496 -1459
rect 499 -1460 500 -1459
rect 947 -1460 948 -1459
rect 996 -1460 997 -1459
rect 1073 -1460 1074 -1459
rect 16 -1462 17 -1461
rect 331 -1462 332 -1461
rect 352 -1462 353 -1461
rect 523 -1462 524 -1461
rect 551 -1462 552 -1461
rect 674 -1462 675 -1461
rect 681 -1462 682 -1461
rect 702 -1462 703 -1461
rect 744 -1462 745 -1461
rect 1045 -1462 1046 -1461
rect 1062 -1462 1063 -1461
rect 1073 -1462 1074 -1461
rect 30 -1464 31 -1463
rect 187 -1464 188 -1463
rect 198 -1464 199 -1463
rect 548 -1464 549 -1463
rect 569 -1464 570 -1463
rect 660 -1464 661 -1463
rect 681 -1464 682 -1463
rect 765 -1464 766 -1463
rect 856 -1464 857 -1463
rect 912 -1464 913 -1463
rect 947 -1464 948 -1463
rect 1031 -1464 1032 -1463
rect 23 -1466 24 -1465
rect 198 -1466 199 -1465
rect 257 -1466 258 -1465
rect 261 -1466 262 -1465
rect 289 -1466 290 -1465
rect 411 -1466 412 -1465
rect 415 -1466 416 -1465
rect 429 -1466 430 -1465
rect 436 -1466 437 -1465
rect 506 -1466 507 -1465
rect 516 -1466 517 -1465
rect 758 -1466 759 -1465
rect 765 -1466 766 -1465
rect 835 -1466 836 -1465
rect 856 -1466 857 -1465
rect 961 -1466 962 -1465
rect 1017 -1466 1018 -1465
rect 1020 -1466 1021 -1465
rect 23 -1468 24 -1467
rect 254 -1468 255 -1467
rect 292 -1468 293 -1467
rect 359 -1468 360 -1467
rect 387 -1468 388 -1467
rect 499 -1468 500 -1467
rect 502 -1468 503 -1467
rect 695 -1468 696 -1467
rect 747 -1468 748 -1467
rect 877 -1468 878 -1467
rect 884 -1468 885 -1467
rect 1010 -1468 1011 -1467
rect 1017 -1468 1018 -1467
rect 1038 -1468 1039 -1467
rect 33 -1470 34 -1469
rect 716 -1470 717 -1469
rect 758 -1470 759 -1469
rect 786 -1470 787 -1469
rect 835 -1470 836 -1469
rect 954 -1470 955 -1469
rect 1020 -1470 1021 -1469
rect 1038 -1470 1039 -1469
rect 44 -1472 45 -1471
rect 110 -1472 111 -1471
rect 114 -1472 115 -1471
rect 268 -1472 269 -1471
rect 310 -1472 311 -1471
rect 509 -1472 510 -1471
rect 541 -1472 542 -1471
rect 548 -1472 549 -1471
rect 569 -1472 570 -1471
rect 663 -1472 664 -1471
rect 695 -1472 696 -1471
rect 919 -1472 920 -1471
rect 933 -1472 934 -1471
rect 961 -1472 962 -1471
rect 30 -1474 31 -1473
rect 44 -1474 45 -1473
rect 51 -1474 52 -1473
rect 215 -1474 216 -1473
rect 254 -1474 255 -1473
rect 296 -1474 297 -1473
rect 310 -1474 311 -1473
rect 327 -1474 328 -1473
rect 331 -1474 332 -1473
rect 373 -1474 374 -1473
rect 387 -1474 388 -1473
rect 478 -1474 479 -1473
rect 485 -1474 486 -1473
rect 667 -1474 668 -1473
rect 730 -1474 731 -1473
rect 919 -1474 920 -1473
rect 954 -1474 955 -1473
rect 1094 -1474 1095 -1473
rect 2 -1476 3 -1475
rect 215 -1476 216 -1475
rect 296 -1476 297 -1475
rect 513 -1476 514 -1475
rect 541 -1476 542 -1475
rect 639 -1476 640 -1475
rect 730 -1476 731 -1475
rect 751 -1476 752 -1475
rect 786 -1476 787 -1475
rect 891 -1476 892 -1475
rect 912 -1476 913 -1475
rect 989 -1476 990 -1475
rect 1094 -1476 1095 -1475
rect 1108 -1476 1109 -1475
rect 2 -1478 3 -1477
rect 96 -1478 97 -1477
rect 103 -1478 104 -1477
rect 674 -1478 675 -1477
rect 688 -1478 689 -1477
rect 989 -1478 990 -1477
rect 51 -1480 52 -1479
rect 324 -1480 325 -1479
rect 345 -1480 346 -1479
rect 415 -1480 416 -1479
rect 422 -1480 423 -1479
rect 506 -1480 507 -1479
rect 576 -1480 577 -1479
rect 821 -1480 822 -1479
rect 859 -1480 860 -1479
rect 933 -1480 934 -1479
rect 37 -1482 38 -1481
rect 324 -1482 325 -1481
rect 373 -1482 374 -1481
rect 380 -1482 381 -1481
rect 394 -1482 395 -1481
rect 404 -1482 405 -1481
rect 408 -1482 409 -1481
rect 744 -1482 745 -1481
rect 821 -1482 822 -1481
rect 905 -1482 906 -1481
rect 9 -1484 10 -1483
rect 37 -1484 38 -1483
rect 65 -1484 66 -1483
rect 191 -1484 192 -1483
rect 233 -1484 234 -1483
rect 751 -1484 752 -1483
rect 863 -1484 864 -1483
rect 1045 -1484 1046 -1483
rect 58 -1486 59 -1485
rect 191 -1486 192 -1485
rect 226 -1486 227 -1485
rect 233 -1486 234 -1485
rect 366 -1486 367 -1485
rect 380 -1486 381 -1485
rect 401 -1486 402 -1485
rect 614 -1486 615 -1485
rect 639 -1486 640 -1485
rect 709 -1486 710 -1485
rect 807 -1486 808 -1485
rect 863 -1486 864 -1485
rect 870 -1486 871 -1485
rect 891 -1486 892 -1485
rect 58 -1488 59 -1487
rect 142 -1488 143 -1487
rect 163 -1488 164 -1487
rect 180 -1488 181 -1487
rect 226 -1488 227 -1487
rect 289 -1488 290 -1487
rect 422 -1488 423 -1487
rect 670 -1488 671 -1487
rect 807 -1488 808 -1487
rect 940 -1488 941 -1487
rect 65 -1490 66 -1489
rect 450 -1490 451 -1489
rect 464 -1490 465 -1489
rect 611 -1490 612 -1489
rect 870 -1490 871 -1489
rect 968 -1490 969 -1489
rect 72 -1492 73 -1491
rect 268 -1492 269 -1491
rect 432 -1492 433 -1491
rect 716 -1492 717 -1491
rect 877 -1492 878 -1491
rect 982 -1492 983 -1491
rect 72 -1494 73 -1493
rect 219 -1494 220 -1493
rect 439 -1494 440 -1493
rect 814 -1494 815 -1493
rect 884 -1494 885 -1493
rect 898 -1494 899 -1493
rect 940 -1494 941 -1493
rect 1024 -1494 1025 -1493
rect 79 -1496 80 -1495
rect 334 -1496 335 -1495
rect 443 -1496 444 -1495
rect 471 -1496 472 -1495
rect 485 -1496 486 -1495
rect 793 -1496 794 -1495
rect 814 -1496 815 -1495
rect 828 -1496 829 -1495
rect 968 -1496 969 -1495
rect 1003 -1496 1004 -1495
rect 1024 -1496 1025 -1495
rect 1080 -1496 1081 -1495
rect 79 -1498 80 -1497
rect 247 -1498 248 -1497
rect 443 -1498 444 -1497
rect 562 -1498 563 -1497
rect 590 -1498 591 -1497
rect 604 -1498 605 -1497
rect 793 -1498 794 -1497
rect 849 -1498 850 -1497
rect 982 -1498 983 -1497
rect 1052 -1498 1053 -1497
rect 86 -1500 87 -1499
rect 145 -1500 146 -1499
rect 163 -1500 164 -1499
rect 520 -1500 521 -1499
rect 534 -1500 535 -1499
rect 590 -1500 591 -1499
rect 597 -1500 598 -1499
rect 646 -1500 647 -1499
rect 779 -1500 780 -1499
rect 849 -1500 850 -1499
rect 1003 -1500 1004 -1499
rect 1066 -1500 1067 -1499
rect 86 -1502 87 -1501
rect 149 -1502 150 -1501
rect 166 -1502 167 -1501
rect 632 -1502 633 -1501
rect 646 -1502 647 -1501
rect 737 -1502 738 -1501
rect 772 -1502 773 -1501
rect 779 -1502 780 -1501
rect 828 -1502 829 -1501
rect 842 -1502 843 -1501
rect 107 -1504 108 -1503
rect 170 -1504 171 -1503
rect 177 -1504 178 -1503
rect 492 -1504 493 -1503
rect 534 -1504 535 -1503
rect 709 -1504 710 -1503
rect 842 -1504 843 -1503
rect 926 -1504 927 -1503
rect 93 -1506 94 -1505
rect 107 -1506 108 -1505
rect 114 -1506 115 -1505
rect 691 -1506 692 -1505
rect 705 -1506 706 -1505
rect 926 -1506 927 -1505
rect 93 -1508 94 -1507
rect 600 -1508 601 -1507
rect 677 -1508 678 -1507
rect 737 -1508 738 -1507
rect 121 -1510 122 -1509
rect 579 -1510 580 -1509
rect 691 -1510 692 -1509
rect 800 -1510 801 -1509
rect 124 -1512 125 -1511
rect 240 -1512 241 -1511
rect 247 -1512 248 -1511
rect 618 -1512 619 -1511
rect 800 -1512 801 -1511
rect 975 -1512 976 -1511
rect 128 -1514 129 -1513
rect 261 -1514 262 -1513
rect 366 -1514 367 -1513
rect 562 -1514 563 -1513
rect 618 -1514 619 -1513
rect 723 -1514 724 -1513
rect 128 -1516 129 -1515
rect 184 -1516 185 -1515
rect 212 -1516 213 -1515
rect 975 -1516 976 -1515
rect 100 -1518 101 -1517
rect 212 -1518 213 -1517
rect 219 -1518 220 -1517
rect 408 -1518 409 -1517
rect 450 -1518 451 -1517
rect 537 -1518 538 -1517
rect 555 -1518 556 -1517
rect 905 -1518 906 -1517
rect 135 -1520 136 -1519
rect 352 -1520 353 -1519
rect 359 -1520 360 -1519
rect 723 -1520 724 -1519
rect 135 -1522 136 -1521
rect 338 -1522 339 -1521
rect 457 -1522 458 -1521
rect 632 -1522 633 -1521
rect 149 -1524 150 -1523
rect 625 -1524 626 -1523
rect 156 -1526 157 -1525
rect 170 -1526 171 -1525
rect 177 -1526 178 -1525
rect 394 -1526 395 -1525
rect 457 -1526 458 -1525
rect 576 -1526 577 -1525
rect 625 -1526 626 -1525
rect 653 -1526 654 -1525
rect 156 -1528 157 -1527
rect 898 -1528 899 -1527
rect 184 -1530 185 -1529
rect 205 -1530 206 -1529
rect 240 -1530 241 -1529
rect 317 -1530 318 -1529
rect 338 -1530 339 -1529
rect 1031 -1530 1032 -1529
rect 194 -1532 195 -1531
rect 653 -1532 654 -1531
rect 205 -1534 206 -1533
rect 345 -1534 346 -1533
rect 527 -1534 528 -1533
rect 555 -1534 556 -1533
rect 275 -1536 276 -1535
rect 317 -1536 318 -1535
rect 527 -1536 528 -1535
rect 583 -1536 584 -1535
rect 513 -1538 514 -1537
rect 583 -1538 584 -1537
rect 2 -1549 3 -1548
rect 247 -1549 248 -1548
rect 254 -1549 255 -1548
rect 289 -1549 290 -1548
rect 352 -1549 353 -1548
rect 359 -1549 360 -1548
rect 376 -1549 377 -1548
rect 436 -1549 437 -1548
rect 457 -1549 458 -1548
rect 919 -1549 920 -1548
rect 940 -1549 941 -1548
rect 1010 -1549 1011 -1548
rect 1034 -1549 1035 -1548
rect 1038 -1549 1039 -1548
rect 1045 -1549 1046 -1548
rect 1101 -1549 1102 -1548
rect 5 -1551 6 -1550
rect 100 -1551 101 -1550
rect 145 -1551 146 -1550
rect 1052 -1551 1053 -1550
rect 1059 -1551 1060 -1550
rect 1108 -1551 1109 -1550
rect 9 -1553 10 -1552
rect 250 -1553 251 -1552
rect 261 -1553 262 -1552
rect 436 -1553 437 -1552
rect 464 -1553 465 -1552
rect 695 -1553 696 -1552
rect 772 -1553 773 -1552
rect 891 -1553 892 -1552
rect 975 -1553 976 -1552
rect 1045 -1553 1046 -1552
rect 1094 -1553 1095 -1552
rect 1115 -1553 1116 -1552
rect 9 -1555 10 -1554
rect 485 -1555 486 -1554
rect 513 -1555 514 -1554
rect 670 -1555 671 -1554
rect 674 -1555 675 -1554
rect 1017 -1555 1018 -1554
rect 1073 -1555 1074 -1554
rect 1094 -1555 1095 -1554
rect 30 -1557 31 -1556
rect 149 -1557 150 -1556
rect 156 -1557 157 -1556
rect 184 -1557 185 -1556
rect 198 -1557 199 -1556
rect 261 -1557 262 -1556
rect 268 -1557 269 -1556
rect 534 -1557 535 -1556
rect 562 -1557 563 -1556
rect 905 -1557 906 -1556
rect 926 -1557 927 -1556
rect 1017 -1557 1018 -1556
rect 33 -1559 34 -1558
rect 40 -1559 41 -1558
rect 51 -1559 52 -1558
rect 460 -1559 461 -1558
rect 471 -1559 472 -1558
rect 751 -1559 752 -1558
rect 821 -1559 822 -1558
rect 891 -1559 892 -1558
rect 989 -1559 990 -1558
rect 1073 -1559 1074 -1558
rect 37 -1561 38 -1560
rect 653 -1561 654 -1560
rect 660 -1561 661 -1560
rect 758 -1561 759 -1560
rect 821 -1561 822 -1560
rect 1069 -1561 1070 -1560
rect 37 -1563 38 -1562
rect 44 -1563 45 -1562
rect 51 -1563 52 -1562
rect 425 -1563 426 -1562
rect 478 -1563 479 -1562
rect 499 -1563 500 -1562
rect 520 -1563 521 -1562
rect 618 -1563 619 -1562
rect 625 -1563 626 -1562
rect 772 -1563 773 -1562
rect 835 -1563 836 -1562
rect 926 -1563 927 -1562
rect 961 -1563 962 -1562
rect 989 -1563 990 -1562
rect 996 -1563 997 -1562
rect 1080 -1563 1081 -1562
rect 65 -1565 66 -1564
rect 499 -1565 500 -1564
rect 534 -1565 535 -1564
rect 898 -1565 899 -1564
rect 16 -1567 17 -1566
rect 65 -1567 66 -1566
rect 72 -1567 73 -1566
rect 520 -1567 521 -1566
rect 565 -1567 566 -1566
rect 1024 -1567 1025 -1566
rect 16 -1569 17 -1568
rect 222 -1569 223 -1568
rect 268 -1569 269 -1568
rect 338 -1569 339 -1568
rect 359 -1569 360 -1568
rect 677 -1569 678 -1568
rect 716 -1569 717 -1568
rect 751 -1569 752 -1568
rect 814 -1569 815 -1568
rect 898 -1569 899 -1568
rect 982 -1569 983 -1568
rect 1024 -1569 1025 -1568
rect 72 -1571 73 -1570
rect 86 -1571 87 -1570
rect 93 -1571 94 -1570
rect 569 -1571 570 -1570
rect 576 -1571 577 -1570
rect 688 -1571 689 -1570
rect 716 -1571 717 -1570
rect 744 -1571 745 -1570
rect 765 -1571 766 -1570
rect 814 -1571 815 -1570
rect 859 -1571 860 -1570
rect 1003 -1571 1004 -1570
rect 79 -1573 80 -1572
rect 149 -1573 150 -1572
rect 163 -1573 164 -1572
rect 471 -1573 472 -1572
rect 478 -1573 479 -1572
rect 674 -1573 675 -1572
rect 684 -1573 685 -1572
rect 744 -1573 745 -1572
rect 765 -1573 766 -1572
rect 863 -1573 864 -1572
rect 870 -1573 871 -1572
rect 919 -1573 920 -1572
rect 933 -1573 934 -1572
rect 1003 -1573 1004 -1572
rect 79 -1575 80 -1574
rect 275 -1575 276 -1574
rect 282 -1575 283 -1574
rect 292 -1575 293 -1574
rect 345 -1575 346 -1574
rect 863 -1575 864 -1574
rect 884 -1575 885 -1574
rect 975 -1575 976 -1574
rect 86 -1577 87 -1576
rect 114 -1577 115 -1576
rect 121 -1577 122 -1576
rect 156 -1577 157 -1576
rect 163 -1577 164 -1576
rect 450 -1577 451 -1576
rect 464 -1577 465 -1576
rect 618 -1577 619 -1576
rect 625 -1577 626 -1576
rect 1038 -1577 1039 -1576
rect 96 -1579 97 -1578
rect 516 -1579 517 -1578
rect 527 -1579 528 -1578
rect 576 -1579 577 -1578
rect 590 -1579 591 -1578
rect 961 -1579 962 -1578
rect 968 -1579 969 -1578
rect 982 -1579 983 -1578
rect 100 -1581 101 -1580
rect 107 -1581 108 -1580
rect 121 -1581 122 -1580
rect 135 -1581 136 -1580
rect 166 -1581 167 -1580
rect 485 -1581 486 -1580
rect 506 -1581 507 -1580
rect 527 -1581 528 -1580
rect 583 -1581 584 -1580
rect 590 -1581 591 -1580
rect 593 -1581 594 -1580
rect 702 -1581 703 -1580
rect 723 -1581 724 -1580
rect 835 -1581 836 -1580
rect 912 -1581 913 -1580
rect 968 -1581 969 -1580
rect 107 -1583 108 -1582
rect 310 -1583 311 -1582
rect 331 -1583 332 -1582
rect 450 -1583 451 -1582
rect 597 -1583 598 -1582
rect 1087 -1583 1088 -1582
rect 128 -1585 129 -1584
rect 145 -1585 146 -1584
rect 177 -1585 178 -1584
rect 401 -1585 402 -1584
rect 597 -1585 598 -1584
rect 604 -1585 605 -1584
rect 611 -1585 612 -1584
rect 677 -1585 678 -1584
rect 723 -1585 724 -1584
rect 730 -1585 731 -1584
rect 793 -1585 794 -1584
rect 870 -1585 871 -1584
rect 114 -1587 115 -1586
rect 611 -1587 612 -1586
rect 614 -1587 615 -1586
rect 940 -1587 941 -1586
rect 128 -1589 129 -1588
rect 352 -1589 353 -1588
rect 366 -1589 367 -1588
rect 401 -1589 402 -1588
rect 429 -1589 430 -1588
rect 604 -1589 605 -1588
rect 632 -1589 633 -1588
rect 905 -1589 906 -1588
rect 180 -1591 181 -1590
rect 422 -1591 423 -1590
rect 457 -1591 458 -1590
rect 793 -1591 794 -1590
rect 800 -1591 801 -1590
rect 933 -1591 934 -1590
rect 201 -1593 202 -1592
rect 681 -1593 682 -1592
rect 730 -1593 731 -1592
rect 849 -1593 850 -1592
rect 205 -1595 206 -1594
rect 208 -1595 209 -1594
rect 212 -1595 213 -1594
rect 229 -1595 230 -1594
rect 233 -1595 234 -1594
rect 506 -1595 507 -1594
rect 635 -1595 636 -1594
rect 702 -1595 703 -1594
rect 800 -1595 801 -1594
rect 1062 -1595 1063 -1594
rect 191 -1597 192 -1596
rect 212 -1597 213 -1596
rect 219 -1597 220 -1596
rect 254 -1597 255 -1596
rect 278 -1597 279 -1596
rect 849 -1597 850 -1596
rect 58 -1599 59 -1598
rect 191 -1599 192 -1598
rect 226 -1599 227 -1598
rect 345 -1599 346 -1598
rect 366 -1599 367 -1598
rect 467 -1599 468 -1598
rect 639 -1599 640 -1598
rect 653 -1599 654 -1598
rect 663 -1599 664 -1598
rect 807 -1599 808 -1598
rect 828 -1599 829 -1598
rect 884 -1599 885 -1598
rect 44 -1601 45 -1600
rect 226 -1601 227 -1600
rect 233 -1601 234 -1600
rect 387 -1601 388 -1600
rect 394 -1601 395 -1600
rect 562 -1601 563 -1600
rect 639 -1601 640 -1600
rect 1031 -1601 1032 -1600
rect 58 -1603 59 -1602
rect 695 -1603 696 -1602
rect 737 -1603 738 -1602
rect 807 -1603 808 -1602
rect 947 -1603 948 -1602
rect 1031 -1603 1032 -1602
rect 240 -1605 241 -1604
rect 331 -1605 332 -1604
rect 355 -1605 356 -1604
rect 394 -1605 395 -1604
rect 408 -1605 409 -1604
rect 429 -1605 430 -1604
rect 646 -1605 647 -1604
rect 912 -1605 913 -1604
rect 947 -1605 948 -1604
rect 954 -1605 955 -1604
rect 240 -1607 241 -1606
rect 317 -1607 318 -1606
rect 324 -1607 325 -1606
rect 632 -1607 633 -1606
rect 667 -1607 668 -1606
rect 779 -1607 780 -1606
rect 877 -1607 878 -1606
rect 954 -1607 955 -1606
rect 282 -1609 283 -1608
rect 586 -1609 587 -1608
rect 709 -1609 710 -1608
rect 877 -1609 878 -1608
rect 303 -1611 304 -1610
rect 317 -1611 318 -1610
rect 373 -1611 374 -1610
rect 387 -1611 388 -1610
rect 408 -1611 409 -1610
rect 415 -1611 416 -1610
rect 492 -1611 493 -1610
rect 646 -1611 647 -1610
rect 737 -1611 738 -1610
rect 786 -1611 787 -1610
rect 23 -1613 24 -1612
rect 492 -1613 493 -1612
rect 523 -1613 524 -1612
rect 709 -1613 710 -1612
rect 758 -1613 759 -1612
rect 779 -1613 780 -1612
rect 786 -1613 787 -1612
rect 856 -1613 857 -1612
rect 23 -1615 24 -1614
rect 296 -1615 297 -1614
rect 310 -1615 311 -1614
rect 327 -1615 328 -1614
rect 338 -1615 339 -1614
rect 373 -1615 374 -1614
rect 415 -1615 416 -1614
rect 569 -1615 570 -1614
rect 775 -1615 776 -1614
rect 828 -1615 829 -1614
rect 856 -1615 857 -1614
rect 996 -1615 997 -1614
rect 296 -1617 297 -1616
rect 380 -1617 381 -1616
rect 537 -1617 538 -1616
rect 667 -1617 668 -1616
rect 380 -1619 381 -1618
rect 443 -1619 444 -1618
rect 443 -1621 444 -1620
rect 541 -1621 542 -1620
rect 541 -1623 542 -1622
rect 555 -1623 556 -1622
rect 548 -1625 549 -1624
rect 555 -1625 556 -1624
rect 82 -1627 83 -1626
rect 548 -1627 549 -1626
rect 9 -1638 10 -1637
rect 341 -1638 342 -1637
rect 355 -1638 356 -1637
rect 604 -1638 605 -1637
rect 607 -1638 608 -1637
rect 926 -1638 927 -1637
rect 1059 -1638 1060 -1637
rect 1108 -1638 1109 -1637
rect 23 -1640 24 -1639
rect 26 -1640 27 -1639
rect 37 -1640 38 -1639
rect 40 -1640 41 -1639
rect 58 -1640 59 -1639
rect 695 -1640 696 -1639
rect 779 -1640 780 -1639
rect 884 -1640 885 -1639
rect 1066 -1640 1067 -1639
rect 1094 -1640 1095 -1639
rect 23 -1642 24 -1641
rect 142 -1642 143 -1641
rect 149 -1642 150 -1641
rect 306 -1642 307 -1641
rect 313 -1642 314 -1641
rect 485 -1642 486 -1641
rect 523 -1642 524 -1641
rect 660 -1642 661 -1641
rect 674 -1642 675 -1641
rect 989 -1642 990 -1641
rect 1069 -1642 1070 -1641
rect 1115 -1642 1116 -1641
rect 37 -1644 38 -1643
rect 198 -1644 199 -1643
rect 222 -1644 223 -1643
rect 520 -1644 521 -1643
rect 534 -1644 535 -1643
rect 576 -1644 577 -1643
rect 583 -1644 584 -1643
rect 947 -1644 948 -1643
rect 1094 -1644 1095 -1643
rect 1101 -1644 1102 -1643
rect 58 -1646 59 -1645
rect 100 -1646 101 -1645
rect 114 -1646 115 -1645
rect 198 -1646 199 -1645
rect 247 -1646 248 -1645
rect 324 -1646 325 -1645
rect 376 -1646 377 -1645
rect 828 -1646 829 -1645
rect 835 -1646 836 -1645
rect 884 -1646 885 -1645
rect 947 -1646 948 -1645
rect 1073 -1646 1074 -1645
rect 51 -1648 52 -1647
rect 114 -1648 115 -1647
rect 135 -1648 136 -1647
rect 443 -1648 444 -1647
rect 450 -1648 451 -1647
rect 485 -1648 486 -1647
rect 572 -1648 573 -1647
rect 912 -1648 913 -1647
rect 16 -1650 17 -1649
rect 135 -1650 136 -1649
rect 138 -1650 139 -1649
rect 331 -1650 332 -1649
rect 383 -1650 384 -1649
rect 761 -1650 762 -1649
rect 786 -1650 787 -1649
rect 828 -1650 829 -1649
rect 912 -1650 913 -1649
rect 996 -1650 997 -1649
rect 61 -1652 62 -1651
rect 663 -1652 664 -1651
rect 684 -1652 685 -1651
rect 891 -1652 892 -1651
rect 65 -1654 66 -1653
rect 100 -1654 101 -1653
rect 142 -1654 143 -1653
rect 177 -1654 178 -1653
rect 187 -1654 188 -1653
rect 506 -1654 507 -1653
rect 586 -1654 587 -1653
rect 1087 -1654 1088 -1653
rect 40 -1656 41 -1655
rect 51 -1656 52 -1655
rect 79 -1656 80 -1655
rect 380 -1656 381 -1655
rect 394 -1656 395 -1655
rect 446 -1656 447 -1655
rect 450 -1656 451 -1655
rect 590 -1656 591 -1655
rect 611 -1656 612 -1655
rect 656 -1656 657 -1655
rect 691 -1656 692 -1655
rect 716 -1656 717 -1655
rect 730 -1656 731 -1655
rect 835 -1656 836 -1655
rect 891 -1656 892 -1655
rect 1010 -1656 1011 -1655
rect 82 -1658 83 -1657
rect 436 -1658 437 -1657
rect 460 -1658 461 -1657
rect 821 -1658 822 -1657
rect 93 -1660 94 -1659
rect 128 -1660 129 -1659
rect 149 -1660 150 -1659
rect 226 -1660 227 -1659
rect 254 -1660 255 -1659
rect 331 -1660 332 -1659
rect 380 -1660 381 -1659
rect 758 -1660 759 -1659
rect 786 -1660 787 -1659
rect 870 -1660 871 -1659
rect 54 -1662 55 -1661
rect 128 -1662 129 -1661
rect 159 -1662 160 -1661
rect 457 -1662 458 -1661
rect 506 -1662 507 -1661
rect 541 -1662 542 -1661
rect 590 -1662 591 -1661
rect 597 -1662 598 -1661
rect 614 -1662 615 -1661
rect 898 -1662 899 -1661
rect 96 -1664 97 -1663
rect 107 -1664 108 -1663
rect 170 -1664 171 -1663
rect 362 -1664 363 -1663
rect 401 -1664 402 -1663
rect 625 -1664 626 -1663
rect 639 -1664 640 -1663
rect 660 -1664 661 -1663
rect 667 -1664 668 -1663
rect 758 -1664 759 -1663
rect 765 -1664 766 -1663
rect 870 -1664 871 -1663
rect 898 -1664 899 -1663
rect 961 -1664 962 -1663
rect 72 -1666 73 -1665
rect 107 -1666 108 -1665
rect 156 -1666 157 -1665
rect 170 -1666 171 -1665
rect 191 -1666 192 -1665
rect 863 -1666 864 -1665
rect 961 -1666 962 -1665
rect 982 -1666 983 -1665
rect 72 -1668 73 -1667
rect 86 -1668 87 -1667
rect 191 -1668 192 -1667
rect 205 -1668 206 -1667
rect 226 -1668 227 -1667
rect 240 -1668 241 -1667
rect 254 -1668 255 -1667
rect 261 -1668 262 -1667
rect 296 -1668 297 -1667
rect 327 -1668 328 -1667
rect 387 -1668 388 -1667
rect 401 -1668 402 -1667
rect 422 -1668 423 -1667
rect 674 -1668 675 -1667
rect 681 -1668 682 -1667
rect 765 -1668 766 -1667
rect 821 -1668 822 -1667
rect 919 -1668 920 -1667
rect 86 -1670 87 -1669
rect 212 -1670 213 -1669
rect 240 -1670 241 -1669
rect 366 -1670 367 -1669
rect 387 -1670 388 -1669
rect 569 -1670 570 -1669
rect 597 -1670 598 -1669
rect 653 -1670 654 -1669
rect 695 -1670 696 -1669
rect 751 -1670 752 -1669
rect 842 -1670 843 -1669
rect 863 -1670 864 -1669
rect 919 -1670 920 -1669
rect 1031 -1670 1032 -1669
rect 65 -1672 66 -1671
rect 653 -1672 654 -1671
rect 702 -1672 703 -1671
rect 779 -1672 780 -1671
rect 842 -1672 843 -1671
rect 954 -1672 955 -1671
rect 163 -1674 164 -1673
rect 261 -1674 262 -1673
rect 296 -1674 297 -1673
rect 310 -1674 311 -1673
rect 317 -1674 318 -1673
rect 355 -1674 356 -1673
rect 366 -1674 367 -1673
rect 492 -1674 493 -1673
rect 618 -1674 619 -1673
rect 1062 -1674 1063 -1673
rect 163 -1676 164 -1675
rect 376 -1676 377 -1675
rect 422 -1676 423 -1675
rect 537 -1676 538 -1675
rect 618 -1676 619 -1675
rect 688 -1676 689 -1675
rect 702 -1676 703 -1675
rect 807 -1676 808 -1675
rect 954 -1676 955 -1675
rect 1080 -1676 1081 -1675
rect 201 -1678 202 -1677
rect 394 -1678 395 -1677
rect 425 -1678 426 -1677
rect 905 -1678 906 -1677
rect 205 -1680 206 -1679
rect 289 -1680 290 -1679
rect 317 -1680 318 -1679
rect 359 -1680 360 -1679
rect 429 -1680 430 -1679
rect 436 -1680 437 -1679
rect 457 -1680 458 -1679
rect 464 -1680 465 -1679
rect 471 -1680 472 -1679
rect 667 -1680 668 -1679
rect 716 -1680 717 -1679
rect 793 -1680 794 -1679
rect 807 -1680 808 -1679
rect 975 -1680 976 -1679
rect 212 -1682 213 -1681
rect 415 -1682 416 -1681
rect 464 -1682 465 -1681
rect 513 -1682 514 -1681
rect 625 -1682 626 -1681
rect 709 -1682 710 -1681
rect 730 -1682 731 -1681
rect 933 -1682 934 -1681
rect 233 -1684 234 -1683
rect 310 -1684 311 -1683
rect 327 -1684 328 -1683
rect 849 -1684 850 -1683
rect 905 -1684 906 -1683
rect 940 -1684 941 -1683
rect 184 -1686 185 -1685
rect 849 -1686 850 -1685
rect 933 -1686 934 -1685
rect 1045 -1686 1046 -1685
rect 44 -1688 45 -1687
rect 184 -1688 185 -1687
rect 233 -1688 234 -1687
rect 338 -1688 339 -1687
rect 359 -1688 360 -1687
rect 569 -1688 570 -1687
rect 632 -1688 633 -1687
rect 681 -1688 682 -1687
rect 709 -1688 710 -1687
rect 737 -1688 738 -1687
rect 744 -1688 745 -1687
rect 793 -1688 794 -1687
rect 940 -1688 941 -1687
rect 1038 -1688 1039 -1687
rect 44 -1690 45 -1689
rect 68 -1690 69 -1689
rect 268 -1690 269 -1689
rect 289 -1690 290 -1689
rect 373 -1690 374 -1689
rect 429 -1690 430 -1689
rect 471 -1690 472 -1689
rect 499 -1690 500 -1689
rect 513 -1690 514 -1689
rect 562 -1690 563 -1689
rect 639 -1690 640 -1689
rect 646 -1690 647 -1689
rect 737 -1690 738 -1689
rect 877 -1690 878 -1689
rect 268 -1692 269 -1691
rect 275 -1692 276 -1691
rect 373 -1692 374 -1691
rect 772 -1692 773 -1691
rect 877 -1692 878 -1691
rect 1052 -1692 1053 -1691
rect 415 -1694 416 -1693
rect 527 -1694 528 -1693
rect 646 -1694 647 -1693
rect 677 -1694 678 -1693
rect 723 -1694 724 -1693
rect 772 -1694 773 -1693
rect 408 -1696 409 -1695
rect 527 -1696 528 -1695
rect 723 -1696 724 -1695
rect 814 -1696 815 -1695
rect 408 -1698 409 -1697
rect 579 -1698 580 -1697
rect 744 -1698 745 -1697
rect 800 -1698 801 -1697
rect 478 -1700 479 -1699
rect 541 -1700 542 -1699
rect 751 -1700 752 -1699
rect 1024 -1700 1025 -1699
rect 30 -1702 31 -1701
rect 478 -1702 479 -1701
rect 481 -1702 482 -1701
rect 562 -1702 563 -1701
rect 800 -1702 801 -1701
rect 968 -1702 969 -1701
rect 30 -1704 31 -1703
rect 121 -1704 122 -1703
rect 488 -1704 489 -1703
rect 632 -1704 633 -1703
rect 968 -1704 969 -1703
rect 1003 -1704 1004 -1703
rect 121 -1706 122 -1705
rect 282 -1706 283 -1705
rect 499 -1706 500 -1705
rect 548 -1706 549 -1705
rect 282 -1708 283 -1707
rect 303 -1708 304 -1707
rect 548 -1708 549 -1707
rect 555 -1708 556 -1707
rect 275 -1710 276 -1709
rect 303 -1710 304 -1709
rect 555 -1710 556 -1709
rect 856 -1710 857 -1709
rect 856 -1712 857 -1711
rect 1017 -1712 1018 -1711
rect 2 -1723 3 -1722
rect 212 -1723 213 -1722
rect 254 -1723 255 -1722
rect 324 -1723 325 -1722
rect 338 -1723 339 -1722
rect 607 -1723 608 -1722
rect 653 -1723 654 -1722
rect 828 -1723 829 -1722
rect 849 -1723 850 -1722
rect 1017 -1723 1018 -1722
rect 1052 -1723 1053 -1722
rect 1069 -1723 1070 -1722
rect 16 -1725 17 -1724
rect 37 -1725 38 -1724
rect 51 -1725 52 -1724
rect 93 -1725 94 -1724
rect 100 -1725 101 -1724
rect 138 -1725 139 -1724
rect 159 -1725 160 -1724
rect 240 -1725 241 -1724
rect 261 -1725 262 -1724
rect 849 -1725 850 -1724
rect 870 -1725 871 -1724
rect 908 -1725 909 -1724
rect 919 -1725 920 -1724
rect 996 -1725 997 -1724
rect 1055 -1725 1056 -1724
rect 1087 -1725 1088 -1724
rect 30 -1727 31 -1726
rect 222 -1727 223 -1726
rect 226 -1727 227 -1726
rect 261 -1727 262 -1726
rect 275 -1727 276 -1726
rect 324 -1727 325 -1726
rect 359 -1727 360 -1726
rect 520 -1727 521 -1726
rect 527 -1727 528 -1726
rect 730 -1727 731 -1726
rect 758 -1727 759 -1726
rect 807 -1727 808 -1726
rect 817 -1727 818 -1726
rect 933 -1727 934 -1726
rect 940 -1727 941 -1726
rect 982 -1727 983 -1726
rect 23 -1729 24 -1728
rect 222 -1729 223 -1728
rect 233 -1729 234 -1728
rect 254 -1729 255 -1728
rect 275 -1729 276 -1728
rect 282 -1729 283 -1728
rect 296 -1729 297 -1728
rect 303 -1729 304 -1728
rect 366 -1729 367 -1728
rect 432 -1729 433 -1728
rect 436 -1729 437 -1728
rect 523 -1729 524 -1728
rect 527 -1729 528 -1728
rect 597 -1729 598 -1728
rect 632 -1729 633 -1728
rect 919 -1729 920 -1728
rect 926 -1729 927 -1728
rect 961 -1729 962 -1728
rect 30 -1731 31 -1730
rect 677 -1731 678 -1730
rect 681 -1731 682 -1730
rect 814 -1731 815 -1730
rect 828 -1731 829 -1730
rect 863 -1731 864 -1730
rect 877 -1731 878 -1730
rect 1003 -1731 1004 -1730
rect 37 -1733 38 -1732
rect 44 -1733 45 -1732
rect 65 -1733 66 -1732
rect 457 -1733 458 -1732
rect 478 -1733 479 -1732
rect 751 -1733 752 -1732
rect 761 -1733 762 -1732
rect 1045 -1733 1046 -1732
rect 44 -1735 45 -1734
rect 121 -1735 122 -1734
rect 212 -1735 213 -1734
rect 317 -1735 318 -1734
rect 366 -1735 367 -1734
rect 380 -1735 381 -1734
rect 408 -1735 409 -1734
rect 653 -1735 654 -1734
rect 660 -1735 661 -1734
rect 989 -1735 990 -1734
rect 65 -1737 66 -1736
rect 205 -1737 206 -1736
rect 219 -1737 220 -1736
rect 317 -1737 318 -1736
rect 380 -1737 381 -1736
rect 464 -1737 465 -1736
rect 495 -1737 496 -1736
rect 499 -1737 500 -1736
rect 534 -1737 535 -1736
rect 660 -1737 661 -1736
rect 674 -1737 675 -1736
rect 856 -1737 857 -1736
rect 863 -1737 864 -1736
rect 912 -1737 913 -1736
rect 926 -1737 927 -1736
rect 947 -1737 948 -1736
rect 954 -1737 955 -1736
rect 1024 -1737 1025 -1736
rect 79 -1739 80 -1738
rect 383 -1739 384 -1738
rect 408 -1739 409 -1738
rect 502 -1739 503 -1738
rect 506 -1739 507 -1738
rect 534 -1739 535 -1738
rect 586 -1739 587 -1738
rect 751 -1739 752 -1738
rect 793 -1739 794 -1738
rect 912 -1739 913 -1738
rect 929 -1739 930 -1738
rect 961 -1739 962 -1738
rect 79 -1741 80 -1740
rect 355 -1741 356 -1740
rect 425 -1741 426 -1740
rect 632 -1741 633 -1740
rect 667 -1741 668 -1740
rect 856 -1741 857 -1740
rect 891 -1741 892 -1740
rect 940 -1741 941 -1740
rect 947 -1741 948 -1740
rect 968 -1741 969 -1740
rect 86 -1743 87 -1742
rect 373 -1743 374 -1742
rect 443 -1743 444 -1742
rect 1031 -1743 1032 -1742
rect 86 -1745 87 -1744
rect 107 -1745 108 -1744
rect 121 -1745 122 -1744
rect 376 -1745 377 -1744
rect 443 -1745 444 -1744
rect 579 -1745 580 -1744
rect 597 -1745 598 -1744
rect 625 -1745 626 -1744
rect 667 -1745 668 -1744
rect 772 -1745 773 -1744
rect 842 -1745 843 -1744
rect 877 -1745 878 -1744
rect 891 -1745 892 -1744
rect 898 -1745 899 -1744
rect 905 -1745 906 -1744
rect 1038 -1745 1039 -1744
rect 100 -1747 101 -1746
rect 289 -1747 290 -1746
rect 296 -1747 297 -1746
rect 418 -1747 419 -1746
rect 450 -1747 451 -1746
rect 583 -1747 584 -1746
rect 670 -1747 671 -1746
rect 898 -1747 899 -1746
rect 107 -1749 108 -1748
rect 142 -1749 143 -1748
rect 156 -1749 157 -1748
rect 674 -1749 675 -1748
rect 681 -1749 682 -1748
rect 709 -1749 710 -1748
rect 716 -1749 717 -1748
rect 1059 -1749 1060 -1748
rect 135 -1751 136 -1750
rect 793 -1751 794 -1750
rect 800 -1751 801 -1750
rect 905 -1751 906 -1750
rect 23 -1753 24 -1752
rect 135 -1753 136 -1752
rect 142 -1753 143 -1752
rect 191 -1753 192 -1752
rect 198 -1753 199 -1752
rect 499 -1753 500 -1752
rect 506 -1753 507 -1752
rect 646 -1753 647 -1752
rect 688 -1753 689 -1752
rect 786 -1753 787 -1752
rect 156 -1755 157 -1754
rect 387 -1755 388 -1754
rect 450 -1755 451 -1754
rect 520 -1755 521 -1754
rect 569 -1755 570 -1754
rect 646 -1755 647 -1754
rect 688 -1755 689 -1754
rect 821 -1755 822 -1754
rect 163 -1757 164 -1756
rect 716 -1757 717 -1756
rect 723 -1757 724 -1756
rect 821 -1757 822 -1756
rect 149 -1759 150 -1758
rect 723 -1759 724 -1758
rect 730 -1759 731 -1758
rect 835 -1759 836 -1758
rect 149 -1761 150 -1760
rect 345 -1761 346 -1760
rect 348 -1761 349 -1760
rect 786 -1761 787 -1760
rect 163 -1763 164 -1762
rect 184 -1763 185 -1762
rect 191 -1763 192 -1762
rect 691 -1763 692 -1762
rect 702 -1763 703 -1762
rect 870 -1763 871 -1762
rect 114 -1765 115 -1764
rect 184 -1765 185 -1764
rect 198 -1765 199 -1764
rect 1010 -1765 1011 -1764
rect 226 -1767 227 -1766
rect 425 -1767 426 -1766
rect 457 -1767 458 -1766
rect 611 -1767 612 -1766
rect 625 -1767 626 -1766
rect 800 -1767 801 -1766
rect 233 -1769 234 -1768
rect 310 -1769 311 -1768
rect 373 -1769 374 -1768
rect 488 -1769 489 -1768
rect 576 -1769 577 -1768
rect 968 -1769 969 -1768
rect 128 -1771 129 -1770
rect 310 -1771 311 -1770
rect 387 -1771 388 -1770
rect 429 -1771 430 -1770
rect 464 -1771 465 -1770
rect 513 -1771 514 -1770
rect 611 -1771 612 -1770
rect 975 -1771 976 -1770
rect 128 -1773 129 -1772
rect 247 -1773 248 -1772
rect 268 -1773 269 -1772
rect 303 -1773 304 -1772
rect 306 -1773 307 -1772
rect 436 -1773 437 -1772
rect 485 -1773 486 -1772
rect 576 -1773 577 -1772
rect 639 -1773 640 -1772
rect 702 -1773 703 -1772
rect 737 -1773 738 -1772
rect 772 -1773 773 -1772
rect 240 -1775 241 -1774
rect 530 -1775 531 -1774
rect 618 -1775 619 -1774
rect 639 -1775 640 -1774
rect 695 -1775 696 -1774
rect 737 -1775 738 -1774
rect 744 -1775 745 -1774
rect 807 -1775 808 -1774
rect 268 -1777 269 -1776
rect 331 -1777 332 -1776
rect 352 -1777 353 -1776
rect 485 -1777 486 -1776
rect 492 -1777 493 -1776
rect 744 -1777 745 -1776
rect 765 -1777 766 -1776
rect 835 -1777 836 -1776
rect 58 -1779 59 -1778
rect 331 -1779 332 -1778
rect 352 -1779 353 -1778
rect 569 -1779 570 -1778
rect 600 -1779 601 -1778
rect 695 -1779 696 -1778
rect 712 -1779 713 -1778
rect 765 -1779 766 -1778
rect 58 -1781 59 -1780
rect 72 -1781 73 -1780
rect 282 -1781 283 -1780
rect 401 -1781 402 -1780
rect 415 -1781 416 -1780
rect 492 -1781 493 -1780
rect 72 -1783 73 -1782
rect 247 -1783 248 -1782
rect 289 -1783 290 -1782
rect 341 -1783 342 -1782
rect 362 -1783 363 -1782
rect 618 -1783 619 -1782
rect 394 -1785 395 -1784
rect 513 -1785 514 -1784
rect 394 -1787 395 -1786
rect 530 -1787 531 -1786
rect 401 -1789 402 -1788
rect 555 -1789 556 -1788
rect 415 -1791 416 -1790
rect 471 -1791 472 -1790
rect 555 -1791 556 -1790
rect 590 -1791 591 -1790
rect 429 -1793 430 -1792
rect 954 -1793 955 -1792
rect 471 -1795 472 -1794
rect 562 -1795 563 -1794
rect 590 -1795 591 -1794
rect 604 -1795 605 -1794
rect 541 -1797 542 -1796
rect 562 -1797 563 -1796
rect 604 -1797 605 -1796
rect 842 -1797 843 -1796
rect 541 -1799 542 -1798
rect 548 -1799 549 -1798
rect 548 -1801 549 -1800
rect 884 -1801 885 -1800
rect 117 -1803 118 -1802
rect 884 -1803 885 -1802
rect 2 -1814 3 -1813
rect 425 -1814 426 -1813
rect 443 -1814 444 -1813
rect 453 -1814 454 -1813
rect 499 -1814 500 -1813
rect 870 -1814 871 -1813
rect 933 -1814 934 -1813
rect 947 -1814 948 -1813
rect 1010 -1814 1011 -1813
rect 1052 -1814 1053 -1813
rect 1087 -1814 1088 -1813
rect 1101 -1814 1102 -1813
rect 5 -1816 6 -1815
rect 527 -1816 528 -1815
rect 604 -1816 605 -1815
rect 702 -1816 703 -1815
rect 709 -1816 710 -1815
rect 996 -1816 997 -1815
rect 1017 -1816 1018 -1815
rect 1073 -1816 1074 -1815
rect 1087 -1816 1088 -1815
rect 1094 -1816 1095 -1815
rect 37 -1818 38 -1817
rect 40 -1818 41 -1817
rect 54 -1818 55 -1817
rect 72 -1818 73 -1817
rect 79 -1818 80 -1817
rect 432 -1818 433 -1817
rect 443 -1818 444 -1817
rect 492 -1818 493 -1817
rect 502 -1818 503 -1817
rect 653 -1818 654 -1817
rect 667 -1818 668 -1817
rect 758 -1818 759 -1817
rect 912 -1818 913 -1817
rect 933 -1818 934 -1817
rect 975 -1818 976 -1817
rect 996 -1818 997 -1817
rect 1045 -1818 1046 -1817
rect 1055 -1818 1056 -1817
rect 47 -1820 48 -1819
rect 72 -1820 73 -1819
rect 93 -1820 94 -1819
rect 849 -1820 850 -1819
rect 891 -1820 892 -1819
rect 912 -1820 913 -1819
rect 926 -1820 927 -1819
rect 1017 -1820 1018 -1819
rect 103 -1822 104 -1821
rect 373 -1822 374 -1821
rect 387 -1822 388 -1821
rect 635 -1822 636 -1821
rect 646 -1822 647 -1821
rect 870 -1822 871 -1821
rect 891 -1822 892 -1821
rect 940 -1822 941 -1821
rect 954 -1822 955 -1821
rect 975 -1822 976 -1821
rect 114 -1824 115 -1823
rect 261 -1824 262 -1823
rect 268 -1824 269 -1823
rect 362 -1824 363 -1823
rect 373 -1824 374 -1823
rect 712 -1824 713 -1823
rect 733 -1824 734 -1823
rect 905 -1824 906 -1823
rect 919 -1824 920 -1823
rect 940 -1824 941 -1823
rect 93 -1826 94 -1825
rect 114 -1826 115 -1825
rect 121 -1826 122 -1825
rect 184 -1826 185 -1825
rect 198 -1826 199 -1825
rect 793 -1826 794 -1825
rect 863 -1826 864 -1825
rect 926 -1826 927 -1825
rect 121 -1828 122 -1827
rect 583 -1828 584 -1827
rect 590 -1828 591 -1827
rect 646 -1828 647 -1827
rect 688 -1828 689 -1827
rect 1069 -1828 1070 -1827
rect 124 -1830 125 -1829
rect 219 -1830 220 -1829
rect 226 -1830 227 -1829
rect 418 -1830 419 -1829
rect 429 -1830 430 -1829
rect 947 -1830 948 -1829
rect 135 -1832 136 -1831
rect 1010 -1832 1011 -1831
rect 135 -1834 136 -1833
rect 191 -1834 192 -1833
rect 194 -1834 195 -1833
rect 590 -1834 591 -1833
rect 614 -1834 615 -1833
rect 821 -1834 822 -1833
rect 877 -1834 878 -1833
rect 905 -1834 906 -1833
rect 163 -1836 164 -1835
rect 352 -1836 353 -1835
rect 366 -1836 367 -1835
rect 877 -1836 878 -1835
rect 884 -1836 885 -1835
rect 919 -1836 920 -1835
rect 163 -1838 164 -1837
rect 551 -1838 552 -1837
rect 569 -1838 570 -1837
rect 709 -1838 710 -1837
rect 737 -1838 738 -1837
rect 849 -1838 850 -1837
rect 898 -1838 899 -1837
rect 954 -1838 955 -1837
rect 198 -1840 199 -1839
rect 359 -1840 360 -1839
rect 394 -1840 395 -1839
rect 604 -1840 605 -1839
rect 628 -1840 629 -1839
rect 681 -1840 682 -1839
rect 695 -1840 696 -1839
rect 702 -1840 703 -1839
rect 723 -1840 724 -1839
rect 737 -1840 738 -1839
rect 751 -1840 752 -1839
rect 758 -1840 759 -1839
rect 765 -1840 766 -1839
rect 898 -1840 899 -1839
rect 201 -1842 202 -1841
rect 268 -1842 269 -1841
rect 282 -1842 283 -1841
rect 387 -1842 388 -1841
rect 415 -1842 416 -1841
rect 751 -1842 752 -1841
rect 772 -1842 773 -1841
rect 863 -1842 864 -1841
rect 208 -1844 209 -1843
rect 233 -1844 234 -1843
rect 250 -1844 251 -1843
rect 618 -1844 619 -1843
rect 695 -1844 696 -1843
rect 716 -1844 717 -1843
rect 723 -1844 724 -1843
rect 800 -1844 801 -1843
rect 814 -1844 815 -1843
rect 821 -1844 822 -1843
rect 842 -1844 843 -1843
rect 884 -1844 885 -1843
rect 226 -1846 227 -1845
rect 558 -1846 559 -1845
rect 576 -1846 577 -1845
rect 793 -1846 794 -1845
rect 800 -1846 801 -1845
rect 807 -1846 808 -1845
rect 814 -1846 815 -1845
rect 1059 -1846 1060 -1845
rect 233 -1848 234 -1847
rect 471 -1848 472 -1847
rect 481 -1848 482 -1847
rect 716 -1848 717 -1847
rect 730 -1848 731 -1847
rect 772 -1848 773 -1847
rect 786 -1848 787 -1847
rect 842 -1848 843 -1847
rect 1031 -1848 1032 -1847
rect 1059 -1848 1060 -1847
rect 254 -1850 255 -1849
rect 359 -1850 360 -1849
rect 366 -1850 367 -1849
rect 576 -1850 577 -1849
rect 583 -1850 584 -1849
rect 625 -1850 626 -1849
rect 691 -1850 692 -1849
rect 807 -1850 808 -1849
rect 989 -1850 990 -1849
rect 1031 -1850 1032 -1849
rect 100 -1852 101 -1851
rect 254 -1852 255 -1851
rect 261 -1852 262 -1851
rect 436 -1852 437 -1851
rect 457 -1852 458 -1851
rect 681 -1852 682 -1851
rect 744 -1852 745 -1851
rect 765 -1852 766 -1851
rect 779 -1852 780 -1851
rect 786 -1852 787 -1851
rect 961 -1852 962 -1851
rect 989 -1852 990 -1851
rect 100 -1854 101 -1853
rect 205 -1854 206 -1853
rect 282 -1854 283 -1853
rect 408 -1854 409 -1853
rect 418 -1854 419 -1853
rect 429 -1854 430 -1853
rect 436 -1854 437 -1853
rect 670 -1854 671 -1853
rect 835 -1854 836 -1853
rect 961 -1854 962 -1853
rect 149 -1856 150 -1855
rect 457 -1856 458 -1855
rect 485 -1856 486 -1855
rect 653 -1856 654 -1855
rect 23 -1858 24 -1857
rect 485 -1858 486 -1857
rect 488 -1858 489 -1857
rect 744 -1858 745 -1857
rect 23 -1860 24 -1859
rect 310 -1860 311 -1859
rect 317 -1860 318 -1859
rect 345 -1860 346 -1859
rect 352 -1860 353 -1859
rect 464 -1860 465 -1859
rect 492 -1860 493 -1859
rect 506 -1860 507 -1859
rect 520 -1860 521 -1859
rect 856 -1860 857 -1859
rect 65 -1862 66 -1861
rect 310 -1862 311 -1861
rect 317 -1862 318 -1861
rect 355 -1862 356 -1861
rect 394 -1862 395 -1861
rect 670 -1862 671 -1861
rect 65 -1864 66 -1863
rect 82 -1864 83 -1863
rect 205 -1864 206 -1863
rect 240 -1864 241 -1863
rect 296 -1864 297 -1863
rect 523 -1864 524 -1863
rect 562 -1864 563 -1863
rect 625 -1864 626 -1863
rect 632 -1864 633 -1863
rect 856 -1864 857 -1863
rect 79 -1866 80 -1865
rect 520 -1866 521 -1865
rect 534 -1866 535 -1865
rect 562 -1866 563 -1865
rect 569 -1866 570 -1865
rect 730 -1866 731 -1865
rect 117 -1868 118 -1867
rect 240 -1868 241 -1867
rect 303 -1868 304 -1867
rect 380 -1868 381 -1867
rect 408 -1868 409 -1867
rect 446 -1868 447 -1867
rect 450 -1868 451 -1867
rect 464 -1868 465 -1867
rect 621 -1868 622 -1867
rect 835 -1868 836 -1867
rect 117 -1870 118 -1869
rect 338 -1870 339 -1869
rect 450 -1870 451 -1869
rect 597 -1870 598 -1869
rect 632 -1870 633 -1869
rect 1038 -1870 1039 -1869
rect 16 -1872 17 -1871
rect 338 -1872 339 -1871
rect 453 -1872 454 -1871
rect 506 -1872 507 -1871
rect 639 -1872 640 -1871
rect 779 -1872 780 -1871
rect 1003 -1872 1004 -1871
rect 1038 -1872 1039 -1871
rect 128 -1874 129 -1873
rect 296 -1874 297 -1873
rect 306 -1874 307 -1873
rect 674 -1874 675 -1873
rect 982 -1874 983 -1873
rect 1003 -1874 1004 -1873
rect 86 -1876 87 -1875
rect 128 -1876 129 -1875
rect 177 -1876 178 -1875
rect 534 -1876 535 -1875
rect 548 -1876 549 -1875
rect 674 -1876 675 -1875
rect 86 -1878 87 -1877
rect 247 -1878 248 -1877
rect 289 -1878 290 -1877
rect 380 -1878 381 -1877
rect 422 -1878 423 -1877
rect 982 -1878 983 -1877
rect 9 -1880 10 -1879
rect 422 -1880 423 -1879
rect 513 -1880 514 -1879
rect 639 -1880 640 -1879
rect 9 -1882 10 -1881
rect 16 -1882 17 -1881
rect 142 -1882 143 -1881
rect 177 -1882 178 -1881
rect 212 -1882 213 -1881
rect 247 -1882 248 -1881
rect 275 -1882 276 -1881
rect 289 -1882 290 -1881
rect 324 -1882 325 -1881
rect 369 -1882 370 -1881
rect 513 -1882 514 -1881
rect 541 -1882 542 -1881
rect 96 -1884 97 -1883
rect 142 -1884 143 -1883
rect 156 -1884 157 -1883
rect 324 -1884 325 -1883
rect 331 -1884 332 -1883
rect 471 -1884 472 -1883
rect 30 -1886 31 -1885
rect 156 -1886 157 -1885
rect 170 -1886 171 -1885
rect 212 -1886 213 -1885
rect 331 -1886 332 -1885
rect 478 -1886 479 -1885
rect 30 -1888 31 -1887
rect 44 -1888 45 -1887
rect 107 -1888 108 -1887
rect 275 -1888 276 -1887
rect 390 -1888 391 -1887
rect 541 -1888 542 -1887
rect 44 -1890 45 -1889
rect 1045 -1890 1046 -1889
rect 51 -1892 52 -1891
rect 107 -1892 108 -1891
rect 170 -1892 171 -1891
rect 348 -1892 349 -1891
rect 478 -1892 479 -1891
rect 660 -1892 661 -1891
rect 51 -1894 52 -1893
rect 68 -1894 69 -1893
rect 551 -1894 552 -1893
rect 660 -1894 661 -1893
rect 2 -1905 3 -1904
rect 527 -1905 528 -1904
rect 530 -1905 531 -1904
rect 1031 -1905 1032 -1904
rect 1073 -1905 1074 -1904
rect 1108 -1905 1109 -1904
rect 9 -1907 10 -1906
rect 40 -1907 41 -1906
rect 44 -1907 45 -1906
rect 128 -1907 129 -1906
rect 142 -1907 143 -1906
rect 191 -1907 192 -1906
rect 194 -1907 195 -1906
rect 492 -1907 493 -1906
rect 502 -1907 503 -1906
rect 534 -1907 535 -1906
rect 551 -1907 552 -1906
rect 849 -1907 850 -1906
rect 1003 -1907 1004 -1906
rect 1031 -1907 1032 -1906
rect 1045 -1907 1046 -1906
rect 1073 -1907 1074 -1906
rect 1080 -1907 1081 -1906
rect 1087 -1907 1088 -1906
rect 1101 -1907 1102 -1906
rect 1115 -1907 1116 -1906
rect 9 -1909 10 -1908
rect 100 -1909 101 -1908
rect 114 -1909 115 -1908
rect 135 -1909 136 -1908
rect 149 -1909 150 -1908
rect 268 -1909 269 -1908
rect 296 -1909 297 -1908
rect 366 -1909 367 -1908
rect 369 -1909 370 -1908
rect 702 -1909 703 -1908
rect 821 -1909 822 -1908
rect 824 -1909 825 -1908
rect 842 -1909 843 -1908
rect 1066 -1909 1067 -1908
rect 16 -1911 17 -1910
rect 481 -1911 482 -1910
rect 485 -1911 486 -1910
rect 695 -1911 696 -1910
rect 702 -1911 703 -1910
rect 1097 -1911 1098 -1910
rect 19 -1913 20 -1912
rect 422 -1913 423 -1912
rect 443 -1913 444 -1912
rect 604 -1913 605 -1912
rect 618 -1913 619 -1912
rect 919 -1913 920 -1912
rect 968 -1913 969 -1912
rect 1003 -1913 1004 -1912
rect 1024 -1913 1025 -1912
rect 1087 -1913 1088 -1912
rect 33 -1915 34 -1914
rect 1045 -1915 1046 -1914
rect 37 -1917 38 -1916
rect 394 -1917 395 -1916
rect 450 -1917 451 -1916
rect 457 -1917 458 -1916
rect 471 -1917 472 -1916
rect 492 -1917 493 -1916
rect 516 -1917 517 -1916
rect 870 -1917 871 -1916
rect 968 -1917 969 -1916
rect 996 -1917 997 -1916
rect 47 -1919 48 -1918
rect 975 -1919 976 -1918
rect 51 -1921 52 -1920
rect 58 -1921 59 -1920
rect 65 -1921 66 -1920
rect 72 -1921 73 -1920
rect 75 -1921 76 -1920
rect 499 -1921 500 -1920
rect 527 -1921 528 -1920
rect 1038 -1921 1039 -1920
rect 58 -1923 59 -1922
rect 394 -1923 395 -1922
rect 453 -1923 454 -1922
rect 1066 -1923 1067 -1922
rect 82 -1925 83 -1924
rect 247 -1925 248 -1924
rect 324 -1925 325 -1924
rect 604 -1925 605 -1924
rect 618 -1925 619 -1924
rect 856 -1925 857 -1924
rect 870 -1925 871 -1924
rect 933 -1925 934 -1924
rect 947 -1925 948 -1924
rect 975 -1925 976 -1924
rect 93 -1927 94 -1926
rect 534 -1927 535 -1926
rect 555 -1927 556 -1926
rect 744 -1927 745 -1926
rect 768 -1927 769 -1926
rect 919 -1927 920 -1926
rect 926 -1927 927 -1926
rect 947 -1927 948 -1926
rect 954 -1927 955 -1926
rect 996 -1927 997 -1926
rect 93 -1929 94 -1928
rect 219 -1929 220 -1928
rect 222 -1929 223 -1928
rect 289 -1929 290 -1928
rect 324 -1929 325 -1928
rect 464 -1929 465 -1928
rect 471 -1929 472 -1928
rect 506 -1929 507 -1928
rect 558 -1929 559 -1928
rect 842 -1929 843 -1928
rect 856 -1929 857 -1928
rect 1069 -1929 1070 -1928
rect 100 -1931 101 -1930
rect 345 -1931 346 -1930
rect 348 -1931 349 -1930
rect 408 -1931 409 -1930
rect 485 -1931 486 -1930
rect 576 -1931 577 -1930
rect 621 -1931 622 -1930
rect 793 -1931 794 -1930
rect 821 -1931 822 -1930
rect 828 -1931 829 -1930
rect 912 -1931 913 -1930
rect 933 -1931 934 -1930
rect 940 -1931 941 -1930
rect 954 -1931 955 -1930
rect 124 -1933 125 -1932
rect 1059 -1933 1060 -1932
rect 128 -1935 129 -1934
rect 376 -1935 377 -1934
rect 387 -1935 388 -1934
rect 401 -1935 402 -1934
rect 506 -1935 507 -1934
rect 737 -1935 738 -1934
rect 824 -1935 825 -1934
rect 828 -1935 829 -1934
rect 835 -1935 836 -1934
rect 940 -1935 941 -1934
rect 1010 -1935 1011 -1934
rect 1059 -1935 1060 -1934
rect 152 -1937 153 -1936
rect 877 -1937 878 -1936
rect 898 -1937 899 -1936
rect 912 -1937 913 -1936
rect 23 -1939 24 -1938
rect 898 -1939 899 -1938
rect 44 -1941 45 -1940
rect 152 -1941 153 -1940
rect 156 -1941 157 -1940
rect 835 -1941 836 -1940
rect 877 -1941 878 -1940
rect 891 -1941 892 -1940
rect 107 -1943 108 -1942
rect 156 -1943 157 -1942
rect 159 -1943 160 -1942
rect 1024 -1943 1025 -1942
rect 107 -1945 108 -1944
rect 142 -1945 143 -1944
rect 184 -1945 185 -1944
rect 268 -1945 269 -1944
rect 338 -1945 339 -1944
rect 457 -1945 458 -1944
rect 576 -1945 577 -1944
rect 611 -1945 612 -1944
rect 621 -1945 622 -1944
rect 1052 -1945 1053 -1944
rect 184 -1947 185 -1946
rect 366 -1947 367 -1946
rect 369 -1947 370 -1946
rect 408 -1947 409 -1946
rect 583 -1947 584 -1946
rect 611 -1947 612 -1946
rect 632 -1947 633 -1946
rect 1038 -1947 1039 -1946
rect 198 -1949 199 -1948
rect 289 -1949 290 -1948
rect 338 -1949 339 -1948
rect 646 -1949 647 -1948
rect 660 -1949 661 -1948
rect 793 -1949 794 -1948
rect 1017 -1949 1018 -1948
rect 1052 -1949 1053 -1948
rect 198 -1951 199 -1950
rect 282 -1951 283 -1950
rect 345 -1951 346 -1950
rect 401 -1951 402 -1950
rect 569 -1951 570 -1950
rect 583 -1951 584 -1950
rect 635 -1951 636 -1950
rect 723 -1951 724 -1950
rect 989 -1951 990 -1950
rect 1017 -1951 1018 -1950
rect 23 -1953 24 -1952
rect 723 -1953 724 -1952
rect 807 -1953 808 -1952
rect 989 -1953 990 -1952
rect 54 -1955 55 -1954
rect 569 -1955 570 -1954
rect 635 -1955 636 -1954
rect 772 -1955 773 -1954
rect 807 -1955 808 -1954
rect 884 -1955 885 -1954
rect 54 -1957 55 -1956
rect 226 -1957 227 -1956
rect 229 -1957 230 -1956
rect 296 -1957 297 -1956
rect 352 -1957 353 -1956
rect 415 -1957 416 -1956
rect 646 -1957 647 -1956
rect 905 -1957 906 -1956
rect 180 -1959 181 -1958
rect 415 -1959 416 -1958
rect 625 -1959 626 -1958
rect 905 -1959 906 -1958
rect 117 -1961 118 -1960
rect 625 -1961 626 -1960
rect 660 -1961 661 -1960
rect 779 -1961 780 -1960
rect 863 -1961 864 -1960
rect 884 -1961 885 -1960
rect 208 -1963 209 -1962
rect 982 -1963 983 -1962
rect 149 -1965 150 -1964
rect 982 -1965 983 -1964
rect 222 -1967 223 -1966
rect 261 -1967 262 -1966
rect 275 -1967 276 -1966
rect 282 -1967 283 -1966
rect 331 -1967 332 -1966
rect 352 -1967 353 -1966
rect 359 -1967 360 -1966
rect 1010 -1967 1011 -1966
rect 163 -1969 164 -1968
rect 275 -1969 276 -1968
rect 331 -1969 332 -1968
rect 373 -1969 374 -1968
rect 390 -1969 391 -1968
rect 891 -1969 892 -1968
rect 163 -1971 164 -1970
rect 530 -1971 531 -1970
rect 670 -1971 671 -1970
rect 849 -1971 850 -1970
rect 240 -1973 241 -1972
rect 422 -1973 423 -1972
rect 681 -1973 682 -1972
rect 737 -1973 738 -1972
rect 751 -1973 752 -1972
rect 863 -1973 864 -1972
rect 240 -1975 241 -1974
rect 254 -1975 255 -1974
rect 359 -1975 360 -1974
rect 380 -1975 381 -1974
rect 667 -1975 668 -1974
rect 681 -1975 682 -1974
rect 688 -1975 689 -1974
rect 961 -1975 962 -1974
rect 86 -1977 87 -1976
rect 380 -1977 381 -1976
rect 520 -1977 521 -1976
rect 667 -1977 668 -1976
rect 674 -1977 675 -1976
rect 961 -1977 962 -1976
rect 61 -1979 62 -1978
rect 520 -1979 521 -1978
rect 597 -1979 598 -1978
rect 688 -1979 689 -1978
rect 695 -1979 696 -1978
rect 709 -1979 710 -1978
rect 751 -1979 752 -1978
rect 814 -1979 815 -1978
rect 233 -1981 234 -1980
rect 597 -1981 598 -1980
rect 649 -1981 650 -1980
rect 814 -1981 815 -1980
rect 212 -1983 213 -1982
rect 233 -1983 234 -1982
rect 247 -1983 248 -1982
rect 730 -1983 731 -1982
rect 758 -1983 759 -1982
rect 772 -1983 773 -1982
rect 121 -1985 122 -1984
rect 212 -1985 213 -1984
rect 254 -1985 255 -1984
rect 303 -1985 304 -1984
rect 373 -1985 374 -1984
rect 464 -1985 465 -1984
rect 653 -1985 654 -1984
rect 674 -1985 675 -1984
rect 709 -1985 710 -1984
rect 716 -1985 717 -1984
rect 730 -1985 731 -1984
rect 800 -1985 801 -1984
rect 121 -1987 122 -1986
rect 205 -1987 206 -1986
rect 303 -1987 304 -1986
rect 310 -1987 311 -1986
rect 548 -1987 549 -1986
rect 716 -1987 717 -1986
rect 758 -1987 759 -1986
rect 765 -1987 766 -1986
rect 170 -1989 171 -1988
rect 800 -1989 801 -1988
rect 170 -1991 171 -1990
rect 177 -1991 178 -1990
rect 205 -1991 206 -1990
rect 499 -1991 500 -1990
rect 548 -1991 549 -1990
rect 1104 -1991 1105 -1990
rect 310 -1993 311 -1992
rect 541 -1993 542 -1992
rect 639 -1993 640 -1992
rect 653 -1993 654 -1992
rect 317 -1995 318 -1994
rect 765 -1995 766 -1994
rect 317 -1997 318 -1996
rect 436 -1997 437 -1996
rect 513 -1997 514 -1996
rect 541 -1997 542 -1996
rect 590 -1997 591 -1996
rect 639 -1997 640 -1996
rect 261 -1999 262 -1998
rect 436 -1999 437 -1998
rect 2 -2010 3 -2009
rect 222 -2010 223 -2009
rect 229 -2010 230 -2009
rect 373 -2010 374 -2009
rect 376 -2010 377 -2009
rect 898 -2010 899 -2009
rect 926 -2010 927 -2009
rect 933 -2010 934 -2009
rect 943 -2010 944 -2009
rect 1017 -2010 1018 -2009
rect 1080 -2010 1081 -2009
rect 1094 -2010 1095 -2009
rect 1104 -2010 1105 -2009
rect 1108 -2010 1109 -2009
rect 1115 -2010 1116 -2009
rect 1122 -2010 1123 -2009
rect 9 -2012 10 -2011
rect 23 -2012 24 -2011
rect 33 -2012 34 -2011
rect 1024 -2012 1025 -2011
rect 1038 -2012 1039 -2011
rect 1080 -2012 1081 -2011
rect 9 -2014 10 -2013
rect 163 -2014 164 -2013
rect 170 -2014 171 -2013
rect 226 -2014 227 -2013
rect 275 -2014 276 -2013
rect 436 -2014 437 -2013
rect 439 -2014 440 -2013
rect 1066 -2014 1067 -2013
rect 1073 -2014 1074 -2013
rect 1108 -2014 1109 -2013
rect 16 -2016 17 -2015
rect 345 -2016 346 -2015
rect 348 -2016 349 -2015
rect 800 -2016 801 -2015
rect 807 -2016 808 -2015
rect 933 -2016 934 -2015
rect 982 -2016 983 -2015
rect 1017 -2016 1018 -2015
rect 1031 -2016 1032 -2015
rect 1038 -2016 1039 -2015
rect 1045 -2016 1046 -2015
rect 1073 -2016 1074 -2015
rect 16 -2018 17 -2017
rect 100 -2018 101 -2017
rect 107 -2018 108 -2017
rect 583 -2018 584 -2017
rect 593 -2018 594 -2017
rect 961 -2018 962 -2017
rect 996 -2018 997 -2017
rect 1024 -2018 1025 -2017
rect 1059 -2018 1060 -2017
rect 1094 -2018 1095 -2017
rect 51 -2020 52 -2019
rect 835 -2020 836 -2019
rect 863 -2020 864 -2019
rect 898 -2020 899 -2019
rect 929 -2020 930 -2019
rect 968 -2020 969 -2019
rect 1003 -2020 1004 -2019
rect 1045 -2020 1046 -2019
rect 54 -2022 55 -2021
rect 345 -2022 346 -2021
rect 380 -2022 381 -2021
rect 460 -2022 461 -2021
rect 464 -2022 465 -2021
rect 646 -2022 647 -2021
rect 688 -2022 689 -2021
rect 779 -2022 780 -2021
rect 782 -2022 783 -2021
rect 821 -2022 822 -2021
rect 835 -2022 836 -2021
rect 912 -2022 913 -2021
rect 940 -2022 941 -2021
rect 961 -2022 962 -2021
rect 975 -2022 976 -2021
rect 1003 -2022 1004 -2021
rect 1010 -2022 1011 -2021
rect 1066 -2022 1067 -2021
rect 37 -2024 38 -2023
rect 380 -2024 381 -2023
rect 394 -2024 395 -2023
rect 646 -2024 647 -2023
rect 691 -2024 692 -2023
rect 1059 -2024 1060 -2023
rect 37 -2026 38 -2025
rect 177 -2026 178 -2025
rect 180 -2026 181 -2025
rect 233 -2026 234 -2025
rect 275 -2026 276 -2025
rect 471 -2026 472 -2025
rect 502 -2026 503 -2025
rect 905 -2026 906 -2025
rect 954 -2026 955 -2025
rect 982 -2026 983 -2025
rect 44 -2028 45 -2027
rect 464 -2028 465 -2027
rect 471 -2028 472 -2027
rect 530 -2028 531 -2027
rect 569 -2028 570 -2027
rect 632 -2028 633 -2027
rect 716 -2028 717 -2027
rect 905 -2028 906 -2027
rect 44 -2030 45 -2029
rect 212 -2030 213 -2029
rect 222 -2030 223 -2029
rect 604 -2030 605 -2029
rect 611 -2030 612 -2029
rect 1115 -2030 1116 -2029
rect 58 -2032 59 -2031
rect 75 -2032 76 -2031
rect 79 -2032 80 -2031
rect 170 -2032 171 -2031
rect 177 -2032 178 -2031
rect 282 -2032 283 -2031
rect 324 -2032 325 -2031
rect 355 -2032 356 -2031
rect 394 -2032 395 -2031
rect 418 -2032 419 -2031
rect 478 -2032 479 -2031
rect 604 -2032 605 -2031
rect 625 -2032 626 -2031
rect 1031 -2032 1032 -2031
rect 58 -2034 59 -2033
rect 849 -2034 850 -2033
rect 870 -2034 871 -2033
rect 975 -2034 976 -2033
rect 65 -2036 66 -2035
rect 366 -2036 367 -2035
rect 408 -2036 409 -2035
rect 534 -2036 535 -2035
rect 579 -2036 580 -2035
rect 779 -2036 780 -2035
rect 821 -2036 822 -2035
rect 828 -2036 829 -2035
rect 842 -2036 843 -2035
rect 863 -2036 864 -2035
rect 877 -2036 878 -2035
rect 996 -2036 997 -2035
rect 65 -2038 66 -2037
rect 128 -2038 129 -2037
rect 135 -2038 136 -2037
rect 492 -2038 493 -2037
rect 513 -2038 514 -2037
rect 723 -2038 724 -2037
rect 744 -2038 745 -2037
rect 772 -2038 773 -2037
rect 842 -2038 843 -2037
rect 891 -2038 892 -2037
rect 51 -2040 52 -2039
rect 135 -2040 136 -2039
rect 149 -2040 150 -2039
rect 527 -2040 528 -2039
rect 534 -2040 535 -2039
rect 562 -2040 563 -2039
rect 667 -2040 668 -2039
rect 870 -2040 871 -2039
rect 884 -2040 885 -2039
rect 1010 -2040 1011 -2039
rect 72 -2042 73 -2041
rect 107 -2042 108 -2041
rect 110 -2042 111 -2041
rect 156 -2042 157 -2041
rect 184 -2042 185 -2041
rect 635 -2042 636 -2041
rect 695 -2042 696 -2041
rect 723 -2042 724 -2041
rect 751 -2042 752 -2041
rect 772 -2042 773 -2041
rect 891 -2042 892 -2041
rect 989 -2042 990 -2041
rect 75 -2044 76 -2043
rect 590 -2044 591 -2043
rect 695 -2044 696 -2043
rect 730 -2044 731 -2043
rect 758 -2044 759 -2043
rect 807 -2044 808 -2043
rect 79 -2046 80 -2045
rect 422 -2046 423 -2045
rect 429 -2046 430 -2045
rect 478 -2046 479 -2045
rect 492 -2046 493 -2045
rect 499 -2046 500 -2045
rect 506 -2046 507 -2045
rect 744 -2046 745 -2045
rect 761 -2046 762 -2045
rect 1087 -2046 1088 -2045
rect 86 -2048 87 -2047
rect 800 -2048 801 -2047
rect 814 -2048 815 -2047
rect 1087 -2048 1088 -2047
rect 86 -2050 87 -2049
rect 751 -2050 752 -2049
rect 765 -2050 766 -2049
rect 1052 -2050 1053 -2049
rect 96 -2052 97 -2051
rect 793 -2052 794 -2051
rect 100 -2054 101 -2053
rect 114 -2054 115 -2053
rect 117 -2054 118 -2053
rect 163 -2054 164 -2053
rect 184 -2054 185 -2053
rect 618 -2054 619 -2053
rect 688 -2054 689 -2053
rect 793 -2054 794 -2053
rect 114 -2056 115 -2055
rect 373 -2056 374 -2055
rect 401 -2056 402 -2055
rect 422 -2056 423 -2055
rect 443 -2056 444 -2055
rect 667 -2056 668 -2055
rect 709 -2056 710 -2055
rect 730 -2056 731 -2055
rect 768 -2056 769 -2055
rect 884 -2056 885 -2055
rect 121 -2058 122 -2057
rect 205 -2058 206 -2057
rect 226 -2058 227 -2057
rect 614 -2058 615 -2057
rect 618 -2058 619 -2057
rect 681 -2058 682 -2057
rect 786 -2058 787 -2057
rect 814 -2058 815 -2057
rect 82 -2060 83 -2059
rect 121 -2060 122 -2059
rect 128 -2060 129 -2059
rect 331 -2060 332 -2059
rect 338 -2060 339 -2059
rect 527 -2060 528 -2059
rect 555 -2060 556 -2059
rect 765 -2060 766 -2059
rect 110 -2062 111 -2061
rect 338 -2062 339 -2061
rect 366 -2062 367 -2061
rect 548 -2062 549 -2061
rect 572 -2062 573 -2061
rect 786 -2062 787 -2061
rect 138 -2064 139 -2063
rect 681 -2064 682 -2063
rect 138 -2066 139 -2065
rect 912 -2066 913 -2065
rect 142 -2068 143 -2067
rect 156 -2068 157 -2067
rect 198 -2068 199 -2067
rect 233 -2068 234 -2067
rect 247 -2068 248 -2067
rect 429 -2068 430 -2067
rect 443 -2068 444 -2067
rect 597 -2068 598 -2067
rect 674 -2068 675 -2067
rect 709 -2068 710 -2067
rect 26 -2070 27 -2069
rect 597 -2070 598 -2069
rect 89 -2072 90 -2071
rect 198 -2072 199 -2071
rect 247 -2072 248 -2071
rect 296 -2072 297 -2071
rect 310 -2072 311 -2071
rect 590 -2072 591 -2071
rect 89 -2074 90 -2073
rect 737 -2074 738 -2073
rect 149 -2076 150 -2075
rect 212 -2076 213 -2075
rect 254 -2076 255 -2075
rect 499 -2076 500 -2075
rect 516 -2076 517 -2075
rect 989 -2076 990 -2075
rect 152 -2078 153 -2077
rect 191 -2078 192 -2077
rect 240 -2078 241 -2077
rect 254 -2078 255 -2077
rect 282 -2078 283 -2077
rect 352 -2078 353 -2077
rect 369 -2078 370 -2077
rect 828 -2078 829 -2077
rect 152 -2080 153 -2079
rect 968 -2080 969 -2079
rect 191 -2082 192 -2081
rect 268 -2082 269 -2081
rect 289 -2082 290 -2081
rect 310 -2082 311 -2081
rect 324 -2082 325 -2081
rect 352 -2082 353 -2081
rect 387 -2082 388 -2081
rect 401 -2082 402 -2081
rect 411 -2082 412 -2081
rect 954 -2082 955 -2081
rect 240 -2084 241 -2083
rect 450 -2084 451 -2083
rect 457 -2084 458 -2083
rect 506 -2084 507 -2083
rect 520 -2084 521 -2083
rect 562 -2084 563 -2083
rect 576 -2084 577 -2083
rect 674 -2084 675 -2083
rect 737 -2084 738 -2083
rect 877 -2084 878 -2083
rect 142 -2086 143 -2085
rect 450 -2086 451 -2085
rect 541 -2086 542 -2085
rect 555 -2086 556 -2085
rect 268 -2088 269 -2087
rect 453 -2088 454 -2087
rect 541 -2088 542 -2087
rect 758 -2088 759 -2087
rect 289 -2090 290 -2089
rect 856 -2090 857 -2089
rect 296 -2092 297 -2091
rect 303 -2092 304 -2091
rect 317 -2092 318 -2091
rect 387 -2092 388 -2091
rect 411 -2092 412 -2091
rect 639 -2092 640 -2091
rect 303 -2094 304 -2093
rect 649 -2094 650 -2093
rect 317 -2096 318 -2095
rect 359 -2096 360 -2095
rect 415 -2096 416 -2095
rect 583 -2096 584 -2095
rect 639 -2096 640 -2095
rect 856 -2096 857 -2095
rect 261 -2098 262 -2097
rect 359 -2098 360 -2097
rect 415 -2098 416 -2097
rect 849 -2098 850 -2097
rect 93 -2100 94 -2099
rect 261 -2100 262 -2099
rect 331 -2100 332 -2099
rect 642 -2100 643 -2099
rect 93 -2102 94 -2101
rect 1101 -2102 1102 -2101
rect 341 -2104 342 -2103
rect 520 -2104 521 -2103
rect 548 -2104 549 -2103
rect 660 -2104 661 -2103
rect 716 -2104 717 -2103
rect 1101 -2104 1102 -2103
rect 485 -2106 486 -2105
rect 660 -2106 661 -2105
rect 485 -2108 486 -2107
rect 702 -2108 703 -2107
rect 653 -2110 654 -2109
rect 702 -2110 703 -2109
rect 653 -2112 654 -2111
rect 1052 -2112 1053 -2111
rect 9 -2123 10 -2122
rect 397 -2123 398 -2122
rect 401 -2123 402 -2122
rect 418 -2123 419 -2122
rect 432 -2123 433 -2122
rect 604 -2123 605 -2122
rect 611 -2123 612 -2122
rect 1115 -2123 1116 -2122
rect 9 -2125 10 -2124
rect 254 -2125 255 -2124
rect 275 -2125 276 -2124
rect 415 -2125 416 -2124
rect 436 -2125 437 -2124
rect 579 -2125 580 -2124
rect 590 -2125 591 -2124
rect 628 -2125 629 -2124
rect 642 -2125 643 -2124
rect 1010 -2125 1011 -2124
rect 1052 -2125 1053 -2124
rect 1055 -2125 1056 -2124
rect 1101 -2125 1102 -2124
rect 1122 -2125 1123 -2124
rect 16 -2127 17 -2126
rect 457 -2127 458 -2126
rect 485 -2127 486 -2126
rect 499 -2127 500 -2126
rect 523 -2127 524 -2126
rect 807 -2127 808 -2126
rect 873 -2127 874 -2126
rect 961 -2127 962 -2126
rect 16 -2129 17 -2128
rect 89 -2129 90 -2128
rect 93 -2129 94 -2128
rect 275 -2129 276 -2128
rect 282 -2129 283 -2128
rect 338 -2129 339 -2128
rect 359 -2129 360 -2128
rect 569 -2129 570 -2128
rect 576 -2129 577 -2128
rect 982 -2129 983 -2128
rect 23 -2131 24 -2130
rect 149 -2131 150 -2130
rect 152 -2131 153 -2130
rect 366 -2131 367 -2130
rect 373 -2131 374 -2130
rect 450 -2131 451 -2130
rect 485 -2131 486 -2130
rect 541 -2131 542 -2130
rect 548 -2131 549 -2130
rect 562 -2131 563 -2130
rect 565 -2131 566 -2130
rect 1017 -2131 1018 -2130
rect 23 -2133 24 -2132
rect 583 -2133 584 -2132
rect 604 -2133 605 -2132
rect 1045 -2133 1046 -2132
rect 30 -2135 31 -2134
rect 40 -2135 41 -2134
rect 58 -2135 59 -2134
rect 170 -2135 171 -2134
rect 173 -2135 174 -2134
rect 345 -2135 346 -2134
rect 366 -2135 367 -2134
rect 380 -2135 381 -2134
rect 394 -2135 395 -2134
rect 583 -2135 584 -2134
rect 611 -2135 612 -2134
rect 709 -2135 710 -2134
rect 730 -2135 731 -2134
rect 733 -2135 734 -2134
rect 737 -2135 738 -2134
rect 996 -2135 997 -2134
rect 1017 -2135 1018 -2134
rect 1094 -2135 1095 -2134
rect 51 -2137 52 -2136
rect 380 -2137 381 -2136
rect 401 -2137 402 -2136
rect 670 -2137 671 -2136
rect 684 -2137 685 -2136
rect 975 -2137 976 -2136
rect 982 -2137 983 -2136
rect 1087 -2137 1088 -2136
rect 51 -2139 52 -2138
rect 338 -2139 339 -2138
rect 376 -2139 377 -2138
rect 408 -2139 409 -2138
rect 415 -2139 416 -2138
rect 698 -2139 699 -2138
rect 723 -2139 724 -2138
rect 737 -2139 738 -2138
rect 807 -2139 808 -2138
rect 877 -2139 878 -2138
rect 940 -2139 941 -2138
rect 954 -2139 955 -2138
rect 961 -2139 962 -2138
rect 1024 -2139 1025 -2138
rect 1038 -2139 1039 -2138
rect 1045 -2139 1046 -2138
rect 58 -2141 59 -2140
rect 387 -2141 388 -2140
rect 408 -2141 409 -2140
rect 492 -2141 493 -2140
rect 530 -2141 531 -2140
rect 989 -2141 990 -2140
rect 61 -2143 62 -2142
rect 541 -2143 542 -2142
rect 548 -2143 549 -2142
rect 551 -2143 552 -2142
rect 555 -2143 556 -2142
rect 572 -2143 573 -2142
rect 593 -2143 594 -2142
rect 1024 -2143 1025 -2142
rect 72 -2145 73 -2144
rect 506 -2145 507 -2144
rect 534 -2145 535 -2144
rect 600 -2145 601 -2144
rect 625 -2145 626 -2144
rect 1003 -2145 1004 -2144
rect 75 -2147 76 -2146
rect 1010 -2147 1011 -2146
rect 75 -2149 76 -2148
rect 660 -2149 661 -2148
rect 691 -2149 692 -2148
rect 814 -2149 815 -2148
rect 891 -2149 892 -2148
rect 954 -2149 955 -2148
rect 989 -2149 990 -2148
rect 1108 -2149 1109 -2148
rect 79 -2151 80 -2150
rect 800 -2151 801 -2150
rect 814 -2151 815 -2150
rect 828 -2151 829 -2150
rect 835 -2151 836 -2150
rect 891 -2151 892 -2150
rect 947 -2151 948 -2150
rect 996 -2151 997 -2150
rect 1003 -2151 1004 -2150
rect 1080 -2151 1081 -2150
rect 79 -2153 80 -2152
rect 191 -2153 192 -2152
rect 219 -2153 220 -2152
rect 341 -2153 342 -2152
rect 443 -2153 444 -2152
rect 509 -2153 510 -2152
rect 534 -2153 535 -2152
rect 667 -2153 668 -2152
rect 695 -2153 696 -2152
rect 877 -2153 878 -2152
rect 947 -2153 948 -2152
rect 968 -2153 969 -2152
rect 86 -2155 87 -2154
rect 471 -2155 472 -2154
rect 527 -2155 528 -2154
rect 968 -2155 969 -2154
rect 72 -2157 73 -2156
rect 86 -2157 87 -2156
rect 93 -2157 94 -2156
rect 191 -2157 192 -2156
rect 226 -2157 227 -2156
rect 576 -2157 577 -2156
rect 625 -2157 626 -2156
rect 702 -2157 703 -2156
rect 730 -2157 731 -2156
rect 842 -2157 843 -2156
rect 96 -2159 97 -2158
rect 597 -2159 598 -2158
rect 653 -2159 654 -2158
rect 695 -2159 696 -2158
rect 702 -2159 703 -2158
rect 772 -2159 773 -2158
rect 786 -2159 787 -2158
rect 800 -2159 801 -2158
rect 828 -2159 829 -2158
rect 863 -2159 864 -2158
rect 107 -2161 108 -2160
rect 289 -2161 290 -2160
rect 317 -2161 318 -2160
rect 387 -2161 388 -2160
rect 443 -2161 444 -2160
rect 464 -2161 465 -2160
rect 471 -2161 472 -2160
rect 761 -2161 762 -2160
rect 765 -2161 766 -2160
rect 772 -2161 773 -2160
rect 779 -2161 780 -2160
rect 786 -2161 787 -2160
rect 835 -2161 836 -2160
rect 870 -2161 871 -2160
rect 37 -2163 38 -2162
rect 779 -2163 780 -2162
rect 863 -2163 864 -2162
rect 905 -2163 906 -2162
rect 44 -2165 45 -2164
rect 289 -2165 290 -2164
rect 320 -2165 321 -2164
rect 975 -2165 976 -2164
rect 44 -2167 45 -2166
rect 212 -2167 213 -2166
rect 226 -2167 227 -2166
rect 303 -2167 304 -2166
rect 324 -2167 325 -2166
rect 359 -2167 360 -2166
rect 453 -2167 454 -2166
rect 1038 -2167 1039 -2166
rect 107 -2169 108 -2168
rect 166 -2169 167 -2168
rect 177 -2169 178 -2168
rect 282 -2169 283 -2168
rect 303 -2169 304 -2168
rect 429 -2169 430 -2168
rect 464 -2169 465 -2168
rect 478 -2169 479 -2168
rect 527 -2169 528 -2168
rect 726 -2169 727 -2168
rect 744 -2169 745 -2168
rect 842 -2169 843 -2168
rect 905 -2169 906 -2168
rect 1031 -2169 1032 -2168
rect 65 -2171 66 -2170
rect 177 -2171 178 -2170
rect 198 -2171 199 -2170
rect 324 -2171 325 -2170
rect 345 -2171 346 -2170
rect 429 -2171 430 -2170
rect 555 -2171 556 -2170
rect 632 -2171 633 -2170
rect 656 -2171 657 -2170
rect 1073 -2171 1074 -2170
rect 65 -2173 66 -2172
rect 268 -2173 269 -2172
rect 422 -2173 423 -2172
rect 478 -2173 479 -2172
rect 597 -2173 598 -2172
rect 933 -2173 934 -2172
rect 110 -2175 111 -2174
rect 590 -2175 591 -2174
rect 632 -2175 633 -2174
rect 646 -2175 647 -2174
rect 660 -2175 661 -2174
rect 681 -2175 682 -2174
rect 733 -2175 734 -2174
rect 744 -2175 745 -2174
rect 751 -2175 752 -2174
rect 765 -2175 766 -2174
rect 114 -2177 115 -2176
rect 121 -2177 122 -2176
rect 128 -2177 129 -2176
rect 135 -2177 136 -2176
rect 138 -2177 139 -2176
rect 856 -2177 857 -2176
rect 82 -2179 83 -2178
rect 128 -2179 129 -2178
rect 142 -2179 143 -2178
rect 502 -2179 503 -2178
rect 513 -2179 514 -2178
rect 751 -2179 752 -2178
rect 117 -2181 118 -2180
rect 793 -2181 794 -2180
rect 142 -2183 143 -2182
rect 240 -2183 241 -2182
rect 261 -2183 262 -2182
rect 341 -2183 342 -2182
rect 422 -2183 423 -2182
rect 740 -2183 741 -2182
rect 149 -2185 150 -2184
rect 156 -2185 157 -2184
rect 163 -2185 164 -2184
rect 254 -2185 255 -2184
rect 261 -2185 262 -2184
rect 296 -2185 297 -2184
rect 436 -2185 437 -2184
rect 933 -2185 934 -2184
rect 121 -2187 122 -2186
rect 296 -2187 297 -2186
rect 513 -2187 514 -2186
rect 723 -2187 724 -2186
rect 124 -2189 125 -2188
rect 156 -2189 157 -2188
rect 184 -2189 185 -2188
rect 240 -2189 241 -2188
rect 268 -2189 269 -2188
rect 331 -2189 332 -2188
rect 639 -2189 640 -2188
rect 793 -2189 794 -2188
rect 2 -2191 3 -2190
rect 639 -2191 640 -2190
rect 646 -2191 647 -2190
rect 674 -2191 675 -2190
rect 688 -2191 689 -2190
rect 856 -2191 857 -2190
rect 2 -2193 3 -2192
rect 758 -2193 759 -2192
rect 124 -2195 125 -2194
rect 1031 -2195 1032 -2194
rect 198 -2197 199 -2196
rect 355 -2197 356 -2196
rect 667 -2197 668 -2196
rect 1066 -2197 1067 -2196
rect 212 -2199 213 -2198
rect 292 -2199 293 -2198
rect 310 -2199 311 -2198
rect 331 -2199 332 -2198
rect 674 -2199 675 -2198
rect 716 -2199 717 -2198
rect 758 -2199 759 -2198
rect 912 -2199 913 -2198
rect 233 -2201 234 -2200
rect 439 -2201 440 -2200
rect 618 -2201 619 -2200
rect 716 -2201 717 -2200
rect 912 -2201 913 -2200
rect 919 -2201 920 -2200
rect 205 -2203 206 -2202
rect 233 -2203 234 -2202
rect 247 -2203 248 -2202
rect 310 -2203 311 -2202
rect 520 -2203 521 -2202
rect 618 -2203 619 -2202
rect 919 -2203 920 -2202
rect 926 -2203 927 -2202
rect 205 -2205 206 -2204
rect 492 -2205 493 -2204
rect 520 -2205 521 -2204
rect 709 -2205 710 -2204
rect 926 -2205 927 -2204
rect 1059 -2205 1060 -2204
rect 247 -2207 248 -2206
rect 607 -2207 608 -2206
rect 9 -2218 10 -2217
rect 205 -2218 206 -2217
rect 208 -2218 209 -2217
rect 639 -2218 640 -2217
rect 653 -2218 654 -2217
rect 670 -2218 671 -2217
rect 691 -2218 692 -2217
rect 863 -2218 864 -2217
rect 870 -2218 871 -2217
rect 968 -2218 969 -2217
rect 9 -2220 10 -2219
rect 338 -2220 339 -2219
rect 341 -2220 342 -2219
rect 485 -2220 486 -2219
rect 488 -2220 489 -2219
rect 779 -2220 780 -2219
rect 856 -2220 857 -2219
rect 929 -2220 930 -2219
rect 16 -2222 17 -2221
rect 103 -2222 104 -2221
rect 121 -2222 122 -2221
rect 254 -2222 255 -2221
rect 282 -2222 283 -2221
rect 317 -2222 318 -2221
rect 348 -2222 349 -2221
rect 366 -2222 367 -2221
rect 373 -2222 374 -2221
rect 471 -2222 472 -2221
rect 485 -2222 486 -2221
rect 688 -2222 689 -2221
rect 695 -2222 696 -2221
rect 982 -2222 983 -2221
rect 30 -2224 31 -2223
rect 345 -2224 346 -2223
rect 355 -2224 356 -2223
rect 387 -2224 388 -2223
rect 394 -2224 395 -2223
rect 1031 -2224 1032 -2223
rect 44 -2226 45 -2225
rect 383 -2226 384 -2225
rect 387 -2226 388 -2225
rect 422 -2226 423 -2225
rect 436 -2226 437 -2225
rect 681 -2226 682 -2225
rect 695 -2226 696 -2225
rect 737 -2226 738 -2225
rect 768 -2226 769 -2225
rect 800 -2226 801 -2225
rect 856 -2226 857 -2225
rect 1017 -2226 1018 -2225
rect 37 -2228 38 -2227
rect 44 -2228 45 -2227
rect 51 -2228 52 -2227
rect 191 -2228 192 -2227
rect 194 -2228 195 -2227
rect 212 -2228 213 -2227
rect 215 -2228 216 -2227
rect 296 -2228 297 -2227
rect 310 -2228 311 -2227
rect 338 -2228 339 -2227
rect 359 -2228 360 -2227
rect 394 -2228 395 -2227
rect 401 -2228 402 -2227
rect 422 -2228 423 -2227
rect 439 -2228 440 -2227
rect 1010 -2228 1011 -2227
rect 30 -2230 31 -2229
rect 51 -2230 52 -2229
rect 93 -2230 94 -2229
rect 173 -2230 174 -2229
rect 177 -2230 178 -2229
rect 303 -2230 304 -2229
rect 317 -2230 318 -2229
rect 324 -2230 325 -2229
rect 331 -2230 332 -2229
rect 355 -2230 356 -2229
rect 359 -2230 360 -2229
rect 579 -2230 580 -2229
rect 590 -2230 591 -2229
rect 835 -2230 836 -2229
rect 863 -2230 864 -2229
rect 1024 -2230 1025 -2229
rect 23 -2232 24 -2231
rect 303 -2232 304 -2231
rect 331 -2232 332 -2231
rect 499 -2232 500 -2231
rect 502 -2232 503 -2231
rect 520 -2232 521 -2231
rect 548 -2232 549 -2231
rect 569 -2232 570 -2231
rect 572 -2232 573 -2231
rect 702 -2232 703 -2231
rect 723 -2232 724 -2231
rect 814 -2232 815 -2231
rect 835 -2232 836 -2231
rect 961 -2232 962 -2231
rect 23 -2234 24 -2233
rect 163 -2234 164 -2233
rect 166 -2234 167 -2233
rect 544 -2234 545 -2233
rect 576 -2234 577 -2233
rect 639 -2234 640 -2233
rect 653 -2234 654 -2233
rect 709 -2234 710 -2233
rect 723 -2234 724 -2233
rect 772 -2234 773 -2233
rect 779 -2234 780 -2233
rect 793 -2234 794 -2233
rect 800 -2234 801 -2233
rect 912 -2234 913 -2233
rect 922 -2234 923 -2233
rect 996 -2234 997 -2233
rect 37 -2236 38 -2235
rect 142 -2236 143 -2235
rect 156 -2236 157 -2235
rect 184 -2236 185 -2235
rect 201 -2236 202 -2235
rect 565 -2236 566 -2235
rect 590 -2236 591 -2235
rect 632 -2236 633 -2235
rect 667 -2236 668 -2235
rect 730 -2236 731 -2235
rect 737 -2236 738 -2235
rect 786 -2236 787 -2235
rect 793 -2236 794 -2235
rect 940 -2236 941 -2235
rect 961 -2236 962 -2235
rect 1003 -2236 1004 -2235
rect 2 -2238 3 -2237
rect 142 -2238 143 -2237
rect 170 -2238 171 -2237
rect 275 -2238 276 -2237
rect 282 -2238 283 -2237
rect 397 -2238 398 -2237
rect 401 -2238 402 -2237
rect 492 -2238 493 -2237
rect 506 -2238 507 -2237
rect 555 -2238 556 -2237
rect 597 -2238 598 -2237
rect 716 -2238 717 -2237
rect 726 -2238 727 -2237
rect 1045 -2238 1046 -2237
rect 2 -2240 3 -2239
rect 114 -2240 115 -2239
rect 121 -2240 122 -2239
rect 583 -2240 584 -2239
rect 604 -2240 605 -2239
rect 618 -2240 619 -2239
rect 681 -2240 682 -2239
rect 730 -2240 731 -2239
rect 758 -2240 759 -2239
rect 786 -2240 787 -2239
rect 814 -2240 815 -2239
rect 828 -2240 829 -2239
rect 940 -2240 941 -2239
rect 989 -2240 990 -2239
rect 79 -2242 80 -2241
rect 163 -2242 164 -2241
rect 198 -2242 199 -2241
rect 275 -2242 276 -2241
rect 296 -2242 297 -2241
rect 327 -2242 328 -2241
rect 408 -2242 409 -2241
rect 509 -2242 510 -2241
rect 513 -2242 514 -2241
rect 632 -2242 633 -2241
rect 698 -2242 699 -2241
rect 905 -2242 906 -2241
rect 93 -2244 94 -2243
rect 107 -2244 108 -2243
rect 114 -2244 115 -2243
rect 128 -2244 129 -2243
rect 135 -2244 136 -2243
rect 292 -2244 293 -2243
rect 380 -2244 381 -2243
rect 408 -2244 409 -2243
rect 429 -2244 430 -2243
rect 513 -2244 514 -2243
rect 527 -2244 528 -2243
rect 555 -2244 556 -2243
rect 583 -2244 584 -2243
rect 842 -2244 843 -2243
rect 100 -2246 101 -2245
rect 107 -2246 108 -2245
rect 135 -2246 136 -2245
rect 149 -2246 150 -2245
rect 156 -2246 157 -2245
rect 198 -2246 199 -2245
rect 205 -2246 206 -2245
rect 219 -2246 220 -2245
rect 226 -2246 227 -2245
rect 380 -2246 381 -2245
rect 429 -2246 430 -2245
rect 541 -2246 542 -2245
rect 548 -2246 549 -2245
rect 576 -2246 577 -2245
rect 604 -2246 605 -2245
rect 646 -2246 647 -2245
rect 709 -2246 710 -2245
rect 765 -2246 766 -2245
rect 772 -2246 773 -2245
rect 849 -2246 850 -2245
rect 65 -2248 66 -2247
rect 149 -2248 150 -2247
rect 212 -2248 213 -2247
rect 268 -2248 269 -2247
rect 450 -2248 451 -2247
rect 562 -2248 563 -2247
rect 618 -2248 619 -2247
rect 625 -2248 626 -2247
rect 646 -2248 647 -2247
rect 684 -2248 685 -2247
rect 716 -2248 717 -2247
rect 891 -2248 892 -2247
rect 33 -2250 34 -2249
rect 268 -2250 269 -2249
rect 450 -2250 451 -2249
rect 744 -2250 745 -2249
rect 758 -2250 759 -2249
rect 821 -2250 822 -2249
rect 828 -2250 829 -2249
rect 933 -2250 934 -2249
rect 65 -2252 66 -2251
rect 187 -2252 188 -2251
rect 226 -2252 227 -2251
rect 289 -2252 290 -2251
rect 352 -2252 353 -2251
rect 744 -2252 745 -2251
rect 821 -2252 822 -2251
rect 975 -2252 976 -2251
rect 72 -2254 73 -2253
rect 219 -2254 220 -2253
rect 240 -2254 241 -2253
rect 324 -2254 325 -2253
rect 352 -2254 353 -2253
rect 464 -2254 465 -2253
rect 467 -2254 468 -2253
rect 527 -2254 528 -2253
rect 541 -2254 542 -2253
rect 877 -2254 878 -2253
rect 891 -2254 892 -2253
rect 1038 -2254 1039 -2253
rect 240 -2256 241 -2255
rect 415 -2256 416 -2255
rect 457 -2256 458 -2255
rect 481 -2256 482 -2255
rect 593 -2256 594 -2255
rect 625 -2256 626 -2255
rect 684 -2256 685 -2255
rect 702 -2256 703 -2255
rect 842 -2256 843 -2255
rect 919 -2256 920 -2255
rect 968 -2256 969 -2255
rect 975 -2256 976 -2255
rect 58 -2258 59 -2257
rect 415 -2258 416 -2257
rect 443 -2258 444 -2257
rect 457 -2258 458 -2257
rect 471 -2258 472 -2257
rect 611 -2258 612 -2257
rect 849 -2258 850 -2257
rect 898 -2258 899 -2257
rect 912 -2258 913 -2257
rect 933 -2258 934 -2257
rect 16 -2260 17 -2259
rect 58 -2260 59 -2259
rect 254 -2260 255 -2259
rect 369 -2260 370 -2259
rect 443 -2260 444 -2259
rect 674 -2260 675 -2259
rect 877 -2260 878 -2259
rect 926 -2260 927 -2259
rect 261 -2262 262 -2261
rect 310 -2262 311 -2261
rect 478 -2262 479 -2261
rect 674 -2262 675 -2261
rect 233 -2264 234 -2263
rect 261 -2264 262 -2263
rect 478 -2264 479 -2263
rect 492 -2264 493 -2263
rect 534 -2264 535 -2263
rect 898 -2264 899 -2263
rect 233 -2266 234 -2265
rect 523 -2266 524 -2265
rect 611 -2266 612 -2265
rect 660 -2266 661 -2265
rect 502 -2268 503 -2267
rect 534 -2268 535 -2267
rect 660 -2268 661 -2267
rect 751 -2268 752 -2267
rect 751 -2270 752 -2269
rect 807 -2270 808 -2269
rect 807 -2272 808 -2271
rect 947 -2272 948 -2271
rect 947 -2274 948 -2273
rect 954 -2274 955 -2273
rect 464 -2276 465 -2275
rect 954 -2276 955 -2275
rect 2 -2287 3 -2286
rect 51 -2287 52 -2286
rect 58 -2287 59 -2286
rect 275 -2287 276 -2286
rect 303 -2287 304 -2286
rect 478 -2287 479 -2286
rect 481 -2287 482 -2286
rect 891 -2287 892 -2286
rect 905 -2287 906 -2286
rect 933 -2287 934 -2286
rect 2 -2289 3 -2288
rect 30 -2289 31 -2288
rect 44 -2289 45 -2288
rect 54 -2289 55 -2288
rect 58 -2289 59 -2288
rect 436 -2289 437 -2288
rect 450 -2289 451 -2288
rect 467 -2289 468 -2288
rect 499 -2289 500 -2288
rect 611 -2289 612 -2288
rect 642 -2289 643 -2288
rect 800 -2289 801 -2288
rect 877 -2289 878 -2288
rect 891 -2289 892 -2288
rect 908 -2289 909 -2288
rect 947 -2289 948 -2288
rect 9 -2291 10 -2290
rect 128 -2291 129 -2290
rect 191 -2291 192 -2290
rect 212 -2291 213 -2290
rect 226 -2291 227 -2290
rect 345 -2291 346 -2290
rect 376 -2291 377 -2290
rect 646 -2291 647 -2290
rect 684 -2291 685 -2290
rect 835 -2291 836 -2290
rect 877 -2291 878 -2290
rect 954 -2291 955 -2290
rect 12 -2293 13 -2292
rect 215 -2293 216 -2292
rect 268 -2293 269 -2292
rect 488 -2293 489 -2292
rect 502 -2293 503 -2292
rect 723 -2293 724 -2292
rect 765 -2293 766 -2292
rect 828 -2293 829 -2292
rect 884 -2293 885 -2292
rect 912 -2293 913 -2292
rect 922 -2293 923 -2292
rect 929 -2293 930 -2292
rect 947 -2293 948 -2292
rect 961 -2293 962 -2292
rect 16 -2295 17 -2294
rect 485 -2295 486 -2294
rect 534 -2295 535 -2294
rect 565 -2295 566 -2294
rect 576 -2295 577 -2294
rect 856 -2295 857 -2294
rect 926 -2295 927 -2294
rect 975 -2295 976 -2294
rect 16 -2297 17 -2296
rect 233 -2297 234 -2296
rect 268 -2297 269 -2296
rect 296 -2297 297 -2296
rect 303 -2297 304 -2296
rect 415 -2297 416 -2296
rect 436 -2297 437 -2296
rect 457 -2297 458 -2296
rect 464 -2297 465 -2296
rect 562 -2297 563 -2296
rect 583 -2297 584 -2296
rect 660 -2297 661 -2296
rect 723 -2297 724 -2296
rect 821 -2297 822 -2296
rect 842 -2297 843 -2296
rect 884 -2297 885 -2296
rect 23 -2299 24 -2298
rect 51 -2299 52 -2298
rect 61 -2299 62 -2298
rect 705 -2299 706 -2298
rect 768 -2299 769 -2298
rect 849 -2299 850 -2298
rect 856 -2299 857 -2298
rect 898 -2299 899 -2298
rect 23 -2301 24 -2300
rect 282 -2301 283 -2300
rect 296 -2301 297 -2300
rect 464 -2301 465 -2300
rect 467 -2301 468 -2300
rect 471 -2301 472 -2300
rect 520 -2301 521 -2300
rect 576 -2301 577 -2300
rect 597 -2301 598 -2300
rect 646 -2301 647 -2300
rect 779 -2301 780 -2300
rect 828 -2301 829 -2300
rect 849 -2301 850 -2300
rect 901 -2301 902 -2300
rect 30 -2303 31 -2302
rect 229 -2303 230 -2302
rect 233 -2303 234 -2302
rect 261 -2303 262 -2302
rect 275 -2303 276 -2302
rect 362 -2303 363 -2302
rect 373 -2303 374 -2302
rect 485 -2303 486 -2302
rect 562 -2303 563 -2302
rect 758 -2303 759 -2302
rect 786 -2303 787 -2302
rect 821 -2303 822 -2302
rect 44 -2305 45 -2304
rect 779 -2305 780 -2304
rect 793 -2305 794 -2304
rect 842 -2305 843 -2304
rect 47 -2307 48 -2306
rect 131 -2307 132 -2306
rect 163 -2307 164 -2306
rect 191 -2307 192 -2306
rect 261 -2307 262 -2306
rect 289 -2307 290 -2306
rect 310 -2307 311 -2306
rect 334 -2307 335 -2306
rect 341 -2307 342 -2306
rect 716 -2307 717 -2306
rect 793 -2307 794 -2306
rect 863 -2307 864 -2306
rect 65 -2309 66 -2308
rect 310 -2309 311 -2308
rect 313 -2309 314 -2308
rect 786 -2309 787 -2308
rect 800 -2309 801 -2308
rect 814 -2309 815 -2308
rect 65 -2311 66 -2310
rect 100 -2311 101 -2310
rect 107 -2311 108 -2310
rect 625 -2311 626 -2310
rect 667 -2311 668 -2310
rect 814 -2311 815 -2310
rect 72 -2313 73 -2312
rect 177 -2313 178 -2312
rect 282 -2313 283 -2312
rect 408 -2313 409 -2312
rect 415 -2313 416 -2312
rect 716 -2313 717 -2312
rect 72 -2315 73 -2314
rect 79 -2315 80 -2314
rect 82 -2315 83 -2314
rect 86 -2315 87 -2314
rect 93 -2315 94 -2314
rect 103 -2315 104 -2314
rect 107 -2315 108 -2314
rect 110 -2315 111 -2314
rect 114 -2315 115 -2314
rect 198 -2315 199 -2314
rect 289 -2315 290 -2314
rect 338 -2315 339 -2314
rect 355 -2315 356 -2314
rect 471 -2315 472 -2314
rect 537 -2315 538 -2314
rect 758 -2315 759 -2314
rect 79 -2317 80 -2316
rect 149 -2317 150 -2316
rect 163 -2317 164 -2316
rect 338 -2317 339 -2316
rect 355 -2317 356 -2316
rect 660 -2317 661 -2316
rect 681 -2317 682 -2316
rect 863 -2317 864 -2316
rect 86 -2319 87 -2318
rect 541 -2319 542 -2318
rect 586 -2319 587 -2318
rect 667 -2319 668 -2318
rect 93 -2321 94 -2320
rect 523 -2321 524 -2320
rect 597 -2321 598 -2320
rect 604 -2321 605 -2320
rect 611 -2321 612 -2320
rect 632 -2321 633 -2320
rect 100 -2323 101 -2322
rect 422 -2323 423 -2322
rect 450 -2323 451 -2322
rect 730 -2323 731 -2322
rect 114 -2325 115 -2324
rect 135 -2325 136 -2324
rect 149 -2325 150 -2324
rect 184 -2325 185 -2324
rect 198 -2325 199 -2324
rect 205 -2325 206 -2324
rect 317 -2325 318 -2324
rect 397 -2325 398 -2324
rect 401 -2325 402 -2324
rect 541 -2325 542 -2324
rect 625 -2325 626 -2324
rect 688 -2325 689 -2324
rect 54 -2327 55 -2326
rect 135 -2327 136 -2326
rect 142 -2327 143 -2326
rect 184 -2327 185 -2326
rect 205 -2327 206 -2326
rect 348 -2327 349 -2326
rect 359 -2327 360 -2326
rect 730 -2327 731 -2326
rect 128 -2329 129 -2328
rect 240 -2329 241 -2328
rect 317 -2329 318 -2328
rect 674 -2329 675 -2328
rect 688 -2329 689 -2328
rect 695 -2329 696 -2328
rect 142 -2331 143 -2330
rect 156 -2331 157 -2330
rect 177 -2331 178 -2330
rect 247 -2331 248 -2330
rect 324 -2331 325 -2330
rect 443 -2331 444 -2330
rect 513 -2331 514 -2330
rect 632 -2331 633 -2330
rect 674 -2331 675 -2330
rect 709 -2331 710 -2330
rect 37 -2333 38 -2332
rect 156 -2333 157 -2332
rect 180 -2333 181 -2332
rect 695 -2333 696 -2332
rect 702 -2333 703 -2332
rect 709 -2333 710 -2332
rect 37 -2335 38 -2334
rect 110 -2335 111 -2334
rect 121 -2335 122 -2334
rect 247 -2335 248 -2334
rect 254 -2335 255 -2334
rect 513 -2335 514 -2334
rect 702 -2335 703 -2334
rect 751 -2335 752 -2334
rect 121 -2337 122 -2336
rect 292 -2337 293 -2336
rect 359 -2337 360 -2336
rect 394 -2337 395 -2336
rect 401 -2337 402 -2336
rect 653 -2337 654 -2336
rect 737 -2337 738 -2336
rect 751 -2337 752 -2336
rect 240 -2339 241 -2338
rect 527 -2339 528 -2338
rect 737 -2339 738 -2338
rect 744 -2339 745 -2338
rect 254 -2341 255 -2340
rect 579 -2341 580 -2340
rect 744 -2341 745 -2340
rect 772 -2341 773 -2340
rect 352 -2343 353 -2342
rect 527 -2343 528 -2342
rect 772 -2343 773 -2342
rect 870 -2343 871 -2342
rect 366 -2345 367 -2344
rect 604 -2345 605 -2344
rect 870 -2345 871 -2344
rect 940 -2345 941 -2344
rect 170 -2347 171 -2346
rect 366 -2347 367 -2346
rect 380 -2347 381 -2346
rect 681 -2347 682 -2346
rect 159 -2349 160 -2348
rect 170 -2349 171 -2348
rect 331 -2349 332 -2348
rect 380 -2349 381 -2348
rect 383 -2349 384 -2348
rect 408 -2349 409 -2348
rect 422 -2349 423 -2348
rect 429 -2349 430 -2348
rect 443 -2349 444 -2348
rect 548 -2349 549 -2348
rect 373 -2351 374 -2350
rect 429 -2351 430 -2350
rect 492 -2351 493 -2350
rect 653 -2351 654 -2350
rect 394 -2353 395 -2352
rect 835 -2353 836 -2352
rect 492 -2355 493 -2354
rect 555 -2355 556 -2354
rect 548 -2357 549 -2356
rect 590 -2357 591 -2356
rect 544 -2359 545 -2358
rect 590 -2359 591 -2358
rect 555 -2361 556 -2360
rect 807 -2361 808 -2360
rect 583 -2363 584 -2362
rect 807 -2363 808 -2362
rect 16 -2374 17 -2373
rect 138 -2374 139 -2373
rect 156 -2374 157 -2373
rect 215 -2374 216 -2373
rect 226 -2374 227 -2373
rect 667 -2374 668 -2373
rect 702 -2374 703 -2373
rect 709 -2374 710 -2373
rect 726 -2374 727 -2373
rect 821 -2374 822 -2373
rect 940 -2374 941 -2373
rect 947 -2374 948 -2373
rect 23 -2376 24 -2375
rect 219 -2376 220 -2375
rect 240 -2376 241 -2375
rect 558 -2376 559 -2375
rect 569 -2376 570 -2375
rect 667 -2376 668 -2375
rect 709 -2376 710 -2375
rect 765 -2376 766 -2375
rect 772 -2376 773 -2375
rect 828 -2376 829 -2375
rect 30 -2378 31 -2377
rect 156 -2378 157 -2377
rect 177 -2378 178 -2377
rect 226 -2378 227 -2377
rect 233 -2378 234 -2377
rect 240 -2378 241 -2377
rect 247 -2378 248 -2377
rect 352 -2378 353 -2377
rect 376 -2378 377 -2377
rect 758 -2378 759 -2377
rect 761 -2378 762 -2377
rect 842 -2378 843 -2377
rect 2 -2380 3 -2379
rect 30 -2380 31 -2379
rect 44 -2380 45 -2379
rect 61 -2380 62 -2379
rect 93 -2380 94 -2379
rect 208 -2380 209 -2379
rect 212 -2380 213 -2379
rect 373 -2380 374 -2379
rect 404 -2380 405 -2379
rect 779 -2380 780 -2379
rect 828 -2380 829 -2379
rect 877 -2380 878 -2379
rect 37 -2382 38 -2381
rect 93 -2382 94 -2381
rect 100 -2382 101 -2381
rect 359 -2382 360 -2381
rect 411 -2382 412 -2381
rect 436 -2382 437 -2381
rect 457 -2382 458 -2381
rect 576 -2382 577 -2381
rect 583 -2382 584 -2381
rect 660 -2382 661 -2381
rect 723 -2382 724 -2381
rect 765 -2382 766 -2381
rect 772 -2382 773 -2381
rect 793 -2382 794 -2381
rect 51 -2384 52 -2383
rect 730 -2384 731 -2383
rect 751 -2384 752 -2383
rect 754 -2384 755 -2383
rect 100 -2386 101 -2385
rect 149 -2386 150 -2385
rect 177 -2386 178 -2385
rect 254 -2386 255 -2385
rect 268 -2386 269 -2385
rect 289 -2386 290 -2385
rect 303 -2386 304 -2385
rect 418 -2386 419 -2385
rect 460 -2386 461 -2385
rect 506 -2386 507 -2385
rect 520 -2386 521 -2385
rect 548 -2386 549 -2385
rect 555 -2386 556 -2385
rect 625 -2386 626 -2385
rect 639 -2386 640 -2385
rect 688 -2386 689 -2385
rect 723 -2386 724 -2385
rect 849 -2386 850 -2385
rect 107 -2388 108 -2387
rect 450 -2388 451 -2387
rect 464 -2388 465 -2387
rect 506 -2388 507 -2387
rect 523 -2388 524 -2387
rect 611 -2388 612 -2387
rect 618 -2388 619 -2387
rect 628 -2388 629 -2387
rect 639 -2388 640 -2387
rect 835 -2388 836 -2387
rect 107 -2390 108 -2389
rect 149 -2390 150 -2389
rect 163 -2390 164 -2389
rect 289 -2390 290 -2389
rect 310 -2390 311 -2389
rect 604 -2390 605 -2389
rect 611 -2390 612 -2389
rect 674 -2390 675 -2389
rect 114 -2392 115 -2391
rect 152 -2392 153 -2391
rect 163 -2392 164 -2391
rect 184 -2392 185 -2391
rect 205 -2392 206 -2391
rect 247 -2392 248 -2391
rect 275 -2392 276 -2391
rect 397 -2392 398 -2391
rect 408 -2392 409 -2391
rect 436 -2392 437 -2391
rect 450 -2392 451 -2391
rect 471 -2392 472 -2391
rect 481 -2392 482 -2391
rect 716 -2392 717 -2391
rect 114 -2394 115 -2393
rect 170 -2394 171 -2393
rect 184 -2394 185 -2393
rect 222 -2394 223 -2393
rect 233 -2394 234 -2393
rect 387 -2394 388 -2393
rect 408 -2394 409 -2393
rect 646 -2394 647 -2393
rect 660 -2394 661 -2393
rect 737 -2394 738 -2393
rect 121 -2396 122 -2395
rect 271 -2396 272 -2395
rect 275 -2396 276 -2395
rect 422 -2396 423 -2395
rect 464 -2396 465 -2395
rect 814 -2396 815 -2395
rect 65 -2398 66 -2397
rect 121 -2398 122 -2397
rect 135 -2398 136 -2397
rect 303 -2398 304 -2397
rect 310 -2398 311 -2397
rect 355 -2398 356 -2397
rect 380 -2398 381 -2397
rect 604 -2398 605 -2397
rect 618 -2398 619 -2397
rect 695 -2398 696 -2397
rect 716 -2398 717 -2397
rect 807 -2398 808 -2397
rect 170 -2400 171 -2399
rect 191 -2400 192 -2399
rect 219 -2400 220 -2399
rect 548 -2400 549 -2399
rect 551 -2400 552 -2399
rect 646 -2400 647 -2399
rect 674 -2400 675 -2399
rect 786 -2400 787 -2399
rect 807 -2400 808 -2399
rect 863 -2400 864 -2399
rect 191 -2402 192 -2401
rect 198 -2402 199 -2401
rect 282 -2402 283 -2401
rect 457 -2402 458 -2401
rect 471 -2402 472 -2401
rect 562 -2402 563 -2401
rect 737 -2402 738 -2401
rect 744 -2402 745 -2401
rect 128 -2404 129 -2403
rect 282 -2404 283 -2403
rect 313 -2404 314 -2403
rect 541 -2404 542 -2403
rect 744 -2404 745 -2403
rect 856 -2404 857 -2403
rect 128 -2406 129 -2405
rect 296 -2406 297 -2405
rect 324 -2406 325 -2405
rect 341 -2406 342 -2405
rect 345 -2406 346 -2405
rect 422 -2406 423 -2405
rect 527 -2406 528 -2405
rect 569 -2406 570 -2405
rect 79 -2408 80 -2407
rect 296 -2408 297 -2407
rect 317 -2408 318 -2407
rect 345 -2408 346 -2407
rect 527 -2408 528 -2407
rect 590 -2408 591 -2407
rect 58 -2410 59 -2409
rect 79 -2410 80 -2409
rect 198 -2410 199 -2409
rect 222 -2410 223 -2409
rect 317 -2410 318 -2409
rect 544 -2410 545 -2409
rect 58 -2412 59 -2411
rect 65 -2412 66 -2411
rect 324 -2412 325 -2411
rect 415 -2412 416 -2411
rect 534 -2412 535 -2411
rect 597 -2412 598 -2411
rect 331 -2414 332 -2413
rect 380 -2414 381 -2413
rect 415 -2414 416 -2413
rect 429 -2414 430 -2413
rect 499 -2414 500 -2413
rect 534 -2414 535 -2413
rect 597 -2414 598 -2413
rect 681 -2414 682 -2413
rect 331 -2416 332 -2415
rect 366 -2416 367 -2415
rect 429 -2416 430 -2415
rect 590 -2416 591 -2415
rect 653 -2416 654 -2415
rect 681 -2416 682 -2415
rect 334 -2418 335 -2417
rect 387 -2418 388 -2417
rect 401 -2418 402 -2417
rect 653 -2418 654 -2417
rect 254 -2420 255 -2419
rect 334 -2420 335 -2419
rect 338 -2420 339 -2419
rect 513 -2420 514 -2419
rect 366 -2422 367 -2421
rect 485 -2422 486 -2421
rect 499 -2422 500 -2421
rect 632 -2422 633 -2421
rect 401 -2424 402 -2423
rect 492 -2424 493 -2423
rect 513 -2424 514 -2423
rect 565 -2424 566 -2423
rect 443 -2426 444 -2425
rect 492 -2426 493 -2425
rect 394 -2428 395 -2427
rect 443 -2428 444 -2427
rect 488 -2428 489 -2427
rect 632 -2428 633 -2427
rect 65 -2439 66 -2438
rect 72 -2439 73 -2438
rect 79 -2439 80 -2438
rect 264 -2439 265 -2438
rect 268 -2439 269 -2438
rect 408 -2439 409 -2438
rect 422 -2439 423 -2438
rect 464 -2439 465 -2438
rect 471 -2439 472 -2438
rect 583 -2439 584 -2438
rect 590 -2439 591 -2438
rect 593 -2439 594 -2438
rect 625 -2439 626 -2438
rect 716 -2439 717 -2438
rect 730 -2439 731 -2438
rect 737 -2439 738 -2438
rect 754 -2439 755 -2438
rect 807 -2439 808 -2438
rect 926 -2439 927 -2438
rect 933 -2439 934 -2438
rect 93 -2441 94 -2440
rect 131 -2441 132 -2440
rect 135 -2441 136 -2440
rect 142 -2441 143 -2440
rect 170 -2441 171 -2440
rect 215 -2441 216 -2440
rect 233 -2441 234 -2440
rect 369 -2441 370 -2440
rect 401 -2441 402 -2440
rect 471 -2441 472 -2440
rect 474 -2441 475 -2440
rect 481 -2441 482 -2440
rect 485 -2441 486 -2440
rect 604 -2441 605 -2440
rect 625 -2441 626 -2440
rect 660 -2441 661 -2440
rect 681 -2441 682 -2440
rect 688 -2441 689 -2440
rect 695 -2441 696 -2440
rect 702 -2441 703 -2440
rect 716 -2441 717 -2440
rect 726 -2441 727 -2440
rect 730 -2441 731 -2440
rect 733 -2441 734 -2440
rect 779 -2441 780 -2440
rect 828 -2441 829 -2440
rect 100 -2443 101 -2442
rect 156 -2443 157 -2442
rect 191 -2443 192 -2442
rect 208 -2443 209 -2442
rect 240 -2443 241 -2442
rect 257 -2443 258 -2442
rect 275 -2443 276 -2442
rect 331 -2443 332 -2442
rect 334 -2443 335 -2442
rect 390 -2443 391 -2442
rect 408 -2443 409 -2442
rect 415 -2443 416 -2442
rect 422 -2443 423 -2442
rect 478 -2443 479 -2442
rect 502 -2443 503 -2442
rect 569 -2443 570 -2442
rect 576 -2443 577 -2442
rect 653 -2443 654 -2442
rect 660 -2443 661 -2442
rect 667 -2443 668 -2442
rect 681 -2443 682 -2442
rect 709 -2443 710 -2442
rect 100 -2445 101 -2444
rect 117 -2445 118 -2444
rect 121 -2445 122 -2444
rect 219 -2445 220 -2444
rect 226 -2445 227 -2444
rect 275 -2445 276 -2444
rect 296 -2445 297 -2444
rect 597 -2445 598 -2444
rect 604 -2445 605 -2444
rect 611 -2445 612 -2444
rect 642 -2445 643 -2444
rect 646 -2445 647 -2444
rect 709 -2445 710 -2444
rect 744 -2445 745 -2444
rect 107 -2447 108 -2446
rect 121 -2447 122 -2446
rect 128 -2447 129 -2446
rect 219 -2447 220 -2446
rect 226 -2447 227 -2446
rect 261 -2447 262 -2446
rect 310 -2447 311 -2446
rect 488 -2447 489 -2446
rect 506 -2447 507 -2446
rect 600 -2447 601 -2446
rect 611 -2447 612 -2446
rect 632 -2447 633 -2446
rect 114 -2449 115 -2448
rect 233 -2449 234 -2448
rect 254 -2449 255 -2448
rect 268 -2449 269 -2448
rect 317 -2449 318 -2448
rect 432 -2449 433 -2448
rect 443 -2449 444 -2448
rect 478 -2449 479 -2448
rect 499 -2449 500 -2448
rect 506 -2449 507 -2448
rect 513 -2449 514 -2448
rect 579 -2449 580 -2448
rect 107 -2451 108 -2450
rect 114 -2451 115 -2450
rect 149 -2451 150 -2450
rect 170 -2451 171 -2450
rect 191 -2451 192 -2450
rect 198 -2451 199 -2450
rect 222 -2451 223 -2450
rect 310 -2451 311 -2450
rect 345 -2451 346 -2450
rect 401 -2451 402 -2450
rect 443 -2451 444 -2450
rect 450 -2451 451 -2450
rect 457 -2451 458 -2450
rect 492 -2451 493 -2450
rect 513 -2451 514 -2450
rect 534 -2451 535 -2450
rect 541 -2451 542 -2450
rect 562 -2451 563 -2450
rect 569 -2451 570 -2450
rect 618 -2451 619 -2450
rect 86 -2453 87 -2452
rect 450 -2453 451 -2452
rect 460 -2453 461 -2452
rect 520 -2453 521 -2452
rect 527 -2453 528 -2452
rect 551 -2453 552 -2452
rect 555 -2453 556 -2452
rect 576 -2453 577 -2452
rect 152 -2455 153 -2454
rect 198 -2455 199 -2454
rect 282 -2455 283 -2454
rect 317 -2455 318 -2454
rect 331 -2455 332 -2454
rect 345 -2455 346 -2454
rect 348 -2455 349 -2454
rect 387 -2455 388 -2454
rect 534 -2455 535 -2454
rect 674 -2455 675 -2454
rect 163 -2457 164 -2456
rect 240 -2457 241 -2456
rect 289 -2457 290 -2456
rect 432 -2457 433 -2456
rect 548 -2457 549 -2456
rect 639 -2457 640 -2456
rect 674 -2457 675 -2456
rect 758 -2457 759 -2456
rect 163 -2459 164 -2458
rect 184 -2459 185 -2458
rect 212 -2459 213 -2458
rect 282 -2459 283 -2458
rect 352 -2459 353 -2458
rect 394 -2459 395 -2458
rect 639 -2459 640 -2458
rect 723 -2459 724 -2458
rect 737 -2459 738 -2458
rect 758 -2459 759 -2458
rect 184 -2461 185 -2460
rect 205 -2461 206 -2460
rect 247 -2461 248 -2460
rect 289 -2461 290 -2460
rect 324 -2461 325 -2460
rect 352 -2461 353 -2460
rect 359 -2461 360 -2460
rect 467 -2461 468 -2460
rect 723 -2461 724 -2460
rect 761 -2461 762 -2460
rect 177 -2463 178 -2462
rect 247 -2463 248 -2462
rect 338 -2463 339 -2462
rect 359 -2463 360 -2462
rect 366 -2463 367 -2462
rect 415 -2463 416 -2462
rect 761 -2463 762 -2462
rect 772 -2463 773 -2462
rect 159 -2465 160 -2464
rect 177 -2465 178 -2464
rect 299 -2465 300 -2464
rect 338 -2465 339 -2464
rect 387 -2465 388 -2464
rect 436 -2465 437 -2464
rect 380 -2467 381 -2466
rect 436 -2467 437 -2466
rect 373 -2469 374 -2468
rect 380 -2469 381 -2468
rect 394 -2469 395 -2468
rect 397 -2469 398 -2468
rect 65 -2480 66 -2479
rect 72 -2480 73 -2479
rect 86 -2480 87 -2479
rect 96 -2480 97 -2479
rect 100 -2480 101 -2479
rect 110 -2480 111 -2479
rect 114 -2480 115 -2479
rect 121 -2480 122 -2479
rect 131 -2480 132 -2479
rect 135 -2480 136 -2479
rect 142 -2480 143 -2479
rect 170 -2480 171 -2479
rect 177 -2480 178 -2479
rect 187 -2480 188 -2479
rect 198 -2480 199 -2479
rect 212 -2480 213 -2479
rect 219 -2480 220 -2479
rect 254 -2480 255 -2479
rect 282 -2480 283 -2479
rect 362 -2480 363 -2479
rect 376 -2480 377 -2479
rect 422 -2480 423 -2479
rect 432 -2480 433 -2479
rect 457 -2480 458 -2479
rect 467 -2480 468 -2479
rect 478 -2480 479 -2479
rect 502 -2480 503 -2479
rect 513 -2480 514 -2479
rect 523 -2480 524 -2479
rect 541 -2480 542 -2479
rect 576 -2480 577 -2479
rect 586 -2480 587 -2479
rect 590 -2480 591 -2479
rect 625 -2480 626 -2479
rect 667 -2480 668 -2479
rect 681 -2480 682 -2479
rect 744 -2480 745 -2479
rect 751 -2480 752 -2479
rect 758 -2480 759 -2479
rect 765 -2480 766 -2479
rect 933 -2480 934 -2479
rect 936 -2480 937 -2479
rect 940 -2480 941 -2479
rect 947 -2480 948 -2479
rect 100 -2482 101 -2481
rect 121 -2482 122 -2481
rect 138 -2482 139 -2481
rect 219 -2482 220 -2481
rect 226 -2482 227 -2481
rect 229 -2482 230 -2481
rect 247 -2482 248 -2481
rect 324 -2482 325 -2481
rect 338 -2482 339 -2481
rect 404 -2482 405 -2481
rect 450 -2482 451 -2481
rect 548 -2482 549 -2481
rect 597 -2482 598 -2481
rect 674 -2482 675 -2481
rect 681 -2482 682 -2481
rect 688 -2482 689 -2481
rect 758 -2482 759 -2481
rect 761 -2482 762 -2481
rect 107 -2484 108 -2483
rect 114 -2484 115 -2483
rect 149 -2484 150 -2483
rect 163 -2484 164 -2483
rect 177 -2484 178 -2483
rect 191 -2484 192 -2483
rect 226 -2484 227 -2483
rect 261 -2484 262 -2483
rect 275 -2484 276 -2483
rect 324 -2484 325 -2483
rect 359 -2484 360 -2483
rect 373 -2484 374 -2483
rect 401 -2484 402 -2483
rect 422 -2484 423 -2483
rect 443 -2484 444 -2483
rect 450 -2484 451 -2483
rect 471 -2484 472 -2483
rect 527 -2484 528 -2483
rect 688 -2484 689 -2483
rect 695 -2484 696 -2483
rect 159 -2486 160 -2485
rect 170 -2486 171 -2485
rect 233 -2486 234 -2485
rect 261 -2486 262 -2485
rect 271 -2486 272 -2485
rect 275 -2486 276 -2485
rect 296 -2486 297 -2485
rect 303 -2486 304 -2485
rect 310 -2486 311 -2485
rect 366 -2486 367 -2485
rect 401 -2486 402 -2485
rect 537 -2486 538 -2485
rect 695 -2486 696 -2485
rect 709 -2486 710 -2485
rect 229 -2488 230 -2487
rect 233 -2488 234 -2487
rect 236 -2488 237 -2487
rect 310 -2488 311 -2487
rect 359 -2488 360 -2487
rect 408 -2488 409 -2487
rect 415 -2488 416 -2487
rect 443 -2488 444 -2487
rect 506 -2488 507 -2487
rect 520 -2488 521 -2487
rect 523 -2488 524 -2487
rect 527 -2488 528 -2487
rect 709 -2488 710 -2487
rect 716 -2488 717 -2487
rect 240 -2490 241 -2489
rect 296 -2490 297 -2489
rect 303 -2490 304 -2489
rect 331 -2490 332 -2489
rect 408 -2490 409 -2489
rect 436 -2490 437 -2489
rect 520 -2490 521 -2489
rect 569 -2490 570 -2489
rect 716 -2490 717 -2489
rect 723 -2490 724 -2489
rect 247 -2492 248 -2491
rect 268 -2492 269 -2491
rect 317 -2492 318 -2491
rect 331 -2492 332 -2491
rect 723 -2492 724 -2491
rect 737 -2492 738 -2491
rect 289 -2494 290 -2493
rect 317 -2494 318 -2493
rect 201 -2496 202 -2495
rect 289 -2496 290 -2495
rect 5 -2507 6 -2506
rect 9 -2507 10 -2506
rect 86 -2507 87 -2506
rect 103 -2507 104 -2506
rect 107 -2507 108 -2506
rect 121 -2507 122 -2506
rect 142 -2507 143 -2506
rect 194 -2507 195 -2506
rect 201 -2507 202 -2506
rect 205 -2507 206 -2506
rect 219 -2507 220 -2506
rect 240 -2507 241 -2506
rect 247 -2507 248 -2506
rect 271 -2507 272 -2506
rect 275 -2507 276 -2506
rect 282 -2507 283 -2506
rect 285 -2507 286 -2506
rect 317 -2507 318 -2506
rect 331 -2507 332 -2506
rect 345 -2507 346 -2506
rect 352 -2507 353 -2506
rect 362 -2507 363 -2506
rect 380 -2507 381 -2506
rect 383 -2507 384 -2506
rect 387 -2507 388 -2506
rect 408 -2507 409 -2506
rect 450 -2507 451 -2506
rect 457 -2507 458 -2506
rect 523 -2507 524 -2506
rect 527 -2507 528 -2506
rect 597 -2507 598 -2506
rect 604 -2507 605 -2506
rect 660 -2507 661 -2506
rect 663 -2507 664 -2506
rect 681 -2507 682 -2506
rect 702 -2507 703 -2506
rect 709 -2507 710 -2506
rect 712 -2507 713 -2506
rect 723 -2507 724 -2506
rect 730 -2507 731 -2506
rect 740 -2507 741 -2506
rect 751 -2507 752 -2506
rect 887 -2507 888 -2506
rect 891 -2507 892 -2506
rect 933 -2507 934 -2506
rect 940 -2507 941 -2506
rect 943 -2507 944 -2506
rect 947 -2507 948 -2506
rect 100 -2509 101 -2508
rect 107 -2509 108 -2508
rect 114 -2509 115 -2508
rect 117 -2509 118 -2508
rect 149 -2509 150 -2508
rect 166 -2509 167 -2508
rect 184 -2509 185 -2508
rect 187 -2509 188 -2508
rect 191 -2509 192 -2508
rect 226 -2509 227 -2508
rect 229 -2509 230 -2508
rect 233 -2509 234 -2508
rect 254 -2509 255 -2508
rect 278 -2509 279 -2508
rect 289 -2509 290 -2508
rect 303 -2509 304 -2508
rect 394 -2509 395 -2508
rect 397 -2509 398 -2508
rect 404 -2509 405 -2508
rect 418 -2509 419 -2508
rect 443 -2509 444 -2508
rect 450 -2509 451 -2508
rect 604 -2509 605 -2508
rect 611 -2509 612 -2508
rect 695 -2509 696 -2508
rect 705 -2509 706 -2508
rect 744 -2509 745 -2508
rect 758 -2509 759 -2508
rect 156 -2511 157 -2510
rect 159 -2511 160 -2510
rect 163 -2511 164 -2510
rect 170 -2511 171 -2510
rect 177 -2511 178 -2510
rect 191 -2511 192 -2510
rect 212 -2511 213 -2510
rect 226 -2511 227 -2510
rect 261 -2511 262 -2510
rect 268 -2511 269 -2510
rect 296 -2511 297 -2510
rect 310 -2511 311 -2510
rect 401 -2511 402 -2510
rect 404 -2511 405 -2510
rect 163 -2513 164 -2512
rect 180 -2513 181 -2512
rect 299 -2513 300 -2512
rect 341 -2513 342 -2512
rect 310 -2515 311 -2514
rect 324 -2515 325 -2514
rect 5 -2526 6 -2525
rect 9 -2526 10 -2525
rect 100 -2526 101 -2525
rect 107 -2526 108 -2525
rect 114 -2526 115 -2525
rect 124 -2526 125 -2525
rect 163 -2526 164 -2525
rect 170 -2526 171 -2525
rect 180 -2526 181 -2525
rect 184 -2526 185 -2525
rect 191 -2526 192 -2525
rect 198 -2526 199 -2525
rect 292 -2526 293 -2525
rect 296 -2526 297 -2525
rect 303 -2526 304 -2525
rect 310 -2526 311 -2525
rect 341 -2526 342 -2525
rect 345 -2526 346 -2525
rect 450 -2526 451 -2525
rect 457 -2526 458 -2525
rect 597 -2526 598 -2525
rect 604 -2526 605 -2525
rect 663 -2526 664 -2525
rect 667 -2526 668 -2525
rect 716 -2526 717 -2525
rect 723 -2526 724 -2525
rect 730 -2526 731 -2525
rect 740 -2526 741 -2525
rect 121 -2528 122 -2527
rect 131 -2528 132 -2527
<< metal2 >>
rect 93 -3 94 1
rect 100 -3 101 1
rect 107 -3 108 1
rect 128 -3 129 1
rect 205 -3 206 1
rect 212 -3 213 1
rect 215 -3 216 1
rect 236 -3 237 1
rect 240 -3 241 1
rect 247 -3 248 1
rect 261 -3 262 1
rect 268 -3 269 1
rect 324 -3 325 1
rect 334 -3 335 1
rect 429 -3 430 1
rect 450 -3 451 1
rect 464 -3 465 1
rect 488 -3 489 1
rect 530 -3 531 1
rect 534 -3 535 1
rect 583 -3 584 1
rect 597 -3 598 1
rect 660 -3 661 1
rect 667 -3 668 1
rect 117 -3 118 -1
rect 121 -3 122 -1
rect 226 -3 227 -1
rect 233 -3 234 -1
rect 86 -13 87 -11
rect 103 -22 104 -12
rect 117 -22 118 -12
rect 128 -13 129 -11
rect 135 -22 136 -12
rect 145 -13 146 -11
rect 173 -22 174 -12
rect 198 -22 199 -12
rect 205 -13 206 -11
rect 215 -22 216 -12
rect 226 -13 227 -11
rect 250 -13 251 -11
rect 254 -22 255 -12
rect 268 -13 269 -11
rect 289 -22 290 -12
rect 306 -22 307 -12
rect 310 -22 311 -12
rect 324 -13 325 -11
rect 348 -22 349 -12
rect 359 -22 360 -12
rect 373 -22 374 -12
rect 446 -22 447 -12
rect 450 -13 451 -11
rect 464 -13 465 -11
rect 485 -13 486 -11
rect 527 -22 528 -12
rect 534 -13 535 -11
rect 541 -22 542 -12
rect 548 -13 549 -11
rect 569 -22 570 -12
rect 590 -13 591 -11
rect 604 -22 605 -12
rect 607 -13 608 -11
rect 618 -22 619 -12
rect 667 -13 668 -11
rect 674 -22 675 -12
rect 89 -15 90 -11
rect 100 -15 101 -11
rect 177 -22 178 -14
rect 212 -22 213 -14
rect 219 -15 220 -11
rect 226 -22 227 -14
rect 233 -22 234 -14
rect 247 -22 248 -14
rect 257 -15 258 -11
rect 275 -22 276 -14
rect 317 -22 318 -14
rect 331 -22 332 -14
rect 415 -22 416 -14
rect 429 -15 430 -11
rect 453 -22 454 -14
rect 471 -22 472 -14
rect 492 -22 493 -14
rect 513 -22 514 -14
rect 562 -22 563 -14
rect 576 -22 577 -14
rect 597 -15 598 -11
rect 611 -22 612 -14
rect 93 -17 94 -11
rect 107 -17 108 -11
rect 184 -22 185 -16
rect 205 -22 206 -16
rect 219 -22 220 -16
rect 222 -17 223 -11
rect 240 -17 241 -11
rect 240 -22 241 -16
rect 240 -17 241 -11
rect 240 -22 241 -16
rect 261 -22 262 -16
rect 282 -17 283 -11
rect 324 -22 325 -16
rect 341 -17 342 -11
rect 429 -22 430 -16
rect 439 -22 440 -16
rect 506 -22 507 -16
rect 509 -17 510 -11
rect 100 -22 101 -18
rect 121 -19 122 -11
rect 236 -22 237 -18
rect 282 -22 283 -18
rect 268 -22 269 -20
rect 303 -22 304 -20
rect 86 -53 87 -31
rect 103 -32 104 -30
rect 114 -53 115 -31
rect 187 -53 188 -31
rect 191 -53 192 -31
rect 219 -32 220 -30
rect 226 -32 227 -30
rect 229 -50 230 -31
rect 247 -32 248 -30
rect 352 -53 353 -31
rect 359 -32 360 -30
rect 408 -53 409 -31
rect 415 -32 416 -30
rect 422 -32 423 -30
rect 429 -32 430 -30
rect 436 -53 437 -31
rect 446 -32 447 -30
rect 499 -53 500 -31
rect 506 -32 507 -30
rect 506 -53 507 -31
rect 506 -32 507 -30
rect 506 -53 507 -31
rect 520 -32 521 -30
rect 534 -53 535 -31
rect 551 -53 552 -31
rect 562 -53 563 -31
rect 569 -32 570 -30
rect 597 -53 598 -31
rect 604 -32 605 -30
rect 639 -53 640 -31
rect 663 -53 664 -31
rect 667 -53 668 -31
rect 674 -32 675 -30
rect 702 -53 703 -31
rect 765 -53 766 -31
rect 842 -53 843 -31
rect 93 -53 94 -33
rect 100 -34 101 -30
rect 121 -53 122 -33
rect 135 -34 136 -30
rect 163 -53 164 -33
rect 236 -53 237 -33
rect 247 -53 248 -33
rect 254 -34 255 -30
rect 275 -34 276 -30
rect 345 -53 346 -33
rect 366 -53 367 -33
rect 373 -34 374 -30
rect 383 -34 384 -30
rect 394 -53 395 -33
rect 471 -34 472 -30
rect 520 -53 521 -33
rect 527 -34 528 -30
rect 590 -53 591 -33
rect 611 -34 612 -30
rect 653 -53 654 -33
rect 677 -53 678 -33
rect 681 -53 682 -33
rect 128 -53 129 -35
rect 145 -53 146 -35
rect 177 -36 178 -30
rect 194 -36 195 -30
rect 198 -36 199 -30
rect 205 -53 206 -35
rect 212 -36 213 -30
rect 275 -53 276 -35
rect 282 -36 283 -30
rect 303 -53 304 -35
rect 313 -53 314 -35
rect 317 -36 318 -30
rect 338 -36 339 -30
rect 338 -53 339 -35
rect 338 -36 339 -30
rect 338 -53 339 -35
rect 341 -53 342 -35
rect 422 -53 423 -35
rect 464 -36 465 -30
rect 611 -53 612 -35
rect 618 -36 619 -30
rect 646 -53 647 -35
rect 135 -53 136 -37
rect 268 -38 269 -30
rect 282 -53 283 -37
rect 348 -38 349 -30
rect 373 -53 374 -37
rect 443 -53 444 -37
rect 464 -53 465 -37
rect 625 -53 626 -37
rect 156 -53 157 -39
rect 177 -53 178 -39
rect 184 -40 185 -30
rect 219 -53 220 -39
rect 226 -53 227 -39
rect 261 -40 262 -30
rect 268 -53 269 -39
rect 289 -40 290 -30
rect 296 -40 297 -30
rect 429 -53 430 -39
rect 471 -53 472 -39
rect 586 -53 587 -39
rect 198 -53 199 -41
rect 331 -53 332 -41
rect 383 -53 384 -41
rect 485 -53 486 -41
rect 527 -53 528 -41
rect 632 -53 633 -41
rect 201 -53 202 -43
rect 254 -53 255 -43
rect 289 -53 290 -43
rect 324 -44 325 -30
rect 387 -53 388 -43
rect 467 -44 468 -30
rect 478 -53 479 -43
rect 492 -44 493 -30
rect 541 -44 542 -30
rect 569 -53 570 -43
rect 576 -44 577 -30
rect 576 -53 577 -43
rect 576 -44 577 -30
rect 576 -53 577 -43
rect 173 -53 174 -45
rect 324 -53 325 -45
rect 513 -46 514 -30
rect 541 -53 542 -45
rect 555 -46 556 -30
rect 604 -53 605 -45
rect 212 -53 213 -47
rect 299 -53 300 -47
rect 310 -48 311 -30
rect 317 -53 318 -47
rect 555 -53 556 -47
rect 772 -53 773 -47
rect 261 -53 262 -49
rect 250 -53 251 -51
rect 401 -53 402 -51
rect 30 -122 31 -62
rect 152 -122 153 -62
rect 159 -122 160 -62
rect 250 -63 251 -61
rect 317 -63 318 -61
rect 338 -122 339 -62
rect 429 -63 430 -61
rect 821 -122 822 -62
rect 842 -63 843 -61
rect 877 -122 878 -62
rect 58 -122 59 -64
rect 107 -122 108 -64
rect 114 -65 115 -61
rect 173 -65 174 -61
rect 198 -122 199 -64
rect 205 -65 206 -61
rect 219 -65 220 -61
rect 229 -122 230 -64
rect 233 -65 234 -61
rect 345 -65 346 -61
rect 394 -65 395 -61
rect 429 -122 430 -64
rect 450 -122 451 -64
rect 467 -65 468 -61
rect 471 -65 472 -61
rect 474 -81 475 -64
rect 485 -65 486 -61
rect 513 -122 514 -64
rect 530 -65 531 -61
rect 688 -122 689 -64
rect 702 -65 703 -61
rect 779 -122 780 -64
rect 37 -122 38 -66
rect 173 -122 174 -66
rect 219 -122 220 -66
rect 278 -122 279 -66
rect 317 -122 318 -66
rect 716 -122 717 -66
rect 772 -67 773 -61
rect 870 -122 871 -66
rect 61 -122 62 -68
rect 320 -122 321 -68
rect 324 -69 325 -61
rect 380 -69 381 -61
rect 457 -122 458 -68
rect 555 -69 556 -61
rect 583 -69 584 -61
rect 793 -122 794 -68
rect 65 -122 66 -70
rect 93 -71 94 -61
rect 100 -122 101 -70
rect 205 -122 206 -70
rect 233 -122 234 -70
rect 387 -71 388 -61
rect 464 -122 465 -70
rect 478 -71 479 -61
rect 485 -122 486 -70
rect 499 -71 500 -61
rect 502 -122 503 -70
rect 807 -122 808 -70
rect 72 -122 73 -72
rect 128 -73 129 -61
rect 142 -122 143 -72
rect 243 -73 244 -61
rect 254 -73 255 -61
rect 555 -122 556 -72
rect 590 -73 591 -61
rect 772 -122 773 -72
rect 79 -122 80 -74
rect 86 -75 87 -61
rect 93 -122 94 -74
rect 303 -75 304 -61
rect 331 -75 332 -61
rect 695 -122 696 -74
rect 702 -122 703 -74
rect 765 -75 766 -61
rect 86 -122 87 -76
rect 282 -77 283 -61
rect 289 -77 290 -61
rect 324 -122 325 -76
rect 331 -122 332 -76
rect 352 -77 353 -61
rect 376 -122 377 -76
rect 478 -122 479 -76
rect 495 -77 496 -61
rect 828 -122 829 -76
rect 103 -122 104 -78
rect 282 -122 283 -78
rect 380 -122 381 -78
rect 408 -79 409 -61
rect 471 -122 472 -78
rect 492 -79 493 -61
rect 506 -79 507 -61
rect 509 -122 510 -78
rect 548 -79 549 -61
rect 618 -122 619 -78
rect 625 -79 626 -61
rect 814 -122 815 -78
rect 117 -122 118 -80
rect 170 -81 171 -61
rect 240 -81 241 -61
rect 408 -122 409 -80
rect 492 -122 493 -80
rect 569 -81 570 -61
rect 625 -122 626 -80
rect 632 -81 633 -61
rect 786 -122 787 -80
rect 51 -122 52 -82
rect 240 -122 241 -82
rect 261 -83 262 -61
rect 303 -122 304 -82
rect 355 -122 356 -82
rect 632 -122 633 -82
rect 639 -83 640 -61
rect 744 -122 745 -82
rect 121 -85 122 -61
rect 254 -122 255 -84
rect 268 -85 269 -61
rect 289 -122 290 -84
rect 387 -122 388 -84
rect 835 -122 836 -84
rect 121 -122 122 -86
rect 163 -87 164 -61
rect 247 -122 248 -86
rect 261 -122 262 -86
rect 268 -122 269 -86
rect 373 -87 374 -61
rect 397 -122 398 -86
rect 548 -122 549 -86
rect 586 -87 587 -61
rect 590 -122 591 -86
rect 604 -87 605 -61
rect 737 -122 738 -86
rect 128 -122 129 -88
rect 674 -122 675 -88
rect 681 -89 682 -61
rect 730 -122 731 -88
rect 149 -91 150 -61
rect 156 -91 157 -61
rect 163 -122 164 -90
rect 418 -91 419 -61
rect 527 -122 528 -90
rect 586 -122 587 -90
rect 597 -91 598 -61
rect 681 -122 682 -90
rect 709 -122 710 -90
rect 842 -122 843 -90
rect 401 -93 402 -61
rect 569 -122 570 -92
rect 576 -93 577 -61
rect 597 -122 598 -92
rect 611 -93 612 -61
rect 723 -122 724 -92
rect 366 -95 367 -61
rect 401 -122 402 -94
rect 443 -95 444 -61
rect 611 -122 612 -94
rect 646 -95 647 -61
rect 758 -122 759 -94
rect 359 -97 360 -61
rect 646 -122 647 -96
rect 653 -97 654 -61
rect 751 -122 752 -96
rect 226 -99 227 -61
rect 359 -122 360 -98
rect 436 -99 437 -61
rect 443 -122 444 -98
rect 520 -99 521 -61
rect 653 -122 654 -98
rect 660 -99 661 -61
rect 765 -122 766 -98
rect 177 -101 178 -61
rect 226 -122 227 -100
rect 310 -101 311 -61
rect 520 -122 521 -100
rect 534 -101 535 -61
rect 639 -122 640 -100
rect 667 -101 668 -61
rect 800 -122 801 -100
rect 156 -122 157 -102
rect 667 -122 668 -102
rect 177 -122 178 -104
rect 212 -105 213 -61
rect 310 -122 311 -104
rect 341 -105 342 -61
rect 415 -122 416 -104
rect 436 -122 437 -104
rect 499 -122 500 -104
rect 534 -122 535 -104
rect 541 -105 542 -61
rect 604 -122 605 -104
rect 191 -107 192 -61
rect 212 -122 213 -106
rect 422 -107 423 -61
rect 541 -122 542 -106
rect 562 -107 563 -61
rect 576 -122 577 -106
rect 47 -122 48 -108
rect 422 -122 423 -108
rect 191 -122 192 -110
rect 390 -122 391 -110
rect 296 -113 297 -61
rect 562 -122 563 -112
rect 275 -115 276 -61
rect 296 -122 297 -114
rect 184 -117 185 -61
rect 275 -122 276 -116
rect 135 -119 136 -61
rect 184 -122 185 -118
rect 135 -122 136 -120
rect 366 -122 367 -120
rect 23 -211 24 -131
rect 121 -132 122 -130
rect 128 -132 129 -130
rect 208 -211 209 -131
rect 226 -132 227 -130
rect 688 -132 689 -130
rect 723 -132 724 -130
rect 863 -211 864 -131
rect 870 -132 871 -130
rect 954 -211 955 -131
rect 1108 -132 1109 -130
rect 1108 -211 1109 -131
rect 1108 -132 1109 -130
rect 1108 -211 1109 -131
rect 30 -134 31 -130
rect 135 -134 136 -130
rect 145 -211 146 -133
rect 415 -211 416 -133
rect 436 -134 437 -130
rect 436 -211 437 -133
rect 436 -134 437 -130
rect 436 -211 437 -133
rect 499 -134 500 -130
rect 639 -134 640 -130
rect 751 -134 752 -130
rect 870 -211 871 -133
rect 877 -134 878 -130
rect 912 -211 913 -133
rect 30 -211 31 -135
rect 163 -136 164 -130
rect 170 -136 171 -130
rect 828 -136 829 -130
rect 37 -138 38 -130
rect 100 -211 101 -137
rect 149 -138 150 -130
rect 177 -138 178 -130
rect 250 -211 251 -137
rect 835 -138 836 -130
rect 37 -211 38 -139
rect 205 -140 206 -130
rect 275 -140 276 -130
rect 310 -140 311 -130
rect 317 -140 318 -130
rect 492 -140 493 -130
rect 509 -140 510 -130
rect 737 -140 738 -130
rect 765 -140 766 -130
rect 891 -211 892 -139
rect 44 -211 45 -141
rect 142 -142 143 -130
rect 156 -142 157 -130
rect 821 -142 822 -130
rect 51 -144 52 -130
rect 275 -211 276 -143
rect 299 -211 300 -143
rect 352 -144 353 -130
rect 362 -211 363 -143
rect 919 -211 920 -143
rect 51 -211 52 -145
rect 124 -211 125 -145
rect 142 -211 143 -145
rect 373 -211 374 -145
rect 376 -146 377 -130
rect 569 -146 570 -130
rect 579 -211 580 -145
rect 758 -146 759 -130
rect 772 -146 773 -130
rect 905 -211 906 -145
rect 58 -148 59 -130
rect 646 -148 647 -130
rect 660 -148 661 -130
rect 758 -211 759 -147
rect 779 -148 780 -130
rect 884 -211 885 -147
rect 65 -150 66 -130
rect 114 -150 115 -130
rect 117 -150 118 -130
rect 156 -211 157 -149
rect 159 -150 160 -130
rect 348 -150 349 -130
rect 352 -211 353 -149
rect 541 -150 542 -130
rect 548 -150 549 -130
rect 849 -211 850 -149
rect 79 -152 80 -130
rect 674 -152 675 -130
rect 681 -152 682 -130
rect 779 -211 780 -151
rect 786 -152 787 -130
rect 926 -211 927 -151
rect 79 -211 80 -153
rect 152 -154 153 -130
rect 163 -211 164 -153
rect 198 -154 199 -130
rect 310 -211 311 -153
rect 471 -154 472 -130
rect 495 -211 496 -153
rect 660 -211 661 -153
rect 667 -154 668 -130
rect 765 -211 766 -153
rect 793 -154 794 -130
rect 933 -211 934 -153
rect 86 -156 87 -130
rect 397 -156 398 -130
rect 418 -156 419 -130
rect 639 -211 640 -155
rect 695 -156 696 -130
rect 821 -211 822 -155
rect 89 -211 90 -157
rect 128 -211 129 -157
rect 152 -211 153 -157
rect 856 -211 857 -157
rect 114 -211 115 -159
rect 180 -211 181 -159
rect 198 -211 199 -159
rect 212 -160 213 -130
rect 317 -211 318 -159
rect 408 -160 409 -130
rect 422 -160 423 -130
rect 499 -211 500 -159
rect 513 -160 514 -130
rect 541 -211 542 -159
rect 583 -160 584 -130
rect 898 -211 899 -159
rect 170 -211 171 -161
rect 215 -211 216 -161
rect 320 -162 321 -130
rect 401 -162 402 -130
rect 429 -162 430 -130
rect 513 -211 514 -161
rect 520 -162 521 -130
rect 548 -211 549 -161
rect 583 -211 584 -161
rect 730 -162 731 -130
rect 737 -211 738 -161
rect 877 -211 878 -161
rect 173 -164 174 -130
rect 457 -164 458 -130
rect 464 -164 465 -130
rect 471 -211 472 -163
rect 492 -211 493 -163
rect 695 -211 696 -163
rect 702 -164 703 -130
rect 772 -211 773 -163
rect 800 -164 801 -130
rect 940 -211 941 -163
rect 212 -211 213 -165
rect 303 -166 304 -130
rect 324 -166 325 -130
rect 355 -166 356 -130
rect 359 -166 360 -130
rect 408 -211 409 -165
rect 443 -166 444 -130
rect 786 -211 787 -165
rect 814 -166 815 -130
rect 947 -211 948 -165
rect 65 -211 66 -167
rect 359 -211 360 -167
rect 380 -168 381 -130
rect 464 -211 465 -167
rect 506 -168 507 -130
rect 800 -211 801 -167
rect 93 -170 94 -130
rect 380 -211 381 -169
rect 387 -211 388 -169
rect 429 -211 430 -169
rect 520 -211 521 -169
rect 835 -211 836 -169
rect 93 -211 94 -171
rect 184 -172 185 -130
rect 219 -172 220 -130
rect 303 -211 304 -171
rect 324 -211 325 -171
rect 688 -211 689 -171
rect 709 -172 710 -130
rect 751 -211 752 -171
rect 135 -211 136 -173
rect 219 -211 220 -173
rect 261 -174 262 -130
rect 506 -211 507 -173
rect 523 -211 524 -173
rect 723 -211 724 -173
rect 107 -176 108 -130
rect 261 -211 262 -175
rect 327 -211 328 -175
rect 338 -176 339 -130
rect 345 -176 346 -130
rect 422 -211 423 -175
rect 534 -176 535 -130
rect 569 -211 570 -175
rect 590 -176 591 -130
rect 646 -211 647 -175
rect 716 -176 717 -130
rect 828 -211 829 -175
rect 184 -211 185 -177
rect 191 -178 192 -130
rect 268 -178 269 -130
rect 338 -211 339 -177
rect 348 -211 349 -177
rect 527 -178 528 -130
rect 597 -178 598 -130
rect 730 -211 731 -177
rect 72 -180 73 -130
rect 597 -211 598 -179
rect 611 -180 612 -130
rect 667 -211 668 -179
rect 72 -211 73 -181
rect 702 -211 703 -181
rect 191 -211 192 -183
rect 229 -184 230 -130
rect 268 -211 269 -183
rect 289 -184 290 -130
rect 331 -184 332 -130
rect 443 -211 444 -183
rect 450 -184 451 -130
rect 534 -211 535 -183
rect 555 -184 556 -130
rect 611 -211 612 -183
rect 618 -184 619 -130
rect 709 -211 710 -183
rect 205 -211 206 -185
rect 289 -211 290 -185
rect 334 -211 335 -185
rect 842 -186 843 -130
rect 366 -188 367 -130
rect 450 -211 451 -187
rect 478 -188 479 -130
rect 555 -211 556 -187
rect 618 -211 619 -187
rect 842 -211 843 -187
rect 296 -190 297 -130
rect 366 -211 367 -189
rect 394 -190 395 -130
rect 681 -211 682 -189
rect 282 -192 283 -130
rect 394 -211 395 -191
rect 401 -211 402 -191
rect 674 -211 675 -191
rect 240 -194 241 -130
rect 282 -211 283 -193
rect 296 -211 297 -193
rect 590 -211 591 -193
rect 625 -194 626 -130
rect 793 -211 794 -193
rect 240 -211 241 -195
rect 254 -196 255 -130
rect 478 -211 479 -195
rect 562 -196 563 -130
rect 625 -211 626 -195
rect 814 -211 815 -195
rect 233 -198 234 -130
rect 254 -211 255 -197
rect 345 -211 346 -197
rect 562 -211 563 -197
rect 632 -198 633 -130
rect 716 -211 717 -197
rect 58 -211 59 -199
rect 233 -211 234 -199
rect 485 -200 486 -130
rect 527 -211 528 -199
rect 604 -200 605 -130
rect 632 -211 633 -199
rect 110 -211 111 -201
rect 485 -211 486 -201
rect 576 -202 577 -130
rect 604 -211 605 -201
rect 576 -211 577 -203
rect 744 -204 745 -130
rect 653 -206 654 -130
rect 744 -211 745 -205
rect 653 -211 654 -207
rect 807 -208 808 -130
rect 656 -211 657 -209
rect 807 -211 808 -209
rect 16 -294 17 -220
rect 702 -221 703 -219
rect 723 -221 724 -219
rect 908 -294 909 -220
rect 1108 -221 1109 -219
rect 1108 -294 1109 -220
rect 1108 -221 1109 -219
rect 1108 -294 1109 -220
rect 23 -223 24 -219
rect 208 -223 209 -219
rect 261 -223 262 -219
rect 345 -294 346 -222
rect 352 -223 353 -219
rect 387 -223 388 -219
rect 401 -223 402 -219
rect 828 -223 829 -219
rect 887 -294 888 -222
rect 912 -223 913 -219
rect 23 -294 24 -224
rect 79 -225 80 -219
rect 114 -225 115 -219
rect 233 -294 234 -224
rect 254 -225 255 -219
rect 387 -294 388 -224
rect 471 -225 472 -219
rect 492 -294 493 -224
rect 495 -225 496 -219
rect 905 -225 906 -219
rect 30 -227 31 -219
rect 362 -227 363 -219
rect 366 -227 367 -219
rect 404 -227 405 -219
rect 502 -294 503 -226
rect 555 -227 556 -219
rect 579 -227 580 -219
rect 926 -227 927 -219
rect 30 -294 31 -228
rect 156 -229 157 -219
rect 163 -229 164 -219
rect 222 -229 223 -219
rect 296 -294 297 -228
rect 394 -294 395 -228
rect 555 -294 556 -228
rect 611 -229 612 -219
rect 618 -229 619 -219
rect 863 -229 864 -219
rect 44 -231 45 -219
rect 138 -294 139 -230
rect 142 -231 143 -219
rect 534 -231 535 -219
rect 604 -231 605 -219
rect 604 -294 605 -230
rect 604 -231 605 -219
rect 604 -294 605 -230
rect 611 -294 612 -230
rect 667 -231 668 -219
rect 674 -231 675 -219
rect 905 -294 906 -230
rect 51 -233 52 -219
rect 254 -294 255 -232
rect 299 -233 300 -219
rect 401 -294 402 -232
rect 621 -233 622 -219
rect 898 -233 899 -219
rect 51 -294 52 -234
rect 58 -235 59 -219
rect 65 -235 66 -219
rect 261 -294 262 -234
rect 299 -294 300 -234
rect 408 -235 409 -219
rect 618 -294 619 -234
rect 898 -294 899 -234
rect 58 -294 59 -236
rect 467 -294 468 -236
rect 625 -294 626 -236
rect 660 -237 661 -219
rect 663 -294 664 -236
rect 667 -294 668 -236
rect 674 -294 675 -236
rect 688 -237 689 -219
rect 702 -294 703 -236
rect 779 -237 780 -219
rect 807 -237 808 -219
rect 863 -294 864 -236
rect 65 -294 66 -238
rect 107 -294 108 -238
rect 121 -239 122 -219
rect 562 -239 563 -219
rect 628 -239 629 -219
rect 933 -239 934 -219
rect 68 -294 69 -240
rect 366 -294 367 -240
rect 408 -294 409 -240
rect 436 -241 437 -219
rect 541 -241 542 -219
rect 562 -294 563 -240
rect 639 -241 640 -219
rect 912 -294 913 -240
rect 72 -243 73 -219
rect 303 -243 304 -219
rect 317 -243 318 -219
rect 471 -294 472 -242
rect 541 -294 542 -242
rect 548 -243 549 -219
rect 597 -243 598 -219
rect 639 -294 640 -242
rect 646 -243 647 -219
rect 646 -294 647 -242
rect 646 -243 647 -219
rect 646 -294 647 -242
rect 653 -243 654 -219
rect 947 -243 948 -219
rect 72 -294 73 -244
rect 338 -245 339 -219
rect 359 -245 360 -219
rect 478 -245 479 -219
rect 527 -245 528 -219
rect 548 -294 549 -244
rect 597 -294 598 -244
rect 709 -245 710 -219
rect 723 -294 724 -244
rect 730 -245 731 -219
rect 737 -294 738 -244
rect 744 -245 745 -219
rect 800 -245 801 -219
rect 807 -294 808 -244
rect 828 -294 829 -244
rect 884 -245 885 -219
rect 79 -294 80 -246
rect 114 -294 115 -246
rect 121 -294 122 -246
rect 170 -247 171 -219
rect 177 -247 178 -219
rect 275 -247 276 -219
rect 289 -247 290 -219
rect 303 -294 304 -246
rect 317 -294 318 -246
rect 534 -294 535 -246
rect 653 -294 654 -246
rect 716 -247 717 -219
rect 730 -294 731 -246
rect 772 -247 773 -219
rect 93 -249 94 -219
rect 275 -294 276 -248
rect 324 -249 325 -219
rect 849 -249 850 -219
rect 100 -251 101 -219
rect 156 -294 157 -250
rect 170 -294 171 -250
rect 856 -251 857 -219
rect 100 -294 101 -252
rect 149 -253 150 -219
rect 173 -294 174 -252
rect 289 -294 290 -252
rect 324 -294 325 -252
rect 520 -253 521 -219
rect 688 -294 689 -252
rect 751 -253 752 -219
rect 814 -253 815 -219
rect 849 -294 850 -252
rect 856 -294 857 -252
rect 919 -253 920 -219
rect 117 -294 118 -254
rect 149 -294 150 -254
rect 177 -294 178 -254
rect 184 -255 185 -219
rect 194 -294 195 -254
rect 506 -255 507 -219
rect 695 -255 696 -219
rect 800 -294 801 -254
rect 814 -294 815 -254
rect 835 -255 836 -219
rect 919 -294 920 -254
rect 954 -255 955 -219
rect 93 -294 94 -256
rect 184 -294 185 -256
rect 198 -257 199 -219
rect 226 -294 227 -256
rect 240 -257 241 -219
rect 695 -294 696 -256
rect 709 -294 710 -256
rect 758 -257 759 -219
rect 37 -259 38 -219
rect 240 -294 241 -258
rect 331 -259 332 -219
rect 464 -259 465 -219
rect 485 -259 486 -219
rect 772 -294 773 -258
rect 37 -294 38 -260
rect 247 -261 248 -219
rect 331 -294 332 -260
rect 569 -261 570 -219
rect 740 -261 741 -219
rect 779 -294 780 -260
rect 47 -294 48 -262
rect 198 -294 199 -262
rect 205 -263 206 -219
rect 205 -294 206 -262
rect 205 -263 206 -219
rect 205 -294 206 -262
rect 219 -263 220 -219
rect 478 -294 479 -262
rect 485 -294 486 -262
rect 940 -263 941 -219
rect 135 -265 136 -219
rect 166 -294 167 -264
rect 219 -294 220 -264
rect 229 -265 230 -219
rect 247 -294 248 -264
rect 268 -265 269 -219
rect 338 -294 339 -264
rect 380 -265 381 -219
rect 397 -265 398 -219
rect 835 -294 836 -264
rect 86 -294 87 -266
rect 135 -294 136 -266
rect 142 -294 143 -266
rect 212 -267 213 -219
rect 282 -267 283 -219
rect 380 -294 381 -266
rect 436 -294 437 -266
rect 786 -267 787 -219
rect 128 -269 129 -219
rect 268 -294 269 -268
rect 282 -294 283 -268
rect 355 -294 356 -268
rect 362 -294 363 -268
rect 590 -269 591 -219
rect 744 -294 745 -268
rect 765 -269 766 -219
rect 191 -271 192 -219
rect 212 -294 213 -270
rect 450 -271 451 -219
rect 527 -294 528 -270
rect 583 -271 584 -219
rect 786 -294 787 -270
rect 191 -294 192 -272
rect 429 -273 430 -219
rect 443 -273 444 -219
rect 583 -294 584 -272
rect 590 -294 591 -272
rect 632 -273 633 -219
rect 751 -294 752 -272
rect 821 -273 822 -219
rect 334 -275 335 -219
rect 429 -294 430 -274
rect 488 -294 489 -274
rect 716 -294 717 -274
rect 758 -294 759 -274
rect 793 -275 794 -219
rect 821 -294 822 -274
rect 842 -275 843 -219
rect 415 -277 416 -219
rect 443 -294 444 -276
rect 506 -294 507 -276
rect 513 -277 514 -219
rect 632 -294 633 -276
rect 681 -277 682 -219
rect 793 -294 794 -276
rect 870 -277 871 -219
rect 152 -279 153 -219
rect 513 -294 514 -278
rect 842 -294 843 -278
rect 877 -279 878 -219
rect 257 -294 258 -280
rect 681 -294 682 -280
rect 870 -294 871 -280
rect 891 -281 892 -219
rect 310 -283 311 -219
rect 415 -294 416 -282
rect 422 -283 423 -219
rect 450 -294 451 -282
rect 576 -283 577 -219
rect 877 -294 878 -282
rect 310 -294 311 -284
rect 520 -294 521 -284
rect 373 -287 374 -219
rect 422 -294 423 -286
rect 457 -287 458 -219
rect 576 -294 577 -286
rect 373 -294 374 -288
rect 765 -294 766 -288
rect 457 -294 458 -290
rect 499 -291 500 -219
rect 499 -294 500 -292
rect 569 -294 570 -292
rect 16 -304 17 -302
rect 184 -304 185 -302
rect 240 -304 241 -302
rect 474 -389 475 -303
rect 492 -304 493 -302
rect 520 -389 521 -303
rect 523 -304 524 -302
rect 856 -304 857 -302
rect 863 -304 864 -302
rect 905 -389 906 -303
rect 1108 -304 1109 -302
rect 1108 -389 1109 -303
rect 1108 -304 1109 -302
rect 1108 -389 1109 -303
rect 23 -306 24 -302
rect 100 -306 101 -302
rect 110 -389 111 -305
rect 121 -306 122 -302
rect 124 -389 125 -305
rect 131 -306 132 -302
rect 159 -389 160 -305
rect 250 -389 251 -305
rect 254 -389 255 -305
rect 387 -306 388 -302
rect 394 -389 395 -305
rect 884 -306 885 -302
rect 898 -389 899 -305
rect 912 -306 913 -302
rect 23 -389 24 -307
rect 208 -308 209 -302
rect 233 -308 234 -302
rect 240 -389 241 -307
rect 247 -308 248 -302
rect 320 -308 321 -302
rect 352 -308 353 -302
rect 467 -308 468 -302
rect 544 -389 545 -307
rect 653 -308 654 -302
rect 660 -389 661 -307
rect 744 -308 745 -302
rect 800 -308 801 -302
rect 880 -389 881 -307
rect 30 -310 31 -302
rect 352 -389 353 -309
rect 355 -310 356 -302
rect 506 -310 507 -302
rect 516 -389 517 -309
rect 744 -389 745 -309
rect 835 -310 836 -302
rect 887 -389 888 -309
rect 37 -312 38 -302
rect 96 -389 97 -311
rect 100 -389 101 -311
rect 198 -312 199 -302
rect 233 -389 234 -311
rect 628 -389 629 -311
rect 681 -312 682 -302
rect 933 -389 934 -311
rect 37 -389 38 -313
rect 299 -314 300 -302
rect 306 -389 307 -313
rect 800 -389 801 -313
rect 807 -314 808 -302
rect 835 -389 836 -313
rect 863 -389 864 -313
rect 870 -314 871 -302
rect 877 -314 878 -302
rect 891 -389 892 -313
rect 44 -389 45 -315
rect 103 -316 104 -302
rect 117 -316 118 -302
rect 156 -316 157 -302
rect 170 -316 171 -302
rect 541 -316 542 -302
rect 625 -316 626 -302
rect 653 -389 654 -315
rect 786 -316 787 -302
rect 870 -389 871 -315
rect 877 -389 878 -315
rect 919 -316 920 -302
rect 47 -318 48 -302
rect 555 -318 556 -302
rect 646 -318 647 -302
rect 681 -389 682 -317
rect 716 -318 717 -302
rect 786 -389 787 -317
rect 793 -318 794 -302
rect 807 -389 808 -317
rect 58 -320 59 -302
rect 401 -320 402 -302
rect 422 -320 423 -302
rect 488 -320 489 -302
rect 541 -389 542 -319
rect 723 -320 724 -302
rect 730 -320 731 -302
rect 793 -389 794 -319
rect 58 -389 59 -321
rect 86 -322 87 -302
rect 128 -322 129 -302
rect 135 -322 136 -302
rect 149 -322 150 -302
rect 198 -389 199 -321
rect 261 -322 262 -302
rect 261 -389 262 -321
rect 261 -322 262 -302
rect 261 -389 262 -321
rect 268 -322 269 -302
rect 499 -389 500 -321
rect 576 -322 577 -302
rect 716 -389 717 -321
rect 65 -324 66 -302
rect 373 -324 374 -302
rect 439 -324 440 -302
rect 737 -324 738 -302
rect 9 -389 10 -325
rect 65 -389 66 -325
rect 68 -326 69 -302
rect 751 -326 752 -302
rect 68 -389 69 -327
rect 86 -389 87 -327
rect 128 -389 129 -327
rect 163 -328 164 -302
rect 173 -328 174 -302
rect 639 -328 640 -302
rect 702 -328 703 -302
rect 751 -389 752 -327
rect 79 -330 80 -302
rect 114 -389 115 -329
rect 135 -389 136 -329
rect 723 -389 724 -329
rect 79 -389 80 -331
rect 849 -332 850 -302
rect 82 -389 83 -333
rect 506 -389 507 -333
rect 527 -334 528 -302
rect 576 -389 577 -333
rect 597 -334 598 -302
rect 730 -389 731 -333
rect 842 -334 843 -302
rect 849 -389 850 -333
rect 149 -389 150 -335
rect 219 -336 220 -302
rect 268 -389 269 -335
rect 275 -336 276 -302
rect 296 -336 297 -302
rect 443 -336 444 -302
rect 464 -336 465 -302
rect 772 -336 773 -302
rect 16 -389 17 -337
rect 219 -389 220 -337
rect 275 -389 276 -337
rect 485 -338 486 -302
rect 513 -338 514 -302
rect 527 -389 528 -337
rect 583 -338 584 -302
rect 597 -389 598 -337
rect 618 -338 619 -302
rect 639 -389 640 -337
rect 674 -338 675 -302
rect 702 -389 703 -337
rect 709 -338 710 -302
rect 737 -389 738 -337
rect 772 -389 773 -337
rect 779 -338 780 -302
rect 163 -389 164 -339
rect 187 -389 188 -339
rect 191 -340 192 -302
rect 401 -389 402 -339
rect 404 -340 405 -302
rect 618 -389 619 -339
rect 667 -340 668 -302
rect 674 -389 675 -339
rect 688 -340 689 -302
rect 842 -389 843 -339
rect 170 -389 171 -341
rect 191 -389 192 -341
rect 205 -342 206 -302
rect 583 -389 584 -341
rect 709 -389 710 -341
rect 894 -342 895 -302
rect 173 -389 174 -343
rect 331 -344 332 -302
rect 345 -344 346 -302
rect 688 -389 689 -343
rect 779 -389 780 -343
rect 828 -344 829 -302
rect 72 -346 73 -302
rect 345 -389 346 -345
rect 359 -346 360 -302
rect 670 -389 671 -345
rect 814 -346 815 -302
rect 828 -389 829 -345
rect 72 -389 73 -347
rect 121 -389 122 -347
rect 177 -348 178 -302
rect 177 -389 178 -347
rect 177 -348 178 -302
rect 177 -389 178 -347
rect 205 -389 206 -347
rect 215 -389 216 -347
rect 289 -348 290 -302
rect 296 -389 297 -347
rect 310 -348 311 -302
rect 387 -389 388 -347
rect 408 -348 409 -302
rect 485 -389 486 -347
rect 513 -389 514 -347
rect 590 -348 591 -302
rect 814 -389 815 -347
rect 821 -348 822 -302
rect 194 -350 195 -302
rect 821 -389 822 -349
rect 226 -352 227 -302
rect 289 -389 290 -351
rect 310 -389 311 -351
rect 415 -352 416 -302
rect 443 -389 444 -351
rect 695 -352 696 -302
rect 212 -354 213 -302
rect 226 -389 227 -353
rect 247 -389 248 -353
rect 415 -389 416 -353
rect 450 -354 451 -302
rect 464 -389 465 -353
rect 471 -354 472 -302
rect 646 -389 647 -353
rect 257 -389 258 -355
rect 408 -389 409 -355
rect 562 -356 563 -302
rect 590 -389 591 -355
rect 632 -356 633 -302
rect 695 -389 696 -355
rect 264 -389 265 -357
rect 562 -389 563 -357
rect 604 -358 605 -302
rect 632 -389 633 -357
rect 282 -360 283 -302
rect 450 -389 451 -359
rect 142 -362 143 -302
rect 282 -389 283 -361
rect 317 -389 318 -361
rect 611 -362 612 -302
rect 107 -364 108 -302
rect 142 -389 143 -363
rect 320 -389 321 -363
rect 422 -389 423 -363
rect 429 -364 430 -302
rect 604 -389 605 -363
rect 107 -389 108 -365
rect 856 -389 857 -365
rect 324 -368 325 -302
rect 429 -389 430 -367
rect 534 -368 535 -302
rect 611 -389 612 -367
rect 324 -389 325 -369
rect 765 -370 766 -302
rect 331 -389 332 -371
rect 884 -389 885 -371
rect 341 -389 342 -373
rect 359 -389 360 -373
rect 366 -374 367 -302
rect 555 -389 556 -373
rect 758 -374 759 -302
rect 765 -389 766 -373
rect 303 -376 304 -302
rect 366 -389 367 -375
rect 373 -389 374 -375
rect 457 -376 458 -302
rect 534 -389 535 -375
rect 569 -376 570 -302
rect 51 -378 52 -302
rect 303 -389 304 -377
rect 338 -378 339 -302
rect 457 -389 458 -377
rect 548 -378 549 -302
rect 569 -389 570 -377
rect 51 -389 52 -379
rect 93 -380 94 -302
rect 380 -380 381 -302
rect 548 -389 549 -379
rect 436 -382 437 -302
rect 758 -389 759 -381
rect 397 -384 398 -302
rect 436 -389 437 -383
rect 397 -389 398 -385
rect 478 -386 479 -302
rect 166 -388 167 -302
rect 478 -389 479 -387
rect 2 -478 3 -398
rect 579 -478 580 -398
rect 611 -399 612 -397
rect 996 -478 997 -398
rect 1108 -399 1109 -397
rect 1115 -478 1116 -398
rect 9 -401 10 -397
rect 30 -401 31 -397
rect 44 -401 45 -397
rect 138 -401 139 -397
rect 145 -478 146 -400
rect 443 -401 444 -397
rect 464 -401 465 -397
rect 464 -478 465 -400
rect 464 -401 465 -397
rect 464 -478 465 -400
rect 474 -401 475 -397
rect 842 -401 843 -397
rect 849 -401 850 -397
rect 975 -478 976 -400
rect 982 -478 983 -400
rect 1031 -478 1032 -400
rect 16 -478 17 -402
rect 100 -403 101 -397
rect 107 -478 108 -402
rect 331 -403 332 -397
rect 338 -478 339 -402
rect 366 -403 367 -397
rect 380 -403 381 -397
rect 513 -478 514 -402
rect 569 -403 570 -397
rect 611 -478 612 -402
rect 628 -403 629 -397
rect 870 -403 871 -397
rect 884 -403 885 -397
rect 898 -403 899 -397
rect 905 -403 906 -397
rect 905 -478 906 -402
rect 905 -403 906 -397
rect 905 -478 906 -402
rect 933 -403 934 -397
rect 1045 -478 1046 -402
rect 23 -405 24 -397
rect 156 -405 157 -397
rect 170 -405 171 -397
rect 800 -405 801 -397
rect 807 -405 808 -397
rect 954 -478 955 -404
rect 989 -478 990 -404
rect 1038 -478 1039 -404
rect 23 -478 24 -406
rect 51 -407 52 -397
rect 58 -407 59 -397
rect 366 -478 367 -406
rect 380 -478 381 -406
rect 506 -407 507 -397
rect 569 -478 570 -406
rect 821 -407 822 -397
rect 828 -407 829 -397
rect 926 -478 927 -406
rect 37 -409 38 -397
rect 331 -478 332 -408
rect 341 -409 342 -397
rect 401 -409 402 -397
rect 422 -409 423 -397
rect 443 -478 444 -408
rect 474 -478 475 -408
rect 1024 -478 1025 -408
rect 44 -478 45 -410
rect 275 -411 276 -397
rect 296 -411 297 -397
rect 303 -478 304 -410
rect 306 -411 307 -397
rect 807 -478 808 -410
rect 863 -411 864 -397
rect 1010 -478 1011 -410
rect 51 -478 52 -412
rect 310 -413 311 -397
rect 327 -413 328 -397
rect 688 -413 689 -397
rect 702 -413 703 -397
rect 828 -478 829 -412
rect 835 -413 836 -397
rect 863 -478 864 -412
rect 891 -413 892 -397
rect 1017 -478 1018 -412
rect 65 -478 66 -414
rect 583 -415 584 -397
rect 625 -415 626 -397
rect 933 -478 934 -414
rect 79 -417 80 -397
rect 352 -417 353 -397
rect 383 -417 384 -397
rect 548 -417 549 -397
rect 572 -478 573 -416
rect 961 -478 962 -416
rect 79 -478 80 -418
rect 128 -419 129 -397
rect 135 -478 136 -418
rect 520 -419 521 -397
rect 576 -419 577 -397
rect 625 -478 626 -418
rect 635 -478 636 -418
rect 793 -419 794 -397
rect 814 -419 815 -397
rect 891 -478 892 -418
rect 82 -421 83 -397
rect 702 -478 703 -420
rect 709 -421 710 -397
rect 800 -478 801 -420
rect 96 -423 97 -397
rect 821 -478 822 -422
rect 100 -478 101 -424
rect 422 -478 423 -424
rect 478 -425 479 -397
rect 583 -478 584 -424
rect 632 -425 633 -397
rect 709 -478 710 -424
rect 723 -425 724 -397
rect 842 -478 843 -424
rect 114 -478 115 -426
rect 471 -427 472 -397
rect 485 -427 486 -397
rect 548 -478 549 -426
rect 576 -478 577 -426
rect 849 -478 850 -426
rect 117 -429 118 -397
rect 856 -429 857 -397
rect 121 -431 122 -397
rect 387 -431 388 -397
rect 397 -478 398 -430
rect 646 -431 647 -397
rect 667 -431 668 -397
rect 856 -478 857 -430
rect 86 -433 87 -397
rect 387 -478 388 -432
rect 401 -478 402 -432
rect 499 -433 500 -397
rect 506 -478 507 -432
rect 558 -478 559 -432
rect 590 -433 591 -397
rect 646 -478 647 -432
rect 667 -478 668 -432
rect 751 -433 752 -397
rect 765 -433 766 -397
rect 898 -478 899 -432
rect 72 -435 73 -397
rect 86 -478 87 -434
rect 121 -478 122 -434
rect 163 -435 164 -397
rect 170 -478 171 -434
rect 261 -435 262 -397
rect 264 -435 265 -397
rect 562 -435 563 -397
rect 590 -478 591 -434
rect 604 -435 605 -397
rect 681 -435 682 -397
rect 765 -478 766 -434
rect 772 -435 773 -397
rect 912 -478 913 -434
rect 72 -478 73 -436
rect 131 -478 132 -436
rect 149 -437 150 -397
rect 163 -478 164 -436
rect 184 -437 185 -397
rect 618 -437 619 -397
rect 639 -437 640 -397
rect 772 -478 773 -436
rect 786 -437 787 -397
rect 947 -478 948 -436
rect 61 -478 62 -438
rect 618 -478 619 -438
rect 653 -439 654 -397
rect 786 -478 787 -438
rect 149 -478 150 -440
rect 373 -441 374 -397
rect 408 -441 409 -397
rect 520 -478 521 -440
rect 534 -441 535 -397
rect 604 -478 605 -440
rect 688 -478 689 -440
rect 870 -478 871 -440
rect 12 -478 13 -442
rect 408 -478 409 -442
rect 429 -443 430 -397
rect 485 -478 486 -442
rect 492 -443 493 -397
rect 919 -478 920 -442
rect 156 -478 157 -444
rect 177 -445 178 -397
rect 184 -478 185 -444
rect 191 -445 192 -397
rect 198 -445 199 -397
rect 261 -478 262 -444
rect 268 -445 269 -397
rect 320 -445 321 -397
rect 327 -478 328 -444
rect 457 -445 458 -397
rect 460 -478 461 -444
rect 751 -478 752 -444
rect 177 -478 178 -446
rect 212 -478 213 -446
rect 219 -447 220 -397
rect 296 -478 297 -446
rect 352 -478 353 -446
rect 1003 -478 1004 -446
rect 180 -478 181 -448
rect 219 -478 220 -448
rect 233 -449 234 -397
rect 310 -478 311 -448
rect 373 -478 374 -448
rect 527 -449 528 -397
rect 534 -478 535 -448
rect 660 -449 661 -397
rect 716 -449 717 -397
rect 723 -478 724 -448
rect 730 -449 731 -397
rect 884 -478 885 -448
rect 187 -451 188 -397
rect 415 -451 416 -397
rect 425 -478 426 -450
rect 660 -478 661 -450
rect 695 -451 696 -397
rect 730 -478 731 -450
rect 737 -451 738 -397
rect 968 -478 969 -450
rect 191 -478 192 -452
rect 877 -453 878 -397
rect 198 -478 199 -454
rect 226 -455 227 -397
rect 233 -478 234 -454
rect 394 -455 395 -397
rect 429 -478 430 -454
rect 436 -455 437 -397
rect 450 -455 451 -397
rect 527 -478 528 -454
rect 597 -455 598 -397
rect 716 -478 717 -454
rect 744 -455 745 -397
rect 835 -478 836 -454
rect 205 -457 206 -397
rect 226 -478 227 -456
rect 247 -457 248 -397
rect 268 -478 269 -456
rect 275 -478 276 -456
rect 502 -478 503 -456
rect 516 -457 517 -397
rect 737 -478 738 -456
rect 758 -457 759 -397
rect 877 -478 878 -456
rect 93 -459 94 -397
rect 205 -478 206 -458
rect 240 -459 241 -397
rect 247 -478 248 -458
rect 250 -459 251 -397
rect 289 -459 290 -397
rect 317 -459 318 -397
rect 436 -478 437 -458
rect 457 -478 458 -458
rect 940 -478 941 -458
rect 93 -478 94 -460
rect 124 -478 125 -460
rect 142 -461 143 -397
rect 240 -478 241 -460
rect 254 -461 255 -397
rect 1034 -478 1035 -460
rect 68 -478 69 -462
rect 254 -478 255 -462
rect 282 -463 283 -397
rect 383 -478 384 -462
rect 481 -478 482 -462
rect 653 -478 654 -462
rect 674 -463 675 -397
rect 744 -478 745 -462
rect 110 -465 111 -397
rect 317 -478 318 -464
rect 359 -465 360 -397
rect 450 -478 451 -464
rect 495 -465 496 -397
rect 793 -478 794 -464
rect 142 -478 143 -466
rect 681 -478 682 -466
rect 695 -478 696 -466
rect 779 -467 780 -397
rect 173 -469 174 -397
rect 289 -478 290 -468
rect 345 -469 346 -397
rect 359 -478 360 -468
rect 499 -478 500 -468
rect 597 -478 598 -468
rect 30 -478 31 -470
rect 345 -478 346 -470
rect 541 -471 542 -397
rect 674 -478 675 -470
rect 324 -473 325 -397
rect 541 -478 542 -472
rect 544 -473 545 -397
rect 758 -478 759 -472
rect 37 -478 38 -474
rect 324 -478 325 -474
rect 555 -475 556 -397
rect 779 -478 780 -474
rect 492 -478 493 -476
rect 555 -478 556 -476
rect 9 -595 10 -487
rect 632 -488 633 -486
rect 646 -488 647 -486
rect 646 -595 647 -487
rect 646 -488 647 -486
rect 646 -595 647 -487
rect 814 -488 815 -486
rect 1031 -595 1032 -487
rect 1111 -595 1112 -487
rect 1122 -595 1123 -487
rect 30 -490 31 -486
rect 33 -496 34 -489
rect 44 -490 45 -486
rect 282 -490 283 -486
rect 285 -490 286 -486
rect 618 -490 619 -486
rect 765 -490 766 -486
rect 814 -595 815 -489
rect 817 -490 818 -486
rect 835 -490 836 -486
rect 954 -490 955 -486
rect 1038 -595 1039 -489
rect 1115 -490 1116 -486
rect 1129 -595 1130 -489
rect 23 -492 24 -486
rect 618 -595 619 -491
rect 772 -492 773 -486
rect 835 -595 836 -491
rect 975 -492 976 -486
rect 1052 -595 1053 -491
rect 30 -595 31 -493
rect 212 -494 213 -486
rect 296 -494 297 -486
rect 355 -494 356 -486
rect 373 -494 374 -486
rect 530 -595 531 -493
rect 555 -494 556 -486
rect 912 -494 913 -486
rect 1010 -494 1011 -486
rect 1059 -595 1060 -493
rect 212 -595 213 -495
rect 296 -595 297 -495
rect 310 -496 311 -486
rect 317 -496 318 -486
rect 1073 -595 1074 -495
rect 37 -498 38 -486
rect 282 -595 283 -497
rect 310 -595 311 -497
rect 492 -498 493 -486
rect 499 -595 500 -497
rect 551 -595 552 -497
rect 565 -498 566 -486
rect 968 -498 969 -486
rect 1017 -498 1018 -486
rect 1066 -595 1067 -497
rect 44 -595 45 -499
rect 401 -500 402 -486
rect 415 -500 416 -486
rect 765 -595 766 -499
rect 842 -500 843 -486
rect 1017 -595 1018 -499
rect 1024 -500 1025 -486
rect 1094 -595 1095 -499
rect 16 -502 17 -486
rect 415 -595 416 -501
rect 422 -502 423 -486
rect 604 -502 605 -486
rect 709 -502 710 -486
rect 772 -595 773 -501
rect 863 -502 864 -486
rect 975 -595 976 -501
rect 1045 -502 1046 -486
rect 1115 -595 1116 -501
rect 16 -595 17 -503
rect 352 -504 353 -486
rect 359 -504 360 -486
rect 373 -595 374 -503
rect 397 -504 398 -486
rect 807 -504 808 -486
rect 926 -504 927 -486
rect 968 -595 969 -503
rect 982 -504 983 -486
rect 1045 -595 1046 -503
rect 58 -595 59 -505
rect 72 -506 73 -486
rect 79 -506 80 -486
rect 142 -506 143 -486
rect 149 -506 150 -486
rect 394 -595 395 -505
rect 401 -595 402 -505
rect 418 -506 419 -486
rect 425 -506 426 -486
rect 996 -506 997 -486
rect 61 -508 62 -486
rect 639 -595 640 -507
rect 695 -508 696 -486
rect 926 -595 927 -507
rect 940 -508 941 -486
rect 1010 -595 1011 -507
rect 26 -595 27 -509
rect 940 -595 941 -509
rect 65 -595 66 -511
rect 303 -512 304 -486
rect 327 -512 328 -486
rect 422 -595 423 -511
rect 443 -512 444 -486
rect 478 -595 479 -511
rect 481 -512 482 -486
rect 779 -512 780 -486
rect 800 -512 801 -486
rect 863 -595 864 -511
rect 891 -512 892 -486
rect 982 -595 983 -511
rect 72 -595 73 -513
rect 583 -514 584 -486
rect 597 -514 598 -486
rect 842 -595 843 -513
rect 856 -514 857 -486
rect 891 -595 892 -513
rect 919 -514 920 -486
rect 996 -595 997 -513
rect 79 -595 80 -515
rect 93 -516 94 -486
rect 96 -595 97 -515
rect 240 -516 241 -486
rect 261 -516 262 -486
rect 317 -595 318 -515
rect 338 -516 339 -486
rect 460 -516 461 -486
rect 464 -516 465 -486
rect 471 -516 472 -486
rect 474 -595 475 -515
rect 590 -516 591 -486
rect 597 -595 598 -515
rect 828 -516 829 -486
rect 877 -516 878 -486
rect 919 -595 920 -515
rect 51 -518 52 -486
rect 471 -595 472 -517
rect 485 -518 486 -486
rect 492 -595 493 -517
rect 502 -518 503 -486
rect 730 -518 731 -486
rect 758 -518 759 -486
rect 807 -595 808 -517
rect 51 -595 52 -519
rect 331 -520 332 -486
rect 341 -595 342 -519
rect 632 -595 633 -519
rect 712 -595 713 -519
rect 828 -595 829 -519
rect 100 -522 101 -486
rect 359 -595 360 -521
rect 383 -522 384 -486
rect 856 -595 857 -521
rect 2 -524 3 -486
rect 100 -595 101 -523
rect 114 -524 115 -486
rect 380 -595 381 -523
rect 436 -524 437 -486
rect 485 -595 486 -523
rect 506 -524 507 -486
rect 590 -595 591 -523
rect 600 -595 601 -523
rect 954 -595 955 -523
rect 114 -595 115 -525
rect 208 -526 209 -486
rect 261 -595 262 -525
rect 268 -526 269 -486
rect 271 -595 272 -525
rect 779 -595 780 -525
rect 121 -595 122 -527
rect 562 -528 563 -486
rect 569 -528 570 -486
rect 604 -595 605 -527
rect 716 -528 717 -486
rect 800 -595 801 -527
rect 128 -530 129 -486
rect 387 -530 388 -486
rect 457 -530 458 -486
rect 884 -530 885 -486
rect 107 -532 108 -486
rect 387 -595 388 -531
rect 429 -532 430 -486
rect 457 -595 458 -531
rect 506 -595 507 -531
rect 660 -532 661 -486
rect 758 -595 759 -531
rect 849 -532 850 -486
rect 107 -595 108 -533
rect 821 -534 822 -486
rect 128 -595 129 -535
rect 205 -595 206 -535
rect 303 -595 304 -535
rect 436 -595 437 -535
rect 523 -595 524 -535
rect 898 -536 899 -486
rect 135 -538 136 -486
rect 429 -595 430 -537
rect 534 -538 535 -486
rect 709 -595 710 -537
rect 723 -538 724 -486
rect 898 -595 899 -537
rect 135 -595 136 -539
rect 254 -540 255 -486
rect 324 -540 325 -486
rect 884 -595 885 -539
rect 142 -595 143 -541
rect 275 -542 276 -486
rect 324 -595 325 -541
rect 450 -542 451 -486
rect 534 -595 535 -541
rect 695 -595 696 -541
rect 723 -595 724 -541
rect 786 -542 787 -486
rect 145 -544 146 -486
rect 240 -595 241 -543
rect 247 -544 248 -486
rect 254 -595 255 -543
rect 275 -595 276 -543
rect 289 -544 290 -486
rect 331 -595 332 -543
rect 684 -595 685 -543
rect 688 -544 689 -486
rect 786 -595 787 -543
rect 138 -595 139 -545
rect 289 -595 290 -545
rect 345 -595 346 -545
rect 681 -546 682 -486
rect 744 -546 745 -486
rect 821 -595 822 -545
rect 149 -595 150 -547
rect 233 -548 234 -486
rect 247 -595 248 -547
rect 268 -595 269 -547
rect 348 -548 349 -486
rect 674 -548 675 -486
rect 681 -595 682 -547
rect 933 -548 934 -486
rect 86 -550 87 -486
rect 233 -595 234 -549
rect 348 -595 349 -549
rect 443 -595 444 -549
rect 450 -595 451 -549
rect 464 -595 465 -549
rect 527 -550 528 -486
rect 674 -595 675 -549
rect 702 -550 703 -486
rect 744 -595 745 -549
rect 751 -550 752 -486
rect 849 -595 850 -549
rect 86 -595 87 -551
rect 170 -552 171 -486
rect 180 -595 181 -551
rect 226 -552 227 -486
rect 366 -552 367 -486
rect 660 -595 661 -551
rect 93 -595 94 -553
rect 933 -595 934 -553
rect 156 -556 157 -486
rect 352 -595 353 -555
rect 527 -595 528 -555
rect 583 -595 584 -555
rect 611 -556 612 -486
rect 702 -595 703 -555
rect 156 -595 157 -557
rect 215 -595 216 -557
rect 537 -558 538 -486
rect 877 -595 878 -557
rect 163 -560 164 -486
rect 170 -595 171 -559
rect 191 -560 192 -486
rect 226 -595 227 -559
rect 537 -595 538 -559
rect 667 -560 668 -486
rect 163 -595 164 -561
rect 366 -595 367 -561
rect 541 -562 542 -486
rect 751 -595 752 -561
rect 166 -595 167 -563
rect 1024 -595 1025 -563
rect 184 -566 185 -486
rect 191 -595 192 -565
rect 198 -566 199 -486
rect 1080 -595 1081 -565
rect 184 -595 185 -567
rect 219 -568 220 -486
rect 513 -568 514 -486
rect 541 -595 542 -567
rect 555 -595 556 -567
rect 565 -595 566 -567
rect 572 -568 573 -486
rect 793 -568 794 -486
rect 198 -595 199 -569
rect 208 -595 209 -569
rect 219 -595 220 -569
rect 611 -595 612 -569
rect 625 -570 626 -486
rect 716 -595 717 -569
rect 737 -570 738 -486
rect 793 -595 794 -569
rect 408 -572 409 -486
rect 737 -595 738 -571
rect 408 -595 409 -573
rect 576 -595 577 -573
rect 579 -595 580 -573
rect 912 -595 913 -573
rect 513 -595 514 -575
rect 520 -576 521 -486
rect 562 -595 563 -575
rect 1087 -595 1088 -575
rect 625 -595 626 -577
rect 653 -578 654 -486
rect 548 -580 549 -486
rect 653 -595 654 -579
rect 548 -595 549 -581
rect 1003 -582 1004 -486
rect 635 -584 636 -486
rect 667 -595 668 -583
rect 989 -584 990 -486
rect 1003 -595 1004 -583
rect 642 -586 643 -486
rect 688 -595 689 -585
rect 961 -586 962 -486
rect 989 -595 990 -585
rect 905 -588 906 -486
rect 961 -595 962 -587
rect 905 -595 906 -589
rect 947 -590 948 -486
rect 870 -592 871 -486
rect 947 -595 948 -591
rect 572 -595 573 -593
rect 870 -595 871 -593
rect 2 -605 3 -603
rect 233 -605 234 -603
rect 240 -605 241 -603
rect 240 -696 241 -604
rect 240 -605 241 -603
rect 240 -696 241 -604
rect 254 -605 255 -603
rect 268 -605 269 -603
rect 289 -605 290 -603
rect 534 -605 535 -603
rect 544 -696 545 -604
rect 1010 -605 1011 -603
rect 1111 -696 1112 -604
rect 1143 -696 1144 -604
rect 2 -696 3 -606
rect 107 -607 108 -603
rect 121 -607 122 -603
rect 268 -696 269 -606
rect 303 -607 304 -603
rect 303 -696 304 -606
rect 303 -607 304 -603
rect 303 -696 304 -606
rect 310 -607 311 -603
rect 523 -607 524 -603
rect 534 -696 535 -606
rect 646 -607 647 -603
rect 684 -607 685 -603
rect 1052 -607 1053 -603
rect 1115 -607 1116 -603
rect 1150 -696 1151 -606
rect 5 -609 6 -603
rect 527 -696 528 -608
rect 548 -609 549 -603
rect 898 -609 899 -603
rect 989 -609 990 -603
rect 1052 -696 1053 -608
rect 1101 -609 1102 -603
rect 1115 -696 1116 -608
rect 1122 -609 1123 -603
rect 1122 -696 1123 -608
rect 1122 -609 1123 -603
rect 1122 -696 1123 -608
rect 1129 -609 1130 -603
rect 1157 -696 1158 -608
rect 9 -611 10 -603
rect 212 -611 213 -603
rect 338 -611 339 -603
rect 751 -611 752 -603
rect 779 -611 780 -603
rect 779 -696 780 -610
rect 779 -611 780 -603
rect 779 -696 780 -610
rect 793 -611 794 -603
rect 793 -696 794 -610
rect 793 -611 794 -603
rect 793 -696 794 -610
rect 898 -696 899 -610
rect 1045 -611 1046 -603
rect 1094 -611 1095 -603
rect 1101 -696 1102 -610
rect 1129 -696 1130 -610
rect 1139 -696 1140 -610
rect 16 -613 17 -603
rect 348 -613 349 -603
rect 362 -696 363 -612
rect 576 -613 577 -603
rect 579 -613 580 -603
rect 1038 -613 1039 -603
rect 1066 -613 1067 -603
rect 1094 -696 1095 -612
rect 16 -696 17 -614
rect 65 -615 66 -603
rect 72 -615 73 -603
rect 516 -696 517 -614
rect 541 -615 542 -603
rect 576 -696 577 -614
rect 604 -615 605 -603
rect 1108 -615 1109 -603
rect 23 -696 24 -616
rect 128 -617 129 -603
rect 135 -617 136 -603
rect 212 -696 213 -616
rect 338 -696 339 -616
rect 457 -617 458 -603
rect 460 -696 461 -616
rect 842 -617 843 -603
rect 926 -617 927 -603
rect 1066 -696 1067 -616
rect 26 -619 27 -603
rect 58 -619 59 -603
rect 65 -696 66 -618
rect 296 -619 297 -603
rect 341 -619 342 -603
rect 611 -619 612 -603
rect 709 -696 710 -618
rect 786 -619 787 -603
rect 926 -696 927 -618
rect 933 -619 934 -603
rect 961 -619 962 -603
rect 989 -696 990 -618
rect 1024 -619 1025 -603
rect 1045 -696 1046 -618
rect 37 -621 38 -603
rect 618 -621 619 -603
rect 712 -621 713 -603
rect 1087 -621 1088 -603
rect 47 -696 48 -622
rect 345 -623 346 -603
rect 366 -623 367 -603
rect 565 -696 566 -622
rect 569 -623 570 -603
rect 737 -623 738 -603
rect 786 -696 787 -622
rect 975 -623 976 -603
rect 1031 -623 1032 -603
rect 1087 -696 1088 -622
rect 51 -625 52 -603
rect 233 -696 234 -624
rect 292 -696 293 -624
rect 611 -696 612 -624
rect 618 -696 619 -624
rect 744 -625 745 -603
rect 905 -625 906 -603
rect 975 -696 976 -624
rect 982 -625 983 -603
rect 1031 -696 1032 -624
rect 44 -627 45 -603
rect 51 -696 52 -626
rect 58 -696 59 -626
rect 170 -627 171 -603
rect 173 -696 174 -626
rect 660 -627 661 -603
rect 730 -696 731 -626
rect 807 -627 808 -603
rect 870 -627 871 -603
rect 905 -696 906 -626
rect 912 -627 913 -603
rect 961 -696 962 -626
rect 968 -627 969 -603
rect 982 -696 983 -626
rect 40 -629 41 -603
rect 660 -696 661 -628
rect 726 -696 727 -628
rect 968 -696 969 -628
rect 44 -696 45 -630
rect 765 -631 766 -603
rect 933 -696 934 -630
rect 940 -631 941 -603
rect 72 -696 73 -632
rect 79 -633 80 -603
rect 86 -633 87 -603
rect 215 -633 216 -603
rect 296 -696 297 -632
rect 597 -633 598 -603
rect 604 -696 605 -632
rect 835 -633 836 -603
rect 940 -696 941 -632
rect 947 -633 948 -603
rect 86 -696 87 -634
rect 142 -635 143 -603
rect 156 -635 157 -603
rect 254 -696 255 -634
rect 317 -635 318 -603
rect 345 -696 346 -634
rect 359 -635 360 -603
rect 366 -696 367 -634
rect 373 -635 374 -603
rect 373 -696 374 -634
rect 373 -635 374 -603
rect 373 -696 374 -634
rect 380 -635 381 -603
rect 383 -645 384 -634
rect 394 -635 395 -603
rect 541 -696 542 -634
rect 548 -696 549 -634
rect 555 -635 556 -603
rect 562 -635 563 -603
rect 1017 -635 1018 -603
rect 37 -696 38 -636
rect 359 -696 360 -636
rect 380 -696 381 -636
rect 387 -637 388 -603
rect 394 -696 395 -636
rect 450 -637 451 -603
rect 453 -696 454 -636
rect 485 -637 486 -603
rect 513 -637 514 -603
rect 569 -696 570 -636
rect 572 -637 573 -603
rect 863 -637 864 -603
rect 947 -696 948 -636
rect 954 -637 955 -603
rect 1003 -637 1004 -603
rect 1017 -696 1018 -636
rect 93 -639 94 -603
rect 1073 -639 1074 -603
rect 93 -696 94 -640
rect 219 -641 220 -603
rect 313 -696 314 -640
rect 317 -696 318 -640
rect 387 -696 388 -640
rect 590 -641 591 -603
rect 597 -696 598 -640
rect 688 -641 689 -603
rect 765 -696 766 -640
rect 772 -641 773 -603
rect 828 -641 829 -603
rect 835 -696 836 -640
rect 863 -696 864 -640
rect 919 -641 920 -603
rect 1059 -641 1060 -603
rect 1073 -696 1074 -640
rect 100 -643 101 -603
rect 996 -643 997 -603
rect 100 -696 101 -644
rect 131 -696 132 -644
rect 135 -696 136 -644
rect 222 -645 223 -603
rect 590 -696 591 -644
rect 625 -645 626 -603
rect 919 -696 920 -644
rect 107 -696 108 -646
rect 184 -647 185 -603
rect 201 -696 202 -646
rect 639 -647 640 -603
rect 688 -696 689 -646
rect 733 -647 734 -603
rect 789 -696 790 -646
rect 996 -696 997 -646
rect 114 -649 115 -603
rect 807 -696 808 -648
rect 117 -696 118 -650
rect 156 -696 157 -650
rect 163 -651 164 -603
rect 282 -651 283 -603
rect 401 -651 402 -603
rect 485 -696 486 -650
rect 495 -696 496 -650
rect 639 -696 640 -650
rect 723 -651 724 -603
rect 828 -696 829 -650
rect 128 -696 129 -652
rect 1038 -696 1039 -652
rect 138 -655 139 -603
rect 800 -655 801 -603
rect 142 -696 143 -656
rect 149 -657 150 -603
rect 163 -696 164 -656
rect 261 -657 262 -603
rect 275 -657 276 -603
rect 282 -696 283 -656
rect 408 -657 409 -603
rect 555 -696 556 -656
rect 562 -696 563 -656
rect 842 -696 843 -656
rect 30 -659 31 -603
rect 149 -696 150 -658
rect 177 -659 178 -603
rect 1003 -696 1004 -658
rect 30 -696 31 -660
rect 82 -696 83 -660
rect 124 -696 125 -660
rect 261 -696 262 -660
rect 275 -696 276 -660
rect 457 -696 458 -660
rect 467 -661 468 -603
rect 653 -661 654 -603
rect 723 -696 724 -660
rect 912 -696 913 -660
rect 177 -696 178 -662
rect 191 -663 192 -603
rect 205 -663 206 -603
rect 352 -663 353 -603
rect 408 -696 409 -662
rect 478 -663 479 -603
rect 513 -696 514 -662
rect 646 -696 647 -662
rect 653 -696 654 -662
rect 702 -663 703 -603
rect 800 -696 801 -662
rect 814 -663 815 -603
rect 184 -696 185 -664
rect 198 -665 199 -603
rect 205 -696 206 -664
rect 324 -665 325 -603
rect 352 -696 353 -664
rect 492 -665 493 -603
rect 520 -665 521 -603
rect 870 -696 871 -664
rect 219 -696 220 -666
rect 247 -667 248 -603
rect 415 -667 416 -603
rect 436 -696 437 -666
rect 439 -667 440 -603
rect 1010 -696 1011 -666
rect 191 -696 192 -668
rect 247 -696 248 -668
rect 415 -696 416 -668
rect 478 -696 479 -668
rect 492 -696 493 -668
rect 674 -669 675 -603
rect 702 -696 703 -668
rect 856 -669 857 -603
rect 226 -671 227 -603
rect 401 -696 402 -670
rect 429 -671 430 -603
rect 625 -696 626 -670
rect 632 -671 633 -603
rect 954 -696 955 -670
rect 422 -673 423 -603
rect 429 -696 430 -672
rect 443 -673 444 -603
rect 520 -696 521 -672
rect 551 -673 552 -603
rect 737 -696 738 -672
rect 775 -696 776 -672
rect 814 -696 815 -672
rect 856 -696 857 -672
rect 891 -673 892 -603
rect 324 -696 325 -674
rect 443 -696 444 -674
rect 450 -696 451 -674
rect 681 -696 682 -674
rect 884 -675 885 -603
rect 891 -696 892 -674
rect 422 -696 423 -676
rect 506 -677 507 -603
rect 583 -677 584 -603
rect 632 -696 633 -676
rect 674 -696 675 -676
rect 695 -677 696 -603
rect 877 -677 878 -603
rect 884 -696 885 -676
rect 103 -679 104 -603
rect 506 -696 507 -678
rect 583 -696 584 -678
rect 607 -696 608 -678
rect 667 -679 668 -603
rect 695 -696 696 -678
rect 849 -679 850 -603
rect 877 -696 878 -678
rect 467 -696 468 -680
rect 1024 -696 1025 -680
rect 471 -683 472 -603
rect 751 -696 752 -682
rect 849 -696 850 -682
rect 1080 -683 1081 -603
rect 471 -696 472 -684
rect 499 -685 500 -603
rect 667 -696 668 -684
rect 758 -685 759 -603
rect 474 -687 475 -603
rect 1059 -696 1060 -686
rect 481 -696 482 -688
rect 499 -696 500 -688
rect 758 -696 759 -688
rect 821 -689 822 -603
rect 716 -691 717 -603
rect 821 -696 822 -690
rect 331 -693 332 -603
rect 716 -696 717 -692
rect 331 -696 332 -694
rect 1080 -696 1081 -694
rect 2 -706 3 -704
rect 114 -706 115 -704
rect 128 -773 129 -705
rect 156 -706 157 -704
rect 208 -706 209 -704
rect 292 -706 293 -704
rect 310 -706 311 -704
rect 485 -706 486 -704
rect 513 -706 514 -704
rect 891 -706 892 -704
rect 936 -773 937 -705
rect 968 -706 969 -704
rect 1080 -706 1081 -704
rect 1143 -706 1144 -704
rect 16 -708 17 -704
rect 369 -773 370 -707
rect 373 -708 374 -704
rect 373 -773 374 -707
rect 373 -708 374 -704
rect 373 -773 374 -707
rect 443 -708 444 -704
rect 772 -708 773 -704
rect 775 -708 776 -704
rect 1031 -708 1032 -704
rect 1083 -708 1084 -704
rect 1150 -708 1151 -704
rect 30 -710 31 -704
rect 198 -710 199 -704
rect 268 -710 269 -704
rect 271 -750 272 -709
rect 282 -710 283 -704
rect 282 -773 283 -709
rect 282 -710 283 -704
rect 282 -773 283 -709
rect 292 -773 293 -709
rect 401 -710 402 -704
rect 446 -710 447 -704
rect 821 -710 822 -704
rect 880 -773 881 -709
rect 884 -710 885 -704
rect 891 -773 892 -709
rect 1010 -710 1011 -704
rect 1031 -773 1032 -709
rect 1129 -710 1130 -704
rect 44 -773 45 -711
rect 51 -712 52 -704
rect 58 -712 59 -704
rect 289 -712 290 -704
rect 327 -773 328 -711
rect 422 -712 423 -704
rect 436 -712 437 -704
rect 446 -773 447 -711
rect 450 -773 451 -711
rect 590 -712 591 -704
rect 604 -773 605 -711
rect 800 -712 801 -704
rect 821 -773 822 -711
rect 870 -712 871 -704
rect 884 -773 885 -711
rect 947 -712 948 -704
rect 968 -773 969 -711
rect 1101 -712 1102 -704
rect 1111 -712 1112 -704
rect 1157 -712 1158 -704
rect 51 -773 52 -713
rect 156 -773 157 -713
rect 177 -714 178 -704
rect 198 -773 199 -713
rect 268 -773 269 -713
rect 275 -714 276 -704
rect 289 -773 290 -713
rect 471 -714 472 -704
rect 478 -714 479 -704
rect 919 -714 920 -704
rect 1122 -714 1123 -704
rect 1122 -773 1123 -713
rect 1122 -714 1123 -704
rect 1122 -773 1123 -713
rect 58 -773 59 -715
rect 296 -716 297 -704
rect 317 -716 318 -704
rect 422 -773 423 -715
rect 436 -773 437 -715
rect 443 -773 444 -715
rect 453 -716 454 -704
rect 569 -716 570 -704
rect 590 -773 591 -715
rect 940 -716 941 -704
rect 72 -718 73 -704
rect 72 -773 73 -717
rect 72 -718 73 -704
rect 72 -773 73 -717
rect 82 -718 83 -704
rect 89 -773 90 -717
rect 114 -773 115 -717
rect 135 -718 136 -704
rect 142 -718 143 -704
rect 159 -773 160 -717
rect 163 -718 164 -704
rect 177 -773 178 -717
rect 233 -718 234 -704
rect 296 -773 297 -717
rect 317 -773 318 -717
rect 394 -718 395 -704
rect 401 -773 402 -717
rect 499 -718 500 -704
rect 516 -718 517 -704
rect 716 -718 717 -704
rect 723 -718 724 -704
rect 954 -718 955 -704
rect 121 -720 122 -704
rect 478 -773 479 -719
rect 485 -773 486 -719
rect 583 -720 584 -704
rect 639 -720 640 -704
rect 663 -773 664 -719
rect 705 -773 706 -719
rect 912 -720 913 -704
rect 919 -773 920 -719
rect 1003 -720 1004 -704
rect 93 -722 94 -704
rect 121 -773 122 -721
rect 131 -722 132 -704
rect 345 -722 346 -704
rect 352 -722 353 -704
rect 460 -722 461 -704
rect 467 -722 468 -704
rect 807 -722 808 -704
rect 870 -773 871 -721
rect 898 -722 899 -704
rect 912 -773 913 -721
rect 996 -722 997 -704
rect 1003 -773 1004 -721
rect 1045 -722 1046 -704
rect 93 -773 94 -723
rect 331 -724 332 -704
rect 338 -724 339 -704
rect 492 -773 493 -723
rect 541 -773 542 -723
rect 646 -724 647 -704
rect 653 -724 654 -704
rect 667 -773 668 -723
rect 688 -724 689 -704
rect 807 -773 808 -723
rect 877 -724 878 -704
rect 898 -773 899 -723
rect 940 -773 941 -723
rect 989 -724 990 -704
rect 996 -773 997 -723
rect 1017 -724 1018 -704
rect 135 -773 136 -725
rect 152 -773 153 -725
rect 163 -773 164 -725
rect 184 -726 185 -704
rect 205 -726 206 -704
rect 331 -773 332 -725
rect 352 -773 353 -725
rect 380 -726 381 -704
rect 457 -726 458 -704
rect 618 -726 619 -704
rect 639 -773 640 -725
rect 674 -726 675 -704
rect 688 -773 689 -725
rect 709 -726 710 -704
rect 716 -773 717 -725
rect 1052 -726 1053 -704
rect 142 -773 143 -727
rect 149 -728 150 -704
rect 173 -773 174 -727
rect 460 -773 461 -727
rect 471 -773 472 -727
rect 506 -728 507 -704
rect 513 -773 514 -727
rect 618 -773 619 -727
rect 646 -773 647 -727
rect 681 -728 682 -704
rect 709 -773 710 -727
rect 730 -728 731 -704
rect 737 -728 738 -704
rect 744 -773 745 -727
rect 747 -728 748 -704
rect 800 -773 801 -727
rect 989 -773 990 -727
rect 1094 -728 1095 -704
rect 65 -730 66 -704
rect 149 -773 150 -729
rect 184 -773 185 -729
rect 387 -730 388 -704
rect 457 -773 458 -729
rect 933 -730 934 -704
rect 37 -732 38 -704
rect 65 -773 66 -731
rect 226 -732 227 -704
rect 338 -773 339 -731
rect 359 -732 360 -704
rect 366 -732 367 -704
rect 380 -773 381 -731
rect 537 -773 538 -731
rect 544 -732 545 -704
rect 1038 -732 1039 -704
rect 30 -773 31 -733
rect 37 -773 38 -733
rect 226 -773 227 -733
rect 726 -734 727 -704
rect 730 -773 731 -733
rect 793 -734 794 -704
rect 863 -734 864 -704
rect 933 -773 934 -733
rect 233 -773 234 -735
rect 254 -736 255 -704
rect 261 -736 262 -704
rect 499 -773 500 -735
rect 506 -773 507 -735
rect 520 -736 521 -704
rect 555 -736 556 -704
rect 569 -773 570 -735
rect 583 -773 584 -735
rect 719 -773 720 -735
rect 723 -773 724 -735
rect 765 -736 766 -704
rect 775 -773 776 -735
rect 975 -736 976 -704
rect 79 -738 80 -704
rect 765 -773 766 -737
rect 786 -738 787 -704
rect 961 -738 962 -704
rect 79 -773 80 -739
rect 86 -740 87 -704
rect 240 -740 241 -704
rect 254 -773 255 -739
rect 261 -773 262 -739
rect 408 -740 409 -704
rect 464 -740 465 -704
rect 520 -773 521 -739
rect 534 -740 535 -704
rect 555 -773 556 -739
rect 562 -740 563 -704
rect 737 -773 738 -739
rect 751 -740 752 -704
rect 950 -773 951 -739
rect 954 -773 955 -739
rect 975 -773 976 -739
rect 23 -742 24 -704
rect 86 -773 87 -741
rect 240 -773 241 -741
rect 303 -742 304 -704
rect 310 -773 311 -741
rect 345 -773 346 -741
rect 362 -742 363 -704
rect 429 -742 430 -704
rect 495 -742 496 -704
rect 674 -773 675 -741
rect 681 -773 682 -741
rect 695 -742 696 -704
rect 702 -742 703 -704
rect 751 -773 752 -741
rect 758 -742 759 -704
rect 772 -773 773 -741
rect 786 -773 787 -741
rect 814 -742 815 -704
rect 856 -742 857 -704
rect 863 -773 864 -741
rect 23 -773 24 -743
rect 124 -744 125 -704
rect 219 -744 220 -704
rect 303 -773 304 -743
rect 324 -744 325 -704
rect 359 -773 360 -743
rect 387 -773 388 -743
rect 415 -744 416 -704
rect 534 -773 535 -743
rect 562 -773 563 -743
rect 597 -744 598 -704
rect 961 -773 962 -743
rect 100 -746 101 -704
rect 429 -773 430 -745
rect 597 -773 598 -745
rect 835 -746 836 -704
rect 856 -773 857 -745
rect 926 -746 927 -704
rect 100 -773 101 -747
rect 191 -748 192 -704
rect 208 -773 209 -747
rect 415 -773 416 -747
rect 653 -773 654 -747
rect 1066 -748 1067 -704
rect 107 -750 108 -704
rect 191 -773 192 -749
rect 212 -750 213 -704
rect 219 -773 220 -749
rect 275 -773 276 -749
rect 324 -773 325 -749
rect 394 -773 395 -749
rect 408 -773 409 -749
rect 548 -750 549 -704
rect 656 -773 657 -749
rect 695 -773 696 -749
rect 702 -773 703 -749
rect 1073 -750 1074 -704
rect 107 -773 108 -751
rect 247 -752 248 -704
rect 548 -773 549 -751
rect 660 -752 661 -704
rect 758 -773 759 -751
rect 1059 -752 1060 -704
rect 103 -773 104 -753
rect 247 -773 248 -753
rect 660 -773 661 -753
rect 828 -754 829 -704
rect 835 -773 836 -753
rect 982 -754 983 -704
rect 170 -756 171 -704
rect 212 -773 213 -755
rect 814 -773 815 -755
rect 905 -756 906 -704
rect 926 -773 927 -755
rect 1115 -756 1116 -704
rect 9 -758 10 -704
rect 170 -773 171 -757
rect 828 -773 829 -757
rect 842 -758 843 -704
rect 849 -758 850 -704
rect 905 -773 906 -757
rect 982 -773 983 -757
rect 1087 -758 1088 -704
rect 527 -760 528 -704
rect 842 -773 843 -759
rect 849 -773 850 -759
rect 1024 -760 1025 -704
rect 527 -773 528 -761
rect 576 -762 577 -704
rect 576 -773 577 -763
rect 611 -764 612 -704
rect 611 -773 612 -765
rect 625 -766 626 -704
rect 625 -773 626 -767
rect 632 -768 633 -704
rect 632 -773 633 -769
rect 779 -770 780 -704
rect 761 -773 762 -771
rect 779 -773 780 -771
rect 2 -860 3 -782
rect 156 -783 157 -781
rect 173 -783 174 -781
rect 467 -783 468 -781
rect 492 -783 493 -781
rect 1017 -860 1018 -782
rect 1087 -860 1088 -782
rect 1094 -860 1095 -782
rect 1108 -860 1109 -782
rect 1153 -860 1154 -782
rect 16 -860 17 -784
rect 184 -785 185 -781
rect 194 -860 195 -784
rect 394 -785 395 -781
rect 408 -785 409 -781
rect 492 -860 493 -784
rect 499 -785 500 -781
rect 663 -785 664 -781
rect 667 -785 668 -781
rect 716 -860 717 -784
rect 719 -785 720 -781
rect 744 -785 745 -781
rect 779 -785 780 -781
rect 1045 -860 1046 -784
rect 1122 -785 1123 -781
rect 1143 -860 1144 -784
rect 23 -787 24 -781
rect 138 -787 139 -781
rect 149 -860 150 -786
rect 268 -787 269 -781
rect 275 -787 276 -781
rect 275 -860 276 -786
rect 275 -787 276 -781
rect 275 -860 276 -786
rect 289 -860 290 -786
rect 345 -787 346 -781
rect 355 -860 356 -786
rect 954 -860 955 -786
rect 957 -787 958 -781
rect 996 -787 997 -781
rect 1010 -787 1011 -781
rect 1066 -860 1067 -786
rect 1139 -860 1140 -786
rect 1150 -860 1151 -786
rect 23 -860 24 -788
rect 86 -789 87 -781
rect 107 -789 108 -781
rect 327 -860 328 -788
rect 341 -860 342 -788
rect 352 -789 353 -781
rect 373 -789 374 -781
rect 373 -860 374 -788
rect 373 -789 374 -781
rect 373 -860 374 -788
rect 408 -860 409 -788
rect 481 -860 482 -788
rect 506 -789 507 -781
rect 534 -789 535 -781
rect 537 -789 538 -781
rect 632 -789 633 -781
rect 646 -789 647 -781
rect 1101 -860 1102 -788
rect 30 -860 31 -790
rect 502 -860 503 -790
rect 548 -791 549 -781
rect 667 -860 668 -790
rect 674 -791 675 -781
rect 933 -860 934 -790
rect 947 -791 948 -781
rect 1003 -791 1004 -781
rect 37 -793 38 -781
rect 37 -860 38 -792
rect 37 -793 38 -781
rect 37 -860 38 -792
rect 40 -860 41 -792
rect 618 -793 619 -781
rect 621 -793 622 -781
rect 870 -793 871 -781
rect 884 -793 885 -781
rect 1003 -860 1004 -792
rect 44 -795 45 -781
rect 44 -860 45 -794
rect 44 -795 45 -781
rect 44 -860 45 -794
rect 51 -795 52 -781
rect 170 -860 171 -794
rect 177 -795 178 -781
rect 184 -860 185 -794
rect 198 -795 199 -781
rect 205 -860 206 -794
rect 208 -795 209 -781
rect 240 -795 241 -781
rect 247 -795 248 -781
rect 506 -860 507 -794
rect 513 -795 514 -781
rect 548 -860 549 -794
rect 562 -795 563 -781
rect 618 -860 619 -794
rect 625 -795 626 -781
rect 625 -860 626 -794
rect 625 -795 626 -781
rect 625 -860 626 -794
rect 653 -795 654 -781
rect 842 -795 843 -781
rect 866 -860 867 -794
rect 1052 -860 1053 -794
rect 51 -860 52 -796
rect 460 -797 461 -781
rect 464 -797 465 -781
rect 758 -860 759 -796
rect 768 -860 769 -796
rect 1010 -860 1011 -796
rect 58 -799 59 -781
rect 530 -799 531 -781
rect 541 -799 542 -781
rect 842 -860 843 -798
rect 912 -799 913 -781
rect 996 -860 997 -798
rect 58 -860 59 -800
rect 261 -801 262 -781
rect 268 -860 269 -800
rect 450 -801 451 -781
rect 453 -860 454 -800
rect 905 -801 906 -781
rect 961 -801 962 -781
rect 1073 -860 1074 -800
rect 65 -803 66 -781
rect 100 -860 101 -802
rect 128 -803 129 -781
rect 513 -860 514 -802
rect 569 -803 570 -781
rect 569 -860 570 -802
rect 569 -803 570 -781
rect 569 -860 570 -802
rect 583 -803 584 -781
rect 583 -860 584 -802
rect 583 -803 584 -781
rect 583 -860 584 -802
rect 593 -860 594 -802
rect 1059 -860 1060 -802
rect 65 -860 66 -804
rect 72 -805 73 -781
rect 75 -860 76 -804
rect 107 -860 108 -804
rect 128 -860 129 -804
rect 226 -805 227 -781
rect 240 -860 241 -804
rect 499 -860 500 -804
rect 604 -805 605 -781
rect 632 -860 633 -804
rect 653 -860 654 -804
rect 1122 -860 1123 -804
rect 86 -860 87 -806
rect 114 -807 115 -781
rect 156 -860 157 -806
rect 324 -807 325 -781
rect 345 -860 346 -806
rect 415 -807 416 -781
rect 422 -807 423 -781
rect 450 -860 451 -806
rect 457 -807 458 -781
rect 926 -807 927 -781
rect 982 -807 983 -781
rect 1024 -860 1025 -806
rect 114 -860 115 -808
rect 296 -809 297 -781
rect 310 -860 311 -808
rect 338 -809 339 -781
rect 359 -809 360 -781
rect 464 -860 465 -808
rect 478 -809 479 -781
rect 674 -860 675 -808
rect 737 -809 738 -781
rect 1038 -860 1039 -808
rect 93 -811 94 -781
rect 296 -860 297 -810
rect 313 -811 314 -781
rect 520 -811 521 -781
rect 527 -811 528 -781
rect 982 -860 983 -810
rect 989 -811 990 -781
rect 1115 -860 1116 -810
rect 93 -860 94 -812
rect 331 -813 332 -781
rect 380 -813 381 -781
rect 527 -860 528 -812
rect 607 -860 608 -812
rect 870 -860 871 -812
rect 877 -813 878 -781
rect 989 -860 990 -812
rect 152 -815 153 -781
rect 359 -860 360 -814
rect 383 -860 384 -814
rect 534 -860 535 -814
rect 614 -860 615 -814
rect 849 -815 850 -781
rect 898 -815 899 -781
rect 905 -860 906 -814
rect 926 -860 927 -814
rect 1031 -815 1032 -781
rect 177 -860 178 -816
rect 292 -817 293 -781
rect 317 -817 318 -781
rect 415 -860 416 -816
rect 422 -860 423 -816
rect 436 -817 437 -781
rect 443 -817 444 -781
rect 590 -817 591 -781
rect 656 -817 657 -781
rect 705 -817 706 -781
rect 744 -860 745 -816
rect 936 -817 937 -781
rect 142 -819 143 -781
rect 443 -860 444 -818
rect 457 -860 458 -818
rect 485 -819 486 -781
rect 495 -819 496 -781
rect 646 -860 647 -818
rect 656 -860 657 -818
rect 947 -860 948 -818
rect 142 -860 143 -820
rect 233 -821 234 -781
rect 254 -821 255 -781
rect 331 -860 332 -820
rect 387 -821 388 -781
rect 541 -860 542 -820
rect 660 -821 661 -781
rect 1080 -860 1081 -820
rect 121 -823 122 -781
rect 254 -860 255 -822
rect 317 -860 318 -822
rect 366 -823 367 -781
rect 387 -860 388 -822
rect 429 -823 430 -781
rect 436 -860 437 -822
rect 702 -823 703 -781
rect 751 -823 752 -781
rect 849 -860 850 -822
rect 863 -823 864 -781
rect 1031 -860 1032 -822
rect 79 -825 80 -781
rect 121 -860 122 -824
rect 198 -860 199 -824
rect 212 -825 213 -781
rect 222 -860 223 -824
rect 247 -860 248 -824
rect 261 -860 262 -824
rect 366 -860 367 -824
rect 401 -825 402 -781
rect 702 -860 703 -824
rect 751 -860 752 -824
rect 940 -825 941 -781
rect 212 -860 213 -826
rect 226 -860 227 -826
rect 233 -860 234 -826
rect 446 -827 447 -781
rect 471 -827 472 -781
rect 485 -860 486 -826
rect 520 -860 521 -826
rect 775 -827 776 -781
rect 779 -860 780 -826
rect 821 -827 822 -781
rect 828 -827 829 -781
rect 877 -860 878 -826
rect 324 -860 325 -828
rect 737 -860 738 -828
rect 765 -829 766 -781
rect 961 -860 962 -828
rect 401 -860 402 -830
rect 635 -860 636 -830
rect 660 -860 661 -830
rect 681 -831 682 -781
rect 723 -831 724 -781
rect 821 -860 822 -830
rect 828 -860 829 -830
rect 975 -831 976 -781
rect 135 -833 136 -781
rect 681 -860 682 -832
rect 772 -833 773 -781
rect 912 -860 913 -832
rect 135 -860 136 -834
rect 163 -835 164 -781
rect 471 -860 472 -834
rect 611 -835 612 -781
rect 688 -835 689 -781
rect 772 -860 773 -834
rect 793 -835 794 -781
rect 919 -835 920 -781
rect 163 -860 164 -836
rect 219 -837 220 -781
rect 478 -860 479 -836
rect 597 -837 598 -781
rect 604 -860 605 -836
rect 975 -860 976 -836
rect 219 -860 220 -838
rect 303 -839 304 -781
rect 555 -839 556 -781
rect 723 -860 724 -838
rect 730 -839 731 -781
rect 793 -860 794 -838
rect 807 -839 808 -781
rect 919 -860 920 -838
rect 282 -841 283 -781
rect 303 -860 304 -840
rect 555 -860 556 -840
rect 800 -841 801 -781
rect 814 -841 815 -781
rect 898 -860 899 -840
rect 191 -843 192 -781
rect 282 -860 283 -842
rect 565 -860 566 -842
rect 765 -860 766 -842
rect 786 -843 787 -781
rect 814 -860 815 -842
rect 835 -843 836 -781
rect 884 -860 885 -842
rect 103 -845 104 -781
rect 835 -860 836 -844
rect 863 -860 864 -844
rect 968 -845 969 -781
rect 82 -860 83 -846
rect 968 -860 969 -846
rect 576 -849 577 -781
rect 597 -860 598 -848
rect 611 -860 612 -848
rect 940 -860 941 -848
rect 352 -860 353 -850
rect 576 -860 577 -850
rect 579 -860 580 -850
rect 807 -860 808 -850
rect 639 -853 640 -781
rect 688 -860 689 -852
rect 695 -853 696 -781
rect 730 -860 731 -852
rect 786 -860 787 -852
rect 856 -853 857 -781
rect 338 -860 339 -854
rect 695 -860 696 -854
rect 709 -855 710 -781
rect 800 -860 801 -854
rect 856 -860 857 -854
rect 891 -855 892 -781
rect 369 -857 370 -781
rect 891 -860 892 -856
rect 394 -860 395 -858
rect 639 -860 640 -858
rect 709 -860 710 -858
rect 796 -859 797 -781
rect 9 -961 10 -869
rect 149 -870 150 -868
rect 184 -870 185 -868
rect 184 -961 185 -869
rect 184 -870 185 -868
rect 184 -961 185 -869
rect 198 -870 199 -868
rect 219 -961 220 -869
rect 222 -870 223 -868
rect 282 -870 283 -868
rect 303 -870 304 -868
rect 303 -961 304 -869
rect 303 -870 304 -868
rect 303 -961 304 -869
rect 317 -870 318 -868
rect 432 -870 433 -868
rect 481 -870 482 -868
rect 870 -870 871 -868
rect 940 -870 941 -868
rect 940 -961 941 -869
rect 940 -870 941 -868
rect 940 -961 941 -869
rect 954 -870 955 -868
rect 954 -961 955 -869
rect 954 -870 955 -868
rect 954 -961 955 -869
rect 968 -870 969 -868
rect 968 -961 969 -869
rect 968 -870 969 -868
rect 968 -961 969 -869
rect 982 -870 983 -868
rect 1150 -961 1151 -869
rect 12 -872 13 -868
rect 380 -872 381 -868
rect 383 -872 384 -868
rect 544 -872 545 -868
rect 555 -872 556 -868
rect 1101 -872 1102 -868
rect 16 -874 17 -868
rect 152 -961 153 -873
rect 170 -874 171 -868
rect 380 -961 381 -873
rect 394 -874 395 -868
rect 912 -874 913 -868
rect 989 -874 990 -868
rect 1101 -961 1102 -873
rect 30 -876 31 -868
rect 429 -876 430 -868
rect 492 -876 493 -868
rect 579 -876 580 -868
rect 583 -876 584 -868
rect 653 -961 654 -875
rect 768 -876 769 -868
rect 1031 -876 1032 -868
rect 1052 -876 1053 -868
rect 1157 -961 1158 -875
rect 30 -961 31 -877
rect 75 -878 76 -868
rect 79 -878 80 -868
rect 765 -961 766 -877
rect 779 -878 780 -868
rect 870 -961 871 -877
rect 912 -961 913 -877
rect 933 -878 934 -868
rect 1017 -878 1018 -868
rect 1129 -878 1130 -868
rect 44 -880 45 -868
rect 44 -961 45 -879
rect 44 -880 45 -868
rect 44 -961 45 -879
rect 58 -880 59 -868
rect 446 -961 447 -879
rect 478 -961 479 -879
rect 492 -961 493 -879
rect 537 -961 538 -879
rect 919 -880 920 -868
rect 933 -961 934 -879
rect 947 -880 948 -868
rect 1087 -880 1088 -868
rect 1094 -961 1095 -879
rect 1097 -880 1098 -868
rect 1143 -880 1144 -868
rect 16 -961 17 -881
rect 58 -961 59 -881
rect 65 -882 66 -868
rect 82 -882 83 -868
rect 93 -882 94 -868
rect 502 -961 503 -881
rect 565 -882 566 -868
rect 702 -882 703 -868
rect 709 -882 710 -868
rect 1052 -961 1053 -881
rect 1115 -882 1116 -868
rect 1129 -961 1130 -881
rect 72 -884 73 -868
rect 1136 -884 1137 -868
rect 75 -961 76 -885
rect 86 -886 87 -868
rect 93 -961 94 -885
rect 156 -886 157 -868
rect 170 -961 171 -885
rect 453 -886 454 -868
rect 572 -961 573 -885
rect 821 -886 822 -868
rect 856 -886 857 -868
rect 982 -961 983 -885
rect 1108 -886 1109 -868
rect 1115 -961 1116 -885
rect 79 -961 80 -887
rect 548 -888 549 -868
rect 576 -888 577 -868
rect 1087 -961 1088 -887
rect 1108 -961 1109 -887
rect 1122 -888 1123 -868
rect 86 -961 87 -889
rect 128 -890 129 -868
rect 135 -890 136 -868
rect 191 -890 192 -868
rect 198 -961 199 -889
rect 205 -890 206 -868
rect 229 -890 230 -868
rect 555 -961 556 -889
rect 562 -890 563 -868
rect 1122 -961 1123 -889
rect 51 -892 52 -868
rect 128 -961 129 -891
rect 135 -961 136 -891
rect 268 -892 269 -868
rect 275 -892 276 -868
rect 275 -961 276 -891
rect 275 -892 276 -868
rect 275 -961 276 -891
rect 310 -892 311 -868
rect 317 -961 318 -891
rect 324 -892 325 -868
rect 499 -892 500 -868
rect 548 -961 549 -891
rect 698 -961 699 -891
rect 730 -892 731 -868
rect 821 -961 822 -891
rect 905 -892 906 -868
rect 1143 -961 1144 -891
rect 51 -961 52 -893
rect 415 -894 416 -868
rect 418 -961 419 -893
rect 1038 -894 1039 -868
rect 82 -961 83 -895
rect 191 -961 192 -895
rect 261 -961 262 -895
rect 579 -961 580 -895
rect 590 -896 591 -868
rect 1073 -896 1074 -868
rect 114 -898 115 -868
rect 355 -898 356 -868
rect 359 -898 360 -868
rect 369 -942 370 -897
rect 394 -961 395 -897
rect 422 -898 423 -868
rect 439 -961 440 -897
rect 1031 -961 1032 -897
rect 1073 -961 1074 -897
rect 1080 -898 1081 -868
rect 114 -961 115 -899
rect 240 -900 241 -868
rect 268 -961 269 -899
rect 299 -961 300 -899
rect 310 -961 311 -899
rect 614 -900 615 -868
rect 635 -900 636 -868
rect 1003 -900 1004 -868
rect 1010 -900 1011 -868
rect 1038 -961 1039 -899
rect 142 -902 143 -868
rect 226 -902 227 -868
rect 240 -961 241 -901
rect 345 -902 346 -868
rect 359 -961 360 -901
rect 751 -902 752 -868
rect 758 -902 759 -868
rect 779 -961 780 -901
rect 891 -902 892 -868
rect 905 -961 906 -901
rect 919 -961 920 -901
rect 926 -902 927 -868
rect 947 -961 948 -901
rect 1024 -902 1025 -868
rect 142 -961 143 -903
rect 212 -904 213 -868
rect 226 -961 227 -903
rect 450 -904 451 -868
rect 562 -961 563 -903
rect 597 -904 598 -868
rect 604 -904 605 -868
rect 1017 -961 1018 -903
rect 149 -961 150 -905
rect 583 -961 584 -905
rect 604 -961 605 -905
rect 618 -906 619 -868
rect 639 -906 640 -868
rect 863 -961 864 -905
rect 898 -906 899 -868
rect 926 -961 927 -905
rect 961 -906 962 -868
rect 1010 -961 1011 -905
rect 156 -961 157 -907
rect 401 -908 402 -868
rect 408 -908 409 -868
rect 429 -961 430 -907
rect 443 -908 444 -868
rect 709 -961 710 -907
rect 723 -908 724 -868
rect 730 -961 731 -907
rect 751 -961 752 -907
rect 828 -908 829 -868
rect 961 -961 962 -907
rect 975 -908 976 -868
rect 996 -908 997 -868
rect 1003 -961 1004 -907
rect 163 -910 164 -868
rect 212 -961 213 -909
rect 254 -910 255 -868
rect 597 -961 598 -909
rect 611 -910 612 -868
rect 660 -910 661 -868
rect 674 -910 675 -868
rect 1080 -961 1081 -909
rect 121 -912 122 -868
rect 254 -961 255 -911
rect 324 -961 325 -911
rect 506 -912 507 -868
rect 534 -912 535 -868
rect 618 -961 619 -911
rect 625 -912 626 -868
rect 674 -961 675 -911
rect 695 -912 696 -868
rect 702 -961 703 -911
rect 716 -912 717 -868
rect 723 -961 724 -911
rect 793 -912 794 -868
rect 1024 -961 1025 -911
rect 2 -914 3 -868
rect 793 -961 794 -913
rect 807 -914 808 -868
rect 828 -961 829 -913
rect 884 -914 885 -868
rect 975 -961 976 -913
rect 100 -916 101 -868
rect 121 -961 122 -915
rect 163 -961 164 -915
rect 415 -961 416 -915
rect 443 -961 444 -915
rect 989 -961 990 -915
rect 65 -961 66 -917
rect 100 -961 101 -917
rect 177 -918 178 -868
rect 205 -961 206 -917
rect 331 -918 332 -868
rect 397 -918 398 -868
rect 408 -961 409 -917
rect 457 -918 458 -868
rect 481 -961 482 -917
rect 639 -961 640 -917
rect 646 -918 647 -868
rect 660 -961 661 -917
rect 716 -961 717 -917
rect 800 -918 801 -868
rect 807 -961 808 -917
rect 835 -918 836 -868
rect 877 -918 878 -868
rect 884 -961 885 -917
rect 289 -920 290 -868
rect 331 -961 332 -919
rect 338 -920 339 -868
rect 527 -920 528 -868
rect 541 -920 542 -868
rect 996 -961 997 -919
rect 107 -922 108 -868
rect 338 -961 339 -921
rect 341 -922 342 -868
rect 422 -961 423 -921
rect 450 -961 451 -921
rect 485 -922 486 -868
rect 506 -961 507 -921
rect 1059 -922 1060 -868
rect 107 -961 108 -923
rect 194 -924 195 -868
rect 289 -961 290 -923
rect 436 -924 437 -868
rect 457 -961 458 -923
rect 688 -924 689 -868
rect 814 -924 815 -868
rect 835 -961 836 -923
rect 849 -924 850 -868
rect 877 -961 878 -923
rect 1059 -961 1060 -923
rect 1066 -924 1067 -868
rect 72 -961 73 -925
rect 1066 -961 1067 -925
rect 345 -961 346 -927
rect 464 -928 465 -868
rect 471 -928 472 -868
rect 814 -961 815 -927
rect 352 -930 353 -868
rect 646 -961 647 -929
rect 688 -961 689 -929
rect 786 -930 787 -868
rect 362 -961 363 -931
rect 401 -961 402 -931
rect 464 -961 465 -931
rect 527 -961 528 -931
rect 541 -961 542 -931
rect 1045 -932 1046 -868
rect 366 -934 367 -868
rect 576 -961 577 -933
rect 593 -934 594 -868
rect 800 -961 801 -933
rect 352 -961 353 -935
rect 593 -961 594 -935
rect 614 -961 615 -935
rect 758 -961 759 -935
rect 366 -961 367 -937
rect 373 -938 374 -868
rect 485 -961 486 -937
rect 558 -938 559 -868
rect 569 -938 570 -868
rect 891 -961 892 -937
rect 177 -961 178 -939
rect 569 -961 570 -939
rect 621 -961 622 -939
rect 1045 -961 1046 -939
rect 471 -961 472 -941
rect 513 -942 514 -868
rect 849 -961 850 -941
rect 373 -961 374 -943
rect 544 -961 545 -943
rect 625 -961 626 -943
rect 842 -944 843 -868
rect 513 -961 514 -945
rect 520 -946 521 -868
rect 632 -946 633 -868
rect 898 -961 899 -945
rect 23 -948 24 -868
rect 520 -961 521 -947
rect 632 -961 633 -947
rect 1136 -961 1137 -947
rect 23 -961 24 -949
rect 387 -950 388 -868
rect 681 -950 682 -868
rect 842 -961 843 -949
rect 247 -952 248 -868
rect 387 -961 388 -951
rect 667 -952 668 -868
rect 681 -961 682 -951
rect 744 -952 745 -868
rect 786 -961 787 -951
rect 233 -954 234 -868
rect 247 -961 248 -953
rect 667 -961 668 -953
rect 772 -954 773 -868
rect 233 -961 234 -955
rect 296 -956 297 -868
rect 691 -961 692 -955
rect 772 -961 773 -955
rect 737 -958 738 -868
rect 744 -961 745 -957
rect 37 -961 38 -959
rect 737 -961 738 -959
rect 9 -971 10 -969
rect 282 -971 283 -969
rect 285 -971 286 -969
rect 310 -971 311 -969
rect 359 -1076 360 -970
rect 726 -1076 727 -970
rect 859 -971 860 -969
rect 961 -971 962 -969
rect 9 -1076 10 -972
rect 485 -973 486 -969
rect 541 -1076 542 -972
rect 1136 -973 1137 -969
rect 16 -975 17 -969
rect 597 -975 598 -969
rect 607 -1076 608 -974
rect 905 -975 906 -969
rect 16 -1076 17 -976
rect 166 -1076 167 -976
rect 184 -977 185 -969
rect 184 -1076 185 -976
rect 184 -977 185 -969
rect 184 -1076 185 -976
rect 194 -1076 195 -976
rect 380 -977 381 -969
rect 401 -977 402 -969
rect 464 -1076 465 -976
rect 467 -977 468 -969
rect 765 -977 766 -969
rect 23 -979 24 -969
rect 436 -979 437 -969
rect 439 -979 440 -969
rect 688 -1076 689 -978
rect 691 -979 692 -969
rect 961 -1076 962 -978
rect 23 -1076 24 -980
rect 390 -1076 391 -980
rect 436 -1076 437 -980
rect 558 -1076 559 -980
rect 569 -981 570 -969
rect 1115 -981 1116 -969
rect 30 -983 31 -969
rect 33 -987 34 -982
rect 37 -983 38 -969
rect 254 -983 255 -969
rect 271 -1076 272 -982
rect 324 -983 325 -969
rect 362 -983 363 -969
rect 628 -983 629 -969
rect 632 -1076 633 -982
rect 982 -983 983 -969
rect 30 -1076 31 -984
rect 653 -985 654 -969
rect 695 -1076 696 -984
rect 828 -985 829 -969
rect 982 -1076 983 -984
rect 1045 -985 1046 -969
rect 653 -1076 654 -986
rect 698 -987 699 -969
rect 1052 -987 1053 -969
rect 37 -1076 38 -988
rect 44 -989 45 -969
rect 65 -989 66 -969
rect 933 -989 934 -969
rect 1045 -1076 1046 -988
rect 1073 -989 1074 -969
rect 44 -1076 45 -990
rect 527 -991 528 -969
rect 569 -1076 570 -990
rect 926 -991 927 -969
rect 933 -1076 934 -990
rect 996 -991 997 -969
rect 1052 -1076 1053 -990
rect 1101 -991 1102 -969
rect 2 -993 3 -969
rect 926 -1076 927 -992
rect 68 -995 69 -969
rect 415 -995 416 -969
rect 422 -995 423 -969
rect 527 -1076 528 -994
rect 576 -1076 577 -994
rect 674 -995 675 -969
rect 786 -995 787 -969
rect 1073 -1076 1074 -994
rect 68 -1076 69 -996
rect 338 -997 339 -969
rect 380 -1076 381 -996
rect 513 -997 514 -969
rect 579 -997 580 -969
rect 1024 -997 1025 -969
rect 72 -999 73 -969
rect 86 -999 87 -969
rect 114 -999 115 -969
rect 401 -1076 402 -998
rect 415 -1076 416 -998
rect 520 -999 521 -969
rect 590 -999 591 -969
rect 667 -999 668 -969
rect 674 -1076 675 -998
rect 779 -999 780 -969
rect 786 -1076 787 -998
rect 912 -999 913 -969
rect 1024 -1076 1025 -998
rect 1122 -999 1123 -969
rect 72 -1076 73 -1000
rect 93 -1001 94 -969
rect 114 -1076 115 -1000
rect 275 -1001 276 -969
rect 282 -1076 283 -1000
rect 709 -1001 710 -969
rect 779 -1076 780 -1000
rect 940 -1001 941 -969
rect 82 -1003 83 -969
rect 555 -1003 556 -969
rect 590 -1076 591 -1002
rect 681 -1003 682 -969
rect 709 -1076 710 -1002
rect 863 -1003 864 -969
rect 912 -1076 913 -1002
rect 1031 -1003 1032 -969
rect 82 -1076 83 -1004
rect 793 -1005 794 -969
rect 842 -1005 843 -969
rect 940 -1076 941 -1004
rect 1010 -1005 1011 -969
rect 1031 -1076 1032 -1004
rect 86 -1076 87 -1006
rect 205 -1007 206 -969
rect 219 -1007 220 -969
rect 219 -1076 220 -1006
rect 219 -1007 220 -969
rect 219 -1076 220 -1006
rect 229 -1076 230 -1006
rect 233 -1007 234 -969
rect 240 -1007 241 -969
rect 506 -1007 507 -969
rect 513 -1076 514 -1006
rect 604 -1007 605 -969
rect 614 -1007 615 -969
rect 716 -1007 717 -969
rect 793 -1076 794 -1006
rect 884 -1007 885 -969
rect 1010 -1076 1011 -1006
rect 1041 -1076 1042 -1006
rect 93 -1076 94 -1008
rect 107 -1009 108 -969
rect 135 -1009 136 -969
rect 418 -1009 419 -969
rect 443 -1076 444 -1008
rect 450 -1009 451 -969
rect 471 -1009 472 -969
rect 681 -1076 682 -1008
rect 716 -1076 717 -1008
rect 821 -1009 822 -969
rect 842 -1076 843 -1008
rect 898 -1009 899 -969
rect 58 -1011 59 -969
rect 821 -1076 822 -1010
rect 863 -1076 864 -1010
rect 968 -1011 969 -969
rect 58 -1076 59 -1012
rect 75 -1013 76 -969
rect 107 -1076 108 -1012
rect 121 -1013 122 -969
rect 135 -1076 136 -1012
rect 226 -1013 227 -969
rect 233 -1076 234 -1012
rect 429 -1013 430 -969
rect 450 -1076 451 -1012
rect 702 -1013 703 -969
rect 884 -1076 885 -1012
rect 975 -1013 976 -969
rect 121 -1076 122 -1014
rect 163 -1015 164 -969
rect 191 -1015 192 -969
rect 422 -1076 423 -1014
rect 471 -1076 472 -1014
rect 488 -1076 489 -1014
rect 492 -1015 493 -969
rect 506 -1076 507 -1014
rect 520 -1076 521 -1014
rect 544 -1015 545 -969
rect 548 -1015 549 -969
rect 702 -1076 703 -1014
rect 898 -1076 899 -1014
rect 1017 -1015 1018 -969
rect 149 -1076 150 -1016
rect 212 -1017 213 -969
rect 240 -1076 241 -1016
rect 457 -1017 458 -969
rect 474 -1017 475 -969
rect 1017 -1076 1018 -1016
rect 163 -1076 164 -1018
rect 205 -1076 206 -1018
rect 254 -1076 255 -1018
rect 740 -1076 741 -1018
rect 947 -1019 948 -969
rect 968 -1076 969 -1018
rect 975 -1076 976 -1018
rect 1038 -1019 1039 -969
rect 191 -1076 192 -1020
rect 296 -1076 297 -1020
rect 303 -1021 304 -969
rect 548 -1076 549 -1020
rect 555 -1076 556 -1020
rect 807 -1021 808 -969
rect 856 -1021 857 -969
rect 947 -1076 948 -1020
rect 177 -1023 178 -969
rect 303 -1076 304 -1022
rect 306 -1023 307 -969
rect 583 -1023 584 -969
rect 593 -1023 594 -969
rect 1080 -1023 1081 -969
rect 177 -1076 178 -1024
rect 373 -1025 374 -969
rect 408 -1025 409 -969
rect 429 -1076 430 -1024
rect 446 -1025 447 -969
rect 807 -1076 808 -1024
rect 1080 -1076 1081 -1024
rect 1094 -1025 1095 -969
rect 268 -1027 269 -969
rect 324 -1076 325 -1026
rect 331 -1027 332 -969
rect 373 -1076 374 -1026
rect 408 -1076 409 -1026
rect 492 -1076 493 -1026
rect 502 -1027 503 -969
rect 996 -1076 997 -1026
rect 142 -1029 143 -969
rect 268 -1076 269 -1028
rect 275 -1076 276 -1028
rect 394 -1029 395 -969
rect 457 -1076 458 -1028
rect 737 -1029 738 -969
rect 51 -1031 52 -969
rect 394 -1076 395 -1030
rect 478 -1031 479 -969
rect 1087 -1031 1088 -969
rect 2 -1076 3 -1032
rect 51 -1076 52 -1032
rect 100 -1033 101 -969
rect 142 -1076 143 -1032
rect 156 -1033 157 -969
rect 478 -1076 479 -1032
rect 481 -1033 482 -969
rect 814 -1033 815 -969
rect 156 -1076 157 -1034
rect 247 -1035 248 -969
rect 289 -1035 290 -969
rect 331 -1076 332 -1034
rect 338 -1076 339 -1034
rect 397 -1076 398 -1034
rect 583 -1076 584 -1034
rect 891 -1035 892 -969
rect 247 -1076 248 -1036
rect 317 -1037 318 -969
rect 600 -1076 601 -1036
rect 765 -1076 766 -1036
rect 891 -1076 892 -1036
rect 1003 -1037 1004 -969
rect 289 -1076 290 -1038
rect 345 -1039 346 -969
rect 618 -1039 619 -969
rect 828 -1076 829 -1038
rect 1003 -1076 1004 -1038
rect 1066 -1039 1067 -969
rect 261 -1041 262 -969
rect 345 -1076 346 -1040
rect 562 -1041 563 -969
rect 618 -1076 619 -1040
rect 621 -1041 622 -969
rect 870 -1041 871 -969
rect 919 -1041 920 -969
rect 1066 -1076 1067 -1040
rect 261 -1076 262 -1042
rect 352 -1043 353 -969
rect 499 -1043 500 -969
rect 919 -1076 920 -1042
rect 310 -1076 311 -1044
rect 387 -1045 388 -969
rect 562 -1076 563 -1044
rect 572 -1045 573 -969
rect 635 -1045 636 -969
rect 751 -1045 752 -969
rect 870 -1076 871 -1044
rect 989 -1045 990 -969
rect 317 -1076 318 -1046
rect 534 -1047 535 -969
rect 572 -1076 573 -1046
rect 905 -1076 906 -1046
rect 989 -1076 990 -1046
rect 1108 -1047 1109 -969
rect 352 -1076 353 -1048
rect 366 -1049 367 -969
rect 387 -1076 388 -1048
rect 639 -1049 640 -969
rect 667 -1076 668 -1048
rect 772 -1049 773 -969
rect 128 -1051 129 -969
rect 366 -1076 367 -1050
rect 495 -1076 496 -1050
rect 639 -1076 640 -1050
rect 737 -1076 738 -1050
rect 1129 -1051 1130 -969
rect 128 -1076 129 -1052
rect 170 -1053 171 -969
rect 534 -1076 535 -1052
rect 646 -1053 647 -969
rect 751 -1076 752 -1052
rect 835 -1053 836 -969
rect 1129 -1076 1130 -1052
rect 1157 -1053 1158 -969
rect 170 -1076 171 -1054
rect 198 -1055 199 -969
rect 611 -1055 612 -969
rect 646 -1076 647 -1054
rect 800 -1055 801 -969
rect 835 -1076 836 -1054
rect 198 -1076 199 -1056
rect 849 -1057 850 -969
rect 611 -1076 612 -1058
rect 723 -1059 724 -969
rect 744 -1059 745 -969
rect 800 -1076 801 -1058
rect 849 -1076 850 -1058
rect 954 -1059 955 -969
rect 625 -1061 626 -969
rect 772 -1076 773 -1060
rect 954 -1076 955 -1060
rect 1059 -1061 1060 -969
rect 502 -1076 503 -1062
rect 625 -1076 626 -1062
rect 635 -1076 636 -1062
rect 856 -1076 857 -1062
rect 723 -1076 724 -1064
rect 1143 -1065 1144 -969
rect 730 -1067 731 -969
rect 744 -1076 745 -1066
rect 1143 -1076 1144 -1066
rect 1150 -1067 1151 -969
rect 660 -1069 661 -969
rect 730 -1076 731 -1068
rect 660 -1076 661 -1070
rect 758 -1071 759 -969
rect 758 -1076 759 -1072
rect 877 -1073 878 -969
rect 604 -1076 605 -1074
rect 877 -1076 878 -1074
rect 5 -1165 6 -1085
rect 348 -1165 349 -1085
rect 366 -1086 367 -1084
rect 369 -1106 370 -1085
rect 390 -1086 391 -1084
rect 898 -1086 899 -1084
rect 947 -1086 948 -1084
rect 1038 -1086 1039 -1084
rect 1041 -1086 1042 -1084
rect 1066 -1086 1067 -1084
rect 1076 -1165 1077 -1085
rect 1080 -1086 1081 -1084
rect 1122 -1165 1123 -1085
rect 1129 -1086 1130 -1084
rect 1143 -1086 1144 -1084
rect 1150 -1165 1151 -1085
rect 9 -1088 10 -1084
rect 467 -1165 468 -1087
rect 488 -1088 489 -1084
rect 520 -1088 521 -1084
rect 523 -1165 524 -1087
rect 828 -1088 829 -1084
rect 905 -1088 906 -1084
rect 947 -1165 948 -1087
rect 968 -1088 969 -1084
rect 968 -1165 969 -1087
rect 968 -1088 969 -1084
rect 968 -1165 969 -1087
rect 996 -1088 997 -1084
rect 1059 -1088 1060 -1084
rect 9 -1165 10 -1089
rect 30 -1090 31 -1084
rect 40 -1165 41 -1089
rect 898 -1165 899 -1089
rect 982 -1090 983 -1084
rect 996 -1165 997 -1089
rect 1031 -1090 1032 -1084
rect 1066 -1165 1067 -1089
rect 16 -1092 17 -1084
rect 495 -1092 496 -1084
rect 506 -1092 507 -1084
rect 506 -1165 507 -1091
rect 506 -1092 507 -1084
rect 506 -1165 507 -1091
rect 513 -1092 514 -1084
rect 691 -1165 692 -1091
rect 723 -1165 724 -1091
rect 751 -1092 752 -1084
rect 779 -1092 780 -1084
rect 828 -1165 829 -1091
rect 856 -1092 857 -1084
rect 905 -1165 906 -1091
rect 926 -1092 927 -1084
rect 982 -1165 983 -1091
rect 1017 -1092 1018 -1084
rect 1031 -1165 1032 -1091
rect 1045 -1092 1046 -1084
rect 1045 -1165 1046 -1091
rect 1045 -1092 1046 -1084
rect 1045 -1165 1046 -1091
rect 1052 -1092 1053 -1084
rect 1052 -1165 1053 -1091
rect 1052 -1092 1053 -1084
rect 1052 -1165 1053 -1091
rect 51 -1094 52 -1084
rect 58 -1094 59 -1084
rect 61 -1165 62 -1093
rect 198 -1094 199 -1084
rect 212 -1094 213 -1084
rect 800 -1094 801 -1084
rect 817 -1094 818 -1084
rect 954 -1094 955 -1084
rect 1010 -1094 1011 -1084
rect 1017 -1165 1018 -1093
rect 51 -1165 52 -1095
rect 275 -1096 276 -1084
rect 324 -1096 325 -1084
rect 408 -1096 409 -1084
rect 418 -1165 419 -1095
rect 989 -1096 990 -1084
rect 1003 -1096 1004 -1084
rect 1010 -1165 1011 -1095
rect 65 -1098 66 -1084
rect 156 -1098 157 -1084
rect 166 -1098 167 -1084
rect 702 -1098 703 -1084
rect 740 -1165 741 -1097
rect 779 -1165 780 -1097
rect 789 -1165 790 -1097
rect 863 -1098 864 -1084
rect 926 -1165 927 -1097
rect 933 -1098 934 -1084
rect 940 -1098 941 -1084
rect 1003 -1165 1004 -1097
rect 65 -1165 66 -1099
rect 72 -1100 73 -1084
rect 79 -1100 80 -1084
rect 205 -1100 206 -1084
rect 212 -1165 213 -1099
rect 219 -1100 220 -1084
rect 268 -1165 269 -1099
rect 331 -1100 332 -1084
rect 366 -1165 367 -1099
rect 394 -1100 395 -1084
rect 397 -1100 398 -1084
rect 443 -1100 444 -1084
rect 450 -1100 451 -1084
rect 513 -1165 514 -1099
rect 527 -1100 528 -1084
rect 635 -1100 636 -1084
rect 639 -1100 640 -1084
rect 702 -1165 703 -1099
rect 751 -1165 752 -1099
rect 814 -1100 815 -1084
rect 835 -1100 836 -1084
rect 856 -1165 857 -1099
rect 870 -1100 871 -1084
rect 940 -1165 941 -1099
rect 975 -1100 976 -1084
rect 989 -1165 990 -1099
rect 68 -1102 69 -1084
rect 502 -1102 503 -1084
rect 541 -1102 542 -1084
rect 954 -1165 955 -1101
rect 79 -1165 80 -1103
rect 93 -1104 94 -1084
rect 100 -1104 101 -1084
rect 107 -1165 108 -1103
rect 114 -1104 115 -1084
rect 198 -1165 199 -1103
rect 205 -1165 206 -1103
rect 261 -1104 262 -1084
rect 324 -1165 325 -1103
rect 1038 -1165 1039 -1103
rect 93 -1165 94 -1105
rect 285 -1106 286 -1084
rect 331 -1165 332 -1105
rect 352 -1106 353 -1084
rect 394 -1165 395 -1105
rect 401 -1106 402 -1084
rect 520 -1165 521 -1105
rect 544 -1106 545 -1084
rect 821 -1106 822 -1084
rect 835 -1165 836 -1105
rect 842 -1106 843 -1084
rect 884 -1106 885 -1084
rect 933 -1165 934 -1105
rect 72 -1165 73 -1107
rect 352 -1165 353 -1107
rect 355 -1165 356 -1107
rect 821 -1165 822 -1107
rect 842 -1165 843 -1107
rect 1041 -1165 1042 -1107
rect 100 -1165 101 -1109
rect 142 -1110 143 -1084
rect 149 -1110 150 -1084
rect 156 -1165 157 -1109
rect 170 -1110 171 -1084
rect 219 -1165 220 -1109
rect 254 -1110 255 -1084
rect 401 -1165 402 -1109
rect 415 -1110 416 -1084
rect 443 -1165 444 -1109
rect 450 -1165 451 -1109
rect 737 -1110 738 -1084
rect 765 -1110 766 -1084
rect 800 -1165 801 -1109
rect 919 -1110 920 -1084
rect 975 -1165 976 -1109
rect 23 -1112 24 -1084
rect 170 -1165 171 -1111
rect 177 -1112 178 -1084
rect 411 -1165 412 -1111
rect 422 -1112 423 -1084
rect 527 -1165 528 -1111
rect 555 -1112 556 -1084
rect 744 -1112 745 -1084
rect 765 -1165 766 -1111
rect 1073 -1112 1074 -1084
rect 23 -1165 24 -1113
rect 37 -1114 38 -1084
rect 103 -1114 104 -1084
rect 688 -1114 689 -1084
rect 744 -1165 745 -1113
rect 758 -1114 759 -1084
rect 772 -1114 773 -1084
rect 884 -1165 885 -1113
rect 891 -1114 892 -1084
rect 919 -1165 920 -1113
rect 114 -1165 115 -1115
rect 128 -1116 129 -1084
rect 152 -1165 153 -1115
rect 313 -1165 314 -1115
rect 383 -1165 384 -1115
rect 1059 -1165 1060 -1115
rect 177 -1165 178 -1117
rect 303 -1118 304 -1084
rect 429 -1118 430 -1084
rect 429 -1165 430 -1117
rect 429 -1118 430 -1084
rect 429 -1165 430 -1117
rect 436 -1118 437 -1084
rect 541 -1165 542 -1117
rect 555 -1165 556 -1117
rect 1024 -1118 1025 -1084
rect 184 -1120 185 -1084
rect 261 -1165 262 -1119
rect 296 -1120 297 -1084
rect 422 -1165 423 -1119
rect 492 -1165 493 -1119
rect 733 -1165 734 -1119
rect 793 -1120 794 -1084
rect 793 -1165 794 -1119
rect 793 -1120 794 -1084
rect 793 -1165 794 -1119
rect 891 -1165 892 -1119
rect 912 -1120 913 -1084
rect 121 -1122 122 -1084
rect 296 -1165 297 -1121
rect 303 -1165 304 -1121
rect 345 -1122 346 -1084
rect 380 -1122 381 -1084
rect 436 -1165 437 -1121
rect 499 -1122 500 -1084
rect 863 -1165 864 -1121
rect 877 -1122 878 -1084
rect 912 -1165 913 -1121
rect 30 -1165 31 -1123
rect 345 -1165 346 -1123
rect 373 -1124 374 -1084
rect 380 -1165 381 -1123
rect 499 -1165 500 -1123
rect 1073 -1165 1074 -1123
rect 44 -1126 45 -1084
rect 373 -1165 374 -1125
rect 502 -1165 503 -1125
rect 786 -1126 787 -1084
rect 44 -1165 45 -1127
rect 572 -1128 573 -1084
rect 576 -1128 577 -1084
rect 597 -1128 598 -1084
rect 607 -1128 608 -1084
rect 618 -1128 619 -1084
rect 632 -1128 633 -1084
rect 758 -1165 759 -1127
rect 110 -1130 111 -1084
rect 877 -1165 878 -1129
rect 121 -1165 122 -1131
rect 289 -1132 290 -1084
rect 387 -1132 388 -1084
rect 632 -1165 633 -1131
rect 639 -1165 640 -1131
rect 709 -1132 710 -1084
rect 163 -1165 164 -1133
rect 289 -1165 290 -1133
rect 481 -1165 482 -1133
rect 786 -1165 787 -1133
rect 184 -1165 185 -1135
rect 408 -1165 409 -1135
rect 565 -1165 566 -1135
rect 814 -1165 815 -1135
rect 191 -1138 192 -1084
rect 275 -1165 276 -1137
rect 569 -1165 570 -1137
rect 611 -1138 612 -1084
rect 618 -1165 619 -1137
rect 646 -1138 647 -1084
rect 653 -1138 654 -1084
rect 772 -1165 773 -1137
rect 86 -1140 87 -1084
rect 191 -1165 192 -1139
rect 215 -1140 216 -1084
rect 485 -1140 486 -1084
rect 558 -1140 559 -1084
rect 646 -1165 647 -1139
rect 667 -1140 668 -1084
rect 667 -1165 668 -1139
rect 667 -1140 668 -1084
rect 667 -1165 668 -1139
rect 684 -1140 685 -1084
rect 961 -1140 962 -1084
rect 86 -1165 87 -1141
rect 317 -1142 318 -1084
rect 415 -1165 416 -1141
rect 611 -1165 612 -1141
rect 709 -1165 710 -1141
rect 716 -1142 717 -1084
rect 849 -1142 850 -1084
rect 961 -1165 962 -1141
rect 54 -1144 55 -1084
rect 716 -1165 717 -1143
rect 807 -1144 808 -1084
rect 849 -1165 850 -1143
rect 128 -1165 129 -1145
rect 558 -1165 559 -1145
rect 583 -1146 584 -1084
rect 681 -1146 682 -1084
rect 226 -1148 227 -1084
rect 387 -1165 388 -1147
rect 471 -1148 472 -1084
rect 681 -1165 682 -1147
rect 135 -1150 136 -1084
rect 226 -1165 227 -1149
rect 240 -1150 241 -1084
rect 576 -1165 577 -1149
rect 586 -1150 587 -1084
rect 870 -1165 871 -1149
rect 135 -1165 136 -1151
rect 534 -1152 535 -1084
rect 562 -1152 563 -1084
rect 583 -1165 584 -1151
rect 590 -1152 591 -1084
rect 590 -1165 591 -1151
rect 590 -1152 591 -1084
rect 590 -1165 591 -1151
rect 604 -1152 605 -1084
rect 653 -1165 654 -1151
rect 240 -1165 241 -1153
rect 338 -1154 339 -1084
rect 457 -1154 458 -1084
rect 471 -1165 472 -1153
rect 478 -1154 479 -1084
rect 485 -1165 486 -1153
rect 534 -1165 535 -1153
rect 695 -1154 696 -1084
rect 247 -1156 248 -1084
rect 254 -1165 255 -1155
rect 310 -1156 311 -1084
rect 338 -1165 339 -1155
rect 359 -1156 360 -1084
rect 457 -1165 458 -1155
rect 548 -1156 549 -1084
rect 604 -1165 605 -1155
rect 625 -1156 626 -1084
rect 807 -1165 808 -1155
rect 233 -1158 234 -1084
rect 247 -1165 248 -1157
rect 317 -1165 318 -1157
rect 464 -1158 465 -1084
rect 548 -1165 549 -1157
rect 660 -1158 661 -1084
rect 674 -1158 675 -1084
rect 695 -1165 696 -1157
rect 37 -1165 38 -1159
rect 233 -1165 234 -1159
rect 282 -1165 283 -1159
rect 674 -1165 675 -1159
rect 464 -1165 465 -1161
rect 625 -1165 626 -1161
rect 660 -1165 661 -1161
rect 730 -1162 731 -1084
rect 730 -1165 731 -1163
rect 1024 -1165 1025 -1163
rect 2 -1248 3 -1174
rect 145 -1175 146 -1173
rect 149 -1248 150 -1174
rect 205 -1175 206 -1173
rect 226 -1175 227 -1173
rect 310 -1175 311 -1173
rect 313 -1175 314 -1173
rect 821 -1175 822 -1173
rect 835 -1175 836 -1173
rect 835 -1248 836 -1174
rect 835 -1175 836 -1173
rect 835 -1248 836 -1174
rect 982 -1175 983 -1173
rect 1073 -1248 1074 -1174
rect 1115 -1248 1116 -1174
rect 1122 -1175 1123 -1173
rect 1129 -1248 1130 -1174
rect 1157 -1248 1158 -1174
rect 16 -1177 17 -1173
rect 275 -1177 276 -1173
rect 303 -1177 304 -1173
rect 408 -1248 409 -1176
rect 460 -1248 461 -1176
rect 471 -1177 472 -1173
rect 485 -1177 486 -1173
rect 488 -1205 489 -1176
rect 506 -1177 507 -1173
rect 520 -1248 521 -1176
rect 558 -1177 559 -1173
rect 695 -1177 696 -1173
rect 730 -1177 731 -1173
rect 933 -1177 934 -1173
rect 989 -1177 990 -1173
rect 1080 -1248 1081 -1176
rect 1150 -1177 1151 -1173
rect 1164 -1248 1165 -1176
rect 16 -1248 17 -1178
rect 380 -1179 381 -1173
rect 383 -1179 384 -1173
rect 478 -1179 479 -1173
rect 485 -1248 486 -1178
rect 604 -1179 605 -1173
rect 653 -1179 654 -1173
rect 730 -1248 731 -1178
rect 751 -1179 752 -1173
rect 856 -1248 857 -1178
rect 863 -1179 864 -1173
rect 933 -1248 934 -1178
rect 996 -1179 997 -1173
rect 1087 -1248 1088 -1178
rect 19 -1181 20 -1173
rect 247 -1181 248 -1173
rect 310 -1248 311 -1180
rect 317 -1181 318 -1173
rect 331 -1181 332 -1173
rect 355 -1181 356 -1173
rect 359 -1181 360 -1173
rect 821 -1248 822 -1180
rect 912 -1181 913 -1173
rect 989 -1248 990 -1180
rect 1003 -1181 1004 -1173
rect 1094 -1248 1095 -1180
rect 23 -1183 24 -1173
rect 37 -1183 38 -1173
rect 58 -1183 59 -1173
rect 940 -1183 941 -1173
rect 947 -1183 948 -1173
rect 1003 -1248 1004 -1182
rect 1017 -1183 1018 -1173
rect 1108 -1248 1109 -1182
rect 23 -1248 24 -1184
rect 362 -1185 363 -1173
rect 380 -1248 381 -1184
rect 401 -1185 402 -1173
rect 443 -1185 444 -1173
rect 471 -1248 472 -1184
rect 478 -1248 479 -1184
rect 537 -1248 538 -1184
rect 562 -1185 563 -1173
rect 807 -1185 808 -1173
rect 877 -1185 878 -1173
rect 940 -1248 941 -1184
rect 1031 -1185 1032 -1173
rect 1143 -1248 1144 -1184
rect 37 -1248 38 -1186
rect 352 -1187 353 -1173
rect 366 -1187 367 -1173
rect 401 -1248 402 -1186
rect 429 -1187 430 -1173
rect 443 -1248 444 -1186
rect 464 -1187 465 -1173
rect 667 -1187 668 -1173
rect 681 -1187 682 -1173
rect 751 -1248 752 -1186
rect 758 -1187 759 -1173
rect 807 -1248 808 -1186
rect 884 -1187 885 -1173
rect 947 -1248 948 -1186
rect 1041 -1187 1042 -1173
rect 1066 -1187 1067 -1173
rect 44 -1189 45 -1173
rect 366 -1248 367 -1188
rect 394 -1189 395 -1173
rect 418 -1189 419 -1173
rect 429 -1248 430 -1188
rect 642 -1248 643 -1188
rect 656 -1248 657 -1188
rect 1136 -1248 1137 -1188
rect 44 -1248 45 -1190
rect 65 -1191 66 -1173
rect 96 -1248 97 -1190
rect 527 -1191 528 -1173
rect 534 -1191 535 -1173
rect 758 -1248 759 -1190
rect 786 -1191 787 -1173
rect 968 -1191 969 -1173
rect 1045 -1191 1046 -1173
rect 1101 -1248 1102 -1190
rect 58 -1248 59 -1192
rect 128 -1193 129 -1173
rect 135 -1193 136 -1173
rect 481 -1193 482 -1173
rect 506 -1248 507 -1192
rect 1024 -1193 1025 -1173
rect 1052 -1193 1053 -1173
rect 1122 -1248 1123 -1192
rect 61 -1195 62 -1173
rect 135 -1248 136 -1194
rect 142 -1195 143 -1173
rect 415 -1195 416 -1173
rect 513 -1195 514 -1173
rect 604 -1248 605 -1194
rect 681 -1248 682 -1194
rect 961 -1195 962 -1173
rect 1059 -1195 1060 -1173
rect 1150 -1248 1151 -1194
rect 65 -1248 66 -1196
rect 194 -1248 195 -1196
rect 198 -1197 199 -1173
rect 285 -1197 286 -1173
rect 289 -1197 290 -1173
rect 352 -1248 353 -1196
rect 394 -1248 395 -1196
rect 555 -1197 556 -1173
rect 562 -1248 563 -1196
rect 576 -1197 577 -1173
rect 597 -1197 598 -1173
rect 660 -1197 661 -1173
rect 688 -1197 689 -1173
rect 1024 -1248 1025 -1196
rect 100 -1199 101 -1173
rect 107 -1199 108 -1173
rect 121 -1199 122 -1173
rect 359 -1248 360 -1198
rect 415 -1248 416 -1198
rect 502 -1199 503 -1173
rect 523 -1199 524 -1173
rect 1066 -1248 1067 -1198
rect 100 -1248 101 -1200
rect 114 -1201 115 -1173
rect 121 -1248 122 -1200
rect 611 -1201 612 -1173
rect 688 -1248 689 -1200
rect 716 -1201 717 -1173
rect 733 -1201 734 -1173
rect 863 -1248 864 -1200
rect 891 -1201 892 -1173
rect 1017 -1248 1018 -1200
rect 79 -1203 80 -1173
rect 114 -1248 115 -1202
rect 128 -1248 129 -1202
rect 177 -1203 178 -1173
rect 184 -1203 185 -1173
rect 205 -1248 206 -1202
rect 222 -1203 223 -1173
rect 275 -1248 276 -1202
rect 296 -1203 297 -1173
rect 331 -1248 332 -1202
rect 345 -1203 346 -1173
rect 772 -1203 773 -1173
rect 786 -1248 787 -1202
rect 1010 -1203 1011 -1173
rect 79 -1248 80 -1204
rect 450 -1205 451 -1173
rect 513 -1248 514 -1204
rect 527 -1248 528 -1204
rect 632 -1205 633 -1173
rect 695 -1248 696 -1204
rect 765 -1205 766 -1173
rect 789 -1205 790 -1173
rect 1031 -1248 1032 -1204
rect 107 -1248 108 -1206
rect 324 -1207 325 -1173
rect 345 -1248 346 -1206
rect 373 -1207 374 -1173
rect 422 -1207 423 -1173
rect 772 -1248 773 -1206
rect 859 -1207 860 -1173
rect 1052 -1248 1053 -1206
rect 72 -1209 73 -1173
rect 324 -1248 325 -1208
rect 373 -1248 374 -1208
rect 814 -1209 815 -1173
rect 905 -1209 906 -1173
rect 961 -1248 962 -1208
rect 975 -1209 976 -1173
rect 1059 -1248 1060 -1208
rect 142 -1248 143 -1210
rect 369 -1248 370 -1210
rect 422 -1248 423 -1210
rect 492 -1211 493 -1173
rect 555 -1248 556 -1210
rect 1118 -1248 1119 -1210
rect 152 -1213 153 -1173
rect 464 -1248 465 -1212
rect 569 -1213 570 -1173
rect 611 -1248 612 -1212
rect 702 -1213 703 -1173
rect 891 -1248 892 -1212
rect 898 -1213 899 -1173
rect 975 -1248 976 -1212
rect 93 -1215 94 -1173
rect 702 -1248 703 -1214
rect 716 -1248 717 -1214
rect 877 -1248 878 -1214
rect 919 -1215 920 -1173
rect 996 -1248 997 -1214
rect 156 -1217 157 -1173
rect 219 -1248 220 -1216
rect 233 -1217 234 -1173
rect 884 -1248 885 -1216
rect 926 -1217 927 -1173
rect 1010 -1248 1011 -1216
rect 86 -1219 87 -1173
rect 233 -1248 234 -1218
rect 240 -1219 241 -1173
rect 296 -1248 297 -1218
rect 436 -1219 437 -1173
rect 450 -1248 451 -1218
rect 467 -1219 468 -1173
rect 569 -1248 570 -1218
rect 576 -1248 577 -1218
rect 590 -1219 591 -1173
rect 670 -1248 671 -1218
rect 919 -1248 920 -1218
rect 954 -1219 955 -1173
rect 1045 -1248 1046 -1218
rect 51 -1221 52 -1173
rect 436 -1248 437 -1220
rect 583 -1221 584 -1173
rect 590 -1248 591 -1220
rect 719 -1248 720 -1220
rect 954 -1248 955 -1220
rect 51 -1248 52 -1222
rect 268 -1223 269 -1173
rect 723 -1223 724 -1173
rect 765 -1248 766 -1222
rect 828 -1223 829 -1173
rect 898 -1248 899 -1222
rect 86 -1248 87 -1224
rect 170 -1225 171 -1173
rect 177 -1248 178 -1224
rect 387 -1225 388 -1173
rect 646 -1225 647 -1173
rect 723 -1248 724 -1224
rect 737 -1225 738 -1173
rect 912 -1248 913 -1224
rect 9 -1227 10 -1173
rect 170 -1248 171 -1226
rect 184 -1248 185 -1226
rect 261 -1227 262 -1173
rect 268 -1248 269 -1226
rect 282 -1227 283 -1173
rect 387 -1248 388 -1226
rect 625 -1227 626 -1173
rect 744 -1227 745 -1173
rect 814 -1248 815 -1226
rect 849 -1227 850 -1173
rect 926 -1248 927 -1226
rect 9 -1248 10 -1228
rect 30 -1229 31 -1173
rect 93 -1248 94 -1228
rect 583 -1248 584 -1228
rect 618 -1229 619 -1173
rect 646 -1248 647 -1228
rect 709 -1229 710 -1173
rect 744 -1248 745 -1228
rect 779 -1229 780 -1173
rect 849 -1248 850 -1228
rect 870 -1229 871 -1173
rect 905 -1248 906 -1228
rect 30 -1248 31 -1230
rect 289 -1248 290 -1230
rect 492 -1248 493 -1230
rect 737 -1248 738 -1230
rect 779 -1248 780 -1230
rect 793 -1231 794 -1173
rect 800 -1231 801 -1173
rect 870 -1248 871 -1230
rect 159 -1248 160 -1232
rect 600 -1233 601 -1173
rect 625 -1248 626 -1232
rect 667 -1248 668 -1232
rect 674 -1233 675 -1173
rect 709 -1248 710 -1232
rect 800 -1248 801 -1232
rect 1038 -1233 1039 -1173
rect 163 -1235 164 -1173
rect 982 -1248 983 -1234
rect 163 -1248 164 -1236
rect 212 -1237 213 -1173
rect 240 -1248 241 -1236
rect 348 -1237 349 -1173
rect 541 -1237 542 -1173
rect 618 -1248 619 -1236
rect 639 -1237 640 -1173
rect 793 -1248 794 -1236
rect 968 -1248 969 -1236
rect 1038 -1248 1039 -1236
rect 191 -1239 192 -1173
rect 226 -1248 227 -1238
rect 247 -1248 248 -1238
rect 303 -1248 304 -1238
rect 509 -1248 510 -1238
rect 541 -1248 542 -1238
rect 548 -1239 549 -1173
rect 674 -1248 675 -1238
rect 201 -1248 202 -1240
rect 317 -1248 318 -1240
rect 499 -1241 500 -1173
rect 548 -1248 549 -1240
rect 600 -1248 601 -1240
rect 842 -1241 843 -1173
rect 212 -1248 213 -1242
rect 271 -1248 272 -1242
rect 282 -1248 283 -1242
rect 338 -1243 339 -1173
rect 457 -1243 458 -1173
rect 499 -1248 500 -1242
rect 705 -1248 706 -1242
rect 842 -1248 843 -1242
rect 254 -1245 255 -1173
rect 261 -1248 262 -1244
rect 338 -1248 339 -1244
rect 684 -1248 685 -1244
rect 254 -1248 255 -1246
rect 376 -1248 377 -1246
rect 457 -1248 458 -1246
rect 660 -1248 661 -1246
rect 2 -1258 3 -1256
rect 72 -1258 73 -1256
rect 159 -1258 160 -1256
rect 387 -1258 388 -1256
rect 404 -1341 405 -1257
rect 527 -1258 528 -1256
rect 534 -1258 535 -1256
rect 618 -1258 619 -1256
rect 632 -1258 633 -1256
rect 814 -1258 815 -1256
rect 821 -1258 822 -1256
rect 1132 -1258 1133 -1256
rect 1164 -1258 1165 -1256
rect 1171 -1341 1172 -1257
rect 2 -1341 3 -1259
rect 51 -1260 52 -1256
rect 72 -1341 73 -1259
rect 268 -1260 269 -1256
rect 282 -1260 283 -1256
rect 303 -1260 304 -1256
rect 317 -1260 318 -1256
rect 439 -1341 440 -1259
rect 443 -1260 444 -1256
rect 446 -1286 447 -1259
rect 485 -1260 486 -1256
rect 702 -1341 703 -1259
rect 705 -1260 706 -1256
rect 1017 -1260 1018 -1256
rect 1024 -1260 1025 -1256
rect 1027 -1260 1028 -1256
rect 1122 -1260 1123 -1256
rect 1129 -1341 1130 -1259
rect 1157 -1260 1158 -1256
rect 1164 -1341 1165 -1259
rect 44 -1262 45 -1256
rect 215 -1341 216 -1261
rect 219 -1262 220 -1256
rect 219 -1341 220 -1261
rect 219 -1262 220 -1256
rect 219 -1341 220 -1261
rect 226 -1262 227 -1256
rect 226 -1341 227 -1261
rect 226 -1262 227 -1256
rect 226 -1341 227 -1261
rect 233 -1262 234 -1256
rect 292 -1262 293 -1256
rect 303 -1341 304 -1261
rect 555 -1262 556 -1256
rect 572 -1341 573 -1261
rect 870 -1262 871 -1256
rect 968 -1262 969 -1256
rect 1101 -1262 1102 -1256
rect 1122 -1341 1123 -1261
rect 1143 -1262 1144 -1256
rect 33 -1341 34 -1263
rect 44 -1341 45 -1263
rect 51 -1341 52 -1263
rect 170 -1264 171 -1256
rect 191 -1264 192 -1256
rect 1073 -1264 1074 -1256
rect 1143 -1341 1144 -1263
rect 1150 -1264 1151 -1256
rect 47 -1266 48 -1256
rect 1073 -1341 1074 -1265
rect 142 -1268 143 -1256
rect 814 -1341 815 -1267
rect 828 -1268 829 -1256
rect 877 -1268 878 -1256
rect 968 -1341 969 -1267
rect 982 -1268 983 -1256
rect 1024 -1341 1025 -1267
rect 1038 -1268 1039 -1256
rect 1052 -1268 1053 -1256
rect 1101 -1341 1102 -1267
rect 142 -1341 143 -1269
rect 212 -1270 213 -1256
rect 233 -1341 234 -1269
rect 296 -1270 297 -1256
rect 317 -1341 318 -1269
rect 411 -1341 412 -1269
rect 443 -1341 444 -1269
rect 464 -1270 465 -1256
rect 471 -1270 472 -1256
rect 485 -1341 486 -1269
rect 492 -1270 493 -1256
rect 604 -1270 605 -1256
rect 618 -1341 619 -1269
rect 674 -1270 675 -1256
rect 684 -1341 685 -1269
rect 961 -1270 962 -1256
rect 9 -1272 10 -1256
rect 212 -1341 213 -1271
rect 240 -1272 241 -1256
rect 369 -1272 370 -1256
rect 408 -1272 409 -1256
rect 506 -1272 507 -1256
rect 523 -1341 524 -1271
rect 898 -1272 899 -1256
rect 905 -1272 906 -1256
rect 961 -1341 962 -1271
rect 9 -1341 10 -1273
rect 254 -1274 255 -1256
rect 261 -1274 262 -1256
rect 271 -1274 272 -1256
rect 282 -1341 283 -1273
rect 660 -1274 661 -1256
rect 667 -1274 668 -1256
rect 989 -1274 990 -1256
rect 16 -1276 17 -1256
rect 604 -1341 605 -1275
rect 632 -1341 633 -1275
rect 751 -1276 752 -1256
rect 786 -1341 787 -1275
rect 807 -1276 808 -1256
rect 828 -1341 829 -1275
rect 1010 -1276 1011 -1256
rect 16 -1341 17 -1277
rect 180 -1341 181 -1277
rect 191 -1341 192 -1277
rect 205 -1278 206 -1256
rect 261 -1341 262 -1277
rect 537 -1341 538 -1277
rect 555 -1341 556 -1277
rect 562 -1278 563 -1256
rect 569 -1278 570 -1256
rect 982 -1341 983 -1277
rect 1010 -1341 1011 -1277
rect 1080 -1278 1081 -1256
rect 114 -1280 115 -1256
rect 240 -1341 241 -1279
rect 268 -1341 269 -1279
rect 338 -1280 339 -1256
rect 359 -1280 360 -1256
rect 387 -1341 388 -1279
rect 436 -1280 437 -1256
rect 807 -1341 808 -1279
rect 831 -1280 832 -1256
rect 1087 -1280 1088 -1256
rect 58 -1282 59 -1256
rect 359 -1341 360 -1281
rect 464 -1341 465 -1281
rect 471 -1341 472 -1281
rect 513 -1282 514 -1256
rect 534 -1341 535 -1281
rect 737 -1282 738 -1256
rect 751 -1341 752 -1281
rect 849 -1282 850 -1256
rect 877 -1341 878 -1281
rect 891 -1282 892 -1256
rect 1066 -1282 1067 -1256
rect 1087 -1341 1088 -1281
rect 58 -1341 59 -1283
rect 194 -1284 195 -1256
rect 205 -1341 206 -1283
rect 247 -1284 248 -1256
rect 289 -1284 290 -1256
rect 373 -1341 374 -1283
rect 457 -1284 458 -1256
rect 1052 -1341 1053 -1283
rect 86 -1286 87 -1256
rect 114 -1341 115 -1285
rect 135 -1286 136 -1256
rect 289 -1341 290 -1285
rect 296 -1341 297 -1285
rect 429 -1286 430 -1256
rect 457 -1341 458 -1285
rect 562 -1341 563 -1285
rect 576 -1286 577 -1256
rect 597 -1286 598 -1256
rect 600 -1286 601 -1256
rect 912 -1286 913 -1256
rect 1027 -1341 1028 -1285
rect 1038 -1341 1039 -1285
rect 1045 -1286 1046 -1256
rect 1066 -1341 1067 -1285
rect 86 -1341 87 -1287
rect 100 -1288 101 -1256
rect 107 -1288 108 -1256
rect 135 -1341 136 -1287
rect 156 -1288 157 -1256
rect 870 -1341 871 -1287
rect 891 -1341 892 -1287
rect 947 -1288 948 -1256
rect 1003 -1288 1004 -1256
rect 1045 -1341 1046 -1287
rect 26 -1341 27 -1289
rect 156 -1341 157 -1289
rect 163 -1290 164 -1256
rect 254 -1341 255 -1289
rect 275 -1290 276 -1256
rect 429 -1341 430 -1289
rect 478 -1290 479 -1256
rect 737 -1341 738 -1289
rect 796 -1341 797 -1289
rect 856 -1290 857 -1256
rect 912 -1341 913 -1289
rect 933 -1290 934 -1256
rect 947 -1341 948 -1289
rect 989 -1341 990 -1289
rect 1003 -1341 1004 -1289
rect 1031 -1290 1032 -1256
rect 37 -1292 38 -1256
rect 275 -1341 276 -1291
rect 324 -1292 325 -1256
rect 569 -1341 570 -1291
rect 590 -1292 591 -1256
rect 674 -1341 675 -1291
rect 688 -1292 689 -1256
rect 821 -1341 822 -1291
rect 835 -1292 836 -1256
rect 905 -1341 906 -1291
rect 933 -1341 934 -1291
rect 954 -1292 955 -1256
rect 1031 -1341 1032 -1291
rect 1136 -1292 1137 -1256
rect 37 -1341 38 -1293
rect 184 -1294 185 -1256
rect 247 -1341 248 -1293
rect 394 -1294 395 -1256
rect 408 -1341 409 -1293
rect 576 -1341 577 -1293
rect 607 -1341 608 -1293
rect 1080 -1341 1081 -1293
rect 1136 -1341 1137 -1293
rect 1157 -1341 1158 -1293
rect 100 -1341 101 -1295
rect 310 -1296 311 -1256
rect 324 -1341 325 -1295
rect 422 -1296 423 -1256
rect 495 -1296 496 -1256
rect 688 -1341 689 -1295
rect 716 -1341 717 -1295
rect 1115 -1296 1116 -1256
rect 107 -1341 108 -1297
rect 128 -1298 129 -1256
rect 170 -1341 171 -1297
rect 635 -1298 636 -1256
rect 639 -1298 640 -1256
rect 1017 -1341 1018 -1297
rect 1108 -1298 1109 -1256
rect 1115 -1341 1116 -1297
rect 30 -1300 31 -1256
rect 128 -1341 129 -1299
rect 184 -1341 185 -1299
rect 187 -1300 188 -1256
rect 310 -1341 311 -1299
rect 415 -1300 416 -1256
rect 499 -1300 500 -1256
rect 527 -1341 528 -1299
rect 541 -1300 542 -1256
rect 590 -1341 591 -1299
rect 621 -1341 622 -1299
rect 831 -1341 832 -1299
rect 849 -1341 850 -1299
rect 975 -1300 976 -1256
rect 1094 -1300 1095 -1256
rect 1108 -1341 1109 -1299
rect 65 -1302 66 -1256
rect 415 -1341 416 -1301
rect 513 -1341 514 -1301
rect 520 -1302 521 -1256
rect 642 -1302 643 -1256
rect 1059 -1302 1060 -1256
rect 121 -1304 122 -1256
rect 639 -1341 640 -1303
rect 646 -1304 647 -1256
rect 667 -1341 668 -1303
rect 670 -1304 671 -1256
rect 765 -1304 766 -1256
rect 779 -1304 780 -1256
rect 835 -1341 836 -1303
rect 842 -1304 843 -1256
rect 1094 -1341 1095 -1303
rect 79 -1306 80 -1256
rect 121 -1341 122 -1305
rect 338 -1341 339 -1305
rect 628 -1341 629 -1305
rect 646 -1341 647 -1305
rect 758 -1306 759 -1256
rect 772 -1306 773 -1256
rect 779 -1341 780 -1305
rect 800 -1306 801 -1256
rect 898 -1341 899 -1305
rect 940 -1306 941 -1256
rect 954 -1341 955 -1305
rect 975 -1341 976 -1305
rect 996 -1306 997 -1256
rect 79 -1341 80 -1307
rect 96 -1341 97 -1307
rect 345 -1308 346 -1256
rect 499 -1341 500 -1307
rect 506 -1341 507 -1307
rect 772 -1341 773 -1307
rect 842 -1341 843 -1307
rect 863 -1308 864 -1256
rect 198 -1310 199 -1256
rect 345 -1341 346 -1309
rect 348 -1341 349 -1309
rect 1059 -1341 1060 -1309
rect 177 -1312 178 -1256
rect 198 -1341 199 -1311
rect 352 -1312 353 -1256
rect 422 -1341 423 -1311
rect 436 -1341 437 -1311
rect 940 -1341 941 -1311
rect 352 -1341 353 -1313
rect 380 -1314 381 -1256
rect 394 -1341 395 -1313
rect 541 -1341 542 -1313
rect 597 -1341 598 -1313
rect 996 -1341 997 -1313
rect 366 -1316 367 -1256
rect 765 -1341 766 -1315
rect 856 -1341 857 -1315
rect 919 -1316 920 -1256
rect 23 -1341 24 -1317
rect 919 -1341 920 -1317
rect 331 -1320 332 -1256
rect 366 -1341 367 -1319
rect 380 -1341 381 -1319
rect 401 -1320 402 -1256
rect 520 -1341 521 -1319
rect 660 -1341 661 -1319
rect 709 -1320 710 -1256
rect 800 -1341 801 -1319
rect 149 -1322 150 -1256
rect 331 -1341 332 -1321
rect 401 -1341 402 -1321
rect 460 -1322 461 -1256
rect 625 -1322 626 -1256
rect 709 -1341 710 -1321
rect 723 -1322 724 -1256
rect 863 -1341 864 -1321
rect 149 -1341 150 -1323
rect 681 -1341 682 -1323
rect 695 -1324 696 -1256
rect 723 -1341 724 -1323
rect 733 -1341 734 -1323
rect 884 -1324 885 -1256
rect 103 -1341 104 -1325
rect 695 -1341 696 -1325
rect 744 -1326 745 -1256
rect 758 -1341 759 -1325
rect 884 -1341 885 -1325
rect 926 -1326 927 -1256
rect 460 -1341 461 -1327
rect 509 -1328 510 -1256
rect 544 -1341 545 -1327
rect 926 -1341 927 -1327
rect 653 -1330 654 -1256
rect 789 -1330 790 -1256
rect 492 -1341 493 -1331
rect 653 -1341 654 -1331
rect 656 -1332 657 -1256
rect 793 -1332 794 -1256
rect 548 -1334 549 -1256
rect 793 -1341 794 -1333
rect 548 -1341 549 -1335
rect 583 -1336 584 -1256
rect 730 -1336 731 -1256
rect 744 -1341 745 -1335
rect 583 -1341 584 -1337
rect 611 -1338 612 -1256
rect 478 -1341 479 -1339
rect 611 -1341 612 -1339
rect 2 -1351 3 -1349
rect 432 -1448 433 -1350
rect 436 -1448 437 -1350
rect 688 -1351 689 -1349
rect 733 -1351 734 -1349
rect 1045 -1351 1046 -1349
rect 1101 -1351 1102 -1349
rect 1150 -1351 1151 -1349
rect 1153 -1351 1154 -1349
rect 1164 -1351 1165 -1349
rect 2 -1448 3 -1352
rect 121 -1353 122 -1349
rect 135 -1353 136 -1349
rect 334 -1448 335 -1352
rect 359 -1353 360 -1349
rect 523 -1353 524 -1349
rect 527 -1353 528 -1349
rect 947 -1448 948 -1352
rect 950 -1353 951 -1349
rect 1129 -1353 1130 -1349
rect 1136 -1353 1137 -1349
rect 1171 -1353 1172 -1349
rect 9 -1355 10 -1349
rect 163 -1355 164 -1349
rect 215 -1355 216 -1349
rect 415 -1355 416 -1349
rect 506 -1355 507 -1349
rect 541 -1448 542 -1354
rect 544 -1355 545 -1349
rect 646 -1355 647 -1349
rect 688 -1448 689 -1354
rect 975 -1355 976 -1349
rect 996 -1448 997 -1354
rect 1066 -1355 1067 -1349
rect 16 -1357 17 -1349
rect 411 -1357 412 -1349
rect 506 -1448 507 -1356
rect 632 -1357 633 -1349
rect 681 -1357 682 -1349
rect 975 -1448 976 -1356
rect 1031 -1357 1032 -1349
rect 1066 -1448 1067 -1356
rect 23 -1448 24 -1358
rect 446 -1448 447 -1358
rect 513 -1359 514 -1349
rect 513 -1448 514 -1358
rect 513 -1359 514 -1349
rect 513 -1448 514 -1358
rect 520 -1448 521 -1358
rect 842 -1359 843 -1349
rect 919 -1359 920 -1349
rect 919 -1448 920 -1358
rect 919 -1359 920 -1349
rect 919 -1448 920 -1358
rect 940 -1359 941 -1349
rect 940 -1448 941 -1358
rect 940 -1359 941 -1349
rect 940 -1448 941 -1358
rect 1031 -1448 1032 -1358
rect 1094 -1359 1095 -1349
rect 26 -1361 27 -1349
rect 240 -1361 241 -1349
rect 275 -1361 276 -1349
rect 527 -1448 528 -1360
rect 537 -1361 538 -1349
rect 898 -1361 899 -1349
rect 1045 -1448 1046 -1360
rect 1143 -1361 1144 -1349
rect 33 -1363 34 -1349
rect 58 -1363 59 -1349
rect 65 -1363 66 -1349
rect 485 -1363 486 -1349
rect 562 -1363 563 -1349
rect 646 -1448 647 -1362
rect 681 -1448 682 -1362
rect 751 -1363 752 -1349
rect 772 -1363 773 -1349
rect 905 -1363 906 -1349
rect 44 -1365 45 -1349
rect 68 -1365 69 -1349
rect 93 -1365 94 -1349
rect 107 -1365 108 -1349
rect 121 -1448 122 -1364
rect 1080 -1365 1081 -1349
rect 44 -1448 45 -1366
rect 86 -1367 87 -1349
rect 100 -1367 101 -1349
rect 205 -1367 206 -1349
rect 212 -1367 213 -1349
rect 1094 -1448 1095 -1366
rect 16 -1448 17 -1368
rect 100 -1448 101 -1368
rect 103 -1369 104 -1349
rect 275 -1448 276 -1368
rect 289 -1448 290 -1368
rect 422 -1369 423 -1349
rect 485 -1448 486 -1368
rect 674 -1369 675 -1349
rect 751 -1448 752 -1368
rect 758 -1369 759 -1349
rect 772 -1448 773 -1368
rect 835 -1369 836 -1349
rect 842 -1448 843 -1368
rect 856 -1369 857 -1349
rect 898 -1448 899 -1368
rect 1024 -1369 1025 -1349
rect 51 -1371 52 -1349
rect 460 -1371 461 -1349
rect 492 -1448 493 -1370
rect 1080 -1448 1081 -1370
rect 51 -1448 52 -1372
rect 352 -1373 353 -1349
rect 359 -1448 360 -1372
rect 380 -1373 381 -1349
rect 387 -1373 388 -1349
rect 905 -1448 906 -1372
rect 58 -1448 59 -1374
rect 247 -1375 248 -1349
rect 268 -1375 269 -1349
rect 380 -1448 381 -1374
rect 387 -1448 388 -1374
rect 499 -1375 500 -1349
rect 600 -1448 601 -1374
rect 1052 -1375 1053 -1349
rect 65 -1448 66 -1376
rect 114 -1377 115 -1349
rect 128 -1377 129 -1349
rect 240 -1448 241 -1376
rect 247 -1448 248 -1376
rect 296 -1377 297 -1349
rect 303 -1377 304 -1349
rect 495 -1377 496 -1349
rect 569 -1377 570 -1349
rect 1052 -1448 1053 -1376
rect 37 -1379 38 -1349
rect 128 -1448 129 -1378
rect 135 -1448 136 -1378
rect 331 -1379 332 -1349
rect 366 -1379 367 -1349
rect 366 -1448 367 -1378
rect 366 -1379 367 -1349
rect 366 -1448 367 -1378
rect 373 -1379 374 -1349
rect 373 -1448 374 -1378
rect 373 -1379 374 -1349
rect 373 -1448 374 -1378
rect 394 -1379 395 -1349
rect 394 -1448 395 -1378
rect 394 -1379 395 -1349
rect 394 -1448 395 -1378
rect 408 -1379 409 -1349
rect 450 -1379 451 -1349
rect 611 -1379 612 -1349
rect 968 -1379 969 -1349
rect 37 -1448 38 -1380
rect 324 -1381 325 -1349
rect 331 -1448 332 -1380
rect 415 -1448 416 -1380
rect 422 -1448 423 -1380
rect 569 -1448 570 -1380
rect 611 -1448 612 -1380
rect 695 -1381 696 -1349
rect 758 -1448 759 -1380
rect 821 -1381 822 -1349
rect 828 -1381 829 -1349
rect 1108 -1381 1109 -1349
rect 72 -1383 73 -1349
rect 86 -1448 87 -1382
rect 103 -1448 104 -1382
rect 177 -1383 178 -1349
rect 187 -1448 188 -1382
rect 408 -1448 409 -1382
rect 443 -1383 444 -1349
rect 450 -1448 451 -1382
rect 509 -1448 510 -1382
rect 968 -1448 969 -1382
rect 1108 -1448 1109 -1382
rect 1157 -1383 1158 -1349
rect 72 -1448 73 -1384
rect 555 -1385 556 -1349
rect 614 -1385 615 -1349
rect 814 -1385 815 -1349
rect 821 -1448 822 -1384
rect 877 -1385 878 -1349
rect 79 -1387 80 -1349
rect 555 -1448 556 -1386
rect 625 -1387 626 -1349
rect 954 -1387 955 -1349
rect 79 -1448 80 -1388
rect 198 -1389 199 -1349
rect 226 -1389 227 -1349
rect 348 -1389 349 -1349
rect 618 -1389 619 -1349
rect 625 -1448 626 -1388
rect 632 -1448 633 -1388
rect 653 -1389 654 -1349
rect 660 -1389 661 -1349
rect 835 -1448 836 -1388
rect 849 -1389 850 -1349
rect 954 -1448 955 -1388
rect 110 -1448 111 -1390
rect 1024 -1448 1025 -1390
rect 149 -1393 150 -1349
rect 404 -1448 405 -1392
rect 653 -1448 654 -1392
rect 807 -1393 808 -1349
rect 814 -1448 815 -1392
rect 1062 -1448 1063 -1392
rect 149 -1448 150 -1394
rect 317 -1395 318 -1349
rect 324 -1448 325 -1394
rect 429 -1395 430 -1349
rect 660 -1448 661 -1394
rect 667 -1395 668 -1349
rect 674 -1448 675 -1394
rect 716 -1395 717 -1349
rect 775 -1395 776 -1349
rect 786 -1395 787 -1349
rect 828 -1448 829 -1394
rect 933 -1395 934 -1349
rect 156 -1397 157 -1349
rect 730 -1448 731 -1396
rect 786 -1448 787 -1396
rect 870 -1397 871 -1349
rect 877 -1448 878 -1396
rect 912 -1397 913 -1349
rect 933 -1448 934 -1396
rect 1087 -1397 1088 -1349
rect 156 -1448 157 -1398
rect 261 -1399 262 -1349
rect 282 -1399 283 -1349
rect 667 -1448 668 -1398
rect 695 -1448 696 -1398
rect 723 -1399 724 -1349
rect 856 -1448 857 -1398
rect 1059 -1399 1060 -1349
rect 163 -1448 164 -1400
rect 184 -1401 185 -1349
rect 191 -1401 192 -1349
rect 205 -1448 206 -1400
rect 219 -1401 220 -1349
rect 282 -1448 283 -1400
rect 292 -1401 293 -1349
rect 495 -1448 496 -1400
rect 716 -1448 717 -1400
rect 765 -1401 766 -1349
rect 870 -1448 871 -1400
rect 884 -1401 885 -1349
rect 912 -1448 913 -1400
rect 1010 -1401 1011 -1349
rect 177 -1448 178 -1402
rect 352 -1448 353 -1402
rect 534 -1403 535 -1349
rect 884 -1448 885 -1402
rect 926 -1403 927 -1349
rect 1087 -1448 1088 -1402
rect 194 -1448 195 -1404
rect 268 -1448 269 -1404
rect 296 -1448 297 -1404
rect 502 -1448 503 -1404
rect 723 -1448 724 -1404
rect 737 -1405 738 -1349
rect 765 -1448 766 -1404
rect 779 -1405 780 -1349
rect 891 -1405 892 -1349
rect 926 -1448 927 -1404
rect 961 -1405 962 -1349
rect 1010 -1448 1011 -1404
rect 198 -1448 199 -1406
rect 604 -1407 605 -1349
rect 737 -1448 738 -1406
rect 744 -1407 745 -1349
rect 779 -1448 780 -1406
rect 800 -1407 801 -1349
rect 961 -1448 962 -1406
rect 982 -1407 983 -1349
rect 30 -1409 31 -1349
rect 800 -1448 801 -1408
rect 982 -1448 983 -1408
rect 989 -1409 990 -1349
rect 30 -1448 31 -1410
rect 142 -1411 143 -1349
rect 219 -1448 220 -1410
rect 233 -1411 234 -1349
rect 254 -1411 255 -1349
rect 261 -1448 262 -1410
rect 310 -1411 311 -1349
rect 439 -1411 440 -1349
rect 471 -1411 472 -1349
rect 534 -1448 535 -1410
rect 604 -1448 605 -1410
rect 709 -1411 710 -1349
rect 793 -1411 794 -1349
rect 891 -1448 892 -1410
rect 989 -1448 990 -1410
rect 1003 -1411 1004 -1349
rect 93 -1448 94 -1412
rect 744 -1448 745 -1412
rect 1003 -1448 1004 -1412
rect 1073 -1413 1074 -1349
rect 142 -1448 143 -1414
rect 170 -1415 171 -1349
rect 226 -1448 227 -1414
rect 457 -1415 458 -1349
rect 464 -1415 465 -1349
rect 471 -1448 472 -1414
rect 639 -1415 640 -1349
rect 709 -1448 710 -1414
rect 1073 -1448 1074 -1414
rect 1122 -1415 1123 -1349
rect 96 -1417 97 -1349
rect 170 -1448 171 -1416
rect 233 -1448 234 -1416
rect 401 -1417 402 -1349
rect 457 -1448 458 -1416
rect 691 -1448 692 -1416
rect 702 -1417 703 -1349
rect 793 -1448 794 -1416
rect 254 -1448 255 -1418
rect 849 -1448 850 -1418
rect 303 -1448 304 -1420
rect 439 -1448 440 -1420
rect 464 -1448 465 -1420
rect 576 -1421 577 -1349
rect 702 -1448 703 -1420
rect 807 -1448 808 -1420
rect 310 -1448 311 -1422
rect 597 -1423 598 -1349
rect 317 -1448 318 -1424
rect 579 -1448 580 -1424
rect 338 -1427 339 -1349
rect 618 -1448 619 -1426
rect 338 -1448 339 -1428
rect 488 -1448 489 -1428
rect 499 -1448 500 -1428
rect 639 -1448 640 -1428
rect 401 -1448 402 -1430
rect 562 -1448 563 -1430
rect 576 -1448 577 -1430
rect 863 -1431 864 -1349
rect 345 -1433 346 -1349
rect 863 -1448 864 -1432
rect 345 -1448 346 -1434
rect 478 -1435 479 -1349
rect 478 -1448 479 -1436
rect 590 -1437 591 -1349
rect 583 -1439 584 -1349
rect 590 -1448 591 -1438
rect 548 -1441 549 -1349
rect 583 -1448 584 -1440
rect 548 -1448 549 -1442
rect 1017 -1443 1018 -1349
rect 1017 -1448 1018 -1444
rect 1038 -1445 1039 -1349
rect 1038 -1448 1039 -1446
rect 1115 -1447 1116 -1349
rect 9 -1458 10 -1456
rect 467 -1539 468 -1457
rect 481 -1539 482 -1457
rect 604 -1458 605 -1456
rect 611 -1458 612 -1456
rect 996 -1458 997 -1456
rect 1010 -1458 1011 -1456
rect 1059 -1539 1060 -1457
rect 16 -1460 17 -1456
rect 495 -1460 496 -1456
rect 499 -1460 500 -1456
rect 947 -1460 948 -1456
rect 996 -1539 997 -1459
rect 1073 -1460 1074 -1456
rect 16 -1539 17 -1461
rect 331 -1462 332 -1456
rect 352 -1462 353 -1456
rect 523 -1539 524 -1461
rect 551 -1462 552 -1456
rect 674 -1462 675 -1456
rect 681 -1462 682 -1456
rect 702 -1539 703 -1461
rect 744 -1462 745 -1456
rect 1045 -1462 1046 -1456
rect 1062 -1462 1063 -1456
rect 1073 -1539 1074 -1461
rect 30 -1464 31 -1456
rect 187 -1464 188 -1456
rect 198 -1464 199 -1456
rect 548 -1464 549 -1456
rect 569 -1464 570 -1456
rect 660 -1464 661 -1456
rect 681 -1539 682 -1463
rect 765 -1464 766 -1456
rect 856 -1464 857 -1456
rect 912 -1464 913 -1456
rect 947 -1539 948 -1463
rect 1031 -1464 1032 -1456
rect 23 -1466 24 -1456
rect 198 -1539 199 -1465
rect 257 -1466 258 -1456
rect 261 -1466 262 -1456
rect 282 -1466 283 -1456
rect 282 -1539 283 -1465
rect 282 -1466 283 -1456
rect 282 -1539 283 -1465
rect 289 -1466 290 -1456
rect 411 -1466 412 -1456
rect 415 -1466 416 -1456
rect 429 -1539 430 -1465
rect 436 -1539 437 -1465
rect 506 -1466 507 -1456
rect 516 -1539 517 -1465
rect 758 -1466 759 -1456
rect 765 -1539 766 -1465
rect 835 -1466 836 -1456
rect 856 -1539 857 -1465
rect 961 -1466 962 -1456
rect 1017 -1466 1018 -1456
rect 1020 -1470 1021 -1465
rect 23 -1539 24 -1467
rect 254 -1468 255 -1456
rect 292 -1539 293 -1467
rect 359 -1468 360 -1456
rect 387 -1468 388 -1456
rect 499 -1539 500 -1467
rect 502 -1468 503 -1456
rect 695 -1468 696 -1456
rect 747 -1468 748 -1456
rect 877 -1468 878 -1456
rect 884 -1468 885 -1456
rect 1010 -1539 1011 -1467
rect 1017 -1539 1018 -1467
rect 1038 -1468 1039 -1456
rect 33 -1539 34 -1469
rect 716 -1470 717 -1456
rect 758 -1539 759 -1469
rect 786 -1470 787 -1456
rect 835 -1539 836 -1469
rect 954 -1470 955 -1456
rect 1038 -1539 1039 -1469
rect 44 -1472 45 -1456
rect 110 -1472 111 -1456
rect 114 -1472 115 -1456
rect 268 -1472 269 -1456
rect 303 -1472 304 -1456
rect 303 -1539 304 -1471
rect 303 -1472 304 -1456
rect 303 -1539 304 -1471
rect 310 -1472 311 -1456
rect 509 -1472 510 -1456
rect 541 -1472 542 -1456
rect 548 -1539 549 -1471
rect 569 -1539 570 -1471
rect 663 -1539 664 -1471
rect 695 -1539 696 -1471
rect 919 -1472 920 -1456
rect 933 -1472 934 -1456
rect 961 -1539 962 -1471
rect 30 -1539 31 -1473
rect 44 -1539 45 -1473
rect 51 -1474 52 -1456
rect 215 -1474 216 -1456
rect 254 -1539 255 -1473
rect 296 -1474 297 -1456
rect 310 -1539 311 -1473
rect 327 -1539 328 -1473
rect 331 -1539 332 -1473
rect 373 -1474 374 -1456
rect 387 -1539 388 -1473
rect 478 -1539 479 -1473
rect 485 -1474 486 -1456
rect 667 -1474 668 -1456
rect 730 -1474 731 -1456
rect 919 -1539 920 -1473
rect 954 -1539 955 -1473
rect 1094 -1474 1095 -1456
rect 2 -1476 3 -1456
rect 215 -1539 216 -1475
rect 296 -1539 297 -1475
rect 513 -1476 514 -1456
rect 541 -1539 542 -1475
rect 639 -1476 640 -1456
rect 730 -1539 731 -1475
rect 751 -1476 752 -1456
rect 786 -1539 787 -1475
rect 891 -1476 892 -1456
rect 912 -1539 913 -1475
rect 989 -1476 990 -1456
rect 1094 -1539 1095 -1475
rect 1108 -1476 1109 -1456
rect 2 -1539 3 -1477
rect 96 -1539 97 -1477
rect 103 -1478 104 -1456
rect 674 -1539 675 -1477
rect 688 -1539 689 -1477
rect 989 -1539 990 -1477
rect 51 -1539 52 -1479
rect 324 -1480 325 -1456
rect 345 -1480 346 -1456
rect 415 -1539 416 -1479
rect 422 -1480 423 -1456
rect 506 -1539 507 -1479
rect 576 -1480 577 -1456
rect 821 -1480 822 -1456
rect 859 -1480 860 -1456
rect 933 -1539 934 -1479
rect 37 -1482 38 -1456
rect 324 -1539 325 -1481
rect 373 -1539 374 -1481
rect 380 -1482 381 -1456
rect 394 -1482 395 -1456
rect 404 -1482 405 -1456
rect 408 -1482 409 -1456
rect 744 -1539 745 -1481
rect 821 -1539 822 -1481
rect 905 -1482 906 -1456
rect 9 -1539 10 -1483
rect 37 -1539 38 -1483
rect 65 -1484 66 -1456
rect 191 -1484 192 -1456
rect 233 -1484 234 -1456
rect 751 -1539 752 -1483
rect 863 -1484 864 -1456
rect 1045 -1539 1046 -1483
rect 58 -1486 59 -1456
rect 191 -1539 192 -1485
rect 226 -1486 227 -1456
rect 233 -1539 234 -1485
rect 366 -1486 367 -1456
rect 380 -1539 381 -1485
rect 401 -1539 402 -1485
rect 614 -1486 615 -1456
rect 639 -1539 640 -1485
rect 709 -1486 710 -1456
rect 807 -1486 808 -1456
rect 863 -1539 864 -1485
rect 870 -1486 871 -1456
rect 891 -1539 892 -1485
rect 58 -1539 59 -1487
rect 142 -1488 143 -1456
rect 163 -1488 164 -1456
rect 180 -1488 181 -1456
rect 226 -1539 227 -1487
rect 289 -1539 290 -1487
rect 422 -1539 423 -1487
rect 670 -1539 671 -1487
rect 807 -1539 808 -1487
rect 940 -1488 941 -1456
rect 65 -1539 66 -1489
rect 450 -1490 451 -1456
rect 464 -1490 465 -1456
rect 611 -1539 612 -1489
rect 870 -1539 871 -1489
rect 968 -1490 969 -1456
rect 72 -1492 73 -1456
rect 268 -1539 269 -1491
rect 432 -1492 433 -1456
rect 716 -1539 717 -1491
rect 877 -1539 878 -1491
rect 982 -1492 983 -1456
rect 72 -1539 73 -1493
rect 219 -1494 220 -1456
rect 439 -1494 440 -1456
rect 814 -1494 815 -1456
rect 884 -1539 885 -1493
rect 898 -1494 899 -1456
rect 940 -1539 941 -1493
rect 1024 -1494 1025 -1456
rect 79 -1496 80 -1456
rect 334 -1496 335 -1456
rect 443 -1496 444 -1456
rect 471 -1496 472 -1456
rect 485 -1539 486 -1495
rect 793 -1496 794 -1456
rect 814 -1539 815 -1495
rect 828 -1496 829 -1456
rect 968 -1539 969 -1495
rect 1003 -1496 1004 -1456
rect 1024 -1539 1025 -1495
rect 1080 -1496 1081 -1456
rect 79 -1539 80 -1497
rect 247 -1498 248 -1456
rect 443 -1539 444 -1497
rect 562 -1498 563 -1456
rect 590 -1498 591 -1456
rect 604 -1539 605 -1497
rect 793 -1539 794 -1497
rect 849 -1498 850 -1456
rect 982 -1539 983 -1497
rect 1052 -1498 1053 -1456
rect 86 -1500 87 -1456
rect 145 -1539 146 -1499
rect 163 -1539 164 -1499
rect 520 -1500 521 -1456
rect 534 -1500 535 -1456
rect 590 -1539 591 -1499
rect 597 -1539 598 -1499
rect 646 -1500 647 -1456
rect 779 -1500 780 -1456
rect 849 -1539 850 -1499
rect 1003 -1539 1004 -1499
rect 1066 -1500 1067 -1456
rect 86 -1539 87 -1501
rect 149 -1502 150 -1456
rect 166 -1539 167 -1501
rect 632 -1502 633 -1456
rect 646 -1539 647 -1501
rect 737 -1502 738 -1456
rect 772 -1502 773 -1456
rect 779 -1539 780 -1501
rect 828 -1539 829 -1501
rect 842 -1502 843 -1456
rect 107 -1504 108 -1456
rect 170 -1504 171 -1456
rect 177 -1504 178 -1456
rect 492 -1539 493 -1503
rect 534 -1539 535 -1503
rect 709 -1539 710 -1503
rect 842 -1539 843 -1503
rect 926 -1504 927 -1456
rect 93 -1506 94 -1456
rect 107 -1539 108 -1505
rect 114 -1539 115 -1505
rect 691 -1506 692 -1456
rect 705 -1506 706 -1456
rect 926 -1539 927 -1505
rect 93 -1539 94 -1507
rect 600 -1508 601 -1456
rect 677 -1539 678 -1507
rect 737 -1539 738 -1507
rect 121 -1539 122 -1509
rect 579 -1510 580 -1456
rect 691 -1539 692 -1509
rect 800 -1510 801 -1456
rect 124 -1512 125 -1456
rect 240 -1512 241 -1456
rect 247 -1539 248 -1511
rect 618 -1512 619 -1456
rect 800 -1539 801 -1511
rect 975 -1512 976 -1456
rect 128 -1514 129 -1456
rect 261 -1539 262 -1513
rect 366 -1539 367 -1513
rect 562 -1539 563 -1513
rect 618 -1539 619 -1513
rect 723 -1514 724 -1456
rect 128 -1539 129 -1515
rect 184 -1516 185 -1456
rect 212 -1516 213 -1456
rect 975 -1539 976 -1515
rect 100 -1539 101 -1517
rect 212 -1539 213 -1517
rect 219 -1539 220 -1517
rect 408 -1539 409 -1517
rect 450 -1539 451 -1517
rect 537 -1539 538 -1517
rect 555 -1518 556 -1456
rect 905 -1539 906 -1517
rect 135 -1520 136 -1456
rect 352 -1539 353 -1519
rect 359 -1539 360 -1519
rect 723 -1539 724 -1519
rect 135 -1539 136 -1521
rect 338 -1522 339 -1456
rect 457 -1522 458 -1456
rect 632 -1539 633 -1521
rect 149 -1539 150 -1523
rect 625 -1524 626 -1456
rect 156 -1526 157 -1456
rect 170 -1539 171 -1525
rect 177 -1539 178 -1525
rect 394 -1539 395 -1525
rect 457 -1539 458 -1525
rect 576 -1539 577 -1525
rect 625 -1539 626 -1525
rect 653 -1526 654 -1456
rect 156 -1539 157 -1527
rect 898 -1539 899 -1527
rect 184 -1539 185 -1529
rect 205 -1530 206 -1456
rect 240 -1539 241 -1529
rect 317 -1530 318 -1456
rect 338 -1539 339 -1529
rect 1031 -1539 1032 -1529
rect 194 -1532 195 -1456
rect 653 -1539 654 -1531
rect 205 -1539 206 -1533
rect 345 -1539 346 -1533
rect 527 -1534 528 -1456
rect 555 -1539 556 -1533
rect 275 -1536 276 -1456
rect 317 -1539 318 -1535
rect 527 -1539 528 -1535
rect 583 -1536 584 -1456
rect 513 -1539 514 -1537
rect 583 -1539 584 -1537
rect 2 -1549 3 -1547
rect 247 -1628 248 -1548
rect 254 -1549 255 -1547
rect 289 -1628 290 -1548
rect 352 -1549 353 -1547
rect 359 -1549 360 -1547
rect 376 -1628 377 -1548
rect 436 -1549 437 -1547
rect 457 -1549 458 -1547
rect 919 -1549 920 -1547
rect 940 -1549 941 -1547
rect 1010 -1628 1011 -1548
rect 1034 -1549 1035 -1547
rect 1038 -1549 1039 -1547
rect 1045 -1549 1046 -1547
rect 1101 -1628 1102 -1548
rect 5 -1628 6 -1550
rect 100 -1551 101 -1547
rect 145 -1551 146 -1547
rect 1052 -1628 1053 -1550
rect 1059 -1551 1060 -1547
rect 1108 -1628 1109 -1550
rect 9 -1553 10 -1547
rect 250 -1553 251 -1547
rect 261 -1553 262 -1547
rect 436 -1628 437 -1552
rect 464 -1553 465 -1547
rect 695 -1553 696 -1547
rect 772 -1553 773 -1547
rect 891 -1553 892 -1547
rect 975 -1553 976 -1547
rect 1045 -1628 1046 -1552
rect 1094 -1553 1095 -1547
rect 1115 -1628 1116 -1552
rect 9 -1628 10 -1554
rect 485 -1555 486 -1547
rect 513 -1628 514 -1554
rect 670 -1555 671 -1547
rect 674 -1555 675 -1547
rect 1017 -1555 1018 -1547
rect 1073 -1555 1074 -1547
rect 1094 -1628 1095 -1554
rect 30 -1628 31 -1556
rect 149 -1557 150 -1547
rect 156 -1557 157 -1547
rect 184 -1557 185 -1547
rect 198 -1557 199 -1547
rect 261 -1628 262 -1556
rect 268 -1557 269 -1547
rect 534 -1557 535 -1547
rect 562 -1557 563 -1547
rect 905 -1557 906 -1547
rect 926 -1557 927 -1547
rect 1017 -1628 1018 -1556
rect 33 -1559 34 -1547
rect 40 -1559 41 -1547
rect 51 -1559 52 -1547
rect 460 -1559 461 -1547
rect 471 -1559 472 -1547
rect 751 -1559 752 -1547
rect 821 -1559 822 -1547
rect 891 -1628 892 -1558
rect 989 -1559 990 -1547
rect 1073 -1628 1074 -1558
rect 37 -1561 38 -1547
rect 653 -1561 654 -1547
rect 660 -1628 661 -1560
rect 758 -1561 759 -1547
rect 821 -1628 822 -1560
rect 1069 -1628 1070 -1560
rect 37 -1628 38 -1562
rect 44 -1563 45 -1547
rect 51 -1628 52 -1562
rect 425 -1628 426 -1562
rect 478 -1563 479 -1547
rect 499 -1563 500 -1547
rect 520 -1563 521 -1547
rect 618 -1563 619 -1547
rect 625 -1563 626 -1547
rect 772 -1628 773 -1562
rect 835 -1563 836 -1547
rect 926 -1628 927 -1562
rect 961 -1563 962 -1547
rect 989 -1628 990 -1562
rect 996 -1563 997 -1547
rect 1080 -1628 1081 -1562
rect 65 -1565 66 -1547
rect 499 -1628 500 -1564
rect 534 -1628 535 -1564
rect 898 -1565 899 -1547
rect 16 -1567 17 -1547
rect 65 -1628 66 -1566
rect 72 -1567 73 -1547
rect 520 -1628 521 -1566
rect 565 -1567 566 -1547
rect 1024 -1567 1025 -1547
rect 16 -1628 17 -1568
rect 222 -1628 223 -1568
rect 268 -1628 269 -1568
rect 338 -1569 339 -1547
rect 359 -1628 360 -1568
rect 677 -1569 678 -1547
rect 716 -1569 717 -1547
rect 751 -1628 752 -1568
rect 814 -1569 815 -1547
rect 898 -1628 899 -1568
rect 982 -1569 983 -1547
rect 1024 -1628 1025 -1568
rect 72 -1628 73 -1570
rect 86 -1571 87 -1547
rect 93 -1628 94 -1570
rect 569 -1571 570 -1547
rect 576 -1571 577 -1547
rect 688 -1628 689 -1570
rect 716 -1628 717 -1570
rect 744 -1571 745 -1547
rect 765 -1571 766 -1547
rect 814 -1628 815 -1570
rect 842 -1571 843 -1547
rect 842 -1628 843 -1570
rect 842 -1571 843 -1547
rect 842 -1628 843 -1570
rect 859 -1628 860 -1570
rect 1003 -1571 1004 -1547
rect 79 -1573 80 -1547
rect 149 -1628 150 -1572
rect 163 -1573 164 -1547
rect 471 -1628 472 -1572
rect 478 -1628 479 -1572
rect 674 -1628 675 -1572
rect 684 -1628 685 -1572
rect 744 -1628 745 -1572
rect 765 -1628 766 -1572
rect 863 -1573 864 -1547
rect 870 -1573 871 -1547
rect 919 -1628 920 -1572
rect 933 -1573 934 -1547
rect 1003 -1628 1004 -1572
rect 79 -1628 80 -1574
rect 275 -1628 276 -1574
rect 282 -1575 283 -1547
rect 292 -1575 293 -1547
rect 345 -1575 346 -1547
rect 863 -1628 864 -1574
rect 884 -1575 885 -1547
rect 975 -1628 976 -1574
rect 86 -1628 87 -1576
rect 114 -1577 115 -1547
rect 121 -1577 122 -1547
rect 156 -1628 157 -1576
rect 163 -1628 164 -1576
rect 450 -1577 451 -1547
rect 464 -1628 465 -1576
rect 618 -1628 619 -1576
rect 625 -1628 626 -1576
rect 1038 -1628 1039 -1576
rect 96 -1628 97 -1578
rect 516 -1579 517 -1547
rect 527 -1579 528 -1547
rect 576 -1628 577 -1578
rect 590 -1579 591 -1547
rect 961 -1628 962 -1578
rect 968 -1579 969 -1547
rect 982 -1628 983 -1578
rect 100 -1628 101 -1580
rect 107 -1581 108 -1547
rect 121 -1628 122 -1580
rect 135 -1581 136 -1547
rect 166 -1581 167 -1547
rect 485 -1628 486 -1580
rect 506 -1581 507 -1547
rect 527 -1628 528 -1580
rect 583 -1581 584 -1547
rect 590 -1628 591 -1580
rect 593 -1581 594 -1547
rect 702 -1581 703 -1547
rect 723 -1581 724 -1547
rect 835 -1628 836 -1580
rect 912 -1581 913 -1547
rect 968 -1628 969 -1580
rect 107 -1628 108 -1582
rect 310 -1583 311 -1547
rect 331 -1583 332 -1547
rect 450 -1628 451 -1582
rect 597 -1583 598 -1547
rect 1087 -1628 1088 -1582
rect 128 -1585 129 -1547
rect 145 -1628 146 -1584
rect 170 -1585 171 -1547
rect 170 -1628 171 -1584
rect 170 -1585 171 -1547
rect 170 -1628 171 -1584
rect 177 -1628 178 -1584
rect 401 -1585 402 -1547
rect 597 -1628 598 -1584
rect 604 -1585 605 -1547
rect 611 -1585 612 -1547
rect 677 -1628 678 -1584
rect 723 -1628 724 -1584
rect 730 -1585 731 -1547
rect 793 -1585 794 -1547
rect 870 -1628 871 -1584
rect 114 -1628 115 -1586
rect 611 -1628 612 -1586
rect 614 -1628 615 -1586
rect 940 -1628 941 -1586
rect 128 -1628 129 -1588
rect 352 -1628 353 -1588
rect 366 -1589 367 -1547
rect 401 -1628 402 -1588
rect 429 -1589 430 -1547
rect 604 -1628 605 -1588
rect 632 -1589 633 -1547
rect 905 -1628 906 -1588
rect 180 -1591 181 -1547
rect 422 -1591 423 -1547
rect 457 -1628 458 -1590
rect 793 -1628 794 -1590
rect 800 -1591 801 -1547
rect 933 -1628 934 -1590
rect 201 -1628 202 -1592
rect 681 -1593 682 -1547
rect 730 -1628 731 -1592
rect 849 -1593 850 -1547
rect 205 -1628 206 -1594
rect 208 -1595 209 -1547
rect 212 -1595 213 -1547
rect 229 -1628 230 -1594
rect 233 -1595 234 -1547
rect 506 -1628 507 -1594
rect 635 -1628 636 -1594
rect 702 -1628 703 -1594
rect 800 -1628 801 -1594
rect 1062 -1628 1063 -1594
rect 191 -1597 192 -1547
rect 212 -1628 213 -1596
rect 219 -1597 220 -1547
rect 254 -1628 255 -1596
rect 278 -1597 279 -1547
rect 849 -1628 850 -1596
rect 58 -1599 59 -1547
rect 191 -1628 192 -1598
rect 226 -1599 227 -1547
rect 345 -1628 346 -1598
rect 366 -1628 367 -1598
rect 467 -1599 468 -1547
rect 639 -1599 640 -1547
rect 653 -1628 654 -1598
rect 663 -1599 664 -1547
rect 807 -1599 808 -1547
rect 828 -1599 829 -1547
rect 884 -1628 885 -1598
rect 44 -1628 45 -1600
rect 226 -1628 227 -1600
rect 233 -1628 234 -1600
rect 387 -1601 388 -1547
rect 394 -1601 395 -1547
rect 562 -1628 563 -1600
rect 639 -1628 640 -1600
rect 1031 -1601 1032 -1547
rect 58 -1628 59 -1602
rect 695 -1628 696 -1602
rect 737 -1603 738 -1547
rect 807 -1628 808 -1602
rect 947 -1603 948 -1547
rect 1031 -1628 1032 -1602
rect 240 -1605 241 -1547
rect 331 -1628 332 -1604
rect 355 -1628 356 -1604
rect 394 -1628 395 -1604
rect 408 -1605 409 -1547
rect 429 -1628 430 -1604
rect 646 -1605 647 -1547
rect 912 -1628 913 -1604
rect 947 -1628 948 -1604
rect 954 -1605 955 -1547
rect 240 -1628 241 -1606
rect 317 -1607 318 -1547
rect 324 -1607 325 -1547
rect 632 -1628 633 -1606
rect 667 -1607 668 -1547
rect 779 -1607 780 -1547
rect 877 -1607 878 -1547
rect 954 -1628 955 -1606
rect 282 -1628 283 -1608
rect 586 -1628 587 -1608
rect 709 -1609 710 -1547
rect 877 -1628 878 -1608
rect 303 -1611 304 -1547
rect 317 -1628 318 -1610
rect 373 -1611 374 -1547
rect 387 -1628 388 -1610
rect 408 -1628 409 -1610
rect 415 -1611 416 -1547
rect 492 -1611 493 -1547
rect 646 -1628 647 -1610
rect 737 -1628 738 -1610
rect 786 -1611 787 -1547
rect 23 -1613 24 -1547
rect 492 -1628 493 -1612
rect 523 -1613 524 -1547
rect 709 -1628 710 -1612
rect 758 -1628 759 -1612
rect 779 -1628 780 -1612
rect 786 -1628 787 -1612
rect 856 -1613 857 -1547
rect 23 -1628 24 -1614
rect 296 -1615 297 -1547
rect 310 -1628 311 -1614
rect 327 -1628 328 -1614
rect 338 -1628 339 -1614
rect 373 -1628 374 -1614
rect 415 -1628 416 -1614
rect 569 -1628 570 -1614
rect 775 -1615 776 -1547
rect 828 -1628 829 -1614
rect 856 -1628 857 -1614
rect 996 -1628 997 -1614
rect 296 -1628 297 -1616
rect 380 -1617 381 -1547
rect 537 -1617 538 -1547
rect 667 -1628 668 -1616
rect 380 -1628 381 -1618
rect 443 -1619 444 -1547
rect 443 -1628 444 -1620
rect 541 -1621 542 -1547
rect 541 -1628 542 -1622
rect 555 -1623 556 -1547
rect 548 -1625 549 -1547
rect 555 -1628 556 -1624
rect 82 -1628 83 -1626
rect 548 -1628 549 -1626
rect 9 -1638 10 -1636
rect 341 -1713 342 -1637
rect 345 -1638 346 -1636
rect 345 -1713 346 -1637
rect 345 -1638 346 -1636
rect 345 -1713 346 -1637
rect 355 -1638 356 -1636
rect 604 -1638 605 -1636
rect 607 -1713 608 -1637
rect 926 -1638 927 -1636
rect 1059 -1638 1060 -1636
rect 1108 -1638 1109 -1636
rect 23 -1640 24 -1636
rect 26 -1656 27 -1639
rect 37 -1640 38 -1636
rect 40 -1656 41 -1639
rect 58 -1640 59 -1636
rect 695 -1640 696 -1636
rect 779 -1640 780 -1636
rect 884 -1640 885 -1636
rect 1066 -1713 1067 -1639
rect 1094 -1640 1095 -1636
rect 23 -1713 24 -1641
rect 142 -1642 143 -1636
rect 149 -1642 150 -1636
rect 306 -1642 307 -1636
rect 313 -1713 314 -1641
rect 485 -1642 486 -1636
rect 523 -1713 524 -1641
rect 660 -1642 661 -1636
rect 674 -1642 675 -1636
rect 989 -1642 990 -1636
rect 1069 -1642 1070 -1636
rect 1115 -1642 1116 -1636
rect 37 -1713 38 -1643
rect 198 -1644 199 -1636
rect 222 -1644 223 -1636
rect 520 -1644 521 -1636
rect 534 -1713 535 -1643
rect 576 -1644 577 -1636
rect 583 -1644 584 -1636
rect 947 -1644 948 -1636
rect 1094 -1713 1095 -1643
rect 1101 -1644 1102 -1636
rect 58 -1713 59 -1645
rect 100 -1646 101 -1636
rect 114 -1646 115 -1636
rect 198 -1713 199 -1645
rect 247 -1713 248 -1645
rect 324 -1646 325 -1636
rect 376 -1646 377 -1636
rect 828 -1646 829 -1636
rect 835 -1646 836 -1636
rect 884 -1713 885 -1645
rect 947 -1713 948 -1645
rect 1073 -1646 1074 -1636
rect 51 -1648 52 -1636
rect 114 -1713 115 -1647
rect 135 -1648 136 -1636
rect 443 -1713 444 -1647
rect 450 -1648 451 -1636
rect 485 -1713 486 -1647
rect 572 -1648 573 -1636
rect 912 -1648 913 -1636
rect 16 -1650 17 -1636
rect 135 -1713 136 -1649
rect 138 -1650 139 -1636
rect 331 -1650 332 -1636
rect 383 -1713 384 -1649
rect 761 -1713 762 -1649
rect 786 -1650 787 -1636
rect 828 -1713 829 -1649
rect 912 -1713 913 -1649
rect 996 -1650 997 -1636
rect 61 -1652 62 -1636
rect 663 -1713 664 -1651
rect 684 -1652 685 -1636
rect 891 -1652 892 -1636
rect 65 -1654 66 -1636
rect 100 -1713 101 -1653
rect 142 -1713 143 -1653
rect 177 -1654 178 -1636
rect 187 -1654 188 -1636
rect 506 -1654 507 -1636
rect 586 -1713 587 -1653
rect 1087 -1654 1088 -1636
rect 51 -1713 52 -1655
rect 79 -1713 80 -1655
rect 380 -1656 381 -1636
rect 394 -1656 395 -1636
rect 446 -1656 447 -1636
rect 450 -1713 451 -1655
rect 590 -1656 591 -1636
rect 611 -1713 612 -1655
rect 656 -1713 657 -1655
rect 691 -1713 692 -1655
rect 716 -1656 717 -1636
rect 730 -1656 731 -1636
rect 835 -1713 836 -1655
rect 891 -1713 892 -1655
rect 1010 -1656 1011 -1636
rect 82 -1658 83 -1636
rect 436 -1658 437 -1636
rect 460 -1658 461 -1636
rect 821 -1658 822 -1636
rect 93 -1713 94 -1659
rect 128 -1660 129 -1636
rect 149 -1713 150 -1659
rect 226 -1660 227 -1636
rect 254 -1660 255 -1636
rect 331 -1713 332 -1659
rect 380 -1713 381 -1659
rect 758 -1660 759 -1636
rect 786 -1713 787 -1659
rect 870 -1660 871 -1636
rect 54 -1713 55 -1661
rect 128 -1713 129 -1661
rect 159 -1713 160 -1661
rect 457 -1662 458 -1636
rect 506 -1713 507 -1661
rect 541 -1662 542 -1636
rect 590 -1713 591 -1661
rect 597 -1662 598 -1636
rect 614 -1662 615 -1636
rect 898 -1662 899 -1636
rect 96 -1664 97 -1636
rect 107 -1664 108 -1636
rect 170 -1664 171 -1636
rect 362 -1713 363 -1663
rect 401 -1664 402 -1636
rect 625 -1664 626 -1636
rect 639 -1664 640 -1636
rect 660 -1713 661 -1663
rect 667 -1664 668 -1636
rect 758 -1713 759 -1663
rect 765 -1664 766 -1636
rect 870 -1713 871 -1663
rect 898 -1713 899 -1663
rect 961 -1664 962 -1636
rect 72 -1666 73 -1636
rect 107 -1713 108 -1665
rect 156 -1666 157 -1636
rect 170 -1713 171 -1665
rect 191 -1666 192 -1636
rect 863 -1666 864 -1636
rect 961 -1713 962 -1665
rect 982 -1666 983 -1636
rect 72 -1713 73 -1667
rect 86 -1668 87 -1636
rect 191 -1713 192 -1667
rect 205 -1668 206 -1636
rect 226 -1713 227 -1667
rect 240 -1668 241 -1636
rect 254 -1713 255 -1667
rect 261 -1668 262 -1636
rect 296 -1668 297 -1636
rect 327 -1668 328 -1636
rect 387 -1668 388 -1636
rect 401 -1713 402 -1667
rect 422 -1668 423 -1636
rect 674 -1713 675 -1667
rect 681 -1668 682 -1636
rect 765 -1713 766 -1667
rect 821 -1713 822 -1667
rect 919 -1668 920 -1636
rect 86 -1713 87 -1669
rect 212 -1670 213 -1636
rect 240 -1713 241 -1669
rect 366 -1670 367 -1636
rect 387 -1713 388 -1669
rect 569 -1670 570 -1636
rect 597 -1713 598 -1669
rect 653 -1670 654 -1636
rect 695 -1713 696 -1669
rect 751 -1670 752 -1636
rect 842 -1670 843 -1636
rect 863 -1713 864 -1669
rect 919 -1713 920 -1669
rect 1031 -1670 1032 -1636
rect 65 -1713 66 -1671
rect 653 -1713 654 -1671
rect 702 -1672 703 -1636
rect 779 -1713 780 -1671
rect 842 -1713 843 -1671
rect 954 -1672 955 -1636
rect 163 -1674 164 -1636
rect 261 -1713 262 -1673
rect 296 -1713 297 -1673
rect 310 -1674 311 -1636
rect 317 -1674 318 -1636
rect 355 -1713 356 -1673
rect 366 -1713 367 -1673
rect 492 -1674 493 -1636
rect 618 -1674 619 -1636
rect 1062 -1674 1063 -1636
rect 163 -1713 164 -1675
rect 376 -1713 377 -1675
rect 422 -1713 423 -1675
rect 537 -1676 538 -1636
rect 618 -1713 619 -1675
rect 688 -1676 689 -1636
rect 702 -1713 703 -1675
rect 807 -1676 808 -1636
rect 954 -1713 955 -1675
rect 1080 -1676 1081 -1636
rect 201 -1678 202 -1636
rect 394 -1713 395 -1677
rect 425 -1678 426 -1636
rect 905 -1678 906 -1636
rect 205 -1713 206 -1679
rect 289 -1680 290 -1636
rect 317 -1713 318 -1679
rect 359 -1680 360 -1636
rect 429 -1680 430 -1636
rect 436 -1713 437 -1679
rect 457 -1713 458 -1679
rect 464 -1680 465 -1636
rect 471 -1680 472 -1636
rect 667 -1713 668 -1679
rect 716 -1713 717 -1679
rect 793 -1680 794 -1636
rect 807 -1713 808 -1679
rect 975 -1680 976 -1636
rect 212 -1713 213 -1681
rect 415 -1682 416 -1636
rect 464 -1713 465 -1681
rect 513 -1682 514 -1636
rect 625 -1713 626 -1681
rect 709 -1682 710 -1636
rect 730 -1713 731 -1681
rect 933 -1682 934 -1636
rect 233 -1684 234 -1636
rect 310 -1713 311 -1683
rect 327 -1713 328 -1683
rect 849 -1684 850 -1636
rect 905 -1713 906 -1683
rect 940 -1684 941 -1636
rect 184 -1686 185 -1636
rect 849 -1713 850 -1685
rect 933 -1713 934 -1685
rect 1045 -1686 1046 -1636
rect 44 -1688 45 -1636
rect 184 -1713 185 -1687
rect 233 -1713 234 -1687
rect 338 -1688 339 -1636
rect 359 -1713 360 -1687
rect 569 -1713 570 -1687
rect 632 -1688 633 -1636
rect 681 -1713 682 -1687
rect 709 -1713 710 -1687
rect 737 -1688 738 -1636
rect 744 -1688 745 -1636
rect 793 -1713 794 -1687
rect 940 -1713 941 -1687
rect 1038 -1688 1039 -1636
rect 44 -1713 45 -1689
rect 68 -1713 69 -1689
rect 268 -1690 269 -1636
rect 289 -1713 290 -1689
rect 373 -1690 374 -1636
rect 429 -1713 430 -1689
rect 471 -1713 472 -1689
rect 499 -1690 500 -1636
rect 513 -1713 514 -1689
rect 562 -1690 563 -1636
rect 639 -1713 640 -1689
rect 646 -1690 647 -1636
rect 737 -1713 738 -1689
rect 877 -1690 878 -1636
rect 268 -1713 269 -1691
rect 275 -1692 276 -1636
rect 373 -1713 374 -1691
rect 772 -1692 773 -1636
rect 877 -1713 878 -1691
rect 1052 -1692 1053 -1636
rect 415 -1713 416 -1693
rect 527 -1694 528 -1636
rect 646 -1713 647 -1693
rect 677 -1694 678 -1636
rect 723 -1694 724 -1636
rect 772 -1713 773 -1693
rect 408 -1696 409 -1636
rect 527 -1713 528 -1695
rect 723 -1713 724 -1695
rect 814 -1696 815 -1636
rect 408 -1713 409 -1697
rect 579 -1713 580 -1697
rect 744 -1713 745 -1697
rect 800 -1698 801 -1636
rect 478 -1700 479 -1636
rect 541 -1713 542 -1699
rect 751 -1713 752 -1699
rect 1024 -1700 1025 -1636
rect 30 -1702 31 -1636
rect 478 -1713 479 -1701
rect 481 -1713 482 -1701
rect 562 -1713 563 -1701
rect 800 -1713 801 -1701
rect 968 -1702 969 -1636
rect 30 -1713 31 -1703
rect 121 -1704 122 -1636
rect 488 -1713 489 -1703
rect 632 -1713 633 -1703
rect 968 -1713 969 -1703
rect 1003 -1704 1004 -1636
rect 121 -1713 122 -1705
rect 282 -1706 283 -1636
rect 499 -1713 500 -1705
rect 548 -1706 549 -1636
rect 282 -1713 283 -1707
rect 303 -1708 304 -1636
rect 548 -1713 549 -1707
rect 555 -1708 556 -1636
rect 275 -1713 276 -1709
rect 303 -1713 304 -1709
rect 555 -1713 556 -1709
rect 856 -1710 857 -1636
rect 856 -1713 857 -1711
rect 1017 -1712 1018 -1636
rect 2 -1804 3 -1722
rect 212 -1723 213 -1721
rect 254 -1723 255 -1721
rect 324 -1723 325 -1721
rect 338 -1804 339 -1722
rect 607 -1723 608 -1721
rect 653 -1723 654 -1721
rect 828 -1723 829 -1721
rect 849 -1723 850 -1721
rect 1017 -1804 1018 -1722
rect 1052 -1804 1053 -1722
rect 1069 -1723 1070 -1721
rect 1094 -1723 1095 -1721
rect 1094 -1804 1095 -1722
rect 1094 -1723 1095 -1721
rect 1094 -1804 1095 -1722
rect 16 -1804 17 -1724
rect 37 -1725 38 -1721
rect 51 -1804 52 -1724
rect 93 -1725 94 -1721
rect 100 -1725 101 -1721
rect 138 -1804 139 -1724
rect 159 -1725 160 -1721
rect 240 -1725 241 -1721
rect 261 -1725 262 -1721
rect 849 -1804 850 -1724
rect 870 -1725 871 -1721
rect 908 -1725 909 -1721
rect 919 -1725 920 -1721
rect 996 -1804 997 -1724
rect 1055 -1804 1056 -1724
rect 1087 -1804 1088 -1724
rect 30 -1727 31 -1721
rect 222 -1727 223 -1721
rect 226 -1727 227 -1721
rect 261 -1804 262 -1726
rect 275 -1727 276 -1721
rect 324 -1804 325 -1726
rect 359 -1804 360 -1726
rect 520 -1727 521 -1721
rect 527 -1727 528 -1721
rect 730 -1727 731 -1721
rect 758 -1804 759 -1726
rect 807 -1727 808 -1721
rect 817 -1727 818 -1721
rect 933 -1727 934 -1721
rect 940 -1727 941 -1721
rect 982 -1804 983 -1726
rect 23 -1729 24 -1721
rect 222 -1804 223 -1728
rect 233 -1729 234 -1721
rect 254 -1804 255 -1728
rect 275 -1804 276 -1728
rect 282 -1729 283 -1721
rect 296 -1729 297 -1721
rect 303 -1729 304 -1721
rect 366 -1729 367 -1721
rect 432 -1804 433 -1728
rect 436 -1729 437 -1721
rect 523 -1729 524 -1721
rect 527 -1804 528 -1728
rect 597 -1729 598 -1721
rect 632 -1729 633 -1721
rect 919 -1804 920 -1728
rect 926 -1729 927 -1721
rect 961 -1729 962 -1721
rect 30 -1804 31 -1730
rect 677 -1731 678 -1721
rect 681 -1731 682 -1721
rect 814 -1804 815 -1730
rect 828 -1804 829 -1730
rect 863 -1731 864 -1721
rect 877 -1731 878 -1721
rect 1003 -1804 1004 -1730
rect 37 -1804 38 -1732
rect 44 -1733 45 -1721
rect 65 -1733 66 -1721
rect 457 -1733 458 -1721
rect 478 -1804 479 -1732
rect 751 -1733 752 -1721
rect 761 -1733 762 -1721
rect 1045 -1804 1046 -1732
rect 44 -1804 45 -1734
rect 121 -1735 122 -1721
rect 170 -1735 171 -1721
rect 170 -1804 171 -1734
rect 170 -1735 171 -1721
rect 170 -1804 171 -1734
rect 177 -1735 178 -1721
rect 177 -1804 178 -1734
rect 177 -1735 178 -1721
rect 177 -1804 178 -1734
rect 212 -1804 213 -1734
rect 317 -1735 318 -1721
rect 366 -1804 367 -1734
rect 380 -1735 381 -1721
rect 408 -1735 409 -1721
rect 653 -1804 654 -1734
rect 660 -1735 661 -1721
rect 989 -1804 990 -1734
rect 65 -1804 66 -1736
rect 205 -1737 206 -1721
rect 219 -1804 220 -1736
rect 317 -1804 318 -1736
rect 380 -1804 381 -1736
rect 464 -1737 465 -1721
rect 495 -1737 496 -1721
rect 499 -1737 500 -1721
rect 534 -1737 535 -1721
rect 660 -1804 661 -1736
rect 674 -1737 675 -1721
rect 856 -1737 857 -1721
rect 863 -1804 864 -1736
rect 912 -1737 913 -1721
rect 926 -1804 927 -1736
rect 947 -1737 948 -1721
rect 954 -1737 955 -1721
rect 1024 -1804 1025 -1736
rect 79 -1739 80 -1721
rect 383 -1739 384 -1721
rect 408 -1804 409 -1738
rect 502 -1804 503 -1738
rect 506 -1739 507 -1721
rect 534 -1804 535 -1738
rect 586 -1739 587 -1721
rect 751 -1804 752 -1738
rect 779 -1739 780 -1721
rect 779 -1804 780 -1738
rect 779 -1739 780 -1721
rect 779 -1804 780 -1738
rect 793 -1739 794 -1721
rect 912 -1804 913 -1738
rect 929 -1739 930 -1721
rect 961 -1804 962 -1738
rect 79 -1804 80 -1740
rect 355 -1741 356 -1721
rect 425 -1741 426 -1721
rect 632 -1804 633 -1740
rect 667 -1741 668 -1721
rect 856 -1804 857 -1740
rect 891 -1741 892 -1721
rect 940 -1804 941 -1740
rect 947 -1804 948 -1740
rect 968 -1741 969 -1721
rect 86 -1743 87 -1721
rect 373 -1743 374 -1721
rect 443 -1743 444 -1721
rect 1031 -1804 1032 -1742
rect 86 -1804 87 -1744
rect 107 -1745 108 -1721
rect 121 -1804 122 -1744
rect 376 -1745 377 -1721
rect 443 -1804 444 -1744
rect 579 -1745 580 -1721
rect 597 -1804 598 -1744
rect 625 -1745 626 -1721
rect 667 -1804 668 -1744
rect 772 -1745 773 -1721
rect 842 -1745 843 -1721
rect 877 -1804 878 -1744
rect 891 -1804 892 -1744
rect 898 -1745 899 -1721
rect 905 -1745 906 -1721
rect 1038 -1804 1039 -1744
rect 100 -1804 101 -1746
rect 289 -1747 290 -1721
rect 296 -1804 297 -1746
rect 418 -1804 419 -1746
rect 450 -1747 451 -1721
rect 583 -1804 584 -1746
rect 670 -1804 671 -1746
rect 898 -1804 899 -1746
rect 107 -1804 108 -1748
rect 142 -1749 143 -1721
rect 156 -1749 157 -1721
rect 674 -1804 675 -1748
rect 681 -1804 682 -1748
rect 709 -1749 710 -1721
rect 716 -1749 717 -1721
rect 1059 -1804 1060 -1748
rect 135 -1751 136 -1721
rect 793 -1804 794 -1750
rect 800 -1751 801 -1721
rect 905 -1804 906 -1750
rect 23 -1804 24 -1752
rect 135 -1804 136 -1752
rect 142 -1804 143 -1752
rect 191 -1753 192 -1721
rect 198 -1753 199 -1721
rect 499 -1804 500 -1752
rect 506 -1804 507 -1752
rect 646 -1753 647 -1721
rect 688 -1753 689 -1721
rect 786 -1753 787 -1721
rect 156 -1804 157 -1754
rect 387 -1755 388 -1721
rect 450 -1804 451 -1754
rect 520 -1804 521 -1754
rect 569 -1755 570 -1721
rect 646 -1804 647 -1754
rect 688 -1804 689 -1754
rect 821 -1755 822 -1721
rect 163 -1757 164 -1721
rect 716 -1804 717 -1756
rect 723 -1757 724 -1721
rect 821 -1804 822 -1756
rect 149 -1759 150 -1721
rect 723 -1804 724 -1758
rect 730 -1804 731 -1758
rect 835 -1759 836 -1721
rect 149 -1804 150 -1760
rect 345 -1761 346 -1721
rect 348 -1804 349 -1760
rect 786 -1804 787 -1760
rect 163 -1804 164 -1762
rect 184 -1763 185 -1721
rect 191 -1804 192 -1762
rect 691 -1804 692 -1762
rect 702 -1763 703 -1721
rect 870 -1804 871 -1762
rect 114 -1765 115 -1721
rect 184 -1804 185 -1764
rect 198 -1804 199 -1764
rect 1010 -1804 1011 -1764
rect 226 -1804 227 -1766
rect 425 -1804 426 -1766
rect 457 -1804 458 -1766
rect 611 -1767 612 -1721
rect 625 -1804 626 -1766
rect 800 -1804 801 -1766
rect 233 -1804 234 -1768
rect 310 -1769 311 -1721
rect 373 -1804 374 -1768
rect 488 -1769 489 -1721
rect 576 -1769 577 -1721
rect 968 -1804 969 -1768
rect 128 -1771 129 -1721
rect 310 -1804 311 -1770
rect 387 -1804 388 -1770
rect 429 -1771 430 -1721
rect 464 -1804 465 -1770
rect 513 -1771 514 -1721
rect 611 -1804 612 -1770
rect 975 -1804 976 -1770
rect 128 -1804 129 -1772
rect 247 -1773 248 -1721
rect 268 -1773 269 -1721
rect 303 -1804 304 -1772
rect 306 -1804 307 -1772
rect 436 -1804 437 -1772
rect 485 -1773 486 -1721
rect 576 -1804 577 -1772
rect 639 -1773 640 -1721
rect 702 -1804 703 -1772
rect 737 -1773 738 -1721
rect 772 -1804 773 -1772
rect 240 -1804 241 -1774
rect 530 -1775 531 -1721
rect 618 -1775 619 -1721
rect 639 -1804 640 -1774
rect 695 -1775 696 -1721
rect 737 -1804 738 -1774
rect 744 -1775 745 -1721
rect 807 -1804 808 -1774
rect 268 -1804 269 -1776
rect 331 -1777 332 -1721
rect 352 -1777 353 -1721
rect 485 -1804 486 -1776
rect 492 -1777 493 -1721
rect 744 -1804 745 -1776
rect 765 -1777 766 -1721
rect 835 -1804 836 -1776
rect 58 -1779 59 -1721
rect 331 -1804 332 -1778
rect 352 -1804 353 -1778
rect 569 -1804 570 -1778
rect 600 -1804 601 -1778
rect 695 -1804 696 -1778
rect 712 -1804 713 -1778
rect 765 -1804 766 -1778
rect 58 -1804 59 -1780
rect 72 -1781 73 -1721
rect 282 -1804 283 -1780
rect 401 -1781 402 -1721
rect 415 -1781 416 -1721
rect 492 -1804 493 -1780
rect 72 -1804 73 -1782
rect 247 -1804 248 -1782
rect 289 -1804 290 -1782
rect 341 -1783 342 -1721
rect 362 -1783 363 -1721
rect 618 -1804 619 -1782
rect 394 -1785 395 -1721
rect 513 -1804 514 -1784
rect 394 -1804 395 -1786
rect 530 -1804 531 -1786
rect 401 -1804 402 -1788
rect 555 -1789 556 -1721
rect 415 -1804 416 -1790
rect 471 -1791 472 -1721
rect 555 -1804 556 -1790
rect 590 -1791 591 -1721
rect 429 -1804 430 -1792
rect 954 -1804 955 -1792
rect 471 -1804 472 -1794
rect 562 -1795 563 -1721
rect 590 -1804 591 -1794
rect 604 -1795 605 -1721
rect 541 -1797 542 -1721
rect 562 -1804 563 -1796
rect 604 -1804 605 -1796
rect 842 -1804 843 -1796
rect 541 -1804 542 -1798
rect 548 -1799 549 -1721
rect 548 -1804 549 -1800
rect 884 -1801 885 -1721
rect 117 -1804 118 -1802
rect 884 -1804 885 -1802
rect 2 -1814 3 -1812
rect 425 -1814 426 -1812
rect 443 -1814 444 -1812
rect 453 -1872 454 -1813
rect 499 -1814 500 -1812
rect 870 -1814 871 -1812
rect 933 -1814 934 -1812
rect 947 -1814 948 -1812
rect 968 -1814 969 -1812
rect 968 -1895 969 -1813
rect 968 -1814 969 -1812
rect 968 -1895 969 -1813
rect 1010 -1814 1011 -1812
rect 1052 -1895 1053 -1813
rect 1087 -1814 1088 -1812
rect 1101 -1895 1102 -1813
rect 5 -1895 6 -1815
rect 527 -1816 528 -1812
rect 555 -1816 556 -1812
rect 555 -1895 556 -1815
rect 555 -1816 556 -1812
rect 555 -1895 556 -1815
rect 604 -1816 605 -1812
rect 702 -1816 703 -1812
rect 709 -1816 710 -1812
rect 996 -1816 997 -1812
rect 1017 -1816 1018 -1812
rect 1073 -1895 1074 -1815
rect 1087 -1895 1088 -1815
rect 1094 -1816 1095 -1812
rect 37 -1818 38 -1812
rect 40 -1895 41 -1817
rect 54 -1895 55 -1817
rect 72 -1818 73 -1812
rect 79 -1818 80 -1812
rect 432 -1818 433 -1812
rect 443 -1895 444 -1817
rect 492 -1818 493 -1812
rect 502 -1895 503 -1817
rect 653 -1818 654 -1812
rect 667 -1895 668 -1817
rect 758 -1818 759 -1812
rect 828 -1818 829 -1812
rect 828 -1895 829 -1817
rect 828 -1818 829 -1812
rect 828 -1895 829 -1817
rect 912 -1818 913 -1812
rect 933 -1895 934 -1817
rect 975 -1818 976 -1812
rect 996 -1895 997 -1817
rect 1024 -1818 1025 -1812
rect 1024 -1895 1025 -1817
rect 1024 -1818 1025 -1812
rect 1024 -1895 1025 -1817
rect 1045 -1818 1046 -1812
rect 1055 -1818 1056 -1812
rect 47 -1895 48 -1819
rect 72 -1895 73 -1819
rect 93 -1820 94 -1812
rect 849 -1820 850 -1812
rect 891 -1820 892 -1812
rect 912 -1895 913 -1819
rect 926 -1820 927 -1812
rect 1017 -1895 1018 -1819
rect 58 -1822 59 -1812
rect 58 -1895 59 -1821
rect 58 -1822 59 -1812
rect 58 -1895 59 -1821
rect 103 -1822 104 -1812
rect 373 -1822 374 -1812
rect 387 -1822 388 -1812
rect 635 -1895 636 -1821
rect 646 -1822 647 -1812
rect 870 -1895 871 -1821
rect 891 -1895 892 -1821
rect 940 -1822 941 -1812
rect 954 -1822 955 -1812
rect 975 -1895 976 -1821
rect 114 -1824 115 -1812
rect 261 -1824 262 -1812
rect 268 -1824 269 -1812
rect 362 -1895 363 -1823
rect 373 -1895 374 -1823
rect 712 -1824 713 -1812
rect 733 -1895 734 -1823
rect 905 -1824 906 -1812
rect 919 -1824 920 -1812
rect 940 -1895 941 -1823
rect 93 -1895 94 -1825
rect 114 -1895 115 -1825
rect 121 -1826 122 -1812
rect 184 -1895 185 -1825
rect 198 -1826 199 -1812
rect 793 -1826 794 -1812
rect 863 -1826 864 -1812
rect 926 -1895 927 -1825
rect 121 -1895 122 -1827
rect 583 -1828 584 -1812
rect 590 -1828 591 -1812
rect 646 -1895 647 -1827
rect 688 -1895 689 -1827
rect 1069 -1895 1070 -1827
rect 124 -1895 125 -1829
rect 219 -1830 220 -1812
rect 226 -1830 227 -1812
rect 418 -1830 419 -1812
rect 429 -1830 430 -1812
rect 947 -1895 948 -1829
rect 135 -1832 136 -1812
rect 1010 -1895 1011 -1831
rect 135 -1895 136 -1833
rect 191 -1834 192 -1812
rect 194 -1895 195 -1833
rect 590 -1895 591 -1833
rect 611 -1834 612 -1812
rect 611 -1895 612 -1833
rect 611 -1834 612 -1812
rect 611 -1895 612 -1833
rect 614 -1834 615 -1812
rect 821 -1834 822 -1812
rect 877 -1834 878 -1812
rect 905 -1895 906 -1833
rect 163 -1836 164 -1812
rect 352 -1836 353 -1812
rect 366 -1836 367 -1812
rect 877 -1895 878 -1835
rect 884 -1836 885 -1812
rect 919 -1895 920 -1835
rect 163 -1895 164 -1837
rect 551 -1838 552 -1812
rect 569 -1838 570 -1812
rect 709 -1895 710 -1837
rect 737 -1838 738 -1812
rect 849 -1895 850 -1837
rect 898 -1838 899 -1812
rect 954 -1895 955 -1837
rect 198 -1895 199 -1839
rect 359 -1840 360 -1812
rect 394 -1840 395 -1812
rect 604 -1895 605 -1839
rect 628 -1840 629 -1812
rect 681 -1840 682 -1812
rect 695 -1840 696 -1812
rect 702 -1895 703 -1839
rect 723 -1840 724 -1812
rect 737 -1895 738 -1839
rect 751 -1840 752 -1812
rect 758 -1895 759 -1839
rect 765 -1840 766 -1812
rect 898 -1895 899 -1839
rect 201 -1842 202 -1812
rect 268 -1895 269 -1841
rect 282 -1842 283 -1812
rect 387 -1895 388 -1841
rect 401 -1842 402 -1812
rect 401 -1895 402 -1841
rect 401 -1842 402 -1812
rect 401 -1895 402 -1841
rect 415 -1842 416 -1812
rect 751 -1895 752 -1841
rect 772 -1842 773 -1812
rect 863 -1895 864 -1841
rect 208 -1844 209 -1812
rect 233 -1844 234 -1812
rect 250 -1844 251 -1812
rect 618 -1844 619 -1812
rect 695 -1895 696 -1843
rect 716 -1844 717 -1812
rect 723 -1895 724 -1843
rect 800 -1844 801 -1812
rect 814 -1844 815 -1812
rect 821 -1895 822 -1843
rect 842 -1844 843 -1812
rect 884 -1895 885 -1843
rect 226 -1895 227 -1845
rect 558 -1895 559 -1845
rect 576 -1846 577 -1812
rect 793 -1895 794 -1845
rect 800 -1895 801 -1845
rect 807 -1846 808 -1812
rect 814 -1895 815 -1845
rect 1059 -1846 1060 -1812
rect 233 -1895 234 -1847
rect 471 -1848 472 -1812
rect 481 -1895 482 -1847
rect 716 -1895 717 -1847
rect 730 -1848 731 -1812
rect 772 -1895 773 -1847
rect 786 -1848 787 -1812
rect 842 -1895 843 -1847
rect 1031 -1848 1032 -1812
rect 1059 -1895 1060 -1847
rect 254 -1850 255 -1812
rect 359 -1895 360 -1849
rect 366 -1895 367 -1849
rect 576 -1895 577 -1849
rect 583 -1895 584 -1849
rect 625 -1850 626 -1812
rect 691 -1850 692 -1812
rect 807 -1895 808 -1849
rect 989 -1850 990 -1812
rect 1031 -1895 1032 -1849
rect 100 -1852 101 -1812
rect 254 -1895 255 -1851
rect 261 -1895 262 -1851
rect 436 -1852 437 -1812
rect 457 -1852 458 -1812
rect 681 -1895 682 -1851
rect 744 -1852 745 -1812
rect 765 -1895 766 -1851
rect 779 -1852 780 -1812
rect 786 -1895 787 -1851
rect 961 -1852 962 -1812
rect 989 -1895 990 -1851
rect 100 -1895 101 -1853
rect 205 -1854 206 -1812
rect 282 -1895 283 -1853
rect 408 -1854 409 -1812
rect 418 -1895 419 -1853
rect 429 -1895 430 -1853
rect 436 -1895 437 -1853
rect 670 -1854 671 -1812
rect 835 -1854 836 -1812
rect 961 -1895 962 -1853
rect 149 -1856 150 -1812
rect 457 -1895 458 -1855
rect 485 -1856 486 -1812
rect 653 -1895 654 -1855
rect 23 -1858 24 -1812
rect 485 -1895 486 -1857
rect 488 -1895 489 -1857
rect 744 -1895 745 -1857
rect 23 -1895 24 -1859
rect 310 -1860 311 -1812
rect 317 -1860 318 -1812
rect 345 -1895 346 -1859
rect 352 -1895 353 -1859
rect 464 -1860 465 -1812
rect 492 -1895 493 -1859
rect 506 -1860 507 -1812
rect 520 -1860 521 -1812
rect 856 -1860 857 -1812
rect 65 -1862 66 -1812
rect 310 -1895 311 -1861
rect 317 -1895 318 -1861
rect 355 -1862 356 -1812
rect 394 -1895 395 -1861
rect 670 -1895 671 -1861
rect 65 -1895 66 -1863
rect 82 -1895 83 -1863
rect 205 -1895 206 -1863
rect 240 -1864 241 -1812
rect 296 -1864 297 -1812
rect 523 -1864 524 -1812
rect 562 -1864 563 -1812
rect 625 -1895 626 -1863
rect 632 -1864 633 -1812
rect 856 -1895 857 -1863
rect 79 -1895 80 -1865
rect 520 -1895 521 -1865
rect 534 -1866 535 -1812
rect 562 -1895 563 -1865
rect 569 -1895 570 -1865
rect 730 -1895 731 -1865
rect 117 -1868 118 -1812
rect 240 -1895 241 -1867
rect 303 -1895 304 -1867
rect 380 -1868 381 -1812
rect 408 -1895 409 -1867
rect 446 -1895 447 -1867
rect 450 -1868 451 -1812
rect 464 -1895 465 -1867
rect 621 -1895 622 -1867
rect 835 -1895 836 -1867
rect 117 -1895 118 -1869
rect 338 -1870 339 -1812
rect 450 -1895 451 -1869
rect 597 -1895 598 -1869
rect 632 -1895 633 -1869
rect 1038 -1870 1039 -1812
rect 16 -1872 17 -1812
rect 338 -1895 339 -1871
rect 506 -1895 507 -1871
rect 639 -1872 640 -1812
rect 779 -1895 780 -1871
rect 1003 -1872 1004 -1812
rect 1038 -1895 1039 -1871
rect 128 -1874 129 -1812
rect 296 -1895 297 -1873
rect 306 -1874 307 -1812
rect 674 -1874 675 -1812
rect 982 -1874 983 -1812
rect 1003 -1895 1004 -1873
rect 86 -1876 87 -1812
rect 128 -1895 129 -1875
rect 177 -1876 178 -1812
rect 534 -1895 535 -1875
rect 548 -1895 549 -1875
rect 674 -1895 675 -1875
rect 86 -1895 87 -1877
rect 247 -1878 248 -1812
rect 289 -1878 290 -1812
rect 380 -1895 381 -1877
rect 422 -1878 423 -1812
rect 982 -1895 983 -1877
rect 9 -1880 10 -1812
rect 422 -1895 423 -1879
rect 513 -1880 514 -1812
rect 639 -1895 640 -1879
rect 9 -1895 10 -1881
rect 16 -1895 17 -1881
rect 142 -1882 143 -1812
rect 177 -1895 178 -1881
rect 212 -1882 213 -1812
rect 247 -1895 248 -1881
rect 275 -1882 276 -1812
rect 289 -1895 290 -1881
rect 324 -1882 325 -1812
rect 369 -1895 370 -1881
rect 513 -1895 514 -1881
rect 541 -1882 542 -1812
rect 96 -1884 97 -1812
rect 142 -1895 143 -1883
rect 156 -1884 157 -1812
rect 324 -1895 325 -1883
rect 331 -1884 332 -1812
rect 471 -1895 472 -1883
rect 30 -1886 31 -1812
rect 156 -1895 157 -1885
rect 170 -1886 171 -1812
rect 212 -1895 213 -1885
rect 331 -1895 332 -1885
rect 478 -1886 479 -1812
rect 30 -1895 31 -1887
rect 44 -1888 45 -1812
rect 107 -1888 108 -1812
rect 275 -1895 276 -1887
rect 390 -1895 391 -1887
rect 541 -1895 542 -1887
rect 44 -1895 45 -1889
rect 1045 -1895 1046 -1889
rect 51 -1892 52 -1812
rect 107 -1895 108 -1891
rect 170 -1895 171 -1891
rect 348 -1892 349 -1812
rect 478 -1895 479 -1891
rect 660 -1892 661 -1812
rect 51 -1895 52 -1893
rect 68 -1895 69 -1893
rect 551 -1895 552 -1893
rect 660 -1895 661 -1893
rect 2 -2000 3 -1904
rect 527 -1905 528 -1903
rect 530 -1905 531 -1903
rect 1031 -1905 1032 -1903
rect 1073 -1905 1074 -1903
rect 1108 -2000 1109 -1904
rect 9 -1907 10 -1903
rect 40 -1907 41 -1903
rect 44 -1907 45 -1903
rect 128 -1907 129 -1903
rect 142 -1907 143 -1903
rect 191 -2000 192 -1906
rect 194 -1907 195 -1903
rect 492 -1907 493 -1903
rect 502 -1907 503 -1903
rect 534 -1907 535 -1903
rect 551 -1907 552 -1903
rect 849 -1907 850 -1903
rect 1003 -1907 1004 -1903
rect 1031 -2000 1032 -1906
rect 1045 -1907 1046 -1903
rect 1073 -2000 1074 -1906
rect 1080 -2000 1081 -1906
rect 1087 -1907 1088 -1903
rect 1101 -1907 1102 -1903
rect 1115 -2000 1116 -1906
rect 9 -2000 10 -1908
rect 100 -1909 101 -1903
rect 114 -2000 115 -1908
rect 135 -1909 136 -1903
rect 149 -1909 150 -1903
rect 268 -1909 269 -1903
rect 296 -1909 297 -1903
rect 366 -1909 367 -1903
rect 369 -1909 370 -1903
rect 702 -1909 703 -1903
rect 786 -1909 787 -1903
rect 786 -2000 787 -1908
rect 786 -1909 787 -1903
rect 786 -2000 787 -1908
rect 821 -1909 822 -1903
rect 824 -1935 825 -1908
rect 842 -1909 843 -1903
rect 1066 -1909 1067 -1903
rect 16 -2000 17 -1910
rect 481 -1911 482 -1903
rect 485 -1911 486 -1903
rect 695 -1911 696 -1903
rect 702 -2000 703 -1910
rect 1097 -2000 1098 -1910
rect 19 -1913 20 -1903
rect 422 -1913 423 -1903
rect 429 -1913 430 -1903
rect 429 -2000 430 -1912
rect 429 -1913 430 -1903
rect 429 -2000 430 -1912
rect 443 -2000 444 -1912
rect 604 -1913 605 -1903
rect 618 -1913 619 -1903
rect 919 -1913 920 -1903
rect 968 -1913 969 -1903
rect 1003 -2000 1004 -1912
rect 1024 -1913 1025 -1903
rect 1087 -2000 1088 -1912
rect 30 -1915 31 -1903
rect 30 -2000 31 -1914
rect 30 -1915 31 -1903
rect 30 -2000 31 -1914
rect 33 -2000 34 -1914
rect 1045 -2000 1046 -1914
rect 37 -2000 38 -1916
rect 394 -1917 395 -1903
rect 450 -2000 451 -1916
rect 457 -1917 458 -1903
rect 471 -1917 472 -1903
rect 492 -2000 493 -1916
rect 516 -2000 517 -1916
rect 870 -1917 871 -1903
rect 968 -2000 969 -1916
rect 996 -1917 997 -1903
rect 47 -1919 48 -1903
rect 975 -1919 976 -1903
rect 51 -1921 52 -1903
rect 58 -1921 59 -1903
rect 65 -2000 66 -1920
rect 72 -1921 73 -1903
rect 75 -2000 76 -1920
rect 499 -1921 500 -1903
rect 527 -2000 528 -1920
rect 1038 -1921 1039 -1903
rect 58 -2000 59 -1922
rect 394 -2000 395 -1922
rect 453 -1923 454 -1903
rect 1066 -2000 1067 -1922
rect 82 -1925 83 -1903
rect 247 -1925 248 -1903
rect 324 -1925 325 -1903
rect 604 -2000 605 -1924
rect 618 -2000 619 -1924
rect 856 -1925 857 -1903
rect 870 -2000 871 -1924
rect 933 -1925 934 -1903
rect 947 -1925 948 -1903
rect 975 -2000 976 -1924
rect 93 -1927 94 -1903
rect 534 -2000 535 -1926
rect 555 -2000 556 -1926
rect 744 -1927 745 -1903
rect 768 -2000 769 -1926
rect 919 -2000 920 -1926
rect 926 -1927 927 -1903
rect 947 -2000 948 -1926
rect 954 -1927 955 -1903
rect 996 -2000 997 -1926
rect 93 -2000 94 -1928
rect 219 -2000 220 -1928
rect 222 -1929 223 -1903
rect 289 -1929 290 -1903
rect 324 -2000 325 -1928
rect 464 -1929 465 -1903
rect 471 -2000 472 -1928
rect 506 -1929 507 -1903
rect 558 -1929 559 -1903
rect 842 -2000 843 -1928
rect 856 -2000 857 -1928
rect 1069 -1929 1070 -1903
rect 100 -2000 101 -1930
rect 345 -1931 346 -1903
rect 348 -2000 349 -1930
rect 408 -1931 409 -1903
rect 478 -1931 479 -1903
rect 478 -2000 479 -1930
rect 478 -1931 479 -1903
rect 478 -2000 479 -1930
rect 485 -2000 486 -1930
rect 576 -1931 577 -1903
rect 621 -1931 622 -1903
rect 793 -1931 794 -1903
rect 821 -2000 822 -1930
rect 828 -1931 829 -1903
rect 912 -1931 913 -1903
rect 933 -2000 934 -1930
rect 940 -1931 941 -1903
rect 954 -2000 955 -1930
rect 124 -1933 125 -1903
rect 1059 -1933 1060 -1903
rect 128 -2000 129 -1934
rect 376 -2000 377 -1934
rect 387 -2000 388 -1934
rect 401 -1935 402 -1903
rect 506 -2000 507 -1934
rect 737 -1935 738 -1903
rect 828 -2000 829 -1934
rect 835 -1935 836 -1903
rect 940 -2000 941 -1934
rect 1010 -1935 1011 -1903
rect 1059 -2000 1060 -1934
rect 152 -1937 153 -1903
rect 877 -1937 878 -1903
rect 898 -1937 899 -1903
rect 912 -2000 913 -1936
rect 23 -1939 24 -1903
rect 898 -2000 899 -1938
rect 44 -2000 45 -1940
rect 152 -2000 153 -1940
rect 156 -1941 157 -1903
rect 835 -2000 836 -1940
rect 877 -2000 878 -1940
rect 891 -1941 892 -1903
rect 107 -1943 108 -1903
rect 156 -2000 157 -1942
rect 159 -1943 160 -1903
rect 1024 -2000 1025 -1942
rect 107 -2000 108 -1944
rect 142 -2000 143 -1944
rect 184 -1945 185 -1903
rect 268 -2000 269 -1944
rect 338 -1945 339 -1903
rect 457 -2000 458 -1944
rect 562 -1945 563 -1903
rect 562 -2000 563 -1944
rect 562 -1945 563 -1903
rect 562 -2000 563 -1944
rect 576 -2000 577 -1944
rect 611 -1945 612 -1903
rect 621 -2000 622 -1944
rect 1052 -1945 1053 -1903
rect 184 -2000 185 -1946
rect 366 -2000 367 -1946
rect 369 -2000 370 -1946
rect 408 -2000 409 -1946
rect 583 -1947 584 -1903
rect 611 -2000 612 -1946
rect 632 -1947 633 -1903
rect 1038 -2000 1039 -1946
rect 198 -1949 199 -1903
rect 289 -2000 290 -1948
rect 338 -2000 339 -1948
rect 646 -1949 647 -1903
rect 660 -1949 661 -1903
rect 793 -2000 794 -1948
rect 1017 -1949 1018 -1903
rect 1052 -2000 1053 -1948
rect 198 -2000 199 -1950
rect 282 -1951 283 -1903
rect 345 -2000 346 -1950
rect 401 -2000 402 -1950
rect 569 -1951 570 -1903
rect 583 -2000 584 -1950
rect 635 -1951 636 -1903
rect 723 -1951 724 -1903
rect 989 -1951 990 -1903
rect 1017 -2000 1018 -1950
rect 23 -2000 24 -1952
rect 723 -2000 724 -1952
rect 807 -1953 808 -1903
rect 989 -2000 990 -1952
rect 54 -1955 55 -1903
rect 569 -2000 570 -1954
rect 635 -2000 636 -1954
rect 772 -1955 773 -1903
rect 807 -2000 808 -1954
rect 884 -1955 885 -1903
rect 54 -2000 55 -1956
rect 226 -1957 227 -1903
rect 229 -2000 230 -1956
rect 296 -2000 297 -1956
rect 352 -1957 353 -1903
rect 415 -1957 416 -1903
rect 646 -2000 647 -1956
rect 905 -1957 906 -1903
rect 180 -2000 181 -1958
rect 415 -2000 416 -1958
rect 625 -1959 626 -1903
rect 905 -2000 906 -1958
rect 117 -1961 118 -1903
rect 625 -2000 626 -1960
rect 660 -2000 661 -1960
rect 779 -1961 780 -1903
rect 863 -1961 864 -1903
rect 884 -2000 885 -1960
rect 208 -2000 209 -1962
rect 982 -1963 983 -1903
rect 149 -2000 150 -1964
rect 982 -2000 983 -1964
rect 222 -2000 223 -1966
rect 261 -1967 262 -1903
rect 275 -1967 276 -1903
rect 282 -2000 283 -1966
rect 331 -1967 332 -1903
rect 352 -2000 353 -1966
rect 359 -1967 360 -1903
rect 1010 -2000 1011 -1966
rect 163 -1969 164 -1903
rect 275 -2000 276 -1968
rect 331 -2000 332 -1968
rect 373 -1969 374 -1903
rect 390 -1969 391 -1903
rect 891 -2000 892 -1968
rect 163 -2000 164 -1970
rect 530 -2000 531 -1970
rect 670 -1971 671 -1903
rect 849 -2000 850 -1970
rect 240 -1973 241 -1903
rect 422 -2000 423 -1972
rect 681 -1973 682 -1903
rect 737 -2000 738 -1972
rect 751 -1973 752 -1903
rect 863 -2000 864 -1972
rect 240 -2000 241 -1974
rect 254 -1975 255 -1903
rect 359 -2000 360 -1974
rect 380 -1975 381 -1903
rect 667 -1975 668 -1903
rect 681 -2000 682 -1974
rect 688 -1975 689 -1903
rect 961 -1975 962 -1903
rect 86 -1977 87 -1903
rect 380 -2000 381 -1976
rect 520 -1977 521 -1903
rect 667 -2000 668 -1976
rect 674 -1977 675 -1903
rect 961 -2000 962 -1976
rect 61 -2000 62 -1978
rect 520 -2000 521 -1978
rect 597 -1979 598 -1903
rect 688 -2000 689 -1978
rect 695 -2000 696 -1978
rect 709 -1979 710 -1903
rect 751 -2000 752 -1978
rect 814 -1979 815 -1903
rect 233 -1981 234 -1903
rect 597 -2000 598 -1980
rect 649 -2000 650 -1980
rect 814 -2000 815 -1980
rect 212 -1983 213 -1903
rect 233 -2000 234 -1982
rect 247 -2000 248 -1982
rect 730 -1983 731 -1903
rect 758 -1983 759 -1903
rect 772 -2000 773 -1982
rect 121 -1985 122 -1903
rect 212 -2000 213 -1984
rect 254 -2000 255 -1984
rect 303 -1985 304 -1903
rect 373 -2000 374 -1984
rect 464 -2000 465 -1984
rect 653 -1985 654 -1903
rect 674 -2000 675 -1984
rect 709 -2000 710 -1984
rect 716 -1985 717 -1903
rect 730 -2000 731 -1984
rect 800 -1985 801 -1903
rect 121 -2000 122 -1986
rect 205 -1987 206 -1903
rect 303 -2000 304 -1986
rect 310 -1987 311 -1903
rect 548 -1987 549 -1903
rect 716 -2000 717 -1986
rect 758 -2000 759 -1986
rect 765 -1987 766 -1903
rect 170 -1989 171 -1903
rect 800 -2000 801 -1988
rect 170 -2000 171 -1990
rect 177 -1991 178 -1903
rect 205 -2000 206 -1990
rect 499 -2000 500 -1990
rect 548 -2000 549 -1990
rect 1104 -2000 1105 -1990
rect 310 -2000 311 -1992
rect 541 -1993 542 -1903
rect 639 -1993 640 -1903
rect 653 -2000 654 -1992
rect 317 -1995 318 -1903
rect 765 -2000 766 -1994
rect 317 -2000 318 -1996
rect 436 -1997 437 -1903
rect 513 -1997 514 -1903
rect 541 -2000 542 -1996
rect 590 -1997 591 -1903
rect 639 -2000 640 -1996
rect 261 -2000 262 -1998
rect 436 -2000 437 -1998
rect 2 -2113 3 -2009
rect 222 -2010 223 -2008
rect 229 -2010 230 -2008
rect 373 -2010 374 -2008
rect 376 -2010 377 -2008
rect 898 -2010 899 -2008
rect 919 -2010 920 -2008
rect 919 -2113 920 -2009
rect 919 -2010 920 -2008
rect 919 -2113 920 -2009
rect 926 -2113 927 -2009
rect 933 -2010 934 -2008
rect 943 -2113 944 -2009
rect 1017 -2010 1018 -2008
rect 1080 -2010 1081 -2008
rect 1094 -2010 1095 -2008
rect 1104 -2010 1105 -2008
rect 1108 -2010 1109 -2008
rect 1115 -2010 1116 -2008
rect 1122 -2113 1123 -2009
rect 9 -2012 10 -2008
rect 23 -2113 24 -2011
rect 30 -2012 31 -2008
rect 30 -2113 31 -2011
rect 30 -2012 31 -2008
rect 30 -2113 31 -2011
rect 33 -2012 34 -2008
rect 1024 -2012 1025 -2008
rect 1038 -2012 1039 -2008
rect 1080 -2113 1081 -2011
rect 9 -2113 10 -2013
rect 163 -2014 164 -2008
rect 170 -2014 171 -2008
rect 226 -2014 227 -2008
rect 275 -2014 276 -2008
rect 436 -2113 437 -2013
rect 439 -2014 440 -2008
rect 1066 -2014 1067 -2008
rect 1073 -2014 1074 -2008
rect 1108 -2113 1109 -2013
rect 16 -2016 17 -2008
rect 345 -2016 346 -2008
rect 348 -2016 349 -2008
rect 800 -2016 801 -2008
rect 807 -2016 808 -2008
rect 933 -2113 934 -2015
rect 947 -2016 948 -2008
rect 947 -2113 948 -2015
rect 947 -2016 948 -2008
rect 947 -2113 948 -2015
rect 982 -2016 983 -2008
rect 1017 -2113 1018 -2015
rect 1031 -2016 1032 -2008
rect 1038 -2113 1039 -2015
rect 1045 -2016 1046 -2008
rect 1073 -2113 1074 -2015
rect 16 -2113 17 -2017
rect 100 -2018 101 -2008
rect 107 -2018 108 -2008
rect 583 -2018 584 -2008
rect 593 -2018 594 -2008
rect 961 -2018 962 -2008
rect 996 -2018 997 -2008
rect 1024 -2113 1025 -2017
rect 1059 -2018 1060 -2008
rect 1094 -2113 1095 -2017
rect 51 -2020 52 -2008
rect 835 -2020 836 -2008
rect 863 -2020 864 -2008
rect 898 -2113 899 -2019
rect 929 -2020 930 -2008
rect 968 -2020 969 -2008
rect 1003 -2020 1004 -2008
rect 1045 -2113 1046 -2019
rect 54 -2022 55 -2008
rect 345 -2113 346 -2021
rect 380 -2022 381 -2008
rect 460 -2113 461 -2021
rect 464 -2022 465 -2008
rect 646 -2022 647 -2008
rect 688 -2022 689 -2008
rect 779 -2022 780 -2008
rect 782 -2022 783 -2008
rect 821 -2022 822 -2008
rect 835 -2113 836 -2021
rect 912 -2022 913 -2008
rect 940 -2022 941 -2008
rect 961 -2113 962 -2021
rect 975 -2022 976 -2008
rect 1003 -2113 1004 -2021
rect 1010 -2022 1011 -2008
rect 1066 -2113 1067 -2021
rect 37 -2024 38 -2008
rect 380 -2113 381 -2023
rect 394 -2024 395 -2008
rect 646 -2113 647 -2023
rect 691 -2113 692 -2023
rect 1059 -2113 1060 -2023
rect 37 -2113 38 -2025
rect 177 -2026 178 -2008
rect 180 -2026 181 -2008
rect 233 -2026 234 -2008
rect 275 -2113 276 -2025
rect 471 -2026 472 -2008
rect 502 -2113 503 -2025
rect 905 -2026 906 -2008
rect 954 -2026 955 -2008
rect 982 -2113 983 -2025
rect 44 -2028 45 -2008
rect 464 -2113 465 -2027
rect 471 -2113 472 -2027
rect 530 -2028 531 -2008
rect 569 -2028 570 -2008
rect 632 -2113 633 -2027
rect 716 -2028 717 -2008
rect 905 -2113 906 -2027
rect 44 -2113 45 -2029
rect 212 -2030 213 -2008
rect 222 -2113 223 -2029
rect 604 -2030 605 -2008
rect 611 -2030 612 -2008
rect 1115 -2113 1116 -2029
rect 58 -2032 59 -2008
rect 75 -2032 76 -2008
rect 79 -2032 80 -2008
rect 170 -2113 171 -2031
rect 177 -2113 178 -2031
rect 282 -2032 283 -2008
rect 324 -2032 325 -2008
rect 355 -2113 356 -2031
rect 394 -2113 395 -2031
rect 418 -2113 419 -2031
rect 478 -2032 479 -2008
rect 604 -2113 605 -2031
rect 625 -2032 626 -2008
rect 1031 -2113 1032 -2031
rect 58 -2113 59 -2033
rect 849 -2034 850 -2008
rect 870 -2034 871 -2008
rect 975 -2113 976 -2033
rect 65 -2036 66 -2008
rect 366 -2036 367 -2008
rect 408 -2036 409 -2008
rect 534 -2036 535 -2008
rect 579 -2113 580 -2035
rect 779 -2113 780 -2035
rect 821 -2113 822 -2035
rect 828 -2036 829 -2008
rect 842 -2036 843 -2008
rect 863 -2113 864 -2035
rect 877 -2036 878 -2008
rect 996 -2113 997 -2035
rect 65 -2113 66 -2037
rect 128 -2038 129 -2008
rect 135 -2038 136 -2008
rect 492 -2038 493 -2008
rect 513 -2113 514 -2037
rect 723 -2038 724 -2008
rect 744 -2038 745 -2008
rect 772 -2038 773 -2008
rect 842 -2113 843 -2037
rect 891 -2038 892 -2008
rect 51 -2113 52 -2039
rect 135 -2113 136 -2039
rect 149 -2040 150 -2008
rect 527 -2040 528 -2008
rect 534 -2113 535 -2039
rect 562 -2040 563 -2008
rect 667 -2040 668 -2008
rect 870 -2113 871 -2039
rect 884 -2040 885 -2008
rect 1010 -2113 1011 -2039
rect 72 -2113 73 -2041
rect 107 -2113 108 -2041
rect 110 -2042 111 -2008
rect 156 -2042 157 -2008
rect 184 -2042 185 -2008
rect 635 -2042 636 -2008
rect 695 -2042 696 -2008
rect 723 -2113 724 -2041
rect 751 -2042 752 -2008
rect 772 -2113 773 -2041
rect 891 -2113 892 -2041
rect 989 -2042 990 -2008
rect 75 -2113 76 -2043
rect 590 -2044 591 -2008
rect 695 -2113 696 -2043
rect 730 -2044 731 -2008
rect 758 -2044 759 -2008
rect 807 -2113 808 -2043
rect 79 -2113 80 -2045
rect 422 -2046 423 -2008
rect 429 -2046 430 -2008
rect 478 -2113 479 -2045
rect 492 -2113 493 -2045
rect 499 -2046 500 -2008
rect 506 -2046 507 -2008
rect 744 -2113 745 -2045
rect 761 -2113 762 -2045
rect 1087 -2046 1088 -2008
rect 86 -2048 87 -2008
rect 800 -2113 801 -2047
rect 814 -2048 815 -2008
rect 1087 -2113 1088 -2047
rect 86 -2113 87 -2049
rect 751 -2113 752 -2049
rect 765 -2050 766 -2008
rect 1052 -2050 1053 -2008
rect 96 -2113 97 -2051
rect 793 -2052 794 -2008
rect 100 -2113 101 -2053
rect 114 -2054 115 -2008
rect 117 -2113 118 -2053
rect 163 -2113 164 -2053
rect 184 -2113 185 -2053
rect 618 -2054 619 -2008
rect 688 -2113 689 -2053
rect 793 -2113 794 -2053
rect 114 -2113 115 -2055
rect 373 -2113 374 -2055
rect 401 -2056 402 -2008
rect 422 -2113 423 -2055
rect 443 -2056 444 -2008
rect 667 -2113 668 -2055
rect 709 -2056 710 -2008
rect 730 -2113 731 -2055
rect 768 -2056 769 -2008
rect 884 -2113 885 -2055
rect 121 -2058 122 -2008
rect 205 -2113 206 -2057
rect 226 -2113 227 -2057
rect 614 -2113 615 -2057
rect 618 -2113 619 -2057
rect 681 -2058 682 -2008
rect 786 -2058 787 -2008
rect 814 -2113 815 -2057
rect 82 -2113 83 -2059
rect 121 -2113 122 -2059
rect 128 -2113 129 -2059
rect 331 -2060 332 -2008
rect 338 -2060 339 -2008
rect 527 -2113 528 -2059
rect 555 -2060 556 -2008
rect 765 -2113 766 -2059
rect 110 -2113 111 -2061
rect 338 -2113 339 -2061
rect 366 -2113 367 -2061
rect 548 -2062 549 -2008
rect 572 -2113 573 -2061
rect 786 -2113 787 -2061
rect 138 -2064 139 -2008
rect 681 -2113 682 -2063
rect 138 -2113 139 -2065
rect 912 -2113 913 -2065
rect 142 -2068 143 -2008
rect 156 -2113 157 -2067
rect 198 -2068 199 -2008
rect 233 -2113 234 -2067
rect 247 -2068 248 -2008
rect 429 -2113 430 -2067
rect 443 -2113 444 -2067
rect 597 -2068 598 -2008
rect 674 -2068 675 -2008
rect 709 -2113 710 -2067
rect 26 -2070 27 -2008
rect 597 -2113 598 -2069
rect 89 -2072 90 -2008
rect 198 -2113 199 -2071
rect 247 -2113 248 -2071
rect 296 -2072 297 -2008
rect 310 -2072 311 -2008
rect 590 -2113 591 -2071
rect 89 -2113 90 -2073
rect 737 -2074 738 -2008
rect 149 -2113 150 -2075
rect 212 -2113 213 -2075
rect 254 -2076 255 -2008
rect 499 -2113 500 -2075
rect 516 -2076 517 -2008
rect 989 -2113 990 -2075
rect 152 -2078 153 -2008
rect 191 -2078 192 -2008
rect 240 -2078 241 -2008
rect 254 -2113 255 -2077
rect 282 -2113 283 -2077
rect 352 -2078 353 -2008
rect 369 -2078 370 -2008
rect 828 -2113 829 -2077
rect 152 -2113 153 -2079
rect 968 -2113 969 -2079
rect 191 -2113 192 -2081
rect 268 -2082 269 -2008
rect 289 -2082 290 -2008
rect 310 -2113 311 -2081
rect 324 -2113 325 -2081
rect 352 -2113 353 -2081
rect 387 -2082 388 -2008
rect 401 -2113 402 -2081
rect 411 -2082 412 -2008
rect 954 -2113 955 -2081
rect 240 -2113 241 -2083
rect 450 -2084 451 -2008
rect 457 -2084 458 -2008
rect 506 -2113 507 -2083
rect 520 -2084 521 -2008
rect 562 -2113 563 -2083
rect 576 -2084 577 -2008
rect 674 -2113 675 -2083
rect 737 -2113 738 -2083
rect 877 -2113 878 -2083
rect 142 -2113 143 -2085
rect 450 -2113 451 -2085
rect 541 -2086 542 -2008
rect 555 -2113 556 -2085
rect 268 -2113 269 -2087
rect 453 -2113 454 -2087
rect 541 -2113 542 -2087
rect 758 -2113 759 -2087
rect 289 -2113 290 -2089
rect 856 -2090 857 -2008
rect 296 -2113 297 -2091
rect 303 -2092 304 -2008
rect 317 -2092 318 -2008
rect 387 -2113 388 -2091
rect 411 -2113 412 -2091
rect 639 -2092 640 -2008
rect 303 -2113 304 -2093
rect 649 -2094 650 -2008
rect 317 -2113 318 -2095
rect 359 -2096 360 -2008
rect 415 -2096 416 -2008
rect 583 -2113 584 -2095
rect 639 -2113 640 -2095
rect 856 -2113 857 -2095
rect 261 -2098 262 -2008
rect 359 -2113 360 -2097
rect 415 -2113 416 -2097
rect 849 -2113 850 -2097
rect 93 -2100 94 -2008
rect 261 -2113 262 -2099
rect 331 -2113 332 -2099
rect 642 -2113 643 -2099
rect 93 -2113 94 -2101
rect 1101 -2102 1102 -2008
rect 341 -2113 342 -2103
rect 520 -2113 521 -2103
rect 548 -2113 549 -2103
rect 660 -2104 661 -2008
rect 716 -2113 717 -2103
rect 1101 -2113 1102 -2103
rect 485 -2106 486 -2008
rect 660 -2113 661 -2105
rect 485 -2113 486 -2107
rect 702 -2108 703 -2008
rect 653 -2110 654 -2008
rect 702 -2113 703 -2109
rect 653 -2113 654 -2111
rect 1052 -2113 1053 -2111
rect 9 -2123 10 -2121
rect 397 -2208 398 -2122
rect 401 -2123 402 -2121
rect 418 -2123 419 -2121
rect 432 -2208 433 -2122
rect 604 -2123 605 -2121
rect 611 -2123 612 -2121
rect 1115 -2123 1116 -2121
rect 9 -2208 10 -2124
rect 254 -2125 255 -2121
rect 275 -2125 276 -2121
rect 415 -2125 416 -2121
rect 436 -2125 437 -2121
rect 579 -2125 580 -2121
rect 590 -2125 591 -2121
rect 628 -2125 629 -2121
rect 642 -2125 643 -2121
rect 1010 -2125 1011 -2121
rect 1052 -2125 1053 -2121
rect 1055 -2208 1056 -2124
rect 1101 -2125 1102 -2121
rect 1122 -2125 1123 -2121
rect 16 -2127 17 -2121
rect 457 -2208 458 -2126
rect 485 -2127 486 -2121
rect 499 -2208 500 -2126
rect 523 -2208 524 -2126
rect 807 -2127 808 -2121
rect 821 -2127 822 -2121
rect 821 -2208 822 -2126
rect 821 -2127 822 -2121
rect 821 -2208 822 -2126
rect 849 -2127 850 -2121
rect 849 -2208 850 -2126
rect 849 -2127 850 -2121
rect 849 -2208 850 -2126
rect 873 -2208 874 -2126
rect 961 -2127 962 -2121
rect 16 -2208 17 -2128
rect 89 -2129 90 -2121
rect 93 -2129 94 -2121
rect 275 -2208 276 -2128
rect 282 -2129 283 -2121
rect 338 -2129 339 -2121
rect 359 -2129 360 -2121
rect 569 -2129 570 -2121
rect 576 -2129 577 -2121
rect 982 -2129 983 -2121
rect 23 -2131 24 -2121
rect 149 -2131 150 -2121
rect 152 -2131 153 -2121
rect 366 -2131 367 -2121
rect 373 -2131 374 -2121
rect 450 -2208 451 -2130
rect 485 -2208 486 -2130
rect 541 -2131 542 -2121
rect 548 -2131 549 -2121
rect 562 -2131 563 -2121
rect 565 -2208 566 -2130
rect 1017 -2131 1018 -2121
rect 23 -2208 24 -2132
rect 583 -2133 584 -2121
rect 604 -2208 605 -2132
rect 1045 -2133 1046 -2121
rect 30 -2135 31 -2121
rect 40 -2208 41 -2134
rect 58 -2135 59 -2121
rect 170 -2135 171 -2121
rect 173 -2208 174 -2134
rect 345 -2135 346 -2121
rect 366 -2208 367 -2134
rect 380 -2135 381 -2121
rect 394 -2135 395 -2121
rect 583 -2208 584 -2134
rect 611 -2208 612 -2134
rect 709 -2135 710 -2121
rect 730 -2135 731 -2121
rect 733 -2175 734 -2134
rect 737 -2135 738 -2121
rect 996 -2135 997 -2121
rect 1017 -2208 1018 -2134
rect 1094 -2135 1095 -2121
rect 51 -2137 52 -2121
rect 380 -2208 381 -2136
rect 401 -2208 402 -2136
rect 670 -2208 671 -2136
rect 684 -2208 685 -2136
rect 975 -2137 976 -2121
rect 982 -2208 983 -2136
rect 1087 -2137 1088 -2121
rect 51 -2208 52 -2138
rect 338 -2208 339 -2138
rect 376 -2208 377 -2138
rect 408 -2139 409 -2121
rect 415 -2208 416 -2138
rect 698 -2208 699 -2138
rect 723 -2139 724 -2121
rect 737 -2208 738 -2138
rect 807 -2208 808 -2138
rect 877 -2139 878 -2121
rect 884 -2139 885 -2121
rect 884 -2208 885 -2138
rect 884 -2139 885 -2121
rect 884 -2208 885 -2138
rect 898 -2139 899 -2121
rect 898 -2208 899 -2138
rect 898 -2139 899 -2121
rect 898 -2208 899 -2138
rect 940 -2208 941 -2138
rect 954 -2139 955 -2121
rect 961 -2208 962 -2138
rect 1024 -2139 1025 -2121
rect 1038 -2139 1039 -2121
rect 1045 -2208 1046 -2138
rect 58 -2208 59 -2140
rect 387 -2141 388 -2121
rect 408 -2208 409 -2140
rect 492 -2141 493 -2121
rect 530 -2141 531 -2121
rect 989 -2141 990 -2121
rect 61 -2143 62 -2121
rect 541 -2208 542 -2142
rect 548 -2208 549 -2142
rect 551 -2143 552 -2121
rect 555 -2143 556 -2121
rect 572 -2208 573 -2142
rect 593 -2208 594 -2142
rect 1024 -2208 1025 -2142
rect 72 -2145 73 -2121
rect 506 -2145 507 -2121
rect 534 -2145 535 -2121
rect 600 -2208 601 -2144
rect 625 -2145 626 -2121
rect 1003 -2145 1004 -2121
rect 75 -2147 76 -2121
rect 1010 -2208 1011 -2146
rect 75 -2208 76 -2148
rect 660 -2149 661 -2121
rect 691 -2149 692 -2121
rect 814 -2149 815 -2121
rect 891 -2149 892 -2121
rect 954 -2208 955 -2148
rect 989 -2208 990 -2148
rect 1108 -2149 1109 -2121
rect 79 -2151 80 -2121
rect 800 -2151 801 -2121
rect 814 -2208 815 -2150
rect 828 -2151 829 -2121
rect 835 -2151 836 -2121
rect 891 -2208 892 -2150
rect 947 -2151 948 -2121
rect 996 -2208 997 -2150
rect 1003 -2208 1004 -2150
rect 1080 -2151 1081 -2121
rect 79 -2208 80 -2152
rect 191 -2153 192 -2121
rect 219 -2208 220 -2152
rect 341 -2153 342 -2121
rect 443 -2153 444 -2121
rect 509 -2208 510 -2152
rect 534 -2208 535 -2152
rect 667 -2153 668 -2121
rect 695 -2153 696 -2121
rect 877 -2208 878 -2152
rect 947 -2208 948 -2152
rect 968 -2153 969 -2121
rect 86 -2155 87 -2121
rect 471 -2155 472 -2121
rect 527 -2155 528 -2121
rect 968 -2208 969 -2154
rect 72 -2208 73 -2156
rect 86 -2208 87 -2156
rect 93 -2208 94 -2156
rect 191 -2208 192 -2156
rect 226 -2157 227 -2121
rect 576 -2208 577 -2156
rect 625 -2208 626 -2156
rect 702 -2157 703 -2121
rect 730 -2208 731 -2156
rect 842 -2157 843 -2121
rect 96 -2159 97 -2121
rect 597 -2159 598 -2121
rect 653 -2208 654 -2158
rect 695 -2208 696 -2158
rect 702 -2208 703 -2158
rect 772 -2159 773 -2121
rect 786 -2159 787 -2121
rect 800 -2208 801 -2158
rect 828 -2208 829 -2158
rect 863 -2159 864 -2121
rect 100 -2161 101 -2121
rect 100 -2208 101 -2160
rect 100 -2161 101 -2121
rect 100 -2208 101 -2160
rect 107 -2161 108 -2121
rect 289 -2161 290 -2121
rect 317 -2161 318 -2121
rect 387 -2208 388 -2160
rect 443 -2208 444 -2160
rect 464 -2161 465 -2121
rect 471 -2208 472 -2160
rect 761 -2161 762 -2121
rect 765 -2161 766 -2121
rect 772 -2208 773 -2160
rect 779 -2161 780 -2121
rect 786 -2208 787 -2160
rect 835 -2208 836 -2160
rect 870 -2161 871 -2121
rect 37 -2163 38 -2121
rect 779 -2208 780 -2162
rect 863 -2208 864 -2162
rect 905 -2163 906 -2121
rect 44 -2165 45 -2121
rect 289 -2208 290 -2164
rect 320 -2208 321 -2164
rect 975 -2208 976 -2164
rect 44 -2208 45 -2166
rect 212 -2167 213 -2121
rect 226 -2208 227 -2166
rect 303 -2167 304 -2121
rect 324 -2167 325 -2121
rect 359 -2208 360 -2166
rect 453 -2167 454 -2121
rect 1038 -2208 1039 -2166
rect 107 -2208 108 -2168
rect 166 -2208 167 -2168
rect 177 -2169 178 -2121
rect 282 -2208 283 -2168
rect 303 -2208 304 -2168
rect 429 -2169 430 -2121
rect 464 -2208 465 -2168
rect 478 -2169 479 -2121
rect 527 -2208 528 -2168
rect 726 -2208 727 -2168
rect 744 -2169 745 -2121
rect 842 -2208 843 -2168
rect 905 -2208 906 -2168
rect 1031 -2169 1032 -2121
rect 65 -2171 66 -2121
rect 177 -2208 178 -2170
rect 198 -2171 199 -2121
rect 324 -2208 325 -2170
rect 345 -2208 346 -2170
rect 429 -2208 430 -2170
rect 555 -2208 556 -2170
rect 632 -2171 633 -2121
rect 656 -2171 657 -2121
rect 1073 -2171 1074 -2121
rect 65 -2208 66 -2172
rect 268 -2173 269 -2121
rect 422 -2173 423 -2121
rect 478 -2208 479 -2172
rect 597 -2208 598 -2172
rect 933 -2173 934 -2121
rect 110 -2175 111 -2121
rect 590 -2208 591 -2174
rect 632 -2208 633 -2174
rect 646 -2175 647 -2121
rect 660 -2208 661 -2174
rect 681 -2175 682 -2121
rect 744 -2208 745 -2174
rect 751 -2175 752 -2121
rect 765 -2208 766 -2174
rect 114 -2208 115 -2176
rect 121 -2177 122 -2121
rect 128 -2177 129 -2121
rect 135 -2208 136 -2176
rect 138 -2177 139 -2121
rect 856 -2177 857 -2121
rect 82 -2179 83 -2121
rect 128 -2208 129 -2178
rect 142 -2179 143 -2121
rect 502 -2208 503 -2178
rect 513 -2179 514 -2121
rect 751 -2208 752 -2178
rect 117 -2181 118 -2121
rect 793 -2181 794 -2121
rect 142 -2208 143 -2182
rect 240 -2183 241 -2121
rect 261 -2183 262 -2121
rect 341 -2208 342 -2182
rect 422 -2208 423 -2182
rect 740 -2183 741 -2121
rect 149 -2208 150 -2184
rect 156 -2185 157 -2121
rect 163 -2185 164 -2121
rect 254 -2208 255 -2184
rect 261 -2208 262 -2184
rect 296 -2185 297 -2121
rect 436 -2208 437 -2184
rect 933 -2208 934 -2184
rect 121 -2208 122 -2186
rect 296 -2208 297 -2186
rect 513 -2208 514 -2186
rect 723 -2208 724 -2186
rect 124 -2189 125 -2121
rect 156 -2208 157 -2188
rect 184 -2189 185 -2121
rect 240 -2208 241 -2188
rect 268 -2208 269 -2188
rect 331 -2189 332 -2121
rect 639 -2189 640 -2121
rect 793 -2208 794 -2188
rect 2 -2191 3 -2121
rect 639 -2208 640 -2190
rect 646 -2208 647 -2190
rect 674 -2191 675 -2121
rect 688 -2208 689 -2190
rect 856 -2208 857 -2190
rect 2 -2208 3 -2192
rect 758 -2193 759 -2121
rect 124 -2208 125 -2194
rect 1031 -2208 1032 -2194
rect 198 -2208 199 -2196
rect 355 -2208 356 -2196
rect 667 -2208 668 -2196
rect 1066 -2197 1067 -2121
rect 212 -2208 213 -2198
rect 292 -2199 293 -2121
rect 310 -2199 311 -2121
rect 331 -2208 332 -2198
rect 674 -2208 675 -2198
rect 716 -2199 717 -2121
rect 758 -2208 759 -2198
rect 912 -2199 913 -2121
rect 233 -2201 234 -2121
rect 439 -2208 440 -2200
rect 618 -2201 619 -2121
rect 716 -2208 717 -2200
rect 912 -2208 913 -2200
rect 919 -2201 920 -2121
rect 205 -2203 206 -2121
rect 233 -2208 234 -2202
rect 247 -2203 248 -2121
rect 310 -2208 311 -2202
rect 520 -2203 521 -2121
rect 618 -2208 619 -2202
rect 919 -2208 920 -2202
rect 926 -2203 927 -2121
rect 205 -2208 206 -2204
rect 492 -2208 493 -2204
rect 520 -2208 521 -2204
rect 709 -2208 710 -2204
rect 926 -2208 927 -2204
rect 1059 -2205 1060 -2121
rect 247 -2208 248 -2206
rect 607 -2208 608 -2206
rect 9 -2218 10 -2216
rect 205 -2218 206 -2216
rect 208 -2218 209 -2216
rect 639 -2218 640 -2216
rect 653 -2218 654 -2216
rect 670 -2218 671 -2216
rect 691 -2218 692 -2216
rect 863 -2218 864 -2216
rect 870 -2277 871 -2217
rect 968 -2218 969 -2216
rect 9 -2277 10 -2219
rect 338 -2220 339 -2216
rect 341 -2220 342 -2216
rect 485 -2220 486 -2216
rect 488 -2277 489 -2219
rect 779 -2220 780 -2216
rect 856 -2220 857 -2216
rect 929 -2277 930 -2219
rect 16 -2222 17 -2216
rect 103 -2277 104 -2221
rect 121 -2222 122 -2216
rect 254 -2222 255 -2216
rect 282 -2222 283 -2216
rect 317 -2222 318 -2216
rect 348 -2277 349 -2221
rect 366 -2222 367 -2216
rect 373 -2277 374 -2221
rect 471 -2222 472 -2216
rect 485 -2277 486 -2221
rect 688 -2277 689 -2221
rect 695 -2222 696 -2216
rect 982 -2222 983 -2216
rect 30 -2224 31 -2216
rect 345 -2224 346 -2216
rect 355 -2224 356 -2216
rect 387 -2224 388 -2216
rect 394 -2224 395 -2216
rect 1031 -2224 1032 -2216
rect 44 -2226 45 -2216
rect 383 -2277 384 -2225
rect 387 -2277 388 -2225
rect 422 -2226 423 -2216
rect 436 -2277 437 -2225
rect 681 -2226 682 -2216
rect 695 -2277 696 -2225
rect 737 -2226 738 -2216
rect 768 -2277 769 -2225
rect 800 -2226 801 -2216
rect 856 -2277 857 -2225
rect 1017 -2226 1018 -2216
rect 37 -2228 38 -2216
rect 44 -2277 45 -2227
rect 51 -2228 52 -2216
rect 191 -2277 192 -2227
rect 194 -2228 195 -2216
rect 212 -2228 213 -2216
rect 215 -2277 216 -2227
rect 296 -2228 297 -2216
rect 310 -2228 311 -2216
rect 338 -2277 339 -2227
rect 359 -2228 360 -2216
rect 394 -2277 395 -2227
rect 401 -2228 402 -2216
rect 422 -2277 423 -2227
rect 439 -2228 440 -2216
rect 1010 -2228 1011 -2216
rect 30 -2277 31 -2229
rect 51 -2277 52 -2229
rect 86 -2230 87 -2216
rect 86 -2277 87 -2229
rect 86 -2230 87 -2216
rect 86 -2277 87 -2229
rect 93 -2230 94 -2216
rect 173 -2230 174 -2216
rect 177 -2277 178 -2229
rect 303 -2230 304 -2216
rect 317 -2277 318 -2229
rect 324 -2230 325 -2216
rect 331 -2230 332 -2216
rect 355 -2277 356 -2229
rect 359 -2277 360 -2229
rect 579 -2277 580 -2229
rect 590 -2230 591 -2216
rect 835 -2230 836 -2216
rect 863 -2277 864 -2229
rect 1024 -2230 1025 -2216
rect 23 -2232 24 -2216
rect 303 -2277 304 -2231
rect 331 -2277 332 -2231
rect 499 -2277 500 -2231
rect 502 -2232 503 -2216
rect 520 -2277 521 -2231
rect 548 -2232 549 -2216
rect 569 -2277 570 -2231
rect 572 -2232 573 -2216
rect 702 -2232 703 -2216
rect 723 -2232 724 -2216
rect 814 -2232 815 -2216
rect 835 -2277 836 -2231
rect 961 -2232 962 -2216
rect 23 -2277 24 -2233
rect 163 -2234 164 -2216
rect 166 -2234 167 -2216
rect 544 -2277 545 -2233
rect 576 -2234 577 -2216
rect 639 -2277 640 -2233
rect 653 -2277 654 -2233
rect 709 -2234 710 -2216
rect 723 -2277 724 -2233
rect 772 -2234 773 -2216
rect 779 -2277 780 -2233
rect 793 -2234 794 -2216
rect 800 -2277 801 -2233
rect 912 -2234 913 -2216
rect 922 -2277 923 -2233
rect 996 -2234 997 -2216
rect 37 -2277 38 -2235
rect 142 -2236 143 -2216
rect 156 -2236 157 -2216
rect 184 -2277 185 -2235
rect 201 -2277 202 -2235
rect 565 -2236 566 -2216
rect 590 -2277 591 -2235
rect 632 -2236 633 -2216
rect 667 -2277 668 -2235
rect 730 -2236 731 -2216
rect 737 -2277 738 -2235
rect 786 -2236 787 -2216
rect 793 -2277 794 -2235
rect 940 -2236 941 -2216
rect 961 -2277 962 -2235
rect 1003 -2236 1004 -2216
rect 2 -2238 3 -2216
rect 142 -2277 143 -2237
rect 170 -2277 171 -2237
rect 275 -2238 276 -2216
rect 282 -2277 283 -2237
rect 397 -2238 398 -2216
rect 401 -2277 402 -2237
rect 492 -2238 493 -2216
rect 506 -2277 507 -2237
rect 555 -2238 556 -2216
rect 597 -2277 598 -2237
rect 716 -2238 717 -2216
rect 726 -2238 727 -2216
rect 1045 -2238 1046 -2216
rect 2 -2277 3 -2239
rect 114 -2240 115 -2216
rect 121 -2277 122 -2239
rect 583 -2240 584 -2216
rect 604 -2240 605 -2216
rect 618 -2240 619 -2216
rect 681 -2277 682 -2239
rect 730 -2277 731 -2239
rect 758 -2240 759 -2216
rect 786 -2277 787 -2239
rect 814 -2277 815 -2239
rect 828 -2240 829 -2216
rect 884 -2240 885 -2216
rect 884 -2277 885 -2239
rect 884 -2240 885 -2216
rect 884 -2277 885 -2239
rect 940 -2277 941 -2239
rect 989 -2240 990 -2216
rect 79 -2242 80 -2216
rect 163 -2277 164 -2241
rect 198 -2242 199 -2216
rect 275 -2277 276 -2241
rect 296 -2277 297 -2241
rect 327 -2277 328 -2241
rect 408 -2242 409 -2216
rect 509 -2242 510 -2216
rect 513 -2242 514 -2216
rect 632 -2277 633 -2241
rect 698 -2242 699 -2216
rect 905 -2242 906 -2216
rect 93 -2277 94 -2243
rect 107 -2244 108 -2216
rect 114 -2277 115 -2243
rect 128 -2244 129 -2216
rect 135 -2244 136 -2216
rect 292 -2277 293 -2243
rect 380 -2244 381 -2216
rect 408 -2277 409 -2243
rect 429 -2244 430 -2216
rect 513 -2277 514 -2243
rect 527 -2244 528 -2216
rect 555 -2277 556 -2243
rect 583 -2277 584 -2243
rect 842 -2244 843 -2216
rect 100 -2246 101 -2216
rect 107 -2277 108 -2245
rect 135 -2277 136 -2245
rect 149 -2246 150 -2216
rect 156 -2277 157 -2245
rect 198 -2277 199 -2245
rect 205 -2277 206 -2245
rect 219 -2246 220 -2216
rect 226 -2246 227 -2216
rect 380 -2277 381 -2245
rect 429 -2277 430 -2245
rect 541 -2246 542 -2216
rect 548 -2277 549 -2245
rect 576 -2277 577 -2245
rect 604 -2277 605 -2245
rect 646 -2246 647 -2216
rect 709 -2277 710 -2245
rect 765 -2246 766 -2216
rect 772 -2277 773 -2245
rect 849 -2246 850 -2216
rect 65 -2248 66 -2216
rect 149 -2277 150 -2247
rect 212 -2277 213 -2247
rect 268 -2248 269 -2216
rect 450 -2248 451 -2216
rect 562 -2277 563 -2247
rect 618 -2277 619 -2247
rect 625 -2248 626 -2216
rect 646 -2277 647 -2247
rect 684 -2248 685 -2216
rect 716 -2277 717 -2247
rect 891 -2248 892 -2216
rect 33 -2250 34 -2216
rect 268 -2277 269 -2249
rect 450 -2277 451 -2249
rect 744 -2250 745 -2216
rect 758 -2277 759 -2249
rect 821 -2250 822 -2216
rect 828 -2277 829 -2249
rect 933 -2250 934 -2216
rect 65 -2277 66 -2251
rect 187 -2252 188 -2216
rect 226 -2277 227 -2251
rect 289 -2252 290 -2216
rect 352 -2252 353 -2216
rect 744 -2277 745 -2251
rect 821 -2277 822 -2251
rect 975 -2252 976 -2216
rect 72 -2277 73 -2253
rect 219 -2277 220 -2253
rect 240 -2254 241 -2216
rect 324 -2277 325 -2253
rect 352 -2277 353 -2253
rect 464 -2254 465 -2216
rect 467 -2277 468 -2253
rect 527 -2277 528 -2253
rect 541 -2277 542 -2253
rect 877 -2254 878 -2216
rect 891 -2277 892 -2253
rect 1038 -2254 1039 -2216
rect 240 -2277 241 -2255
rect 415 -2256 416 -2216
rect 457 -2256 458 -2216
rect 481 -2277 482 -2255
rect 593 -2256 594 -2216
rect 625 -2277 626 -2255
rect 684 -2277 685 -2255
rect 702 -2277 703 -2255
rect 842 -2277 843 -2255
rect 919 -2256 920 -2216
rect 968 -2277 969 -2255
rect 975 -2277 976 -2255
rect 58 -2258 59 -2216
rect 415 -2277 416 -2257
rect 443 -2258 444 -2216
rect 457 -2277 458 -2257
rect 471 -2277 472 -2257
rect 611 -2258 612 -2216
rect 849 -2277 850 -2257
rect 898 -2258 899 -2216
rect 912 -2277 913 -2257
rect 933 -2277 934 -2257
rect 16 -2277 17 -2259
rect 58 -2277 59 -2259
rect 247 -2260 248 -2216
rect 247 -2277 248 -2259
rect 247 -2260 248 -2216
rect 247 -2277 248 -2259
rect 254 -2277 255 -2259
rect 369 -2277 370 -2259
rect 443 -2277 444 -2259
rect 674 -2260 675 -2216
rect 877 -2277 878 -2259
rect 926 -2260 927 -2216
rect 261 -2262 262 -2216
rect 310 -2277 311 -2261
rect 478 -2262 479 -2216
rect 674 -2277 675 -2261
rect 233 -2264 234 -2216
rect 261 -2277 262 -2263
rect 478 -2277 479 -2263
rect 492 -2277 493 -2263
rect 534 -2264 535 -2216
rect 898 -2277 899 -2263
rect 233 -2277 234 -2265
rect 523 -2266 524 -2216
rect 611 -2277 612 -2265
rect 660 -2266 661 -2216
rect 502 -2277 503 -2267
rect 534 -2277 535 -2267
rect 660 -2277 661 -2267
rect 751 -2268 752 -2216
rect 751 -2277 752 -2269
rect 807 -2270 808 -2216
rect 807 -2277 808 -2271
rect 947 -2272 948 -2216
rect 947 -2277 948 -2273
rect 954 -2274 955 -2216
rect 464 -2277 465 -2275
rect 954 -2277 955 -2275
rect 2 -2287 3 -2285
rect 51 -2287 52 -2285
rect 58 -2287 59 -2285
rect 275 -2287 276 -2285
rect 303 -2287 304 -2285
rect 478 -2364 479 -2286
rect 481 -2287 482 -2285
rect 891 -2287 892 -2285
rect 905 -2287 906 -2285
rect 933 -2287 934 -2285
rect 2 -2364 3 -2288
rect 30 -2289 31 -2285
rect 44 -2289 45 -2285
rect 54 -2289 55 -2285
rect 58 -2364 59 -2288
rect 436 -2289 437 -2285
rect 450 -2289 451 -2285
rect 467 -2289 468 -2285
rect 499 -2364 500 -2288
rect 611 -2289 612 -2285
rect 618 -2289 619 -2285
rect 618 -2364 619 -2288
rect 618 -2289 619 -2285
rect 618 -2364 619 -2288
rect 639 -2289 640 -2285
rect 639 -2364 640 -2288
rect 639 -2289 640 -2285
rect 639 -2364 640 -2288
rect 642 -2364 643 -2288
rect 800 -2289 801 -2285
rect 877 -2289 878 -2285
rect 891 -2364 892 -2288
rect 908 -2289 909 -2285
rect 947 -2289 948 -2285
rect 9 -2291 10 -2285
rect 128 -2291 129 -2285
rect 191 -2291 192 -2285
rect 212 -2364 213 -2290
rect 226 -2291 227 -2285
rect 345 -2364 346 -2290
rect 376 -2364 377 -2290
rect 646 -2291 647 -2285
rect 684 -2291 685 -2285
rect 835 -2291 836 -2285
rect 877 -2364 878 -2290
rect 954 -2291 955 -2285
rect 12 -2364 13 -2292
rect 215 -2293 216 -2285
rect 268 -2293 269 -2285
rect 488 -2293 489 -2285
rect 502 -2293 503 -2285
rect 723 -2293 724 -2285
rect 765 -2364 766 -2292
rect 828 -2293 829 -2285
rect 884 -2293 885 -2285
rect 912 -2293 913 -2285
rect 922 -2293 923 -2285
rect 929 -2364 930 -2292
rect 947 -2364 948 -2292
rect 961 -2293 962 -2285
rect 16 -2295 17 -2285
rect 485 -2295 486 -2285
rect 506 -2295 507 -2285
rect 506 -2364 507 -2294
rect 506 -2295 507 -2285
rect 506 -2364 507 -2294
rect 534 -2295 535 -2285
rect 565 -2364 566 -2294
rect 569 -2295 570 -2285
rect 569 -2364 570 -2294
rect 569 -2295 570 -2285
rect 569 -2364 570 -2294
rect 576 -2295 577 -2285
rect 856 -2295 857 -2285
rect 926 -2295 927 -2285
rect 975 -2295 976 -2285
rect 16 -2364 17 -2296
rect 233 -2297 234 -2285
rect 268 -2364 269 -2296
rect 296 -2297 297 -2285
rect 303 -2364 304 -2296
rect 415 -2297 416 -2285
rect 436 -2364 437 -2296
rect 457 -2297 458 -2285
rect 464 -2297 465 -2285
rect 562 -2297 563 -2285
rect 583 -2297 584 -2285
rect 660 -2297 661 -2285
rect 723 -2364 724 -2296
rect 821 -2297 822 -2285
rect 842 -2297 843 -2285
rect 884 -2364 885 -2296
rect 23 -2299 24 -2285
rect 51 -2364 52 -2298
rect 61 -2299 62 -2285
rect 705 -2364 706 -2298
rect 768 -2299 769 -2285
rect 849 -2299 850 -2285
rect 856 -2364 857 -2298
rect 898 -2299 899 -2285
rect 23 -2364 24 -2300
rect 282 -2301 283 -2285
rect 296 -2364 297 -2300
rect 464 -2364 465 -2300
rect 467 -2364 468 -2300
rect 471 -2301 472 -2285
rect 520 -2301 521 -2285
rect 576 -2364 577 -2300
rect 597 -2301 598 -2285
rect 646 -2364 647 -2300
rect 779 -2301 780 -2285
rect 828 -2364 829 -2300
rect 849 -2364 850 -2300
rect 901 -2301 902 -2285
rect 30 -2364 31 -2302
rect 229 -2364 230 -2302
rect 233 -2364 234 -2302
rect 261 -2303 262 -2285
rect 275 -2364 276 -2302
rect 362 -2364 363 -2302
rect 373 -2303 374 -2285
rect 485 -2364 486 -2302
rect 562 -2364 563 -2302
rect 758 -2303 759 -2285
rect 786 -2303 787 -2285
rect 821 -2364 822 -2302
rect 44 -2364 45 -2304
rect 779 -2364 780 -2304
rect 793 -2305 794 -2285
rect 842 -2364 843 -2304
rect 47 -2364 48 -2306
rect 131 -2307 132 -2285
rect 163 -2307 164 -2285
rect 191 -2364 192 -2306
rect 261 -2364 262 -2306
rect 289 -2307 290 -2285
rect 310 -2307 311 -2285
rect 334 -2364 335 -2306
rect 341 -2364 342 -2306
rect 716 -2307 717 -2285
rect 793 -2364 794 -2306
rect 863 -2307 864 -2285
rect 65 -2309 66 -2285
rect 310 -2364 311 -2308
rect 313 -2364 314 -2308
rect 786 -2364 787 -2308
rect 800 -2364 801 -2308
rect 814 -2309 815 -2285
rect 65 -2364 66 -2310
rect 100 -2311 101 -2285
rect 107 -2311 108 -2285
rect 625 -2311 626 -2285
rect 667 -2311 668 -2285
rect 814 -2364 815 -2310
rect 72 -2313 73 -2285
rect 177 -2313 178 -2285
rect 282 -2364 283 -2312
rect 408 -2313 409 -2285
rect 415 -2364 416 -2312
rect 716 -2364 717 -2312
rect 72 -2364 73 -2314
rect 79 -2315 80 -2285
rect 82 -2315 83 -2285
rect 86 -2315 87 -2285
rect 93 -2315 94 -2285
rect 103 -2315 104 -2285
rect 107 -2364 108 -2314
rect 110 -2315 111 -2285
rect 114 -2315 115 -2285
rect 198 -2315 199 -2285
rect 289 -2364 290 -2314
rect 338 -2315 339 -2285
rect 355 -2315 356 -2285
rect 471 -2364 472 -2314
rect 537 -2364 538 -2314
rect 758 -2364 759 -2314
rect 79 -2364 80 -2316
rect 149 -2317 150 -2285
rect 163 -2364 164 -2316
rect 338 -2364 339 -2316
rect 355 -2364 356 -2316
rect 660 -2364 661 -2316
rect 681 -2317 682 -2285
rect 863 -2364 864 -2316
rect 86 -2364 87 -2318
rect 541 -2319 542 -2285
rect 586 -2364 587 -2318
rect 667 -2364 668 -2318
rect 93 -2364 94 -2320
rect 523 -2364 524 -2320
rect 597 -2364 598 -2320
rect 604 -2321 605 -2285
rect 611 -2364 612 -2320
rect 632 -2321 633 -2285
rect 100 -2364 101 -2322
rect 422 -2323 423 -2285
rect 450 -2364 451 -2322
rect 730 -2323 731 -2285
rect 114 -2364 115 -2324
rect 135 -2325 136 -2285
rect 149 -2364 150 -2324
rect 184 -2325 185 -2285
rect 198 -2364 199 -2324
rect 205 -2325 206 -2285
rect 317 -2325 318 -2285
rect 397 -2364 398 -2324
rect 401 -2325 402 -2285
rect 541 -2364 542 -2324
rect 625 -2364 626 -2324
rect 688 -2325 689 -2285
rect 54 -2364 55 -2326
rect 135 -2364 136 -2326
rect 142 -2327 143 -2285
rect 184 -2364 185 -2326
rect 205 -2364 206 -2326
rect 348 -2327 349 -2285
rect 359 -2327 360 -2285
rect 730 -2364 731 -2326
rect 128 -2364 129 -2328
rect 240 -2329 241 -2285
rect 317 -2364 318 -2328
rect 674 -2329 675 -2285
rect 688 -2364 689 -2328
rect 695 -2329 696 -2285
rect 142 -2364 143 -2330
rect 156 -2331 157 -2285
rect 177 -2364 178 -2330
rect 247 -2331 248 -2285
rect 324 -2364 325 -2330
rect 443 -2331 444 -2285
rect 513 -2331 514 -2285
rect 632 -2364 633 -2330
rect 674 -2364 675 -2330
rect 709 -2331 710 -2285
rect 37 -2333 38 -2285
rect 156 -2364 157 -2332
rect 180 -2333 181 -2285
rect 695 -2364 696 -2332
rect 702 -2333 703 -2285
rect 709 -2364 710 -2332
rect 37 -2364 38 -2334
rect 110 -2364 111 -2334
rect 121 -2335 122 -2285
rect 247 -2364 248 -2334
rect 254 -2335 255 -2285
rect 513 -2364 514 -2334
rect 702 -2364 703 -2334
rect 751 -2335 752 -2285
rect 121 -2364 122 -2336
rect 292 -2337 293 -2285
rect 359 -2364 360 -2336
rect 394 -2337 395 -2285
rect 401 -2364 402 -2336
rect 653 -2337 654 -2285
rect 737 -2337 738 -2285
rect 751 -2364 752 -2336
rect 240 -2364 241 -2338
rect 527 -2339 528 -2285
rect 737 -2364 738 -2338
rect 744 -2339 745 -2285
rect 254 -2364 255 -2340
rect 579 -2341 580 -2285
rect 744 -2364 745 -2340
rect 772 -2341 773 -2285
rect 352 -2343 353 -2285
rect 527 -2364 528 -2342
rect 772 -2364 773 -2342
rect 870 -2343 871 -2285
rect 366 -2345 367 -2285
rect 604 -2364 605 -2344
rect 870 -2364 871 -2344
rect 940 -2345 941 -2285
rect 170 -2347 171 -2285
rect 366 -2364 367 -2346
rect 380 -2347 381 -2285
rect 681 -2364 682 -2346
rect 159 -2364 160 -2348
rect 170 -2364 171 -2348
rect 331 -2349 332 -2285
rect 380 -2364 381 -2348
rect 383 -2349 384 -2285
rect 408 -2364 409 -2348
rect 422 -2364 423 -2348
rect 429 -2349 430 -2285
rect 443 -2364 444 -2348
rect 548 -2349 549 -2285
rect 373 -2364 374 -2350
rect 429 -2364 430 -2350
rect 492 -2351 493 -2285
rect 653 -2364 654 -2350
rect 387 -2353 388 -2285
rect 387 -2364 388 -2352
rect 387 -2353 388 -2285
rect 387 -2364 388 -2352
rect 394 -2364 395 -2352
rect 835 -2364 836 -2352
rect 492 -2364 493 -2354
rect 555 -2355 556 -2285
rect 548 -2364 549 -2356
rect 590 -2357 591 -2285
rect 544 -2359 545 -2285
rect 590 -2364 591 -2358
rect 555 -2364 556 -2360
rect 807 -2361 808 -2285
rect 583 -2364 584 -2362
rect 807 -2364 808 -2362
rect 16 -2374 17 -2372
rect 138 -2429 139 -2373
rect 142 -2374 143 -2372
rect 142 -2429 143 -2373
rect 142 -2374 143 -2372
rect 142 -2429 143 -2373
rect 156 -2374 157 -2372
rect 215 -2429 216 -2373
rect 226 -2374 227 -2372
rect 667 -2374 668 -2372
rect 702 -2429 703 -2373
rect 709 -2374 710 -2372
rect 726 -2429 727 -2373
rect 821 -2374 822 -2372
rect 884 -2374 885 -2372
rect 884 -2429 885 -2373
rect 884 -2374 885 -2372
rect 884 -2429 885 -2373
rect 891 -2374 892 -2372
rect 891 -2429 892 -2373
rect 891 -2374 892 -2372
rect 891 -2429 892 -2373
rect 926 -2374 927 -2372
rect 926 -2429 927 -2373
rect 926 -2374 927 -2372
rect 926 -2429 927 -2373
rect 940 -2429 941 -2373
rect 947 -2374 948 -2372
rect 23 -2376 24 -2372
rect 219 -2376 220 -2372
rect 240 -2376 241 -2372
rect 558 -2376 559 -2372
rect 569 -2376 570 -2372
rect 667 -2429 668 -2375
rect 709 -2429 710 -2375
rect 765 -2376 766 -2372
rect 772 -2376 773 -2372
rect 828 -2376 829 -2372
rect 30 -2378 31 -2372
rect 156 -2429 157 -2377
rect 177 -2378 178 -2372
rect 226 -2429 227 -2377
rect 233 -2378 234 -2372
rect 240 -2429 241 -2377
rect 247 -2378 248 -2372
rect 352 -2429 353 -2377
rect 376 -2429 377 -2377
rect 758 -2378 759 -2372
rect 761 -2429 762 -2377
rect 842 -2378 843 -2372
rect 2 -2380 3 -2372
rect 30 -2429 31 -2379
rect 44 -2380 45 -2372
rect 61 -2429 62 -2379
rect 72 -2380 73 -2372
rect 72 -2429 73 -2379
rect 72 -2380 73 -2372
rect 72 -2429 73 -2379
rect 86 -2380 87 -2372
rect 86 -2429 87 -2379
rect 86 -2380 87 -2372
rect 86 -2429 87 -2379
rect 93 -2380 94 -2372
rect 208 -2429 209 -2379
rect 212 -2380 213 -2372
rect 373 -2429 374 -2379
rect 404 -2380 405 -2372
rect 779 -2380 780 -2372
rect 828 -2429 829 -2379
rect 877 -2380 878 -2372
rect 37 -2382 38 -2372
rect 93 -2429 94 -2381
rect 100 -2382 101 -2372
rect 359 -2429 360 -2381
rect 411 -2429 412 -2381
rect 436 -2382 437 -2372
rect 457 -2382 458 -2372
rect 576 -2382 577 -2372
rect 583 -2429 584 -2381
rect 660 -2382 661 -2372
rect 723 -2382 724 -2372
rect 765 -2429 766 -2381
rect 772 -2429 773 -2381
rect 793 -2382 794 -2372
rect 51 -2384 52 -2372
rect 730 -2384 731 -2372
rect 751 -2384 752 -2372
rect 754 -2429 755 -2383
rect 100 -2429 101 -2385
rect 149 -2386 150 -2372
rect 177 -2429 178 -2385
rect 254 -2386 255 -2372
rect 261 -2386 262 -2372
rect 261 -2429 262 -2385
rect 261 -2386 262 -2372
rect 261 -2429 262 -2385
rect 268 -2429 269 -2385
rect 289 -2386 290 -2372
rect 303 -2386 304 -2372
rect 418 -2386 419 -2372
rect 460 -2429 461 -2385
rect 506 -2386 507 -2372
rect 520 -2429 521 -2385
rect 548 -2386 549 -2372
rect 555 -2429 556 -2385
rect 625 -2386 626 -2372
rect 639 -2386 640 -2372
rect 688 -2386 689 -2372
rect 723 -2429 724 -2385
rect 849 -2386 850 -2372
rect 107 -2388 108 -2372
rect 450 -2388 451 -2372
rect 464 -2388 465 -2372
rect 506 -2429 507 -2387
rect 523 -2388 524 -2372
rect 611 -2388 612 -2372
rect 618 -2388 619 -2372
rect 628 -2429 629 -2387
rect 639 -2429 640 -2387
rect 835 -2388 836 -2372
rect 107 -2429 108 -2389
rect 149 -2429 150 -2389
rect 163 -2390 164 -2372
rect 289 -2429 290 -2389
rect 310 -2390 311 -2372
rect 604 -2390 605 -2372
rect 611 -2429 612 -2389
rect 674 -2390 675 -2372
rect 114 -2392 115 -2372
rect 152 -2429 153 -2391
rect 163 -2429 164 -2391
rect 184 -2392 185 -2372
rect 205 -2392 206 -2372
rect 247 -2429 248 -2391
rect 275 -2392 276 -2372
rect 397 -2429 398 -2391
rect 408 -2392 409 -2372
rect 436 -2429 437 -2391
rect 450 -2429 451 -2391
rect 471 -2392 472 -2372
rect 481 -2429 482 -2391
rect 716 -2392 717 -2372
rect 114 -2429 115 -2393
rect 170 -2394 171 -2372
rect 184 -2429 185 -2393
rect 222 -2394 223 -2372
rect 233 -2429 234 -2393
rect 387 -2394 388 -2372
rect 408 -2429 409 -2393
rect 646 -2394 647 -2372
rect 660 -2429 661 -2393
rect 737 -2394 738 -2372
rect 121 -2396 122 -2372
rect 271 -2396 272 -2372
rect 275 -2429 276 -2395
rect 422 -2396 423 -2372
rect 464 -2429 465 -2395
rect 814 -2396 815 -2372
rect 65 -2398 66 -2372
rect 121 -2429 122 -2397
rect 135 -2398 136 -2372
rect 303 -2429 304 -2397
rect 310 -2429 311 -2397
rect 355 -2398 356 -2372
rect 380 -2398 381 -2372
rect 604 -2429 605 -2397
rect 618 -2429 619 -2397
rect 695 -2398 696 -2372
rect 716 -2429 717 -2397
rect 807 -2398 808 -2372
rect 170 -2429 171 -2399
rect 191 -2400 192 -2372
rect 219 -2429 220 -2399
rect 548 -2429 549 -2399
rect 551 -2429 552 -2399
rect 646 -2429 647 -2399
rect 674 -2429 675 -2399
rect 786 -2400 787 -2372
rect 807 -2429 808 -2399
rect 863 -2400 864 -2372
rect 191 -2429 192 -2401
rect 198 -2402 199 -2372
rect 282 -2402 283 -2372
rect 457 -2429 458 -2401
rect 471 -2429 472 -2401
rect 562 -2429 563 -2401
rect 737 -2429 738 -2401
rect 744 -2402 745 -2372
rect 128 -2404 129 -2372
rect 282 -2429 283 -2403
rect 313 -2404 314 -2372
rect 541 -2404 542 -2372
rect 744 -2429 745 -2403
rect 856 -2404 857 -2372
rect 128 -2429 129 -2405
rect 296 -2406 297 -2372
rect 324 -2406 325 -2372
rect 341 -2406 342 -2372
rect 345 -2406 346 -2372
rect 422 -2429 423 -2405
rect 527 -2406 528 -2372
rect 569 -2429 570 -2405
rect 79 -2408 80 -2372
rect 296 -2429 297 -2407
rect 317 -2408 318 -2372
rect 345 -2429 346 -2407
rect 527 -2429 528 -2407
rect 590 -2408 591 -2372
rect 58 -2410 59 -2372
rect 79 -2429 80 -2409
rect 198 -2429 199 -2409
rect 222 -2429 223 -2409
rect 317 -2429 318 -2409
rect 544 -2429 545 -2409
rect 58 -2429 59 -2411
rect 65 -2429 66 -2411
rect 324 -2429 325 -2411
rect 415 -2412 416 -2372
rect 534 -2412 535 -2372
rect 597 -2412 598 -2372
rect 331 -2414 332 -2372
rect 380 -2429 381 -2413
rect 415 -2429 416 -2413
rect 429 -2414 430 -2372
rect 499 -2414 500 -2372
rect 534 -2429 535 -2413
rect 597 -2429 598 -2413
rect 681 -2414 682 -2372
rect 331 -2429 332 -2415
rect 366 -2416 367 -2372
rect 429 -2429 430 -2415
rect 590 -2429 591 -2415
rect 653 -2416 654 -2372
rect 681 -2429 682 -2415
rect 334 -2418 335 -2372
rect 387 -2429 388 -2417
rect 401 -2418 402 -2372
rect 653 -2429 654 -2417
rect 254 -2429 255 -2419
rect 334 -2429 335 -2419
rect 338 -2429 339 -2419
rect 513 -2420 514 -2372
rect 366 -2429 367 -2421
rect 485 -2422 486 -2372
rect 499 -2429 500 -2421
rect 632 -2422 633 -2372
rect 401 -2429 402 -2423
rect 492 -2424 493 -2372
rect 513 -2429 514 -2423
rect 565 -2424 566 -2372
rect 443 -2426 444 -2372
rect 492 -2429 493 -2425
rect 394 -2429 395 -2427
rect 443 -2429 444 -2427
rect 488 -2429 489 -2427
rect 632 -2429 633 -2427
rect 65 -2439 66 -2437
rect 72 -2470 73 -2438
rect 79 -2439 80 -2437
rect 264 -2470 265 -2438
rect 268 -2439 269 -2437
rect 408 -2439 409 -2437
rect 422 -2439 423 -2437
rect 464 -2439 465 -2437
rect 471 -2439 472 -2437
rect 583 -2439 584 -2437
rect 590 -2439 591 -2437
rect 593 -2470 594 -2438
rect 625 -2439 626 -2437
rect 716 -2439 717 -2437
rect 730 -2439 731 -2437
rect 737 -2439 738 -2437
rect 754 -2439 755 -2437
rect 807 -2439 808 -2437
rect 884 -2439 885 -2437
rect 884 -2470 885 -2438
rect 884 -2439 885 -2437
rect 884 -2470 885 -2438
rect 891 -2439 892 -2437
rect 891 -2470 892 -2438
rect 891 -2439 892 -2437
rect 891 -2470 892 -2438
rect 926 -2439 927 -2437
rect 933 -2470 934 -2438
rect 940 -2439 941 -2437
rect 940 -2470 941 -2438
rect 940 -2439 941 -2437
rect 940 -2470 941 -2438
rect 93 -2441 94 -2437
rect 131 -2470 132 -2440
rect 135 -2470 136 -2440
rect 142 -2441 143 -2437
rect 170 -2441 171 -2437
rect 215 -2441 216 -2437
rect 233 -2441 234 -2437
rect 369 -2470 370 -2440
rect 401 -2441 402 -2437
rect 471 -2470 472 -2440
rect 474 -2441 475 -2437
rect 481 -2441 482 -2437
rect 485 -2441 486 -2437
rect 604 -2441 605 -2437
rect 625 -2470 626 -2440
rect 660 -2441 661 -2437
rect 681 -2441 682 -2437
rect 688 -2470 689 -2440
rect 695 -2470 696 -2440
rect 702 -2441 703 -2437
rect 716 -2470 717 -2440
rect 726 -2441 727 -2437
rect 730 -2470 731 -2440
rect 733 -2441 734 -2437
rect 765 -2441 766 -2437
rect 765 -2470 766 -2440
rect 765 -2441 766 -2437
rect 765 -2470 766 -2440
rect 779 -2441 780 -2437
rect 828 -2441 829 -2437
rect 100 -2443 101 -2437
rect 156 -2443 157 -2437
rect 191 -2443 192 -2437
rect 208 -2443 209 -2437
rect 240 -2443 241 -2437
rect 257 -2470 258 -2442
rect 275 -2443 276 -2437
rect 331 -2443 332 -2437
rect 334 -2443 335 -2437
rect 390 -2470 391 -2442
rect 408 -2470 409 -2442
rect 415 -2443 416 -2437
rect 422 -2470 423 -2442
rect 478 -2443 479 -2437
rect 502 -2470 503 -2442
rect 569 -2443 570 -2437
rect 576 -2443 577 -2437
rect 653 -2443 654 -2437
rect 660 -2470 661 -2442
rect 667 -2443 668 -2437
rect 681 -2470 682 -2442
rect 709 -2443 710 -2437
rect 100 -2470 101 -2444
rect 117 -2470 118 -2444
rect 121 -2445 122 -2437
rect 219 -2445 220 -2437
rect 226 -2445 227 -2437
rect 275 -2470 276 -2444
rect 296 -2445 297 -2437
rect 597 -2445 598 -2437
rect 604 -2470 605 -2444
rect 611 -2445 612 -2437
rect 642 -2470 643 -2444
rect 646 -2445 647 -2437
rect 709 -2470 710 -2444
rect 744 -2445 745 -2437
rect 107 -2447 108 -2437
rect 121 -2470 122 -2446
rect 128 -2447 129 -2437
rect 219 -2470 220 -2446
rect 226 -2470 227 -2446
rect 261 -2447 262 -2437
rect 303 -2447 304 -2437
rect 303 -2470 304 -2446
rect 303 -2447 304 -2437
rect 303 -2470 304 -2446
rect 310 -2447 311 -2437
rect 488 -2447 489 -2437
rect 506 -2447 507 -2437
rect 600 -2470 601 -2446
rect 611 -2470 612 -2446
rect 632 -2447 633 -2437
rect 114 -2449 115 -2437
rect 233 -2470 234 -2448
rect 254 -2449 255 -2437
rect 268 -2470 269 -2448
rect 317 -2449 318 -2437
rect 432 -2449 433 -2437
rect 443 -2449 444 -2437
rect 478 -2470 479 -2448
rect 499 -2449 500 -2437
rect 506 -2470 507 -2448
rect 513 -2449 514 -2437
rect 579 -2449 580 -2437
rect 107 -2470 108 -2450
rect 114 -2470 115 -2450
rect 149 -2451 150 -2437
rect 170 -2470 171 -2450
rect 191 -2470 192 -2450
rect 198 -2451 199 -2437
rect 222 -2451 223 -2437
rect 310 -2470 311 -2450
rect 345 -2451 346 -2437
rect 401 -2470 402 -2450
rect 443 -2470 444 -2450
rect 450 -2451 451 -2437
rect 457 -2470 458 -2450
rect 492 -2451 493 -2437
rect 513 -2470 514 -2450
rect 534 -2451 535 -2437
rect 541 -2470 542 -2450
rect 562 -2451 563 -2437
rect 569 -2470 570 -2450
rect 618 -2451 619 -2437
rect 86 -2453 87 -2437
rect 450 -2470 451 -2452
rect 460 -2453 461 -2437
rect 520 -2453 521 -2437
rect 527 -2453 528 -2437
rect 551 -2453 552 -2437
rect 555 -2453 556 -2437
rect 576 -2470 577 -2452
rect 152 -2455 153 -2437
rect 198 -2470 199 -2454
rect 282 -2455 283 -2437
rect 317 -2470 318 -2454
rect 331 -2470 332 -2454
rect 345 -2470 346 -2454
rect 348 -2470 349 -2454
rect 387 -2455 388 -2437
rect 534 -2470 535 -2454
rect 674 -2455 675 -2437
rect 163 -2457 164 -2437
rect 240 -2470 241 -2456
rect 289 -2457 290 -2437
rect 432 -2470 433 -2456
rect 548 -2470 549 -2456
rect 639 -2457 640 -2437
rect 674 -2470 675 -2456
rect 758 -2457 759 -2437
rect 163 -2470 164 -2458
rect 184 -2459 185 -2437
rect 212 -2459 213 -2437
rect 282 -2470 283 -2458
rect 352 -2459 353 -2437
rect 394 -2459 395 -2437
rect 639 -2470 640 -2458
rect 723 -2459 724 -2437
rect 737 -2470 738 -2458
rect 758 -2470 759 -2458
rect 184 -2470 185 -2460
rect 205 -2470 206 -2460
rect 247 -2461 248 -2437
rect 289 -2470 290 -2460
rect 324 -2461 325 -2437
rect 352 -2470 353 -2460
rect 359 -2461 360 -2437
rect 467 -2461 468 -2437
rect 723 -2470 724 -2460
rect 761 -2461 762 -2437
rect 177 -2463 178 -2437
rect 247 -2470 248 -2462
rect 338 -2463 339 -2437
rect 359 -2470 360 -2462
rect 366 -2463 367 -2437
rect 415 -2470 416 -2462
rect 761 -2470 762 -2462
rect 772 -2463 773 -2437
rect 159 -2465 160 -2437
rect 177 -2470 178 -2464
rect 299 -2470 300 -2464
rect 338 -2470 339 -2464
rect 387 -2470 388 -2464
rect 436 -2465 437 -2437
rect 380 -2467 381 -2437
rect 436 -2470 437 -2466
rect 373 -2470 374 -2468
rect 380 -2470 381 -2468
rect 394 -2470 395 -2468
rect 397 -2469 398 -2437
rect 5 -2480 6 -2478
rect 5 -2497 6 -2479
rect 5 -2480 6 -2478
rect 5 -2497 6 -2479
rect 65 -2480 66 -2478
rect 72 -2480 73 -2478
rect 86 -2497 87 -2479
rect 96 -2497 97 -2479
rect 100 -2480 101 -2478
rect 110 -2497 111 -2479
rect 114 -2480 115 -2478
rect 121 -2480 122 -2478
rect 131 -2480 132 -2478
rect 135 -2480 136 -2478
rect 142 -2497 143 -2479
rect 170 -2480 171 -2478
rect 177 -2480 178 -2478
rect 187 -2480 188 -2478
rect 198 -2480 199 -2478
rect 212 -2497 213 -2479
rect 219 -2480 220 -2478
rect 254 -2497 255 -2479
rect 282 -2480 283 -2478
rect 362 -2497 363 -2479
rect 376 -2480 377 -2478
rect 422 -2480 423 -2478
rect 432 -2480 433 -2478
rect 457 -2480 458 -2478
rect 467 -2480 468 -2478
rect 478 -2480 479 -2478
rect 502 -2480 503 -2478
rect 513 -2480 514 -2478
rect 523 -2480 524 -2478
rect 541 -2480 542 -2478
rect 576 -2480 577 -2478
rect 586 -2480 587 -2478
rect 590 -2480 591 -2478
rect 625 -2480 626 -2478
rect 660 -2480 661 -2478
rect 660 -2497 661 -2479
rect 660 -2480 661 -2478
rect 660 -2497 661 -2479
rect 667 -2497 668 -2479
rect 681 -2480 682 -2478
rect 730 -2480 731 -2478
rect 730 -2497 731 -2479
rect 730 -2480 731 -2478
rect 730 -2497 731 -2479
rect 744 -2497 745 -2479
rect 751 -2497 752 -2479
rect 758 -2480 759 -2478
rect 765 -2480 766 -2478
rect 884 -2480 885 -2478
rect 884 -2497 885 -2479
rect 884 -2480 885 -2478
rect 884 -2497 885 -2479
rect 891 -2480 892 -2478
rect 891 -2497 892 -2479
rect 891 -2480 892 -2478
rect 891 -2497 892 -2479
rect 933 -2497 934 -2479
rect 936 -2480 937 -2478
rect 940 -2480 941 -2478
rect 947 -2497 948 -2479
rect 100 -2497 101 -2481
rect 121 -2497 122 -2481
rect 138 -2497 139 -2481
rect 219 -2497 220 -2481
rect 226 -2482 227 -2478
rect 229 -2488 230 -2481
rect 247 -2482 248 -2478
rect 324 -2482 325 -2478
rect 338 -2482 339 -2478
rect 404 -2497 405 -2481
rect 450 -2482 451 -2478
rect 548 -2482 549 -2478
rect 597 -2482 598 -2478
rect 674 -2482 675 -2478
rect 681 -2497 682 -2481
rect 688 -2482 689 -2478
rect 758 -2497 759 -2481
rect 761 -2482 762 -2478
rect 107 -2484 108 -2478
rect 114 -2497 115 -2483
rect 149 -2497 150 -2483
rect 163 -2484 164 -2478
rect 177 -2497 178 -2483
rect 191 -2484 192 -2478
rect 205 -2484 206 -2478
rect 205 -2497 206 -2483
rect 205 -2484 206 -2478
rect 205 -2497 206 -2483
rect 226 -2497 227 -2483
rect 261 -2484 262 -2478
rect 275 -2484 276 -2478
rect 324 -2497 325 -2483
rect 352 -2484 353 -2478
rect 352 -2497 353 -2483
rect 352 -2484 353 -2478
rect 352 -2497 353 -2483
rect 359 -2484 360 -2478
rect 373 -2484 374 -2478
rect 380 -2484 381 -2478
rect 380 -2497 381 -2483
rect 380 -2484 381 -2478
rect 380 -2497 381 -2483
rect 394 -2484 395 -2478
rect 394 -2497 395 -2483
rect 394 -2484 395 -2478
rect 394 -2497 395 -2483
rect 401 -2484 402 -2478
rect 422 -2497 423 -2483
rect 443 -2484 444 -2478
rect 450 -2497 451 -2483
rect 471 -2484 472 -2478
rect 527 -2484 528 -2478
rect 604 -2484 605 -2478
rect 604 -2497 605 -2483
rect 604 -2484 605 -2478
rect 604 -2497 605 -2483
rect 611 -2484 612 -2478
rect 611 -2497 612 -2483
rect 611 -2484 612 -2478
rect 611 -2497 612 -2483
rect 688 -2497 689 -2483
rect 695 -2484 696 -2478
rect 159 -2497 160 -2485
rect 170 -2497 171 -2485
rect 233 -2486 234 -2478
rect 261 -2497 262 -2485
rect 271 -2497 272 -2485
rect 275 -2497 276 -2485
rect 296 -2486 297 -2478
rect 303 -2486 304 -2478
rect 310 -2486 311 -2478
rect 366 -2486 367 -2478
rect 401 -2497 402 -2485
rect 537 -2486 538 -2478
rect 695 -2497 696 -2485
rect 709 -2486 710 -2478
rect 233 -2497 234 -2487
rect 236 -2488 237 -2478
rect 310 -2497 311 -2487
rect 359 -2497 360 -2487
rect 408 -2488 409 -2478
rect 415 -2488 416 -2478
rect 443 -2497 444 -2487
rect 506 -2488 507 -2478
rect 520 -2488 521 -2478
rect 523 -2497 524 -2487
rect 527 -2497 528 -2487
rect 709 -2497 710 -2487
rect 716 -2488 717 -2478
rect 240 -2497 241 -2489
rect 296 -2497 297 -2489
rect 303 -2497 304 -2489
rect 331 -2490 332 -2478
rect 408 -2497 409 -2489
rect 436 -2490 437 -2478
rect 520 -2497 521 -2489
rect 569 -2490 570 -2478
rect 716 -2497 717 -2489
rect 723 -2490 724 -2478
rect 247 -2497 248 -2491
rect 268 -2492 269 -2478
rect 317 -2492 318 -2478
rect 331 -2497 332 -2491
rect 723 -2497 724 -2491
rect 737 -2492 738 -2478
rect 289 -2494 290 -2478
rect 317 -2497 318 -2493
rect 201 -2497 202 -2495
rect 289 -2497 290 -2495
rect 5 -2507 6 -2505
rect 9 -2516 10 -2506
rect 86 -2507 87 -2505
rect 103 -2507 104 -2505
rect 107 -2507 108 -2505
rect 121 -2507 122 -2505
rect 142 -2507 143 -2505
rect 194 -2507 195 -2505
rect 201 -2507 202 -2505
rect 205 -2507 206 -2505
rect 219 -2507 220 -2505
rect 240 -2507 241 -2505
rect 247 -2507 248 -2505
rect 271 -2516 272 -2506
rect 275 -2507 276 -2505
rect 282 -2507 283 -2505
rect 285 -2516 286 -2506
rect 317 -2507 318 -2505
rect 331 -2507 332 -2505
rect 345 -2516 346 -2506
rect 352 -2507 353 -2505
rect 362 -2516 363 -2506
rect 380 -2507 381 -2505
rect 383 -2516 384 -2506
rect 387 -2507 388 -2505
rect 408 -2507 409 -2505
rect 450 -2507 451 -2505
rect 457 -2516 458 -2506
rect 523 -2516 524 -2506
rect 527 -2507 528 -2505
rect 597 -2516 598 -2506
rect 604 -2507 605 -2505
rect 660 -2507 661 -2505
rect 663 -2516 664 -2506
rect 667 -2507 668 -2505
rect 667 -2516 668 -2506
rect 667 -2507 668 -2505
rect 667 -2516 668 -2506
rect 681 -2507 682 -2505
rect 702 -2507 703 -2505
rect 709 -2507 710 -2505
rect 712 -2516 713 -2506
rect 716 -2507 717 -2505
rect 716 -2516 717 -2506
rect 716 -2507 717 -2505
rect 716 -2516 717 -2506
rect 723 -2507 724 -2505
rect 730 -2516 731 -2506
rect 740 -2507 741 -2505
rect 751 -2507 752 -2505
rect 887 -2507 888 -2505
rect 891 -2507 892 -2505
rect 933 -2507 934 -2505
rect 940 -2507 941 -2505
rect 943 -2507 944 -2505
rect 947 -2507 948 -2505
rect 100 -2509 101 -2505
rect 107 -2516 108 -2508
rect 114 -2516 115 -2508
rect 117 -2509 118 -2505
rect 149 -2509 150 -2505
rect 166 -2509 167 -2505
rect 184 -2516 185 -2508
rect 187 -2509 188 -2505
rect 191 -2509 192 -2505
rect 226 -2509 227 -2505
rect 229 -2516 230 -2508
rect 233 -2509 234 -2505
rect 254 -2509 255 -2505
rect 278 -2516 279 -2508
rect 289 -2509 290 -2505
rect 303 -2509 304 -2505
rect 394 -2509 395 -2505
rect 397 -2516 398 -2508
rect 404 -2509 405 -2505
rect 418 -2509 419 -2505
rect 443 -2509 444 -2505
rect 450 -2516 451 -2508
rect 604 -2516 605 -2508
rect 611 -2509 612 -2505
rect 688 -2509 689 -2505
rect 688 -2516 689 -2508
rect 688 -2509 689 -2505
rect 688 -2516 689 -2508
rect 695 -2509 696 -2505
rect 705 -2509 706 -2505
rect 744 -2509 745 -2505
rect 758 -2509 759 -2505
rect 156 -2511 157 -2505
rect 159 -2516 160 -2510
rect 163 -2511 164 -2505
rect 170 -2511 171 -2505
rect 177 -2511 178 -2505
rect 191 -2516 192 -2510
rect 212 -2511 213 -2505
rect 226 -2516 227 -2510
rect 261 -2511 262 -2505
rect 268 -2511 269 -2505
rect 296 -2516 297 -2510
rect 310 -2511 311 -2505
rect 401 -2511 402 -2505
rect 404 -2516 405 -2510
rect 163 -2516 164 -2512
rect 180 -2516 181 -2512
rect 299 -2513 300 -2505
rect 341 -2516 342 -2512
rect 310 -2516 311 -2514
rect 324 -2515 325 -2505
rect 5 -2526 6 -2524
rect 9 -2526 10 -2524
rect 100 -2526 101 -2524
rect 107 -2526 108 -2524
rect 114 -2526 115 -2524
rect 124 -2526 125 -2524
rect 163 -2526 164 -2524
rect 170 -2526 171 -2524
rect 180 -2526 181 -2524
rect 184 -2526 185 -2524
rect 191 -2526 192 -2524
rect 198 -2526 199 -2524
rect 292 -2526 293 -2524
rect 296 -2526 297 -2524
rect 303 -2526 304 -2524
rect 310 -2526 311 -2524
rect 341 -2526 342 -2524
rect 345 -2526 346 -2524
rect 450 -2526 451 -2524
rect 457 -2526 458 -2524
rect 597 -2526 598 -2524
rect 604 -2526 605 -2524
rect 663 -2526 664 -2524
rect 667 -2526 668 -2524
rect 716 -2526 717 -2524
rect 723 -2526 724 -2524
rect 730 -2526 731 -2524
rect 740 -2526 741 -2524
rect 121 -2528 122 -2524
rect 131 -2528 132 -2524
<< labels >>
rlabel pdiffusion 3 -8 3 -8 0 cellNo=39
rlabel pdiffusion 10 -8 10 -8 0 cellNo=557
rlabel pdiffusion 17 -8 17 -8 0 cellNo=73
rlabel pdiffusion 24 -8 24 -8 0 cellNo=710
rlabel pdiffusion 31 -8 31 -8 0 cellNo=178
rlabel pdiffusion 38 -8 38 -8 0 cellNo=970
rlabel pdiffusion 87 -8 87 -8 0 cellNo=1000
rlabel pdiffusion 94 -8 94 -8 0 feedthrough
rlabel pdiffusion 101 -8 101 -8 0 cellNo=731
rlabel pdiffusion 108 -8 108 -8 0 cellNo=816
rlabel pdiffusion 115 -8 115 -8 0 cellNo=369
rlabel pdiffusion 122 -8 122 -8 0 feedthrough
rlabel pdiffusion 129 -8 129 -8 0 feedthrough
rlabel pdiffusion 143 -8 143 -8 0 cellNo=518
rlabel pdiffusion 206 -8 206 -8 0 feedthrough
rlabel pdiffusion 213 -8 213 -8 0 cellNo=590
rlabel pdiffusion 220 -8 220 -8 0 cellNo=988
rlabel pdiffusion 227 -8 227 -8 0 feedthrough
rlabel pdiffusion 234 -8 234 -8 0 cellNo=313
rlabel pdiffusion 241 -8 241 -8 0 feedthrough
rlabel pdiffusion 248 -8 248 -8 0 cellNo=53
rlabel pdiffusion 255 -8 255 -8 0 cellNo=110
rlabel pdiffusion 262 -8 262 -8 0 cellNo=189
rlabel pdiffusion 269 -8 269 -8 0 feedthrough
rlabel pdiffusion 283 -8 283 -8 0 cellNo=691
rlabel pdiffusion 325 -8 325 -8 0 feedthrough
rlabel pdiffusion 332 -8 332 -8 0 cellNo=277
rlabel pdiffusion 339 -8 339 -8 0 cellNo=406
rlabel pdiffusion 430 -8 430 -8 0 feedthrough
rlabel pdiffusion 451 -8 451 -8 0 cellNo=390
rlabel pdiffusion 465 -8 465 -8 0 feedthrough
rlabel pdiffusion 486 -8 486 -8 0 cellNo=907
rlabel pdiffusion 507 -8 507 -8 0 cellNo=449
rlabel pdiffusion 528 -8 528 -8 0 cellNo=612
rlabel pdiffusion 535 -8 535 -8 0 feedthrough
rlabel pdiffusion 549 -8 549 -8 0 cellNo=662
rlabel pdiffusion 584 -8 584 -8 0 cellNo=430
rlabel pdiffusion 591 -8 591 -8 0 cellNo=695
rlabel pdiffusion 598 -8 598 -8 0 feedthrough
rlabel pdiffusion 605 -8 605 -8 0 cellNo=375
rlabel pdiffusion 661 -8 661 -8 0 cellNo=788
rlabel pdiffusion 668 -8 668 -8 0 feedthrough
rlabel pdiffusion 3 -27 3 -27 0 cellNo=129
rlabel pdiffusion 10 -27 10 -27 0 cellNo=159
rlabel pdiffusion 17 -27 17 -27 0 cellNo=316
rlabel pdiffusion 24 -27 24 -27 0 cellNo=175
rlabel pdiffusion 31 -27 31 -27 0 cellNo=302
rlabel pdiffusion 101 -27 101 -27 0 cellNo=549
rlabel pdiffusion 115 -27 115 -27 0 cellNo=100
rlabel pdiffusion 136 -27 136 -27 0 feedthrough
rlabel pdiffusion 171 -27 171 -27 0 cellNo=876
rlabel pdiffusion 178 -27 178 -27 0 feedthrough
rlabel pdiffusion 185 -27 185 -27 0 feedthrough
rlabel pdiffusion 192 -27 192 -27 0 cellNo=273
rlabel pdiffusion 199 -27 199 -27 0 feedthrough
rlabel pdiffusion 206 -27 206 -27 0 cellNo=31
rlabel pdiffusion 213 -27 213 -27 0 cellNo=637
rlabel pdiffusion 220 -27 220 -27 0 feedthrough
rlabel pdiffusion 227 -27 227 -27 0 feedthrough
rlabel pdiffusion 234 -27 234 -27 0 cellNo=832
rlabel pdiffusion 241 -27 241 -27 0 cellNo=344
rlabel pdiffusion 248 -27 248 -27 0 feedthrough
rlabel pdiffusion 255 -27 255 -27 0 feedthrough
rlabel pdiffusion 262 -27 262 -27 0 feedthrough
rlabel pdiffusion 269 -27 269 -27 0 feedthrough
rlabel pdiffusion 276 -27 276 -27 0 feedthrough
rlabel pdiffusion 283 -27 283 -27 0 feedthrough
rlabel pdiffusion 290 -27 290 -27 0 feedthrough
rlabel pdiffusion 297 -27 297 -27 0 cellNo=609
rlabel pdiffusion 304 -27 304 -27 0 cellNo=761
rlabel pdiffusion 311 -27 311 -27 0 feedthrough
rlabel pdiffusion 318 -27 318 -27 0 feedthrough
rlabel pdiffusion 325 -27 325 -27 0 feedthrough
rlabel pdiffusion 332 -27 332 -27 0 cellNo=397
rlabel pdiffusion 339 -27 339 -27 0 cellNo=328
rlabel pdiffusion 346 -27 346 -27 0 cellNo=845
rlabel pdiffusion 360 -27 360 -27 0 feedthrough
rlabel pdiffusion 374 -27 374 -27 0 feedthrough
rlabel pdiffusion 381 -27 381 -27 0 cellNo=982
rlabel pdiffusion 416 -27 416 -27 0 feedthrough
rlabel pdiffusion 423 -27 423 -27 0 cellNo=725
rlabel pdiffusion 430 -27 430 -27 0 feedthrough
rlabel pdiffusion 437 -27 437 -27 0 cellNo=782
rlabel pdiffusion 444 -27 444 -27 0 cellNo=969
rlabel pdiffusion 451 -27 451 -27 0 cellNo=329
rlabel pdiffusion 465 -27 465 -27 0 cellNo=868
rlabel pdiffusion 472 -27 472 -27 0 feedthrough
rlabel pdiffusion 493 -27 493 -27 0 feedthrough
rlabel pdiffusion 507 -27 507 -27 0 feedthrough
rlabel pdiffusion 514 -27 514 -27 0 cellNo=567
rlabel pdiffusion 521 -27 521 -27 0 cellNo=528
rlabel pdiffusion 528 -27 528 -27 0 feedthrough
rlabel pdiffusion 542 -27 542 -27 0 feedthrough
rlabel pdiffusion 556 -27 556 -27 0 cellNo=86
rlabel pdiffusion 563 -27 563 -27 0 cellNo=994
rlabel pdiffusion 570 -27 570 -27 0 feedthrough
rlabel pdiffusion 577 -27 577 -27 0 feedthrough
rlabel pdiffusion 605 -27 605 -27 0 feedthrough
rlabel pdiffusion 612 -27 612 -27 0 feedthrough
rlabel pdiffusion 619 -27 619 -27 0 feedthrough
rlabel pdiffusion 675 -27 675 -27 0 feedthrough
rlabel pdiffusion 3 -58 3 -58 0 cellNo=121
rlabel pdiffusion 10 -58 10 -58 0 cellNo=680
rlabel pdiffusion 17 -58 17 -58 0 cellNo=171
rlabel pdiffusion 24 -58 24 -58 0 cellNo=295
rlabel pdiffusion 87 -58 87 -58 0 feedthrough
rlabel pdiffusion 94 -58 94 -58 0 feedthrough
rlabel pdiffusion 115 -58 115 -58 0 feedthrough
rlabel pdiffusion 122 -58 122 -58 0 feedthrough
rlabel pdiffusion 129 -58 129 -58 0 feedthrough
rlabel pdiffusion 136 -58 136 -58 0 feedthrough
rlabel pdiffusion 143 -58 143 -58 0 cellNo=949
rlabel pdiffusion 150 -58 150 -58 0 cellNo=435
rlabel pdiffusion 157 -58 157 -58 0 feedthrough
rlabel pdiffusion 164 -58 164 -58 0 feedthrough
rlabel pdiffusion 171 -58 171 -58 0 cellNo=486
rlabel pdiffusion 178 -58 178 -58 0 cellNo=573
rlabel pdiffusion 185 -58 185 -58 0 cellNo=824
rlabel pdiffusion 192 -58 192 -58 0 feedthrough
rlabel pdiffusion 199 -58 199 -58 0 cellNo=880
rlabel pdiffusion 206 -58 206 -58 0 feedthrough
rlabel pdiffusion 213 -58 213 -58 0 feedthrough
rlabel pdiffusion 220 -58 220 -58 0 feedthrough
rlabel pdiffusion 227 -58 227 -58 0 feedthrough
rlabel pdiffusion 234 -58 234 -58 0 cellNo=732
rlabel pdiffusion 241 -58 241 -58 0 cellNo=106
rlabel pdiffusion 248 -58 248 -58 0 cellNo=339
rlabel pdiffusion 255 -58 255 -58 0 feedthrough
rlabel pdiffusion 262 -58 262 -58 0 feedthrough
rlabel pdiffusion 269 -58 269 -58 0 feedthrough
rlabel pdiffusion 276 -58 276 -58 0 cellNo=179
rlabel pdiffusion 283 -58 283 -58 0 feedthrough
rlabel pdiffusion 290 -58 290 -58 0 feedthrough
rlabel pdiffusion 297 -58 297 -58 0 cellNo=542
rlabel pdiffusion 304 -58 304 -58 0 feedthrough
rlabel pdiffusion 311 -58 311 -58 0 cellNo=162
rlabel pdiffusion 318 -58 318 -58 0 feedthrough
rlabel pdiffusion 325 -58 325 -58 0 feedthrough
rlabel pdiffusion 332 -58 332 -58 0 feedthrough
rlabel pdiffusion 339 -58 339 -58 0 cellNo=158
rlabel pdiffusion 346 -58 346 -58 0 feedthrough
rlabel pdiffusion 353 -58 353 -58 0 feedthrough
rlabel pdiffusion 360 -58 360 -58 0 cellNo=251
rlabel pdiffusion 367 -58 367 -58 0 feedthrough
rlabel pdiffusion 374 -58 374 -58 0 cellNo=623
rlabel pdiffusion 381 -58 381 -58 0 cellNo=27
rlabel pdiffusion 388 -58 388 -58 0 feedthrough
rlabel pdiffusion 395 -58 395 -58 0 feedthrough
rlabel pdiffusion 402 -58 402 -58 0 feedthrough
rlabel pdiffusion 409 -58 409 -58 0 feedthrough
rlabel pdiffusion 416 -58 416 -58 0 cellNo=50
rlabel pdiffusion 423 -58 423 -58 0 feedthrough
rlabel pdiffusion 430 -58 430 -58 0 feedthrough
rlabel pdiffusion 437 -58 437 -58 0 feedthrough
rlabel pdiffusion 444 -58 444 -58 0 feedthrough
rlabel pdiffusion 465 -58 465 -58 0 cellNo=878
rlabel pdiffusion 472 -58 472 -58 0 feedthrough
rlabel pdiffusion 479 -58 479 -58 0 feedthrough
rlabel pdiffusion 486 -58 486 -58 0 feedthrough
rlabel pdiffusion 493 -58 493 -58 0 cellNo=44
rlabel pdiffusion 500 -58 500 -58 0 feedthrough
rlabel pdiffusion 507 -58 507 -58 0 feedthrough
rlabel pdiffusion 521 -58 521 -58 0 feedthrough
rlabel pdiffusion 528 -58 528 -58 0 cellNo=392
rlabel pdiffusion 535 -58 535 -58 0 feedthrough
rlabel pdiffusion 542 -58 542 -58 0 feedthrough
rlabel pdiffusion 549 -58 549 -58 0 cellNo=320
rlabel pdiffusion 556 -58 556 -58 0 cellNo=318
rlabel pdiffusion 563 -58 563 -58 0 feedthrough
rlabel pdiffusion 570 -58 570 -58 0 feedthrough
rlabel pdiffusion 577 -58 577 -58 0 feedthrough
rlabel pdiffusion 584 -58 584 -58 0 cellNo=770
rlabel pdiffusion 591 -58 591 -58 0 feedthrough
rlabel pdiffusion 598 -58 598 -58 0 feedthrough
rlabel pdiffusion 605 -58 605 -58 0 feedthrough
rlabel pdiffusion 612 -58 612 -58 0 feedthrough
rlabel pdiffusion 626 -58 626 -58 0 feedthrough
rlabel pdiffusion 633 -58 633 -58 0 feedthrough
rlabel pdiffusion 640 -58 640 -58 0 feedthrough
rlabel pdiffusion 647 -58 647 -58 0 feedthrough
rlabel pdiffusion 654 -58 654 -58 0 feedthrough
rlabel pdiffusion 661 -58 661 -58 0 cellNo=900
rlabel pdiffusion 668 -58 668 -58 0 feedthrough
rlabel pdiffusion 675 -58 675 -58 0 cellNo=42
rlabel pdiffusion 682 -58 682 -58 0 feedthrough
rlabel pdiffusion 703 -58 703 -58 0 feedthrough
rlabel pdiffusion 766 -58 766 -58 0 cellNo=234
rlabel pdiffusion 773 -58 773 -58 0 feedthrough
rlabel pdiffusion 843 -58 843 -58 0 feedthrough
rlabel pdiffusion 3 -127 3 -127 0 cellNo=92
rlabel pdiffusion 10 -127 10 -127 0 cellNo=148
rlabel pdiffusion 17 -127 17 -127 0 cellNo=225
rlabel pdiffusion 24 -127 24 -127 0 cellNo=899
rlabel pdiffusion 31 -127 31 -127 0 feedthrough
rlabel pdiffusion 38 -127 38 -127 0 feedthrough
rlabel pdiffusion 45 -127 45 -127 0 cellNo=540
rlabel pdiffusion 52 -127 52 -127 0 cellNo=942
rlabel pdiffusion 59 -127 59 -127 0 cellNo=463
rlabel pdiffusion 66 -127 66 -127 0 feedthrough
rlabel pdiffusion 73 -127 73 -127 0 feedthrough
rlabel pdiffusion 80 -127 80 -127 0 cellNo=335
rlabel pdiffusion 87 -127 87 -127 0 feedthrough
rlabel pdiffusion 94 -127 94 -127 0 feedthrough
rlabel pdiffusion 101 -127 101 -127 0 cellNo=850
rlabel pdiffusion 108 -127 108 -127 0 feedthrough
rlabel pdiffusion 115 -127 115 -127 0 cellNo=774
rlabel pdiffusion 122 -127 122 -127 0 feedthrough
rlabel pdiffusion 129 -127 129 -127 0 cellNo=651
rlabel pdiffusion 136 -127 136 -127 0 cellNo=357
rlabel pdiffusion 143 -127 143 -127 0 feedthrough
rlabel pdiffusion 150 -127 150 -127 0 cellNo=510
rlabel pdiffusion 157 -127 157 -127 0 cellNo=746
rlabel pdiffusion 164 -127 164 -127 0 feedthrough
rlabel pdiffusion 171 -127 171 -127 0 cellNo=686
rlabel pdiffusion 178 -127 178 -127 0 feedthrough
rlabel pdiffusion 185 -127 185 -127 0 feedthrough
rlabel pdiffusion 192 -127 192 -127 0 feedthrough
rlabel pdiffusion 199 -127 199 -127 0 feedthrough
rlabel pdiffusion 206 -127 206 -127 0 feedthrough
rlabel pdiffusion 213 -127 213 -127 0 feedthrough
rlabel pdiffusion 220 -127 220 -127 0 feedthrough
rlabel pdiffusion 227 -127 227 -127 0 cellNo=213
rlabel pdiffusion 234 -127 234 -127 0 feedthrough
rlabel pdiffusion 241 -127 241 -127 0 feedthrough
rlabel pdiffusion 248 -127 248 -127 0 cellNo=212
rlabel pdiffusion 255 -127 255 -127 0 feedthrough
rlabel pdiffusion 262 -127 262 -127 0 feedthrough
rlabel pdiffusion 269 -127 269 -127 0 feedthrough
rlabel pdiffusion 276 -127 276 -127 0 cellNo=400
rlabel pdiffusion 283 -127 283 -127 0 feedthrough
rlabel pdiffusion 290 -127 290 -127 0 feedthrough
rlabel pdiffusion 297 -127 297 -127 0 feedthrough
rlabel pdiffusion 304 -127 304 -127 0 feedthrough
rlabel pdiffusion 311 -127 311 -127 0 feedthrough
rlabel pdiffusion 318 -127 318 -127 0 cellNo=786
rlabel pdiffusion 325 -127 325 -127 0 feedthrough
rlabel pdiffusion 332 -127 332 -127 0 feedthrough
rlabel pdiffusion 339 -127 339 -127 0 feedthrough
rlabel pdiffusion 346 -127 346 -127 0 cellNo=652
rlabel pdiffusion 353 -127 353 -127 0 cellNo=977
rlabel pdiffusion 360 -127 360 -127 0 feedthrough
rlabel pdiffusion 367 -127 367 -127 0 feedthrough
rlabel pdiffusion 374 -127 374 -127 0 cellNo=182
rlabel pdiffusion 381 -127 381 -127 0 feedthrough
rlabel pdiffusion 388 -127 388 -127 0 cellNo=967
rlabel pdiffusion 395 -127 395 -127 0 cellNo=513
rlabel pdiffusion 402 -127 402 -127 0 feedthrough
rlabel pdiffusion 409 -127 409 -127 0 feedthrough
rlabel pdiffusion 416 -127 416 -127 0 cellNo=618
rlabel pdiffusion 423 -127 423 -127 0 feedthrough
rlabel pdiffusion 430 -127 430 -127 0 feedthrough
rlabel pdiffusion 437 -127 437 -127 0 feedthrough
rlabel pdiffusion 444 -127 444 -127 0 feedthrough
rlabel pdiffusion 451 -127 451 -127 0 feedthrough
rlabel pdiffusion 458 -127 458 -127 0 feedthrough
rlabel pdiffusion 465 -127 465 -127 0 feedthrough
rlabel pdiffusion 472 -127 472 -127 0 feedthrough
rlabel pdiffusion 479 -127 479 -127 0 feedthrough
rlabel pdiffusion 486 -127 486 -127 0 feedthrough
rlabel pdiffusion 493 -127 493 -127 0 feedthrough
rlabel pdiffusion 500 -127 500 -127 0 cellNo=511
rlabel pdiffusion 507 -127 507 -127 0 cellNo=592
rlabel pdiffusion 514 -127 514 -127 0 feedthrough
rlabel pdiffusion 521 -127 521 -127 0 feedthrough
rlabel pdiffusion 528 -127 528 -127 0 feedthrough
rlabel pdiffusion 535 -127 535 -127 0 feedthrough
rlabel pdiffusion 542 -127 542 -127 0 feedthrough
rlabel pdiffusion 549 -127 549 -127 0 feedthrough
rlabel pdiffusion 556 -127 556 -127 0 feedthrough
rlabel pdiffusion 563 -127 563 -127 0 feedthrough
rlabel pdiffusion 570 -127 570 -127 0 feedthrough
rlabel pdiffusion 577 -127 577 -127 0 feedthrough
rlabel pdiffusion 584 -127 584 -127 0 cellNo=735
rlabel pdiffusion 591 -127 591 -127 0 feedthrough
rlabel pdiffusion 598 -127 598 -127 0 feedthrough
rlabel pdiffusion 605 -127 605 -127 0 feedthrough
rlabel pdiffusion 612 -127 612 -127 0 feedthrough
rlabel pdiffusion 619 -127 619 -127 0 feedthrough
rlabel pdiffusion 626 -127 626 -127 0 feedthrough
rlabel pdiffusion 633 -127 633 -127 0 feedthrough
rlabel pdiffusion 640 -127 640 -127 0 feedthrough
rlabel pdiffusion 647 -127 647 -127 0 feedthrough
rlabel pdiffusion 654 -127 654 -127 0 feedthrough
rlabel pdiffusion 661 -127 661 -127 0 cellNo=160
rlabel pdiffusion 668 -127 668 -127 0 feedthrough
rlabel pdiffusion 675 -127 675 -127 0 feedthrough
rlabel pdiffusion 682 -127 682 -127 0 feedthrough
rlabel pdiffusion 689 -127 689 -127 0 feedthrough
rlabel pdiffusion 696 -127 696 -127 0 feedthrough
rlabel pdiffusion 703 -127 703 -127 0 feedthrough
rlabel pdiffusion 710 -127 710 -127 0 feedthrough
rlabel pdiffusion 717 -127 717 -127 0 feedthrough
rlabel pdiffusion 724 -127 724 -127 0 feedthrough
rlabel pdiffusion 731 -127 731 -127 0 feedthrough
rlabel pdiffusion 738 -127 738 -127 0 feedthrough
rlabel pdiffusion 745 -127 745 -127 0 feedthrough
rlabel pdiffusion 752 -127 752 -127 0 feedthrough
rlabel pdiffusion 759 -127 759 -127 0 feedthrough
rlabel pdiffusion 766 -127 766 -127 0 feedthrough
rlabel pdiffusion 773 -127 773 -127 0 feedthrough
rlabel pdiffusion 780 -127 780 -127 0 feedthrough
rlabel pdiffusion 787 -127 787 -127 0 feedthrough
rlabel pdiffusion 794 -127 794 -127 0 feedthrough
rlabel pdiffusion 801 -127 801 -127 0 feedthrough
rlabel pdiffusion 808 -127 808 -127 0 feedthrough
rlabel pdiffusion 815 -127 815 -127 0 feedthrough
rlabel pdiffusion 822 -127 822 -127 0 feedthrough
rlabel pdiffusion 829 -127 829 -127 0 feedthrough
rlabel pdiffusion 836 -127 836 -127 0 feedthrough
rlabel pdiffusion 843 -127 843 -127 0 cellNo=332
rlabel pdiffusion 871 -127 871 -127 0 feedthrough
rlabel pdiffusion 878 -127 878 -127 0 feedthrough
rlabel pdiffusion 1109 -127 1109 -127 0 cellNo=897
rlabel pdiffusion 3 -216 3 -216 0 cellNo=133
rlabel pdiffusion 10 -216 10 -216 0 cellNo=190
rlabel pdiffusion 17 -216 17 -216 0 cellNo=768
rlabel pdiffusion 24 -216 24 -216 0 feedthrough
rlabel pdiffusion 31 -216 31 -216 0 feedthrough
rlabel pdiffusion 38 -216 38 -216 0 feedthrough
rlabel pdiffusion 45 -216 45 -216 0 feedthrough
rlabel pdiffusion 52 -216 52 -216 0 feedthrough
rlabel pdiffusion 59 -216 59 -216 0 feedthrough
rlabel pdiffusion 66 -216 66 -216 0 feedthrough
rlabel pdiffusion 73 -216 73 -216 0 cellNo=56
rlabel pdiffusion 80 -216 80 -216 0 feedthrough
rlabel pdiffusion 87 -216 87 -216 0 cellNo=745
rlabel pdiffusion 94 -216 94 -216 0 feedthrough
rlabel pdiffusion 101 -216 101 -216 0 feedthrough
rlabel pdiffusion 108 -216 108 -216 0 cellNo=219
rlabel pdiffusion 115 -216 115 -216 0 feedthrough
rlabel pdiffusion 122 -216 122 -216 0 cellNo=249
rlabel pdiffusion 129 -216 129 -216 0 feedthrough
rlabel pdiffusion 136 -216 136 -216 0 feedthrough
rlabel pdiffusion 143 -216 143 -216 0 cellNo=314
rlabel pdiffusion 150 -216 150 -216 0 cellNo=708
rlabel pdiffusion 157 -216 157 -216 0 feedthrough
rlabel pdiffusion 164 -216 164 -216 0 feedthrough
rlabel pdiffusion 171 -216 171 -216 0 feedthrough
rlabel pdiffusion 178 -216 178 -216 0 cellNo=644
rlabel pdiffusion 185 -216 185 -216 0 feedthrough
rlabel pdiffusion 192 -216 192 -216 0 feedthrough
rlabel pdiffusion 199 -216 199 -216 0 feedthrough
rlabel pdiffusion 206 -216 206 -216 0 cellNo=634
rlabel pdiffusion 213 -216 213 -216 0 cellNo=436
rlabel pdiffusion 220 -216 220 -216 0 cellNo=393
rlabel pdiffusion 227 -216 227 -216 0 cellNo=751
rlabel pdiffusion 234 -216 234 -216 0 cellNo=152
rlabel pdiffusion 241 -216 241 -216 0 feedthrough
rlabel pdiffusion 248 -216 248 -216 0 cellNo=217
rlabel pdiffusion 255 -216 255 -216 0 feedthrough
rlabel pdiffusion 262 -216 262 -216 0 feedthrough
rlabel pdiffusion 269 -216 269 -216 0 feedthrough
rlabel pdiffusion 276 -216 276 -216 0 feedthrough
rlabel pdiffusion 283 -216 283 -216 0 feedthrough
rlabel pdiffusion 290 -216 290 -216 0 feedthrough
rlabel pdiffusion 297 -216 297 -216 0 cellNo=765
rlabel pdiffusion 304 -216 304 -216 0 feedthrough
rlabel pdiffusion 311 -216 311 -216 0 feedthrough
rlabel pdiffusion 318 -216 318 -216 0 feedthrough
rlabel pdiffusion 325 -216 325 -216 0 cellNo=257
rlabel pdiffusion 332 -216 332 -216 0 cellNo=935
rlabel pdiffusion 339 -216 339 -216 0 feedthrough
rlabel pdiffusion 346 -216 346 -216 0 cellNo=617
rlabel pdiffusion 353 -216 353 -216 0 feedthrough
rlabel pdiffusion 360 -216 360 -216 0 cellNo=727
rlabel pdiffusion 367 -216 367 -216 0 feedthrough
rlabel pdiffusion 374 -216 374 -216 0 feedthrough
rlabel pdiffusion 381 -216 381 -216 0 feedthrough
rlabel pdiffusion 388 -216 388 -216 0 cellNo=512
rlabel pdiffusion 395 -216 395 -216 0 cellNo=524
rlabel pdiffusion 402 -216 402 -216 0 cellNo=443
rlabel pdiffusion 409 -216 409 -216 0 feedthrough
rlabel pdiffusion 416 -216 416 -216 0 feedthrough
rlabel pdiffusion 423 -216 423 -216 0 feedthrough
rlabel pdiffusion 430 -216 430 -216 0 feedthrough
rlabel pdiffusion 437 -216 437 -216 0 feedthrough
rlabel pdiffusion 444 -216 444 -216 0 feedthrough
rlabel pdiffusion 451 -216 451 -216 0 feedthrough
rlabel pdiffusion 458 -216 458 -216 0 cellNo=779
rlabel pdiffusion 465 -216 465 -216 0 feedthrough
rlabel pdiffusion 472 -216 472 -216 0 feedthrough
rlabel pdiffusion 479 -216 479 -216 0 feedthrough
rlabel pdiffusion 486 -216 486 -216 0 feedthrough
rlabel pdiffusion 493 -216 493 -216 0 cellNo=596
rlabel pdiffusion 500 -216 500 -216 0 feedthrough
rlabel pdiffusion 507 -216 507 -216 0 feedthrough
rlabel pdiffusion 514 -216 514 -216 0 feedthrough
rlabel pdiffusion 521 -216 521 -216 0 cellNo=299
rlabel pdiffusion 528 -216 528 -216 0 feedthrough
rlabel pdiffusion 535 -216 535 -216 0 feedthrough
rlabel pdiffusion 542 -216 542 -216 0 feedthrough
rlabel pdiffusion 549 -216 549 -216 0 feedthrough
rlabel pdiffusion 556 -216 556 -216 0 feedthrough
rlabel pdiffusion 563 -216 563 -216 0 feedthrough
rlabel pdiffusion 570 -216 570 -216 0 feedthrough
rlabel pdiffusion 577 -216 577 -216 0 cellNo=94
rlabel pdiffusion 584 -216 584 -216 0 feedthrough
rlabel pdiffusion 591 -216 591 -216 0 feedthrough
rlabel pdiffusion 598 -216 598 -216 0 feedthrough
rlabel pdiffusion 605 -216 605 -216 0 feedthrough
rlabel pdiffusion 612 -216 612 -216 0 feedthrough
rlabel pdiffusion 619 -216 619 -216 0 cellNo=144
rlabel pdiffusion 626 -216 626 -216 0 cellNo=324
rlabel pdiffusion 633 -216 633 -216 0 feedthrough
rlabel pdiffusion 640 -216 640 -216 0 feedthrough
rlabel pdiffusion 647 -216 647 -216 0 feedthrough
rlabel pdiffusion 654 -216 654 -216 0 cellNo=205
rlabel pdiffusion 661 -216 661 -216 0 feedthrough
rlabel pdiffusion 668 -216 668 -216 0 feedthrough
rlabel pdiffusion 675 -216 675 -216 0 feedthrough
rlabel pdiffusion 682 -216 682 -216 0 feedthrough
rlabel pdiffusion 689 -216 689 -216 0 feedthrough
rlabel pdiffusion 696 -216 696 -216 0 feedthrough
rlabel pdiffusion 703 -216 703 -216 0 feedthrough
rlabel pdiffusion 710 -216 710 -216 0 feedthrough
rlabel pdiffusion 717 -216 717 -216 0 feedthrough
rlabel pdiffusion 724 -216 724 -216 0 feedthrough
rlabel pdiffusion 731 -216 731 -216 0 feedthrough
rlabel pdiffusion 738 -216 738 -216 0 cellNo=793
rlabel pdiffusion 745 -216 745 -216 0 feedthrough
rlabel pdiffusion 752 -216 752 -216 0 feedthrough
rlabel pdiffusion 759 -216 759 -216 0 feedthrough
rlabel pdiffusion 766 -216 766 -216 0 feedthrough
rlabel pdiffusion 773 -216 773 -216 0 feedthrough
rlabel pdiffusion 780 -216 780 -216 0 feedthrough
rlabel pdiffusion 787 -216 787 -216 0 feedthrough
rlabel pdiffusion 794 -216 794 -216 0 feedthrough
rlabel pdiffusion 801 -216 801 -216 0 feedthrough
rlabel pdiffusion 808 -216 808 -216 0 feedthrough
rlabel pdiffusion 815 -216 815 -216 0 feedthrough
rlabel pdiffusion 822 -216 822 -216 0 feedthrough
rlabel pdiffusion 829 -216 829 -216 0 feedthrough
rlabel pdiffusion 836 -216 836 -216 0 feedthrough
rlabel pdiffusion 843 -216 843 -216 0 feedthrough
rlabel pdiffusion 850 -216 850 -216 0 feedthrough
rlabel pdiffusion 857 -216 857 -216 0 feedthrough
rlabel pdiffusion 864 -216 864 -216 0 feedthrough
rlabel pdiffusion 871 -216 871 -216 0 feedthrough
rlabel pdiffusion 878 -216 878 -216 0 feedthrough
rlabel pdiffusion 885 -216 885 -216 0 feedthrough
rlabel pdiffusion 892 -216 892 -216 0 feedthrough
rlabel pdiffusion 899 -216 899 -216 0 feedthrough
rlabel pdiffusion 906 -216 906 -216 0 feedthrough
rlabel pdiffusion 913 -216 913 -216 0 feedthrough
rlabel pdiffusion 920 -216 920 -216 0 feedthrough
rlabel pdiffusion 927 -216 927 -216 0 feedthrough
rlabel pdiffusion 934 -216 934 -216 0 feedthrough
rlabel pdiffusion 941 -216 941 -216 0 feedthrough
rlabel pdiffusion 948 -216 948 -216 0 feedthrough
rlabel pdiffusion 955 -216 955 -216 0 feedthrough
rlabel pdiffusion 1109 -216 1109 -216 0 feedthrough
rlabel pdiffusion 3 -299 3 -299 0 cellNo=556
rlabel pdiffusion 10 -299 10 -299 0 cellNo=696
rlabel pdiffusion 17 -299 17 -299 0 feedthrough
rlabel pdiffusion 24 -299 24 -299 0 feedthrough
rlabel pdiffusion 31 -299 31 -299 0 feedthrough
rlabel pdiffusion 38 -299 38 -299 0 feedthrough
rlabel pdiffusion 45 -299 45 -299 0 cellNo=11
rlabel pdiffusion 52 -299 52 -299 0 feedthrough
rlabel pdiffusion 59 -299 59 -299 0 feedthrough
rlabel pdiffusion 66 -299 66 -299 0 cellNo=194
rlabel pdiffusion 73 -299 73 -299 0 feedthrough
rlabel pdiffusion 80 -299 80 -299 0 feedthrough
rlabel pdiffusion 87 -299 87 -299 0 feedthrough
rlabel pdiffusion 94 -299 94 -299 0 feedthrough
rlabel pdiffusion 101 -299 101 -299 0 cellNo=222
rlabel pdiffusion 108 -299 108 -299 0 feedthrough
rlabel pdiffusion 115 -299 115 -299 0 cellNo=909
rlabel pdiffusion 122 -299 122 -299 0 cellNo=240
rlabel pdiffusion 129 -299 129 -299 0 cellNo=738
rlabel pdiffusion 136 -299 136 -299 0 cellNo=368
rlabel pdiffusion 143 -299 143 -299 0 feedthrough
rlabel pdiffusion 150 -299 150 -299 0 feedthrough
rlabel pdiffusion 157 -299 157 -299 0 feedthrough
rlabel pdiffusion 164 -299 164 -299 0 cellNo=223
rlabel pdiffusion 171 -299 171 -299 0 cellNo=514
rlabel pdiffusion 178 -299 178 -299 0 feedthrough
rlabel pdiffusion 185 -299 185 -299 0 cellNo=754
rlabel pdiffusion 192 -299 192 -299 0 cellNo=871
rlabel pdiffusion 199 -299 199 -299 0 feedthrough
rlabel pdiffusion 206 -299 206 -299 0 cellNo=59
rlabel pdiffusion 213 -299 213 -299 0 feedthrough
rlabel pdiffusion 220 -299 220 -299 0 feedthrough
rlabel pdiffusion 227 -299 227 -299 0 feedthrough
rlabel pdiffusion 234 -299 234 -299 0 feedthrough
rlabel pdiffusion 241 -299 241 -299 0 feedthrough
rlabel pdiffusion 248 -299 248 -299 0 feedthrough
rlabel pdiffusion 255 -299 255 -299 0 cellNo=191
rlabel pdiffusion 262 -299 262 -299 0 feedthrough
rlabel pdiffusion 269 -299 269 -299 0 feedthrough
rlabel pdiffusion 276 -299 276 -299 0 feedthrough
rlabel pdiffusion 283 -299 283 -299 0 feedthrough
rlabel pdiffusion 290 -299 290 -299 0 feedthrough
rlabel pdiffusion 297 -299 297 -299 0 cellNo=559
rlabel pdiffusion 304 -299 304 -299 0 feedthrough
rlabel pdiffusion 311 -299 311 -299 0 feedthrough
rlabel pdiffusion 318 -299 318 -299 0 cellNo=520
rlabel pdiffusion 325 -299 325 -299 0 feedthrough
rlabel pdiffusion 332 -299 332 -299 0 feedthrough
rlabel pdiffusion 339 -299 339 -299 0 feedthrough
rlabel pdiffusion 346 -299 346 -299 0 feedthrough
rlabel pdiffusion 353 -299 353 -299 0 cellNo=229
rlabel pdiffusion 360 -299 360 -299 0 cellNo=376
rlabel pdiffusion 367 -299 367 -299 0 feedthrough
rlabel pdiffusion 374 -299 374 -299 0 cellNo=131
rlabel pdiffusion 381 -299 381 -299 0 feedthrough
rlabel pdiffusion 388 -299 388 -299 0 feedthrough
rlabel pdiffusion 395 -299 395 -299 0 cellNo=703
rlabel pdiffusion 402 -299 402 -299 0 cellNo=169
rlabel pdiffusion 409 -299 409 -299 0 feedthrough
rlabel pdiffusion 416 -299 416 -299 0 feedthrough
rlabel pdiffusion 423 -299 423 -299 0 feedthrough
rlabel pdiffusion 430 -299 430 -299 0 feedthrough
rlabel pdiffusion 437 -299 437 -299 0 cellNo=48
rlabel pdiffusion 444 -299 444 -299 0 feedthrough
rlabel pdiffusion 451 -299 451 -299 0 feedthrough
rlabel pdiffusion 458 -299 458 -299 0 feedthrough
rlabel pdiffusion 465 -299 465 -299 0 cellNo=461
rlabel pdiffusion 472 -299 472 -299 0 feedthrough
rlabel pdiffusion 479 -299 479 -299 0 feedthrough
rlabel pdiffusion 486 -299 486 -299 0 cellNo=619
rlabel pdiffusion 493 -299 493 -299 0 feedthrough
rlabel pdiffusion 500 -299 500 -299 0 cellNo=576
rlabel pdiffusion 507 -299 507 -299 0 feedthrough
rlabel pdiffusion 514 -299 514 -299 0 feedthrough
rlabel pdiffusion 521 -299 521 -299 0 cellNo=456
rlabel pdiffusion 528 -299 528 -299 0 feedthrough
rlabel pdiffusion 535 -299 535 -299 0 feedthrough
rlabel pdiffusion 542 -299 542 -299 0 feedthrough
rlabel pdiffusion 549 -299 549 -299 0 feedthrough
rlabel pdiffusion 556 -299 556 -299 0 feedthrough
rlabel pdiffusion 563 -299 563 -299 0 feedthrough
rlabel pdiffusion 570 -299 570 -299 0 feedthrough
rlabel pdiffusion 577 -299 577 -299 0 feedthrough
rlabel pdiffusion 584 -299 584 -299 0 feedthrough
rlabel pdiffusion 591 -299 591 -299 0 feedthrough
rlabel pdiffusion 598 -299 598 -299 0 feedthrough
rlabel pdiffusion 605 -299 605 -299 0 feedthrough
rlabel pdiffusion 612 -299 612 -299 0 feedthrough
rlabel pdiffusion 619 -299 619 -299 0 feedthrough
rlabel pdiffusion 626 -299 626 -299 0 feedthrough
rlabel pdiffusion 633 -299 633 -299 0 feedthrough
rlabel pdiffusion 640 -299 640 -299 0 feedthrough
rlabel pdiffusion 647 -299 647 -299 0 feedthrough
rlabel pdiffusion 654 -299 654 -299 0 feedthrough
rlabel pdiffusion 661 -299 661 -299 0 cellNo=853
rlabel pdiffusion 668 -299 668 -299 0 feedthrough
rlabel pdiffusion 675 -299 675 -299 0 feedthrough
rlabel pdiffusion 682 -299 682 -299 0 feedthrough
rlabel pdiffusion 689 -299 689 -299 0 feedthrough
rlabel pdiffusion 696 -299 696 -299 0 feedthrough
rlabel pdiffusion 703 -299 703 -299 0 feedthrough
rlabel pdiffusion 710 -299 710 -299 0 feedthrough
rlabel pdiffusion 717 -299 717 -299 0 feedthrough
rlabel pdiffusion 724 -299 724 -299 0 feedthrough
rlabel pdiffusion 731 -299 731 -299 0 feedthrough
rlabel pdiffusion 738 -299 738 -299 0 feedthrough
rlabel pdiffusion 745 -299 745 -299 0 feedthrough
rlabel pdiffusion 752 -299 752 -299 0 feedthrough
rlabel pdiffusion 759 -299 759 -299 0 feedthrough
rlabel pdiffusion 766 -299 766 -299 0 feedthrough
rlabel pdiffusion 773 -299 773 -299 0 feedthrough
rlabel pdiffusion 780 -299 780 -299 0 feedthrough
rlabel pdiffusion 787 -299 787 -299 0 feedthrough
rlabel pdiffusion 794 -299 794 -299 0 feedthrough
rlabel pdiffusion 801 -299 801 -299 0 feedthrough
rlabel pdiffusion 808 -299 808 -299 0 feedthrough
rlabel pdiffusion 815 -299 815 -299 0 feedthrough
rlabel pdiffusion 822 -299 822 -299 0 feedthrough
rlabel pdiffusion 829 -299 829 -299 0 feedthrough
rlabel pdiffusion 836 -299 836 -299 0 feedthrough
rlabel pdiffusion 843 -299 843 -299 0 feedthrough
rlabel pdiffusion 850 -299 850 -299 0 feedthrough
rlabel pdiffusion 857 -299 857 -299 0 feedthrough
rlabel pdiffusion 864 -299 864 -299 0 feedthrough
rlabel pdiffusion 871 -299 871 -299 0 feedthrough
rlabel pdiffusion 878 -299 878 -299 0 feedthrough
rlabel pdiffusion 885 -299 885 -299 0 cellNo=308
rlabel pdiffusion 892 -299 892 -299 0 cellNo=278
rlabel pdiffusion 899 -299 899 -299 0 cellNo=720
rlabel pdiffusion 906 -299 906 -299 0 cellNo=515
rlabel pdiffusion 913 -299 913 -299 0 feedthrough
rlabel pdiffusion 920 -299 920 -299 0 feedthrough
rlabel pdiffusion 1109 -299 1109 -299 0 feedthrough
rlabel pdiffusion 3 -394 3 -394 0 cellNo=448
rlabel pdiffusion 10 -394 10 -394 0 feedthrough
rlabel pdiffusion 17 -394 17 -394 0 cellNo=377
rlabel pdiffusion 24 -394 24 -394 0 feedthrough
rlabel pdiffusion 31 -394 31 -394 0 cellNo=307
rlabel pdiffusion 38 -394 38 -394 0 feedthrough
rlabel pdiffusion 45 -394 45 -394 0 feedthrough
rlabel pdiffusion 52 -394 52 -394 0 feedthrough
rlabel pdiffusion 59 -394 59 -394 0 feedthrough
rlabel pdiffusion 66 -394 66 -394 0 cellNo=224
rlabel pdiffusion 73 -394 73 -394 0 feedthrough
rlabel pdiffusion 80 -394 80 -394 0 cellNo=156
rlabel pdiffusion 87 -394 87 -394 0 feedthrough
rlabel pdiffusion 94 -394 94 -394 0 cellNo=927
rlabel pdiffusion 101 -394 101 -394 0 feedthrough
rlabel pdiffusion 108 -394 108 -394 0 cellNo=565
rlabel pdiffusion 115 -394 115 -394 0 cellNo=125
rlabel pdiffusion 122 -394 122 -394 0 cellNo=370
rlabel pdiffusion 129 -394 129 -394 0 feedthrough
rlabel pdiffusion 136 -394 136 -394 0 cellNo=33
rlabel pdiffusion 143 -394 143 -394 0 feedthrough
rlabel pdiffusion 150 -394 150 -394 0 feedthrough
rlabel pdiffusion 157 -394 157 -394 0 cellNo=407
rlabel pdiffusion 164 -394 164 -394 0 feedthrough
rlabel pdiffusion 171 -394 171 -394 0 cellNo=233
rlabel pdiffusion 178 -394 178 -394 0 feedthrough
rlabel pdiffusion 185 -394 185 -394 0 cellNo=993
rlabel pdiffusion 192 -394 192 -394 0 feedthrough
rlabel pdiffusion 199 -394 199 -394 0 feedthrough
rlabel pdiffusion 206 -394 206 -394 0 feedthrough
rlabel pdiffusion 213 -394 213 -394 0 cellNo=747
rlabel pdiffusion 220 -394 220 -394 0 feedthrough
rlabel pdiffusion 227 -394 227 -394 0 feedthrough
rlabel pdiffusion 234 -394 234 -394 0 feedthrough
rlabel pdiffusion 241 -394 241 -394 0 feedthrough
rlabel pdiffusion 248 -394 248 -394 0 cellNo=107
rlabel pdiffusion 255 -394 255 -394 0 cellNo=840
rlabel pdiffusion 262 -394 262 -394 0 cellNo=72
rlabel pdiffusion 269 -394 269 -394 0 feedthrough
rlabel pdiffusion 276 -394 276 -394 0 feedthrough
rlabel pdiffusion 283 -394 283 -394 0 feedthrough
rlabel pdiffusion 290 -394 290 -394 0 feedthrough
rlabel pdiffusion 297 -394 297 -394 0 feedthrough
rlabel pdiffusion 304 -394 304 -394 0 cellNo=418
rlabel pdiffusion 311 -394 311 -394 0 feedthrough
rlabel pdiffusion 318 -394 318 -394 0 cellNo=142
rlabel pdiffusion 325 -394 325 -394 0 cellNo=268
rlabel pdiffusion 332 -394 332 -394 0 feedthrough
rlabel pdiffusion 339 -394 339 -394 0 cellNo=315
rlabel pdiffusion 346 -394 346 -394 0 feedthrough
rlabel pdiffusion 353 -394 353 -394 0 feedthrough
rlabel pdiffusion 360 -394 360 -394 0 feedthrough
rlabel pdiffusion 367 -394 367 -394 0 feedthrough
rlabel pdiffusion 374 -394 374 -394 0 cellNo=97
rlabel pdiffusion 381 -394 381 -394 0 cellNo=575
rlabel pdiffusion 388 -394 388 -394 0 feedthrough
rlabel pdiffusion 395 -394 395 -394 0 cellNo=752
rlabel pdiffusion 402 -394 402 -394 0 feedthrough
rlabel pdiffusion 409 -394 409 -394 0 feedthrough
rlabel pdiffusion 416 -394 416 -394 0 feedthrough
rlabel pdiffusion 423 -394 423 -394 0 feedthrough
rlabel pdiffusion 430 -394 430 -394 0 feedthrough
rlabel pdiffusion 437 -394 437 -394 0 feedthrough
rlabel pdiffusion 444 -394 444 -394 0 feedthrough
rlabel pdiffusion 451 -394 451 -394 0 feedthrough
rlabel pdiffusion 458 -394 458 -394 0 feedthrough
rlabel pdiffusion 465 -394 465 -394 0 feedthrough
rlabel pdiffusion 472 -394 472 -394 0 cellNo=679
rlabel pdiffusion 479 -394 479 -394 0 feedthrough
rlabel pdiffusion 486 -394 486 -394 0 feedthrough
rlabel pdiffusion 493 -394 493 -394 0 cellNo=464
rlabel pdiffusion 500 -394 500 -394 0 feedthrough
rlabel pdiffusion 507 -394 507 -394 0 feedthrough
rlabel pdiffusion 514 -394 514 -394 0 cellNo=161
rlabel pdiffusion 521 -394 521 -394 0 feedthrough
rlabel pdiffusion 528 -394 528 -394 0 feedthrough
rlabel pdiffusion 535 -394 535 -394 0 feedthrough
rlabel pdiffusion 542 -394 542 -394 0 cellNo=264
rlabel pdiffusion 549 -394 549 -394 0 feedthrough
rlabel pdiffusion 556 -394 556 -394 0 feedthrough
rlabel pdiffusion 563 -394 563 -394 0 feedthrough
rlabel pdiffusion 570 -394 570 -394 0 feedthrough
rlabel pdiffusion 577 -394 577 -394 0 feedthrough
rlabel pdiffusion 584 -394 584 -394 0 feedthrough
rlabel pdiffusion 591 -394 591 -394 0 feedthrough
rlabel pdiffusion 598 -394 598 -394 0 feedthrough
rlabel pdiffusion 605 -394 605 -394 0 feedthrough
rlabel pdiffusion 612 -394 612 -394 0 feedthrough
rlabel pdiffusion 619 -394 619 -394 0 feedthrough
rlabel pdiffusion 626 -394 626 -394 0 cellNo=943
rlabel pdiffusion 633 -394 633 -394 0 feedthrough
rlabel pdiffusion 640 -394 640 -394 0 feedthrough
rlabel pdiffusion 647 -394 647 -394 0 feedthrough
rlabel pdiffusion 654 -394 654 -394 0 feedthrough
rlabel pdiffusion 661 -394 661 -394 0 feedthrough
rlabel pdiffusion 668 -394 668 -394 0 cellNo=604
rlabel pdiffusion 675 -394 675 -394 0 feedthrough
rlabel pdiffusion 682 -394 682 -394 0 feedthrough
rlabel pdiffusion 689 -394 689 -394 0 feedthrough
rlabel pdiffusion 696 -394 696 -394 0 feedthrough
rlabel pdiffusion 703 -394 703 -394 0 feedthrough
rlabel pdiffusion 710 -394 710 -394 0 feedthrough
rlabel pdiffusion 717 -394 717 -394 0 feedthrough
rlabel pdiffusion 724 -394 724 -394 0 feedthrough
rlabel pdiffusion 731 -394 731 -394 0 feedthrough
rlabel pdiffusion 738 -394 738 -394 0 feedthrough
rlabel pdiffusion 745 -394 745 -394 0 feedthrough
rlabel pdiffusion 752 -394 752 -394 0 feedthrough
rlabel pdiffusion 759 -394 759 -394 0 feedthrough
rlabel pdiffusion 766 -394 766 -394 0 feedthrough
rlabel pdiffusion 773 -394 773 -394 0 feedthrough
rlabel pdiffusion 780 -394 780 -394 0 feedthrough
rlabel pdiffusion 787 -394 787 -394 0 feedthrough
rlabel pdiffusion 794 -394 794 -394 0 feedthrough
rlabel pdiffusion 801 -394 801 -394 0 feedthrough
rlabel pdiffusion 808 -394 808 -394 0 feedthrough
rlabel pdiffusion 815 -394 815 -394 0 feedthrough
rlabel pdiffusion 822 -394 822 -394 0 feedthrough
rlabel pdiffusion 829 -394 829 -394 0 feedthrough
rlabel pdiffusion 836 -394 836 -394 0 feedthrough
rlabel pdiffusion 843 -394 843 -394 0 feedthrough
rlabel pdiffusion 850 -394 850 -394 0 feedthrough
rlabel pdiffusion 857 -394 857 -394 0 feedthrough
rlabel pdiffusion 864 -394 864 -394 0 feedthrough
rlabel pdiffusion 871 -394 871 -394 0 feedthrough
rlabel pdiffusion 878 -394 878 -394 0 cellNo=230
rlabel pdiffusion 885 -394 885 -394 0 cellNo=506
rlabel pdiffusion 892 -394 892 -394 0 feedthrough
rlabel pdiffusion 899 -394 899 -394 0 feedthrough
rlabel pdiffusion 906 -394 906 -394 0 feedthrough
rlabel pdiffusion 934 -394 934 -394 0 feedthrough
rlabel pdiffusion 1109 -394 1109 -394 0 feedthrough
rlabel pdiffusion 3 -483 3 -483 0 feedthrough
rlabel pdiffusion 10 -483 10 -483 0 cellNo=262
rlabel pdiffusion 17 -483 17 -483 0 feedthrough
rlabel pdiffusion 24 -483 24 -483 0 feedthrough
rlabel pdiffusion 31 -483 31 -483 0 feedthrough
rlabel pdiffusion 38 -483 38 -483 0 feedthrough
rlabel pdiffusion 45 -483 45 -483 0 feedthrough
rlabel pdiffusion 52 -483 52 -483 0 feedthrough
rlabel pdiffusion 59 -483 59 -483 0 cellNo=25
rlabel pdiffusion 66 -483 66 -483 0 cellNo=327
rlabel pdiffusion 73 -483 73 -483 0 feedthrough
rlabel pdiffusion 80 -483 80 -483 0 feedthrough
rlabel pdiffusion 87 -483 87 -483 0 feedthrough
rlabel pdiffusion 94 -483 94 -483 0 feedthrough
rlabel pdiffusion 101 -483 101 -483 0 feedthrough
rlabel pdiffusion 108 -483 108 -483 0 feedthrough
rlabel pdiffusion 115 -483 115 -483 0 feedthrough
rlabel pdiffusion 122 -483 122 -483 0 cellNo=646
rlabel pdiffusion 129 -483 129 -483 0 cellNo=699
rlabel pdiffusion 136 -483 136 -483 0 feedthrough
rlabel pdiffusion 143 -483 143 -483 0 cellNo=537
rlabel pdiffusion 150 -483 150 -483 0 feedthrough
rlabel pdiffusion 157 -483 157 -483 0 feedthrough
rlabel pdiffusion 164 -483 164 -483 0 feedthrough
rlabel pdiffusion 171 -483 171 -483 0 feedthrough
rlabel pdiffusion 178 -483 178 -483 0 cellNo=678
rlabel pdiffusion 185 -483 185 -483 0 feedthrough
rlabel pdiffusion 192 -483 192 -483 0 feedthrough
rlabel pdiffusion 199 -483 199 -483 0 cellNo=76
rlabel pdiffusion 206 -483 206 -483 0 cellNo=649
rlabel pdiffusion 213 -483 213 -483 0 feedthrough
rlabel pdiffusion 220 -483 220 -483 0 feedthrough
rlabel pdiffusion 227 -483 227 -483 0 feedthrough
rlabel pdiffusion 234 -483 234 -483 0 feedthrough
rlabel pdiffusion 241 -483 241 -483 0 feedthrough
rlabel pdiffusion 248 -483 248 -483 0 feedthrough
rlabel pdiffusion 255 -483 255 -483 0 feedthrough
rlabel pdiffusion 262 -483 262 -483 0 feedthrough
rlabel pdiffusion 269 -483 269 -483 0 feedthrough
rlabel pdiffusion 276 -483 276 -483 0 feedthrough
rlabel pdiffusion 283 -483 283 -483 0 cellNo=19
rlabel pdiffusion 290 -483 290 -483 0 feedthrough
rlabel pdiffusion 297 -483 297 -483 0 feedthrough
rlabel pdiffusion 304 -483 304 -483 0 feedthrough
rlabel pdiffusion 311 -483 311 -483 0 feedthrough
rlabel pdiffusion 318 -483 318 -483 0 feedthrough
rlabel pdiffusion 325 -483 325 -483 0 cellNo=740
rlabel pdiffusion 332 -483 332 -483 0 feedthrough
rlabel pdiffusion 339 -483 339 -483 0 feedthrough
rlabel pdiffusion 346 -483 346 -483 0 cellNo=66
rlabel pdiffusion 353 -483 353 -483 0 cellNo=300
rlabel pdiffusion 360 -483 360 -483 0 feedthrough
rlabel pdiffusion 367 -483 367 -483 0 feedthrough
rlabel pdiffusion 374 -483 374 -483 0 feedthrough
rlabel pdiffusion 381 -483 381 -483 0 cellNo=766
rlabel pdiffusion 388 -483 388 -483 0 feedthrough
rlabel pdiffusion 395 -483 395 -483 0 cellNo=999
rlabel pdiffusion 402 -483 402 -483 0 feedthrough
rlabel pdiffusion 409 -483 409 -483 0 feedthrough
rlabel pdiffusion 416 -483 416 -483 0 cellNo=917
rlabel pdiffusion 423 -483 423 -483 0 cellNo=711
rlabel pdiffusion 430 -483 430 -483 0 feedthrough
rlabel pdiffusion 437 -483 437 -483 0 feedthrough
rlabel pdiffusion 444 -483 444 -483 0 feedthrough
rlabel pdiffusion 451 -483 451 -483 0 feedthrough
rlabel pdiffusion 458 -483 458 -483 0 cellNo=830
rlabel pdiffusion 465 -483 465 -483 0 feedthrough
rlabel pdiffusion 472 -483 472 -483 0 cellNo=60
rlabel pdiffusion 479 -483 479 -483 0 cellNo=616
rlabel pdiffusion 486 -483 486 -483 0 feedthrough
rlabel pdiffusion 493 -483 493 -483 0 feedthrough
rlabel pdiffusion 500 -483 500 -483 0 cellNo=925
rlabel pdiffusion 507 -483 507 -483 0 feedthrough
rlabel pdiffusion 514 -483 514 -483 0 feedthrough
rlabel pdiffusion 521 -483 521 -483 0 feedthrough
rlabel pdiffusion 528 -483 528 -483 0 feedthrough
rlabel pdiffusion 535 -483 535 -483 0 cellNo=57
rlabel pdiffusion 542 -483 542 -483 0 feedthrough
rlabel pdiffusion 549 -483 549 -483 0 feedthrough
rlabel pdiffusion 556 -483 556 -483 0 cellNo=289
rlabel pdiffusion 563 -483 563 -483 0 cellNo=366
rlabel pdiffusion 570 -483 570 -483 0 cellNo=349
rlabel pdiffusion 577 -483 577 -483 0 cellNo=608
rlabel pdiffusion 584 -483 584 -483 0 feedthrough
rlabel pdiffusion 591 -483 591 -483 0 feedthrough
rlabel pdiffusion 598 -483 598 -483 0 feedthrough
rlabel pdiffusion 605 -483 605 -483 0 feedthrough
rlabel pdiffusion 612 -483 612 -483 0 feedthrough
rlabel pdiffusion 619 -483 619 -483 0 feedthrough
rlabel pdiffusion 626 -483 626 -483 0 feedthrough
rlabel pdiffusion 633 -483 633 -483 0 cellNo=581
rlabel pdiffusion 640 -483 640 -483 0 cellNo=760
rlabel pdiffusion 647 -483 647 -483 0 feedthrough
rlabel pdiffusion 654 -483 654 -483 0 feedthrough
rlabel pdiffusion 661 -483 661 -483 0 feedthrough
rlabel pdiffusion 668 -483 668 -483 0 feedthrough
rlabel pdiffusion 675 -483 675 -483 0 feedthrough
rlabel pdiffusion 682 -483 682 -483 0 feedthrough
rlabel pdiffusion 689 -483 689 -483 0 cellNo=384
rlabel pdiffusion 696 -483 696 -483 0 feedthrough
rlabel pdiffusion 703 -483 703 -483 0 feedthrough
rlabel pdiffusion 710 -483 710 -483 0 feedthrough
rlabel pdiffusion 717 -483 717 -483 0 feedthrough
rlabel pdiffusion 724 -483 724 -483 0 feedthrough
rlabel pdiffusion 731 -483 731 -483 0 feedthrough
rlabel pdiffusion 738 -483 738 -483 0 feedthrough
rlabel pdiffusion 745 -483 745 -483 0 feedthrough
rlabel pdiffusion 752 -483 752 -483 0 feedthrough
rlabel pdiffusion 759 -483 759 -483 0 feedthrough
rlabel pdiffusion 766 -483 766 -483 0 feedthrough
rlabel pdiffusion 773 -483 773 -483 0 feedthrough
rlabel pdiffusion 780 -483 780 -483 0 feedthrough
rlabel pdiffusion 787 -483 787 -483 0 feedthrough
rlabel pdiffusion 794 -483 794 -483 0 feedthrough
rlabel pdiffusion 801 -483 801 -483 0 feedthrough
rlabel pdiffusion 808 -483 808 -483 0 feedthrough
rlabel pdiffusion 815 -483 815 -483 0 cellNo=620
rlabel pdiffusion 822 -483 822 -483 0 feedthrough
rlabel pdiffusion 829 -483 829 -483 0 feedthrough
rlabel pdiffusion 836 -483 836 -483 0 feedthrough
rlabel pdiffusion 843 -483 843 -483 0 feedthrough
rlabel pdiffusion 850 -483 850 -483 0 feedthrough
rlabel pdiffusion 857 -483 857 -483 0 feedthrough
rlabel pdiffusion 864 -483 864 -483 0 feedthrough
rlabel pdiffusion 871 -483 871 -483 0 feedthrough
rlabel pdiffusion 878 -483 878 -483 0 feedthrough
rlabel pdiffusion 885 -483 885 -483 0 feedthrough
rlabel pdiffusion 892 -483 892 -483 0 feedthrough
rlabel pdiffusion 899 -483 899 -483 0 feedthrough
rlabel pdiffusion 906 -483 906 -483 0 feedthrough
rlabel pdiffusion 913 -483 913 -483 0 feedthrough
rlabel pdiffusion 920 -483 920 -483 0 feedthrough
rlabel pdiffusion 927 -483 927 -483 0 feedthrough
rlabel pdiffusion 934 -483 934 -483 0 feedthrough
rlabel pdiffusion 941 -483 941 -483 0 feedthrough
rlabel pdiffusion 948 -483 948 -483 0 feedthrough
rlabel pdiffusion 955 -483 955 -483 0 feedthrough
rlabel pdiffusion 962 -483 962 -483 0 feedthrough
rlabel pdiffusion 969 -483 969 -483 0 feedthrough
rlabel pdiffusion 976 -483 976 -483 0 feedthrough
rlabel pdiffusion 983 -483 983 -483 0 feedthrough
rlabel pdiffusion 990 -483 990 -483 0 feedthrough
rlabel pdiffusion 997 -483 997 -483 0 feedthrough
rlabel pdiffusion 1004 -483 1004 -483 0 feedthrough
rlabel pdiffusion 1011 -483 1011 -483 0 feedthrough
rlabel pdiffusion 1018 -483 1018 -483 0 feedthrough
rlabel pdiffusion 1025 -483 1025 -483 0 feedthrough
rlabel pdiffusion 1032 -483 1032 -483 0 cellNo=441
rlabel pdiffusion 1039 -483 1039 -483 0 cellNo=309
rlabel pdiffusion 1046 -483 1046 -483 0 feedthrough
rlabel pdiffusion 1116 -483 1116 -483 0 feedthrough
rlabel pdiffusion 3 -600 3 -600 0 cellNo=929
rlabel pdiffusion 10 -600 10 -600 0 feedthrough
rlabel pdiffusion 17 -600 17 -600 0 feedthrough
rlabel pdiffusion 24 -600 24 -600 0 cellNo=238
rlabel pdiffusion 31 -600 31 -600 0 feedthrough
rlabel pdiffusion 38 -600 38 -600 0 cellNo=545
rlabel pdiffusion 45 -600 45 -600 0 feedthrough
rlabel pdiffusion 52 -600 52 -600 0 feedthrough
rlabel pdiffusion 59 -600 59 -600 0 feedthrough
rlabel pdiffusion 66 -600 66 -600 0 feedthrough
rlabel pdiffusion 73 -600 73 -600 0 feedthrough
rlabel pdiffusion 80 -600 80 -600 0 feedthrough
rlabel pdiffusion 87 -600 87 -600 0 feedthrough
rlabel pdiffusion 94 -600 94 -600 0 cellNo=450
rlabel pdiffusion 101 -600 101 -600 0 cellNo=635
rlabel pdiffusion 108 -600 108 -600 0 cellNo=259
rlabel pdiffusion 115 -600 115 -600 0 feedthrough
rlabel pdiffusion 122 -600 122 -600 0 feedthrough
rlabel pdiffusion 129 -600 129 -600 0 feedthrough
rlabel pdiffusion 136 -600 136 -600 0 cellNo=489
rlabel pdiffusion 143 -600 143 -600 0 feedthrough
rlabel pdiffusion 150 -600 150 -600 0 feedthrough
rlabel pdiffusion 157 -600 157 -600 0 feedthrough
rlabel pdiffusion 164 -600 164 -600 0 cellNo=186
rlabel pdiffusion 171 -600 171 -600 0 feedthrough
rlabel pdiffusion 178 -600 178 -600 0 cellNo=231
rlabel pdiffusion 185 -600 185 -600 0 feedthrough
rlabel pdiffusion 192 -600 192 -600 0 feedthrough
rlabel pdiffusion 199 -600 199 -600 0 feedthrough
rlabel pdiffusion 206 -600 206 -600 0 cellNo=236
rlabel pdiffusion 213 -600 213 -600 0 cellNo=253
rlabel pdiffusion 220 -600 220 -600 0 cellNo=210
rlabel pdiffusion 227 -600 227 -600 0 feedthrough
rlabel pdiffusion 234 -600 234 -600 0 feedthrough
rlabel pdiffusion 241 -600 241 -600 0 feedthrough
rlabel pdiffusion 248 -600 248 -600 0 feedthrough
rlabel pdiffusion 255 -600 255 -600 0 feedthrough
rlabel pdiffusion 262 -600 262 -600 0 feedthrough
rlabel pdiffusion 269 -600 269 -600 0 cellNo=155
rlabel pdiffusion 276 -600 276 -600 0 feedthrough
rlabel pdiffusion 283 -600 283 -600 0 feedthrough
rlabel pdiffusion 290 -600 290 -600 0 feedthrough
rlabel pdiffusion 297 -600 297 -600 0 feedthrough
rlabel pdiffusion 304 -600 304 -600 0 feedthrough
rlabel pdiffusion 311 -600 311 -600 0 feedthrough
rlabel pdiffusion 318 -600 318 -600 0 feedthrough
rlabel pdiffusion 325 -600 325 -600 0 feedthrough
rlabel pdiffusion 332 -600 332 -600 0 feedthrough
rlabel pdiffusion 339 -600 339 -600 0 cellNo=682
rlabel pdiffusion 346 -600 346 -600 0 cellNo=8
rlabel pdiffusion 353 -600 353 -600 0 feedthrough
rlabel pdiffusion 360 -600 360 -600 0 feedthrough
rlabel pdiffusion 367 -600 367 -600 0 feedthrough
rlabel pdiffusion 374 -600 374 -600 0 feedthrough
rlabel pdiffusion 381 -600 381 -600 0 feedthrough
rlabel pdiffusion 388 -600 388 -600 0 feedthrough
rlabel pdiffusion 395 -600 395 -600 0 feedthrough
rlabel pdiffusion 402 -600 402 -600 0 feedthrough
rlabel pdiffusion 409 -600 409 -600 0 feedthrough
rlabel pdiffusion 416 -600 416 -600 0 feedthrough
rlabel pdiffusion 423 -600 423 -600 0 feedthrough
rlabel pdiffusion 430 -600 430 -600 0 feedthrough
rlabel pdiffusion 437 -600 437 -600 0 cellNo=232
rlabel pdiffusion 444 -600 444 -600 0 feedthrough
rlabel pdiffusion 451 -600 451 -600 0 feedthrough
rlabel pdiffusion 458 -600 458 -600 0 feedthrough
rlabel pdiffusion 465 -600 465 -600 0 cellNo=83
rlabel pdiffusion 472 -600 472 -600 0 cellNo=867
rlabel pdiffusion 479 -600 479 -600 0 feedthrough
rlabel pdiffusion 486 -600 486 -600 0 feedthrough
rlabel pdiffusion 493 -600 493 -600 0 feedthrough
rlabel pdiffusion 500 -600 500 -600 0 feedthrough
rlabel pdiffusion 507 -600 507 -600 0 feedthrough
rlabel pdiffusion 514 -600 514 -600 0 feedthrough
rlabel pdiffusion 521 -600 521 -600 0 cellNo=643
rlabel pdiffusion 528 -600 528 -600 0 cellNo=272
rlabel pdiffusion 535 -600 535 -600 0 cellNo=146
rlabel pdiffusion 542 -600 542 -600 0 feedthrough
rlabel pdiffusion 549 -600 549 -600 0 cellNo=597
rlabel pdiffusion 556 -600 556 -600 0 feedthrough
rlabel pdiffusion 563 -600 563 -600 0 cellNo=758
rlabel pdiffusion 570 -600 570 -600 0 cellNo=507
rlabel pdiffusion 577 -600 577 -600 0 cellNo=2
rlabel pdiffusion 584 -600 584 -600 0 feedthrough
rlabel pdiffusion 591 -600 591 -600 0 feedthrough
rlabel pdiffusion 598 -600 598 -600 0 cellNo=214
rlabel pdiffusion 605 -600 605 -600 0 feedthrough
rlabel pdiffusion 612 -600 612 -600 0 feedthrough
rlabel pdiffusion 619 -600 619 -600 0 feedthrough
rlabel pdiffusion 626 -600 626 -600 0 feedthrough
rlabel pdiffusion 633 -600 633 -600 0 cellNo=173
rlabel pdiffusion 640 -600 640 -600 0 feedthrough
rlabel pdiffusion 647 -600 647 -600 0 feedthrough
rlabel pdiffusion 654 -600 654 -600 0 feedthrough
rlabel pdiffusion 661 -600 661 -600 0 feedthrough
rlabel pdiffusion 668 -600 668 -600 0 feedthrough
rlabel pdiffusion 675 -600 675 -600 0 feedthrough
rlabel pdiffusion 682 -600 682 -600 0 cellNo=812
rlabel pdiffusion 689 -600 689 -600 0 feedthrough
rlabel pdiffusion 696 -600 696 -600 0 feedthrough
rlabel pdiffusion 703 -600 703 -600 0 feedthrough
rlabel pdiffusion 710 -600 710 -600 0 cellNo=276
rlabel pdiffusion 717 -600 717 -600 0 feedthrough
rlabel pdiffusion 724 -600 724 -600 0 feedthrough
rlabel pdiffusion 731 -600 731 -600 0 cellNo=551
rlabel pdiffusion 738 -600 738 -600 0 feedthrough
rlabel pdiffusion 745 -600 745 -600 0 feedthrough
rlabel pdiffusion 752 -600 752 -600 0 feedthrough
rlabel pdiffusion 759 -600 759 -600 0 feedthrough
rlabel pdiffusion 766 -600 766 -600 0 feedthrough
rlabel pdiffusion 773 -600 773 -600 0 feedthrough
rlabel pdiffusion 780 -600 780 -600 0 feedthrough
rlabel pdiffusion 787 -600 787 -600 0 feedthrough
rlabel pdiffusion 794 -600 794 -600 0 feedthrough
rlabel pdiffusion 801 -600 801 -600 0 feedthrough
rlabel pdiffusion 808 -600 808 -600 0 feedthrough
rlabel pdiffusion 815 -600 815 -600 0 feedthrough
rlabel pdiffusion 822 -600 822 -600 0 feedthrough
rlabel pdiffusion 829 -600 829 -600 0 feedthrough
rlabel pdiffusion 836 -600 836 -600 0 feedthrough
rlabel pdiffusion 843 -600 843 -600 0 feedthrough
rlabel pdiffusion 850 -600 850 -600 0 feedthrough
rlabel pdiffusion 857 -600 857 -600 0 feedthrough
rlabel pdiffusion 864 -600 864 -600 0 feedthrough
rlabel pdiffusion 871 -600 871 -600 0 feedthrough
rlabel pdiffusion 878 -600 878 -600 0 feedthrough
rlabel pdiffusion 885 -600 885 -600 0 feedthrough
rlabel pdiffusion 892 -600 892 -600 0 feedthrough
rlabel pdiffusion 899 -600 899 -600 0 feedthrough
rlabel pdiffusion 906 -600 906 -600 0 feedthrough
rlabel pdiffusion 913 -600 913 -600 0 feedthrough
rlabel pdiffusion 920 -600 920 -600 0 feedthrough
rlabel pdiffusion 927 -600 927 -600 0 feedthrough
rlabel pdiffusion 934 -600 934 -600 0 feedthrough
rlabel pdiffusion 941 -600 941 -600 0 feedthrough
rlabel pdiffusion 948 -600 948 -600 0 feedthrough
rlabel pdiffusion 955 -600 955 -600 0 feedthrough
rlabel pdiffusion 962 -600 962 -600 0 feedthrough
rlabel pdiffusion 969 -600 969 -600 0 feedthrough
rlabel pdiffusion 976 -600 976 -600 0 feedthrough
rlabel pdiffusion 983 -600 983 -600 0 feedthrough
rlabel pdiffusion 990 -600 990 -600 0 feedthrough
rlabel pdiffusion 997 -600 997 -600 0 feedthrough
rlabel pdiffusion 1004 -600 1004 -600 0 feedthrough
rlabel pdiffusion 1011 -600 1011 -600 0 feedthrough
rlabel pdiffusion 1018 -600 1018 -600 0 feedthrough
rlabel pdiffusion 1025 -600 1025 -600 0 feedthrough
rlabel pdiffusion 1032 -600 1032 -600 0 feedthrough
rlabel pdiffusion 1039 -600 1039 -600 0 feedthrough
rlabel pdiffusion 1046 -600 1046 -600 0 feedthrough
rlabel pdiffusion 1053 -600 1053 -600 0 feedthrough
rlabel pdiffusion 1060 -600 1060 -600 0 feedthrough
rlabel pdiffusion 1067 -600 1067 -600 0 feedthrough
rlabel pdiffusion 1074 -600 1074 -600 0 feedthrough
rlabel pdiffusion 1081 -600 1081 -600 0 feedthrough
rlabel pdiffusion 1088 -600 1088 -600 0 feedthrough
rlabel pdiffusion 1095 -600 1095 -600 0 feedthrough
rlabel pdiffusion 1102 -600 1102 -600 0 cellNo=624
rlabel pdiffusion 1109 -600 1109 -600 0 cellNo=32
rlabel pdiffusion 1116 -600 1116 -600 0 feedthrough
rlabel pdiffusion 1123 -600 1123 -600 0 feedthrough
rlabel pdiffusion 1130 -600 1130 -600 0 feedthrough
rlabel pdiffusion 3 -701 3 -701 0 feedthrough
rlabel pdiffusion 10 -701 10 -701 0 cellNo=111
rlabel pdiffusion 17 -701 17 -701 0 feedthrough
rlabel pdiffusion 24 -701 24 -701 0 feedthrough
rlabel pdiffusion 31 -701 31 -701 0 feedthrough
rlabel pdiffusion 38 -701 38 -701 0 feedthrough
rlabel pdiffusion 45 -701 45 -701 0 cellNo=286
rlabel pdiffusion 52 -701 52 -701 0 feedthrough
rlabel pdiffusion 59 -701 59 -701 0 feedthrough
rlabel pdiffusion 66 -701 66 -701 0 feedthrough
rlabel pdiffusion 73 -701 73 -701 0 feedthrough
rlabel pdiffusion 80 -701 80 -701 0 cellNo=817
rlabel pdiffusion 87 -701 87 -701 0 feedthrough
rlabel pdiffusion 94 -701 94 -701 0 feedthrough
rlabel pdiffusion 101 -701 101 -701 0 feedthrough
rlabel pdiffusion 108 -701 108 -701 0 feedthrough
rlabel pdiffusion 115 -701 115 -701 0 cellNo=260
rlabel pdiffusion 122 -701 122 -701 0 cellNo=409
rlabel pdiffusion 129 -701 129 -701 0 cellNo=451
rlabel pdiffusion 136 -701 136 -701 0 feedthrough
rlabel pdiffusion 143 -701 143 -701 0 feedthrough
rlabel pdiffusion 150 -701 150 -701 0 feedthrough
rlabel pdiffusion 157 -701 157 -701 0 feedthrough
rlabel pdiffusion 164 -701 164 -701 0 feedthrough
rlabel pdiffusion 171 -701 171 -701 0 cellNo=715
rlabel pdiffusion 178 -701 178 -701 0 feedthrough
rlabel pdiffusion 185 -701 185 -701 0 feedthrough
rlabel pdiffusion 192 -701 192 -701 0 cellNo=333
rlabel pdiffusion 199 -701 199 -701 0 cellNo=800
rlabel pdiffusion 206 -701 206 -701 0 cellNo=906
rlabel pdiffusion 213 -701 213 -701 0 feedthrough
rlabel pdiffusion 220 -701 220 -701 0 feedthrough
rlabel pdiffusion 227 -701 227 -701 0 cellNo=490
rlabel pdiffusion 234 -701 234 -701 0 feedthrough
rlabel pdiffusion 241 -701 241 -701 0 feedthrough
rlabel pdiffusion 248 -701 248 -701 0 feedthrough
rlabel pdiffusion 255 -701 255 -701 0 feedthrough
rlabel pdiffusion 262 -701 262 -701 0 feedthrough
rlabel pdiffusion 269 -701 269 -701 0 feedthrough
rlabel pdiffusion 276 -701 276 -701 0 feedthrough
rlabel pdiffusion 283 -701 283 -701 0 feedthrough
rlabel pdiffusion 290 -701 290 -701 0 cellNo=440
rlabel pdiffusion 297 -701 297 -701 0 feedthrough
rlabel pdiffusion 304 -701 304 -701 0 feedthrough
rlabel pdiffusion 311 -701 311 -701 0 cellNo=284
rlabel pdiffusion 318 -701 318 -701 0 feedthrough
rlabel pdiffusion 325 -701 325 -701 0 feedthrough
rlabel pdiffusion 332 -701 332 -701 0 feedthrough
rlabel pdiffusion 339 -701 339 -701 0 feedthrough
rlabel pdiffusion 346 -701 346 -701 0 feedthrough
rlabel pdiffusion 353 -701 353 -701 0 feedthrough
rlabel pdiffusion 360 -701 360 -701 0 cellNo=882
rlabel pdiffusion 367 -701 367 -701 0 feedthrough
rlabel pdiffusion 374 -701 374 -701 0 feedthrough
rlabel pdiffusion 381 -701 381 -701 0 feedthrough
rlabel pdiffusion 388 -701 388 -701 0 feedthrough
rlabel pdiffusion 395 -701 395 -701 0 feedthrough
rlabel pdiffusion 402 -701 402 -701 0 feedthrough
rlabel pdiffusion 409 -701 409 -701 0 feedthrough
rlabel pdiffusion 416 -701 416 -701 0 feedthrough
rlabel pdiffusion 423 -701 423 -701 0 feedthrough
rlabel pdiffusion 430 -701 430 -701 0 feedthrough
rlabel pdiffusion 437 -701 437 -701 0 feedthrough
rlabel pdiffusion 444 -701 444 -701 0 cellNo=911
rlabel pdiffusion 451 -701 451 -701 0 cellNo=547
rlabel pdiffusion 458 -701 458 -701 0 cellNo=466
rlabel pdiffusion 465 -701 465 -701 0 cellNo=802
rlabel pdiffusion 472 -701 472 -701 0 feedthrough
rlabel pdiffusion 479 -701 479 -701 0 cellNo=462
rlabel pdiffusion 486 -701 486 -701 0 feedthrough
rlabel pdiffusion 493 -701 493 -701 0 cellNo=250
rlabel pdiffusion 500 -701 500 -701 0 feedthrough
rlabel pdiffusion 507 -701 507 -701 0 feedthrough
rlabel pdiffusion 514 -701 514 -701 0 cellNo=245
rlabel pdiffusion 521 -701 521 -701 0 feedthrough
rlabel pdiffusion 528 -701 528 -701 0 feedthrough
rlabel pdiffusion 535 -701 535 -701 0 feedthrough
rlabel pdiffusion 542 -701 542 -701 0 cellNo=861
rlabel pdiffusion 549 -701 549 -701 0 feedthrough
rlabel pdiffusion 556 -701 556 -701 0 feedthrough
rlabel pdiffusion 563 -701 563 -701 0 cellNo=803
rlabel pdiffusion 570 -701 570 -701 0 feedthrough
rlabel pdiffusion 577 -701 577 -701 0 feedthrough
rlabel pdiffusion 584 -701 584 -701 0 feedthrough
rlabel pdiffusion 591 -701 591 -701 0 feedthrough
rlabel pdiffusion 598 -701 598 -701 0 feedthrough
rlabel pdiffusion 605 -701 605 -701 0 cellNo=103
rlabel pdiffusion 612 -701 612 -701 0 feedthrough
rlabel pdiffusion 619 -701 619 -701 0 feedthrough
rlabel pdiffusion 626 -701 626 -701 0 feedthrough
rlabel pdiffusion 633 -701 633 -701 0 feedthrough
rlabel pdiffusion 640 -701 640 -701 0 feedthrough
rlabel pdiffusion 647 -701 647 -701 0 feedthrough
rlabel pdiffusion 654 -701 654 -701 0 feedthrough
rlabel pdiffusion 661 -701 661 -701 0 feedthrough
rlabel pdiffusion 668 -701 668 -701 0 cellNo=321
rlabel pdiffusion 675 -701 675 -701 0 feedthrough
rlabel pdiffusion 682 -701 682 -701 0 feedthrough
rlabel pdiffusion 689 -701 689 -701 0 feedthrough
rlabel pdiffusion 696 -701 696 -701 0 feedthrough
rlabel pdiffusion 703 -701 703 -701 0 feedthrough
rlabel pdiffusion 710 -701 710 -701 0 feedthrough
rlabel pdiffusion 717 -701 717 -701 0 feedthrough
rlabel pdiffusion 724 -701 724 -701 0 cellNo=981
rlabel pdiffusion 731 -701 731 -701 0 feedthrough
rlabel pdiffusion 738 -701 738 -701 0 feedthrough
rlabel pdiffusion 745 -701 745 -701 0 cellNo=509
rlabel pdiffusion 752 -701 752 -701 0 feedthrough
rlabel pdiffusion 759 -701 759 -701 0 feedthrough
rlabel pdiffusion 766 -701 766 -701 0 feedthrough
rlabel pdiffusion 773 -701 773 -701 0 cellNo=481
rlabel pdiffusion 780 -701 780 -701 0 feedthrough
rlabel pdiffusion 787 -701 787 -701 0 cellNo=28
rlabel pdiffusion 794 -701 794 -701 0 feedthrough
rlabel pdiffusion 801 -701 801 -701 0 feedthrough
rlabel pdiffusion 808 -701 808 -701 0 feedthrough
rlabel pdiffusion 815 -701 815 -701 0 feedthrough
rlabel pdiffusion 822 -701 822 -701 0 feedthrough
rlabel pdiffusion 829 -701 829 -701 0 feedthrough
rlabel pdiffusion 836 -701 836 -701 0 feedthrough
rlabel pdiffusion 843 -701 843 -701 0 feedthrough
rlabel pdiffusion 850 -701 850 -701 0 feedthrough
rlabel pdiffusion 857 -701 857 -701 0 feedthrough
rlabel pdiffusion 864 -701 864 -701 0 feedthrough
rlabel pdiffusion 871 -701 871 -701 0 feedthrough
rlabel pdiffusion 878 -701 878 -701 0 feedthrough
rlabel pdiffusion 885 -701 885 -701 0 feedthrough
rlabel pdiffusion 892 -701 892 -701 0 feedthrough
rlabel pdiffusion 899 -701 899 -701 0 feedthrough
rlabel pdiffusion 906 -701 906 -701 0 feedthrough
rlabel pdiffusion 913 -701 913 -701 0 feedthrough
rlabel pdiffusion 920 -701 920 -701 0 feedthrough
rlabel pdiffusion 927 -701 927 -701 0 feedthrough
rlabel pdiffusion 934 -701 934 -701 0 feedthrough
rlabel pdiffusion 941 -701 941 -701 0 feedthrough
rlabel pdiffusion 948 -701 948 -701 0 feedthrough
rlabel pdiffusion 955 -701 955 -701 0 feedthrough
rlabel pdiffusion 962 -701 962 -701 0 feedthrough
rlabel pdiffusion 969 -701 969 -701 0 feedthrough
rlabel pdiffusion 976 -701 976 -701 0 feedthrough
rlabel pdiffusion 983 -701 983 -701 0 feedthrough
rlabel pdiffusion 990 -701 990 -701 0 feedthrough
rlabel pdiffusion 997 -701 997 -701 0 feedthrough
rlabel pdiffusion 1004 -701 1004 -701 0 feedthrough
rlabel pdiffusion 1011 -701 1011 -701 0 feedthrough
rlabel pdiffusion 1018 -701 1018 -701 0 feedthrough
rlabel pdiffusion 1025 -701 1025 -701 0 feedthrough
rlabel pdiffusion 1032 -701 1032 -701 0 feedthrough
rlabel pdiffusion 1039 -701 1039 -701 0 feedthrough
rlabel pdiffusion 1046 -701 1046 -701 0 feedthrough
rlabel pdiffusion 1053 -701 1053 -701 0 feedthrough
rlabel pdiffusion 1060 -701 1060 -701 0 feedthrough
rlabel pdiffusion 1067 -701 1067 -701 0 feedthrough
rlabel pdiffusion 1074 -701 1074 -701 0 feedthrough
rlabel pdiffusion 1081 -701 1081 -701 0 cellNo=380
rlabel pdiffusion 1088 -701 1088 -701 0 feedthrough
rlabel pdiffusion 1095 -701 1095 -701 0 feedthrough
rlabel pdiffusion 1102 -701 1102 -701 0 feedthrough
rlabel pdiffusion 1109 -701 1109 -701 0 cellNo=585
rlabel pdiffusion 1116 -701 1116 -701 0 feedthrough
rlabel pdiffusion 1123 -701 1123 -701 0 feedthrough
rlabel pdiffusion 1130 -701 1130 -701 0 feedthrough
rlabel pdiffusion 1137 -701 1137 -701 0 cellNo=656
rlabel pdiffusion 1144 -701 1144 -701 0 feedthrough
rlabel pdiffusion 1151 -701 1151 -701 0 feedthrough
rlabel pdiffusion 1158 -701 1158 -701 0 feedthrough
rlabel pdiffusion 24 -778 24 -778 0 feedthrough
rlabel pdiffusion 31 -778 31 -778 0 cellNo=472
rlabel pdiffusion 38 -778 38 -778 0 feedthrough
rlabel pdiffusion 45 -778 45 -778 0 feedthrough
rlabel pdiffusion 52 -778 52 -778 0 feedthrough
rlabel pdiffusion 59 -778 59 -778 0 feedthrough
rlabel pdiffusion 66 -778 66 -778 0 feedthrough
rlabel pdiffusion 73 -778 73 -778 0 feedthrough
rlabel pdiffusion 80 -778 80 -778 0 feedthrough
rlabel pdiffusion 87 -778 87 -778 0 cellNo=849
rlabel pdiffusion 94 -778 94 -778 0 feedthrough
rlabel pdiffusion 101 -778 101 -778 0 cellNo=85
rlabel pdiffusion 108 -778 108 -778 0 feedthrough
rlabel pdiffusion 115 -778 115 -778 0 feedthrough
rlabel pdiffusion 122 -778 122 -778 0 feedthrough
rlabel pdiffusion 129 -778 129 -778 0 feedthrough
rlabel pdiffusion 136 -778 136 -778 0 cellNo=787
rlabel pdiffusion 143 -778 143 -778 0 feedthrough
rlabel pdiffusion 150 -778 150 -778 0 cellNo=360
rlabel pdiffusion 157 -778 157 -778 0 cellNo=258
rlabel pdiffusion 164 -778 164 -778 0 feedthrough
rlabel pdiffusion 171 -778 171 -778 0 cellNo=323
rlabel pdiffusion 178 -778 178 -778 0 feedthrough
rlabel pdiffusion 185 -778 185 -778 0 feedthrough
rlabel pdiffusion 192 -778 192 -778 0 feedthrough
rlabel pdiffusion 199 -778 199 -778 0 feedthrough
rlabel pdiffusion 206 -778 206 -778 0 cellNo=980
rlabel pdiffusion 213 -778 213 -778 0 feedthrough
rlabel pdiffusion 220 -778 220 -778 0 feedthrough
rlabel pdiffusion 227 -778 227 -778 0 feedthrough
rlabel pdiffusion 234 -778 234 -778 0 feedthrough
rlabel pdiffusion 241 -778 241 -778 0 feedthrough
rlabel pdiffusion 248 -778 248 -778 0 feedthrough
rlabel pdiffusion 255 -778 255 -778 0 feedthrough
rlabel pdiffusion 262 -778 262 -778 0 feedthrough
rlabel pdiffusion 269 -778 269 -778 0 feedthrough
rlabel pdiffusion 276 -778 276 -778 0 feedthrough
rlabel pdiffusion 283 -778 283 -778 0 feedthrough
rlabel pdiffusion 290 -778 290 -778 0 cellNo=605
rlabel pdiffusion 297 -778 297 -778 0 feedthrough
rlabel pdiffusion 304 -778 304 -778 0 feedthrough
rlabel pdiffusion 311 -778 311 -778 0 cellNo=280
rlabel pdiffusion 318 -778 318 -778 0 feedthrough
rlabel pdiffusion 325 -778 325 -778 0 cellNo=266
rlabel pdiffusion 332 -778 332 -778 0 feedthrough
rlabel pdiffusion 339 -778 339 -778 0 feedthrough
rlabel pdiffusion 346 -778 346 -778 0 feedthrough
rlabel pdiffusion 353 -778 353 -778 0 feedthrough
rlabel pdiffusion 360 -778 360 -778 0 feedthrough
rlabel pdiffusion 367 -778 367 -778 0 cellNo=987
rlabel pdiffusion 374 -778 374 -778 0 feedthrough
rlabel pdiffusion 381 -778 381 -778 0 feedthrough
rlabel pdiffusion 388 -778 388 -778 0 feedthrough
rlabel pdiffusion 395 -778 395 -778 0 feedthrough
rlabel pdiffusion 402 -778 402 -778 0 feedthrough
rlabel pdiffusion 409 -778 409 -778 0 feedthrough
rlabel pdiffusion 416 -778 416 -778 0 feedthrough
rlabel pdiffusion 423 -778 423 -778 0 feedthrough
rlabel pdiffusion 430 -778 430 -778 0 feedthrough
rlabel pdiffusion 437 -778 437 -778 0 feedthrough
rlabel pdiffusion 444 -778 444 -778 0 cellNo=373
rlabel pdiffusion 451 -778 451 -778 0 feedthrough
rlabel pdiffusion 458 -778 458 -778 0 cellNo=798
rlabel pdiffusion 465 -778 465 -778 0 cellNo=586
rlabel pdiffusion 472 -778 472 -778 0 feedthrough
rlabel pdiffusion 479 -778 479 -778 0 feedthrough
rlabel pdiffusion 486 -778 486 -778 0 feedthrough
rlabel pdiffusion 493 -778 493 -778 0 cellNo=963
rlabel pdiffusion 500 -778 500 -778 0 feedthrough
rlabel pdiffusion 507 -778 507 -778 0 feedthrough
rlabel pdiffusion 514 -778 514 -778 0 feedthrough
rlabel pdiffusion 521 -778 521 -778 0 feedthrough
rlabel pdiffusion 528 -778 528 -778 0 cellNo=465
rlabel pdiffusion 535 -778 535 -778 0 cellNo=628
rlabel pdiffusion 542 -778 542 -778 0 feedthrough
rlabel pdiffusion 549 -778 549 -778 0 feedthrough
rlabel pdiffusion 556 -778 556 -778 0 feedthrough
rlabel pdiffusion 563 -778 563 -778 0 feedthrough
rlabel pdiffusion 570 -778 570 -778 0 feedthrough
rlabel pdiffusion 577 -778 577 -778 0 feedthrough
rlabel pdiffusion 584 -778 584 -778 0 feedthrough
rlabel pdiffusion 591 -778 591 -778 0 feedthrough
rlabel pdiffusion 598 -778 598 -778 0 feedthrough
rlabel pdiffusion 605 -778 605 -778 0 feedthrough
rlabel pdiffusion 612 -778 612 -778 0 feedthrough
rlabel pdiffusion 619 -778 619 -778 0 cellNo=687
rlabel pdiffusion 626 -778 626 -778 0 feedthrough
rlabel pdiffusion 633 -778 633 -778 0 feedthrough
rlabel pdiffusion 640 -778 640 -778 0 feedthrough
rlabel pdiffusion 647 -778 647 -778 0 feedthrough
rlabel pdiffusion 654 -778 654 -778 0 cellNo=645
rlabel pdiffusion 661 -778 661 -778 0 cellNo=502
rlabel pdiffusion 668 -778 668 -778 0 feedthrough
rlabel pdiffusion 675 -778 675 -778 0 feedthrough
rlabel pdiffusion 682 -778 682 -778 0 feedthrough
rlabel pdiffusion 689 -778 689 -778 0 feedthrough
rlabel pdiffusion 696 -778 696 -778 0 feedthrough
rlabel pdiffusion 703 -778 703 -778 0 cellNo=17
rlabel pdiffusion 710 -778 710 -778 0 feedthrough
rlabel pdiffusion 717 -778 717 -778 0 cellNo=403
rlabel pdiffusion 724 -778 724 -778 0 feedthrough
rlabel pdiffusion 731 -778 731 -778 0 feedthrough
rlabel pdiffusion 738 -778 738 -778 0 feedthrough
rlabel pdiffusion 745 -778 745 -778 0 feedthrough
rlabel pdiffusion 752 -778 752 -778 0 feedthrough
rlabel pdiffusion 759 -778 759 -778 0 cellNo=21
rlabel pdiffusion 766 -778 766 -778 0 feedthrough
rlabel pdiffusion 773 -778 773 -778 0 cellNo=756
rlabel pdiffusion 780 -778 780 -778 0 feedthrough
rlabel pdiffusion 787 -778 787 -778 0 feedthrough
rlabel pdiffusion 794 -778 794 -778 0 cellNo=447
rlabel pdiffusion 801 -778 801 -778 0 feedthrough
rlabel pdiffusion 808 -778 808 -778 0 feedthrough
rlabel pdiffusion 815 -778 815 -778 0 feedthrough
rlabel pdiffusion 822 -778 822 -778 0 feedthrough
rlabel pdiffusion 829 -778 829 -778 0 feedthrough
rlabel pdiffusion 836 -778 836 -778 0 feedthrough
rlabel pdiffusion 843 -778 843 -778 0 feedthrough
rlabel pdiffusion 850 -778 850 -778 0 feedthrough
rlabel pdiffusion 857 -778 857 -778 0 feedthrough
rlabel pdiffusion 864 -778 864 -778 0 feedthrough
rlabel pdiffusion 871 -778 871 -778 0 feedthrough
rlabel pdiffusion 878 -778 878 -778 0 cellNo=168
rlabel pdiffusion 885 -778 885 -778 0 feedthrough
rlabel pdiffusion 892 -778 892 -778 0 feedthrough
rlabel pdiffusion 899 -778 899 -778 0 feedthrough
rlabel pdiffusion 906 -778 906 -778 0 feedthrough
rlabel pdiffusion 913 -778 913 -778 0 feedthrough
rlabel pdiffusion 920 -778 920 -778 0 feedthrough
rlabel pdiffusion 927 -778 927 -778 0 feedthrough
rlabel pdiffusion 934 -778 934 -778 0 cellNo=20
rlabel pdiffusion 941 -778 941 -778 0 cellNo=419
rlabel pdiffusion 948 -778 948 -778 0 cellNo=170
rlabel pdiffusion 955 -778 955 -778 0 cellNo=297
rlabel pdiffusion 962 -778 962 -778 0 feedthrough
rlabel pdiffusion 969 -778 969 -778 0 feedthrough
rlabel pdiffusion 976 -778 976 -778 0 feedthrough
rlabel pdiffusion 983 -778 983 -778 0 feedthrough
rlabel pdiffusion 990 -778 990 -778 0 feedthrough
rlabel pdiffusion 997 -778 997 -778 0 feedthrough
rlabel pdiffusion 1004 -778 1004 -778 0 feedthrough
rlabel pdiffusion 1011 -778 1011 -778 0 cellNo=423
rlabel pdiffusion 1032 -778 1032 -778 0 feedthrough
rlabel pdiffusion 1123 -778 1123 -778 0 feedthrough
rlabel pdiffusion 3 -865 3 -865 0 feedthrough
rlabel pdiffusion 10 -865 10 -865 0 cellNo=68
rlabel pdiffusion 17 -865 17 -865 0 feedthrough
rlabel pdiffusion 24 -865 24 -865 0 feedthrough
rlabel pdiffusion 31 -865 31 -865 0 feedthrough
rlabel pdiffusion 38 -865 38 -865 0 cellNo=174
rlabel pdiffusion 45 -865 45 -865 0 feedthrough
rlabel pdiffusion 52 -865 52 -865 0 feedthrough
rlabel pdiffusion 59 -865 59 -865 0 feedthrough
rlabel pdiffusion 66 -865 66 -865 0 feedthrough
rlabel pdiffusion 73 -865 73 -865 0 cellNo=653
rlabel pdiffusion 80 -865 80 -865 0 cellNo=831
rlabel pdiffusion 87 -865 87 -865 0 feedthrough
rlabel pdiffusion 94 -865 94 -865 0 feedthrough
rlabel pdiffusion 101 -865 101 -865 0 feedthrough
rlabel pdiffusion 108 -865 108 -865 0 feedthrough
rlabel pdiffusion 115 -865 115 -865 0 feedthrough
rlabel pdiffusion 122 -865 122 -865 0 feedthrough
rlabel pdiffusion 129 -865 129 -865 0 feedthrough
rlabel pdiffusion 136 -865 136 -865 0 feedthrough
rlabel pdiffusion 143 -865 143 -865 0 feedthrough
rlabel pdiffusion 150 -865 150 -865 0 feedthrough
rlabel pdiffusion 157 -865 157 -865 0 feedthrough
rlabel pdiffusion 164 -865 164 -865 0 feedthrough
rlabel pdiffusion 171 -865 171 -865 0 feedthrough
rlabel pdiffusion 178 -865 178 -865 0 feedthrough
rlabel pdiffusion 185 -865 185 -865 0 feedthrough
rlabel pdiffusion 192 -865 192 -865 0 cellNo=874
rlabel pdiffusion 199 -865 199 -865 0 feedthrough
rlabel pdiffusion 206 -865 206 -865 0 feedthrough
rlabel pdiffusion 213 -865 213 -865 0 feedthrough
rlabel pdiffusion 220 -865 220 -865 0 cellNo=700
rlabel pdiffusion 227 -865 227 -865 0 cellNo=714
rlabel pdiffusion 234 -865 234 -865 0 feedthrough
rlabel pdiffusion 241 -865 241 -865 0 feedthrough
rlabel pdiffusion 248 -865 248 -865 0 feedthrough
rlabel pdiffusion 255 -865 255 -865 0 feedthrough
rlabel pdiffusion 262 -865 262 -865 0 cellNo=116
rlabel pdiffusion 269 -865 269 -865 0 feedthrough
rlabel pdiffusion 276 -865 276 -865 0 feedthrough
rlabel pdiffusion 283 -865 283 -865 0 feedthrough
rlabel pdiffusion 290 -865 290 -865 0 feedthrough
rlabel pdiffusion 297 -865 297 -865 0 feedthrough
rlabel pdiffusion 304 -865 304 -865 0 feedthrough
rlabel pdiffusion 311 -865 311 -865 0 feedthrough
rlabel pdiffusion 318 -865 318 -865 0 feedthrough
rlabel pdiffusion 325 -865 325 -865 0 cellNo=140
rlabel pdiffusion 332 -865 332 -865 0 feedthrough
rlabel pdiffusion 339 -865 339 -865 0 cellNo=362
rlabel pdiffusion 346 -865 346 -865 0 feedthrough
rlabel pdiffusion 353 -865 353 -865 0 cellNo=858
rlabel pdiffusion 360 -865 360 -865 0 feedthrough
rlabel pdiffusion 367 -865 367 -865 0 feedthrough
rlabel pdiffusion 374 -865 374 -865 0 feedthrough
rlabel pdiffusion 381 -865 381 -865 0 cellNo=371
rlabel pdiffusion 388 -865 388 -865 0 feedthrough
rlabel pdiffusion 395 -865 395 -865 0 cellNo=117
rlabel pdiffusion 402 -865 402 -865 0 feedthrough
rlabel pdiffusion 409 -865 409 -865 0 feedthrough
rlabel pdiffusion 416 -865 416 -865 0 feedthrough
rlabel pdiffusion 423 -865 423 -865 0 feedthrough
rlabel pdiffusion 430 -865 430 -865 0 cellNo=478
rlabel pdiffusion 437 -865 437 -865 0 feedthrough
rlabel pdiffusion 444 -865 444 -865 0 feedthrough
rlabel pdiffusion 451 -865 451 -865 0 cellNo=594
rlabel pdiffusion 458 -865 458 -865 0 feedthrough
rlabel pdiffusion 465 -865 465 -865 0 feedthrough
rlabel pdiffusion 472 -865 472 -865 0 feedthrough
rlabel pdiffusion 479 -865 479 -865 0 cellNo=193
rlabel pdiffusion 486 -865 486 -865 0 feedthrough
rlabel pdiffusion 493 -865 493 -865 0 feedthrough
rlabel pdiffusion 500 -865 500 -865 0 cellNo=730
rlabel pdiffusion 507 -865 507 -865 0 feedthrough
rlabel pdiffusion 514 -865 514 -865 0 feedthrough
rlabel pdiffusion 521 -865 521 -865 0 feedthrough
rlabel pdiffusion 528 -865 528 -865 0 feedthrough
rlabel pdiffusion 535 -865 535 -865 0 feedthrough
rlabel pdiffusion 542 -865 542 -865 0 cellNo=427
rlabel pdiffusion 549 -865 549 -865 0 feedthrough
rlabel pdiffusion 556 -865 556 -865 0 cellNo=12
rlabel pdiffusion 563 -865 563 -865 0 cellNo=613
rlabel pdiffusion 570 -865 570 -865 0 feedthrough
rlabel pdiffusion 577 -865 577 -865 0 cellNo=208
rlabel pdiffusion 584 -865 584 -865 0 feedthrough
rlabel pdiffusion 591 -865 591 -865 0 cellNo=52
rlabel pdiffusion 598 -865 598 -865 0 feedthrough
rlabel pdiffusion 605 -865 605 -865 0 cellNo=666
rlabel pdiffusion 612 -865 612 -865 0 cellNo=621
rlabel pdiffusion 619 -865 619 -865 0 feedthrough
rlabel pdiffusion 626 -865 626 -865 0 feedthrough
rlabel pdiffusion 633 -865 633 -865 0 cellNo=342
rlabel pdiffusion 640 -865 640 -865 0 feedthrough
rlabel pdiffusion 647 -865 647 -865 0 feedthrough
rlabel pdiffusion 654 -865 654 -865 0 cellNo=777
rlabel pdiffusion 661 -865 661 -865 0 feedthrough
rlabel pdiffusion 668 -865 668 -865 0 feedthrough
rlabel pdiffusion 675 -865 675 -865 0 feedthrough
rlabel pdiffusion 682 -865 682 -865 0 feedthrough
rlabel pdiffusion 689 -865 689 -865 0 feedthrough
rlabel pdiffusion 696 -865 696 -865 0 feedthrough
rlabel pdiffusion 703 -865 703 -865 0 feedthrough
rlabel pdiffusion 710 -865 710 -865 0 feedthrough
rlabel pdiffusion 717 -865 717 -865 0 feedthrough
rlabel pdiffusion 724 -865 724 -865 0 feedthrough
rlabel pdiffusion 731 -865 731 -865 0 feedthrough
rlabel pdiffusion 738 -865 738 -865 0 feedthrough
rlabel pdiffusion 745 -865 745 -865 0 feedthrough
rlabel pdiffusion 752 -865 752 -865 0 feedthrough
rlabel pdiffusion 759 -865 759 -865 0 feedthrough
rlabel pdiffusion 766 -865 766 -865 0 cellNo=252
rlabel pdiffusion 773 -865 773 -865 0 feedthrough
rlabel pdiffusion 780 -865 780 -865 0 feedthrough
rlabel pdiffusion 787 -865 787 -865 0 feedthrough
rlabel pdiffusion 794 -865 794 -865 0 feedthrough
rlabel pdiffusion 801 -865 801 -865 0 feedthrough
rlabel pdiffusion 808 -865 808 -865 0 feedthrough
rlabel pdiffusion 815 -865 815 -865 0 feedthrough
rlabel pdiffusion 822 -865 822 -865 0 feedthrough
rlabel pdiffusion 829 -865 829 -865 0 feedthrough
rlabel pdiffusion 836 -865 836 -865 0 feedthrough
rlabel pdiffusion 843 -865 843 -865 0 feedthrough
rlabel pdiffusion 850 -865 850 -865 0 feedthrough
rlabel pdiffusion 857 -865 857 -865 0 feedthrough
rlabel pdiffusion 864 -865 864 -865 0 cellNo=663
rlabel pdiffusion 871 -865 871 -865 0 feedthrough
rlabel pdiffusion 878 -865 878 -865 0 feedthrough
rlabel pdiffusion 885 -865 885 -865 0 feedthrough
rlabel pdiffusion 892 -865 892 -865 0 feedthrough
rlabel pdiffusion 899 -865 899 -865 0 feedthrough
rlabel pdiffusion 906 -865 906 -865 0 feedthrough
rlabel pdiffusion 913 -865 913 -865 0 feedthrough
rlabel pdiffusion 920 -865 920 -865 0 feedthrough
rlabel pdiffusion 927 -865 927 -865 0 feedthrough
rlabel pdiffusion 934 -865 934 -865 0 feedthrough
rlabel pdiffusion 941 -865 941 -865 0 feedthrough
rlabel pdiffusion 948 -865 948 -865 0 feedthrough
rlabel pdiffusion 955 -865 955 -865 0 feedthrough
rlabel pdiffusion 962 -865 962 -865 0 feedthrough
rlabel pdiffusion 969 -865 969 -865 0 feedthrough
rlabel pdiffusion 976 -865 976 -865 0 feedthrough
rlabel pdiffusion 983 -865 983 -865 0 feedthrough
rlabel pdiffusion 990 -865 990 -865 0 feedthrough
rlabel pdiffusion 997 -865 997 -865 0 feedthrough
rlabel pdiffusion 1004 -865 1004 -865 0 feedthrough
rlabel pdiffusion 1011 -865 1011 -865 0 feedthrough
rlabel pdiffusion 1018 -865 1018 -865 0 feedthrough
rlabel pdiffusion 1025 -865 1025 -865 0 feedthrough
rlabel pdiffusion 1032 -865 1032 -865 0 feedthrough
rlabel pdiffusion 1039 -865 1039 -865 0 feedthrough
rlabel pdiffusion 1046 -865 1046 -865 0 feedthrough
rlabel pdiffusion 1053 -865 1053 -865 0 feedthrough
rlabel pdiffusion 1060 -865 1060 -865 0 feedthrough
rlabel pdiffusion 1067 -865 1067 -865 0 feedthrough
rlabel pdiffusion 1074 -865 1074 -865 0 feedthrough
rlabel pdiffusion 1081 -865 1081 -865 0 feedthrough
rlabel pdiffusion 1088 -865 1088 -865 0 feedthrough
rlabel pdiffusion 1095 -865 1095 -865 0 cellNo=799
rlabel pdiffusion 1102 -865 1102 -865 0 feedthrough
rlabel pdiffusion 1109 -865 1109 -865 0 feedthrough
rlabel pdiffusion 1116 -865 1116 -865 0 feedthrough
rlabel pdiffusion 1123 -865 1123 -865 0 feedthrough
rlabel pdiffusion 1130 -865 1130 -865 0 cellNo=408
rlabel pdiffusion 1137 -865 1137 -865 0 cellNo=532
rlabel pdiffusion 1144 -865 1144 -865 0 feedthrough
rlabel pdiffusion 1151 -865 1151 -865 0 cellNo=521
rlabel pdiffusion 3 -966 3 -966 0 cellNo=494
rlabel pdiffusion 10 -966 10 -966 0 feedthrough
rlabel pdiffusion 17 -966 17 -966 0 cellNo=626
rlabel pdiffusion 24 -966 24 -966 0 feedthrough
rlabel pdiffusion 31 -966 31 -966 0 cellNo=47
rlabel pdiffusion 38 -966 38 -966 0 cellNo=163
rlabel pdiffusion 45 -966 45 -966 0 feedthrough
rlabel pdiffusion 52 -966 52 -966 0 feedthrough
rlabel pdiffusion 59 -966 59 -966 0 feedthrough
rlabel pdiffusion 66 -966 66 -966 0 cellNo=164
rlabel pdiffusion 73 -966 73 -966 0 cellNo=404
rlabel pdiffusion 80 -966 80 -966 0 cellNo=961
rlabel pdiffusion 87 -966 87 -966 0 feedthrough
rlabel pdiffusion 94 -966 94 -966 0 feedthrough
rlabel pdiffusion 101 -966 101 -966 0 feedthrough
rlabel pdiffusion 108 -966 108 -966 0 feedthrough
rlabel pdiffusion 115 -966 115 -966 0 feedthrough
rlabel pdiffusion 122 -966 122 -966 0 feedthrough
rlabel pdiffusion 129 -966 129 -966 0 feedthrough
rlabel pdiffusion 136 -966 136 -966 0 feedthrough
rlabel pdiffusion 143 -966 143 -966 0 feedthrough
rlabel pdiffusion 150 -966 150 -966 0 cellNo=431
rlabel pdiffusion 157 -966 157 -966 0 feedthrough
rlabel pdiffusion 164 -966 164 -966 0 feedthrough
rlabel pdiffusion 171 -966 171 -966 0 feedthrough
rlabel pdiffusion 178 -966 178 -966 0 feedthrough
rlabel pdiffusion 185 -966 185 -966 0 feedthrough
rlabel pdiffusion 192 -966 192 -966 0 feedthrough
rlabel pdiffusion 199 -966 199 -966 0 feedthrough
rlabel pdiffusion 206 -966 206 -966 0 feedthrough
rlabel pdiffusion 213 -966 213 -966 0 feedthrough
rlabel pdiffusion 220 -966 220 -966 0 feedthrough
rlabel pdiffusion 227 -966 227 -966 0 feedthrough
rlabel pdiffusion 234 -966 234 -966 0 feedthrough
rlabel pdiffusion 241 -966 241 -966 0 feedthrough
rlabel pdiffusion 248 -966 248 -966 0 feedthrough
rlabel pdiffusion 255 -966 255 -966 0 feedthrough
rlabel pdiffusion 262 -966 262 -966 0 feedthrough
rlabel pdiffusion 269 -966 269 -966 0 feedthrough
rlabel pdiffusion 276 -966 276 -966 0 feedthrough
rlabel pdiffusion 283 -966 283 -966 0 cellNo=976
rlabel pdiffusion 290 -966 290 -966 0 feedthrough
rlabel pdiffusion 297 -966 297 -966 0 cellNo=606
rlabel pdiffusion 304 -966 304 -966 0 cellNo=750
rlabel pdiffusion 311 -966 311 -966 0 feedthrough
rlabel pdiffusion 318 -966 318 -966 0 feedthrough
rlabel pdiffusion 325 -966 325 -966 0 feedthrough
rlabel pdiffusion 332 -966 332 -966 0 feedthrough
rlabel pdiffusion 339 -966 339 -966 0 feedthrough
rlabel pdiffusion 346 -966 346 -966 0 feedthrough
rlabel pdiffusion 353 -966 353 -966 0 feedthrough
rlabel pdiffusion 360 -966 360 -966 0 cellNo=54
rlabel pdiffusion 367 -966 367 -966 0 feedthrough
rlabel pdiffusion 374 -966 374 -966 0 feedthrough
rlabel pdiffusion 381 -966 381 -966 0 feedthrough
rlabel pdiffusion 388 -966 388 -966 0 feedthrough
rlabel pdiffusion 395 -966 395 -966 0 feedthrough
rlabel pdiffusion 402 -966 402 -966 0 feedthrough
rlabel pdiffusion 409 -966 409 -966 0 feedthrough
rlabel pdiffusion 416 -966 416 -966 0 cellNo=550
rlabel pdiffusion 423 -966 423 -966 0 feedthrough
rlabel pdiffusion 430 -966 430 -966 0 feedthrough
rlabel pdiffusion 437 -966 437 -966 0 cellNo=374
rlabel pdiffusion 444 -966 444 -966 0 cellNo=872
rlabel pdiffusion 451 -966 451 -966 0 feedthrough
rlabel pdiffusion 458 -966 458 -966 0 feedthrough
rlabel pdiffusion 465 -966 465 -966 0 cellNo=508
rlabel pdiffusion 472 -966 472 -966 0 cellNo=432
rlabel pdiffusion 479 -966 479 -966 0 cellNo=274
rlabel pdiffusion 486 -966 486 -966 0 feedthrough
rlabel pdiffusion 493 -966 493 -966 0 feedthrough
rlabel pdiffusion 500 -966 500 -966 0 cellNo=112
rlabel pdiffusion 507 -966 507 -966 0 cellNo=487
rlabel pdiffusion 514 -966 514 -966 0 feedthrough
rlabel pdiffusion 521 -966 521 -966 0 feedthrough
rlabel pdiffusion 528 -966 528 -966 0 feedthrough
rlabel pdiffusion 535 -966 535 -966 0 cellNo=157
rlabel pdiffusion 542 -966 542 -966 0 cellNo=589
rlabel pdiffusion 549 -966 549 -966 0 feedthrough
rlabel pdiffusion 556 -966 556 -966 0 feedthrough
rlabel pdiffusion 563 -966 563 -966 0 feedthrough
rlabel pdiffusion 570 -966 570 -966 0 cellNo=848
rlabel pdiffusion 577 -966 577 -966 0 cellNo=572
rlabel pdiffusion 584 -966 584 -966 0 feedthrough
rlabel pdiffusion 591 -966 591 -966 0 cellNo=525
rlabel pdiffusion 598 -966 598 -966 0 feedthrough
rlabel pdiffusion 605 -966 605 -966 0 feedthrough
rlabel pdiffusion 612 -966 612 -966 0 cellNo=202
rlabel pdiffusion 619 -966 619 -966 0 cellNo=673
rlabel pdiffusion 626 -966 626 -966 0 cellNo=185
rlabel pdiffusion 633 -966 633 -966 0 cellNo=712
rlabel pdiffusion 640 -966 640 -966 0 feedthrough
rlabel pdiffusion 647 -966 647 -966 0 feedthrough
rlabel pdiffusion 654 -966 654 -966 0 feedthrough
rlabel pdiffusion 661 -966 661 -966 0 feedthrough
rlabel pdiffusion 668 -966 668 -966 0 feedthrough
rlabel pdiffusion 675 -966 675 -966 0 feedthrough
rlabel pdiffusion 682 -966 682 -966 0 feedthrough
rlabel pdiffusion 689 -966 689 -966 0 cellNo=215
rlabel pdiffusion 696 -966 696 -966 0 cellNo=467
rlabel pdiffusion 703 -966 703 -966 0 feedthrough
rlabel pdiffusion 710 -966 710 -966 0 feedthrough
rlabel pdiffusion 717 -966 717 -966 0 feedthrough
rlabel pdiffusion 724 -966 724 -966 0 feedthrough
rlabel pdiffusion 731 -966 731 -966 0 feedthrough
rlabel pdiffusion 738 -966 738 -966 0 feedthrough
rlabel pdiffusion 745 -966 745 -966 0 feedthrough
rlabel pdiffusion 752 -966 752 -966 0 feedthrough
rlabel pdiffusion 759 -966 759 -966 0 feedthrough
rlabel pdiffusion 766 -966 766 -966 0 feedthrough
rlabel pdiffusion 773 -966 773 -966 0 feedthrough
rlabel pdiffusion 780 -966 780 -966 0 feedthrough
rlabel pdiffusion 787 -966 787 -966 0 feedthrough
rlabel pdiffusion 794 -966 794 -966 0 feedthrough
rlabel pdiffusion 801 -966 801 -966 0 feedthrough
rlabel pdiffusion 808 -966 808 -966 0 feedthrough
rlabel pdiffusion 815 -966 815 -966 0 feedthrough
rlabel pdiffusion 822 -966 822 -966 0 feedthrough
rlabel pdiffusion 829 -966 829 -966 0 feedthrough
rlabel pdiffusion 836 -966 836 -966 0 feedthrough
rlabel pdiffusion 843 -966 843 -966 0 feedthrough
rlabel pdiffusion 850 -966 850 -966 0 feedthrough
rlabel pdiffusion 857 -966 857 -966 0 cellNo=91
rlabel pdiffusion 864 -966 864 -966 0 feedthrough
rlabel pdiffusion 871 -966 871 -966 0 feedthrough
rlabel pdiffusion 878 -966 878 -966 0 feedthrough
rlabel pdiffusion 885 -966 885 -966 0 feedthrough
rlabel pdiffusion 892 -966 892 -966 0 feedthrough
rlabel pdiffusion 899 -966 899 -966 0 feedthrough
rlabel pdiffusion 906 -966 906 -966 0 feedthrough
rlabel pdiffusion 913 -966 913 -966 0 feedthrough
rlabel pdiffusion 920 -966 920 -966 0 feedthrough
rlabel pdiffusion 927 -966 927 -966 0 feedthrough
rlabel pdiffusion 934 -966 934 -966 0 feedthrough
rlabel pdiffusion 941 -966 941 -966 0 feedthrough
rlabel pdiffusion 948 -966 948 -966 0 feedthrough
rlabel pdiffusion 955 -966 955 -966 0 feedthrough
rlabel pdiffusion 962 -966 962 -966 0 feedthrough
rlabel pdiffusion 969 -966 969 -966 0 feedthrough
rlabel pdiffusion 976 -966 976 -966 0 feedthrough
rlabel pdiffusion 983 -966 983 -966 0 feedthrough
rlabel pdiffusion 990 -966 990 -966 0 feedthrough
rlabel pdiffusion 997 -966 997 -966 0 feedthrough
rlabel pdiffusion 1004 -966 1004 -966 0 feedthrough
rlabel pdiffusion 1011 -966 1011 -966 0 feedthrough
rlabel pdiffusion 1018 -966 1018 -966 0 feedthrough
rlabel pdiffusion 1025 -966 1025 -966 0 feedthrough
rlabel pdiffusion 1032 -966 1032 -966 0 feedthrough
rlabel pdiffusion 1039 -966 1039 -966 0 feedthrough
rlabel pdiffusion 1046 -966 1046 -966 0 feedthrough
rlabel pdiffusion 1053 -966 1053 -966 0 feedthrough
rlabel pdiffusion 1060 -966 1060 -966 0 feedthrough
rlabel pdiffusion 1067 -966 1067 -966 0 feedthrough
rlabel pdiffusion 1074 -966 1074 -966 0 feedthrough
rlabel pdiffusion 1081 -966 1081 -966 0 feedthrough
rlabel pdiffusion 1088 -966 1088 -966 0 feedthrough
rlabel pdiffusion 1095 -966 1095 -966 0 feedthrough
rlabel pdiffusion 1102 -966 1102 -966 0 feedthrough
rlabel pdiffusion 1109 -966 1109 -966 0 feedthrough
rlabel pdiffusion 1116 -966 1116 -966 0 feedthrough
rlabel pdiffusion 1123 -966 1123 -966 0 feedthrough
rlabel pdiffusion 1130 -966 1130 -966 0 feedthrough
rlabel pdiffusion 1137 -966 1137 -966 0 feedthrough
rlabel pdiffusion 1144 -966 1144 -966 0 feedthrough
rlabel pdiffusion 1151 -966 1151 -966 0 feedthrough
rlabel pdiffusion 1158 -966 1158 -966 0 feedthrough
rlabel pdiffusion 3 -1081 3 -1081 0 cellNo=209
rlabel pdiffusion 10 -1081 10 -1081 0 feedthrough
rlabel pdiffusion 17 -1081 17 -1081 0 feedthrough
rlabel pdiffusion 24 -1081 24 -1081 0 feedthrough
rlabel pdiffusion 31 -1081 31 -1081 0 feedthrough
rlabel pdiffusion 38 -1081 38 -1081 0 feedthrough
rlabel pdiffusion 45 -1081 45 -1081 0 feedthrough
rlabel pdiffusion 52 -1081 52 -1081 0 cellNo=381
rlabel pdiffusion 59 -1081 59 -1081 0 feedthrough
rlabel pdiffusion 66 -1081 66 -1081 0 cellNo=311
rlabel pdiffusion 73 -1081 73 -1081 0 feedthrough
rlabel pdiffusion 80 -1081 80 -1081 0 cellNo=292
rlabel pdiffusion 87 -1081 87 -1081 0 feedthrough
rlabel pdiffusion 94 -1081 94 -1081 0 feedthrough
rlabel pdiffusion 101 -1081 101 -1081 0 cellNo=723
rlabel pdiffusion 108 -1081 108 -1081 0 cellNo=411
rlabel pdiffusion 115 -1081 115 -1081 0 feedthrough
rlabel pdiffusion 122 -1081 122 -1081 0 feedthrough
rlabel pdiffusion 129 -1081 129 -1081 0 feedthrough
rlabel pdiffusion 136 -1081 136 -1081 0 feedthrough
rlabel pdiffusion 143 -1081 143 -1081 0 feedthrough
rlabel pdiffusion 150 -1081 150 -1081 0 feedthrough
rlabel pdiffusion 157 -1081 157 -1081 0 feedthrough
rlabel pdiffusion 164 -1081 164 -1081 0 cellNo=598
rlabel pdiffusion 171 -1081 171 -1081 0 feedthrough
rlabel pdiffusion 178 -1081 178 -1081 0 feedthrough
rlabel pdiffusion 185 -1081 185 -1081 0 feedthrough
rlabel pdiffusion 192 -1081 192 -1081 0 cellNo=884
rlabel pdiffusion 199 -1081 199 -1081 0 cellNo=886
rlabel pdiffusion 206 -1081 206 -1081 0 feedthrough
rlabel pdiffusion 213 -1081 213 -1081 0 cellNo=989
rlabel pdiffusion 220 -1081 220 -1081 0 feedthrough
rlabel pdiffusion 227 -1081 227 -1081 0 cellNo=438
rlabel pdiffusion 234 -1081 234 -1081 0 feedthrough
rlabel pdiffusion 241 -1081 241 -1081 0 feedthrough
rlabel pdiffusion 248 -1081 248 -1081 0 feedthrough
rlabel pdiffusion 255 -1081 255 -1081 0 feedthrough
rlabel pdiffusion 262 -1081 262 -1081 0 feedthrough
rlabel pdiffusion 269 -1081 269 -1081 0 cellNo=684
rlabel pdiffusion 276 -1081 276 -1081 0 feedthrough
rlabel pdiffusion 283 -1081 283 -1081 0 cellNo=811
rlabel pdiffusion 290 -1081 290 -1081 0 feedthrough
rlabel pdiffusion 297 -1081 297 -1081 0 feedthrough
rlabel pdiffusion 304 -1081 304 -1081 0 feedthrough
rlabel pdiffusion 311 -1081 311 -1081 0 feedthrough
rlabel pdiffusion 318 -1081 318 -1081 0 feedthrough
rlabel pdiffusion 325 -1081 325 -1081 0 cellNo=356
rlabel pdiffusion 332 -1081 332 -1081 0 feedthrough
rlabel pdiffusion 339 -1081 339 -1081 0 feedthrough
rlabel pdiffusion 346 -1081 346 -1081 0 feedthrough
rlabel pdiffusion 353 -1081 353 -1081 0 feedthrough
rlabel pdiffusion 360 -1081 360 -1081 0 feedthrough
rlabel pdiffusion 367 -1081 367 -1081 0 feedthrough
rlabel pdiffusion 374 -1081 374 -1081 0 feedthrough
rlabel pdiffusion 381 -1081 381 -1081 0 feedthrough
rlabel pdiffusion 388 -1081 388 -1081 0 cellNo=826
rlabel pdiffusion 395 -1081 395 -1081 0 cellNo=526
rlabel pdiffusion 402 -1081 402 -1081 0 feedthrough
rlabel pdiffusion 409 -1081 409 -1081 0 feedthrough
rlabel pdiffusion 416 -1081 416 -1081 0 feedthrough
rlabel pdiffusion 423 -1081 423 -1081 0 feedthrough
rlabel pdiffusion 430 -1081 430 -1081 0 feedthrough
rlabel pdiffusion 437 -1081 437 -1081 0 feedthrough
rlabel pdiffusion 444 -1081 444 -1081 0 feedthrough
rlabel pdiffusion 451 -1081 451 -1081 0 feedthrough
rlabel pdiffusion 458 -1081 458 -1081 0 feedthrough
rlabel pdiffusion 465 -1081 465 -1081 0 feedthrough
rlabel pdiffusion 472 -1081 472 -1081 0 feedthrough
rlabel pdiffusion 479 -1081 479 -1081 0 feedthrough
rlabel pdiffusion 486 -1081 486 -1081 0 cellNo=702
rlabel pdiffusion 493 -1081 493 -1081 0 cellNo=717
rlabel pdiffusion 500 -1081 500 -1081 0 cellNo=317
rlabel pdiffusion 507 -1081 507 -1081 0 feedthrough
rlabel pdiffusion 514 -1081 514 -1081 0 feedthrough
rlabel pdiffusion 521 -1081 521 -1081 0 feedthrough
rlabel pdiffusion 528 -1081 528 -1081 0 feedthrough
rlabel pdiffusion 535 -1081 535 -1081 0 feedthrough
rlabel pdiffusion 542 -1081 542 -1081 0 cellNo=890
rlabel pdiffusion 549 -1081 549 -1081 0 feedthrough
rlabel pdiffusion 556 -1081 556 -1081 0 cellNo=734
rlabel pdiffusion 563 -1081 563 -1081 0 feedthrough
rlabel pdiffusion 570 -1081 570 -1081 0 cellNo=41
rlabel pdiffusion 577 -1081 577 -1081 0 feedthrough
rlabel pdiffusion 584 -1081 584 -1081 0 cellNo=130
rlabel pdiffusion 591 -1081 591 -1081 0 feedthrough
rlabel pdiffusion 598 -1081 598 -1081 0 cellNo=503
rlabel pdiffusion 605 -1081 605 -1081 0 cellNo=343
rlabel pdiffusion 612 -1081 612 -1081 0 feedthrough
rlabel pdiffusion 619 -1081 619 -1081 0 feedthrough
rlabel pdiffusion 626 -1081 626 -1081 0 feedthrough
rlabel pdiffusion 633 -1081 633 -1081 0 cellNo=568
rlabel pdiffusion 640 -1081 640 -1081 0 feedthrough
rlabel pdiffusion 647 -1081 647 -1081 0 feedthrough
rlabel pdiffusion 654 -1081 654 -1081 0 feedthrough
rlabel pdiffusion 661 -1081 661 -1081 0 feedthrough
rlabel pdiffusion 668 -1081 668 -1081 0 feedthrough
rlabel pdiffusion 675 -1081 675 -1081 0 feedthrough
rlabel pdiffusion 682 -1081 682 -1081 0 cellNo=681
rlabel pdiffusion 689 -1081 689 -1081 0 feedthrough
rlabel pdiffusion 696 -1081 696 -1081 0 feedthrough
rlabel pdiffusion 703 -1081 703 -1081 0 feedthrough
rlabel pdiffusion 710 -1081 710 -1081 0 feedthrough
rlabel pdiffusion 717 -1081 717 -1081 0 feedthrough
rlabel pdiffusion 724 -1081 724 -1081 0 cellNo=36
rlabel pdiffusion 731 -1081 731 -1081 0 feedthrough
rlabel pdiffusion 738 -1081 738 -1081 0 cellNo=815
rlabel pdiffusion 745 -1081 745 -1081 0 feedthrough
rlabel pdiffusion 752 -1081 752 -1081 0 feedthrough
rlabel pdiffusion 759 -1081 759 -1081 0 feedthrough
rlabel pdiffusion 766 -1081 766 -1081 0 feedthrough
rlabel pdiffusion 773 -1081 773 -1081 0 feedthrough
rlabel pdiffusion 780 -1081 780 -1081 0 feedthrough
rlabel pdiffusion 787 -1081 787 -1081 0 feedthrough
rlabel pdiffusion 794 -1081 794 -1081 0 feedthrough
rlabel pdiffusion 801 -1081 801 -1081 0 feedthrough
rlabel pdiffusion 808 -1081 808 -1081 0 feedthrough
rlabel pdiffusion 815 -1081 815 -1081 0 cellNo=283
rlabel pdiffusion 822 -1081 822 -1081 0 feedthrough
rlabel pdiffusion 829 -1081 829 -1081 0 feedthrough
rlabel pdiffusion 836 -1081 836 -1081 0 feedthrough
rlabel pdiffusion 843 -1081 843 -1081 0 feedthrough
rlabel pdiffusion 850 -1081 850 -1081 0 feedthrough
rlabel pdiffusion 857 -1081 857 -1081 0 feedthrough
rlabel pdiffusion 864 -1081 864 -1081 0 feedthrough
rlabel pdiffusion 871 -1081 871 -1081 0 feedthrough
rlabel pdiffusion 878 -1081 878 -1081 0 feedthrough
rlabel pdiffusion 885 -1081 885 -1081 0 feedthrough
rlabel pdiffusion 892 -1081 892 -1081 0 feedthrough
rlabel pdiffusion 899 -1081 899 -1081 0 feedthrough
rlabel pdiffusion 906 -1081 906 -1081 0 feedthrough
rlabel pdiffusion 913 -1081 913 -1081 0 feedthrough
rlabel pdiffusion 920 -1081 920 -1081 0 feedthrough
rlabel pdiffusion 927 -1081 927 -1081 0 feedthrough
rlabel pdiffusion 934 -1081 934 -1081 0 feedthrough
rlabel pdiffusion 941 -1081 941 -1081 0 feedthrough
rlabel pdiffusion 948 -1081 948 -1081 0 feedthrough
rlabel pdiffusion 955 -1081 955 -1081 0 feedthrough
rlabel pdiffusion 962 -1081 962 -1081 0 feedthrough
rlabel pdiffusion 969 -1081 969 -1081 0 feedthrough
rlabel pdiffusion 976 -1081 976 -1081 0 feedthrough
rlabel pdiffusion 983 -1081 983 -1081 0 feedthrough
rlabel pdiffusion 990 -1081 990 -1081 0 feedthrough
rlabel pdiffusion 997 -1081 997 -1081 0 feedthrough
rlabel pdiffusion 1004 -1081 1004 -1081 0 feedthrough
rlabel pdiffusion 1011 -1081 1011 -1081 0 feedthrough
rlabel pdiffusion 1018 -1081 1018 -1081 0 feedthrough
rlabel pdiffusion 1025 -1081 1025 -1081 0 feedthrough
rlabel pdiffusion 1032 -1081 1032 -1081 0 feedthrough
rlabel pdiffusion 1039 -1081 1039 -1081 0 cellNo=248
rlabel pdiffusion 1046 -1081 1046 -1081 0 feedthrough
rlabel pdiffusion 1053 -1081 1053 -1081 0 feedthrough
rlabel pdiffusion 1060 -1081 1060 -1081 0 cellNo=631
rlabel pdiffusion 1067 -1081 1067 -1081 0 feedthrough
rlabel pdiffusion 1074 -1081 1074 -1081 0 feedthrough
rlabel pdiffusion 1081 -1081 1081 -1081 0 feedthrough
rlabel pdiffusion 1130 -1081 1130 -1081 0 feedthrough
rlabel pdiffusion 1144 -1081 1144 -1081 0 feedthrough
rlabel pdiffusion 3 -1170 3 -1170 0 cellNo=578
rlabel pdiffusion 10 -1170 10 -1170 0 feedthrough
rlabel pdiffusion 17 -1170 17 -1170 0 cellNo=496
rlabel pdiffusion 24 -1170 24 -1170 0 feedthrough
rlabel pdiffusion 31 -1170 31 -1170 0 feedthrough
rlabel pdiffusion 38 -1170 38 -1170 0 cellNo=263
rlabel pdiffusion 45 -1170 45 -1170 0 feedthrough
rlabel pdiffusion 52 -1170 52 -1170 0 feedthrough
rlabel pdiffusion 59 -1170 59 -1170 0 cellNo=10
rlabel pdiffusion 66 -1170 66 -1170 0 feedthrough
rlabel pdiffusion 73 -1170 73 -1170 0 feedthrough
rlabel pdiffusion 80 -1170 80 -1170 0 feedthrough
rlabel pdiffusion 87 -1170 87 -1170 0 feedthrough
rlabel pdiffusion 94 -1170 94 -1170 0 feedthrough
rlabel pdiffusion 101 -1170 101 -1170 0 cellNo=147
rlabel pdiffusion 108 -1170 108 -1170 0 feedthrough
rlabel pdiffusion 115 -1170 115 -1170 0 feedthrough
rlabel pdiffusion 122 -1170 122 -1170 0 feedthrough
rlabel pdiffusion 129 -1170 129 -1170 0 feedthrough
rlabel pdiffusion 136 -1170 136 -1170 0 feedthrough
rlabel pdiffusion 143 -1170 143 -1170 0 cellNo=26
rlabel pdiffusion 150 -1170 150 -1170 0 cellNo=90
rlabel pdiffusion 157 -1170 157 -1170 0 feedthrough
rlabel pdiffusion 164 -1170 164 -1170 0 cellNo=346
rlabel pdiffusion 171 -1170 171 -1170 0 cellNo=226
rlabel pdiffusion 178 -1170 178 -1170 0 feedthrough
rlabel pdiffusion 185 -1170 185 -1170 0 feedthrough
rlabel pdiffusion 192 -1170 192 -1170 0 feedthrough
rlabel pdiffusion 199 -1170 199 -1170 0 feedthrough
rlabel pdiffusion 206 -1170 206 -1170 0 feedthrough
rlabel pdiffusion 213 -1170 213 -1170 0 feedthrough
rlabel pdiffusion 220 -1170 220 -1170 0 cellNo=571
rlabel pdiffusion 227 -1170 227 -1170 0 feedthrough
rlabel pdiffusion 234 -1170 234 -1170 0 feedthrough
rlabel pdiffusion 241 -1170 241 -1170 0 feedthrough
rlabel pdiffusion 248 -1170 248 -1170 0 feedthrough
rlabel pdiffusion 255 -1170 255 -1170 0 feedthrough
rlabel pdiffusion 262 -1170 262 -1170 0 feedthrough
rlabel pdiffusion 269 -1170 269 -1170 0 feedthrough
rlabel pdiffusion 276 -1170 276 -1170 0 feedthrough
rlabel pdiffusion 283 -1170 283 -1170 0 cellNo=398
rlabel pdiffusion 290 -1170 290 -1170 0 feedthrough
rlabel pdiffusion 297 -1170 297 -1170 0 feedthrough
rlabel pdiffusion 304 -1170 304 -1170 0 feedthrough
rlabel pdiffusion 311 -1170 311 -1170 0 cellNo=529
rlabel pdiffusion 318 -1170 318 -1170 0 feedthrough
rlabel pdiffusion 325 -1170 325 -1170 0 feedthrough
rlabel pdiffusion 332 -1170 332 -1170 0 feedthrough
rlabel pdiffusion 339 -1170 339 -1170 0 feedthrough
rlabel pdiffusion 346 -1170 346 -1170 0 cellNo=389
rlabel pdiffusion 353 -1170 353 -1170 0 cellNo=145
rlabel pdiffusion 360 -1170 360 -1170 0 cellNo=895
rlabel pdiffusion 367 -1170 367 -1170 0 feedthrough
rlabel pdiffusion 374 -1170 374 -1170 0 feedthrough
rlabel pdiffusion 381 -1170 381 -1170 0 cellNo=337
rlabel pdiffusion 388 -1170 388 -1170 0 feedthrough
rlabel pdiffusion 395 -1170 395 -1170 0 feedthrough
rlabel pdiffusion 402 -1170 402 -1170 0 feedthrough
rlabel pdiffusion 409 -1170 409 -1170 0 cellNo=228
rlabel pdiffusion 416 -1170 416 -1170 0 cellNo=207
rlabel pdiffusion 423 -1170 423 -1170 0 feedthrough
rlabel pdiffusion 430 -1170 430 -1170 0 feedthrough
rlabel pdiffusion 437 -1170 437 -1170 0 feedthrough
rlabel pdiffusion 444 -1170 444 -1170 0 feedthrough
rlabel pdiffusion 451 -1170 451 -1170 0 feedthrough
rlabel pdiffusion 458 -1170 458 -1170 0 feedthrough
rlabel pdiffusion 465 -1170 465 -1170 0 cellNo=88
rlabel pdiffusion 472 -1170 472 -1170 0 feedthrough
rlabel pdiffusion 479 -1170 479 -1170 0 cellNo=877
rlabel pdiffusion 486 -1170 486 -1170 0 feedthrough
rlabel pdiffusion 493 -1170 493 -1170 0 feedthrough
rlabel pdiffusion 500 -1170 500 -1170 0 cellNo=87
rlabel pdiffusion 507 -1170 507 -1170 0 feedthrough
rlabel pdiffusion 514 -1170 514 -1170 0 feedthrough
rlabel pdiffusion 521 -1170 521 -1170 0 cellNo=804
rlabel pdiffusion 528 -1170 528 -1170 0 feedthrough
rlabel pdiffusion 535 -1170 535 -1170 0 feedthrough
rlabel pdiffusion 542 -1170 542 -1170 0 feedthrough
rlabel pdiffusion 549 -1170 549 -1170 0 feedthrough
rlabel pdiffusion 556 -1170 556 -1170 0 cellNo=866
rlabel pdiffusion 563 -1170 563 -1170 0 cellNo=844
rlabel pdiffusion 570 -1170 570 -1170 0 feedthrough
rlabel pdiffusion 577 -1170 577 -1170 0 feedthrough
rlabel pdiffusion 584 -1170 584 -1170 0 feedthrough
rlabel pdiffusion 591 -1170 591 -1170 0 feedthrough
rlabel pdiffusion 598 -1170 598 -1170 0 cellNo=310
rlabel pdiffusion 605 -1170 605 -1170 0 feedthrough
rlabel pdiffusion 612 -1170 612 -1170 0 feedthrough
rlabel pdiffusion 619 -1170 619 -1170 0 feedthrough
rlabel pdiffusion 626 -1170 626 -1170 0 feedthrough
rlabel pdiffusion 633 -1170 633 -1170 0 feedthrough
rlabel pdiffusion 640 -1170 640 -1170 0 feedthrough
rlabel pdiffusion 647 -1170 647 -1170 0 feedthrough
rlabel pdiffusion 654 -1170 654 -1170 0 feedthrough
rlabel pdiffusion 661 -1170 661 -1170 0 feedthrough
rlabel pdiffusion 668 -1170 668 -1170 0 feedthrough
rlabel pdiffusion 675 -1170 675 -1170 0 feedthrough
rlabel pdiffusion 682 -1170 682 -1170 0 feedthrough
rlabel pdiffusion 689 -1170 689 -1170 0 cellNo=81
rlabel pdiffusion 696 -1170 696 -1170 0 feedthrough
rlabel pdiffusion 703 -1170 703 -1170 0 feedthrough
rlabel pdiffusion 710 -1170 710 -1170 0 feedthrough
rlabel pdiffusion 717 -1170 717 -1170 0 feedthrough
rlabel pdiffusion 724 -1170 724 -1170 0 feedthrough
rlabel pdiffusion 731 -1170 731 -1170 0 cellNo=991
rlabel pdiffusion 738 -1170 738 -1170 0 cellNo=80
rlabel pdiffusion 745 -1170 745 -1170 0 feedthrough
rlabel pdiffusion 752 -1170 752 -1170 0 feedthrough
rlabel pdiffusion 759 -1170 759 -1170 0 feedthrough
rlabel pdiffusion 766 -1170 766 -1170 0 feedthrough
rlabel pdiffusion 773 -1170 773 -1170 0 feedthrough
rlabel pdiffusion 780 -1170 780 -1170 0 feedthrough
rlabel pdiffusion 787 -1170 787 -1170 0 cellNo=847
rlabel pdiffusion 794 -1170 794 -1170 0 feedthrough
rlabel pdiffusion 801 -1170 801 -1170 0 feedthrough
rlabel pdiffusion 808 -1170 808 -1170 0 feedthrough
rlabel pdiffusion 815 -1170 815 -1170 0 feedthrough
rlabel pdiffusion 822 -1170 822 -1170 0 feedthrough
rlabel pdiffusion 829 -1170 829 -1170 0 feedthrough
rlabel pdiffusion 836 -1170 836 -1170 0 feedthrough
rlabel pdiffusion 843 -1170 843 -1170 0 feedthrough
rlabel pdiffusion 850 -1170 850 -1170 0 feedthrough
rlabel pdiffusion 857 -1170 857 -1170 0 cellNo=62
rlabel pdiffusion 864 -1170 864 -1170 0 feedthrough
rlabel pdiffusion 871 -1170 871 -1170 0 feedthrough
rlabel pdiffusion 878 -1170 878 -1170 0 feedthrough
rlabel pdiffusion 885 -1170 885 -1170 0 feedthrough
rlabel pdiffusion 892 -1170 892 -1170 0 feedthrough
rlabel pdiffusion 899 -1170 899 -1170 0 feedthrough
rlabel pdiffusion 906 -1170 906 -1170 0 feedthrough
rlabel pdiffusion 913 -1170 913 -1170 0 feedthrough
rlabel pdiffusion 920 -1170 920 -1170 0 feedthrough
rlabel pdiffusion 927 -1170 927 -1170 0 feedthrough
rlabel pdiffusion 934 -1170 934 -1170 0 feedthrough
rlabel pdiffusion 941 -1170 941 -1170 0 feedthrough
rlabel pdiffusion 948 -1170 948 -1170 0 feedthrough
rlabel pdiffusion 955 -1170 955 -1170 0 feedthrough
rlabel pdiffusion 962 -1170 962 -1170 0 feedthrough
rlabel pdiffusion 969 -1170 969 -1170 0 feedthrough
rlabel pdiffusion 976 -1170 976 -1170 0 feedthrough
rlabel pdiffusion 983 -1170 983 -1170 0 feedthrough
rlabel pdiffusion 990 -1170 990 -1170 0 feedthrough
rlabel pdiffusion 997 -1170 997 -1170 0 feedthrough
rlabel pdiffusion 1004 -1170 1004 -1170 0 feedthrough
rlabel pdiffusion 1011 -1170 1011 -1170 0 feedthrough
rlabel pdiffusion 1018 -1170 1018 -1170 0 feedthrough
rlabel pdiffusion 1025 -1170 1025 -1170 0 feedthrough
rlabel pdiffusion 1032 -1170 1032 -1170 0 feedthrough
rlabel pdiffusion 1039 -1170 1039 -1170 0 cellNo=291
rlabel pdiffusion 1046 -1170 1046 -1170 0 feedthrough
rlabel pdiffusion 1053 -1170 1053 -1170 0 feedthrough
rlabel pdiffusion 1060 -1170 1060 -1170 0 feedthrough
rlabel pdiffusion 1067 -1170 1067 -1170 0 feedthrough
rlabel pdiffusion 1074 -1170 1074 -1170 0 cellNo=825
rlabel pdiffusion 1123 -1170 1123 -1170 0 feedthrough
rlabel pdiffusion 1151 -1170 1151 -1170 0 feedthrough
rlabel pdiffusion 3 -1253 3 -1253 0 feedthrough
rlabel pdiffusion 10 -1253 10 -1253 0 feedthrough
rlabel pdiffusion 17 -1253 17 -1253 0 feedthrough
rlabel pdiffusion 24 -1253 24 -1253 0 cellNo=405
rlabel pdiffusion 31 -1253 31 -1253 0 feedthrough
rlabel pdiffusion 38 -1253 38 -1253 0 feedthrough
rlabel pdiffusion 45 -1253 45 -1253 0 cellNo=425
rlabel pdiffusion 52 -1253 52 -1253 0 feedthrough
rlabel pdiffusion 59 -1253 59 -1253 0 feedthrough
rlabel pdiffusion 66 -1253 66 -1253 0 feedthrough
rlabel pdiffusion 73 -1253 73 -1253 0 cellNo=46
rlabel pdiffusion 80 -1253 80 -1253 0 feedthrough
rlabel pdiffusion 87 -1253 87 -1253 0 feedthrough
rlabel pdiffusion 94 -1253 94 -1253 0 cellNo=301
rlabel pdiffusion 101 -1253 101 -1253 0 feedthrough
rlabel pdiffusion 108 -1253 108 -1253 0 feedthrough
rlabel pdiffusion 115 -1253 115 -1253 0 feedthrough
rlabel pdiffusion 122 -1253 122 -1253 0 feedthrough
rlabel pdiffusion 129 -1253 129 -1253 0 feedthrough
rlabel pdiffusion 136 -1253 136 -1253 0 feedthrough
rlabel pdiffusion 143 -1253 143 -1253 0 feedthrough
rlabel pdiffusion 150 -1253 150 -1253 0 feedthrough
rlabel pdiffusion 157 -1253 157 -1253 0 cellNo=241
rlabel pdiffusion 164 -1253 164 -1253 0 feedthrough
rlabel pdiffusion 171 -1253 171 -1253 0 feedthrough
rlabel pdiffusion 178 -1253 178 -1253 0 feedthrough
rlabel pdiffusion 185 -1253 185 -1253 0 cellNo=78
rlabel pdiffusion 192 -1253 192 -1253 0 cellNo=34
rlabel pdiffusion 199 -1253 199 -1253 0 cellNo=395
rlabel pdiffusion 206 -1253 206 -1253 0 feedthrough
rlabel pdiffusion 213 -1253 213 -1253 0 feedthrough
rlabel pdiffusion 220 -1253 220 -1253 0 feedthrough
rlabel pdiffusion 227 -1253 227 -1253 0 feedthrough
rlabel pdiffusion 234 -1253 234 -1253 0 feedthrough
rlabel pdiffusion 241 -1253 241 -1253 0 feedthrough
rlabel pdiffusion 248 -1253 248 -1253 0 feedthrough
rlabel pdiffusion 255 -1253 255 -1253 0 feedthrough
rlabel pdiffusion 262 -1253 262 -1253 0 feedthrough
rlabel pdiffusion 269 -1253 269 -1253 0 cellNo=499
rlabel pdiffusion 276 -1253 276 -1253 0 feedthrough
rlabel pdiffusion 283 -1253 283 -1253 0 feedthrough
rlabel pdiffusion 290 -1253 290 -1253 0 cellNo=446
rlabel pdiffusion 297 -1253 297 -1253 0 feedthrough
rlabel pdiffusion 304 -1253 304 -1253 0 cellNo=290
rlabel pdiffusion 311 -1253 311 -1253 0 feedthrough
rlabel pdiffusion 318 -1253 318 -1253 0 feedthrough
rlabel pdiffusion 325 -1253 325 -1253 0 feedthrough
rlabel pdiffusion 332 -1253 332 -1253 0 feedthrough
rlabel pdiffusion 339 -1253 339 -1253 0 feedthrough
rlabel pdiffusion 346 -1253 346 -1253 0 feedthrough
rlabel pdiffusion 353 -1253 353 -1253 0 feedthrough
rlabel pdiffusion 360 -1253 360 -1253 0 cellNo=108
rlabel pdiffusion 367 -1253 367 -1253 0 cellNo=79
rlabel pdiffusion 374 -1253 374 -1253 0 cellNo=964
rlabel pdiffusion 381 -1253 381 -1253 0 feedthrough
rlabel pdiffusion 388 -1253 388 -1253 0 feedthrough
rlabel pdiffusion 395 -1253 395 -1253 0 feedthrough
rlabel pdiffusion 402 -1253 402 -1253 0 feedthrough
rlabel pdiffusion 409 -1253 409 -1253 0 feedthrough
rlabel pdiffusion 416 -1253 416 -1253 0 feedthrough
rlabel pdiffusion 423 -1253 423 -1253 0 feedthrough
rlabel pdiffusion 430 -1253 430 -1253 0 feedthrough
rlabel pdiffusion 437 -1253 437 -1253 0 cellNo=200
rlabel pdiffusion 444 -1253 444 -1253 0 feedthrough
rlabel pdiffusion 451 -1253 451 -1253 0 feedthrough
rlabel pdiffusion 458 -1253 458 -1253 0 cellNo=584
rlabel pdiffusion 465 -1253 465 -1253 0 feedthrough
rlabel pdiffusion 472 -1253 472 -1253 0 feedthrough
rlabel pdiffusion 479 -1253 479 -1253 0 feedthrough
rlabel pdiffusion 486 -1253 486 -1253 0 feedthrough
rlabel pdiffusion 493 -1253 493 -1253 0 cellNo=615
rlabel pdiffusion 500 -1253 500 -1253 0 feedthrough
rlabel pdiffusion 507 -1253 507 -1253 0 cellNo=721
rlabel pdiffusion 514 -1253 514 -1253 0 feedthrough
rlabel pdiffusion 521 -1253 521 -1253 0 feedthrough
rlabel pdiffusion 528 -1253 528 -1253 0 feedthrough
rlabel pdiffusion 535 -1253 535 -1253 0 cellNo=654
rlabel pdiffusion 542 -1253 542 -1253 0 feedthrough
rlabel pdiffusion 549 -1253 549 -1253 0 feedthrough
rlabel pdiffusion 556 -1253 556 -1253 0 feedthrough
rlabel pdiffusion 563 -1253 563 -1253 0 feedthrough
rlabel pdiffusion 570 -1253 570 -1253 0 feedthrough
rlabel pdiffusion 577 -1253 577 -1253 0 feedthrough
rlabel pdiffusion 584 -1253 584 -1253 0 feedthrough
rlabel pdiffusion 591 -1253 591 -1253 0 feedthrough
rlabel pdiffusion 598 -1253 598 -1253 0 cellNo=966
rlabel pdiffusion 605 -1253 605 -1253 0 feedthrough
rlabel pdiffusion 612 -1253 612 -1253 0 feedthrough
rlabel pdiffusion 619 -1253 619 -1253 0 feedthrough
rlabel pdiffusion 626 -1253 626 -1253 0 feedthrough
rlabel pdiffusion 633 -1253 633 -1253 0 cellNo=387
rlabel pdiffusion 640 -1253 640 -1253 0 cellNo=501
rlabel pdiffusion 647 -1253 647 -1253 0 feedthrough
rlabel pdiffusion 654 -1253 654 -1253 0 cellNo=625
rlabel pdiffusion 661 -1253 661 -1253 0 feedthrough
rlabel pdiffusion 668 -1253 668 -1253 0 cellNo=640
rlabel pdiffusion 675 -1253 675 -1253 0 feedthrough
rlabel pdiffusion 682 -1253 682 -1253 0 cellNo=184
rlabel pdiffusion 689 -1253 689 -1253 0 feedthrough
rlabel pdiffusion 696 -1253 696 -1253 0 feedthrough
rlabel pdiffusion 703 -1253 703 -1253 0 cellNo=433
rlabel pdiffusion 710 -1253 710 -1253 0 feedthrough
rlabel pdiffusion 717 -1253 717 -1253 0 cellNo=995
rlabel pdiffusion 724 -1253 724 -1253 0 feedthrough
rlabel pdiffusion 731 -1253 731 -1253 0 feedthrough
rlabel pdiffusion 738 -1253 738 -1253 0 feedthrough
rlabel pdiffusion 745 -1253 745 -1253 0 feedthrough
rlabel pdiffusion 752 -1253 752 -1253 0 feedthrough
rlabel pdiffusion 759 -1253 759 -1253 0 feedthrough
rlabel pdiffusion 766 -1253 766 -1253 0 feedthrough
rlabel pdiffusion 773 -1253 773 -1253 0 feedthrough
rlabel pdiffusion 780 -1253 780 -1253 0 feedthrough
rlabel pdiffusion 787 -1253 787 -1253 0 cellNo=698
rlabel pdiffusion 794 -1253 794 -1253 0 feedthrough
rlabel pdiffusion 801 -1253 801 -1253 0 feedthrough
rlabel pdiffusion 808 -1253 808 -1253 0 feedthrough
rlabel pdiffusion 815 -1253 815 -1253 0 feedthrough
rlabel pdiffusion 822 -1253 822 -1253 0 feedthrough
rlabel pdiffusion 829 -1253 829 -1253 0 cellNo=5
rlabel pdiffusion 836 -1253 836 -1253 0 feedthrough
rlabel pdiffusion 843 -1253 843 -1253 0 feedthrough
rlabel pdiffusion 850 -1253 850 -1253 0 feedthrough
rlabel pdiffusion 857 -1253 857 -1253 0 feedthrough
rlabel pdiffusion 864 -1253 864 -1253 0 feedthrough
rlabel pdiffusion 871 -1253 871 -1253 0 feedthrough
rlabel pdiffusion 878 -1253 878 -1253 0 feedthrough
rlabel pdiffusion 885 -1253 885 -1253 0 feedthrough
rlabel pdiffusion 892 -1253 892 -1253 0 feedthrough
rlabel pdiffusion 899 -1253 899 -1253 0 feedthrough
rlabel pdiffusion 906 -1253 906 -1253 0 feedthrough
rlabel pdiffusion 913 -1253 913 -1253 0 feedthrough
rlabel pdiffusion 920 -1253 920 -1253 0 feedthrough
rlabel pdiffusion 927 -1253 927 -1253 0 feedthrough
rlabel pdiffusion 934 -1253 934 -1253 0 feedthrough
rlabel pdiffusion 941 -1253 941 -1253 0 feedthrough
rlabel pdiffusion 948 -1253 948 -1253 0 feedthrough
rlabel pdiffusion 955 -1253 955 -1253 0 feedthrough
rlabel pdiffusion 962 -1253 962 -1253 0 feedthrough
rlabel pdiffusion 969 -1253 969 -1253 0 cellNo=492
rlabel pdiffusion 976 -1253 976 -1253 0 feedthrough
rlabel pdiffusion 983 -1253 983 -1253 0 feedthrough
rlabel pdiffusion 990 -1253 990 -1253 0 feedthrough
rlabel pdiffusion 997 -1253 997 -1253 0 feedthrough
rlabel pdiffusion 1004 -1253 1004 -1253 0 feedthrough
rlabel pdiffusion 1011 -1253 1011 -1253 0 feedthrough
rlabel pdiffusion 1018 -1253 1018 -1253 0 feedthrough
rlabel pdiffusion 1025 -1253 1025 -1253 0 feedthrough
rlabel pdiffusion 1032 -1253 1032 -1253 0 feedthrough
rlabel pdiffusion 1039 -1253 1039 -1253 0 feedthrough
rlabel pdiffusion 1046 -1253 1046 -1253 0 feedthrough
rlabel pdiffusion 1053 -1253 1053 -1253 0 feedthrough
rlabel pdiffusion 1060 -1253 1060 -1253 0 feedthrough
rlabel pdiffusion 1067 -1253 1067 -1253 0 feedthrough
rlabel pdiffusion 1074 -1253 1074 -1253 0 feedthrough
rlabel pdiffusion 1081 -1253 1081 -1253 0 feedthrough
rlabel pdiffusion 1088 -1253 1088 -1253 0 feedthrough
rlabel pdiffusion 1095 -1253 1095 -1253 0 feedthrough
rlabel pdiffusion 1102 -1253 1102 -1253 0 feedthrough
rlabel pdiffusion 1109 -1253 1109 -1253 0 feedthrough
rlabel pdiffusion 1116 -1253 1116 -1253 0 cellNo=227
rlabel pdiffusion 1123 -1253 1123 -1253 0 feedthrough
rlabel pdiffusion 1130 -1253 1130 -1253 0 cellNo=622
rlabel pdiffusion 1137 -1253 1137 -1253 0 feedthrough
rlabel pdiffusion 1144 -1253 1144 -1253 0 feedthrough
rlabel pdiffusion 1151 -1253 1151 -1253 0 feedthrough
rlabel pdiffusion 1158 -1253 1158 -1253 0 feedthrough
rlabel pdiffusion 1165 -1253 1165 -1253 0 feedthrough
rlabel pdiffusion 3 -1346 3 -1346 0 feedthrough
rlabel pdiffusion 10 -1346 10 -1346 0 feedthrough
rlabel pdiffusion 17 -1346 17 -1346 0 feedthrough
rlabel pdiffusion 24 -1346 24 -1346 0 cellNo=743
rlabel pdiffusion 31 -1346 31 -1346 0 cellNo=552
rlabel pdiffusion 38 -1346 38 -1346 0 feedthrough
rlabel pdiffusion 45 -1346 45 -1346 0 feedthrough
rlabel pdiffusion 52 -1346 52 -1346 0 feedthrough
rlabel pdiffusion 59 -1346 59 -1346 0 feedthrough
rlabel pdiffusion 66 -1346 66 -1346 0 cellNo=444
rlabel pdiffusion 73 -1346 73 -1346 0 feedthrough
rlabel pdiffusion 80 -1346 80 -1346 0 feedthrough
rlabel pdiffusion 87 -1346 87 -1346 0 feedthrough
rlabel pdiffusion 94 -1346 94 -1346 0 cellNo=655
rlabel pdiffusion 101 -1346 101 -1346 0 cellNo=873
rlabel pdiffusion 108 -1346 108 -1346 0 feedthrough
rlabel pdiffusion 115 -1346 115 -1346 0 feedthrough
rlabel pdiffusion 122 -1346 122 -1346 0 feedthrough
rlabel pdiffusion 129 -1346 129 -1346 0 feedthrough
rlabel pdiffusion 136 -1346 136 -1346 0 feedthrough
rlabel pdiffusion 143 -1346 143 -1346 0 feedthrough
rlabel pdiffusion 150 -1346 150 -1346 0 feedthrough
rlabel pdiffusion 157 -1346 157 -1346 0 feedthrough
rlabel pdiffusion 164 -1346 164 -1346 0 cellNo=582
rlabel pdiffusion 171 -1346 171 -1346 0 feedthrough
rlabel pdiffusion 178 -1346 178 -1346 0 cellNo=89
rlabel pdiffusion 185 -1346 185 -1346 0 feedthrough
rlabel pdiffusion 192 -1346 192 -1346 0 feedthrough
rlabel pdiffusion 199 -1346 199 -1346 0 feedthrough
rlabel pdiffusion 206 -1346 206 -1346 0 feedthrough
rlabel pdiffusion 213 -1346 213 -1346 0 cellNo=183
rlabel pdiffusion 220 -1346 220 -1346 0 feedthrough
rlabel pdiffusion 227 -1346 227 -1346 0 feedthrough
rlabel pdiffusion 234 -1346 234 -1346 0 feedthrough
rlabel pdiffusion 241 -1346 241 -1346 0 feedthrough
rlabel pdiffusion 248 -1346 248 -1346 0 feedthrough
rlabel pdiffusion 255 -1346 255 -1346 0 feedthrough
rlabel pdiffusion 262 -1346 262 -1346 0 feedthrough
rlabel pdiffusion 269 -1346 269 -1346 0 feedthrough
rlabel pdiffusion 276 -1346 276 -1346 0 feedthrough
rlabel pdiffusion 283 -1346 283 -1346 0 feedthrough
rlabel pdiffusion 290 -1346 290 -1346 0 cellNo=165
rlabel pdiffusion 297 -1346 297 -1346 0 feedthrough
rlabel pdiffusion 304 -1346 304 -1346 0 feedthrough
rlabel pdiffusion 311 -1346 311 -1346 0 feedthrough
rlabel pdiffusion 318 -1346 318 -1346 0 feedthrough
rlabel pdiffusion 325 -1346 325 -1346 0 feedthrough
rlabel pdiffusion 332 -1346 332 -1346 0 feedthrough
rlabel pdiffusion 339 -1346 339 -1346 0 feedthrough
rlabel pdiffusion 346 -1346 346 -1346 0 cellNo=18
rlabel pdiffusion 353 -1346 353 -1346 0 feedthrough
rlabel pdiffusion 360 -1346 360 -1346 0 feedthrough
rlabel pdiffusion 367 -1346 367 -1346 0 feedthrough
rlabel pdiffusion 374 -1346 374 -1346 0 feedthrough
rlabel pdiffusion 381 -1346 381 -1346 0 feedthrough
rlabel pdiffusion 388 -1346 388 -1346 0 feedthrough
rlabel pdiffusion 395 -1346 395 -1346 0 feedthrough
rlabel pdiffusion 402 -1346 402 -1346 0 cellNo=71
rlabel pdiffusion 409 -1346 409 -1346 0 cellNo=306
rlabel pdiffusion 416 -1346 416 -1346 0 feedthrough
rlabel pdiffusion 423 -1346 423 -1346 0 feedthrough
rlabel pdiffusion 430 -1346 430 -1346 0 feedthrough
rlabel pdiffusion 437 -1346 437 -1346 0 cellNo=14
rlabel pdiffusion 444 -1346 444 -1346 0 feedthrough
rlabel pdiffusion 451 -1346 451 -1346 0 feedthrough
rlabel pdiffusion 458 -1346 458 -1346 0 cellNo=187
rlabel pdiffusion 465 -1346 465 -1346 0 feedthrough
rlabel pdiffusion 472 -1346 472 -1346 0 feedthrough
rlabel pdiffusion 479 -1346 479 -1346 0 feedthrough
rlabel pdiffusion 486 -1346 486 -1346 0 feedthrough
rlabel pdiffusion 493 -1346 493 -1346 0 cellNo=560
rlabel pdiffusion 500 -1346 500 -1346 0 feedthrough
rlabel pdiffusion 507 -1346 507 -1346 0 feedthrough
rlabel pdiffusion 514 -1346 514 -1346 0 feedthrough
rlabel pdiffusion 521 -1346 521 -1346 0 cellNo=417
rlabel pdiffusion 528 -1346 528 -1346 0 feedthrough
rlabel pdiffusion 535 -1346 535 -1346 0 cellNo=132
rlabel pdiffusion 542 -1346 542 -1346 0 cellNo=439
rlabel pdiffusion 549 -1346 549 -1346 0 feedthrough
rlabel pdiffusion 556 -1346 556 -1346 0 feedthrough
rlabel pdiffusion 563 -1346 563 -1346 0 feedthrough
rlabel pdiffusion 570 -1346 570 -1346 0 cellNo=127
rlabel pdiffusion 577 -1346 577 -1346 0 feedthrough
rlabel pdiffusion 584 -1346 584 -1346 0 feedthrough
rlabel pdiffusion 591 -1346 591 -1346 0 feedthrough
rlabel pdiffusion 598 -1346 598 -1346 0 feedthrough
rlabel pdiffusion 605 -1346 605 -1346 0 cellNo=864
rlabel pdiffusion 612 -1346 612 -1346 0 cellNo=859
rlabel pdiffusion 619 -1346 619 -1346 0 cellNo=113
rlabel pdiffusion 626 -1346 626 -1346 0 cellNo=924
rlabel pdiffusion 633 -1346 633 -1346 0 feedthrough
rlabel pdiffusion 640 -1346 640 -1346 0 feedthrough
rlabel pdiffusion 647 -1346 647 -1346 0 feedthrough
rlabel pdiffusion 654 -1346 654 -1346 0 feedthrough
rlabel pdiffusion 661 -1346 661 -1346 0 feedthrough
rlabel pdiffusion 668 -1346 668 -1346 0 feedthrough
rlabel pdiffusion 675 -1346 675 -1346 0 feedthrough
rlabel pdiffusion 682 -1346 682 -1346 0 cellNo=460
rlabel pdiffusion 689 -1346 689 -1346 0 feedthrough
rlabel pdiffusion 696 -1346 696 -1346 0 feedthrough
rlabel pdiffusion 703 -1346 703 -1346 0 feedthrough
rlabel pdiffusion 710 -1346 710 -1346 0 feedthrough
rlabel pdiffusion 717 -1346 717 -1346 0 feedthrough
rlabel pdiffusion 724 -1346 724 -1346 0 feedthrough
rlabel pdiffusion 731 -1346 731 -1346 0 cellNo=795
rlabel pdiffusion 738 -1346 738 -1346 0 feedthrough
rlabel pdiffusion 745 -1346 745 -1346 0 feedthrough
rlabel pdiffusion 752 -1346 752 -1346 0 feedthrough
rlabel pdiffusion 759 -1346 759 -1346 0 feedthrough
rlabel pdiffusion 766 -1346 766 -1346 0 feedthrough
rlabel pdiffusion 773 -1346 773 -1346 0 cellNo=860
rlabel pdiffusion 780 -1346 780 -1346 0 feedthrough
rlabel pdiffusion 787 -1346 787 -1346 0 feedthrough
rlabel pdiffusion 794 -1346 794 -1346 0 cellNo=841
rlabel pdiffusion 801 -1346 801 -1346 0 feedthrough
rlabel pdiffusion 808 -1346 808 -1346 0 feedthrough
rlabel pdiffusion 815 -1346 815 -1346 0 feedthrough
rlabel pdiffusion 822 -1346 822 -1346 0 feedthrough
rlabel pdiffusion 829 -1346 829 -1346 0 cellNo=43
rlabel pdiffusion 836 -1346 836 -1346 0 feedthrough
rlabel pdiffusion 843 -1346 843 -1346 0 feedthrough
rlabel pdiffusion 850 -1346 850 -1346 0 feedthrough
rlabel pdiffusion 857 -1346 857 -1346 0 feedthrough
rlabel pdiffusion 864 -1346 864 -1346 0 feedthrough
rlabel pdiffusion 871 -1346 871 -1346 0 feedthrough
rlabel pdiffusion 878 -1346 878 -1346 0 feedthrough
rlabel pdiffusion 885 -1346 885 -1346 0 feedthrough
rlabel pdiffusion 892 -1346 892 -1346 0 feedthrough
rlabel pdiffusion 899 -1346 899 -1346 0 feedthrough
rlabel pdiffusion 906 -1346 906 -1346 0 feedthrough
rlabel pdiffusion 913 -1346 913 -1346 0 feedthrough
rlabel pdiffusion 920 -1346 920 -1346 0 feedthrough
rlabel pdiffusion 927 -1346 927 -1346 0 feedthrough
rlabel pdiffusion 934 -1346 934 -1346 0 feedthrough
rlabel pdiffusion 941 -1346 941 -1346 0 feedthrough
rlabel pdiffusion 948 -1346 948 -1346 0 cellNo=104
rlabel pdiffusion 955 -1346 955 -1346 0 feedthrough
rlabel pdiffusion 962 -1346 962 -1346 0 feedthrough
rlabel pdiffusion 969 -1346 969 -1346 0 feedthrough
rlabel pdiffusion 976 -1346 976 -1346 0 feedthrough
rlabel pdiffusion 983 -1346 983 -1346 0 feedthrough
rlabel pdiffusion 990 -1346 990 -1346 0 feedthrough
rlabel pdiffusion 997 -1346 997 -1346 0 cellNo=354
rlabel pdiffusion 1004 -1346 1004 -1346 0 feedthrough
rlabel pdiffusion 1011 -1346 1011 -1346 0 feedthrough
rlabel pdiffusion 1018 -1346 1018 -1346 0 feedthrough
rlabel pdiffusion 1025 -1346 1025 -1346 0 feedthrough
rlabel pdiffusion 1032 -1346 1032 -1346 0 feedthrough
rlabel pdiffusion 1039 -1346 1039 -1346 0 feedthrough
rlabel pdiffusion 1046 -1346 1046 -1346 0 feedthrough
rlabel pdiffusion 1053 -1346 1053 -1346 0 feedthrough
rlabel pdiffusion 1060 -1346 1060 -1346 0 feedthrough
rlabel pdiffusion 1067 -1346 1067 -1346 0 feedthrough
rlabel pdiffusion 1074 -1346 1074 -1346 0 feedthrough
rlabel pdiffusion 1081 -1346 1081 -1346 0 feedthrough
rlabel pdiffusion 1088 -1346 1088 -1346 0 feedthrough
rlabel pdiffusion 1095 -1346 1095 -1346 0 feedthrough
rlabel pdiffusion 1102 -1346 1102 -1346 0 feedthrough
rlabel pdiffusion 1109 -1346 1109 -1346 0 feedthrough
rlabel pdiffusion 1116 -1346 1116 -1346 0 feedthrough
rlabel pdiffusion 1123 -1346 1123 -1346 0 feedthrough
rlabel pdiffusion 1130 -1346 1130 -1346 0 feedthrough
rlabel pdiffusion 1137 -1346 1137 -1346 0 cellNo=365
rlabel pdiffusion 1144 -1346 1144 -1346 0 feedthrough
rlabel pdiffusion 1151 -1346 1151 -1346 0 cellNo=852
rlabel pdiffusion 1158 -1346 1158 -1346 0 feedthrough
rlabel pdiffusion 1165 -1346 1165 -1346 0 feedthrough
rlabel pdiffusion 1172 -1346 1172 -1346 0 feedthrough
rlabel pdiffusion 3 -1453 3 -1453 0 feedthrough
rlabel pdiffusion 10 -1453 10 -1453 0 cellNo=198
rlabel pdiffusion 17 -1453 17 -1453 0 feedthrough
rlabel pdiffusion 24 -1453 24 -1453 0 feedthrough
rlabel pdiffusion 31 -1453 31 -1453 0 feedthrough
rlabel pdiffusion 38 -1453 38 -1453 0 feedthrough
rlabel pdiffusion 45 -1453 45 -1453 0 feedthrough
rlabel pdiffusion 52 -1453 52 -1453 0 feedthrough
rlabel pdiffusion 59 -1453 59 -1453 0 feedthrough
rlabel pdiffusion 66 -1453 66 -1453 0 feedthrough
rlabel pdiffusion 73 -1453 73 -1453 0 feedthrough
rlabel pdiffusion 80 -1453 80 -1453 0 feedthrough
rlabel pdiffusion 87 -1453 87 -1453 0 feedthrough
rlabel pdiffusion 94 -1453 94 -1453 0 feedthrough
rlabel pdiffusion 101 -1453 101 -1453 0 cellNo=527
rlabel pdiffusion 108 -1453 108 -1453 0 cellNo=243
rlabel pdiffusion 115 -1453 115 -1453 0 cellNo=287
rlabel pdiffusion 122 -1453 122 -1453 0 cellNo=77
rlabel pdiffusion 129 -1453 129 -1453 0 feedthrough
rlabel pdiffusion 136 -1453 136 -1453 0 feedthrough
rlabel pdiffusion 143 -1453 143 -1453 0 feedthrough
rlabel pdiffusion 150 -1453 150 -1453 0 feedthrough
rlabel pdiffusion 157 -1453 157 -1453 0 feedthrough
rlabel pdiffusion 164 -1453 164 -1453 0 feedthrough
rlabel pdiffusion 171 -1453 171 -1453 0 feedthrough
rlabel pdiffusion 178 -1453 178 -1453 0 cellNo=954
rlabel pdiffusion 185 -1453 185 -1453 0 cellNo=469
rlabel pdiffusion 192 -1453 192 -1453 0 cellNo=579
rlabel pdiffusion 199 -1453 199 -1453 0 feedthrough
rlabel pdiffusion 206 -1453 206 -1453 0 feedthrough
rlabel pdiffusion 213 -1453 213 -1453 0 cellNo=563
rlabel pdiffusion 220 -1453 220 -1453 0 feedthrough
rlabel pdiffusion 227 -1453 227 -1453 0 feedthrough
rlabel pdiffusion 234 -1453 234 -1453 0 feedthrough
rlabel pdiffusion 241 -1453 241 -1453 0 feedthrough
rlabel pdiffusion 248 -1453 248 -1453 0 feedthrough
rlabel pdiffusion 255 -1453 255 -1453 0 cellNo=150
rlabel pdiffusion 262 -1453 262 -1453 0 feedthrough
rlabel pdiffusion 269 -1453 269 -1453 0 feedthrough
rlabel pdiffusion 276 -1453 276 -1453 0 feedthrough
rlabel pdiffusion 283 -1453 283 -1453 0 feedthrough
rlabel pdiffusion 290 -1453 290 -1453 0 feedthrough
rlabel pdiffusion 297 -1453 297 -1453 0 feedthrough
rlabel pdiffusion 304 -1453 304 -1453 0 feedthrough
rlabel pdiffusion 311 -1453 311 -1453 0 feedthrough
rlabel pdiffusion 318 -1453 318 -1453 0 feedthrough
rlabel pdiffusion 325 -1453 325 -1453 0 feedthrough
rlabel pdiffusion 332 -1453 332 -1453 0 cellNo=883
rlabel pdiffusion 339 -1453 339 -1453 0 feedthrough
rlabel pdiffusion 346 -1453 346 -1453 0 feedthrough
rlabel pdiffusion 353 -1453 353 -1453 0 feedthrough
rlabel pdiffusion 360 -1453 360 -1453 0 feedthrough
rlabel pdiffusion 367 -1453 367 -1453 0 feedthrough
rlabel pdiffusion 374 -1453 374 -1453 0 feedthrough
rlabel pdiffusion 381 -1453 381 -1453 0 feedthrough
rlabel pdiffusion 388 -1453 388 -1453 0 feedthrough
rlabel pdiffusion 395 -1453 395 -1453 0 feedthrough
rlabel pdiffusion 402 -1453 402 -1453 0 cellNo=345
rlabel pdiffusion 409 -1453 409 -1453 0 cellNo=569
rlabel pdiffusion 416 -1453 416 -1453 0 feedthrough
rlabel pdiffusion 423 -1453 423 -1453 0 feedthrough
rlabel pdiffusion 430 -1453 430 -1453 0 cellNo=166
rlabel pdiffusion 437 -1453 437 -1453 0 cellNo=833
rlabel pdiffusion 444 -1453 444 -1453 0 cellNo=82
rlabel pdiffusion 451 -1453 451 -1453 0 feedthrough
rlabel pdiffusion 458 -1453 458 -1453 0 feedthrough
rlabel pdiffusion 465 -1453 465 -1453 0 feedthrough
rlabel pdiffusion 472 -1453 472 -1453 0 feedthrough
rlabel pdiffusion 479 -1453 479 -1453 0 cellNo=119
rlabel pdiffusion 486 -1453 486 -1453 0 cellNo=627
rlabel pdiffusion 493 -1453 493 -1453 0 cellNo=474
rlabel pdiffusion 500 -1453 500 -1453 0 cellNo=555
rlabel pdiffusion 507 -1453 507 -1453 0 cellNo=401
rlabel pdiffusion 514 -1453 514 -1453 0 feedthrough
rlabel pdiffusion 521 -1453 521 -1453 0 feedthrough
rlabel pdiffusion 528 -1453 528 -1453 0 feedthrough
rlabel pdiffusion 535 -1453 535 -1453 0 feedthrough
rlabel pdiffusion 542 -1453 542 -1453 0 feedthrough
rlabel pdiffusion 549 -1453 549 -1453 0 cellNo=636
rlabel pdiffusion 556 -1453 556 -1453 0 feedthrough
rlabel pdiffusion 563 -1453 563 -1453 0 feedthrough
rlabel pdiffusion 570 -1453 570 -1453 0 cellNo=744
rlabel pdiffusion 577 -1453 577 -1453 0 cellNo=661
rlabel pdiffusion 584 -1453 584 -1453 0 feedthrough
rlabel pdiffusion 591 -1453 591 -1453 0 feedthrough
rlabel pdiffusion 598 -1453 598 -1453 0 cellNo=726
rlabel pdiffusion 605 -1453 605 -1453 0 feedthrough
rlabel pdiffusion 612 -1453 612 -1453 0 cellNo=851
rlabel pdiffusion 619 -1453 619 -1453 0 feedthrough
rlabel pdiffusion 626 -1453 626 -1453 0 feedthrough
rlabel pdiffusion 633 -1453 633 -1453 0 feedthrough
rlabel pdiffusion 640 -1453 640 -1453 0 feedthrough
rlabel pdiffusion 647 -1453 647 -1453 0 feedthrough
rlabel pdiffusion 654 -1453 654 -1453 0 feedthrough
rlabel pdiffusion 661 -1453 661 -1453 0 feedthrough
rlabel pdiffusion 668 -1453 668 -1453 0 feedthrough
rlabel pdiffusion 675 -1453 675 -1453 0 feedthrough
rlabel pdiffusion 682 -1453 682 -1453 0 feedthrough
rlabel pdiffusion 689 -1453 689 -1453 0 cellNo=665
rlabel pdiffusion 696 -1453 696 -1453 0 feedthrough
rlabel pdiffusion 703 -1453 703 -1453 0 cellNo=475
rlabel pdiffusion 710 -1453 710 -1453 0 feedthrough
rlabel pdiffusion 717 -1453 717 -1453 0 feedthrough
rlabel pdiffusion 724 -1453 724 -1453 0 feedthrough
rlabel pdiffusion 731 -1453 731 -1453 0 feedthrough
rlabel pdiffusion 738 -1453 738 -1453 0 feedthrough
rlabel pdiffusion 745 -1453 745 -1453 0 cellNo=305
rlabel pdiffusion 752 -1453 752 -1453 0 feedthrough
rlabel pdiffusion 759 -1453 759 -1453 0 feedthrough
rlabel pdiffusion 766 -1453 766 -1453 0 feedthrough
rlabel pdiffusion 773 -1453 773 -1453 0 feedthrough
rlabel pdiffusion 780 -1453 780 -1453 0 feedthrough
rlabel pdiffusion 787 -1453 787 -1453 0 feedthrough
rlabel pdiffusion 794 -1453 794 -1453 0 feedthrough
rlabel pdiffusion 801 -1453 801 -1453 0 feedthrough
rlabel pdiffusion 808 -1453 808 -1453 0 feedthrough
rlabel pdiffusion 815 -1453 815 -1453 0 feedthrough
rlabel pdiffusion 822 -1453 822 -1453 0 feedthrough
rlabel pdiffusion 829 -1453 829 -1453 0 feedthrough
rlabel pdiffusion 836 -1453 836 -1453 0 feedthrough
rlabel pdiffusion 843 -1453 843 -1453 0 feedthrough
rlabel pdiffusion 850 -1453 850 -1453 0 feedthrough
rlabel pdiffusion 857 -1453 857 -1453 0 cellNo=962
rlabel pdiffusion 864 -1453 864 -1453 0 feedthrough
rlabel pdiffusion 871 -1453 871 -1453 0 feedthrough
rlabel pdiffusion 878 -1453 878 -1453 0 feedthrough
rlabel pdiffusion 885 -1453 885 -1453 0 feedthrough
rlabel pdiffusion 892 -1453 892 -1453 0 feedthrough
rlabel pdiffusion 899 -1453 899 -1453 0 feedthrough
rlabel pdiffusion 906 -1453 906 -1453 0 feedthrough
rlabel pdiffusion 913 -1453 913 -1453 0 feedthrough
rlabel pdiffusion 920 -1453 920 -1453 0 feedthrough
rlabel pdiffusion 927 -1453 927 -1453 0 feedthrough
rlabel pdiffusion 934 -1453 934 -1453 0 feedthrough
rlabel pdiffusion 941 -1453 941 -1453 0 feedthrough
rlabel pdiffusion 948 -1453 948 -1453 0 feedthrough
rlabel pdiffusion 955 -1453 955 -1453 0 feedthrough
rlabel pdiffusion 962 -1453 962 -1453 0 feedthrough
rlabel pdiffusion 969 -1453 969 -1453 0 feedthrough
rlabel pdiffusion 976 -1453 976 -1453 0 feedthrough
rlabel pdiffusion 983 -1453 983 -1453 0 feedthrough
rlabel pdiffusion 990 -1453 990 -1453 0 feedthrough
rlabel pdiffusion 997 -1453 997 -1453 0 feedthrough
rlabel pdiffusion 1004 -1453 1004 -1453 0 feedthrough
rlabel pdiffusion 1011 -1453 1011 -1453 0 feedthrough
rlabel pdiffusion 1018 -1453 1018 -1453 0 feedthrough
rlabel pdiffusion 1025 -1453 1025 -1453 0 feedthrough
rlabel pdiffusion 1032 -1453 1032 -1453 0 feedthrough
rlabel pdiffusion 1039 -1453 1039 -1453 0 feedthrough
rlabel pdiffusion 1046 -1453 1046 -1453 0 feedthrough
rlabel pdiffusion 1053 -1453 1053 -1453 0 feedthrough
rlabel pdiffusion 1060 -1453 1060 -1453 0 cellNo=98
rlabel pdiffusion 1067 -1453 1067 -1453 0 feedthrough
rlabel pdiffusion 1074 -1453 1074 -1453 0 feedthrough
rlabel pdiffusion 1081 -1453 1081 -1453 0 feedthrough
rlabel pdiffusion 1088 -1453 1088 -1453 0 cellNo=968
rlabel pdiffusion 1095 -1453 1095 -1453 0 feedthrough
rlabel pdiffusion 1109 -1453 1109 -1453 0 feedthrough
rlabel pdiffusion 3 -1544 3 -1544 0 feedthrough
rlabel pdiffusion 10 -1544 10 -1544 0 feedthrough
rlabel pdiffusion 17 -1544 17 -1544 0 feedthrough
rlabel pdiffusion 24 -1544 24 -1544 0 feedthrough
rlabel pdiffusion 31 -1544 31 -1544 0 cellNo=854
rlabel pdiffusion 38 -1544 38 -1544 0 cellNo=650
rlabel pdiffusion 45 -1544 45 -1544 0 feedthrough
rlabel pdiffusion 52 -1544 52 -1544 0 feedthrough
rlabel pdiffusion 59 -1544 59 -1544 0 feedthrough
rlabel pdiffusion 66 -1544 66 -1544 0 feedthrough
rlabel pdiffusion 73 -1544 73 -1544 0 feedthrough
rlabel pdiffusion 80 -1544 80 -1544 0 feedthrough
rlabel pdiffusion 87 -1544 87 -1544 0 feedthrough
rlabel pdiffusion 94 -1544 94 -1544 0 cellNo=420
rlabel pdiffusion 101 -1544 101 -1544 0 feedthrough
rlabel pdiffusion 108 -1544 108 -1544 0 feedthrough
rlabel pdiffusion 115 -1544 115 -1544 0 feedthrough
rlabel pdiffusion 122 -1544 122 -1544 0 feedthrough
rlabel pdiffusion 129 -1544 129 -1544 0 feedthrough
rlabel pdiffusion 136 -1544 136 -1544 0 feedthrough
rlabel pdiffusion 143 -1544 143 -1544 0 cellNo=105
rlabel pdiffusion 150 -1544 150 -1544 0 feedthrough
rlabel pdiffusion 157 -1544 157 -1544 0 cellNo=120
rlabel pdiffusion 164 -1544 164 -1544 0 cellNo=641
rlabel pdiffusion 171 -1544 171 -1544 0 feedthrough
rlabel pdiffusion 178 -1544 178 -1544 0 cellNo=154
rlabel pdiffusion 185 -1544 185 -1544 0 feedthrough
rlabel pdiffusion 192 -1544 192 -1544 0 feedthrough
rlabel pdiffusion 199 -1544 199 -1544 0 feedthrough
rlabel pdiffusion 206 -1544 206 -1544 0 cellNo=167
rlabel pdiffusion 213 -1544 213 -1544 0 cellNo=722
rlabel pdiffusion 220 -1544 220 -1544 0 cellNo=905
rlabel pdiffusion 227 -1544 227 -1544 0 feedthrough
rlabel pdiffusion 234 -1544 234 -1544 0 feedthrough
rlabel pdiffusion 241 -1544 241 -1544 0 feedthrough
rlabel pdiffusion 248 -1544 248 -1544 0 cellNo=382
rlabel pdiffusion 255 -1544 255 -1544 0 feedthrough
rlabel pdiffusion 262 -1544 262 -1544 0 feedthrough
rlabel pdiffusion 269 -1544 269 -1544 0 feedthrough
rlabel pdiffusion 276 -1544 276 -1544 0 cellNo=946
rlabel pdiffusion 283 -1544 283 -1544 0 feedthrough
rlabel pdiffusion 290 -1544 290 -1544 0 cellNo=239
rlabel pdiffusion 297 -1544 297 -1544 0 feedthrough
rlabel pdiffusion 304 -1544 304 -1544 0 feedthrough
rlabel pdiffusion 311 -1544 311 -1544 0 feedthrough
rlabel pdiffusion 318 -1544 318 -1544 0 feedthrough
rlabel pdiffusion 325 -1544 325 -1544 0 cellNo=904
rlabel pdiffusion 332 -1544 332 -1544 0 feedthrough
rlabel pdiffusion 339 -1544 339 -1544 0 feedthrough
rlabel pdiffusion 346 -1544 346 -1544 0 feedthrough
rlabel pdiffusion 353 -1544 353 -1544 0 feedthrough
rlabel pdiffusion 360 -1544 360 -1544 0 cellNo=372
rlabel pdiffusion 367 -1544 367 -1544 0 feedthrough
rlabel pdiffusion 374 -1544 374 -1544 0 feedthrough
rlabel pdiffusion 381 -1544 381 -1544 0 feedthrough
rlabel pdiffusion 388 -1544 388 -1544 0 feedthrough
rlabel pdiffusion 395 -1544 395 -1544 0 feedthrough
rlabel pdiffusion 402 -1544 402 -1544 0 feedthrough
rlabel pdiffusion 409 -1544 409 -1544 0 feedthrough
rlabel pdiffusion 416 -1544 416 -1544 0 feedthrough
rlabel pdiffusion 423 -1544 423 -1544 0 feedthrough
rlabel pdiffusion 430 -1544 430 -1544 0 feedthrough
rlabel pdiffusion 437 -1544 437 -1544 0 feedthrough
rlabel pdiffusion 444 -1544 444 -1544 0 feedthrough
rlabel pdiffusion 451 -1544 451 -1544 0 feedthrough
rlabel pdiffusion 458 -1544 458 -1544 0 cellNo=947
rlabel pdiffusion 465 -1544 465 -1544 0 cellNo=561
rlabel pdiffusion 472 -1544 472 -1544 0 cellNo=351
rlabel pdiffusion 479 -1544 479 -1544 0 cellNo=188
rlabel pdiffusion 486 -1544 486 -1544 0 cellNo=479
rlabel pdiffusion 493 -1544 493 -1544 0 feedthrough
rlabel pdiffusion 500 -1544 500 -1544 0 feedthrough
rlabel pdiffusion 507 -1544 507 -1544 0 feedthrough
rlabel pdiffusion 514 -1544 514 -1544 0 cellNo=998
rlabel pdiffusion 521 -1544 521 -1544 0 cellNo=204
rlabel pdiffusion 528 -1544 528 -1544 0 feedthrough
rlabel pdiffusion 535 -1544 535 -1544 0 cellNo=30
rlabel pdiffusion 542 -1544 542 -1544 0 feedthrough
rlabel pdiffusion 549 -1544 549 -1544 0 feedthrough
rlabel pdiffusion 556 -1544 556 -1544 0 feedthrough
rlabel pdiffusion 563 -1544 563 -1544 0 cellNo=544
rlabel pdiffusion 570 -1544 570 -1544 0 feedthrough
rlabel pdiffusion 577 -1544 577 -1544 0 feedthrough
rlabel pdiffusion 584 -1544 584 -1544 0 feedthrough
rlabel pdiffusion 591 -1544 591 -1544 0 cellNo=275
rlabel pdiffusion 598 -1544 598 -1544 0 feedthrough
rlabel pdiffusion 605 -1544 605 -1544 0 feedthrough
rlabel pdiffusion 612 -1544 612 -1544 0 feedthrough
rlabel pdiffusion 619 -1544 619 -1544 0 feedthrough
rlabel pdiffusion 626 -1544 626 -1544 0 feedthrough
rlabel pdiffusion 633 -1544 633 -1544 0 feedthrough
rlabel pdiffusion 640 -1544 640 -1544 0 feedthrough
rlabel pdiffusion 647 -1544 647 -1544 0 feedthrough
rlabel pdiffusion 654 -1544 654 -1544 0 feedthrough
rlabel pdiffusion 661 -1544 661 -1544 0 cellNo=785
rlabel pdiffusion 668 -1544 668 -1544 0 cellNo=265
rlabel pdiffusion 675 -1544 675 -1544 0 cellNo=69
rlabel pdiffusion 682 -1544 682 -1544 0 feedthrough
rlabel pdiffusion 689 -1544 689 -1544 0 cellNo=517
rlabel pdiffusion 696 -1544 696 -1544 0 feedthrough
rlabel pdiffusion 703 -1544 703 -1544 0 feedthrough
rlabel pdiffusion 710 -1544 710 -1544 0 feedthrough
rlabel pdiffusion 717 -1544 717 -1544 0 feedthrough
rlabel pdiffusion 724 -1544 724 -1544 0 feedthrough
rlabel pdiffusion 731 -1544 731 -1544 0 feedthrough
rlabel pdiffusion 738 -1544 738 -1544 0 feedthrough
rlabel pdiffusion 745 -1544 745 -1544 0 feedthrough
rlabel pdiffusion 752 -1544 752 -1544 0 feedthrough
rlabel pdiffusion 759 -1544 759 -1544 0 feedthrough
rlabel pdiffusion 766 -1544 766 -1544 0 feedthrough
rlabel pdiffusion 773 -1544 773 -1544 0 cellNo=350
rlabel pdiffusion 780 -1544 780 -1544 0 feedthrough
rlabel pdiffusion 787 -1544 787 -1544 0 feedthrough
rlabel pdiffusion 794 -1544 794 -1544 0 feedthrough
rlabel pdiffusion 801 -1544 801 -1544 0 feedthrough
rlabel pdiffusion 808 -1544 808 -1544 0 feedthrough
rlabel pdiffusion 815 -1544 815 -1544 0 feedthrough
rlabel pdiffusion 822 -1544 822 -1544 0 feedthrough
rlabel pdiffusion 829 -1544 829 -1544 0 feedthrough
rlabel pdiffusion 836 -1544 836 -1544 0 feedthrough
rlabel pdiffusion 843 -1544 843 -1544 0 feedthrough
rlabel pdiffusion 850 -1544 850 -1544 0 feedthrough
rlabel pdiffusion 857 -1544 857 -1544 0 feedthrough
rlabel pdiffusion 864 -1544 864 -1544 0 feedthrough
rlabel pdiffusion 871 -1544 871 -1544 0 feedthrough
rlabel pdiffusion 878 -1544 878 -1544 0 feedthrough
rlabel pdiffusion 885 -1544 885 -1544 0 feedthrough
rlabel pdiffusion 892 -1544 892 -1544 0 feedthrough
rlabel pdiffusion 899 -1544 899 -1544 0 feedthrough
rlabel pdiffusion 906 -1544 906 -1544 0 feedthrough
rlabel pdiffusion 913 -1544 913 -1544 0 feedthrough
rlabel pdiffusion 920 -1544 920 -1544 0 feedthrough
rlabel pdiffusion 927 -1544 927 -1544 0 feedthrough
rlabel pdiffusion 934 -1544 934 -1544 0 feedthrough
rlabel pdiffusion 941 -1544 941 -1544 0 feedthrough
rlabel pdiffusion 948 -1544 948 -1544 0 feedthrough
rlabel pdiffusion 955 -1544 955 -1544 0 feedthrough
rlabel pdiffusion 962 -1544 962 -1544 0 feedthrough
rlabel pdiffusion 969 -1544 969 -1544 0 feedthrough
rlabel pdiffusion 976 -1544 976 -1544 0 feedthrough
rlabel pdiffusion 983 -1544 983 -1544 0 feedthrough
rlabel pdiffusion 990 -1544 990 -1544 0 feedthrough
rlabel pdiffusion 997 -1544 997 -1544 0 feedthrough
rlabel pdiffusion 1004 -1544 1004 -1544 0 feedthrough
rlabel pdiffusion 1011 -1544 1011 -1544 0 cellNo=956
rlabel pdiffusion 1018 -1544 1018 -1544 0 feedthrough
rlabel pdiffusion 1025 -1544 1025 -1544 0 feedthrough
rlabel pdiffusion 1032 -1544 1032 -1544 0 cellNo=386
rlabel pdiffusion 1039 -1544 1039 -1544 0 feedthrough
rlabel pdiffusion 1046 -1544 1046 -1544 0 feedthrough
rlabel pdiffusion 1060 -1544 1060 -1544 0 feedthrough
rlabel pdiffusion 1074 -1544 1074 -1544 0 feedthrough
rlabel pdiffusion 1095 -1544 1095 -1544 0 feedthrough
rlabel pdiffusion 3 -1633 3 -1633 0 cellNo=181
rlabel pdiffusion 10 -1633 10 -1633 0 feedthrough
rlabel pdiffusion 17 -1633 17 -1633 0 feedthrough
rlabel pdiffusion 24 -1633 24 -1633 0 feedthrough
rlabel pdiffusion 31 -1633 31 -1633 0 feedthrough
rlabel pdiffusion 38 -1633 38 -1633 0 feedthrough
rlabel pdiffusion 45 -1633 45 -1633 0 feedthrough
rlabel pdiffusion 52 -1633 52 -1633 0 feedthrough
rlabel pdiffusion 59 -1633 59 -1633 0 cellNo=206
rlabel pdiffusion 66 -1633 66 -1633 0 feedthrough
rlabel pdiffusion 73 -1633 73 -1633 0 feedthrough
rlabel pdiffusion 80 -1633 80 -1633 0 cellNo=421
rlabel pdiffusion 87 -1633 87 -1633 0 feedthrough
rlabel pdiffusion 94 -1633 94 -1633 0 cellNo=516
rlabel pdiffusion 101 -1633 101 -1633 0 feedthrough
rlabel pdiffusion 108 -1633 108 -1633 0 feedthrough
rlabel pdiffusion 115 -1633 115 -1633 0 feedthrough
rlabel pdiffusion 122 -1633 122 -1633 0 feedthrough
rlabel pdiffusion 129 -1633 129 -1633 0 feedthrough
rlabel pdiffusion 136 -1633 136 -1633 0 cellNo=282
rlabel pdiffusion 143 -1633 143 -1633 0 cellNo=593
rlabel pdiffusion 150 -1633 150 -1633 0 feedthrough
rlabel pdiffusion 157 -1633 157 -1633 0 feedthrough
rlabel pdiffusion 164 -1633 164 -1633 0 feedthrough
rlabel pdiffusion 171 -1633 171 -1633 0 feedthrough
rlabel pdiffusion 178 -1633 178 -1633 0 feedthrough
rlabel pdiffusion 185 -1633 185 -1633 0 cellNo=973
rlabel pdiffusion 192 -1633 192 -1633 0 cellNo=546
rlabel pdiffusion 199 -1633 199 -1633 0 cellNo=937
rlabel pdiffusion 206 -1633 206 -1633 0 feedthrough
rlabel pdiffusion 213 -1633 213 -1633 0 feedthrough
rlabel pdiffusion 220 -1633 220 -1633 0 cellNo=602
rlabel pdiffusion 227 -1633 227 -1633 0 cellNo=709
rlabel pdiffusion 234 -1633 234 -1633 0 feedthrough
rlabel pdiffusion 241 -1633 241 -1633 0 feedthrough
rlabel pdiffusion 248 -1633 248 -1633 0 cellNo=807
rlabel pdiffusion 255 -1633 255 -1633 0 feedthrough
rlabel pdiffusion 262 -1633 262 -1633 0 feedthrough
rlabel pdiffusion 269 -1633 269 -1633 0 feedthrough
rlabel pdiffusion 276 -1633 276 -1633 0 feedthrough
rlabel pdiffusion 283 -1633 283 -1633 0 feedthrough
rlabel pdiffusion 290 -1633 290 -1633 0 feedthrough
rlabel pdiffusion 297 -1633 297 -1633 0 feedthrough
rlabel pdiffusion 304 -1633 304 -1633 0 cellNo=894
rlabel pdiffusion 311 -1633 311 -1633 0 feedthrough
rlabel pdiffusion 318 -1633 318 -1633 0 feedthrough
rlabel pdiffusion 325 -1633 325 -1633 0 cellNo=237
rlabel pdiffusion 332 -1633 332 -1633 0 feedthrough
rlabel pdiffusion 339 -1633 339 -1633 0 feedthrough
rlabel pdiffusion 346 -1633 346 -1633 0 feedthrough
rlabel pdiffusion 353 -1633 353 -1633 0 cellNo=452
rlabel pdiffusion 360 -1633 360 -1633 0 feedthrough
rlabel pdiffusion 367 -1633 367 -1633 0 feedthrough
rlabel pdiffusion 374 -1633 374 -1633 0 cellNo=399
rlabel pdiffusion 381 -1633 381 -1633 0 feedthrough
rlabel pdiffusion 388 -1633 388 -1633 0 feedthrough
rlabel pdiffusion 395 -1633 395 -1633 0 feedthrough
rlabel pdiffusion 402 -1633 402 -1633 0 feedthrough
rlabel pdiffusion 409 -1633 409 -1633 0 feedthrough
rlabel pdiffusion 416 -1633 416 -1633 0 feedthrough
rlabel pdiffusion 423 -1633 423 -1633 0 cellNo=814
rlabel pdiffusion 430 -1633 430 -1633 0 feedthrough
rlabel pdiffusion 437 -1633 437 -1633 0 feedthrough
rlabel pdiffusion 444 -1633 444 -1633 0 cellNo=944
rlabel pdiffusion 451 -1633 451 -1633 0 feedthrough
rlabel pdiffusion 458 -1633 458 -1633 0 cellNo=577
rlabel pdiffusion 465 -1633 465 -1633 0 cellNo=124
rlabel pdiffusion 472 -1633 472 -1633 0 feedthrough
rlabel pdiffusion 479 -1633 479 -1633 0 feedthrough
rlabel pdiffusion 486 -1633 486 -1633 0 feedthrough
rlabel pdiffusion 493 -1633 493 -1633 0 feedthrough
rlabel pdiffusion 500 -1633 500 -1633 0 feedthrough
rlabel pdiffusion 507 -1633 507 -1633 0 feedthrough
rlabel pdiffusion 514 -1633 514 -1633 0 feedthrough
rlabel pdiffusion 521 -1633 521 -1633 0 feedthrough
rlabel pdiffusion 528 -1633 528 -1633 0 feedthrough
rlabel pdiffusion 535 -1633 535 -1633 0 cellNo=199
rlabel pdiffusion 542 -1633 542 -1633 0 feedthrough
rlabel pdiffusion 549 -1633 549 -1633 0 feedthrough
rlabel pdiffusion 556 -1633 556 -1633 0 feedthrough
rlabel pdiffusion 563 -1633 563 -1633 0 feedthrough
rlabel pdiffusion 570 -1633 570 -1633 0 cellNo=930
rlabel pdiffusion 577 -1633 577 -1633 0 feedthrough
rlabel pdiffusion 584 -1633 584 -1633 0 cellNo=484
rlabel pdiffusion 591 -1633 591 -1633 0 feedthrough
rlabel pdiffusion 598 -1633 598 -1633 0 feedthrough
rlabel pdiffusion 605 -1633 605 -1633 0 feedthrough
rlabel pdiffusion 612 -1633 612 -1633 0 cellNo=477
rlabel pdiffusion 619 -1633 619 -1633 0 feedthrough
rlabel pdiffusion 626 -1633 626 -1633 0 cellNo=566
rlabel pdiffusion 633 -1633 633 -1633 0 cellNo=355
rlabel pdiffusion 640 -1633 640 -1633 0 feedthrough
rlabel pdiffusion 647 -1633 647 -1633 0 feedthrough
rlabel pdiffusion 654 -1633 654 -1633 0 feedthrough
rlabel pdiffusion 661 -1633 661 -1633 0 feedthrough
rlabel pdiffusion 668 -1633 668 -1633 0 feedthrough
rlabel pdiffusion 675 -1633 675 -1633 0 cellNo=358
rlabel pdiffusion 682 -1633 682 -1633 0 cellNo=737
rlabel pdiffusion 689 -1633 689 -1633 0 feedthrough
rlabel pdiffusion 696 -1633 696 -1633 0 feedthrough
rlabel pdiffusion 703 -1633 703 -1633 0 feedthrough
rlabel pdiffusion 710 -1633 710 -1633 0 feedthrough
rlabel pdiffusion 717 -1633 717 -1633 0 feedthrough
rlabel pdiffusion 724 -1633 724 -1633 0 feedthrough
rlabel pdiffusion 731 -1633 731 -1633 0 feedthrough
rlabel pdiffusion 738 -1633 738 -1633 0 feedthrough
rlabel pdiffusion 745 -1633 745 -1633 0 feedthrough
rlabel pdiffusion 752 -1633 752 -1633 0 feedthrough
rlabel pdiffusion 759 -1633 759 -1633 0 feedthrough
rlabel pdiffusion 766 -1633 766 -1633 0 feedthrough
rlabel pdiffusion 773 -1633 773 -1633 0 feedthrough
rlabel pdiffusion 780 -1633 780 -1633 0 cellNo=595
rlabel pdiffusion 787 -1633 787 -1633 0 feedthrough
rlabel pdiffusion 794 -1633 794 -1633 0 feedthrough
rlabel pdiffusion 801 -1633 801 -1633 0 feedthrough
rlabel pdiffusion 808 -1633 808 -1633 0 feedthrough
rlabel pdiffusion 815 -1633 815 -1633 0 feedthrough
rlabel pdiffusion 822 -1633 822 -1633 0 feedthrough
rlabel pdiffusion 829 -1633 829 -1633 0 feedthrough
rlabel pdiffusion 836 -1633 836 -1633 0 feedthrough
rlabel pdiffusion 843 -1633 843 -1633 0 feedthrough
rlabel pdiffusion 850 -1633 850 -1633 0 feedthrough
rlabel pdiffusion 857 -1633 857 -1633 0 cellNo=918
rlabel pdiffusion 864 -1633 864 -1633 0 feedthrough
rlabel pdiffusion 871 -1633 871 -1633 0 feedthrough
rlabel pdiffusion 878 -1633 878 -1633 0 feedthrough
rlabel pdiffusion 885 -1633 885 -1633 0 feedthrough
rlabel pdiffusion 892 -1633 892 -1633 0 feedthrough
rlabel pdiffusion 899 -1633 899 -1633 0 feedthrough
rlabel pdiffusion 906 -1633 906 -1633 0 feedthrough
rlabel pdiffusion 913 -1633 913 -1633 0 feedthrough
rlabel pdiffusion 920 -1633 920 -1633 0 feedthrough
rlabel pdiffusion 927 -1633 927 -1633 0 feedthrough
rlabel pdiffusion 934 -1633 934 -1633 0 feedthrough
rlabel pdiffusion 941 -1633 941 -1633 0 feedthrough
rlabel pdiffusion 948 -1633 948 -1633 0 feedthrough
rlabel pdiffusion 955 -1633 955 -1633 0 feedthrough
rlabel pdiffusion 962 -1633 962 -1633 0 feedthrough
rlabel pdiffusion 969 -1633 969 -1633 0 feedthrough
rlabel pdiffusion 976 -1633 976 -1633 0 feedthrough
rlabel pdiffusion 983 -1633 983 -1633 0 feedthrough
rlabel pdiffusion 990 -1633 990 -1633 0 feedthrough
rlabel pdiffusion 997 -1633 997 -1633 0 feedthrough
rlabel pdiffusion 1004 -1633 1004 -1633 0 feedthrough
rlabel pdiffusion 1011 -1633 1011 -1633 0 feedthrough
rlabel pdiffusion 1018 -1633 1018 -1633 0 feedthrough
rlabel pdiffusion 1025 -1633 1025 -1633 0 feedthrough
rlabel pdiffusion 1032 -1633 1032 -1633 0 feedthrough
rlabel pdiffusion 1039 -1633 1039 -1633 0 feedthrough
rlabel pdiffusion 1046 -1633 1046 -1633 0 feedthrough
rlabel pdiffusion 1053 -1633 1053 -1633 0 feedthrough
rlabel pdiffusion 1060 -1633 1060 -1633 0 cellNo=591
rlabel pdiffusion 1067 -1633 1067 -1633 0 cellNo=933
rlabel pdiffusion 1074 -1633 1074 -1633 0 feedthrough
rlabel pdiffusion 1081 -1633 1081 -1633 0 feedthrough
rlabel pdiffusion 1088 -1633 1088 -1633 0 feedthrough
rlabel pdiffusion 1095 -1633 1095 -1633 0 feedthrough
rlabel pdiffusion 1102 -1633 1102 -1633 0 feedthrough
rlabel pdiffusion 1109 -1633 1109 -1633 0 feedthrough
rlabel pdiffusion 1116 -1633 1116 -1633 0 feedthrough
rlabel pdiffusion 24 -1718 24 -1718 0 feedthrough
rlabel pdiffusion 31 -1718 31 -1718 0 feedthrough
rlabel pdiffusion 38 -1718 38 -1718 0 feedthrough
rlabel pdiffusion 45 -1718 45 -1718 0 feedthrough
rlabel pdiffusion 52 -1718 52 -1718 0 cellNo=603
rlabel pdiffusion 59 -1718 59 -1718 0 feedthrough
rlabel pdiffusion 66 -1718 66 -1718 0 cellNo=724
rlabel pdiffusion 73 -1718 73 -1718 0 feedthrough
rlabel pdiffusion 80 -1718 80 -1718 0 feedthrough
rlabel pdiffusion 87 -1718 87 -1718 0 feedthrough
rlabel pdiffusion 94 -1718 94 -1718 0 feedthrough
rlabel pdiffusion 101 -1718 101 -1718 0 feedthrough
rlabel pdiffusion 108 -1718 108 -1718 0 feedthrough
rlabel pdiffusion 115 -1718 115 -1718 0 feedthrough
rlabel pdiffusion 122 -1718 122 -1718 0 feedthrough
rlabel pdiffusion 129 -1718 129 -1718 0 feedthrough
rlabel pdiffusion 136 -1718 136 -1718 0 feedthrough
rlabel pdiffusion 143 -1718 143 -1718 0 feedthrough
rlabel pdiffusion 150 -1718 150 -1718 0 feedthrough
rlabel pdiffusion 157 -1718 157 -1718 0 cellNo=657
rlabel pdiffusion 164 -1718 164 -1718 0 feedthrough
rlabel pdiffusion 171 -1718 171 -1718 0 feedthrough
rlabel pdiffusion 178 -1718 178 -1718 0 feedthrough
rlabel pdiffusion 185 -1718 185 -1718 0 feedthrough
rlabel pdiffusion 192 -1718 192 -1718 0 feedthrough
rlabel pdiffusion 199 -1718 199 -1718 0 feedthrough
rlabel pdiffusion 206 -1718 206 -1718 0 feedthrough
rlabel pdiffusion 213 -1718 213 -1718 0 feedthrough
rlabel pdiffusion 220 -1718 220 -1718 0 cellNo=298
rlabel pdiffusion 227 -1718 227 -1718 0 feedthrough
rlabel pdiffusion 234 -1718 234 -1718 0 feedthrough
rlabel pdiffusion 241 -1718 241 -1718 0 feedthrough
rlabel pdiffusion 248 -1718 248 -1718 0 feedthrough
rlabel pdiffusion 255 -1718 255 -1718 0 feedthrough
rlabel pdiffusion 262 -1718 262 -1718 0 feedthrough
rlabel pdiffusion 269 -1718 269 -1718 0 feedthrough
rlabel pdiffusion 276 -1718 276 -1718 0 feedthrough
rlabel pdiffusion 283 -1718 283 -1718 0 feedthrough
rlabel pdiffusion 290 -1718 290 -1718 0 feedthrough
rlabel pdiffusion 297 -1718 297 -1718 0 feedthrough
rlabel pdiffusion 304 -1718 304 -1718 0 cellNo=326
rlabel pdiffusion 311 -1718 311 -1718 0 cellNo=984
rlabel pdiffusion 318 -1718 318 -1718 0 feedthrough
rlabel pdiffusion 325 -1718 325 -1718 0 cellNo=893
rlabel pdiffusion 332 -1718 332 -1718 0 feedthrough
rlabel pdiffusion 339 -1718 339 -1718 0 cellNo=599
rlabel pdiffusion 346 -1718 346 -1718 0 feedthrough
rlabel pdiffusion 353 -1718 353 -1718 0 cellNo=912
rlabel pdiffusion 360 -1718 360 -1718 0 cellNo=836
rlabel pdiffusion 367 -1718 367 -1718 0 feedthrough
rlabel pdiffusion 374 -1718 374 -1718 0 cellNo=639
rlabel pdiffusion 381 -1718 381 -1718 0 cellNo=806
rlabel pdiffusion 388 -1718 388 -1718 0 feedthrough
rlabel pdiffusion 395 -1718 395 -1718 0 feedthrough
rlabel pdiffusion 402 -1718 402 -1718 0 feedthrough
rlabel pdiffusion 409 -1718 409 -1718 0 feedthrough
rlabel pdiffusion 416 -1718 416 -1718 0 feedthrough
rlabel pdiffusion 423 -1718 423 -1718 0 cellNo=543
rlabel pdiffusion 430 -1718 430 -1718 0 cellNo=151
rlabel pdiffusion 437 -1718 437 -1718 0 feedthrough
rlabel pdiffusion 444 -1718 444 -1718 0 feedthrough
rlabel pdiffusion 451 -1718 451 -1718 0 feedthrough
rlabel pdiffusion 458 -1718 458 -1718 0 feedthrough
rlabel pdiffusion 465 -1718 465 -1718 0 feedthrough
rlabel pdiffusion 472 -1718 472 -1718 0 feedthrough
rlabel pdiffusion 479 -1718 479 -1718 0 cellNo=138
rlabel pdiffusion 486 -1718 486 -1718 0 cellNo=294
rlabel pdiffusion 493 -1718 493 -1718 0 cellNo=902
rlabel pdiffusion 500 -1718 500 -1718 0 feedthrough
rlabel pdiffusion 507 -1718 507 -1718 0 feedthrough
rlabel pdiffusion 514 -1718 514 -1718 0 feedthrough
rlabel pdiffusion 521 -1718 521 -1718 0 cellNo=459
rlabel pdiffusion 528 -1718 528 -1718 0 cellNo=201
rlabel pdiffusion 535 -1718 535 -1718 0 feedthrough
rlabel pdiffusion 542 -1718 542 -1718 0 feedthrough
rlabel pdiffusion 549 -1718 549 -1718 0 feedthrough
rlabel pdiffusion 556 -1718 556 -1718 0 feedthrough
rlabel pdiffusion 563 -1718 563 -1718 0 feedthrough
rlabel pdiffusion 570 -1718 570 -1718 0 feedthrough
rlabel pdiffusion 577 -1718 577 -1718 0 cellNo=776
rlabel pdiffusion 584 -1718 584 -1718 0 cellNo=771
rlabel pdiffusion 591 -1718 591 -1718 0 feedthrough
rlabel pdiffusion 598 -1718 598 -1718 0 feedthrough
rlabel pdiffusion 605 -1718 605 -1718 0 cellNo=216
rlabel pdiffusion 612 -1718 612 -1718 0 feedthrough
rlabel pdiffusion 619 -1718 619 -1718 0 feedthrough
rlabel pdiffusion 626 -1718 626 -1718 0 feedthrough
rlabel pdiffusion 633 -1718 633 -1718 0 feedthrough
rlabel pdiffusion 640 -1718 640 -1718 0 feedthrough
rlabel pdiffusion 647 -1718 647 -1718 0 feedthrough
rlabel pdiffusion 654 -1718 654 -1718 0 cellNo=135
rlabel pdiffusion 661 -1718 661 -1718 0 cellNo=338
rlabel pdiffusion 668 -1718 668 -1718 0 feedthrough
rlabel pdiffusion 675 -1718 675 -1718 0 cellNo=58
rlabel pdiffusion 682 -1718 682 -1718 0 feedthrough
rlabel pdiffusion 689 -1718 689 -1718 0 cellNo=442
rlabel pdiffusion 696 -1718 696 -1718 0 feedthrough
rlabel pdiffusion 703 -1718 703 -1718 0 feedthrough
rlabel pdiffusion 710 -1718 710 -1718 0 feedthrough
rlabel pdiffusion 717 -1718 717 -1718 0 feedthrough
rlabel pdiffusion 724 -1718 724 -1718 0 feedthrough
rlabel pdiffusion 731 -1718 731 -1718 0 feedthrough
rlabel pdiffusion 738 -1718 738 -1718 0 feedthrough
rlabel pdiffusion 745 -1718 745 -1718 0 feedthrough
rlabel pdiffusion 752 -1718 752 -1718 0 cellNo=95
rlabel pdiffusion 759 -1718 759 -1718 0 cellNo=548
rlabel pdiffusion 766 -1718 766 -1718 0 feedthrough
rlabel pdiffusion 773 -1718 773 -1718 0 feedthrough
rlabel pdiffusion 780 -1718 780 -1718 0 feedthrough
rlabel pdiffusion 787 -1718 787 -1718 0 feedthrough
rlabel pdiffusion 794 -1718 794 -1718 0 feedthrough
rlabel pdiffusion 801 -1718 801 -1718 0 feedthrough
rlabel pdiffusion 808 -1718 808 -1718 0 feedthrough
rlabel pdiffusion 815 -1718 815 -1718 0 cellNo=683
rlabel pdiffusion 822 -1718 822 -1718 0 feedthrough
rlabel pdiffusion 829 -1718 829 -1718 0 feedthrough
rlabel pdiffusion 836 -1718 836 -1718 0 feedthrough
rlabel pdiffusion 843 -1718 843 -1718 0 feedthrough
rlabel pdiffusion 850 -1718 850 -1718 0 feedthrough
rlabel pdiffusion 857 -1718 857 -1718 0 feedthrough
rlabel pdiffusion 864 -1718 864 -1718 0 feedthrough
rlabel pdiffusion 871 -1718 871 -1718 0 feedthrough
rlabel pdiffusion 878 -1718 878 -1718 0 feedthrough
rlabel pdiffusion 885 -1718 885 -1718 0 feedthrough
rlabel pdiffusion 892 -1718 892 -1718 0 feedthrough
rlabel pdiffusion 899 -1718 899 -1718 0 feedthrough
rlabel pdiffusion 906 -1718 906 -1718 0 cellNo=938
rlabel pdiffusion 913 -1718 913 -1718 0 feedthrough
rlabel pdiffusion 920 -1718 920 -1718 0 feedthrough
rlabel pdiffusion 927 -1718 927 -1718 0 cellNo=978
rlabel pdiffusion 934 -1718 934 -1718 0 feedthrough
rlabel pdiffusion 941 -1718 941 -1718 0 feedthrough
rlabel pdiffusion 948 -1718 948 -1718 0 feedthrough
rlabel pdiffusion 955 -1718 955 -1718 0 feedthrough
rlabel pdiffusion 962 -1718 962 -1718 0 feedthrough
rlabel pdiffusion 969 -1718 969 -1718 0 feedthrough
rlabel pdiffusion 1067 -1718 1067 -1718 0 cellNo=633
rlabel pdiffusion 1095 -1718 1095 -1718 0 feedthrough
rlabel pdiffusion 3 -1809 3 -1809 0 feedthrough
rlabel pdiffusion 10 -1809 10 -1809 0 cellNo=742
rlabel pdiffusion 17 -1809 17 -1809 0 feedthrough
rlabel pdiffusion 24 -1809 24 -1809 0 feedthrough
rlabel pdiffusion 31 -1809 31 -1809 0 feedthrough
rlabel pdiffusion 38 -1809 38 -1809 0 feedthrough
rlabel pdiffusion 45 -1809 45 -1809 0 feedthrough
rlabel pdiffusion 52 -1809 52 -1809 0 feedthrough
rlabel pdiffusion 59 -1809 59 -1809 0 feedthrough
rlabel pdiffusion 66 -1809 66 -1809 0 feedthrough
rlabel pdiffusion 73 -1809 73 -1809 0 feedthrough
rlabel pdiffusion 80 -1809 80 -1809 0 feedthrough
rlabel pdiffusion 87 -1809 87 -1809 0 feedthrough
rlabel pdiffusion 94 -1809 94 -1809 0 cellNo=176
rlabel pdiffusion 101 -1809 101 -1809 0 cellNo=396
rlabel pdiffusion 108 -1809 108 -1809 0 cellNo=196
rlabel pdiffusion 115 -1809 115 -1809 0 cellNo=971
rlabel pdiffusion 122 -1809 122 -1809 0 feedthrough
rlabel pdiffusion 129 -1809 129 -1809 0 feedthrough
rlabel pdiffusion 136 -1809 136 -1809 0 cellNo=114
rlabel pdiffusion 143 -1809 143 -1809 0 feedthrough
rlabel pdiffusion 150 -1809 150 -1809 0 cellNo=180
rlabel pdiffusion 157 -1809 157 -1809 0 feedthrough
rlabel pdiffusion 164 -1809 164 -1809 0 feedthrough
rlabel pdiffusion 171 -1809 171 -1809 0 feedthrough
rlabel pdiffusion 178 -1809 178 -1809 0 feedthrough
rlabel pdiffusion 185 -1809 185 -1809 0 cellNo=614
rlabel pdiffusion 192 -1809 192 -1809 0 feedthrough
rlabel pdiffusion 199 -1809 199 -1809 0 cellNo=891
rlabel pdiffusion 206 -1809 206 -1809 0 cellNo=211
rlabel pdiffusion 213 -1809 213 -1809 0 feedthrough
rlabel pdiffusion 220 -1809 220 -1809 0 cellNo=972
rlabel pdiffusion 227 -1809 227 -1809 0 feedthrough
rlabel pdiffusion 234 -1809 234 -1809 0 feedthrough
rlabel pdiffusion 241 -1809 241 -1809 0 feedthrough
rlabel pdiffusion 248 -1809 248 -1809 0 cellNo=729
rlabel pdiffusion 255 -1809 255 -1809 0 feedthrough
rlabel pdiffusion 262 -1809 262 -1809 0 feedthrough
rlabel pdiffusion 269 -1809 269 -1809 0 feedthrough
rlabel pdiffusion 276 -1809 276 -1809 0 feedthrough
rlabel pdiffusion 283 -1809 283 -1809 0 feedthrough
rlabel pdiffusion 290 -1809 290 -1809 0 feedthrough
rlabel pdiffusion 297 -1809 297 -1809 0 feedthrough
rlabel pdiffusion 304 -1809 304 -1809 0 cellNo=648
rlabel pdiffusion 311 -1809 311 -1809 0 feedthrough
rlabel pdiffusion 318 -1809 318 -1809 0 feedthrough
rlabel pdiffusion 325 -1809 325 -1809 0 feedthrough
rlabel pdiffusion 332 -1809 332 -1809 0 feedthrough
rlabel pdiffusion 339 -1809 339 -1809 0 feedthrough
rlabel pdiffusion 346 -1809 346 -1809 0 cellNo=670
rlabel pdiffusion 353 -1809 353 -1809 0 cellNo=570
rlabel pdiffusion 360 -1809 360 -1809 0 feedthrough
rlabel pdiffusion 367 -1809 367 -1809 0 feedthrough
rlabel pdiffusion 374 -1809 374 -1809 0 feedthrough
rlabel pdiffusion 381 -1809 381 -1809 0 feedthrough
rlabel pdiffusion 388 -1809 388 -1809 0 feedthrough
rlabel pdiffusion 395 -1809 395 -1809 0 feedthrough
rlabel pdiffusion 402 -1809 402 -1809 0 feedthrough
rlabel pdiffusion 409 -1809 409 -1809 0 feedthrough
rlabel pdiffusion 416 -1809 416 -1809 0 cellNo=139
rlabel pdiffusion 423 -1809 423 -1809 0 cellNo=379
rlabel pdiffusion 430 -1809 430 -1809 0 cellNo=672
rlabel pdiffusion 437 -1809 437 -1809 0 feedthrough
rlabel pdiffusion 444 -1809 444 -1809 0 feedthrough
rlabel pdiffusion 451 -1809 451 -1809 0 feedthrough
rlabel pdiffusion 458 -1809 458 -1809 0 feedthrough
rlabel pdiffusion 465 -1809 465 -1809 0 feedthrough
rlabel pdiffusion 472 -1809 472 -1809 0 feedthrough
rlabel pdiffusion 479 -1809 479 -1809 0 feedthrough
rlabel pdiffusion 486 -1809 486 -1809 0 feedthrough
rlabel pdiffusion 493 -1809 493 -1809 0 feedthrough
rlabel pdiffusion 500 -1809 500 -1809 0 cellNo=664
rlabel pdiffusion 507 -1809 507 -1809 0 feedthrough
rlabel pdiffusion 514 -1809 514 -1809 0 feedthrough
rlabel pdiffusion 521 -1809 521 -1809 0 cellNo=553
rlabel pdiffusion 528 -1809 528 -1809 0 cellNo=580
rlabel pdiffusion 535 -1809 535 -1809 0 feedthrough
rlabel pdiffusion 542 -1809 542 -1809 0 feedthrough
rlabel pdiffusion 549 -1809 549 -1809 0 cellNo=694
rlabel pdiffusion 556 -1809 556 -1809 0 feedthrough
rlabel pdiffusion 563 -1809 563 -1809 0 feedthrough
rlabel pdiffusion 570 -1809 570 -1809 0 feedthrough
rlabel pdiffusion 577 -1809 577 -1809 0 feedthrough
rlabel pdiffusion 584 -1809 584 -1809 0 feedthrough
rlabel pdiffusion 591 -1809 591 -1809 0 feedthrough
rlabel pdiffusion 598 -1809 598 -1809 0 cellNo=951
rlabel pdiffusion 605 -1809 605 -1809 0 cellNo=896
rlabel pdiffusion 612 -1809 612 -1809 0 cellNo=539
rlabel pdiffusion 619 -1809 619 -1809 0 feedthrough
rlabel pdiffusion 626 -1809 626 -1809 0 cellNo=394
rlabel pdiffusion 633 -1809 633 -1809 0 feedthrough
rlabel pdiffusion 640 -1809 640 -1809 0 feedthrough
rlabel pdiffusion 647 -1809 647 -1809 0 feedthrough
rlabel pdiffusion 654 -1809 654 -1809 0 feedthrough
rlabel pdiffusion 661 -1809 661 -1809 0 feedthrough
rlabel pdiffusion 668 -1809 668 -1809 0 cellNo=197
rlabel pdiffusion 675 -1809 675 -1809 0 feedthrough
rlabel pdiffusion 682 -1809 682 -1809 0 feedthrough
rlabel pdiffusion 689 -1809 689 -1809 0 cellNo=149
rlabel pdiffusion 696 -1809 696 -1809 0 feedthrough
rlabel pdiffusion 703 -1809 703 -1809 0 feedthrough
rlabel pdiffusion 710 -1809 710 -1809 0 cellNo=675
rlabel pdiffusion 717 -1809 717 -1809 0 feedthrough
rlabel pdiffusion 724 -1809 724 -1809 0 feedthrough
rlabel pdiffusion 731 -1809 731 -1809 0 feedthrough
rlabel pdiffusion 738 -1809 738 -1809 0 feedthrough
rlabel pdiffusion 745 -1809 745 -1809 0 feedthrough
rlabel pdiffusion 752 -1809 752 -1809 0 feedthrough
rlabel pdiffusion 759 -1809 759 -1809 0 feedthrough
rlabel pdiffusion 766 -1809 766 -1809 0 cellNo=975
rlabel pdiffusion 773 -1809 773 -1809 0 feedthrough
rlabel pdiffusion 780 -1809 780 -1809 0 feedthrough
rlabel pdiffusion 787 -1809 787 -1809 0 feedthrough
rlabel pdiffusion 794 -1809 794 -1809 0 feedthrough
rlabel pdiffusion 801 -1809 801 -1809 0 feedthrough
rlabel pdiffusion 808 -1809 808 -1809 0 feedthrough
rlabel pdiffusion 815 -1809 815 -1809 0 feedthrough
rlabel pdiffusion 822 -1809 822 -1809 0 feedthrough
rlabel pdiffusion 829 -1809 829 -1809 0 feedthrough
rlabel pdiffusion 836 -1809 836 -1809 0 feedthrough
rlabel pdiffusion 843 -1809 843 -1809 0 feedthrough
rlabel pdiffusion 850 -1809 850 -1809 0 feedthrough
rlabel pdiffusion 857 -1809 857 -1809 0 feedthrough
rlabel pdiffusion 864 -1809 864 -1809 0 feedthrough
rlabel pdiffusion 871 -1809 871 -1809 0 feedthrough
rlabel pdiffusion 878 -1809 878 -1809 0 feedthrough
rlabel pdiffusion 885 -1809 885 -1809 0 feedthrough
rlabel pdiffusion 892 -1809 892 -1809 0 feedthrough
rlabel pdiffusion 899 -1809 899 -1809 0 feedthrough
rlabel pdiffusion 906 -1809 906 -1809 0 feedthrough
rlabel pdiffusion 913 -1809 913 -1809 0 feedthrough
rlabel pdiffusion 920 -1809 920 -1809 0 feedthrough
rlabel pdiffusion 927 -1809 927 -1809 0 feedthrough
rlabel pdiffusion 934 -1809 934 -1809 0 cellNo=136
rlabel pdiffusion 941 -1809 941 -1809 0 feedthrough
rlabel pdiffusion 948 -1809 948 -1809 0 feedthrough
rlabel pdiffusion 955 -1809 955 -1809 0 feedthrough
rlabel pdiffusion 962 -1809 962 -1809 0 feedthrough
rlabel pdiffusion 969 -1809 969 -1809 0 feedthrough
rlabel pdiffusion 976 -1809 976 -1809 0 feedthrough
rlabel pdiffusion 983 -1809 983 -1809 0 feedthrough
rlabel pdiffusion 990 -1809 990 -1809 0 feedthrough
rlabel pdiffusion 997 -1809 997 -1809 0 feedthrough
rlabel pdiffusion 1004 -1809 1004 -1809 0 feedthrough
rlabel pdiffusion 1011 -1809 1011 -1809 0 feedthrough
rlabel pdiffusion 1018 -1809 1018 -1809 0 feedthrough
rlabel pdiffusion 1025 -1809 1025 -1809 0 feedthrough
rlabel pdiffusion 1032 -1809 1032 -1809 0 feedthrough
rlabel pdiffusion 1039 -1809 1039 -1809 0 feedthrough
rlabel pdiffusion 1046 -1809 1046 -1809 0 feedthrough
rlabel pdiffusion 1053 -1809 1053 -1809 0 cellNo=269
rlabel pdiffusion 1060 -1809 1060 -1809 0 feedthrough
rlabel pdiffusion 1088 -1809 1088 -1809 0 feedthrough
rlabel pdiffusion 1095 -1809 1095 -1809 0 feedthrough
rlabel pdiffusion 3 -1900 3 -1900 0 cellNo=336
rlabel pdiffusion 10 -1900 10 -1900 0 feedthrough
rlabel pdiffusion 17 -1900 17 -1900 0 cellNo=564
rlabel pdiffusion 24 -1900 24 -1900 0 cellNo=997
rlabel pdiffusion 31 -1900 31 -1900 0 feedthrough
rlabel pdiffusion 38 -1900 38 -1900 0 cellNo=554
rlabel pdiffusion 45 -1900 45 -1900 0 cellNo=101
rlabel pdiffusion 52 -1900 52 -1900 0 cellNo=781
rlabel pdiffusion 59 -1900 59 -1900 0 feedthrough
rlabel pdiffusion 66 -1900 66 -1900 0 cellNo=334
rlabel pdiffusion 73 -1900 73 -1900 0 feedthrough
rlabel pdiffusion 80 -1900 80 -1900 0 cellNo=685
rlabel pdiffusion 87 -1900 87 -1900 0 feedthrough
rlabel pdiffusion 94 -1900 94 -1900 0 feedthrough
rlabel pdiffusion 101 -1900 101 -1900 0 feedthrough
rlabel pdiffusion 108 -1900 108 -1900 0 feedthrough
rlabel pdiffusion 115 -1900 115 -1900 0 cellNo=137
rlabel pdiffusion 122 -1900 122 -1900 0 cellNo=668
rlabel pdiffusion 129 -1900 129 -1900 0 feedthrough
rlabel pdiffusion 136 -1900 136 -1900 0 feedthrough
rlabel pdiffusion 143 -1900 143 -1900 0 feedthrough
rlabel pdiffusion 150 -1900 150 -1900 0 cellNo=887
rlabel pdiffusion 157 -1900 157 -1900 0 cellNo=919
rlabel pdiffusion 164 -1900 164 -1900 0 feedthrough
rlabel pdiffusion 171 -1900 171 -1900 0 feedthrough
rlabel pdiffusion 178 -1900 178 -1900 0 feedthrough
rlabel pdiffusion 185 -1900 185 -1900 0 feedthrough
rlabel pdiffusion 192 -1900 192 -1900 0 cellNo=783
rlabel pdiffusion 199 -1900 199 -1900 0 feedthrough
rlabel pdiffusion 206 -1900 206 -1900 0 feedthrough
rlabel pdiffusion 213 -1900 213 -1900 0 feedthrough
rlabel pdiffusion 220 -1900 220 -1900 0 cellNo=143
rlabel pdiffusion 227 -1900 227 -1900 0 feedthrough
rlabel pdiffusion 234 -1900 234 -1900 0 feedthrough
rlabel pdiffusion 241 -1900 241 -1900 0 feedthrough
rlabel pdiffusion 248 -1900 248 -1900 0 feedthrough
rlabel pdiffusion 255 -1900 255 -1900 0 feedthrough
rlabel pdiffusion 262 -1900 262 -1900 0 feedthrough
rlabel pdiffusion 269 -1900 269 -1900 0 feedthrough
rlabel pdiffusion 276 -1900 276 -1900 0 feedthrough
rlabel pdiffusion 283 -1900 283 -1900 0 feedthrough
rlabel pdiffusion 290 -1900 290 -1900 0 feedthrough
rlabel pdiffusion 297 -1900 297 -1900 0 feedthrough
rlabel pdiffusion 304 -1900 304 -1900 0 feedthrough
rlabel pdiffusion 311 -1900 311 -1900 0 feedthrough
rlabel pdiffusion 318 -1900 318 -1900 0 feedthrough
rlabel pdiffusion 325 -1900 325 -1900 0 feedthrough
rlabel pdiffusion 332 -1900 332 -1900 0 feedthrough
rlabel pdiffusion 339 -1900 339 -1900 0 feedthrough
rlabel pdiffusion 346 -1900 346 -1900 0 feedthrough
rlabel pdiffusion 353 -1900 353 -1900 0 feedthrough
rlabel pdiffusion 360 -1900 360 -1900 0 cellNo=498
rlabel pdiffusion 367 -1900 367 -1900 0 cellNo=304
rlabel pdiffusion 374 -1900 374 -1900 0 feedthrough
rlabel pdiffusion 381 -1900 381 -1900 0 feedthrough
rlabel pdiffusion 388 -1900 388 -1900 0 cellNo=118
rlabel pdiffusion 395 -1900 395 -1900 0 feedthrough
rlabel pdiffusion 402 -1900 402 -1900 0 feedthrough
rlabel pdiffusion 409 -1900 409 -1900 0 feedthrough
rlabel pdiffusion 416 -1900 416 -1900 0 cellNo=218
rlabel pdiffusion 423 -1900 423 -1900 0 feedthrough
rlabel pdiffusion 430 -1900 430 -1900 0 feedthrough
rlabel pdiffusion 437 -1900 437 -1900 0 feedthrough
rlabel pdiffusion 444 -1900 444 -1900 0 cellNo=716
rlabel pdiffusion 451 -1900 451 -1900 0 cellNo=629
rlabel pdiffusion 458 -1900 458 -1900 0 feedthrough
rlabel pdiffusion 465 -1900 465 -1900 0 feedthrough
rlabel pdiffusion 472 -1900 472 -1900 0 feedthrough
rlabel pdiffusion 479 -1900 479 -1900 0 cellNo=885
rlabel pdiffusion 486 -1900 486 -1900 0 cellNo=415
rlabel pdiffusion 493 -1900 493 -1900 0 feedthrough
rlabel pdiffusion 500 -1900 500 -1900 0 cellNo=965
rlabel pdiffusion 507 -1900 507 -1900 0 feedthrough
rlabel pdiffusion 514 -1900 514 -1900 0 feedthrough
rlabel pdiffusion 521 -1900 521 -1900 0 feedthrough
rlabel pdiffusion 528 -1900 528 -1900 0 cellNo=773
rlabel pdiffusion 535 -1900 535 -1900 0 feedthrough
rlabel pdiffusion 542 -1900 542 -1900 0 feedthrough
rlabel pdiffusion 549 -1900 549 -1900 0 cellNo=348
rlabel pdiffusion 556 -1900 556 -1900 0 cellNo=921
rlabel pdiffusion 563 -1900 563 -1900 0 feedthrough
rlabel pdiffusion 570 -1900 570 -1900 0 feedthrough
rlabel pdiffusion 577 -1900 577 -1900 0 feedthrough
rlabel pdiffusion 584 -1900 584 -1900 0 feedthrough
rlabel pdiffusion 591 -1900 591 -1900 0 feedthrough
rlabel pdiffusion 598 -1900 598 -1900 0 feedthrough
rlabel pdiffusion 605 -1900 605 -1900 0 feedthrough
rlabel pdiffusion 612 -1900 612 -1900 0 feedthrough
rlabel pdiffusion 619 -1900 619 -1900 0 cellNo=172
rlabel pdiffusion 626 -1900 626 -1900 0 feedthrough
rlabel pdiffusion 633 -1900 633 -1900 0 cellNo=434
rlabel pdiffusion 640 -1900 640 -1900 0 feedthrough
rlabel pdiffusion 647 -1900 647 -1900 0 feedthrough
rlabel pdiffusion 654 -1900 654 -1900 0 feedthrough
rlabel pdiffusion 661 -1900 661 -1900 0 feedthrough
rlabel pdiffusion 668 -1900 668 -1900 0 cellNo=523
rlabel pdiffusion 675 -1900 675 -1900 0 feedthrough
rlabel pdiffusion 682 -1900 682 -1900 0 feedthrough
rlabel pdiffusion 689 -1900 689 -1900 0 cellNo=3
rlabel pdiffusion 696 -1900 696 -1900 0 feedthrough
rlabel pdiffusion 703 -1900 703 -1900 0 feedthrough
rlabel pdiffusion 710 -1900 710 -1900 0 feedthrough
rlabel pdiffusion 717 -1900 717 -1900 0 feedthrough
rlabel pdiffusion 724 -1900 724 -1900 0 feedthrough
rlabel pdiffusion 731 -1900 731 -1900 0 cellNo=757
rlabel pdiffusion 738 -1900 738 -1900 0 feedthrough
rlabel pdiffusion 745 -1900 745 -1900 0 feedthrough
rlabel pdiffusion 752 -1900 752 -1900 0 feedthrough
rlabel pdiffusion 759 -1900 759 -1900 0 feedthrough
rlabel pdiffusion 766 -1900 766 -1900 0 feedthrough
rlabel pdiffusion 773 -1900 773 -1900 0 feedthrough
rlabel pdiffusion 780 -1900 780 -1900 0 feedthrough
rlabel pdiffusion 787 -1900 787 -1900 0 feedthrough
rlabel pdiffusion 794 -1900 794 -1900 0 feedthrough
rlabel pdiffusion 801 -1900 801 -1900 0 feedthrough
rlabel pdiffusion 808 -1900 808 -1900 0 feedthrough
rlabel pdiffusion 815 -1900 815 -1900 0 feedthrough
rlabel pdiffusion 822 -1900 822 -1900 0 feedthrough
rlabel pdiffusion 829 -1900 829 -1900 0 feedthrough
rlabel pdiffusion 836 -1900 836 -1900 0 feedthrough
rlabel pdiffusion 843 -1900 843 -1900 0 feedthrough
rlabel pdiffusion 850 -1900 850 -1900 0 feedthrough
rlabel pdiffusion 857 -1900 857 -1900 0 feedthrough
rlabel pdiffusion 864 -1900 864 -1900 0 feedthrough
rlabel pdiffusion 871 -1900 871 -1900 0 feedthrough
rlabel pdiffusion 878 -1900 878 -1900 0 feedthrough
rlabel pdiffusion 885 -1900 885 -1900 0 feedthrough
rlabel pdiffusion 892 -1900 892 -1900 0 feedthrough
rlabel pdiffusion 899 -1900 899 -1900 0 feedthrough
rlabel pdiffusion 906 -1900 906 -1900 0 feedthrough
rlabel pdiffusion 913 -1900 913 -1900 0 feedthrough
rlabel pdiffusion 920 -1900 920 -1900 0 feedthrough
rlabel pdiffusion 927 -1900 927 -1900 0 feedthrough
rlabel pdiffusion 934 -1900 934 -1900 0 feedthrough
rlabel pdiffusion 941 -1900 941 -1900 0 feedthrough
rlabel pdiffusion 948 -1900 948 -1900 0 feedthrough
rlabel pdiffusion 955 -1900 955 -1900 0 feedthrough
rlabel pdiffusion 962 -1900 962 -1900 0 feedthrough
rlabel pdiffusion 969 -1900 969 -1900 0 feedthrough
rlabel pdiffusion 976 -1900 976 -1900 0 feedthrough
rlabel pdiffusion 983 -1900 983 -1900 0 feedthrough
rlabel pdiffusion 990 -1900 990 -1900 0 feedthrough
rlabel pdiffusion 997 -1900 997 -1900 0 feedthrough
rlabel pdiffusion 1004 -1900 1004 -1900 0 feedthrough
rlabel pdiffusion 1011 -1900 1011 -1900 0 feedthrough
rlabel pdiffusion 1018 -1900 1018 -1900 0 feedthrough
rlabel pdiffusion 1025 -1900 1025 -1900 0 feedthrough
rlabel pdiffusion 1032 -1900 1032 -1900 0 feedthrough
rlabel pdiffusion 1039 -1900 1039 -1900 0 feedthrough
rlabel pdiffusion 1046 -1900 1046 -1900 0 feedthrough
rlabel pdiffusion 1053 -1900 1053 -1900 0 feedthrough
rlabel pdiffusion 1060 -1900 1060 -1900 0 feedthrough
rlabel pdiffusion 1067 -1900 1067 -1900 0 cellNo=319
rlabel pdiffusion 1074 -1900 1074 -1900 0 feedthrough
rlabel pdiffusion 1088 -1900 1088 -1900 0 feedthrough
rlabel pdiffusion 1102 -1900 1102 -1900 0 feedthrough
rlabel pdiffusion 3 -2005 3 -2005 0 cellNo=437
rlabel pdiffusion 10 -2005 10 -2005 0 feedthrough
rlabel pdiffusion 17 -2005 17 -2005 0 feedthrough
rlabel pdiffusion 24 -2005 24 -2005 0 cellNo=928
rlabel pdiffusion 31 -2005 31 -2005 0 cellNo=413
rlabel pdiffusion 38 -2005 38 -2005 0 feedthrough
rlabel pdiffusion 45 -2005 45 -2005 0 feedthrough
rlabel pdiffusion 52 -2005 52 -2005 0 cellNo=920
rlabel pdiffusion 59 -2005 59 -2005 0 cellNo=51
rlabel pdiffusion 66 -2005 66 -2005 0 feedthrough
rlabel pdiffusion 73 -2005 73 -2005 0 cellNo=915
rlabel pdiffusion 80 -2005 80 -2005 0 cellNo=713
rlabel pdiffusion 87 -2005 87 -2005 0 cellNo=340
rlabel pdiffusion 94 -2005 94 -2005 0 feedthrough
rlabel pdiffusion 101 -2005 101 -2005 0 feedthrough
rlabel pdiffusion 108 -2005 108 -2005 0 cellNo=1
rlabel pdiffusion 115 -2005 115 -2005 0 feedthrough
rlabel pdiffusion 122 -2005 122 -2005 0 feedthrough
rlabel pdiffusion 129 -2005 129 -2005 0 feedthrough
rlabel pdiffusion 136 -2005 136 -2005 0 cellNo=347
rlabel pdiffusion 143 -2005 143 -2005 0 feedthrough
rlabel pdiffusion 150 -2005 150 -2005 0 cellNo=410
rlabel pdiffusion 157 -2005 157 -2005 0 feedthrough
rlabel pdiffusion 164 -2005 164 -2005 0 feedthrough
rlabel pdiffusion 171 -2005 171 -2005 0 feedthrough
rlabel pdiffusion 178 -2005 178 -2005 0 cellNo=153
rlabel pdiffusion 185 -2005 185 -2005 0 feedthrough
rlabel pdiffusion 192 -2005 192 -2005 0 feedthrough
rlabel pdiffusion 199 -2005 199 -2005 0 feedthrough
rlabel pdiffusion 206 -2005 206 -2005 0 cellNo=865
rlabel pdiffusion 213 -2005 213 -2005 0 feedthrough
rlabel pdiffusion 220 -2005 220 -2005 0 cellNo=65
rlabel pdiffusion 227 -2005 227 -2005 0 cellNo=677
rlabel pdiffusion 234 -2005 234 -2005 0 feedthrough
rlabel pdiffusion 241 -2005 241 -2005 0 feedthrough
rlabel pdiffusion 248 -2005 248 -2005 0 feedthrough
rlabel pdiffusion 255 -2005 255 -2005 0 feedthrough
rlabel pdiffusion 262 -2005 262 -2005 0 feedthrough
rlabel pdiffusion 269 -2005 269 -2005 0 feedthrough
rlabel pdiffusion 276 -2005 276 -2005 0 feedthrough
rlabel pdiffusion 283 -2005 283 -2005 0 feedthrough
rlabel pdiffusion 290 -2005 290 -2005 0 feedthrough
rlabel pdiffusion 297 -2005 297 -2005 0 feedthrough
rlabel pdiffusion 304 -2005 304 -2005 0 feedthrough
rlabel pdiffusion 311 -2005 311 -2005 0 feedthrough
rlabel pdiffusion 318 -2005 318 -2005 0 feedthrough
rlabel pdiffusion 325 -2005 325 -2005 0 feedthrough
rlabel pdiffusion 332 -2005 332 -2005 0 feedthrough
rlabel pdiffusion 339 -2005 339 -2005 0 feedthrough
rlabel pdiffusion 346 -2005 346 -2005 0 cellNo=426
rlabel pdiffusion 353 -2005 353 -2005 0 feedthrough
rlabel pdiffusion 360 -2005 360 -2005 0 feedthrough
rlabel pdiffusion 367 -2005 367 -2005 0 cellNo=4
rlabel pdiffusion 374 -2005 374 -2005 0 cellNo=534
rlabel pdiffusion 381 -2005 381 -2005 0 feedthrough
rlabel pdiffusion 388 -2005 388 -2005 0 feedthrough
rlabel pdiffusion 395 -2005 395 -2005 0 feedthrough
rlabel pdiffusion 402 -2005 402 -2005 0 feedthrough
rlabel pdiffusion 409 -2005 409 -2005 0 cellNo=823
rlabel pdiffusion 416 -2005 416 -2005 0 feedthrough
rlabel pdiffusion 423 -2005 423 -2005 0 feedthrough
rlabel pdiffusion 430 -2005 430 -2005 0 feedthrough
rlabel pdiffusion 437 -2005 437 -2005 0 cellNo=35
rlabel pdiffusion 444 -2005 444 -2005 0 feedthrough
rlabel pdiffusion 451 -2005 451 -2005 0 feedthrough
rlabel pdiffusion 458 -2005 458 -2005 0 feedthrough
rlabel pdiffusion 465 -2005 465 -2005 0 feedthrough
rlabel pdiffusion 472 -2005 472 -2005 0 feedthrough
rlabel pdiffusion 479 -2005 479 -2005 0 feedthrough
rlabel pdiffusion 486 -2005 486 -2005 0 feedthrough
rlabel pdiffusion 493 -2005 493 -2005 0 feedthrough
rlabel pdiffusion 500 -2005 500 -2005 0 feedthrough
rlabel pdiffusion 507 -2005 507 -2005 0 feedthrough
rlabel pdiffusion 514 -2005 514 -2005 0 cellNo=805
rlabel pdiffusion 521 -2005 521 -2005 0 feedthrough
rlabel pdiffusion 528 -2005 528 -2005 0 cellNo=325
rlabel pdiffusion 535 -2005 535 -2005 0 feedthrough
rlabel pdiffusion 542 -2005 542 -2005 0 feedthrough
rlabel pdiffusion 549 -2005 549 -2005 0 feedthrough
rlabel pdiffusion 556 -2005 556 -2005 0 feedthrough
rlabel pdiffusion 563 -2005 563 -2005 0 feedthrough
rlabel pdiffusion 570 -2005 570 -2005 0 feedthrough
rlabel pdiffusion 577 -2005 577 -2005 0 feedthrough
rlabel pdiffusion 584 -2005 584 -2005 0 feedthrough
rlabel pdiffusion 591 -2005 591 -2005 0 cellNo=134
rlabel pdiffusion 598 -2005 598 -2005 0 feedthrough
rlabel pdiffusion 605 -2005 605 -2005 0 feedthrough
rlabel pdiffusion 612 -2005 612 -2005 0 feedthrough
rlabel pdiffusion 619 -2005 619 -2005 0 cellNo=870
rlabel pdiffusion 626 -2005 626 -2005 0 feedthrough
rlabel pdiffusion 633 -2005 633 -2005 0 cellNo=385
rlabel pdiffusion 640 -2005 640 -2005 0 feedthrough
rlabel pdiffusion 647 -2005 647 -2005 0 cellNo=16
rlabel pdiffusion 654 -2005 654 -2005 0 feedthrough
rlabel pdiffusion 661 -2005 661 -2005 0 feedthrough
rlabel pdiffusion 668 -2005 668 -2005 0 feedthrough
rlabel pdiffusion 675 -2005 675 -2005 0 feedthrough
rlabel pdiffusion 682 -2005 682 -2005 0 feedthrough
rlabel pdiffusion 689 -2005 689 -2005 0 feedthrough
rlabel pdiffusion 696 -2005 696 -2005 0 feedthrough
rlabel pdiffusion 703 -2005 703 -2005 0 feedthrough
rlabel pdiffusion 710 -2005 710 -2005 0 feedthrough
rlabel pdiffusion 717 -2005 717 -2005 0 feedthrough
rlabel pdiffusion 724 -2005 724 -2005 0 feedthrough
rlabel pdiffusion 731 -2005 731 -2005 0 feedthrough
rlabel pdiffusion 738 -2005 738 -2005 0 feedthrough
rlabel pdiffusion 745 -2005 745 -2005 0 cellNo=733
rlabel pdiffusion 752 -2005 752 -2005 0 feedthrough
rlabel pdiffusion 759 -2005 759 -2005 0 feedthrough
rlabel pdiffusion 766 -2005 766 -2005 0 cellNo=429
rlabel pdiffusion 773 -2005 773 -2005 0 feedthrough
rlabel pdiffusion 780 -2005 780 -2005 0 cellNo=775
rlabel pdiffusion 787 -2005 787 -2005 0 feedthrough
rlabel pdiffusion 794 -2005 794 -2005 0 feedthrough
rlabel pdiffusion 801 -2005 801 -2005 0 feedthrough
rlabel pdiffusion 808 -2005 808 -2005 0 feedthrough
rlabel pdiffusion 815 -2005 815 -2005 0 feedthrough
rlabel pdiffusion 822 -2005 822 -2005 0 feedthrough
rlabel pdiffusion 829 -2005 829 -2005 0 feedthrough
rlabel pdiffusion 836 -2005 836 -2005 0 feedthrough
rlabel pdiffusion 843 -2005 843 -2005 0 feedthrough
rlabel pdiffusion 850 -2005 850 -2005 0 feedthrough
rlabel pdiffusion 857 -2005 857 -2005 0 feedthrough
rlabel pdiffusion 864 -2005 864 -2005 0 feedthrough
rlabel pdiffusion 871 -2005 871 -2005 0 feedthrough
rlabel pdiffusion 878 -2005 878 -2005 0 feedthrough
rlabel pdiffusion 885 -2005 885 -2005 0 feedthrough
rlabel pdiffusion 892 -2005 892 -2005 0 feedthrough
rlabel pdiffusion 899 -2005 899 -2005 0 feedthrough
rlabel pdiffusion 906 -2005 906 -2005 0 feedthrough
rlabel pdiffusion 913 -2005 913 -2005 0 feedthrough
rlabel pdiffusion 920 -2005 920 -2005 0 feedthrough
rlabel pdiffusion 927 -2005 927 -2005 0 cellNo=445
rlabel pdiffusion 934 -2005 934 -2005 0 feedthrough
rlabel pdiffusion 941 -2005 941 -2005 0 feedthrough
rlabel pdiffusion 948 -2005 948 -2005 0 feedthrough
rlabel pdiffusion 955 -2005 955 -2005 0 feedthrough
rlabel pdiffusion 962 -2005 962 -2005 0 feedthrough
rlabel pdiffusion 969 -2005 969 -2005 0 feedthrough
rlabel pdiffusion 976 -2005 976 -2005 0 feedthrough
rlabel pdiffusion 983 -2005 983 -2005 0 feedthrough
rlabel pdiffusion 990 -2005 990 -2005 0 feedthrough
rlabel pdiffusion 997 -2005 997 -2005 0 feedthrough
rlabel pdiffusion 1004 -2005 1004 -2005 0 feedthrough
rlabel pdiffusion 1011 -2005 1011 -2005 0 feedthrough
rlabel pdiffusion 1018 -2005 1018 -2005 0 feedthrough
rlabel pdiffusion 1025 -2005 1025 -2005 0 feedthrough
rlabel pdiffusion 1032 -2005 1032 -2005 0 feedthrough
rlabel pdiffusion 1039 -2005 1039 -2005 0 feedthrough
rlabel pdiffusion 1046 -2005 1046 -2005 0 feedthrough
rlabel pdiffusion 1053 -2005 1053 -2005 0 feedthrough
rlabel pdiffusion 1060 -2005 1060 -2005 0 feedthrough
rlabel pdiffusion 1067 -2005 1067 -2005 0 feedthrough
rlabel pdiffusion 1074 -2005 1074 -2005 0 feedthrough
rlabel pdiffusion 1081 -2005 1081 -2005 0 feedthrough
rlabel pdiffusion 1088 -2005 1088 -2005 0 feedthrough
rlabel pdiffusion 1095 -2005 1095 -2005 0 cellNo=791
rlabel pdiffusion 1102 -2005 1102 -2005 0 cellNo=837
rlabel pdiffusion 1109 -2005 1109 -2005 0 feedthrough
rlabel pdiffusion 1116 -2005 1116 -2005 0 feedthrough
rlabel pdiffusion 3 -2118 3 -2118 0 feedthrough
rlabel pdiffusion 10 -2118 10 -2118 0 feedthrough
rlabel pdiffusion 17 -2118 17 -2118 0 feedthrough
rlabel pdiffusion 24 -2118 24 -2118 0 feedthrough
rlabel pdiffusion 31 -2118 31 -2118 0 feedthrough
rlabel pdiffusion 38 -2118 38 -2118 0 feedthrough
rlabel pdiffusion 45 -2118 45 -2118 0 feedthrough
rlabel pdiffusion 52 -2118 52 -2118 0 feedthrough
rlabel pdiffusion 59 -2118 59 -2118 0 cellNo=957
rlabel pdiffusion 66 -2118 66 -2118 0 feedthrough
rlabel pdiffusion 73 -2118 73 -2118 0 cellNo=898
rlabel pdiffusion 80 -2118 80 -2118 0 cellNo=778
rlabel pdiffusion 87 -2118 87 -2118 0 cellNo=378
rlabel pdiffusion 94 -2118 94 -2118 0 cellNo=707
rlabel pdiffusion 101 -2118 101 -2118 0 feedthrough
rlabel pdiffusion 108 -2118 108 -2118 0 cellNo=128
rlabel pdiffusion 115 -2118 115 -2118 0 cellNo=505
rlabel pdiffusion 122 -2118 122 -2118 0 cellNo=763
rlabel pdiffusion 129 -2118 129 -2118 0 feedthrough
rlabel pdiffusion 136 -2118 136 -2118 0 cellNo=939
rlabel pdiffusion 143 -2118 143 -2118 0 feedthrough
rlabel pdiffusion 150 -2118 150 -2118 0 cellNo=424
rlabel pdiffusion 157 -2118 157 -2118 0 feedthrough
rlabel pdiffusion 164 -2118 164 -2118 0 feedthrough
rlabel pdiffusion 171 -2118 171 -2118 0 feedthrough
rlabel pdiffusion 178 -2118 178 -2118 0 feedthrough
rlabel pdiffusion 185 -2118 185 -2118 0 feedthrough
rlabel pdiffusion 192 -2118 192 -2118 0 feedthrough
rlabel pdiffusion 199 -2118 199 -2118 0 feedthrough
rlabel pdiffusion 206 -2118 206 -2118 0 feedthrough
rlabel pdiffusion 213 -2118 213 -2118 0 feedthrough
rlabel pdiffusion 220 -2118 220 -2118 0 cellNo=829
rlabel pdiffusion 227 -2118 227 -2118 0 feedthrough
rlabel pdiffusion 234 -2118 234 -2118 0 feedthrough
rlabel pdiffusion 241 -2118 241 -2118 0 feedthrough
rlabel pdiffusion 248 -2118 248 -2118 0 feedthrough
rlabel pdiffusion 255 -2118 255 -2118 0 feedthrough
rlabel pdiffusion 262 -2118 262 -2118 0 feedthrough
rlabel pdiffusion 269 -2118 269 -2118 0 feedthrough
rlabel pdiffusion 276 -2118 276 -2118 0 feedthrough
rlabel pdiffusion 283 -2118 283 -2118 0 feedthrough
rlabel pdiffusion 290 -2118 290 -2118 0 cellNo=267
rlabel pdiffusion 297 -2118 297 -2118 0 feedthrough
rlabel pdiffusion 304 -2118 304 -2118 0 feedthrough
rlabel pdiffusion 311 -2118 311 -2118 0 feedthrough
rlabel pdiffusion 318 -2118 318 -2118 0 feedthrough
rlabel pdiffusion 325 -2118 325 -2118 0 feedthrough
rlabel pdiffusion 332 -2118 332 -2118 0 feedthrough
rlabel pdiffusion 339 -2118 339 -2118 0 cellNo=839
rlabel pdiffusion 346 -2118 346 -2118 0 feedthrough
rlabel pdiffusion 353 -2118 353 -2118 0 cellNo=522
rlabel pdiffusion 360 -2118 360 -2118 0 feedthrough
rlabel pdiffusion 367 -2118 367 -2118 0 feedthrough
rlabel pdiffusion 374 -2118 374 -2118 0 feedthrough
rlabel pdiffusion 381 -2118 381 -2118 0 feedthrough
rlabel pdiffusion 388 -2118 388 -2118 0 feedthrough
rlabel pdiffusion 395 -2118 395 -2118 0 feedthrough
rlabel pdiffusion 402 -2118 402 -2118 0 feedthrough
rlabel pdiffusion 409 -2118 409 -2118 0 cellNo=531
rlabel pdiffusion 416 -2118 416 -2118 0 cellNo=482
rlabel pdiffusion 423 -2118 423 -2118 0 feedthrough
rlabel pdiffusion 430 -2118 430 -2118 0 feedthrough
rlabel pdiffusion 437 -2118 437 -2118 0 feedthrough
rlabel pdiffusion 444 -2118 444 -2118 0 feedthrough
rlabel pdiffusion 451 -2118 451 -2118 0 cellNo=607
rlabel pdiffusion 458 -2118 458 -2118 0 cellNo=497
rlabel pdiffusion 465 -2118 465 -2118 0 feedthrough
rlabel pdiffusion 472 -2118 472 -2118 0 feedthrough
rlabel pdiffusion 479 -2118 479 -2118 0 feedthrough
rlabel pdiffusion 486 -2118 486 -2118 0 feedthrough
rlabel pdiffusion 493 -2118 493 -2118 0 feedthrough
rlabel pdiffusion 500 -2118 500 -2118 0 cellNo=792
rlabel pdiffusion 507 -2118 507 -2118 0 feedthrough
rlabel pdiffusion 514 -2118 514 -2118 0 feedthrough
rlabel pdiffusion 521 -2118 521 -2118 0 feedthrough
rlabel pdiffusion 528 -2118 528 -2118 0 cellNo=945
rlabel pdiffusion 535 -2118 535 -2118 0 feedthrough
rlabel pdiffusion 542 -2118 542 -2118 0 feedthrough
rlabel pdiffusion 549 -2118 549 -2118 0 cellNo=741
rlabel pdiffusion 556 -2118 556 -2118 0 feedthrough
rlabel pdiffusion 563 -2118 563 -2118 0 feedthrough
rlabel pdiffusion 570 -2118 570 -2118 0 cellNo=495
rlabel pdiffusion 577 -2118 577 -2118 0 cellNo=690
rlabel pdiffusion 584 -2118 584 -2118 0 feedthrough
rlabel pdiffusion 591 -2118 591 -2118 0 feedthrough
rlabel pdiffusion 598 -2118 598 -2118 0 feedthrough
rlabel pdiffusion 605 -2118 605 -2118 0 feedthrough
rlabel pdiffusion 612 -2118 612 -2118 0 cellNo=857
rlabel pdiffusion 619 -2118 619 -2118 0 feedthrough
rlabel pdiffusion 626 -2118 626 -2118 0 cellNo=485
rlabel pdiffusion 633 -2118 633 -2118 0 feedthrough
rlabel pdiffusion 640 -2118 640 -2118 0 cellNo=979
rlabel pdiffusion 647 -2118 647 -2118 0 feedthrough
rlabel pdiffusion 654 -2118 654 -2118 0 cellNo=530
rlabel pdiffusion 661 -2118 661 -2118 0 feedthrough
rlabel pdiffusion 668 -2118 668 -2118 0 feedthrough
rlabel pdiffusion 675 -2118 675 -2118 0 feedthrough
rlabel pdiffusion 682 -2118 682 -2118 0 feedthrough
rlabel pdiffusion 689 -2118 689 -2118 0 cellNo=341
rlabel pdiffusion 696 -2118 696 -2118 0 feedthrough
rlabel pdiffusion 703 -2118 703 -2118 0 feedthrough
rlabel pdiffusion 710 -2118 710 -2118 0 feedthrough
rlabel pdiffusion 717 -2118 717 -2118 0 feedthrough
rlabel pdiffusion 724 -2118 724 -2118 0 feedthrough
rlabel pdiffusion 731 -2118 731 -2118 0 feedthrough
rlabel pdiffusion 738 -2118 738 -2118 0 cellNo=493
rlabel pdiffusion 745 -2118 745 -2118 0 feedthrough
rlabel pdiffusion 752 -2118 752 -2118 0 feedthrough
rlabel pdiffusion 759 -2118 759 -2118 0 cellNo=630
rlabel pdiffusion 766 -2118 766 -2118 0 feedthrough
rlabel pdiffusion 773 -2118 773 -2118 0 feedthrough
rlabel pdiffusion 780 -2118 780 -2118 0 feedthrough
rlabel pdiffusion 787 -2118 787 -2118 0 feedthrough
rlabel pdiffusion 794 -2118 794 -2118 0 feedthrough
rlabel pdiffusion 801 -2118 801 -2118 0 feedthrough
rlabel pdiffusion 808 -2118 808 -2118 0 feedthrough
rlabel pdiffusion 815 -2118 815 -2118 0 feedthrough
rlabel pdiffusion 822 -2118 822 -2118 0 feedthrough
rlabel pdiffusion 829 -2118 829 -2118 0 feedthrough
rlabel pdiffusion 836 -2118 836 -2118 0 feedthrough
rlabel pdiffusion 843 -2118 843 -2118 0 feedthrough
rlabel pdiffusion 850 -2118 850 -2118 0 feedthrough
rlabel pdiffusion 857 -2118 857 -2118 0 feedthrough
rlabel pdiffusion 864 -2118 864 -2118 0 feedthrough
rlabel pdiffusion 871 -2118 871 -2118 0 feedthrough
rlabel pdiffusion 878 -2118 878 -2118 0 feedthrough
rlabel pdiffusion 885 -2118 885 -2118 0 feedthrough
rlabel pdiffusion 892 -2118 892 -2118 0 feedthrough
rlabel pdiffusion 899 -2118 899 -2118 0 feedthrough
rlabel pdiffusion 906 -2118 906 -2118 0 feedthrough
rlabel pdiffusion 913 -2118 913 -2118 0 feedthrough
rlabel pdiffusion 920 -2118 920 -2118 0 feedthrough
rlabel pdiffusion 927 -2118 927 -2118 0 feedthrough
rlabel pdiffusion 934 -2118 934 -2118 0 feedthrough
rlabel pdiffusion 941 -2118 941 -2118 0 cellNo=473
rlabel pdiffusion 948 -2118 948 -2118 0 feedthrough
rlabel pdiffusion 955 -2118 955 -2118 0 feedthrough
rlabel pdiffusion 962 -2118 962 -2118 0 feedthrough
rlabel pdiffusion 969 -2118 969 -2118 0 feedthrough
rlabel pdiffusion 976 -2118 976 -2118 0 feedthrough
rlabel pdiffusion 983 -2118 983 -2118 0 feedthrough
rlabel pdiffusion 990 -2118 990 -2118 0 feedthrough
rlabel pdiffusion 997 -2118 997 -2118 0 feedthrough
rlabel pdiffusion 1004 -2118 1004 -2118 0 feedthrough
rlabel pdiffusion 1011 -2118 1011 -2118 0 feedthrough
rlabel pdiffusion 1018 -2118 1018 -2118 0 feedthrough
rlabel pdiffusion 1025 -2118 1025 -2118 0 feedthrough
rlabel pdiffusion 1032 -2118 1032 -2118 0 feedthrough
rlabel pdiffusion 1039 -2118 1039 -2118 0 feedthrough
rlabel pdiffusion 1046 -2118 1046 -2118 0 feedthrough
rlabel pdiffusion 1053 -2118 1053 -2118 0 feedthrough
rlabel pdiffusion 1060 -2118 1060 -2118 0 feedthrough
rlabel pdiffusion 1067 -2118 1067 -2118 0 feedthrough
rlabel pdiffusion 1074 -2118 1074 -2118 0 feedthrough
rlabel pdiffusion 1081 -2118 1081 -2118 0 feedthrough
rlabel pdiffusion 1088 -2118 1088 -2118 0 feedthrough
rlabel pdiffusion 1095 -2118 1095 -2118 0 feedthrough
rlabel pdiffusion 1102 -2118 1102 -2118 0 cellNo=363
rlabel pdiffusion 1109 -2118 1109 -2118 0 feedthrough
rlabel pdiffusion 1116 -2118 1116 -2118 0 feedthrough
rlabel pdiffusion 1123 -2118 1123 -2118 0 feedthrough
rlabel pdiffusion 3 -2213 3 -2213 0 feedthrough
rlabel pdiffusion 10 -2213 10 -2213 0 feedthrough
rlabel pdiffusion 17 -2213 17 -2213 0 feedthrough
rlabel pdiffusion 24 -2213 24 -2213 0 feedthrough
rlabel pdiffusion 31 -2213 31 -2213 0 cellNo=84
rlabel pdiffusion 38 -2213 38 -2213 0 cellNo=749
rlabel pdiffusion 45 -2213 45 -2213 0 feedthrough
rlabel pdiffusion 52 -2213 52 -2213 0 feedthrough
rlabel pdiffusion 59 -2213 59 -2213 0 feedthrough
rlabel pdiffusion 66 -2213 66 -2213 0 feedthrough
rlabel pdiffusion 73 -2213 73 -2213 0 cellNo=910
rlabel pdiffusion 80 -2213 80 -2213 0 feedthrough
rlabel pdiffusion 87 -2213 87 -2213 0 feedthrough
rlabel pdiffusion 94 -2213 94 -2213 0 feedthrough
rlabel pdiffusion 101 -2213 101 -2213 0 feedthrough
rlabel pdiffusion 108 -2213 108 -2213 0 feedthrough
rlabel pdiffusion 115 -2213 115 -2213 0 feedthrough
rlabel pdiffusion 122 -2213 122 -2213 0 cellNo=416
rlabel pdiffusion 129 -2213 129 -2213 0 feedthrough
rlabel pdiffusion 136 -2213 136 -2213 0 feedthrough
rlabel pdiffusion 143 -2213 143 -2213 0 feedthrough
rlabel pdiffusion 150 -2213 150 -2213 0 feedthrough
rlabel pdiffusion 157 -2213 157 -2213 0 feedthrough
rlabel pdiffusion 164 -2213 164 -2213 0 cellNo=402
rlabel pdiffusion 171 -2213 171 -2213 0 cellNo=936
rlabel pdiffusion 178 -2213 178 -2213 0 cellNo=533
rlabel pdiffusion 185 -2213 185 -2213 0 cellNo=203
rlabel pdiffusion 192 -2213 192 -2213 0 cellNo=454
rlabel pdiffusion 199 -2213 199 -2213 0 feedthrough
rlabel pdiffusion 206 -2213 206 -2213 0 cellNo=948
rlabel pdiffusion 213 -2213 213 -2213 0 feedthrough
rlabel pdiffusion 220 -2213 220 -2213 0 feedthrough
rlabel pdiffusion 227 -2213 227 -2213 0 feedthrough
rlabel pdiffusion 234 -2213 234 -2213 0 feedthrough
rlabel pdiffusion 241 -2213 241 -2213 0 feedthrough
rlabel pdiffusion 248 -2213 248 -2213 0 feedthrough
rlabel pdiffusion 255 -2213 255 -2213 0 feedthrough
rlabel pdiffusion 262 -2213 262 -2213 0 feedthrough
rlabel pdiffusion 269 -2213 269 -2213 0 feedthrough
rlabel pdiffusion 276 -2213 276 -2213 0 feedthrough
rlabel pdiffusion 283 -2213 283 -2213 0 feedthrough
rlabel pdiffusion 290 -2213 290 -2213 0 feedthrough
rlabel pdiffusion 297 -2213 297 -2213 0 feedthrough
rlabel pdiffusion 304 -2213 304 -2213 0 feedthrough
rlabel pdiffusion 311 -2213 311 -2213 0 feedthrough
rlabel pdiffusion 318 -2213 318 -2213 0 cellNo=359
rlabel pdiffusion 325 -2213 325 -2213 0 feedthrough
rlabel pdiffusion 332 -2213 332 -2213 0 feedthrough
rlabel pdiffusion 339 -2213 339 -2213 0 cellNo=813
rlabel pdiffusion 346 -2213 346 -2213 0 feedthrough
rlabel pdiffusion 353 -2213 353 -2213 0 cellNo=923
rlabel pdiffusion 360 -2213 360 -2213 0 feedthrough
rlabel pdiffusion 367 -2213 367 -2213 0 feedthrough
rlabel pdiffusion 374 -2213 374 -2213 0 cellNo=535
rlabel pdiffusion 381 -2213 381 -2213 0 feedthrough
rlabel pdiffusion 388 -2213 388 -2213 0 feedthrough
rlabel pdiffusion 395 -2213 395 -2213 0 cellNo=834
rlabel pdiffusion 402 -2213 402 -2213 0 feedthrough
rlabel pdiffusion 409 -2213 409 -2213 0 feedthrough
rlabel pdiffusion 416 -2213 416 -2213 0 feedthrough
rlabel pdiffusion 423 -2213 423 -2213 0 feedthrough
rlabel pdiffusion 430 -2213 430 -2213 0 cellNo=388
rlabel pdiffusion 437 -2213 437 -2213 0 cellNo=587
rlabel pdiffusion 444 -2213 444 -2213 0 feedthrough
rlabel pdiffusion 451 -2213 451 -2213 0 feedthrough
rlabel pdiffusion 458 -2213 458 -2213 0 feedthrough
rlabel pdiffusion 465 -2213 465 -2213 0 feedthrough
rlabel pdiffusion 472 -2213 472 -2213 0 feedthrough
rlabel pdiffusion 479 -2213 479 -2213 0 feedthrough
rlabel pdiffusion 486 -2213 486 -2213 0 feedthrough
rlabel pdiffusion 493 -2213 493 -2213 0 feedthrough
rlabel pdiffusion 500 -2213 500 -2213 0 cellNo=40
rlabel pdiffusion 507 -2213 507 -2213 0 cellNo=959
rlabel pdiffusion 514 -2213 514 -2213 0 feedthrough
rlabel pdiffusion 521 -2213 521 -2213 0 cellNo=960
rlabel pdiffusion 528 -2213 528 -2213 0 feedthrough
rlabel pdiffusion 535 -2213 535 -2213 0 feedthrough
rlabel pdiffusion 542 -2213 542 -2213 0 feedthrough
rlabel pdiffusion 549 -2213 549 -2213 0 feedthrough
rlabel pdiffusion 556 -2213 556 -2213 0 feedthrough
rlabel pdiffusion 563 -2213 563 -2213 0 cellNo=660
rlabel pdiffusion 570 -2213 570 -2213 0 cellNo=748
rlabel pdiffusion 577 -2213 577 -2213 0 feedthrough
rlabel pdiffusion 584 -2213 584 -2213 0 feedthrough
rlabel pdiffusion 591 -2213 591 -2213 0 cellNo=221
rlabel pdiffusion 598 -2213 598 -2213 0 cellNo=64
rlabel pdiffusion 605 -2213 605 -2213 0 cellNo=468
rlabel pdiffusion 612 -2213 612 -2213 0 feedthrough
rlabel pdiffusion 619 -2213 619 -2213 0 feedthrough
rlabel pdiffusion 626 -2213 626 -2213 0 feedthrough
rlabel pdiffusion 633 -2213 633 -2213 0 feedthrough
rlabel pdiffusion 640 -2213 640 -2213 0 feedthrough
rlabel pdiffusion 647 -2213 647 -2213 0 feedthrough
rlabel pdiffusion 654 -2213 654 -2213 0 feedthrough
rlabel pdiffusion 661 -2213 661 -2213 0 feedthrough
rlabel pdiffusion 668 -2213 668 -2213 0 cellNo=536
rlabel pdiffusion 675 -2213 675 -2213 0 feedthrough
rlabel pdiffusion 682 -2213 682 -2213 0 cellNo=49
rlabel pdiffusion 689 -2213 689 -2213 0 cellNo=940
rlabel pdiffusion 696 -2213 696 -2213 0 cellNo=790
rlabel pdiffusion 703 -2213 703 -2213 0 feedthrough
rlabel pdiffusion 710 -2213 710 -2213 0 feedthrough
rlabel pdiffusion 717 -2213 717 -2213 0 feedthrough
rlabel pdiffusion 724 -2213 724 -2213 0 cellNo=122
rlabel pdiffusion 731 -2213 731 -2213 0 feedthrough
rlabel pdiffusion 738 -2213 738 -2213 0 feedthrough
rlabel pdiffusion 745 -2213 745 -2213 0 feedthrough
rlabel pdiffusion 752 -2213 752 -2213 0 feedthrough
rlabel pdiffusion 759 -2213 759 -2213 0 feedthrough
rlabel pdiffusion 766 -2213 766 -2213 0 feedthrough
rlabel pdiffusion 773 -2213 773 -2213 0 feedthrough
rlabel pdiffusion 780 -2213 780 -2213 0 feedthrough
rlabel pdiffusion 787 -2213 787 -2213 0 feedthrough
rlabel pdiffusion 794 -2213 794 -2213 0 feedthrough
rlabel pdiffusion 801 -2213 801 -2213 0 feedthrough
rlabel pdiffusion 808 -2213 808 -2213 0 feedthrough
rlabel pdiffusion 815 -2213 815 -2213 0 feedthrough
rlabel pdiffusion 822 -2213 822 -2213 0 feedthrough
rlabel pdiffusion 829 -2213 829 -2213 0 feedthrough
rlabel pdiffusion 836 -2213 836 -2213 0 feedthrough
rlabel pdiffusion 843 -2213 843 -2213 0 feedthrough
rlabel pdiffusion 850 -2213 850 -2213 0 feedthrough
rlabel pdiffusion 857 -2213 857 -2213 0 feedthrough
rlabel pdiffusion 864 -2213 864 -2213 0 feedthrough
rlabel pdiffusion 871 -2213 871 -2213 0 cellNo=235
rlabel pdiffusion 878 -2213 878 -2213 0 feedthrough
rlabel pdiffusion 885 -2213 885 -2213 0 feedthrough
rlabel pdiffusion 892 -2213 892 -2213 0 feedthrough
rlabel pdiffusion 899 -2213 899 -2213 0 feedthrough
rlabel pdiffusion 906 -2213 906 -2213 0 feedthrough
rlabel pdiffusion 913 -2213 913 -2213 0 feedthrough
rlabel pdiffusion 920 -2213 920 -2213 0 feedthrough
rlabel pdiffusion 927 -2213 927 -2213 0 feedthrough
rlabel pdiffusion 934 -2213 934 -2213 0 feedthrough
rlabel pdiffusion 941 -2213 941 -2213 0 feedthrough
rlabel pdiffusion 948 -2213 948 -2213 0 feedthrough
rlabel pdiffusion 955 -2213 955 -2213 0 feedthrough
rlabel pdiffusion 962 -2213 962 -2213 0 feedthrough
rlabel pdiffusion 969 -2213 969 -2213 0 feedthrough
rlabel pdiffusion 976 -2213 976 -2213 0 feedthrough
rlabel pdiffusion 983 -2213 983 -2213 0 feedthrough
rlabel pdiffusion 990 -2213 990 -2213 0 feedthrough
rlabel pdiffusion 997 -2213 997 -2213 0 feedthrough
rlabel pdiffusion 1004 -2213 1004 -2213 0 feedthrough
rlabel pdiffusion 1011 -2213 1011 -2213 0 feedthrough
rlabel pdiffusion 1018 -2213 1018 -2213 0 feedthrough
rlabel pdiffusion 1025 -2213 1025 -2213 0 feedthrough
rlabel pdiffusion 1032 -2213 1032 -2213 0 feedthrough
rlabel pdiffusion 1039 -2213 1039 -2213 0 feedthrough
rlabel pdiffusion 1046 -2213 1046 -2213 0 feedthrough
rlabel pdiffusion 1053 -2213 1053 -2213 0 cellNo=922
rlabel pdiffusion 3 -2282 3 -2282 0 feedthrough
rlabel pdiffusion 10 -2282 10 -2282 0 feedthrough
rlabel pdiffusion 17 -2282 17 -2282 0 feedthrough
rlabel pdiffusion 24 -2282 24 -2282 0 feedthrough
rlabel pdiffusion 31 -2282 31 -2282 0 feedthrough
rlabel pdiffusion 38 -2282 38 -2282 0 feedthrough
rlabel pdiffusion 45 -2282 45 -2282 0 feedthrough
rlabel pdiffusion 52 -2282 52 -2282 0 cellNo=476
rlabel pdiffusion 59 -2282 59 -2282 0 cellNo=279
rlabel pdiffusion 66 -2282 66 -2282 0 feedthrough
rlabel pdiffusion 73 -2282 73 -2282 0 feedthrough
rlabel pdiffusion 80 -2282 80 -2282 0 cellNo=414
rlabel pdiffusion 87 -2282 87 -2282 0 feedthrough
rlabel pdiffusion 94 -2282 94 -2282 0 feedthrough
rlabel pdiffusion 101 -2282 101 -2282 0 cellNo=810
rlabel pdiffusion 108 -2282 108 -2282 0 cellNo=638
rlabel pdiffusion 115 -2282 115 -2282 0 feedthrough
rlabel pdiffusion 122 -2282 122 -2282 0 feedthrough
rlabel pdiffusion 129 -2282 129 -2282 0 cellNo=102
rlabel pdiffusion 136 -2282 136 -2282 0 feedthrough
rlabel pdiffusion 143 -2282 143 -2282 0 feedthrough
rlabel pdiffusion 150 -2282 150 -2282 0 feedthrough
rlabel pdiffusion 157 -2282 157 -2282 0 feedthrough
rlabel pdiffusion 164 -2282 164 -2282 0 feedthrough
rlabel pdiffusion 171 -2282 171 -2282 0 feedthrough
rlabel pdiffusion 178 -2282 178 -2282 0 cellNo=504
rlabel pdiffusion 185 -2282 185 -2282 0 feedthrough
rlabel pdiffusion 192 -2282 192 -2282 0 feedthrough
rlabel pdiffusion 199 -2282 199 -2282 0 cellNo=470
rlabel pdiffusion 206 -2282 206 -2282 0 feedthrough
rlabel pdiffusion 213 -2282 213 -2282 0 cellNo=671
rlabel pdiffusion 220 -2282 220 -2282 0 cellNo=256
rlabel pdiffusion 227 -2282 227 -2282 0 feedthrough
rlabel pdiffusion 234 -2282 234 -2282 0 feedthrough
rlabel pdiffusion 241 -2282 241 -2282 0 feedthrough
rlabel pdiffusion 248 -2282 248 -2282 0 feedthrough
rlabel pdiffusion 255 -2282 255 -2282 0 feedthrough
rlabel pdiffusion 262 -2282 262 -2282 0 feedthrough
rlabel pdiffusion 269 -2282 269 -2282 0 feedthrough
rlabel pdiffusion 276 -2282 276 -2282 0 feedthrough
rlabel pdiffusion 283 -2282 283 -2282 0 feedthrough
rlabel pdiffusion 290 -2282 290 -2282 0 cellNo=74
rlabel pdiffusion 297 -2282 297 -2282 0 feedthrough
rlabel pdiffusion 304 -2282 304 -2282 0 feedthrough
rlabel pdiffusion 311 -2282 311 -2282 0 feedthrough
rlabel pdiffusion 318 -2282 318 -2282 0 feedthrough
rlabel pdiffusion 325 -2282 325 -2282 0 cellNo=693
rlabel pdiffusion 332 -2282 332 -2282 0 feedthrough
rlabel pdiffusion 339 -2282 339 -2282 0 feedthrough
rlabel pdiffusion 346 -2282 346 -2282 0 cellNo=519
rlabel pdiffusion 353 -2282 353 -2282 0 cellNo=990
rlabel pdiffusion 360 -2282 360 -2282 0 feedthrough
rlabel pdiffusion 367 -2282 367 -2282 0 cellNo=706
rlabel pdiffusion 374 -2282 374 -2282 0 feedthrough
rlabel pdiffusion 381 -2282 381 -2282 0 cellNo=177
rlabel pdiffusion 388 -2282 388 -2282 0 feedthrough
rlabel pdiffusion 395 -2282 395 -2282 0 feedthrough
rlabel pdiffusion 402 -2282 402 -2282 0 feedthrough
rlabel pdiffusion 409 -2282 409 -2282 0 feedthrough
rlabel pdiffusion 416 -2282 416 -2282 0 feedthrough
rlabel pdiffusion 423 -2282 423 -2282 0 feedthrough
rlabel pdiffusion 430 -2282 430 -2282 0 feedthrough
rlabel pdiffusion 437 -2282 437 -2282 0 feedthrough
rlabel pdiffusion 444 -2282 444 -2282 0 feedthrough
rlabel pdiffusion 451 -2282 451 -2282 0 feedthrough
rlabel pdiffusion 458 -2282 458 -2282 0 feedthrough
rlabel pdiffusion 465 -2282 465 -2282 0 cellNo=123
rlabel pdiffusion 472 -2282 472 -2282 0 feedthrough
rlabel pdiffusion 479 -2282 479 -2282 0 cellNo=285
rlabel pdiffusion 486 -2282 486 -2282 0 cellNo=352
rlabel pdiffusion 493 -2282 493 -2282 0 feedthrough
rlabel pdiffusion 500 -2282 500 -2282 0 cellNo=632
rlabel pdiffusion 507 -2282 507 -2282 0 feedthrough
rlabel pdiffusion 514 -2282 514 -2282 0 feedthrough
rlabel pdiffusion 521 -2282 521 -2282 0 feedthrough
rlabel pdiffusion 528 -2282 528 -2282 0 feedthrough
rlabel pdiffusion 535 -2282 535 -2282 0 feedthrough
rlabel pdiffusion 542 -2282 542 -2282 0 cellNo=658
rlabel pdiffusion 549 -2282 549 -2282 0 feedthrough
rlabel pdiffusion 556 -2282 556 -2282 0 feedthrough
rlabel pdiffusion 563 -2282 563 -2282 0 feedthrough
rlabel pdiffusion 570 -2282 570 -2282 0 feedthrough
rlabel pdiffusion 577 -2282 577 -2282 0 cellNo=705
rlabel pdiffusion 584 -2282 584 -2282 0 cellNo=676
rlabel pdiffusion 591 -2282 591 -2282 0 feedthrough
rlabel pdiffusion 598 -2282 598 -2282 0 feedthrough
rlabel pdiffusion 605 -2282 605 -2282 0 feedthrough
rlabel pdiffusion 612 -2282 612 -2282 0 feedthrough
rlabel pdiffusion 619 -2282 619 -2282 0 feedthrough
rlabel pdiffusion 626 -2282 626 -2282 0 feedthrough
rlabel pdiffusion 633 -2282 633 -2282 0 feedthrough
rlabel pdiffusion 640 -2282 640 -2282 0 feedthrough
rlabel pdiffusion 647 -2282 647 -2282 0 feedthrough
rlabel pdiffusion 654 -2282 654 -2282 0 feedthrough
rlabel pdiffusion 661 -2282 661 -2282 0 feedthrough
rlabel pdiffusion 668 -2282 668 -2282 0 feedthrough
rlabel pdiffusion 675 -2282 675 -2282 0 feedthrough
rlabel pdiffusion 682 -2282 682 -2282 0 cellNo=303
rlabel pdiffusion 689 -2282 689 -2282 0 feedthrough
rlabel pdiffusion 696 -2282 696 -2282 0 feedthrough
rlabel pdiffusion 703 -2282 703 -2282 0 feedthrough
rlabel pdiffusion 710 -2282 710 -2282 0 feedthrough
rlabel pdiffusion 717 -2282 717 -2282 0 cellNo=688
rlabel pdiffusion 724 -2282 724 -2282 0 feedthrough
rlabel pdiffusion 731 -2282 731 -2282 0 feedthrough
rlabel pdiffusion 738 -2282 738 -2282 0 feedthrough
rlabel pdiffusion 745 -2282 745 -2282 0 feedthrough
rlabel pdiffusion 752 -2282 752 -2282 0 feedthrough
rlabel pdiffusion 759 -2282 759 -2282 0 feedthrough
rlabel pdiffusion 766 -2282 766 -2282 0 cellNo=952
rlabel pdiffusion 773 -2282 773 -2282 0 feedthrough
rlabel pdiffusion 780 -2282 780 -2282 0 feedthrough
rlabel pdiffusion 787 -2282 787 -2282 0 feedthrough
rlabel pdiffusion 794 -2282 794 -2282 0 feedthrough
rlabel pdiffusion 801 -2282 801 -2282 0 feedthrough
rlabel pdiffusion 808 -2282 808 -2282 0 feedthrough
rlabel pdiffusion 815 -2282 815 -2282 0 feedthrough
rlabel pdiffusion 822 -2282 822 -2282 0 feedthrough
rlabel pdiffusion 829 -2282 829 -2282 0 feedthrough
rlabel pdiffusion 836 -2282 836 -2282 0 feedthrough
rlabel pdiffusion 843 -2282 843 -2282 0 feedthrough
rlabel pdiffusion 850 -2282 850 -2282 0 feedthrough
rlabel pdiffusion 857 -2282 857 -2282 0 feedthrough
rlabel pdiffusion 864 -2282 864 -2282 0 feedthrough
rlabel pdiffusion 871 -2282 871 -2282 0 feedthrough
rlabel pdiffusion 878 -2282 878 -2282 0 feedthrough
rlabel pdiffusion 885 -2282 885 -2282 0 feedthrough
rlabel pdiffusion 892 -2282 892 -2282 0 feedthrough
rlabel pdiffusion 899 -2282 899 -2282 0 cellNo=115
rlabel pdiffusion 906 -2282 906 -2282 0 cellNo=412
rlabel pdiffusion 913 -2282 913 -2282 0 cellNo=797
rlabel pdiffusion 920 -2282 920 -2282 0 cellNo=109
rlabel pdiffusion 927 -2282 927 -2282 0 cellNo=759
rlabel pdiffusion 934 -2282 934 -2282 0 feedthrough
rlabel pdiffusion 941 -2282 941 -2282 0 feedthrough
rlabel pdiffusion 948 -2282 948 -2282 0 feedthrough
rlabel pdiffusion 955 -2282 955 -2282 0 feedthrough
rlabel pdiffusion 962 -2282 962 -2282 0 feedthrough
rlabel pdiffusion 969 -2282 969 -2282 0 cellNo=642
rlabel pdiffusion 976 -2282 976 -2282 0 feedthrough
rlabel pdiffusion 3 -2369 3 -2369 0 feedthrough
rlabel pdiffusion 10 -2369 10 -2369 0 cellNo=701
rlabel pdiffusion 17 -2369 17 -2369 0 feedthrough
rlabel pdiffusion 24 -2369 24 -2369 0 feedthrough
rlabel pdiffusion 31 -2369 31 -2369 0 feedthrough
rlabel pdiffusion 38 -2369 38 -2369 0 feedthrough
rlabel pdiffusion 45 -2369 45 -2369 0 cellNo=903
rlabel pdiffusion 52 -2369 52 -2369 0 cellNo=931
rlabel pdiffusion 59 -2369 59 -2369 0 feedthrough
rlabel pdiffusion 66 -2369 66 -2369 0 feedthrough
rlabel pdiffusion 73 -2369 73 -2369 0 feedthrough
rlabel pdiffusion 80 -2369 80 -2369 0 feedthrough
rlabel pdiffusion 87 -2369 87 -2369 0 feedthrough
rlabel pdiffusion 94 -2369 94 -2369 0 cellNo=293
rlabel pdiffusion 101 -2369 101 -2369 0 feedthrough
rlabel pdiffusion 108 -2369 108 -2369 0 cellNo=789
rlabel pdiffusion 115 -2369 115 -2369 0 feedthrough
rlabel pdiffusion 122 -2369 122 -2369 0 feedthrough
rlabel pdiffusion 129 -2369 129 -2369 0 feedthrough
rlabel pdiffusion 136 -2369 136 -2369 0 feedthrough
rlabel pdiffusion 143 -2369 143 -2369 0 feedthrough
rlabel pdiffusion 150 -2369 150 -2369 0 feedthrough
rlabel pdiffusion 157 -2369 157 -2369 0 cellNo=862
rlabel pdiffusion 164 -2369 164 -2369 0 feedthrough
rlabel pdiffusion 171 -2369 171 -2369 0 feedthrough
rlabel pdiffusion 178 -2369 178 -2369 0 feedthrough
rlabel pdiffusion 185 -2369 185 -2369 0 feedthrough
rlabel pdiffusion 192 -2369 192 -2369 0 feedthrough
rlabel pdiffusion 199 -2369 199 -2369 0 feedthrough
rlabel pdiffusion 206 -2369 206 -2369 0 feedthrough
rlabel pdiffusion 213 -2369 213 -2369 0 feedthrough
rlabel pdiffusion 220 -2369 220 -2369 0 cellNo=767
rlabel pdiffusion 227 -2369 227 -2369 0 cellNo=312
rlabel pdiffusion 234 -2369 234 -2369 0 feedthrough
rlabel pdiffusion 241 -2369 241 -2369 0 feedthrough
rlabel pdiffusion 248 -2369 248 -2369 0 feedthrough
rlabel pdiffusion 255 -2369 255 -2369 0 feedthrough
rlabel pdiffusion 262 -2369 262 -2369 0 feedthrough
rlabel pdiffusion 269 -2369 269 -2369 0 cellNo=126
rlabel pdiffusion 276 -2369 276 -2369 0 feedthrough
rlabel pdiffusion 283 -2369 283 -2369 0 feedthrough
rlabel pdiffusion 290 -2369 290 -2369 0 feedthrough
rlabel pdiffusion 297 -2369 297 -2369 0 feedthrough
rlabel pdiffusion 304 -2369 304 -2369 0 feedthrough
rlabel pdiffusion 311 -2369 311 -2369 0 cellNo=244
rlabel pdiffusion 318 -2369 318 -2369 0 feedthrough
rlabel pdiffusion 325 -2369 325 -2369 0 feedthrough
rlabel pdiffusion 332 -2369 332 -2369 0 cellNo=889
rlabel pdiffusion 339 -2369 339 -2369 0 cellNo=99
rlabel pdiffusion 346 -2369 346 -2369 0 feedthrough
rlabel pdiffusion 353 -2369 353 -2369 0 cellNo=422
rlabel pdiffusion 360 -2369 360 -2369 0 cellNo=932
rlabel pdiffusion 367 -2369 367 -2369 0 feedthrough
rlabel pdiffusion 374 -2369 374 -2369 0 cellNo=391
rlabel pdiffusion 381 -2369 381 -2369 0 feedthrough
rlabel pdiffusion 388 -2369 388 -2369 0 feedthrough
rlabel pdiffusion 395 -2369 395 -2369 0 cellNo=364
rlabel pdiffusion 402 -2369 402 -2369 0 cellNo=96
rlabel pdiffusion 409 -2369 409 -2369 0 feedthrough
rlabel pdiffusion 416 -2369 416 -2369 0 cellNo=220
rlabel pdiffusion 423 -2369 423 -2369 0 feedthrough
rlabel pdiffusion 430 -2369 430 -2369 0 feedthrough
rlabel pdiffusion 437 -2369 437 -2369 0 feedthrough
rlabel pdiffusion 444 -2369 444 -2369 0 feedthrough
rlabel pdiffusion 451 -2369 451 -2369 0 feedthrough
rlabel pdiffusion 458 -2369 458 -2369 0 cellNo=574
rlabel pdiffusion 465 -2369 465 -2369 0 cellNo=697
rlabel pdiffusion 472 -2369 472 -2369 0 feedthrough
rlabel pdiffusion 479 -2369 479 -2369 0 cellNo=753
rlabel pdiffusion 486 -2369 486 -2369 0 feedthrough
rlabel pdiffusion 493 -2369 493 -2369 0 feedthrough
rlabel pdiffusion 500 -2369 500 -2369 0 feedthrough
rlabel pdiffusion 507 -2369 507 -2369 0 feedthrough
rlabel pdiffusion 514 -2369 514 -2369 0 feedthrough
rlabel pdiffusion 521 -2369 521 -2369 0 cellNo=986
rlabel pdiffusion 528 -2369 528 -2369 0 feedthrough
rlabel pdiffusion 535 -2369 535 -2369 0 cellNo=718
rlabel pdiffusion 542 -2369 542 -2369 0 feedthrough
rlabel pdiffusion 549 -2369 549 -2369 0 feedthrough
rlabel pdiffusion 556 -2369 556 -2369 0 cellNo=93
rlabel pdiffusion 563 -2369 563 -2369 0 cellNo=55
rlabel pdiffusion 570 -2369 570 -2369 0 feedthrough
rlabel pdiffusion 577 -2369 577 -2369 0 feedthrough
rlabel pdiffusion 584 -2369 584 -2369 0 cellNo=762
rlabel pdiffusion 591 -2369 591 -2369 0 feedthrough
rlabel pdiffusion 598 -2369 598 -2369 0 feedthrough
rlabel pdiffusion 605 -2369 605 -2369 0 feedthrough
rlabel pdiffusion 612 -2369 612 -2369 0 feedthrough
rlabel pdiffusion 619 -2369 619 -2369 0 feedthrough
rlabel pdiffusion 626 -2369 626 -2369 0 feedthrough
rlabel pdiffusion 633 -2369 633 -2369 0 feedthrough
rlabel pdiffusion 640 -2369 640 -2369 0 cellNo=916
rlabel pdiffusion 647 -2369 647 -2369 0 feedthrough
rlabel pdiffusion 654 -2369 654 -2369 0 feedthrough
rlabel pdiffusion 661 -2369 661 -2369 0 feedthrough
rlabel pdiffusion 668 -2369 668 -2369 0 feedthrough
rlabel pdiffusion 675 -2369 675 -2369 0 feedthrough
rlabel pdiffusion 682 -2369 682 -2369 0 feedthrough
rlabel pdiffusion 689 -2369 689 -2369 0 feedthrough
rlabel pdiffusion 696 -2369 696 -2369 0 feedthrough
rlabel pdiffusion 703 -2369 703 -2369 0 cellNo=558
rlabel pdiffusion 710 -2369 710 -2369 0 feedthrough
rlabel pdiffusion 717 -2369 717 -2369 0 feedthrough
rlabel pdiffusion 724 -2369 724 -2369 0 feedthrough
rlabel pdiffusion 731 -2369 731 -2369 0 feedthrough
rlabel pdiffusion 738 -2369 738 -2369 0 feedthrough
rlabel pdiffusion 745 -2369 745 -2369 0 feedthrough
rlabel pdiffusion 752 -2369 752 -2369 0 feedthrough
rlabel pdiffusion 759 -2369 759 -2369 0 feedthrough
rlabel pdiffusion 766 -2369 766 -2369 0 feedthrough
rlabel pdiffusion 773 -2369 773 -2369 0 cellNo=769
rlabel pdiffusion 780 -2369 780 -2369 0 feedthrough
rlabel pdiffusion 787 -2369 787 -2369 0 feedthrough
rlabel pdiffusion 794 -2369 794 -2369 0 feedthrough
rlabel pdiffusion 801 -2369 801 -2369 0 cellNo=322
rlabel pdiffusion 808 -2369 808 -2369 0 feedthrough
rlabel pdiffusion 815 -2369 815 -2369 0 feedthrough
rlabel pdiffusion 822 -2369 822 -2369 0 feedthrough
rlabel pdiffusion 829 -2369 829 -2369 0 feedthrough
rlabel pdiffusion 836 -2369 836 -2369 0 feedthrough
rlabel pdiffusion 843 -2369 843 -2369 0 feedthrough
rlabel pdiffusion 850 -2369 850 -2369 0 feedthrough
rlabel pdiffusion 857 -2369 857 -2369 0 feedthrough
rlabel pdiffusion 864 -2369 864 -2369 0 feedthrough
rlabel pdiffusion 871 -2369 871 -2369 0 cellNo=953
rlabel pdiffusion 878 -2369 878 -2369 0 feedthrough
rlabel pdiffusion 885 -2369 885 -2369 0 feedthrough
rlabel pdiffusion 892 -2369 892 -2369 0 feedthrough
rlabel pdiffusion 927 -2369 927 -2369 0 cellNo=383
rlabel pdiffusion 948 -2369 948 -2369 0 feedthrough
rlabel pdiffusion 31 -2434 31 -2434 0 cellNo=242
rlabel pdiffusion 59 -2434 59 -2434 0 cellNo=611
rlabel pdiffusion 66 -2434 66 -2434 0 feedthrough
rlabel pdiffusion 73 -2434 73 -2434 0 cellNo=195
rlabel pdiffusion 80 -2434 80 -2434 0 feedthrough
rlabel pdiffusion 87 -2434 87 -2434 0 feedthrough
rlabel pdiffusion 94 -2434 94 -2434 0 feedthrough
rlabel pdiffusion 101 -2434 101 -2434 0 feedthrough
rlabel pdiffusion 108 -2434 108 -2434 0 feedthrough
rlabel pdiffusion 115 -2434 115 -2434 0 feedthrough
rlabel pdiffusion 122 -2434 122 -2434 0 feedthrough
rlabel pdiffusion 129 -2434 129 -2434 0 feedthrough
rlabel pdiffusion 136 -2434 136 -2434 0 cellNo=480
rlabel pdiffusion 143 -2434 143 -2434 0 feedthrough
rlabel pdiffusion 150 -2434 150 -2434 0 cellNo=63
rlabel pdiffusion 157 -2434 157 -2434 0 cellNo=458
rlabel pdiffusion 164 -2434 164 -2434 0 feedthrough
rlabel pdiffusion 171 -2434 171 -2434 0 feedthrough
rlabel pdiffusion 178 -2434 178 -2434 0 feedthrough
rlabel pdiffusion 185 -2434 185 -2434 0 cellNo=331
rlabel pdiffusion 192 -2434 192 -2434 0 feedthrough
rlabel pdiffusion 199 -2434 199 -2434 0 feedthrough
rlabel pdiffusion 206 -2434 206 -2434 0 cellNo=704
rlabel pdiffusion 213 -2434 213 -2434 0 cellNo=827
rlabel pdiffusion 220 -2434 220 -2434 0 cellNo=22
rlabel pdiffusion 227 -2434 227 -2434 0 feedthrough
rlabel pdiffusion 234 -2434 234 -2434 0 feedthrough
rlabel pdiffusion 241 -2434 241 -2434 0 feedthrough
rlabel pdiffusion 248 -2434 248 -2434 0 feedthrough
rlabel pdiffusion 255 -2434 255 -2434 0 feedthrough
rlabel pdiffusion 262 -2434 262 -2434 0 feedthrough
rlabel pdiffusion 269 -2434 269 -2434 0 feedthrough
rlabel pdiffusion 276 -2434 276 -2434 0 feedthrough
rlabel pdiffusion 283 -2434 283 -2434 0 feedthrough
rlabel pdiffusion 290 -2434 290 -2434 0 feedthrough
rlabel pdiffusion 297 -2434 297 -2434 0 cellNo=719
rlabel pdiffusion 304 -2434 304 -2434 0 feedthrough
rlabel pdiffusion 311 -2434 311 -2434 0 feedthrough
rlabel pdiffusion 318 -2434 318 -2434 0 feedthrough
rlabel pdiffusion 325 -2434 325 -2434 0 feedthrough
rlabel pdiffusion 332 -2434 332 -2434 0 cellNo=296
rlabel pdiffusion 339 -2434 339 -2434 0 feedthrough
rlabel pdiffusion 346 -2434 346 -2434 0 feedthrough
rlabel pdiffusion 353 -2434 353 -2434 0 feedthrough
rlabel pdiffusion 360 -2434 360 -2434 0 feedthrough
rlabel pdiffusion 367 -2434 367 -2434 0 feedthrough
rlabel pdiffusion 374 -2434 374 -2434 0 cellNo=974
rlabel pdiffusion 381 -2434 381 -2434 0 feedthrough
rlabel pdiffusion 388 -2434 388 -2434 0 feedthrough
rlabel pdiffusion 395 -2434 395 -2434 0 cellNo=822
rlabel pdiffusion 402 -2434 402 -2434 0 feedthrough
rlabel pdiffusion 409 -2434 409 -2434 0 cellNo=820
rlabel pdiffusion 416 -2434 416 -2434 0 feedthrough
rlabel pdiffusion 423 -2434 423 -2434 0 feedthrough
rlabel pdiffusion 430 -2434 430 -2434 0 cellNo=38
rlabel pdiffusion 437 -2434 437 -2434 0 feedthrough
rlabel pdiffusion 444 -2434 444 -2434 0 feedthrough
rlabel pdiffusion 451 -2434 451 -2434 0 feedthrough
rlabel pdiffusion 458 -2434 458 -2434 0 cellNo=246
rlabel pdiffusion 465 -2434 465 -2434 0 cellNo=914
rlabel pdiffusion 472 -2434 472 -2434 0 cellNo=875
rlabel pdiffusion 479 -2434 479 -2434 0 cellNo=6
rlabel pdiffusion 486 -2434 486 -2434 0 cellNo=23
rlabel pdiffusion 493 -2434 493 -2434 0 feedthrough
rlabel pdiffusion 500 -2434 500 -2434 0 feedthrough
rlabel pdiffusion 507 -2434 507 -2434 0 feedthrough
rlabel pdiffusion 514 -2434 514 -2434 0 feedthrough
rlabel pdiffusion 521 -2434 521 -2434 0 feedthrough
rlabel pdiffusion 528 -2434 528 -2434 0 feedthrough
rlabel pdiffusion 535 -2434 535 -2434 0 feedthrough
rlabel pdiffusion 542 -2434 542 -2434 0 cellNo=483
rlabel pdiffusion 549 -2434 549 -2434 0 cellNo=288
rlabel pdiffusion 556 -2434 556 -2434 0 feedthrough
rlabel pdiffusion 563 -2434 563 -2434 0 feedthrough
rlabel pdiffusion 570 -2434 570 -2434 0 feedthrough
rlabel pdiffusion 577 -2434 577 -2434 0 cellNo=808
rlabel pdiffusion 584 -2434 584 -2434 0 feedthrough
rlabel pdiffusion 591 -2434 591 -2434 0 feedthrough
rlabel pdiffusion 598 -2434 598 -2434 0 feedthrough
rlabel pdiffusion 605 -2434 605 -2434 0 feedthrough
rlabel pdiffusion 612 -2434 612 -2434 0 feedthrough
rlabel pdiffusion 619 -2434 619 -2434 0 feedthrough
rlabel pdiffusion 626 -2434 626 -2434 0 cellNo=647
rlabel pdiffusion 633 -2434 633 -2434 0 feedthrough
rlabel pdiffusion 640 -2434 640 -2434 0 feedthrough
rlabel pdiffusion 647 -2434 647 -2434 0 feedthrough
rlabel pdiffusion 654 -2434 654 -2434 0 feedthrough
rlabel pdiffusion 661 -2434 661 -2434 0 feedthrough
rlabel pdiffusion 668 -2434 668 -2434 0 feedthrough
rlabel pdiffusion 675 -2434 675 -2434 0 feedthrough
rlabel pdiffusion 682 -2434 682 -2434 0 feedthrough
rlabel pdiffusion 703 -2434 703 -2434 0 feedthrough
rlabel pdiffusion 710 -2434 710 -2434 0 feedthrough
rlabel pdiffusion 717 -2434 717 -2434 0 feedthrough
rlabel pdiffusion 724 -2434 724 -2434 0 cellNo=271
rlabel pdiffusion 731 -2434 731 -2434 0 cellNo=692
rlabel pdiffusion 738 -2434 738 -2434 0 feedthrough
rlabel pdiffusion 745 -2434 745 -2434 0 feedthrough
rlabel pdiffusion 752 -2434 752 -2434 0 cellNo=583
rlabel pdiffusion 759 -2434 759 -2434 0 cellNo=610
rlabel pdiffusion 766 -2434 766 -2434 0 feedthrough
rlabel pdiffusion 773 -2434 773 -2434 0 feedthrough
rlabel pdiffusion 780 -2434 780 -2434 0 cellNo=453
rlabel pdiffusion 808 -2434 808 -2434 0 feedthrough
rlabel pdiffusion 829 -2434 829 -2434 0 feedthrough
rlabel pdiffusion 885 -2434 885 -2434 0 feedthrough
rlabel pdiffusion 892 -2434 892 -2434 0 feedthrough
rlabel pdiffusion 927 -2434 927 -2434 0 feedthrough
rlabel pdiffusion 941 -2434 941 -2434 0 feedthrough
rlabel pdiffusion 3 -2475 3 -2475 0 cellNo=996
rlabel pdiffusion 66 -2475 66 -2475 0 cellNo=24
rlabel pdiffusion 73 -2475 73 -2475 0 feedthrough
rlabel pdiffusion 101 -2475 101 -2475 0 feedthrough
rlabel pdiffusion 108 -2475 108 -2475 0 feedthrough
rlabel pdiffusion 115 -2475 115 -2475 0 cellNo=254
rlabel pdiffusion 122 -2475 122 -2475 0 feedthrough
rlabel pdiffusion 129 -2475 129 -2475 0 cellNo=901
rlabel pdiffusion 136 -2475 136 -2475 0 feedthrough
rlabel pdiffusion 164 -2475 164 -2475 0 feedthrough
rlabel pdiffusion 171 -2475 171 -2475 0 feedthrough
rlabel pdiffusion 178 -2475 178 -2475 0 feedthrough
rlabel pdiffusion 185 -2475 185 -2475 0 cellNo=908
rlabel pdiffusion 192 -2475 192 -2475 0 feedthrough
rlabel pdiffusion 199 -2475 199 -2475 0 feedthrough
rlabel pdiffusion 206 -2475 206 -2475 0 feedthrough
rlabel pdiffusion 220 -2475 220 -2475 0 feedthrough
rlabel pdiffusion 227 -2475 227 -2475 0 feedthrough
rlabel pdiffusion 234 -2475 234 -2475 0 cellNo=601
rlabel pdiffusion 241 -2475 241 -2475 0 cellNo=261
rlabel pdiffusion 248 -2475 248 -2475 0 feedthrough
rlabel pdiffusion 255 -2475 255 -2475 0 cellNo=141
rlabel pdiffusion 262 -2475 262 -2475 0 cellNo=801
rlabel pdiffusion 269 -2475 269 -2475 0 feedthrough
rlabel pdiffusion 276 -2475 276 -2475 0 feedthrough
rlabel pdiffusion 283 -2475 283 -2475 0 feedthrough
rlabel pdiffusion 290 -2475 290 -2475 0 feedthrough
rlabel pdiffusion 297 -2475 297 -2475 0 cellNo=13
rlabel pdiffusion 304 -2475 304 -2475 0 feedthrough
rlabel pdiffusion 311 -2475 311 -2475 0 feedthrough
rlabel pdiffusion 318 -2475 318 -2475 0 feedthrough
rlabel pdiffusion 325 -2475 325 -2475 0 cellNo=270
rlabel pdiffusion 332 -2475 332 -2475 0 feedthrough
rlabel pdiffusion 339 -2475 339 -2475 0 feedthrough
rlabel pdiffusion 346 -2475 346 -2475 0 cellNo=500
rlabel pdiffusion 353 -2475 353 -2475 0 feedthrough
rlabel pdiffusion 360 -2475 360 -2475 0 feedthrough
rlabel pdiffusion 367 -2475 367 -2475 0 cellNo=934
rlabel pdiffusion 374 -2475 374 -2475 0 cellNo=828
rlabel pdiffusion 381 -2475 381 -2475 0 feedthrough
rlabel pdiffusion 388 -2475 388 -2475 0 cellNo=29
rlabel pdiffusion 395 -2475 395 -2475 0 feedthrough
rlabel pdiffusion 402 -2475 402 -2475 0 feedthrough
rlabel pdiffusion 409 -2475 409 -2475 0 feedthrough
rlabel pdiffusion 416 -2475 416 -2475 0 feedthrough
rlabel pdiffusion 423 -2475 423 -2475 0 feedthrough
rlabel pdiffusion 430 -2475 430 -2475 0 cellNo=689
rlabel pdiffusion 437 -2475 437 -2475 0 feedthrough
rlabel pdiffusion 444 -2475 444 -2475 0 feedthrough
rlabel pdiffusion 451 -2475 451 -2475 0 cellNo=835
rlabel pdiffusion 458 -2475 458 -2475 0 feedthrough
rlabel pdiffusion 465 -2475 465 -2475 0 cellNo=75
rlabel pdiffusion 472 -2475 472 -2475 0 feedthrough
rlabel pdiffusion 479 -2475 479 -2475 0 feedthrough
rlabel pdiffusion 500 -2475 500 -2475 0 cellNo=667
rlabel pdiffusion 507 -2475 507 -2475 0 feedthrough
rlabel pdiffusion 514 -2475 514 -2475 0 feedthrough
rlabel pdiffusion 521 -2475 521 -2475 0 cellNo=926
rlabel pdiffusion 528 -2475 528 -2475 0 cellNo=330
rlabel pdiffusion 535 -2475 535 -2475 0 cellNo=838
rlabel pdiffusion 542 -2475 542 -2475 0 feedthrough
rlabel pdiffusion 549 -2475 549 -2475 0 feedthrough
rlabel pdiffusion 570 -2475 570 -2475 0 feedthrough
rlabel pdiffusion 577 -2475 577 -2475 0 feedthrough
rlabel pdiffusion 584 -2475 584 -2475 0 cellNo=457
rlabel pdiffusion 591 -2475 591 -2475 0 cellNo=879
rlabel pdiffusion 598 -2475 598 -2475 0 cellNo=562
rlabel pdiffusion 605 -2475 605 -2475 0 feedthrough
rlabel pdiffusion 612 -2475 612 -2475 0 feedthrough
rlabel pdiffusion 626 -2475 626 -2475 0 feedthrough
rlabel pdiffusion 640 -2475 640 -2475 0 cellNo=728
rlabel pdiffusion 661 -2475 661 -2475 0 feedthrough
rlabel pdiffusion 675 -2475 675 -2475 0 feedthrough
rlabel pdiffusion 682 -2475 682 -2475 0 feedthrough
rlabel pdiffusion 689 -2475 689 -2475 0 feedthrough
rlabel pdiffusion 696 -2475 696 -2475 0 cellNo=45
rlabel pdiffusion 710 -2475 710 -2475 0 feedthrough
rlabel pdiffusion 717 -2475 717 -2475 0 feedthrough
rlabel pdiffusion 724 -2475 724 -2475 0 feedthrough
rlabel pdiffusion 731 -2475 731 -2475 0 feedthrough
rlabel pdiffusion 738 -2475 738 -2475 0 feedthrough
rlabel pdiffusion 759 -2475 759 -2475 0 cellNo=796
rlabel pdiffusion 766 -2475 766 -2475 0 feedthrough
rlabel pdiffusion 885 -2475 885 -2475 0 feedthrough
rlabel pdiffusion 892 -2475 892 -2475 0 feedthrough
rlabel pdiffusion 934 -2475 934 -2475 0 cellNo=455
rlabel pdiffusion 941 -2475 941 -2475 0 feedthrough
rlabel pdiffusion 3 -2502 3 -2502 0 cellNo=955
rlabel pdiffusion 87 -2502 87 -2502 0 feedthrough
rlabel pdiffusion 94 -2502 94 -2502 0 cellNo=674
rlabel pdiffusion 101 -2502 101 -2502 0 cellNo=9
rlabel pdiffusion 108 -2502 108 -2502 0 cellNo=794
rlabel pdiffusion 115 -2502 115 -2502 0 cellNo=67
rlabel pdiffusion 122 -2502 122 -2502 0 feedthrough
rlabel pdiffusion 136 -2502 136 -2502 0 cellNo=856
rlabel pdiffusion 143 -2502 143 -2502 0 feedthrough
rlabel pdiffusion 150 -2502 150 -2502 0 feedthrough
rlabel pdiffusion 157 -2502 157 -2502 0 cellNo=353
rlabel pdiffusion 164 -2502 164 -2502 0 cellNo=843
rlabel pdiffusion 171 -2502 171 -2502 0 feedthrough
rlabel pdiffusion 178 -2502 178 -2502 0 feedthrough
rlabel pdiffusion 185 -2502 185 -2502 0 cellNo=659
rlabel pdiffusion 192 -2502 192 -2502 0 cellNo=588
rlabel pdiffusion 199 -2502 199 -2502 0 cellNo=281
rlabel pdiffusion 206 -2502 206 -2502 0 feedthrough
rlabel pdiffusion 213 -2502 213 -2502 0 feedthrough
rlabel pdiffusion 220 -2502 220 -2502 0 cellNo=7
rlabel pdiffusion 227 -2502 227 -2502 0 feedthrough
rlabel pdiffusion 234 -2502 234 -2502 0 feedthrough
rlabel pdiffusion 241 -2502 241 -2502 0 feedthrough
rlabel pdiffusion 248 -2502 248 -2502 0 feedthrough
rlabel pdiffusion 255 -2502 255 -2502 0 feedthrough
rlabel pdiffusion 262 -2502 262 -2502 0 feedthrough
rlabel pdiffusion 269 -2502 269 -2502 0 cellNo=70
rlabel pdiffusion 276 -2502 276 -2502 0 feedthrough
rlabel pdiffusion 283 -2502 283 -2502 0 cellNo=913
rlabel pdiffusion 290 -2502 290 -2502 0 feedthrough
rlabel pdiffusion 297 -2502 297 -2502 0 cellNo=255
rlabel pdiffusion 304 -2502 304 -2502 0 cellNo=821
rlabel pdiffusion 311 -2502 311 -2502 0 feedthrough
rlabel pdiffusion 318 -2502 318 -2502 0 feedthrough
rlabel pdiffusion 325 -2502 325 -2502 0 feedthrough
rlabel pdiffusion 332 -2502 332 -2502 0 feedthrough
rlabel pdiffusion 353 -2502 353 -2502 0 feedthrough
rlabel pdiffusion 360 -2502 360 -2502 0 cellNo=892
rlabel pdiffusion 381 -2502 381 -2502 0 feedthrough
rlabel pdiffusion 388 -2502 388 -2502 0 cellNo=367
rlabel pdiffusion 395 -2502 395 -2502 0 feedthrough
rlabel pdiffusion 402 -2502 402 -2502 0 cellNo=491
rlabel pdiffusion 409 -2502 409 -2502 0 feedthrough
rlabel pdiffusion 416 -2502 416 -2502 0 cellNo=247
rlabel pdiffusion 423 -2502 423 -2502 0 cellNo=992
rlabel pdiffusion 444 -2502 444 -2502 0 feedthrough
rlabel pdiffusion 451 -2502 451 -2502 0 feedthrough
rlabel pdiffusion 521 -2502 521 -2502 0 cellNo=736
rlabel pdiffusion 528 -2502 528 -2502 0 feedthrough
rlabel pdiffusion 605 -2502 605 -2502 0 feedthrough
rlabel pdiffusion 612 -2502 612 -2502 0 feedthrough
rlabel pdiffusion 661 -2502 661 -2502 0 feedthrough
rlabel pdiffusion 668 -2502 668 -2502 0 feedthrough
rlabel pdiffusion 682 -2502 682 -2502 0 feedthrough
rlabel pdiffusion 689 -2502 689 -2502 0 feedthrough
rlabel pdiffusion 696 -2502 696 -2502 0 feedthrough
rlabel pdiffusion 703 -2502 703 -2502 0 cellNo=15
rlabel pdiffusion 710 -2502 710 -2502 0 feedthrough
rlabel pdiffusion 717 -2502 717 -2502 0 feedthrough
rlabel pdiffusion 724 -2502 724 -2502 0 feedthrough
rlabel pdiffusion 731 -2502 731 -2502 0 cellNo=541
rlabel pdiffusion 738 -2502 738 -2502 0 cellNo=488
rlabel pdiffusion 745 -2502 745 -2502 0 cellNo=888
rlabel pdiffusion 752 -2502 752 -2502 0 feedthrough
rlabel pdiffusion 759 -2502 759 -2502 0 feedthrough
rlabel pdiffusion 885 -2502 885 -2502 0 cellNo=818
rlabel pdiffusion 892 -2502 892 -2502 0 feedthrough
rlabel pdiffusion 934 -2502 934 -2502 0 feedthrough
rlabel pdiffusion 941 -2502 941 -2502 0 cellNo=772
rlabel pdiffusion 948 -2502 948 -2502 0 feedthrough
rlabel pdiffusion 3 -2521 3 -2521 0 cellNo=846
rlabel pdiffusion 10 -2521 10 -2521 0 feedthrough
rlabel pdiffusion 101 -2521 101 -2521 0 cellNo=739
rlabel pdiffusion 108 -2521 108 -2521 0 feedthrough
rlabel pdiffusion 115 -2521 115 -2521 0 feedthrough
rlabel pdiffusion 122 -2521 122 -2521 0 cellNo=600
rlabel pdiffusion 129 -2521 129 -2521 0 cellNo=784
rlabel pdiffusion 157 -2521 157 -2521 0 cellNo=37
rlabel pdiffusion 164 -2521 164 -2521 0 feedthrough
rlabel pdiffusion 171 -2521 171 -2521 0 cellNo=669
rlabel pdiffusion 178 -2521 178 -2521 0 cellNo=809
rlabel pdiffusion 185 -2521 185 -2521 0 feedthrough
rlabel pdiffusion 192 -2521 192 -2521 0 feedthrough
rlabel pdiffusion 199 -2521 199 -2521 0 cellNo=855
rlabel pdiffusion 227 -2521 227 -2521 0 cellNo=950
rlabel pdiffusion 269 -2521 269 -2521 0 cellNo=61
rlabel pdiffusion 276 -2521 276 -2521 0 cellNo=471
rlabel pdiffusion 283 -2521 283 -2521 0 cellNo=842
rlabel pdiffusion 290 -2521 290 -2521 0 cellNo=780
rlabel pdiffusion 297 -2521 297 -2521 0 feedthrough
rlabel pdiffusion 304 -2521 304 -2521 0 cellNo=755
rlabel pdiffusion 311 -2521 311 -2521 0 feedthrough
rlabel pdiffusion 339 -2521 339 -2521 0 cellNo=881
rlabel pdiffusion 346 -2521 346 -2521 0 feedthrough
rlabel pdiffusion 360 -2521 360 -2521 0 cellNo=538
rlabel pdiffusion 381 -2521 381 -2521 0 cellNo=958
rlabel pdiffusion 395 -2521 395 -2521 0 cellNo=428
rlabel pdiffusion 402 -2521 402 -2521 0 cellNo=941
rlabel pdiffusion 451 -2521 451 -2521 0 feedthrough
rlabel pdiffusion 458 -2521 458 -2521 0 cellNo=863
rlabel pdiffusion 521 -2521 521 -2521 0 cellNo=361
rlabel pdiffusion 598 -2521 598 -2521 0 cellNo=983
rlabel pdiffusion 605 -2521 605 -2521 0 feedthrough
rlabel pdiffusion 661 -2521 661 -2521 0 cellNo=819
rlabel pdiffusion 668 -2521 668 -2521 0 feedthrough
rlabel pdiffusion 689 -2521 689 -2521 0 cellNo=764
rlabel pdiffusion 710 -2521 710 -2521 0 cellNo=192
rlabel pdiffusion 717 -2521 717 -2521 0 feedthrough
rlabel pdiffusion 724 -2521 724 -2521 0 cellNo=985
rlabel pdiffusion 731 -2521 731 -2521 0 feedthrough
rlabel pdiffusion 738 -2521 738 -2521 0 cellNo=869
rlabel polysilicon 86 -10 86 -10 0 3
rlabel polysilicon 89 -10 89 -10 0 4
rlabel polysilicon 93 -4 93 -4 0 1
rlabel polysilicon 93 -10 93 -10 0 3
rlabel polysilicon 100 -4 100 -4 0 1
rlabel polysilicon 100 -10 100 -10 0 3
rlabel polysilicon 107 -4 107 -4 0 1
rlabel polysilicon 107 -10 107 -10 0 3
rlabel polysilicon 117 -4 117 -4 0 2
rlabel polysilicon 121 -4 121 -4 0 1
rlabel polysilicon 121 -10 121 -10 0 3
rlabel polysilicon 128 -4 128 -4 0 1
rlabel polysilicon 128 -10 128 -10 0 3
rlabel polysilicon 145 -10 145 -10 0 4
rlabel polysilicon 205 -4 205 -4 0 1
rlabel polysilicon 205 -10 205 -10 0 3
rlabel polysilicon 212 -4 212 -4 0 1
rlabel polysilicon 215 -4 215 -4 0 2
rlabel polysilicon 219 -10 219 -10 0 3
rlabel polysilicon 222 -10 222 -10 0 4
rlabel polysilicon 226 -4 226 -4 0 1
rlabel polysilicon 226 -10 226 -10 0 3
rlabel polysilicon 233 -4 233 -4 0 1
rlabel polysilicon 236 -4 236 -4 0 2
rlabel polysilicon 240 -4 240 -4 0 1
rlabel polysilicon 240 -10 240 -10 0 3
rlabel polysilicon 247 -4 247 -4 0 1
rlabel polysilicon 250 -10 250 -10 0 4
rlabel polysilicon 257 -10 257 -10 0 4
rlabel polysilicon 261 -4 261 -4 0 1
rlabel polysilicon 268 -4 268 -4 0 1
rlabel polysilicon 268 -10 268 -10 0 3
rlabel polysilicon 282 -10 282 -10 0 3
rlabel polysilicon 324 -4 324 -4 0 1
rlabel polysilicon 324 -10 324 -10 0 3
rlabel polysilicon 334 -4 334 -4 0 2
rlabel polysilicon 341 -10 341 -10 0 4
rlabel polysilicon 429 -4 429 -4 0 1
rlabel polysilicon 429 -10 429 -10 0 3
rlabel polysilicon 450 -4 450 -4 0 1
rlabel polysilicon 450 -10 450 -10 0 3
rlabel polysilicon 464 -4 464 -4 0 1
rlabel polysilicon 464 -10 464 -10 0 3
rlabel polysilicon 488 -4 488 -4 0 2
rlabel polysilicon 485 -10 485 -10 0 3
rlabel polysilicon 509 -10 509 -10 0 4
rlabel polysilicon 530 -4 530 -4 0 2
rlabel polysilicon 534 -4 534 -4 0 1
rlabel polysilicon 534 -10 534 -10 0 3
rlabel polysilicon 548 -10 548 -10 0 3
rlabel polysilicon 583 -4 583 -4 0 1
rlabel polysilicon 590 -10 590 -10 0 3
rlabel polysilicon 597 -4 597 -4 0 1
rlabel polysilicon 597 -10 597 -10 0 3
rlabel polysilicon 607 -10 607 -10 0 4
rlabel polysilicon 660 -4 660 -4 0 1
rlabel polysilicon 667 -4 667 -4 0 1
rlabel polysilicon 667 -10 667 -10 0 3
rlabel polysilicon 100 -23 100 -23 0 1
rlabel polysilicon 103 -23 103 -23 0 2
rlabel polysilicon 100 -29 100 -29 0 3
rlabel polysilicon 103 -29 103 -29 0 4
rlabel polysilicon 117 -23 117 -23 0 2
rlabel polysilicon 135 -23 135 -23 0 1
rlabel polysilicon 135 -29 135 -29 0 3
rlabel polysilicon 173 -23 173 -23 0 2
rlabel polysilicon 177 -23 177 -23 0 1
rlabel polysilicon 177 -29 177 -29 0 3
rlabel polysilicon 184 -23 184 -23 0 1
rlabel polysilicon 184 -29 184 -29 0 3
rlabel polysilicon 194 -29 194 -29 0 4
rlabel polysilicon 198 -23 198 -23 0 1
rlabel polysilicon 198 -29 198 -29 0 3
rlabel polysilicon 205 -23 205 -23 0 1
rlabel polysilicon 212 -23 212 -23 0 1
rlabel polysilicon 215 -23 215 -23 0 2
rlabel polysilicon 212 -29 212 -29 0 3
rlabel polysilicon 219 -23 219 -23 0 1
rlabel polysilicon 219 -29 219 -29 0 3
rlabel polysilicon 226 -23 226 -23 0 1
rlabel polysilicon 226 -29 226 -29 0 3
rlabel polysilicon 233 -23 233 -23 0 1
rlabel polysilicon 236 -23 236 -23 0 2
rlabel polysilicon 240 -23 240 -23 0 1
rlabel polysilicon 247 -23 247 -23 0 1
rlabel polysilicon 247 -29 247 -29 0 3
rlabel polysilicon 254 -23 254 -23 0 1
rlabel polysilicon 254 -29 254 -29 0 3
rlabel polysilicon 261 -23 261 -23 0 1
rlabel polysilicon 261 -29 261 -29 0 3
rlabel polysilicon 268 -23 268 -23 0 1
rlabel polysilicon 268 -29 268 -29 0 3
rlabel polysilicon 275 -23 275 -23 0 1
rlabel polysilicon 275 -29 275 -29 0 3
rlabel polysilicon 282 -23 282 -23 0 1
rlabel polysilicon 282 -29 282 -29 0 3
rlabel polysilicon 289 -23 289 -23 0 1
rlabel polysilicon 289 -29 289 -29 0 3
rlabel polysilicon 296 -29 296 -29 0 3
rlabel polysilicon 303 -23 303 -23 0 1
rlabel polysilicon 306 -23 306 -23 0 2
rlabel polysilicon 310 -23 310 -23 0 1
rlabel polysilicon 310 -29 310 -29 0 3
rlabel polysilicon 317 -23 317 -23 0 1
rlabel polysilicon 317 -29 317 -29 0 3
rlabel polysilicon 324 -23 324 -23 0 1
rlabel polysilicon 324 -29 324 -29 0 3
rlabel polysilicon 331 -23 331 -23 0 1
rlabel polysilicon 338 -29 338 -29 0 3
rlabel polysilicon 348 -23 348 -23 0 2
rlabel polysilicon 348 -29 348 -29 0 4
rlabel polysilicon 359 -23 359 -23 0 1
rlabel polysilicon 359 -29 359 -29 0 3
rlabel polysilicon 373 -23 373 -23 0 1
rlabel polysilicon 373 -29 373 -29 0 3
rlabel polysilicon 383 -29 383 -29 0 4
rlabel polysilicon 415 -23 415 -23 0 1
rlabel polysilicon 415 -29 415 -29 0 3
rlabel polysilicon 422 -29 422 -29 0 3
rlabel polysilicon 429 -23 429 -23 0 1
rlabel polysilicon 429 -29 429 -29 0 3
rlabel polysilicon 439 -23 439 -23 0 2
rlabel polysilicon 446 -23 446 -23 0 2
rlabel polysilicon 446 -29 446 -29 0 4
rlabel polysilicon 453 -23 453 -23 0 2
rlabel polysilicon 464 -29 464 -29 0 3
rlabel polysilicon 467 -29 467 -29 0 4
rlabel polysilicon 471 -23 471 -23 0 1
rlabel polysilicon 471 -29 471 -29 0 3
rlabel polysilicon 492 -23 492 -23 0 1
rlabel polysilicon 492 -29 492 -29 0 3
rlabel polysilicon 506 -23 506 -23 0 1
rlabel polysilicon 506 -29 506 -29 0 3
rlabel polysilicon 513 -23 513 -23 0 1
rlabel polysilicon 513 -29 513 -29 0 3
rlabel polysilicon 520 -29 520 -29 0 3
rlabel polysilicon 527 -23 527 -23 0 1
rlabel polysilicon 527 -29 527 -29 0 3
rlabel polysilicon 541 -23 541 -23 0 1
rlabel polysilicon 541 -29 541 -29 0 3
rlabel polysilicon 555 -29 555 -29 0 3
rlabel polysilicon 562 -23 562 -23 0 1
rlabel polysilicon 569 -23 569 -23 0 1
rlabel polysilicon 569 -29 569 -29 0 3
rlabel polysilicon 576 -23 576 -23 0 1
rlabel polysilicon 576 -29 576 -29 0 3
rlabel polysilicon 604 -23 604 -23 0 1
rlabel polysilicon 604 -29 604 -29 0 3
rlabel polysilicon 611 -23 611 -23 0 1
rlabel polysilicon 611 -29 611 -29 0 3
rlabel polysilicon 618 -23 618 -23 0 1
rlabel polysilicon 618 -29 618 -29 0 3
rlabel polysilicon 674 -23 674 -23 0 1
rlabel polysilicon 674 -29 674 -29 0 3
rlabel polysilicon 86 -54 86 -54 0 1
rlabel polysilicon 86 -60 86 -60 0 3
rlabel polysilicon 93 -54 93 -54 0 1
rlabel polysilicon 93 -60 93 -60 0 3
rlabel polysilicon 114 -54 114 -54 0 1
rlabel polysilicon 114 -60 114 -60 0 3
rlabel polysilicon 121 -54 121 -54 0 1
rlabel polysilicon 121 -60 121 -60 0 3
rlabel polysilicon 128 -54 128 -54 0 1
rlabel polysilicon 128 -60 128 -60 0 3
rlabel polysilicon 135 -54 135 -54 0 1
rlabel polysilicon 135 -60 135 -60 0 3
rlabel polysilicon 145 -54 145 -54 0 2
rlabel polysilicon 149 -60 149 -60 0 3
rlabel polysilicon 156 -54 156 -54 0 1
rlabel polysilicon 156 -60 156 -60 0 3
rlabel polysilicon 163 -54 163 -54 0 1
rlabel polysilicon 163 -60 163 -60 0 3
rlabel polysilicon 173 -54 173 -54 0 2
rlabel polysilicon 170 -60 170 -60 0 3
rlabel polysilicon 173 -60 173 -60 0 4
rlabel polysilicon 177 -54 177 -54 0 1
rlabel polysilicon 177 -60 177 -60 0 3
rlabel polysilicon 187 -54 187 -54 0 2
rlabel polysilicon 184 -60 184 -60 0 3
rlabel polysilicon 191 -54 191 -54 0 1
rlabel polysilicon 191 -60 191 -60 0 3
rlabel polysilicon 198 -54 198 -54 0 1
rlabel polysilicon 201 -54 201 -54 0 2
rlabel polysilicon 205 -54 205 -54 0 1
rlabel polysilicon 205 -60 205 -60 0 3
rlabel polysilicon 212 -54 212 -54 0 1
rlabel polysilicon 212 -60 212 -60 0 3
rlabel polysilicon 219 -54 219 -54 0 1
rlabel polysilicon 219 -60 219 -60 0 3
rlabel polysilicon 226 -54 226 -54 0 1
rlabel polysilicon 226 -60 226 -60 0 3
rlabel polysilicon 236 -54 236 -54 0 2
rlabel polysilicon 233 -60 233 -60 0 3
rlabel polysilicon 240 -60 240 -60 0 3
rlabel polysilicon 243 -60 243 -60 0 4
rlabel polysilicon 247 -54 247 -54 0 1
rlabel polysilicon 250 -54 250 -54 0 2
rlabel polysilicon 250 -60 250 -60 0 4
rlabel polysilicon 254 -54 254 -54 0 1
rlabel polysilicon 254 -60 254 -60 0 3
rlabel polysilicon 261 -54 261 -54 0 1
rlabel polysilicon 261 -60 261 -60 0 3
rlabel polysilicon 268 -54 268 -54 0 1
rlabel polysilicon 268 -60 268 -60 0 3
rlabel polysilicon 275 -54 275 -54 0 1
rlabel polysilicon 275 -60 275 -60 0 3
rlabel polysilicon 282 -54 282 -54 0 1
rlabel polysilicon 282 -60 282 -60 0 3
rlabel polysilicon 289 -54 289 -54 0 1
rlabel polysilicon 289 -60 289 -60 0 3
rlabel polysilicon 299 -54 299 -54 0 2
rlabel polysilicon 296 -60 296 -60 0 3
rlabel polysilicon 303 -54 303 -54 0 1
rlabel polysilicon 303 -60 303 -60 0 3
rlabel polysilicon 313 -54 313 -54 0 2
rlabel polysilicon 310 -60 310 -60 0 3
rlabel polysilicon 317 -54 317 -54 0 1
rlabel polysilicon 317 -60 317 -60 0 3
rlabel polysilicon 324 -54 324 -54 0 1
rlabel polysilicon 324 -60 324 -60 0 3
rlabel polysilicon 331 -54 331 -54 0 1
rlabel polysilicon 331 -60 331 -60 0 3
rlabel polysilicon 338 -54 338 -54 0 1
rlabel polysilicon 341 -54 341 -54 0 2
rlabel polysilicon 341 -60 341 -60 0 4
rlabel polysilicon 345 -54 345 -54 0 1
rlabel polysilicon 345 -60 345 -60 0 3
rlabel polysilicon 352 -54 352 -54 0 1
rlabel polysilicon 352 -60 352 -60 0 3
rlabel polysilicon 359 -60 359 -60 0 3
rlabel polysilicon 366 -54 366 -54 0 1
rlabel polysilicon 366 -60 366 -60 0 3
rlabel polysilicon 373 -54 373 -54 0 1
rlabel polysilicon 373 -60 373 -60 0 3
rlabel polysilicon 383 -54 383 -54 0 2
rlabel polysilicon 380 -60 380 -60 0 3
rlabel polysilicon 387 -54 387 -54 0 1
rlabel polysilicon 387 -60 387 -60 0 3
rlabel polysilicon 394 -54 394 -54 0 1
rlabel polysilicon 394 -60 394 -60 0 3
rlabel polysilicon 401 -54 401 -54 0 1
rlabel polysilicon 401 -60 401 -60 0 3
rlabel polysilicon 408 -54 408 -54 0 1
rlabel polysilicon 408 -60 408 -60 0 3
rlabel polysilicon 418 -60 418 -60 0 4
rlabel polysilicon 422 -54 422 -54 0 1
rlabel polysilicon 422 -60 422 -60 0 3
rlabel polysilicon 429 -54 429 -54 0 1
rlabel polysilicon 429 -60 429 -60 0 3
rlabel polysilicon 436 -54 436 -54 0 1
rlabel polysilicon 436 -60 436 -60 0 3
rlabel polysilicon 443 -54 443 -54 0 1
rlabel polysilicon 443 -60 443 -60 0 3
rlabel polysilicon 464 -54 464 -54 0 1
rlabel polysilicon 467 -60 467 -60 0 4
rlabel polysilicon 471 -54 471 -54 0 1
rlabel polysilicon 471 -60 471 -60 0 3
rlabel polysilicon 478 -54 478 -54 0 1
rlabel polysilicon 478 -60 478 -60 0 3
rlabel polysilicon 485 -54 485 -54 0 1
rlabel polysilicon 485 -60 485 -60 0 3
rlabel polysilicon 492 -60 492 -60 0 3
rlabel polysilicon 495 -60 495 -60 0 4
rlabel polysilicon 499 -54 499 -54 0 1
rlabel polysilicon 499 -60 499 -60 0 3
rlabel polysilicon 506 -54 506 -54 0 1
rlabel polysilicon 506 -60 506 -60 0 3
rlabel polysilicon 520 -54 520 -54 0 1
rlabel polysilicon 520 -60 520 -60 0 3
rlabel polysilicon 527 -54 527 -54 0 1
rlabel polysilicon 530 -60 530 -60 0 4
rlabel polysilicon 534 -54 534 -54 0 1
rlabel polysilicon 534 -60 534 -60 0 3
rlabel polysilicon 541 -54 541 -54 0 1
rlabel polysilicon 541 -60 541 -60 0 3
rlabel polysilicon 551 -54 551 -54 0 2
rlabel polysilicon 548 -60 548 -60 0 3
rlabel polysilicon 555 -54 555 -54 0 1
rlabel polysilicon 555 -60 555 -60 0 3
rlabel polysilicon 562 -54 562 -54 0 1
rlabel polysilicon 562 -60 562 -60 0 3
rlabel polysilicon 569 -54 569 -54 0 1
rlabel polysilicon 569 -60 569 -60 0 3
rlabel polysilicon 576 -54 576 -54 0 1
rlabel polysilicon 576 -60 576 -60 0 3
rlabel polysilicon 586 -54 586 -54 0 2
rlabel polysilicon 583 -60 583 -60 0 3
rlabel polysilicon 586 -60 586 -60 0 4
rlabel polysilicon 590 -54 590 -54 0 1
rlabel polysilicon 590 -60 590 -60 0 3
rlabel polysilicon 597 -54 597 -54 0 1
rlabel polysilicon 597 -60 597 -60 0 3
rlabel polysilicon 604 -54 604 -54 0 1
rlabel polysilicon 604 -60 604 -60 0 3
rlabel polysilicon 611 -54 611 -54 0 1
rlabel polysilicon 611 -60 611 -60 0 3
rlabel polysilicon 625 -54 625 -54 0 1
rlabel polysilicon 625 -60 625 -60 0 3
rlabel polysilicon 632 -54 632 -54 0 1
rlabel polysilicon 632 -60 632 -60 0 3
rlabel polysilicon 639 -54 639 -54 0 1
rlabel polysilicon 639 -60 639 -60 0 3
rlabel polysilicon 646 -54 646 -54 0 1
rlabel polysilicon 646 -60 646 -60 0 3
rlabel polysilicon 653 -54 653 -54 0 1
rlabel polysilicon 653 -60 653 -60 0 3
rlabel polysilicon 663 -54 663 -54 0 2
rlabel polysilicon 660 -60 660 -60 0 3
rlabel polysilicon 667 -54 667 -54 0 1
rlabel polysilicon 667 -60 667 -60 0 3
rlabel polysilicon 677 -54 677 -54 0 2
rlabel polysilicon 681 -54 681 -54 0 1
rlabel polysilicon 681 -60 681 -60 0 3
rlabel polysilicon 702 -54 702 -54 0 1
rlabel polysilicon 702 -60 702 -60 0 3
rlabel polysilicon 765 -54 765 -54 0 1
rlabel polysilicon 765 -60 765 -60 0 3
rlabel polysilicon 772 -54 772 -54 0 1
rlabel polysilicon 772 -60 772 -60 0 3
rlabel polysilicon 842 -54 842 -54 0 1
rlabel polysilicon 842 -60 842 -60 0 3
rlabel polysilicon 30 -123 30 -123 0 1
rlabel polysilicon 30 -129 30 -129 0 3
rlabel polysilicon 37 -123 37 -123 0 1
rlabel polysilicon 37 -129 37 -129 0 3
rlabel polysilicon 47 -123 47 -123 0 2
rlabel polysilicon 51 -123 51 -123 0 1
rlabel polysilicon 51 -129 51 -129 0 3
rlabel polysilicon 58 -123 58 -123 0 1
rlabel polysilicon 61 -123 61 -123 0 2
rlabel polysilicon 58 -129 58 -129 0 3
rlabel polysilicon 65 -123 65 -123 0 1
rlabel polysilicon 65 -129 65 -129 0 3
rlabel polysilicon 72 -123 72 -123 0 1
rlabel polysilicon 72 -129 72 -129 0 3
rlabel polysilicon 79 -123 79 -123 0 1
rlabel polysilicon 79 -129 79 -129 0 3
rlabel polysilicon 86 -123 86 -123 0 1
rlabel polysilicon 86 -129 86 -129 0 3
rlabel polysilicon 93 -123 93 -123 0 1
rlabel polysilicon 93 -129 93 -129 0 3
rlabel polysilicon 100 -123 100 -123 0 1
rlabel polysilicon 103 -123 103 -123 0 2
rlabel polysilicon 107 -123 107 -123 0 1
rlabel polysilicon 107 -129 107 -129 0 3
rlabel polysilicon 117 -123 117 -123 0 2
rlabel polysilicon 114 -129 114 -129 0 3
rlabel polysilicon 117 -129 117 -129 0 4
rlabel polysilicon 121 -123 121 -123 0 1
rlabel polysilicon 121 -129 121 -129 0 3
rlabel polysilicon 128 -123 128 -123 0 1
rlabel polysilicon 128 -129 128 -129 0 3
rlabel polysilicon 135 -123 135 -123 0 1
rlabel polysilicon 135 -129 135 -129 0 3
rlabel polysilicon 142 -123 142 -123 0 1
rlabel polysilicon 142 -129 142 -129 0 3
rlabel polysilicon 152 -123 152 -123 0 2
rlabel polysilicon 149 -129 149 -129 0 3
rlabel polysilicon 152 -129 152 -129 0 4
rlabel polysilicon 156 -123 156 -123 0 1
rlabel polysilicon 159 -123 159 -123 0 2
rlabel polysilicon 156 -129 156 -129 0 3
rlabel polysilicon 159 -129 159 -129 0 4
rlabel polysilicon 163 -123 163 -123 0 1
rlabel polysilicon 163 -129 163 -129 0 3
rlabel polysilicon 173 -123 173 -123 0 2
rlabel polysilicon 170 -129 170 -129 0 3
rlabel polysilicon 173 -129 173 -129 0 4
rlabel polysilicon 177 -123 177 -123 0 1
rlabel polysilicon 177 -129 177 -129 0 3
rlabel polysilicon 184 -123 184 -123 0 1
rlabel polysilicon 184 -129 184 -129 0 3
rlabel polysilicon 191 -123 191 -123 0 1
rlabel polysilicon 191 -129 191 -129 0 3
rlabel polysilicon 198 -123 198 -123 0 1
rlabel polysilicon 198 -129 198 -129 0 3
rlabel polysilicon 205 -123 205 -123 0 1
rlabel polysilicon 205 -129 205 -129 0 3
rlabel polysilicon 212 -123 212 -123 0 1
rlabel polysilicon 212 -129 212 -129 0 3
rlabel polysilicon 219 -123 219 -123 0 1
rlabel polysilicon 219 -129 219 -129 0 3
rlabel polysilicon 226 -123 226 -123 0 1
rlabel polysilicon 229 -123 229 -123 0 2
rlabel polysilicon 226 -129 226 -129 0 3
rlabel polysilicon 229 -129 229 -129 0 4
rlabel polysilicon 233 -123 233 -123 0 1
rlabel polysilicon 233 -129 233 -129 0 3
rlabel polysilicon 240 -123 240 -123 0 1
rlabel polysilicon 240 -129 240 -129 0 3
rlabel polysilicon 247 -123 247 -123 0 1
rlabel polysilicon 254 -123 254 -123 0 1
rlabel polysilicon 254 -129 254 -129 0 3
rlabel polysilicon 261 -123 261 -123 0 1
rlabel polysilicon 261 -129 261 -129 0 3
rlabel polysilicon 268 -123 268 -123 0 1
rlabel polysilicon 268 -129 268 -129 0 3
rlabel polysilicon 275 -123 275 -123 0 1
rlabel polysilicon 278 -123 278 -123 0 2
rlabel polysilicon 275 -129 275 -129 0 3
rlabel polysilicon 282 -123 282 -123 0 1
rlabel polysilicon 282 -129 282 -129 0 3
rlabel polysilicon 289 -123 289 -123 0 1
rlabel polysilicon 289 -129 289 -129 0 3
rlabel polysilicon 296 -123 296 -123 0 1
rlabel polysilicon 296 -129 296 -129 0 3
rlabel polysilicon 303 -123 303 -123 0 1
rlabel polysilicon 303 -129 303 -129 0 3
rlabel polysilicon 310 -123 310 -123 0 1
rlabel polysilicon 310 -129 310 -129 0 3
rlabel polysilicon 317 -123 317 -123 0 1
rlabel polysilicon 320 -123 320 -123 0 2
rlabel polysilicon 317 -129 317 -129 0 3
rlabel polysilicon 320 -129 320 -129 0 4
rlabel polysilicon 324 -123 324 -123 0 1
rlabel polysilicon 324 -129 324 -129 0 3
rlabel polysilicon 331 -123 331 -123 0 1
rlabel polysilicon 331 -129 331 -129 0 3
rlabel polysilicon 338 -123 338 -123 0 1
rlabel polysilicon 338 -129 338 -129 0 3
rlabel polysilicon 345 -129 345 -129 0 3
rlabel polysilicon 348 -129 348 -129 0 4
rlabel polysilicon 355 -123 355 -123 0 2
rlabel polysilicon 352 -129 352 -129 0 3
rlabel polysilicon 355 -129 355 -129 0 4
rlabel polysilicon 359 -123 359 -123 0 1
rlabel polysilicon 359 -129 359 -129 0 3
rlabel polysilicon 366 -123 366 -123 0 1
rlabel polysilicon 366 -129 366 -129 0 3
rlabel polysilicon 376 -123 376 -123 0 2
rlabel polysilicon 376 -129 376 -129 0 4
rlabel polysilicon 380 -123 380 -123 0 1
rlabel polysilicon 380 -129 380 -129 0 3
rlabel polysilicon 387 -123 387 -123 0 1
rlabel polysilicon 390 -123 390 -123 0 2
rlabel polysilicon 397 -123 397 -123 0 2
rlabel polysilicon 394 -129 394 -129 0 3
rlabel polysilicon 397 -129 397 -129 0 4
rlabel polysilicon 401 -123 401 -123 0 1
rlabel polysilicon 401 -129 401 -129 0 3
rlabel polysilicon 408 -123 408 -123 0 1
rlabel polysilicon 408 -129 408 -129 0 3
rlabel polysilicon 415 -123 415 -123 0 1
rlabel polysilicon 418 -129 418 -129 0 4
rlabel polysilicon 422 -123 422 -123 0 1
rlabel polysilicon 422 -129 422 -129 0 3
rlabel polysilicon 429 -123 429 -123 0 1
rlabel polysilicon 429 -129 429 -129 0 3
rlabel polysilicon 436 -123 436 -123 0 1
rlabel polysilicon 436 -129 436 -129 0 3
rlabel polysilicon 443 -123 443 -123 0 1
rlabel polysilicon 443 -129 443 -129 0 3
rlabel polysilicon 450 -123 450 -123 0 1
rlabel polysilicon 450 -129 450 -129 0 3
rlabel polysilicon 457 -123 457 -123 0 1
rlabel polysilicon 457 -129 457 -129 0 3
rlabel polysilicon 464 -123 464 -123 0 1
rlabel polysilicon 464 -129 464 -129 0 3
rlabel polysilicon 471 -123 471 -123 0 1
rlabel polysilicon 471 -129 471 -129 0 3
rlabel polysilicon 478 -123 478 -123 0 1
rlabel polysilicon 478 -129 478 -129 0 3
rlabel polysilicon 485 -123 485 -123 0 1
rlabel polysilicon 485 -129 485 -129 0 3
rlabel polysilicon 492 -123 492 -123 0 1
rlabel polysilicon 492 -129 492 -129 0 3
rlabel polysilicon 499 -123 499 -123 0 1
rlabel polysilicon 502 -123 502 -123 0 2
rlabel polysilicon 499 -129 499 -129 0 3
rlabel polysilicon 509 -123 509 -123 0 2
rlabel polysilicon 506 -129 506 -129 0 3
rlabel polysilicon 509 -129 509 -129 0 4
rlabel polysilicon 513 -123 513 -123 0 1
rlabel polysilicon 513 -129 513 -129 0 3
rlabel polysilicon 520 -123 520 -123 0 1
rlabel polysilicon 520 -129 520 -129 0 3
rlabel polysilicon 527 -123 527 -123 0 1
rlabel polysilicon 527 -129 527 -129 0 3
rlabel polysilicon 534 -123 534 -123 0 1
rlabel polysilicon 534 -129 534 -129 0 3
rlabel polysilicon 541 -123 541 -123 0 1
rlabel polysilicon 541 -129 541 -129 0 3
rlabel polysilicon 548 -123 548 -123 0 1
rlabel polysilicon 548 -129 548 -129 0 3
rlabel polysilicon 555 -123 555 -123 0 1
rlabel polysilicon 555 -129 555 -129 0 3
rlabel polysilicon 562 -123 562 -123 0 1
rlabel polysilicon 562 -129 562 -129 0 3
rlabel polysilicon 569 -123 569 -123 0 1
rlabel polysilicon 569 -129 569 -129 0 3
rlabel polysilicon 576 -123 576 -123 0 1
rlabel polysilicon 576 -129 576 -129 0 3
rlabel polysilicon 586 -123 586 -123 0 2
rlabel polysilicon 583 -129 583 -129 0 3
rlabel polysilicon 590 -123 590 -123 0 1
rlabel polysilicon 590 -129 590 -129 0 3
rlabel polysilicon 597 -123 597 -123 0 1
rlabel polysilicon 597 -129 597 -129 0 3
rlabel polysilicon 604 -123 604 -123 0 1
rlabel polysilicon 604 -129 604 -129 0 3
rlabel polysilicon 611 -123 611 -123 0 1
rlabel polysilicon 611 -129 611 -129 0 3
rlabel polysilicon 618 -123 618 -123 0 1
rlabel polysilicon 618 -129 618 -129 0 3
rlabel polysilicon 625 -123 625 -123 0 1
rlabel polysilicon 625 -129 625 -129 0 3
rlabel polysilicon 632 -123 632 -123 0 1
rlabel polysilicon 632 -129 632 -129 0 3
rlabel polysilicon 639 -123 639 -123 0 1
rlabel polysilicon 639 -129 639 -129 0 3
rlabel polysilicon 646 -123 646 -123 0 1
rlabel polysilicon 646 -129 646 -129 0 3
rlabel polysilicon 653 -123 653 -123 0 1
rlabel polysilicon 653 -129 653 -129 0 3
rlabel polysilicon 660 -129 660 -129 0 3
rlabel polysilicon 667 -123 667 -123 0 1
rlabel polysilicon 667 -129 667 -129 0 3
rlabel polysilicon 674 -123 674 -123 0 1
rlabel polysilicon 674 -129 674 -129 0 3
rlabel polysilicon 681 -123 681 -123 0 1
rlabel polysilicon 681 -129 681 -129 0 3
rlabel polysilicon 688 -123 688 -123 0 1
rlabel polysilicon 688 -129 688 -129 0 3
rlabel polysilicon 695 -123 695 -123 0 1
rlabel polysilicon 695 -129 695 -129 0 3
rlabel polysilicon 702 -123 702 -123 0 1
rlabel polysilicon 702 -129 702 -129 0 3
rlabel polysilicon 709 -123 709 -123 0 1
rlabel polysilicon 709 -129 709 -129 0 3
rlabel polysilicon 716 -123 716 -123 0 1
rlabel polysilicon 716 -129 716 -129 0 3
rlabel polysilicon 723 -123 723 -123 0 1
rlabel polysilicon 723 -129 723 -129 0 3
rlabel polysilicon 730 -123 730 -123 0 1
rlabel polysilicon 730 -129 730 -129 0 3
rlabel polysilicon 737 -123 737 -123 0 1
rlabel polysilicon 737 -129 737 -129 0 3
rlabel polysilicon 744 -123 744 -123 0 1
rlabel polysilicon 744 -129 744 -129 0 3
rlabel polysilicon 751 -123 751 -123 0 1
rlabel polysilicon 751 -129 751 -129 0 3
rlabel polysilicon 758 -123 758 -123 0 1
rlabel polysilicon 758 -129 758 -129 0 3
rlabel polysilicon 765 -123 765 -123 0 1
rlabel polysilicon 765 -129 765 -129 0 3
rlabel polysilicon 772 -123 772 -123 0 1
rlabel polysilicon 772 -129 772 -129 0 3
rlabel polysilicon 779 -123 779 -123 0 1
rlabel polysilicon 779 -129 779 -129 0 3
rlabel polysilicon 786 -123 786 -123 0 1
rlabel polysilicon 786 -129 786 -129 0 3
rlabel polysilicon 793 -123 793 -123 0 1
rlabel polysilicon 793 -129 793 -129 0 3
rlabel polysilicon 800 -123 800 -123 0 1
rlabel polysilicon 800 -129 800 -129 0 3
rlabel polysilicon 807 -123 807 -123 0 1
rlabel polysilicon 807 -129 807 -129 0 3
rlabel polysilicon 814 -123 814 -123 0 1
rlabel polysilicon 814 -129 814 -129 0 3
rlabel polysilicon 821 -123 821 -123 0 1
rlabel polysilicon 821 -129 821 -129 0 3
rlabel polysilicon 828 -123 828 -123 0 1
rlabel polysilicon 828 -129 828 -129 0 3
rlabel polysilicon 835 -123 835 -123 0 1
rlabel polysilicon 835 -129 835 -129 0 3
rlabel polysilicon 842 -123 842 -123 0 1
rlabel polysilicon 842 -129 842 -129 0 3
rlabel polysilicon 870 -123 870 -123 0 1
rlabel polysilicon 870 -129 870 -129 0 3
rlabel polysilicon 877 -123 877 -123 0 1
rlabel polysilicon 877 -129 877 -129 0 3
rlabel polysilicon 1108 -129 1108 -129 0 3
rlabel polysilicon 23 -212 23 -212 0 1
rlabel polysilicon 23 -218 23 -218 0 3
rlabel polysilicon 30 -212 30 -212 0 1
rlabel polysilicon 30 -218 30 -218 0 3
rlabel polysilicon 37 -212 37 -212 0 1
rlabel polysilicon 37 -218 37 -218 0 3
rlabel polysilicon 44 -212 44 -212 0 1
rlabel polysilicon 44 -218 44 -218 0 3
rlabel polysilicon 51 -212 51 -212 0 1
rlabel polysilicon 51 -218 51 -218 0 3
rlabel polysilicon 58 -212 58 -212 0 1
rlabel polysilicon 58 -218 58 -218 0 3
rlabel polysilicon 65 -212 65 -212 0 1
rlabel polysilicon 65 -218 65 -218 0 3
rlabel polysilicon 72 -212 72 -212 0 1
rlabel polysilicon 72 -218 72 -218 0 3
rlabel polysilicon 79 -212 79 -212 0 1
rlabel polysilicon 79 -218 79 -218 0 3
rlabel polysilicon 89 -212 89 -212 0 2
rlabel polysilicon 93 -212 93 -212 0 1
rlabel polysilicon 93 -218 93 -218 0 3
rlabel polysilicon 100 -212 100 -212 0 1
rlabel polysilicon 100 -218 100 -218 0 3
rlabel polysilicon 110 -212 110 -212 0 2
rlabel polysilicon 114 -212 114 -212 0 1
rlabel polysilicon 114 -218 114 -218 0 3
rlabel polysilicon 124 -212 124 -212 0 2
rlabel polysilicon 121 -218 121 -218 0 3
rlabel polysilicon 128 -212 128 -212 0 1
rlabel polysilicon 128 -218 128 -218 0 3
rlabel polysilicon 135 -212 135 -212 0 1
rlabel polysilicon 135 -218 135 -218 0 3
rlabel polysilicon 142 -212 142 -212 0 1
rlabel polysilicon 145 -212 145 -212 0 2
rlabel polysilicon 142 -218 142 -218 0 3
rlabel polysilicon 152 -212 152 -212 0 2
rlabel polysilicon 149 -218 149 -218 0 3
rlabel polysilicon 152 -218 152 -218 0 4
rlabel polysilicon 156 -212 156 -212 0 1
rlabel polysilicon 156 -218 156 -218 0 3
rlabel polysilicon 163 -212 163 -212 0 1
rlabel polysilicon 163 -218 163 -218 0 3
rlabel polysilicon 170 -212 170 -212 0 1
rlabel polysilicon 170 -218 170 -218 0 3
rlabel polysilicon 180 -212 180 -212 0 2
rlabel polysilicon 177 -218 177 -218 0 3
rlabel polysilicon 184 -212 184 -212 0 1
rlabel polysilicon 184 -218 184 -218 0 3
rlabel polysilicon 191 -212 191 -212 0 1
rlabel polysilicon 191 -218 191 -218 0 3
rlabel polysilicon 198 -212 198 -212 0 1
rlabel polysilicon 198 -218 198 -218 0 3
rlabel polysilicon 205 -212 205 -212 0 1
rlabel polysilicon 208 -212 208 -212 0 2
rlabel polysilicon 205 -218 205 -218 0 3
rlabel polysilicon 208 -218 208 -218 0 4
rlabel polysilicon 212 -212 212 -212 0 1
rlabel polysilicon 215 -212 215 -212 0 2
rlabel polysilicon 212 -218 212 -218 0 3
rlabel polysilicon 219 -212 219 -212 0 1
rlabel polysilicon 219 -218 219 -218 0 3
rlabel polysilicon 222 -218 222 -218 0 4
rlabel polysilicon 229 -218 229 -218 0 4
rlabel polysilicon 233 -212 233 -212 0 1
rlabel polysilicon 240 -212 240 -212 0 1
rlabel polysilicon 240 -218 240 -218 0 3
rlabel polysilicon 250 -212 250 -212 0 2
rlabel polysilicon 247 -218 247 -218 0 3
rlabel polysilicon 254 -212 254 -212 0 1
rlabel polysilicon 254 -218 254 -218 0 3
rlabel polysilicon 261 -212 261 -212 0 1
rlabel polysilicon 261 -218 261 -218 0 3
rlabel polysilicon 268 -212 268 -212 0 1
rlabel polysilicon 268 -218 268 -218 0 3
rlabel polysilicon 275 -212 275 -212 0 1
rlabel polysilicon 275 -218 275 -218 0 3
rlabel polysilicon 282 -212 282 -212 0 1
rlabel polysilicon 282 -218 282 -218 0 3
rlabel polysilicon 289 -212 289 -212 0 1
rlabel polysilicon 289 -218 289 -218 0 3
rlabel polysilicon 296 -212 296 -212 0 1
rlabel polysilicon 299 -212 299 -212 0 2
rlabel polysilicon 299 -218 299 -218 0 4
rlabel polysilicon 303 -212 303 -212 0 1
rlabel polysilicon 303 -218 303 -218 0 3
rlabel polysilicon 310 -212 310 -212 0 1
rlabel polysilicon 310 -218 310 -218 0 3
rlabel polysilicon 317 -212 317 -212 0 1
rlabel polysilicon 317 -218 317 -218 0 3
rlabel polysilicon 324 -212 324 -212 0 1
rlabel polysilicon 327 -212 327 -212 0 2
rlabel polysilicon 324 -218 324 -218 0 3
rlabel polysilicon 334 -212 334 -212 0 2
rlabel polysilicon 331 -218 331 -218 0 3
rlabel polysilicon 334 -218 334 -218 0 4
rlabel polysilicon 338 -212 338 -212 0 1
rlabel polysilicon 338 -218 338 -218 0 3
rlabel polysilicon 345 -212 345 -212 0 1
rlabel polysilicon 348 -212 348 -212 0 2
rlabel polysilicon 352 -212 352 -212 0 1
rlabel polysilicon 352 -218 352 -218 0 3
rlabel polysilicon 359 -212 359 -212 0 1
rlabel polysilicon 362 -212 362 -212 0 2
rlabel polysilicon 359 -218 359 -218 0 3
rlabel polysilicon 362 -218 362 -218 0 4
rlabel polysilicon 366 -212 366 -212 0 1
rlabel polysilicon 366 -218 366 -218 0 3
rlabel polysilicon 373 -212 373 -212 0 1
rlabel polysilicon 373 -218 373 -218 0 3
rlabel polysilicon 380 -212 380 -212 0 1
rlabel polysilicon 380 -218 380 -218 0 3
rlabel polysilicon 387 -212 387 -212 0 1
rlabel polysilicon 387 -218 387 -218 0 3
rlabel polysilicon 394 -212 394 -212 0 1
rlabel polysilicon 397 -218 397 -218 0 4
rlabel polysilicon 401 -212 401 -212 0 1
rlabel polysilicon 401 -218 401 -218 0 3
rlabel polysilicon 404 -218 404 -218 0 4
rlabel polysilicon 408 -212 408 -212 0 1
rlabel polysilicon 408 -218 408 -218 0 3
rlabel polysilicon 415 -212 415 -212 0 1
rlabel polysilicon 415 -218 415 -218 0 3
rlabel polysilicon 422 -212 422 -212 0 1
rlabel polysilicon 422 -218 422 -218 0 3
rlabel polysilicon 429 -212 429 -212 0 1
rlabel polysilicon 429 -218 429 -218 0 3
rlabel polysilicon 436 -212 436 -212 0 1
rlabel polysilicon 436 -218 436 -218 0 3
rlabel polysilicon 443 -212 443 -212 0 1
rlabel polysilicon 443 -218 443 -218 0 3
rlabel polysilicon 450 -212 450 -212 0 1
rlabel polysilicon 450 -218 450 -218 0 3
rlabel polysilicon 457 -218 457 -218 0 3
rlabel polysilicon 464 -212 464 -212 0 1
rlabel polysilicon 464 -218 464 -218 0 3
rlabel polysilicon 471 -212 471 -212 0 1
rlabel polysilicon 471 -218 471 -218 0 3
rlabel polysilicon 478 -212 478 -212 0 1
rlabel polysilicon 478 -218 478 -218 0 3
rlabel polysilicon 485 -212 485 -212 0 1
rlabel polysilicon 485 -218 485 -218 0 3
rlabel polysilicon 492 -212 492 -212 0 1
rlabel polysilicon 495 -212 495 -212 0 2
rlabel polysilicon 495 -218 495 -218 0 4
rlabel polysilicon 499 -212 499 -212 0 1
rlabel polysilicon 499 -218 499 -218 0 3
rlabel polysilicon 506 -212 506 -212 0 1
rlabel polysilicon 506 -218 506 -218 0 3
rlabel polysilicon 513 -212 513 -212 0 1
rlabel polysilicon 513 -218 513 -218 0 3
rlabel polysilicon 520 -212 520 -212 0 1
rlabel polysilicon 523 -212 523 -212 0 2
rlabel polysilicon 520 -218 520 -218 0 3
rlabel polysilicon 527 -212 527 -212 0 1
rlabel polysilicon 527 -218 527 -218 0 3
rlabel polysilicon 534 -212 534 -212 0 1
rlabel polysilicon 534 -218 534 -218 0 3
rlabel polysilicon 541 -212 541 -212 0 1
rlabel polysilicon 541 -218 541 -218 0 3
rlabel polysilicon 548 -212 548 -212 0 1
rlabel polysilicon 548 -218 548 -218 0 3
rlabel polysilicon 555 -212 555 -212 0 1
rlabel polysilicon 555 -218 555 -218 0 3
rlabel polysilicon 562 -212 562 -212 0 1
rlabel polysilicon 562 -218 562 -218 0 3
rlabel polysilicon 569 -212 569 -212 0 1
rlabel polysilicon 569 -218 569 -218 0 3
rlabel polysilicon 576 -212 576 -212 0 1
rlabel polysilicon 579 -212 579 -212 0 2
rlabel polysilicon 576 -218 576 -218 0 3
rlabel polysilicon 579 -218 579 -218 0 4
rlabel polysilicon 583 -212 583 -212 0 1
rlabel polysilicon 583 -218 583 -218 0 3
rlabel polysilicon 590 -212 590 -212 0 1
rlabel polysilicon 590 -218 590 -218 0 3
rlabel polysilicon 597 -212 597 -212 0 1
rlabel polysilicon 597 -218 597 -218 0 3
rlabel polysilicon 604 -212 604 -212 0 1
rlabel polysilicon 604 -218 604 -218 0 3
rlabel polysilicon 611 -212 611 -212 0 1
rlabel polysilicon 611 -218 611 -218 0 3
rlabel polysilicon 618 -212 618 -212 0 1
rlabel polysilicon 618 -218 618 -218 0 3
rlabel polysilicon 621 -218 621 -218 0 4
rlabel polysilicon 625 -212 625 -212 0 1
rlabel polysilicon 628 -218 628 -218 0 4
rlabel polysilicon 632 -212 632 -212 0 1
rlabel polysilicon 632 -218 632 -218 0 3
rlabel polysilicon 639 -212 639 -212 0 1
rlabel polysilicon 639 -218 639 -218 0 3
rlabel polysilicon 646 -212 646 -212 0 1
rlabel polysilicon 646 -218 646 -218 0 3
rlabel polysilicon 653 -212 653 -212 0 1
rlabel polysilicon 656 -212 656 -212 0 2
rlabel polysilicon 653 -218 653 -218 0 3
rlabel polysilicon 660 -212 660 -212 0 1
rlabel polysilicon 660 -218 660 -218 0 3
rlabel polysilicon 667 -212 667 -212 0 1
rlabel polysilicon 667 -218 667 -218 0 3
rlabel polysilicon 674 -212 674 -212 0 1
rlabel polysilicon 674 -218 674 -218 0 3
rlabel polysilicon 681 -212 681 -212 0 1
rlabel polysilicon 681 -218 681 -218 0 3
rlabel polysilicon 688 -212 688 -212 0 1
rlabel polysilicon 688 -218 688 -218 0 3
rlabel polysilicon 695 -212 695 -212 0 1
rlabel polysilicon 695 -218 695 -218 0 3
rlabel polysilicon 702 -212 702 -212 0 1
rlabel polysilicon 702 -218 702 -218 0 3
rlabel polysilicon 709 -212 709 -212 0 1
rlabel polysilicon 709 -218 709 -218 0 3
rlabel polysilicon 716 -212 716 -212 0 1
rlabel polysilicon 716 -218 716 -218 0 3
rlabel polysilicon 723 -212 723 -212 0 1
rlabel polysilicon 723 -218 723 -218 0 3
rlabel polysilicon 730 -212 730 -212 0 1
rlabel polysilicon 730 -218 730 -218 0 3
rlabel polysilicon 737 -212 737 -212 0 1
rlabel polysilicon 740 -218 740 -218 0 4
rlabel polysilicon 744 -212 744 -212 0 1
rlabel polysilicon 744 -218 744 -218 0 3
rlabel polysilicon 751 -212 751 -212 0 1
rlabel polysilicon 751 -218 751 -218 0 3
rlabel polysilicon 758 -212 758 -212 0 1
rlabel polysilicon 758 -218 758 -218 0 3
rlabel polysilicon 765 -212 765 -212 0 1
rlabel polysilicon 765 -218 765 -218 0 3
rlabel polysilicon 772 -212 772 -212 0 1
rlabel polysilicon 772 -218 772 -218 0 3
rlabel polysilicon 779 -212 779 -212 0 1
rlabel polysilicon 779 -218 779 -218 0 3
rlabel polysilicon 786 -212 786 -212 0 1
rlabel polysilicon 786 -218 786 -218 0 3
rlabel polysilicon 793 -212 793 -212 0 1
rlabel polysilicon 793 -218 793 -218 0 3
rlabel polysilicon 800 -212 800 -212 0 1
rlabel polysilicon 800 -218 800 -218 0 3
rlabel polysilicon 807 -212 807 -212 0 1
rlabel polysilicon 807 -218 807 -218 0 3
rlabel polysilicon 814 -212 814 -212 0 1
rlabel polysilicon 814 -218 814 -218 0 3
rlabel polysilicon 821 -212 821 -212 0 1
rlabel polysilicon 821 -218 821 -218 0 3
rlabel polysilicon 828 -212 828 -212 0 1
rlabel polysilicon 828 -218 828 -218 0 3
rlabel polysilicon 835 -212 835 -212 0 1
rlabel polysilicon 835 -218 835 -218 0 3
rlabel polysilicon 842 -212 842 -212 0 1
rlabel polysilicon 842 -218 842 -218 0 3
rlabel polysilicon 849 -212 849 -212 0 1
rlabel polysilicon 849 -218 849 -218 0 3
rlabel polysilicon 856 -212 856 -212 0 1
rlabel polysilicon 856 -218 856 -218 0 3
rlabel polysilicon 863 -212 863 -212 0 1
rlabel polysilicon 863 -218 863 -218 0 3
rlabel polysilicon 870 -212 870 -212 0 1
rlabel polysilicon 870 -218 870 -218 0 3
rlabel polysilicon 877 -212 877 -212 0 1
rlabel polysilicon 877 -218 877 -218 0 3
rlabel polysilicon 884 -212 884 -212 0 1
rlabel polysilicon 884 -218 884 -218 0 3
rlabel polysilicon 891 -212 891 -212 0 1
rlabel polysilicon 891 -218 891 -218 0 3
rlabel polysilicon 898 -212 898 -212 0 1
rlabel polysilicon 898 -218 898 -218 0 3
rlabel polysilicon 905 -212 905 -212 0 1
rlabel polysilicon 905 -218 905 -218 0 3
rlabel polysilicon 912 -212 912 -212 0 1
rlabel polysilicon 912 -218 912 -218 0 3
rlabel polysilicon 919 -212 919 -212 0 1
rlabel polysilicon 919 -218 919 -218 0 3
rlabel polysilicon 926 -212 926 -212 0 1
rlabel polysilicon 926 -218 926 -218 0 3
rlabel polysilicon 933 -212 933 -212 0 1
rlabel polysilicon 933 -218 933 -218 0 3
rlabel polysilicon 940 -212 940 -212 0 1
rlabel polysilicon 940 -218 940 -218 0 3
rlabel polysilicon 947 -212 947 -212 0 1
rlabel polysilicon 947 -218 947 -218 0 3
rlabel polysilicon 954 -212 954 -212 0 1
rlabel polysilicon 954 -218 954 -218 0 3
rlabel polysilicon 1108 -212 1108 -212 0 1
rlabel polysilicon 1108 -218 1108 -218 0 3
rlabel polysilicon 16 -295 16 -295 0 1
rlabel polysilicon 16 -301 16 -301 0 3
rlabel polysilicon 23 -295 23 -295 0 1
rlabel polysilicon 23 -301 23 -301 0 3
rlabel polysilicon 30 -295 30 -295 0 1
rlabel polysilicon 30 -301 30 -301 0 3
rlabel polysilicon 37 -295 37 -295 0 1
rlabel polysilicon 37 -301 37 -301 0 3
rlabel polysilicon 47 -295 47 -295 0 2
rlabel polysilicon 47 -301 47 -301 0 4
rlabel polysilicon 51 -295 51 -295 0 1
rlabel polysilicon 51 -301 51 -301 0 3
rlabel polysilicon 58 -295 58 -295 0 1
rlabel polysilicon 58 -301 58 -301 0 3
rlabel polysilicon 65 -295 65 -295 0 1
rlabel polysilicon 68 -295 68 -295 0 2
rlabel polysilicon 65 -301 65 -301 0 3
rlabel polysilicon 68 -301 68 -301 0 4
rlabel polysilicon 72 -295 72 -295 0 1
rlabel polysilicon 72 -301 72 -301 0 3
rlabel polysilicon 79 -295 79 -295 0 1
rlabel polysilicon 79 -301 79 -301 0 3
rlabel polysilicon 86 -295 86 -295 0 1
rlabel polysilicon 86 -301 86 -301 0 3
rlabel polysilicon 93 -295 93 -295 0 1
rlabel polysilicon 93 -301 93 -301 0 3
rlabel polysilicon 100 -295 100 -295 0 1
rlabel polysilicon 100 -301 100 -301 0 3
rlabel polysilicon 103 -301 103 -301 0 4
rlabel polysilicon 107 -295 107 -295 0 1
rlabel polysilicon 107 -301 107 -301 0 3
rlabel polysilicon 114 -295 114 -295 0 1
rlabel polysilicon 117 -295 117 -295 0 2
rlabel polysilicon 117 -301 117 -301 0 4
rlabel polysilicon 121 -295 121 -295 0 1
rlabel polysilicon 121 -301 121 -301 0 3
rlabel polysilicon 128 -301 128 -301 0 3
rlabel polysilicon 131 -301 131 -301 0 4
rlabel polysilicon 135 -295 135 -295 0 1
rlabel polysilicon 138 -295 138 -295 0 2
rlabel polysilicon 135 -301 135 -301 0 3
rlabel polysilicon 142 -295 142 -295 0 1
rlabel polysilicon 142 -301 142 -301 0 3
rlabel polysilicon 149 -295 149 -295 0 1
rlabel polysilicon 149 -301 149 -301 0 3
rlabel polysilicon 156 -295 156 -295 0 1
rlabel polysilicon 156 -301 156 -301 0 3
rlabel polysilicon 166 -295 166 -295 0 2
rlabel polysilicon 163 -301 163 -301 0 3
rlabel polysilicon 166 -301 166 -301 0 4
rlabel polysilicon 170 -295 170 -295 0 1
rlabel polysilicon 173 -295 173 -295 0 2
rlabel polysilicon 170 -301 170 -301 0 3
rlabel polysilicon 173 -301 173 -301 0 4
rlabel polysilicon 177 -295 177 -295 0 1
rlabel polysilicon 177 -301 177 -301 0 3
rlabel polysilicon 184 -295 184 -295 0 1
rlabel polysilicon 184 -301 184 -301 0 3
rlabel polysilicon 191 -295 191 -295 0 1
rlabel polysilicon 194 -295 194 -295 0 2
rlabel polysilicon 191 -301 191 -301 0 3
rlabel polysilicon 194 -301 194 -301 0 4
rlabel polysilicon 198 -295 198 -295 0 1
rlabel polysilicon 198 -301 198 -301 0 3
rlabel polysilicon 205 -295 205 -295 0 1
rlabel polysilicon 205 -301 205 -301 0 3
rlabel polysilicon 208 -301 208 -301 0 4
rlabel polysilicon 212 -295 212 -295 0 1
rlabel polysilicon 212 -301 212 -301 0 3
rlabel polysilicon 219 -295 219 -295 0 1
rlabel polysilicon 219 -301 219 -301 0 3
rlabel polysilicon 226 -295 226 -295 0 1
rlabel polysilicon 226 -301 226 -301 0 3
rlabel polysilicon 233 -295 233 -295 0 1
rlabel polysilicon 233 -301 233 -301 0 3
rlabel polysilicon 240 -295 240 -295 0 1
rlabel polysilicon 240 -301 240 -301 0 3
rlabel polysilicon 247 -295 247 -295 0 1
rlabel polysilicon 247 -301 247 -301 0 3
rlabel polysilicon 254 -295 254 -295 0 1
rlabel polysilicon 257 -295 257 -295 0 2
rlabel polysilicon 261 -295 261 -295 0 1
rlabel polysilicon 261 -301 261 -301 0 3
rlabel polysilicon 268 -295 268 -295 0 1
rlabel polysilicon 268 -301 268 -301 0 3
rlabel polysilicon 275 -295 275 -295 0 1
rlabel polysilicon 275 -301 275 -301 0 3
rlabel polysilicon 282 -295 282 -295 0 1
rlabel polysilicon 282 -301 282 -301 0 3
rlabel polysilicon 289 -295 289 -295 0 1
rlabel polysilicon 289 -301 289 -301 0 3
rlabel polysilicon 296 -295 296 -295 0 1
rlabel polysilicon 299 -295 299 -295 0 2
rlabel polysilicon 296 -301 296 -301 0 3
rlabel polysilicon 299 -301 299 -301 0 4
rlabel polysilicon 303 -295 303 -295 0 1
rlabel polysilicon 303 -301 303 -301 0 3
rlabel polysilicon 310 -295 310 -295 0 1
rlabel polysilicon 310 -301 310 -301 0 3
rlabel polysilicon 317 -295 317 -295 0 1
rlabel polysilicon 320 -301 320 -301 0 4
rlabel polysilicon 324 -295 324 -295 0 1
rlabel polysilicon 324 -301 324 -301 0 3
rlabel polysilicon 331 -295 331 -295 0 1
rlabel polysilicon 331 -301 331 -301 0 3
rlabel polysilicon 338 -295 338 -295 0 1
rlabel polysilicon 338 -301 338 -301 0 3
rlabel polysilicon 345 -295 345 -295 0 1
rlabel polysilicon 345 -301 345 -301 0 3
rlabel polysilicon 355 -295 355 -295 0 2
rlabel polysilicon 352 -301 352 -301 0 3
rlabel polysilicon 355 -301 355 -301 0 4
rlabel polysilicon 362 -295 362 -295 0 2
rlabel polysilicon 359 -301 359 -301 0 3
rlabel polysilicon 366 -295 366 -295 0 1
rlabel polysilicon 366 -301 366 -301 0 3
rlabel polysilicon 373 -295 373 -295 0 1
rlabel polysilicon 373 -301 373 -301 0 3
rlabel polysilicon 380 -295 380 -295 0 1
rlabel polysilicon 380 -301 380 -301 0 3
rlabel polysilicon 387 -295 387 -295 0 1
rlabel polysilicon 387 -301 387 -301 0 3
rlabel polysilicon 394 -295 394 -295 0 1
rlabel polysilicon 397 -301 397 -301 0 4
rlabel polysilicon 401 -295 401 -295 0 1
rlabel polysilicon 401 -301 401 -301 0 3
rlabel polysilicon 404 -301 404 -301 0 4
rlabel polysilicon 408 -295 408 -295 0 1
rlabel polysilicon 408 -301 408 -301 0 3
rlabel polysilicon 415 -295 415 -295 0 1
rlabel polysilicon 415 -301 415 -301 0 3
rlabel polysilicon 422 -295 422 -295 0 1
rlabel polysilicon 422 -301 422 -301 0 3
rlabel polysilicon 429 -295 429 -295 0 1
rlabel polysilicon 429 -301 429 -301 0 3
rlabel polysilicon 436 -295 436 -295 0 1
rlabel polysilicon 436 -301 436 -301 0 3
rlabel polysilicon 439 -301 439 -301 0 4
rlabel polysilicon 443 -295 443 -295 0 1
rlabel polysilicon 443 -301 443 -301 0 3
rlabel polysilicon 450 -295 450 -295 0 1
rlabel polysilicon 450 -301 450 -301 0 3
rlabel polysilicon 457 -295 457 -295 0 1
rlabel polysilicon 457 -301 457 -301 0 3
rlabel polysilicon 467 -295 467 -295 0 2
rlabel polysilicon 464 -301 464 -301 0 3
rlabel polysilicon 467 -301 467 -301 0 4
rlabel polysilicon 471 -295 471 -295 0 1
rlabel polysilicon 471 -301 471 -301 0 3
rlabel polysilicon 478 -295 478 -295 0 1
rlabel polysilicon 478 -301 478 -301 0 3
rlabel polysilicon 485 -295 485 -295 0 1
rlabel polysilicon 488 -295 488 -295 0 2
rlabel polysilicon 485 -301 485 -301 0 3
rlabel polysilicon 488 -301 488 -301 0 4
rlabel polysilicon 492 -295 492 -295 0 1
rlabel polysilicon 492 -301 492 -301 0 3
rlabel polysilicon 499 -295 499 -295 0 1
rlabel polysilicon 502 -295 502 -295 0 2
rlabel polysilicon 506 -295 506 -295 0 1
rlabel polysilicon 506 -301 506 -301 0 3
rlabel polysilicon 513 -295 513 -295 0 1
rlabel polysilicon 513 -301 513 -301 0 3
rlabel polysilicon 520 -295 520 -295 0 1
rlabel polysilicon 523 -301 523 -301 0 4
rlabel polysilicon 527 -295 527 -295 0 1
rlabel polysilicon 527 -301 527 -301 0 3
rlabel polysilicon 534 -295 534 -295 0 1
rlabel polysilicon 534 -301 534 -301 0 3
rlabel polysilicon 541 -295 541 -295 0 1
rlabel polysilicon 541 -301 541 -301 0 3
rlabel polysilicon 548 -295 548 -295 0 1
rlabel polysilicon 548 -301 548 -301 0 3
rlabel polysilicon 555 -295 555 -295 0 1
rlabel polysilicon 555 -301 555 -301 0 3
rlabel polysilicon 562 -295 562 -295 0 1
rlabel polysilicon 562 -301 562 -301 0 3
rlabel polysilicon 569 -295 569 -295 0 1
rlabel polysilicon 569 -301 569 -301 0 3
rlabel polysilicon 576 -295 576 -295 0 1
rlabel polysilicon 576 -301 576 -301 0 3
rlabel polysilicon 583 -295 583 -295 0 1
rlabel polysilicon 583 -301 583 -301 0 3
rlabel polysilicon 590 -295 590 -295 0 1
rlabel polysilicon 590 -301 590 -301 0 3
rlabel polysilicon 597 -295 597 -295 0 1
rlabel polysilicon 597 -301 597 -301 0 3
rlabel polysilicon 604 -295 604 -295 0 1
rlabel polysilicon 604 -301 604 -301 0 3
rlabel polysilicon 611 -295 611 -295 0 1
rlabel polysilicon 611 -301 611 -301 0 3
rlabel polysilicon 618 -295 618 -295 0 1
rlabel polysilicon 618 -301 618 -301 0 3
rlabel polysilicon 625 -295 625 -295 0 1
rlabel polysilicon 625 -301 625 -301 0 3
rlabel polysilicon 632 -295 632 -295 0 1
rlabel polysilicon 632 -301 632 -301 0 3
rlabel polysilicon 639 -295 639 -295 0 1
rlabel polysilicon 639 -301 639 -301 0 3
rlabel polysilicon 646 -295 646 -295 0 1
rlabel polysilicon 646 -301 646 -301 0 3
rlabel polysilicon 653 -295 653 -295 0 1
rlabel polysilicon 653 -301 653 -301 0 3
rlabel polysilicon 663 -295 663 -295 0 2
rlabel polysilicon 667 -295 667 -295 0 1
rlabel polysilicon 667 -301 667 -301 0 3
rlabel polysilicon 674 -295 674 -295 0 1
rlabel polysilicon 674 -301 674 -301 0 3
rlabel polysilicon 681 -295 681 -295 0 1
rlabel polysilicon 681 -301 681 -301 0 3
rlabel polysilicon 688 -295 688 -295 0 1
rlabel polysilicon 688 -301 688 -301 0 3
rlabel polysilicon 695 -295 695 -295 0 1
rlabel polysilicon 695 -301 695 -301 0 3
rlabel polysilicon 702 -295 702 -295 0 1
rlabel polysilicon 702 -301 702 -301 0 3
rlabel polysilicon 709 -295 709 -295 0 1
rlabel polysilicon 709 -301 709 -301 0 3
rlabel polysilicon 716 -295 716 -295 0 1
rlabel polysilicon 716 -301 716 -301 0 3
rlabel polysilicon 723 -295 723 -295 0 1
rlabel polysilicon 723 -301 723 -301 0 3
rlabel polysilicon 730 -295 730 -295 0 1
rlabel polysilicon 730 -301 730 -301 0 3
rlabel polysilicon 737 -295 737 -295 0 1
rlabel polysilicon 737 -301 737 -301 0 3
rlabel polysilicon 744 -295 744 -295 0 1
rlabel polysilicon 744 -301 744 -301 0 3
rlabel polysilicon 751 -295 751 -295 0 1
rlabel polysilicon 751 -301 751 -301 0 3
rlabel polysilicon 758 -295 758 -295 0 1
rlabel polysilicon 758 -301 758 -301 0 3
rlabel polysilicon 765 -295 765 -295 0 1
rlabel polysilicon 765 -301 765 -301 0 3
rlabel polysilicon 772 -295 772 -295 0 1
rlabel polysilicon 772 -301 772 -301 0 3
rlabel polysilicon 779 -295 779 -295 0 1
rlabel polysilicon 779 -301 779 -301 0 3
rlabel polysilicon 786 -295 786 -295 0 1
rlabel polysilicon 786 -301 786 -301 0 3
rlabel polysilicon 793 -295 793 -295 0 1
rlabel polysilicon 793 -301 793 -301 0 3
rlabel polysilicon 800 -295 800 -295 0 1
rlabel polysilicon 800 -301 800 -301 0 3
rlabel polysilicon 807 -295 807 -295 0 1
rlabel polysilicon 807 -301 807 -301 0 3
rlabel polysilicon 814 -295 814 -295 0 1
rlabel polysilicon 814 -301 814 -301 0 3
rlabel polysilicon 821 -295 821 -295 0 1
rlabel polysilicon 821 -301 821 -301 0 3
rlabel polysilicon 828 -295 828 -295 0 1
rlabel polysilicon 828 -301 828 -301 0 3
rlabel polysilicon 835 -295 835 -295 0 1
rlabel polysilicon 835 -301 835 -301 0 3
rlabel polysilicon 842 -295 842 -295 0 1
rlabel polysilicon 842 -301 842 -301 0 3
rlabel polysilicon 849 -295 849 -295 0 1
rlabel polysilicon 849 -301 849 -301 0 3
rlabel polysilicon 856 -295 856 -295 0 1
rlabel polysilicon 856 -301 856 -301 0 3
rlabel polysilicon 863 -295 863 -295 0 1
rlabel polysilicon 863 -301 863 -301 0 3
rlabel polysilicon 870 -295 870 -295 0 1
rlabel polysilicon 870 -301 870 -301 0 3
rlabel polysilicon 877 -295 877 -295 0 1
rlabel polysilicon 877 -301 877 -301 0 3
rlabel polysilicon 887 -295 887 -295 0 2
rlabel polysilicon 884 -301 884 -301 0 3
rlabel polysilicon 894 -301 894 -301 0 4
rlabel polysilicon 898 -295 898 -295 0 1
rlabel polysilicon 905 -295 905 -295 0 1
rlabel polysilicon 908 -295 908 -295 0 2
rlabel polysilicon 912 -295 912 -295 0 1
rlabel polysilicon 912 -301 912 -301 0 3
rlabel polysilicon 919 -295 919 -295 0 1
rlabel polysilicon 919 -301 919 -301 0 3
rlabel polysilicon 1108 -295 1108 -295 0 1
rlabel polysilicon 1108 -301 1108 -301 0 3
rlabel polysilicon 9 -390 9 -390 0 1
rlabel polysilicon 9 -396 9 -396 0 3
rlabel polysilicon 16 -390 16 -390 0 1
rlabel polysilicon 23 -390 23 -390 0 1
rlabel polysilicon 23 -396 23 -396 0 3
rlabel polysilicon 30 -396 30 -396 0 3
rlabel polysilicon 37 -390 37 -390 0 1
rlabel polysilicon 37 -396 37 -396 0 3
rlabel polysilicon 44 -390 44 -390 0 1
rlabel polysilicon 44 -396 44 -396 0 3
rlabel polysilicon 51 -390 51 -390 0 1
rlabel polysilicon 51 -396 51 -396 0 3
rlabel polysilicon 58 -390 58 -390 0 1
rlabel polysilicon 58 -396 58 -396 0 3
rlabel polysilicon 65 -390 65 -390 0 1
rlabel polysilicon 68 -390 68 -390 0 2
rlabel polysilicon 72 -390 72 -390 0 1
rlabel polysilicon 72 -396 72 -396 0 3
rlabel polysilicon 79 -390 79 -390 0 1
rlabel polysilicon 82 -390 82 -390 0 2
rlabel polysilicon 79 -396 79 -396 0 3
rlabel polysilicon 82 -396 82 -396 0 4
rlabel polysilicon 86 -390 86 -390 0 1
rlabel polysilicon 86 -396 86 -396 0 3
rlabel polysilicon 96 -390 96 -390 0 2
rlabel polysilicon 93 -396 93 -396 0 3
rlabel polysilicon 96 -396 96 -396 0 4
rlabel polysilicon 100 -390 100 -390 0 1
rlabel polysilicon 100 -396 100 -396 0 3
rlabel polysilicon 107 -390 107 -390 0 1
rlabel polysilicon 110 -390 110 -390 0 2
rlabel polysilicon 110 -396 110 -396 0 4
rlabel polysilicon 114 -390 114 -390 0 1
rlabel polysilicon 117 -396 117 -396 0 4
rlabel polysilicon 121 -390 121 -390 0 1
rlabel polysilicon 124 -390 124 -390 0 2
rlabel polysilicon 121 -396 121 -396 0 3
rlabel polysilicon 128 -390 128 -390 0 1
rlabel polysilicon 128 -396 128 -396 0 3
rlabel polysilicon 135 -390 135 -390 0 1
rlabel polysilicon 138 -396 138 -396 0 4
rlabel polysilicon 142 -390 142 -390 0 1
rlabel polysilicon 142 -396 142 -396 0 3
rlabel polysilicon 149 -390 149 -390 0 1
rlabel polysilicon 149 -396 149 -396 0 3
rlabel polysilicon 159 -390 159 -390 0 2
rlabel polysilicon 156 -396 156 -396 0 3
rlabel polysilicon 163 -390 163 -390 0 1
rlabel polysilicon 163 -396 163 -396 0 3
rlabel polysilicon 170 -390 170 -390 0 1
rlabel polysilicon 173 -390 173 -390 0 2
rlabel polysilicon 170 -396 170 -396 0 3
rlabel polysilicon 173 -396 173 -396 0 4
rlabel polysilicon 177 -390 177 -390 0 1
rlabel polysilicon 177 -396 177 -396 0 3
rlabel polysilicon 187 -390 187 -390 0 2
rlabel polysilicon 184 -396 184 -396 0 3
rlabel polysilicon 187 -396 187 -396 0 4
rlabel polysilicon 191 -390 191 -390 0 1
rlabel polysilicon 191 -396 191 -396 0 3
rlabel polysilicon 198 -390 198 -390 0 1
rlabel polysilicon 198 -396 198 -396 0 3
rlabel polysilicon 205 -390 205 -390 0 1
rlabel polysilicon 205 -396 205 -396 0 3
rlabel polysilicon 215 -390 215 -390 0 2
rlabel polysilicon 219 -390 219 -390 0 1
rlabel polysilicon 219 -396 219 -396 0 3
rlabel polysilicon 226 -390 226 -390 0 1
rlabel polysilicon 226 -396 226 -396 0 3
rlabel polysilicon 233 -390 233 -390 0 1
rlabel polysilicon 233 -396 233 -396 0 3
rlabel polysilicon 240 -390 240 -390 0 1
rlabel polysilicon 240 -396 240 -396 0 3
rlabel polysilicon 247 -390 247 -390 0 1
rlabel polysilicon 250 -390 250 -390 0 2
rlabel polysilicon 247 -396 247 -396 0 3
rlabel polysilicon 250 -396 250 -396 0 4
rlabel polysilicon 254 -390 254 -390 0 1
rlabel polysilicon 257 -390 257 -390 0 2
rlabel polysilicon 254 -396 254 -396 0 3
rlabel polysilicon 261 -390 261 -390 0 1
rlabel polysilicon 264 -390 264 -390 0 2
rlabel polysilicon 261 -396 261 -396 0 3
rlabel polysilicon 264 -396 264 -396 0 4
rlabel polysilicon 268 -390 268 -390 0 1
rlabel polysilicon 268 -396 268 -396 0 3
rlabel polysilicon 275 -390 275 -390 0 1
rlabel polysilicon 275 -396 275 -396 0 3
rlabel polysilicon 282 -390 282 -390 0 1
rlabel polysilicon 282 -396 282 -396 0 3
rlabel polysilicon 289 -390 289 -390 0 1
rlabel polysilicon 289 -396 289 -396 0 3
rlabel polysilicon 296 -390 296 -390 0 1
rlabel polysilicon 296 -396 296 -396 0 3
rlabel polysilicon 303 -390 303 -390 0 1
rlabel polysilicon 306 -390 306 -390 0 2
rlabel polysilicon 306 -396 306 -396 0 4
rlabel polysilicon 310 -390 310 -390 0 1
rlabel polysilicon 310 -396 310 -396 0 3
rlabel polysilicon 317 -390 317 -390 0 1
rlabel polysilicon 320 -390 320 -390 0 2
rlabel polysilicon 317 -396 317 -396 0 3
rlabel polysilicon 320 -396 320 -396 0 4
rlabel polysilicon 324 -390 324 -390 0 1
rlabel polysilicon 324 -396 324 -396 0 3
rlabel polysilicon 327 -396 327 -396 0 4
rlabel polysilicon 331 -390 331 -390 0 1
rlabel polysilicon 331 -396 331 -396 0 3
rlabel polysilicon 341 -390 341 -390 0 2
rlabel polysilicon 341 -396 341 -396 0 4
rlabel polysilicon 345 -390 345 -390 0 1
rlabel polysilicon 345 -396 345 -396 0 3
rlabel polysilicon 352 -390 352 -390 0 1
rlabel polysilicon 352 -396 352 -396 0 3
rlabel polysilicon 359 -390 359 -390 0 1
rlabel polysilicon 359 -396 359 -396 0 3
rlabel polysilicon 366 -390 366 -390 0 1
rlabel polysilicon 366 -396 366 -396 0 3
rlabel polysilicon 373 -390 373 -390 0 1
rlabel polysilicon 373 -396 373 -396 0 3
rlabel polysilicon 380 -396 380 -396 0 3
rlabel polysilicon 383 -396 383 -396 0 4
rlabel polysilicon 387 -390 387 -390 0 1
rlabel polysilicon 387 -396 387 -396 0 3
rlabel polysilicon 394 -390 394 -390 0 1
rlabel polysilicon 397 -390 397 -390 0 2
rlabel polysilicon 394 -396 394 -396 0 3
rlabel polysilicon 401 -390 401 -390 0 1
rlabel polysilicon 401 -396 401 -396 0 3
rlabel polysilicon 408 -390 408 -390 0 1
rlabel polysilicon 408 -396 408 -396 0 3
rlabel polysilicon 415 -390 415 -390 0 1
rlabel polysilicon 415 -396 415 -396 0 3
rlabel polysilicon 422 -390 422 -390 0 1
rlabel polysilicon 422 -396 422 -396 0 3
rlabel polysilicon 429 -390 429 -390 0 1
rlabel polysilicon 429 -396 429 -396 0 3
rlabel polysilicon 436 -390 436 -390 0 1
rlabel polysilicon 436 -396 436 -396 0 3
rlabel polysilicon 443 -390 443 -390 0 1
rlabel polysilicon 443 -396 443 -396 0 3
rlabel polysilicon 450 -390 450 -390 0 1
rlabel polysilicon 450 -396 450 -396 0 3
rlabel polysilicon 457 -390 457 -390 0 1
rlabel polysilicon 457 -396 457 -396 0 3
rlabel polysilicon 464 -390 464 -390 0 1
rlabel polysilicon 464 -396 464 -396 0 3
rlabel polysilicon 474 -390 474 -390 0 2
rlabel polysilicon 471 -396 471 -396 0 3
rlabel polysilicon 474 -396 474 -396 0 4
rlabel polysilicon 478 -390 478 -390 0 1
rlabel polysilicon 478 -396 478 -396 0 3
rlabel polysilicon 485 -390 485 -390 0 1
rlabel polysilicon 485 -396 485 -396 0 3
rlabel polysilicon 492 -396 492 -396 0 3
rlabel polysilicon 495 -396 495 -396 0 4
rlabel polysilicon 499 -390 499 -390 0 1
rlabel polysilicon 499 -396 499 -396 0 3
rlabel polysilicon 506 -390 506 -390 0 1
rlabel polysilicon 506 -396 506 -396 0 3
rlabel polysilicon 513 -390 513 -390 0 1
rlabel polysilicon 516 -390 516 -390 0 2
rlabel polysilicon 516 -396 516 -396 0 4
rlabel polysilicon 520 -390 520 -390 0 1
rlabel polysilicon 520 -396 520 -396 0 3
rlabel polysilicon 527 -390 527 -390 0 1
rlabel polysilicon 527 -396 527 -396 0 3
rlabel polysilicon 534 -390 534 -390 0 1
rlabel polysilicon 534 -396 534 -396 0 3
rlabel polysilicon 541 -390 541 -390 0 1
rlabel polysilicon 544 -390 544 -390 0 2
rlabel polysilicon 541 -396 541 -396 0 3
rlabel polysilicon 544 -396 544 -396 0 4
rlabel polysilicon 548 -390 548 -390 0 1
rlabel polysilicon 548 -396 548 -396 0 3
rlabel polysilicon 555 -390 555 -390 0 1
rlabel polysilicon 555 -396 555 -396 0 3
rlabel polysilicon 562 -390 562 -390 0 1
rlabel polysilicon 562 -396 562 -396 0 3
rlabel polysilicon 569 -390 569 -390 0 1
rlabel polysilicon 569 -396 569 -396 0 3
rlabel polysilicon 576 -390 576 -390 0 1
rlabel polysilicon 576 -396 576 -396 0 3
rlabel polysilicon 583 -390 583 -390 0 1
rlabel polysilicon 583 -396 583 -396 0 3
rlabel polysilicon 590 -390 590 -390 0 1
rlabel polysilicon 590 -396 590 -396 0 3
rlabel polysilicon 597 -390 597 -390 0 1
rlabel polysilicon 597 -396 597 -396 0 3
rlabel polysilicon 604 -390 604 -390 0 1
rlabel polysilicon 604 -396 604 -396 0 3
rlabel polysilicon 611 -390 611 -390 0 1
rlabel polysilicon 611 -396 611 -396 0 3
rlabel polysilicon 618 -390 618 -390 0 1
rlabel polysilicon 618 -396 618 -396 0 3
rlabel polysilicon 628 -390 628 -390 0 2
rlabel polysilicon 625 -396 625 -396 0 3
rlabel polysilicon 628 -396 628 -396 0 4
rlabel polysilicon 632 -390 632 -390 0 1
rlabel polysilicon 632 -396 632 -396 0 3
rlabel polysilicon 639 -390 639 -390 0 1
rlabel polysilicon 639 -396 639 -396 0 3
rlabel polysilicon 646 -390 646 -390 0 1
rlabel polysilicon 646 -396 646 -396 0 3
rlabel polysilicon 653 -390 653 -390 0 1
rlabel polysilicon 653 -396 653 -396 0 3
rlabel polysilicon 660 -390 660 -390 0 1
rlabel polysilicon 660 -396 660 -396 0 3
rlabel polysilicon 670 -390 670 -390 0 2
rlabel polysilicon 667 -396 667 -396 0 3
rlabel polysilicon 674 -390 674 -390 0 1
rlabel polysilicon 674 -396 674 -396 0 3
rlabel polysilicon 681 -390 681 -390 0 1
rlabel polysilicon 681 -396 681 -396 0 3
rlabel polysilicon 688 -390 688 -390 0 1
rlabel polysilicon 688 -396 688 -396 0 3
rlabel polysilicon 695 -390 695 -390 0 1
rlabel polysilicon 695 -396 695 -396 0 3
rlabel polysilicon 702 -390 702 -390 0 1
rlabel polysilicon 702 -396 702 -396 0 3
rlabel polysilicon 709 -390 709 -390 0 1
rlabel polysilicon 709 -396 709 -396 0 3
rlabel polysilicon 716 -390 716 -390 0 1
rlabel polysilicon 716 -396 716 -396 0 3
rlabel polysilicon 723 -390 723 -390 0 1
rlabel polysilicon 723 -396 723 -396 0 3
rlabel polysilicon 730 -390 730 -390 0 1
rlabel polysilicon 730 -396 730 -396 0 3
rlabel polysilicon 737 -390 737 -390 0 1
rlabel polysilicon 737 -396 737 -396 0 3
rlabel polysilicon 744 -390 744 -390 0 1
rlabel polysilicon 744 -396 744 -396 0 3
rlabel polysilicon 751 -390 751 -390 0 1
rlabel polysilicon 751 -396 751 -396 0 3
rlabel polysilicon 758 -390 758 -390 0 1
rlabel polysilicon 758 -396 758 -396 0 3
rlabel polysilicon 765 -390 765 -390 0 1
rlabel polysilicon 765 -396 765 -396 0 3
rlabel polysilicon 772 -390 772 -390 0 1
rlabel polysilicon 772 -396 772 -396 0 3
rlabel polysilicon 779 -390 779 -390 0 1
rlabel polysilicon 779 -396 779 -396 0 3
rlabel polysilicon 786 -390 786 -390 0 1
rlabel polysilicon 786 -396 786 -396 0 3
rlabel polysilicon 793 -390 793 -390 0 1
rlabel polysilicon 793 -396 793 -396 0 3
rlabel polysilicon 800 -390 800 -390 0 1
rlabel polysilicon 800 -396 800 -396 0 3
rlabel polysilicon 807 -390 807 -390 0 1
rlabel polysilicon 807 -396 807 -396 0 3
rlabel polysilicon 814 -390 814 -390 0 1
rlabel polysilicon 814 -396 814 -396 0 3
rlabel polysilicon 821 -390 821 -390 0 1
rlabel polysilicon 821 -396 821 -396 0 3
rlabel polysilicon 828 -390 828 -390 0 1
rlabel polysilicon 828 -396 828 -396 0 3
rlabel polysilicon 835 -390 835 -390 0 1
rlabel polysilicon 835 -396 835 -396 0 3
rlabel polysilicon 842 -390 842 -390 0 1
rlabel polysilicon 842 -396 842 -396 0 3
rlabel polysilicon 849 -390 849 -390 0 1
rlabel polysilicon 849 -396 849 -396 0 3
rlabel polysilicon 856 -390 856 -390 0 1
rlabel polysilicon 856 -396 856 -396 0 3
rlabel polysilicon 863 -390 863 -390 0 1
rlabel polysilicon 863 -396 863 -396 0 3
rlabel polysilicon 870 -390 870 -390 0 1
rlabel polysilicon 870 -396 870 -396 0 3
rlabel polysilicon 877 -390 877 -390 0 1
rlabel polysilicon 880 -390 880 -390 0 2
rlabel polysilicon 877 -396 877 -396 0 3
rlabel polysilicon 884 -390 884 -390 0 1
rlabel polysilicon 887 -390 887 -390 0 2
rlabel polysilicon 884 -396 884 -396 0 3
rlabel polysilicon 891 -390 891 -390 0 1
rlabel polysilicon 891 -396 891 -396 0 3
rlabel polysilicon 898 -390 898 -390 0 1
rlabel polysilicon 898 -396 898 -396 0 3
rlabel polysilicon 905 -390 905 -390 0 1
rlabel polysilicon 905 -396 905 -396 0 3
rlabel polysilicon 933 -390 933 -390 0 1
rlabel polysilicon 933 -396 933 -396 0 3
rlabel polysilicon 1108 -390 1108 -390 0 1
rlabel polysilicon 1108 -396 1108 -396 0 3
rlabel polysilicon 2 -479 2 -479 0 1
rlabel polysilicon 2 -485 2 -485 0 3
rlabel polysilicon 12 -479 12 -479 0 2
rlabel polysilicon 16 -479 16 -479 0 1
rlabel polysilicon 16 -485 16 -485 0 3
rlabel polysilicon 23 -479 23 -479 0 1
rlabel polysilicon 23 -485 23 -485 0 3
rlabel polysilicon 30 -479 30 -479 0 1
rlabel polysilicon 30 -485 30 -485 0 3
rlabel polysilicon 37 -479 37 -479 0 1
rlabel polysilicon 37 -485 37 -485 0 3
rlabel polysilicon 44 -479 44 -479 0 1
rlabel polysilicon 44 -485 44 -485 0 3
rlabel polysilicon 51 -479 51 -479 0 1
rlabel polysilicon 51 -485 51 -485 0 3
rlabel polysilicon 61 -479 61 -479 0 2
rlabel polysilicon 61 -485 61 -485 0 4
rlabel polysilicon 65 -479 65 -479 0 1
rlabel polysilicon 68 -479 68 -479 0 2
rlabel polysilicon 72 -479 72 -479 0 1
rlabel polysilicon 72 -485 72 -485 0 3
rlabel polysilicon 79 -479 79 -479 0 1
rlabel polysilicon 79 -485 79 -485 0 3
rlabel polysilicon 86 -479 86 -479 0 1
rlabel polysilicon 86 -485 86 -485 0 3
rlabel polysilicon 93 -479 93 -479 0 1
rlabel polysilicon 93 -485 93 -485 0 3
rlabel polysilicon 100 -479 100 -479 0 1
rlabel polysilicon 100 -485 100 -485 0 3
rlabel polysilicon 107 -479 107 -479 0 1
rlabel polysilicon 107 -485 107 -485 0 3
rlabel polysilicon 114 -479 114 -479 0 1
rlabel polysilicon 114 -485 114 -485 0 3
rlabel polysilicon 121 -479 121 -479 0 1
rlabel polysilicon 124 -479 124 -479 0 2
rlabel polysilicon 131 -479 131 -479 0 2
rlabel polysilicon 128 -485 128 -485 0 3
rlabel polysilicon 135 -479 135 -479 0 1
rlabel polysilicon 135 -485 135 -485 0 3
rlabel polysilicon 142 -479 142 -479 0 1
rlabel polysilicon 145 -479 145 -479 0 2
rlabel polysilicon 142 -485 142 -485 0 3
rlabel polysilicon 145 -485 145 -485 0 4
rlabel polysilicon 149 -479 149 -479 0 1
rlabel polysilicon 149 -485 149 -485 0 3
rlabel polysilicon 156 -479 156 -479 0 1
rlabel polysilicon 156 -485 156 -485 0 3
rlabel polysilicon 163 -479 163 -479 0 1
rlabel polysilicon 163 -485 163 -485 0 3
rlabel polysilicon 170 -479 170 -479 0 1
rlabel polysilicon 170 -485 170 -485 0 3
rlabel polysilicon 177 -479 177 -479 0 1
rlabel polysilicon 180 -479 180 -479 0 2
rlabel polysilicon 184 -479 184 -479 0 1
rlabel polysilicon 184 -485 184 -485 0 3
rlabel polysilicon 191 -479 191 -479 0 1
rlabel polysilicon 191 -485 191 -485 0 3
rlabel polysilicon 198 -479 198 -479 0 1
rlabel polysilicon 198 -485 198 -485 0 3
rlabel polysilicon 205 -479 205 -479 0 1
rlabel polysilicon 208 -485 208 -485 0 4
rlabel polysilicon 212 -479 212 -479 0 1
rlabel polysilicon 212 -485 212 -485 0 3
rlabel polysilicon 219 -479 219 -479 0 1
rlabel polysilicon 219 -485 219 -485 0 3
rlabel polysilicon 226 -479 226 -479 0 1
rlabel polysilicon 226 -485 226 -485 0 3
rlabel polysilicon 233 -479 233 -479 0 1
rlabel polysilicon 233 -485 233 -485 0 3
rlabel polysilicon 240 -479 240 -479 0 1
rlabel polysilicon 240 -485 240 -485 0 3
rlabel polysilicon 247 -479 247 -479 0 1
rlabel polysilicon 247 -485 247 -485 0 3
rlabel polysilicon 254 -479 254 -479 0 1
rlabel polysilicon 254 -485 254 -485 0 3
rlabel polysilicon 261 -479 261 -479 0 1
rlabel polysilicon 261 -485 261 -485 0 3
rlabel polysilicon 268 -479 268 -479 0 1
rlabel polysilicon 268 -485 268 -485 0 3
rlabel polysilicon 275 -479 275 -479 0 1
rlabel polysilicon 275 -485 275 -485 0 3
rlabel polysilicon 282 -485 282 -485 0 3
rlabel polysilicon 285 -485 285 -485 0 4
rlabel polysilicon 289 -479 289 -479 0 1
rlabel polysilicon 289 -485 289 -485 0 3
rlabel polysilicon 296 -479 296 -479 0 1
rlabel polysilicon 296 -485 296 -485 0 3
rlabel polysilicon 303 -479 303 -479 0 1
rlabel polysilicon 303 -485 303 -485 0 3
rlabel polysilicon 310 -479 310 -479 0 1
rlabel polysilicon 310 -485 310 -485 0 3
rlabel polysilicon 317 -479 317 -479 0 1
rlabel polysilicon 317 -485 317 -485 0 3
rlabel polysilicon 324 -479 324 -479 0 1
rlabel polysilicon 327 -479 327 -479 0 2
rlabel polysilicon 324 -485 324 -485 0 3
rlabel polysilicon 327 -485 327 -485 0 4
rlabel polysilicon 331 -479 331 -479 0 1
rlabel polysilicon 331 -485 331 -485 0 3
rlabel polysilicon 338 -479 338 -479 0 1
rlabel polysilicon 338 -485 338 -485 0 3
rlabel polysilicon 345 -479 345 -479 0 1
rlabel polysilicon 348 -485 348 -485 0 4
rlabel polysilicon 352 -479 352 -479 0 1
rlabel polysilicon 352 -485 352 -485 0 3
rlabel polysilicon 355 -485 355 -485 0 4
rlabel polysilicon 359 -479 359 -479 0 1
rlabel polysilicon 359 -485 359 -485 0 3
rlabel polysilicon 366 -479 366 -479 0 1
rlabel polysilicon 366 -485 366 -485 0 3
rlabel polysilicon 373 -479 373 -479 0 1
rlabel polysilicon 373 -485 373 -485 0 3
rlabel polysilicon 380 -479 380 -479 0 1
rlabel polysilicon 383 -479 383 -479 0 2
rlabel polysilicon 383 -485 383 -485 0 4
rlabel polysilicon 387 -479 387 -479 0 1
rlabel polysilicon 387 -485 387 -485 0 3
rlabel polysilicon 397 -479 397 -479 0 2
rlabel polysilicon 397 -485 397 -485 0 4
rlabel polysilicon 401 -479 401 -479 0 1
rlabel polysilicon 401 -485 401 -485 0 3
rlabel polysilicon 408 -479 408 -479 0 1
rlabel polysilicon 408 -485 408 -485 0 3
rlabel polysilicon 415 -485 415 -485 0 3
rlabel polysilicon 418 -485 418 -485 0 4
rlabel polysilicon 422 -479 422 -479 0 1
rlabel polysilicon 425 -479 425 -479 0 2
rlabel polysilicon 422 -485 422 -485 0 3
rlabel polysilicon 425 -485 425 -485 0 4
rlabel polysilicon 429 -479 429 -479 0 1
rlabel polysilicon 429 -485 429 -485 0 3
rlabel polysilicon 436 -479 436 -479 0 1
rlabel polysilicon 436 -485 436 -485 0 3
rlabel polysilicon 443 -479 443 -479 0 1
rlabel polysilicon 443 -485 443 -485 0 3
rlabel polysilicon 450 -479 450 -479 0 1
rlabel polysilicon 450 -485 450 -485 0 3
rlabel polysilicon 457 -479 457 -479 0 1
rlabel polysilicon 460 -479 460 -479 0 2
rlabel polysilicon 457 -485 457 -485 0 3
rlabel polysilicon 460 -485 460 -485 0 4
rlabel polysilicon 464 -479 464 -479 0 1
rlabel polysilicon 464 -485 464 -485 0 3
rlabel polysilicon 474 -479 474 -479 0 2
rlabel polysilicon 471 -485 471 -485 0 3
rlabel polysilicon 481 -479 481 -479 0 2
rlabel polysilicon 481 -485 481 -485 0 4
rlabel polysilicon 485 -479 485 -479 0 1
rlabel polysilicon 485 -485 485 -485 0 3
rlabel polysilicon 492 -479 492 -479 0 1
rlabel polysilicon 492 -485 492 -485 0 3
rlabel polysilicon 499 -479 499 -479 0 1
rlabel polysilicon 502 -479 502 -479 0 2
rlabel polysilicon 502 -485 502 -485 0 4
rlabel polysilicon 506 -479 506 -479 0 1
rlabel polysilicon 506 -485 506 -485 0 3
rlabel polysilicon 513 -479 513 -479 0 1
rlabel polysilicon 513 -485 513 -485 0 3
rlabel polysilicon 520 -479 520 -479 0 1
rlabel polysilicon 520 -485 520 -485 0 3
rlabel polysilicon 527 -479 527 -479 0 1
rlabel polysilicon 527 -485 527 -485 0 3
rlabel polysilicon 534 -479 534 -479 0 1
rlabel polysilicon 534 -485 534 -485 0 3
rlabel polysilicon 537 -485 537 -485 0 4
rlabel polysilicon 541 -479 541 -479 0 1
rlabel polysilicon 541 -485 541 -485 0 3
rlabel polysilicon 548 -479 548 -479 0 1
rlabel polysilicon 548 -485 548 -485 0 3
rlabel polysilicon 555 -479 555 -479 0 1
rlabel polysilicon 558 -479 558 -479 0 2
rlabel polysilicon 555 -485 555 -485 0 3
rlabel polysilicon 562 -485 562 -485 0 3
rlabel polysilicon 565 -485 565 -485 0 4
rlabel polysilicon 569 -479 569 -479 0 1
rlabel polysilicon 572 -479 572 -479 0 2
rlabel polysilicon 569 -485 569 -485 0 3
rlabel polysilicon 572 -485 572 -485 0 4
rlabel polysilicon 576 -479 576 -479 0 1
rlabel polysilicon 579 -479 579 -479 0 2
rlabel polysilicon 583 -479 583 -479 0 1
rlabel polysilicon 583 -485 583 -485 0 3
rlabel polysilicon 590 -479 590 -479 0 1
rlabel polysilicon 590 -485 590 -485 0 3
rlabel polysilicon 597 -479 597 -479 0 1
rlabel polysilicon 597 -485 597 -485 0 3
rlabel polysilicon 604 -479 604 -479 0 1
rlabel polysilicon 604 -485 604 -485 0 3
rlabel polysilicon 611 -479 611 -479 0 1
rlabel polysilicon 611 -485 611 -485 0 3
rlabel polysilicon 618 -479 618 -479 0 1
rlabel polysilicon 618 -485 618 -485 0 3
rlabel polysilicon 625 -479 625 -479 0 1
rlabel polysilicon 625 -485 625 -485 0 3
rlabel polysilicon 635 -479 635 -479 0 2
rlabel polysilicon 632 -485 632 -485 0 3
rlabel polysilicon 635 -485 635 -485 0 4
rlabel polysilicon 642 -485 642 -485 0 4
rlabel polysilicon 646 -479 646 -479 0 1
rlabel polysilicon 646 -485 646 -485 0 3
rlabel polysilicon 653 -479 653 -479 0 1
rlabel polysilicon 653 -485 653 -485 0 3
rlabel polysilicon 660 -479 660 -479 0 1
rlabel polysilicon 660 -485 660 -485 0 3
rlabel polysilicon 667 -479 667 -479 0 1
rlabel polysilicon 667 -485 667 -485 0 3
rlabel polysilicon 674 -479 674 -479 0 1
rlabel polysilicon 674 -485 674 -485 0 3
rlabel polysilicon 681 -479 681 -479 0 1
rlabel polysilicon 681 -485 681 -485 0 3
rlabel polysilicon 688 -479 688 -479 0 1
rlabel polysilicon 688 -485 688 -485 0 3
rlabel polysilicon 695 -479 695 -479 0 1
rlabel polysilicon 695 -485 695 -485 0 3
rlabel polysilicon 702 -479 702 -479 0 1
rlabel polysilicon 702 -485 702 -485 0 3
rlabel polysilicon 709 -479 709 -479 0 1
rlabel polysilicon 709 -485 709 -485 0 3
rlabel polysilicon 716 -479 716 -479 0 1
rlabel polysilicon 716 -485 716 -485 0 3
rlabel polysilicon 723 -479 723 -479 0 1
rlabel polysilicon 723 -485 723 -485 0 3
rlabel polysilicon 730 -479 730 -479 0 1
rlabel polysilicon 730 -485 730 -485 0 3
rlabel polysilicon 737 -479 737 -479 0 1
rlabel polysilicon 737 -485 737 -485 0 3
rlabel polysilicon 744 -479 744 -479 0 1
rlabel polysilicon 744 -485 744 -485 0 3
rlabel polysilicon 751 -479 751 -479 0 1
rlabel polysilicon 751 -485 751 -485 0 3
rlabel polysilicon 758 -479 758 -479 0 1
rlabel polysilicon 758 -485 758 -485 0 3
rlabel polysilicon 765 -479 765 -479 0 1
rlabel polysilicon 765 -485 765 -485 0 3
rlabel polysilicon 772 -479 772 -479 0 1
rlabel polysilicon 772 -485 772 -485 0 3
rlabel polysilicon 779 -479 779 -479 0 1
rlabel polysilicon 779 -485 779 -485 0 3
rlabel polysilicon 786 -479 786 -479 0 1
rlabel polysilicon 786 -485 786 -485 0 3
rlabel polysilicon 793 -479 793 -479 0 1
rlabel polysilicon 793 -485 793 -485 0 3
rlabel polysilicon 800 -479 800 -479 0 1
rlabel polysilicon 800 -485 800 -485 0 3
rlabel polysilicon 807 -479 807 -479 0 1
rlabel polysilicon 807 -485 807 -485 0 3
rlabel polysilicon 814 -485 814 -485 0 3
rlabel polysilicon 817 -485 817 -485 0 4
rlabel polysilicon 821 -479 821 -479 0 1
rlabel polysilicon 821 -485 821 -485 0 3
rlabel polysilicon 828 -479 828 -479 0 1
rlabel polysilicon 828 -485 828 -485 0 3
rlabel polysilicon 835 -479 835 -479 0 1
rlabel polysilicon 835 -485 835 -485 0 3
rlabel polysilicon 842 -479 842 -479 0 1
rlabel polysilicon 842 -485 842 -485 0 3
rlabel polysilicon 849 -479 849 -479 0 1
rlabel polysilicon 849 -485 849 -485 0 3
rlabel polysilicon 856 -479 856 -479 0 1
rlabel polysilicon 856 -485 856 -485 0 3
rlabel polysilicon 863 -479 863 -479 0 1
rlabel polysilicon 863 -485 863 -485 0 3
rlabel polysilicon 870 -479 870 -479 0 1
rlabel polysilicon 870 -485 870 -485 0 3
rlabel polysilicon 877 -479 877 -479 0 1
rlabel polysilicon 877 -485 877 -485 0 3
rlabel polysilicon 884 -479 884 -479 0 1
rlabel polysilicon 884 -485 884 -485 0 3
rlabel polysilicon 891 -479 891 -479 0 1
rlabel polysilicon 891 -485 891 -485 0 3
rlabel polysilicon 898 -479 898 -479 0 1
rlabel polysilicon 898 -485 898 -485 0 3
rlabel polysilicon 905 -479 905 -479 0 1
rlabel polysilicon 905 -485 905 -485 0 3
rlabel polysilicon 912 -479 912 -479 0 1
rlabel polysilicon 912 -485 912 -485 0 3
rlabel polysilicon 919 -479 919 -479 0 1
rlabel polysilicon 919 -485 919 -485 0 3
rlabel polysilicon 926 -479 926 -479 0 1
rlabel polysilicon 926 -485 926 -485 0 3
rlabel polysilicon 933 -479 933 -479 0 1
rlabel polysilicon 933 -485 933 -485 0 3
rlabel polysilicon 940 -479 940 -479 0 1
rlabel polysilicon 940 -485 940 -485 0 3
rlabel polysilicon 947 -479 947 -479 0 1
rlabel polysilicon 947 -485 947 -485 0 3
rlabel polysilicon 954 -479 954 -479 0 1
rlabel polysilicon 954 -485 954 -485 0 3
rlabel polysilicon 961 -479 961 -479 0 1
rlabel polysilicon 961 -485 961 -485 0 3
rlabel polysilicon 968 -479 968 -479 0 1
rlabel polysilicon 968 -485 968 -485 0 3
rlabel polysilicon 975 -479 975 -479 0 1
rlabel polysilicon 975 -485 975 -485 0 3
rlabel polysilicon 982 -479 982 -479 0 1
rlabel polysilicon 982 -485 982 -485 0 3
rlabel polysilicon 989 -479 989 -479 0 1
rlabel polysilicon 989 -485 989 -485 0 3
rlabel polysilicon 996 -479 996 -479 0 1
rlabel polysilicon 996 -485 996 -485 0 3
rlabel polysilicon 1003 -479 1003 -479 0 1
rlabel polysilicon 1003 -485 1003 -485 0 3
rlabel polysilicon 1010 -479 1010 -479 0 1
rlabel polysilicon 1010 -485 1010 -485 0 3
rlabel polysilicon 1017 -479 1017 -479 0 1
rlabel polysilicon 1017 -485 1017 -485 0 3
rlabel polysilicon 1024 -479 1024 -479 0 1
rlabel polysilicon 1024 -485 1024 -485 0 3
rlabel polysilicon 1031 -479 1031 -479 0 1
rlabel polysilicon 1034 -479 1034 -479 0 2
rlabel polysilicon 1038 -479 1038 -479 0 1
rlabel polysilicon 1045 -479 1045 -479 0 1
rlabel polysilicon 1045 -485 1045 -485 0 3
rlabel polysilicon 1115 -479 1115 -479 0 1
rlabel polysilicon 1115 -485 1115 -485 0 3
rlabel polysilicon 2 -602 2 -602 0 3
rlabel polysilicon 5 -602 5 -602 0 4
rlabel polysilicon 9 -596 9 -596 0 1
rlabel polysilicon 9 -602 9 -602 0 3
rlabel polysilicon 16 -596 16 -596 0 1
rlabel polysilicon 16 -602 16 -602 0 3
rlabel polysilicon 26 -596 26 -596 0 2
rlabel polysilicon 26 -602 26 -602 0 4
rlabel polysilicon 30 -596 30 -596 0 1
rlabel polysilicon 30 -602 30 -602 0 3
rlabel polysilicon 37 -602 37 -602 0 3
rlabel polysilicon 40 -602 40 -602 0 4
rlabel polysilicon 44 -596 44 -596 0 1
rlabel polysilicon 44 -602 44 -602 0 3
rlabel polysilicon 51 -596 51 -596 0 1
rlabel polysilicon 51 -602 51 -602 0 3
rlabel polysilicon 58 -596 58 -596 0 1
rlabel polysilicon 58 -602 58 -602 0 3
rlabel polysilicon 65 -596 65 -596 0 1
rlabel polysilicon 65 -602 65 -602 0 3
rlabel polysilicon 72 -596 72 -596 0 1
rlabel polysilicon 72 -602 72 -602 0 3
rlabel polysilicon 79 -596 79 -596 0 1
rlabel polysilicon 79 -602 79 -602 0 3
rlabel polysilicon 86 -596 86 -596 0 1
rlabel polysilicon 86 -602 86 -602 0 3
rlabel polysilicon 93 -596 93 -596 0 1
rlabel polysilicon 96 -596 96 -596 0 2
rlabel polysilicon 93 -602 93 -602 0 3
rlabel polysilicon 100 -596 100 -596 0 1
rlabel polysilicon 100 -602 100 -602 0 3
rlabel polysilicon 103 -602 103 -602 0 4
rlabel polysilicon 107 -596 107 -596 0 1
rlabel polysilicon 107 -602 107 -602 0 3
rlabel polysilicon 114 -596 114 -596 0 1
rlabel polysilicon 114 -602 114 -602 0 3
rlabel polysilicon 121 -596 121 -596 0 1
rlabel polysilicon 121 -602 121 -602 0 3
rlabel polysilicon 128 -596 128 -596 0 1
rlabel polysilicon 128 -602 128 -602 0 3
rlabel polysilicon 135 -596 135 -596 0 1
rlabel polysilicon 138 -596 138 -596 0 2
rlabel polysilicon 135 -602 135 -602 0 3
rlabel polysilicon 138 -602 138 -602 0 4
rlabel polysilicon 142 -596 142 -596 0 1
rlabel polysilicon 142 -602 142 -602 0 3
rlabel polysilicon 149 -596 149 -596 0 1
rlabel polysilicon 149 -602 149 -602 0 3
rlabel polysilicon 156 -596 156 -596 0 1
rlabel polysilicon 156 -602 156 -602 0 3
rlabel polysilicon 163 -596 163 -596 0 1
rlabel polysilicon 166 -596 166 -596 0 2
rlabel polysilicon 163 -602 163 -602 0 3
rlabel polysilicon 170 -596 170 -596 0 1
rlabel polysilicon 170 -602 170 -602 0 3
rlabel polysilicon 180 -596 180 -596 0 2
rlabel polysilicon 177 -602 177 -602 0 3
rlabel polysilicon 184 -596 184 -596 0 1
rlabel polysilicon 184 -602 184 -602 0 3
rlabel polysilicon 191 -596 191 -596 0 1
rlabel polysilicon 191 -602 191 -602 0 3
rlabel polysilicon 198 -596 198 -596 0 1
rlabel polysilicon 198 -602 198 -602 0 3
rlabel polysilicon 205 -596 205 -596 0 1
rlabel polysilicon 208 -596 208 -596 0 2
rlabel polysilicon 205 -602 205 -602 0 3
rlabel polysilicon 212 -596 212 -596 0 1
rlabel polysilicon 215 -596 215 -596 0 2
rlabel polysilicon 212 -602 212 -602 0 3
rlabel polysilicon 215 -602 215 -602 0 4
rlabel polysilicon 219 -596 219 -596 0 1
rlabel polysilicon 219 -602 219 -602 0 3
rlabel polysilicon 222 -602 222 -602 0 4
rlabel polysilicon 226 -596 226 -596 0 1
rlabel polysilicon 226 -602 226 -602 0 3
rlabel polysilicon 233 -596 233 -596 0 1
rlabel polysilicon 233 -602 233 -602 0 3
rlabel polysilicon 240 -596 240 -596 0 1
rlabel polysilicon 240 -602 240 -602 0 3
rlabel polysilicon 247 -596 247 -596 0 1
rlabel polysilicon 247 -602 247 -602 0 3
rlabel polysilicon 254 -596 254 -596 0 1
rlabel polysilicon 254 -602 254 -602 0 3
rlabel polysilicon 261 -596 261 -596 0 1
rlabel polysilicon 261 -602 261 -602 0 3
rlabel polysilicon 268 -596 268 -596 0 1
rlabel polysilicon 271 -596 271 -596 0 2
rlabel polysilicon 268 -602 268 -602 0 3
rlabel polysilicon 275 -596 275 -596 0 1
rlabel polysilicon 275 -602 275 -602 0 3
rlabel polysilicon 282 -596 282 -596 0 1
rlabel polysilicon 282 -602 282 -602 0 3
rlabel polysilicon 289 -596 289 -596 0 1
rlabel polysilicon 289 -602 289 -602 0 3
rlabel polysilicon 296 -596 296 -596 0 1
rlabel polysilicon 296 -602 296 -602 0 3
rlabel polysilicon 303 -596 303 -596 0 1
rlabel polysilicon 303 -602 303 -602 0 3
rlabel polysilicon 310 -596 310 -596 0 1
rlabel polysilicon 310 -602 310 -602 0 3
rlabel polysilicon 317 -596 317 -596 0 1
rlabel polysilicon 317 -602 317 -602 0 3
rlabel polysilicon 324 -596 324 -596 0 1
rlabel polysilicon 324 -602 324 -602 0 3
rlabel polysilicon 331 -596 331 -596 0 1
rlabel polysilicon 331 -602 331 -602 0 3
rlabel polysilicon 341 -596 341 -596 0 2
rlabel polysilicon 338 -602 338 -602 0 3
rlabel polysilicon 341 -602 341 -602 0 4
rlabel polysilicon 345 -596 345 -596 0 1
rlabel polysilicon 348 -596 348 -596 0 2
rlabel polysilicon 345 -602 345 -602 0 3
rlabel polysilicon 348 -602 348 -602 0 4
rlabel polysilicon 352 -596 352 -596 0 1
rlabel polysilicon 352 -602 352 -602 0 3
rlabel polysilicon 359 -596 359 -596 0 1
rlabel polysilicon 359 -602 359 -602 0 3
rlabel polysilicon 366 -596 366 -596 0 1
rlabel polysilicon 366 -602 366 -602 0 3
rlabel polysilicon 373 -596 373 -596 0 1
rlabel polysilicon 373 -602 373 -602 0 3
rlabel polysilicon 380 -596 380 -596 0 1
rlabel polysilicon 380 -602 380 -602 0 3
rlabel polysilicon 387 -596 387 -596 0 1
rlabel polysilicon 387 -602 387 -602 0 3
rlabel polysilicon 394 -596 394 -596 0 1
rlabel polysilicon 394 -602 394 -602 0 3
rlabel polysilicon 401 -596 401 -596 0 1
rlabel polysilicon 401 -602 401 -602 0 3
rlabel polysilicon 408 -596 408 -596 0 1
rlabel polysilicon 408 -602 408 -602 0 3
rlabel polysilicon 415 -596 415 -596 0 1
rlabel polysilicon 415 -602 415 -602 0 3
rlabel polysilicon 422 -596 422 -596 0 1
rlabel polysilicon 422 -602 422 -602 0 3
rlabel polysilicon 429 -596 429 -596 0 1
rlabel polysilicon 429 -602 429 -602 0 3
rlabel polysilicon 436 -596 436 -596 0 1
rlabel polysilicon 439 -602 439 -602 0 4
rlabel polysilicon 443 -596 443 -596 0 1
rlabel polysilicon 443 -602 443 -602 0 3
rlabel polysilicon 450 -596 450 -596 0 1
rlabel polysilicon 450 -602 450 -602 0 3
rlabel polysilicon 457 -596 457 -596 0 1
rlabel polysilicon 457 -602 457 -602 0 3
rlabel polysilicon 464 -596 464 -596 0 1
rlabel polysilicon 467 -602 467 -602 0 4
rlabel polysilicon 471 -596 471 -596 0 1
rlabel polysilicon 474 -596 474 -596 0 2
rlabel polysilicon 471 -602 471 -602 0 3
rlabel polysilicon 474 -602 474 -602 0 4
rlabel polysilicon 478 -596 478 -596 0 1
rlabel polysilicon 478 -602 478 -602 0 3
rlabel polysilicon 485 -596 485 -596 0 1
rlabel polysilicon 485 -602 485 -602 0 3
rlabel polysilicon 492 -596 492 -596 0 1
rlabel polysilicon 492 -602 492 -602 0 3
rlabel polysilicon 499 -596 499 -596 0 1
rlabel polysilicon 499 -602 499 -602 0 3
rlabel polysilicon 506 -596 506 -596 0 1
rlabel polysilicon 506 -602 506 -602 0 3
rlabel polysilicon 513 -596 513 -596 0 1
rlabel polysilicon 513 -602 513 -602 0 3
rlabel polysilicon 523 -596 523 -596 0 2
rlabel polysilicon 520 -602 520 -602 0 3
rlabel polysilicon 523 -602 523 -602 0 4
rlabel polysilicon 527 -596 527 -596 0 1
rlabel polysilicon 530 -596 530 -596 0 2
rlabel polysilicon 534 -596 534 -596 0 1
rlabel polysilicon 537 -596 537 -596 0 2
rlabel polysilicon 534 -602 534 -602 0 3
rlabel polysilicon 541 -596 541 -596 0 1
rlabel polysilicon 541 -602 541 -602 0 3
rlabel polysilicon 548 -596 548 -596 0 1
rlabel polysilicon 551 -596 551 -596 0 2
rlabel polysilicon 548 -602 548 -602 0 3
rlabel polysilicon 551 -602 551 -602 0 4
rlabel polysilicon 555 -596 555 -596 0 1
rlabel polysilicon 555 -602 555 -602 0 3
rlabel polysilicon 562 -596 562 -596 0 1
rlabel polysilicon 565 -596 565 -596 0 2
rlabel polysilicon 562 -602 562 -602 0 3
rlabel polysilicon 572 -596 572 -596 0 2
rlabel polysilicon 569 -602 569 -602 0 3
rlabel polysilicon 572 -602 572 -602 0 4
rlabel polysilicon 576 -596 576 -596 0 1
rlabel polysilicon 579 -596 579 -596 0 2
rlabel polysilicon 576 -602 576 -602 0 3
rlabel polysilicon 579 -602 579 -602 0 4
rlabel polysilicon 583 -596 583 -596 0 1
rlabel polysilicon 583 -602 583 -602 0 3
rlabel polysilicon 590 -596 590 -596 0 1
rlabel polysilicon 590 -602 590 -602 0 3
rlabel polysilicon 597 -596 597 -596 0 1
rlabel polysilicon 600 -596 600 -596 0 2
rlabel polysilicon 597 -602 597 -602 0 3
rlabel polysilicon 604 -596 604 -596 0 1
rlabel polysilicon 604 -602 604 -602 0 3
rlabel polysilicon 611 -596 611 -596 0 1
rlabel polysilicon 611 -602 611 -602 0 3
rlabel polysilicon 618 -596 618 -596 0 1
rlabel polysilicon 618 -602 618 -602 0 3
rlabel polysilicon 625 -596 625 -596 0 1
rlabel polysilicon 625 -602 625 -602 0 3
rlabel polysilicon 632 -596 632 -596 0 1
rlabel polysilicon 632 -602 632 -602 0 3
rlabel polysilicon 639 -596 639 -596 0 1
rlabel polysilicon 639 -602 639 -602 0 3
rlabel polysilicon 646 -596 646 -596 0 1
rlabel polysilicon 646 -602 646 -602 0 3
rlabel polysilicon 653 -596 653 -596 0 1
rlabel polysilicon 653 -602 653 -602 0 3
rlabel polysilicon 660 -596 660 -596 0 1
rlabel polysilicon 660 -602 660 -602 0 3
rlabel polysilicon 667 -596 667 -596 0 1
rlabel polysilicon 667 -602 667 -602 0 3
rlabel polysilicon 674 -596 674 -596 0 1
rlabel polysilicon 674 -602 674 -602 0 3
rlabel polysilicon 681 -596 681 -596 0 1
rlabel polysilicon 684 -596 684 -596 0 2
rlabel polysilicon 684 -602 684 -602 0 4
rlabel polysilicon 688 -596 688 -596 0 1
rlabel polysilicon 688 -602 688 -602 0 3
rlabel polysilicon 695 -596 695 -596 0 1
rlabel polysilicon 695 -602 695 -602 0 3
rlabel polysilicon 702 -596 702 -596 0 1
rlabel polysilicon 702 -602 702 -602 0 3
rlabel polysilicon 709 -596 709 -596 0 1
rlabel polysilicon 712 -596 712 -596 0 2
rlabel polysilicon 712 -602 712 -602 0 4
rlabel polysilicon 716 -596 716 -596 0 1
rlabel polysilicon 716 -602 716 -602 0 3
rlabel polysilicon 723 -596 723 -596 0 1
rlabel polysilicon 723 -602 723 -602 0 3
rlabel polysilicon 733 -602 733 -602 0 4
rlabel polysilicon 737 -596 737 -596 0 1
rlabel polysilicon 737 -602 737 -602 0 3
rlabel polysilicon 744 -596 744 -596 0 1
rlabel polysilicon 744 -602 744 -602 0 3
rlabel polysilicon 751 -596 751 -596 0 1
rlabel polysilicon 751 -602 751 -602 0 3
rlabel polysilicon 758 -596 758 -596 0 1
rlabel polysilicon 758 -602 758 -602 0 3
rlabel polysilicon 765 -596 765 -596 0 1
rlabel polysilicon 765 -602 765 -602 0 3
rlabel polysilicon 772 -596 772 -596 0 1
rlabel polysilicon 772 -602 772 -602 0 3
rlabel polysilicon 779 -596 779 -596 0 1
rlabel polysilicon 779 -602 779 -602 0 3
rlabel polysilicon 786 -596 786 -596 0 1
rlabel polysilicon 786 -602 786 -602 0 3
rlabel polysilicon 793 -596 793 -596 0 1
rlabel polysilicon 793 -602 793 -602 0 3
rlabel polysilicon 800 -596 800 -596 0 1
rlabel polysilicon 800 -602 800 -602 0 3
rlabel polysilicon 807 -596 807 -596 0 1
rlabel polysilicon 807 -602 807 -602 0 3
rlabel polysilicon 814 -596 814 -596 0 1
rlabel polysilicon 814 -602 814 -602 0 3
rlabel polysilicon 821 -596 821 -596 0 1
rlabel polysilicon 821 -602 821 -602 0 3
rlabel polysilicon 828 -596 828 -596 0 1
rlabel polysilicon 828 -602 828 -602 0 3
rlabel polysilicon 835 -596 835 -596 0 1
rlabel polysilicon 835 -602 835 -602 0 3
rlabel polysilicon 842 -596 842 -596 0 1
rlabel polysilicon 842 -602 842 -602 0 3
rlabel polysilicon 849 -596 849 -596 0 1
rlabel polysilicon 849 -602 849 -602 0 3
rlabel polysilicon 856 -596 856 -596 0 1
rlabel polysilicon 856 -602 856 -602 0 3
rlabel polysilicon 863 -596 863 -596 0 1
rlabel polysilicon 863 -602 863 -602 0 3
rlabel polysilicon 870 -596 870 -596 0 1
rlabel polysilicon 870 -602 870 -602 0 3
rlabel polysilicon 877 -596 877 -596 0 1
rlabel polysilicon 877 -602 877 -602 0 3
rlabel polysilicon 884 -596 884 -596 0 1
rlabel polysilicon 884 -602 884 -602 0 3
rlabel polysilicon 891 -596 891 -596 0 1
rlabel polysilicon 891 -602 891 -602 0 3
rlabel polysilicon 898 -596 898 -596 0 1
rlabel polysilicon 898 -602 898 -602 0 3
rlabel polysilicon 905 -596 905 -596 0 1
rlabel polysilicon 905 -602 905 -602 0 3
rlabel polysilicon 912 -596 912 -596 0 1
rlabel polysilicon 912 -602 912 -602 0 3
rlabel polysilicon 919 -596 919 -596 0 1
rlabel polysilicon 919 -602 919 -602 0 3
rlabel polysilicon 926 -596 926 -596 0 1
rlabel polysilicon 926 -602 926 -602 0 3
rlabel polysilicon 933 -596 933 -596 0 1
rlabel polysilicon 933 -602 933 -602 0 3
rlabel polysilicon 940 -596 940 -596 0 1
rlabel polysilicon 940 -602 940 -602 0 3
rlabel polysilicon 947 -596 947 -596 0 1
rlabel polysilicon 947 -602 947 -602 0 3
rlabel polysilicon 954 -596 954 -596 0 1
rlabel polysilicon 954 -602 954 -602 0 3
rlabel polysilicon 961 -596 961 -596 0 1
rlabel polysilicon 961 -602 961 -602 0 3
rlabel polysilicon 968 -596 968 -596 0 1
rlabel polysilicon 968 -602 968 -602 0 3
rlabel polysilicon 975 -596 975 -596 0 1
rlabel polysilicon 975 -602 975 -602 0 3
rlabel polysilicon 982 -596 982 -596 0 1
rlabel polysilicon 982 -602 982 -602 0 3
rlabel polysilicon 989 -596 989 -596 0 1
rlabel polysilicon 989 -602 989 -602 0 3
rlabel polysilicon 996 -596 996 -596 0 1
rlabel polysilicon 996 -602 996 -602 0 3
rlabel polysilicon 1003 -596 1003 -596 0 1
rlabel polysilicon 1003 -602 1003 -602 0 3
rlabel polysilicon 1010 -596 1010 -596 0 1
rlabel polysilicon 1010 -602 1010 -602 0 3
rlabel polysilicon 1017 -596 1017 -596 0 1
rlabel polysilicon 1017 -602 1017 -602 0 3
rlabel polysilicon 1024 -596 1024 -596 0 1
rlabel polysilicon 1024 -602 1024 -602 0 3
rlabel polysilicon 1031 -596 1031 -596 0 1
rlabel polysilicon 1031 -602 1031 -602 0 3
rlabel polysilicon 1038 -596 1038 -596 0 1
rlabel polysilicon 1038 -602 1038 -602 0 3
rlabel polysilicon 1045 -596 1045 -596 0 1
rlabel polysilicon 1045 -602 1045 -602 0 3
rlabel polysilicon 1052 -596 1052 -596 0 1
rlabel polysilicon 1052 -602 1052 -602 0 3
rlabel polysilicon 1059 -596 1059 -596 0 1
rlabel polysilicon 1059 -602 1059 -602 0 3
rlabel polysilicon 1066 -596 1066 -596 0 1
rlabel polysilicon 1066 -602 1066 -602 0 3
rlabel polysilicon 1073 -596 1073 -596 0 1
rlabel polysilicon 1073 -602 1073 -602 0 3
rlabel polysilicon 1080 -596 1080 -596 0 1
rlabel polysilicon 1080 -602 1080 -602 0 3
rlabel polysilicon 1087 -596 1087 -596 0 1
rlabel polysilicon 1087 -602 1087 -602 0 3
rlabel polysilicon 1094 -596 1094 -596 0 1
rlabel polysilicon 1094 -602 1094 -602 0 3
rlabel polysilicon 1101 -602 1101 -602 0 3
rlabel polysilicon 1111 -596 1111 -596 0 2
rlabel polysilicon 1108 -602 1108 -602 0 3
rlabel polysilicon 1115 -596 1115 -596 0 1
rlabel polysilicon 1115 -602 1115 -602 0 3
rlabel polysilicon 1122 -596 1122 -596 0 1
rlabel polysilicon 1122 -602 1122 -602 0 3
rlabel polysilicon 1129 -596 1129 -596 0 1
rlabel polysilicon 1129 -602 1129 -602 0 3
rlabel polysilicon 2 -697 2 -697 0 1
rlabel polysilicon 2 -703 2 -703 0 3
rlabel polysilicon 9 -703 9 -703 0 3
rlabel polysilicon 16 -697 16 -697 0 1
rlabel polysilicon 16 -703 16 -703 0 3
rlabel polysilicon 23 -697 23 -697 0 1
rlabel polysilicon 23 -703 23 -703 0 3
rlabel polysilicon 30 -697 30 -697 0 1
rlabel polysilicon 30 -703 30 -703 0 3
rlabel polysilicon 37 -697 37 -697 0 1
rlabel polysilicon 37 -703 37 -703 0 3
rlabel polysilicon 44 -697 44 -697 0 1
rlabel polysilicon 47 -697 47 -697 0 2
rlabel polysilicon 51 -697 51 -697 0 1
rlabel polysilicon 51 -703 51 -703 0 3
rlabel polysilicon 58 -697 58 -697 0 1
rlabel polysilicon 58 -703 58 -703 0 3
rlabel polysilicon 65 -697 65 -697 0 1
rlabel polysilicon 65 -703 65 -703 0 3
rlabel polysilicon 72 -697 72 -697 0 1
rlabel polysilicon 72 -703 72 -703 0 3
rlabel polysilicon 82 -697 82 -697 0 2
rlabel polysilicon 79 -703 79 -703 0 3
rlabel polysilicon 82 -703 82 -703 0 4
rlabel polysilicon 86 -697 86 -697 0 1
rlabel polysilicon 86 -703 86 -703 0 3
rlabel polysilicon 93 -697 93 -697 0 1
rlabel polysilicon 93 -703 93 -703 0 3
rlabel polysilicon 100 -697 100 -697 0 1
rlabel polysilicon 100 -703 100 -703 0 3
rlabel polysilicon 107 -697 107 -697 0 1
rlabel polysilicon 107 -703 107 -703 0 3
rlabel polysilicon 117 -697 117 -697 0 2
rlabel polysilicon 114 -703 114 -703 0 3
rlabel polysilicon 124 -697 124 -697 0 2
rlabel polysilicon 121 -703 121 -703 0 3
rlabel polysilicon 124 -703 124 -703 0 4
rlabel polysilicon 128 -697 128 -697 0 1
rlabel polysilicon 131 -697 131 -697 0 2
rlabel polysilicon 131 -703 131 -703 0 4
rlabel polysilicon 135 -697 135 -697 0 1
rlabel polysilicon 135 -703 135 -703 0 3
rlabel polysilicon 142 -697 142 -697 0 1
rlabel polysilicon 142 -703 142 -703 0 3
rlabel polysilicon 149 -697 149 -697 0 1
rlabel polysilicon 149 -703 149 -703 0 3
rlabel polysilicon 156 -697 156 -697 0 1
rlabel polysilicon 156 -703 156 -703 0 3
rlabel polysilicon 163 -697 163 -697 0 1
rlabel polysilicon 163 -703 163 -703 0 3
rlabel polysilicon 173 -697 173 -697 0 2
rlabel polysilicon 170 -703 170 -703 0 3
rlabel polysilicon 177 -697 177 -697 0 1
rlabel polysilicon 177 -703 177 -703 0 3
rlabel polysilicon 184 -697 184 -697 0 1
rlabel polysilicon 184 -703 184 -703 0 3
rlabel polysilicon 191 -697 191 -697 0 1
rlabel polysilicon 191 -703 191 -703 0 3
rlabel polysilicon 201 -697 201 -697 0 2
rlabel polysilicon 198 -703 198 -703 0 3
rlabel polysilicon 205 -697 205 -697 0 1
rlabel polysilicon 205 -703 205 -703 0 3
rlabel polysilicon 208 -703 208 -703 0 4
rlabel polysilicon 212 -697 212 -697 0 1
rlabel polysilicon 212 -703 212 -703 0 3
rlabel polysilicon 219 -697 219 -697 0 1
rlabel polysilicon 219 -703 219 -703 0 3
rlabel polysilicon 226 -703 226 -703 0 3
rlabel polysilicon 233 -697 233 -697 0 1
rlabel polysilicon 233 -703 233 -703 0 3
rlabel polysilicon 240 -697 240 -697 0 1
rlabel polysilicon 240 -703 240 -703 0 3
rlabel polysilicon 247 -697 247 -697 0 1
rlabel polysilicon 247 -703 247 -703 0 3
rlabel polysilicon 254 -697 254 -697 0 1
rlabel polysilicon 254 -703 254 -703 0 3
rlabel polysilicon 261 -697 261 -697 0 1
rlabel polysilicon 261 -703 261 -703 0 3
rlabel polysilicon 268 -697 268 -697 0 1
rlabel polysilicon 268 -703 268 -703 0 3
rlabel polysilicon 275 -697 275 -697 0 1
rlabel polysilicon 275 -703 275 -703 0 3
rlabel polysilicon 282 -697 282 -697 0 1
rlabel polysilicon 282 -703 282 -703 0 3
rlabel polysilicon 292 -697 292 -697 0 2
rlabel polysilicon 289 -703 289 -703 0 3
rlabel polysilicon 292 -703 292 -703 0 4
rlabel polysilicon 296 -697 296 -697 0 1
rlabel polysilicon 296 -703 296 -703 0 3
rlabel polysilicon 303 -697 303 -697 0 1
rlabel polysilicon 303 -703 303 -703 0 3
rlabel polysilicon 313 -697 313 -697 0 2
rlabel polysilicon 310 -703 310 -703 0 3
rlabel polysilicon 317 -697 317 -697 0 1
rlabel polysilicon 317 -703 317 -703 0 3
rlabel polysilicon 324 -697 324 -697 0 1
rlabel polysilicon 324 -703 324 -703 0 3
rlabel polysilicon 331 -697 331 -697 0 1
rlabel polysilicon 331 -703 331 -703 0 3
rlabel polysilicon 338 -697 338 -697 0 1
rlabel polysilicon 338 -703 338 -703 0 3
rlabel polysilicon 345 -697 345 -697 0 1
rlabel polysilicon 345 -703 345 -703 0 3
rlabel polysilicon 352 -697 352 -697 0 1
rlabel polysilicon 352 -703 352 -703 0 3
rlabel polysilicon 359 -697 359 -697 0 1
rlabel polysilicon 362 -697 362 -697 0 2
rlabel polysilicon 359 -703 359 -703 0 3
rlabel polysilicon 362 -703 362 -703 0 4
rlabel polysilicon 366 -697 366 -697 0 1
rlabel polysilicon 366 -703 366 -703 0 3
rlabel polysilicon 373 -697 373 -697 0 1
rlabel polysilicon 373 -703 373 -703 0 3
rlabel polysilicon 380 -697 380 -697 0 1
rlabel polysilicon 380 -703 380 -703 0 3
rlabel polysilicon 387 -697 387 -697 0 1
rlabel polysilicon 387 -703 387 -703 0 3
rlabel polysilicon 394 -697 394 -697 0 1
rlabel polysilicon 394 -703 394 -703 0 3
rlabel polysilicon 401 -697 401 -697 0 1
rlabel polysilicon 401 -703 401 -703 0 3
rlabel polysilicon 408 -697 408 -697 0 1
rlabel polysilicon 408 -703 408 -703 0 3
rlabel polysilicon 415 -697 415 -697 0 1
rlabel polysilicon 415 -703 415 -703 0 3
rlabel polysilicon 422 -697 422 -697 0 1
rlabel polysilicon 422 -703 422 -703 0 3
rlabel polysilicon 429 -697 429 -697 0 1
rlabel polysilicon 429 -703 429 -703 0 3
rlabel polysilicon 436 -697 436 -697 0 1
rlabel polysilicon 436 -703 436 -703 0 3
rlabel polysilicon 443 -697 443 -697 0 1
rlabel polysilicon 443 -703 443 -703 0 3
rlabel polysilicon 446 -703 446 -703 0 4
rlabel polysilicon 450 -697 450 -697 0 1
rlabel polysilicon 453 -697 453 -697 0 2
rlabel polysilicon 453 -703 453 -703 0 4
rlabel polysilicon 457 -697 457 -697 0 1
rlabel polysilicon 460 -697 460 -697 0 2
rlabel polysilicon 457 -703 457 -703 0 3
rlabel polysilicon 460 -703 460 -703 0 4
rlabel polysilicon 467 -697 467 -697 0 2
rlabel polysilicon 464 -703 464 -703 0 3
rlabel polysilicon 467 -703 467 -703 0 4
rlabel polysilicon 471 -697 471 -697 0 1
rlabel polysilicon 471 -703 471 -703 0 3
rlabel polysilicon 478 -697 478 -697 0 1
rlabel polysilicon 481 -697 481 -697 0 2
rlabel polysilicon 478 -703 478 -703 0 3
rlabel polysilicon 485 -697 485 -697 0 1
rlabel polysilicon 485 -703 485 -703 0 3
rlabel polysilicon 492 -697 492 -697 0 1
rlabel polysilicon 495 -697 495 -697 0 2
rlabel polysilicon 495 -703 495 -703 0 4
rlabel polysilicon 499 -697 499 -697 0 1
rlabel polysilicon 499 -703 499 -703 0 3
rlabel polysilicon 506 -697 506 -697 0 1
rlabel polysilicon 506 -703 506 -703 0 3
rlabel polysilicon 513 -697 513 -697 0 1
rlabel polysilicon 516 -697 516 -697 0 2
rlabel polysilicon 513 -703 513 -703 0 3
rlabel polysilicon 516 -703 516 -703 0 4
rlabel polysilicon 520 -697 520 -697 0 1
rlabel polysilicon 520 -703 520 -703 0 3
rlabel polysilicon 527 -697 527 -697 0 1
rlabel polysilicon 527 -703 527 -703 0 3
rlabel polysilicon 534 -697 534 -697 0 1
rlabel polysilicon 534 -703 534 -703 0 3
rlabel polysilicon 541 -697 541 -697 0 1
rlabel polysilicon 544 -697 544 -697 0 2
rlabel polysilicon 544 -703 544 -703 0 4
rlabel polysilicon 548 -697 548 -697 0 1
rlabel polysilicon 548 -703 548 -703 0 3
rlabel polysilicon 555 -697 555 -697 0 1
rlabel polysilicon 555 -703 555 -703 0 3
rlabel polysilicon 562 -697 562 -697 0 1
rlabel polysilicon 565 -697 565 -697 0 2
rlabel polysilicon 562 -703 562 -703 0 3
rlabel polysilicon 569 -697 569 -697 0 1
rlabel polysilicon 569 -703 569 -703 0 3
rlabel polysilicon 576 -697 576 -697 0 1
rlabel polysilicon 576 -703 576 -703 0 3
rlabel polysilicon 583 -697 583 -697 0 1
rlabel polysilicon 583 -703 583 -703 0 3
rlabel polysilicon 590 -697 590 -697 0 1
rlabel polysilicon 590 -703 590 -703 0 3
rlabel polysilicon 597 -697 597 -697 0 1
rlabel polysilicon 597 -703 597 -703 0 3
rlabel polysilicon 604 -697 604 -697 0 1
rlabel polysilicon 607 -697 607 -697 0 2
rlabel polysilicon 611 -697 611 -697 0 1
rlabel polysilicon 611 -703 611 -703 0 3
rlabel polysilicon 618 -697 618 -697 0 1
rlabel polysilicon 618 -703 618 -703 0 3
rlabel polysilicon 625 -697 625 -697 0 1
rlabel polysilicon 625 -703 625 -703 0 3
rlabel polysilicon 632 -697 632 -697 0 1
rlabel polysilicon 632 -703 632 -703 0 3
rlabel polysilicon 639 -697 639 -697 0 1
rlabel polysilicon 639 -703 639 -703 0 3
rlabel polysilicon 646 -697 646 -697 0 1
rlabel polysilicon 646 -703 646 -703 0 3
rlabel polysilicon 653 -697 653 -697 0 1
rlabel polysilicon 653 -703 653 -703 0 3
rlabel polysilicon 660 -697 660 -697 0 1
rlabel polysilicon 660 -703 660 -703 0 3
rlabel polysilicon 667 -697 667 -697 0 1
rlabel polysilicon 674 -697 674 -697 0 1
rlabel polysilicon 674 -703 674 -703 0 3
rlabel polysilicon 681 -697 681 -697 0 1
rlabel polysilicon 681 -703 681 -703 0 3
rlabel polysilicon 688 -697 688 -697 0 1
rlabel polysilicon 688 -703 688 -703 0 3
rlabel polysilicon 695 -697 695 -697 0 1
rlabel polysilicon 695 -703 695 -703 0 3
rlabel polysilicon 702 -697 702 -697 0 1
rlabel polysilicon 702 -703 702 -703 0 3
rlabel polysilicon 709 -697 709 -697 0 1
rlabel polysilicon 709 -703 709 -703 0 3
rlabel polysilicon 716 -697 716 -697 0 1
rlabel polysilicon 716 -703 716 -703 0 3
rlabel polysilicon 723 -697 723 -697 0 1
rlabel polysilicon 726 -697 726 -697 0 2
rlabel polysilicon 723 -703 723 -703 0 3
rlabel polysilicon 726 -703 726 -703 0 4
rlabel polysilicon 730 -697 730 -697 0 1
rlabel polysilicon 730 -703 730 -703 0 3
rlabel polysilicon 737 -697 737 -697 0 1
rlabel polysilicon 737 -703 737 -703 0 3
rlabel polysilicon 747 -703 747 -703 0 4
rlabel polysilicon 751 -697 751 -697 0 1
rlabel polysilicon 751 -703 751 -703 0 3
rlabel polysilicon 758 -697 758 -697 0 1
rlabel polysilicon 758 -703 758 -703 0 3
rlabel polysilicon 765 -697 765 -697 0 1
rlabel polysilicon 765 -703 765 -703 0 3
rlabel polysilicon 775 -697 775 -697 0 2
rlabel polysilicon 772 -703 772 -703 0 3
rlabel polysilicon 775 -703 775 -703 0 4
rlabel polysilicon 779 -697 779 -697 0 1
rlabel polysilicon 779 -703 779 -703 0 3
rlabel polysilicon 786 -697 786 -697 0 1
rlabel polysilicon 789 -697 789 -697 0 2
rlabel polysilicon 786 -703 786 -703 0 3
rlabel polysilicon 793 -697 793 -697 0 1
rlabel polysilicon 793 -703 793 -703 0 3
rlabel polysilicon 800 -697 800 -697 0 1
rlabel polysilicon 800 -703 800 -703 0 3
rlabel polysilicon 807 -697 807 -697 0 1
rlabel polysilicon 807 -703 807 -703 0 3
rlabel polysilicon 814 -697 814 -697 0 1
rlabel polysilicon 814 -703 814 -703 0 3
rlabel polysilicon 821 -697 821 -697 0 1
rlabel polysilicon 821 -703 821 -703 0 3
rlabel polysilicon 828 -697 828 -697 0 1
rlabel polysilicon 828 -703 828 -703 0 3
rlabel polysilicon 835 -697 835 -697 0 1
rlabel polysilicon 835 -703 835 -703 0 3
rlabel polysilicon 842 -697 842 -697 0 1
rlabel polysilicon 842 -703 842 -703 0 3
rlabel polysilicon 849 -697 849 -697 0 1
rlabel polysilicon 849 -703 849 -703 0 3
rlabel polysilicon 856 -697 856 -697 0 1
rlabel polysilicon 856 -703 856 -703 0 3
rlabel polysilicon 863 -697 863 -697 0 1
rlabel polysilicon 863 -703 863 -703 0 3
rlabel polysilicon 870 -697 870 -697 0 1
rlabel polysilicon 870 -703 870 -703 0 3
rlabel polysilicon 877 -697 877 -697 0 1
rlabel polysilicon 877 -703 877 -703 0 3
rlabel polysilicon 884 -697 884 -697 0 1
rlabel polysilicon 884 -703 884 -703 0 3
rlabel polysilicon 891 -697 891 -697 0 1
rlabel polysilicon 891 -703 891 -703 0 3
rlabel polysilicon 898 -697 898 -697 0 1
rlabel polysilicon 898 -703 898 -703 0 3
rlabel polysilicon 905 -697 905 -697 0 1
rlabel polysilicon 905 -703 905 -703 0 3
rlabel polysilicon 912 -697 912 -697 0 1
rlabel polysilicon 912 -703 912 -703 0 3
rlabel polysilicon 919 -697 919 -697 0 1
rlabel polysilicon 919 -703 919 -703 0 3
rlabel polysilicon 926 -697 926 -697 0 1
rlabel polysilicon 926 -703 926 -703 0 3
rlabel polysilicon 933 -697 933 -697 0 1
rlabel polysilicon 933 -703 933 -703 0 3
rlabel polysilicon 940 -697 940 -697 0 1
rlabel polysilicon 940 -703 940 -703 0 3
rlabel polysilicon 947 -697 947 -697 0 1
rlabel polysilicon 947 -703 947 -703 0 3
rlabel polysilicon 954 -697 954 -697 0 1
rlabel polysilicon 954 -703 954 -703 0 3
rlabel polysilicon 961 -697 961 -697 0 1
rlabel polysilicon 961 -703 961 -703 0 3
rlabel polysilicon 968 -697 968 -697 0 1
rlabel polysilicon 968 -703 968 -703 0 3
rlabel polysilicon 975 -697 975 -697 0 1
rlabel polysilicon 975 -703 975 -703 0 3
rlabel polysilicon 982 -697 982 -697 0 1
rlabel polysilicon 982 -703 982 -703 0 3
rlabel polysilicon 989 -697 989 -697 0 1
rlabel polysilicon 989 -703 989 -703 0 3
rlabel polysilicon 996 -697 996 -697 0 1
rlabel polysilicon 996 -703 996 -703 0 3
rlabel polysilicon 1003 -697 1003 -697 0 1
rlabel polysilicon 1003 -703 1003 -703 0 3
rlabel polysilicon 1010 -697 1010 -697 0 1
rlabel polysilicon 1010 -703 1010 -703 0 3
rlabel polysilicon 1017 -697 1017 -697 0 1
rlabel polysilicon 1017 -703 1017 -703 0 3
rlabel polysilicon 1024 -697 1024 -697 0 1
rlabel polysilicon 1024 -703 1024 -703 0 3
rlabel polysilicon 1031 -697 1031 -697 0 1
rlabel polysilicon 1031 -703 1031 -703 0 3
rlabel polysilicon 1038 -697 1038 -697 0 1
rlabel polysilicon 1038 -703 1038 -703 0 3
rlabel polysilicon 1045 -697 1045 -697 0 1
rlabel polysilicon 1045 -703 1045 -703 0 3
rlabel polysilicon 1052 -697 1052 -697 0 1
rlabel polysilicon 1052 -703 1052 -703 0 3
rlabel polysilicon 1059 -697 1059 -697 0 1
rlabel polysilicon 1059 -703 1059 -703 0 3
rlabel polysilicon 1066 -697 1066 -697 0 1
rlabel polysilicon 1066 -703 1066 -703 0 3
rlabel polysilicon 1073 -697 1073 -697 0 1
rlabel polysilicon 1073 -703 1073 -703 0 3
rlabel polysilicon 1080 -697 1080 -697 0 1
rlabel polysilicon 1080 -703 1080 -703 0 3
rlabel polysilicon 1083 -703 1083 -703 0 4
rlabel polysilicon 1087 -697 1087 -697 0 1
rlabel polysilicon 1087 -703 1087 -703 0 3
rlabel polysilicon 1094 -697 1094 -697 0 1
rlabel polysilicon 1094 -703 1094 -703 0 3
rlabel polysilicon 1101 -697 1101 -697 0 1
rlabel polysilicon 1101 -703 1101 -703 0 3
rlabel polysilicon 1111 -697 1111 -697 0 2
rlabel polysilicon 1111 -703 1111 -703 0 4
rlabel polysilicon 1115 -697 1115 -697 0 1
rlabel polysilicon 1115 -703 1115 -703 0 3
rlabel polysilicon 1122 -697 1122 -697 0 1
rlabel polysilicon 1122 -703 1122 -703 0 3
rlabel polysilicon 1129 -697 1129 -697 0 1
rlabel polysilicon 1129 -703 1129 -703 0 3
rlabel polysilicon 1139 -697 1139 -697 0 2
rlabel polysilicon 1143 -697 1143 -697 0 1
rlabel polysilicon 1143 -703 1143 -703 0 3
rlabel polysilicon 1150 -697 1150 -697 0 1
rlabel polysilicon 1150 -703 1150 -703 0 3
rlabel polysilicon 1157 -697 1157 -697 0 1
rlabel polysilicon 1157 -703 1157 -703 0 3
rlabel polysilicon 23 -774 23 -774 0 1
rlabel polysilicon 23 -780 23 -780 0 3
rlabel polysilicon 30 -774 30 -774 0 1
rlabel polysilicon 37 -774 37 -774 0 1
rlabel polysilicon 37 -780 37 -780 0 3
rlabel polysilicon 44 -774 44 -774 0 1
rlabel polysilicon 44 -780 44 -780 0 3
rlabel polysilicon 51 -774 51 -774 0 1
rlabel polysilicon 51 -780 51 -780 0 3
rlabel polysilicon 58 -774 58 -774 0 1
rlabel polysilicon 58 -780 58 -780 0 3
rlabel polysilicon 65 -774 65 -774 0 1
rlabel polysilicon 65 -780 65 -780 0 3
rlabel polysilicon 72 -774 72 -774 0 1
rlabel polysilicon 72 -780 72 -780 0 3
rlabel polysilicon 79 -774 79 -774 0 1
rlabel polysilicon 79 -780 79 -780 0 3
rlabel polysilicon 86 -774 86 -774 0 1
rlabel polysilicon 89 -774 89 -774 0 2
rlabel polysilicon 86 -780 86 -780 0 3
rlabel polysilicon 93 -774 93 -774 0 1
rlabel polysilicon 93 -780 93 -780 0 3
rlabel polysilicon 100 -774 100 -774 0 1
rlabel polysilicon 103 -774 103 -774 0 2
rlabel polysilicon 103 -780 103 -780 0 4
rlabel polysilicon 107 -774 107 -774 0 1
rlabel polysilicon 107 -780 107 -780 0 3
rlabel polysilicon 114 -774 114 -774 0 1
rlabel polysilicon 114 -780 114 -780 0 3
rlabel polysilicon 121 -774 121 -774 0 1
rlabel polysilicon 121 -780 121 -780 0 3
rlabel polysilicon 128 -774 128 -774 0 1
rlabel polysilicon 128 -780 128 -780 0 3
rlabel polysilicon 135 -774 135 -774 0 1
rlabel polysilicon 135 -780 135 -780 0 3
rlabel polysilicon 138 -780 138 -780 0 4
rlabel polysilicon 142 -774 142 -774 0 1
rlabel polysilicon 142 -780 142 -780 0 3
rlabel polysilicon 149 -774 149 -774 0 1
rlabel polysilicon 152 -774 152 -774 0 2
rlabel polysilicon 152 -780 152 -780 0 4
rlabel polysilicon 156 -774 156 -774 0 1
rlabel polysilicon 159 -774 159 -774 0 2
rlabel polysilicon 156 -780 156 -780 0 3
rlabel polysilicon 163 -774 163 -774 0 1
rlabel polysilicon 163 -780 163 -780 0 3
rlabel polysilicon 170 -774 170 -774 0 1
rlabel polysilicon 173 -774 173 -774 0 2
rlabel polysilicon 173 -780 173 -780 0 4
rlabel polysilicon 177 -774 177 -774 0 1
rlabel polysilicon 177 -780 177 -780 0 3
rlabel polysilicon 184 -774 184 -774 0 1
rlabel polysilicon 184 -780 184 -780 0 3
rlabel polysilicon 191 -774 191 -774 0 1
rlabel polysilicon 191 -780 191 -780 0 3
rlabel polysilicon 198 -774 198 -774 0 1
rlabel polysilicon 198 -780 198 -780 0 3
rlabel polysilicon 208 -774 208 -774 0 2
rlabel polysilicon 208 -780 208 -780 0 4
rlabel polysilicon 212 -774 212 -774 0 1
rlabel polysilicon 212 -780 212 -780 0 3
rlabel polysilicon 219 -774 219 -774 0 1
rlabel polysilicon 219 -780 219 -780 0 3
rlabel polysilicon 226 -774 226 -774 0 1
rlabel polysilicon 226 -780 226 -780 0 3
rlabel polysilicon 233 -774 233 -774 0 1
rlabel polysilicon 233 -780 233 -780 0 3
rlabel polysilicon 240 -774 240 -774 0 1
rlabel polysilicon 240 -780 240 -780 0 3
rlabel polysilicon 247 -774 247 -774 0 1
rlabel polysilicon 247 -780 247 -780 0 3
rlabel polysilicon 254 -774 254 -774 0 1
rlabel polysilicon 254 -780 254 -780 0 3
rlabel polysilicon 261 -774 261 -774 0 1
rlabel polysilicon 261 -780 261 -780 0 3
rlabel polysilicon 268 -774 268 -774 0 1
rlabel polysilicon 268 -780 268 -780 0 3
rlabel polysilicon 275 -774 275 -774 0 1
rlabel polysilicon 275 -780 275 -780 0 3
rlabel polysilicon 282 -774 282 -774 0 1
rlabel polysilicon 282 -780 282 -780 0 3
rlabel polysilicon 289 -774 289 -774 0 1
rlabel polysilicon 292 -774 292 -774 0 2
rlabel polysilicon 292 -780 292 -780 0 4
rlabel polysilicon 296 -774 296 -774 0 1
rlabel polysilicon 296 -780 296 -780 0 3
rlabel polysilicon 303 -774 303 -774 0 1
rlabel polysilicon 303 -780 303 -780 0 3
rlabel polysilicon 310 -774 310 -774 0 1
rlabel polysilicon 313 -780 313 -780 0 4
rlabel polysilicon 317 -774 317 -774 0 1
rlabel polysilicon 317 -780 317 -780 0 3
rlabel polysilicon 324 -774 324 -774 0 1
rlabel polysilicon 327 -774 327 -774 0 2
rlabel polysilicon 324 -780 324 -780 0 3
rlabel polysilicon 331 -774 331 -774 0 1
rlabel polysilicon 331 -780 331 -780 0 3
rlabel polysilicon 338 -774 338 -774 0 1
rlabel polysilicon 338 -780 338 -780 0 3
rlabel polysilicon 345 -774 345 -774 0 1
rlabel polysilicon 345 -780 345 -780 0 3
rlabel polysilicon 352 -774 352 -774 0 1
rlabel polysilicon 352 -780 352 -780 0 3
rlabel polysilicon 359 -774 359 -774 0 1
rlabel polysilicon 359 -780 359 -780 0 3
rlabel polysilicon 369 -774 369 -774 0 2
rlabel polysilicon 366 -780 366 -780 0 3
rlabel polysilicon 369 -780 369 -780 0 4
rlabel polysilicon 373 -774 373 -774 0 1
rlabel polysilicon 373 -780 373 -780 0 3
rlabel polysilicon 380 -774 380 -774 0 1
rlabel polysilicon 380 -780 380 -780 0 3
rlabel polysilicon 387 -774 387 -774 0 1
rlabel polysilicon 387 -780 387 -780 0 3
rlabel polysilicon 394 -774 394 -774 0 1
rlabel polysilicon 394 -780 394 -780 0 3
rlabel polysilicon 401 -774 401 -774 0 1
rlabel polysilicon 401 -780 401 -780 0 3
rlabel polysilicon 408 -774 408 -774 0 1
rlabel polysilicon 408 -780 408 -780 0 3
rlabel polysilicon 415 -774 415 -774 0 1
rlabel polysilicon 415 -780 415 -780 0 3
rlabel polysilicon 422 -774 422 -774 0 1
rlabel polysilicon 422 -780 422 -780 0 3
rlabel polysilicon 429 -774 429 -774 0 1
rlabel polysilicon 429 -780 429 -780 0 3
rlabel polysilicon 436 -774 436 -774 0 1
rlabel polysilicon 436 -780 436 -780 0 3
rlabel polysilicon 443 -774 443 -774 0 1
rlabel polysilicon 446 -774 446 -774 0 2
rlabel polysilicon 443 -780 443 -780 0 3
rlabel polysilicon 446 -780 446 -780 0 4
rlabel polysilicon 450 -774 450 -774 0 1
rlabel polysilicon 450 -780 450 -780 0 3
rlabel polysilicon 457 -774 457 -774 0 1
rlabel polysilicon 460 -774 460 -774 0 2
rlabel polysilicon 457 -780 457 -780 0 3
rlabel polysilicon 460 -780 460 -780 0 4
rlabel polysilicon 464 -780 464 -780 0 3
rlabel polysilicon 467 -780 467 -780 0 4
rlabel polysilicon 471 -774 471 -774 0 1
rlabel polysilicon 471 -780 471 -780 0 3
rlabel polysilicon 478 -774 478 -774 0 1
rlabel polysilicon 478 -780 478 -780 0 3
rlabel polysilicon 485 -774 485 -774 0 1
rlabel polysilicon 485 -780 485 -780 0 3
rlabel polysilicon 492 -774 492 -774 0 1
rlabel polysilicon 492 -780 492 -780 0 3
rlabel polysilicon 495 -780 495 -780 0 4
rlabel polysilicon 499 -774 499 -774 0 1
rlabel polysilicon 499 -780 499 -780 0 3
rlabel polysilicon 506 -774 506 -774 0 1
rlabel polysilicon 506 -780 506 -780 0 3
rlabel polysilicon 513 -774 513 -774 0 1
rlabel polysilicon 513 -780 513 -780 0 3
rlabel polysilicon 520 -774 520 -774 0 1
rlabel polysilicon 520 -780 520 -780 0 3
rlabel polysilicon 527 -774 527 -774 0 1
rlabel polysilicon 527 -780 527 -780 0 3
rlabel polysilicon 530 -780 530 -780 0 4
rlabel polysilicon 534 -774 534 -774 0 1
rlabel polysilicon 537 -774 537 -774 0 2
rlabel polysilicon 534 -780 534 -780 0 3
rlabel polysilicon 537 -780 537 -780 0 4
rlabel polysilicon 541 -774 541 -774 0 1
rlabel polysilicon 541 -780 541 -780 0 3
rlabel polysilicon 548 -774 548 -774 0 1
rlabel polysilicon 548 -780 548 -780 0 3
rlabel polysilicon 555 -774 555 -774 0 1
rlabel polysilicon 555 -780 555 -780 0 3
rlabel polysilicon 562 -774 562 -774 0 1
rlabel polysilicon 562 -780 562 -780 0 3
rlabel polysilicon 569 -774 569 -774 0 1
rlabel polysilicon 569 -780 569 -780 0 3
rlabel polysilicon 576 -774 576 -774 0 1
rlabel polysilicon 576 -780 576 -780 0 3
rlabel polysilicon 583 -774 583 -774 0 1
rlabel polysilicon 583 -780 583 -780 0 3
rlabel polysilicon 590 -774 590 -774 0 1
rlabel polysilicon 590 -780 590 -780 0 3
rlabel polysilicon 597 -774 597 -774 0 1
rlabel polysilicon 597 -780 597 -780 0 3
rlabel polysilicon 604 -774 604 -774 0 1
rlabel polysilicon 604 -780 604 -780 0 3
rlabel polysilicon 611 -774 611 -774 0 1
rlabel polysilicon 611 -780 611 -780 0 3
rlabel polysilicon 618 -774 618 -774 0 1
rlabel polysilicon 618 -780 618 -780 0 3
rlabel polysilicon 621 -780 621 -780 0 4
rlabel polysilicon 625 -774 625 -774 0 1
rlabel polysilicon 625 -780 625 -780 0 3
rlabel polysilicon 632 -774 632 -774 0 1
rlabel polysilicon 632 -780 632 -780 0 3
rlabel polysilicon 639 -774 639 -774 0 1
rlabel polysilicon 639 -780 639 -780 0 3
rlabel polysilicon 646 -774 646 -774 0 1
rlabel polysilicon 646 -780 646 -780 0 3
rlabel polysilicon 653 -774 653 -774 0 1
rlabel polysilicon 656 -774 656 -774 0 2
rlabel polysilicon 653 -780 653 -780 0 3
rlabel polysilicon 656 -780 656 -780 0 4
rlabel polysilicon 660 -774 660 -774 0 1
rlabel polysilicon 663 -774 663 -774 0 2
rlabel polysilicon 660 -780 660 -780 0 3
rlabel polysilicon 663 -780 663 -780 0 4
rlabel polysilicon 667 -774 667 -774 0 1
rlabel polysilicon 667 -780 667 -780 0 3
rlabel polysilicon 674 -774 674 -774 0 1
rlabel polysilicon 674 -780 674 -780 0 3
rlabel polysilicon 681 -774 681 -774 0 1
rlabel polysilicon 681 -780 681 -780 0 3
rlabel polysilicon 688 -774 688 -774 0 1
rlabel polysilicon 688 -780 688 -780 0 3
rlabel polysilicon 695 -774 695 -774 0 1
rlabel polysilicon 695 -780 695 -780 0 3
rlabel polysilicon 702 -774 702 -774 0 1
rlabel polysilicon 705 -774 705 -774 0 2
rlabel polysilicon 702 -780 702 -780 0 3
rlabel polysilicon 705 -780 705 -780 0 4
rlabel polysilicon 709 -774 709 -774 0 1
rlabel polysilicon 709 -780 709 -780 0 3
rlabel polysilicon 716 -774 716 -774 0 1
rlabel polysilicon 719 -774 719 -774 0 2
rlabel polysilicon 719 -780 719 -780 0 4
rlabel polysilicon 723 -774 723 -774 0 1
rlabel polysilicon 723 -780 723 -780 0 3
rlabel polysilicon 730 -774 730 -774 0 1
rlabel polysilicon 730 -780 730 -780 0 3
rlabel polysilicon 737 -774 737 -774 0 1
rlabel polysilicon 737 -780 737 -780 0 3
rlabel polysilicon 744 -774 744 -774 0 1
rlabel polysilicon 744 -780 744 -780 0 3
rlabel polysilicon 751 -774 751 -774 0 1
rlabel polysilicon 751 -780 751 -780 0 3
rlabel polysilicon 758 -774 758 -774 0 1
rlabel polysilicon 761 -774 761 -774 0 2
rlabel polysilicon 765 -774 765 -774 0 1
rlabel polysilicon 765 -780 765 -780 0 3
rlabel polysilicon 772 -774 772 -774 0 1
rlabel polysilicon 775 -774 775 -774 0 2
rlabel polysilicon 772 -780 772 -780 0 3
rlabel polysilicon 775 -780 775 -780 0 4
rlabel polysilicon 779 -774 779 -774 0 1
rlabel polysilicon 779 -780 779 -780 0 3
rlabel polysilicon 786 -774 786 -774 0 1
rlabel polysilicon 786 -780 786 -780 0 3
rlabel polysilicon 793 -780 793 -780 0 3
rlabel polysilicon 796 -780 796 -780 0 4
rlabel polysilicon 800 -774 800 -774 0 1
rlabel polysilicon 800 -780 800 -780 0 3
rlabel polysilicon 807 -774 807 -774 0 1
rlabel polysilicon 807 -780 807 -780 0 3
rlabel polysilicon 814 -774 814 -774 0 1
rlabel polysilicon 814 -780 814 -780 0 3
rlabel polysilicon 821 -774 821 -774 0 1
rlabel polysilicon 821 -780 821 -780 0 3
rlabel polysilicon 828 -774 828 -774 0 1
rlabel polysilicon 828 -780 828 -780 0 3
rlabel polysilicon 835 -774 835 -774 0 1
rlabel polysilicon 835 -780 835 -780 0 3
rlabel polysilicon 842 -774 842 -774 0 1
rlabel polysilicon 842 -780 842 -780 0 3
rlabel polysilicon 849 -774 849 -774 0 1
rlabel polysilicon 849 -780 849 -780 0 3
rlabel polysilicon 856 -774 856 -774 0 1
rlabel polysilicon 856 -780 856 -780 0 3
rlabel polysilicon 863 -774 863 -774 0 1
rlabel polysilicon 863 -780 863 -780 0 3
rlabel polysilicon 870 -774 870 -774 0 1
rlabel polysilicon 870 -780 870 -780 0 3
rlabel polysilicon 880 -774 880 -774 0 2
rlabel polysilicon 877 -780 877 -780 0 3
rlabel polysilicon 884 -774 884 -774 0 1
rlabel polysilicon 884 -780 884 -780 0 3
rlabel polysilicon 891 -774 891 -774 0 1
rlabel polysilicon 891 -780 891 -780 0 3
rlabel polysilicon 898 -774 898 -774 0 1
rlabel polysilicon 898 -780 898 -780 0 3
rlabel polysilicon 905 -774 905 -774 0 1
rlabel polysilicon 905 -780 905 -780 0 3
rlabel polysilicon 912 -774 912 -774 0 1
rlabel polysilicon 912 -780 912 -780 0 3
rlabel polysilicon 919 -774 919 -774 0 1
rlabel polysilicon 919 -780 919 -780 0 3
rlabel polysilicon 926 -774 926 -774 0 1
rlabel polysilicon 926 -780 926 -780 0 3
rlabel polysilicon 933 -774 933 -774 0 1
rlabel polysilicon 936 -774 936 -774 0 2
rlabel polysilicon 936 -780 936 -780 0 4
rlabel polysilicon 940 -774 940 -774 0 1
rlabel polysilicon 940 -780 940 -780 0 3
rlabel polysilicon 950 -774 950 -774 0 2
rlabel polysilicon 947 -780 947 -780 0 3
rlabel polysilicon 954 -774 954 -774 0 1
rlabel polysilicon 957 -780 957 -780 0 4
rlabel polysilicon 961 -774 961 -774 0 1
rlabel polysilicon 961 -780 961 -780 0 3
rlabel polysilicon 968 -774 968 -774 0 1
rlabel polysilicon 968 -780 968 -780 0 3
rlabel polysilicon 975 -774 975 -774 0 1
rlabel polysilicon 975 -780 975 -780 0 3
rlabel polysilicon 982 -774 982 -774 0 1
rlabel polysilicon 982 -780 982 -780 0 3
rlabel polysilicon 989 -774 989 -774 0 1
rlabel polysilicon 989 -780 989 -780 0 3
rlabel polysilicon 996 -774 996 -774 0 1
rlabel polysilicon 996 -780 996 -780 0 3
rlabel polysilicon 1003 -774 1003 -774 0 1
rlabel polysilicon 1003 -780 1003 -780 0 3
rlabel polysilicon 1010 -780 1010 -780 0 3
rlabel polysilicon 1031 -774 1031 -774 0 1
rlabel polysilicon 1031 -780 1031 -780 0 3
rlabel polysilicon 1122 -774 1122 -774 0 1
rlabel polysilicon 1122 -780 1122 -780 0 3
rlabel polysilicon 2 -861 2 -861 0 1
rlabel polysilicon 2 -867 2 -867 0 3
rlabel polysilicon 12 -867 12 -867 0 4
rlabel polysilicon 16 -861 16 -861 0 1
rlabel polysilicon 16 -867 16 -867 0 3
rlabel polysilicon 23 -861 23 -861 0 1
rlabel polysilicon 23 -867 23 -867 0 3
rlabel polysilicon 30 -861 30 -861 0 1
rlabel polysilicon 30 -867 30 -867 0 3
rlabel polysilicon 37 -861 37 -861 0 1
rlabel polysilicon 40 -861 40 -861 0 2
rlabel polysilicon 44 -861 44 -861 0 1
rlabel polysilicon 44 -867 44 -867 0 3
rlabel polysilicon 51 -861 51 -861 0 1
rlabel polysilicon 51 -867 51 -867 0 3
rlabel polysilicon 58 -861 58 -861 0 1
rlabel polysilicon 58 -867 58 -867 0 3
rlabel polysilicon 65 -861 65 -861 0 1
rlabel polysilicon 65 -867 65 -867 0 3
rlabel polysilicon 75 -861 75 -861 0 2
rlabel polysilicon 72 -867 72 -867 0 3
rlabel polysilicon 75 -867 75 -867 0 4
rlabel polysilicon 82 -861 82 -861 0 2
rlabel polysilicon 79 -867 79 -867 0 3
rlabel polysilicon 82 -867 82 -867 0 4
rlabel polysilicon 86 -861 86 -861 0 1
rlabel polysilicon 86 -867 86 -867 0 3
rlabel polysilicon 93 -861 93 -861 0 1
rlabel polysilicon 93 -867 93 -867 0 3
rlabel polysilicon 100 -861 100 -861 0 1
rlabel polysilicon 100 -867 100 -867 0 3
rlabel polysilicon 107 -861 107 -861 0 1
rlabel polysilicon 107 -867 107 -867 0 3
rlabel polysilicon 114 -861 114 -861 0 1
rlabel polysilicon 114 -867 114 -867 0 3
rlabel polysilicon 121 -861 121 -861 0 1
rlabel polysilicon 121 -867 121 -867 0 3
rlabel polysilicon 128 -861 128 -861 0 1
rlabel polysilicon 128 -867 128 -867 0 3
rlabel polysilicon 135 -861 135 -861 0 1
rlabel polysilicon 135 -867 135 -867 0 3
rlabel polysilicon 142 -861 142 -861 0 1
rlabel polysilicon 142 -867 142 -867 0 3
rlabel polysilicon 149 -861 149 -861 0 1
rlabel polysilicon 149 -867 149 -867 0 3
rlabel polysilicon 156 -861 156 -861 0 1
rlabel polysilicon 156 -867 156 -867 0 3
rlabel polysilicon 163 -861 163 -861 0 1
rlabel polysilicon 163 -867 163 -867 0 3
rlabel polysilicon 170 -861 170 -861 0 1
rlabel polysilicon 170 -867 170 -867 0 3
rlabel polysilicon 177 -861 177 -861 0 1
rlabel polysilicon 177 -867 177 -867 0 3
rlabel polysilicon 184 -861 184 -861 0 1
rlabel polysilicon 184 -867 184 -867 0 3
rlabel polysilicon 194 -861 194 -861 0 2
rlabel polysilicon 191 -867 191 -867 0 3
rlabel polysilicon 194 -867 194 -867 0 4
rlabel polysilicon 198 -861 198 -861 0 1
rlabel polysilicon 198 -867 198 -867 0 3
rlabel polysilicon 205 -861 205 -861 0 1
rlabel polysilicon 205 -867 205 -867 0 3
rlabel polysilicon 212 -861 212 -861 0 1
rlabel polysilicon 212 -867 212 -867 0 3
rlabel polysilicon 219 -861 219 -861 0 1
rlabel polysilicon 222 -861 222 -861 0 2
rlabel polysilicon 222 -867 222 -867 0 4
rlabel polysilicon 226 -861 226 -861 0 1
rlabel polysilicon 226 -867 226 -867 0 3
rlabel polysilicon 229 -867 229 -867 0 4
rlabel polysilicon 233 -861 233 -861 0 1
rlabel polysilicon 233 -867 233 -867 0 3
rlabel polysilicon 240 -861 240 -861 0 1
rlabel polysilicon 240 -867 240 -867 0 3
rlabel polysilicon 247 -861 247 -861 0 1
rlabel polysilicon 247 -867 247 -867 0 3
rlabel polysilicon 254 -861 254 -861 0 1
rlabel polysilicon 254 -867 254 -867 0 3
rlabel polysilicon 261 -861 261 -861 0 1
rlabel polysilicon 268 -861 268 -861 0 1
rlabel polysilicon 268 -867 268 -867 0 3
rlabel polysilicon 275 -861 275 -861 0 1
rlabel polysilicon 275 -867 275 -867 0 3
rlabel polysilicon 282 -861 282 -861 0 1
rlabel polysilicon 282 -867 282 -867 0 3
rlabel polysilicon 289 -861 289 -861 0 1
rlabel polysilicon 289 -867 289 -867 0 3
rlabel polysilicon 296 -861 296 -861 0 1
rlabel polysilicon 296 -867 296 -867 0 3
rlabel polysilicon 303 -861 303 -861 0 1
rlabel polysilicon 303 -867 303 -867 0 3
rlabel polysilicon 310 -861 310 -861 0 1
rlabel polysilicon 310 -867 310 -867 0 3
rlabel polysilicon 317 -861 317 -861 0 1
rlabel polysilicon 317 -867 317 -867 0 3
rlabel polysilicon 324 -861 324 -861 0 1
rlabel polysilicon 327 -861 327 -861 0 2
rlabel polysilicon 324 -867 324 -867 0 3
rlabel polysilicon 331 -861 331 -861 0 1
rlabel polysilicon 331 -867 331 -867 0 3
rlabel polysilicon 338 -861 338 -861 0 1
rlabel polysilicon 341 -861 341 -861 0 2
rlabel polysilicon 338 -867 338 -867 0 3
rlabel polysilicon 341 -867 341 -867 0 4
rlabel polysilicon 345 -861 345 -861 0 1
rlabel polysilicon 345 -867 345 -867 0 3
rlabel polysilicon 352 -861 352 -861 0 1
rlabel polysilicon 355 -861 355 -861 0 2
rlabel polysilicon 352 -867 352 -867 0 3
rlabel polysilicon 355 -867 355 -867 0 4
rlabel polysilicon 359 -861 359 -861 0 1
rlabel polysilicon 359 -867 359 -867 0 3
rlabel polysilicon 366 -861 366 -861 0 1
rlabel polysilicon 366 -867 366 -867 0 3
rlabel polysilicon 373 -861 373 -861 0 1
rlabel polysilicon 373 -867 373 -867 0 3
rlabel polysilicon 383 -861 383 -861 0 2
rlabel polysilicon 380 -867 380 -867 0 3
rlabel polysilicon 383 -867 383 -867 0 4
rlabel polysilicon 387 -861 387 -861 0 1
rlabel polysilicon 387 -867 387 -867 0 3
rlabel polysilicon 394 -861 394 -861 0 1
rlabel polysilicon 394 -867 394 -867 0 3
rlabel polysilicon 397 -867 397 -867 0 4
rlabel polysilicon 401 -861 401 -861 0 1
rlabel polysilicon 401 -867 401 -867 0 3
rlabel polysilicon 408 -861 408 -861 0 1
rlabel polysilicon 408 -867 408 -867 0 3
rlabel polysilicon 415 -861 415 -861 0 1
rlabel polysilicon 415 -867 415 -867 0 3
rlabel polysilicon 422 -861 422 -861 0 1
rlabel polysilicon 422 -867 422 -867 0 3
rlabel polysilicon 429 -867 429 -867 0 3
rlabel polysilicon 432 -867 432 -867 0 4
rlabel polysilicon 436 -861 436 -861 0 1
rlabel polysilicon 436 -867 436 -867 0 3
rlabel polysilicon 443 -861 443 -861 0 1
rlabel polysilicon 443 -867 443 -867 0 3
rlabel polysilicon 450 -861 450 -861 0 1
rlabel polysilicon 453 -861 453 -861 0 2
rlabel polysilicon 450 -867 450 -867 0 3
rlabel polysilicon 453 -867 453 -867 0 4
rlabel polysilicon 457 -861 457 -861 0 1
rlabel polysilicon 457 -867 457 -867 0 3
rlabel polysilicon 464 -861 464 -861 0 1
rlabel polysilicon 464 -867 464 -867 0 3
rlabel polysilicon 471 -861 471 -861 0 1
rlabel polysilicon 471 -867 471 -867 0 3
rlabel polysilicon 478 -861 478 -861 0 1
rlabel polysilicon 481 -861 481 -861 0 2
rlabel polysilicon 481 -867 481 -867 0 4
rlabel polysilicon 485 -861 485 -861 0 1
rlabel polysilicon 485 -867 485 -867 0 3
rlabel polysilicon 492 -861 492 -861 0 1
rlabel polysilicon 492 -867 492 -867 0 3
rlabel polysilicon 499 -861 499 -861 0 1
rlabel polysilicon 502 -861 502 -861 0 2
rlabel polysilicon 499 -867 499 -867 0 3
rlabel polysilicon 506 -861 506 -861 0 1
rlabel polysilicon 506 -867 506 -867 0 3
rlabel polysilicon 513 -861 513 -861 0 1
rlabel polysilicon 513 -867 513 -867 0 3
rlabel polysilicon 520 -861 520 -861 0 1
rlabel polysilicon 520 -867 520 -867 0 3
rlabel polysilicon 527 -861 527 -861 0 1
rlabel polysilicon 527 -867 527 -867 0 3
rlabel polysilicon 534 -861 534 -861 0 1
rlabel polysilicon 534 -867 534 -867 0 3
rlabel polysilicon 541 -861 541 -861 0 1
rlabel polysilicon 541 -867 541 -867 0 3
rlabel polysilicon 544 -867 544 -867 0 4
rlabel polysilicon 548 -861 548 -861 0 1
rlabel polysilicon 548 -867 548 -867 0 3
rlabel polysilicon 555 -861 555 -861 0 1
rlabel polysilicon 555 -867 555 -867 0 3
rlabel polysilicon 558 -867 558 -867 0 4
rlabel polysilicon 565 -861 565 -861 0 2
rlabel polysilicon 562 -867 562 -867 0 3
rlabel polysilicon 565 -867 565 -867 0 4
rlabel polysilicon 569 -861 569 -861 0 1
rlabel polysilicon 569 -867 569 -867 0 3
rlabel polysilicon 576 -861 576 -861 0 1
rlabel polysilicon 579 -861 579 -861 0 2
rlabel polysilicon 576 -867 576 -867 0 3
rlabel polysilicon 579 -867 579 -867 0 4
rlabel polysilicon 583 -861 583 -861 0 1
rlabel polysilicon 583 -867 583 -867 0 3
rlabel polysilicon 593 -861 593 -861 0 2
rlabel polysilicon 590 -867 590 -867 0 3
rlabel polysilicon 593 -867 593 -867 0 4
rlabel polysilicon 597 -861 597 -861 0 1
rlabel polysilicon 597 -867 597 -867 0 3
rlabel polysilicon 604 -861 604 -861 0 1
rlabel polysilicon 607 -861 607 -861 0 2
rlabel polysilicon 604 -867 604 -867 0 3
rlabel polysilicon 611 -861 611 -861 0 1
rlabel polysilicon 614 -861 614 -861 0 2
rlabel polysilicon 611 -867 611 -867 0 3
rlabel polysilicon 614 -867 614 -867 0 4
rlabel polysilicon 618 -861 618 -861 0 1
rlabel polysilicon 618 -867 618 -867 0 3
rlabel polysilicon 625 -861 625 -861 0 1
rlabel polysilicon 625 -867 625 -867 0 3
rlabel polysilicon 632 -861 632 -861 0 1
rlabel polysilicon 635 -861 635 -861 0 2
rlabel polysilicon 632 -867 632 -867 0 3
rlabel polysilicon 635 -867 635 -867 0 4
rlabel polysilicon 639 -861 639 -861 0 1
rlabel polysilicon 639 -867 639 -867 0 3
rlabel polysilicon 646 -861 646 -861 0 1
rlabel polysilicon 646 -867 646 -867 0 3
rlabel polysilicon 653 -861 653 -861 0 1
rlabel polysilicon 656 -861 656 -861 0 2
rlabel polysilicon 660 -861 660 -861 0 1
rlabel polysilicon 660 -867 660 -867 0 3
rlabel polysilicon 667 -861 667 -861 0 1
rlabel polysilicon 667 -867 667 -867 0 3
rlabel polysilicon 674 -861 674 -861 0 1
rlabel polysilicon 674 -867 674 -867 0 3
rlabel polysilicon 681 -861 681 -861 0 1
rlabel polysilicon 681 -867 681 -867 0 3
rlabel polysilicon 688 -861 688 -861 0 1
rlabel polysilicon 688 -867 688 -867 0 3
rlabel polysilicon 695 -861 695 -861 0 1
rlabel polysilicon 695 -867 695 -867 0 3
rlabel polysilicon 702 -861 702 -861 0 1
rlabel polysilicon 702 -867 702 -867 0 3
rlabel polysilicon 709 -861 709 -861 0 1
rlabel polysilicon 709 -867 709 -867 0 3
rlabel polysilicon 716 -861 716 -861 0 1
rlabel polysilicon 716 -867 716 -867 0 3
rlabel polysilicon 723 -861 723 -861 0 1
rlabel polysilicon 723 -867 723 -867 0 3
rlabel polysilicon 730 -861 730 -861 0 1
rlabel polysilicon 730 -867 730 -867 0 3
rlabel polysilicon 737 -861 737 -861 0 1
rlabel polysilicon 737 -867 737 -867 0 3
rlabel polysilicon 744 -861 744 -861 0 1
rlabel polysilicon 744 -867 744 -867 0 3
rlabel polysilicon 751 -861 751 -861 0 1
rlabel polysilicon 751 -867 751 -867 0 3
rlabel polysilicon 758 -861 758 -861 0 1
rlabel polysilicon 758 -867 758 -867 0 3
rlabel polysilicon 765 -861 765 -861 0 1
rlabel polysilicon 768 -861 768 -861 0 2
rlabel polysilicon 768 -867 768 -867 0 4
rlabel polysilicon 772 -861 772 -861 0 1
rlabel polysilicon 772 -867 772 -867 0 3
rlabel polysilicon 779 -861 779 -861 0 1
rlabel polysilicon 779 -867 779 -867 0 3
rlabel polysilicon 786 -861 786 -861 0 1
rlabel polysilicon 786 -867 786 -867 0 3
rlabel polysilicon 793 -861 793 -861 0 1
rlabel polysilicon 793 -867 793 -867 0 3
rlabel polysilicon 800 -861 800 -861 0 1
rlabel polysilicon 800 -867 800 -867 0 3
rlabel polysilicon 807 -861 807 -861 0 1
rlabel polysilicon 807 -867 807 -867 0 3
rlabel polysilicon 814 -861 814 -861 0 1
rlabel polysilicon 814 -867 814 -867 0 3
rlabel polysilicon 821 -861 821 -861 0 1
rlabel polysilicon 821 -867 821 -867 0 3
rlabel polysilicon 828 -861 828 -861 0 1
rlabel polysilicon 828 -867 828 -867 0 3
rlabel polysilicon 835 -861 835 -861 0 1
rlabel polysilicon 835 -867 835 -867 0 3
rlabel polysilicon 842 -861 842 -861 0 1
rlabel polysilicon 842 -867 842 -867 0 3
rlabel polysilicon 849 -861 849 -861 0 1
rlabel polysilicon 849 -867 849 -867 0 3
rlabel polysilicon 856 -861 856 -861 0 1
rlabel polysilicon 856 -867 856 -867 0 3
rlabel polysilicon 863 -861 863 -861 0 1
rlabel polysilicon 866 -861 866 -861 0 2
rlabel polysilicon 870 -861 870 -861 0 1
rlabel polysilicon 870 -867 870 -867 0 3
rlabel polysilicon 877 -861 877 -861 0 1
rlabel polysilicon 877 -867 877 -867 0 3
rlabel polysilicon 884 -861 884 -861 0 1
rlabel polysilicon 884 -867 884 -867 0 3
rlabel polysilicon 891 -861 891 -861 0 1
rlabel polysilicon 891 -867 891 -867 0 3
rlabel polysilicon 898 -861 898 -861 0 1
rlabel polysilicon 898 -867 898 -867 0 3
rlabel polysilicon 905 -861 905 -861 0 1
rlabel polysilicon 905 -867 905 -867 0 3
rlabel polysilicon 912 -861 912 -861 0 1
rlabel polysilicon 912 -867 912 -867 0 3
rlabel polysilicon 919 -861 919 -861 0 1
rlabel polysilicon 919 -867 919 -867 0 3
rlabel polysilicon 926 -861 926 -861 0 1
rlabel polysilicon 926 -867 926 -867 0 3
rlabel polysilicon 933 -861 933 -861 0 1
rlabel polysilicon 933 -867 933 -867 0 3
rlabel polysilicon 940 -861 940 -861 0 1
rlabel polysilicon 940 -867 940 -867 0 3
rlabel polysilicon 947 -861 947 -861 0 1
rlabel polysilicon 947 -867 947 -867 0 3
rlabel polysilicon 954 -861 954 -861 0 1
rlabel polysilicon 954 -867 954 -867 0 3
rlabel polysilicon 961 -861 961 -861 0 1
rlabel polysilicon 961 -867 961 -867 0 3
rlabel polysilicon 968 -861 968 -861 0 1
rlabel polysilicon 968 -867 968 -867 0 3
rlabel polysilicon 975 -861 975 -861 0 1
rlabel polysilicon 975 -867 975 -867 0 3
rlabel polysilicon 982 -861 982 -861 0 1
rlabel polysilicon 982 -867 982 -867 0 3
rlabel polysilicon 989 -861 989 -861 0 1
rlabel polysilicon 989 -867 989 -867 0 3
rlabel polysilicon 996 -861 996 -861 0 1
rlabel polysilicon 996 -867 996 -867 0 3
rlabel polysilicon 1003 -861 1003 -861 0 1
rlabel polysilicon 1003 -867 1003 -867 0 3
rlabel polysilicon 1010 -861 1010 -861 0 1
rlabel polysilicon 1010 -867 1010 -867 0 3
rlabel polysilicon 1017 -861 1017 -861 0 1
rlabel polysilicon 1017 -867 1017 -867 0 3
rlabel polysilicon 1024 -861 1024 -861 0 1
rlabel polysilicon 1024 -867 1024 -867 0 3
rlabel polysilicon 1031 -861 1031 -861 0 1
rlabel polysilicon 1031 -867 1031 -867 0 3
rlabel polysilicon 1038 -861 1038 -861 0 1
rlabel polysilicon 1038 -867 1038 -867 0 3
rlabel polysilicon 1045 -861 1045 -861 0 1
rlabel polysilicon 1045 -867 1045 -867 0 3
rlabel polysilicon 1052 -861 1052 -861 0 1
rlabel polysilicon 1052 -867 1052 -867 0 3
rlabel polysilicon 1059 -861 1059 -861 0 1
rlabel polysilicon 1059 -867 1059 -867 0 3
rlabel polysilicon 1066 -861 1066 -861 0 1
rlabel polysilicon 1066 -867 1066 -867 0 3
rlabel polysilicon 1073 -861 1073 -861 0 1
rlabel polysilicon 1073 -867 1073 -867 0 3
rlabel polysilicon 1080 -861 1080 -861 0 1
rlabel polysilicon 1080 -867 1080 -867 0 3
rlabel polysilicon 1087 -861 1087 -861 0 1
rlabel polysilicon 1087 -867 1087 -867 0 3
rlabel polysilicon 1094 -861 1094 -861 0 1
rlabel polysilicon 1097 -867 1097 -867 0 4
rlabel polysilicon 1101 -861 1101 -861 0 1
rlabel polysilicon 1101 -867 1101 -867 0 3
rlabel polysilicon 1108 -861 1108 -861 0 1
rlabel polysilicon 1108 -867 1108 -867 0 3
rlabel polysilicon 1115 -861 1115 -861 0 1
rlabel polysilicon 1115 -867 1115 -867 0 3
rlabel polysilicon 1122 -861 1122 -861 0 1
rlabel polysilicon 1122 -867 1122 -867 0 3
rlabel polysilicon 1129 -867 1129 -867 0 3
rlabel polysilicon 1139 -861 1139 -861 0 2
rlabel polysilicon 1136 -867 1136 -867 0 3
rlabel polysilicon 1143 -861 1143 -861 0 1
rlabel polysilicon 1143 -867 1143 -867 0 3
rlabel polysilicon 1150 -861 1150 -861 0 1
rlabel polysilicon 1153 -861 1153 -861 0 2
rlabel polysilicon 2 -968 2 -968 0 3
rlabel polysilicon 9 -962 9 -962 0 1
rlabel polysilicon 9 -968 9 -968 0 3
rlabel polysilicon 16 -962 16 -962 0 1
rlabel polysilicon 16 -968 16 -968 0 3
rlabel polysilicon 23 -962 23 -962 0 1
rlabel polysilicon 23 -968 23 -968 0 3
rlabel polysilicon 30 -962 30 -962 0 1
rlabel polysilicon 30 -968 30 -968 0 3
rlabel polysilicon 37 -962 37 -962 0 1
rlabel polysilicon 37 -968 37 -968 0 3
rlabel polysilicon 44 -962 44 -962 0 1
rlabel polysilicon 44 -968 44 -968 0 3
rlabel polysilicon 51 -962 51 -962 0 1
rlabel polysilicon 51 -968 51 -968 0 3
rlabel polysilicon 58 -962 58 -962 0 1
rlabel polysilicon 58 -968 58 -968 0 3
rlabel polysilicon 65 -962 65 -962 0 1
rlabel polysilicon 65 -968 65 -968 0 3
rlabel polysilicon 68 -968 68 -968 0 4
rlabel polysilicon 72 -962 72 -962 0 1
rlabel polysilicon 75 -962 75 -962 0 2
rlabel polysilicon 72 -968 72 -968 0 3
rlabel polysilicon 75 -968 75 -968 0 4
rlabel polysilicon 79 -962 79 -962 0 1
rlabel polysilicon 82 -962 82 -962 0 2
rlabel polysilicon 82 -968 82 -968 0 4
rlabel polysilicon 86 -962 86 -962 0 1
rlabel polysilicon 86 -968 86 -968 0 3
rlabel polysilicon 93 -962 93 -962 0 1
rlabel polysilicon 93 -968 93 -968 0 3
rlabel polysilicon 100 -962 100 -962 0 1
rlabel polysilicon 100 -968 100 -968 0 3
rlabel polysilicon 107 -962 107 -962 0 1
rlabel polysilicon 107 -968 107 -968 0 3
rlabel polysilicon 114 -962 114 -962 0 1
rlabel polysilicon 114 -968 114 -968 0 3
rlabel polysilicon 121 -962 121 -962 0 1
rlabel polysilicon 121 -968 121 -968 0 3
rlabel polysilicon 128 -962 128 -962 0 1
rlabel polysilicon 128 -968 128 -968 0 3
rlabel polysilicon 135 -962 135 -962 0 1
rlabel polysilicon 135 -968 135 -968 0 3
rlabel polysilicon 142 -962 142 -962 0 1
rlabel polysilicon 142 -968 142 -968 0 3
rlabel polysilicon 149 -962 149 -962 0 1
rlabel polysilicon 152 -962 152 -962 0 2
rlabel polysilicon 156 -962 156 -962 0 1
rlabel polysilicon 156 -968 156 -968 0 3
rlabel polysilicon 163 -962 163 -962 0 1
rlabel polysilicon 163 -968 163 -968 0 3
rlabel polysilicon 170 -962 170 -962 0 1
rlabel polysilicon 170 -968 170 -968 0 3
rlabel polysilicon 177 -962 177 -962 0 1
rlabel polysilicon 177 -968 177 -968 0 3
rlabel polysilicon 184 -962 184 -962 0 1
rlabel polysilicon 184 -968 184 -968 0 3
rlabel polysilicon 191 -962 191 -962 0 1
rlabel polysilicon 191 -968 191 -968 0 3
rlabel polysilicon 198 -962 198 -962 0 1
rlabel polysilicon 198 -968 198 -968 0 3
rlabel polysilicon 205 -962 205 -962 0 1
rlabel polysilicon 205 -968 205 -968 0 3
rlabel polysilicon 212 -962 212 -962 0 1
rlabel polysilicon 212 -968 212 -968 0 3
rlabel polysilicon 219 -962 219 -962 0 1
rlabel polysilicon 219 -968 219 -968 0 3
rlabel polysilicon 226 -962 226 -962 0 1
rlabel polysilicon 226 -968 226 -968 0 3
rlabel polysilicon 233 -962 233 -962 0 1
rlabel polysilicon 233 -968 233 -968 0 3
rlabel polysilicon 240 -962 240 -962 0 1
rlabel polysilicon 240 -968 240 -968 0 3
rlabel polysilicon 247 -962 247 -962 0 1
rlabel polysilicon 247 -968 247 -968 0 3
rlabel polysilicon 254 -962 254 -962 0 1
rlabel polysilicon 254 -968 254 -968 0 3
rlabel polysilicon 261 -962 261 -962 0 1
rlabel polysilicon 261 -968 261 -968 0 3
rlabel polysilicon 268 -962 268 -962 0 1
rlabel polysilicon 268 -968 268 -968 0 3
rlabel polysilicon 275 -962 275 -962 0 1
rlabel polysilicon 275 -968 275 -968 0 3
rlabel polysilicon 282 -968 282 -968 0 3
rlabel polysilicon 285 -968 285 -968 0 4
rlabel polysilicon 289 -962 289 -962 0 1
rlabel polysilicon 289 -968 289 -968 0 3
rlabel polysilicon 299 -962 299 -962 0 2
rlabel polysilicon 303 -962 303 -962 0 1
rlabel polysilicon 303 -968 303 -968 0 3
rlabel polysilicon 306 -968 306 -968 0 4
rlabel polysilicon 310 -962 310 -962 0 1
rlabel polysilicon 310 -968 310 -968 0 3
rlabel polysilicon 317 -962 317 -962 0 1
rlabel polysilicon 317 -968 317 -968 0 3
rlabel polysilicon 324 -962 324 -962 0 1
rlabel polysilicon 324 -968 324 -968 0 3
rlabel polysilicon 331 -962 331 -962 0 1
rlabel polysilicon 331 -968 331 -968 0 3
rlabel polysilicon 338 -962 338 -962 0 1
rlabel polysilicon 338 -968 338 -968 0 3
rlabel polysilicon 345 -962 345 -962 0 1
rlabel polysilicon 345 -968 345 -968 0 3
rlabel polysilicon 352 -962 352 -962 0 1
rlabel polysilicon 352 -968 352 -968 0 3
rlabel polysilicon 359 -962 359 -962 0 1
rlabel polysilicon 362 -962 362 -962 0 2
rlabel polysilicon 362 -968 362 -968 0 4
rlabel polysilicon 366 -962 366 -962 0 1
rlabel polysilicon 366 -968 366 -968 0 3
rlabel polysilicon 373 -962 373 -962 0 1
rlabel polysilicon 373 -968 373 -968 0 3
rlabel polysilicon 380 -962 380 -962 0 1
rlabel polysilicon 380 -968 380 -968 0 3
rlabel polysilicon 387 -962 387 -962 0 1
rlabel polysilicon 387 -968 387 -968 0 3
rlabel polysilicon 394 -962 394 -962 0 1
rlabel polysilicon 394 -968 394 -968 0 3
rlabel polysilicon 401 -962 401 -962 0 1
rlabel polysilicon 401 -968 401 -968 0 3
rlabel polysilicon 408 -962 408 -962 0 1
rlabel polysilicon 408 -968 408 -968 0 3
rlabel polysilicon 415 -962 415 -962 0 1
rlabel polysilicon 418 -962 418 -962 0 2
rlabel polysilicon 415 -968 415 -968 0 3
rlabel polysilicon 418 -968 418 -968 0 4
rlabel polysilicon 422 -962 422 -962 0 1
rlabel polysilicon 422 -968 422 -968 0 3
rlabel polysilicon 429 -962 429 -962 0 1
rlabel polysilicon 429 -968 429 -968 0 3
rlabel polysilicon 439 -962 439 -962 0 2
rlabel polysilicon 436 -968 436 -968 0 3
rlabel polysilicon 439 -968 439 -968 0 4
rlabel polysilicon 443 -962 443 -962 0 1
rlabel polysilicon 446 -962 446 -962 0 2
rlabel polysilicon 446 -968 446 -968 0 4
rlabel polysilicon 450 -962 450 -962 0 1
rlabel polysilicon 450 -968 450 -968 0 3
rlabel polysilicon 457 -962 457 -962 0 1
rlabel polysilicon 457 -968 457 -968 0 3
rlabel polysilicon 464 -962 464 -962 0 1
rlabel polysilicon 467 -968 467 -968 0 4
rlabel polysilicon 471 -962 471 -962 0 1
rlabel polysilicon 471 -968 471 -968 0 3
rlabel polysilicon 474 -968 474 -968 0 4
rlabel polysilicon 478 -962 478 -962 0 1
rlabel polysilicon 481 -962 481 -962 0 2
rlabel polysilicon 478 -968 478 -968 0 3
rlabel polysilicon 481 -968 481 -968 0 4
rlabel polysilicon 485 -962 485 -962 0 1
rlabel polysilicon 485 -968 485 -968 0 3
rlabel polysilicon 492 -962 492 -962 0 1
rlabel polysilicon 492 -968 492 -968 0 3
rlabel polysilicon 502 -962 502 -962 0 2
rlabel polysilicon 499 -968 499 -968 0 3
rlabel polysilicon 502 -968 502 -968 0 4
rlabel polysilicon 506 -962 506 -962 0 1
rlabel polysilicon 506 -968 506 -968 0 3
rlabel polysilicon 513 -962 513 -962 0 1
rlabel polysilicon 513 -968 513 -968 0 3
rlabel polysilicon 520 -962 520 -962 0 1
rlabel polysilicon 520 -968 520 -968 0 3
rlabel polysilicon 527 -962 527 -962 0 1
rlabel polysilicon 527 -968 527 -968 0 3
rlabel polysilicon 537 -962 537 -962 0 2
rlabel polysilicon 534 -968 534 -968 0 3
rlabel polysilicon 541 -962 541 -962 0 1
rlabel polysilicon 544 -962 544 -962 0 2
rlabel polysilicon 544 -968 544 -968 0 4
rlabel polysilicon 548 -962 548 -962 0 1
rlabel polysilicon 548 -968 548 -968 0 3
rlabel polysilicon 555 -962 555 -962 0 1
rlabel polysilicon 555 -968 555 -968 0 3
rlabel polysilicon 562 -962 562 -962 0 1
rlabel polysilicon 562 -968 562 -968 0 3
rlabel polysilicon 569 -962 569 -962 0 1
rlabel polysilicon 572 -962 572 -962 0 2
rlabel polysilicon 569 -968 569 -968 0 3
rlabel polysilicon 572 -968 572 -968 0 4
rlabel polysilicon 576 -962 576 -962 0 1
rlabel polysilicon 579 -962 579 -962 0 2
rlabel polysilicon 579 -968 579 -968 0 4
rlabel polysilicon 583 -962 583 -962 0 1
rlabel polysilicon 583 -968 583 -968 0 3
rlabel polysilicon 593 -962 593 -962 0 2
rlabel polysilicon 590 -968 590 -968 0 3
rlabel polysilicon 593 -968 593 -968 0 4
rlabel polysilicon 597 -962 597 -962 0 1
rlabel polysilicon 597 -968 597 -968 0 3
rlabel polysilicon 604 -962 604 -962 0 1
rlabel polysilicon 604 -968 604 -968 0 3
rlabel polysilicon 614 -962 614 -962 0 2
rlabel polysilicon 611 -968 611 -968 0 3
rlabel polysilicon 614 -968 614 -968 0 4
rlabel polysilicon 618 -962 618 -962 0 1
rlabel polysilicon 621 -962 621 -962 0 2
rlabel polysilicon 618 -968 618 -968 0 3
rlabel polysilicon 621 -968 621 -968 0 4
rlabel polysilicon 625 -962 625 -962 0 1
rlabel polysilicon 625 -968 625 -968 0 3
rlabel polysilicon 628 -968 628 -968 0 4
rlabel polysilicon 632 -962 632 -962 0 1
rlabel polysilicon 635 -968 635 -968 0 4
rlabel polysilicon 639 -962 639 -962 0 1
rlabel polysilicon 639 -968 639 -968 0 3
rlabel polysilicon 646 -962 646 -962 0 1
rlabel polysilicon 646 -968 646 -968 0 3
rlabel polysilicon 653 -962 653 -962 0 1
rlabel polysilicon 653 -968 653 -968 0 3
rlabel polysilicon 660 -962 660 -962 0 1
rlabel polysilicon 660 -968 660 -968 0 3
rlabel polysilicon 667 -962 667 -962 0 1
rlabel polysilicon 667 -968 667 -968 0 3
rlabel polysilicon 674 -962 674 -962 0 1
rlabel polysilicon 674 -968 674 -968 0 3
rlabel polysilicon 681 -962 681 -962 0 1
rlabel polysilicon 681 -968 681 -968 0 3
rlabel polysilicon 688 -962 688 -962 0 1
rlabel polysilicon 691 -962 691 -962 0 2
rlabel polysilicon 691 -968 691 -968 0 4
rlabel polysilicon 698 -962 698 -962 0 2
rlabel polysilicon 698 -968 698 -968 0 4
rlabel polysilicon 702 -962 702 -962 0 1
rlabel polysilicon 702 -968 702 -968 0 3
rlabel polysilicon 709 -962 709 -962 0 1
rlabel polysilicon 709 -968 709 -968 0 3
rlabel polysilicon 716 -962 716 -962 0 1
rlabel polysilicon 716 -968 716 -968 0 3
rlabel polysilicon 723 -962 723 -962 0 1
rlabel polysilicon 723 -968 723 -968 0 3
rlabel polysilicon 730 -962 730 -962 0 1
rlabel polysilicon 730 -968 730 -968 0 3
rlabel polysilicon 737 -962 737 -962 0 1
rlabel polysilicon 737 -968 737 -968 0 3
rlabel polysilicon 744 -962 744 -962 0 1
rlabel polysilicon 744 -968 744 -968 0 3
rlabel polysilicon 751 -962 751 -962 0 1
rlabel polysilicon 751 -968 751 -968 0 3
rlabel polysilicon 758 -962 758 -962 0 1
rlabel polysilicon 758 -968 758 -968 0 3
rlabel polysilicon 765 -962 765 -962 0 1
rlabel polysilicon 765 -968 765 -968 0 3
rlabel polysilicon 772 -962 772 -962 0 1
rlabel polysilicon 772 -968 772 -968 0 3
rlabel polysilicon 779 -962 779 -962 0 1
rlabel polysilicon 779 -968 779 -968 0 3
rlabel polysilicon 786 -962 786 -962 0 1
rlabel polysilicon 786 -968 786 -968 0 3
rlabel polysilicon 793 -962 793 -962 0 1
rlabel polysilicon 793 -968 793 -968 0 3
rlabel polysilicon 800 -962 800 -962 0 1
rlabel polysilicon 800 -968 800 -968 0 3
rlabel polysilicon 807 -962 807 -962 0 1
rlabel polysilicon 807 -968 807 -968 0 3
rlabel polysilicon 814 -962 814 -962 0 1
rlabel polysilicon 814 -968 814 -968 0 3
rlabel polysilicon 821 -962 821 -962 0 1
rlabel polysilicon 821 -968 821 -968 0 3
rlabel polysilicon 828 -962 828 -962 0 1
rlabel polysilicon 828 -968 828 -968 0 3
rlabel polysilicon 835 -962 835 -962 0 1
rlabel polysilicon 835 -968 835 -968 0 3
rlabel polysilicon 842 -962 842 -962 0 1
rlabel polysilicon 842 -968 842 -968 0 3
rlabel polysilicon 849 -962 849 -962 0 1
rlabel polysilicon 849 -968 849 -968 0 3
rlabel polysilicon 856 -968 856 -968 0 3
rlabel polysilicon 859 -968 859 -968 0 4
rlabel polysilicon 863 -962 863 -962 0 1
rlabel polysilicon 863 -968 863 -968 0 3
rlabel polysilicon 870 -962 870 -962 0 1
rlabel polysilicon 870 -968 870 -968 0 3
rlabel polysilicon 877 -962 877 -962 0 1
rlabel polysilicon 877 -968 877 -968 0 3
rlabel polysilicon 884 -962 884 -962 0 1
rlabel polysilicon 884 -968 884 -968 0 3
rlabel polysilicon 891 -962 891 -962 0 1
rlabel polysilicon 891 -968 891 -968 0 3
rlabel polysilicon 898 -962 898 -962 0 1
rlabel polysilicon 898 -968 898 -968 0 3
rlabel polysilicon 905 -962 905 -962 0 1
rlabel polysilicon 905 -968 905 -968 0 3
rlabel polysilicon 912 -962 912 -962 0 1
rlabel polysilicon 912 -968 912 -968 0 3
rlabel polysilicon 919 -962 919 -962 0 1
rlabel polysilicon 919 -968 919 -968 0 3
rlabel polysilicon 926 -962 926 -962 0 1
rlabel polysilicon 926 -968 926 -968 0 3
rlabel polysilicon 933 -962 933 -962 0 1
rlabel polysilicon 933 -968 933 -968 0 3
rlabel polysilicon 940 -962 940 -962 0 1
rlabel polysilicon 940 -968 940 -968 0 3
rlabel polysilicon 947 -962 947 -962 0 1
rlabel polysilicon 947 -968 947 -968 0 3
rlabel polysilicon 954 -962 954 -962 0 1
rlabel polysilicon 954 -968 954 -968 0 3
rlabel polysilicon 961 -962 961 -962 0 1
rlabel polysilicon 961 -968 961 -968 0 3
rlabel polysilicon 968 -962 968 -962 0 1
rlabel polysilicon 968 -968 968 -968 0 3
rlabel polysilicon 975 -962 975 -962 0 1
rlabel polysilicon 975 -968 975 -968 0 3
rlabel polysilicon 982 -962 982 -962 0 1
rlabel polysilicon 982 -968 982 -968 0 3
rlabel polysilicon 989 -962 989 -962 0 1
rlabel polysilicon 989 -968 989 -968 0 3
rlabel polysilicon 996 -962 996 -962 0 1
rlabel polysilicon 996 -968 996 -968 0 3
rlabel polysilicon 1003 -962 1003 -962 0 1
rlabel polysilicon 1003 -968 1003 -968 0 3
rlabel polysilicon 1010 -962 1010 -962 0 1
rlabel polysilicon 1010 -968 1010 -968 0 3
rlabel polysilicon 1017 -962 1017 -962 0 1
rlabel polysilicon 1017 -968 1017 -968 0 3
rlabel polysilicon 1024 -962 1024 -962 0 1
rlabel polysilicon 1024 -968 1024 -968 0 3
rlabel polysilicon 1031 -962 1031 -962 0 1
rlabel polysilicon 1031 -968 1031 -968 0 3
rlabel polysilicon 1038 -962 1038 -962 0 1
rlabel polysilicon 1038 -968 1038 -968 0 3
rlabel polysilicon 1045 -962 1045 -962 0 1
rlabel polysilicon 1045 -968 1045 -968 0 3
rlabel polysilicon 1052 -962 1052 -962 0 1
rlabel polysilicon 1052 -968 1052 -968 0 3
rlabel polysilicon 1059 -962 1059 -962 0 1
rlabel polysilicon 1059 -968 1059 -968 0 3
rlabel polysilicon 1066 -962 1066 -962 0 1
rlabel polysilicon 1066 -968 1066 -968 0 3
rlabel polysilicon 1073 -962 1073 -962 0 1
rlabel polysilicon 1073 -968 1073 -968 0 3
rlabel polysilicon 1080 -962 1080 -962 0 1
rlabel polysilicon 1080 -968 1080 -968 0 3
rlabel polysilicon 1087 -962 1087 -962 0 1
rlabel polysilicon 1087 -968 1087 -968 0 3
rlabel polysilicon 1094 -962 1094 -962 0 1
rlabel polysilicon 1094 -968 1094 -968 0 3
rlabel polysilicon 1101 -962 1101 -962 0 1
rlabel polysilicon 1101 -968 1101 -968 0 3
rlabel polysilicon 1108 -962 1108 -962 0 1
rlabel polysilicon 1108 -968 1108 -968 0 3
rlabel polysilicon 1115 -962 1115 -962 0 1
rlabel polysilicon 1115 -968 1115 -968 0 3
rlabel polysilicon 1122 -962 1122 -962 0 1
rlabel polysilicon 1122 -968 1122 -968 0 3
rlabel polysilicon 1129 -962 1129 -962 0 1
rlabel polysilicon 1129 -968 1129 -968 0 3
rlabel polysilicon 1136 -962 1136 -962 0 1
rlabel polysilicon 1136 -968 1136 -968 0 3
rlabel polysilicon 1143 -962 1143 -962 0 1
rlabel polysilicon 1143 -968 1143 -968 0 3
rlabel polysilicon 1150 -962 1150 -962 0 1
rlabel polysilicon 1150 -968 1150 -968 0 3
rlabel polysilicon 1157 -962 1157 -962 0 1
rlabel polysilicon 1157 -968 1157 -968 0 3
rlabel polysilicon 2 -1077 2 -1077 0 1
rlabel polysilicon 9 -1077 9 -1077 0 1
rlabel polysilicon 9 -1083 9 -1083 0 3
rlabel polysilicon 16 -1077 16 -1077 0 1
rlabel polysilicon 16 -1083 16 -1083 0 3
rlabel polysilicon 23 -1077 23 -1077 0 1
rlabel polysilicon 23 -1083 23 -1083 0 3
rlabel polysilicon 30 -1077 30 -1077 0 1
rlabel polysilicon 30 -1083 30 -1083 0 3
rlabel polysilicon 37 -1077 37 -1077 0 1
rlabel polysilicon 37 -1083 37 -1083 0 3
rlabel polysilicon 44 -1077 44 -1077 0 1
rlabel polysilicon 44 -1083 44 -1083 0 3
rlabel polysilicon 51 -1077 51 -1077 0 1
rlabel polysilicon 51 -1083 51 -1083 0 3
rlabel polysilicon 54 -1083 54 -1083 0 4
rlabel polysilicon 58 -1077 58 -1077 0 1
rlabel polysilicon 58 -1083 58 -1083 0 3
rlabel polysilicon 68 -1077 68 -1077 0 2
rlabel polysilicon 65 -1083 65 -1083 0 3
rlabel polysilicon 68 -1083 68 -1083 0 4
rlabel polysilicon 72 -1077 72 -1077 0 1
rlabel polysilicon 72 -1083 72 -1083 0 3
rlabel polysilicon 82 -1077 82 -1077 0 2
rlabel polysilicon 79 -1083 79 -1083 0 3
rlabel polysilicon 86 -1077 86 -1077 0 1
rlabel polysilicon 86 -1083 86 -1083 0 3
rlabel polysilicon 93 -1077 93 -1077 0 1
rlabel polysilicon 93 -1083 93 -1083 0 3
rlabel polysilicon 100 -1083 100 -1083 0 3
rlabel polysilicon 103 -1083 103 -1083 0 4
rlabel polysilicon 107 -1077 107 -1077 0 1
rlabel polysilicon 110 -1083 110 -1083 0 4
rlabel polysilicon 114 -1077 114 -1077 0 1
rlabel polysilicon 114 -1083 114 -1083 0 3
rlabel polysilicon 121 -1077 121 -1077 0 1
rlabel polysilicon 121 -1083 121 -1083 0 3
rlabel polysilicon 128 -1077 128 -1077 0 1
rlabel polysilicon 128 -1083 128 -1083 0 3
rlabel polysilicon 135 -1077 135 -1077 0 1
rlabel polysilicon 135 -1083 135 -1083 0 3
rlabel polysilicon 142 -1077 142 -1077 0 1
rlabel polysilicon 142 -1083 142 -1083 0 3
rlabel polysilicon 149 -1077 149 -1077 0 1
rlabel polysilicon 149 -1083 149 -1083 0 3
rlabel polysilicon 156 -1077 156 -1077 0 1
rlabel polysilicon 156 -1083 156 -1083 0 3
rlabel polysilicon 163 -1077 163 -1077 0 1
rlabel polysilicon 166 -1077 166 -1077 0 2
rlabel polysilicon 166 -1083 166 -1083 0 4
rlabel polysilicon 170 -1077 170 -1077 0 1
rlabel polysilicon 170 -1083 170 -1083 0 3
rlabel polysilicon 177 -1077 177 -1077 0 1
rlabel polysilicon 177 -1083 177 -1083 0 3
rlabel polysilicon 184 -1077 184 -1077 0 1
rlabel polysilicon 184 -1083 184 -1083 0 3
rlabel polysilicon 191 -1077 191 -1077 0 1
rlabel polysilicon 194 -1077 194 -1077 0 2
rlabel polysilicon 191 -1083 191 -1083 0 3
rlabel polysilicon 198 -1077 198 -1077 0 1
rlabel polysilicon 198 -1083 198 -1083 0 3
rlabel polysilicon 205 -1077 205 -1077 0 1
rlabel polysilicon 205 -1083 205 -1083 0 3
rlabel polysilicon 212 -1083 212 -1083 0 3
rlabel polysilicon 215 -1083 215 -1083 0 4
rlabel polysilicon 219 -1077 219 -1077 0 1
rlabel polysilicon 219 -1083 219 -1083 0 3
rlabel polysilicon 229 -1077 229 -1077 0 2
rlabel polysilicon 226 -1083 226 -1083 0 3
rlabel polysilicon 233 -1077 233 -1077 0 1
rlabel polysilicon 233 -1083 233 -1083 0 3
rlabel polysilicon 240 -1077 240 -1077 0 1
rlabel polysilicon 240 -1083 240 -1083 0 3
rlabel polysilicon 247 -1077 247 -1077 0 1
rlabel polysilicon 247 -1083 247 -1083 0 3
rlabel polysilicon 254 -1077 254 -1077 0 1
rlabel polysilicon 254 -1083 254 -1083 0 3
rlabel polysilicon 261 -1077 261 -1077 0 1
rlabel polysilicon 261 -1083 261 -1083 0 3
rlabel polysilicon 268 -1077 268 -1077 0 1
rlabel polysilicon 271 -1077 271 -1077 0 2
rlabel polysilicon 275 -1077 275 -1077 0 1
rlabel polysilicon 275 -1083 275 -1083 0 3
rlabel polysilicon 282 -1077 282 -1077 0 1
rlabel polysilicon 285 -1083 285 -1083 0 4
rlabel polysilicon 289 -1077 289 -1077 0 1
rlabel polysilicon 289 -1083 289 -1083 0 3
rlabel polysilicon 296 -1077 296 -1077 0 1
rlabel polysilicon 296 -1083 296 -1083 0 3
rlabel polysilicon 303 -1077 303 -1077 0 1
rlabel polysilicon 303 -1083 303 -1083 0 3
rlabel polysilicon 310 -1077 310 -1077 0 1
rlabel polysilicon 310 -1083 310 -1083 0 3
rlabel polysilicon 317 -1077 317 -1077 0 1
rlabel polysilicon 317 -1083 317 -1083 0 3
rlabel polysilicon 324 -1077 324 -1077 0 1
rlabel polysilicon 324 -1083 324 -1083 0 3
rlabel polysilicon 331 -1077 331 -1077 0 1
rlabel polysilicon 331 -1083 331 -1083 0 3
rlabel polysilicon 338 -1077 338 -1077 0 1
rlabel polysilicon 338 -1083 338 -1083 0 3
rlabel polysilicon 345 -1077 345 -1077 0 1
rlabel polysilicon 345 -1083 345 -1083 0 3
rlabel polysilicon 352 -1077 352 -1077 0 1
rlabel polysilicon 352 -1083 352 -1083 0 3
rlabel polysilicon 359 -1077 359 -1077 0 1
rlabel polysilicon 359 -1083 359 -1083 0 3
rlabel polysilicon 366 -1077 366 -1077 0 1
rlabel polysilicon 366 -1083 366 -1083 0 3
rlabel polysilicon 373 -1077 373 -1077 0 1
rlabel polysilicon 373 -1083 373 -1083 0 3
rlabel polysilicon 380 -1077 380 -1077 0 1
rlabel polysilicon 380 -1083 380 -1083 0 3
rlabel polysilicon 387 -1077 387 -1077 0 1
rlabel polysilicon 390 -1077 390 -1077 0 2
rlabel polysilicon 387 -1083 387 -1083 0 3
rlabel polysilicon 390 -1083 390 -1083 0 4
rlabel polysilicon 394 -1077 394 -1077 0 1
rlabel polysilicon 397 -1077 397 -1077 0 2
rlabel polysilicon 394 -1083 394 -1083 0 3
rlabel polysilicon 397 -1083 397 -1083 0 4
rlabel polysilicon 401 -1077 401 -1077 0 1
rlabel polysilicon 401 -1083 401 -1083 0 3
rlabel polysilicon 408 -1077 408 -1077 0 1
rlabel polysilicon 408 -1083 408 -1083 0 3
rlabel polysilicon 415 -1077 415 -1077 0 1
rlabel polysilicon 415 -1083 415 -1083 0 3
rlabel polysilicon 422 -1077 422 -1077 0 1
rlabel polysilicon 422 -1083 422 -1083 0 3
rlabel polysilicon 429 -1077 429 -1077 0 1
rlabel polysilicon 429 -1083 429 -1083 0 3
rlabel polysilicon 436 -1077 436 -1077 0 1
rlabel polysilicon 436 -1083 436 -1083 0 3
rlabel polysilicon 443 -1077 443 -1077 0 1
rlabel polysilicon 443 -1083 443 -1083 0 3
rlabel polysilicon 450 -1077 450 -1077 0 1
rlabel polysilicon 450 -1083 450 -1083 0 3
rlabel polysilicon 457 -1077 457 -1077 0 1
rlabel polysilicon 457 -1083 457 -1083 0 3
rlabel polysilicon 464 -1077 464 -1077 0 1
rlabel polysilicon 464 -1083 464 -1083 0 3
rlabel polysilicon 471 -1077 471 -1077 0 1
rlabel polysilicon 471 -1083 471 -1083 0 3
rlabel polysilicon 478 -1077 478 -1077 0 1
rlabel polysilicon 478 -1083 478 -1083 0 3
rlabel polysilicon 488 -1077 488 -1077 0 2
rlabel polysilicon 485 -1083 485 -1083 0 3
rlabel polysilicon 488 -1083 488 -1083 0 4
rlabel polysilicon 492 -1077 492 -1077 0 1
rlabel polysilicon 495 -1077 495 -1077 0 2
rlabel polysilicon 495 -1083 495 -1083 0 4
rlabel polysilicon 502 -1077 502 -1077 0 2
rlabel polysilicon 499 -1083 499 -1083 0 3
rlabel polysilicon 502 -1083 502 -1083 0 4
rlabel polysilicon 506 -1077 506 -1077 0 1
rlabel polysilicon 506 -1083 506 -1083 0 3
rlabel polysilicon 513 -1077 513 -1077 0 1
rlabel polysilicon 513 -1083 513 -1083 0 3
rlabel polysilicon 520 -1077 520 -1077 0 1
rlabel polysilicon 520 -1083 520 -1083 0 3
rlabel polysilicon 527 -1077 527 -1077 0 1
rlabel polysilicon 527 -1083 527 -1083 0 3
rlabel polysilicon 534 -1077 534 -1077 0 1
rlabel polysilicon 534 -1083 534 -1083 0 3
rlabel polysilicon 541 -1077 541 -1077 0 1
rlabel polysilicon 541 -1083 541 -1083 0 3
rlabel polysilicon 544 -1083 544 -1083 0 4
rlabel polysilicon 548 -1077 548 -1077 0 1
rlabel polysilicon 548 -1083 548 -1083 0 3
rlabel polysilicon 555 -1077 555 -1077 0 1
rlabel polysilicon 558 -1077 558 -1077 0 2
rlabel polysilicon 555 -1083 555 -1083 0 3
rlabel polysilicon 558 -1083 558 -1083 0 4
rlabel polysilicon 562 -1077 562 -1077 0 1
rlabel polysilicon 562 -1083 562 -1083 0 3
rlabel polysilicon 569 -1077 569 -1077 0 1
rlabel polysilicon 572 -1077 572 -1077 0 2
rlabel polysilicon 572 -1083 572 -1083 0 4
rlabel polysilicon 576 -1077 576 -1077 0 1
rlabel polysilicon 576 -1083 576 -1083 0 3
rlabel polysilicon 583 -1077 583 -1077 0 1
rlabel polysilicon 583 -1083 583 -1083 0 3
rlabel polysilicon 586 -1083 586 -1083 0 4
rlabel polysilicon 590 -1077 590 -1077 0 1
rlabel polysilicon 590 -1083 590 -1083 0 3
rlabel polysilicon 600 -1077 600 -1077 0 2
rlabel polysilicon 597 -1083 597 -1083 0 3
rlabel polysilicon 604 -1077 604 -1077 0 1
rlabel polysilicon 607 -1077 607 -1077 0 2
rlabel polysilicon 604 -1083 604 -1083 0 3
rlabel polysilicon 607 -1083 607 -1083 0 4
rlabel polysilicon 611 -1077 611 -1077 0 1
rlabel polysilicon 611 -1083 611 -1083 0 3
rlabel polysilicon 618 -1077 618 -1077 0 1
rlabel polysilicon 618 -1083 618 -1083 0 3
rlabel polysilicon 625 -1077 625 -1077 0 1
rlabel polysilicon 625 -1083 625 -1083 0 3
rlabel polysilicon 632 -1077 632 -1077 0 1
rlabel polysilicon 635 -1077 635 -1077 0 2
rlabel polysilicon 632 -1083 632 -1083 0 3
rlabel polysilicon 635 -1083 635 -1083 0 4
rlabel polysilicon 639 -1077 639 -1077 0 1
rlabel polysilicon 639 -1083 639 -1083 0 3
rlabel polysilicon 646 -1077 646 -1077 0 1
rlabel polysilicon 646 -1083 646 -1083 0 3
rlabel polysilicon 653 -1077 653 -1077 0 1
rlabel polysilicon 653 -1083 653 -1083 0 3
rlabel polysilicon 660 -1077 660 -1077 0 1
rlabel polysilicon 660 -1083 660 -1083 0 3
rlabel polysilicon 667 -1077 667 -1077 0 1
rlabel polysilicon 667 -1083 667 -1083 0 3
rlabel polysilicon 674 -1077 674 -1077 0 1
rlabel polysilicon 674 -1083 674 -1083 0 3
rlabel polysilicon 681 -1077 681 -1077 0 1
rlabel polysilicon 681 -1083 681 -1083 0 3
rlabel polysilicon 684 -1083 684 -1083 0 4
rlabel polysilicon 688 -1077 688 -1077 0 1
rlabel polysilicon 688 -1083 688 -1083 0 3
rlabel polysilicon 695 -1077 695 -1077 0 1
rlabel polysilicon 695 -1083 695 -1083 0 3
rlabel polysilicon 702 -1077 702 -1077 0 1
rlabel polysilicon 702 -1083 702 -1083 0 3
rlabel polysilicon 709 -1077 709 -1077 0 1
rlabel polysilicon 709 -1083 709 -1083 0 3
rlabel polysilicon 716 -1077 716 -1077 0 1
rlabel polysilicon 716 -1083 716 -1083 0 3
rlabel polysilicon 723 -1077 723 -1077 0 1
rlabel polysilicon 726 -1077 726 -1077 0 2
rlabel polysilicon 730 -1077 730 -1077 0 1
rlabel polysilicon 730 -1083 730 -1083 0 3
rlabel polysilicon 737 -1077 737 -1077 0 1
rlabel polysilicon 740 -1077 740 -1077 0 2
rlabel polysilicon 737 -1083 737 -1083 0 3
rlabel polysilicon 744 -1077 744 -1077 0 1
rlabel polysilicon 744 -1083 744 -1083 0 3
rlabel polysilicon 751 -1077 751 -1077 0 1
rlabel polysilicon 751 -1083 751 -1083 0 3
rlabel polysilicon 758 -1077 758 -1077 0 1
rlabel polysilicon 758 -1083 758 -1083 0 3
rlabel polysilicon 765 -1077 765 -1077 0 1
rlabel polysilicon 765 -1083 765 -1083 0 3
rlabel polysilicon 772 -1077 772 -1077 0 1
rlabel polysilicon 772 -1083 772 -1083 0 3
rlabel polysilicon 779 -1077 779 -1077 0 1
rlabel polysilicon 779 -1083 779 -1083 0 3
rlabel polysilicon 786 -1077 786 -1077 0 1
rlabel polysilicon 786 -1083 786 -1083 0 3
rlabel polysilicon 793 -1077 793 -1077 0 1
rlabel polysilicon 793 -1083 793 -1083 0 3
rlabel polysilicon 800 -1077 800 -1077 0 1
rlabel polysilicon 800 -1083 800 -1083 0 3
rlabel polysilicon 807 -1077 807 -1077 0 1
rlabel polysilicon 807 -1083 807 -1083 0 3
rlabel polysilicon 814 -1083 814 -1083 0 3
rlabel polysilicon 817 -1083 817 -1083 0 4
rlabel polysilicon 821 -1077 821 -1077 0 1
rlabel polysilicon 821 -1083 821 -1083 0 3
rlabel polysilicon 828 -1077 828 -1077 0 1
rlabel polysilicon 828 -1083 828 -1083 0 3
rlabel polysilicon 835 -1077 835 -1077 0 1
rlabel polysilicon 835 -1083 835 -1083 0 3
rlabel polysilicon 842 -1077 842 -1077 0 1
rlabel polysilicon 842 -1083 842 -1083 0 3
rlabel polysilicon 849 -1077 849 -1077 0 1
rlabel polysilicon 849 -1083 849 -1083 0 3
rlabel polysilicon 856 -1077 856 -1077 0 1
rlabel polysilicon 856 -1083 856 -1083 0 3
rlabel polysilicon 863 -1077 863 -1077 0 1
rlabel polysilicon 863 -1083 863 -1083 0 3
rlabel polysilicon 870 -1077 870 -1077 0 1
rlabel polysilicon 870 -1083 870 -1083 0 3
rlabel polysilicon 877 -1077 877 -1077 0 1
rlabel polysilicon 877 -1083 877 -1083 0 3
rlabel polysilicon 884 -1077 884 -1077 0 1
rlabel polysilicon 884 -1083 884 -1083 0 3
rlabel polysilicon 891 -1077 891 -1077 0 1
rlabel polysilicon 891 -1083 891 -1083 0 3
rlabel polysilicon 898 -1077 898 -1077 0 1
rlabel polysilicon 898 -1083 898 -1083 0 3
rlabel polysilicon 905 -1077 905 -1077 0 1
rlabel polysilicon 905 -1083 905 -1083 0 3
rlabel polysilicon 912 -1077 912 -1077 0 1
rlabel polysilicon 912 -1083 912 -1083 0 3
rlabel polysilicon 919 -1077 919 -1077 0 1
rlabel polysilicon 919 -1083 919 -1083 0 3
rlabel polysilicon 926 -1077 926 -1077 0 1
rlabel polysilicon 926 -1083 926 -1083 0 3
rlabel polysilicon 933 -1077 933 -1077 0 1
rlabel polysilicon 933 -1083 933 -1083 0 3
rlabel polysilicon 940 -1077 940 -1077 0 1
rlabel polysilicon 940 -1083 940 -1083 0 3
rlabel polysilicon 947 -1077 947 -1077 0 1
rlabel polysilicon 947 -1083 947 -1083 0 3
rlabel polysilicon 954 -1077 954 -1077 0 1
rlabel polysilicon 954 -1083 954 -1083 0 3
rlabel polysilicon 961 -1077 961 -1077 0 1
rlabel polysilicon 961 -1083 961 -1083 0 3
rlabel polysilicon 968 -1077 968 -1077 0 1
rlabel polysilicon 968 -1083 968 -1083 0 3
rlabel polysilicon 975 -1077 975 -1077 0 1
rlabel polysilicon 975 -1083 975 -1083 0 3
rlabel polysilicon 982 -1077 982 -1077 0 1
rlabel polysilicon 982 -1083 982 -1083 0 3
rlabel polysilicon 989 -1077 989 -1077 0 1
rlabel polysilicon 989 -1083 989 -1083 0 3
rlabel polysilicon 996 -1077 996 -1077 0 1
rlabel polysilicon 996 -1083 996 -1083 0 3
rlabel polysilicon 1003 -1077 1003 -1077 0 1
rlabel polysilicon 1003 -1083 1003 -1083 0 3
rlabel polysilicon 1010 -1077 1010 -1077 0 1
rlabel polysilicon 1010 -1083 1010 -1083 0 3
rlabel polysilicon 1017 -1077 1017 -1077 0 1
rlabel polysilicon 1017 -1083 1017 -1083 0 3
rlabel polysilicon 1024 -1077 1024 -1077 0 1
rlabel polysilicon 1024 -1083 1024 -1083 0 3
rlabel polysilicon 1031 -1077 1031 -1077 0 1
rlabel polysilicon 1031 -1083 1031 -1083 0 3
rlabel polysilicon 1041 -1077 1041 -1077 0 2
rlabel polysilicon 1038 -1083 1038 -1083 0 3
rlabel polysilicon 1041 -1083 1041 -1083 0 4
rlabel polysilicon 1045 -1077 1045 -1077 0 1
rlabel polysilicon 1045 -1083 1045 -1083 0 3
rlabel polysilicon 1052 -1077 1052 -1077 0 1
rlabel polysilicon 1052 -1083 1052 -1083 0 3
rlabel polysilicon 1059 -1083 1059 -1083 0 3
rlabel polysilicon 1066 -1077 1066 -1077 0 1
rlabel polysilicon 1066 -1083 1066 -1083 0 3
rlabel polysilicon 1073 -1077 1073 -1077 0 1
rlabel polysilicon 1073 -1083 1073 -1083 0 3
rlabel polysilicon 1080 -1077 1080 -1077 0 1
rlabel polysilicon 1080 -1083 1080 -1083 0 3
rlabel polysilicon 1129 -1077 1129 -1077 0 1
rlabel polysilicon 1129 -1083 1129 -1083 0 3
rlabel polysilicon 1143 -1077 1143 -1077 0 1
rlabel polysilicon 1143 -1083 1143 -1083 0 3
rlabel polysilicon 5 -1166 5 -1166 0 2
rlabel polysilicon 9 -1166 9 -1166 0 1
rlabel polysilicon 9 -1172 9 -1172 0 3
rlabel polysilicon 16 -1172 16 -1172 0 3
rlabel polysilicon 19 -1172 19 -1172 0 4
rlabel polysilicon 23 -1166 23 -1166 0 1
rlabel polysilicon 23 -1172 23 -1172 0 3
rlabel polysilicon 30 -1166 30 -1166 0 1
rlabel polysilicon 30 -1172 30 -1172 0 3
rlabel polysilicon 37 -1166 37 -1166 0 1
rlabel polysilicon 40 -1166 40 -1166 0 2
rlabel polysilicon 37 -1172 37 -1172 0 3
rlabel polysilicon 44 -1166 44 -1166 0 1
rlabel polysilicon 44 -1172 44 -1172 0 3
rlabel polysilicon 51 -1166 51 -1166 0 1
rlabel polysilicon 51 -1172 51 -1172 0 3
rlabel polysilicon 61 -1166 61 -1166 0 2
rlabel polysilicon 58 -1172 58 -1172 0 3
rlabel polysilicon 61 -1172 61 -1172 0 4
rlabel polysilicon 65 -1166 65 -1166 0 1
rlabel polysilicon 65 -1172 65 -1172 0 3
rlabel polysilicon 72 -1166 72 -1166 0 1
rlabel polysilicon 72 -1172 72 -1172 0 3
rlabel polysilicon 79 -1166 79 -1166 0 1
rlabel polysilicon 79 -1172 79 -1172 0 3
rlabel polysilicon 86 -1166 86 -1166 0 1
rlabel polysilicon 86 -1172 86 -1172 0 3
rlabel polysilicon 93 -1166 93 -1166 0 1
rlabel polysilicon 93 -1172 93 -1172 0 3
rlabel polysilicon 100 -1166 100 -1166 0 1
rlabel polysilicon 100 -1172 100 -1172 0 3
rlabel polysilicon 107 -1166 107 -1166 0 1
rlabel polysilicon 107 -1172 107 -1172 0 3
rlabel polysilicon 114 -1166 114 -1166 0 1
rlabel polysilicon 114 -1172 114 -1172 0 3
rlabel polysilicon 121 -1166 121 -1166 0 1
rlabel polysilicon 121 -1172 121 -1172 0 3
rlabel polysilicon 128 -1166 128 -1166 0 1
rlabel polysilicon 128 -1172 128 -1172 0 3
rlabel polysilicon 135 -1166 135 -1166 0 1
rlabel polysilicon 135 -1172 135 -1172 0 3
rlabel polysilicon 142 -1172 142 -1172 0 3
rlabel polysilicon 145 -1172 145 -1172 0 4
rlabel polysilicon 152 -1166 152 -1166 0 2
rlabel polysilicon 152 -1172 152 -1172 0 4
rlabel polysilicon 156 -1166 156 -1166 0 1
rlabel polysilicon 156 -1172 156 -1172 0 3
rlabel polysilicon 163 -1166 163 -1166 0 1
rlabel polysilicon 163 -1172 163 -1172 0 3
rlabel polysilicon 170 -1166 170 -1166 0 1
rlabel polysilicon 170 -1172 170 -1172 0 3
rlabel polysilicon 177 -1166 177 -1166 0 1
rlabel polysilicon 177 -1172 177 -1172 0 3
rlabel polysilicon 184 -1166 184 -1166 0 1
rlabel polysilicon 184 -1172 184 -1172 0 3
rlabel polysilicon 191 -1166 191 -1166 0 1
rlabel polysilicon 191 -1172 191 -1172 0 3
rlabel polysilicon 198 -1166 198 -1166 0 1
rlabel polysilicon 198 -1172 198 -1172 0 3
rlabel polysilicon 205 -1166 205 -1166 0 1
rlabel polysilicon 205 -1172 205 -1172 0 3
rlabel polysilicon 212 -1166 212 -1166 0 1
rlabel polysilicon 212 -1172 212 -1172 0 3
rlabel polysilicon 219 -1166 219 -1166 0 1
rlabel polysilicon 222 -1172 222 -1172 0 4
rlabel polysilicon 226 -1166 226 -1166 0 1
rlabel polysilicon 226 -1172 226 -1172 0 3
rlabel polysilicon 233 -1166 233 -1166 0 1
rlabel polysilicon 233 -1172 233 -1172 0 3
rlabel polysilicon 240 -1166 240 -1166 0 1
rlabel polysilicon 240 -1172 240 -1172 0 3
rlabel polysilicon 247 -1166 247 -1166 0 1
rlabel polysilicon 247 -1172 247 -1172 0 3
rlabel polysilicon 254 -1166 254 -1166 0 1
rlabel polysilicon 254 -1172 254 -1172 0 3
rlabel polysilicon 261 -1166 261 -1166 0 1
rlabel polysilicon 261 -1172 261 -1172 0 3
rlabel polysilicon 268 -1166 268 -1166 0 1
rlabel polysilicon 268 -1172 268 -1172 0 3
rlabel polysilicon 275 -1166 275 -1166 0 1
rlabel polysilicon 275 -1172 275 -1172 0 3
rlabel polysilicon 282 -1166 282 -1166 0 1
rlabel polysilicon 282 -1172 282 -1172 0 3
rlabel polysilicon 285 -1172 285 -1172 0 4
rlabel polysilicon 289 -1166 289 -1166 0 1
rlabel polysilicon 289 -1172 289 -1172 0 3
rlabel polysilicon 296 -1166 296 -1166 0 1
rlabel polysilicon 296 -1172 296 -1172 0 3
rlabel polysilicon 303 -1166 303 -1166 0 1
rlabel polysilicon 303 -1172 303 -1172 0 3
rlabel polysilicon 313 -1166 313 -1166 0 2
rlabel polysilicon 310 -1172 310 -1172 0 3
rlabel polysilicon 313 -1172 313 -1172 0 4
rlabel polysilicon 317 -1166 317 -1166 0 1
rlabel polysilicon 317 -1172 317 -1172 0 3
rlabel polysilicon 324 -1166 324 -1166 0 1
rlabel polysilicon 324 -1172 324 -1172 0 3
rlabel polysilicon 331 -1166 331 -1166 0 1
rlabel polysilicon 331 -1172 331 -1172 0 3
rlabel polysilicon 338 -1166 338 -1166 0 1
rlabel polysilicon 338 -1172 338 -1172 0 3
rlabel polysilicon 345 -1166 345 -1166 0 1
rlabel polysilicon 348 -1166 348 -1166 0 2
rlabel polysilicon 345 -1172 345 -1172 0 3
rlabel polysilicon 348 -1172 348 -1172 0 4
rlabel polysilicon 352 -1166 352 -1166 0 1
rlabel polysilicon 355 -1166 355 -1166 0 2
rlabel polysilicon 352 -1172 352 -1172 0 3
rlabel polysilicon 355 -1172 355 -1172 0 4
rlabel polysilicon 359 -1172 359 -1172 0 3
rlabel polysilicon 362 -1172 362 -1172 0 4
rlabel polysilicon 366 -1166 366 -1166 0 1
rlabel polysilicon 366 -1172 366 -1172 0 3
rlabel polysilicon 373 -1166 373 -1166 0 1
rlabel polysilicon 373 -1172 373 -1172 0 3
rlabel polysilicon 380 -1166 380 -1166 0 1
rlabel polysilicon 383 -1166 383 -1166 0 2
rlabel polysilicon 380 -1172 380 -1172 0 3
rlabel polysilicon 383 -1172 383 -1172 0 4
rlabel polysilicon 387 -1166 387 -1166 0 1
rlabel polysilicon 387 -1172 387 -1172 0 3
rlabel polysilicon 394 -1166 394 -1166 0 1
rlabel polysilicon 394 -1172 394 -1172 0 3
rlabel polysilicon 401 -1166 401 -1166 0 1
rlabel polysilicon 401 -1172 401 -1172 0 3
rlabel polysilicon 408 -1166 408 -1166 0 1
rlabel polysilicon 411 -1166 411 -1166 0 2
rlabel polysilicon 415 -1166 415 -1166 0 1
rlabel polysilicon 418 -1166 418 -1166 0 2
rlabel polysilicon 415 -1172 415 -1172 0 3
rlabel polysilicon 418 -1172 418 -1172 0 4
rlabel polysilicon 422 -1166 422 -1166 0 1
rlabel polysilicon 422 -1172 422 -1172 0 3
rlabel polysilicon 429 -1166 429 -1166 0 1
rlabel polysilicon 429 -1172 429 -1172 0 3
rlabel polysilicon 436 -1166 436 -1166 0 1
rlabel polysilicon 436 -1172 436 -1172 0 3
rlabel polysilicon 443 -1166 443 -1166 0 1
rlabel polysilicon 443 -1172 443 -1172 0 3
rlabel polysilicon 450 -1166 450 -1166 0 1
rlabel polysilicon 450 -1172 450 -1172 0 3
rlabel polysilicon 457 -1166 457 -1166 0 1
rlabel polysilicon 457 -1172 457 -1172 0 3
rlabel polysilicon 464 -1166 464 -1166 0 1
rlabel polysilicon 467 -1166 467 -1166 0 2
rlabel polysilicon 464 -1172 464 -1172 0 3
rlabel polysilicon 467 -1172 467 -1172 0 4
rlabel polysilicon 471 -1166 471 -1166 0 1
rlabel polysilicon 471 -1172 471 -1172 0 3
rlabel polysilicon 481 -1166 481 -1166 0 2
rlabel polysilicon 478 -1172 478 -1172 0 3
rlabel polysilicon 481 -1172 481 -1172 0 4
rlabel polysilicon 485 -1166 485 -1166 0 1
rlabel polysilicon 485 -1172 485 -1172 0 3
rlabel polysilicon 492 -1166 492 -1166 0 1
rlabel polysilicon 492 -1172 492 -1172 0 3
rlabel polysilicon 499 -1166 499 -1166 0 1
rlabel polysilicon 502 -1166 502 -1166 0 2
rlabel polysilicon 499 -1172 499 -1172 0 3
rlabel polysilicon 502 -1172 502 -1172 0 4
rlabel polysilicon 506 -1166 506 -1166 0 1
rlabel polysilicon 506 -1172 506 -1172 0 3
rlabel polysilicon 513 -1166 513 -1166 0 1
rlabel polysilicon 513 -1172 513 -1172 0 3
rlabel polysilicon 520 -1166 520 -1166 0 1
rlabel polysilicon 523 -1166 523 -1166 0 2
rlabel polysilicon 523 -1172 523 -1172 0 4
rlabel polysilicon 527 -1166 527 -1166 0 1
rlabel polysilicon 527 -1172 527 -1172 0 3
rlabel polysilicon 534 -1166 534 -1166 0 1
rlabel polysilicon 534 -1172 534 -1172 0 3
rlabel polysilicon 541 -1166 541 -1166 0 1
rlabel polysilicon 541 -1172 541 -1172 0 3
rlabel polysilicon 548 -1166 548 -1166 0 1
rlabel polysilicon 548 -1172 548 -1172 0 3
rlabel polysilicon 555 -1166 555 -1166 0 1
rlabel polysilicon 558 -1166 558 -1166 0 2
rlabel polysilicon 555 -1172 555 -1172 0 3
rlabel polysilicon 558 -1172 558 -1172 0 4
rlabel polysilicon 565 -1166 565 -1166 0 2
rlabel polysilicon 562 -1172 562 -1172 0 3
rlabel polysilicon 569 -1166 569 -1166 0 1
rlabel polysilicon 569 -1172 569 -1172 0 3
rlabel polysilicon 576 -1166 576 -1166 0 1
rlabel polysilicon 576 -1172 576 -1172 0 3
rlabel polysilicon 583 -1166 583 -1166 0 1
rlabel polysilicon 583 -1172 583 -1172 0 3
rlabel polysilicon 590 -1166 590 -1166 0 1
rlabel polysilicon 590 -1172 590 -1172 0 3
rlabel polysilicon 597 -1172 597 -1172 0 3
rlabel polysilicon 600 -1172 600 -1172 0 4
rlabel polysilicon 604 -1166 604 -1166 0 1
rlabel polysilicon 604 -1172 604 -1172 0 3
rlabel polysilicon 611 -1166 611 -1166 0 1
rlabel polysilicon 611 -1172 611 -1172 0 3
rlabel polysilicon 618 -1166 618 -1166 0 1
rlabel polysilicon 618 -1172 618 -1172 0 3
rlabel polysilicon 625 -1166 625 -1166 0 1
rlabel polysilicon 625 -1172 625 -1172 0 3
rlabel polysilicon 632 -1166 632 -1166 0 1
rlabel polysilicon 632 -1172 632 -1172 0 3
rlabel polysilicon 639 -1166 639 -1166 0 1
rlabel polysilicon 639 -1172 639 -1172 0 3
rlabel polysilicon 646 -1166 646 -1166 0 1
rlabel polysilicon 646 -1172 646 -1172 0 3
rlabel polysilicon 653 -1166 653 -1166 0 1
rlabel polysilicon 653 -1172 653 -1172 0 3
rlabel polysilicon 660 -1166 660 -1166 0 1
rlabel polysilicon 660 -1172 660 -1172 0 3
rlabel polysilicon 667 -1166 667 -1166 0 1
rlabel polysilicon 667 -1172 667 -1172 0 3
rlabel polysilicon 674 -1166 674 -1166 0 1
rlabel polysilicon 674 -1172 674 -1172 0 3
rlabel polysilicon 681 -1166 681 -1166 0 1
rlabel polysilicon 681 -1172 681 -1172 0 3
rlabel polysilicon 691 -1166 691 -1166 0 2
rlabel polysilicon 688 -1172 688 -1172 0 3
rlabel polysilicon 695 -1166 695 -1166 0 1
rlabel polysilicon 695 -1172 695 -1172 0 3
rlabel polysilicon 702 -1166 702 -1166 0 1
rlabel polysilicon 702 -1172 702 -1172 0 3
rlabel polysilicon 709 -1166 709 -1166 0 1
rlabel polysilicon 709 -1172 709 -1172 0 3
rlabel polysilicon 716 -1166 716 -1166 0 1
rlabel polysilicon 716 -1172 716 -1172 0 3
rlabel polysilicon 723 -1166 723 -1166 0 1
rlabel polysilicon 723 -1172 723 -1172 0 3
rlabel polysilicon 730 -1166 730 -1166 0 1
rlabel polysilicon 733 -1166 733 -1166 0 2
rlabel polysilicon 730 -1172 730 -1172 0 3
rlabel polysilicon 733 -1172 733 -1172 0 4
rlabel polysilicon 740 -1166 740 -1166 0 2
rlabel polysilicon 737 -1172 737 -1172 0 3
rlabel polysilicon 744 -1166 744 -1166 0 1
rlabel polysilicon 744 -1172 744 -1172 0 3
rlabel polysilicon 751 -1166 751 -1166 0 1
rlabel polysilicon 751 -1172 751 -1172 0 3
rlabel polysilicon 758 -1166 758 -1166 0 1
rlabel polysilicon 758 -1172 758 -1172 0 3
rlabel polysilicon 765 -1166 765 -1166 0 1
rlabel polysilicon 765 -1172 765 -1172 0 3
rlabel polysilicon 772 -1166 772 -1166 0 1
rlabel polysilicon 772 -1172 772 -1172 0 3
rlabel polysilicon 779 -1166 779 -1166 0 1
rlabel polysilicon 779 -1172 779 -1172 0 3
rlabel polysilicon 786 -1166 786 -1166 0 1
rlabel polysilicon 789 -1166 789 -1166 0 2
rlabel polysilicon 786 -1172 786 -1172 0 3
rlabel polysilicon 789 -1172 789 -1172 0 4
rlabel polysilicon 793 -1166 793 -1166 0 1
rlabel polysilicon 793 -1172 793 -1172 0 3
rlabel polysilicon 800 -1166 800 -1166 0 1
rlabel polysilicon 800 -1172 800 -1172 0 3
rlabel polysilicon 807 -1166 807 -1166 0 1
rlabel polysilicon 807 -1172 807 -1172 0 3
rlabel polysilicon 814 -1166 814 -1166 0 1
rlabel polysilicon 814 -1172 814 -1172 0 3
rlabel polysilicon 821 -1166 821 -1166 0 1
rlabel polysilicon 821 -1172 821 -1172 0 3
rlabel polysilicon 828 -1166 828 -1166 0 1
rlabel polysilicon 828 -1172 828 -1172 0 3
rlabel polysilicon 835 -1166 835 -1166 0 1
rlabel polysilicon 835 -1172 835 -1172 0 3
rlabel polysilicon 842 -1166 842 -1166 0 1
rlabel polysilicon 842 -1172 842 -1172 0 3
rlabel polysilicon 849 -1166 849 -1166 0 1
rlabel polysilicon 849 -1172 849 -1172 0 3
rlabel polysilicon 856 -1166 856 -1166 0 1
rlabel polysilicon 859 -1172 859 -1172 0 4
rlabel polysilicon 863 -1166 863 -1166 0 1
rlabel polysilicon 863 -1172 863 -1172 0 3
rlabel polysilicon 870 -1166 870 -1166 0 1
rlabel polysilicon 870 -1172 870 -1172 0 3
rlabel polysilicon 877 -1166 877 -1166 0 1
rlabel polysilicon 877 -1172 877 -1172 0 3
rlabel polysilicon 884 -1166 884 -1166 0 1
rlabel polysilicon 884 -1172 884 -1172 0 3
rlabel polysilicon 891 -1166 891 -1166 0 1
rlabel polysilicon 891 -1172 891 -1172 0 3
rlabel polysilicon 898 -1166 898 -1166 0 1
rlabel polysilicon 898 -1172 898 -1172 0 3
rlabel polysilicon 905 -1166 905 -1166 0 1
rlabel polysilicon 905 -1172 905 -1172 0 3
rlabel polysilicon 912 -1166 912 -1166 0 1
rlabel polysilicon 912 -1172 912 -1172 0 3
rlabel polysilicon 919 -1166 919 -1166 0 1
rlabel polysilicon 919 -1172 919 -1172 0 3
rlabel polysilicon 926 -1166 926 -1166 0 1
rlabel polysilicon 926 -1172 926 -1172 0 3
rlabel polysilicon 933 -1166 933 -1166 0 1
rlabel polysilicon 933 -1172 933 -1172 0 3
rlabel polysilicon 940 -1166 940 -1166 0 1
rlabel polysilicon 940 -1172 940 -1172 0 3
rlabel polysilicon 947 -1166 947 -1166 0 1
rlabel polysilicon 947 -1172 947 -1172 0 3
rlabel polysilicon 954 -1166 954 -1166 0 1
rlabel polysilicon 954 -1172 954 -1172 0 3
rlabel polysilicon 961 -1166 961 -1166 0 1
rlabel polysilicon 961 -1172 961 -1172 0 3
rlabel polysilicon 968 -1166 968 -1166 0 1
rlabel polysilicon 968 -1172 968 -1172 0 3
rlabel polysilicon 975 -1166 975 -1166 0 1
rlabel polysilicon 975 -1172 975 -1172 0 3
rlabel polysilicon 982 -1166 982 -1166 0 1
rlabel polysilicon 982 -1172 982 -1172 0 3
rlabel polysilicon 989 -1166 989 -1166 0 1
rlabel polysilicon 989 -1172 989 -1172 0 3
rlabel polysilicon 996 -1166 996 -1166 0 1
rlabel polysilicon 996 -1172 996 -1172 0 3
rlabel polysilicon 1003 -1166 1003 -1166 0 1
rlabel polysilicon 1003 -1172 1003 -1172 0 3
rlabel polysilicon 1010 -1166 1010 -1166 0 1
rlabel polysilicon 1010 -1172 1010 -1172 0 3
rlabel polysilicon 1017 -1166 1017 -1166 0 1
rlabel polysilicon 1017 -1172 1017 -1172 0 3
rlabel polysilicon 1024 -1166 1024 -1166 0 1
rlabel polysilicon 1024 -1172 1024 -1172 0 3
rlabel polysilicon 1031 -1166 1031 -1166 0 1
rlabel polysilicon 1031 -1172 1031 -1172 0 3
rlabel polysilicon 1038 -1166 1038 -1166 0 1
rlabel polysilicon 1041 -1166 1041 -1166 0 2
rlabel polysilicon 1038 -1172 1038 -1172 0 3
rlabel polysilicon 1041 -1172 1041 -1172 0 4
rlabel polysilicon 1045 -1166 1045 -1166 0 1
rlabel polysilicon 1045 -1172 1045 -1172 0 3
rlabel polysilicon 1052 -1166 1052 -1166 0 1
rlabel polysilicon 1052 -1172 1052 -1172 0 3
rlabel polysilicon 1059 -1166 1059 -1166 0 1
rlabel polysilicon 1059 -1172 1059 -1172 0 3
rlabel polysilicon 1066 -1166 1066 -1166 0 1
rlabel polysilicon 1066 -1172 1066 -1172 0 3
rlabel polysilicon 1073 -1166 1073 -1166 0 1
rlabel polysilicon 1076 -1166 1076 -1166 0 2
rlabel polysilicon 1122 -1166 1122 -1166 0 1
rlabel polysilicon 1122 -1172 1122 -1172 0 3
rlabel polysilicon 1150 -1166 1150 -1166 0 1
rlabel polysilicon 1150 -1172 1150 -1172 0 3
rlabel polysilicon 2 -1249 2 -1249 0 1
rlabel polysilicon 2 -1255 2 -1255 0 3
rlabel polysilicon 9 -1249 9 -1249 0 1
rlabel polysilicon 9 -1255 9 -1255 0 3
rlabel polysilicon 16 -1249 16 -1249 0 1
rlabel polysilicon 16 -1255 16 -1255 0 3
rlabel polysilicon 23 -1249 23 -1249 0 1
rlabel polysilicon 30 -1249 30 -1249 0 1
rlabel polysilicon 30 -1255 30 -1255 0 3
rlabel polysilicon 37 -1249 37 -1249 0 1
rlabel polysilicon 37 -1255 37 -1255 0 3
rlabel polysilicon 44 -1249 44 -1249 0 1
rlabel polysilicon 44 -1255 44 -1255 0 3
rlabel polysilicon 47 -1255 47 -1255 0 4
rlabel polysilicon 51 -1249 51 -1249 0 1
rlabel polysilicon 51 -1255 51 -1255 0 3
rlabel polysilicon 58 -1249 58 -1249 0 1
rlabel polysilicon 58 -1255 58 -1255 0 3
rlabel polysilicon 65 -1249 65 -1249 0 1
rlabel polysilicon 65 -1255 65 -1255 0 3
rlabel polysilicon 72 -1255 72 -1255 0 3
rlabel polysilicon 79 -1249 79 -1249 0 1
rlabel polysilicon 79 -1255 79 -1255 0 3
rlabel polysilicon 86 -1249 86 -1249 0 1
rlabel polysilicon 86 -1255 86 -1255 0 3
rlabel polysilicon 93 -1249 93 -1249 0 1
rlabel polysilicon 96 -1249 96 -1249 0 2
rlabel polysilicon 100 -1249 100 -1249 0 1
rlabel polysilicon 100 -1255 100 -1255 0 3
rlabel polysilicon 107 -1249 107 -1249 0 1
rlabel polysilicon 107 -1255 107 -1255 0 3
rlabel polysilicon 114 -1249 114 -1249 0 1
rlabel polysilicon 114 -1255 114 -1255 0 3
rlabel polysilicon 121 -1249 121 -1249 0 1
rlabel polysilicon 121 -1255 121 -1255 0 3
rlabel polysilicon 128 -1249 128 -1249 0 1
rlabel polysilicon 128 -1255 128 -1255 0 3
rlabel polysilicon 135 -1249 135 -1249 0 1
rlabel polysilicon 135 -1255 135 -1255 0 3
rlabel polysilicon 142 -1249 142 -1249 0 1
rlabel polysilicon 142 -1255 142 -1255 0 3
rlabel polysilicon 149 -1249 149 -1249 0 1
rlabel polysilicon 149 -1255 149 -1255 0 3
rlabel polysilicon 159 -1249 159 -1249 0 2
rlabel polysilicon 156 -1255 156 -1255 0 3
rlabel polysilicon 159 -1255 159 -1255 0 4
rlabel polysilicon 163 -1249 163 -1249 0 1
rlabel polysilicon 163 -1255 163 -1255 0 3
rlabel polysilicon 170 -1249 170 -1249 0 1
rlabel polysilicon 170 -1255 170 -1255 0 3
rlabel polysilicon 177 -1249 177 -1249 0 1
rlabel polysilicon 177 -1255 177 -1255 0 3
rlabel polysilicon 184 -1249 184 -1249 0 1
rlabel polysilicon 184 -1255 184 -1255 0 3
rlabel polysilicon 187 -1255 187 -1255 0 4
rlabel polysilicon 194 -1249 194 -1249 0 2
rlabel polysilicon 191 -1255 191 -1255 0 3
rlabel polysilicon 194 -1255 194 -1255 0 4
rlabel polysilicon 201 -1249 201 -1249 0 2
rlabel polysilicon 198 -1255 198 -1255 0 3
rlabel polysilicon 205 -1249 205 -1249 0 1
rlabel polysilicon 205 -1255 205 -1255 0 3
rlabel polysilicon 212 -1249 212 -1249 0 1
rlabel polysilicon 212 -1255 212 -1255 0 3
rlabel polysilicon 219 -1249 219 -1249 0 1
rlabel polysilicon 219 -1255 219 -1255 0 3
rlabel polysilicon 226 -1249 226 -1249 0 1
rlabel polysilicon 226 -1255 226 -1255 0 3
rlabel polysilicon 233 -1249 233 -1249 0 1
rlabel polysilicon 233 -1255 233 -1255 0 3
rlabel polysilicon 240 -1249 240 -1249 0 1
rlabel polysilicon 240 -1255 240 -1255 0 3
rlabel polysilicon 247 -1249 247 -1249 0 1
rlabel polysilicon 247 -1255 247 -1255 0 3
rlabel polysilicon 254 -1249 254 -1249 0 1
rlabel polysilicon 254 -1255 254 -1255 0 3
rlabel polysilicon 261 -1249 261 -1249 0 1
rlabel polysilicon 261 -1255 261 -1255 0 3
rlabel polysilicon 268 -1249 268 -1249 0 1
rlabel polysilicon 271 -1249 271 -1249 0 2
rlabel polysilicon 268 -1255 268 -1255 0 3
rlabel polysilicon 271 -1255 271 -1255 0 4
rlabel polysilicon 275 -1249 275 -1249 0 1
rlabel polysilicon 275 -1255 275 -1255 0 3
rlabel polysilicon 282 -1249 282 -1249 0 1
rlabel polysilicon 282 -1255 282 -1255 0 3
rlabel polysilicon 289 -1249 289 -1249 0 1
rlabel polysilicon 289 -1255 289 -1255 0 3
rlabel polysilicon 292 -1255 292 -1255 0 4
rlabel polysilicon 296 -1249 296 -1249 0 1
rlabel polysilicon 296 -1255 296 -1255 0 3
rlabel polysilicon 303 -1249 303 -1249 0 1
rlabel polysilicon 303 -1255 303 -1255 0 3
rlabel polysilicon 310 -1249 310 -1249 0 1
rlabel polysilicon 310 -1255 310 -1255 0 3
rlabel polysilicon 317 -1249 317 -1249 0 1
rlabel polysilicon 317 -1255 317 -1255 0 3
rlabel polysilicon 324 -1249 324 -1249 0 1
rlabel polysilicon 324 -1255 324 -1255 0 3
rlabel polysilicon 331 -1249 331 -1249 0 1
rlabel polysilicon 331 -1255 331 -1255 0 3
rlabel polysilicon 338 -1249 338 -1249 0 1
rlabel polysilicon 338 -1255 338 -1255 0 3
rlabel polysilicon 345 -1249 345 -1249 0 1
rlabel polysilicon 345 -1255 345 -1255 0 3
rlabel polysilicon 352 -1249 352 -1249 0 1
rlabel polysilicon 352 -1255 352 -1255 0 3
rlabel polysilicon 359 -1249 359 -1249 0 1
rlabel polysilicon 359 -1255 359 -1255 0 3
rlabel polysilicon 366 -1249 366 -1249 0 1
rlabel polysilicon 369 -1249 369 -1249 0 2
rlabel polysilicon 366 -1255 366 -1255 0 3
rlabel polysilicon 369 -1255 369 -1255 0 4
rlabel polysilicon 373 -1249 373 -1249 0 1
rlabel polysilicon 376 -1249 376 -1249 0 2
rlabel polysilicon 380 -1249 380 -1249 0 1
rlabel polysilicon 380 -1255 380 -1255 0 3
rlabel polysilicon 387 -1249 387 -1249 0 1
rlabel polysilicon 387 -1255 387 -1255 0 3
rlabel polysilicon 394 -1249 394 -1249 0 1
rlabel polysilicon 394 -1255 394 -1255 0 3
rlabel polysilicon 401 -1249 401 -1249 0 1
rlabel polysilicon 401 -1255 401 -1255 0 3
rlabel polysilicon 408 -1249 408 -1249 0 1
rlabel polysilicon 408 -1255 408 -1255 0 3
rlabel polysilicon 415 -1249 415 -1249 0 1
rlabel polysilicon 415 -1255 415 -1255 0 3
rlabel polysilicon 422 -1249 422 -1249 0 1
rlabel polysilicon 422 -1255 422 -1255 0 3
rlabel polysilicon 429 -1249 429 -1249 0 1
rlabel polysilicon 429 -1255 429 -1255 0 3
rlabel polysilicon 436 -1249 436 -1249 0 1
rlabel polysilicon 436 -1255 436 -1255 0 3
rlabel polysilicon 443 -1249 443 -1249 0 1
rlabel polysilicon 443 -1255 443 -1255 0 3
rlabel polysilicon 450 -1249 450 -1249 0 1
rlabel polysilicon 457 -1249 457 -1249 0 1
rlabel polysilicon 460 -1249 460 -1249 0 2
rlabel polysilicon 457 -1255 457 -1255 0 3
rlabel polysilicon 460 -1255 460 -1255 0 4
rlabel polysilicon 464 -1249 464 -1249 0 1
rlabel polysilicon 464 -1255 464 -1255 0 3
rlabel polysilicon 471 -1249 471 -1249 0 1
rlabel polysilicon 471 -1255 471 -1255 0 3
rlabel polysilicon 478 -1249 478 -1249 0 1
rlabel polysilicon 478 -1255 478 -1255 0 3
rlabel polysilicon 485 -1249 485 -1249 0 1
rlabel polysilicon 485 -1255 485 -1255 0 3
rlabel polysilicon 492 -1249 492 -1249 0 1
rlabel polysilicon 492 -1255 492 -1255 0 3
rlabel polysilicon 495 -1255 495 -1255 0 4
rlabel polysilicon 499 -1249 499 -1249 0 1
rlabel polysilicon 499 -1255 499 -1255 0 3
rlabel polysilicon 506 -1249 506 -1249 0 1
rlabel polysilicon 509 -1249 509 -1249 0 2
rlabel polysilicon 506 -1255 506 -1255 0 3
rlabel polysilicon 509 -1255 509 -1255 0 4
rlabel polysilicon 513 -1249 513 -1249 0 1
rlabel polysilicon 513 -1255 513 -1255 0 3
rlabel polysilicon 520 -1249 520 -1249 0 1
rlabel polysilicon 520 -1255 520 -1255 0 3
rlabel polysilicon 527 -1249 527 -1249 0 1
rlabel polysilicon 527 -1255 527 -1255 0 3
rlabel polysilicon 537 -1249 537 -1249 0 2
rlabel polysilicon 534 -1255 534 -1255 0 3
rlabel polysilicon 541 -1249 541 -1249 0 1
rlabel polysilicon 541 -1255 541 -1255 0 3
rlabel polysilicon 548 -1249 548 -1249 0 1
rlabel polysilicon 548 -1255 548 -1255 0 3
rlabel polysilicon 555 -1249 555 -1249 0 1
rlabel polysilicon 555 -1255 555 -1255 0 3
rlabel polysilicon 562 -1249 562 -1249 0 1
rlabel polysilicon 562 -1255 562 -1255 0 3
rlabel polysilicon 569 -1249 569 -1249 0 1
rlabel polysilicon 569 -1255 569 -1255 0 3
rlabel polysilicon 576 -1249 576 -1249 0 1
rlabel polysilicon 576 -1255 576 -1255 0 3
rlabel polysilicon 583 -1249 583 -1249 0 1
rlabel polysilicon 583 -1255 583 -1255 0 3
rlabel polysilicon 590 -1249 590 -1249 0 1
rlabel polysilicon 590 -1255 590 -1255 0 3
rlabel polysilicon 600 -1249 600 -1249 0 2
rlabel polysilicon 597 -1255 597 -1255 0 3
rlabel polysilicon 600 -1255 600 -1255 0 4
rlabel polysilicon 604 -1249 604 -1249 0 1
rlabel polysilicon 604 -1255 604 -1255 0 3
rlabel polysilicon 611 -1249 611 -1249 0 1
rlabel polysilicon 611 -1255 611 -1255 0 3
rlabel polysilicon 618 -1249 618 -1249 0 1
rlabel polysilicon 618 -1255 618 -1255 0 3
rlabel polysilicon 625 -1249 625 -1249 0 1
rlabel polysilicon 625 -1255 625 -1255 0 3
rlabel polysilicon 632 -1255 632 -1255 0 3
rlabel polysilicon 635 -1255 635 -1255 0 4
rlabel polysilicon 642 -1249 642 -1249 0 2
rlabel polysilicon 639 -1255 639 -1255 0 3
rlabel polysilicon 642 -1255 642 -1255 0 4
rlabel polysilicon 646 -1249 646 -1249 0 1
rlabel polysilicon 646 -1255 646 -1255 0 3
rlabel polysilicon 656 -1249 656 -1249 0 2
rlabel polysilicon 653 -1255 653 -1255 0 3
rlabel polysilicon 656 -1255 656 -1255 0 4
rlabel polysilicon 660 -1249 660 -1249 0 1
rlabel polysilicon 660 -1255 660 -1255 0 3
rlabel polysilicon 667 -1249 667 -1249 0 1
rlabel polysilicon 670 -1249 670 -1249 0 2
rlabel polysilicon 667 -1255 667 -1255 0 3
rlabel polysilicon 670 -1255 670 -1255 0 4
rlabel polysilicon 674 -1249 674 -1249 0 1
rlabel polysilicon 674 -1255 674 -1255 0 3
rlabel polysilicon 681 -1249 681 -1249 0 1
rlabel polysilicon 684 -1249 684 -1249 0 2
rlabel polysilicon 688 -1249 688 -1249 0 1
rlabel polysilicon 688 -1255 688 -1255 0 3
rlabel polysilicon 695 -1249 695 -1249 0 1
rlabel polysilicon 695 -1255 695 -1255 0 3
rlabel polysilicon 702 -1249 702 -1249 0 1
rlabel polysilicon 705 -1249 705 -1249 0 2
rlabel polysilicon 705 -1255 705 -1255 0 4
rlabel polysilicon 709 -1249 709 -1249 0 1
rlabel polysilicon 709 -1255 709 -1255 0 3
rlabel polysilicon 716 -1249 716 -1249 0 1
rlabel polysilicon 719 -1249 719 -1249 0 2
rlabel polysilicon 723 -1249 723 -1249 0 1
rlabel polysilicon 723 -1255 723 -1255 0 3
rlabel polysilicon 730 -1249 730 -1249 0 1
rlabel polysilicon 730 -1255 730 -1255 0 3
rlabel polysilicon 737 -1249 737 -1249 0 1
rlabel polysilicon 737 -1255 737 -1255 0 3
rlabel polysilicon 744 -1249 744 -1249 0 1
rlabel polysilicon 744 -1255 744 -1255 0 3
rlabel polysilicon 751 -1249 751 -1249 0 1
rlabel polysilicon 751 -1255 751 -1255 0 3
rlabel polysilicon 758 -1249 758 -1249 0 1
rlabel polysilicon 758 -1255 758 -1255 0 3
rlabel polysilicon 765 -1249 765 -1249 0 1
rlabel polysilicon 765 -1255 765 -1255 0 3
rlabel polysilicon 772 -1249 772 -1249 0 1
rlabel polysilicon 772 -1255 772 -1255 0 3
rlabel polysilicon 779 -1249 779 -1249 0 1
rlabel polysilicon 779 -1255 779 -1255 0 3
rlabel polysilicon 786 -1249 786 -1249 0 1
rlabel polysilicon 789 -1255 789 -1255 0 4
rlabel polysilicon 793 -1249 793 -1249 0 1
rlabel polysilicon 793 -1255 793 -1255 0 3
rlabel polysilicon 800 -1249 800 -1249 0 1
rlabel polysilicon 800 -1255 800 -1255 0 3
rlabel polysilicon 807 -1249 807 -1249 0 1
rlabel polysilicon 807 -1255 807 -1255 0 3
rlabel polysilicon 814 -1249 814 -1249 0 1
rlabel polysilicon 814 -1255 814 -1255 0 3
rlabel polysilicon 821 -1249 821 -1249 0 1
rlabel polysilicon 821 -1255 821 -1255 0 3
rlabel polysilicon 828 -1255 828 -1255 0 3
rlabel polysilicon 831 -1255 831 -1255 0 4
rlabel polysilicon 835 -1249 835 -1249 0 1
rlabel polysilicon 835 -1255 835 -1255 0 3
rlabel polysilicon 842 -1249 842 -1249 0 1
rlabel polysilicon 842 -1255 842 -1255 0 3
rlabel polysilicon 849 -1249 849 -1249 0 1
rlabel polysilicon 849 -1255 849 -1255 0 3
rlabel polysilicon 856 -1249 856 -1249 0 1
rlabel polysilicon 856 -1255 856 -1255 0 3
rlabel polysilicon 863 -1249 863 -1249 0 1
rlabel polysilicon 863 -1255 863 -1255 0 3
rlabel polysilicon 870 -1249 870 -1249 0 1
rlabel polysilicon 870 -1255 870 -1255 0 3
rlabel polysilicon 877 -1249 877 -1249 0 1
rlabel polysilicon 877 -1255 877 -1255 0 3
rlabel polysilicon 884 -1249 884 -1249 0 1
rlabel polysilicon 884 -1255 884 -1255 0 3
rlabel polysilicon 891 -1249 891 -1249 0 1
rlabel polysilicon 891 -1255 891 -1255 0 3
rlabel polysilicon 898 -1249 898 -1249 0 1
rlabel polysilicon 898 -1255 898 -1255 0 3
rlabel polysilicon 905 -1249 905 -1249 0 1
rlabel polysilicon 905 -1255 905 -1255 0 3
rlabel polysilicon 912 -1249 912 -1249 0 1
rlabel polysilicon 912 -1255 912 -1255 0 3
rlabel polysilicon 919 -1249 919 -1249 0 1
rlabel polysilicon 919 -1255 919 -1255 0 3
rlabel polysilicon 926 -1249 926 -1249 0 1
rlabel polysilicon 926 -1255 926 -1255 0 3
rlabel polysilicon 933 -1249 933 -1249 0 1
rlabel polysilicon 933 -1255 933 -1255 0 3
rlabel polysilicon 940 -1249 940 -1249 0 1
rlabel polysilicon 940 -1255 940 -1255 0 3
rlabel polysilicon 947 -1249 947 -1249 0 1
rlabel polysilicon 947 -1255 947 -1255 0 3
rlabel polysilicon 954 -1249 954 -1249 0 1
rlabel polysilicon 954 -1255 954 -1255 0 3
rlabel polysilicon 961 -1249 961 -1249 0 1
rlabel polysilicon 961 -1255 961 -1255 0 3
rlabel polysilicon 968 -1249 968 -1249 0 1
rlabel polysilicon 968 -1255 968 -1255 0 3
rlabel polysilicon 975 -1249 975 -1249 0 1
rlabel polysilicon 975 -1255 975 -1255 0 3
rlabel polysilicon 982 -1249 982 -1249 0 1
rlabel polysilicon 982 -1255 982 -1255 0 3
rlabel polysilicon 989 -1249 989 -1249 0 1
rlabel polysilicon 989 -1255 989 -1255 0 3
rlabel polysilicon 996 -1249 996 -1249 0 1
rlabel polysilicon 996 -1255 996 -1255 0 3
rlabel polysilicon 1003 -1249 1003 -1249 0 1
rlabel polysilicon 1003 -1255 1003 -1255 0 3
rlabel polysilicon 1010 -1249 1010 -1249 0 1
rlabel polysilicon 1010 -1255 1010 -1255 0 3
rlabel polysilicon 1017 -1249 1017 -1249 0 1
rlabel polysilicon 1017 -1255 1017 -1255 0 3
rlabel polysilicon 1024 -1249 1024 -1249 0 1
rlabel polysilicon 1024 -1255 1024 -1255 0 3
rlabel polysilicon 1027 -1255 1027 -1255 0 4
rlabel polysilicon 1031 -1249 1031 -1249 0 1
rlabel polysilicon 1031 -1255 1031 -1255 0 3
rlabel polysilicon 1038 -1249 1038 -1249 0 1
rlabel polysilicon 1038 -1255 1038 -1255 0 3
rlabel polysilicon 1045 -1249 1045 -1249 0 1
rlabel polysilicon 1045 -1255 1045 -1255 0 3
rlabel polysilicon 1052 -1249 1052 -1249 0 1
rlabel polysilicon 1052 -1255 1052 -1255 0 3
rlabel polysilicon 1059 -1249 1059 -1249 0 1
rlabel polysilicon 1059 -1255 1059 -1255 0 3
rlabel polysilicon 1066 -1249 1066 -1249 0 1
rlabel polysilicon 1066 -1255 1066 -1255 0 3
rlabel polysilicon 1073 -1249 1073 -1249 0 1
rlabel polysilicon 1073 -1255 1073 -1255 0 3
rlabel polysilicon 1080 -1249 1080 -1249 0 1
rlabel polysilicon 1080 -1255 1080 -1255 0 3
rlabel polysilicon 1087 -1249 1087 -1249 0 1
rlabel polysilicon 1087 -1255 1087 -1255 0 3
rlabel polysilicon 1094 -1249 1094 -1249 0 1
rlabel polysilicon 1094 -1255 1094 -1255 0 3
rlabel polysilicon 1101 -1249 1101 -1249 0 1
rlabel polysilicon 1101 -1255 1101 -1255 0 3
rlabel polysilicon 1108 -1249 1108 -1249 0 1
rlabel polysilicon 1108 -1255 1108 -1255 0 3
rlabel polysilicon 1115 -1249 1115 -1249 0 1
rlabel polysilicon 1118 -1249 1118 -1249 0 2
rlabel polysilicon 1115 -1255 1115 -1255 0 3
rlabel polysilicon 1122 -1249 1122 -1249 0 1
rlabel polysilicon 1122 -1255 1122 -1255 0 3
rlabel polysilicon 1129 -1249 1129 -1249 0 1
rlabel polysilicon 1132 -1255 1132 -1255 0 4
rlabel polysilicon 1136 -1249 1136 -1249 0 1
rlabel polysilicon 1136 -1255 1136 -1255 0 3
rlabel polysilicon 1143 -1249 1143 -1249 0 1
rlabel polysilicon 1143 -1255 1143 -1255 0 3
rlabel polysilicon 1150 -1249 1150 -1249 0 1
rlabel polysilicon 1150 -1255 1150 -1255 0 3
rlabel polysilicon 1157 -1249 1157 -1249 0 1
rlabel polysilicon 1157 -1255 1157 -1255 0 3
rlabel polysilicon 1164 -1249 1164 -1249 0 1
rlabel polysilicon 1164 -1255 1164 -1255 0 3
rlabel polysilicon 2 -1342 2 -1342 0 1
rlabel polysilicon 2 -1348 2 -1348 0 3
rlabel polysilicon 9 -1342 9 -1342 0 1
rlabel polysilicon 9 -1348 9 -1348 0 3
rlabel polysilicon 16 -1342 16 -1342 0 1
rlabel polysilicon 16 -1348 16 -1348 0 3
rlabel polysilicon 23 -1342 23 -1342 0 1
rlabel polysilicon 26 -1342 26 -1342 0 2
rlabel polysilicon 26 -1348 26 -1348 0 4
rlabel polysilicon 33 -1342 33 -1342 0 2
rlabel polysilicon 30 -1348 30 -1348 0 3
rlabel polysilicon 33 -1348 33 -1348 0 4
rlabel polysilicon 37 -1342 37 -1342 0 1
rlabel polysilicon 37 -1348 37 -1348 0 3
rlabel polysilicon 44 -1342 44 -1342 0 1
rlabel polysilicon 44 -1348 44 -1348 0 3
rlabel polysilicon 51 -1342 51 -1342 0 1
rlabel polysilicon 51 -1348 51 -1348 0 3
rlabel polysilicon 58 -1342 58 -1342 0 1
rlabel polysilicon 58 -1348 58 -1348 0 3
rlabel polysilicon 65 -1348 65 -1348 0 3
rlabel polysilicon 68 -1348 68 -1348 0 4
rlabel polysilicon 72 -1342 72 -1342 0 1
rlabel polysilicon 72 -1348 72 -1348 0 3
rlabel polysilicon 79 -1342 79 -1342 0 1
rlabel polysilicon 79 -1348 79 -1348 0 3
rlabel polysilicon 86 -1342 86 -1342 0 1
rlabel polysilicon 86 -1348 86 -1348 0 3
rlabel polysilicon 96 -1342 96 -1342 0 2
rlabel polysilicon 93 -1348 93 -1348 0 3
rlabel polysilicon 96 -1348 96 -1348 0 4
rlabel polysilicon 100 -1342 100 -1342 0 1
rlabel polysilicon 103 -1342 103 -1342 0 2
rlabel polysilicon 100 -1348 100 -1348 0 3
rlabel polysilicon 103 -1348 103 -1348 0 4
rlabel polysilicon 107 -1342 107 -1342 0 1
rlabel polysilicon 107 -1348 107 -1348 0 3
rlabel polysilicon 114 -1342 114 -1342 0 1
rlabel polysilicon 114 -1348 114 -1348 0 3
rlabel polysilicon 121 -1342 121 -1342 0 1
rlabel polysilicon 121 -1348 121 -1348 0 3
rlabel polysilicon 128 -1342 128 -1342 0 1
rlabel polysilicon 128 -1348 128 -1348 0 3
rlabel polysilicon 135 -1342 135 -1342 0 1
rlabel polysilicon 135 -1348 135 -1348 0 3
rlabel polysilicon 142 -1342 142 -1342 0 1
rlabel polysilicon 142 -1348 142 -1348 0 3
rlabel polysilicon 149 -1342 149 -1342 0 1
rlabel polysilicon 149 -1348 149 -1348 0 3
rlabel polysilicon 156 -1342 156 -1342 0 1
rlabel polysilicon 156 -1348 156 -1348 0 3
rlabel polysilicon 163 -1348 163 -1348 0 3
rlabel polysilicon 170 -1342 170 -1342 0 1
rlabel polysilicon 170 -1348 170 -1348 0 3
rlabel polysilicon 180 -1342 180 -1342 0 2
rlabel polysilicon 177 -1348 177 -1348 0 3
rlabel polysilicon 184 -1342 184 -1342 0 1
rlabel polysilicon 184 -1348 184 -1348 0 3
rlabel polysilicon 191 -1342 191 -1342 0 1
rlabel polysilicon 191 -1348 191 -1348 0 3
rlabel polysilicon 198 -1342 198 -1342 0 1
rlabel polysilicon 198 -1348 198 -1348 0 3
rlabel polysilicon 205 -1342 205 -1342 0 1
rlabel polysilicon 205 -1348 205 -1348 0 3
rlabel polysilicon 212 -1342 212 -1342 0 1
rlabel polysilicon 215 -1342 215 -1342 0 2
rlabel polysilicon 212 -1348 212 -1348 0 3
rlabel polysilicon 215 -1348 215 -1348 0 4
rlabel polysilicon 219 -1342 219 -1342 0 1
rlabel polysilicon 219 -1348 219 -1348 0 3
rlabel polysilicon 226 -1342 226 -1342 0 1
rlabel polysilicon 226 -1348 226 -1348 0 3
rlabel polysilicon 233 -1342 233 -1342 0 1
rlabel polysilicon 233 -1348 233 -1348 0 3
rlabel polysilicon 240 -1342 240 -1342 0 1
rlabel polysilicon 240 -1348 240 -1348 0 3
rlabel polysilicon 247 -1342 247 -1342 0 1
rlabel polysilicon 247 -1348 247 -1348 0 3
rlabel polysilicon 254 -1342 254 -1342 0 1
rlabel polysilicon 254 -1348 254 -1348 0 3
rlabel polysilicon 261 -1342 261 -1342 0 1
rlabel polysilicon 261 -1348 261 -1348 0 3
rlabel polysilicon 268 -1342 268 -1342 0 1
rlabel polysilicon 268 -1348 268 -1348 0 3
rlabel polysilicon 275 -1342 275 -1342 0 1
rlabel polysilicon 275 -1348 275 -1348 0 3
rlabel polysilicon 282 -1342 282 -1342 0 1
rlabel polysilicon 282 -1348 282 -1348 0 3
rlabel polysilicon 289 -1342 289 -1342 0 1
rlabel polysilicon 292 -1348 292 -1348 0 4
rlabel polysilicon 296 -1342 296 -1342 0 1
rlabel polysilicon 296 -1348 296 -1348 0 3
rlabel polysilicon 303 -1342 303 -1342 0 1
rlabel polysilicon 303 -1348 303 -1348 0 3
rlabel polysilicon 310 -1342 310 -1342 0 1
rlabel polysilicon 310 -1348 310 -1348 0 3
rlabel polysilicon 317 -1342 317 -1342 0 1
rlabel polysilicon 317 -1348 317 -1348 0 3
rlabel polysilicon 324 -1342 324 -1342 0 1
rlabel polysilicon 324 -1348 324 -1348 0 3
rlabel polysilicon 331 -1342 331 -1342 0 1
rlabel polysilicon 331 -1348 331 -1348 0 3
rlabel polysilicon 338 -1342 338 -1342 0 1
rlabel polysilicon 338 -1348 338 -1348 0 3
rlabel polysilicon 345 -1342 345 -1342 0 1
rlabel polysilicon 348 -1342 348 -1342 0 2
rlabel polysilicon 345 -1348 345 -1348 0 3
rlabel polysilicon 348 -1348 348 -1348 0 4
rlabel polysilicon 352 -1342 352 -1342 0 1
rlabel polysilicon 352 -1348 352 -1348 0 3
rlabel polysilicon 359 -1342 359 -1342 0 1
rlabel polysilicon 359 -1348 359 -1348 0 3
rlabel polysilicon 366 -1342 366 -1342 0 1
rlabel polysilicon 366 -1348 366 -1348 0 3
rlabel polysilicon 373 -1342 373 -1342 0 1
rlabel polysilicon 373 -1348 373 -1348 0 3
rlabel polysilicon 380 -1342 380 -1342 0 1
rlabel polysilicon 380 -1348 380 -1348 0 3
rlabel polysilicon 387 -1342 387 -1342 0 1
rlabel polysilicon 387 -1348 387 -1348 0 3
rlabel polysilicon 394 -1342 394 -1342 0 1
rlabel polysilicon 394 -1348 394 -1348 0 3
rlabel polysilicon 401 -1342 401 -1342 0 1
rlabel polysilicon 404 -1342 404 -1342 0 2
rlabel polysilicon 401 -1348 401 -1348 0 3
rlabel polysilicon 408 -1342 408 -1342 0 1
rlabel polysilicon 411 -1342 411 -1342 0 2
rlabel polysilicon 408 -1348 408 -1348 0 3
rlabel polysilicon 411 -1348 411 -1348 0 4
rlabel polysilicon 415 -1342 415 -1342 0 1
rlabel polysilicon 415 -1348 415 -1348 0 3
rlabel polysilicon 422 -1342 422 -1342 0 1
rlabel polysilicon 422 -1348 422 -1348 0 3
rlabel polysilicon 429 -1342 429 -1342 0 1
rlabel polysilicon 429 -1348 429 -1348 0 3
rlabel polysilicon 436 -1342 436 -1342 0 1
rlabel polysilicon 439 -1342 439 -1342 0 2
rlabel polysilicon 439 -1348 439 -1348 0 4
rlabel polysilicon 443 -1342 443 -1342 0 1
rlabel polysilicon 443 -1348 443 -1348 0 3
rlabel polysilicon 450 -1348 450 -1348 0 3
rlabel polysilicon 457 -1342 457 -1342 0 1
rlabel polysilicon 460 -1342 460 -1342 0 2
rlabel polysilicon 457 -1348 457 -1348 0 3
rlabel polysilicon 460 -1348 460 -1348 0 4
rlabel polysilicon 464 -1342 464 -1342 0 1
rlabel polysilicon 464 -1348 464 -1348 0 3
rlabel polysilicon 471 -1342 471 -1342 0 1
rlabel polysilicon 471 -1348 471 -1348 0 3
rlabel polysilicon 478 -1342 478 -1342 0 1
rlabel polysilicon 478 -1348 478 -1348 0 3
rlabel polysilicon 485 -1342 485 -1342 0 1
rlabel polysilicon 485 -1348 485 -1348 0 3
rlabel polysilicon 492 -1342 492 -1342 0 1
rlabel polysilicon 495 -1348 495 -1348 0 4
rlabel polysilicon 499 -1342 499 -1342 0 1
rlabel polysilicon 499 -1348 499 -1348 0 3
rlabel polysilicon 506 -1342 506 -1342 0 1
rlabel polysilicon 506 -1348 506 -1348 0 3
rlabel polysilicon 513 -1342 513 -1342 0 1
rlabel polysilicon 513 -1348 513 -1348 0 3
rlabel polysilicon 520 -1342 520 -1342 0 1
rlabel polysilicon 523 -1342 523 -1342 0 2
rlabel polysilicon 523 -1348 523 -1348 0 4
rlabel polysilicon 527 -1342 527 -1342 0 1
rlabel polysilicon 527 -1348 527 -1348 0 3
rlabel polysilicon 534 -1342 534 -1342 0 1
rlabel polysilicon 537 -1342 537 -1342 0 2
rlabel polysilicon 534 -1348 534 -1348 0 3
rlabel polysilicon 537 -1348 537 -1348 0 4
rlabel polysilicon 541 -1342 541 -1342 0 1
rlabel polysilicon 544 -1342 544 -1342 0 2
rlabel polysilicon 544 -1348 544 -1348 0 4
rlabel polysilicon 548 -1342 548 -1342 0 1
rlabel polysilicon 548 -1348 548 -1348 0 3
rlabel polysilicon 555 -1342 555 -1342 0 1
rlabel polysilicon 555 -1348 555 -1348 0 3
rlabel polysilicon 562 -1342 562 -1342 0 1
rlabel polysilicon 562 -1348 562 -1348 0 3
rlabel polysilicon 569 -1342 569 -1342 0 1
rlabel polysilicon 572 -1342 572 -1342 0 2
rlabel polysilicon 569 -1348 569 -1348 0 3
rlabel polysilicon 576 -1342 576 -1342 0 1
rlabel polysilicon 576 -1348 576 -1348 0 3
rlabel polysilicon 583 -1342 583 -1342 0 1
rlabel polysilicon 583 -1348 583 -1348 0 3
rlabel polysilicon 590 -1342 590 -1342 0 1
rlabel polysilicon 590 -1348 590 -1348 0 3
rlabel polysilicon 597 -1342 597 -1342 0 1
rlabel polysilicon 597 -1348 597 -1348 0 3
rlabel polysilicon 604 -1342 604 -1342 0 1
rlabel polysilicon 607 -1342 607 -1342 0 2
rlabel polysilicon 604 -1348 604 -1348 0 3
rlabel polysilicon 611 -1342 611 -1342 0 1
rlabel polysilicon 611 -1348 611 -1348 0 3
rlabel polysilicon 614 -1348 614 -1348 0 4
rlabel polysilicon 618 -1342 618 -1342 0 1
rlabel polysilicon 621 -1342 621 -1342 0 2
rlabel polysilicon 618 -1348 618 -1348 0 3
rlabel polysilicon 628 -1342 628 -1342 0 2
rlabel polysilicon 625 -1348 625 -1348 0 3
rlabel polysilicon 632 -1342 632 -1342 0 1
rlabel polysilicon 632 -1348 632 -1348 0 3
rlabel polysilicon 639 -1342 639 -1342 0 1
rlabel polysilicon 639 -1348 639 -1348 0 3
rlabel polysilicon 646 -1342 646 -1342 0 1
rlabel polysilicon 646 -1348 646 -1348 0 3
rlabel polysilicon 653 -1342 653 -1342 0 1
rlabel polysilicon 653 -1348 653 -1348 0 3
rlabel polysilicon 660 -1342 660 -1342 0 1
rlabel polysilicon 660 -1348 660 -1348 0 3
rlabel polysilicon 667 -1342 667 -1342 0 1
rlabel polysilicon 667 -1348 667 -1348 0 3
rlabel polysilicon 674 -1342 674 -1342 0 1
rlabel polysilicon 674 -1348 674 -1348 0 3
rlabel polysilicon 681 -1342 681 -1342 0 1
rlabel polysilicon 684 -1342 684 -1342 0 2
rlabel polysilicon 681 -1348 681 -1348 0 3
rlabel polysilicon 688 -1342 688 -1342 0 1
rlabel polysilicon 688 -1348 688 -1348 0 3
rlabel polysilicon 695 -1342 695 -1342 0 1
rlabel polysilicon 695 -1348 695 -1348 0 3
rlabel polysilicon 702 -1342 702 -1342 0 1
rlabel polysilicon 702 -1348 702 -1348 0 3
rlabel polysilicon 709 -1342 709 -1342 0 1
rlabel polysilicon 709 -1348 709 -1348 0 3
rlabel polysilicon 716 -1342 716 -1342 0 1
rlabel polysilicon 716 -1348 716 -1348 0 3
rlabel polysilicon 723 -1342 723 -1342 0 1
rlabel polysilicon 723 -1348 723 -1348 0 3
rlabel polysilicon 733 -1342 733 -1342 0 2
rlabel polysilicon 733 -1348 733 -1348 0 4
rlabel polysilicon 737 -1342 737 -1342 0 1
rlabel polysilicon 737 -1348 737 -1348 0 3
rlabel polysilicon 744 -1342 744 -1342 0 1
rlabel polysilicon 744 -1348 744 -1348 0 3
rlabel polysilicon 751 -1342 751 -1342 0 1
rlabel polysilicon 751 -1348 751 -1348 0 3
rlabel polysilicon 758 -1342 758 -1342 0 1
rlabel polysilicon 758 -1348 758 -1348 0 3
rlabel polysilicon 765 -1342 765 -1342 0 1
rlabel polysilicon 765 -1348 765 -1348 0 3
rlabel polysilicon 772 -1342 772 -1342 0 1
rlabel polysilicon 772 -1348 772 -1348 0 3
rlabel polysilicon 775 -1348 775 -1348 0 4
rlabel polysilicon 779 -1342 779 -1342 0 1
rlabel polysilicon 779 -1348 779 -1348 0 3
rlabel polysilicon 786 -1342 786 -1342 0 1
rlabel polysilicon 786 -1348 786 -1348 0 3
rlabel polysilicon 793 -1342 793 -1342 0 1
rlabel polysilicon 796 -1342 796 -1342 0 2
rlabel polysilicon 793 -1348 793 -1348 0 3
rlabel polysilicon 800 -1342 800 -1342 0 1
rlabel polysilicon 800 -1348 800 -1348 0 3
rlabel polysilicon 807 -1342 807 -1342 0 1
rlabel polysilicon 807 -1348 807 -1348 0 3
rlabel polysilicon 814 -1342 814 -1342 0 1
rlabel polysilicon 814 -1348 814 -1348 0 3
rlabel polysilicon 821 -1342 821 -1342 0 1
rlabel polysilicon 821 -1348 821 -1348 0 3
rlabel polysilicon 828 -1342 828 -1342 0 1
rlabel polysilicon 831 -1342 831 -1342 0 2
rlabel polysilicon 828 -1348 828 -1348 0 3
rlabel polysilicon 835 -1342 835 -1342 0 1
rlabel polysilicon 835 -1348 835 -1348 0 3
rlabel polysilicon 842 -1342 842 -1342 0 1
rlabel polysilicon 842 -1348 842 -1348 0 3
rlabel polysilicon 849 -1342 849 -1342 0 1
rlabel polysilicon 849 -1348 849 -1348 0 3
rlabel polysilicon 856 -1342 856 -1342 0 1
rlabel polysilicon 856 -1348 856 -1348 0 3
rlabel polysilicon 863 -1342 863 -1342 0 1
rlabel polysilicon 863 -1348 863 -1348 0 3
rlabel polysilicon 870 -1342 870 -1342 0 1
rlabel polysilicon 870 -1348 870 -1348 0 3
rlabel polysilicon 877 -1342 877 -1342 0 1
rlabel polysilicon 877 -1348 877 -1348 0 3
rlabel polysilicon 884 -1342 884 -1342 0 1
rlabel polysilicon 884 -1348 884 -1348 0 3
rlabel polysilicon 891 -1342 891 -1342 0 1
rlabel polysilicon 891 -1348 891 -1348 0 3
rlabel polysilicon 898 -1342 898 -1342 0 1
rlabel polysilicon 898 -1348 898 -1348 0 3
rlabel polysilicon 905 -1342 905 -1342 0 1
rlabel polysilicon 905 -1348 905 -1348 0 3
rlabel polysilicon 912 -1342 912 -1342 0 1
rlabel polysilicon 912 -1348 912 -1348 0 3
rlabel polysilicon 919 -1342 919 -1342 0 1
rlabel polysilicon 919 -1348 919 -1348 0 3
rlabel polysilicon 926 -1342 926 -1342 0 1
rlabel polysilicon 926 -1348 926 -1348 0 3
rlabel polysilicon 933 -1342 933 -1342 0 1
rlabel polysilicon 933 -1348 933 -1348 0 3
rlabel polysilicon 940 -1342 940 -1342 0 1
rlabel polysilicon 940 -1348 940 -1348 0 3
rlabel polysilicon 947 -1342 947 -1342 0 1
rlabel polysilicon 950 -1348 950 -1348 0 4
rlabel polysilicon 954 -1342 954 -1342 0 1
rlabel polysilicon 954 -1348 954 -1348 0 3
rlabel polysilicon 961 -1342 961 -1342 0 1
rlabel polysilicon 961 -1348 961 -1348 0 3
rlabel polysilicon 968 -1342 968 -1342 0 1
rlabel polysilicon 968 -1348 968 -1348 0 3
rlabel polysilicon 975 -1342 975 -1342 0 1
rlabel polysilicon 975 -1348 975 -1348 0 3
rlabel polysilicon 982 -1342 982 -1342 0 1
rlabel polysilicon 982 -1348 982 -1348 0 3
rlabel polysilicon 989 -1342 989 -1342 0 1
rlabel polysilicon 989 -1348 989 -1348 0 3
rlabel polysilicon 996 -1342 996 -1342 0 1
rlabel polysilicon 1003 -1342 1003 -1342 0 1
rlabel polysilicon 1003 -1348 1003 -1348 0 3
rlabel polysilicon 1010 -1342 1010 -1342 0 1
rlabel polysilicon 1010 -1348 1010 -1348 0 3
rlabel polysilicon 1017 -1342 1017 -1342 0 1
rlabel polysilicon 1017 -1348 1017 -1348 0 3
rlabel polysilicon 1024 -1342 1024 -1342 0 1
rlabel polysilicon 1027 -1342 1027 -1342 0 2
rlabel polysilicon 1024 -1348 1024 -1348 0 3
rlabel polysilicon 1031 -1342 1031 -1342 0 1
rlabel polysilicon 1031 -1348 1031 -1348 0 3
rlabel polysilicon 1038 -1342 1038 -1342 0 1
rlabel polysilicon 1038 -1348 1038 -1348 0 3
rlabel polysilicon 1045 -1342 1045 -1342 0 1
rlabel polysilicon 1045 -1348 1045 -1348 0 3
rlabel polysilicon 1052 -1342 1052 -1342 0 1
rlabel polysilicon 1052 -1348 1052 -1348 0 3
rlabel polysilicon 1059 -1342 1059 -1342 0 1
rlabel polysilicon 1059 -1348 1059 -1348 0 3
rlabel polysilicon 1066 -1342 1066 -1342 0 1
rlabel polysilicon 1066 -1348 1066 -1348 0 3
rlabel polysilicon 1073 -1342 1073 -1342 0 1
rlabel polysilicon 1073 -1348 1073 -1348 0 3
rlabel polysilicon 1080 -1342 1080 -1342 0 1
rlabel polysilicon 1080 -1348 1080 -1348 0 3
rlabel polysilicon 1087 -1342 1087 -1342 0 1
rlabel polysilicon 1087 -1348 1087 -1348 0 3
rlabel polysilicon 1094 -1342 1094 -1342 0 1
rlabel polysilicon 1094 -1348 1094 -1348 0 3
rlabel polysilicon 1101 -1342 1101 -1342 0 1
rlabel polysilicon 1101 -1348 1101 -1348 0 3
rlabel polysilicon 1108 -1342 1108 -1342 0 1
rlabel polysilicon 1108 -1348 1108 -1348 0 3
rlabel polysilicon 1115 -1342 1115 -1342 0 1
rlabel polysilicon 1115 -1348 1115 -1348 0 3
rlabel polysilicon 1122 -1342 1122 -1342 0 1
rlabel polysilicon 1122 -1348 1122 -1348 0 3
rlabel polysilicon 1129 -1342 1129 -1342 0 1
rlabel polysilicon 1129 -1348 1129 -1348 0 3
rlabel polysilicon 1136 -1342 1136 -1342 0 1
rlabel polysilicon 1136 -1348 1136 -1348 0 3
rlabel polysilicon 1143 -1342 1143 -1342 0 1
rlabel polysilicon 1143 -1348 1143 -1348 0 3
rlabel polysilicon 1150 -1348 1150 -1348 0 3
rlabel polysilicon 1153 -1348 1153 -1348 0 4
rlabel polysilicon 1157 -1342 1157 -1342 0 1
rlabel polysilicon 1157 -1348 1157 -1348 0 3
rlabel polysilicon 1164 -1342 1164 -1342 0 1
rlabel polysilicon 1164 -1348 1164 -1348 0 3
rlabel polysilicon 1171 -1342 1171 -1342 0 1
rlabel polysilicon 1171 -1348 1171 -1348 0 3
rlabel polysilicon 2 -1449 2 -1449 0 1
rlabel polysilicon 2 -1455 2 -1455 0 3
rlabel polysilicon 9 -1455 9 -1455 0 3
rlabel polysilicon 16 -1449 16 -1449 0 1
rlabel polysilicon 16 -1455 16 -1455 0 3
rlabel polysilicon 23 -1449 23 -1449 0 1
rlabel polysilicon 23 -1455 23 -1455 0 3
rlabel polysilicon 30 -1449 30 -1449 0 1
rlabel polysilicon 30 -1455 30 -1455 0 3
rlabel polysilicon 37 -1449 37 -1449 0 1
rlabel polysilicon 37 -1455 37 -1455 0 3
rlabel polysilicon 44 -1449 44 -1449 0 1
rlabel polysilicon 44 -1455 44 -1455 0 3
rlabel polysilicon 51 -1449 51 -1449 0 1
rlabel polysilicon 51 -1455 51 -1455 0 3
rlabel polysilicon 58 -1449 58 -1449 0 1
rlabel polysilicon 58 -1455 58 -1455 0 3
rlabel polysilicon 65 -1449 65 -1449 0 1
rlabel polysilicon 65 -1455 65 -1455 0 3
rlabel polysilicon 72 -1449 72 -1449 0 1
rlabel polysilicon 72 -1455 72 -1455 0 3
rlabel polysilicon 79 -1449 79 -1449 0 1
rlabel polysilicon 79 -1455 79 -1455 0 3
rlabel polysilicon 86 -1449 86 -1449 0 1
rlabel polysilicon 86 -1455 86 -1455 0 3
rlabel polysilicon 93 -1449 93 -1449 0 1
rlabel polysilicon 93 -1455 93 -1455 0 3
rlabel polysilicon 100 -1449 100 -1449 0 1
rlabel polysilicon 103 -1449 103 -1449 0 2
rlabel polysilicon 103 -1455 103 -1455 0 4
rlabel polysilicon 110 -1449 110 -1449 0 2
rlabel polysilicon 107 -1455 107 -1455 0 3
rlabel polysilicon 110 -1455 110 -1455 0 4
rlabel polysilicon 114 -1455 114 -1455 0 3
rlabel polysilicon 121 -1449 121 -1449 0 1
rlabel polysilicon 124 -1455 124 -1455 0 4
rlabel polysilicon 128 -1449 128 -1449 0 1
rlabel polysilicon 128 -1455 128 -1455 0 3
rlabel polysilicon 135 -1449 135 -1449 0 1
rlabel polysilicon 135 -1455 135 -1455 0 3
rlabel polysilicon 142 -1449 142 -1449 0 1
rlabel polysilicon 142 -1455 142 -1455 0 3
rlabel polysilicon 149 -1449 149 -1449 0 1
rlabel polysilicon 149 -1455 149 -1455 0 3
rlabel polysilicon 156 -1449 156 -1449 0 1
rlabel polysilicon 156 -1455 156 -1455 0 3
rlabel polysilicon 163 -1449 163 -1449 0 1
rlabel polysilicon 163 -1455 163 -1455 0 3
rlabel polysilicon 170 -1449 170 -1449 0 1
rlabel polysilicon 170 -1455 170 -1455 0 3
rlabel polysilicon 177 -1449 177 -1449 0 1
rlabel polysilicon 177 -1455 177 -1455 0 3
rlabel polysilicon 180 -1455 180 -1455 0 4
rlabel polysilicon 187 -1449 187 -1449 0 2
rlabel polysilicon 184 -1455 184 -1455 0 3
rlabel polysilicon 187 -1455 187 -1455 0 4
rlabel polysilicon 194 -1449 194 -1449 0 2
rlabel polysilicon 191 -1455 191 -1455 0 3
rlabel polysilicon 194 -1455 194 -1455 0 4
rlabel polysilicon 198 -1449 198 -1449 0 1
rlabel polysilicon 198 -1455 198 -1455 0 3
rlabel polysilicon 205 -1449 205 -1449 0 1
rlabel polysilicon 205 -1455 205 -1455 0 3
rlabel polysilicon 212 -1455 212 -1455 0 3
rlabel polysilicon 215 -1455 215 -1455 0 4
rlabel polysilicon 219 -1449 219 -1449 0 1
rlabel polysilicon 219 -1455 219 -1455 0 3
rlabel polysilicon 226 -1449 226 -1449 0 1
rlabel polysilicon 226 -1455 226 -1455 0 3
rlabel polysilicon 233 -1449 233 -1449 0 1
rlabel polysilicon 233 -1455 233 -1455 0 3
rlabel polysilicon 240 -1449 240 -1449 0 1
rlabel polysilicon 240 -1455 240 -1455 0 3
rlabel polysilicon 247 -1449 247 -1449 0 1
rlabel polysilicon 247 -1455 247 -1455 0 3
rlabel polysilicon 254 -1449 254 -1449 0 1
rlabel polysilicon 254 -1455 254 -1455 0 3
rlabel polysilicon 257 -1455 257 -1455 0 4
rlabel polysilicon 261 -1449 261 -1449 0 1
rlabel polysilicon 261 -1455 261 -1455 0 3
rlabel polysilicon 268 -1449 268 -1449 0 1
rlabel polysilicon 268 -1455 268 -1455 0 3
rlabel polysilicon 275 -1449 275 -1449 0 1
rlabel polysilicon 275 -1455 275 -1455 0 3
rlabel polysilicon 282 -1449 282 -1449 0 1
rlabel polysilicon 282 -1455 282 -1455 0 3
rlabel polysilicon 289 -1449 289 -1449 0 1
rlabel polysilicon 289 -1455 289 -1455 0 3
rlabel polysilicon 296 -1449 296 -1449 0 1
rlabel polysilicon 296 -1455 296 -1455 0 3
rlabel polysilicon 303 -1449 303 -1449 0 1
rlabel polysilicon 303 -1455 303 -1455 0 3
rlabel polysilicon 310 -1449 310 -1449 0 1
rlabel polysilicon 310 -1455 310 -1455 0 3
rlabel polysilicon 317 -1449 317 -1449 0 1
rlabel polysilicon 317 -1455 317 -1455 0 3
rlabel polysilicon 324 -1449 324 -1449 0 1
rlabel polysilicon 324 -1455 324 -1455 0 3
rlabel polysilicon 331 -1449 331 -1449 0 1
rlabel polysilicon 334 -1449 334 -1449 0 2
rlabel polysilicon 331 -1455 331 -1455 0 3
rlabel polysilicon 334 -1455 334 -1455 0 4
rlabel polysilicon 338 -1449 338 -1449 0 1
rlabel polysilicon 338 -1455 338 -1455 0 3
rlabel polysilicon 345 -1449 345 -1449 0 1
rlabel polysilicon 345 -1455 345 -1455 0 3
rlabel polysilicon 352 -1449 352 -1449 0 1
rlabel polysilicon 352 -1455 352 -1455 0 3
rlabel polysilicon 359 -1449 359 -1449 0 1
rlabel polysilicon 359 -1455 359 -1455 0 3
rlabel polysilicon 366 -1449 366 -1449 0 1
rlabel polysilicon 366 -1455 366 -1455 0 3
rlabel polysilicon 373 -1449 373 -1449 0 1
rlabel polysilicon 373 -1455 373 -1455 0 3
rlabel polysilicon 380 -1449 380 -1449 0 1
rlabel polysilicon 380 -1455 380 -1455 0 3
rlabel polysilicon 387 -1449 387 -1449 0 1
rlabel polysilicon 387 -1455 387 -1455 0 3
rlabel polysilicon 394 -1449 394 -1449 0 1
rlabel polysilicon 394 -1455 394 -1455 0 3
rlabel polysilicon 401 -1449 401 -1449 0 1
rlabel polysilicon 404 -1449 404 -1449 0 2
rlabel polysilicon 404 -1455 404 -1455 0 4
rlabel polysilicon 408 -1449 408 -1449 0 1
rlabel polysilicon 408 -1455 408 -1455 0 3
rlabel polysilicon 411 -1455 411 -1455 0 4
rlabel polysilicon 415 -1449 415 -1449 0 1
rlabel polysilicon 415 -1455 415 -1455 0 3
rlabel polysilicon 422 -1449 422 -1449 0 1
rlabel polysilicon 422 -1455 422 -1455 0 3
rlabel polysilicon 432 -1449 432 -1449 0 2
rlabel polysilicon 432 -1455 432 -1455 0 4
rlabel polysilicon 436 -1449 436 -1449 0 1
rlabel polysilicon 439 -1449 439 -1449 0 2
rlabel polysilicon 439 -1455 439 -1455 0 4
rlabel polysilicon 446 -1449 446 -1449 0 2
rlabel polysilicon 443 -1455 443 -1455 0 3
rlabel polysilicon 450 -1449 450 -1449 0 1
rlabel polysilicon 450 -1455 450 -1455 0 3
rlabel polysilicon 457 -1449 457 -1449 0 1
rlabel polysilicon 457 -1455 457 -1455 0 3
rlabel polysilicon 464 -1449 464 -1449 0 1
rlabel polysilicon 464 -1455 464 -1455 0 3
rlabel polysilicon 471 -1449 471 -1449 0 1
rlabel polysilicon 471 -1455 471 -1455 0 3
rlabel polysilicon 478 -1449 478 -1449 0 1
rlabel polysilicon 485 -1449 485 -1449 0 1
rlabel polysilicon 488 -1449 488 -1449 0 2
rlabel polysilicon 485 -1455 485 -1455 0 3
rlabel polysilicon 492 -1449 492 -1449 0 1
rlabel polysilicon 495 -1449 495 -1449 0 2
rlabel polysilicon 495 -1455 495 -1455 0 4
rlabel polysilicon 499 -1449 499 -1449 0 1
rlabel polysilicon 502 -1449 502 -1449 0 2
rlabel polysilicon 499 -1455 499 -1455 0 3
rlabel polysilicon 502 -1455 502 -1455 0 4
rlabel polysilicon 506 -1449 506 -1449 0 1
rlabel polysilicon 509 -1449 509 -1449 0 2
rlabel polysilicon 506 -1455 506 -1455 0 3
rlabel polysilicon 509 -1455 509 -1455 0 4
rlabel polysilicon 513 -1449 513 -1449 0 1
rlabel polysilicon 513 -1455 513 -1455 0 3
rlabel polysilicon 520 -1449 520 -1449 0 1
rlabel polysilicon 520 -1455 520 -1455 0 3
rlabel polysilicon 527 -1449 527 -1449 0 1
rlabel polysilicon 527 -1455 527 -1455 0 3
rlabel polysilicon 534 -1449 534 -1449 0 1
rlabel polysilicon 534 -1455 534 -1455 0 3
rlabel polysilicon 541 -1449 541 -1449 0 1
rlabel polysilicon 541 -1455 541 -1455 0 3
rlabel polysilicon 548 -1449 548 -1449 0 1
rlabel polysilicon 548 -1455 548 -1455 0 3
rlabel polysilicon 551 -1455 551 -1455 0 4
rlabel polysilicon 555 -1449 555 -1449 0 1
rlabel polysilicon 555 -1455 555 -1455 0 3
rlabel polysilicon 562 -1449 562 -1449 0 1
rlabel polysilicon 562 -1455 562 -1455 0 3
rlabel polysilicon 569 -1449 569 -1449 0 1
rlabel polysilicon 569 -1455 569 -1455 0 3
rlabel polysilicon 576 -1449 576 -1449 0 1
rlabel polysilicon 579 -1449 579 -1449 0 2
rlabel polysilicon 576 -1455 576 -1455 0 3
rlabel polysilicon 579 -1455 579 -1455 0 4
rlabel polysilicon 583 -1449 583 -1449 0 1
rlabel polysilicon 583 -1455 583 -1455 0 3
rlabel polysilicon 590 -1449 590 -1449 0 1
rlabel polysilicon 590 -1455 590 -1455 0 3
rlabel polysilicon 600 -1449 600 -1449 0 2
rlabel polysilicon 600 -1455 600 -1455 0 4
rlabel polysilicon 604 -1449 604 -1449 0 1
rlabel polysilicon 604 -1455 604 -1455 0 3
rlabel polysilicon 611 -1449 611 -1449 0 1
rlabel polysilicon 611 -1455 611 -1455 0 3
rlabel polysilicon 614 -1455 614 -1455 0 4
rlabel polysilicon 618 -1449 618 -1449 0 1
rlabel polysilicon 618 -1455 618 -1455 0 3
rlabel polysilicon 625 -1449 625 -1449 0 1
rlabel polysilicon 625 -1455 625 -1455 0 3
rlabel polysilicon 632 -1449 632 -1449 0 1
rlabel polysilicon 632 -1455 632 -1455 0 3
rlabel polysilicon 639 -1449 639 -1449 0 1
rlabel polysilicon 639 -1455 639 -1455 0 3
rlabel polysilicon 646 -1449 646 -1449 0 1
rlabel polysilicon 646 -1455 646 -1455 0 3
rlabel polysilicon 653 -1449 653 -1449 0 1
rlabel polysilicon 653 -1455 653 -1455 0 3
rlabel polysilicon 660 -1449 660 -1449 0 1
rlabel polysilicon 660 -1455 660 -1455 0 3
rlabel polysilicon 667 -1449 667 -1449 0 1
rlabel polysilicon 667 -1455 667 -1455 0 3
rlabel polysilicon 674 -1449 674 -1449 0 1
rlabel polysilicon 674 -1455 674 -1455 0 3
rlabel polysilicon 681 -1449 681 -1449 0 1
rlabel polysilicon 681 -1455 681 -1455 0 3
rlabel polysilicon 688 -1449 688 -1449 0 1
rlabel polysilicon 691 -1449 691 -1449 0 2
rlabel polysilicon 691 -1455 691 -1455 0 4
rlabel polysilicon 695 -1449 695 -1449 0 1
rlabel polysilicon 695 -1455 695 -1455 0 3
rlabel polysilicon 702 -1449 702 -1449 0 1
rlabel polysilicon 705 -1455 705 -1455 0 4
rlabel polysilicon 709 -1449 709 -1449 0 1
rlabel polysilicon 709 -1455 709 -1455 0 3
rlabel polysilicon 716 -1449 716 -1449 0 1
rlabel polysilicon 716 -1455 716 -1455 0 3
rlabel polysilicon 723 -1449 723 -1449 0 1
rlabel polysilicon 723 -1455 723 -1455 0 3
rlabel polysilicon 730 -1449 730 -1449 0 1
rlabel polysilicon 730 -1455 730 -1455 0 3
rlabel polysilicon 737 -1449 737 -1449 0 1
rlabel polysilicon 737 -1455 737 -1455 0 3
rlabel polysilicon 744 -1449 744 -1449 0 1
rlabel polysilicon 744 -1455 744 -1455 0 3
rlabel polysilicon 747 -1455 747 -1455 0 4
rlabel polysilicon 751 -1449 751 -1449 0 1
rlabel polysilicon 751 -1455 751 -1455 0 3
rlabel polysilicon 758 -1449 758 -1449 0 1
rlabel polysilicon 758 -1455 758 -1455 0 3
rlabel polysilicon 765 -1449 765 -1449 0 1
rlabel polysilicon 765 -1455 765 -1455 0 3
rlabel polysilicon 772 -1449 772 -1449 0 1
rlabel polysilicon 772 -1455 772 -1455 0 3
rlabel polysilicon 779 -1449 779 -1449 0 1
rlabel polysilicon 779 -1455 779 -1455 0 3
rlabel polysilicon 786 -1449 786 -1449 0 1
rlabel polysilicon 786 -1455 786 -1455 0 3
rlabel polysilicon 793 -1449 793 -1449 0 1
rlabel polysilicon 793 -1455 793 -1455 0 3
rlabel polysilicon 800 -1449 800 -1449 0 1
rlabel polysilicon 800 -1455 800 -1455 0 3
rlabel polysilicon 807 -1449 807 -1449 0 1
rlabel polysilicon 807 -1455 807 -1455 0 3
rlabel polysilicon 814 -1449 814 -1449 0 1
rlabel polysilicon 814 -1455 814 -1455 0 3
rlabel polysilicon 821 -1449 821 -1449 0 1
rlabel polysilicon 821 -1455 821 -1455 0 3
rlabel polysilicon 828 -1449 828 -1449 0 1
rlabel polysilicon 828 -1455 828 -1455 0 3
rlabel polysilicon 835 -1449 835 -1449 0 1
rlabel polysilicon 835 -1455 835 -1455 0 3
rlabel polysilicon 842 -1449 842 -1449 0 1
rlabel polysilicon 842 -1455 842 -1455 0 3
rlabel polysilicon 849 -1449 849 -1449 0 1
rlabel polysilicon 849 -1455 849 -1455 0 3
rlabel polysilicon 856 -1449 856 -1449 0 1
rlabel polysilicon 856 -1455 856 -1455 0 3
rlabel polysilicon 859 -1455 859 -1455 0 4
rlabel polysilicon 863 -1449 863 -1449 0 1
rlabel polysilicon 863 -1455 863 -1455 0 3
rlabel polysilicon 870 -1449 870 -1449 0 1
rlabel polysilicon 870 -1455 870 -1455 0 3
rlabel polysilicon 877 -1449 877 -1449 0 1
rlabel polysilicon 877 -1455 877 -1455 0 3
rlabel polysilicon 884 -1449 884 -1449 0 1
rlabel polysilicon 884 -1455 884 -1455 0 3
rlabel polysilicon 891 -1449 891 -1449 0 1
rlabel polysilicon 891 -1455 891 -1455 0 3
rlabel polysilicon 898 -1449 898 -1449 0 1
rlabel polysilicon 898 -1455 898 -1455 0 3
rlabel polysilicon 905 -1449 905 -1449 0 1
rlabel polysilicon 905 -1455 905 -1455 0 3
rlabel polysilicon 912 -1449 912 -1449 0 1
rlabel polysilicon 912 -1455 912 -1455 0 3
rlabel polysilicon 919 -1449 919 -1449 0 1
rlabel polysilicon 919 -1455 919 -1455 0 3
rlabel polysilicon 926 -1449 926 -1449 0 1
rlabel polysilicon 926 -1455 926 -1455 0 3
rlabel polysilicon 933 -1449 933 -1449 0 1
rlabel polysilicon 933 -1455 933 -1455 0 3
rlabel polysilicon 940 -1449 940 -1449 0 1
rlabel polysilicon 940 -1455 940 -1455 0 3
rlabel polysilicon 947 -1449 947 -1449 0 1
rlabel polysilicon 947 -1455 947 -1455 0 3
rlabel polysilicon 954 -1449 954 -1449 0 1
rlabel polysilicon 954 -1455 954 -1455 0 3
rlabel polysilicon 961 -1449 961 -1449 0 1
rlabel polysilicon 961 -1455 961 -1455 0 3
rlabel polysilicon 968 -1449 968 -1449 0 1
rlabel polysilicon 968 -1455 968 -1455 0 3
rlabel polysilicon 975 -1449 975 -1449 0 1
rlabel polysilicon 975 -1455 975 -1455 0 3
rlabel polysilicon 982 -1449 982 -1449 0 1
rlabel polysilicon 982 -1455 982 -1455 0 3
rlabel polysilicon 989 -1449 989 -1449 0 1
rlabel polysilicon 989 -1455 989 -1455 0 3
rlabel polysilicon 996 -1449 996 -1449 0 1
rlabel polysilicon 996 -1455 996 -1455 0 3
rlabel polysilicon 1003 -1449 1003 -1449 0 1
rlabel polysilicon 1003 -1455 1003 -1455 0 3
rlabel polysilicon 1010 -1449 1010 -1449 0 1
rlabel polysilicon 1010 -1455 1010 -1455 0 3
rlabel polysilicon 1017 -1449 1017 -1449 0 1
rlabel polysilicon 1017 -1455 1017 -1455 0 3
rlabel polysilicon 1024 -1449 1024 -1449 0 1
rlabel polysilicon 1024 -1455 1024 -1455 0 3
rlabel polysilicon 1031 -1449 1031 -1449 0 1
rlabel polysilicon 1031 -1455 1031 -1455 0 3
rlabel polysilicon 1038 -1449 1038 -1449 0 1
rlabel polysilicon 1038 -1455 1038 -1455 0 3
rlabel polysilicon 1045 -1449 1045 -1449 0 1
rlabel polysilicon 1045 -1455 1045 -1455 0 3
rlabel polysilicon 1052 -1449 1052 -1449 0 1
rlabel polysilicon 1052 -1455 1052 -1455 0 3
rlabel polysilicon 1062 -1449 1062 -1449 0 2
rlabel polysilicon 1062 -1455 1062 -1455 0 4
rlabel polysilicon 1066 -1449 1066 -1449 0 1
rlabel polysilicon 1066 -1455 1066 -1455 0 3
rlabel polysilicon 1073 -1449 1073 -1449 0 1
rlabel polysilicon 1073 -1455 1073 -1455 0 3
rlabel polysilicon 1080 -1449 1080 -1449 0 1
rlabel polysilicon 1080 -1455 1080 -1455 0 3
rlabel polysilicon 1087 -1449 1087 -1449 0 1
rlabel polysilicon 1094 -1449 1094 -1449 0 1
rlabel polysilicon 1094 -1455 1094 -1455 0 3
rlabel polysilicon 1108 -1449 1108 -1449 0 1
rlabel polysilicon 1108 -1455 1108 -1455 0 3
rlabel polysilicon 2 -1540 2 -1540 0 1
rlabel polysilicon 2 -1546 2 -1546 0 3
rlabel polysilicon 9 -1540 9 -1540 0 1
rlabel polysilicon 9 -1546 9 -1546 0 3
rlabel polysilicon 16 -1540 16 -1540 0 1
rlabel polysilicon 16 -1546 16 -1546 0 3
rlabel polysilicon 23 -1540 23 -1540 0 1
rlabel polysilicon 23 -1546 23 -1546 0 3
rlabel polysilicon 30 -1540 30 -1540 0 1
rlabel polysilicon 33 -1540 33 -1540 0 2
rlabel polysilicon 33 -1546 33 -1546 0 4
rlabel polysilicon 37 -1540 37 -1540 0 1
rlabel polysilicon 37 -1546 37 -1546 0 3
rlabel polysilicon 40 -1546 40 -1546 0 4
rlabel polysilicon 44 -1540 44 -1540 0 1
rlabel polysilicon 44 -1546 44 -1546 0 3
rlabel polysilicon 51 -1540 51 -1540 0 1
rlabel polysilicon 51 -1546 51 -1546 0 3
rlabel polysilicon 58 -1540 58 -1540 0 1
rlabel polysilicon 58 -1546 58 -1546 0 3
rlabel polysilicon 65 -1540 65 -1540 0 1
rlabel polysilicon 65 -1546 65 -1546 0 3
rlabel polysilicon 72 -1540 72 -1540 0 1
rlabel polysilicon 72 -1546 72 -1546 0 3
rlabel polysilicon 79 -1540 79 -1540 0 1
rlabel polysilicon 79 -1546 79 -1546 0 3
rlabel polysilicon 86 -1540 86 -1540 0 1
rlabel polysilicon 86 -1546 86 -1546 0 3
rlabel polysilicon 93 -1540 93 -1540 0 1
rlabel polysilicon 96 -1540 96 -1540 0 2
rlabel polysilicon 100 -1540 100 -1540 0 1
rlabel polysilicon 100 -1546 100 -1546 0 3
rlabel polysilicon 107 -1540 107 -1540 0 1
rlabel polysilicon 107 -1546 107 -1546 0 3
rlabel polysilicon 114 -1540 114 -1540 0 1
rlabel polysilicon 114 -1546 114 -1546 0 3
rlabel polysilicon 121 -1540 121 -1540 0 1
rlabel polysilicon 121 -1546 121 -1546 0 3
rlabel polysilicon 128 -1540 128 -1540 0 1
rlabel polysilicon 128 -1546 128 -1546 0 3
rlabel polysilicon 135 -1540 135 -1540 0 1
rlabel polysilicon 135 -1546 135 -1546 0 3
rlabel polysilicon 145 -1540 145 -1540 0 2
rlabel polysilicon 145 -1546 145 -1546 0 4
rlabel polysilicon 149 -1540 149 -1540 0 1
rlabel polysilicon 149 -1546 149 -1546 0 3
rlabel polysilicon 156 -1540 156 -1540 0 1
rlabel polysilicon 156 -1546 156 -1546 0 3
rlabel polysilicon 163 -1540 163 -1540 0 1
rlabel polysilicon 166 -1540 166 -1540 0 2
rlabel polysilicon 163 -1546 163 -1546 0 3
rlabel polysilicon 166 -1546 166 -1546 0 4
rlabel polysilicon 170 -1540 170 -1540 0 1
rlabel polysilicon 170 -1546 170 -1546 0 3
rlabel polysilicon 177 -1540 177 -1540 0 1
rlabel polysilicon 180 -1546 180 -1546 0 4
rlabel polysilicon 184 -1540 184 -1540 0 1
rlabel polysilicon 184 -1546 184 -1546 0 3
rlabel polysilicon 191 -1540 191 -1540 0 1
rlabel polysilicon 191 -1546 191 -1546 0 3
rlabel polysilicon 198 -1540 198 -1540 0 1
rlabel polysilicon 198 -1546 198 -1546 0 3
rlabel polysilicon 205 -1540 205 -1540 0 1
rlabel polysilicon 208 -1546 208 -1546 0 4
rlabel polysilicon 212 -1540 212 -1540 0 1
rlabel polysilicon 215 -1540 215 -1540 0 2
rlabel polysilicon 212 -1546 212 -1546 0 3
rlabel polysilicon 219 -1540 219 -1540 0 1
rlabel polysilicon 219 -1546 219 -1546 0 3
rlabel polysilicon 226 -1540 226 -1540 0 1
rlabel polysilicon 226 -1546 226 -1546 0 3
rlabel polysilicon 233 -1540 233 -1540 0 1
rlabel polysilicon 233 -1546 233 -1546 0 3
rlabel polysilicon 240 -1540 240 -1540 0 1
rlabel polysilicon 240 -1546 240 -1546 0 3
rlabel polysilicon 247 -1540 247 -1540 0 1
rlabel polysilicon 250 -1546 250 -1546 0 4
rlabel polysilicon 254 -1540 254 -1540 0 1
rlabel polysilicon 254 -1546 254 -1546 0 3
rlabel polysilicon 261 -1540 261 -1540 0 1
rlabel polysilicon 261 -1546 261 -1546 0 3
rlabel polysilicon 268 -1540 268 -1540 0 1
rlabel polysilicon 268 -1546 268 -1546 0 3
rlabel polysilicon 278 -1546 278 -1546 0 4
rlabel polysilicon 282 -1540 282 -1540 0 1
rlabel polysilicon 282 -1546 282 -1546 0 3
rlabel polysilicon 289 -1540 289 -1540 0 1
rlabel polysilicon 292 -1540 292 -1540 0 2
rlabel polysilicon 292 -1546 292 -1546 0 4
rlabel polysilicon 296 -1540 296 -1540 0 1
rlabel polysilicon 296 -1546 296 -1546 0 3
rlabel polysilicon 303 -1540 303 -1540 0 1
rlabel polysilicon 303 -1546 303 -1546 0 3
rlabel polysilicon 310 -1540 310 -1540 0 1
rlabel polysilicon 310 -1546 310 -1546 0 3
rlabel polysilicon 317 -1540 317 -1540 0 1
rlabel polysilicon 317 -1546 317 -1546 0 3
rlabel polysilicon 324 -1540 324 -1540 0 1
rlabel polysilicon 327 -1540 327 -1540 0 2
rlabel polysilicon 324 -1546 324 -1546 0 3
rlabel polysilicon 331 -1540 331 -1540 0 1
rlabel polysilicon 331 -1546 331 -1546 0 3
rlabel polysilicon 338 -1540 338 -1540 0 1
rlabel polysilicon 338 -1546 338 -1546 0 3
rlabel polysilicon 345 -1540 345 -1540 0 1
rlabel polysilicon 345 -1546 345 -1546 0 3
rlabel polysilicon 352 -1540 352 -1540 0 1
rlabel polysilicon 352 -1546 352 -1546 0 3
rlabel polysilicon 359 -1540 359 -1540 0 1
rlabel polysilicon 359 -1546 359 -1546 0 3
rlabel polysilicon 366 -1540 366 -1540 0 1
rlabel polysilicon 366 -1546 366 -1546 0 3
rlabel polysilicon 373 -1540 373 -1540 0 1
rlabel polysilicon 373 -1546 373 -1546 0 3
rlabel polysilicon 380 -1540 380 -1540 0 1
rlabel polysilicon 380 -1546 380 -1546 0 3
rlabel polysilicon 387 -1540 387 -1540 0 1
rlabel polysilicon 387 -1546 387 -1546 0 3
rlabel polysilicon 394 -1540 394 -1540 0 1
rlabel polysilicon 394 -1546 394 -1546 0 3
rlabel polysilicon 401 -1540 401 -1540 0 1
rlabel polysilicon 401 -1546 401 -1546 0 3
rlabel polysilicon 408 -1540 408 -1540 0 1
rlabel polysilicon 408 -1546 408 -1546 0 3
rlabel polysilicon 415 -1540 415 -1540 0 1
rlabel polysilicon 415 -1546 415 -1546 0 3
rlabel polysilicon 422 -1540 422 -1540 0 1
rlabel polysilicon 422 -1546 422 -1546 0 3
rlabel polysilicon 429 -1540 429 -1540 0 1
rlabel polysilicon 429 -1546 429 -1546 0 3
rlabel polysilicon 436 -1540 436 -1540 0 1
rlabel polysilicon 436 -1546 436 -1546 0 3
rlabel polysilicon 443 -1540 443 -1540 0 1
rlabel polysilicon 443 -1546 443 -1546 0 3
rlabel polysilicon 450 -1540 450 -1540 0 1
rlabel polysilicon 450 -1546 450 -1546 0 3
rlabel polysilicon 457 -1540 457 -1540 0 1
rlabel polysilicon 457 -1546 457 -1546 0 3
rlabel polysilicon 460 -1546 460 -1546 0 4
rlabel polysilicon 467 -1540 467 -1540 0 2
rlabel polysilicon 464 -1546 464 -1546 0 3
rlabel polysilicon 467 -1546 467 -1546 0 4
rlabel polysilicon 471 -1546 471 -1546 0 3
rlabel polysilicon 478 -1540 478 -1540 0 1
rlabel polysilicon 481 -1540 481 -1540 0 2
rlabel polysilicon 478 -1546 478 -1546 0 3
rlabel polysilicon 485 -1540 485 -1540 0 1
rlabel polysilicon 485 -1546 485 -1546 0 3
rlabel polysilicon 492 -1540 492 -1540 0 1
rlabel polysilicon 492 -1546 492 -1546 0 3
rlabel polysilicon 499 -1540 499 -1540 0 1
rlabel polysilicon 499 -1546 499 -1546 0 3
rlabel polysilicon 506 -1540 506 -1540 0 1
rlabel polysilicon 506 -1546 506 -1546 0 3
rlabel polysilicon 513 -1540 513 -1540 0 1
rlabel polysilicon 516 -1540 516 -1540 0 2
rlabel polysilicon 516 -1546 516 -1546 0 4
rlabel polysilicon 523 -1540 523 -1540 0 2
rlabel polysilicon 520 -1546 520 -1546 0 3
rlabel polysilicon 523 -1546 523 -1546 0 4
rlabel polysilicon 527 -1540 527 -1540 0 1
rlabel polysilicon 527 -1546 527 -1546 0 3
rlabel polysilicon 534 -1540 534 -1540 0 1
rlabel polysilicon 537 -1540 537 -1540 0 2
rlabel polysilicon 534 -1546 534 -1546 0 3
rlabel polysilicon 537 -1546 537 -1546 0 4
rlabel polysilicon 541 -1540 541 -1540 0 1
rlabel polysilicon 541 -1546 541 -1546 0 3
rlabel polysilicon 548 -1540 548 -1540 0 1
rlabel polysilicon 548 -1546 548 -1546 0 3
rlabel polysilicon 555 -1540 555 -1540 0 1
rlabel polysilicon 555 -1546 555 -1546 0 3
rlabel polysilicon 562 -1540 562 -1540 0 1
rlabel polysilicon 562 -1546 562 -1546 0 3
rlabel polysilicon 565 -1546 565 -1546 0 4
rlabel polysilicon 569 -1540 569 -1540 0 1
rlabel polysilicon 569 -1546 569 -1546 0 3
rlabel polysilicon 576 -1540 576 -1540 0 1
rlabel polysilicon 576 -1546 576 -1546 0 3
rlabel polysilicon 583 -1540 583 -1540 0 1
rlabel polysilicon 583 -1546 583 -1546 0 3
rlabel polysilicon 590 -1540 590 -1540 0 1
rlabel polysilicon 590 -1546 590 -1546 0 3
rlabel polysilicon 593 -1546 593 -1546 0 4
rlabel polysilicon 597 -1540 597 -1540 0 1
rlabel polysilicon 597 -1546 597 -1546 0 3
rlabel polysilicon 604 -1540 604 -1540 0 1
rlabel polysilicon 604 -1546 604 -1546 0 3
rlabel polysilicon 611 -1540 611 -1540 0 1
rlabel polysilicon 611 -1546 611 -1546 0 3
rlabel polysilicon 618 -1540 618 -1540 0 1
rlabel polysilicon 618 -1546 618 -1546 0 3
rlabel polysilicon 625 -1540 625 -1540 0 1
rlabel polysilicon 625 -1546 625 -1546 0 3
rlabel polysilicon 632 -1540 632 -1540 0 1
rlabel polysilicon 632 -1546 632 -1546 0 3
rlabel polysilicon 639 -1540 639 -1540 0 1
rlabel polysilicon 639 -1546 639 -1546 0 3
rlabel polysilicon 646 -1540 646 -1540 0 1
rlabel polysilicon 646 -1546 646 -1546 0 3
rlabel polysilicon 653 -1540 653 -1540 0 1
rlabel polysilicon 653 -1546 653 -1546 0 3
rlabel polysilicon 663 -1540 663 -1540 0 2
rlabel polysilicon 663 -1546 663 -1546 0 4
rlabel polysilicon 670 -1540 670 -1540 0 2
rlabel polysilicon 667 -1546 667 -1546 0 3
rlabel polysilicon 670 -1546 670 -1546 0 4
rlabel polysilicon 674 -1540 674 -1540 0 1
rlabel polysilicon 677 -1540 677 -1540 0 2
rlabel polysilicon 674 -1546 674 -1546 0 3
rlabel polysilicon 677 -1546 677 -1546 0 4
rlabel polysilicon 681 -1540 681 -1540 0 1
rlabel polysilicon 681 -1546 681 -1546 0 3
rlabel polysilicon 688 -1540 688 -1540 0 1
rlabel polysilicon 691 -1540 691 -1540 0 2
rlabel polysilicon 695 -1540 695 -1540 0 1
rlabel polysilicon 695 -1546 695 -1546 0 3
rlabel polysilicon 702 -1540 702 -1540 0 1
rlabel polysilicon 702 -1546 702 -1546 0 3
rlabel polysilicon 709 -1540 709 -1540 0 1
rlabel polysilicon 709 -1546 709 -1546 0 3
rlabel polysilicon 716 -1540 716 -1540 0 1
rlabel polysilicon 716 -1546 716 -1546 0 3
rlabel polysilicon 723 -1540 723 -1540 0 1
rlabel polysilicon 723 -1546 723 -1546 0 3
rlabel polysilicon 730 -1540 730 -1540 0 1
rlabel polysilicon 730 -1546 730 -1546 0 3
rlabel polysilicon 737 -1540 737 -1540 0 1
rlabel polysilicon 737 -1546 737 -1546 0 3
rlabel polysilicon 744 -1540 744 -1540 0 1
rlabel polysilicon 744 -1546 744 -1546 0 3
rlabel polysilicon 751 -1540 751 -1540 0 1
rlabel polysilicon 751 -1546 751 -1546 0 3
rlabel polysilicon 758 -1540 758 -1540 0 1
rlabel polysilicon 758 -1546 758 -1546 0 3
rlabel polysilicon 765 -1540 765 -1540 0 1
rlabel polysilicon 765 -1546 765 -1546 0 3
rlabel polysilicon 772 -1546 772 -1546 0 3
rlabel polysilicon 775 -1546 775 -1546 0 4
rlabel polysilicon 779 -1540 779 -1540 0 1
rlabel polysilicon 779 -1546 779 -1546 0 3
rlabel polysilicon 786 -1540 786 -1540 0 1
rlabel polysilicon 786 -1546 786 -1546 0 3
rlabel polysilicon 793 -1540 793 -1540 0 1
rlabel polysilicon 793 -1546 793 -1546 0 3
rlabel polysilicon 800 -1540 800 -1540 0 1
rlabel polysilicon 800 -1546 800 -1546 0 3
rlabel polysilicon 807 -1540 807 -1540 0 1
rlabel polysilicon 807 -1546 807 -1546 0 3
rlabel polysilicon 814 -1540 814 -1540 0 1
rlabel polysilicon 814 -1546 814 -1546 0 3
rlabel polysilicon 821 -1540 821 -1540 0 1
rlabel polysilicon 821 -1546 821 -1546 0 3
rlabel polysilicon 828 -1540 828 -1540 0 1
rlabel polysilicon 828 -1546 828 -1546 0 3
rlabel polysilicon 835 -1540 835 -1540 0 1
rlabel polysilicon 835 -1546 835 -1546 0 3
rlabel polysilicon 842 -1540 842 -1540 0 1
rlabel polysilicon 842 -1546 842 -1546 0 3
rlabel polysilicon 849 -1540 849 -1540 0 1
rlabel polysilicon 849 -1546 849 -1546 0 3
rlabel polysilicon 856 -1540 856 -1540 0 1
rlabel polysilicon 856 -1546 856 -1546 0 3
rlabel polysilicon 863 -1540 863 -1540 0 1
rlabel polysilicon 863 -1546 863 -1546 0 3
rlabel polysilicon 870 -1540 870 -1540 0 1
rlabel polysilicon 870 -1546 870 -1546 0 3
rlabel polysilicon 877 -1540 877 -1540 0 1
rlabel polysilicon 877 -1546 877 -1546 0 3
rlabel polysilicon 884 -1540 884 -1540 0 1
rlabel polysilicon 884 -1546 884 -1546 0 3
rlabel polysilicon 891 -1540 891 -1540 0 1
rlabel polysilicon 891 -1546 891 -1546 0 3
rlabel polysilicon 898 -1540 898 -1540 0 1
rlabel polysilicon 898 -1546 898 -1546 0 3
rlabel polysilicon 905 -1540 905 -1540 0 1
rlabel polysilicon 905 -1546 905 -1546 0 3
rlabel polysilicon 912 -1540 912 -1540 0 1
rlabel polysilicon 912 -1546 912 -1546 0 3
rlabel polysilicon 919 -1540 919 -1540 0 1
rlabel polysilicon 919 -1546 919 -1546 0 3
rlabel polysilicon 926 -1540 926 -1540 0 1
rlabel polysilicon 926 -1546 926 -1546 0 3
rlabel polysilicon 933 -1540 933 -1540 0 1
rlabel polysilicon 933 -1546 933 -1546 0 3
rlabel polysilicon 940 -1540 940 -1540 0 1
rlabel polysilicon 940 -1546 940 -1546 0 3
rlabel polysilicon 947 -1540 947 -1540 0 1
rlabel polysilicon 947 -1546 947 -1546 0 3
rlabel polysilicon 954 -1540 954 -1540 0 1
rlabel polysilicon 954 -1546 954 -1546 0 3
rlabel polysilicon 961 -1540 961 -1540 0 1
rlabel polysilicon 961 -1546 961 -1546 0 3
rlabel polysilicon 968 -1540 968 -1540 0 1
rlabel polysilicon 968 -1546 968 -1546 0 3
rlabel polysilicon 975 -1540 975 -1540 0 1
rlabel polysilicon 975 -1546 975 -1546 0 3
rlabel polysilicon 982 -1540 982 -1540 0 1
rlabel polysilicon 982 -1546 982 -1546 0 3
rlabel polysilicon 989 -1540 989 -1540 0 1
rlabel polysilicon 989 -1546 989 -1546 0 3
rlabel polysilicon 996 -1540 996 -1540 0 1
rlabel polysilicon 996 -1546 996 -1546 0 3
rlabel polysilicon 1003 -1540 1003 -1540 0 1
rlabel polysilicon 1003 -1546 1003 -1546 0 3
rlabel polysilicon 1010 -1540 1010 -1540 0 1
rlabel polysilicon 1017 -1540 1017 -1540 0 1
rlabel polysilicon 1017 -1546 1017 -1546 0 3
rlabel polysilicon 1024 -1540 1024 -1540 0 1
rlabel polysilicon 1024 -1546 1024 -1546 0 3
rlabel polysilicon 1031 -1540 1031 -1540 0 1
rlabel polysilicon 1031 -1546 1031 -1546 0 3
rlabel polysilicon 1034 -1546 1034 -1546 0 4
rlabel polysilicon 1038 -1540 1038 -1540 0 1
rlabel polysilicon 1038 -1546 1038 -1546 0 3
rlabel polysilicon 1045 -1540 1045 -1540 0 1
rlabel polysilicon 1045 -1546 1045 -1546 0 3
rlabel polysilicon 1059 -1540 1059 -1540 0 1
rlabel polysilicon 1059 -1546 1059 -1546 0 3
rlabel polysilicon 1073 -1540 1073 -1540 0 1
rlabel polysilicon 1073 -1546 1073 -1546 0 3
rlabel polysilicon 1094 -1540 1094 -1540 0 1
rlabel polysilicon 1094 -1546 1094 -1546 0 3
rlabel polysilicon 5 -1629 5 -1629 0 2
rlabel polysilicon 9 -1629 9 -1629 0 1
rlabel polysilicon 9 -1635 9 -1635 0 3
rlabel polysilicon 16 -1629 16 -1629 0 1
rlabel polysilicon 16 -1635 16 -1635 0 3
rlabel polysilicon 23 -1629 23 -1629 0 1
rlabel polysilicon 23 -1635 23 -1635 0 3
rlabel polysilicon 30 -1629 30 -1629 0 1
rlabel polysilicon 30 -1635 30 -1635 0 3
rlabel polysilicon 37 -1629 37 -1629 0 1
rlabel polysilicon 37 -1635 37 -1635 0 3
rlabel polysilicon 44 -1629 44 -1629 0 1
rlabel polysilicon 44 -1635 44 -1635 0 3
rlabel polysilicon 51 -1629 51 -1629 0 1
rlabel polysilicon 51 -1635 51 -1635 0 3
rlabel polysilicon 58 -1629 58 -1629 0 1
rlabel polysilicon 58 -1635 58 -1635 0 3
rlabel polysilicon 61 -1635 61 -1635 0 4
rlabel polysilicon 65 -1629 65 -1629 0 1
rlabel polysilicon 65 -1635 65 -1635 0 3
rlabel polysilicon 72 -1629 72 -1629 0 1
rlabel polysilicon 72 -1635 72 -1635 0 3
rlabel polysilicon 79 -1629 79 -1629 0 1
rlabel polysilicon 82 -1629 82 -1629 0 2
rlabel polysilicon 82 -1635 82 -1635 0 4
rlabel polysilicon 86 -1629 86 -1629 0 1
rlabel polysilicon 86 -1635 86 -1635 0 3
rlabel polysilicon 93 -1629 93 -1629 0 1
rlabel polysilicon 96 -1629 96 -1629 0 2
rlabel polysilicon 96 -1635 96 -1635 0 4
rlabel polysilicon 100 -1629 100 -1629 0 1
rlabel polysilicon 100 -1635 100 -1635 0 3
rlabel polysilicon 107 -1629 107 -1629 0 1
rlabel polysilicon 107 -1635 107 -1635 0 3
rlabel polysilicon 114 -1629 114 -1629 0 1
rlabel polysilicon 114 -1635 114 -1635 0 3
rlabel polysilicon 121 -1629 121 -1629 0 1
rlabel polysilicon 121 -1635 121 -1635 0 3
rlabel polysilicon 128 -1629 128 -1629 0 1
rlabel polysilicon 128 -1635 128 -1635 0 3
rlabel polysilicon 135 -1635 135 -1635 0 3
rlabel polysilicon 138 -1635 138 -1635 0 4
rlabel polysilicon 145 -1629 145 -1629 0 2
rlabel polysilicon 142 -1635 142 -1635 0 3
rlabel polysilicon 149 -1629 149 -1629 0 1
rlabel polysilicon 149 -1635 149 -1635 0 3
rlabel polysilicon 156 -1629 156 -1629 0 1
rlabel polysilicon 156 -1635 156 -1635 0 3
rlabel polysilicon 163 -1629 163 -1629 0 1
rlabel polysilicon 163 -1635 163 -1635 0 3
rlabel polysilicon 170 -1629 170 -1629 0 1
rlabel polysilicon 170 -1635 170 -1635 0 3
rlabel polysilicon 177 -1629 177 -1629 0 1
rlabel polysilicon 177 -1635 177 -1635 0 3
rlabel polysilicon 184 -1635 184 -1635 0 3
rlabel polysilicon 187 -1635 187 -1635 0 4
rlabel polysilicon 191 -1629 191 -1629 0 1
rlabel polysilicon 191 -1635 191 -1635 0 3
rlabel polysilicon 201 -1629 201 -1629 0 2
rlabel polysilicon 198 -1635 198 -1635 0 3
rlabel polysilicon 201 -1635 201 -1635 0 4
rlabel polysilicon 205 -1629 205 -1629 0 1
rlabel polysilicon 205 -1635 205 -1635 0 3
rlabel polysilicon 212 -1629 212 -1629 0 1
rlabel polysilicon 212 -1635 212 -1635 0 3
rlabel polysilicon 222 -1629 222 -1629 0 2
rlabel polysilicon 222 -1635 222 -1635 0 4
rlabel polysilicon 226 -1629 226 -1629 0 1
rlabel polysilicon 229 -1629 229 -1629 0 2
rlabel polysilicon 226 -1635 226 -1635 0 3
rlabel polysilicon 233 -1629 233 -1629 0 1
rlabel polysilicon 233 -1635 233 -1635 0 3
rlabel polysilicon 240 -1629 240 -1629 0 1
rlabel polysilicon 240 -1635 240 -1635 0 3
rlabel polysilicon 247 -1629 247 -1629 0 1
rlabel polysilicon 254 -1629 254 -1629 0 1
rlabel polysilicon 254 -1635 254 -1635 0 3
rlabel polysilicon 261 -1629 261 -1629 0 1
rlabel polysilicon 261 -1635 261 -1635 0 3
rlabel polysilicon 268 -1629 268 -1629 0 1
rlabel polysilicon 268 -1635 268 -1635 0 3
rlabel polysilicon 275 -1629 275 -1629 0 1
rlabel polysilicon 275 -1635 275 -1635 0 3
rlabel polysilicon 282 -1629 282 -1629 0 1
rlabel polysilicon 282 -1635 282 -1635 0 3
rlabel polysilicon 289 -1629 289 -1629 0 1
rlabel polysilicon 289 -1635 289 -1635 0 3
rlabel polysilicon 296 -1629 296 -1629 0 1
rlabel polysilicon 296 -1635 296 -1635 0 3
rlabel polysilicon 303 -1635 303 -1635 0 3
rlabel polysilicon 306 -1635 306 -1635 0 4
rlabel polysilicon 310 -1629 310 -1629 0 1
rlabel polysilicon 310 -1635 310 -1635 0 3
rlabel polysilicon 317 -1629 317 -1629 0 1
rlabel polysilicon 317 -1635 317 -1635 0 3
rlabel polysilicon 327 -1629 327 -1629 0 2
rlabel polysilicon 324 -1635 324 -1635 0 3
rlabel polysilicon 327 -1635 327 -1635 0 4
rlabel polysilicon 331 -1629 331 -1629 0 1
rlabel polysilicon 331 -1635 331 -1635 0 3
rlabel polysilicon 338 -1629 338 -1629 0 1
rlabel polysilicon 338 -1635 338 -1635 0 3
rlabel polysilicon 345 -1629 345 -1629 0 1
rlabel polysilicon 345 -1635 345 -1635 0 3
rlabel polysilicon 352 -1629 352 -1629 0 1
rlabel polysilicon 355 -1629 355 -1629 0 2
rlabel polysilicon 355 -1635 355 -1635 0 4
rlabel polysilicon 359 -1629 359 -1629 0 1
rlabel polysilicon 359 -1635 359 -1635 0 3
rlabel polysilicon 366 -1629 366 -1629 0 1
rlabel polysilicon 366 -1635 366 -1635 0 3
rlabel polysilicon 373 -1629 373 -1629 0 1
rlabel polysilicon 376 -1629 376 -1629 0 2
rlabel polysilicon 373 -1635 373 -1635 0 3
rlabel polysilicon 376 -1635 376 -1635 0 4
rlabel polysilicon 380 -1629 380 -1629 0 1
rlabel polysilicon 380 -1635 380 -1635 0 3
rlabel polysilicon 387 -1629 387 -1629 0 1
rlabel polysilicon 387 -1635 387 -1635 0 3
rlabel polysilicon 394 -1629 394 -1629 0 1
rlabel polysilicon 394 -1635 394 -1635 0 3
rlabel polysilicon 401 -1629 401 -1629 0 1
rlabel polysilicon 401 -1635 401 -1635 0 3
rlabel polysilicon 408 -1629 408 -1629 0 1
rlabel polysilicon 408 -1635 408 -1635 0 3
rlabel polysilicon 415 -1629 415 -1629 0 1
rlabel polysilicon 415 -1635 415 -1635 0 3
rlabel polysilicon 425 -1629 425 -1629 0 2
rlabel polysilicon 422 -1635 422 -1635 0 3
rlabel polysilicon 425 -1635 425 -1635 0 4
rlabel polysilicon 429 -1629 429 -1629 0 1
rlabel polysilicon 429 -1635 429 -1635 0 3
rlabel polysilicon 436 -1629 436 -1629 0 1
rlabel polysilicon 436 -1635 436 -1635 0 3
rlabel polysilicon 443 -1629 443 -1629 0 1
rlabel polysilicon 446 -1635 446 -1635 0 4
rlabel polysilicon 450 -1629 450 -1629 0 1
rlabel polysilicon 450 -1635 450 -1635 0 3
rlabel polysilicon 457 -1629 457 -1629 0 1
rlabel polysilicon 457 -1635 457 -1635 0 3
rlabel polysilicon 460 -1635 460 -1635 0 4
rlabel polysilicon 464 -1629 464 -1629 0 1
rlabel polysilicon 464 -1635 464 -1635 0 3
rlabel polysilicon 471 -1629 471 -1629 0 1
rlabel polysilicon 471 -1635 471 -1635 0 3
rlabel polysilicon 478 -1629 478 -1629 0 1
rlabel polysilicon 478 -1635 478 -1635 0 3
rlabel polysilicon 485 -1629 485 -1629 0 1
rlabel polysilicon 485 -1635 485 -1635 0 3
rlabel polysilicon 492 -1629 492 -1629 0 1
rlabel polysilicon 492 -1635 492 -1635 0 3
rlabel polysilicon 499 -1629 499 -1629 0 1
rlabel polysilicon 499 -1635 499 -1635 0 3
rlabel polysilicon 506 -1629 506 -1629 0 1
rlabel polysilicon 506 -1635 506 -1635 0 3
rlabel polysilicon 513 -1629 513 -1629 0 1
rlabel polysilicon 513 -1635 513 -1635 0 3
rlabel polysilicon 520 -1629 520 -1629 0 1
rlabel polysilicon 520 -1635 520 -1635 0 3
rlabel polysilicon 527 -1629 527 -1629 0 1
rlabel polysilicon 527 -1635 527 -1635 0 3
rlabel polysilicon 534 -1629 534 -1629 0 1
rlabel polysilicon 537 -1635 537 -1635 0 4
rlabel polysilicon 541 -1629 541 -1629 0 1
rlabel polysilicon 541 -1635 541 -1635 0 3
rlabel polysilicon 548 -1629 548 -1629 0 1
rlabel polysilicon 548 -1635 548 -1635 0 3
rlabel polysilicon 555 -1629 555 -1629 0 1
rlabel polysilicon 555 -1635 555 -1635 0 3
rlabel polysilicon 562 -1629 562 -1629 0 1
rlabel polysilicon 562 -1635 562 -1635 0 3
rlabel polysilicon 569 -1629 569 -1629 0 1
rlabel polysilicon 569 -1635 569 -1635 0 3
rlabel polysilicon 572 -1635 572 -1635 0 4
rlabel polysilicon 576 -1629 576 -1629 0 1
rlabel polysilicon 576 -1635 576 -1635 0 3
rlabel polysilicon 586 -1629 586 -1629 0 2
rlabel polysilicon 583 -1635 583 -1635 0 3
rlabel polysilicon 590 -1629 590 -1629 0 1
rlabel polysilicon 590 -1635 590 -1635 0 3
rlabel polysilicon 597 -1629 597 -1629 0 1
rlabel polysilicon 597 -1635 597 -1635 0 3
rlabel polysilicon 604 -1629 604 -1629 0 1
rlabel polysilicon 604 -1635 604 -1635 0 3
rlabel polysilicon 611 -1629 611 -1629 0 1
rlabel polysilicon 614 -1629 614 -1629 0 2
rlabel polysilicon 614 -1635 614 -1635 0 4
rlabel polysilicon 618 -1629 618 -1629 0 1
rlabel polysilicon 618 -1635 618 -1635 0 3
rlabel polysilicon 625 -1629 625 -1629 0 1
rlabel polysilicon 625 -1635 625 -1635 0 3
rlabel polysilicon 632 -1629 632 -1629 0 1
rlabel polysilicon 635 -1629 635 -1629 0 2
rlabel polysilicon 632 -1635 632 -1635 0 3
rlabel polysilicon 639 -1629 639 -1629 0 1
rlabel polysilicon 639 -1635 639 -1635 0 3
rlabel polysilicon 646 -1629 646 -1629 0 1
rlabel polysilicon 646 -1635 646 -1635 0 3
rlabel polysilicon 653 -1629 653 -1629 0 1
rlabel polysilicon 653 -1635 653 -1635 0 3
rlabel polysilicon 660 -1629 660 -1629 0 1
rlabel polysilicon 660 -1635 660 -1635 0 3
rlabel polysilicon 667 -1629 667 -1629 0 1
rlabel polysilicon 667 -1635 667 -1635 0 3
rlabel polysilicon 674 -1629 674 -1629 0 1
rlabel polysilicon 677 -1629 677 -1629 0 2
rlabel polysilicon 674 -1635 674 -1635 0 3
rlabel polysilicon 677 -1635 677 -1635 0 4
rlabel polysilicon 684 -1629 684 -1629 0 2
rlabel polysilicon 681 -1635 681 -1635 0 3
rlabel polysilicon 684 -1635 684 -1635 0 4
rlabel polysilicon 688 -1629 688 -1629 0 1
rlabel polysilicon 688 -1635 688 -1635 0 3
rlabel polysilicon 695 -1629 695 -1629 0 1
rlabel polysilicon 695 -1635 695 -1635 0 3
rlabel polysilicon 702 -1629 702 -1629 0 1
rlabel polysilicon 702 -1635 702 -1635 0 3
rlabel polysilicon 709 -1629 709 -1629 0 1
rlabel polysilicon 709 -1635 709 -1635 0 3
rlabel polysilicon 716 -1629 716 -1629 0 1
rlabel polysilicon 716 -1635 716 -1635 0 3
rlabel polysilicon 723 -1629 723 -1629 0 1
rlabel polysilicon 723 -1635 723 -1635 0 3
rlabel polysilicon 730 -1629 730 -1629 0 1
rlabel polysilicon 730 -1635 730 -1635 0 3
rlabel polysilicon 737 -1629 737 -1629 0 1
rlabel polysilicon 737 -1635 737 -1635 0 3
rlabel polysilicon 744 -1629 744 -1629 0 1
rlabel polysilicon 744 -1635 744 -1635 0 3
rlabel polysilicon 751 -1629 751 -1629 0 1
rlabel polysilicon 751 -1635 751 -1635 0 3
rlabel polysilicon 758 -1629 758 -1629 0 1
rlabel polysilicon 758 -1635 758 -1635 0 3
rlabel polysilicon 765 -1629 765 -1629 0 1
rlabel polysilicon 765 -1635 765 -1635 0 3
rlabel polysilicon 772 -1629 772 -1629 0 1
rlabel polysilicon 772 -1635 772 -1635 0 3
rlabel polysilicon 779 -1629 779 -1629 0 1
rlabel polysilicon 779 -1635 779 -1635 0 3
rlabel polysilicon 786 -1629 786 -1629 0 1
rlabel polysilicon 786 -1635 786 -1635 0 3
rlabel polysilicon 793 -1629 793 -1629 0 1
rlabel polysilicon 793 -1635 793 -1635 0 3
rlabel polysilicon 800 -1629 800 -1629 0 1
rlabel polysilicon 800 -1635 800 -1635 0 3
rlabel polysilicon 807 -1629 807 -1629 0 1
rlabel polysilicon 807 -1635 807 -1635 0 3
rlabel polysilicon 814 -1629 814 -1629 0 1
rlabel polysilicon 814 -1635 814 -1635 0 3
rlabel polysilicon 821 -1629 821 -1629 0 1
rlabel polysilicon 821 -1635 821 -1635 0 3
rlabel polysilicon 828 -1629 828 -1629 0 1
rlabel polysilicon 828 -1635 828 -1635 0 3
rlabel polysilicon 835 -1629 835 -1629 0 1
rlabel polysilicon 835 -1635 835 -1635 0 3
rlabel polysilicon 842 -1629 842 -1629 0 1
rlabel polysilicon 842 -1635 842 -1635 0 3
rlabel polysilicon 849 -1629 849 -1629 0 1
rlabel polysilicon 849 -1635 849 -1635 0 3
rlabel polysilicon 856 -1629 856 -1629 0 1
rlabel polysilicon 859 -1629 859 -1629 0 2
rlabel polysilicon 856 -1635 856 -1635 0 3
rlabel polysilicon 863 -1629 863 -1629 0 1
rlabel polysilicon 863 -1635 863 -1635 0 3
rlabel polysilicon 870 -1629 870 -1629 0 1
rlabel polysilicon 870 -1635 870 -1635 0 3
rlabel polysilicon 877 -1629 877 -1629 0 1
rlabel polysilicon 877 -1635 877 -1635 0 3
rlabel polysilicon 884 -1629 884 -1629 0 1
rlabel polysilicon 884 -1635 884 -1635 0 3
rlabel polysilicon 891 -1629 891 -1629 0 1
rlabel polysilicon 891 -1635 891 -1635 0 3
rlabel polysilicon 898 -1629 898 -1629 0 1
rlabel polysilicon 898 -1635 898 -1635 0 3
rlabel polysilicon 905 -1629 905 -1629 0 1
rlabel polysilicon 905 -1635 905 -1635 0 3
rlabel polysilicon 912 -1629 912 -1629 0 1
rlabel polysilicon 912 -1635 912 -1635 0 3
rlabel polysilicon 919 -1629 919 -1629 0 1
rlabel polysilicon 919 -1635 919 -1635 0 3
rlabel polysilicon 926 -1629 926 -1629 0 1
rlabel polysilicon 926 -1635 926 -1635 0 3
rlabel polysilicon 933 -1629 933 -1629 0 1
rlabel polysilicon 933 -1635 933 -1635 0 3
rlabel polysilicon 940 -1629 940 -1629 0 1
rlabel polysilicon 940 -1635 940 -1635 0 3
rlabel polysilicon 947 -1629 947 -1629 0 1
rlabel polysilicon 947 -1635 947 -1635 0 3
rlabel polysilicon 954 -1629 954 -1629 0 1
rlabel polysilicon 954 -1635 954 -1635 0 3
rlabel polysilicon 961 -1629 961 -1629 0 1
rlabel polysilicon 961 -1635 961 -1635 0 3
rlabel polysilicon 968 -1629 968 -1629 0 1
rlabel polysilicon 968 -1635 968 -1635 0 3
rlabel polysilicon 975 -1629 975 -1629 0 1
rlabel polysilicon 975 -1635 975 -1635 0 3
rlabel polysilicon 982 -1629 982 -1629 0 1
rlabel polysilicon 982 -1635 982 -1635 0 3
rlabel polysilicon 989 -1629 989 -1629 0 1
rlabel polysilicon 989 -1635 989 -1635 0 3
rlabel polysilicon 996 -1629 996 -1629 0 1
rlabel polysilicon 996 -1635 996 -1635 0 3
rlabel polysilicon 1003 -1629 1003 -1629 0 1
rlabel polysilicon 1003 -1635 1003 -1635 0 3
rlabel polysilicon 1010 -1629 1010 -1629 0 1
rlabel polysilicon 1010 -1635 1010 -1635 0 3
rlabel polysilicon 1017 -1629 1017 -1629 0 1
rlabel polysilicon 1017 -1635 1017 -1635 0 3
rlabel polysilicon 1024 -1629 1024 -1629 0 1
rlabel polysilicon 1024 -1635 1024 -1635 0 3
rlabel polysilicon 1031 -1629 1031 -1629 0 1
rlabel polysilicon 1031 -1635 1031 -1635 0 3
rlabel polysilicon 1038 -1629 1038 -1629 0 1
rlabel polysilicon 1038 -1635 1038 -1635 0 3
rlabel polysilicon 1045 -1629 1045 -1629 0 1
rlabel polysilicon 1045 -1635 1045 -1635 0 3
rlabel polysilicon 1052 -1629 1052 -1629 0 1
rlabel polysilicon 1052 -1635 1052 -1635 0 3
rlabel polysilicon 1062 -1629 1062 -1629 0 2
rlabel polysilicon 1059 -1635 1059 -1635 0 3
rlabel polysilicon 1062 -1635 1062 -1635 0 4
rlabel polysilicon 1069 -1629 1069 -1629 0 2
rlabel polysilicon 1069 -1635 1069 -1635 0 4
rlabel polysilicon 1073 -1629 1073 -1629 0 1
rlabel polysilicon 1073 -1635 1073 -1635 0 3
rlabel polysilicon 1080 -1629 1080 -1629 0 1
rlabel polysilicon 1080 -1635 1080 -1635 0 3
rlabel polysilicon 1087 -1629 1087 -1629 0 1
rlabel polysilicon 1087 -1635 1087 -1635 0 3
rlabel polysilicon 1094 -1629 1094 -1629 0 1
rlabel polysilicon 1094 -1635 1094 -1635 0 3
rlabel polysilicon 1101 -1629 1101 -1629 0 1
rlabel polysilicon 1101 -1635 1101 -1635 0 3
rlabel polysilicon 1108 -1629 1108 -1629 0 1
rlabel polysilicon 1108 -1635 1108 -1635 0 3
rlabel polysilicon 1115 -1629 1115 -1629 0 1
rlabel polysilicon 1115 -1635 1115 -1635 0 3
rlabel polysilicon 23 -1714 23 -1714 0 1
rlabel polysilicon 23 -1720 23 -1720 0 3
rlabel polysilicon 30 -1714 30 -1714 0 1
rlabel polysilicon 30 -1720 30 -1720 0 3
rlabel polysilicon 37 -1714 37 -1714 0 1
rlabel polysilicon 37 -1720 37 -1720 0 3
rlabel polysilicon 44 -1714 44 -1714 0 1
rlabel polysilicon 44 -1720 44 -1720 0 3
rlabel polysilicon 51 -1714 51 -1714 0 1
rlabel polysilicon 54 -1714 54 -1714 0 2
rlabel polysilicon 58 -1714 58 -1714 0 1
rlabel polysilicon 58 -1720 58 -1720 0 3
rlabel polysilicon 65 -1714 65 -1714 0 1
rlabel polysilicon 68 -1714 68 -1714 0 2
rlabel polysilicon 65 -1720 65 -1720 0 3
rlabel polysilicon 72 -1714 72 -1714 0 1
rlabel polysilicon 72 -1720 72 -1720 0 3
rlabel polysilicon 79 -1714 79 -1714 0 1
rlabel polysilicon 79 -1720 79 -1720 0 3
rlabel polysilicon 86 -1714 86 -1714 0 1
rlabel polysilicon 86 -1720 86 -1720 0 3
rlabel polysilicon 93 -1714 93 -1714 0 1
rlabel polysilicon 93 -1720 93 -1720 0 3
rlabel polysilicon 100 -1714 100 -1714 0 1
rlabel polysilicon 100 -1720 100 -1720 0 3
rlabel polysilicon 107 -1714 107 -1714 0 1
rlabel polysilicon 107 -1720 107 -1720 0 3
rlabel polysilicon 114 -1714 114 -1714 0 1
rlabel polysilicon 114 -1720 114 -1720 0 3
rlabel polysilicon 121 -1714 121 -1714 0 1
rlabel polysilicon 121 -1720 121 -1720 0 3
rlabel polysilicon 128 -1714 128 -1714 0 1
rlabel polysilicon 128 -1720 128 -1720 0 3
rlabel polysilicon 135 -1714 135 -1714 0 1
rlabel polysilicon 135 -1720 135 -1720 0 3
rlabel polysilicon 142 -1714 142 -1714 0 1
rlabel polysilicon 142 -1720 142 -1720 0 3
rlabel polysilicon 149 -1714 149 -1714 0 1
rlabel polysilicon 149 -1720 149 -1720 0 3
rlabel polysilicon 159 -1714 159 -1714 0 2
rlabel polysilicon 156 -1720 156 -1720 0 3
rlabel polysilicon 159 -1720 159 -1720 0 4
rlabel polysilicon 163 -1714 163 -1714 0 1
rlabel polysilicon 163 -1720 163 -1720 0 3
rlabel polysilicon 170 -1714 170 -1714 0 1
rlabel polysilicon 170 -1720 170 -1720 0 3
rlabel polysilicon 177 -1714 177 -1714 0 1
rlabel polysilicon 177 -1720 177 -1720 0 3
rlabel polysilicon 184 -1714 184 -1714 0 1
rlabel polysilicon 184 -1720 184 -1720 0 3
rlabel polysilicon 191 -1714 191 -1714 0 1
rlabel polysilicon 191 -1720 191 -1720 0 3
rlabel polysilicon 198 -1714 198 -1714 0 1
rlabel polysilicon 198 -1720 198 -1720 0 3
rlabel polysilicon 205 -1714 205 -1714 0 1
rlabel polysilicon 205 -1720 205 -1720 0 3
rlabel polysilicon 212 -1714 212 -1714 0 1
rlabel polysilicon 212 -1720 212 -1720 0 3
rlabel polysilicon 222 -1720 222 -1720 0 4
rlabel polysilicon 226 -1714 226 -1714 0 1
rlabel polysilicon 226 -1720 226 -1720 0 3
rlabel polysilicon 233 -1714 233 -1714 0 1
rlabel polysilicon 233 -1720 233 -1720 0 3
rlabel polysilicon 240 -1714 240 -1714 0 1
rlabel polysilicon 240 -1720 240 -1720 0 3
rlabel polysilicon 247 -1714 247 -1714 0 1
rlabel polysilicon 247 -1720 247 -1720 0 3
rlabel polysilicon 254 -1714 254 -1714 0 1
rlabel polysilicon 254 -1720 254 -1720 0 3
rlabel polysilicon 261 -1714 261 -1714 0 1
rlabel polysilicon 261 -1720 261 -1720 0 3
rlabel polysilicon 268 -1714 268 -1714 0 1
rlabel polysilicon 268 -1720 268 -1720 0 3
rlabel polysilicon 275 -1714 275 -1714 0 1
rlabel polysilicon 275 -1720 275 -1720 0 3
rlabel polysilicon 282 -1714 282 -1714 0 1
rlabel polysilicon 282 -1720 282 -1720 0 3
rlabel polysilicon 289 -1714 289 -1714 0 1
rlabel polysilicon 289 -1720 289 -1720 0 3
rlabel polysilicon 296 -1714 296 -1714 0 1
rlabel polysilicon 296 -1720 296 -1720 0 3
rlabel polysilicon 303 -1714 303 -1714 0 1
rlabel polysilicon 303 -1720 303 -1720 0 3
rlabel polysilicon 310 -1714 310 -1714 0 1
rlabel polysilicon 313 -1714 313 -1714 0 2
rlabel polysilicon 310 -1720 310 -1720 0 3
rlabel polysilicon 317 -1714 317 -1714 0 1
rlabel polysilicon 317 -1720 317 -1720 0 3
rlabel polysilicon 327 -1714 327 -1714 0 2
rlabel polysilicon 324 -1720 324 -1720 0 3
rlabel polysilicon 331 -1714 331 -1714 0 1
rlabel polysilicon 331 -1720 331 -1720 0 3
rlabel polysilicon 341 -1714 341 -1714 0 2
rlabel polysilicon 341 -1720 341 -1720 0 4
rlabel polysilicon 345 -1714 345 -1714 0 1
rlabel polysilicon 345 -1720 345 -1720 0 3
rlabel polysilicon 355 -1714 355 -1714 0 2
rlabel polysilicon 352 -1720 352 -1720 0 3
rlabel polysilicon 355 -1720 355 -1720 0 4
rlabel polysilicon 359 -1714 359 -1714 0 1
rlabel polysilicon 362 -1714 362 -1714 0 2
rlabel polysilicon 362 -1720 362 -1720 0 4
rlabel polysilicon 366 -1714 366 -1714 0 1
rlabel polysilicon 366 -1720 366 -1720 0 3
rlabel polysilicon 373 -1714 373 -1714 0 1
rlabel polysilicon 376 -1714 376 -1714 0 2
rlabel polysilicon 373 -1720 373 -1720 0 3
rlabel polysilicon 376 -1720 376 -1720 0 4
rlabel polysilicon 380 -1714 380 -1714 0 1
rlabel polysilicon 383 -1714 383 -1714 0 2
rlabel polysilicon 380 -1720 380 -1720 0 3
rlabel polysilicon 383 -1720 383 -1720 0 4
rlabel polysilicon 387 -1714 387 -1714 0 1
rlabel polysilicon 387 -1720 387 -1720 0 3
rlabel polysilicon 394 -1714 394 -1714 0 1
rlabel polysilicon 394 -1720 394 -1720 0 3
rlabel polysilicon 401 -1714 401 -1714 0 1
rlabel polysilicon 401 -1720 401 -1720 0 3
rlabel polysilicon 408 -1714 408 -1714 0 1
rlabel polysilicon 408 -1720 408 -1720 0 3
rlabel polysilicon 415 -1714 415 -1714 0 1
rlabel polysilicon 415 -1720 415 -1720 0 3
rlabel polysilicon 422 -1714 422 -1714 0 1
rlabel polysilicon 425 -1720 425 -1720 0 4
rlabel polysilicon 429 -1714 429 -1714 0 1
rlabel polysilicon 429 -1720 429 -1720 0 3
rlabel polysilicon 436 -1714 436 -1714 0 1
rlabel polysilicon 436 -1720 436 -1720 0 3
rlabel polysilicon 443 -1714 443 -1714 0 1
rlabel polysilicon 443 -1720 443 -1720 0 3
rlabel polysilicon 450 -1714 450 -1714 0 1
rlabel polysilicon 450 -1720 450 -1720 0 3
rlabel polysilicon 457 -1714 457 -1714 0 1
rlabel polysilicon 457 -1720 457 -1720 0 3
rlabel polysilicon 464 -1714 464 -1714 0 1
rlabel polysilicon 464 -1720 464 -1720 0 3
rlabel polysilicon 471 -1714 471 -1714 0 1
rlabel polysilicon 471 -1720 471 -1720 0 3
rlabel polysilicon 478 -1714 478 -1714 0 1
rlabel polysilicon 481 -1714 481 -1714 0 2
rlabel polysilicon 485 -1714 485 -1714 0 1
rlabel polysilicon 488 -1714 488 -1714 0 2
rlabel polysilicon 485 -1720 485 -1720 0 3
rlabel polysilicon 488 -1720 488 -1720 0 4
rlabel polysilicon 492 -1720 492 -1720 0 3
rlabel polysilicon 495 -1720 495 -1720 0 4
rlabel polysilicon 499 -1714 499 -1714 0 1
rlabel polysilicon 499 -1720 499 -1720 0 3
rlabel polysilicon 506 -1714 506 -1714 0 1
rlabel polysilicon 506 -1720 506 -1720 0 3
rlabel polysilicon 513 -1714 513 -1714 0 1
rlabel polysilicon 513 -1720 513 -1720 0 3
rlabel polysilicon 523 -1714 523 -1714 0 2
rlabel polysilicon 520 -1720 520 -1720 0 3
rlabel polysilicon 523 -1720 523 -1720 0 4
rlabel polysilicon 527 -1714 527 -1714 0 1
rlabel polysilicon 527 -1720 527 -1720 0 3
rlabel polysilicon 530 -1720 530 -1720 0 4
rlabel polysilicon 534 -1714 534 -1714 0 1
rlabel polysilicon 534 -1720 534 -1720 0 3
rlabel polysilicon 541 -1714 541 -1714 0 1
rlabel polysilicon 541 -1720 541 -1720 0 3
rlabel polysilicon 548 -1714 548 -1714 0 1
rlabel polysilicon 548 -1720 548 -1720 0 3
rlabel polysilicon 555 -1714 555 -1714 0 1
rlabel polysilicon 555 -1720 555 -1720 0 3
rlabel polysilicon 562 -1714 562 -1714 0 1
rlabel polysilicon 562 -1720 562 -1720 0 3
rlabel polysilicon 569 -1714 569 -1714 0 1
rlabel polysilicon 569 -1720 569 -1720 0 3
rlabel polysilicon 579 -1714 579 -1714 0 2
rlabel polysilicon 576 -1720 576 -1720 0 3
rlabel polysilicon 579 -1720 579 -1720 0 4
rlabel polysilicon 586 -1714 586 -1714 0 2
rlabel polysilicon 586 -1720 586 -1720 0 4
rlabel polysilicon 590 -1714 590 -1714 0 1
rlabel polysilicon 590 -1720 590 -1720 0 3
rlabel polysilicon 597 -1714 597 -1714 0 1
rlabel polysilicon 597 -1720 597 -1720 0 3
rlabel polysilicon 607 -1714 607 -1714 0 2
rlabel polysilicon 604 -1720 604 -1720 0 3
rlabel polysilicon 607 -1720 607 -1720 0 4
rlabel polysilicon 611 -1714 611 -1714 0 1
rlabel polysilicon 611 -1720 611 -1720 0 3
rlabel polysilicon 618 -1714 618 -1714 0 1
rlabel polysilicon 618 -1720 618 -1720 0 3
rlabel polysilicon 625 -1714 625 -1714 0 1
rlabel polysilicon 625 -1720 625 -1720 0 3
rlabel polysilicon 632 -1714 632 -1714 0 1
rlabel polysilicon 632 -1720 632 -1720 0 3
rlabel polysilicon 639 -1714 639 -1714 0 1
rlabel polysilicon 639 -1720 639 -1720 0 3
rlabel polysilicon 646 -1714 646 -1714 0 1
rlabel polysilicon 646 -1720 646 -1720 0 3
rlabel polysilicon 653 -1714 653 -1714 0 1
rlabel polysilicon 656 -1714 656 -1714 0 2
rlabel polysilicon 653 -1720 653 -1720 0 3
rlabel polysilicon 660 -1714 660 -1714 0 1
rlabel polysilicon 663 -1714 663 -1714 0 2
rlabel polysilicon 660 -1720 660 -1720 0 3
rlabel polysilicon 667 -1714 667 -1714 0 1
rlabel polysilicon 667 -1720 667 -1720 0 3
rlabel polysilicon 674 -1714 674 -1714 0 1
rlabel polysilicon 674 -1720 674 -1720 0 3
rlabel polysilicon 677 -1720 677 -1720 0 4
rlabel polysilicon 681 -1714 681 -1714 0 1
rlabel polysilicon 681 -1720 681 -1720 0 3
rlabel polysilicon 691 -1714 691 -1714 0 2
rlabel polysilicon 688 -1720 688 -1720 0 3
rlabel polysilicon 695 -1714 695 -1714 0 1
rlabel polysilicon 695 -1720 695 -1720 0 3
rlabel polysilicon 702 -1714 702 -1714 0 1
rlabel polysilicon 702 -1720 702 -1720 0 3
rlabel polysilicon 709 -1714 709 -1714 0 1
rlabel polysilicon 709 -1720 709 -1720 0 3
rlabel polysilicon 716 -1714 716 -1714 0 1
rlabel polysilicon 716 -1720 716 -1720 0 3
rlabel polysilicon 723 -1714 723 -1714 0 1
rlabel polysilicon 723 -1720 723 -1720 0 3
rlabel polysilicon 730 -1714 730 -1714 0 1
rlabel polysilicon 730 -1720 730 -1720 0 3
rlabel polysilicon 737 -1714 737 -1714 0 1
rlabel polysilicon 737 -1720 737 -1720 0 3
rlabel polysilicon 744 -1714 744 -1714 0 1
rlabel polysilicon 744 -1720 744 -1720 0 3
rlabel polysilicon 751 -1714 751 -1714 0 1
rlabel polysilicon 751 -1720 751 -1720 0 3
rlabel polysilicon 758 -1714 758 -1714 0 1
rlabel polysilicon 761 -1714 761 -1714 0 2
rlabel polysilicon 761 -1720 761 -1720 0 4
rlabel polysilicon 765 -1714 765 -1714 0 1
rlabel polysilicon 765 -1720 765 -1720 0 3
rlabel polysilicon 772 -1714 772 -1714 0 1
rlabel polysilicon 772 -1720 772 -1720 0 3
rlabel polysilicon 779 -1714 779 -1714 0 1
rlabel polysilicon 779 -1720 779 -1720 0 3
rlabel polysilicon 786 -1714 786 -1714 0 1
rlabel polysilicon 786 -1720 786 -1720 0 3
rlabel polysilicon 793 -1714 793 -1714 0 1
rlabel polysilicon 793 -1720 793 -1720 0 3
rlabel polysilicon 800 -1714 800 -1714 0 1
rlabel polysilicon 800 -1720 800 -1720 0 3
rlabel polysilicon 807 -1714 807 -1714 0 1
rlabel polysilicon 807 -1720 807 -1720 0 3
rlabel polysilicon 817 -1720 817 -1720 0 4
rlabel polysilicon 821 -1714 821 -1714 0 1
rlabel polysilicon 821 -1720 821 -1720 0 3
rlabel polysilicon 828 -1714 828 -1714 0 1
rlabel polysilicon 828 -1720 828 -1720 0 3
rlabel polysilicon 835 -1714 835 -1714 0 1
rlabel polysilicon 835 -1720 835 -1720 0 3
rlabel polysilicon 842 -1714 842 -1714 0 1
rlabel polysilicon 842 -1720 842 -1720 0 3
rlabel polysilicon 849 -1714 849 -1714 0 1
rlabel polysilicon 849 -1720 849 -1720 0 3
rlabel polysilicon 856 -1714 856 -1714 0 1
rlabel polysilicon 856 -1720 856 -1720 0 3
rlabel polysilicon 863 -1714 863 -1714 0 1
rlabel polysilicon 863 -1720 863 -1720 0 3
rlabel polysilicon 870 -1714 870 -1714 0 1
rlabel polysilicon 870 -1720 870 -1720 0 3
rlabel polysilicon 877 -1714 877 -1714 0 1
rlabel polysilicon 877 -1720 877 -1720 0 3
rlabel polysilicon 884 -1714 884 -1714 0 1
rlabel polysilicon 884 -1720 884 -1720 0 3
rlabel polysilicon 891 -1714 891 -1714 0 1
rlabel polysilicon 891 -1720 891 -1720 0 3
rlabel polysilicon 898 -1714 898 -1714 0 1
rlabel polysilicon 898 -1720 898 -1720 0 3
rlabel polysilicon 905 -1714 905 -1714 0 1
rlabel polysilicon 905 -1720 905 -1720 0 3
rlabel polysilicon 908 -1720 908 -1720 0 4
rlabel polysilicon 912 -1714 912 -1714 0 1
rlabel polysilicon 912 -1720 912 -1720 0 3
rlabel polysilicon 919 -1714 919 -1714 0 1
rlabel polysilicon 919 -1720 919 -1720 0 3
rlabel polysilicon 926 -1720 926 -1720 0 3
rlabel polysilicon 929 -1720 929 -1720 0 4
rlabel polysilicon 933 -1714 933 -1714 0 1
rlabel polysilicon 933 -1720 933 -1720 0 3
rlabel polysilicon 940 -1714 940 -1714 0 1
rlabel polysilicon 940 -1720 940 -1720 0 3
rlabel polysilicon 947 -1714 947 -1714 0 1
rlabel polysilicon 947 -1720 947 -1720 0 3
rlabel polysilicon 954 -1714 954 -1714 0 1
rlabel polysilicon 954 -1720 954 -1720 0 3
rlabel polysilicon 961 -1714 961 -1714 0 1
rlabel polysilicon 961 -1720 961 -1720 0 3
rlabel polysilicon 968 -1714 968 -1714 0 1
rlabel polysilicon 968 -1720 968 -1720 0 3
rlabel polysilicon 1066 -1714 1066 -1714 0 1
rlabel polysilicon 1069 -1720 1069 -1720 0 4
rlabel polysilicon 1094 -1714 1094 -1714 0 1
rlabel polysilicon 1094 -1720 1094 -1720 0 3
rlabel polysilicon 2 -1805 2 -1805 0 1
rlabel polysilicon 2 -1811 2 -1811 0 3
rlabel polysilicon 9 -1811 9 -1811 0 3
rlabel polysilicon 16 -1805 16 -1805 0 1
rlabel polysilicon 16 -1811 16 -1811 0 3
rlabel polysilicon 23 -1805 23 -1805 0 1
rlabel polysilicon 23 -1811 23 -1811 0 3
rlabel polysilicon 30 -1805 30 -1805 0 1
rlabel polysilicon 30 -1811 30 -1811 0 3
rlabel polysilicon 37 -1805 37 -1805 0 1
rlabel polysilicon 37 -1811 37 -1811 0 3
rlabel polysilicon 44 -1805 44 -1805 0 1
rlabel polysilicon 44 -1811 44 -1811 0 3
rlabel polysilicon 51 -1805 51 -1805 0 1
rlabel polysilicon 51 -1811 51 -1811 0 3
rlabel polysilicon 58 -1805 58 -1805 0 1
rlabel polysilicon 58 -1811 58 -1811 0 3
rlabel polysilicon 65 -1805 65 -1805 0 1
rlabel polysilicon 65 -1811 65 -1811 0 3
rlabel polysilicon 72 -1805 72 -1805 0 1
rlabel polysilicon 72 -1811 72 -1811 0 3
rlabel polysilicon 79 -1805 79 -1805 0 1
rlabel polysilicon 79 -1811 79 -1811 0 3
rlabel polysilicon 86 -1805 86 -1805 0 1
rlabel polysilicon 86 -1811 86 -1811 0 3
rlabel polysilicon 93 -1811 93 -1811 0 3
rlabel polysilicon 96 -1811 96 -1811 0 4
rlabel polysilicon 100 -1805 100 -1805 0 1
rlabel polysilicon 100 -1811 100 -1811 0 3
rlabel polysilicon 103 -1811 103 -1811 0 4
rlabel polysilicon 107 -1805 107 -1805 0 1
rlabel polysilicon 107 -1811 107 -1811 0 3
rlabel polysilicon 117 -1805 117 -1805 0 2
rlabel polysilicon 114 -1811 114 -1811 0 3
rlabel polysilicon 117 -1811 117 -1811 0 4
rlabel polysilicon 121 -1805 121 -1805 0 1
rlabel polysilicon 121 -1811 121 -1811 0 3
rlabel polysilicon 128 -1805 128 -1805 0 1
rlabel polysilicon 128 -1811 128 -1811 0 3
rlabel polysilicon 135 -1805 135 -1805 0 1
rlabel polysilicon 138 -1805 138 -1805 0 2
rlabel polysilicon 135 -1811 135 -1811 0 3
rlabel polysilicon 142 -1805 142 -1805 0 1
rlabel polysilicon 142 -1811 142 -1811 0 3
rlabel polysilicon 149 -1805 149 -1805 0 1
rlabel polysilicon 149 -1811 149 -1811 0 3
rlabel polysilicon 156 -1805 156 -1805 0 1
rlabel polysilicon 156 -1811 156 -1811 0 3
rlabel polysilicon 163 -1805 163 -1805 0 1
rlabel polysilicon 163 -1811 163 -1811 0 3
rlabel polysilicon 170 -1805 170 -1805 0 1
rlabel polysilicon 170 -1811 170 -1811 0 3
rlabel polysilicon 177 -1805 177 -1805 0 1
rlabel polysilicon 177 -1811 177 -1811 0 3
rlabel polysilicon 184 -1805 184 -1805 0 1
rlabel polysilicon 191 -1805 191 -1805 0 1
rlabel polysilicon 191 -1811 191 -1811 0 3
rlabel polysilicon 198 -1805 198 -1805 0 1
rlabel polysilicon 198 -1811 198 -1811 0 3
rlabel polysilicon 201 -1811 201 -1811 0 4
rlabel polysilicon 205 -1811 205 -1811 0 3
rlabel polysilicon 208 -1811 208 -1811 0 4
rlabel polysilicon 212 -1805 212 -1805 0 1
rlabel polysilicon 212 -1811 212 -1811 0 3
rlabel polysilicon 219 -1805 219 -1805 0 1
rlabel polysilicon 222 -1805 222 -1805 0 2
rlabel polysilicon 219 -1811 219 -1811 0 3
rlabel polysilicon 226 -1805 226 -1805 0 1
rlabel polysilicon 226 -1811 226 -1811 0 3
rlabel polysilicon 233 -1805 233 -1805 0 1
rlabel polysilicon 233 -1811 233 -1811 0 3
rlabel polysilicon 240 -1805 240 -1805 0 1
rlabel polysilicon 240 -1811 240 -1811 0 3
rlabel polysilicon 247 -1805 247 -1805 0 1
rlabel polysilicon 247 -1811 247 -1811 0 3
rlabel polysilicon 250 -1811 250 -1811 0 4
rlabel polysilicon 254 -1805 254 -1805 0 1
rlabel polysilicon 254 -1811 254 -1811 0 3
rlabel polysilicon 261 -1805 261 -1805 0 1
rlabel polysilicon 261 -1811 261 -1811 0 3
rlabel polysilicon 268 -1805 268 -1805 0 1
rlabel polysilicon 268 -1811 268 -1811 0 3
rlabel polysilicon 275 -1805 275 -1805 0 1
rlabel polysilicon 275 -1811 275 -1811 0 3
rlabel polysilicon 282 -1805 282 -1805 0 1
rlabel polysilicon 282 -1811 282 -1811 0 3
rlabel polysilicon 289 -1805 289 -1805 0 1
rlabel polysilicon 289 -1811 289 -1811 0 3
rlabel polysilicon 296 -1805 296 -1805 0 1
rlabel polysilicon 296 -1811 296 -1811 0 3
rlabel polysilicon 303 -1805 303 -1805 0 1
rlabel polysilicon 306 -1805 306 -1805 0 2
rlabel polysilicon 306 -1811 306 -1811 0 4
rlabel polysilicon 310 -1805 310 -1805 0 1
rlabel polysilicon 310 -1811 310 -1811 0 3
rlabel polysilicon 317 -1805 317 -1805 0 1
rlabel polysilicon 317 -1811 317 -1811 0 3
rlabel polysilicon 324 -1805 324 -1805 0 1
rlabel polysilicon 324 -1811 324 -1811 0 3
rlabel polysilicon 331 -1805 331 -1805 0 1
rlabel polysilicon 331 -1811 331 -1811 0 3
rlabel polysilicon 338 -1805 338 -1805 0 1
rlabel polysilicon 338 -1811 338 -1811 0 3
rlabel polysilicon 348 -1805 348 -1805 0 2
rlabel polysilicon 348 -1811 348 -1811 0 4
rlabel polysilicon 352 -1805 352 -1805 0 1
rlabel polysilicon 352 -1811 352 -1811 0 3
rlabel polysilicon 355 -1811 355 -1811 0 4
rlabel polysilicon 359 -1805 359 -1805 0 1
rlabel polysilicon 359 -1811 359 -1811 0 3
rlabel polysilicon 366 -1805 366 -1805 0 1
rlabel polysilicon 366 -1811 366 -1811 0 3
rlabel polysilicon 373 -1805 373 -1805 0 1
rlabel polysilicon 373 -1811 373 -1811 0 3
rlabel polysilicon 380 -1805 380 -1805 0 1
rlabel polysilicon 380 -1811 380 -1811 0 3
rlabel polysilicon 387 -1805 387 -1805 0 1
rlabel polysilicon 387 -1811 387 -1811 0 3
rlabel polysilicon 394 -1805 394 -1805 0 1
rlabel polysilicon 394 -1811 394 -1811 0 3
rlabel polysilicon 401 -1805 401 -1805 0 1
rlabel polysilicon 401 -1811 401 -1811 0 3
rlabel polysilicon 408 -1805 408 -1805 0 1
rlabel polysilicon 408 -1811 408 -1811 0 3
rlabel polysilicon 415 -1805 415 -1805 0 1
rlabel polysilicon 418 -1805 418 -1805 0 2
rlabel polysilicon 415 -1811 415 -1811 0 3
rlabel polysilicon 418 -1811 418 -1811 0 4
rlabel polysilicon 425 -1805 425 -1805 0 2
rlabel polysilicon 422 -1811 422 -1811 0 3
rlabel polysilicon 425 -1811 425 -1811 0 4
rlabel polysilicon 429 -1805 429 -1805 0 1
rlabel polysilicon 432 -1805 432 -1805 0 2
rlabel polysilicon 429 -1811 429 -1811 0 3
rlabel polysilicon 432 -1811 432 -1811 0 4
rlabel polysilicon 436 -1805 436 -1805 0 1
rlabel polysilicon 436 -1811 436 -1811 0 3
rlabel polysilicon 443 -1805 443 -1805 0 1
rlabel polysilicon 443 -1811 443 -1811 0 3
rlabel polysilicon 450 -1805 450 -1805 0 1
rlabel polysilicon 450 -1811 450 -1811 0 3
rlabel polysilicon 457 -1805 457 -1805 0 1
rlabel polysilicon 457 -1811 457 -1811 0 3
rlabel polysilicon 464 -1805 464 -1805 0 1
rlabel polysilicon 464 -1811 464 -1811 0 3
rlabel polysilicon 471 -1805 471 -1805 0 1
rlabel polysilicon 471 -1811 471 -1811 0 3
rlabel polysilicon 478 -1805 478 -1805 0 1
rlabel polysilicon 478 -1811 478 -1811 0 3
rlabel polysilicon 485 -1805 485 -1805 0 1
rlabel polysilicon 485 -1811 485 -1811 0 3
rlabel polysilicon 492 -1805 492 -1805 0 1
rlabel polysilicon 492 -1811 492 -1811 0 3
rlabel polysilicon 499 -1805 499 -1805 0 1
rlabel polysilicon 502 -1805 502 -1805 0 2
rlabel polysilicon 499 -1811 499 -1811 0 3
rlabel polysilicon 506 -1805 506 -1805 0 1
rlabel polysilicon 506 -1811 506 -1811 0 3
rlabel polysilicon 513 -1805 513 -1805 0 1
rlabel polysilicon 513 -1811 513 -1811 0 3
rlabel polysilicon 520 -1805 520 -1805 0 1
rlabel polysilicon 520 -1811 520 -1811 0 3
rlabel polysilicon 523 -1811 523 -1811 0 4
rlabel polysilicon 527 -1805 527 -1805 0 1
rlabel polysilicon 530 -1805 530 -1805 0 2
rlabel polysilicon 527 -1811 527 -1811 0 3
rlabel polysilicon 534 -1805 534 -1805 0 1
rlabel polysilicon 534 -1811 534 -1811 0 3
rlabel polysilicon 541 -1805 541 -1805 0 1
rlabel polysilicon 541 -1811 541 -1811 0 3
rlabel polysilicon 548 -1805 548 -1805 0 1
rlabel polysilicon 551 -1811 551 -1811 0 4
rlabel polysilicon 555 -1805 555 -1805 0 1
rlabel polysilicon 555 -1811 555 -1811 0 3
rlabel polysilicon 562 -1805 562 -1805 0 1
rlabel polysilicon 562 -1811 562 -1811 0 3
rlabel polysilicon 569 -1805 569 -1805 0 1
rlabel polysilicon 569 -1811 569 -1811 0 3
rlabel polysilicon 576 -1805 576 -1805 0 1
rlabel polysilicon 576 -1811 576 -1811 0 3
rlabel polysilicon 583 -1805 583 -1805 0 1
rlabel polysilicon 583 -1811 583 -1811 0 3
rlabel polysilicon 590 -1805 590 -1805 0 1
rlabel polysilicon 590 -1811 590 -1811 0 3
rlabel polysilicon 597 -1805 597 -1805 0 1
rlabel polysilicon 600 -1805 600 -1805 0 2
rlabel polysilicon 604 -1805 604 -1805 0 1
rlabel polysilicon 604 -1811 604 -1811 0 3
rlabel polysilicon 611 -1805 611 -1805 0 1
rlabel polysilicon 611 -1811 611 -1811 0 3
rlabel polysilicon 614 -1811 614 -1811 0 4
rlabel polysilicon 618 -1805 618 -1805 0 1
rlabel polysilicon 618 -1811 618 -1811 0 3
rlabel polysilicon 625 -1805 625 -1805 0 1
rlabel polysilicon 625 -1811 625 -1811 0 3
rlabel polysilicon 628 -1811 628 -1811 0 4
rlabel polysilicon 632 -1805 632 -1805 0 1
rlabel polysilicon 632 -1811 632 -1811 0 3
rlabel polysilicon 639 -1805 639 -1805 0 1
rlabel polysilicon 639 -1811 639 -1811 0 3
rlabel polysilicon 646 -1805 646 -1805 0 1
rlabel polysilicon 646 -1811 646 -1811 0 3
rlabel polysilicon 653 -1805 653 -1805 0 1
rlabel polysilicon 653 -1811 653 -1811 0 3
rlabel polysilicon 660 -1805 660 -1805 0 1
rlabel polysilicon 660 -1811 660 -1811 0 3
rlabel polysilicon 667 -1805 667 -1805 0 1
rlabel polysilicon 670 -1805 670 -1805 0 2
rlabel polysilicon 670 -1811 670 -1811 0 4
rlabel polysilicon 674 -1805 674 -1805 0 1
rlabel polysilicon 674 -1811 674 -1811 0 3
rlabel polysilicon 681 -1805 681 -1805 0 1
rlabel polysilicon 681 -1811 681 -1811 0 3
rlabel polysilicon 688 -1805 688 -1805 0 1
rlabel polysilicon 691 -1805 691 -1805 0 2
rlabel polysilicon 691 -1811 691 -1811 0 4
rlabel polysilicon 695 -1805 695 -1805 0 1
rlabel polysilicon 695 -1811 695 -1811 0 3
rlabel polysilicon 702 -1805 702 -1805 0 1
rlabel polysilicon 702 -1811 702 -1811 0 3
rlabel polysilicon 712 -1805 712 -1805 0 2
rlabel polysilicon 709 -1811 709 -1811 0 3
rlabel polysilicon 712 -1811 712 -1811 0 4
rlabel polysilicon 716 -1805 716 -1805 0 1
rlabel polysilicon 716 -1811 716 -1811 0 3
rlabel polysilicon 723 -1805 723 -1805 0 1
rlabel polysilicon 723 -1811 723 -1811 0 3
rlabel polysilicon 730 -1805 730 -1805 0 1
rlabel polysilicon 730 -1811 730 -1811 0 3
rlabel polysilicon 737 -1805 737 -1805 0 1
rlabel polysilicon 737 -1811 737 -1811 0 3
rlabel polysilicon 744 -1805 744 -1805 0 1
rlabel polysilicon 744 -1811 744 -1811 0 3
rlabel polysilicon 751 -1805 751 -1805 0 1
rlabel polysilicon 751 -1811 751 -1811 0 3
rlabel polysilicon 758 -1805 758 -1805 0 1
rlabel polysilicon 758 -1811 758 -1811 0 3
rlabel polysilicon 765 -1805 765 -1805 0 1
rlabel polysilicon 765 -1811 765 -1811 0 3
rlabel polysilicon 772 -1805 772 -1805 0 1
rlabel polysilicon 772 -1811 772 -1811 0 3
rlabel polysilicon 779 -1805 779 -1805 0 1
rlabel polysilicon 779 -1811 779 -1811 0 3
rlabel polysilicon 786 -1805 786 -1805 0 1
rlabel polysilicon 786 -1811 786 -1811 0 3
rlabel polysilicon 793 -1805 793 -1805 0 1
rlabel polysilicon 793 -1811 793 -1811 0 3
rlabel polysilicon 800 -1805 800 -1805 0 1
rlabel polysilicon 800 -1811 800 -1811 0 3
rlabel polysilicon 807 -1805 807 -1805 0 1
rlabel polysilicon 807 -1811 807 -1811 0 3
rlabel polysilicon 814 -1805 814 -1805 0 1
rlabel polysilicon 814 -1811 814 -1811 0 3
rlabel polysilicon 821 -1805 821 -1805 0 1
rlabel polysilicon 821 -1811 821 -1811 0 3
rlabel polysilicon 828 -1805 828 -1805 0 1
rlabel polysilicon 828 -1811 828 -1811 0 3
rlabel polysilicon 835 -1805 835 -1805 0 1
rlabel polysilicon 835 -1811 835 -1811 0 3
rlabel polysilicon 842 -1805 842 -1805 0 1
rlabel polysilicon 842 -1811 842 -1811 0 3
rlabel polysilicon 849 -1805 849 -1805 0 1
rlabel polysilicon 849 -1811 849 -1811 0 3
rlabel polysilicon 856 -1805 856 -1805 0 1
rlabel polysilicon 856 -1811 856 -1811 0 3
rlabel polysilicon 863 -1805 863 -1805 0 1
rlabel polysilicon 863 -1811 863 -1811 0 3
rlabel polysilicon 870 -1805 870 -1805 0 1
rlabel polysilicon 870 -1811 870 -1811 0 3
rlabel polysilicon 877 -1805 877 -1805 0 1
rlabel polysilicon 877 -1811 877 -1811 0 3
rlabel polysilicon 884 -1805 884 -1805 0 1
rlabel polysilicon 884 -1811 884 -1811 0 3
rlabel polysilicon 891 -1805 891 -1805 0 1
rlabel polysilicon 891 -1811 891 -1811 0 3
rlabel polysilicon 898 -1805 898 -1805 0 1
rlabel polysilicon 898 -1811 898 -1811 0 3
rlabel polysilicon 905 -1805 905 -1805 0 1
rlabel polysilicon 905 -1811 905 -1811 0 3
rlabel polysilicon 912 -1805 912 -1805 0 1
rlabel polysilicon 912 -1811 912 -1811 0 3
rlabel polysilicon 919 -1805 919 -1805 0 1
rlabel polysilicon 919 -1811 919 -1811 0 3
rlabel polysilicon 926 -1805 926 -1805 0 1
rlabel polysilicon 926 -1811 926 -1811 0 3
rlabel polysilicon 933 -1811 933 -1811 0 3
rlabel polysilicon 940 -1805 940 -1805 0 1
rlabel polysilicon 940 -1811 940 -1811 0 3
rlabel polysilicon 947 -1805 947 -1805 0 1
rlabel polysilicon 947 -1811 947 -1811 0 3
rlabel polysilicon 954 -1805 954 -1805 0 1
rlabel polysilicon 954 -1811 954 -1811 0 3
rlabel polysilicon 961 -1805 961 -1805 0 1
rlabel polysilicon 961 -1811 961 -1811 0 3
rlabel polysilicon 968 -1805 968 -1805 0 1
rlabel polysilicon 968 -1811 968 -1811 0 3
rlabel polysilicon 975 -1805 975 -1805 0 1
rlabel polysilicon 975 -1811 975 -1811 0 3
rlabel polysilicon 982 -1805 982 -1805 0 1
rlabel polysilicon 982 -1811 982 -1811 0 3
rlabel polysilicon 989 -1805 989 -1805 0 1
rlabel polysilicon 989 -1811 989 -1811 0 3
rlabel polysilicon 996 -1805 996 -1805 0 1
rlabel polysilicon 996 -1811 996 -1811 0 3
rlabel polysilicon 1003 -1805 1003 -1805 0 1
rlabel polysilicon 1003 -1811 1003 -1811 0 3
rlabel polysilicon 1010 -1805 1010 -1805 0 1
rlabel polysilicon 1010 -1811 1010 -1811 0 3
rlabel polysilicon 1017 -1805 1017 -1805 0 1
rlabel polysilicon 1017 -1811 1017 -1811 0 3
rlabel polysilicon 1024 -1805 1024 -1805 0 1
rlabel polysilicon 1024 -1811 1024 -1811 0 3
rlabel polysilicon 1031 -1805 1031 -1805 0 1
rlabel polysilicon 1031 -1811 1031 -1811 0 3
rlabel polysilicon 1038 -1805 1038 -1805 0 1
rlabel polysilicon 1038 -1811 1038 -1811 0 3
rlabel polysilicon 1045 -1805 1045 -1805 0 1
rlabel polysilicon 1045 -1811 1045 -1811 0 3
rlabel polysilicon 1052 -1805 1052 -1805 0 1
rlabel polysilicon 1055 -1805 1055 -1805 0 2
rlabel polysilicon 1055 -1811 1055 -1811 0 4
rlabel polysilicon 1059 -1805 1059 -1805 0 1
rlabel polysilicon 1059 -1811 1059 -1811 0 3
rlabel polysilicon 1087 -1805 1087 -1805 0 1
rlabel polysilicon 1087 -1811 1087 -1811 0 3
rlabel polysilicon 1094 -1805 1094 -1805 0 1
rlabel polysilicon 1094 -1811 1094 -1811 0 3
rlabel polysilicon 5 -1896 5 -1896 0 2
rlabel polysilicon 9 -1896 9 -1896 0 1
rlabel polysilicon 9 -1902 9 -1902 0 3
rlabel polysilicon 16 -1896 16 -1896 0 1
rlabel polysilicon 19 -1902 19 -1902 0 4
rlabel polysilicon 23 -1896 23 -1896 0 1
rlabel polysilicon 23 -1902 23 -1902 0 3
rlabel polysilicon 30 -1896 30 -1896 0 1
rlabel polysilicon 30 -1902 30 -1902 0 3
rlabel polysilicon 40 -1896 40 -1896 0 2
rlabel polysilicon 40 -1902 40 -1902 0 4
rlabel polysilicon 44 -1896 44 -1896 0 1
rlabel polysilicon 47 -1896 47 -1896 0 2
rlabel polysilicon 44 -1902 44 -1902 0 3
rlabel polysilicon 47 -1902 47 -1902 0 4
rlabel polysilicon 51 -1896 51 -1896 0 1
rlabel polysilicon 54 -1896 54 -1896 0 2
rlabel polysilicon 51 -1902 51 -1902 0 3
rlabel polysilicon 54 -1902 54 -1902 0 4
rlabel polysilicon 58 -1896 58 -1896 0 1
rlabel polysilicon 58 -1902 58 -1902 0 3
rlabel polysilicon 65 -1896 65 -1896 0 1
rlabel polysilicon 68 -1896 68 -1896 0 2
rlabel polysilicon 72 -1896 72 -1896 0 1
rlabel polysilicon 72 -1902 72 -1902 0 3
rlabel polysilicon 79 -1896 79 -1896 0 1
rlabel polysilicon 82 -1896 82 -1896 0 2
rlabel polysilicon 82 -1902 82 -1902 0 4
rlabel polysilicon 86 -1896 86 -1896 0 1
rlabel polysilicon 86 -1902 86 -1902 0 3
rlabel polysilicon 93 -1896 93 -1896 0 1
rlabel polysilicon 93 -1902 93 -1902 0 3
rlabel polysilicon 100 -1896 100 -1896 0 1
rlabel polysilicon 100 -1902 100 -1902 0 3
rlabel polysilicon 107 -1896 107 -1896 0 1
rlabel polysilicon 107 -1902 107 -1902 0 3
rlabel polysilicon 114 -1896 114 -1896 0 1
rlabel polysilicon 117 -1896 117 -1896 0 2
rlabel polysilicon 117 -1902 117 -1902 0 4
rlabel polysilicon 121 -1896 121 -1896 0 1
rlabel polysilicon 124 -1896 124 -1896 0 2
rlabel polysilicon 121 -1902 121 -1902 0 3
rlabel polysilicon 124 -1902 124 -1902 0 4
rlabel polysilicon 128 -1896 128 -1896 0 1
rlabel polysilicon 128 -1902 128 -1902 0 3
rlabel polysilicon 135 -1896 135 -1896 0 1
rlabel polysilicon 135 -1902 135 -1902 0 3
rlabel polysilicon 142 -1896 142 -1896 0 1
rlabel polysilicon 142 -1902 142 -1902 0 3
rlabel polysilicon 149 -1902 149 -1902 0 3
rlabel polysilicon 152 -1902 152 -1902 0 4
rlabel polysilicon 156 -1896 156 -1896 0 1
rlabel polysilicon 156 -1902 156 -1902 0 3
rlabel polysilicon 159 -1902 159 -1902 0 4
rlabel polysilicon 163 -1896 163 -1896 0 1
rlabel polysilicon 163 -1902 163 -1902 0 3
rlabel polysilicon 170 -1896 170 -1896 0 1
rlabel polysilicon 170 -1902 170 -1902 0 3
rlabel polysilicon 177 -1896 177 -1896 0 1
rlabel polysilicon 177 -1902 177 -1902 0 3
rlabel polysilicon 184 -1896 184 -1896 0 1
rlabel polysilicon 184 -1902 184 -1902 0 3
rlabel polysilicon 194 -1896 194 -1896 0 2
rlabel polysilicon 194 -1902 194 -1902 0 4
rlabel polysilicon 198 -1896 198 -1896 0 1
rlabel polysilicon 198 -1902 198 -1902 0 3
rlabel polysilicon 205 -1896 205 -1896 0 1
rlabel polysilicon 205 -1902 205 -1902 0 3
rlabel polysilicon 212 -1896 212 -1896 0 1
rlabel polysilicon 212 -1902 212 -1902 0 3
rlabel polysilicon 222 -1902 222 -1902 0 4
rlabel polysilicon 226 -1896 226 -1896 0 1
rlabel polysilicon 226 -1902 226 -1902 0 3
rlabel polysilicon 233 -1896 233 -1896 0 1
rlabel polysilicon 233 -1902 233 -1902 0 3
rlabel polysilicon 240 -1896 240 -1896 0 1
rlabel polysilicon 240 -1902 240 -1902 0 3
rlabel polysilicon 247 -1896 247 -1896 0 1
rlabel polysilicon 247 -1902 247 -1902 0 3
rlabel polysilicon 254 -1896 254 -1896 0 1
rlabel polysilicon 254 -1902 254 -1902 0 3
rlabel polysilicon 261 -1896 261 -1896 0 1
rlabel polysilicon 261 -1902 261 -1902 0 3
rlabel polysilicon 268 -1896 268 -1896 0 1
rlabel polysilicon 268 -1902 268 -1902 0 3
rlabel polysilicon 275 -1896 275 -1896 0 1
rlabel polysilicon 275 -1902 275 -1902 0 3
rlabel polysilicon 282 -1896 282 -1896 0 1
rlabel polysilicon 282 -1902 282 -1902 0 3
rlabel polysilicon 289 -1896 289 -1896 0 1
rlabel polysilicon 289 -1902 289 -1902 0 3
rlabel polysilicon 296 -1896 296 -1896 0 1
rlabel polysilicon 296 -1902 296 -1902 0 3
rlabel polysilicon 303 -1896 303 -1896 0 1
rlabel polysilicon 303 -1902 303 -1902 0 3
rlabel polysilicon 310 -1896 310 -1896 0 1
rlabel polysilicon 310 -1902 310 -1902 0 3
rlabel polysilicon 317 -1896 317 -1896 0 1
rlabel polysilicon 317 -1902 317 -1902 0 3
rlabel polysilicon 324 -1896 324 -1896 0 1
rlabel polysilicon 324 -1902 324 -1902 0 3
rlabel polysilicon 331 -1896 331 -1896 0 1
rlabel polysilicon 331 -1902 331 -1902 0 3
rlabel polysilicon 338 -1896 338 -1896 0 1
rlabel polysilicon 338 -1902 338 -1902 0 3
rlabel polysilicon 345 -1896 345 -1896 0 1
rlabel polysilicon 345 -1902 345 -1902 0 3
rlabel polysilicon 352 -1896 352 -1896 0 1
rlabel polysilicon 352 -1902 352 -1902 0 3
rlabel polysilicon 359 -1896 359 -1896 0 1
rlabel polysilicon 362 -1896 362 -1896 0 2
rlabel polysilicon 359 -1902 359 -1902 0 3
rlabel polysilicon 366 -1896 366 -1896 0 1
rlabel polysilicon 369 -1896 369 -1896 0 2
rlabel polysilicon 366 -1902 366 -1902 0 3
rlabel polysilicon 369 -1902 369 -1902 0 4
rlabel polysilicon 373 -1896 373 -1896 0 1
rlabel polysilicon 373 -1902 373 -1902 0 3
rlabel polysilicon 380 -1896 380 -1896 0 1
rlabel polysilicon 380 -1902 380 -1902 0 3
rlabel polysilicon 387 -1896 387 -1896 0 1
rlabel polysilicon 390 -1896 390 -1896 0 2
rlabel polysilicon 390 -1902 390 -1902 0 4
rlabel polysilicon 394 -1896 394 -1896 0 1
rlabel polysilicon 394 -1902 394 -1902 0 3
rlabel polysilicon 401 -1896 401 -1896 0 1
rlabel polysilicon 401 -1902 401 -1902 0 3
rlabel polysilicon 408 -1896 408 -1896 0 1
rlabel polysilicon 408 -1902 408 -1902 0 3
rlabel polysilicon 418 -1896 418 -1896 0 2
rlabel polysilicon 415 -1902 415 -1902 0 3
rlabel polysilicon 422 -1896 422 -1896 0 1
rlabel polysilicon 422 -1902 422 -1902 0 3
rlabel polysilicon 429 -1896 429 -1896 0 1
rlabel polysilicon 429 -1902 429 -1902 0 3
rlabel polysilicon 436 -1896 436 -1896 0 1
rlabel polysilicon 436 -1902 436 -1902 0 3
rlabel polysilicon 443 -1896 443 -1896 0 1
rlabel polysilicon 446 -1896 446 -1896 0 2
rlabel polysilicon 450 -1896 450 -1896 0 1
rlabel polysilicon 453 -1902 453 -1902 0 4
rlabel polysilicon 457 -1896 457 -1896 0 1
rlabel polysilicon 457 -1902 457 -1902 0 3
rlabel polysilicon 464 -1896 464 -1896 0 1
rlabel polysilicon 464 -1902 464 -1902 0 3
rlabel polysilicon 471 -1896 471 -1896 0 1
rlabel polysilicon 471 -1902 471 -1902 0 3
rlabel polysilicon 478 -1896 478 -1896 0 1
rlabel polysilicon 481 -1896 481 -1896 0 2
rlabel polysilicon 478 -1902 478 -1902 0 3
rlabel polysilicon 481 -1902 481 -1902 0 4
rlabel polysilicon 485 -1896 485 -1896 0 1
rlabel polysilicon 488 -1896 488 -1896 0 2
rlabel polysilicon 485 -1902 485 -1902 0 3
rlabel polysilicon 492 -1896 492 -1896 0 1
rlabel polysilicon 492 -1902 492 -1902 0 3
rlabel polysilicon 502 -1896 502 -1896 0 2
rlabel polysilicon 499 -1902 499 -1902 0 3
rlabel polysilicon 502 -1902 502 -1902 0 4
rlabel polysilicon 506 -1896 506 -1896 0 1
rlabel polysilicon 506 -1902 506 -1902 0 3
rlabel polysilicon 513 -1896 513 -1896 0 1
rlabel polysilicon 513 -1902 513 -1902 0 3
rlabel polysilicon 520 -1896 520 -1896 0 1
rlabel polysilicon 520 -1902 520 -1902 0 3
rlabel polysilicon 527 -1902 527 -1902 0 3
rlabel polysilicon 530 -1902 530 -1902 0 4
rlabel polysilicon 534 -1896 534 -1896 0 1
rlabel polysilicon 534 -1902 534 -1902 0 3
rlabel polysilicon 541 -1896 541 -1896 0 1
rlabel polysilicon 541 -1902 541 -1902 0 3
rlabel polysilicon 548 -1896 548 -1896 0 1
rlabel polysilicon 551 -1896 551 -1896 0 2
rlabel polysilicon 548 -1902 548 -1902 0 3
rlabel polysilicon 551 -1902 551 -1902 0 4
rlabel polysilicon 555 -1896 555 -1896 0 1
rlabel polysilicon 558 -1896 558 -1896 0 2
rlabel polysilicon 558 -1902 558 -1902 0 4
rlabel polysilicon 562 -1896 562 -1896 0 1
rlabel polysilicon 562 -1902 562 -1902 0 3
rlabel polysilicon 569 -1896 569 -1896 0 1
rlabel polysilicon 569 -1902 569 -1902 0 3
rlabel polysilicon 576 -1896 576 -1896 0 1
rlabel polysilicon 576 -1902 576 -1902 0 3
rlabel polysilicon 583 -1896 583 -1896 0 1
rlabel polysilicon 583 -1902 583 -1902 0 3
rlabel polysilicon 590 -1896 590 -1896 0 1
rlabel polysilicon 590 -1902 590 -1902 0 3
rlabel polysilicon 597 -1896 597 -1896 0 1
rlabel polysilicon 597 -1902 597 -1902 0 3
rlabel polysilicon 604 -1896 604 -1896 0 1
rlabel polysilicon 604 -1902 604 -1902 0 3
rlabel polysilicon 611 -1896 611 -1896 0 1
rlabel polysilicon 611 -1902 611 -1902 0 3
rlabel polysilicon 621 -1896 621 -1896 0 2
rlabel polysilicon 618 -1902 618 -1902 0 3
rlabel polysilicon 621 -1902 621 -1902 0 4
rlabel polysilicon 625 -1896 625 -1896 0 1
rlabel polysilicon 625 -1902 625 -1902 0 3
rlabel polysilicon 632 -1896 632 -1896 0 1
rlabel polysilicon 635 -1896 635 -1896 0 2
rlabel polysilicon 632 -1902 632 -1902 0 3
rlabel polysilicon 635 -1902 635 -1902 0 4
rlabel polysilicon 639 -1896 639 -1896 0 1
rlabel polysilicon 639 -1902 639 -1902 0 3
rlabel polysilicon 646 -1896 646 -1896 0 1
rlabel polysilicon 646 -1902 646 -1902 0 3
rlabel polysilicon 653 -1896 653 -1896 0 1
rlabel polysilicon 653 -1902 653 -1902 0 3
rlabel polysilicon 660 -1896 660 -1896 0 1
rlabel polysilicon 660 -1902 660 -1902 0 3
rlabel polysilicon 667 -1896 667 -1896 0 1
rlabel polysilicon 670 -1896 670 -1896 0 2
rlabel polysilicon 667 -1902 667 -1902 0 3
rlabel polysilicon 670 -1902 670 -1902 0 4
rlabel polysilicon 674 -1896 674 -1896 0 1
rlabel polysilicon 674 -1902 674 -1902 0 3
rlabel polysilicon 681 -1896 681 -1896 0 1
rlabel polysilicon 681 -1902 681 -1902 0 3
rlabel polysilicon 688 -1896 688 -1896 0 1
rlabel polysilicon 688 -1902 688 -1902 0 3
rlabel polysilicon 695 -1896 695 -1896 0 1
rlabel polysilicon 695 -1902 695 -1902 0 3
rlabel polysilicon 702 -1896 702 -1896 0 1
rlabel polysilicon 702 -1902 702 -1902 0 3
rlabel polysilicon 709 -1896 709 -1896 0 1
rlabel polysilicon 709 -1902 709 -1902 0 3
rlabel polysilicon 716 -1896 716 -1896 0 1
rlabel polysilicon 716 -1902 716 -1902 0 3
rlabel polysilicon 723 -1896 723 -1896 0 1
rlabel polysilicon 723 -1902 723 -1902 0 3
rlabel polysilicon 730 -1896 730 -1896 0 1
rlabel polysilicon 733 -1896 733 -1896 0 2
rlabel polysilicon 730 -1902 730 -1902 0 3
rlabel polysilicon 737 -1896 737 -1896 0 1
rlabel polysilicon 737 -1902 737 -1902 0 3
rlabel polysilicon 744 -1896 744 -1896 0 1
rlabel polysilicon 744 -1902 744 -1902 0 3
rlabel polysilicon 751 -1896 751 -1896 0 1
rlabel polysilicon 751 -1902 751 -1902 0 3
rlabel polysilicon 758 -1896 758 -1896 0 1
rlabel polysilicon 758 -1902 758 -1902 0 3
rlabel polysilicon 765 -1896 765 -1896 0 1
rlabel polysilicon 765 -1902 765 -1902 0 3
rlabel polysilicon 772 -1896 772 -1896 0 1
rlabel polysilicon 772 -1902 772 -1902 0 3
rlabel polysilicon 779 -1896 779 -1896 0 1
rlabel polysilicon 779 -1902 779 -1902 0 3
rlabel polysilicon 786 -1896 786 -1896 0 1
rlabel polysilicon 786 -1902 786 -1902 0 3
rlabel polysilicon 793 -1896 793 -1896 0 1
rlabel polysilicon 793 -1902 793 -1902 0 3
rlabel polysilicon 800 -1896 800 -1896 0 1
rlabel polysilicon 800 -1902 800 -1902 0 3
rlabel polysilicon 807 -1896 807 -1896 0 1
rlabel polysilicon 807 -1902 807 -1902 0 3
rlabel polysilicon 814 -1896 814 -1896 0 1
rlabel polysilicon 814 -1902 814 -1902 0 3
rlabel polysilicon 821 -1896 821 -1896 0 1
rlabel polysilicon 821 -1902 821 -1902 0 3
rlabel polysilicon 828 -1896 828 -1896 0 1
rlabel polysilicon 828 -1902 828 -1902 0 3
rlabel polysilicon 835 -1896 835 -1896 0 1
rlabel polysilicon 835 -1902 835 -1902 0 3
rlabel polysilicon 842 -1896 842 -1896 0 1
rlabel polysilicon 842 -1902 842 -1902 0 3
rlabel polysilicon 849 -1896 849 -1896 0 1
rlabel polysilicon 849 -1902 849 -1902 0 3
rlabel polysilicon 856 -1896 856 -1896 0 1
rlabel polysilicon 856 -1902 856 -1902 0 3
rlabel polysilicon 863 -1896 863 -1896 0 1
rlabel polysilicon 863 -1902 863 -1902 0 3
rlabel polysilicon 870 -1896 870 -1896 0 1
rlabel polysilicon 870 -1902 870 -1902 0 3
rlabel polysilicon 877 -1896 877 -1896 0 1
rlabel polysilicon 877 -1902 877 -1902 0 3
rlabel polysilicon 884 -1896 884 -1896 0 1
rlabel polysilicon 884 -1902 884 -1902 0 3
rlabel polysilicon 891 -1896 891 -1896 0 1
rlabel polysilicon 891 -1902 891 -1902 0 3
rlabel polysilicon 898 -1896 898 -1896 0 1
rlabel polysilicon 898 -1902 898 -1902 0 3
rlabel polysilicon 905 -1896 905 -1896 0 1
rlabel polysilicon 905 -1902 905 -1902 0 3
rlabel polysilicon 912 -1896 912 -1896 0 1
rlabel polysilicon 912 -1902 912 -1902 0 3
rlabel polysilicon 919 -1896 919 -1896 0 1
rlabel polysilicon 919 -1902 919 -1902 0 3
rlabel polysilicon 926 -1896 926 -1896 0 1
rlabel polysilicon 926 -1902 926 -1902 0 3
rlabel polysilicon 933 -1896 933 -1896 0 1
rlabel polysilicon 933 -1902 933 -1902 0 3
rlabel polysilicon 940 -1896 940 -1896 0 1
rlabel polysilicon 940 -1902 940 -1902 0 3
rlabel polysilicon 947 -1896 947 -1896 0 1
rlabel polysilicon 947 -1902 947 -1902 0 3
rlabel polysilicon 954 -1896 954 -1896 0 1
rlabel polysilicon 954 -1902 954 -1902 0 3
rlabel polysilicon 961 -1896 961 -1896 0 1
rlabel polysilicon 961 -1902 961 -1902 0 3
rlabel polysilicon 968 -1896 968 -1896 0 1
rlabel polysilicon 968 -1902 968 -1902 0 3
rlabel polysilicon 975 -1896 975 -1896 0 1
rlabel polysilicon 975 -1902 975 -1902 0 3
rlabel polysilicon 982 -1896 982 -1896 0 1
rlabel polysilicon 982 -1902 982 -1902 0 3
rlabel polysilicon 989 -1896 989 -1896 0 1
rlabel polysilicon 989 -1902 989 -1902 0 3
rlabel polysilicon 996 -1896 996 -1896 0 1
rlabel polysilicon 996 -1902 996 -1902 0 3
rlabel polysilicon 1003 -1896 1003 -1896 0 1
rlabel polysilicon 1003 -1902 1003 -1902 0 3
rlabel polysilicon 1010 -1896 1010 -1896 0 1
rlabel polysilicon 1010 -1902 1010 -1902 0 3
rlabel polysilicon 1017 -1896 1017 -1896 0 1
rlabel polysilicon 1017 -1902 1017 -1902 0 3
rlabel polysilicon 1024 -1896 1024 -1896 0 1
rlabel polysilicon 1024 -1902 1024 -1902 0 3
rlabel polysilicon 1031 -1896 1031 -1896 0 1
rlabel polysilicon 1031 -1902 1031 -1902 0 3
rlabel polysilicon 1038 -1896 1038 -1896 0 1
rlabel polysilicon 1038 -1902 1038 -1902 0 3
rlabel polysilicon 1045 -1896 1045 -1896 0 1
rlabel polysilicon 1045 -1902 1045 -1902 0 3
rlabel polysilicon 1052 -1896 1052 -1896 0 1
rlabel polysilicon 1052 -1902 1052 -1902 0 3
rlabel polysilicon 1059 -1896 1059 -1896 0 1
rlabel polysilicon 1059 -1902 1059 -1902 0 3
rlabel polysilicon 1069 -1896 1069 -1896 0 2
rlabel polysilicon 1066 -1902 1066 -1902 0 3
rlabel polysilicon 1069 -1902 1069 -1902 0 4
rlabel polysilicon 1073 -1896 1073 -1896 0 1
rlabel polysilicon 1073 -1902 1073 -1902 0 3
rlabel polysilicon 1087 -1896 1087 -1896 0 1
rlabel polysilicon 1087 -1902 1087 -1902 0 3
rlabel polysilicon 1101 -1896 1101 -1896 0 1
rlabel polysilicon 1101 -1902 1101 -1902 0 3
rlabel polysilicon 2 -2001 2 -2001 0 1
rlabel polysilicon 9 -2001 9 -2001 0 1
rlabel polysilicon 9 -2007 9 -2007 0 3
rlabel polysilicon 16 -2001 16 -2001 0 1
rlabel polysilicon 16 -2007 16 -2007 0 3
rlabel polysilicon 23 -2001 23 -2001 0 1
rlabel polysilicon 26 -2007 26 -2007 0 4
rlabel polysilicon 30 -2001 30 -2001 0 1
rlabel polysilicon 33 -2001 33 -2001 0 2
rlabel polysilicon 30 -2007 30 -2007 0 3
rlabel polysilicon 33 -2007 33 -2007 0 4
rlabel polysilicon 37 -2001 37 -2001 0 1
rlabel polysilicon 37 -2007 37 -2007 0 3
rlabel polysilicon 44 -2001 44 -2001 0 1
rlabel polysilicon 44 -2007 44 -2007 0 3
rlabel polysilicon 54 -2001 54 -2001 0 2
rlabel polysilicon 51 -2007 51 -2007 0 3
rlabel polysilicon 54 -2007 54 -2007 0 4
rlabel polysilicon 58 -2001 58 -2001 0 1
rlabel polysilicon 61 -2001 61 -2001 0 2
rlabel polysilicon 58 -2007 58 -2007 0 3
rlabel polysilicon 65 -2001 65 -2001 0 1
rlabel polysilicon 65 -2007 65 -2007 0 3
rlabel polysilicon 75 -2001 75 -2001 0 2
rlabel polysilicon 75 -2007 75 -2007 0 4
rlabel polysilicon 79 -2007 79 -2007 0 3
rlabel polysilicon 86 -2007 86 -2007 0 3
rlabel polysilicon 89 -2007 89 -2007 0 4
rlabel polysilicon 93 -2001 93 -2001 0 1
rlabel polysilicon 93 -2007 93 -2007 0 3
rlabel polysilicon 100 -2001 100 -2001 0 1
rlabel polysilicon 100 -2007 100 -2007 0 3
rlabel polysilicon 107 -2001 107 -2001 0 1
rlabel polysilicon 107 -2007 107 -2007 0 3
rlabel polysilicon 110 -2007 110 -2007 0 4
rlabel polysilicon 114 -2001 114 -2001 0 1
rlabel polysilicon 114 -2007 114 -2007 0 3
rlabel polysilicon 121 -2001 121 -2001 0 1
rlabel polysilicon 121 -2007 121 -2007 0 3
rlabel polysilicon 128 -2001 128 -2001 0 1
rlabel polysilicon 128 -2007 128 -2007 0 3
rlabel polysilicon 135 -2007 135 -2007 0 3
rlabel polysilicon 138 -2007 138 -2007 0 4
rlabel polysilicon 142 -2001 142 -2001 0 1
rlabel polysilicon 142 -2007 142 -2007 0 3
rlabel polysilicon 149 -2001 149 -2001 0 1
rlabel polysilicon 152 -2001 152 -2001 0 2
rlabel polysilicon 149 -2007 149 -2007 0 3
rlabel polysilicon 152 -2007 152 -2007 0 4
rlabel polysilicon 156 -2001 156 -2001 0 1
rlabel polysilicon 156 -2007 156 -2007 0 3
rlabel polysilicon 163 -2001 163 -2001 0 1
rlabel polysilicon 163 -2007 163 -2007 0 3
rlabel polysilicon 170 -2001 170 -2001 0 1
rlabel polysilicon 170 -2007 170 -2007 0 3
rlabel polysilicon 180 -2001 180 -2001 0 2
rlabel polysilicon 177 -2007 177 -2007 0 3
rlabel polysilicon 180 -2007 180 -2007 0 4
rlabel polysilicon 184 -2001 184 -2001 0 1
rlabel polysilicon 184 -2007 184 -2007 0 3
rlabel polysilicon 191 -2001 191 -2001 0 1
rlabel polysilicon 191 -2007 191 -2007 0 3
rlabel polysilicon 198 -2001 198 -2001 0 1
rlabel polysilicon 198 -2007 198 -2007 0 3
rlabel polysilicon 205 -2001 205 -2001 0 1
rlabel polysilicon 208 -2001 208 -2001 0 2
rlabel polysilicon 212 -2001 212 -2001 0 1
rlabel polysilicon 212 -2007 212 -2007 0 3
rlabel polysilicon 219 -2001 219 -2001 0 1
rlabel polysilicon 222 -2001 222 -2001 0 2
rlabel polysilicon 222 -2007 222 -2007 0 4
rlabel polysilicon 229 -2001 229 -2001 0 2
rlabel polysilicon 226 -2007 226 -2007 0 3
rlabel polysilicon 229 -2007 229 -2007 0 4
rlabel polysilicon 233 -2001 233 -2001 0 1
rlabel polysilicon 233 -2007 233 -2007 0 3
rlabel polysilicon 240 -2001 240 -2001 0 1
rlabel polysilicon 240 -2007 240 -2007 0 3
rlabel polysilicon 247 -2001 247 -2001 0 1
rlabel polysilicon 247 -2007 247 -2007 0 3
rlabel polysilicon 254 -2001 254 -2001 0 1
rlabel polysilicon 254 -2007 254 -2007 0 3
rlabel polysilicon 261 -2001 261 -2001 0 1
rlabel polysilicon 261 -2007 261 -2007 0 3
rlabel polysilicon 268 -2001 268 -2001 0 1
rlabel polysilicon 268 -2007 268 -2007 0 3
rlabel polysilicon 275 -2001 275 -2001 0 1
rlabel polysilicon 275 -2007 275 -2007 0 3
rlabel polysilicon 282 -2001 282 -2001 0 1
rlabel polysilicon 282 -2007 282 -2007 0 3
rlabel polysilicon 289 -2001 289 -2001 0 1
rlabel polysilicon 289 -2007 289 -2007 0 3
rlabel polysilicon 296 -2001 296 -2001 0 1
rlabel polysilicon 296 -2007 296 -2007 0 3
rlabel polysilicon 303 -2001 303 -2001 0 1
rlabel polysilicon 303 -2007 303 -2007 0 3
rlabel polysilicon 310 -2001 310 -2001 0 1
rlabel polysilicon 310 -2007 310 -2007 0 3
rlabel polysilicon 317 -2001 317 -2001 0 1
rlabel polysilicon 317 -2007 317 -2007 0 3
rlabel polysilicon 324 -2001 324 -2001 0 1
rlabel polysilicon 324 -2007 324 -2007 0 3
rlabel polysilicon 331 -2001 331 -2001 0 1
rlabel polysilicon 331 -2007 331 -2007 0 3
rlabel polysilicon 338 -2001 338 -2001 0 1
rlabel polysilicon 338 -2007 338 -2007 0 3
rlabel polysilicon 345 -2001 345 -2001 0 1
rlabel polysilicon 348 -2001 348 -2001 0 2
rlabel polysilicon 345 -2007 345 -2007 0 3
rlabel polysilicon 348 -2007 348 -2007 0 4
rlabel polysilicon 352 -2001 352 -2001 0 1
rlabel polysilicon 352 -2007 352 -2007 0 3
rlabel polysilicon 359 -2001 359 -2001 0 1
rlabel polysilicon 359 -2007 359 -2007 0 3
rlabel polysilicon 366 -2001 366 -2001 0 1
rlabel polysilicon 369 -2001 369 -2001 0 2
rlabel polysilicon 366 -2007 366 -2007 0 3
rlabel polysilicon 369 -2007 369 -2007 0 4
rlabel polysilicon 373 -2001 373 -2001 0 1
rlabel polysilicon 376 -2001 376 -2001 0 2
rlabel polysilicon 373 -2007 373 -2007 0 3
rlabel polysilicon 376 -2007 376 -2007 0 4
rlabel polysilicon 380 -2001 380 -2001 0 1
rlabel polysilicon 380 -2007 380 -2007 0 3
rlabel polysilicon 387 -2001 387 -2001 0 1
rlabel polysilicon 387 -2007 387 -2007 0 3
rlabel polysilicon 394 -2001 394 -2001 0 1
rlabel polysilicon 394 -2007 394 -2007 0 3
rlabel polysilicon 401 -2001 401 -2001 0 1
rlabel polysilicon 401 -2007 401 -2007 0 3
rlabel polysilicon 408 -2001 408 -2001 0 1
rlabel polysilicon 408 -2007 408 -2007 0 3
rlabel polysilicon 411 -2007 411 -2007 0 4
rlabel polysilicon 415 -2001 415 -2001 0 1
rlabel polysilicon 415 -2007 415 -2007 0 3
rlabel polysilicon 422 -2001 422 -2001 0 1
rlabel polysilicon 422 -2007 422 -2007 0 3
rlabel polysilicon 429 -2001 429 -2001 0 1
rlabel polysilicon 429 -2007 429 -2007 0 3
rlabel polysilicon 436 -2001 436 -2001 0 1
rlabel polysilicon 439 -2007 439 -2007 0 4
rlabel polysilicon 443 -2001 443 -2001 0 1
rlabel polysilicon 443 -2007 443 -2007 0 3
rlabel polysilicon 450 -2001 450 -2001 0 1
rlabel polysilicon 450 -2007 450 -2007 0 3
rlabel polysilicon 457 -2001 457 -2001 0 1
rlabel polysilicon 457 -2007 457 -2007 0 3
rlabel polysilicon 464 -2001 464 -2001 0 1
rlabel polysilicon 464 -2007 464 -2007 0 3
rlabel polysilicon 471 -2001 471 -2001 0 1
rlabel polysilicon 471 -2007 471 -2007 0 3
rlabel polysilicon 478 -2001 478 -2001 0 1
rlabel polysilicon 478 -2007 478 -2007 0 3
rlabel polysilicon 485 -2001 485 -2001 0 1
rlabel polysilicon 485 -2007 485 -2007 0 3
rlabel polysilicon 492 -2001 492 -2001 0 1
rlabel polysilicon 492 -2007 492 -2007 0 3
rlabel polysilicon 499 -2001 499 -2001 0 1
rlabel polysilicon 499 -2007 499 -2007 0 3
rlabel polysilicon 506 -2001 506 -2001 0 1
rlabel polysilicon 506 -2007 506 -2007 0 3
rlabel polysilicon 516 -2001 516 -2001 0 2
rlabel polysilicon 516 -2007 516 -2007 0 4
rlabel polysilicon 520 -2001 520 -2001 0 1
rlabel polysilicon 520 -2007 520 -2007 0 3
rlabel polysilicon 527 -2001 527 -2001 0 1
rlabel polysilicon 530 -2001 530 -2001 0 2
rlabel polysilicon 527 -2007 527 -2007 0 3
rlabel polysilicon 530 -2007 530 -2007 0 4
rlabel polysilicon 534 -2001 534 -2001 0 1
rlabel polysilicon 534 -2007 534 -2007 0 3
rlabel polysilicon 541 -2001 541 -2001 0 1
rlabel polysilicon 541 -2007 541 -2007 0 3
rlabel polysilicon 548 -2001 548 -2001 0 1
rlabel polysilicon 548 -2007 548 -2007 0 3
rlabel polysilicon 555 -2001 555 -2001 0 1
rlabel polysilicon 555 -2007 555 -2007 0 3
rlabel polysilicon 562 -2001 562 -2001 0 1
rlabel polysilicon 562 -2007 562 -2007 0 3
rlabel polysilicon 569 -2001 569 -2001 0 1
rlabel polysilicon 569 -2007 569 -2007 0 3
rlabel polysilicon 576 -2001 576 -2001 0 1
rlabel polysilicon 576 -2007 576 -2007 0 3
rlabel polysilicon 583 -2001 583 -2001 0 1
rlabel polysilicon 583 -2007 583 -2007 0 3
rlabel polysilicon 590 -2007 590 -2007 0 3
rlabel polysilicon 593 -2007 593 -2007 0 4
rlabel polysilicon 597 -2001 597 -2001 0 1
rlabel polysilicon 597 -2007 597 -2007 0 3
rlabel polysilicon 604 -2001 604 -2001 0 1
rlabel polysilicon 604 -2007 604 -2007 0 3
rlabel polysilicon 611 -2001 611 -2001 0 1
rlabel polysilicon 611 -2007 611 -2007 0 3
rlabel polysilicon 618 -2001 618 -2001 0 1
rlabel polysilicon 621 -2001 621 -2001 0 2
rlabel polysilicon 618 -2007 618 -2007 0 3
rlabel polysilicon 625 -2001 625 -2001 0 1
rlabel polysilicon 625 -2007 625 -2007 0 3
rlabel polysilicon 635 -2001 635 -2001 0 2
rlabel polysilicon 635 -2007 635 -2007 0 4
rlabel polysilicon 639 -2001 639 -2001 0 1
rlabel polysilicon 639 -2007 639 -2007 0 3
rlabel polysilicon 646 -2001 646 -2001 0 1
rlabel polysilicon 649 -2001 649 -2001 0 2
rlabel polysilicon 646 -2007 646 -2007 0 3
rlabel polysilicon 649 -2007 649 -2007 0 4
rlabel polysilicon 653 -2001 653 -2001 0 1
rlabel polysilicon 653 -2007 653 -2007 0 3
rlabel polysilicon 660 -2001 660 -2001 0 1
rlabel polysilicon 660 -2007 660 -2007 0 3
rlabel polysilicon 667 -2001 667 -2001 0 1
rlabel polysilicon 667 -2007 667 -2007 0 3
rlabel polysilicon 674 -2001 674 -2001 0 1
rlabel polysilicon 674 -2007 674 -2007 0 3
rlabel polysilicon 681 -2001 681 -2001 0 1
rlabel polysilicon 681 -2007 681 -2007 0 3
rlabel polysilicon 688 -2001 688 -2001 0 1
rlabel polysilicon 688 -2007 688 -2007 0 3
rlabel polysilicon 695 -2001 695 -2001 0 1
rlabel polysilicon 695 -2007 695 -2007 0 3
rlabel polysilicon 702 -2001 702 -2001 0 1
rlabel polysilicon 702 -2007 702 -2007 0 3
rlabel polysilicon 709 -2001 709 -2001 0 1
rlabel polysilicon 709 -2007 709 -2007 0 3
rlabel polysilicon 716 -2001 716 -2001 0 1
rlabel polysilicon 716 -2007 716 -2007 0 3
rlabel polysilicon 723 -2001 723 -2001 0 1
rlabel polysilicon 723 -2007 723 -2007 0 3
rlabel polysilicon 730 -2001 730 -2001 0 1
rlabel polysilicon 730 -2007 730 -2007 0 3
rlabel polysilicon 737 -2001 737 -2001 0 1
rlabel polysilicon 737 -2007 737 -2007 0 3
rlabel polysilicon 744 -2007 744 -2007 0 3
rlabel polysilicon 751 -2001 751 -2001 0 1
rlabel polysilicon 751 -2007 751 -2007 0 3
rlabel polysilicon 758 -2001 758 -2001 0 1
rlabel polysilicon 758 -2007 758 -2007 0 3
rlabel polysilicon 765 -2001 765 -2001 0 1
rlabel polysilicon 768 -2001 768 -2001 0 2
rlabel polysilicon 765 -2007 765 -2007 0 3
rlabel polysilicon 768 -2007 768 -2007 0 4
rlabel polysilicon 772 -2001 772 -2001 0 1
rlabel polysilicon 772 -2007 772 -2007 0 3
rlabel polysilicon 779 -2007 779 -2007 0 3
rlabel polysilicon 782 -2007 782 -2007 0 4
rlabel polysilicon 786 -2001 786 -2001 0 1
rlabel polysilicon 786 -2007 786 -2007 0 3
rlabel polysilicon 793 -2001 793 -2001 0 1
rlabel polysilicon 793 -2007 793 -2007 0 3
rlabel polysilicon 800 -2001 800 -2001 0 1
rlabel polysilicon 800 -2007 800 -2007 0 3
rlabel polysilicon 807 -2001 807 -2001 0 1
rlabel polysilicon 807 -2007 807 -2007 0 3
rlabel polysilicon 814 -2001 814 -2001 0 1
rlabel polysilicon 814 -2007 814 -2007 0 3
rlabel polysilicon 821 -2001 821 -2001 0 1
rlabel polysilicon 821 -2007 821 -2007 0 3
rlabel polysilicon 828 -2001 828 -2001 0 1
rlabel polysilicon 828 -2007 828 -2007 0 3
rlabel polysilicon 835 -2001 835 -2001 0 1
rlabel polysilicon 835 -2007 835 -2007 0 3
rlabel polysilicon 842 -2001 842 -2001 0 1
rlabel polysilicon 842 -2007 842 -2007 0 3
rlabel polysilicon 849 -2001 849 -2001 0 1
rlabel polysilicon 849 -2007 849 -2007 0 3
rlabel polysilicon 856 -2001 856 -2001 0 1
rlabel polysilicon 856 -2007 856 -2007 0 3
rlabel polysilicon 863 -2001 863 -2001 0 1
rlabel polysilicon 863 -2007 863 -2007 0 3
rlabel polysilicon 870 -2001 870 -2001 0 1
rlabel polysilicon 870 -2007 870 -2007 0 3
rlabel polysilicon 877 -2001 877 -2001 0 1
rlabel polysilicon 877 -2007 877 -2007 0 3
rlabel polysilicon 884 -2001 884 -2001 0 1
rlabel polysilicon 884 -2007 884 -2007 0 3
rlabel polysilicon 891 -2001 891 -2001 0 1
rlabel polysilicon 891 -2007 891 -2007 0 3
rlabel polysilicon 898 -2001 898 -2001 0 1
rlabel polysilicon 898 -2007 898 -2007 0 3
rlabel polysilicon 905 -2001 905 -2001 0 1
rlabel polysilicon 905 -2007 905 -2007 0 3
rlabel polysilicon 912 -2001 912 -2001 0 1
rlabel polysilicon 912 -2007 912 -2007 0 3
rlabel polysilicon 919 -2001 919 -2001 0 1
rlabel polysilicon 919 -2007 919 -2007 0 3
rlabel polysilicon 929 -2007 929 -2007 0 4
rlabel polysilicon 933 -2001 933 -2001 0 1
rlabel polysilicon 933 -2007 933 -2007 0 3
rlabel polysilicon 940 -2001 940 -2001 0 1
rlabel polysilicon 940 -2007 940 -2007 0 3
rlabel polysilicon 947 -2001 947 -2001 0 1
rlabel polysilicon 947 -2007 947 -2007 0 3
rlabel polysilicon 954 -2001 954 -2001 0 1
rlabel polysilicon 954 -2007 954 -2007 0 3
rlabel polysilicon 961 -2001 961 -2001 0 1
rlabel polysilicon 961 -2007 961 -2007 0 3
rlabel polysilicon 968 -2001 968 -2001 0 1
rlabel polysilicon 968 -2007 968 -2007 0 3
rlabel polysilicon 975 -2001 975 -2001 0 1
rlabel polysilicon 975 -2007 975 -2007 0 3
rlabel polysilicon 982 -2001 982 -2001 0 1
rlabel polysilicon 982 -2007 982 -2007 0 3
rlabel polysilicon 989 -2001 989 -2001 0 1
rlabel polysilicon 989 -2007 989 -2007 0 3
rlabel polysilicon 996 -2001 996 -2001 0 1
rlabel polysilicon 996 -2007 996 -2007 0 3
rlabel polysilicon 1003 -2001 1003 -2001 0 1
rlabel polysilicon 1003 -2007 1003 -2007 0 3
rlabel polysilicon 1010 -2001 1010 -2001 0 1
rlabel polysilicon 1010 -2007 1010 -2007 0 3
rlabel polysilicon 1017 -2001 1017 -2001 0 1
rlabel polysilicon 1017 -2007 1017 -2007 0 3
rlabel polysilicon 1024 -2001 1024 -2001 0 1
rlabel polysilicon 1024 -2007 1024 -2007 0 3
rlabel polysilicon 1031 -2001 1031 -2001 0 1
rlabel polysilicon 1031 -2007 1031 -2007 0 3
rlabel polysilicon 1038 -2001 1038 -2001 0 1
rlabel polysilicon 1038 -2007 1038 -2007 0 3
rlabel polysilicon 1045 -2001 1045 -2001 0 1
rlabel polysilicon 1045 -2007 1045 -2007 0 3
rlabel polysilicon 1052 -2001 1052 -2001 0 1
rlabel polysilicon 1052 -2007 1052 -2007 0 3
rlabel polysilicon 1059 -2001 1059 -2001 0 1
rlabel polysilicon 1059 -2007 1059 -2007 0 3
rlabel polysilicon 1066 -2001 1066 -2001 0 1
rlabel polysilicon 1066 -2007 1066 -2007 0 3
rlabel polysilicon 1073 -2001 1073 -2001 0 1
rlabel polysilicon 1073 -2007 1073 -2007 0 3
rlabel polysilicon 1080 -2001 1080 -2001 0 1
rlabel polysilicon 1080 -2007 1080 -2007 0 3
rlabel polysilicon 1087 -2001 1087 -2001 0 1
rlabel polysilicon 1087 -2007 1087 -2007 0 3
rlabel polysilicon 1097 -2001 1097 -2001 0 2
rlabel polysilicon 1094 -2007 1094 -2007 0 3
rlabel polysilicon 1104 -2001 1104 -2001 0 2
rlabel polysilicon 1101 -2007 1101 -2007 0 3
rlabel polysilicon 1104 -2007 1104 -2007 0 4
rlabel polysilicon 1108 -2001 1108 -2001 0 1
rlabel polysilicon 1108 -2007 1108 -2007 0 3
rlabel polysilicon 1115 -2001 1115 -2001 0 1
rlabel polysilicon 1115 -2007 1115 -2007 0 3
rlabel polysilicon 2 -2114 2 -2114 0 1
rlabel polysilicon 2 -2120 2 -2120 0 3
rlabel polysilicon 9 -2114 9 -2114 0 1
rlabel polysilicon 9 -2120 9 -2120 0 3
rlabel polysilicon 16 -2114 16 -2114 0 1
rlabel polysilicon 16 -2120 16 -2120 0 3
rlabel polysilicon 23 -2114 23 -2114 0 1
rlabel polysilicon 23 -2120 23 -2120 0 3
rlabel polysilicon 30 -2114 30 -2114 0 1
rlabel polysilicon 30 -2120 30 -2120 0 3
rlabel polysilicon 37 -2114 37 -2114 0 1
rlabel polysilicon 37 -2120 37 -2120 0 3
rlabel polysilicon 44 -2114 44 -2114 0 1
rlabel polysilicon 44 -2120 44 -2120 0 3
rlabel polysilicon 51 -2114 51 -2114 0 1
rlabel polysilicon 51 -2120 51 -2120 0 3
rlabel polysilicon 58 -2114 58 -2114 0 1
rlabel polysilicon 58 -2120 58 -2120 0 3
rlabel polysilicon 61 -2120 61 -2120 0 4
rlabel polysilicon 65 -2114 65 -2114 0 1
rlabel polysilicon 65 -2120 65 -2120 0 3
rlabel polysilicon 72 -2114 72 -2114 0 1
rlabel polysilicon 75 -2114 75 -2114 0 2
rlabel polysilicon 72 -2120 72 -2120 0 3
rlabel polysilicon 75 -2120 75 -2120 0 4
rlabel polysilicon 79 -2114 79 -2114 0 1
rlabel polysilicon 82 -2114 82 -2114 0 2
rlabel polysilicon 79 -2120 79 -2120 0 3
rlabel polysilicon 82 -2120 82 -2120 0 4
rlabel polysilicon 86 -2114 86 -2114 0 1
rlabel polysilicon 89 -2114 89 -2114 0 2
rlabel polysilicon 86 -2120 86 -2120 0 3
rlabel polysilicon 89 -2120 89 -2120 0 4
rlabel polysilicon 93 -2114 93 -2114 0 1
rlabel polysilicon 96 -2114 96 -2114 0 2
rlabel polysilicon 93 -2120 93 -2120 0 3
rlabel polysilicon 96 -2120 96 -2120 0 4
rlabel polysilicon 100 -2114 100 -2114 0 1
rlabel polysilicon 100 -2120 100 -2120 0 3
rlabel polysilicon 107 -2114 107 -2114 0 1
rlabel polysilicon 110 -2114 110 -2114 0 2
rlabel polysilicon 107 -2120 107 -2120 0 3
rlabel polysilicon 110 -2120 110 -2120 0 4
rlabel polysilicon 114 -2114 114 -2114 0 1
rlabel polysilicon 117 -2114 117 -2114 0 2
rlabel polysilicon 117 -2120 117 -2120 0 4
rlabel polysilicon 121 -2114 121 -2114 0 1
rlabel polysilicon 121 -2120 121 -2120 0 3
rlabel polysilicon 124 -2120 124 -2120 0 4
rlabel polysilicon 128 -2114 128 -2114 0 1
rlabel polysilicon 128 -2120 128 -2120 0 3
rlabel polysilicon 135 -2114 135 -2114 0 1
rlabel polysilicon 138 -2114 138 -2114 0 2
rlabel polysilicon 138 -2120 138 -2120 0 4
rlabel polysilicon 142 -2114 142 -2114 0 1
rlabel polysilicon 142 -2120 142 -2120 0 3
rlabel polysilicon 149 -2114 149 -2114 0 1
rlabel polysilicon 152 -2114 152 -2114 0 2
rlabel polysilicon 149 -2120 149 -2120 0 3
rlabel polysilicon 152 -2120 152 -2120 0 4
rlabel polysilicon 156 -2114 156 -2114 0 1
rlabel polysilicon 156 -2120 156 -2120 0 3
rlabel polysilicon 163 -2114 163 -2114 0 1
rlabel polysilicon 163 -2120 163 -2120 0 3
rlabel polysilicon 170 -2114 170 -2114 0 1
rlabel polysilicon 170 -2120 170 -2120 0 3
rlabel polysilicon 177 -2114 177 -2114 0 1
rlabel polysilicon 177 -2120 177 -2120 0 3
rlabel polysilicon 184 -2114 184 -2114 0 1
rlabel polysilicon 184 -2120 184 -2120 0 3
rlabel polysilicon 191 -2114 191 -2114 0 1
rlabel polysilicon 191 -2120 191 -2120 0 3
rlabel polysilicon 198 -2114 198 -2114 0 1
rlabel polysilicon 198 -2120 198 -2120 0 3
rlabel polysilicon 205 -2114 205 -2114 0 1
rlabel polysilicon 205 -2120 205 -2120 0 3
rlabel polysilicon 212 -2114 212 -2114 0 1
rlabel polysilicon 212 -2120 212 -2120 0 3
rlabel polysilicon 222 -2114 222 -2114 0 2
rlabel polysilicon 226 -2114 226 -2114 0 1
rlabel polysilicon 226 -2120 226 -2120 0 3
rlabel polysilicon 233 -2114 233 -2114 0 1
rlabel polysilicon 233 -2120 233 -2120 0 3
rlabel polysilicon 240 -2114 240 -2114 0 1
rlabel polysilicon 240 -2120 240 -2120 0 3
rlabel polysilicon 247 -2114 247 -2114 0 1
rlabel polysilicon 247 -2120 247 -2120 0 3
rlabel polysilicon 254 -2114 254 -2114 0 1
rlabel polysilicon 254 -2120 254 -2120 0 3
rlabel polysilicon 261 -2114 261 -2114 0 1
rlabel polysilicon 261 -2120 261 -2120 0 3
rlabel polysilicon 268 -2114 268 -2114 0 1
rlabel polysilicon 268 -2120 268 -2120 0 3
rlabel polysilicon 275 -2114 275 -2114 0 1
rlabel polysilicon 275 -2120 275 -2120 0 3
rlabel polysilicon 282 -2114 282 -2114 0 1
rlabel polysilicon 282 -2120 282 -2120 0 3
rlabel polysilicon 289 -2114 289 -2114 0 1
rlabel polysilicon 289 -2120 289 -2120 0 3
rlabel polysilicon 292 -2120 292 -2120 0 4
rlabel polysilicon 296 -2114 296 -2114 0 1
rlabel polysilicon 296 -2120 296 -2120 0 3
rlabel polysilicon 303 -2114 303 -2114 0 1
rlabel polysilicon 303 -2120 303 -2120 0 3
rlabel polysilicon 310 -2114 310 -2114 0 1
rlabel polysilicon 310 -2120 310 -2120 0 3
rlabel polysilicon 317 -2114 317 -2114 0 1
rlabel polysilicon 317 -2120 317 -2120 0 3
rlabel polysilicon 324 -2114 324 -2114 0 1
rlabel polysilicon 324 -2120 324 -2120 0 3
rlabel polysilicon 331 -2114 331 -2114 0 1
rlabel polysilicon 331 -2120 331 -2120 0 3
rlabel polysilicon 338 -2114 338 -2114 0 1
rlabel polysilicon 341 -2114 341 -2114 0 2
rlabel polysilicon 338 -2120 338 -2120 0 3
rlabel polysilicon 341 -2120 341 -2120 0 4
rlabel polysilicon 345 -2114 345 -2114 0 1
rlabel polysilicon 345 -2120 345 -2120 0 3
rlabel polysilicon 352 -2114 352 -2114 0 1
rlabel polysilicon 355 -2114 355 -2114 0 2
rlabel polysilicon 359 -2114 359 -2114 0 1
rlabel polysilicon 359 -2120 359 -2120 0 3
rlabel polysilicon 366 -2114 366 -2114 0 1
rlabel polysilicon 366 -2120 366 -2120 0 3
rlabel polysilicon 373 -2114 373 -2114 0 1
rlabel polysilicon 373 -2120 373 -2120 0 3
rlabel polysilicon 380 -2114 380 -2114 0 1
rlabel polysilicon 380 -2120 380 -2120 0 3
rlabel polysilicon 387 -2114 387 -2114 0 1
rlabel polysilicon 387 -2120 387 -2120 0 3
rlabel polysilicon 394 -2114 394 -2114 0 1
rlabel polysilicon 394 -2120 394 -2120 0 3
rlabel polysilicon 401 -2114 401 -2114 0 1
rlabel polysilicon 401 -2120 401 -2120 0 3
rlabel polysilicon 411 -2114 411 -2114 0 2
rlabel polysilicon 408 -2120 408 -2120 0 3
rlabel polysilicon 415 -2114 415 -2114 0 1
rlabel polysilicon 418 -2114 418 -2114 0 2
rlabel polysilicon 415 -2120 415 -2120 0 3
rlabel polysilicon 418 -2120 418 -2120 0 4
rlabel polysilicon 422 -2114 422 -2114 0 1
rlabel polysilicon 422 -2120 422 -2120 0 3
rlabel polysilicon 429 -2114 429 -2114 0 1
rlabel polysilicon 429 -2120 429 -2120 0 3
rlabel polysilicon 436 -2114 436 -2114 0 1
rlabel polysilicon 436 -2120 436 -2120 0 3
rlabel polysilicon 443 -2114 443 -2114 0 1
rlabel polysilicon 443 -2120 443 -2120 0 3
rlabel polysilicon 450 -2114 450 -2114 0 1
rlabel polysilicon 453 -2114 453 -2114 0 2
rlabel polysilicon 453 -2120 453 -2120 0 4
rlabel polysilicon 460 -2114 460 -2114 0 2
rlabel polysilicon 464 -2114 464 -2114 0 1
rlabel polysilicon 464 -2120 464 -2120 0 3
rlabel polysilicon 471 -2114 471 -2114 0 1
rlabel polysilicon 471 -2120 471 -2120 0 3
rlabel polysilicon 478 -2114 478 -2114 0 1
rlabel polysilicon 478 -2120 478 -2120 0 3
rlabel polysilicon 485 -2114 485 -2114 0 1
rlabel polysilicon 485 -2120 485 -2120 0 3
rlabel polysilicon 492 -2114 492 -2114 0 1
rlabel polysilicon 492 -2120 492 -2120 0 3
rlabel polysilicon 499 -2114 499 -2114 0 1
rlabel polysilicon 502 -2114 502 -2114 0 2
rlabel polysilicon 506 -2114 506 -2114 0 1
rlabel polysilicon 506 -2120 506 -2120 0 3
rlabel polysilicon 513 -2114 513 -2114 0 1
rlabel polysilicon 513 -2120 513 -2120 0 3
rlabel polysilicon 520 -2114 520 -2114 0 1
rlabel polysilicon 520 -2120 520 -2120 0 3
rlabel polysilicon 527 -2114 527 -2114 0 1
rlabel polysilicon 527 -2120 527 -2120 0 3
rlabel polysilicon 530 -2120 530 -2120 0 4
rlabel polysilicon 534 -2114 534 -2114 0 1
rlabel polysilicon 534 -2120 534 -2120 0 3
rlabel polysilicon 541 -2114 541 -2114 0 1
rlabel polysilicon 541 -2120 541 -2120 0 3
rlabel polysilicon 548 -2114 548 -2114 0 1
rlabel polysilicon 548 -2120 548 -2120 0 3
rlabel polysilicon 551 -2120 551 -2120 0 4
rlabel polysilicon 555 -2114 555 -2114 0 1
rlabel polysilicon 555 -2120 555 -2120 0 3
rlabel polysilicon 562 -2114 562 -2114 0 1
rlabel polysilicon 562 -2120 562 -2120 0 3
rlabel polysilicon 572 -2114 572 -2114 0 2
rlabel polysilicon 569 -2120 569 -2120 0 3
rlabel polysilicon 579 -2114 579 -2114 0 2
rlabel polysilicon 576 -2120 576 -2120 0 3
rlabel polysilicon 579 -2120 579 -2120 0 4
rlabel polysilicon 583 -2114 583 -2114 0 1
rlabel polysilicon 583 -2120 583 -2120 0 3
rlabel polysilicon 590 -2114 590 -2114 0 1
rlabel polysilicon 590 -2120 590 -2120 0 3
rlabel polysilicon 597 -2114 597 -2114 0 1
rlabel polysilicon 597 -2120 597 -2120 0 3
rlabel polysilicon 604 -2114 604 -2114 0 1
rlabel polysilicon 604 -2120 604 -2120 0 3
rlabel polysilicon 614 -2114 614 -2114 0 2
rlabel polysilicon 611 -2120 611 -2120 0 3
rlabel polysilicon 618 -2114 618 -2114 0 1
rlabel polysilicon 618 -2120 618 -2120 0 3
rlabel polysilicon 625 -2120 625 -2120 0 3
rlabel polysilicon 628 -2120 628 -2120 0 4
rlabel polysilicon 632 -2114 632 -2114 0 1
rlabel polysilicon 632 -2120 632 -2120 0 3
rlabel polysilicon 639 -2114 639 -2114 0 1
rlabel polysilicon 642 -2114 642 -2114 0 2
rlabel polysilicon 639 -2120 639 -2120 0 3
rlabel polysilicon 642 -2120 642 -2120 0 4
rlabel polysilicon 646 -2114 646 -2114 0 1
rlabel polysilicon 646 -2120 646 -2120 0 3
rlabel polysilicon 653 -2114 653 -2114 0 1
rlabel polysilicon 656 -2120 656 -2120 0 4
rlabel polysilicon 660 -2114 660 -2114 0 1
rlabel polysilicon 660 -2120 660 -2120 0 3
rlabel polysilicon 667 -2114 667 -2114 0 1
rlabel polysilicon 667 -2120 667 -2120 0 3
rlabel polysilicon 674 -2114 674 -2114 0 1
rlabel polysilicon 674 -2120 674 -2120 0 3
rlabel polysilicon 681 -2114 681 -2114 0 1
rlabel polysilicon 681 -2120 681 -2120 0 3
rlabel polysilicon 688 -2114 688 -2114 0 1
rlabel polysilicon 691 -2114 691 -2114 0 2
rlabel polysilicon 691 -2120 691 -2120 0 4
rlabel polysilicon 695 -2114 695 -2114 0 1
rlabel polysilicon 695 -2120 695 -2120 0 3
rlabel polysilicon 702 -2114 702 -2114 0 1
rlabel polysilicon 702 -2120 702 -2120 0 3
rlabel polysilicon 709 -2114 709 -2114 0 1
rlabel polysilicon 709 -2120 709 -2120 0 3
rlabel polysilicon 716 -2114 716 -2114 0 1
rlabel polysilicon 716 -2120 716 -2120 0 3
rlabel polysilicon 723 -2114 723 -2114 0 1
rlabel polysilicon 723 -2120 723 -2120 0 3
rlabel polysilicon 730 -2114 730 -2114 0 1
rlabel polysilicon 730 -2120 730 -2120 0 3
rlabel polysilicon 737 -2114 737 -2114 0 1
rlabel polysilicon 737 -2120 737 -2120 0 3
rlabel polysilicon 740 -2120 740 -2120 0 4
rlabel polysilicon 744 -2114 744 -2114 0 1
rlabel polysilicon 744 -2120 744 -2120 0 3
rlabel polysilicon 751 -2114 751 -2114 0 1
rlabel polysilicon 751 -2120 751 -2120 0 3
rlabel polysilicon 758 -2114 758 -2114 0 1
rlabel polysilicon 761 -2114 761 -2114 0 2
rlabel polysilicon 758 -2120 758 -2120 0 3
rlabel polysilicon 761 -2120 761 -2120 0 4
rlabel polysilicon 765 -2114 765 -2114 0 1
rlabel polysilicon 765 -2120 765 -2120 0 3
rlabel polysilicon 772 -2114 772 -2114 0 1
rlabel polysilicon 772 -2120 772 -2120 0 3
rlabel polysilicon 779 -2114 779 -2114 0 1
rlabel polysilicon 779 -2120 779 -2120 0 3
rlabel polysilicon 786 -2114 786 -2114 0 1
rlabel polysilicon 786 -2120 786 -2120 0 3
rlabel polysilicon 793 -2114 793 -2114 0 1
rlabel polysilicon 793 -2120 793 -2120 0 3
rlabel polysilicon 800 -2114 800 -2114 0 1
rlabel polysilicon 800 -2120 800 -2120 0 3
rlabel polysilicon 807 -2114 807 -2114 0 1
rlabel polysilicon 807 -2120 807 -2120 0 3
rlabel polysilicon 814 -2114 814 -2114 0 1
rlabel polysilicon 814 -2120 814 -2120 0 3
rlabel polysilicon 821 -2114 821 -2114 0 1
rlabel polysilicon 821 -2120 821 -2120 0 3
rlabel polysilicon 828 -2114 828 -2114 0 1
rlabel polysilicon 828 -2120 828 -2120 0 3
rlabel polysilicon 835 -2114 835 -2114 0 1
rlabel polysilicon 835 -2120 835 -2120 0 3
rlabel polysilicon 842 -2114 842 -2114 0 1
rlabel polysilicon 842 -2120 842 -2120 0 3
rlabel polysilicon 849 -2114 849 -2114 0 1
rlabel polysilicon 849 -2120 849 -2120 0 3
rlabel polysilicon 856 -2114 856 -2114 0 1
rlabel polysilicon 856 -2120 856 -2120 0 3
rlabel polysilicon 863 -2114 863 -2114 0 1
rlabel polysilicon 863 -2120 863 -2120 0 3
rlabel polysilicon 870 -2114 870 -2114 0 1
rlabel polysilicon 870 -2120 870 -2120 0 3
rlabel polysilicon 877 -2114 877 -2114 0 1
rlabel polysilicon 877 -2120 877 -2120 0 3
rlabel polysilicon 884 -2114 884 -2114 0 1
rlabel polysilicon 884 -2120 884 -2120 0 3
rlabel polysilicon 891 -2114 891 -2114 0 1
rlabel polysilicon 891 -2120 891 -2120 0 3
rlabel polysilicon 898 -2114 898 -2114 0 1
rlabel polysilicon 898 -2120 898 -2120 0 3
rlabel polysilicon 905 -2114 905 -2114 0 1
rlabel polysilicon 905 -2120 905 -2120 0 3
rlabel polysilicon 912 -2114 912 -2114 0 1
rlabel polysilicon 912 -2120 912 -2120 0 3
rlabel polysilicon 919 -2114 919 -2114 0 1
rlabel polysilicon 919 -2120 919 -2120 0 3
rlabel polysilicon 926 -2114 926 -2114 0 1
rlabel polysilicon 926 -2120 926 -2120 0 3
rlabel polysilicon 933 -2114 933 -2114 0 1
rlabel polysilicon 933 -2120 933 -2120 0 3
rlabel polysilicon 943 -2114 943 -2114 0 2
rlabel polysilicon 947 -2114 947 -2114 0 1
rlabel polysilicon 947 -2120 947 -2120 0 3
rlabel polysilicon 954 -2114 954 -2114 0 1
rlabel polysilicon 954 -2120 954 -2120 0 3
rlabel polysilicon 961 -2114 961 -2114 0 1
rlabel polysilicon 961 -2120 961 -2120 0 3
rlabel polysilicon 968 -2114 968 -2114 0 1
rlabel polysilicon 968 -2120 968 -2120 0 3
rlabel polysilicon 975 -2114 975 -2114 0 1
rlabel polysilicon 975 -2120 975 -2120 0 3
rlabel polysilicon 982 -2114 982 -2114 0 1
rlabel polysilicon 982 -2120 982 -2120 0 3
rlabel polysilicon 989 -2114 989 -2114 0 1
rlabel polysilicon 989 -2120 989 -2120 0 3
rlabel polysilicon 996 -2114 996 -2114 0 1
rlabel polysilicon 996 -2120 996 -2120 0 3
rlabel polysilicon 1003 -2114 1003 -2114 0 1
rlabel polysilicon 1003 -2120 1003 -2120 0 3
rlabel polysilicon 1010 -2114 1010 -2114 0 1
rlabel polysilicon 1010 -2120 1010 -2120 0 3
rlabel polysilicon 1017 -2114 1017 -2114 0 1
rlabel polysilicon 1017 -2120 1017 -2120 0 3
rlabel polysilicon 1024 -2114 1024 -2114 0 1
rlabel polysilicon 1024 -2120 1024 -2120 0 3
rlabel polysilicon 1031 -2114 1031 -2114 0 1
rlabel polysilicon 1031 -2120 1031 -2120 0 3
rlabel polysilicon 1038 -2114 1038 -2114 0 1
rlabel polysilicon 1038 -2120 1038 -2120 0 3
rlabel polysilicon 1045 -2114 1045 -2114 0 1
rlabel polysilicon 1045 -2120 1045 -2120 0 3
rlabel polysilicon 1052 -2114 1052 -2114 0 1
rlabel polysilicon 1052 -2120 1052 -2120 0 3
rlabel polysilicon 1059 -2114 1059 -2114 0 1
rlabel polysilicon 1059 -2120 1059 -2120 0 3
rlabel polysilicon 1066 -2114 1066 -2114 0 1
rlabel polysilicon 1066 -2120 1066 -2120 0 3
rlabel polysilicon 1073 -2114 1073 -2114 0 1
rlabel polysilicon 1073 -2120 1073 -2120 0 3
rlabel polysilicon 1080 -2114 1080 -2114 0 1
rlabel polysilicon 1080 -2120 1080 -2120 0 3
rlabel polysilicon 1087 -2114 1087 -2114 0 1
rlabel polysilicon 1087 -2120 1087 -2120 0 3
rlabel polysilicon 1094 -2114 1094 -2114 0 1
rlabel polysilicon 1094 -2120 1094 -2120 0 3
rlabel polysilicon 1101 -2114 1101 -2114 0 1
rlabel polysilicon 1101 -2120 1101 -2120 0 3
rlabel polysilicon 1108 -2114 1108 -2114 0 1
rlabel polysilicon 1108 -2120 1108 -2120 0 3
rlabel polysilicon 1115 -2114 1115 -2114 0 1
rlabel polysilicon 1115 -2120 1115 -2120 0 3
rlabel polysilicon 1122 -2114 1122 -2114 0 1
rlabel polysilicon 1122 -2120 1122 -2120 0 3
rlabel polysilicon 2 -2209 2 -2209 0 1
rlabel polysilicon 2 -2215 2 -2215 0 3
rlabel polysilicon 9 -2209 9 -2209 0 1
rlabel polysilicon 9 -2215 9 -2215 0 3
rlabel polysilicon 16 -2209 16 -2209 0 1
rlabel polysilicon 16 -2215 16 -2215 0 3
rlabel polysilicon 23 -2209 23 -2209 0 1
rlabel polysilicon 23 -2215 23 -2215 0 3
rlabel polysilicon 30 -2215 30 -2215 0 3
rlabel polysilicon 33 -2215 33 -2215 0 4
rlabel polysilicon 40 -2209 40 -2209 0 2
rlabel polysilicon 37 -2215 37 -2215 0 3
rlabel polysilicon 44 -2209 44 -2209 0 1
rlabel polysilicon 44 -2215 44 -2215 0 3
rlabel polysilicon 51 -2209 51 -2209 0 1
rlabel polysilicon 51 -2215 51 -2215 0 3
rlabel polysilicon 58 -2209 58 -2209 0 1
rlabel polysilicon 58 -2215 58 -2215 0 3
rlabel polysilicon 65 -2209 65 -2209 0 1
rlabel polysilicon 65 -2215 65 -2215 0 3
rlabel polysilicon 72 -2209 72 -2209 0 1
rlabel polysilicon 75 -2209 75 -2209 0 2
rlabel polysilicon 79 -2209 79 -2209 0 1
rlabel polysilicon 79 -2215 79 -2215 0 3
rlabel polysilicon 86 -2209 86 -2209 0 1
rlabel polysilicon 86 -2215 86 -2215 0 3
rlabel polysilicon 93 -2209 93 -2209 0 1
rlabel polysilicon 93 -2215 93 -2215 0 3
rlabel polysilicon 100 -2209 100 -2209 0 1
rlabel polysilicon 100 -2215 100 -2215 0 3
rlabel polysilicon 107 -2209 107 -2209 0 1
rlabel polysilicon 107 -2215 107 -2215 0 3
rlabel polysilicon 114 -2209 114 -2209 0 1
rlabel polysilicon 114 -2215 114 -2215 0 3
rlabel polysilicon 121 -2209 121 -2209 0 1
rlabel polysilicon 124 -2209 124 -2209 0 2
rlabel polysilicon 121 -2215 121 -2215 0 3
rlabel polysilicon 128 -2209 128 -2209 0 1
rlabel polysilicon 128 -2215 128 -2215 0 3
rlabel polysilicon 135 -2209 135 -2209 0 1
rlabel polysilicon 135 -2215 135 -2215 0 3
rlabel polysilicon 142 -2209 142 -2209 0 1
rlabel polysilicon 142 -2215 142 -2215 0 3
rlabel polysilicon 149 -2209 149 -2209 0 1
rlabel polysilicon 149 -2215 149 -2215 0 3
rlabel polysilicon 156 -2209 156 -2209 0 1
rlabel polysilicon 156 -2215 156 -2215 0 3
rlabel polysilicon 166 -2209 166 -2209 0 2
rlabel polysilicon 163 -2215 163 -2215 0 3
rlabel polysilicon 166 -2215 166 -2215 0 4
rlabel polysilicon 173 -2209 173 -2209 0 2
rlabel polysilicon 173 -2215 173 -2215 0 4
rlabel polysilicon 177 -2209 177 -2209 0 1
rlabel polysilicon 187 -2215 187 -2215 0 4
rlabel polysilicon 191 -2209 191 -2209 0 1
rlabel polysilicon 194 -2215 194 -2215 0 4
rlabel polysilicon 198 -2209 198 -2209 0 1
rlabel polysilicon 198 -2215 198 -2215 0 3
rlabel polysilicon 205 -2209 205 -2209 0 1
rlabel polysilicon 205 -2215 205 -2215 0 3
rlabel polysilicon 208 -2215 208 -2215 0 4
rlabel polysilicon 212 -2209 212 -2209 0 1
rlabel polysilicon 212 -2215 212 -2215 0 3
rlabel polysilicon 219 -2209 219 -2209 0 1
rlabel polysilicon 219 -2215 219 -2215 0 3
rlabel polysilicon 226 -2209 226 -2209 0 1
rlabel polysilicon 226 -2215 226 -2215 0 3
rlabel polysilicon 233 -2209 233 -2209 0 1
rlabel polysilicon 233 -2215 233 -2215 0 3
rlabel polysilicon 240 -2209 240 -2209 0 1
rlabel polysilicon 240 -2215 240 -2215 0 3
rlabel polysilicon 247 -2209 247 -2209 0 1
rlabel polysilicon 247 -2215 247 -2215 0 3
rlabel polysilicon 254 -2209 254 -2209 0 1
rlabel polysilicon 254 -2215 254 -2215 0 3
rlabel polysilicon 261 -2209 261 -2209 0 1
rlabel polysilicon 261 -2215 261 -2215 0 3
rlabel polysilicon 268 -2209 268 -2209 0 1
rlabel polysilicon 268 -2215 268 -2215 0 3
rlabel polysilicon 275 -2209 275 -2209 0 1
rlabel polysilicon 275 -2215 275 -2215 0 3
rlabel polysilicon 282 -2209 282 -2209 0 1
rlabel polysilicon 282 -2215 282 -2215 0 3
rlabel polysilicon 289 -2209 289 -2209 0 1
rlabel polysilicon 289 -2215 289 -2215 0 3
rlabel polysilicon 296 -2209 296 -2209 0 1
rlabel polysilicon 296 -2215 296 -2215 0 3
rlabel polysilicon 303 -2209 303 -2209 0 1
rlabel polysilicon 303 -2215 303 -2215 0 3
rlabel polysilicon 310 -2209 310 -2209 0 1
rlabel polysilicon 310 -2215 310 -2215 0 3
rlabel polysilicon 320 -2209 320 -2209 0 2
rlabel polysilicon 317 -2215 317 -2215 0 3
rlabel polysilicon 324 -2209 324 -2209 0 1
rlabel polysilicon 324 -2215 324 -2215 0 3
rlabel polysilicon 331 -2209 331 -2209 0 1
rlabel polysilicon 331 -2215 331 -2215 0 3
rlabel polysilicon 338 -2209 338 -2209 0 1
rlabel polysilicon 341 -2209 341 -2209 0 2
rlabel polysilicon 338 -2215 338 -2215 0 3
rlabel polysilicon 341 -2215 341 -2215 0 4
rlabel polysilicon 345 -2209 345 -2209 0 1
rlabel polysilicon 345 -2215 345 -2215 0 3
rlabel polysilicon 355 -2209 355 -2209 0 2
rlabel polysilicon 352 -2215 352 -2215 0 3
rlabel polysilicon 355 -2215 355 -2215 0 4
rlabel polysilicon 359 -2209 359 -2209 0 1
rlabel polysilicon 359 -2215 359 -2215 0 3
rlabel polysilicon 366 -2209 366 -2209 0 1
rlabel polysilicon 366 -2215 366 -2215 0 3
rlabel polysilicon 376 -2209 376 -2209 0 2
rlabel polysilicon 380 -2209 380 -2209 0 1
rlabel polysilicon 380 -2215 380 -2215 0 3
rlabel polysilicon 387 -2209 387 -2209 0 1
rlabel polysilicon 387 -2215 387 -2215 0 3
rlabel polysilicon 397 -2209 397 -2209 0 2
rlabel polysilicon 394 -2215 394 -2215 0 3
rlabel polysilicon 397 -2215 397 -2215 0 4
rlabel polysilicon 401 -2209 401 -2209 0 1
rlabel polysilicon 401 -2215 401 -2215 0 3
rlabel polysilicon 408 -2209 408 -2209 0 1
rlabel polysilicon 408 -2215 408 -2215 0 3
rlabel polysilicon 415 -2209 415 -2209 0 1
rlabel polysilicon 415 -2215 415 -2215 0 3
rlabel polysilicon 422 -2209 422 -2209 0 1
rlabel polysilicon 422 -2215 422 -2215 0 3
rlabel polysilicon 429 -2209 429 -2209 0 1
rlabel polysilicon 432 -2209 432 -2209 0 2
rlabel polysilicon 429 -2215 429 -2215 0 3
rlabel polysilicon 436 -2209 436 -2209 0 1
rlabel polysilicon 439 -2209 439 -2209 0 2
rlabel polysilicon 439 -2215 439 -2215 0 4
rlabel polysilicon 443 -2209 443 -2209 0 1
rlabel polysilicon 443 -2215 443 -2215 0 3
rlabel polysilicon 450 -2209 450 -2209 0 1
rlabel polysilicon 450 -2215 450 -2215 0 3
rlabel polysilicon 457 -2209 457 -2209 0 1
rlabel polysilicon 457 -2215 457 -2215 0 3
rlabel polysilicon 464 -2209 464 -2209 0 1
rlabel polysilicon 464 -2215 464 -2215 0 3
rlabel polysilicon 471 -2209 471 -2209 0 1
rlabel polysilicon 471 -2215 471 -2215 0 3
rlabel polysilicon 478 -2209 478 -2209 0 1
rlabel polysilicon 478 -2215 478 -2215 0 3
rlabel polysilicon 485 -2209 485 -2209 0 1
rlabel polysilicon 485 -2215 485 -2215 0 3
rlabel polysilicon 492 -2209 492 -2209 0 1
rlabel polysilicon 492 -2215 492 -2215 0 3
rlabel polysilicon 499 -2209 499 -2209 0 1
rlabel polysilicon 502 -2209 502 -2209 0 2
rlabel polysilicon 502 -2215 502 -2215 0 4
rlabel polysilicon 509 -2209 509 -2209 0 2
rlabel polysilicon 509 -2215 509 -2215 0 4
rlabel polysilicon 513 -2209 513 -2209 0 1
rlabel polysilicon 513 -2215 513 -2215 0 3
rlabel polysilicon 520 -2209 520 -2209 0 1
rlabel polysilicon 523 -2209 523 -2209 0 2
rlabel polysilicon 523 -2215 523 -2215 0 4
rlabel polysilicon 527 -2209 527 -2209 0 1
rlabel polysilicon 527 -2215 527 -2215 0 3
rlabel polysilicon 534 -2209 534 -2209 0 1
rlabel polysilicon 534 -2215 534 -2215 0 3
rlabel polysilicon 541 -2209 541 -2209 0 1
rlabel polysilicon 541 -2215 541 -2215 0 3
rlabel polysilicon 548 -2209 548 -2209 0 1
rlabel polysilicon 548 -2215 548 -2215 0 3
rlabel polysilicon 555 -2209 555 -2209 0 1
rlabel polysilicon 555 -2215 555 -2215 0 3
rlabel polysilicon 565 -2209 565 -2209 0 2
rlabel polysilicon 565 -2215 565 -2215 0 4
rlabel polysilicon 572 -2209 572 -2209 0 2
rlabel polysilicon 572 -2215 572 -2215 0 4
rlabel polysilicon 576 -2209 576 -2209 0 1
rlabel polysilicon 576 -2215 576 -2215 0 3
rlabel polysilicon 583 -2209 583 -2209 0 1
rlabel polysilicon 583 -2215 583 -2215 0 3
rlabel polysilicon 590 -2209 590 -2209 0 1
rlabel polysilicon 593 -2209 593 -2209 0 2
rlabel polysilicon 590 -2215 590 -2215 0 3
rlabel polysilicon 593 -2215 593 -2215 0 4
rlabel polysilicon 597 -2209 597 -2209 0 1
rlabel polysilicon 600 -2209 600 -2209 0 2
rlabel polysilicon 604 -2209 604 -2209 0 1
rlabel polysilicon 607 -2209 607 -2209 0 2
rlabel polysilicon 604 -2215 604 -2215 0 3
rlabel polysilicon 611 -2209 611 -2209 0 1
rlabel polysilicon 611 -2215 611 -2215 0 3
rlabel polysilicon 618 -2209 618 -2209 0 1
rlabel polysilicon 618 -2215 618 -2215 0 3
rlabel polysilicon 625 -2209 625 -2209 0 1
rlabel polysilicon 625 -2215 625 -2215 0 3
rlabel polysilicon 632 -2209 632 -2209 0 1
rlabel polysilicon 632 -2215 632 -2215 0 3
rlabel polysilicon 639 -2209 639 -2209 0 1
rlabel polysilicon 639 -2215 639 -2215 0 3
rlabel polysilicon 646 -2209 646 -2209 0 1
rlabel polysilicon 646 -2215 646 -2215 0 3
rlabel polysilicon 653 -2209 653 -2209 0 1
rlabel polysilicon 653 -2215 653 -2215 0 3
rlabel polysilicon 660 -2209 660 -2209 0 1
rlabel polysilicon 660 -2215 660 -2215 0 3
rlabel polysilicon 667 -2209 667 -2209 0 1
rlabel polysilicon 670 -2209 670 -2209 0 2
rlabel polysilicon 670 -2215 670 -2215 0 4
rlabel polysilicon 674 -2209 674 -2209 0 1
rlabel polysilicon 674 -2215 674 -2215 0 3
rlabel polysilicon 684 -2209 684 -2209 0 2
rlabel polysilicon 681 -2215 681 -2215 0 3
rlabel polysilicon 684 -2215 684 -2215 0 4
rlabel polysilicon 688 -2209 688 -2209 0 1
rlabel polysilicon 691 -2215 691 -2215 0 4
rlabel polysilicon 695 -2209 695 -2209 0 1
rlabel polysilicon 698 -2209 698 -2209 0 2
rlabel polysilicon 695 -2215 695 -2215 0 3
rlabel polysilicon 698 -2215 698 -2215 0 4
rlabel polysilicon 702 -2209 702 -2209 0 1
rlabel polysilicon 702 -2215 702 -2215 0 3
rlabel polysilicon 709 -2209 709 -2209 0 1
rlabel polysilicon 709 -2215 709 -2215 0 3
rlabel polysilicon 716 -2209 716 -2209 0 1
rlabel polysilicon 716 -2215 716 -2215 0 3
rlabel polysilicon 723 -2209 723 -2209 0 1
rlabel polysilicon 726 -2209 726 -2209 0 2
rlabel polysilicon 723 -2215 723 -2215 0 3
rlabel polysilicon 726 -2215 726 -2215 0 4
rlabel polysilicon 730 -2209 730 -2209 0 1
rlabel polysilicon 730 -2215 730 -2215 0 3
rlabel polysilicon 737 -2209 737 -2209 0 1
rlabel polysilicon 737 -2215 737 -2215 0 3
rlabel polysilicon 744 -2209 744 -2209 0 1
rlabel polysilicon 744 -2215 744 -2215 0 3
rlabel polysilicon 751 -2209 751 -2209 0 1
rlabel polysilicon 751 -2215 751 -2215 0 3
rlabel polysilicon 758 -2209 758 -2209 0 1
rlabel polysilicon 758 -2215 758 -2215 0 3
rlabel polysilicon 765 -2209 765 -2209 0 1
rlabel polysilicon 765 -2215 765 -2215 0 3
rlabel polysilicon 772 -2209 772 -2209 0 1
rlabel polysilicon 772 -2215 772 -2215 0 3
rlabel polysilicon 779 -2209 779 -2209 0 1
rlabel polysilicon 779 -2215 779 -2215 0 3
rlabel polysilicon 786 -2209 786 -2209 0 1
rlabel polysilicon 786 -2215 786 -2215 0 3
rlabel polysilicon 793 -2209 793 -2209 0 1
rlabel polysilicon 793 -2215 793 -2215 0 3
rlabel polysilicon 800 -2209 800 -2209 0 1
rlabel polysilicon 800 -2215 800 -2215 0 3
rlabel polysilicon 807 -2209 807 -2209 0 1
rlabel polysilicon 807 -2215 807 -2215 0 3
rlabel polysilicon 814 -2209 814 -2209 0 1
rlabel polysilicon 814 -2215 814 -2215 0 3
rlabel polysilicon 821 -2209 821 -2209 0 1
rlabel polysilicon 821 -2215 821 -2215 0 3
rlabel polysilicon 828 -2209 828 -2209 0 1
rlabel polysilicon 828 -2215 828 -2215 0 3
rlabel polysilicon 835 -2209 835 -2209 0 1
rlabel polysilicon 835 -2215 835 -2215 0 3
rlabel polysilicon 842 -2209 842 -2209 0 1
rlabel polysilicon 842 -2215 842 -2215 0 3
rlabel polysilicon 849 -2209 849 -2209 0 1
rlabel polysilicon 849 -2215 849 -2215 0 3
rlabel polysilicon 856 -2209 856 -2209 0 1
rlabel polysilicon 856 -2215 856 -2215 0 3
rlabel polysilicon 863 -2209 863 -2209 0 1
rlabel polysilicon 863 -2215 863 -2215 0 3
rlabel polysilicon 873 -2209 873 -2209 0 2
rlabel polysilicon 877 -2209 877 -2209 0 1
rlabel polysilicon 877 -2215 877 -2215 0 3
rlabel polysilicon 884 -2209 884 -2209 0 1
rlabel polysilicon 884 -2215 884 -2215 0 3
rlabel polysilicon 891 -2209 891 -2209 0 1
rlabel polysilicon 891 -2215 891 -2215 0 3
rlabel polysilicon 898 -2209 898 -2209 0 1
rlabel polysilicon 898 -2215 898 -2215 0 3
rlabel polysilicon 905 -2209 905 -2209 0 1
rlabel polysilicon 905 -2215 905 -2215 0 3
rlabel polysilicon 912 -2209 912 -2209 0 1
rlabel polysilicon 912 -2215 912 -2215 0 3
rlabel polysilicon 919 -2209 919 -2209 0 1
rlabel polysilicon 919 -2215 919 -2215 0 3
rlabel polysilicon 926 -2209 926 -2209 0 1
rlabel polysilicon 926 -2215 926 -2215 0 3
rlabel polysilicon 933 -2209 933 -2209 0 1
rlabel polysilicon 933 -2215 933 -2215 0 3
rlabel polysilicon 940 -2209 940 -2209 0 1
rlabel polysilicon 940 -2215 940 -2215 0 3
rlabel polysilicon 947 -2209 947 -2209 0 1
rlabel polysilicon 947 -2215 947 -2215 0 3
rlabel polysilicon 954 -2209 954 -2209 0 1
rlabel polysilicon 954 -2215 954 -2215 0 3
rlabel polysilicon 961 -2209 961 -2209 0 1
rlabel polysilicon 961 -2215 961 -2215 0 3
rlabel polysilicon 968 -2209 968 -2209 0 1
rlabel polysilicon 968 -2215 968 -2215 0 3
rlabel polysilicon 975 -2209 975 -2209 0 1
rlabel polysilicon 975 -2215 975 -2215 0 3
rlabel polysilicon 982 -2209 982 -2209 0 1
rlabel polysilicon 982 -2215 982 -2215 0 3
rlabel polysilicon 989 -2209 989 -2209 0 1
rlabel polysilicon 989 -2215 989 -2215 0 3
rlabel polysilicon 996 -2209 996 -2209 0 1
rlabel polysilicon 996 -2215 996 -2215 0 3
rlabel polysilicon 1003 -2209 1003 -2209 0 1
rlabel polysilicon 1003 -2215 1003 -2215 0 3
rlabel polysilicon 1010 -2209 1010 -2209 0 1
rlabel polysilicon 1010 -2215 1010 -2215 0 3
rlabel polysilicon 1017 -2209 1017 -2209 0 1
rlabel polysilicon 1017 -2215 1017 -2215 0 3
rlabel polysilicon 1024 -2209 1024 -2209 0 1
rlabel polysilicon 1024 -2215 1024 -2215 0 3
rlabel polysilicon 1031 -2209 1031 -2209 0 1
rlabel polysilicon 1031 -2215 1031 -2215 0 3
rlabel polysilicon 1038 -2209 1038 -2209 0 1
rlabel polysilicon 1038 -2215 1038 -2215 0 3
rlabel polysilicon 1045 -2209 1045 -2209 0 1
rlabel polysilicon 1045 -2215 1045 -2215 0 3
rlabel polysilicon 1055 -2209 1055 -2209 0 2
rlabel polysilicon 2 -2278 2 -2278 0 1
rlabel polysilicon 2 -2284 2 -2284 0 3
rlabel polysilicon 9 -2278 9 -2278 0 1
rlabel polysilicon 9 -2284 9 -2284 0 3
rlabel polysilicon 16 -2278 16 -2278 0 1
rlabel polysilicon 16 -2284 16 -2284 0 3
rlabel polysilicon 23 -2278 23 -2278 0 1
rlabel polysilicon 23 -2284 23 -2284 0 3
rlabel polysilicon 30 -2278 30 -2278 0 1
rlabel polysilicon 30 -2284 30 -2284 0 3
rlabel polysilicon 37 -2278 37 -2278 0 1
rlabel polysilicon 37 -2284 37 -2284 0 3
rlabel polysilicon 44 -2278 44 -2278 0 1
rlabel polysilicon 44 -2284 44 -2284 0 3
rlabel polysilicon 51 -2278 51 -2278 0 1
rlabel polysilicon 51 -2284 51 -2284 0 3
rlabel polysilicon 54 -2284 54 -2284 0 4
rlabel polysilicon 58 -2278 58 -2278 0 1
rlabel polysilicon 58 -2284 58 -2284 0 3
rlabel polysilicon 61 -2284 61 -2284 0 4
rlabel polysilicon 65 -2278 65 -2278 0 1
rlabel polysilicon 65 -2284 65 -2284 0 3
rlabel polysilicon 72 -2278 72 -2278 0 1
rlabel polysilicon 72 -2284 72 -2284 0 3
rlabel polysilicon 79 -2284 79 -2284 0 3
rlabel polysilicon 82 -2284 82 -2284 0 4
rlabel polysilicon 86 -2278 86 -2278 0 1
rlabel polysilicon 86 -2284 86 -2284 0 3
rlabel polysilicon 93 -2278 93 -2278 0 1
rlabel polysilicon 93 -2284 93 -2284 0 3
rlabel polysilicon 103 -2278 103 -2278 0 2
rlabel polysilicon 100 -2284 100 -2284 0 3
rlabel polysilicon 103 -2284 103 -2284 0 4
rlabel polysilicon 107 -2278 107 -2278 0 1
rlabel polysilicon 107 -2284 107 -2284 0 3
rlabel polysilicon 110 -2284 110 -2284 0 4
rlabel polysilicon 114 -2278 114 -2278 0 1
rlabel polysilicon 114 -2284 114 -2284 0 3
rlabel polysilicon 121 -2278 121 -2278 0 1
rlabel polysilicon 121 -2284 121 -2284 0 3
rlabel polysilicon 128 -2284 128 -2284 0 3
rlabel polysilicon 131 -2284 131 -2284 0 4
rlabel polysilicon 135 -2278 135 -2278 0 1
rlabel polysilicon 135 -2284 135 -2284 0 3
rlabel polysilicon 142 -2278 142 -2278 0 1
rlabel polysilicon 142 -2284 142 -2284 0 3
rlabel polysilicon 149 -2278 149 -2278 0 1
rlabel polysilicon 149 -2284 149 -2284 0 3
rlabel polysilicon 156 -2278 156 -2278 0 1
rlabel polysilicon 156 -2284 156 -2284 0 3
rlabel polysilicon 163 -2278 163 -2278 0 1
rlabel polysilicon 163 -2284 163 -2284 0 3
rlabel polysilicon 170 -2278 170 -2278 0 1
rlabel polysilicon 170 -2284 170 -2284 0 3
rlabel polysilicon 177 -2278 177 -2278 0 1
rlabel polysilicon 177 -2284 177 -2284 0 3
rlabel polysilicon 180 -2284 180 -2284 0 4
rlabel polysilicon 184 -2278 184 -2278 0 1
rlabel polysilicon 184 -2284 184 -2284 0 3
rlabel polysilicon 191 -2278 191 -2278 0 1
rlabel polysilicon 191 -2284 191 -2284 0 3
rlabel polysilicon 198 -2278 198 -2278 0 1
rlabel polysilicon 201 -2278 201 -2278 0 2
rlabel polysilicon 198 -2284 198 -2284 0 3
rlabel polysilicon 205 -2278 205 -2278 0 1
rlabel polysilicon 205 -2284 205 -2284 0 3
rlabel polysilicon 212 -2278 212 -2278 0 1
rlabel polysilicon 215 -2278 215 -2278 0 2
rlabel polysilicon 215 -2284 215 -2284 0 4
rlabel polysilicon 219 -2278 219 -2278 0 1
rlabel polysilicon 226 -2278 226 -2278 0 1
rlabel polysilicon 226 -2284 226 -2284 0 3
rlabel polysilicon 233 -2278 233 -2278 0 1
rlabel polysilicon 233 -2284 233 -2284 0 3
rlabel polysilicon 240 -2278 240 -2278 0 1
rlabel polysilicon 240 -2284 240 -2284 0 3
rlabel polysilicon 247 -2278 247 -2278 0 1
rlabel polysilicon 247 -2284 247 -2284 0 3
rlabel polysilicon 254 -2278 254 -2278 0 1
rlabel polysilicon 254 -2284 254 -2284 0 3
rlabel polysilicon 261 -2278 261 -2278 0 1
rlabel polysilicon 261 -2284 261 -2284 0 3
rlabel polysilicon 268 -2278 268 -2278 0 1
rlabel polysilicon 268 -2284 268 -2284 0 3
rlabel polysilicon 275 -2278 275 -2278 0 1
rlabel polysilicon 275 -2284 275 -2284 0 3
rlabel polysilicon 282 -2278 282 -2278 0 1
rlabel polysilicon 282 -2284 282 -2284 0 3
rlabel polysilicon 292 -2278 292 -2278 0 2
rlabel polysilicon 289 -2284 289 -2284 0 3
rlabel polysilicon 292 -2284 292 -2284 0 4
rlabel polysilicon 296 -2278 296 -2278 0 1
rlabel polysilicon 296 -2284 296 -2284 0 3
rlabel polysilicon 303 -2278 303 -2278 0 1
rlabel polysilicon 303 -2284 303 -2284 0 3
rlabel polysilicon 310 -2278 310 -2278 0 1
rlabel polysilicon 310 -2284 310 -2284 0 3
rlabel polysilicon 317 -2278 317 -2278 0 1
rlabel polysilicon 317 -2284 317 -2284 0 3
rlabel polysilicon 324 -2278 324 -2278 0 1
rlabel polysilicon 327 -2278 327 -2278 0 2
rlabel polysilicon 331 -2278 331 -2278 0 1
rlabel polysilicon 331 -2284 331 -2284 0 3
rlabel polysilicon 338 -2278 338 -2278 0 1
rlabel polysilicon 338 -2284 338 -2284 0 3
rlabel polysilicon 348 -2278 348 -2278 0 2
rlabel polysilicon 348 -2284 348 -2284 0 4
rlabel polysilicon 352 -2278 352 -2278 0 1
rlabel polysilicon 355 -2278 355 -2278 0 2
rlabel polysilicon 352 -2284 352 -2284 0 3
rlabel polysilicon 355 -2284 355 -2284 0 4
rlabel polysilicon 359 -2278 359 -2278 0 1
rlabel polysilicon 359 -2284 359 -2284 0 3
rlabel polysilicon 369 -2278 369 -2278 0 2
rlabel polysilicon 366 -2284 366 -2284 0 3
rlabel polysilicon 373 -2278 373 -2278 0 1
rlabel polysilicon 373 -2284 373 -2284 0 3
rlabel polysilicon 380 -2278 380 -2278 0 1
rlabel polysilicon 383 -2278 383 -2278 0 2
rlabel polysilicon 380 -2284 380 -2284 0 3
rlabel polysilicon 383 -2284 383 -2284 0 4
rlabel polysilicon 387 -2278 387 -2278 0 1
rlabel polysilicon 387 -2284 387 -2284 0 3
rlabel polysilicon 394 -2278 394 -2278 0 1
rlabel polysilicon 394 -2284 394 -2284 0 3
rlabel polysilicon 401 -2278 401 -2278 0 1
rlabel polysilicon 401 -2284 401 -2284 0 3
rlabel polysilicon 408 -2278 408 -2278 0 1
rlabel polysilicon 408 -2284 408 -2284 0 3
rlabel polysilicon 415 -2278 415 -2278 0 1
rlabel polysilicon 415 -2284 415 -2284 0 3
rlabel polysilicon 422 -2278 422 -2278 0 1
rlabel polysilicon 422 -2284 422 -2284 0 3
rlabel polysilicon 429 -2278 429 -2278 0 1
rlabel polysilicon 429 -2284 429 -2284 0 3
rlabel polysilicon 436 -2278 436 -2278 0 1
rlabel polysilicon 436 -2284 436 -2284 0 3
rlabel polysilicon 443 -2278 443 -2278 0 1
rlabel polysilicon 443 -2284 443 -2284 0 3
rlabel polysilicon 450 -2278 450 -2278 0 1
rlabel polysilicon 450 -2284 450 -2284 0 3
rlabel polysilicon 457 -2278 457 -2278 0 1
rlabel polysilicon 457 -2284 457 -2284 0 3
rlabel polysilicon 464 -2278 464 -2278 0 1
rlabel polysilicon 467 -2278 467 -2278 0 2
rlabel polysilicon 464 -2284 464 -2284 0 3
rlabel polysilicon 467 -2284 467 -2284 0 4
rlabel polysilicon 471 -2278 471 -2278 0 1
rlabel polysilicon 471 -2284 471 -2284 0 3
rlabel polysilicon 478 -2278 478 -2278 0 1
rlabel polysilicon 481 -2278 481 -2278 0 2
rlabel polysilicon 481 -2284 481 -2284 0 4
rlabel polysilicon 485 -2278 485 -2278 0 1
rlabel polysilicon 488 -2278 488 -2278 0 2
rlabel polysilicon 485 -2284 485 -2284 0 3
rlabel polysilicon 488 -2284 488 -2284 0 4
rlabel polysilicon 492 -2278 492 -2278 0 1
rlabel polysilicon 492 -2284 492 -2284 0 3
rlabel polysilicon 499 -2278 499 -2278 0 1
rlabel polysilicon 502 -2278 502 -2278 0 2
rlabel polysilicon 502 -2284 502 -2284 0 4
rlabel polysilicon 506 -2278 506 -2278 0 1
rlabel polysilicon 506 -2284 506 -2284 0 3
rlabel polysilicon 513 -2278 513 -2278 0 1
rlabel polysilicon 513 -2284 513 -2284 0 3
rlabel polysilicon 520 -2278 520 -2278 0 1
rlabel polysilicon 520 -2284 520 -2284 0 3
rlabel polysilicon 527 -2278 527 -2278 0 1
rlabel polysilicon 527 -2284 527 -2284 0 3
rlabel polysilicon 534 -2278 534 -2278 0 1
rlabel polysilicon 534 -2284 534 -2284 0 3
rlabel polysilicon 541 -2278 541 -2278 0 1
rlabel polysilicon 544 -2278 544 -2278 0 2
rlabel polysilicon 541 -2284 541 -2284 0 3
rlabel polysilicon 544 -2284 544 -2284 0 4
rlabel polysilicon 548 -2278 548 -2278 0 1
rlabel polysilicon 548 -2284 548 -2284 0 3
rlabel polysilicon 555 -2278 555 -2278 0 1
rlabel polysilicon 555 -2284 555 -2284 0 3
rlabel polysilicon 562 -2278 562 -2278 0 1
rlabel polysilicon 562 -2284 562 -2284 0 3
rlabel polysilicon 569 -2278 569 -2278 0 1
rlabel polysilicon 569 -2284 569 -2284 0 3
rlabel polysilicon 576 -2278 576 -2278 0 1
rlabel polysilicon 579 -2278 579 -2278 0 2
rlabel polysilicon 576 -2284 576 -2284 0 3
rlabel polysilicon 579 -2284 579 -2284 0 4
rlabel polysilicon 583 -2278 583 -2278 0 1
rlabel polysilicon 583 -2284 583 -2284 0 3
rlabel polysilicon 590 -2278 590 -2278 0 1
rlabel polysilicon 590 -2284 590 -2284 0 3
rlabel polysilicon 597 -2278 597 -2278 0 1
rlabel polysilicon 597 -2284 597 -2284 0 3
rlabel polysilicon 604 -2278 604 -2278 0 1
rlabel polysilicon 604 -2284 604 -2284 0 3
rlabel polysilicon 611 -2278 611 -2278 0 1
rlabel polysilicon 611 -2284 611 -2284 0 3
rlabel polysilicon 618 -2278 618 -2278 0 1
rlabel polysilicon 618 -2284 618 -2284 0 3
rlabel polysilicon 625 -2278 625 -2278 0 1
rlabel polysilicon 625 -2284 625 -2284 0 3
rlabel polysilicon 632 -2278 632 -2278 0 1
rlabel polysilicon 632 -2284 632 -2284 0 3
rlabel polysilicon 639 -2278 639 -2278 0 1
rlabel polysilicon 639 -2284 639 -2284 0 3
rlabel polysilicon 646 -2278 646 -2278 0 1
rlabel polysilicon 646 -2284 646 -2284 0 3
rlabel polysilicon 653 -2278 653 -2278 0 1
rlabel polysilicon 653 -2284 653 -2284 0 3
rlabel polysilicon 660 -2278 660 -2278 0 1
rlabel polysilicon 660 -2284 660 -2284 0 3
rlabel polysilicon 667 -2278 667 -2278 0 1
rlabel polysilicon 667 -2284 667 -2284 0 3
rlabel polysilicon 674 -2278 674 -2278 0 1
rlabel polysilicon 674 -2284 674 -2284 0 3
rlabel polysilicon 681 -2278 681 -2278 0 1
rlabel polysilicon 684 -2278 684 -2278 0 2
rlabel polysilicon 681 -2284 681 -2284 0 3
rlabel polysilicon 684 -2284 684 -2284 0 4
rlabel polysilicon 688 -2278 688 -2278 0 1
rlabel polysilicon 688 -2284 688 -2284 0 3
rlabel polysilicon 695 -2278 695 -2278 0 1
rlabel polysilicon 695 -2284 695 -2284 0 3
rlabel polysilicon 702 -2278 702 -2278 0 1
rlabel polysilicon 702 -2284 702 -2284 0 3
rlabel polysilicon 709 -2278 709 -2278 0 1
rlabel polysilicon 709 -2284 709 -2284 0 3
rlabel polysilicon 716 -2278 716 -2278 0 1
rlabel polysilicon 716 -2284 716 -2284 0 3
rlabel polysilicon 723 -2278 723 -2278 0 1
rlabel polysilicon 723 -2284 723 -2284 0 3
rlabel polysilicon 730 -2278 730 -2278 0 1
rlabel polysilicon 730 -2284 730 -2284 0 3
rlabel polysilicon 737 -2278 737 -2278 0 1
rlabel polysilicon 737 -2284 737 -2284 0 3
rlabel polysilicon 744 -2278 744 -2278 0 1
rlabel polysilicon 744 -2284 744 -2284 0 3
rlabel polysilicon 751 -2278 751 -2278 0 1
rlabel polysilicon 751 -2284 751 -2284 0 3
rlabel polysilicon 758 -2278 758 -2278 0 1
rlabel polysilicon 758 -2284 758 -2284 0 3
rlabel polysilicon 768 -2278 768 -2278 0 2
rlabel polysilicon 768 -2284 768 -2284 0 4
rlabel polysilicon 772 -2278 772 -2278 0 1
rlabel polysilicon 772 -2284 772 -2284 0 3
rlabel polysilicon 779 -2278 779 -2278 0 1
rlabel polysilicon 779 -2284 779 -2284 0 3
rlabel polysilicon 786 -2278 786 -2278 0 1
rlabel polysilicon 786 -2284 786 -2284 0 3
rlabel polysilicon 793 -2278 793 -2278 0 1
rlabel polysilicon 793 -2284 793 -2284 0 3
rlabel polysilicon 800 -2278 800 -2278 0 1
rlabel polysilicon 800 -2284 800 -2284 0 3
rlabel polysilicon 807 -2278 807 -2278 0 1
rlabel polysilicon 807 -2284 807 -2284 0 3
rlabel polysilicon 814 -2278 814 -2278 0 1
rlabel polysilicon 814 -2284 814 -2284 0 3
rlabel polysilicon 821 -2278 821 -2278 0 1
rlabel polysilicon 821 -2284 821 -2284 0 3
rlabel polysilicon 828 -2278 828 -2278 0 1
rlabel polysilicon 828 -2284 828 -2284 0 3
rlabel polysilicon 835 -2278 835 -2278 0 1
rlabel polysilicon 835 -2284 835 -2284 0 3
rlabel polysilicon 842 -2278 842 -2278 0 1
rlabel polysilicon 842 -2284 842 -2284 0 3
rlabel polysilicon 849 -2278 849 -2278 0 1
rlabel polysilicon 849 -2284 849 -2284 0 3
rlabel polysilicon 856 -2278 856 -2278 0 1
rlabel polysilicon 856 -2284 856 -2284 0 3
rlabel polysilicon 863 -2278 863 -2278 0 1
rlabel polysilicon 863 -2284 863 -2284 0 3
rlabel polysilicon 870 -2278 870 -2278 0 1
rlabel polysilicon 870 -2284 870 -2284 0 3
rlabel polysilicon 877 -2278 877 -2278 0 1
rlabel polysilicon 877 -2284 877 -2284 0 3
rlabel polysilicon 884 -2278 884 -2278 0 1
rlabel polysilicon 884 -2284 884 -2284 0 3
rlabel polysilicon 891 -2278 891 -2278 0 1
rlabel polysilicon 891 -2284 891 -2284 0 3
rlabel polysilicon 898 -2278 898 -2278 0 1
rlabel polysilicon 898 -2284 898 -2284 0 3
rlabel polysilicon 901 -2284 901 -2284 0 4
rlabel polysilicon 905 -2284 905 -2284 0 3
rlabel polysilicon 908 -2284 908 -2284 0 4
rlabel polysilicon 912 -2278 912 -2278 0 1
rlabel polysilicon 912 -2284 912 -2284 0 3
rlabel polysilicon 922 -2278 922 -2278 0 2
rlabel polysilicon 922 -2284 922 -2284 0 4
rlabel polysilicon 929 -2278 929 -2278 0 2
rlabel polysilicon 926 -2284 926 -2284 0 3
rlabel polysilicon 933 -2278 933 -2278 0 1
rlabel polysilicon 933 -2284 933 -2284 0 3
rlabel polysilicon 940 -2278 940 -2278 0 1
rlabel polysilicon 940 -2284 940 -2284 0 3
rlabel polysilicon 947 -2278 947 -2278 0 1
rlabel polysilicon 947 -2284 947 -2284 0 3
rlabel polysilicon 954 -2278 954 -2278 0 1
rlabel polysilicon 954 -2284 954 -2284 0 3
rlabel polysilicon 961 -2278 961 -2278 0 1
rlabel polysilicon 961 -2284 961 -2284 0 3
rlabel polysilicon 968 -2278 968 -2278 0 1
rlabel polysilicon 975 -2278 975 -2278 0 1
rlabel polysilicon 975 -2284 975 -2284 0 3
rlabel polysilicon 2 -2365 2 -2365 0 1
rlabel polysilicon 2 -2371 2 -2371 0 3
rlabel polysilicon 12 -2365 12 -2365 0 2
rlabel polysilicon 16 -2365 16 -2365 0 1
rlabel polysilicon 16 -2371 16 -2371 0 3
rlabel polysilicon 23 -2365 23 -2365 0 1
rlabel polysilicon 23 -2371 23 -2371 0 3
rlabel polysilicon 30 -2365 30 -2365 0 1
rlabel polysilicon 30 -2371 30 -2371 0 3
rlabel polysilicon 37 -2365 37 -2365 0 1
rlabel polysilicon 37 -2371 37 -2371 0 3
rlabel polysilicon 44 -2365 44 -2365 0 1
rlabel polysilicon 47 -2365 47 -2365 0 2
rlabel polysilicon 44 -2371 44 -2371 0 3
rlabel polysilicon 51 -2365 51 -2365 0 1
rlabel polysilicon 54 -2365 54 -2365 0 2
rlabel polysilicon 51 -2371 51 -2371 0 3
rlabel polysilicon 58 -2365 58 -2365 0 1
rlabel polysilicon 58 -2371 58 -2371 0 3
rlabel polysilicon 65 -2365 65 -2365 0 1
rlabel polysilicon 65 -2371 65 -2371 0 3
rlabel polysilicon 72 -2365 72 -2365 0 1
rlabel polysilicon 72 -2371 72 -2371 0 3
rlabel polysilicon 79 -2365 79 -2365 0 1
rlabel polysilicon 79 -2371 79 -2371 0 3
rlabel polysilicon 86 -2365 86 -2365 0 1
rlabel polysilicon 86 -2371 86 -2371 0 3
rlabel polysilicon 93 -2365 93 -2365 0 1
rlabel polysilicon 93 -2371 93 -2371 0 3
rlabel polysilicon 100 -2365 100 -2365 0 1
rlabel polysilicon 100 -2371 100 -2371 0 3
rlabel polysilicon 107 -2365 107 -2365 0 1
rlabel polysilicon 110 -2365 110 -2365 0 2
rlabel polysilicon 107 -2371 107 -2371 0 3
rlabel polysilicon 114 -2365 114 -2365 0 1
rlabel polysilicon 114 -2371 114 -2371 0 3
rlabel polysilicon 121 -2365 121 -2365 0 1
rlabel polysilicon 121 -2371 121 -2371 0 3
rlabel polysilicon 128 -2365 128 -2365 0 1
rlabel polysilicon 128 -2371 128 -2371 0 3
rlabel polysilicon 135 -2365 135 -2365 0 1
rlabel polysilicon 135 -2371 135 -2371 0 3
rlabel polysilicon 142 -2365 142 -2365 0 1
rlabel polysilicon 142 -2371 142 -2371 0 3
rlabel polysilicon 149 -2365 149 -2365 0 1
rlabel polysilicon 149 -2371 149 -2371 0 3
rlabel polysilicon 156 -2365 156 -2365 0 1
rlabel polysilicon 159 -2365 159 -2365 0 2
rlabel polysilicon 156 -2371 156 -2371 0 3
rlabel polysilicon 163 -2365 163 -2365 0 1
rlabel polysilicon 163 -2371 163 -2371 0 3
rlabel polysilicon 170 -2365 170 -2365 0 1
rlabel polysilicon 170 -2371 170 -2371 0 3
rlabel polysilicon 177 -2365 177 -2365 0 1
rlabel polysilicon 177 -2371 177 -2371 0 3
rlabel polysilicon 184 -2365 184 -2365 0 1
rlabel polysilicon 184 -2371 184 -2371 0 3
rlabel polysilicon 191 -2365 191 -2365 0 1
rlabel polysilicon 191 -2371 191 -2371 0 3
rlabel polysilicon 198 -2365 198 -2365 0 1
rlabel polysilicon 198 -2371 198 -2371 0 3
rlabel polysilicon 205 -2365 205 -2365 0 1
rlabel polysilicon 205 -2371 205 -2371 0 3
rlabel polysilicon 212 -2365 212 -2365 0 1
rlabel polysilicon 212 -2371 212 -2371 0 3
rlabel polysilicon 219 -2371 219 -2371 0 3
rlabel polysilicon 222 -2371 222 -2371 0 4
rlabel polysilicon 229 -2365 229 -2365 0 2
rlabel polysilicon 226 -2371 226 -2371 0 3
rlabel polysilicon 233 -2365 233 -2365 0 1
rlabel polysilicon 233 -2371 233 -2371 0 3
rlabel polysilicon 240 -2365 240 -2365 0 1
rlabel polysilicon 240 -2371 240 -2371 0 3
rlabel polysilicon 247 -2365 247 -2365 0 1
rlabel polysilicon 247 -2371 247 -2371 0 3
rlabel polysilicon 254 -2365 254 -2365 0 1
rlabel polysilicon 254 -2371 254 -2371 0 3
rlabel polysilicon 261 -2365 261 -2365 0 1
rlabel polysilicon 261 -2371 261 -2371 0 3
rlabel polysilicon 268 -2365 268 -2365 0 1
rlabel polysilicon 271 -2371 271 -2371 0 4
rlabel polysilicon 275 -2365 275 -2365 0 1
rlabel polysilicon 275 -2371 275 -2371 0 3
rlabel polysilicon 282 -2365 282 -2365 0 1
rlabel polysilicon 282 -2371 282 -2371 0 3
rlabel polysilicon 289 -2365 289 -2365 0 1
rlabel polysilicon 289 -2371 289 -2371 0 3
rlabel polysilicon 296 -2365 296 -2365 0 1
rlabel polysilicon 296 -2371 296 -2371 0 3
rlabel polysilicon 303 -2365 303 -2365 0 1
rlabel polysilicon 303 -2371 303 -2371 0 3
rlabel polysilicon 310 -2365 310 -2365 0 1
rlabel polysilicon 313 -2365 313 -2365 0 2
rlabel polysilicon 310 -2371 310 -2371 0 3
rlabel polysilicon 313 -2371 313 -2371 0 4
rlabel polysilicon 317 -2365 317 -2365 0 1
rlabel polysilicon 317 -2371 317 -2371 0 3
rlabel polysilicon 324 -2365 324 -2365 0 1
rlabel polysilicon 324 -2371 324 -2371 0 3
rlabel polysilicon 334 -2365 334 -2365 0 2
rlabel polysilicon 331 -2371 331 -2371 0 3
rlabel polysilicon 334 -2371 334 -2371 0 4
rlabel polysilicon 338 -2365 338 -2365 0 1
rlabel polysilicon 341 -2365 341 -2365 0 2
rlabel polysilicon 341 -2371 341 -2371 0 4
rlabel polysilicon 345 -2365 345 -2365 0 1
rlabel polysilicon 345 -2371 345 -2371 0 3
rlabel polysilicon 355 -2365 355 -2365 0 2
rlabel polysilicon 355 -2371 355 -2371 0 4
rlabel polysilicon 359 -2365 359 -2365 0 1
rlabel polysilicon 362 -2365 362 -2365 0 2
rlabel polysilicon 366 -2365 366 -2365 0 1
rlabel polysilicon 366 -2371 366 -2371 0 3
rlabel polysilicon 373 -2365 373 -2365 0 1
rlabel polysilicon 376 -2365 376 -2365 0 2
rlabel polysilicon 380 -2365 380 -2365 0 1
rlabel polysilicon 380 -2371 380 -2371 0 3
rlabel polysilicon 387 -2365 387 -2365 0 1
rlabel polysilicon 387 -2371 387 -2371 0 3
rlabel polysilicon 394 -2365 394 -2365 0 1
rlabel polysilicon 397 -2365 397 -2365 0 2
rlabel polysilicon 401 -2365 401 -2365 0 1
rlabel polysilicon 401 -2371 401 -2371 0 3
rlabel polysilicon 404 -2371 404 -2371 0 4
rlabel polysilicon 408 -2365 408 -2365 0 1
rlabel polysilicon 408 -2371 408 -2371 0 3
rlabel polysilicon 415 -2365 415 -2365 0 1
rlabel polysilicon 415 -2371 415 -2371 0 3
rlabel polysilicon 418 -2371 418 -2371 0 4
rlabel polysilicon 422 -2365 422 -2365 0 1
rlabel polysilicon 422 -2371 422 -2371 0 3
rlabel polysilicon 429 -2365 429 -2365 0 1
rlabel polysilicon 429 -2371 429 -2371 0 3
rlabel polysilicon 436 -2365 436 -2365 0 1
rlabel polysilicon 436 -2371 436 -2371 0 3
rlabel polysilicon 443 -2365 443 -2365 0 1
rlabel polysilicon 443 -2371 443 -2371 0 3
rlabel polysilicon 450 -2365 450 -2365 0 1
rlabel polysilicon 450 -2371 450 -2371 0 3
rlabel polysilicon 457 -2371 457 -2371 0 3
rlabel polysilicon 464 -2365 464 -2365 0 1
rlabel polysilicon 467 -2365 467 -2365 0 2
rlabel polysilicon 464 -2371 464 -2371 0 3
rlabel polysilicon 471 -2365 471 -2365 0 1
rlabel polysilicon 471 -2371 471 -2371 0 3
rlabel polysilicon 478 -2365 478 -2365 0 1
rlabel polysilicon 485 -2365 485 -2365 0 1
rlabel polysilicon 485 -2371 485 -2371 0 3
rlabel polysilicon 492 -2365 492 -2365 0 1
rlabel polysilicon 492 -2371 492 -2371 0 3
rlabel polysilicon 499 -2365 499 -2365 0 1
rlabel polysilicon 499 -2371 499 -2371 0 3
rlabel polysilicon 506 -2365 506 -2365 0 1
rlabel polysilicon 506 -2371 506 -2371 0 3
rlabel polysilicon 513 -2365 513 -2365 0 1
rlabel polysilicon 513 -2371 513 -2371 0 3
rlabel polysilicon 523 -2365 523 -2365 0 2
rlabel polysilicon 523 -2371 523 -2371 0 4
rlabel polysilicon 527 -2365 527 -2365 0 1
rlabel polysilicon 527 -2371 527 -2371 0 3
rlabel polysilicon 537 -2365 537 -2365 0 2
rlabel polysilicon 534 -2371 534 -2371 0 3
rlabel polysilicon 541 -2365 541 -2365 0 1
rlabel polysilicon 541 -2371 541 -2371 0 3
rlabel polysilicon 548 -2365 548 -2365 0 1
rlabel polysilicon 548 -2371 548 -2371 0 3
rlabel polysilicon 555 -2365 555 -2365 0 1
rlabel polysilicon 558 -2371 558 -2371 0 4
rlabel polysilicon 562 -2365 562 -2365 0 1
rlabel polysilicon 565 -2365 565 -2365 0 2
rlabel polysilicon 565 -2371 565 -2371 0 4
rlabel polysilicon 569 -2365 569 -2365 0 1
rlabel polysilicon 569 -2371 569 -2371 0 3
rlabel polysilicon 576 -2365 576 -2365 0 1
rlabel polysilicon 576 -2371 576 -2371 0 3
rlabel polysilicon 583 -2365 583 -2365 0 1
rlabel polysilicon 586 -2365 586 -2365 0 2
rlabel polysilicon 590 -2365 590 -2365 0 1
rlabel polysilicon 590 -2371 590 -2371 0 3
rlabel polysilicon 597 -2365 597 -2365 0 1
rlabel polysilicon 597 -2371 597 -2371 0 3
rlabel polysilicon 604 -2365 604 -2365 0 1
rlabel polysilicon 604 -2371 604 -2371 0 3
rlabel polysilicon 611 -2365 611 -2365 0 1
rlabel polysilicon 611 -2371 611 -2371 0 3
rlabel polysilicon 618 -2365 618 -2365 0 1
rlabel polysilicon 618 -2371 618 -2371 0 3
rlabel polysilicon 625 -2365 625 -2365 0 1
rlabel polysilicon 625 -2371 625 -2371 0 3
rlabel polysilicon 632 -2365 632 -2365 0 1
rlabel polysilicon 632 -2371 632 -2371 0 3
rlabel polysilicon 639 -2365 639 -2365 0 1
rlabel polysilicon 642 -2365 642 -2365 0 2
rlabel polysilicon 639 -2371 639 -2371 0 3
rlabel polysilicon 646 -2365 646 -2365 0 1
rlabel polysilicon 646 -2371 646 -2371 0 3
rlabel polysilicon 653 -2365 653 -2365 0 1
rlabel polysilicon 653 -2371 653 -2371 0 3
rlabel polysilicon 660 -2365 660 -2365 0 1
rlabel polysilicon 660 -2371 660 -2371 0 3
rlabel polysilicon 667 -2365 667 -2365 0 1
rlabel polysilicon 667 -2371 667 -2371 0 3
rlabel polysilicon 674 -2365 674 -2365 0 1
rlabel polysilicon 674 -2371 674 -2371 0 3
rlabel polysilicon 681 -2365 681 -2365 0 1
rlabel polysilicon 681 -2371 681 -2371 0 3
rlabel polysilicon 688 -2365 688 -2365 0 1
rlabel polysilicon 688 -2371 688 -2371 0 3
rlabel polysilicon 695 -2365 695 -2365 0 1
rlabel polysilicon 695 -2371 695 -2371 0 3
rlabel polysilicon 702 -2365 702 -2365 0 1
rlabel polysilicon 705 -2365 705 -2365 0 2
rlabel polysilicon 709 -2365 709 -2365 0 1
rlabel polysilicon 709 -2371 709 -2371 0 3
rlabel polysilicon 716 -2365 716 -2365 0 1
rlabel polysilicon 716 -2371 716 -2371 0 3
rlabel polysilicon 723 -2365 723 -2365 0 1
rlabel polysilicon 723 -2371 723 -2371 0 3
rlabel polysilicon 730 -2365 730 -2365 0 1
rlabel polysilicon 730 -2371 730 -2371 0 3
rlabel polysilicon 737 -2365 737 -2365 0 1
rlabel polysilicon 737 -2371 737 -2371 0 3
rlabel polysilicon 744 -2365 744 -2365 0 1
rlabel polysilicon 744 -2371 744 -2371 0 3
rlabel polysilicon 751 -2365 751 -2365 0 1
rlabel polysilicon 751 -2371 751 -2371 0 3
rlabel polysilicon 758 -2365 758 -2365 0 1
rlabel polysilicon 758 -2371 758 -2371 0 3
rlabel polysilicon 765 -2365 765 -2365 0 1
rlabel polysilicon 765 -2371 765 -2371 0 3
rlabel polysilicon 772 -2365 772 -2365 0 1
rlabel polysilicon 772 -2371 772 -2371 0 3
rlabel polysilicon 779 -2365 779 -2365 0 1
rlabel polysilicon 779 -2371 779 -2371 0 3
rlabel polysilicon 786 -2365 786 -2365 0 1
rlabel polysilicon 786 -2371 786 -2371 0 3
rlabel polysilicon 793 -2365 793 -2365 0 1
rlabel polysilicon 793 -2371 793 -2371 0 3
rlabel polysilicon 800 -2365 800 -2365 0 1
rlabel polysilicon 807 -2365 807 -2365 0 1
rlabel polysilicon 807 -2371 807 -2371 0 3
rlabel polysilicon 814 -2365 814 -2365 0 1
rlabel polysilicon 814 -2371 814 -2371 0 3
rlabel polysilicon 821 -2365 821 -2365 0 1
rlabel polysilicon 821 -2371 821 -2371 0 3
rlabel polysilicon 828 -2365 828 -2365 0 1
rlabel polysilicon 828 -2371 828 -2371 0 3
rlabel polysilicon 835 -2365 835 -2365 0 1
rlabel polysilicon 835 -2371 835 -2371 0 3
rlabel polysilicon 842 -2365 842 -2365 0 1
rlabel polysilicon 842 -2371 842 -2371 0 3
rlabel polysilicon 849 -2365 849 -2365 0 1
rlabel polysilicon 849 -2371 849 -2371 0 3
rlabel polysilicon 856 -2365 856 -2365 0 1
rlabel polysilicon 856 -2371 856 -2371 0 3
rlabel polysilicon 863 -2365 863 -2365 0 1
rlabel polysilicon 863 -2371 863 -2371 0 3
rlabel polysilicon 870 -2365 870 -2365 0 1
rlabel polysilicon 877 -2365 877 -2365 0 1
rlabel polysilicon 877 -2371 877 -2371 0 3
rlabel polysilicon 884 -2365 884 -2365 0 1
rlabel polysilicon 884 -2371 884 -2371 0 3
rlabel polysilicon 891 -2365 891 -2365 0 1
rlabel polysilicon 891 -2371 891 -2371 0 3
rlabel polysilicon 929 -2365 929 -2365 0 2
rlabel polysilicon 926 -2371 926 -2371 0 3
rlabel polysilicon 947 -2365 947 -2365 0 1
rlabel polysilicon 947 -2371 947 -2371 0 3
rlabel polysilicon 30 -2430 30 -2430 0 1
rlabel polysilicon 58 -2430 58 -2430 0 1
rlabel polysilicon 61 -2430 61 -2430 0 2
rlabel polysilicon 65 -2430 65 -2430 0 1
rlabel polysilicon 65 -2436 65 -2436 0 3
rlabel polysilicon 72 -2430 72 -2430 0 1
rlabel polysilicon 79 -2430 79 -2430 0 1
rlabel polysilicon 79 -2436 79 -2436 0 3
rlabel polysilicon 86 -2430 86 -2430 0 1
rlabel polysilicon 86 -2436 86 -2436 0 3
rlabel polysilicon 93 -2430 93 -2430 0 1
rlabel polysilicon 93 -2436 93 -2436 0 3
rlabel polysilicon 100 -2430 100 -2430 0 1
rlabel polysilicon 100 -2436 100 -2436 0 3
rlabel polysilicon 107 -2430 107 -2430 0 1
rlabel polysilicon 107 -2436 107 -2436 0 3
rlabel polysilicon 114 -2430 114 -2430 0 1
rlabel polysilicon 114 -2436 114 -2436 0 3
rlabel polysilicon 121 -2430 121 -2430 0 1
rlabel polysilicon 121 -2436 121 -2436 0 3
rlabel polysilicon 128 -2430 128 -2430 0 1
rlabel polysilicon 128 -2436 128 -2436 0 3
rlabel polysilicon 138 -2430 138 -2430 0 2
rlabel polysilicon 142 -2430 142 -2430 0 1
rlabel polysilicon 142 -2436 142 -2436 0 3
rlabel polysilicon 149 -2430 149 -2430 0 1
rlabel polysilicon 152 -2430 152 -2430 0 2
rlabel polysilicon 149 -2436 149 -2436 0 3
rlabel polysilicon 152 -2436 152 -2436 0 4
rlabel polysilicon 156 -2430 156 -2430 0 1
rlabel polysilicon 156 -2436 156 -2436 0 3
rlabel polysilicon 159 -2436 159 -2436 0 4
rlabel polysilicon 163 -2430 163 -2430 0 1
rlabel polysilicon 163 -2436 163 -2436 0 3
rlabel polysilicon 170 -2430 170 -2430 0 1
rlabel polysilicon 170 -2436 170 -2436 0 3
rlabel polysilicon 177 -2430 177 -2430 0 1
rlabel polysilicon 177 -2436 177 -2436 0 3
rlabel polysilicon 184 -2430 184 -2430 0 1
rlabel polysilicon 184 -2436 184 -2436 0 3
rlabel polysilicon 191 -2430 191 -2430 0 1
rlabel polysilicon 191 -2436 191 -2436 0 3
rlabel polysilicon 198 -2430 198 -2430 0 1
rlabel polysilicon 198 -2436 198 -2436 0 3
rlabel polysilicon 208 -2430 208 -2430 0 2
rlabel polysilicon 208 -2436 208 -2436 0 4
rlabel polysilicon 215 -2430 215 -2430 0 2
rlabel polysilicon 212 -2436 212 -2436 0 3
rlabel polysilicon 215 -2436 215 -2436 0 4
rlabel polysilicon 219 -2430 219 -2430 0 1
rlabel polysilicon 222 -2430 222 -2430 0 2
rlabel polysilicon 219 -2436 219 -2436 0 3
rlabel polysilicon 222 -2436 222 -2436 0 4
rlabel polysilicon 226 -2430 226 -2430 0 1
rlabel polysilicon 226 -2436 226 -2436 0 3
rlabel polysilicon 233 -2430 233 -2430 0 1
rlabel polysilicon 233 -2436 233 -2436 0 3
rlabel polysilicon 240 -2430 240 -2430 0 1
rlabel polysilicon 240 -2436 240 -2436 0 3
rlabel polysilicon 247 -2430 247 -2430 0 1
rlabel polysilicon 247 -2436 247 -2436 0 3
rlabel polysilicon 254 -2430 254 -2430 0 1
rlabel polysilicon 254 -2436 254 -2436 0 3
rlabel polysilicon 261 -2430 261 -2430 0 1
rlabel polysilicon 261 -2436 261 -2436 0 3
rlabel polysilicon 268 -2430 268 -2430 0 1
rlabel polysilicon 268 -2436 268 -2436 0 3
rlabel polysilicon 275 -2430 275 -2430 0 1
rlabel polysilicon 275 -2436 275 -2436 0 3
rlabel polysilicon 282 -2430 282 -2430 0 1
rlabel polysilicon 282 -2436 282 -2436 0 3
rlabel polysilicon 289 -2430 289 -2430 0 1
rlabel polysilicon 289 -2436 289 -2436 0 3
rlabel polysilicon 296 -2430 296 -2430 0 1
rlabel polysilicon 296 -2436 296 -2436 0 3
rlabel polysilicon 303 -2430 303 -2430 0 1
rlabel polysilicon 303 -2436 303 -2436 0 3
rlabel polysilicon 310 -2430 310 -2430 0 1
rlabel polysilicon 310 -2436 310 -2436 0 3
rlabel polysilicon 317 -2430 317 -2430 0 1
rlabel polysilicon 317 -2436 317 -2436 0 3
rlabel polysilicon 324 -2430 324 -2430 0 1
rlabel polysilicon 324 -2436 324 -2436 0 3
rlabel polysilicon 331 -2430 331 -2430 0 1
rlabel polysilicon 334 -2430 334 -2430 0 2
rlabel polysilicon 331 -2436 331 -2436 0 3
rlabel polysilicon 334 -2436 334 -2436 0 4
rlabel polysilicon 338 -2430 338 -2430 0 1
rlabel polysilicon 338 -2436 338 -2436 0 3
rlabel polysilicon 345 -2430 345 -2430 0 1
rlabel polysilicon 345 -2436 345 -2436 0 3
rlabel polysilicon 352 -2430 352 -2430 0 1
rlabel polysilicon 352 -2436 352 -2436 0 3
rlabel polysilicon 359 -2430 359 -2430 0 1
rlabel polysilicon 359 -2436 359 -2436 0 3
rlabel polysilicon 366 -2430 366 -2430 0 1
rlabel polysilicon 366 -2436 366 -2436 0 3
rlabel polysilicon 373 -2430 373 -2430 0 1
rlabel polysilicon 376 -2430 376 -2430 0 2
rlabel polysilicon 380 -2430 380 -2430 0 1
rlabel polysilicon 380 -2436 380 -2436 0 3
rlabel polysilicon 387 -2430 387 -2430 0 1
rlabel polysilicon 387 -2436 387 -2436 0 3
rlabel polysilicon 394 -2430 394 -2430 0 1
rlabel polysilicon 397 -2430 397 -2430 0 2
rlabel polysilicon 394 -2436 394 -2436 0 3
rlabel polysilicon 397 -2436 397 -2436 0 4
rlabel polysilicon 401 -2430 401 -2430 0 1
rlabel polysilicon 401 -2436 401 -2436 0 3
rlabel polysilicon 408 -2430 408 -2430 0 1
rlabel polysilicon 411 -2430 411 -2430 0 2
rlabel polysilicon 408 -2436 408 -2436 0 3
rlabel polysilicon 415 -2430 415 -2430 0 1
rlabel polysilicon 415 -2436 415 -2436 0 3
rlabel polysilicon 422 -2430 422 -2430 0 1
rlabel polysilicon 422 -2436 422 -2436 0 3
rlabel polysilicon 429 -2430 429 -2430 0 1
rlabel polysilicon 432 -2436 432 -2436 0 4
rlabel polysilicon 436 -2430 436 -2430 0 1
rlabel polysilicon 436 -2436 436 -2436 0 3
rlabel polysilicon 443 -2430 443 -2430 0 1
rlabel polysilicon 443 -2436 443 -2436 0 3
rlabel polysilicon 450 -2430 450 -2430 0 1
rlabel polysilicon 450 -2436 450 -2436 0 3
rlabel polysilicon 457 -2430 457 -2430 0 1
rlabel polysilicon 460 -2430 460 -2430 0 2
rlabel polysilicon 460 -2436 460 -2436 0 4
rlabel polysilicon 464 -2430 464 -2430 0 1
rlabel polysilicon 464 -2436 464 -2436 0 3
rlabel polysilicon 467 -2436 467 -2436 0 4
rlabel polysilicon 471 -2430 471 -2430 0 1
rlabel polysilicon 471 -2436 471 -2436 0 3
rlabel polysilicon 474 -2436 474 -2436 0 4
rlabel polysilicon 481 -2430 481 -2430 0 2
rlabel polysilicon 478 -2436 478 -2436 0 3
rlabel polysilicon 481 -2436 481 -2436 0 4
rlabel polysilicon 488 -2430 488 -2430 0 2
rlabel polysilicon 485 -2436 485 -2436 0 3
rlabel polysilicon 488 -2436 488 -2436 0 4
rlabel polysilicon 492 -2430 492 -2430 0 1
rlabel polysilicon 492 -2436 492 -2436 0 3
rlabel polysilicon 499 -2430 499 -2430 0 1
rlabel polysilicon 499 -2436 499 -2436 0 3
rlabel polysilicon 506 -2430 506 -2430 0 1
rlabel polysilicon 506 -2436 506 -2436 0 3
rlabel polysilicon 513 -2430 513 -2430 0 1
rlabel polysilicon 513 -2436 513 -2436 0 3
rlabel polysilicon 520 -2430 520 -2430 0 1
rlabel polysilicon 520 -2436 520 -2436 0 3
rlabel polysilicon 527 -2430 527 -2430 0 1
rlabel polysilicon 527 -2436 527 -2436 0 3
rlabel polysilicon 534 -2430 534 -2430 0 1
rlabel polysilicon 534 -2436 534 -2436 0 3
rlabel polysilicon 544 -2430 544 -2430 0 2
rlabel polysilicon 548 -2430 548 -2430 0 1
rlabel polysilicon 551 -2430 551 -2430 0 2
rlabel polysilicon 551 -2436 551 -2436 0 4
rlabel polysilicon 555 -2430 555 -2430 0 1
rlabel polysilicon 555 -2436 555 -2436 0 3
rlabel polysilicon 562 -2430 562 -2430 0 1
rlabel polysilicon 562 -2436 562 -2436 0 3
rlabel polysilicon 569 -2430 569 -2430 0 1
rlabel polysilicon 569 -2436 569 -2436 0 3
rlabel polysilicon 576 -2436 576 -2436 0 3
rlabel polysilicon 579 -2436 579 -2436 0 4
rlabel polysilicon 583 -2430 583 -2430 0 1
rlabel polysilicon 583 -2436 583 -2436 0 3
rlabel polysilicon 590 -2430 590 -2430 0 1
rlabel polysilicon 590 -2436 590 -2436 0 3
rlabel polysilicon 597 -2430 597 -2430 0 1
rlabel polysilicon 597 -2436 597 -2436 0 3
rlabel polysilicon 604 -2430 604 -2430 0 1
rlabel polysilicon 604 -2436 604 -2436 0 3
rlabel polysilicon 611 -2430 611 -2430 0 1
rlabel polysilicon 611 -2436 611 -2436 0 3
rlabel polysilicon 618 -2430 618 -2430 0 1
rlabel polysilicon 618 -2436 618 -2436 0 3
rlabel polysilicon 628 -2430 628 -2430 0 2
rlabel polysilicon 625 -2436 625 -2436 0 3
rlabel polysilicon 632 -2430 632 -2430 0 1
rlabel polysilicon 632 -2436 632 -2436 0 3
rlabel polysilicon 639 -2430 639 -2430 0 1
rlabel polysilicon 639 -2436 639 -2436 0 3
rlabel polysilicon 646 -2430 646 -2430 0 1
rlabel polysilicon 646 -2436 646 -2436 0 3
rlabel polysilicon 653 -2430 653 -2430 0 1
rlabel polysilicon 653 -2436 653 -2436 0 3
rlabel polysilicon 660 -2430 660 -2430 0 1
rlabel polysilicon 660 -2436 660 -2436 0 3
rlabel polysilicon 667 -2430 667 -2430 0 1
rlabel polysilicon 667 -2436 667 -2436 0 3
rlabel polysilicon 674 -2430 674 -2430 0 1
rlabel polysilicon 674 -2436 674 -2436 0 3
rlabel polysilicon 681 -2430 681 -2430 0 1
rlabel polysilicon 681 -2436 681 -2436 0 3
rlabel polysilicon 702 -2430 702 -2430 0 1
rlabel polysilicon 702 -2436 702 -2436 0 3
rlabel polysilicon 709 -2430 709 -2430 0 1
rlabel polysilicon 709 -2436 709 -2436 0 3
rlabel polysilicon 716 -2430 716 -2430 0 1
rlabel polysilicon 716 -2436 716 -2436 0 3
rlabel polysilicon 723 -2430 723 -2430 0 1
rlabel polysilicon 726 -2430 726 -2430 0 2
rlabel polysilicon 723 -2436 723 -2436 0 3
rlabel polysilicon 726 -2436 726 -2436 0 4
rlabel polysilicon 730 -2436 730 -2436 0 3
rlabel polysilicon 733 -2436 733 -2436 0 4
rlabel polysilicon 737 -2430 737 -2430 0 1
rlabel polysilicon 737 -2436 737 -2436 0 3
rlabel polysilicon 744 -2430 744 -2430 0 1
rlabel polysilicon 744 -2436 744 -2436 0 3
rlabel polysilicon 754 -2430 754 -2430 0 2
rlabel polysilicon 754 -2436 754 -2436 0 4
rlabel polysilicon 761 -2430 761 -2430 0 2
rlabel polysilicon 758 -2436 758 -2436 0 3
rlabel polysilicon 761 -2436 761 -2436 0 4
rlabel polysilicon 765 -2430 765 -2430 0 1
rlabel polysilicon 765 -2436 765 -2436 0 3
rlabel polysilicon 772 -2430 772 -2430 0 1
rlabel polysilicon 772 -2436 772 -2436 0 3
rlabel polysilicon 779 -2436 779 -2436 0 3
rlabel polysilicon 807 -2430 807 -2430 0 1
rlabel polysilicon 807 -2436 807 -2436 0 3
rlabel polysilicon 828 -2430 828 -2430 0 1
rlabel polysilicon 828 -2436 828 -2436 0 3
rlabel polysilicon 884 -2430 884 -2430 0 1
rlabel polysilicon 884 -2436 884 -2436 0 3
rlabel polysilicon 891 -2430 891 -2430 0 1
rlabel polysilicon 891 -2436 891 -2436 0 3
rlabel polysilicon 926 -2430 926 -2430 0 1
rlabel polysilicon 926 -2436 926 -2436 0 3
rlabel polysilicon 940 -2430 940 -2430 0 1
rlabel polysilicon 940 -2436 940 -2436 0 3
rlabel polysilicon 5 -2477 5 -2477 0 4
rlabel polysilicon 65 -2477 65 -2477 0 3
rlabel polysilicon 72 -2471 72 -2471 0 1
rlabel polysilicon 72 -2477 72 -2477 0 3
rlabel polysilicon 100 -2471 100 -2471 0 1
rlabel polysilicon 100 -2477 100 -2477 0 3
rlabel polysilicon 107 -2471 107 -2471 0 1
rlabel polysilicon 107 -2477 107 -2477 0 3
rlabel polysilicon 114 -2471 114 -2471 0 1
rlabel polysilicon 117 -2471 117 -2471 0 2
rlabel polysilicon 114 -2477 114 -2477 0 3
rlabel polysilicon 121 -2471 121 -2471 0 1
rlabel polysilicon 121 -2477 121 -2477 0 3
rlabel polysilicon 131 -2471 131 -2471 0 2
rlabel polysilicon 131 -2477 131 -2477 0 4
rlabel polysilicon 135 -2471 135 -2471 0 1
rlabel polysilicon 135 -2477 135 -2477 0 3
rlabel polysilicon 163 -2471 163 -2471 0 1
rlabel polysilicon 163 -2477 163 -2477 0 3
rlabel polysilicon 170 -2471 170 -2471 0 1
rlabel polysilicon 170 -2477 170 -2477 0 3
rlabel polysilicon 177 -2471 177 -2471 0 1
rlabel polysilicon 177 -2477 177 -2477 0 3
rlabel polysilicon 184 -2471 184 -2471 0 1
rlabel polysilicon 187 -2477 187 -2477 0 4
rlabel polysilicon 191 -2471 191 -2471 0 1
rlabel polysilicon 191 -2477 191 -2477 0 3
rlabel polysilicon 198 -2471 198 -2471 0 1
rlabel polysilicon 198 -2477 198 -2477 0 3
rlabel polysilicon 205 -2471 205 -2471 0 1
rlabel polysilicon 205 -2477 205 -2477 0 3
rlabel polysilicon 219 -2471 219 -2471 0 1
rlabel polysilicon 219 -2477 219 -2477 0 3
rlabel polysilicon 226 -2471 226 -2471 0 1
rlabel polysilicon 226 -2477 226 -2477 0 3
rlabel polysilicon 233 -2471 233 -2471 0 1
rlabel polysilicon 233 -2477 233 -2477 0 3
rlabel polysilicon 236 -2477 236 -2477 0 4
rlabel polysilicon 240 -2471 240 -2471 0 1
rlabel polysilicon 247 -2471 247 -2471 0 1
rlabel polysilicon 247 -2477 247 -2477 0 3
rlabel polysilicon 257 -2471 257 -2471 0 2
rlabel polysilicon 264 -2471 264 -2471 0 2
rlabel polysilicon 261 -2477 261 -2477 0 3
rlabel polysilicon 268 -2471 268 -2471 0 1
rlabel polysilicon 268 -2477 268 -2477 0 3
rlabel polysilicon 275 -2471 275 -2471 0 1
rlabel polysilicon 275 -2477 275 -2477 0 3
rlabel polysilicon 282 -2471 282 -2471 0 1
rlabel polysilicon 282 -2477 282 -2477 0 3
rlabel polysilicon 289 -2471 289 -2471 0 1
rlabel polysilicon 289 -2477 289 -2477 0 3
rlabel polysilicon 299 -2471 299 -2471 0 2
rlabel polysilicon 296 -2477 296 -2477 0 3
rlabel polysilicon 303 -2471 303 -2471 0 1
rlabel polysilicon 303 -2477 303 -2477 0 3
rlabel polysilicon 310 -2471 310 -2471 0 1
rlabel polysilicon 310 -2477 310 -2477 0 3
rlabel polysilicon 317 -2471 317 -2471 0 1
rlabel polysilicon 317 -2477 317 -2477 0 3
rlabel polysilicon 324 -2477 324 -2477 0 3
rlabel polysilicon 331 -2471 331 -2471 0 1
rlabel polysilicon 331 -2477 331 -2477 0 3
rlabel polysilicon 338 -2471 338 -2471 0 1
rlabel polysilicon 338 -2477 338 -2477 0 3
rlabel polysilicon 345 -2471 345 -2471 0 1
rlabel polysilicon 348 -2471 348 -2471 0 2
rlabel polysilicon 352 -2471 352 -2471 0 1
rlabel polysilicon 352 -2477 352 -2477 0 3
rlabel polysilicon 359 -2471 359 -2471 0 1
rlabel polysilicon 359 -2477 359 -2477 0 3
rlabel polysilicon 369 -2471 369 -2471 0 2
rlabel polysilicon 366 -2477 366 -2477 0 3
rlabel polysilicon 373 -2471 373 -2471 0 1
rlabel polysilicon 373 -2477 373 -2477 0 3
rlabel polysilicon 376 -2477 376 -2477 0 4
rlabel polysilicon 380 -2471 380 -2471 0 1
rlabel polysilicon 380 -2477 380 -2477 0 3
rlabel polysilicon 387 -2471 387 -2471 0 1
rlabel polysilicon 390 -2471 390 -2471 0 2
rlabel polysilicon 394 -2471 394 -2471 0 1
rlabel polysilicon 394 -2477 394 -2477 0 3
rlabel polysilicon 401 -2471 401 -2471 0 1
rlabel polysilicon 401 -2477 401 -2477 0 3
rlabel polysilicon 408 -2471 408 -2471 0 1
rlabel polysilicon 408 -2477 408 -2477 0 3
rlabel polysilicon 415 -2471 415 -2471 0 1
rlabel polysilicon 415 -2477 415 -2477 0 3
rlabel polysilicon 422 -2471 422 -2471 0 1
rlabel polysilicon 422 -2477 422 -2477 0 3
rlabel polysilicon 432 -2471 432 -2471 0 2
rlabel polysilicon 432 -2477 432 -2477 0 4
rlabel polysilicon 436 -2471 436 -2471 0 1
rlabel polysilicon 436 -2477 436 -2477 0 3
rlabel polysilicon 443 -2471 443 -2471 0 1
rlabel polysilicon 443 -2477 443 -2477 0 3
rlabel polysilicon 450 -2471 450 -2471 0 1
rlabel polysilicon 450 -2477 450 -2477 0 3
rlabel polysilicon 457 -2471 457 -2471 0 1
rlabel polysilicon 457 -2477 457 -2477 0 3
rlabel polysilicon 467 -2477 467 -2477 0 4
rlabel polysilicon 471 -2471 471 -2471 0 1
rlabel polysilicon 471 -2477 471 -2477 0 3
rlabel polysilicon 478 -2471 478 -2471 0 1
rlabel polysilicon 478 -2477 478 -2477 0 3
rlabel polysilicon 502 -2471 502 -2471 0 2
rlabel polysilicon 502 -2477 502 -2477 0 4
rlabel polysilicon 506 -2471 506 -2471 0 1
rlabel polysilicon 506 -2477 506 -2477 0 3
rlabel polysilicon 513 -2471 513 -2471 0 1
rlabel polysilicon 513 -2477 513 -2477 0 3
rlabel polysilicon 520 -2477 520 -2477 0 3
rlabel polysilicon 523 -2477 523 -2477 0 4
rlabel polysilicon 527 -2477 527 -2477 0 3
rlabel polysilicon 534 -2471 534 -2471 0 1
rlabel polysilicon 537 -2477 537 -2477 0 4
rlabel polysilicon 541 -2471 541 -2471 0 1
rlabel polysilicon 541 -2477 541 -2477 0 3
rlabel polysilicon 548 -2471 548 -2471 0 1
rlabel polysilicon 548 -2477 548 -2477 0 3
rlabel polysilicon 569 -2471 569 -2471 0 1
rlabel polysilicon 569 -2477 569 -2477 0 3
rlabel polysilicon 576 -2471 576 -2471 0 1
rlabel polysilicon 576 -2477 576 -2477 0 3
rlabel polysilicon 586 -2477 586 -2477 0 4
rlabel polysilicon 593 -2471 593 -2471 0 2
rlabel polysilicon 590 -2477 590 -2477 0 3
rlabel polysilicon 600 -2471 600 -2471 0 2
rlabel polysilicon 597 -2477 597 -2477 0 3
rlabel polysilicon 604 -2471 604 -2471 0 1
rlabel polysilicon 604 -2477 604 -2477 0 3
rlabel polysilicon 611 -2471 611 -2471 0 1
rlabel polysilicon 611 -2477 611 -2477 0 3
rlabel polysilicon 625 -2471 625 -2471 0 1
rlabel polysilicon 625 -2477 625 -2477 0 3
rlabel polysilicon 639 -2471 639 -2471 0 1
rlabel polysilicon 642 -2471 642 -2471 0 2
rlabel polysilicon 660 -2471 660 -2471 0 1
rlabel polysilicon 660 -2477 660 -2477 0 3
rlabel polysilicon 674 -2471 674 -2471 0 1
rlabel polysilicon 674 -2477 674 -2477 0 3
rlabel polysilicon 681 -2471 681 -2471 0 1
rlabel polysilicon 681 -2477 681 -2477 0 3
rlabel polysilicon 688 -2471 688 -2471 0 1
rlabel polysilicon 688 -2477 688 -2477 0 3
rlabel polysilicon 695 -2471 695 -2471 0 1
rlabel polysilicon 695 -2477 695 -2477 0 3
rlabel polysilicon 709 -2471 709 -2471 0 1
rlabel polysilicon 709 -2477 709 -2477 0 3
rlabel polysilicon 716 -2471 716 -2471 0 1
rlabel polysilicon 716 -2477 716 -2477 0 3
rlabel polysilicon 723 -2471 723 -2471 0 1
rlabel polysilicon 723 -2477 723 -2477 0 3
rlabel polysilicon 730 -2471 730 -2471 0 1
rlabel polysilicon 730 -2477 730 -2477 0 3
rlabel polysilicon 737 -2471 737 -2471 0 1
rlabel polysilicon 737 -2477 737 -2477 0 3
rlabel polysilicon 758 -2471 758 -2471 0 1
rlabel polysilicon 761 -2471 761 -2471 0 2
rlabel polysilicon 758 -2477 758 -2477 0 3
rlabel polysilicon 761 -2477 761 -2477 0 4
rlabel polysilicon 765 -2471 765 -2471 0 1
rlabel polysilicon 765 -2477 765 -2477 0 3
rlabel polysilicon 884 -2471 884 -2471 0 1
rlabel polysilicon 884 -2477 884 -2477 0 3
rlabel polysilicon 891 -2471 891 -2471 0 1
rlabel polysilicon 891 -2477 891 -2477 0 3
rlabel polysilicon 933 -2471 933 -2471 0 1
rlabel polysilicon 936 -2477 936 -2477 0 4
rlabel polysilicon 940 -2471 940 -2471 0 1
rlabel polysilicon 940 -2477 940 -2477 0 3
rlabel polysilicon 5 -2498 5 -2498 0 2
rlabel polysilicon 5 -2504 5 -2504 0 4
rlabel polysilicon 86 -2498 86 -2498 0 1
rlabel polysilicon 86 -2504 86 -2504 0 3
rlabel polysilicon 96 -2498 96 -2498 0 2
rlabel polysilicon 100 -2498 100 -2498 0 1
rlabel polysilicon 100 -2504 100 -2504 0 3
rlabel polysilicon 103 -2504 103 -2504 0 4
rlabel polysilicon 110 -2498 110 -2498 0 2
rlabel polysilicon 107 -2504 107 -2504 0 3
rlabel polysilicon 114 -2498 114 -2498 0 1
rlabel polysilicon 117 -2504 117 -2504 0 4
rlabel polysilicon 121 -2498 121 -2498 0 1
rlabel polysilicon 121 -2504 121 -2504 0 3
rlabel polysilicon 138 -2498 138 -2498 0 2
rlabel polysilicon 142 -2498 142 -2498 0 1
rlabel polysilicon 142 -2504 142 -2504 0 3
rlabel polysilicon 149 -2498 149 -2498 0 1
rlabel polysilicon 149 -2504 149 -2504 0 3
rlabel polysilicon 159 -2498 159 -2498 0 2
rlabel polysilicon 156 -2504 156 -2504 0 3
rlabel polysilicon 163 -2504 163 -2504 0 3
rlabel polysilicon 166 -2504 166 -2504 0 4
rlabel polysilicon 170 -2498 170 -2498 0 1
rlabel polysilicon 170 -2504 170 -2504 0 3
rlabel polysilicon 177 -2498 177 -2498 0 1
rlabel polysilicon 177 -2504 177 -2504 0 3
rlabel polysilicon 187 -2504 187 -2504 0 4
rlabel polysilicon 191 -2504 191 -2504 0 3
rlabel polysilicon 194 -2504 194 -2504 0 4
rlabel polysilicon 201 -2498 201 -2498 0 2
rlabel polysilicon 201 -2504 201 -2504 0 4
rlabel polysilicon 205 -2498 205 -2498 0 1
rlabel polysilicon 205 -2504 205 -2504 0 3
rlabel polysilicon 212 -2498 212 -2498 0 1
rlabel polysilicon 212 -2504 212 -2504 0 3
rlabel polysilicon 219 -2498 219 -2498 0 1
rlabel polysilicon 219 -2504 219 -2504 0 3
rlabel polysilicon 226 -2498 226 -2498 0 1
rlabel polysilicon 226 -2504 226 -2504 0 3
rlabel polysilicon 233 -2498 233 -2498 0 1
rlabel polysilicon 233 -2504 233 -2504 0 3
rlabel polysilicon 240 -2498 240 -2498 0 1
rlabel polysilicon 240 -2504 240 -2504 0 3
rlabel polysilicon 247 -2498 247 -2498 0 1
rlabel polysilicon 247 -2504 247 -2504 0 3
rlabel polysilicon 254 -2498 254 -2498 0 1
rlabel polysilicon 254 -2504 254 -2504 0 3
rlabel polysilicon 261 -2498 261 -2498 0 1
rlabel polysilicon 261 -2504 261 -2504 0 3
rlabel polysilicon 271 -2498 271 -2498 0 2
rlabel polysilicon 268 -2504 268 -2504 0 3
rlabel polysilicon 275 -2498 275 -2498 0 1
rlabel polysilicon 275 -2504 275 -2504 0 3
rlabel polysilicon 282 -2504 282 -2504 0 3
rlabel polysilicon 289 -2498 289 -2498 0 1
rlabel polysilicon 289 -2504 289 -2504 0 3
rlabel polysilicon 296 -2498 296 -2498 0 1
rlabel polysilicon 299 -2504 299 -2504 0 4
rlabel polysilicon 303 -2498 303 -2498 0 1
rlabel polysilicon 303 -2504 303 -2504 0 3
rlabel polysilicon 310 -2498 310 -2498 0 1
rlabel polysilicon 310 -2504 310 -2504 0 3
rlabel polysilicon 317 -2498 317 -2498 0 1
rlabel polysilicon 317 -2504 317 -2504 0 3
rlabel polysilicon 324 -2498 324 -2498 0 1
rlabel polysilicon 324 -2504 324 -2504 0 3
rlabel polysilicon 331 -2498 331 -2498 0 1
rlabel polysilicon 331 -2504 331 -2504 0 3
rlabel polysilicon 352 -2498 352 -2498 0 1
rlabel polysilicon 352 -2504 352 -2504 0 3
rlabel polysilicon 359 -2498 359 -2498 0 1
rlabel polysilicon 362 -2498 362 -2498 0 2
rlabel polysilicon 380 -2498 380 -2498 0 1
rlabel polysilicon 380 -2504 380 -2504 0 3
rlabel polysilicon 387 -2504 387 -2504 0 3
rlabel polysilicon 394 -2498 394 -2498 0 1
rlabel polysilicon 394 -2504 394 -2504 0 3
rlabel polysilicon 401 -2498 401 -2498 0 1
rlabel polysilicon 404 -2498 404 -2498 0 2
rlabel polysilicon 401 -2504 401 -2504 0 3
rlabel polysilicon 404 -2504 404 -2504 0 4
rlabel polysilicon 408 -2498 408 -2498 0 1
rlabel polysilicon 408 -2504 408 -2504 0 3
rlabel polysilicon 418 -2504 418 -2504 0 4
rlabel polysilicon 422 -2498 422 -2498 0 1
rlabel polysilicon 443 -2498 443 -2498 0 1
rlabel polysilicon 443 -2504 443 -2504 0 3
rlabel polysilicon 450 -2498 450 -2498 0 1
rlabel polysilicon 450 -2504 450 -2504 0 3
rlabel polysilicon 520 -2498 520 -2498 0 1
rlabel polysilicon 523 -2498 523 -2498 0 2
rlabel polysilicon 527 -2498 527 -2498 0 1
rlabel polysilicon 527 -2504 527 -2504 0 3
rlabel polysilicon 604 -2498 604 -2498 0 1
rlabel polysilicon 604 -2504 604 -2504 0 3
rlabel polysilicon 611 -2498 611 -2498 0 1
rlabel polysilicon 611 -2504 611 -2504 0 3
rlabel polysilicon 660 -2498 660 -2498 0 1
rlabel polysilicon 660 -2504 660 -2504 0 3
rlabel polysilicon 667 -2498 667 -2498 0 1
rlabel polysilicon 667 -2504 667 -2504 0 3
rlabel polysilicon 681 -2498 681 -2498 0 1
rlabel polysilicon 681 -2504 681 -2504 0 3
rlabel polysilicon 688 -2498 688 -2498 0 1
rlabel polysilicon 688 -2504 688 -2504 0 3
rlabel polysilicon 695 -2498 695 -2498 0 1
rlabel polysilicon 695 -2504 695 -2504 0 3
rlabel polysilicon 702 -2504 702 -2504 0 3
rlabel polysilicon 705 -2504 705 -2504 0 4
rlabel polysilicon 709 -2498 709 -2498 0 1
rlabel polysilicon 709 -2504 709 -2504 0 3
rlabel polysilicon 716 -2498 716 -2498 0 1
rlabel polysilicon 716 -2504 716 -2504 0 3
rlabel polysilicon 723 -2498 723 -2498 0 1
rlabel polysilicon 723 -2504 723 -2504 0 3
rlabel polysilicon 730 -2498 730 -2498 0 1
rlabel polysilicon 740 -2504 740 -2504 0 4
rlabel polysilicon 744 -2498 744 -2498 0 1
rlabel polysilicon 744 -2504 744 -2504 0 3
rlabel polysilicon 751 -2498 751 -2498 0 1
rlabel polysilicon 751 -2504 751 -2504 0 3
rlabel polysilicon 758 -2498 758 -2498 0 1
rlabel polysilicon 758 -2504 758 -2504 0 3
rlabel polysilicon 884 -2498 884 -2498 0 1
rlabel polysilicon 887 -2504 887 -2504 0 4
rlabel polysilicon 891 -2498 891 -2498 0 1
rlabel polysilicon 891 -2504 891 -2504 0 3
rlabel polysilicon 933 -2498 933 -2498 0 1
rlabel polysilicon 933 -2504 933 -2504 0 3
rlabel polysilicon 940 -2504 940 -2504 0 3
rlabel polysilicon 943 -2504 943 -2504 0 4
rlabel polysilicon 947 -2498 947 -2498 0 1
rlabel polysilicon 947 -2504 947 -2504 0 3
rlabel polysilicon 5 -2523 5 -2523 0 4
rlabel polysilicon 9 -2517 9 -2517 0 1
rlabel polysilicon 9 -2523 9 -2523 0 3
rlabel polysilicon 100 -2523 100 -2523 0 3
rlabel polysilicon 107 -2517 107 -2517 0 1
rlabel polysilicon 107 -2523 107 -2523 0 3
rlabel polysilicon 114 -2517 114 -2517 0 1
rlabel polysilicon 114 -2523 114 -2523 0 3
rlabel polysilicon 121 -2523 121 -2523 0 3
rlabel polysilicon 124 -2523 124 -2523 0 4
rlabel polysilicon 131 -2523 131 -2523 0 4
rlabel polysilicon 159 -2517 159 -2517 0 2
rlabel polysilicon 163 -2517 163 -2517 0 1
rlabel polysilicon 163 -2523 163 -2523 0 3
rlabel polysilicon 170 -2523 170 -2523 0 3
rlabel polysilicon 180 -2517 180 -2517 0 2
rlabel polysilicon 180 -2523 180 -2523 0 4
rlabel polysilicon 184 -2517 184 -2517 0 1
rlabel polysilicon 184 -2523 184 -2523 0 3
rlabel polysilicon 191 -2517 191 -2517 0 1
rlabel polysilicon 191 -2523 191 -2523 0 3
rlabel polysilicon 198 -2523 198 -2523 0 3
rlabel polysilicon 226 -2517 226 -2517 0 1
rlabel polysilicon 229 -2517 229 -2517 0 2
rlabel polysilicon 271 -2517 271 -2517 0 2
rlabel polysilicon 278 -2517 278 -2517 0 2
rlabel polysilicon 285 -2517 285 -2517 0 2
rlabel polysilicon 292 -2523 292 -2523 0 4
rlabel polysilicon 296 -2517 296 -2517 0 1
rlabel polysilicon 296 -2523 296 -2523 0 3
rlabel polysilicon 303 -2523 303 -2523 0 3
rlabel polysilicon 310 -2517 310 -2517 0 1
rlabel polysilicon 310 -2523 310 -2523 0 3
rlabel polysilicon 341 -2517 341 -2517 0 2
rlabel polysilicon 341 -2523 341 -2523 0 4
rlabel polysilicon 345 -2517 345 -2517 0 1
rlabel polysilicon 345 -2523 345 -2523 0 3
rlabel polysilicon 362 -2517 362 -2517 0 2
rlabel polysilicon 383 -2517 383 -2517 0 2
rlabel polysilicon 397 -2517 397 -2517 0 2
rlabel polysilicon 404 -2517 404 -2517 0 2
rlabel polysilicon 450 -2517 450 -2517 0 1
rlabel polysilicon 450 -2523 450 -2523 0 3
rlabel polysilicon 457 -2517 457 -2517 0 1
rlabel polysilicon 457 -2523 457 -2523 0 3
rlabel polysilicon 523 -2517 523 -2517 0 2
rlabel polysilicon 597 -2517 597 -2517 0 1
rlabel polysilicon 597 -2523 597 -2523 0 3
rlabel polysilicon 604 -2517 604 -2517 0 1
rlabel polysilicon 604 -2523 604 -2523 0 3
rlabel polysilicon 663 -2517 663 -2517 0 2
rlabel polysilicon 663 -2523 663 -2523 0 4
rlabel polysilicon 667 -2517 667 -2517 0 1
rlabel polysilicon 667 -2523 667 -2523 0 3
rlabel polysilicon 688 -2517 688 -2517 0 1
rlabel polysilicon 712 -2517 712 -2517 0 2
rlabel polysilicon 716 -2517 716 -2517 0 1
rlabel polysilicon 716 -2523 716 -2523 0 3
rlabel polysilicon 723 -2523 723 -2523 0 3
rlabel polysilicon 730 -2517 730 -2517 0 1
rlabel polysilicon 730 -2523 730 -2523 0 3
rlabel polysilicon 740 -2523 740 -2523 0 4
rlabel metal2 93 1 93 1 0 net=4475
rlabel metal2 107 1 107 1 0 net=3023
rlabel metal2 205 1 205 1 0 net=6135
rlabel metal2 215 1 215 1 0 net=1006
rlabel metal2 240 1 240 1 0 net=6909
rlabel metal2 261 1 261 1 0 net=4495
rlabel metal2 324 1 324 1 0 net=3651
rlabel metal2 429 1 429 1 0 net=6425
rlabel metal2 464 1 464 1 0 net=5447
rlabel metal2 530 1 530 1 0 net=6287
rlabel metal2 583 1 583 1 0 net=7017
rlabel metal2 660 1 660 1 0 net=7317
rlabel metal2 117 -1 117 -1 0 net=4617
rlabel metal2 226 -1 226 -1 0 net=5669
rlabel metal2 86 -12 86 -12 0 net=779
rlabel metal2 117 -12 117 -12 0 net=3024
rlabel metal2 135 -12 135 -12 0 net=5877
rlabel metal2 173 -12 173 -12 0 net=1453
rlabel metal2 205 -12 205 -12 0 net=6136
rlabel metal2 226 -12 226 -12 0 net=5670
rlabel metal2 254 -12 254 -12 0 net=4497
rlabel metal2 289 -12 289 -12 0 net=2755
rlabel metal2 310 -12 310 -12 0 net=3653
rlabel metal2 348 -12 348 -12 0 net=3845
rlabel metal2 373 -12 373 -12 0 net=4043
rlabel metal2 450 -12 450 -12 0 net=5448
rlabel metal2 485 -12 485 -12 0 net=7291
rlabel metal2 534 -12 534 -12 0 net=6289
rlabel metal2 548 -12 548 -12 0 net=6173
rlabel metal2 590 -12 590 -12 0 net=6889
rlabel metal2 607 -12 607 -12 0 net=7495
rlabel metal2 667 -12 667 -12 0 net=7319
rlabel metal2 89 -14 89 -14 0 net=413
rlabel metal2 177 -14 177 -14 0 net=1427
rlabel metal2 219 -14 219 -14 0 net=2153
rlabel metal2 233 -14 233 -14 0 net=4961
rlabel metal2 257 -14 257 -14 0 net=3971
rlabel metal2 317 -14 317 -14 0 net=7537
rlabel metal2 415 -14 415 -14 0 net=6427
rlabel metal2 453 -14 453 -14 0 net=6009
rlabel metal2 492 -14 492 -14 0 net=4005
rlabel metal2 562 -14 562 -14 0 net=5847
rlabel metal2 597 -14 597 -14 0 net=7019
rlabel metal2 93 -16 93 -16 0 net=4476
rlabel metal2 184 -16 184 -16 0 net=2541
rlabel metal2 219 -16 219 -16 0 net=1853
rlabel metal2 240 -16 240 -16 0 net=6910
rlabel metal2 240 -16 240 -16 0 net=6910
rlabel metal2 261 -16 261 -16 0 net=3573
rlabel metal2 324 -16 324 -16 0 net=1723
rlabel metal2 429 -16 429 -16 0 net=3961
rlabel metal2 506 -16 506 -16 0 net=7091
rlabel metal2 100 -18 100 -18 0 net=4618
rlabel metal2 236 -18 236 -18 0 net=3147
rlabel metal2 268 -20 268 -20 0 net=1241
rlabel metal2 86 -31 86 -31 0 net=3235
rlabel metal2 114 -31 114 -31 0 net=2165
rlabel metal2 191 -31 191 -31 0 net=1855
rlabel metal2 226 -31 226 -31 0 net=2155
rlabel metal2 247 -31 247 -31 0 net=4963
rlabel metal2 359 -31 359 -31 0 net=3847
rlabel metal2 415 -31 415 -31 0 net=6428
rlabel metal2 429 -31 429 -31 0 net=3963
rlabel metal2 446 -31 446 -31 0 net=4335
rlabel metal2 506 -31 506 -31 0 net=7093
rlabel metal2 506 -31 506 -31 0 net=7093
rlabel metal2 520 -31 520 -31 0 net=6649
rlabel metal2 551 -31 551 -31 0 net=4909
rlabel metal2 569 -31 569 -31 0 net=6175
rlabel metal2 604 -31 604 -31 0 net=6891
rlabel metal2 663 -31 663 -31 0 net=7539
rlabel metal2 674 -31 674 -31 0 net=7321
rlabel metal2 765 -31 765 -31 0 net=7199
rlabel metal2 93 -33 93 -33 0 net=3477
rlabel metal2 121 -33 121 -33 0 net=5879
rlabel metal2 163 -33 163 -33 0 net=1763
rlabel metal2 247 -33 247 -33 0 net=4498
rlabel metal2 275 -33 275 -33 0 net=3973
rlabel metal2 366 -33 366 -33 0 net=4045
rlabel metal2 383 -33 383 -33 0 net=4425
rlabel metal2 471 -33 471 -33 0 net=6011
rlabel metal2 527 -33 527 -33 0 net=7293
rlabel metal2 611 -33 611 -33 0 net=7021
rlabel metal2 677 -33 677 -33 0 net=6985
rlabel metal2 128 -35 128 -35 0 net=4891
rlabel metal2 177 -35 177 -35 0 net=1428
rlabel metal2 198 -35 198 -35 0 net=1455
rlabel metal2 212 -35 212 -35 0 net=134
rlabel metal2 282 -35 282 -35 0 net=3149
rlabel metal2 313 -35 313 -35 0 net=7538
rlabel metal2 338 -35 338 -35 0 net=891
rlabel metal2 338 -35 338 -35 0 net=891
rlabel metal2 341 -35 341 -35 0 net=4731
rlabel metal2 464 -35 464 -35 0 net=6931
rlabel metal2 618 -35 618 -35 0 net=7497
rlabel metal2 135 -37 135 -37 0 net=1243
rlabel metal2 282 -37 282 -37 0 net=2533
rlabel metal2 373 -37 373 -37 0 net=5277
rlabel metal2 464 -37 464 -37 0 net=7577
rlabel metal2 156 -39 156 -39 0 net=5527
rlabel metal2 184 -39 184 -39 0 net=2543
rlabel metal2 226 -39 226 -39 0 net=3575
rlabel metal2 268 -39 268 -39 0 net=2757
rlabel metal2 296 -39 296 -39 0 net=7545
rlabel metal2 471 -39 471 -39 0 net=4885
rlabel metal2 198 -41 198 -41 0 net=6525
rlabel metal2 383 -41 383 -41 0 net=4447
rlabel metal2 527 -41 527 -41 0 net=7397
rlabel metal2 201 -43 201 -43 0 net=4941
rlabel metal2 289 -43 289 -43 0 net=1725
rlabel metal2 387 -43 387 -43 0 net=1323
rlabel metal2 478 -43 478 -43 0 net=4007
rlabel metal2 541 -43 541 -43 0 net=6291
rlabel metal2 576 -43 576 -43 0 net=5849
rlabel metal2 576 -43 576 -43 0 net=5849
rlabel metal2 173 -45 173 -45 0 net=3649
rlabel metal2 513 -45 513 -45 0 net=5073
rlabel metal2 555 -45 555 -45 0 net=6763
rlabel metal2 212 -47 212 -47 0 net=3433
rlabel metal2 310 -47 310 -47 0 net=3655
rlabel metal2 555 -47 555 -47 0 net=6823
rlabel metal2 250 -51 250 -51 0 net=5657
rlabel metal2 30 -62 30 -62 0 net=4277
rlabel metal2 159 -62 159 -62 0 net=1193
rlabel metal2 317 -62 317 -62 0 net=3657
rlabel metal2 429 -62 429 -62 0 net=7547
rlabel metal2 842 -62 842 -62 0 net=7201
rlabel metal2 58 -64 58 -64 0 net=3005
rlabel metal2 114 -64 114 -64 0 net=2166
rlabel metal2 198 -64 198 -64 0 net=1457
rlabel metal2 219 -64 219 -64 0 net=2544
rlabel metal2 233 -64 233 -64 0 net=3974
rlabel metal2 394 -64 394 -64 0 net=4427
rlabel metal2 450 -64 450 -64 0 net=4507
rlabel metal2 471 -64 471 -64 0 net=4887
rlabel metal2 485 -64 485 -64 0 net=4449
rlabel metal2 530 -64 530 -64 0 net=2051
rlabel metal2 702 -64 702 -64 0 net=7323
rlabel metal2 37 -66 37 -66 0 net=2013
rlabel metal2 219 -66 219 -66 0 net=1839
rlabel metal2 317 -66 317 -66 0 net=6555
rlabel metal2 772 -66 772 -66 0 net=6825
rlabel metal2 61 -68 61 -68 0 net=653
rlabel metal2 324 -68 324 -68 0 net=3650
rlabel metal2 457 -68 457 -68 0 net=4333
rlabel metal2 583 -68 583 -68 0 net=7403
rlabel metal2 65 -70 65 -70 0 net=3479
rlabel metal2 100 -70 100 -70 0 net=1301
rlabel metal2 233 -70 233 -70 0 net=1325
rlabel metal2 464 -70 464 -70 0 net=4009
rlabel metal2 485 -70 485 -70 0 net=4337
rlabel metal2 502 -70 502 -70 0 net=6895
rlabel metal2 72 -72 72 -72 0 net=4893
rlabel metal2 142 -72 142 -72 0 net=1821
rlabel metal2 254 -72 254 -72 0 net=4943
rlabel metal2 590 -72 590 -72 0 net=7295
rlabel metal2 79 -74 79 -74 0 net=3236
rlabel metal2 93 -74 93 -74 0 net=3151
rlabel metal2 331 -74 331 -74 0 net=6527
rlabel metal2 702 -74 702 -74 0 net=6157
rlabel metal2 86 -76 86 -76 0 net=2535
rlabel metal2 289 -76 289 -76 0 net=1727
rlabel metal2 331 -76 331 -76 0 net=4965
rlabel metal2 376 -76 376 -76 0 net=4519
rlabel metal2 495 -76 495 -76 0 net=7673
rlabel metal2 103 -78 103 -78 0 net=2093
rlabel metal2 380 -78 380 -78 0 net=3849
rlabel metal2 471 -78 471 -78 0 net=3159
rlabel metal2 506 -78 506 -78 0 net=7094
rlabel metal2 548 -78 548 -78 0 net=5701
rlabel metal2 625 -78 625 -78 0 net=7579
rlabel metal2 117 -80 117 -80 0 net=1110
rlabel metal2 240 -80 240 -80 0 net=3863
rlabel metal2 569 -80 569 -80 0 net=6293
rlabel metal2 632 -80 632 -80 0 net=7399
rlabel metal2 51 -82 51 -82 0 net=3327
rlabel metal2 261 -82 261 -82 0 net=2157
rlabel metal2 355 -82 355 -82 0 net=5763
rlabel metal2 639 -82 639 -82 0 net=6893
rlabel metal2 121 -84 121 -84 0 net=5881
rlabel metal2 268 -84 268 -84 0 net=2759
rlabel metal2 387 -84 387 -84 0 net=7751
rlabel metal2 121 -86 121 -86 0 net=1765
rlabel metal2 247 -86 247 -86 0 net=4311
rlabel metal2 268 -86 268 -86 0 net=2343
rlabel metal2 397 -86 397 -86 0 net=4765
rlabel metal2 586 -86 586 -86 0 net=5135
rlabel metal2 604 -86 604 -86 0 net=6765
rlabel metal2 128 -88 128 -88 0 net=6273
rlabel metal2 681 -88 681 -88 0 net=6987
rlabel metal2 149 -90 149 -90 0 net=5528
rlabel metal2 163 -90 163 -90 0 net=2447
rlabel metal2 527 -90 527 -90 0 net=4291
rlabel metal2 597 -90 597 -90 0 net=6177
rlabel metal2 709 -90 709 -90 0 net=6493
rlabel metal2 401 -92 401 -92 0 net=5659
rlabel metal2 576 -92 576 -92 0 net=5851
rlabel metal2 611 -92 611 -92 0 net=6933
rlabel metal2 366 -94 366 -94 0 net=4047
rlabel metal2 443 -94 443 -94 0 net=5279
rlabel metal2 646 -94 646 -94 0 net=7499
rlabel metal2 359 -96 359 -96 0 net=1619
rlabel metal2 653 -96 653 -96 0 net=7023
rlabel metal2 226 -98 226 -98 0 net=3577
rlabel metal2 436 -98 436 -98 0 net=3965
rlabel metal2 520 -98 520 -98 0 net=6013
rlabel metal2 660 -98 660 -98 0 net=7501
rlabel metal2 177 -100 177 -100 0 net=414
rlabel metal2 310 -100 310 -100 0 net=4511
rlabel metal2 534 -100 534 -100 0 net=6651
rlabel metal2 667 -100 667 -100 0 net=7541
rlabel metal2 156 -102 156 -102 0 net=6101
rlabel metal2 177 -104 177 -104 0 net=3435
rlabel metal2 310 -104 310 -104 0 net=5247
rlabel metal2 415 -104 415 -104 0 net=3941
rlabel metal2 499 -104 499 -104 0 net=4581
rlabel metal2 541 -104 541 -104 0 net=5075
rlabel metal2 191 -106 191 -106 0 net=1857
rlabel metal2 422 -106 422 -106 0 net=4733
rlabel metal2 562 -106 562 -106 0 net=4911
rlabel metal2 47 -108 47 -108 0 net=4073
rlabel metal2 191 -110 191 -110 0 net=1711
rlabel metal2 296 -112 296 -112 0 net=5013
rlabel metal2 275 -114 275 -114 0 net=3013
rlabel metal2 184 -116 184 -116 0 net=1154
rlabel metal2 135 -118 135 -118 0 net=1245
rlabel metal2 135 -120 135 -120 0 net=4411
rlabel metal2 23 -131 23 -131 0 net=1767
rlabel metal2 128 -131 128 -131 0 net=395
rlabel metal2 226 -131 226 -131 0 net=2052
rlabel metal2 723 -131 723 -131 0 net=6935
rlabel metal2 870 -131 870 -131 0 net=6827
rlabel metal2 1108 -131 1108 -131 0 net=6769
rlabel metal2 1108 -131 1108 -131 0 net=6769
rlabel metal2 30 -133 30 -133 0 net=4278
rlabel metal2 145 -133 145 -133 0 net=3569
rlabel metal2 436 -133 436 -133 0 net=3943
rlabel metal2 436 -133 436 -133 0 net=3943
rlabel metal2 499 -133 499 -133 0 net=6652
rlabel metal2 751 -133 751 -133 0 net=7025
rlabel metal2 877 -133 877 -133 0 net=7203
rlabel metal2 30 -135 30 -135 0 net=2449
rlabel metal2 170 -135 170 -135 0 net=7674
rlabel metal2 37 -137 37 -137 0 net=2015
rlabel metal2 149 -137 149 -137 0 net=3436
rlabel metal2 250 -137 250 -137 0 net=7752
rlabel metal2 37 -139 37 -139 0 net=1303
rlabel metal2 275 -139 275 -139 0 net=5248
rlabel metal2 317 -139 317 -139 0 net=4888
rlabel metal2 509 -139 509 -139 0 net=6766
rlabel metal2 765 -139 765 -139 0 net=7503
rlabel metal2 44 -141 44 -141 0 net=1823
rlabel metal2 156 -141 156 -141 0 net=7548
rlabel metal2 51 -143 51 -143 0 net=1211
rlabel metal2 299 -143 299 -143 0 net=690
rlabel metal2 362 -143 362 -143 0 net=7583
rlabel metal2 51 -145 51 -145 0 net=2229
rlabel metal2 142 -145 142 -145 0 net=3069
rlabel metal2 376 -145 376 -145 0 net=5660
rlabel metal2 579 -145 579 -145 0 net=7500
rlabel metal2 772 -145 772 -145 0 net=7297
rlabel metal2 58 -147 58 -147 0 net=1620
rlabel metal2 660 -147 660 -147 0 net=6079
rlabel metal2 779 -147 779 -147 0 net=7325
rlabel metal2 65 -149 65 -149 0 net=3480
rlabel metal2 117 -149 117 -149 0 net=5187
rlabel metal2 159 -149 159 -149 0 net=282
rlabel metal2 352 -149 352 -149 0 net=4735
rlabel metal2 548 -149 548 -149 0 net=4767
rlabel metal2 79 -151 79 -151 0 net=6274
rlabel metal2 681 -151 681 -151 0 net=6179
rlabel metal2 786 -151 786 -151 0 net=7401
rlabel metal2 79 -153 79 -153 0 net=3637
rlabel metal2 163 -153 163 -153 0 net=1459
rlabel metal2 310 -153 310 -153 0 net=3161
rlabel metal2 495 -153 495 -153 0 net=5235
rlabel metal2 667 -153 667 -153 0 net=6103
rlabel metal2 793 -153 793 -153 0 net=7405
rlabel metal2 86 -155 86 -155 0 net=2536
rlabel metal2 418 -155 418 -155 0 net=5101
rlabel metal2 695 -155 695 -155 0 net=6529
rlabel metal2 89 -157 89 -157 0 net=3797
rlabel metal2 152 -157 152 -157 0 net=6869
rlabel metal2 114 -159 114 -159 0 net=1291
rlabel metal2 198 -159 198 -159 0 net=1859
rlabel metal2 317 -159 317 -159 0 net=3865
rlabel metal2 422 -159 422 -159 0 net=4075
rlabel metal2 513 -159 513 -159 0 net=4451
rlabel metal2 583 -159 583 -159 0 net=7097
rlabel metal2 170 -161 170 -161 0 net=1499
rlabel metal2 320 -161 320 -161 0 net=4048
rlabel metal2 429 -161 429 -161 0 net=4429
rlabel metal2 520 -161 520 -161 0 net=4513
rlabel metal2 583 -161 583 -161 0 net=6989
rlabel metal2 737 -161 737 -161 0 net=7067
rlabel metal2 173 -163 173 -163 0 net=4334
rlabel metal2 464 -163 464 -163 0 net=4011
rlabel metal2 492 -163 492 -163 0 net=5571
rlabel metal2 702 -163 702 -163 0 net=6159
rlabel metal2 800 -163 800 -163 0 net=7543
rlabel metal2 212 -165 212 -165 0 net=2158
rlabel metal2 324 -165 324 -165 0 net=1728
rlabel metal2 359 -165 359 -165 0 net=3579
rlabel metal2 443 -165 443 -165 0 net=3967
rlabel metal2 814 -165 814 -165 0 net=7581
rlabel metal2 65 -167 65 -167 0 net=3767
rlabel metal2 380 -167 380 -167 0 net=3851
rlabel metal2 506 -167 506 -167 0 net=6387
rlabel metal2 93 -169 93 -169 0 net=3153
rlabel metal2 387 -169 387 -169 0 net=5427
rlabel metal2 520 -169 520 -169 0 net=6575
rlabel metal2 93 -171 93 -171 0 net=1247
rlabel metal2 219 -171 219 -171 0 net=1841
rlabel metal2 324 -171 324 -171 0 net=5495
rlabel metal2 709 -171 709 -171 0 net=6495
rlabel metal2 135 -173 135 -173 0 net=3665
rlabel metal2 261 -173 261 -173 0 net=4313
rlabel metal2 523 -173 523 -173 0 net=5783
rlabel metal2 107 -175 107 -175 0 net=3007
rlabel metal2 327 -175 327 -175 0 net=3658
rlabel metal2 345 -175 345 -175 0 net=3339
rlabel metal2 534 -175 534 -175 0 net=4583
rlabel metal2 590 -175 590 -175 0 net=5137
rlabel metal2 716 -175 716 -175 0 net=6557
rlabel metal2 184 -177 184 -177 0 net=1713
rlabel metal2 268 -177 268 -177 0 net=2345
rlabel metal2 348 -177 348 -177 0 net=4292
rlabel metal2 597 -177 597 -177 0 net=5853
rlabel metal2 72 -179 72 -179 0 net=4895
rlabel metal2 611 -179 611 -179 0 net=5281
rlabel metal2 72 -181 72 -181 0 net=5619
rlabel metal2 191 -183 191 -183 0 net=1693
rlabel metal2 268 -183 268 -183 0 net=2761
rlabel metal2 331 -183 331 -183 0 net=4967
rlabel metal2 450 -183 450 -183 0 net=4509
rlabel metal2 555 -183 555 -183 0 net=4945
rlabel metal2 618 -183 618 -183 0 net=5703
rlabel metal2 205 -185 205 -185 0 net=2253
rlabel metal2 334 -185 334 -185 0 net=1114
rlabel metal2 366 -187 366 -187 0 net=4413
rlabel metal2 478 -187 478 -187 0 net=4521
rlabel metal2 618 -187 618 -187 0 net=6945
rlabel metal2 296 -189 296 -189 0 net=3015
rlabel metal2 394 -189 394 -189 0 net=5457
rlabel metal2 282 -191 282 -191 0 net=2094
rlabel metal2 401 -191 401 -191 0 net=3635
rlabel metal2 240 -193 240 -193 0 net=3329
rlabel metal2 296 -193 296 -193 0 net=4809
rlabel metal2 625 -193 625 -193 0 net=6295
rlabel metal2 240 -195 240 -195 0 net=5883
rlabel metal2 478 -195 478 -195 0 net=5015
rlabel metal2 625 -195 625 -195 0 net=6521
rlabel metal2 233 -197 233 -197 0 net=1327
rlabel metal2 345 -197 345 -197 0 net=4541
rlabel metal2 632 -197 632 -197 0 net=5765
rlabel metal2 58 -199 58 -199 0 net=3291
rlabel metal2 485 -199 485 -199 0 net=4339
rlabel metal2 604 -199 604 -199 0 net=5077
rlabel metal2 110 -201 110 -201 0 net=6191
rlabel metal2 576 -201 576 -201 0 net=4913
rlabel metal2 576 -203 576 -203 0 net=6894
rlabel metal2 653 -205 653 -205 0 net=6015
rlabel metal2 653 -207 653 -207 0 net=6896
rlabel metal2 656 -209 656 -209 0 net=6033
rlabel metal2 16 -220 16 -220 0 net=5621
rlabel metal2 723 -220 723 -220 0 net=5784
rlabel metal2 1108 -220 1108 -220 0 net=6771
rlabel metal2 1108 -220 1108 -220 0 net=6771
rlabel metal2 23 -222 23 -222 0 net=1768
rlabel metal2 261 -222 261 -222 0 net=3009
rlabel metal2 352 -222 352 -222 0 net=4736
rlabel metal2 401 -222 401 -222 0 net=6558
rlabel metal2 887 -222 887 -222 0 net=7204
rlabel metal2 23 -224 23 -224 0 net=3639
rlabel metal2 114 -224 114 -224 0 net=1293
rlabel metal2 254 -224 254 -224 0 net=1329
rlabel metal2 471 -224 471 -224 0 net=4013
rlabel metal2 495 -224 495 -224 0 net=7298
rlabel metal2 30 -226 30 -226 0 net=2450
rlabel metal2 366 -226 366 -226 0 net=3016
rlabel metal2 502 -226 502 -226 0 net=4522
rlabel metal2 579 -226 579 -226 0 net=7402
rlabel metal2 30 -228 30 -228 0 net=5189
rlabel metal2 163 -228 163 -228 0 net=1460
rlabel metal2 296 -228 296 -228 0 net=1113
rlabel metal2 555 -228 555 -228 0 net=4947
rlabel metal2 618 -228 618 -228 0 net=6936
rlabel metal2 44 -230 44 -230 0 net=1824
rlabel metal2 142 -230 142 -230 0 net=4510
rlabel metal2 604 -230 604 -230 0 net=4915
rlabel metal2 604 -230 604 -230 0 net=4915
rlabel metal2 611 -230 611 -230 0 net=5283
rlabel metal2 674 -230 674 -230 0 net=3636
rlabel metal2 51 -232 51 -232 0 net=2230
rlabel metal2 299 -232 299 -232 0 net=612
rlabel metal2 621 -232 621 -232 0 net=7098
rlabel metal2 51 -234 51 -234 0 net=3293
rlabel metal2 65 -234 65 -234 0 net=3769
rlabel metal2 299 -234 299 -234 0 net=3580
rlabel metal2 618 -234 618 -234 0 net=5193
rlabel metal2 58 -236 58 -236 0 net=3581
rlabel metal2 625 -236 625 -236 0 net=5237
rlabel metal2 663 -236 663 -236 0 net=5285
rlabel metal2 674 -236 674 -236 0 net=5497
rlabel metal2 702 -236 702 -236 0 net=6181
rlabel metal2 807 -236 807 -236 0 net=6035
rlabel metal2 65 -238 65 -238 0 net=2701
rlabel metal2 121 -238 121 -238 0 net=4542
rlabel metal2 628 -238 628 -238 0 net=7406
rlabel metal2 68 -240 68 -240 0 net=4133
rlabel metal2 408 -240 408 -240 0 net=3945
rlabel metal2 541 -240 541 -240 0 net=4453
rlabel metal2 639 -240 639 -240 0 net=5103
rlabel metal2 72 -242 72 -242 0 net=1842
rlabel metal2 317 -242 317 -242 0 net=3867
rlabel metal2 541 -242 541 -242 0 net=4515
rlabel metal2 597 -242 597 -242 0 net=4897
rlabel metal2 646 -242 646 -242 0 net=5139
rlabel metal2 646 -242 646 -242 0 net=5139
rlabel metal2 653 -242 653 -242 0 net=7582
rlabel metal2 72 -244 72 -244 0 net=2347
rlabel metal2 359 -244 359 -244 0 net=5016
rlabel metal2 527 -244 527 -244 0 net=4341
rlabel metal2 597 -244 597 -244 0 net=5705
rlabel metal2 723 -244 723 -244 0 net=5855
rlabel metal2 737 -244 737 -244 0 net=6017
rlabel metal2 800 -244 800 -244 0 net=6389
rlabel metal2 828 -244 828 -244 0 net=7327
rlabel metal2 79 -246 79 -246 0 net=4061
rlabel metal2 121 -246 121 -246 0 net=1500
rlabel metal2 177 -246 177 -246 0 net=1212
rlabel metal2 289 -246 289 -246 0 net=2255
rlabel metal2 317 -246 317 -246 0 net=4759
rlabel metal2 653 -246 653 -246 0 net=5767
rlabel metal2 730 -246 730 -246 0 net=6161
rlabel metal2 93 -248 93 -248 0 net=1249
rlabel metal2 324 -248 324 -248 0 net=4768
rlabel metal2 100 -250 100 -250 0 net=2017
rlabel metal2 170 -250 170 -250 0 net=6870
rlabel metal2 100 -252 100 -252 0 net=996
rlabel metal2 173 -252 173 -252 0 net=1895
rlabel metal2 324 -252 324 -252 0 net=3193
rlabel metal2 688 -252 688 -252 0 net=6497
rlabel metal2 814 -252 814 -252 0 net=6523
rlabel metal2 856 -252 856 -252 0 net=7585
rlabel metal2 117 -254 117 -254 0 net=2733
rlabel metal2 177 -254 177 -254 0 net=1715
rlabel metal2 194 -254 194 -254 0 net=4314
rlabel metal2 695 -254 695 -254 0 net=5573
rlabel metal2 814 -254 814 -254 0 net=6577
rlabel metal2 919 -254 919 -254 0 net=6829
rlabel metal2 93 -256 93 -256 0 net=3207
rlabel metal2 198 -256 198 -256 0 net=1861
rlabel metal2 240 -256 240 -256 0 net=5885
rlabel metal2 709 -256 709 -256 0 net=6081
rlabel metal2 37 -258 37 -258 0 net=1305
rlabel metal2 331 -258 331 -258 0 net=3852
rlabel metal2 485 -258 485 -258 0 net=6193
rlabel metal2 37 -260 37 -260 0 net=2651
rlabel metal2 331 -260 331 -260 0 net=4585
rlabel metal2 740 -260 740 -260 0 net=6429
rlabel metal2 47 -262 47 -262 0 net=2493
rlabel metal2 205 -262 205 -262 0 net=818
rlabel metal2 205 -262 205 -262 0 net=818
rlabel metal2 219 -262 219 -262 0 net=2945
rlabel metal2 485 -262 485 -262 0 net=7544
rlabel metal2 135 -264 135 -264 0 net=3666
rlabel metal2 219 -264 219 -264 0 net=1643
rlabel metal2 247 -264 247 -264 0 net=2763
rlabel metal2 338 -264 338 -264 0 net=3155
rlabel metal2 397 -264 397 -264 0 net=7413
rlabel metal2 86 -266 86 -266 0 net=2503
rlabel metal2 142 -266 142 -266 0 net=1825
rlabel metal2 282 -266 282 -266 0 net=3331
rlabel metal2 436 -266 436 -266 0 net=3968
rlabel metal2 128 -268 128 -268 0 net=3799
rlabel metal2 282 -268 282 -268 0 net=3443
rlabel metal2 362 -268 362 -268 0 net=4810
rlabel metal2 744 -268 744 -268 0 net=6105
rlabel metal2 191 -270 191 -270 0 net=1695
rlabel metal2 450 -270 450 -270 0 net=4415
rlabel metal2 583 -270 583 -270 0 net=6991
rlabel metal2 191 -272 191 -272 0 net=5428
rlabel metal2 443 -272 443 -272 0 net=4969
rlabel metal2 590 -272 590 -272 0 net=5079
rlabel metal2 751 -272 751 -272 0 net=6531
rlabel metal2 334 -274 334 -274 0 net=5367
rlabel metal2 488 -274 488 -274 0 net=6845
rlabel metal2 758 -274 758 -274 0 net=6297
rlabel metal2 821 -274 821 -274 0 net=6947
rlabel metal2 415 -276 415 -276 0 net=3571
rlabel metal2 506 -276 506 -276 0 net=4431
rlabel metal2 632 -276 632 -276 0 net=5459
rlabel metal2 793 -276 793 -276 0 net=7027
rlabel metal2 152 -278 152 -278 0 net=4403
rlabel metal2 842 -278 842 -278 0 net=7069
rlabel metal2 257 -280 257 -280 0 net=5639
rlabel metal2 870 -280 870 -280 0 net=7505
rlabel metal2 310 -282 310 -282 0 net=3163
rlabel metal2 422 -282 422 -282 0 net=3341
rlabel metal2 576 -282 576 -282 0 net=7549
rlabel metal2 310 -284 310 -284 0 net=2729
rlabel metal2 373 -286 373 -286 0 net=3071
rlabel metal2 457 -286 457 -286 0 net=5599
rlabel metal2 373 -288 373 -288 0 net=5809
rlabel metal2 457 -290 457 -290 0 net=4077
rlabel metal2 499 -292 499 -292 0 net=5007
rlabel metal2 16 -303 16 -303 0 net=5622
rlabel metal2 240 -303 240 -303 0 net=1306
rlabel metal2 492 -303 492 -303 0 net=4015
rlabel metal2 523 -303 523 -303 0 net=7586
rlabel metal2 863 -303 863 -303 0 net=6037
rlabel metal2 1108 -303 1108 -303 0 net=6773
rlabel metal2 1108 -303 1108 -303 0 net=6773
rlabel metal2 23 -305 23 -305 0 net=3640
rlabel metal2 110 -305 110 -305 0 net=182
rlabel metal2 124 -305 124 -305 0 net=431
rlabel metal2 159 -305 159 -305 0 net=1005
rlabel metal2 254 -305 254 -305 0 net=1330
rlabel metal2 394 -305 394 -305 0 net=384
rlabel metal2 898 -305 898 -305 0 net=5105
rlabel metal2 23 -307 23 -307 0 net=3493
rlabel metal2 233 -307 233 -307 0 net=1295
rlabel metal2 247 -307 247 -307 0 net=2764
rlabel metal2 352 -307 352 -307 0 net=919
rlabel metal2 544 -307 544 -307 0 net=5768
rlabel metal2 660 -307 660 -307 0 net=6107
rlabel metal2 800 -307 800 -307 0 net=5574
rlabel metal2 30 -309 30 -309 0 net=5191
rlabel metal2 355 -309 355 -309 0 net=4432
rlabel metal2 516 -309 516 -309 0 net=6119
rlabel metal2 835 -309 835 -309 0 net=7414
rlabel metal2 37 -311 37 -311 0 net=2652
rlabel metal2 100 -311 100 -311 0 net=2495
rlabel metal2 233 -311 233 -311 0 net=2145
rlabel metal2 681 -311 681 -311 0 net=5641
rlabel metal2 37 -313 37 -313 0 net=2291
rlabel metal2 306 -313 306 -313 0 net=6245
rlabel metal2 807 -313 807 -313 0 net=6391
rlabel metal2 863 -313 863 -313 0 net=7507
rlabel metal2 877 -313 877 -313 0 net=7551
rlabel metal2 44 -315 44 -315 0 net=2141
rlabel metal2 117 -315 117 -315 0 net=2018
rlabel metal2 170 -315 170 -315 0 net=4516
rlabel metal2 625 -315 625 -315 0 net=5239
rlabel metal2 786 -315 786 -315 0 net=6993
rlabel metal2 877 -315 877 -315 0 net=6830
rlabel metal2 47 -317 47 -317 0 net=4948
rlabel metal2 646 -317 646 -317 0 net=5141
rlabel metal2 716 -317 716 -317 0 net=6847
rlabel metal2 793 -317 793 -317 0 net=7029
rlabel metal2 58 -319 58 -319 0 net=3582
rlabel metal2 422 -319 422 -319 0 net=3072
rlabel metal2 541 -319 541 -319 0 net=5856
rlabel metal2 730 -319 730 -319 0 net=6163
rlabel metal2 58 -321 58 -321 0 net=2505
rlabel metal2 128 -321 128 -321 0 net=1133
rlabel metal2 149 -321 149 -321 0 net=2735
rlabel metal2 261 -321 261 -321 0 net=3770
rlabel metal2 261 -321 261 -321 0 net=3770
rlabel metal2 268 -321 268 -321 0 net=3801
rlabel metal2 576 -321 576 -321 0 net=5601
rlabel metal2 65 -323 65 -323 0 net=827
rlabel metal2 439 -323 439 -323 0 net=6018
rlabel metal2 9 -325 9 -325 0 net=2491
rlabel metal2 68 -325 68 -325 0 net=6532
rlabel metal2 68 -327 68 -327 0 net=3937
rlabel metal2 128 -327 128 -327 0 net=2609
rlabel metal2 173 -327 173 -327 0 net=4898
rlabel metal2 702 -327 702 -327 0 net=6183
rlabel metal2 79 -329 79 -329 0 net=4062
rlabel metal2 135 -329 135 -329 0 net=5613
rlabel metal2 79 -331 79 -331 0 net=6524
rlabel metal2 82 -333 82 -333 0 net=2765
rlabel metal2 527 -333 527 -333 0 net=4417
rlabel metal2 597 -333 597 -333 0 net=5707
rlabel metal2 842 -333 842 -333 0 net=7071
rlabel metal2 149 -335 149 -335 0 net=1645
rlabel metal2 268 -335 268 -335 0 net=1251
rlabel metal2 296 -335 296 -335 0 net=3572
rlabel metal2 464 -335 464 -335 0 net=6194
rlabel metal2 16 -337 16 -337 0 net=1507
rlabel metal2 275 -337 275 -337 0 net=2033
rlabel metal2 513 -337 513 -337 0 net=4405
rlabel metal2 583 -337 583 -337 0 net=4971
rlabel metal2 618 -337 618 -337 0 net=5195
rlabel metal2 674 -337 674 -337 0 net=5499
rlabel metal2 709 -337 709 -337 0 net=6083
rlabel metal2 772 -337 772 -337 0 net=6431
rlabel metal2 163 -339 163 -339 0 net=4889
rlabel metal2 191 -339 191 -339 0 net=2907
rlabel metal2 404 -339 404 -339 0 net=4777
rlabel metal2 667 -339 667 -339 0 net=5287
rlabel metal2 688 -339 688 -339 0 net=6499
rlabel metal2 170 -341 170 -341 0 net=1253
rlabel metal2 205 -341 205 -341 0 net=4251
rlabel metal2 709 -341 709 -341 0 net=5343
rlabel metal2 173 -343 173 -343 0 net=4586
rlabel metal2 345 -343 345 -343 0 net=3011
rlabel metal2 779 -343 779 -343 0 net=7329
rlabel metal2 72 -345 72 -345 0 net=2349
rlabel metal2 359 -345 359 -345 0 net=702
rlabel metal2 814 -345 814 -345 0 net=6579
rlabel metal2 72 -347 72 -347 0 net=2875
rlabel metal2 177 -347 177 -347 0 net=1717
rlabel metal2 177 -347 177 -347 0 net=1717
rlabel metal2 205 -347 205 -347 0 net=1361
rlabel metal2 289 -347 289 -347 0 net=1897
rlabel metal2 310 -347 310 -347 0 net=2731
rlabel metal2 408 -347 408 -347 0 net=3947
rlabel metal2 513 -347 513 -347 0 net=5080
rlabel metal2 814 -347 814 -347 0 net=6949
rlabel metal2 194 -349 194 -349 0 net=6309
rlabel metal2 226 -351 226 -351 0 net=1863
rlabel metal2 310 -351 310 -351 0 net=3165
rlabel metal2 443 -351 443 -351 0 net=5887
rlabel metal2 212 -353 212 -353 0 net=1697
rlabel metal2 247 -353 247 -353 0 net=2767
rlabel metal2 450 -353 450 -353 0 net=3343
rlabel metal2 471 -353 471 -353 0 net=3869
rlabel metal2 257 -355 257 -355 0 net=3485
rlabel metal2 562 -355 562 -355 0 net=4455
rlabel metal2 632 -355 632 -355 0 net=5461
rlabel metal2 264 -357 264 -357 0 net=3245
rlabel metal2 604 -357 604 -357 0 net=4917
rlabel metal2 282 -359 282 -359 0 net=3445
rlabel metal2 142 -361 142 -361 0 net=1827
rlabel metal2 317 -361 317 -361 0 net=5284
rlabel metal2 107 -363 107 -363 0 net=2703
rlabel metal2 320 -363 320 -363 0 net=2889
rlabel metal2 429 -363 429 -363 0 net=5369
rlabel metal2 107 -365 107 -365 0 net=6911
rlabel metal2 324 -367 324 -367 0 net=3195
rlabel metal2 534 -367 534 -367 0 net=4761
rlabel metal2 324 -369 324 -369 0 net=5810
rlabel metal2 331 -371 331 -371 0 net=2271
rlabel metal2 341 -373 341 -373 0 net=3771
rlabel metal2 366 -373 366 -373 0 net=4135
rlabel metal2 758 -373 758 -373 0 net=6299
rlabel metal2 303 -375 303 -375 0 net=2257
rlabel metal2 373 -375 373 -375 0 net=4078
rlabel metal2 534 -375 534 -375 0 net=5009
rlabel metal2 51 -377 51 -377 0 net=3294
rlabel metal2 338 -377 338 -377 0 net=3157
rlabel metal2 548 -377 548 -377 0 net=4343
rlabel metal2 51 -379 51 -379 0 net=3209
rlabel metal2 380 -379 380 -379 0 net=3333
rlabel metal2 436 -381 436 -381 0 net=5439
rlabel metal2 397 -383 397 -383 0 net=2747
rlabel metal2 397 -385 397 -385 0 net=2946
rlabel metal2 166 -387 166 -387 0 net=4141
rlabel metal2 2 -398 2 -398 0 net=4707
rlabel metal2 611 -398 611 -398 0 net=4763
rlabel metal2 1108 -398 1108 -398 0 net=6775
rlabel metal2 9 -400 9 -400 0 net=2492
rlabel metal2 44 -400 44 -400 0 net=2142
rlabel metal2 145 -400 145 -400 0 net=5888
rlabel metal2 464 -400 464 -400 0 net=3345
rlabel metal2 464 -400 464 -400 0 net=3345
rlabel metal2 474 -400 474 -400 0 net=6500
rlabel metal2 849 -400 849 -400 0 net=7073
rlabel metal2 982 -400 982 -400 0 net=7463
rlabel metal2 16 -402 16 -402 0 net=2497
rlabel metal2 107 -402 107 -402 0 net=2273
rlabel metal2 338 -402 338 -402 0 net=2259
rlabel metal2 380 -402 380 -402 0 net=3603
rlabel metal2 569 -402 569 -402 0 net=4345
rlabel metal2 628 -402 628 -402 0 net=6994
rlabel metal2 884 -402 884 -402 0 net=5106
rlabel metal2 905 -402 905 -402 0 net=6039
rlabel metal2 905 -402 905 -402 0 net=6039
rlabel metal2 933 -402 933 -402 0 net=5643
rlabel metal2 23 -404 23 -404 0 net=3494
rlabel metal2 170 -404 170 -404 0 net=6246
rlabel metal2 807 -404 807 -404 0 net=7031
rlabel metal2 989 -404 989 -404 0 net=7177
rlabel metal2 23 -406 23 -406 0 net=3211
rlabel metal2 58 -406 58 -406 0 net=2507
rlabel metal2 380 -406 380 -406 0 net=2766
rlabel metal2 569 -406 569 -406 0 net=6310
rlabel metal2 828 -406 828 -406 0 net=6581
rlabel metal2 37 -408 37 -408 0 net=2293
rlabel metal2 341 -408 341 -408 0 net=2908
rlabel metal2 422 -408 422 -408 0 net=2891
rlabel metal2 474 -408 474 -408 0 net=7629
rlabel metal2 44 -410 44 -410 0 net=2035
rlabel metal2 296 -410 296 -410 0 net=1899
rlabel metal2 306 -410 306 -410 0 net=4661
rlabel metal2 863 -410 863 -410 0 net=7509
rlabel metal2 51 -412 51 -412 0 net=3167
rlabel metal2 327 -412 327 -412 0 net=3012
rlabel metal2 702 -412 702 -412 0 net=5501
rlabel metal2 835 -412 835 -412 0 net=6393
rlabel metal2 891 -412 891 -412 0 net=7553
rlabel metal2 65 -414 65 -414 0 net=4252
rlabel metal2 625 -414 625 -414 0 net=7175
rlabel metal2 79 -416 79 -416 0 net=5192
rlabel metal2 383 -416 383 -416 0 net=3334
rlabel metal2 572 -416 572 -416 0 net=7035
rlabel metal2 79 -418 79 -418 0 net=2611
rlabel metal2 135 -418 135 -418 0 net=4017
rlabel metal2 576 -418 576 -418 0 net=4419
rlabel metal2 635 -418 635 -418 0 net=6164
rlabel metal2 814 -418 814 -418 0 net=6951
rlabel metal2 82 -420 82 -420 0 net=4903
rlabel metal2 709 -420 709 -420 0 net=5345
rlabel metal2 96 -422 96 -422 0 net=4929
rlabel metal2 100 -424 100 -424 0 net=2055
rlabel metal2 478 -424 478 -424 0 net=4143
rlabel metal2 632 -424 632 -424 0 net=4919
rlabel metal2 723 -424 723 -424 0 net=5615
rlabel metal2 114 -426 114 -426 0 net=3583
rlabel metal2 485 -426 485 -426 0 net=3949
rlabel metal2 576 -426 576 -426 0 net=5935
rlabel metal2 117 -428 117 -428 0 net=6912
rlabel metal2 121 -430 121 -430 0 net=2732
rlabel metal2 397 -430 397 -430 0 net=3870
rlabel metal2 667 -430 667 -430 0 net=6069
rlabel metal2 86 -432 86 -432 0 net=3939
rlabel metal2 401 -432 401 -432 0 net=3803
rlabel metal2 506 -432 506 -432 0 net=3467
rlabel metal2 590 -432 590 -432 0 net=4457
rlabel metal2 667 -432 667 -432 0 net=6185
rlabel metal2 765 -432 765 -432 0 net=6301
rlabel metal2 72 -434 72 -434 0 net=2877
rlabel metal2 121 -434 121 -434 0 net=4890
rlabel metal2 170 -434 170 -434 0 net=1503
rlabel metal2 264 -434 264 -434 0 net=3246
rlabel metal2 590 -434 590 -434 0 net=5371
rlabel metal2 681 -434 681 -434 0 net=5143
rlabel metal2 772 -434 772 -434 0 net=6433
rlabel metal2 72 -436 72 -436 0 net=3001
rlabel metal2 149 -436 149 -436 0 net=1647
rlabel metal2 184 -436 184 -436 0 net=4778
rlabel metal2 639 -436 639 -436 0 net=5197
rlabel metal2 786 -436 786 -436 0 net=6849
rlabel metal2 61 -438 61 -438 0 net=4241
rlabel metal2 653 -438 653 -438 0 net=5241
rlabel metal2 149 -440 149 -440 0 net=2287
rlabel metal2 408 -440 408 -440 0 net=3487
rlabel metal2 534 -440 534 -440 0 net=5011
rlabel metal2 688 -440 688 -440 0 net=6401
rlabel metal2 12 -442 12 -442 0 net=3915
rlabel metal2 429 -442 429 -442 0 net=3197
rlabel metal2 492 -442 492 -442 0 net=6561
rlabel metal2 156 -444 156 -444 0 net=1719
rlabel metal2 184 -444 184 -444 0 net=1255
rlabel metal2 198 -444 198 -444 0 net=2737
rlabel metal2 268 -444 268 -444 0 net=1252
rlabel metal2 327 -444 327 -444 0 net=3158
rlabel metal2 460 -444 460 -444 0 net=4279
rlabel metal2 177 -446 177 -446 0 net=2679
rlabel metal2 219 -446 219 -446 0 net=1509
rlabel metal2 352 -446 352 -446 0 net=7471
rlabel metal2 180 -448 180 -448 0 net=3295
rlabel metal2 233 -448 233 -448 0 net=2147
rlabel metal2 373 -448 373 -448 0 net=4407
rlabel metal2 534 -448 534 -448 0 net=6108
rlabel metal2 716 -448 716 -448 0 net=5603
rlabel metal2 730 -448 730 -448 0 net=5709
rlabel metal2 187 -450 187 -450 0 net=2768
rlabel metal2 425 -450 425 -450 0 net=4837
rlabel metal2 695 -450 695 -450 0 net=5463
rlabel metal2 737 -450 737 -450 0 net=6085
rlabel metal2 191 -452 191 -452 0 net=1229
rlabel metal2 198 -454 198 -454 0 net=1698
rlabel metal2 233 -454 233 -454 0 net=1235
rlabel metal2 429 -454 429 -454 0 net=2749
rlabel metal2 450 -454 450 -454 0 net=3447
rlabel metal2 597 -454 597 -454 0 net=4973
rlabel metal2 744 -454 744 -454 0 net=6121
rlabel metal2 205 -456 205 -456 0 net=1363
rlabel metal2 247 -456 247 -456 0 net=1741
rlabel metal2 275 -456 275 -456 0 net=1663
rlabel metal2 516 -456 516 -456 0 net=5061
rlabel metal2 758 -456 758 -456 0 net=5441
rlabel metal2 93 -458 93 -458 0 net=292
rlabel metal2 240 -458 240 -458 0 net=1297
rlabel metal2 250 -458 250 -458 0 net=1864
rlabel metal2 317 -458 317 -458 0 net=3481
rlabel metal2 457 -458 457 -458 0 net=6645
rlabel metal2 93 -460 93 -460 0 net=2417
rlabel metal2 142 -460 142 -460 0 net=2705
rlabel metal2 254 -460 254 -460 0 net=109
rlabel metal2 68 -462 68 -462 0 net=4387
rlabel metal2 282 -462 282 -462 0 net=1828
rlabel metal2 481 -462 481 -462 0 net=4567
rlabel metal2 674 -462 674 -462 0 net=5289
rlabel metal2 110 -464 110 -464 0 net=4737
rlabel metal2 359 -464 359 -464 0 net=3773
rlabel metal2 495 -464 495 -464 0 net=4993
rlabel metal2 142 -466 142 -466 0 net=4931
rlabel metal2 695 -466 695 -466 0 net=7331
rlabel metal2 173 -468 173 -468 0 net=1675
rlabel metal2 345 -468 345 -468 0 net=2351
rlabel metal2 499 -468 499 -468 0 net=5201
rlabel metal2 30 -470 30 -470 0 net=2985
rlabel metal2 541 -470 541 -470 0 net=4663
rlabel metal2 324 -472 324 -472 0 net=3619
rlabel metal2 544 -472 544 -472 0 net=5117
rlabel metal2 37 -474 37 -474 0 net=2511
rlabel metal2 555 -474 555 -474 0 net=4137
rlabel metal2 492 -476 492 -476 0 net=3335
rlabel metal2 9 -487 9 -487 0 net=7675
rlabel metal2 646 -487 646 -487 0 net=4459
rlabel metal2 646 -487 646 -487 0 net=4459
rlabel metal2 814 -487 814 -487 0 net=7359
rlabel metal2 1111 -487 1111 -487 0 net=4325
rlabel metal2 30 -489 30 -489 0 net=2986
rlabel metal2 44 -489 44 -489 0 net=2036
rlabel metal2 285 -489 285 -489 0 net=4242
rlabel metal2 765 -489 765 -489 0 net=5145
rlabel metal2 817 -489 817 -489 0 net=6122
rlabel metal2 954 -489 954 -489 0 net=7033
rlabel metal2 1115 -489 1115 -489 0 net=6777
rlabel metal2 23 -491 23 -491 0 net=3213
rlabel metal2 772 -491 772 -491 0 net=5199
rlabel metal2 975 -491 975 -491 0 net=7075
rlabel metal2 30 -493 30 -493 0 net=2681
rlabel metal2 296 -493 296 -493 0 net=1510
rlabel metal2 373 -493 373 -493 0 net=4408
rlabel metal2 555 -493 555 -493 0 net=6434
rlabel metal2 1010 -493 1010 -493 0 net=7511
rlabel metal2 296 -495 296 -495 0 net=2149
rlabel metal2 317 -495 317 -495 0 net=4739
rlabel metal2 37 -497 37 -497 0 net=2513
rlabel metal2 310 -497 310 -497 0 net=3337
rlabel metal2 499 -497 499 -497 0 net=2901
rlabel metal2 565 -497 565 -497 0 net=6086
rlabel metal2 1017 -497 1017 -497 0 net=7555
rlabel metal2 44 -499 44 -499 0 net=3805
rlabel metal2 415 -499 415 -499 0 net=4049
rlabel metal2 842 -499 842 -499 0 net=5617
rlabel metal2 1024 -499 1024 -499 0 net=7631
rlabel metal2 16 -501 16 -501 0 net=2499
rlabel metal2 422 -501 422 -501 0 net=5012
rlabel metal2 709 -501 709 -501 0 net=4921
rlabel metal2 863 -501 863 -501 0 net=6395
rlabel metal2 1045 -501 1045 -501 0 net=5645
rlabel metal2 16 -503 16 -503 0 net=2199
rlabel metal2 359 -503 359 -503 0 net=2353
rlabel metal2 397 -503 397 -503 0 net=4662
rlabel metal2 926 -503 926 -503 0 net=6583
rlabel metal2 982 -503 982 -503 0 net=7465
rlabel metal2 58 -505 58 -505 0 net=3003
rlabel metal2 79 -505 79 -505 0 net=2612
rlabel metal2 149 -505 149 -505 0 net=2289
rlabel metal2 401 -505 401 -505 0 net=2869
rlabel metal2 425 -505 425 -505 0 net=4764
rlabel metal2 61 -507 61 -507 0 net=2053
rlabel metal2 695 -507 695 -507 0 net=7333
rlabel metal2 940 -507 940 -507 0 net=6647
rlabel metal2 26 -509 26 -509 0 net=6341
rlabel metal2 65 -511 65 -511 0 net=1901
rlabel metal2 327 -511 327 -511 0 net=2553
rlabel metal2 443 -511 443 -511 0 net=2893
rlabel metal2 481 -511 481 -511 0 net=4138
rlabel metal2 800 -511 800 -511 0 net=5347
rlabel metal2 891 -511 891 -511 0 net=6953
rlabel metal2 72 -513 72 -513 0 net=4145
rlabel metal2 597 -513 597 -513 0 net=5203
rlabel metal2 856 -513 856 -513 0 net=6071
rlabel metal2 919 -513 919 -513 0 net=6563
rlabel metal2 79 -515 79 -515 0 net=2419
rlabel metal2 96 -515 96 -515 0 net=2706
rlabel metal2 261 -515 261 -515 0 net=2739
rlabel metal2 338 -515 338 -515 0 net=2260
rlabel metal2 464 -515 464 -515 0 net=3346
rlabel metal2 474 -515 474 -515 0 net=5372
rlabel metal2 597 -515 597 -515 0 net=5502
rlabel metal2 877 -515 877 -515 0 net=5443
rlabel metal2 51 -517 51 -517 0 net=3168
rlabel metal2 485 -517 485 -517 0 net=3199
rlabel metal2 502 -517 502 -517 0 net=5464
rlabel metal2 758 -517 758 -517 0 net=5119
rlabel metal2 51 -519 51 -519 0 net=2295
rlabel metal2 341 -519 341 -519 0 net=486
rlabel metal2 712 -519 712 -519 0 net=5465
rlabel metal2 100 -521 100 -521 0 net=2057
rlabel metal2 383 -521 383 -521 0 net=5511
rlabel metal2 2 -523 2 -523 0 net=4708
rlabel metal2 114 -523 114 -523 0 net=3585
rlabel metal2 436 -523 436 -523 0 net=3483
rlabel metal2 506 -523 506 -523 0 net=3469
rlabel metal2 600 -523 600 -523 0 net=6409
rlabel metal2 114 -525 114 -525 0 net=4297
rlabel metal2 261 -525 261 -525 0 net=1743
rlabel metal2 271 -525 271 -525 0 net=4933
rlabel metal2 121 -527 121 -527 0 net=1535
rlabel metal2 569 -527 569 -527 0 net=2943
rlabel metal2 716 -527 716 -527 0 net=4975
rlabel metal2 128 -529 128 -529 0 net=3940
rlabel metal2 457 -529 457 -529 0 net=5710
rlabel metal2 107 -531 107 -531 0 net=2275
rlabel metal2 429 -531 429 -531 0 net=2751
rlabel metal2 506 -531 506 -531 0 net=4839
rlabel metal2 758 -531 758 -531 0 net=5937
rlabel metal2 107 -533 107 -533 0 net=4930
rlabel metal2 128 -535 128 -535 0 net=4477
rlabel metal2 303 -535 303 -535 0 net=2025
rlabel metal2 523 -535 523 -535 0 net=6302
rlabel metal2 135 -537 135 -537 0 net=4019
rlabel metal2 534 -537 534 -537 0 net=784
rlabel metal2 723 -537 723 -537 0 net=5605
rlabel metal2 135 -539 135 -539 0 net=4388
rlabel metal2 324 -539 324 -539 0 net=5625
rlabel metal2 142 -541 142 -541 0 net=1665
rlabel metal2 324 -541 324 -541 0 net=3775
rlabel metal2 534 -541 534 -541 0 net=4205
rlabel metal2 723 -541 723 -541 0 net=5243
rlabel metal2 145 -543 145 -543 0 net=1685
rlabel metal2 247 -543 247 -543 0 net=1299
rlabel metal2 275 -543 275 -543 0 net=1677
rlabel metal2 331 -543 331 -543 0 net=3231
rlabel metal2 688 -543 688 -543 0 net=5051
rlabel metal2 138 -545 138 -545 0 net=1559
rlabel metal2 345 -545 345 -545 0 net=4932
rlabel metal2 744 -545 744 -545 0 net=5291
rlabel metal2 149 -547 149 -547 0 net=1237
rlabel metal2 247 -547 247 -547 0 net=1285
rlabel metal2 348 -547 348 -547 0 net=4664
rlabel metal2 681 -547 681 -547 0 net=7176
rlabel metal2 86 -549 86 -549 0 net=2879
rlabel metal2 348 -549 348 -549 0 net=3175
rlabel metal2 450 -549 450 -549 0 net=2613
rlabel metal2 527 -549 527 -549 0 net=3449
rlabel metal2 702 -549 702 -549 0 net=4905
rlabel metal2 751 -549 751 -549 0 net=4281
rlabel metal2 86 -551 86 -551 0 net=1505
rlabel metal2 180 -551 180 -551 0 net=1364
rlabel metal2 366 -551 366 -551 0 net=2509
rlabel metal2 93 -553 93 -553 0 net=6279
rlabel metal2 156 -555 156 -555 0 net=1721
rlabel metal2 527 -555 527 -555 0 net=4079
rlabel metal2 611 -555 611 -555 0 net=4347
rlabel metal2 156 -557 156 -557 0 net=1793
rlabel metal2 537 -557 537 -557 0 net=5575
rlabel metal2 163 -559 163 -559 0 net=1649
rlabel metal2 191 -559 191 -559 0 net=1231
rlabel metal2 537 -559 537 -559 0 net=6186
rlabel metal2 163 -561 163 -561 0 net=2545
rlabel metal2 541 -561 541 -561 0 net=3621
rlabel metal2 166 -563 166 -563 0 net=7285
rlabel metal2 184 -565 184 -565 0 net=1257
rlabel metal2 198 -565 198 -565 0 net=7623
rlabel metal2 184 -567 184 -567 0 net=3297
rlabel metal2 513 -567 513 -567 0 net=3605
rlabel metal2 555 -567 555 -567 0 net=3373
rlabel metal2 572 -567 572 -567 0 net=4994
rlabel metal2 198 -569 198 -569 0 net=1373
rlabel metal2 219 -569 219 -569 0 net=2251
rlabel metal2 625 -569 625 -569 0 net=4421
rlabel metal2 737 -569 737 -569 0 net=5063
rlabel metal2 408 -571 408 -571 0 net=3917
rlabel metal2 408 -573 408 -573 0 net=3381
rlabel metal2 579 -573 579 -573 0 net=6187
rlabel metal2 513 -575 513 -575 0 net=3489
rlabel metal2 562 -575 562 -575 0 net=7429
rlabel metal2 625 -577 625 -577 0 net=4569
rlabel metal2 548 -579 548 -579 0 net=3951
rlabel metal2 548 -581 548 -581 0 net=7472
rlabel metal2 635 -583 635 -583 0 net=4769
rlabel metal2 989 -583 989 -583 0 net=7179
rlabel metal2 642 -585 642 -585 0 net=4159
rlabel metal2 961 -585 961 -585 0 net=7037
rlabel metal2 905 -587 905 -587 0 net=6041
rlabel metal2 905 -589 905 -589 0 net=6851
rlabel metal2 870 -591 870 -591 0 net=6403
rlabel metal2 572 -593 572 -593 0 net=6023
rlabel metal2 2 -604 2 -604 0 net=2880
rlabel metal2 240 -604 240 -604 0 net=1687
rlabel metal2 240 -604 240 -604 0 net=1687
rlabel metal2 254 -604 254 -604 0 net=1300
rlabel metal2 289 -604 289 -604 0 net=1560
rlabel metal2 544 -604 544 -604 0 net=6648
rlabel metal2 1111 -604 1111 -604 0 net=4657
rlabel metal2 2 -606 2 -606 0 net=5875
rlabel metal2 121 -606 121 -606 0 net=1537
rlabel metal2 303 -606 303 -606 0 net=2027
rlabel metal2 303 -606 303 -606 0 net=2027
rlabel metal2 310 -606 310 -606 0 net=3338
rlabel metal2 534 -606 534 -606 0 net=4461
rlabel metal2 684 -606 684 -606 0 net=7076
rlabel metal2 1115 -606 1115 -606 0 net=5647
rlabel metal2 5 -608 5 -608 0 net=7059
rlabel metal2 548 -608 548 -608 0 net=5606
rlabel metal2 989 -608 989 -608 0 net=7039
rlabel metal2 1101 -608 1101 -608 0 net=7709
rlabel metal2 1122 -608 1122 -608 0 net=4327
rlabel metal2 1122 -608 1122 -608 0 net=4327
rlabel metal2 1129 -608 1129 -608 0 net=6779
rlabel metal2 9 -610 9 -610 0 net=7676
rlabel metal2 338 -610 338 -610 0 net=3622
rlabel metal2 779 -610 779 -610 0 net=4935
rlabel metal2 779 -610 779 -610 0 net=4935
rlabel metal2 793 -610 793 -610 0 net=5065
rlabel metal2 793 -610 793 -610 0 net=5065
rlabel metal2 898 -610 898 -610 0 net=7467
rlabel metal2 1094 -610 1094 -610 0 net=7633
rlabel metal2 1129 -610 1129 -610 0 net=5951
rlabel metal2 16 -612 16 -612 0 net=2200
rlabel metal2 362 -612 362 -612 0 net=810
rlabel metal2 579 -612 579 -612 0 net=7034
rlabel metal2 1066 -612 1066 -612 0 net=7557
rlabel metal2 16 -614 16 -614 0 net=1903
rlabel metal2 72 -614 72 -614 0 net=4146
rlabel metal2 541 -614 541 -614 0 net=3607
rlabel metal2 604 -614 604 -614 0 net=2944
rlabel metal2 23 -616 23 -616 0 net=4479
rlabel metal2 135 -616 135 -616 0 net=1623
rlabel metal2 338 -616 338 -616 0 net=2753
rlabel metal2 460 -616 460 -616 0 net=5204
rlabel metal2 926 -616 926 -616 0 net=7335
rlabel metal2 26 -618 26 -618 0 net=3004
rlabel metal2 65 -618 65 -618 0 net=2151
rlabel metal2 341 -618 341 -618 0 net=2252
rlabel metal2 709 -618 709 -618 0 net=5053
rlabel metal2 926 -618 926 -618 0 net=6281
rlabel metal2 961 -618 961 -618 0 net=6043
rlabel metal2 1024 -618 1024 -618 0 net=7287
rlabel metal2 37 -620 37 -620 0 net=3214
rlabel metal2 712 -620 712 -620 0 net=7430
rlabel metal2 47 -622 47 -622 0 net=376
rlabel metal2 366 -622 366 -622 0 net=2546
rlabel metal2 569 -622 569 -622 0 net=3918
rlabel metal2 786 -622 786 -622 0 net=6396
rlabel metal2 1031 -622 1031 -622 0 net=7361
rlabel metal2 51 -624 51 -624 0 net=2297
rlabel metal2 292 -624 292 -624 0 net=3853
rlabel metal2 618 -624 618 -624 0 net=4907
rlabel metal2 905 -624 905 -624 0 net=6853
rlabel metal2 982 -624 982 -624 0 net=6955
rlabel metal2 44 -626 44 -626 0 net=3807
rlabel metal2 58 -626 58 -626 0 net=1651
rlabel metal2 173 -626 173 -626 0 net=2510
rlabel metal2 730 -626 730 -626 0 net=5121
rlabel metal2 870 -626 870 -626 0 net=6025
rlabel metal2 912 -626 912 -626 0 net=6189
rlabel metal2 968 -626 968 -626 0 net=6585
rlabel metal2 40 -628 40 -628 0 net=4191
rlabel metal2 726 -628 726 -628 0 net=5321
rlabel metal2 44 -630 44 -630 0 net=4050
rlabel metal2 933 -630 933 -630 0 net=6343
rlabel metal2 72 -632 72 -632 0 net=2421
rlabel metal2 86 -632 86 -632 0 net=1506
rlabel metal2 296 -632 296 -632 0 net=2825
rlabel metal2 604 -632 604 -632 0 net=5200
rlabel metal2 940 -632 940 -632 0 net=6405
rlabel metal2 86 -634 86 -634 0 net=1667
rlabel metal2 156 -634 156 -634 0 net=1795
rlabel metal2 317 -634 317 -634 0 net=2741
rlabel metal2 359 -634 359 -634 0 net=2059
rlabel metal2 373 -634 373 -634 0 net=2355
rlabel metal2 373 -634 373 -634 0 net=2355
rlabel metal2 380 -634 380 -634 0 net=3587
rlabel metal2 394 -634 394 -634 0 net=2290
rlabel metal2 548 -634 548 -634 0 net=3375
rlabel metal2 562 -634 562 -634 0 net=5618
rlabel metal2 37 -636 37 -636 0 net=2105
rlabel metal2 380 -636 380 -636 0 net=2277
rlabel metal2 394 -636 394 -636 0 net=2615
rlabel metal2 453 -636 453 -636 0 net=3484
rlabel metal2 513 -636 513 -636 0 net=3491
rlabel metal2 572 -636 572 -636 0 net=5348
rlabel metal2 947 -636 947 -636 0 net=6411
rlabel metal2 1003 -636 1003 -636 0 net=7181
rlabel metal2 93 -638 93 -638 0 net=4740
rlabel metal2 93 -640 93 -640 0 net=3715
rlabel metal2 313 -640 313 -640 0 net=1213
rlabel metal2 387 -640 387 -640 0 net=3471
rlabel metal2 597 -640 597 -640 0 net=4161
rlabel metal2 765 -640 765 -640 0 net=4923
rlabel metal2 828 -640 828 -640 0 net=5467
rlabel metal2 863 -640 863 -640 0 net=5445
rlabel metal2 1059 -640 1059 -640 0 net=7513
rlabel metal2 100 -642 100 -642 0 net=6564
rlabel metal2 100 -644 100 -644 0 net=3511
rlabel metal2 135 -644 135 -644 0 net=2043
rlabel metal2 625 -644 625 -644 0 net=4571
rlabel metal2 107 -646 107 -646 0 net=3299
rlabel metal2 201 -646 201 -646 0 net=2054
rlabel metal2 688 -646 688 -646 0 net=5813
rlabel metal2 789 -646 789 -646 0 net=6709
rlabel metal2 114 -648 114 -648 0 net=4299
rlabel metal2 117 -650 117 -650 0 net=3991
rlabel metal2 163 -650 163 -650 0 net=2514
rlabel metal2 401 -650 401 -650 0 net=2871
rlabel metal2 495 -650 495 -650 0 net=2983
rlabel metal2 723 -650 723 -650 0 net=5245
rlabel metal2 128 -652 128 -652 0 net=6959
rlabel metal2 138 -654 138 -654 0 net=4976
rlabel metal2 142 -656 142 -656 0 net=1239
rlabel metal2 163 -656 163 -656 0 net=1745
rlabel metal2 275 -656 275 -656 0 net=1679
rlabel metal2 408 -656 408 -656 0 net=3383
rlabel metal2 562 -656 562 -656 0 net=5743
rlabel metal2 30 -658 30 -658 0 net=2683
rlabel metal2 177 -658 177 -658 0 net=6755
rlabel metal2 30 -660 30 -660 0 net=3831
rlabel metal2 124 -660 124 -660 0 net=1337
rlabel metal2 275 -660 275 -660 0 net=2079
rlabel metal2 467 -660 467 -660 0 net=3952
rlabel metal2 723 -660 723 -660 0 net=5799
rlabel metal2 177 -662 177 -662 0 net=1259
rlabel metal2 205 -662 205 -662 0 net=1722
rlabel metal2 408 -662 408 -662 0 net=2895
rlabel metal2 513 -662 513 -662 0 net=4125
rlabel metal2 653 -662 653 -662 0 net=4349
rlabel metal2 800 -662 800 -662 0 net=5147
rlabel metal2 184 -664 184 -664 0 net=1375
rlabel metal2 205 -664 205 -664 0 net=3776
rlabel metal2 352 -664 352 -664 0 net=3201
rlabel metal2 520 -664 520 -664 0 net=5825
rlabel metal2 219 -666 219 -666 0 net=1287
rlabel metal2 415 -666 415 -666 0 net=2501
rlabel metal2 439 -666 439 -666 0 net=6913
rlabel metal2 191 -668 191 -668 0 net=1699
rlabel metal2 415 -668 415 -668 0 net=3879
rlabel metal2 492 -668 492 -668 0 net=3450
rlabel metal2 702 -668 702 -668 0 net=5513
rlabel metal2 226 -670 226 -670 0 net=1233
rlabel metal2 429 -670 429 -670 0 net=4021
rlabel metal2 632 -670 632 -670 0 net=6067
rlabel metal2 422 -672 422 -672 0 net=2555
rlabel metal2 443 -672 443 -672 0 net=3177
rlabel metal2 551 -672 551 -672 0 net=4899
rlabel metal2 775 -672 775 -672 0 net=5263
rlabel metal2 856 -672 856 -672 0 net=6073
rlabel metal2 324 -674 324 -674 0 net=2807
rlabel metal2 450 -674 450 -674 0 net=4267
rlabel metal2 884 -674 884 -674 0 net=5627
rlabel metal2 422 -676 422 -676 0 net=4841
rlabel metal2 583 -676 583 -676 0 net=4081
rlabel metal2 674 -676 674 -676 0 net=4207
rlabel metal2 877 -676 877 -676 0 net=5577
rlabel metal2 103 -678 103 -678 0 net=2919
rlabel metal2 583 -678 583 -678 0 net=3525
rlabel metal2 667 -678 667 -678 0 net=4771
rlabel metal2 849 -678 849 -678 0 net=4283
rlabel metal2 467 -680 467 -680 0 net=7195
rlabel metal2 471 -682 471 -682 0 net=4265
rlabel metal2 849 -682 849 -682 0 net=7625
rlabel metal2 471 -684 471 -684 0 net=2903
rlabel metal2 667 -684 667 -684 0 net=5938
rlabel metal2 474 -686 474 -686 0 net=7121
rlabel metal2 481 -688 481 -688 0 net=2819
rlabel metal2 758 -688 758 -688 0 net=5293
rlabel metal2 716 -690 716 -690 0 net=4423
rlabel metal2 331 -692 331 -692 0 net=3233
rlabel metal2 331 -694 331 -694 0 net=1769
rlabel metal2 2 -705 2 -705 0 net=5876
rlabel metal2 128 -705 128 -705 0 net=3993
rlabel metal2 208 -705 208 -705 0 net=152
rlabel metal2 310 -705 310 -705 0 net=2872
rlabel metal2 513 -705 513 -705 0 net=5628
rlabel metal2 936 -705 936 -705 0 net=5322
rlabel metal2 1080 -705 1080 -705 0 net=4658
rlabel metal2 16 -707 16 -707 0 net=1904
rlabel metal2 373 -707 373 -707 0 net=2357
rlabel metal2 373 -707 373 -707 0 net=2357
rlabel metal2 443 -707 443 -707 0 net=439
rlabel metal2 775 -707 775 -707 0 net=6956
rlabel metal2 1083 -707 1083 -707 0 net=5648
rlabel metal2 30 -709 30 -709 0 net=3832
rlabel metal2 268 -709 268 -709 0 net=1539
rlabel metal2 282 -709 282 -709 0 net=1681
rlabel metal2 282 -709 282 -709 0 net=1681
rlabel metal2 292 -709 292 -709 0 net=1234
rlabel metal2 446 -709 446 -709 0 net=4424
rlabel metal2 880 -709 880 -709 0 net=5578
rlabel metal2 891 -709 891 -709 0 net=6915
rlabel metal2 1031 -709 1031 -709 0 net=5953
rlabel metal2 44 -711 44 -711 0 net=3809
rlabel metal2 58 -711 58 -711 0 net=1652
rlabel metal2 327 -711 327 -711 0 net=4842
rlabel metal2 436 -711 436 -711 0 net=2502
rlabel metal2 450 -711 450 -711 0 net=3589
rlabel metal2 604 -711 604 -711 0 net=5149
rlabel metal2 821 -711 821 -711 0 net=5827
rlabel metal2 884 -711 884 -711 0 net=6413
rlabel metal2 968 -711 968 -711 0 net=7635
rlabel metal2 1111 -711 1111 -711 0 net=6780
rlabel metal2 51 -713 51 -713 0 net=4171
rlabel metal2 177 -713 177 -713 0 net=1261
rlabel metal2 268 -713 268 -713 0 net=2081
rlabel metal2 289 -713 289 -713 0 net=2904
rlabel metal2 478 -713 478 -713 0 net=4572
rlabel metal2 1122 -713 1122 -713 0 net=4329
rlabel metal2 1122 -713 1122 -713 0 net=4329
rlabel metal2 58 -715 58 -715 0 net=2827
rlabel metal2 317 -715 317 -715 0 net=1215
rlabel metal2 436 -715 436 -715 0 net=2427
rlabel metal2 453 -715 453 -715 0 net=3492
rlabel metal2 590 -715 590 -715 0 net=6407
rlabel metal2 72 -717 72 -717 0 net=2423
rlabel metal2 72 -717 72 -717 0 net=2423
rlabel metal2 82 -717 82 -717 0 net=473
rlabel metal2 114 -717 114 -717 0 net=2045
rlabel metal2 142 -717 142 -717 0 net=1240
rlabel metal2 163 -717 163 -717 0 net=1747
rlabel metal2 233 -717 233 -717 0 net=2299
rlabel metal2 317 -717 317 -717 0 net=2617
rlabel metal2 401 -717 401 -717 0 net=2821
rlabel metal2 516 -717 516 -717 0 net=3234
rlabel metal2 723 -717 723 -717 0 net=6068
rlabel metal2 121 -719 121 -719 0 net=5315
rlabel metal2 485 -719 485 -719 0 net=3527
rlabel metal2 639 -719 639 -719 0 net=2984
rlabel metal2 705 -719 705 -719 0 net=5800
rlabel metal2 919 -719 919 -719 0 net=6757
rlabel metal2 93 -721 93 -721 0 net=3717
rlabel metal2 131 -721 131 -721 0 net=2742
rlabel metal2 352 -721 352 -721 0 net=3202
rlabel metal2 467 -721 467 -721 0 net=4300
rlabel metal2 870 -721 870 -721 0 net=7469
rlabel metal2 912 -721 912 -721 0 net=6711
rlabel metal2 1003 -721 1003 -721 0 net=7289
rlabel metal2 93 -723 93 -723 0 net=1771
rlabel metal2 338 -723 338 -723 0 net=2754
rlabel metal2 541 -723 541 -723 0 net=4127
rlabel metal2 653 -723 653 -723 0 net=4351
rlabel metal2 688 -723 688 -723 0 net=5815
rlabel metal2 877 -723 877 -723 0 net=4285
rlabel metal2 940 -723 940 -723 0 net=6044
rlabel metal2 996 -723 996 -723 0 net=7183
rlabel metal2 135 -725 135 -725 0 net=404
rlabel metal2 163 -725 163 -725 0 net=1377
rlabel metal2 205 -725 205 -725 0 net=1977
rlabel metal2 352 -725 352 -725 0 net=2279
rlabel metal2 457 -725 457 -725 0 net=4908
rlabel metal2 639 -725 639 -725 0 net=4209
rlabel metal2 688 -725 688 -725 0 net=5055
rlabel metal2 716 -725 716 -725 0 net=7040
rlabel metal2 142 -727 142 -727 0 net=2685
rlabel metal2 173 -727 173 -727 0 net=342
rlabel metal2 471 -727 471 -727 0 net=2921
rlabel metal2 513 -727 513 -727 0 net=3793
rlabel metal2 646 -727 646 -727 0 net=4269
rlabel metal2 709 -727 709 -727 0 net=5123
rlabel metal2 737 -727 737 -727 0 net=4901
rlabel metal2 747 -727 747 -727 0 net=6977
rlabel metal2 989 -727 989 -727 0 net=7559
rlabel metal2 65 -729 65 -729 0 net=2152
rlabel metal2 184 -729 184 -729 0 net=3473
rlabel metal2 457 -729 457 -729 0 net=6344
rlabel metal2 37 -731 37 -731 0 net=2107
rlabel metal2 226 -731 226 -731 0 net=2001
rlabel metal2 359 -731 359 -731 0 net=2060
rlabel metal2 380 -731 380 -731 0 net=2803
rlabel metal2 544 -731 544 -731 0 net=6960
rlabel metal2 30 -733 30 -733 0 net=6351
rlabel metal2 226 -733 226 -733 0 net=2955
rlabel metal2 730 -733 730 -733 0 net=5067
rlabel metal2 863 -733 863 -733 0 net=5446
rlabel metal2 233 -735 233 -735 0 net=1797
rlabel metal2 261 -735 261 -735 0 net=1339
rlabel metal2 506 -735 506 -735 0 net=3179
rlabel metal2 555 -735 555 -735 0 net=3385
rlabel metal2 583 -735 583 -735 0 net=4029
rlabel metal2 723 -735 723 -735 0 net=4925
rlabel metal2 775 -735 775 -735 0 net=6854
rlabel metal2 79 -737 79 -737 0 net=6735
rlabel metal2 786 -737 786 -737 0 net=6190
rlabel metal2 79 -739 79 -739 0 net=1669
rlabel metal2 240 -739 240 -739 0 net=1689
rlabel metal2 261 -739 261 -739 0 net=2897
rlabel metal2 464 -739 464 -739 0 net=3227
rlabel metal2 534 -739 534 -739 0 net=4463
rlabel metal2 562 -739 562 -739 0 net=5363
rlabel metal2 751 -739 751 -739 0 net=4266
rlabel metal2 954 -739 954 -739 0 net=5433
rlabel metal2 23 -741 23 -741 0 net=4480
rlabel metal2 240 -741 240 -741 0 net=2029
rlabel metal2 310 -741 310 -741 0 net=2201
rlabel metal2 362 -741 362 -741 0 net=2556
rlabel metal2 495 -741 495 -741 0 net=6045
rlabel metal2 681 -741 681 -741 0 net=4773
rlabel metal2 702 -741 702 -741 0 net=5515
rlabel metal2 758 -741 758 -741 0 net=5294
rlabel metal2 786 -741 786 -741 0 net=5265
rlabel metal2 856 -741 856 -741 0 net=6075
rlabel metal2 23 -743 23 -743 0 net=4641
rlabel metal2 219 -743 219 -743 0 net=1289
rlabel metal2 324 -743 324 -743 0 net=2809
rlabel metal2 387 -743 387 -743 0 net=3881
rlabel metal2 534 -743 534 -743 0 net=3703
rlabel metal2 597 -743 597 -743 0 net=4163
rlabel metal2 100 -745 100 -745 0 net=3513
rlabel metal2 597 -745 597 -745 0 net=5469
rlabel metal2 856 -745 856 -745 0 net=6283
rlabel metal2 100 -747 100 -747 0 net=117
rlabel metal2 208 -747 208 -747 0 net=3305
rlabel metal2 653 -747 653 -747 0 net=7336
rlabel metal2 107 -749 107 -749 0 net=3301
rlabel metal2 212 -749 212 -749 0 net=1625
rlabel metal2 324 -749 324 -749 0 net=1621
rlabel metal2 408 -749 408 -749 0 net=3377
rlabel metal2 656 -749 656 -749 0 net=5151
rlabel metal2 702 -749 702 -749 0 net=7514
rlabel metal2 107 -751 107 -751 0 net=1701
rlabel metal2 548 -751 548 -751 0 net=4193
rlabel metal2 758 -751 758 -751 0 net=7122
rlabel metal2 103 -753 103 -753 0 net=3285
rlabel metal2 660 -753 660 -753 0 net=5246
rlabel metal2 835 -753 835 -753 0 net=6587
rlabel metal2 170 -755 170 -755 0 net=1519
rlabel metal2 814 -755 814 -755 0 net=6027
rlabel metal2 926 -755 926 -755 0 net=7711
rlabel metal2 9 -757 9 -757 0 net=126
rlabel metal2 828 -757 828 -757 0 net=5745
rlabel metal2 849 -757 849 -757 0 net=7627
rlabel metal2 982 -757 982 -757 0 net=7363
rlabel metal2 527 -759 527 -759 0 net=7061
rlabel metal2 849 -759 849 -759 0 net=7197
rlabel metal2 527 -761 527 -761 0 net=3608
rlabel metal2 576 -763 576 -763 0 net=3855
rlabel metal2 611 -765 611 -765 0 net=4023
rlabel metal2 625 -767 625 -767 0 net=4083
rlabel metal2 632 -769 632 -769 0 net=4937
rlabel metal2 761 -771 761 -771 0 net=7063
rlabel metal2 2 -782 2 -782 0 net=5081
rlabel metal2 173 -782 173 -782 0 net=169
rlabel metal2 492 -782 492 -782 0 net=5487
rlabel metal2 1087 -782 1087 -782 0 net=7431
rlabel metal2 1108 -782 1108 -782 0 net=7487
rlabel metal2 16 -784 16 -784 0 net=3475
rlabel metal2 194 -784 194 -784 0 net=1622
rlabel metal2 408 -784 408 -784 0 net=3379
rlabel metal2 499 -784 499 -784 0 net=1340
rlabel metal2 667 -784 667 -784 0 net=4353
rlabel metal2 719 -784 719 -784 0 net=4902
rlabel metal2 779 -784 779 -784 0 net=7065
rlabel metal2 1122 -784 1122 -784 0 net=4331
rlabel metal2 23 -786 23 -786 0 net=4642
rlabel metal2 149 -786 149 -786 0 net=2083
rlabel metal2 275 -786 275 -786 0 net=1541
rlabel metal2 275 -786 275 -786 0 net=1541
rlabel metal2 289 -786 289 -786 0 net=2203
rlabel metal2 355 -786 355 -786 0 net=6247
rlabel metal2 957 -786 957 -786 0 net=7184
rlabel metal2 1010 -786 1010 -786 0 net=7437
rlabel metal2 1139 -786 1139 -786 0 net=271
rlabel metal2 23 -788 23 -788 0 net=3121
rlabel metal2 107 -788 107 -788 0 net=1702
rlabel metal2 341 -788 341 -788 0 net=2280
rlabel metal2 373 -788 373 -788 0 net=2359
rlabel metal2 373 -788 373 -788 0 net=2359
rlabel metal2 408 -788 408 -788 0 net=2601
rlabel metal2 506 -788 506 -788 0 net=3180
rlabel metal2 537 -788 537 -788 0 net=4938
rlabel metal2 646 -788 646 -788 0 net=4271
rlabel metal2 30 -790 30 -790 0 net=6767
rlabel metal2 548 -790 548 -790 0 net=4195
rlabel metal2 674 -790 674 -790 0 net=6047
rlabel metal2 947 -790 947 -790 0 net=7290
rlabel metal2 37 -792 37 -792 0 net=6352
rlabel metal2 37 -792 37 -792 0 net=6352
rlabel metal2 40 -792 40 -792 0 net=544
rlabel metal2 621 -792 621 -792 0 net=7470
rlabel metal2 884 -792 884 -792 0 net=6415
rlabel metal2 44 -794 44 -794 0 net=3811
rlabel metal2 44 -794 44 -794 0 net=3811
rlabel metal2 51 -794 51 -794 0 net=4173
rlabel metal2 177 -794 177 -794 0 net=1749
rlabel metal2 198 -794 198 -794 0 net=1263
rlabel metal2 208 -794 208 -794 0 net=2030
rlabel metal2 247 -794 247 -794 0 net=3287
rlabel metal2 513 -794 513 -794 0 net=3795
rlabel metal2 562 -794 562 -794 0 net=3705
rlabel metal2 625 -794 625 -794 0 net=4085
rlabel metal2 625 -794 625 -794 0 net=4085
rlabel metal2 653 -794 653 -794 0 net=7062
rlabel metal2 866 -794 866 -794 0 net=7167
rlabel metal2 51 -796 51 -796 0 net=2483
rlabel metal2 464 -796 464 -796 0 net=5023
rlabel metal2 768 -796 768 -796 0 net=7263
rlabel metal2 58 -798 58 -798 0 net=2828
rlabel metal2 541 -798 541 -798 0 net=4129
rlabel metal2 912 -798 912 -798 0 net=6713
rlabel metal2 58 -800 58 -800 0 net=2899
rlabel metal2 268 -800 268 -800 0 net=3591
rlabel metal2 453 -800 453 -800 0 net=7628
rlabel metal2 961 -800 961 -800 0 net=4165
rlabel metal2 65 -802 65 -802 0 net=2109
rlabel metal2 128 -802 128 -802 0 net=3995
rlabel metal2 569 -802 569 -802 0 net=3387
rlabel metal2 569 -802 569 -802 0 net=3387
rlabel metal2 583 -802 583 -802 0 net=4031
rlabel metal2 583 -802 583 -802 0 net=4031
rlabel metal2 593 -802 593 -802 0 net=7373
rlabel metal2 65 -804 65 -804 0 net=2425
rlabel metal2 75 -804 75 -804 0 net=3749
rlabel metal2 128 -804 128 -804 0 net=2957
rlabel metal2 240 -804 240 -804 0 net=2653
rlabel metal2 604 -804 604 -804 0 net=5150
rlabel metal2 653 -804 653 -804 0 net=7677
rlabel metal2 86 -806 86 -806 0 net=2047
rlabel metal2 156 -806 156 -806 0 net=1561
rlabel metal2 345 -806 345 -806 0 net=3307
rlabel metal2 422 -806 422 -806 0 net=1216
rlabel metal2 457 -806 457 -806 0 net=7712
rlabel metal2 982 -806 982 -806 0 net=7365
rlabel metal2 114 -808 114 -808 0 net=2301
rlabel metal2 310 -808 310 -808 0 net=2003
rlabel metal2 359 -808 359 -808 0 net=2811
rlabel metal2 478 -808 478 -808 0 net=5317
rlabel metal2 737 -808 737 -808 0 net=5365
rlabel metal2 93 -810 93 -810 0 net=1773
rlabel metal2 313 -810 313 -810 0 net=3228
rlabel metal2 527 -810 527 -810 0 net=6543
rlabel metal2 989 -810 989 -810 0 net=7561
rlabel metal2 93 -812 93 -812 0 net=1979
rlabel metal2 380 -812 380 -812 0 net=2805
rlabel metal2 607 -812 607 -812 0 net=3923
rlabel metal2 877 -812 877 -812 0 net=7651
rlabel metal2 152 -814 152 -814 0 net=1451
rlabel metal2 383 -814 383 -814 0 net=1847
rlabel metal2 614 -814 614 -814 0 net=7198
rlabel metal2 898 -814 898 -814 0 net=4287
rlabel metal2 926 -814 926 -814 0 net=5955
rlabel metal2 177 -816 177 -816 0 net=1583
rlabel metal2 317 -816 317 -816 0 net=2619
rlabel metal2 422 -816 422 -816 0 net=2429
rlabel metal2 443 -816 443 -816 0 net=6408
rlabel metal2 656 -816 656 -816 0 net=362
rlabel metal2 744 -816 744 -816 0 net=4813
rlabel metal2 142 -818 142 -818 0 net=2687
rlabel metal2 457 -818 457 -818 0 net=3529
rlabel metal2 495 -818 495 -818 0 net=5401
rlabel metal2 656 -818 656 -818 0 net=6195
rlabel metal2 142 -820 142 -820 0 net=1799
rlabel metal2 254 -820 254 -820 0 net=1691
rlabel metal2 387 -820 387 -820 0 net=3882
rlabel metal2 660 -820 660 -820 0 net=7453
rlabel metal2 121 -822 121 -822 0 net=3719
rlabel metal2 317 -822 317 -822 0 net=1709
rlabel metal2 387 -822 387 -822 0 net=3515
rlabel metal2 436 -822 436 -822 0 net=2573
rlabel metal2 751 -822 751 -822 0 net=5517
rlabel metal2 863 -822 863 -822 0 net=6077
rlabel metal2 79 -824 79 -824 0 net=1671
rlabel metal2 198 -824 198 -824 0 net=1521
rlabel metal2 222 -824 222 -824 0 net=2393
rlabel metal2 261 -824 261 -824 0 net=5653
rlabel metal2 401 -824 401 -824 0 net=2823
rlabel metal2 751 -824 751 -824 0 net=4757
rlabel metal2 212 -826 212 -826 0 net=1461
rlabel metal2 233 -826 233 -826 0 net=1315
rlabel metal2 471 -826 471 -826 0 net=2923
rlabel metal2 520 -826 520 -826 0 net=3073
rlabel metal2 779 -826 779 -826 0 net=5829
rlabel metal2 828 -826 828 -826 0 net=5747
rlabel metal2 324 -828 324 -828 0 net=4561
rlabel metal2 765 -828 765 -828 0 net=6737
rlabel metal2 401 -830 401 -830 0 net=2715
rlabel metal2 660 -830 660 -830 0 net=4775
rlabel metal2 723 -830 723 -830 0 net=4927
rlabel metal2 828 -830 828 -830 0 net=5435
rlabel metal2 135 -832 135 -832 0 net=7347
rlabel metal2 772 -832 772 -832 0 net=4977
rlabel metal2 135 -834 135 -834 0 net=1379
rlabel metal2 471 -834 471 -834 0 net=4025
rlabel metal2 688 -834 688 -834 0 net=5057
rlabel metal2 793 -834 793 -834 0 net=6758
rlabel metal2 163 -836 163 -836 0 net=1627
rlabel metal2 478 -836 478 -836 0 net=5470
rlabel metal2 604 -836 604 -836 0 net=6449
rlabel metal2 219 -838 219 -838 0 net=1290
rlabel metal2 555 -838 555 -838 0 net=4465
rlabel metal2 730 -838 730 -838 0 net=5069
rlabel metal2 807 -838 807 -838 0 net=5817
rlabel metal2 282 -840 282 -840 0 net=1683
rlabel metal2 555 -840 555 -840 0 net=6978
rlabel metal2 814 -840 814 -840 0 net=6029
rlabel metal2 191 -842 191 -842 0 net=3303
rlabel metal2 565 -842 565 -842 0 net=365
rlabel metal2 786 -842 786 -842 0 net=5267
rlabel metal2 835 -842 835 -842 0 net=6589
rlabel metal2 103 -844 103 -844 0 net=5489
rlabel metal2 863 -844 863 -844 0 net=7636
rlabel metal2 82 -846 82 -846 0 net=6345
rlabel metal2 576 -848 576 -848 0 net=3857
rlabel metal2 611 -848 611 -848 0 net=6091
rlabel metal2 352 -850 352 -850 0 net=887
rlabel metal2 579 -850 579 -850 0 net=5209
rlabel metal2 639 -852 639 -852 0 net=4211
rlabel metal2 695 -852 695 -852 0 net=5153
rlabel metal2 786 -852 786 -852 0 net=6285
rlabel metal2 338 -854 338 -854 0 net=4301
rlabel metal2 709 -854 709 -854 0 net=5125
rlabel metal2 856 -854 856 -854 0 net=6917
rlabel metal2 369 -856 369 -856 0 net=5991
rlabel metal2 394 -858 394 -858 0 net=5471
rlabel metal2 709 -858 709 -858 0 net=7449
rlabel metal2 9 -869 9 -869 0 net=2085
rlabel metal2 184 -869 184 -869 0 net=1751
rlabel metal2 184 -869 184 -869 0 net=1751
rlabel metal2 198 -869 198 -869 0 net=1523
rlabel metal2 222 -869 222 -869 0 net=3304
rlabel metal2 303 -869 303 -869 0 net=1684
rlabel metal2 303 -869 303 -869 0 net=1684
rlabel metal2 317 -869 317 -869 0 net=1710
rlabel metal2 481 -869 481 -869 0 net=3924
rlabel metal2 940 -869 940 -869 0 net=6093
rlabel metal2 940 -869 940 -869 0 net=6093
rlabel metal2 954 -869 954 -869 0 net=6249
rlabel metal2 954 -869 954 -869 0 net=6249
rlabel metal2 968 -869 968 -869 0 net=6347
rlabel metal2 968 -869 968 -869 0 net=6347
rlabel metal2 982 -869 982 -869 0 net=6545
rlabel metal2 12 -871 12 -871 0 net=902
rlabel metal2 383 -871 383 -871 0 net=910
rlabel metal2 555 -871 555 -871 0 net=4272
rlabel metal2 16 -873 16 -873 0 net=3476
rlabel metal2 170 -873 170 -873 0 net=4175
rlabel metal2 394 -873 394 -873 0 net=4978
rlabel metal2 989 -873 989 -873 0 net=7653
rlabel metal2 30 -875 30 -875 0 net=6768
rlabel metal2 492 -875 492 -875 0 net=3380
rlabel metal2 583 -875 583 -875 0 net=4033
rlabel metal2 768 -875 768 -875 0 net=6078
rlabel metal2 1052 -875 1052 -875 0 net=7169
rlabel metal2 30 -877 30 -877 0 net=48
rlabel metal2 79 -877 79 -877 0 net=5039
rlabel metal2 779 -877 779 -877 0 net=5831
rlabel metal2 912 -877 912 -877 0 net=6049
rlabel metal2 1017 -877 1017 -877 0 net=5488
rlabel metal2 44 -879 44 -879 0 net=3813
rlabel metal2 44 -879 44 -879 0 net=3813
rlabel metal2 58 -879 58 -879 0 net=2900
rlabel metal2 478 -879 478 -879 0 net=3677
rlabel metal2 537 -879 537 -879 0 net=5818
rlabel metal2 933 -879 933 -879 0 net=6197
rlabel metal2 1087 -879 1087 -879 0 net=7433
rlabel metal2 1097 -879 1097 -879 0 net=4332
rlabel metal2 16 -881 16 -881 0 net=5545
rlabel metal2 65 -881 65 -881 0 net=2426
rlabel metal2 93 -881 93 -881 0 net=1980
rlabel metal2 565 -881 565 -881 0 net=2824
rlabel metal2 709 -881 709 -881 0 net=7451
rlabel metal2 1115 -881 1115 -881 0 net=7563
rlabel metal2 72 -883 72 -883 0 net=360
rlabel metal2 75 -885 75 -885 0 net=2048
rlabel metal2 93 -885 93 -885 0 net=1563
rlabel metal2 170 -885 170 -885 0 net=1269
rlabel metal2 572 -885 572 -885 0 net=4928
rlabel metal2 856 -885 856 -885 0 net=6919
rlabel metal2 1108 -885 1108 -885 0 net=7489
rlabel metal2 79 -887 79 -887 0 net=3796
rlabel metal2 576 -887 576 -887 0 net=6087
rlabel metal2 1108 -887 1108 -887 0 net=7679
rlabel metal2 86 -889 86 -889 0 net=2959
rlabel metal2 135 -889 135 -889 0 net=1380
rlabel metal2 198 -889 198 -889 0 net=1265
rlabel metal2 229 -889 229 -889 0 net=2261
rlabel metal2 562 -889 562 -889 0 net=7703
rlabel metal2 51 -891 51 -891 0 net=2485
rlabel metal2 135 -891 135 -891 0 net=3593
rlabel metal2 275 -891 275 -891 0 net=1543
rlabel metal2 275 -891 275 -891 0 net=1543
rlabel metal2 310 -891 310 -891 0 net=2005
rlabel metal2 324 -891 324 -891 0 net=1175
rlabel metal2 548 -891 548 -891 0 net=5733
rlabel metal2 730 -891 730 -891 0 net=5155
rlabel metal2 905 -891 905 -891 0 net=4289
rlabel metal2 51 -893 51 -893 0 net=2621
rlabel metal2 418 -893 418 -893 0 net=5366
rlabel metal2 82 -895 82 -895 0 net=3977
rlabel metal2 261 -895 261 -895 0 net=2067
rlabel metal2 590 -895 590 -895 0 net=4166
rlabel metal2 114 -897 114 -897 0 net=2302
rlabel metal2 359 -897 359 -897 0 net=1452
rlabel metal2 394 -897 394 -897 0 net=2431
rlabel metal2 439 -897 439 -897 0 net=6871
rlabel metal2 1073 -897 1073 -897 0 net=7455
rlabel metal2 114 -899 114 -899 0 net=2655
rlabel metal2 268 -899 268 -899 0 net=2221
rlabel metal2 310 -899 310 -899 0 net=4169
rlabel metal2 635 -899 635 -899 0 net=6416
rlabel metal2 1010 -899 1010 -899 0 net=7265
rlabel metal2 142 -901 142 -901 0 net=1800
rlabel metal2 240 -901 240 -901 0 net=3309
rlabel metal2 359 -901 359 -901 0 net=4758
rlabel metal2 758 -901 758 -901 0 net=5025
rlabel metal2 891 -901 891 -901 0 net=5993
rlabel metal2 919 -901 919 -901 0 net=5957
rlabel metal2 947 -901 947 -901 0 net=7367
rlabel metal2 142 -903 142 -903 0 net=1463
rlabel metal2 226 -903 226 -903 0 net=1217
rlabel metal2 562 -903 562 -903 0 net=3859
rlabel metal2 604 -903 604 -903 0 net=6815
rlabel metal2 149 -905 149 -905 0 net=3601
rlabel metal2 604 -905 604 -905 0 net=3707
rlabel metal2 639 -905 639 -905 0 net=5473
rlabel metal2 898 -905 898 -905 0 net=6031
rlabel metal2 961 -905 961 -905 0 net=6739
rlabel metal2 156 -907 156 -907 0 net=2717
rlabel metal2 408 -907 408 -907 0 net=2603
rlabel metal2 443 -907 443 -907 0 net=2689
rlabel metal2 723 -907 723 -907 0 net=4467
rlabel metal2 751 -907 751 -907 0 net=5437
rlabel metal2 961 -907 961 -907 0 net=6451
rlabel metal2 996 -907 996 -907 0 net=6715
rlabel metal2 163 -909 163 -909 0 net=1629
rlabel metal2 254 -909 254 -909 0 net=3721
rlabel metal2 611 -909 611 -909 0 net=4776
rlabel metal2 674 -909 674 -909 0 net=5319
rlabel metal2 121 -911 121 -911 0 net=1673
rlabel metal2 324 -911 324 -911 0 net=3289
rlabel metal2 534 -911 534 -911 0 net=1848
rlabel metal2 625 -911 625 -911 0 net=4087
rlabel metal2 695 -911 695 -911 0 net=4303
rlabel metal2 716 -911 716 -911 0 net=4355
rlabel metal2 793 -911 793 -911 0 net=5071
rlabel metal2 2 -913 2 -913 0 net=5083
rlabel metal2 807 -913 807 -913 0 net=5211
rlabel metal2 884 -913 884 -913 0 net=6591
rlabel metal2 100 -915 100 -915 0 net=2111
rlabel metal2 163 -915 163 -915 0 net=2467
rlabel metal2 443 -915 443 -915 0 net=6611
rlabel metal2 65 -917 65 -917 0 net=2075
rlabel metal2 177 -917 177 -917 0 net=1585
rlabel metal2 331 -917 331 -917 0 net=1692
rlabel metal2 408 -917 408 -917 0 net=3531
rlabel metal2 481 -917 481 -917 0 net=3777
rlabel metal2 646 -917 646 -917 0 net=5403
rlabel metal2 716 -917 716 -917 0 net=5127
rlabel metal2 807 -917 807 -917 0 net=5491
rlabel metal2 877 -917 877 -917 0 net=5749
rlabel metal2 289 -919 289 -919 0 net=2205
rlabel metal2 338 -919 338 -919 0 net=2806
rlabel metal2 541 -919 541 -919 0 net=6697
rlabel metal2 107 -921 107 -921 0 net=3751
rlabel metal2 341 -921 341 -921 0 net=2597
rlabel metal2 450 -921 450 -921 0 net=2925
rlabel metal2 506 -921 506 -921 0 net=7374
rlabel metal2 107 -923 107 -923 0 net=2769
rlabel metal2 289 -923 289 -923 0 net=2575
rlabel metal2 457 -923 457 -923 0 net=4213
rlabel metal2 814 -923 814 -923 0 net=5269
rlabel metal2 849 -923 849 -923 0 net=5519
rlabel metal2 1059 -923 1059 -923 0 net=7439
rlabel metal2 72 -925 72 -925 0 net=7443
rlabel metal2 345 -927 345 -927 0 net=2813
rlabel metal2 471 -927 471 -927 0 net=4027
rlabel metal2 352 -929 352 -929 0 net=3985
rlabel metal2 688 -929 688 -929 0 net=6286
rlabel metal2 362 -931 362 -931 0 net=3883
rlabel metal2 464 -931 464 -931 0 net=3271
rlabel metal2 541 -931 541 -931 0 net=7066
rlabel metal2 366 -933 366 -933 0 net=5654
rlabel metal2 593 -933 593 -933 0 net=6789
rlabel metal2 352 -935 352 -935 0 net=2169
rlabel metal2 614 -935 614 -935 0 net=4609
rlabel metal2 366 -937 366 -937 0 net=2361
rlabel metal2 485 -937 485 -937 0 net=2829
rlabel metal2 569 -937 569 -937 0 net=3389
rlabel metal2 177 -939 177 -939 0 net=2631
rlabel metal2 621 -939 621 -939 0 net=7337
rlabel metal2 513 -941 513 -941 0 net=3997
rlabel metal2 373 -943 373 -943 0 net=3439
rlabel metal2 625 -943 625 -943 0 net=4130
rlabel metal2 513 -945 513 -945 0 net=3075
rlabel metal2 632 -945 632 -945 0 net=5915
rlabel metal2 23 -947 23 -947 0 net=3123
rlabel metal2 632 -947 632 -947 0 net=2981
rlabel metal2 23 -949 23 -949 0 net=3517
rlabel metal2 681 -949 681 -949 0 net=7349
rlabel metal2 247 -951 247 -951 0 net=2395
rlabel metal2 667 -951 667 -951 0 net=4197
rlabel metal2 744 -951 744 -951 0 net=4815
rlabel metal2 233 -953 233 -953 0 net=1317
rlabel metal2 667 -953 667 -953 0 net=5059
rlabel metal2 233 -955 233 -955 0 net=1775
rlabel metal2 691 -955 691 -955 0 net=4873
rlabel metal2 737 -957 737 -957 0 net=4563
rlabel metal2 37 -959 37 -959 0 net=4501
rlabel metal2 9 -970 9 -970 0 net=2086
rlabel metal2 285 -970 285 -970 0 net=4170
rlabel metal2 359 -970 359 -970 0 net=3609
rlabel metal2 859 -970 859 -970 0 net=6452
rlabel metal2 9 -972 9 -972 0 net=2831
rlabel metal2 541 -972 541 -972 0 net=2982
rlabel metal2 16 -974 16 -974 0 net=3722
rlabel metal2 607 -974 607 -974 0 net=5994
rlabel metal2 16 -976 16 -976 0 net=3711
rlabel metal2 184 -976 184 -976 0 net=1753
rlabel metal2 184 -976 184 -976 0 net=1753
rlabel metal2 194 -976 194 -976 0 net=4176
rlabel metal2 401 -976 401 -976 0 net=3885
rlabel metal2 467 -976 467 -976 0 net=5040
rlabel metal2 23 -978 23 -978 0 net=3518
rlabel metal2 439 -978 439 -978 0 net=4805
rlabel metal2 691 -978 691 -978 0 net=7103
rlabel metal2 23 -980 23 -980 0 net=4167
rlabel metal2 436 -980 436 -980 0 net=4441
rlabel metal2 569 -980 569 -980 0 net=7490
rlabel metal2 30 -982 30 -982 0 net=4869
rlabel metal2 37 -982 37 -982 0 net=1674
rlabel metal2 271 -982 271 -982 0 net=3290
rlabel metal2 362 -982 362 -982 0 net=479
rlabel metal2 632 -982 632 -982 0 net=6920
rlabel metal2 30 -984 30 -984 0 net=4035
rlabel metal2 695 -984 695 -984 0 net=5213
rlabel metal2 982 -984 982 -984 0 net=7339
rlabel metal2 698 -986 698 -986 0 net=7452
rlabel metal2 37 -988 37 -988 0 net=3815
rlabel metal2 65 -988 65 -988 0 net=6198
rlabel metal2 1045 -988 1045 -988 0 net=7457
rlabel metal2 44 -990 44 -990 0 net=3273
rlabel metal2 569 -990 569 -990 0 net=6032
rlabel metal2 933 -990 933 -990 0 net=6699
rlabel metal2 1052 -990 1052 -990 0 net=7655
rlabel metal2 2 -992 2 -992 0 net=7131
rlabel metal2 68 -994 68 -994 0 net=794
rlabel metal2 422 -994 422 -994 0 net=2599
rlabel metal2 576 -994 576 -994 0 net=4089
rlabel metal2 786 -994 786 -994 0 net=4817
rlabel metal2 68 -996 68 -996 0 net=3752
rlabel metal2 380 -996 380 -996 0 net=3077
rlabel metal2 579 -996 579 -996 0 net=5072
rlabel metal2 72 -998 72 -998 0 net=2960
rlabel metal2 114 -998 114 -998 0 net=2657
rlabel metal2 415 -998 415 -998 0 net=3125
rlabel metal2 590 -998 590 -998 0 net=5060
rlabel metal2 674 -998 674 -998 0 net=5027
rlabel metal2 786 -998 786 -998 0 net=6051
rlabel metal2 1024 -998 1024 -998 0 net=7705
rlabel metal2 72 -1000 72 -1000 0 net=1565
rlabel metal2 114 -1000 114 -1000 0 net=1545
rlabel metal2 282 -1000 282 -1000 0 net=2690
rlabel metal2 779 -1000 779 -1000 0 net=6095
rlabel metal2 82 -1002 82 -1002 0 net=2262
rlabel metal2 590 -1002 590 -1002 0 net=4199
rlabel metal2 709 -1002 709 -1002 0 net=5475
rlabel metal2 912 -1002 912 -1002 0 net=6873
rlabel metal2 82 -1004 82 -1004 0 net=5084
rlabel metal2 842 -1004 842 -1004 0 net=7351
rlabel metal2 1010 -1004 1010 -1004 0 net=6741
rlabel metal2 86 -1006 86 -1006 0 net=1587
rlabel metal2 219 -1006 219 -1006 0 net=1525
rlabel metal2 219 -1006 219 -1006 0 net=1525
rlabel metal2 229 -1006 229 -1006 0 net=1776
rlabel metal2 240 -1006 240 -1006 0 net=3310
rlabel metal2 513 -1006 513 -1006 0 net=3709
rlabel metal2 614 -1006 614 -1006 0 net=5128
rlabel metal2 793 -1006 793 -1006 0 net=5751
rlabel metal2 1010 -1006 1010 -1006 0 net=7565
rlabel metal2 93 -1008 93 -1008 0 net=2771
rlabel metal2 135 -1008 135 -1008 0 net=3594
rlabel metal2 443 -1008 443 -1008 0 net=2927
rlabel metal2 471 -1008 471 -1008 0 net=427
rlabel metal2 716 -1008 716 -1008 0 net=5157
rlabel metal2 842 -1008 842 -1008 0 net=5917
rlabel metal2 58 -1010 58 -1010 0 net=5547
rlabel metal2 863 -1010 863 -1010 0 net=6349
rlabel metal2 58 -1012 58 -1012 0 net=3437
rlabel metal2 107 -1012 107 -1012 0 net=2112
rlabel metal2 135 -1012 135 -1012 0 net=1219
rlabel metal2 233 -1012 233 -1012 0 net=2605
rlabel metal2 450 -1012 450 -1012 0 net=4305
rlabel metal2 884 -1012 884 -1012 0 net=6593
rlabel metal2 121 -1014 121 -1014 0 net=2469
rlabel metal2 191 -1014 191 -1014 0 net=3979
rlabel metal2 471 -1014 471 -1014 0 net=5173
rlabel metal2 492 -1014 492 -1014 0 net=3679
rlabel metal2 520 -1014 520 -1014 0 net=4979
rlabel metal2 548 -1014 548 -1014 0 net=5735
rlabel metal2 898 -1014 898 -1014 0 net=6817
rlabel metal2 149 -1016 149 -1016 0 net=1631
rlabel metal2 240 -1016 240 -1016 0 net=4215
rlabel metal2 474 -1016 474 -1016 0 net=7713
rlabel metal2 163 -1018 163 -1018 0 net=5549
rlabel metal2 254 -1018 254 -1018 0 net=2787
rlabel metal2 947 -1018 947 -1018 0 net=7369
rlabel metal2 975 -1018 975 -1018 0 net=7267
rlabel metal2 191 -1020 191 -1020 0 net=5251
rlabel metal2 303 -1020 303 -1020 0 net=4697
rlabel metal2 555 -1020 555 -1020 0 net=5492
rlabel metal2 856 -1020 856 -1020 0 net=6819
rlabel metal2 177 -1022 177 -1022 0 net=2633
rlabel metal2 306 -1022 306 -1022 0 net=3602
rlabel metal2 593 -1022 593 -1022 0 net=5320
rlabel metal2 177 -1024 177 -1024 0 net=3441
rlabel metal2 408 -1024 408 -1024 0 net=3533
rlabel metal2 446 -1024 446 -1024 0 net=6137
rlabel metal2 1080 -1024 1080 -1024 0 net=7435
rlabel metal2 268 -1026 268 -1026 0 net=2222
rlabel metal2 331 -1026 331 -1026 0 net=2207
rlabel metal2 408 -1026 408 -1026 0 net=3723
rlabel metal2 502 -1026 502 -1026 0 net=6995
rlabel metal2 142 -1028 142 -1028 0 net=1464
rlabel metal2 275 -1028 275 -1028 0 net=2433
rlabel metal2 457 -1028 457 -1028 0 net=4503
rlabel metal2 51 -1030 51 -1030 0 net=2622
rlabel metal2 478 -1030 478 -1030 0 net=6088
rlabel metal2 2 -1032 2 -1032 0 net=1050
rlabel metal2 100 -1032 100 -1032 0 net=2077
rlabel metal2 156 -1032 156 -1032 0 net=2719
rlabel metal2 481 -1032 481 -1032 0 net=4028
rlabel metal2 156 -1034 156 -1034 0 net=1319
rlabel metal2 289 -1034 289 -1034 0 net=2577
rlabel metal2 338 -1034 338 -1034 0 net=3051
rlabel metal2 583 -1034 583 -1034 0 net=3390
rlabel metal2 247 -1036 247 -1036 0 net=2007
rlabel metal2 600 -1036 600 -1036 0 net=5777
rlabel metal2 891 -1036 891 -1036 0 net=6717
rlabel metal2 289 -1038 289 -1038 0 net=2815
rlabel metal2 618 -1038 618 -1038 0 net=6659
rlabel metal2 1003 -1038 1003 -1038 0 net=7445
rlabel metal2 261 -1040 261 -1040 0 net=2069
rlabel metal2 562 -1040 562 -1040 0 net=3861
rlabel metal2 621 -1040 621 -1040 0 net=5832
rlabel metal2 919 -1040 919 -1040 0 net=5959
rlabel metal2 261 -1042 261 -1042 0 net=2171
rlabel metal2 499 -1042 499 -1042 0 net=6979
rlabel metal2 310 -1044 310 -1044 0 net=2397
rlabel metal2 562 -1044 562 -1044 0 net=4633
rlabel metal2 635 -1044 635 -1044 0 net=5438
rlabel metal2 870 -1044 870 -1044 0 net=6613
rlabel metal2 317 -1046 317 -1046 0 net=1331
rlabel metal2 572 -1046 572 -1046 0 net=6747
rlabel metal2 989 -1046 989 -1046 0 net=7681
rlabel metal2 352 -1048 352 -1048 0 net=2363
rlabel metal2 387 -1048 387 -1048 0 net=3778
rlabel metal2 667 -1048 667 -1048 0 net=4875
rlabel metal2 128 -1050 128 -1050 0 net=2487
rlabel metal2 495 -1050 495 -1050 0 net=5925
rlabel metal2 737 -1050 737 -1050 0 net=7564
rlabel metal2 128 -1052 128 -1052 0 net=1271
rlabel metal2 534 -1052 534 -1052 0 net=3987
rlabel metal2 751 -1052 751 -1052 0 net=5271
rlabel metal2 1129 -1052 1129 -1052 0 net=7171
rlabel metal2 170 -1054 170 -1054 0 net=1267
rlabel metal2 611 -1054 611 -1054 0 net=4623
rlabel metal2 800 -1054 800 -1054 0 net=6791
rlabel metal2 198 -1056 198 -1056 0 net=3998
rlabel metal2 611 -1058 611 -1058 0 net=4357
rlabel metal2 744 -1058 744 -1058 0 net=4565
rlabel metal2 849 -1058 849 -1058 0 net=6251
rlabel metal2 625 -1060 625 -1060 0 net=6353
rlabel metal2 954 -1060 954 -1060 0 net=7441
rlabel metal2 502 -1062 502 -1062 0 net=5737
rlabel metal2 635 -1062 635 -1062 0 net=6515
rlabel metal2 723 -1064 723 -1064 0 net=4290
rlabel metal2 730 -1066 730 -1066 0 net=4469
rlabel metal2 1143 -1066 1143 -1066 0 net=6547
rlabel metal2 660 -1068 660 -1068 0 net=5405
rlabel metal2 660 -1070 660 -1070 0 net=4611
rlabel metal2 758 -1072 758 -1072 0 net=5521
rlabel metal2 604 -1074 604 -1074 0 net=6639
rlabel metal2 5 -1085 5 -1085 0 net=1194
rlabel metal2 366 -1085 366 -1085 0 net=2489
rlabel metal2 390 -1085 390 -1085 0 net=6818
rlabel metal2 947 -1085 947 -1085 0 net=6820
rlabel metal2 1041 -1085 1041 -1085 0 net=5960
rlabel metal2 1076 -1085 1076 -1085 0 net=7436
rlabel metal2 1122 -1085 1122 -1085 0 net=7173
rlabel metal2 1143 -1085 1143 -1085 0 net=6549
rlabel metal2 9 -1087 9 -1087 0 net=2832
rlabel metal2 488 -1087 488 -1087 0 net=4980
rlabel metal2 523 -1087 523 -1087 0 net=6660
rlabel metal2 905 -1087 905 -1087 0 net=6749
rlabel metal2 968 -1087 968 -1087 0 net=7371
rlabel metal2 968 -1087 968 -1087 0 net=7371
rlabel metal2 996 -1087 996 -1087 0 net=6996
rlabel metal2 9 -1089 9 -1089 0 net=4037
rlabel metal2 40 -1089 40 -1089 0 net=6459
rlabel metal2 982 -1089 982 -1089 0 net=7341
rlabel metal2 1031 -1089 1031 -1089 0 net=6743
rlabel metal2 16 -1091 16 -1091 0 net=3712
rlabel metal2 506 -1091 506 -1091 0 net=3681
rlabel metal2 506 -1091 506 -1091 0 net=3681
rlabel metal2 513 -1091 513 -1091 0 net=3710
rlabel metal2 723 -1091 723 -1091 0 net=5273
rlabel metal2 779 -1091 779 -1091 0 net=6097
rlabel metal2 856 -1091 856 -1091 0 net=6517
rlabel metal2 926 -1091 926 -1091 0 net=7133
rlabel metal2 1017 -1091 1017 -1091 0 net=7715
rlabel metal2 1045 -1091 1045 -1091 0 net=7459
rlabel metal2 1045 -1091 1045 -1091 0 net=7459
rlabel metal2 1052 -1091 1052 -1091 0 net=7657
rlabel metal2 1052 -1091 1052 -1091 0 net=7657
rlabel metal2 51 -1093 51 -1093 0 net=3438
rlabel metal2 61 -1093 61 -1093 0 net=81
rlabel metal2 212 -1093 212 -1093 0 net=4566
rlabel metal2 817 -1093 817 -1093 0 net=7442
rlabel metal2 1010 -1093 1010 -1093 0 net=7567
rlabel metal2 51 -1095 51 -1095 0 net=2435
rlabel metal2 324 -1095 324 -1095 0 net=3724
rlabel metal2 418 -1095 418 -1095 0 net=7682
rlabel metal2 1003 -1095 1003 -1095 0 net=7447
rlabel metal2 65 -1097 65 -1097 0 net=1320
rlabel metal2 166 -1097 166 -1097 0 net=5736
rlabel metal2 740 -1097 740 -1097 0 net=5721
rlabel metal2 789 -1097 789 -1097 0 net=6350
rlabel metal2 926 -1097 926 -1097 0 net=6701
rlabel metal2 940 -1097 940 -1097 0 net=7353
rlabel metal2 65 -1099 65 -1099 0 net=1567
rlabel metal2 79 -1099 79 -1099 0 net=5550
rlabel metal2 212 -1099 212 -1099 0 net=1527
rlabel metal2 268 -1099 268 -1099 0 net=2579
rlabel metal2 366 -1099 366 -1099 0 net=2845
rlabel metal2 397 -1099 397 -1099 0 net=2928
rlabel metal2 450 -1099 450 -1099 0 net=4307
rlabel metal2 527 -1099 527 -1099 0 net=2600
rlabel metal2 639 -1099 639 -1099 0 net=5927
rlabel metal2 751 -1099 751 -1099 0 net=5649
rlabel metal2 835 -1099 835 -1099 0 net=6792
rlabel metal2 870 -1099 870 -1099 0 net=6615
rlabel metal2 975 -1099 975 -1099 0 net=7269
rlabel metal2 68 -1101 68 -1101 0 net=83
rlabel metal2 541 -1101 541 -1101 0 net=6901
rlabel metal2 79 -1103 79 -1103 0 net=2773
rlabel metal2 100 -1103 100 -1103 0 net=5021
rlabel metal2 114 -1103 114 -1103 0 net=1547
rlabel metal2 205 -1103 205 -1103 0 net=2173
rlabel metal2 324 -1103 324 -1103 0 net=5579
rlabel metal2 93 -1105 93 -1105 0 net=4401
rlabel metal2 331 -1105 331 -1105 0 net=2365
rlabel metal2 401 -1105 401 -1105 0 net=2658
rlabel metal2 544 -1105 544 -1105 0 net=5548
rlabel metal2 835 -1105 835 -1105 0 net=5919
rlabel metal2 884 -1105 884 -1105 0 net=6595
rlabel metal2 72 -1107 72 -1107 0 net=3203
rlabel metal2 355 -1107 355 -1107 0 net=5769
rlabel metal2 842 -1107 842 -1107 0 net=5097
rlabel metal2 100 -1109 100 -1109 0 net=2078
rlabel metal2 149 -1109 149 -1109 0 net=1633
rlabel metal2 170 -1109 170 -1109 0 net=1268
rlabel metal2 254 -1109 254 -1109 0 net=2789
rlabel metal2 415 -1109 415 -1109 0 net=3127
rlabel metal2 450 -1109 450 -1109 0 net=3495
rlabel metal2 765 -1109 765 -1109 0 net=5779
rlabel metal2 919 -1109 919 -1109 0 net=6981
rlabel metal2 23 -1111 23 -1111 0 net=4168
rlabel metal2 177 -1111 177 -1111 0 net=3442
rlabel metal2 422 -1111 422 -1111 0 net=3981
rlabel metal2 555 -1111 555 -1111 0 net=4470
rlabel metal2 765 -1111 765 -1111 0 net=4819
rlabel metal2 23 -1113 23 -1113 0 net=3817
rlabel metal2 103 -1113 103 -1113 0 net=4806
rlabel metal2 744 -1113 744 -1113 0 net=5523
rlabel metal2 772 -1113 772 -1113 0 net=6355
rlabel metal2 891 -1113 891 -1113 0 net=6719
rlabel metal2 114 -1115 114 -1115 0 net=1273
rlabel metal2 152 -1115 152 -1115 0 net=213
rlabel metal2 383 -1115 383 -1115 0 net=7743
rlabel metal2 177 -1117 177 -1117 0 net=2635
rlabel metal2 429 -1117 429 -1117 0 net=3535
rlabel metal2 429 -1117 429 -1117 0 net=3535
rlabel metal2 436 -1117 436 -1117 0 net=4443
rlabel metal2 555 -1117 555 -1117 0 net=7706
rlabel metal2 184 -1119 184 -1119 0 net=1755
rlabel metal2 296 -1119 296 -1119 0 net=5253
rlabel metal2 492 -1119 492 -1119 0 net=2881
rlabel metal2 793 -1119 793 -1119 0 net=5753
rlabel metal2 793 -1119 793 -1119 0 net=5753
rlabel metal2 891 -1119 891 -1119 0 net=6875
rlabel metal2 121 -1121 121 -1121 0 net=2471
rlabel metal2 303 -1121 303 -1121 0 net=2071
rlabel metal2 380 -1121 380 -1121 0 net=3079
rlabel metal2 499 -1121 499 -1121 0 net=6165
rlabel metal2 877 -1121 877 -1121 0 net=6641
rlabel metal2 30 -1123 30 -1123 0 net=3065
rlabel metal2 373 -1123 373 -1123 0 net=2208
rlabel metal2 499 -1123 499 -1123 0 net=174
rlabel metal2 44 -1125 44 -1125 0 net=3275
rlabel metal2 502 -1125 502 -1125 0 net=6052
rlabel metal2 44 -1127 44 -1127 0 net=4517
rlabel metal2 576 -1127 576 -1127 0 net=4090
rlabel metal2 607 -1127 607 -1127 0 net=3862
rlabel metal2 632 -1127 632 -1127 0 net=5869
rlabel metal2 110 -1129 110 -1129 0 net=6267
rlabel metal2 121 -1131 121 -1131 0 net=2817
rlabel metal2 387 -1131 387 -1131 0 net=4865
rlabel metal2 639 -1131 639 -1131 0 net=5477
rlabel metal2 163 -1133 163 -1133 0 net=3929
rlabel metal2 481 -1133 481 -1133 0 net=1122
rlabel metal2 184 -1135 184 -1135 0 net=2241
rlabel metal2 565 -1135 565 -1135 0 net=5049
rlabel metal2 191 -1137 191 -1137 0 net=3779
rlabel metal2 569 -1137 569 -1137 0 net=4359
rlabel metal2 618 -1137 618 -1137 0 net=4625
rlabel metal2 653 -1137 653 -1137 0 net=4871
rlabel metal2 86 -1139 86 -1139 0 net=1589
rlabel metal2 215 -1139 215 -1139 0 net=381
rlabel metal2 558 -1139 558 -1139 0 net=4879
rlabel metal2 667 -1139 667 -1139 0 net=4877
rlabel metal2 667 -1139 667 -1139 0 net=4877
rlabel metal2 684 -1139 684 -1139 0 net=7104
rlabel metal2 86 -1141 86 -1141 0 net=1333
rlabel metal2 415 -1141 415 -1141 0 net=4785
rlabel metal2 709 -1141 709 -1141 0 net=5159
rlabel metal2 849 -1141 849 -1141 0 net=6253
rlabel metal2 54 -1143 54 -1143 0 net=5551
rlabel metal2 807 -1143 807 -1143 0 net=6139
rlabel metal2 128 -1145 128 -1145 0 net=2281
rlabel metal2 583 -1145 583 -1145 0 net=905
rlabel metal2 226 -1147 226 -1147 0 net=1465
rlabel metal2 471 -1147 471 -1147 0 net=5175
rlabel metal2 135 -1149 135 -1149 0 net=1221
rlabel metal2 240 -1149 240 -1149 0 net=4217
rlabel metal2 586 -1149 586 -1149 0 net=6055
rlabel metal2 135 -1151 135 -1151 0 net=3989
rlabel metal2 562 -1151 562 -1151 0 net=4635
rlabel metal2 590 -1151 590 -1151 0 net=4201
rlabel metal2 590 -1151 590 -1151 0 net=4201
rlabel metal2 604 -1151 604 -1151 0 net=4995
rlabel metal2 240 -1153 240 -1153 0 net=3053
rlabel metal2 457 -1153 457 -1153 0 net=4505
rlabel metal2 478 -1153 478 -1153 0 net=2721
rlabel metal2 534 -1153 534 -1153 0 net=5215
rlabel metal2 247 -1155 247 -1155 0 net=2009
rlabel metal2 310 -1155 310 -1155 0 net=2399
rlabel metal2 359 -1155 359 -1155 0 net=3611
rlabel metal2 548 -1155 548 -1155 0 net=4699
rlabel metal2 625 -1155 625 -1155 0 net=5739
rlabel metal2 233 -1157 233 -1157 0 net=2607
rlabel metal2 317 -1157 317 -1157 0 net=3887
rlabel metal2 548 -1157 548 -1157 0 net=4613
rlabel metal2 674 -1157 674 -1157 0 net=5029
rlabel metal2 37 -1159 37 -1159 0 net=5961
rlabel metal2 282 -1159 282 -1159 0 net=5409
rlabel metal2 464 -1161 464 -1161 0 net=4861
rlabel metal2 660 -1161 660 -1161 0 net=5407
rlabel metal2 730 -1163 730 -1163 0 net=7663
rlabel metal2 2 -1174 2 -1174 0 net=5111
rlabel metal2 149 -1174 149 -1174 0 net=2175
rlabel metal2 226 -1174 226 -1174 0 net=1222
rlabel metal2 313 -1174 313 -1174 0 net=5770
rlabel metal2 835 -1174 835 -1174 0 net=5921
rlabel metal2 835 -1174 835 -1174 0 net=5921
rlabel metal2 982 -1174 982 -1174 0 net=7135
rlabel metal2 1115 -1174 1115 -1174 0 net=7174
rlabel metal2 1129 -1174 1129 -1174 0 net=3905
rlabel metal2 16 -1176 16 -1176 0 net=3780
rlabel metal2 303 -1176 303 -1176 0 net=2073
rlabel metal2 460 -1176 460 -1176 0 net=4506
rlabel metal2 485 -1176 485 -1176 0 net=2723
rlabel metal2 506 -1176 506 -1176 0 net=3683
rlabel metal2 558 -1176 558 -1176 0 net=5030
rlabel metal2 730 -1176 730 -1176 0 net=6596
rlabel metal2 989 -1176 989 -1176 0 net=7271
rlabel metal2 1150 -1176 1150 -1176 0 net=6551
rlabel metal2 16 -1178 16 -1178 0 net=1549
rlabel metal2 383 -1178 383 -1178 0 net=537
rlabel metal2 485 -1178 485 -1178 0 net=4701
rlabel metal2 653 -1178 653 -1178 0 net=4997
rlabel metal2 751 -1178 751 -1178 0 net=5651
rlabel metal2 863 -1178 863 -1178 0 net=6167
rlabel metal2 996 -1178 996 -1178 0 net=7343
rlabel metal2 19 -1180 19 -1180 0 net=2608
rlabel metal2 310 -1180 310 -1180 0 net=3889
rlabel metal2 331 -1180 331 -1180 0 net=2366
rlabel metal2 359 -1180 359 -1180 0 net=4807
rlabel metal2 912 -1180 912 -1180 0 net=6643
rlabel metal2 1003 -1180 1003 -1180 0 net=7355
rlabel metal2 23 -1182 23 -1182 0 net=3818
rlabel metal2 58 -1182 58 -1182 0 net=6616
rlabel metal2 947 -1182 947 -1182 0 net=6751
rlabel metal2 1017 -1182 1017 -1182 0 net=7569
rlabel metal2 23 -1184 23 -1184 0 net=620
rlabel metal2 380 -1184 380 -1184 0 net=2791
rlabel metal2 443 -1184 443 -1184 0 net=3129
rlabel metal2 478 -1184 478 -1184 0 net=4829
rlabel metal2 562 -1184 562 -1184 0 net=5740
rlabel metal2 877 -1184 877 -1184 0 net=6269
rlabel metal2 1031 -1184 1031 -1184 0 net=7717
rlabel metal2 37 -1186 37 -1186 0 net=3545
rlabel metal2 366 -1186 366 -1186 0 net=2847
rlabel metal2 429 -1186 429 -1186 0 net=3537
rlabel metal2 464 -1186 464 -1186 0 net=4878
rlabel metal2 681 -1186 681 -1186 0 net=5177
rlabel metal2 758 -1186 758 -1186 0 net=5871
rlabel metal2 884 -1186 884 -1186 0 net=6357
rlabel metal2 1041 -1186 1041 -1186 0 net=6744
rlabel metal2 44 -1188 44 -1188 0 net=4518
rlabel metal2 394 -1188 394 -1188 0 net=2490
rlabel metal2 429 -1188 429 -1188 0 net=3037
rlabel metal2 656 -1188 656 -1188 0 net=7665
rlabel metal2 44 -1190 44 -1190 0 net=1568
rlabel metal2 96 -1190 96 -1190 0 net=3982
rlabel metal2 534 -1190 534 -1190 0 net=5217
rlabel metal2 786 -1190 786 -1190 0 net=7372
rlabel metal2 1045 -1190 1045 -1190 0 net=7461
rlabel metal2 58 -1192 58 -1192 0 net=2283
rlabel metal2 135 -1192 135 -1192 0 net=3990
rlabel metal2 506 -1192 506 -1192 0 net=7664
rlabel metal2 1052 -1192 1052 -1192 0 net=7659
rlabel metal2 61 -1194 61 -1194 0 net=2843
rlabel metal2 142 -1194 142 -1194 0 net=466
rlabel metal2 513 -1194 513 -1194 0 net=4309
rlabel metal2 681 -1194 681 -1194 0 net=6254
rlabel metal2 1059 -1194 1059 -1194 0 net=7745
rlabel metal2 65 -1196 65 -1196 0 net=6319
rlabel metal2 198 -1196 198 -1196 0 net=1548
rlabel metal2 289 -1196 289 -1196 0 net=3931
rlabel metal2 394 -1196 394 -1196 0 net=1487
rlabel metal2 562 -1196 562 -1196 0 net=4219
rlabel metal2 597 -1196 597 -1196 0 net=5408
rlabel metal2 688 -1196 688 -1196 0 net=6781
rlabel metal2 100 -1198 100 -1198 0 net=5022
rlabel metal2 121 -1198 121 -1198 0 net=2818
rlabel metal2 415 -1198 415 -1198 0 net=1905
rlabel metal2 523 -1198 523 -1198 0 net=7239
rlabel metal2 100 -1200 100 -1200 0 net=1275
rlabel metal2 121 -1200 121 -1200 0 net=4787
rlabel metal2 688 -1200 688 -1200 0 net=5553
rlabel metal2 733 -1200 733 -1200 0 net=5771
rlabel metal2 891 -1200 891 -1200 0 net=6877
rlabel metal2 79 -1202 79 -1202 0 net=2775
rlabel metal2 128 -1202 128 -1202 0 net=2637
rlabel metal2 184 -1202 184 -1202 0 net=2243
rlabel metal2 222 -1202 222 -1202 0 net=3087
rlabel metal2 296 -1202 296 -1202 0 net=2473
rlabel metal2 345 -1202 345 -1202 0 net=4872
rlabel metal2 786 -1202 786 -1202 0 net=7448
rlabel metal2 79 -1204 79 -1204 0 net=3497
rlabel metal2 527 -1204 527 -1204 0 net=4867
rlabel metal2 695 -1204 695 -1204 0 net=4821
rlabel metal2 789 -1204 789 -1204 0 net=6831
rlabel metal2 107 -1206 107 -1206 0 net=5581
rlabel metal2 345 -1206 345 -1206 0 net=3277
rlabel metal2 422 -1206 422 -1206 0 net=5255
rlabel metal2 859 -1206 859 -1206 0 net=7123
rlabel metal2 72 -1208 72 -1208 0 net=3205
rlabel metal2 373 -1208 373 -1208 0 net=5050
rlabel metal2 905 -1208 905 -1208 0 net=6519
rlabel metal2 975 -1208 975 -1208 0 net=6983
rlabel metal2 142 -1210 142 -1210 0 net=5379
rlabel metal2 422 -1210 422 -1210 0 net=2883
rlabel metal2 555 -1210 555 -1210 0 net=1891
rlabel metal2 152 -1212 152 -1212 0 net=3109
rlabel metal2 569 -1212 569 -1212 0 net=4361
rlabel metal2 702 -1212 702 -1212 0 net=5929
rlabel metal2 898 -1212 898 -1212 0 net=6461
rlabel metal2 93 -1214 93 -1214 0 net=4402
rlabel metal2 716 -1214 716 -1214 0 net=5655
rlabel metal2 919 -1214 919 -1214 0 net=6721
rlabel metal2 156 -1216 156 -1216 0 net=1635
rlabel metal2 233 -1216 233 -1216 0 net=5963
rlabel metal2 926 -1216 926 -1216 0 net=6703
rlabel metal2 86 -1218 86 -1218 0 net=1335
rlabel metal2 240 -1218 240 -1218 0 net=3055
rlabel metal2 436 -1218 436 -1218 0 net=3081
rlabel metal2 467 -1218 467 -1218 0 net=6475
rlabel metal2 576 -1218 576 -1218 0 net=4203
rlabel metal2 670 -1218 670 -1218 0 net=6109
rlabel metal2 954 -1218 954 -1218 0 net=6903
rlabel metal2 51 -1220 51 -1220 0 net=2436
rlabel metal2 583 -1220 583 -1220 0 net=4637
rlabel metal2 719 -1220 719 -1220 0 net=6377
rlabel metal2 51 -1222 51 -1222 0 net=2581
rlabel metal2 723 -1222 723 -1222 0 net=5275
rlabel metal2 828 -1222 828 -1222 0 net=6099
rlabel metal2 86 -1224 86 -1224 0 net=3819
rlabel metal2 177 -1224 177 -1224 0 net=1467
rlabel metal2 646 -1224 646 -1224 0 net=4881
rlabel metal2 737 -1224 737 -1224 0 net=6375
rlabel metal2 9 -1226 9 -1226 0 net=4039
rlabel metal2 184 -1226 184 -1226 0 net=1756
rlabel metal2 268 -1226 268 -1226 0 net=755
rlabel metal2 387 -1226 387 -1226 0 net=4863
rlabel metal2 744 -1226 744 -1226 0 net=5525
rlabel metal2 849 -1226 849 -1226 0 net=6141
rlabel metal2 9 -1228 9 -1228 0 net=3067
rlabel metal2 93 -1228 93 -1228 0 net=4091
rlabel metal2 618 -1228 618 -1228 0 net=4627
rlabel metal2 709 -1228 709 -1228 0 net=5161
rlabel metal2 779 -1228 779 -1228 0 net=5723
rlabel metal2 870 -1228 870 -1228 0 net=6057
rlabel metal2 30 -1230 30 -1230 0 net=1815
rlabel metal2 492 -1230 492 -1230 0 net=5233
rlabel metal2 779 -1230 779 -1230 0 net=5755
rlabel metal2 800 -1230 800 -1230 0 net=5781
rlabel metal2 159 -1232 159 -1232 0 net=738
rlabel metal2 625 -1232 625 -1232 0 net=4779
rlabel metal2 674 -1232 674 -1232 0 net=5411
rlabel metal2 800 -1232 800 -1232 0 net=5429
rlabel metal2 163 -1234 163 -1234 0 net=6571
rlabel metal2 163 -1236 163 -1236 0 net=1529
rlabel metal2 240 -1236 240 -1236 0 net=3871
rlabel metal2 541 -1236 541 -1236 0 net=4445
rlabel metal2 639 -1236 639 -1236 0 net=5479
rlabel metal2 968 -1236 968 -1236 0 net=6855
rlabel metal2 191 -1238 191 -1238 0 net=1591
rlabel metal2 247 -1238 247 -1238 0 net=4001
rlabel metal2 509 -1238 509 -1238 0 net=4433
rlabel metal2 548 -1238 548 -1238 0 net=4615
rlabel metal2 201 -1240 201 -1240 0 net=3843
rlabel metal2 499 -1240 499 -1240 0 net=2539
rlabel metal2 600 -1240 600 -1240 0 net=5098
rlabel metal2 212 -1242 212 -1242 0 net=2591
rlabel metal2 282 -1242 282 -1242 0 net=2401
rlabel metal2 457 -1242 457 -1242 0 net=3613
rlabel metal2 705 -1242 705 -1242 0 net=7249
rlabel metal2 254 -1244 254 -1244 0 net=2011
rlabel metal2 338 -1244 338 -1244 0 net=2309
rlabel metal2 254 -1246 254 -1246 0 net=4619
rlabel metal2 457 -1246 457 -1246 0 net=4679
rlabel metal2 2 -1257 2 -1257 0 net=5112
rlabel metal2 159 -1257 159 -1257 0 net=4864
rlabel metal2 404 -1257 404 -1257 0 net=4868
rlabel metal2 534 -1257 534 -1257 0 net=4446
rlabel metal2 632 -1257 632 -1257 0 net=5526
rlabel metal2 821 -1257 821 -1257 0 net=4808
rlabel metal2 1164 -1257 1164 -1257 0 net=6553
rlabel metal2 2 -1259 2 -1259 0 net=2583
rlabel metal2 72 -1259 72 -1259 0 net=1569
rlabel metal2 282 -1259 282 -1259 0 net=2402
rlabel metal2 317 -1259 317 -1259 0 net=3844
rlabel metal2 443 -1259 443 -1259 0 net=3539
rlabel metal2 485 -1259 485 -1259 0 net=4703
rlabel metal2 705 -1259 705 -1259 0 net=6878
rlabel metal2 1024 -1259 1024 -1259 0 net=6783
rlabel metal2 1122 -1259 1122 -1259 0 net=7661
rlabel metal2 1157 -1259 1157 -1259 0 net=3907
rlabel metal2 44 -1261 44 -1261 0 net=742
rlabel metal2 219 -1261 219 -1261 0 net=1637
rlabel metal2 219 -1261 219 -1261 0 net=1637
rlabel metal2 226 -1261 226 -1261 0 net=1593
rlabel metal2 226 -1261 226 -1261 0 net=1593
rlabel metal2 233 -1261 233 -1261 0 net=1336
rlabel metal2 303 -1261 303 -1261 0 net=1893
rlabel metal2 572 -1261 572 -1261 0 net=5782
rlabel metal2 968 -1261 968 -1261 0 net=7462
rlabel metal2 1122 -1261 1122 -1261 0 net=7719
rlabel metal2 33 -1263 33 -1263 0 net=3565
rlabel metal2 51 -1263 51 -1263 0 net=4041
rlabel metal2 191 -1263 191 -1263 0 net=7136
rlabel metal2 1143 -1263 1143 -1263 0 net=7747
rlabel metal2 47 -1265 47 -1265 0 net=6921
rlabel metal2 142 -1267 142 -1267 0 net=5381
rlabel metal2 828 -1267 828 -1267 0 net=5656
rlabel metal2 968 -1267 968 -1267 0 net=6573
rlabel metal2 1024 -1267 1024 -1267 0 net=6857
rlabel metal2 1052 -1267 1052 -1267 0 net=7125
rlabel metal2 142 -1269 142 -1269 0 net=2593
rlabel metal2 233 -1269 233 -1269 0 net=3057
rlabel metal2 317 -1269 317 -1269 0 net=1959
rlabel metal2 443 -1269 443 -1269 0 net=3111
rlabel metal2 471 -1269 471 -1269 0 net=3131
rlabel metal2 492 -1269 492 -1269 0 net=4310
rlabel metal2 618 -1269 618 -1269 0 net=4616
rlabel metal2 684 -1269 684 -1269 0 net=6520
rlabel metal2 9 -1271 9 -1271 0 net=3068
rlabel metal2 240 -1271 240 -1271 0 net=3872
rlabel metal2 408 -1271 408 -1271 0 net=2074
rlabel metal2 523 -1271 523 -1271 0 net=6100
rlabel metal2 905 -1271 905 -1271 0 net=6059
rlabel metal2 9 -1273 9 -1273 0 net=4621
rlabel metal2 261 -1273 261 -1273 0 net=2012
rlabel metal2 282 -1273 282 -1273 0 net=4681
rlabel metal2 667 -1273 667 -1273 0 net=6644
rlabel metal2 16 -1275 16 -1275 0 net=1550
rlabel metal2 632 -1275 632 -1275 0 net=5179
rlabel metal2 786 -1275 786 -1275 0 net=5873
rlabel metal2 828 -1275 828 -1275 0 net=6704
rlabel metal2 16 -1277 16 -1277 0 net=3825
rlabel metal2 191 -1277 191 -1277 0 net=2245
rlabel metal2 261 -1277 261 -1277 0 net=1551
rlabel metal2 555 -1277 555 -1277 0 net=4221
rlabel metal2 569 -1277 569 -1277 0 net=6477
rlabel metal2 1010 -1277 1010 -1277 0 net=7273
rlabel metal2 114 -1279 114 -1279 0 net=2777
rlabel metal2 268 -1279 268 -1279 0 net=2311
rlabel metal2 359 -1279 359 -1279 0 net=6255
rlabel metal2 436 -1279 436 -1279 0 net=5503
rlabel metal2 831 -1279 831 -1279 0 net=7344
rlabel metal2 58 -1281 58 -1281 0 net=2285
rlabel metal2 471 -1281 471 -1281 0 net=2725
rlabel metal2 534 -1281 534 -1281 0 net=5234
rlabel metal2 751 -1281 751 -1281 0 net=5725
rlabel metal2 877 -1281 877 -1281 0 net=5931
rlabel metal2 1066 -1281 1066 -1281 0 net=7241
rlabel metal2 58 -1283 58 -1283 0 net=3145
rlabel metal2 205 -1283 205 -1283 0 net=4003
rlabel metal2 289 -1283 289 -1283 0 net=2451
rlabel metal2 457 -1283 457 -1283 0 net=6821
rlabel metal2 86 -1285 86 -1285 0 net=3821
rlabel metal2 135 -1285 135 -1285 0 net=2844
rlabel metal2 296 -1285 296 -1285 0 net=3039
rlabel metal2 457 -1285 457 -1285 0 net=4523
rlabel metal2 576 -1285 576 -1285 0 net=4204
rlabel metal2 600 -1285 600 -1285 0 net=6376
rlabel metal2 1027 -1285 1027 -1285 0 net=1
rlabel metal2 1045 -1285 1045 -1285 0 net=6905
rlabel metal2 86 -1287 86 -1287 0 net=1277
rlabel metal2 107 -1287 107 -1287 0 net=5583
rlabel metal2 156 -1287 156 -1287 0 net=5861
rlabel metal2 891 -1287 891 -1287 0 net=6359
rlabel metal2 1003 -1287 1003 -1287 0 net=6753
rlabel metal2 26 -1289 26 -1289 0 net=4987
rlabel metal2 163 -1289 163 -1289 0 net=1531
rlabel metal2 275 -1289 275 -1289 0 net=3089
rlabel metal2 478 -1289 478 -1289 0 net=4831
rlabel metal2 796 -1289 796 -1289 0 net=5652
rlabel metal2 912 -1289 912 -1289 0 net=6169
rlabel metal2 947 -1289 947 -1289 0 net=6675
rlabel metal2 1003 -1289 1003 -1289 0 net=6833
rlabel metal2 37 -1291 37 -1291 0 net=3547
rlabel metal2 324 -1291 324 -1291 0 net=3206
rlabel metal2 590 -1291 590 -1291 0 net=4639
rlabel metal2 688 -1291 688 -1291 0 net=5555
rlabel metal2 835 -1291 835 -1291 0 net=5923
rlabel metal2 933 -1291 933 -1291 0 net=6379
rlabel metal2 1031 -1291 1031 -1291 0 net=7667
rlabel metal2 37 -1293 37 -1293 0 net=2385
rlabel metal2 247 -1293 247 -1293 0 net=1489
rlabel metal2 408 -1293 408 -1293 0 net=4229
rlabel metal2 607 -1293 607 -1293 0 net=6957
rlabel metal2 1136 -1293 1136 -1293 0 net=4709
rlabel metal2 100 -1295 100 -1295 0 net=3890
rlabel metal2 324 -1295 324 -1295 0 net=2885
rlabel metal2 495 -1295 495 -1295 0 net=4685
rlabel metal2 716 -1295 716 -1295 0 net=4717
rlabel metal2 107 -1297 107 -1297 0 net=2639
rlabel metal2 170 -1297 170 -1297 0 net=1885
rlabel metal2 639 -1297 639 -1297 0 net=6725
rlabel metal2 1108 -1297 1108 -1297 0 net=7571
rlabel metal2 30 -1299 30 -1299 0 net=1817
rlabel metal2 184 -1299 184 -1299 0 net=2195
rlabel metal2 310 -1299 310 -1299 0 net=1907
rlabel metal2 499 -1299 499 -1299 0 net=3615
rlabel metal2 541 -1299 541 -1299 0 net=4435
rlabel metal2 621 -1299 621 -1299 0 net=894
rlabel metal2 849 -1299 849 -1299 0 net=6463
rlabel metal2 1094 -1299 1094 -1299 0 net=7357
rlabel metal2 65 -1301 65 -1301 0 net=6321
rlabel metal2 513 -1301 513 -1301 0 net=3685
rlabel metal2 642 -1301 642 -1301 0 net=6984
rlabel metal2 121 -1303 121 -1303 0 net=4789
rlabel metal2 646 -1303 646 -1303 0 net=4629
rlabel metal2 670 -1303 670 -1303 0 net=5276
rlabel metal2 779 -1303 779 -1303 0 net=5757
rlabel metal2 842 -1303 842 -1303 0 net=7251
rlabel metal2 79 -1305 79 -1305 0 net=3499
rlabel metal2 338 -1305 338 -1305 0 net=4545
rlabel metal2 646 -1305 646 -1305 0 net=5219
rlabel metal2 772 -1305 772 -1305 0 net=5257
rlabel metal2 800 -1305 800 -1305 0 net=5431
rlabel metal2 940 -1305 940 -1305 0 net=6271
rlabel metal2 975 -1305 975 -1305 0 net=6723
rlabel metal2 79 -1307 79 -1307 0 net=5041
rlabel metal2 345 -1307 345 -1307 0 net=3279
rlabel metal2 506 -1307 506 -1307 0 net=3415
rlabel metal2 842 -1307 842 -1307 0 net=5773
rlabel metal2 198 -1309 198 -1309 0 net=104
rlabel metal2 348 -1309 348 -1309 0 net=6887
rlabel metal2 177 -1311 177 -1311 0 net=1469
rlabel metal2 352 -1311 352 -1311 0 net=3933
rlabel metal2 436 -1311 436 -1311 0 net=6435
rlabel metal2 352 -1313 352 -1313 0 net=2793
rlabel metal2 394 -1313 394 -1313 0 net=1281
rlabel metal2 597 -1313 597 -1313 0 net=4389
rlabel metal2 366 -1315 366 -1315 0 net=5229
rlabel metal2 856 -1315 856 -1315 0 net=6111
rlabel metal2 23 -1317 23 -1317 0 net=6303
rlabel metal2 331 -1319 331 -1319 0 net=2475
rlabel metal2 380 -1319 380 -1319 0 net=2849
rlabel metal2 520 -1319 520 -1319 0 net=5903
rlabel metal2 709 -1319 709 -1319 0 net=5413
rlabel metal2 149 -1321 149 -1321 0 net=2177
rlabel metal2 401 -1321 401 -1321 0 net=299
rlabel metal2 625 -1321 625 -1321 0 net=4781
rlabel metal2 723 -1321 723 -1321 0 net=4883
rlabel metal2 149 -1323 149 -1323 0 net=2873
rlabel metal2 695 -1323 695 -1323 0 net=4823
rlabel metal2 733 -1323 733 -1323 0 net=5964
rlabel metal2 103 -1325 103 -1325 0 net=4687
rlabel metal2 744 -1325 744 -1325 0 net=5163
rlabel metal2 884 -1325 884 -1325 0 net=6143
rlabel metal2 460 -1327 460 -1327 0 net=298
rlabel metal2 544 -1327 544 -1327 0 net=5711
rlabel metal2 653 -1329 653 -1329 0 net=944
rlabel metal2 492 -1331 492 -1331 0 net=4603
rlabel metal2 656 -1331 656 -1331 0 net=5480
rlabel metal2 548 -1333 548 -1333 0 net=2540
rlabel metal2 548 -1335 548 -1335 0 net=4093
rlabel metal2 730 -1335 730 -1335 0 net=4999
rlabel metal2 583 -1337 583 -1337 0 net=4363
rlabel metal2 478 -1339 478 -1339 0 net=2123
rlabel metal2 2 -1350 2 -1350 0 net=2584
rlabel metal2 436 -1350 436 -1350 0 net=4686
rlabel metal2 733 -1350 733 -1350 0 net=6754
rlabel metal2 1101 -1350 1101 -1350 0 net=7126
rlabel metal2 1153 -1350 1153 -1350 0 net=3908
rlabel metal2 2 -1352 2 -1352 0 net=3501
rlabel metal2 135 -1352 135 -1352 0 net=5584
rlabel metal2 359 -1352 359 -1352 0 net=2286
rlabel metal2 527 -1352 527 -1352 0 net=3617
rlabel metal2 950 -1352 950 -1352 0 net=7662
rlabel metal2 1136 -1352 1136 -1352 0 net=6554
rlabel metal2 9 -1354 9 -1354 0 net=4622
rlabel metal2 215 -1354 215 -1354 0 net=6322
rlabel metal2 506 -1354 506 -1354 0 net=3417
rlabel metal2 544 -1354 544 -1354 0 net=5220
rlabel metal2 688 -1354 688 -1354 0 net=6724
rlabel metal2 996 -1354 996 -1354 0 net=6907
rlabel metal2 16 -1356 16 -1356 0 net=3826
rlabel metal2 506 -1356 506 -1356 0 net=5180
rlabel metal2 681 -1356 681 -1356 0 net=6631
rlabel metal2 1031 -1356 1031 -1356 0 net=7669
rlabel metal2 23 -1358 23 -1358 0 net=1575
rlabel metal2 513 -1358 513 -1358 0 net=3687
rlabel metal2 513 -1358 513 -1358 0 net=3687
rlabel metal2 520 -1358 520 -1358 0 net=5775
rlabel metal2 919 -1358 919 -1358 0 net=6305
rlabel metal2 919 -1358 919 -1358 0 net=6305
rlabel metal2 940 -1358 940 -1358 0 net=6437
rlabel metal2 940 -1358 940 -1358 0 net=6437
rlabel metal2 1031 -1358 1031 -1358 0 net=7253
rlabel metal2 26 -1360 26 -1360 0 net=2778
rlabel metal2 275 -1360 275 -1360 0 net=3549
rlabel metal2 537 -1360 537 -1360 0 net=5432
rlabel metal2 1045 -1360 1045 -1360 0 net=7749
rlabel metal2 33 -1362 33 -1362 0 net=3146
rlabel metal2 65 -1362 65 -1362 0 net=3132
rlabel metal2 562 -1362 562 -1362 0 net=4525
rlabel metal2 681 -1362 681 -1362 0 net=5727
rlabel metal2 772 -1362 772 -1362 0 net=5924
rlabel metal2 44 -1364 44 -1364 0 net=3566
rlabel metal2 93 -1364 93 -1364 0 net=2640
rlabel metal2 121 -1364 121 -1364 0 net=6958
rlabel metal2 44 -1366 44 -1366 0 net=1279
rlabel metal2 100 -1366 100 -1366 0 net=4004
rlabel metal2 212 -1366 212 -1366 0 net=7229
rlabel metal2 16 -1368 16 -1368 0 net=4399
rlabel metal2 103 -1368 103 -1368 0 net=2403
rlabel metal2 289 -1368 289 -1368 0 net=3935
rlabel metal2 485 -1368 485 -1368 0 net=4640
rlabel metal2 751 -1368 751 -1368 0 net=5165
rlabel metal2 772 -1368 772 -1368 0 net=5759
rlabel metal2 842 -1368 842 -1368 0 net=6113
rlabel metal2 898 -1368 898 -1368 0 net=6859
rlabel metal2 51 -1370 51 -1370 0 net=4042
rlabel metal2 492 -1370 492 -1370 0 net=7753
rlabel metal2 51 -1372 51 -1372 0 net=2795
rlabel metal2 359 -1372 359 -1372 0 net=2851
rlabel metal2 387 -1372 387 -1372 0 net=6257
rlabel metal2 58 -1374 58 -1374 0 net=1491
rlabel metal2 268 -1374 268 -1374 0 net=2313
rlabel metal2 387 -1374 387 -1374 0 net=3281
rlabel metal2 600 -1374 600 -1374 0 net=6822
rlabel metal2 65 -1376 65 -1376 0 net=3823
rlabel metal2 128 -1376 128 -1376 0 net=1819
rlabel metal2 247 -1376 247 -1376 0 net=3041
rlabel metal2 303 -1376 303 -1376 0 net=1894
rlabel metal2 569 -1376 569 -1376 0 net=7615
rlabel metal2 37 -1378 37 -1378 0 net=2387
rlabel metal2 135 -1378 135 -1378 0 net=2179
rlabel metal2 366 -1378 366 -1378 0 net=2477
rlabel metal2 366 -1378 366 -1378 0 net=2477
rlabel metal2 373 -1378 373 -1378 0 net=2453
rlabel metal2 373 -1378 373 -1378 0 net=2453
rlabel metal2 394 -1378 394 -1378 0 net=1283
rlabel metal2 394 -1378 394 -1378 0 net=1283
rlabel metal2 408 -1378 408 -1378 0 net=3540
rlabel metal2 611 -1378 611 -1378 0 net=6574
rlabel metal2 37 -1380 37 -1380 0 net=2887
rlabel metal2 331 -1380 331 -1380 0 net=3729
rlabel metal2 422 -1380 422 -1380 0 net=3347
rlabel metal2 611 -1380 611 -1380 0 net=4688
rlabel metal2 758 -1380 758 -1380 0 net=5557
rlabel metal2 828 -1380 828 -1380 0 net=7358
rlabel metal2 72 -1382 72 -1382 0 net=1571
rlabel metal2 103 -1382 103 -1382 0 net=1107
rlabel metal2 187 -1382 187 -1382 0 net=924
rlabel metal2 443 -1382 443 -1382 0 net=3113
rlabel metal2 509 -1382 509 -1382 0 net=6597
rlabel metal2 1108 -1382 1108 -1382 0 net=4711
rlabel metal2 72 -1384 72 -1384 0 net=4223
rlabel metal2 614 -1384 614 -1384 0 net=5382
rlabel metal2 821 -1384 821 -1384 0 net=5933
rlabel metal2 79 -1386 79 -1386 0 net=5043
rlabel metal2 625 -1386 625 -1386 0 net=6272
rlabel metal2 79 -1388 79 -1388 0 net=1471
rlabel metal2 226 -1388 226 -1388 0 net=1594
rlabel metal2 618 -1388 618 -1388 0 net=4393
rlabel metal2 632 -1388 632 -1388 0 net=4605
rlabel metal2 660 -1388 660 -1388 0 net=5905
rlabel metal2 849 -1388 849 -1388 0 net=6465
rlabel metal2 110 -1390 110 -1390 0 net=7105
rlabel metal2 149 -1392 149 -1392 0 net=2874
rlabel metal2 653 -1392 653 -1392 0 net=5505
rlabel metal2 814 -1392 814 -1392 0 net=5047
rlabel metal2 149 -1394 149 -1394 0 net=1961
rlabel metal2 324 -1394 324 -1394 0 net=3091
rlabel metal2 660 -1394 660 -1394 0 net=4631
rlabel metal2 674 -1394 674 -1394 0 net=4719
rlabel metal2 775 -1394 775 -1394 0 net=5874
rlabel metal2 828 -1394 828 -1394 0 net=6381
rlabel metal2 156 -1396 156 -1396 0 net=4989
rlabel metal2 786 -1396 786 -1396 0 net=5863
rlabel metal2 877 -1396 877 -1396 0 net=6171
rlabel metal2 933 -1396 933 -1396 0 net=7243
rlabel metal2 156 -1398 156 -1398 0 net=1553
rlabel metal2 282 -1398 282 -1398 0 net=4683
rlabel metal2 695 -1398 695 -1398 0 net=4825
rlabel metal2 856 -1398 856 -1398 0 net=6888
rlabel metal2 163 -1400 163 -1400 0 net=2197
rlabel metal2 191 -1400 191 -1400 0 net=2247
rlabel metal2 219 -1400 219 -1400 0 net=1639
rlabel metal2 292 -1400 292 -1400 0 net=416
rlabel metal2 716 -1400 716 -1400 0 net=5231
rlabel metal2 870 -1400 870 -1400 0 net=6145
rlabel metal2 912 -1400 912 -1400 0 net=7275
rlabel metal2 177 -1402 177 -1402 0 net=3765
rlabel metal2 534 -1402 534 -1402 0 net=6339
rlabel metal2 926 -1402 926 -1402 0 net=5712
rlabel metal2 194 -1404 194 -1404 0 net=4227
rlabel metal2 296 -1404 296 -1404 0 net=1917
rlabel metal2 723 -1404 723 -1404 0 net=4833
rlabel metal2 765 -1404 765 -1404 0 net=5259
rlabel metal2 891 -1404 891 -1404 0 net=6361
rlabel metal2 961 -1404 961 -1404 0 net=6061
rlabel metal2 198 -1406 198 -1406 0 net=2537
rlabel metal2 737 -1406 737 -1406 0 net=5001
rlabel metal2 779 -1406 779 -1406 0 net=5415
rlabel metal2 961 -1406 961 -1406 0 net=6479
rlabel metal2 30 -1408 30 -1408 0 net=6233
rlabel metal2 982 -1408 982 -1408 0 net=6677
rlabel metal2 30 -1410 30 -1410 0 net=2595
rlabel metal2 219 -1410 219 -1410 0 net=3059
rlabel metal2 254 -1410 254 -1410 0 net=1533
rlabel metal2 310 -1410 310 -1410 0 net=1908
rlabel metal2 471 -1410 471 -1410 0 net=2727
rlabel metal2 604 -1410 604 -1410 0 net=4783
rlabel metal2 793 -1410 793 -1410 0 net=6221
rlabel metal2 989 -1410 989 -1410 0 net=6835
rlabel metal2 93 -1412 93 -1412 0 net=3247
rlabel metal2 1003 -1412 1003 -1412 0 net=6923
rlabel metal2 142 -1414 142 -1414 0 net=1887
rlabel metal2 226 -1414 226 -1414 0 net=1513
rlabel metal2 464 -1414 464 -1414 0 net=3085
rlabel metal2 639 -1414 639 -1414 0 net=4791
rlabel metal2 1073 -1414 1073 -1414 0 net=7721
rlabel metal2 96 -1416 96 -1416 0 net=1937
rlabel metal2 233 -1416 233 -1416 0 net=6019
rlabel metal2 457 -1416 457 -1416 0 net=4981
rlabel metal2 702 -1416 702 -1416 0 net=4705
rlabel metal2 254 -1418 254 -1418 0 net=6199
rlabel metal2 303 -1420 303 -1420 0 net=1787
rlabel metal2 464 -1420 464 -1420 0 net=4231
rlabel metal2 702 -1420 702 -1420 0 net=5661
rlabel metal2 310 -1422 310 -1422 0 net=4391
rlabel metal2 317 -1424 317 -1424 0 net=1757
rlabel metal2 338 -1426 338 -1426 0 net=4547
rlabel metal2 338 -1428 338 -1428 0 net=2133
rlabel metal2 499 -1428 499 -1428 0 net=4437
rlabel metal2 401 -1430 401 -1430 0 net=3781
rlabel metal2 576 -1430 576 -1430 0 net=4884
rlabel metal2 345 -1432 345 -1432 0 net=6207
rlabel metal2 345 -1434 345 -1434 0 net=2125
rlabel metal2 478 -1436 478 -1436 0 net=4436
rlabel metal2 583 -1438 583 -1438 0 net=4365
rlabel metal2 548 -1440 548 -1440 0 net=4095
rlabel metal2 548 -1442 548 -1442 0 net=6726
rlabel metal2 1017 -1444 1017 -1444 0 net=6785
rlabel metal2 1038 -1446 1038 -1446 0 net=7573
rlabel metal2 9 -1457 9 -1457 0 net=21
rlabel metal2 481 -1457 481 -1457 0 net=4784
rlabel metal2 611 -1457 611 -1457 0 net=6908
rlabel metal2 1010 -1457 1010 -1457 0 net=6063
rlabel metal2 16 -1459 16 -1459 0 net=4400
rlabel metal2 499 -1459 499 -1459 0 net=3618
rlabel metal2 996 -1459 996 -1459 0 net=7723
rlabel metal2 16 -1461 16 -1461 0 net=1703
rlabel metal2 352 -1461 352 -1461 0 net=3766
rlabel metal2 551 -1461 551 -1461 0 net=4720
rlabel metal2 681 -1461 681 -1461 0 net=5729
rlabel metal2 744 -1461 744 -1461 0 net=7750
rlabel metal2 1062 -1461 1062 -1461 0 net=5205
rlabel metal2 30 -1463 30 -1463 0 net=2596
rlabel metal2 198 -1463 198 -1463 0 net=2538
rlabel metal2 569 -1463 569 -1463 0 net=4632
rlabel metal2 681 -1463 681 -1463 0 net=5261
rlabel metal2 856 -1463 856 -1463 0 net=7276
rlabel metal2 947 -1463 947 -1463 0 net=7255
rlabel metal2 23 -1465 23 -1465 0 net=1577
rlabel metal2 257 -1465 257 -1465 0 net=1534
rlabel metal2 282 -1465 282 -1465 0 net=1641
rlabel metal2 282 -1465 282 -1465 0 net=1641
rlabel metal2 289 -1465 289 -1465 0 net=3936
rlabel metal2 415 -1465 415 -1465 0 net=3731
rlabel metal2 436 -1465 436 -1465 0 net=3169
rlabel metal2 516 -1465 516 -1465 0 net=5558
rlabel metal2 765 -1465 765 -1465 0 net=5907
rlabel metal2 856 -1465 856 -1465 0 net=6481
rlabel metal2 1017 -1465 1017 -1465 0 net=6787
rlabel metal2 23 -1467 23 -1467 0 net=3017
rlabel metal2 292 -1467 292 -1467 0 net=2852
rlabel metal2 387 -1467 387 -1467 0 net=3283
rlabel metal2 502 -1467 502 -1467 0 net=4826
rlabel metal2 747 -1467 747 -1467 0 net=6172
rlabel metal2 884 -1467 884 -1467 0 net=6340
rlabel metal2 1017 -1467 1017 -1467 0 net=7575
rlabel metal2 33 -1469 33 -1469 0 net=5232
rlabel metal2 758 -1469 758 -1469 0 net=5865
rlabel metal2 835 -1469 835 -1469 0 net=6467
rlabel metal2 44 -1471 44 -1471 0 net=1280
rlabel metal2 114 -1471 114 -1471 0 net=4228
rlabel metal2 303 -1471 303 -1471 0 net=1789
rlabel metal2 303 -1471 303 -1471 0 net=1789
rlabel metal2 310 -1471 310 -1471 0 net=4392
rlabel metal2 541 -1471 541 -1471 0 net=3419
rlabel metal2 569 -1471 569 -1471 0 net=3909
rlabel metal2 695 -1471 695 -1471 0 net=6307
rlabel metal2 933 -1471 933 -1471 0 net=7245
rlabel metal2 30 -1473 30 -1473 0 net=1881
rlabel metal2 51 -1473 51 -1473 0 net=2796
rlabel metal2 254 -1473 254 -1473 0 net=1919
rlabel metal2 310 -1473 310 -1473 0 net=4117
rlabel metal2 331 -1473 331 -1473 0 net=2455
rlabel metal2 387 -1473 387 -1473 0 net=3181
rlabel metal2 485 -1473 485 -1473 0 net=4684
rlabel metal2 730 -1473 730 -1473 0 net=4991
rlabel metal2 954 -1473 954 -1473 0 net=7231
rlabel metal2 2 -1475 2 -1475 0 net=3502
rlabel metal2 296 -1475 296 -1475 0 net=3689
rlabel metal2 541 -1475 541 -1475 0 net=4439
rlabel metal2 730 -1475 730 -1475 0 net=5167
rlabel metal2 786 -1475 786 -1475 0 net=6223
rlabel metal2 912 -1475 912 -1475 0 net=6837
rlabel metal2 1094 -1475 1094 -1475 0 net=4713
rlabel metal2 2 -1477 2 -1477 0 net=5949
rlabel metal2 103 -1477 103 -1477 0 net=538
rlabel metal2 688 -1477 688 -1477 0 net=7683
rlabel metal2 51 -1479 51 -1479 0 net=3093
rlabel metal2 345 -1479 345 -1479 0 net=2127
rlabel metal2 422 -1479 422 -1479 0 net=3349
rlabel metal2 576 -1479 576 -1479 0 net=5934
rlabel metal2 859 -1479 859 -1479 0 net=6997
rlabel metal2 37 -1481 37 -1481 0 net=2888
rlabel metal2 373 -1481 373 -1481 0 net=2315
rlabel metal2 394 -1481 394 -1481 0 net=1284
rlabel metal2 408 -1481 408 -1481 0 net=5819
rlabel metal2 821 -1481 821 -1481 0 net=6259
rlabel metal2 9 -1483 9 -1483 0 net=3505
rlabel metal2 65 -1483 65 -1483 0 net=3824
rlabel metal2 233 -1483 233 -1483 0 net=6021
rlabel metal2 863 -1483 863 -1483 0 net=6209
rlabel metal2 58 -1485 58 -1485 0 net=1493
rlabel metal2 226 -1485 226 -1485 0 net=1515
rlabel metal2 366 -1485 366 -1485 0 net=2479
rlabel metal2 401 -1485 401 -1485 0 net=2781
rlabel metal2 639 -1485 639 -1485 0 net=4793
rlabel metal2 807 -1485 807 -1485 0 net=5663
rlabel metal2 870 -1485 870 -1485 0 net=6147
rlabel metal2 58 -1487 58 -1487 0 net=1889
rlabel metal2 163 -1487 163 -1487 0 net=2198
rlabel metal2 226 -1487 226 -1487 0 net=2113
rlabel metal2 422 -1487 422 -1487 0 net=3713
rlabel metal2 807 -1487 807 -1487 0 net=6439
rlabel metal2 65 -1489 65 -1489 0 net=3115
rlabel metal2 464 -1489 464 -1489 0 net=4233
rlabel metal2 870 -1489 870 -1489 0 net=6599
rlabel metal2 72 -1491 72 -1491 0 net=4225
rlabel metal2 432 -1491 432 -1491 0 net=5561
rlabel metal2 877 -1491 877 -1491 0 net=6679
rlabel metal2 72 -1493 72 -1493 0 net=3061
rlabel metal2 439 -1493 439 -1493 0 net=5048
rlabel metal2 884 -1493 884 -1493 0 net=6861
rlabel metal2 940 -1493 940 -1493 0 net=7107
rlabel metal2 79 -1495 79 -1495 0 net=1472
rlabel metal2 443 -1495 443 -1495 0 net=3086
rlabel metal2 485 -1495 485 -1495 0 net=4706
rlabel metal2 814 -1495 814 -1495 0 net=6383
rlabel metal2 968 -1495 968 -1495 0 net=6925
rlabel metal2 1024 -1495 1024 -1495 0 net=7755
rlabel metal2 79 -1497 79 -1497 0 net=3043
rlabel metal2 443 -1497 443 -1497 0 net=3783
rlabel metal2 590 -1497 590 -1497 0 net=4367
rlabel metal2 793 -1497 793 -1497 0 net=6201
rlabel metal2 982 -1497 982 -1497 0 net=7617
rlabel metal2 86 -1499 86 -1499 0 net=1572
rlabel metal2 163 -1499 163 -1499 0 net=5776
rlabel metal2 534 -1499 534 -1499 0 net=2728
rlabel metal2 597 -1499 597 -1499 0 net=4527
rlabel metal2 779 -1499 779 -1499 0 net=5417
rlabel metal2 1003 -1499 1003 -1499 0 net=7671
rlabel metal2 86 -1501 86 -1501 0 net=1963
rlabel metal2 166 -1501 166 -1501 0 net=4606
rlabel metal2 646 -1501 646 -1501 0 net=5003
rlabel metal2 772 -1501 772 -1501 0 net=5761
rlabel metal2 828 -1501 828 -1501 0 net=6115
rlabel metal2 107 -1503 107 -1503 0 net=1938
rlabel metal2 177 -1503 177 -1503 0 net=4573
rlabel metal2 534 -1503 534 -1503 0 net=6501
rlabel metal2 842 -1503 842 -1503 0 net=6363
rlabel metal2 93 -1505 93 -1505 0 net=3249
rlabel metal2 114 -1505 114 -1505 0 net=1201
rlabel metal2 705 -1505 705 -1505 0 net=7223
rlabel metal2 93 -1507 93 -1507 0 net=948
rlabel metal2 677 -1507 677 -1507 0 net=5713
rlabel metal2 121 -1509 121 -1509 0 net=1729
rlabel metal2 691 -1509 691 -1509 0 net=6234
rlabel metal2 124 -1511 124 -1511 0 net=1820
rlabel metal2 247 -1511 247 -1511 0 net=4548
rlabel metal2 800 -1511 800 -1511 0 net=6633
rlabel metal2 128 -1513 128 -1513 0 net=2389
rlabel metal2 366 -1513 366 -1513 0 net=2191
rlabel metal2 618 -1513 618 -1513 0 net=4835
rlabel metal2 128 -1515 128 -1515 0 net=3221
rlabel metal2 212 -1515 212 -1515 0 net=7531
rlabel metal2 100 -1517 100 -1517 0 net=1473
rlabel metal2 219 -1517 219 -1517 0 net=2797
rlabel metal2 450 -1517 450 -1517 0 net=4845
rlabel metal2 555 -1517 555 -1517 0 net=5045
rlabel metal2 135 -1519 135 -1519 0 net=2181
rlabel metal2 359 -1519 359 -1519 0 net=6149
rlabel metal2 135 -1521 135 -1521 0 net=2135
rlabel metal2 457 -1521 457 -1521 0 net=4983
rlabel metal2 149 -1523 149 -1523 0 net=4395
rlabel metal2 156 -1525 156 -1525 0 net=1555
rlabel metal2 177 -1525 177 -1525 0 net=3667
rlabel metal2 457 -1525 457 -1525 0 net=4949
rlabel metal2 625 -1525 625 -1525 0 net=5507
rlabel metal2 156 -1527 156 -1527 0 net=7381
rlabel metal2 184 -1529 184 -1529 0 net=2249
rlabel metal2 240 -1529 240 -1529 0 net=1759
rlabel metal2 338 -1529 338 -1529 0 net=2659
rlabel metal2 194 -1531 194 -1531 0 net=4071
rlabel metal2 205 -1533 205 -1533 0 net=2547
rlabel metal2 527 -1533 527 -1533 0 net=3551
rlabel metal2 275 -1535 275 -1535 0 net=2405
rlabel metal2 527 -1535 527 -1535 0 net=4097
rlabel metal2 513 -1537 513 -1537 0 net=4181
rlabel metal2 2 -1548 2 -1548 0 net=5950
rlabel metal2 254 -1548 254 -1548 0 net=1921
rlabel metal2 352 -1548 352 -1548 0 net=2182
rlabel metal2 376 -1548 376 -1548 0 net=3170
rlabel metal2 457 -1548 457 -1548 0 net=4992
rlabel metal2 940 -1548 940 -1548 0 net=7109
rlabel metal2 1034 -1548 1034 -1548 0 net=6788
rlabel metal2 1045 -1548 1045 -1548 0 net=6211
rlabel metal2 5 -1550 5 -1550 0 net=1474
rlabel metal2 145 -1550 145 -1550 0 net=7587
rlabel metal2 1059 -1550 1059 -1550 0 net=6065
rlabel metal2 9 -1552 9 -1552 0 net=3506
rlabel metal2 261 -1552 261 -1552 0 net=2391
rlabel metal2 464 -1552 464 -1552 0 net=6308
rlabel metal2 772 -1552 772 -1552 0 net=6148
rlabel metal2 975 -1552 975 -1552 0 net=7533
rlabel metal2 1094 -1552 1094 -1552 0 net=4715
rlabel metal2 9 -1554 9 -1554 0 net=1877
rlabel metal2 513 -1554 513 -1554 0 net=2231
rlabel metal2 674 -1554 674 -1554 0 net=7576
rlabel metal2 1073 -1554 1073 -1554 0 net=5207
rlabel metal2 30 -1556 30 -1556 0 net=4397
rlabel metal2 156 -1556 156 -1556 0 net=2250
rlabel metal2 198 -1556 198 -1556 0 net=1579
rlabel metal2 268 -1556 268 -1556 0 net=4226
rlabel metal2 562 -1556 562 -1556 0 net=5046
rlabel metal2 926 -1556 926 -1556 0 net=7225
rlabel metal2 33 -1558 33 -1558 0 net=882
rlabel metal2 51 -1558 51 -1558 0 net=3094
rlabel metal2 471 -1558 471 -1558 0 net=6022
rlabel metal2 821 -1558 821 -1558 0 net=6261
rlabel metal2 989 -1558 989 -1558 0 net=7685
rlabel metal2 37 -1560 37 -1560 0 net=4072
rlabel metal2 660 -1560 660 -1560 0 net=5867
rlabel metal2 821 -1560 821 -1560 0 net=4843
rlabel metal2 37 -1562 37 -1562 0 net=1883
rlabel metal2 51 -1562 51 -1562 0 net=2119
rlabel metal2 478 -1562 478 -1562 0 net=3284
rlabel metal2 520 -1562 520 -1562 0 net=4836
rlabel metal2 625 -1562 625 -1562 0 net=5509
rlabel metal2 835 -1562 835 -1562 0 net=6469
rlabel metal2 961 -1562 961 -1562 0 net=7247
rlabel metal2 996 -1562 996 -1562 0 net=7725
rlabel metal2 65 -1564 65 -1564 0 net=3117
rlabel metal2 534 -1564 534 -1564 0 net=7382
rlabel metal2 16 -1566 16 -1566 0 net=1705
rlabel metal2 72 -1566 72 -1566 0 net=3063
rlabel metal2 565 -1566 565 -1566 0 net=7756
rlabel metal2 16 -1568 16 -1568 0 net=5801
rlabel metal2 268 -1568 268 -1568 0 net=2661
rlabel metal2 359 -1568 359 -1568 0 net=3237
rlabel metal2 716 -1568 716 -1568 0 net=5563
rlabel metal2 814 -1568 814 -1568 0 net=6385
rlabel metal2 982 -1568 982 -1568 0 net=7619
rlabel metal2 72 -1570 72 -1570 0 net=1965
rlabel metal2 93 -1570 93 -1570 0 net=3910
rlabel metal2 576 -1570 576 -1570 0 net=4951
rlabel metal2 716 -1570 716 -1570 0 net=5821
rlabel metal2 765 -1570 765 -1570 0 net=5909
rlabel metal2 842 -1570 842 -1570 0 net=6365
rlabel metal2 842 -1570 842 -1570 0 net=6365
rlabel metal2 859 -1570 859 -1570 0 net=7672
rlabel metal2 79 -1572 79 -1572 0 net=3045
rlabel metal2 163 -1572 163 -1572 0 net=5985
rlabel metal2 478 -1572 478 -1572 0 net=4483
rlabel metal2 684 -1572 684 -1572 0 net=7005
rlabel metal2 765 -1572 765 -1572 0 net=5665
rlabel metal2 870 -1572 870 -1572 0 net=6601
rlabel metal2 933 -1572 933 -1572 0 net=6999
rlabel metal2 79 -1574 79 -1574 0 net=2529
rlabel metal2 282 -1574 282 -1574 0 net=1642
rlabel metal2 345 -1574 345 -1574 0 net=2549
rlabel metal2 884 -1574 884 -1574 0 net=6863
rlabel metal2 86 -1576 86 -1576 0 net=1203
rlabel metal2 121 -1576 121 -1576 0 net=1731
rlabel metal2 163 -1576 163 -1576 0 net=4847
rlabel metal2 464 -1576 464 -1576 0 net=3983
rlabel metal2 625 -1576 625 -1576 0 net=7415
rlabel metal2 96 -1578 96 -1578 0 net=402
rlabel metal2 527 -1578 527 -1578 0 net=4099
rlabel metal2 590 -1578 590 -1578 0 net=6793
rlabel metal2 968 -1578 968 -1578 0 net=6927
rlabel metal2 100 -1580 100 -1580 0 net=3251
rlabel metal2 121 -1580 121 -1580 0 net=2137
rlabel metal2 166 -1580 166 -1580 0 net=2779
rlabel metal2 506 -1580 506 -1580 0 net=3351
rlabel metal2 583 -1580 583 -1580 0 net=4183
rlabel metal2 593 -1580 593 -1580 0 net=5730
rlabel metal2 723 -1580 723 -1580 0 net=6151
rlabel metal2 912 -1580 912 -1580 0 net=6839
rlabel metal2 107 -1582 107 -1582 0 net=4119
rlabel metal2 331 -1582 331 -1582 0 net=2457
rlabel metal2 597 -1582 597 -1582 0 net=4529
rlabel metal2 128 -1584 128 -1584 0 net=3222
rlabel metal2 170 -1584 170 -1584 0 net=1557
rlabel metal2 170 -1584 170 -1584 0 net=1557
rlabel metal2 177 -1584 177 -1584 0 net=2783
rlabel metal2 597 -1584 597 -1584 0 net=4369
rlabel metal2 611 -1584 611 -1584 0 net=4234
rlabel metal2 723 -1584 723 -1584 0 net=5169
rlabel metal2 793 -1584 793 -1584 0 net=6203
rlabel metal2 114 -1586 114 -1586 0 net=1939
rlabel metal2 614 -1586 614 -1586 0 net=6745
rlabel metal2 128 -1588 128 -1588 0 net=1415
rlabel metal2 366 -1588 366 -1588 0 net=2193
rlabel metal2 429 -1588 429 -1588 0 net=3733
rlabel metal2 632 -1588 632 -1588 0 net=4985
rlabel metal2 180 -1590 180 -1590 0 net=3714
rlabel metal2 457 -1590 457 -1590 0 net=5671
rlabel metal2 800 -1590 800 -1590 0 net=6635
rlabel metal2 201 -1592 201 -1592 0 net=5262
rlabel metal2 730 -1592 730 -1592 0 net=5419
rlabel metal2 205 -1594 205 -1594 0 net=1829
rlabel metal2 212 -1594 212 -1594 0 net=257
rlabel metal2 233 -1594 233 -1594 0 net=1517
rlabel metal2 635 -1594 635 -1594 0 net=5835
rlabel metal2 800 -1594 800 -1594 0 net=5967
rlabel metal2 191 -1596 191 -1596 0 net=1495
rlabel metal2 219 -1596 219 -1596 0 net=2159
rlabel metal2 278 -1596 278 -1596 0 net=5607
rlabel metal2 58 -1598 58 -1598 0 net=1890
rlabel metal2 226 -1598 226 -1598 0 net=2115
rlabel metal2 366 -1598 366 -1598 0 net=2373
rlabel metal2 639 -1598 639 -1598 0 net=4795
rlabel metal2 663 -1598 663 -1598 0 net=6440
rlabel metal2 828 -1598 828 -1598 0 net=6117
rlabel metal2 44 -1600 44 -1600 0 net=2061
rlabel metal2 233 -1600 233 -1600 0 net=3183
rlabel metal2 394 -1600 394 -1600 0 net=3669
rlabel metal2 639 -1600 639 -1600 0 net=4139
rlabel metal2 58 -1602 58 -1602 0 net=4659
rlabel metal2 737 -1602 737 -1602 0 net=5715
rlabel metal2 947 -1602 947 -1602 0 net=7257
rlabel metal2 240 -1604 240 -1604 0 net=1761
rlabel metal2 355 -1604 355 -1604 0 net=2037
rlabel metal2 408 -1604 408 -1604 0 net=2799
rlabel metal2 646 -1604 646 -1604 0 net=5005
rlabel metal2 947 -1604 947 -1604 0 net=7233
rlabel metal2 240 -1606 240 -1606 0 net=2407
rlabel metal2 324 -1606 324 -1606 0 net=561
rlabel metal2 667 -1606 667 -1606 0 net=5762
rlabel metal2 877 -1606 877 -1606 0 net=6681
rlabel metal2 282 -1608 282 -1608 0 net=1987
rlabel metal2 709 -1608 709 -1608 0 net=6503
rlabel metal2 303 -1610 303 -1610 0 net=1791
rlabel metal2 373 -1610 373 -1610 0 net=2317
rlabel metal2 408 -1610 408 -1610 0 net=2129
rlabel metal2 492 -1610 492 -1610 0 net=4575
rlabel metal2 737 -1610 737 -1610 0 net=6225
rlabel metal2 23 -1612 23 -1612 0 net=3019
rlabel metal2 523 -1612 523 -1612 0 net=5017
rlabel metal2 758 -1612 758 -1612 0 net=5341
rlabel metal2 786 -1612 786 -1612 0 net=6483
rlabel metal2 23 -1614 23 -1614 0 net=3691
rlabel metal2 310 -1614 310 -1614 0 net=2225
rlabel metal2 338 -1614 338 -1614 0 net=1995
rlabel metal2 415 -1614 415 -1614 0 net=3461
rlabel metal2 775 -1614 775 -1614 0 net=5731
rlabel metal2 856 -1614 856 -1614 0 net=6961
rlabel metal2 296 -1616 296 -1616 0 net=2481
rlabel metal2 537 -1616 537 -1616 0 net=4409
rlabel metal2 380 -1618 380 -1618 0 net=3785
rlabel metal2 443 -1620 443 -1620 0 net=4440
rlabel metal2 541 -1622 541 -1622 0 net=3553
rlabel metal2 548 -1624 548 -1624 0 net=3421
rlabel metal2 82 -1626 82 -1626 0 net=3507
rlabel metal2 9 -1637 9 -1637 0 net=1878
rlabel metal2 345 -1637 345 -1637 0 net=2117
rlabel metal2 345 -1637 345 -1637 0 net=2117
rlabel metal2 355 -1637 355 -1637 0 net=3734
rlabel metal2 607 -1637 607 -1637 0 net=6470
rlabel metal2 1059 -1637 1059 -1637 0 net=6066
rlabel metal2 23 -1639 23 -1639 0 net=3693
rlabel metal2 37 -1639 37 -1639 0 net=1884
rlabel metal2 58 -1639 58 -1639 0 net=4660
rlabel metal2 779 -1639 779 -1639 0 net=6118
rlabel metal2 1066 -1639 1066 -1639 0 net=5208
rlabel metal2 23 -1641 23 -1641 0 net=6231
rlabel metal2 149 -1641 149 -1641 0 net=3046
rlabel metal2 313 -1641 313 -1641 0 net=2780
rlabel metal2 523 -1641 523 -1641 0 net=5868
rlabel metal2 674 -1641 674 -1641 0 net=7248
rlabel metal2 1069 -1641 1069 -1641 0 net=4716
rlabel metal2 37 -1643 37 -1643 0 net=3261
rlabel metal2 222 -1643 222 -1643 0 net=3064
rlabel metal2 534 -1643 534 -1643 0 net=4101
rlabel metal2 583 -1643 583 -1643 0 net=7234
rlabel metal2 1094 -1643 1094 -1643 0 net=6213
rlabel metal2 58 -1645 58 -1645 0 net=3253
rlabel metal2 114 -1645 114 -1645 0 net=1941
rlabel metal2 247 -1645 247 -1645 0 net=1223
rlabel metal2 376 -1645 376 -1645 0 net=5732
rlabel metal2 835 -1645 835 -1645 0 net=6153
rlabel metal2 947 -1645 947 -1645 0 net=7687
rlabel metal2 51 -1647 51 -1647 0 net=2121
rlabel metal2 135 -1647 135 -1647 0 net=7737
rlabel metal2 450 -1647 450 -1647 0 net=2458
rlabel metal2 572 -1647 572 -1647 0 net=5006
rlabel metal2 16 -1649 16 -1649 0 net=5803
rlabel metal2 138 -1649 138 -1649 0 net=1762
rlabel metal2 383 -1649 383 -1649 0 net=1061
rlabel metal2 786 -1649 786 -1649 0 net=6485
rlabel metal2 912 -1649 912 -1649 0 net=6963
rlabel metal2 61 -1651 61 -1651 0 net=350
rlabel metal2 684 -1651 684 -1651 0 net=6262
rlabel metal2 65 -1653 65 -1653 0 net=1707
rlabel metal2 142 -1653 142 -1653 0 net=2785
rlabel metal2 187 -1653 187 -1653 0 net=1518
rlabel metal2 586 -1653 586 -1653 0 net=4530
rlabel metal2 79 -1655 79 -1655 0 net=3787
rlabel metal2 394 -1655 394 -1655 0 net=2038
rlabel metal2 450 -1655 450 -1655 0 net=4185
rlabel metal2 611 -1655 611 -1655 0 net=5221
rlabel metal2 691 -1655 691 -1655 0 net=5822
rlabel metal2 730 -1655 730 -1655 0 net=5421
rlabel metal2 891 -1655 891 -1655 0 net=7111
rlabel metal2 82 -1657 82 -1657 0 net=2392
rlabel metal2 460 -1657 460 -1657 0 net=4844
rlabel metal2 93 -1659 93 -1659 0 net=1417
rlabel metal2 149 -1659 149 -1659 0 net=5529
rlabel metal2 254 -1659 254 -1659 0 net=2161
rlabel metal2 380 -1659 380 -1659 0 net=5342
rlabel metal2 786 -1659 786 -1659 0 net=6205
rlabel metal2 54 -1661 54 -1661 0 net=4801
rlabel metal2 159 -1661 159 -1661 0 net=380
rlabel metal2 506 -1661 506 -1661 0 net=3555
rlabel metal2 590 -1661 590 -1661 0 net=4371
rlabel metal2 614 -1661 614 -1661 0 net=6386
rlabel metal2 96 -1663 96 -1663 0 net=4120
rlabel metal2 170 -1663 170 -1663 0 net=1558
rlabel metal2 401 -1663 401 -1663 0 net=2194
rlabel metal2 639 -1663 639 -1663 0 net=4140
rlabel metal2 667 -1663 667 -1663 0 net=4410
rlabel metal2 765 -1663 765 -1663 0 net=5667
rlabel metal2 898 -1663 898 -1663 0 net=6795
rlabel metal2 72 -1665 72 -1665 0 net=1967
rlabel metal2 156 -1665 156 -1665 0 net=1733
rlabel metal2 191 -1665 191 -1665 0 net=2550
rlabel metal2 961 -1665 961 -1665 0 net=6929
rlabel metal2 72 -1667 72 -1667 0 net=1205
rlabel metal2 191 -1667 191 -1667 0 net=1831
rlabel metal2 226 -1667 226 -1667 0 net=2409
rlabel metal2 254 -1667 254 -1667 0 net=1581
rlabel metal2 296 -1667 296 -1667 0 net=2482
rlabel metal2 387 -1667 387 -1667 0 net=2319
rlabel metal2 422 -1667 422 -1667 0 net=1038
rlabel metal2 681 -1667 681 -1667 0 net=6653
rlabel metal2 821 -1667 821 -1667 0 net=6603
rlabel metal2 86 -1669 86 -1669 0 net=1497
rlabel metal2 240 -1669 240 -1669 0 net=2375
rlabel metal2 387 -1669 387 -1669 0 net=4063
rlabel metal2 597 -1669 597 -1669 0 net=4797
rlabel metal2 695 -1669 695 -1669 0 net=5565
rlabel metal2 842 -1669 842 -1669 0 net=6367
rlabel metal2 919 -1669 919 -1669 0 net=7259
rlabel metal2 65 -1671 65 -1671 0 net=1168
rlabel metal2 702 -1671 702 -1671 0 net=5837
rlabel metal2 842 -1671 842 -1671 0 net=6683
rlabel metal2 163 -1673 163 -1673 0 net=4849
rlabel metal2 296 -1673 296 -1673 0 net=2227
rlabel metal2 317 -1673 317 -1673 0 net=1792
rlabel metal2 366 -1673 366 -1673 0 net=3021
rlabel metal2 618 -1673 618 -1673 0 net=3984
rlabel metal2 163 -1675 163 -1675 0 net=5323
rlabel metal2 422 -1675 422 -1675 0 net=438
rlabel metal2 618 -1675 618 -1675 0 net=4953
rlabel metal2 702 -1675 702 -1675 0 net=5717
rlabel metal2 954 -1675 954 -1675 0 net=7727
rlabel metal2 201 -1677 201 -1677 0 net=4587
rlabel metal2 425 -1677 425 -1677 0 net=4986
rlabel metal2 205 -1679 205 -1679 0 net=1923
rlabel metal2 317 -1679 317 -1679 0 net=3239
rlabel metal2 429 -1679 429 -1679 0 net=2801
rlabel metal2 457 -1679 457 -1679 0 net=7389
rlabel metal2 471 -1679 471 -1679 0 net=5987
rlabel metal2 716 -1679 716 -1679 0 net=5673
rlabel metal2 807 -1679 807 -1679 0 net=6865
rlabel metal2 212 -1681 212 -1681 0 net=3463
rlabel metal2 464 -1681 464 -1681 0 net=2233
rlabel metal2 625 -1681 625 -1681 0 net=5019
rlabel metal2 730 -1681 730 -1681 0 net=6637
rlabel metal2 233 -1683 233 -1683 0 net=3184
rlabel metal2 327 -1683 327 -1683 0 net=5608
rlabel metal2 905 -1683 905 -1683 0 net=6746
rlabel metal2 184 -1685 184 -1685 0 net=7641
rlabel metal2 933 -1685 933 -1685 0 net=7535
rlabel metal2 44 -1687 44 -1687 0 net=2063
rlabel metal2 233 -1687 233 -1687 0 net=1997
rlabel metal2 359 -1687 359 -1687 0 net=5181
rlabel metal2 632 -1687 632 -1687 0 net=5995
rlabel metal2 709 -1687 709 -1687 0 net=6227
rlabel metal2 744 -1687 744 -1687 0 net=7007
rlabel metal2 940 -1687 940 -1687 0 net=7417
rlabel metal2 44 -1689 44 -1689 0 net=1981
rlabel metal2 268 -1689 268 -1689 0 net=2663
rlabel metal2 373 -1689 373 -1689 0 net=856
rlabel metal2 471 -1689 471 -1689 0 net=3119
rlabel metal2 513 -1689 513 -1689 0 net=3671
rlabel metal2 639 -1689 639 -1689 0 net=4577
rlabel metal2 737 -1689 737 -1689 0 net=6505
rlabel metal2 268 -1691 268 -1691 0 net=2531
rlabel metal2 373 -1691 373 -1691 0 net=5510
rlabel metal2 877 -1691 877 -1691 0 net=7589
rlabel metal2 415 -1693 415 -1693 0 net=3353
rlabel metal2 646 -1693 646 -1693 0 net=5309
rlabel metal2 723 -1693 723 -1693 0 net=5171
rlabel metal2 408 -1695 408 -1695 0 net=2130
rlabel metal2 723 -1695 723 -1695 0 net=5911
rlabel metal2 408 -1697 408 -1697 0 net=4741
rlabel metal2 744 -1697 744 -1697 0 net=5969
rlabel metal2 478 -1699 478 -1699 0 net=4485
rlabel metal2 751 -1699 751 -1699 0 net=7620
rlabel metal2 30 -1701 30 -1701 0 net=4398
rlabel metal2 481 -1701 481 -1701 0 net=4531
rlabel metal2 800 -1701 800 -1701 0 net=6841
rlabel metal2 30 -1703 30 -1703 0 net=2139
rlabel metal2 488 -1703 488 -1703 0 net=7041
rlabel metal2 968 -1703 968 -1703 0 net=7001
rlabel metal2 121 -1705 121 -1705 0 net=1989
rlabel metal2 499 -1705 499 -1705 0 net=3509
rlabel metal2 282 -1707 282 -1707 0 net=2087
rlabel metal2 548 -1707 548 -1707 0 net=3423
rlabel metal2 275 -1709 275 -1709 0 net=1973
rlabel metal2 555 -1709 555 -1709 0 net=2437
rlabel metal2 856 -1711 856 -1711 0 net=7227
rlabel metal2 2 -1722 2 -1722 0 net=3465
rlabel metal2 254 -1722 254 -1722 0 net=1582
rlabel metal2 338 -1722 338 -1722 0 net=1573
rlabel metal2 653 -1722 653 -1722 0 net=6486
rlabel metal2 849 -1722 849 -1722 0 net=7643
rlabel metal2 1052 -1722 1052 -1722 0 net=936
rlabel metal2 1094 -1722 1094 -1722 0 net=6215
rlabel metal2 1094 -1722 1094 -1722 0 net=6215
rlabel metal2 16 -1724 16 -1724 0 net=3263
rlabel metal2 51 -1724 51 -1724 0 net=1419
rlabel metal2 100 -1724 100 -1724 0 net=1708
rlabel metal2 159 -1724 159 -1724 0 net=2376
rlabel metal2 261 -1724 261 -1724 0 net=4851
rlabel metal2 870 -1724 870 -1724 0 net=5668
rlabel metal2 919 -1724 919 -1724 0 net=7261
rlabel metal2 1055 -1724 1055 -1724 0 net=6127
rlabel metal2 30 -1726 30 -1726 0 net=2140
rlabel metal2 226 -1726 226 -1726 0 net=2411
rlabel metal2 275 -1726 275 -1726 0 net=1975
rlabel metal2 359 -1726 359 -1726 0 net=1801
rlabel metal2 527 -1726 527 -1726 0 net=6638
rlabel metal2 758 -1726 758 -1726 0 net=6867
rlabel metal2 817 -1726 817 -1726 0 net=7536
rlabel metal2 940 -1726 940 -1726 0 net=7419
rlabel metal2 23 -1728 23 -1728 0 net=6232
rlabel metal2 233 -1728 233 -1728 0 net=1999
rlabel metal2 275 -1728 275 -1728 0 net=2089
rlabel metal2 296 -1728 296 -1728 0 net=2228
rlabel metal2 366 -1728 366 -1728 0 net=3022
rlabel metal2 436 -1728 436 -1728 0 net=2802
rlabel metal2 527 -1728 527 -1728 0 net=4798
rlabel metal2 632 -1728 632 -1728 0 net=7043
rlabel metal2 926 -1728 926 -1728 0 net=6930
rlabel metal2 30 -1730 30 -1730 0 net=2031
rlabel metal2 681 -1730 681 -1730 0 net=5997
rlabel metal2 828 -1730 828 -1730 0 net=6369
rlabel metal2 877 -1730 877 -1730 0 net=7591
rlabel metal2 37 -1732 37 -1732 0 net=1983
rlabel metal2 65 -1732 65 -1732 0 net=7390
rlabel metal2 478 -1732 478 -1732 0 net=2929
rlabel metal2 761 -1732 761 -1732 0 net=3095
rlabel metal2 44 -1734 44 -1734 0 net=1991
rlabel metal2 170 -1734 170 -1734 0 net=1735
rlabel metal2 170 -1734 170 -1734 0 net=1735
rlabel metal2 177 -1734 177 -1734 0 net=3695
rlabel metal2 177 -1734 177 -1734 0 net=3695
rlabel metal2 212 -1734 212 -1734 0 net=3241
rlabel metal2 366 -1734 366 -1734 0 net=3451
rlabel metal2 408 -1734 408 -1734 0 net=4743
rlabel metal2 660 -1734 660 -1734 0 net=7491
rlabel metal2 65 -1736 65 -1736 0 net=1925
rlabel metal2 219 -1736 219 -1736 0 net=2961
rlabel metal2 380 -1736 380 -1736 0 net=2235
rlabel metal2 495 -1736 495 -1736 0 net=3510
rlabel metal2 534 -1736 534 -1736 0 net=4103
rlabel metal2 674 -1736 674 -1736 0 net=7228
rlabel metal2 863 -1736 863 -1736 0 net=6965
rlabel metal2 926 -1736 926 -1736 0 net=7689
rlabel metal2 954 -1736 954 -1736 0 net=7729
rlabel metal2 79 -1738 79 -1738 0 net=3788
rlabel metal2 408 -1738 408 -1738 0 net=1653
rlabel metal2 506 -1738 506 -1738 0 net=3557
rlabel metal2 586 -1738 586 -1738 0 net=5793
rlabel metal2 779 -1738 779 -1738 0 net=5839
rlabel metal2 779 -1738 779 -1738 0 net=5839
rlabel metal2 793 -1738 793 -1738 0 net=7009
rlabel metal2 929 -1738 929 -1738 0 net=7205
rlabel metal2 79 -1740 79 -1740 0 net=4131
rlabel metal2 425 -1740 425 -1740 0 net=6275
rlabel metal2 667 -1740 667 -1740 0 net=5989
rlabel metal2 891 -1740 891 -1740 0 net=7113
rlabel metal2 947 -1740 947 -1740 0 net=7003
rlabel metal2 86 -1742 86 -1742 0 net=1498
rlabel metal2 443 -1742 443 -1742 0 net=7739
rlabel metal2 86 -1744 86 -1744 0 net=1969
rlabel metal2 121 -1744 121 -1744 0 net=1943
rlabel metal2 443 -1744 443 -1744 0 net=3395
rlabel metal2 597 -1744 597 -1744 0 net=5020
rlabel metal2 667 -1744 667 -1744 0 net=5172
rlabel metal2 842 -1744 842 -1744 0 net=6685
rlabel metal2 891 -1744 891 -1744 0 net=6797
rlabel metal2 905 -1744 905 -1744 0 net=7771
rlabel metal2 100 -1746 100 -1746 0 net=2664
rlabel metal2 296 -1746 296 -1746 0 net=4473
rlabel metal2 450 -1746 450 -1746 0 net=4187
rlabel metal2 670 -1746 670 -1746 0 net=7211
rlabel metal2 107 -1748 107 -1748 0 net=2786
rlabel metal2 156 -1748 156 -1748 0 net=4811
rlabel metal2 681 -1748 681 -1748 0 net=6229
rlabel metal2 716 -1748 716 -1748 0 net=5675
rlabel metal2 135 -1750 135 -1750 0 net=5805
rlabel metal2 800 -1750 800 -1750 0 net=6843
rlabel metal2 23 -1752 23 -1752 0 net=3393
rlabel metal2 142 -1752 142 -1752 0 net=1833
rlabel metal2 198 -1752 198 -1752 0 net=1942
rlabel metal2 506 -1752 506 -1752 0 net=5311
rlabel metal2 688 -1752 688 -1752 0 net=6206
rlabel metal2 156 -1754 156 -1754 0 net=4065
rlabel metal2 450 -1754 450 -1754 0 net=3215
rlabel metal2 569 -1754 569 -1754 0 net=5183
rlabel metal2 688 -1754 688 -1754 0 net=6604
rlabel metal2 163 -1756 163 -1756 0 net=5325
rlabel metal2 723 -1756 723 -1756 0 net=5913
rlabel metal2 149 -1758 149 -1758 0 net=5531
rlabel metal2 730 -1758 730 -1758 0 net=5423
rlabel metal2 149 -1760 149 -1760 0 net=2118
rlabel metal2 348 -1760 348 -1760 0 net=5857
rlabel metal2 163 -1762 163 -1762 0 net=2065
rlabel metal2 191 -1762 191 -1762 0 net=2853
rlabel metal2 702 -1762 702 -1762 0 net=5719
rlabel metal2 114 -1764 114 -1764 0 net=2122
rlabel metal2 198 -1764 198 -1764 0 net=7637
rlabel metal2 226 -1766 226 -1766 0 net=1871
rlabel metal2 457 -1766 457 -1766 0 net=5223
rlabel metal2 625 -1766 625 -1766 0 net=5899
rlabel metal2 233 -1768 233 -1768 0 net=2217
rlabel metal2 373 -1768 373 -1768 0 net=2341
rlabel metal2 576 -1768 576 -1768 0 net=7309
rlabel metal2 128 -1770 128 -1770 0 net=4803
rlabel metal2 387 -1770 387 -1770 0 net=2269
rlabel metal2 464 -1770 464 -1770 0 net=3673
rlabel metal2 611 -1770 611 -1770 0 net=7407
rlabel metal2 128 -1772 128 -1772 0 net=1225
rlabel metal2 268 -1772 268 -1772 0 net=2532
rlabel metal2 306 -1772 306 -1772 0 net=3025
rlabel metal2 485 -1772 485 -1772 0 net=5609
rlabel metal2 639 -1772 639 -1772 0 net=4579
rlabel metal2 737 -1772 737 -1772 0 net=6507
rlabel metal2 240 -1774 240 -1774 0 net=1433
rlabel metal2 618 -1774 618 -1774 0 net=4955
rlabel metal2 695 -1774 695 -1774 0 net=5567
rlabel metal2 744 -1774 744 -1774 0 net=5971
rlabel metal2 268 -1776 268 -1776 0 net=2163
rlabel metal2 352 -1776 352 -1776 0 net=4745
rlabel metal2 492 -1776 492 -1776 0 net=5785
rlabel metal2 765 -1776 765 -1776 0 net=6655
rlabel metal2 58 -1778 58 -1778 0 net=3255
rlabel metal2 352 -1778 352 -1778 0 net=5349
rlabel metal2 600 -1778 600 -1778 0 net=5333
rlabel metal2 712 -1778 712 -1778 0 net=646
rlabel metal2 58 -1780 58 -1780 0 net=1207
rlabel metal2 282 -1780 282 -1780 0 net=2321
rlabel metal2 415 -1780 415 -1780 0 net=3355
rlabel metal2 72 -1782 72 -1782 0 net=3699
rlabel metal2 289 -1782 289 -1782 0 net=2691
rlabel metal2 362 -1782 362 -1782 0 net=4189
rlabel metal2 394 -1784 394 -1784 0 net=4589
rlabel metal2 394 -1786 394 -1786 0 net=4315
rlabel metal2 401 -1788 401 -1788 0 net=2439
rlabel metal2 415 -1790 415 -1790 0 net=3120
rlabel metal2 555 -1790 555 -1790 0 net=4373
rlabel metal2 429 -1792 429 -1792 0 net=7151
rlabel metal2 471 -1794 471 -1794 0 net=4533
rlabel metal2 590 -1794 590 -1794 0 net=4649
rlabel metal2 541 -1796 541 -1796 0 net=4487
rlabel metal2 604 -1796 604 -1796 0 net=6663
rlabel metal2 541 -1798 541 -1798 0 net=3425
rlabel metal2 548 -1800 548 -1800 0 net=6154
rlabel metal2 117 -1802 117 -1802 0 net=6759
rlabel metal2 2 -1813 2 -1813 0 net=3466
rlabel metal2 443 -1813 443 -1813 0 net=3397
rlabel metal2 499 -1813 499 -1813 0 net=5720
rlabel metal2 933 -1813 933 -1813 0 net=7004
rlabel metal2 968 -1813 968 -1813 0 net=7311
rlabel metal2 968 -1813 968 -1813 0 net=7311
rlabel metal2 1010 -1813 1010 -1813 0 net=7639
rlabel metal2 1087 -1813 1087 -1813 0 net=6129
rlabel metal2 5 -1815 5 -1815 0 net=834
rlabel metal2 555 -1815 555 -1815 0 net=4374
rlabel metal2 555 -1815 555 -1815 0 net=4374
rlabel metal2 604 -1815 604 -1815 0 net=4580
rlabel metal2 709 -1815 709 -1815 0 net=7262
rlabel metal2 1017 -1815 1017 -1815 0 net=7645
rlabel metal2 1087 -1815 1087 -1815 0 net=6217
rlabel metal2 37 -1817 37 -1817 0 net=1984
rlabel metal2 54 -1817 54 -1817 0 net=3700
rlabel metal2 79 -1817 79 -1817 0 net=4132
rlabel metal2 443 -1817 443 -1817 0 net=3356
rlabel metal2 502 -1817 502 -1817 0 net=4744
rlabel metal2 667 -1817 667 -1817 0 net=6868
rlabel metal2 828 -1817 828 -1817 0 net=6371
rlabel metal2 828 -1817 828 -1817 0 net=6371
rlabel metal2 912 -1817 912 -1817 0 net=7011
rlabel metal2 975 -1817 975 -1817 0 net=7409
rlabel metal2 1024 -1817 1024 -1817 0 net=7731
rlabel metal2 1024 -1817 1024 -1817 0 net=7731
rlabel metal2 1045 -1817 1045 -1817 0 net=3096
rlabel metal2 47 -1819 47 -1819 0 net=1909
rlabel metal2 93 -1819 93 -1819 0 net=4852
rlabel metal2 891 -1819 891 -1819 0 net=6799
rlabel metal2 926 -1819 926 -1819 0 net=7691
rlabel metal2 58 -1821 58 -1821 0 net=1209
rlabel metal2 58 -1821 58 -1821 0 net=1209
rlabel metal2 103 -1821 103 -1821 0 net=2342
rlabel metal2 387 -1821 387 -1821 0 net=2270
rlabel metal2 646 -1821 646 -1821 0 net=5185
rlabel metal2 891 -1821 891 -1821 0 net=7115
rlabel metal2 954 -1821 954 -1821 0 net=7153
rlabel metal2 114 -1823 114 -1823 0 net=2412
rlabel metal2 268 -1823 268 -1823 0 net=2164
rlabel metal2 373 -1823 373 -1823 0 net=2323
rlabel metal2 733 -1823 733 -1823 0 net=6844
rlabel metal2 919 -1823 919 -1823 0 net=7045
rlabel metal2 93 -1825 93 -1825 0 net=3541
rlabel metal2 121 -1825 121 -1825 0 net=1945
rlabel metal2 198 -1825 198 -1825 0 net=5806
rlabel metal2 863 -1825 863 -1825 0 net=6967
rlabel metal2 121 -1827 121 -1827 0 net=4188
rlabel metal2 590 -1827 590 -1827 0 net=4651
rlabel metal2 688 -1827 688 -1827 0 net=917
rlabel metal2 124 -1829 124 -1829 0 net=1059
rlabel metal2 226 -1829 226 -1829 0 net=1872
rlabel metal2 429 -1829 429 -1829 0 net=7137
rlabel metal2 135 -1831 135 -1831 0 net=7605
rlabel metal2 135 -1833 135 -1833 0 net=2855
rlabel metal2 194 -1833 194 -1833 0 net=4293
rlabel metal2 611 -1833 611 -1833 0 net=4375
rlabel metal2 611 -1833 611 -1833 0 net=4375
rlabel metal2 614 -1833 614 -1833 0 net=5914
rlabel metal2 877 -1833 877 -1833 0 net=6687
rlabel metal2 163 -1835 163 -1835 0 net=2066
rlabel metal2 366 -1835 366 -1835 0 net=3453
rlabel metal2 884 -1835 884 -1835 0 net=6761
rlabel metal2 163 -1837 163 -1837 0 net=1865
rlabel metal2 569 -1837 569 -1837 0 net=5351
rlabel metal2 737 -1837 737 -1837 0 net=5569
rlabel metal2 898 -1837 898 -1837 0 net=7213
rlabel metal2 198 -1839 198 -1839 0 net=1803
rlabel metal2 394 -1839 394 -1839 0 net=4317
rlabel metal2 628 -1839 628 -1839 0 net=6230
rlabel metal2 695 -1839 695 -1839 0 net=5335
rlabel metal2 723 -1839 723 -1839 0 net=5533
rlabel metal2 751 -1839 751 -1839 0 net=5795
rlabel metal2 765 -1839 765 -1839 0 net=6689
rlabel metal2 201 -1841 201 -1841 0 net=1449
rlabel metal2 282 -1841 282 -1841 0 net=2322
rlabel metal2 401 -1841 401 -1841 0 net=2441
rlabel metal2 401 -1841 401 -1841 0 net=2441
rlabel metal2 415 -1841 415 -1841 0 net=6235
rlabel metal2 772 -1841 772 -1841 0 net=6509
rlabel metal2 208 -1843 208 -1843 0 net=2218
rlabel metal2 250 -1843 250 -1843 0 net=4190
rlabel metal2 695 -1843 695 -1843 0 net=5327
rlabel metal2 723 -1843 723 -1843 0 net=5901
rlabel metal2 814 -1843 814 -1843 0 net=5999
rlabel metal2 842 -1843 842 -1843 0 net=6665
rlabel metal2 226 -1845 226 -1845 0 net=5481
rlabel metal2 576 -1845 576 -1845 0 net=5611
rlabel metal2 800 -1845 800 -1845 0 net=5973
rlabel metal2 814 -1845 814 -1845 0 net=5677
rlabel metal2 233 -1847 233 -1847 0 net=4535
rlabel metal2 481 -1847 481 -1847 0 net=5383
rlabel metal2 730 -1847 730 -1847 0 net=5425
rlabel metal2 786 -1847 786 -1847 0 net=5859
rlabel metal2 1031 -1847 1031 -1847 0 net=7741
rlabel metal2 254 -1849 254 -1849 0 net=2000
rlabel metal2 366 -1849 366 -1849 0 net=4153
rlabel metal2 583 -1849 583 -1849 0 net=4147
rlabel metal2 691 -1849 691 -1849 0 net=7185
rlabel metal2 989 -1849 989 -1849 0 net=7493
rlabel metal2 100 -1851 100 -1851 0 net=2947
rlabel metal2 261 -1851 261 -1851 0 net=3027
rlabel metal2 457 -1851 457 -1851 0 net=5225
rlabel metal2 744 -1851 744 -1851 0 net=5787
rlabel metal2 779 -1851 779 -1851 0 net=5841
rlabel metal2 961 -1851 961 -1851 0 net=7207
rlabel metal2 100 -1853 100 -1853 0 net=3595
rlabel metal2 282 -1853 282 -1853 0 net=1655
rlabel metal2 418 -1853 418 -1853 0 net=3029
rlabel metal2 436 -1853 436 -1853 0 net=3311
rlabel metal2 835 -1853 835 -1853 0 net=6657
rlabel metal2 149 -1855 149 -1855 0 net=3099
rlabel metal2 485 -1855 485 -1855 0 net=4747
rlabel metal2 23 -1857 23 -1857 0 net=3394
rlabel metal2 488 -1857 488 -1857 0 net=5629
rlabel metal2 23 -1859 23 -1859 0 net=4804
rlabel metal2 317 -1859 317 -1859 0 net=2963
rlabel metal2 352 -1859 352 -1859 0 net=3675
rlabel metal2 492 -1859 492 -1859 0 net=5313
rlabel metal2 520 -1859 520 -1859 0 net=5990
rlabel metal2 65 -1861 65 -1861 0 net=1927
rlabel metal2 317 -1861 317 -1861 0 net=1425
rlabel metal2 394 -1861 394 -1861 0 net=2565
rlabel metal2 65 -1863 65 -1863 0 net=234
rlabel metal2 205 -1863 205 -1863 0 net=1435
rlabel metal2 296 -1863 296 -1863 0 net=4474
rlabel metal2 562 -1863 562 -1863 0 net=4489
rlabel metal2 632 -1863 632 -1863 0 net=6277
rlabel metal2 79 -1865 79 -1865 0 net=6441
rlabel metal2 534 -1865 534 -1865 0 net=3559
rlabel metal2 569 -1865 569 -1865 0 net=3839
rlabel metal2 117 -1867 117 -1867 0 net=2939
rlabel metal2 303 -1867 303 -1867 0 net=2237
rlabel metal2 408 -1867 408 -1867 0 net=1405
rlabel metal2 450 -1867 450 -1867 0 net=3217
rlabel metal2 621 -1867 621 -1867 0 net=6939
rlabel metal2 117 -1869 117 -1869 0 net=1574
rlabel metal2 450 -1869 450 -1869 0 net=4247
rlabel metal2 632 -1869 632 -1869 0 net=7772
rlabel metal2 16 -1871 16 -1871 0 net=3265
rlabel metal2 639 -1871 639 -1871 0 net=4957
rlabel metal2 1003 -1871 1003 -1871 0 net=7593
rlabel metal2 128 -1873 128 -1873 0 net=1227
rlabel metal2 306 -1873 306 -1873 0 net=4812
rlabel metal2 982 -1873 982 -1873 0 net=7421
rlabel metal2 86 -1875 86 -1875 0 net=1971
rlabel metal2 177 -1875 177 -1875 0 net=3697
rlabel metal2 548 -1875 548 -1875 0 net=6397
rlabel metal2 86 -1877 86 -1877 0 net=5541
rlabel metal2 289 -1877 289 -1877 0 net=2693
rlabel metal2 422 -1877 422 -1877 0 net=7159
rlabel metal2 9 -1879 9 -1879 0 net=2937
rlabel metal2 513 -1879 513 -1879 0 net=4591
rlabel metal2 9 -1881 9 -1881 0 net=2331
rlabel metal2 142 -1881 142 -1881 0 net=1835
rlabel metal2 212 -1881 212 -1881 0 net=3243
rlabel metal2 275 -1881 275 -1881 0 net=2091
rlabel metal2 324 -1881 324 -1881 0 net=1976
rlabel metal2 513 -1881 513 -1881 0 net=3427
rlabel metal2 96 -1883 96 -1883 0 net=2039
rlabel metal2 156 -1883 156 -1883 0 net=4067
rlabel metal2 331 -1883 331 -1883 0 net=3257
rlabel metal2 30 -1885 30 -1885 0 net=2032
rlabel metal2 170 -1885 170 -1885 0 net=1737
rlabel metal2 331 -1885 331 -1885 0 net=2931
rlabel metal2 30 -1887 30 -1887 0 net=1993
rlabel metal2 107 -1887 107 -1887 0 net=1607
rlabel metal2 390 -1887 390 -1887 0 net=3659
rlabel metal2 44 -1889 44 -1889 0 net=7757
rlabel metal2 51 -1891 51 -1891 0 net=1421
rlabel metal2 170 -1891 170 -1891 0 net=5107
rlabel metal2 478 -1891 478 -1891 0 net=4104
rlabel metal2 51 -1893 51 -1893 0 net=593
rlabel metal2 551 -1893 551 -1893 0 net=5697
rlabel metal2 2 -1904 2 -1904 0 net=710
rlabel metal2 530 -1904 530 -1904 0 net=7494
rlabel metal2 1073 -1904 1073 -1904 0 net=7647
rlabel metal2 9 -1906 9 -1906 0 net=2332
rlabel metal2 44 -1906 44 -1906 0 net=1972
rlabel metal2 142 -1906 142 -1906 0 net=2041
rlabel metal2 194 -1906 194 -1906 0 net=5314
rlabel metal2 502 -1906 502 -1906 0 net=3698
rlabel metal2 551 -1906 551 -1906 0 net=5570
rlabel metal2 1003 -1906 1003 -1906 0 net=7423
rlabel metal2 1045 -1906 1045 -1906 0 net=7759
rlabel metal2 1080 -1906 1080 -1906 0 net=6219
rlabel metal2 1101 -1906 1101 -1906 0 net=6131
rlabel metal2 9 -1908 9 -1908 0 net=3597
rlabel metal2 114 -1908 114 -1908 0 net=2857
rlabel metal2 149 -1908 149 -1908 0 net=1450
rlabel metal2 296 -1908 296 -1908 0 net=1228
rlabel metal2 369 -1908 369 -1908 0 net=5336
rlabel metal2 786 -1908 786 -1908 0 net=5843
rlabel metal2 786 -1908 786 -1908 0 net=5843
rlabel metal2 821 -1908 821 -1908 0 net=6001
rlabel metal2 842 -1908 842 -1908 0 net=5860
rlabel metal2 16 -1910 16 -1910 0 net=1985
rlabel metal2 485 -1910 485 -1910 0 net=5328
rlabel metal2 702 -1910 702 -1910 0 net=3047
rlabel metal2 19 -1912 19 -1912 0 net=2938
rlabel metal2 429 -1912 429 -1912 0 net=3031
rlabel metal2 429 -1912 429 -1912 0 net=3031
rlabel metal2 443 -1912 443 -1912 0 net=4319
rlabel metal2 618 -1912 618 -1912 0 net=6762
rlabel metal2 968 -1912 968 -1912 0 net=7313
rlabel metal2 1024 -1912 1024 -1912 0 net=7733
rlabel metal2 30 -1914 30 -1914 0 net=1994
rlabel metal2 30 -1914 30 -1914 0 net=1994
rlabel metal2 33 -1914 33 -1914 0 net=7595
rlabel metal2 37 -1916 37 -1916 0 net=2567
rlabel metal2 450 -1916 450 -1916 0 net=3101
rlabel metal2 471 -1916 471 -1916 0 net=3259
rlabel metal2 516 -1916 516 -1916 0 net=5186
rlabel metal2 968 -1916 968 -1916 0 net=7411
rlabel metal2 47 -1918 47 -1918 0 net=7154
rlabel metal2 51 -1920 51 -1920 0 net=1210
rlabel metal2 65 -1920 65 -1920 0 net=1911
rlabel metal2 75 -1920 75 -1920 0 net=1115
rlabel metal2 527 -1920 527 -1920 0 net=7594
rlabel metal2 58 -1922 58 -1922 0 net=4253
rlabel metal2 453 -1922 453 -1922 0 net=5807
rlabel metal2 82 -1924 82 -1924 0 net=3244
rlabel metal2 324 -1924 324 -1924 0 net=4069
rlabel metal2 618 -1924 618 -1924 0 net=6278
rlabel metal2 870 -1924 870 -1924 0 net=7013
rlabel metal2 947 -1924 947 -1924 0 net=7139
rlabel metal2 93 -1926 93 -1926 0 net=3543
rlabel metal2 555 -1926 555 -1926 0 net=5631
rlabel metal2 768 -1926 768 -1926 0 net=6727
rlabel metal2 926 -1926 926 -1926 0 net=6969
rlabel metal2 954 -1926 954 -1926 0 net=7215
rlabel metal2 93 -1928 93 -1928 0 net=1615
rlabel metal2 222 -1928 222 -1928 0 net=2092
rlabel metal2 324 -1928 324 -1928 0 net=3219
rlabel metal2 471 -1928 471 -1928 0 net=3399
rlabel metal2 558 -1928 558 -1928 0 net=6417
rlabel metal2 856 -1928 856 -1928 0 net=6975
rlabel metal2 100 -1930 100 -1930 0 net=2965
rlabel metal2 348 -1930 348 -1930 0 net=1406
rlabel metal2 478 -1930 478 -1930 0 net=3323
rlabel metal2 478 -1930 478 -1930 0 net=3323
rlabel metal2 485 -1930 485 -1930 0 net=4155
rlabel metal2 621 -1930 621 -1930 0 net=5612
rlabel metal2 821 -1930 821 -1930 0 net=6373
rlabel metal2 912 -1930 912 -1930 0 net=6801
rlabel metal2 940 -1930 940 -1930 0 net=7047
rlabel metal2 124 -1932 124 -1932 0 net=7742
rlabel metal2 128 -1934 128 -1934 0 net=2265
rlabel metal2 387 -1934 387 -1934 0 net=2443
rlabel metal2 506 -1934 506 -1934 0 net=5535
rlabel metal2 835 -1934 835 -1934 0 net=6941
rlabel metal2 1010 -1934 1010 -1934 0 net=7607
rlabel metal2 152 -1936 152 -1936 0 net=3454
rlabel metal2 898 -1936 898 -1936 0 net=6691
rlabel metal2 23 -1938 23 -1938 0 net=6487
rlabel metal2 44 -1940 44 -1940 0 net=3133
rlabel metal2 156 -1940 156 -1940 0 net=5833
rlabel metal2 877 -1940 877 -1940 0 net=7117
rlabel metal2 107 -1942 107 -1942 0 net=1423
rlabel metal2 159 -1942 159 -1942 0 net=4607
rlabel metal2 107 -1944 107 -1944 0 net=2095
rlabel metal2 184 -1944 184 -1944 0 net=1947
rlabel metal2 338 -1944 338 -1944 0 net=3267
rlabel metal2 562 -1944 562 -1944 0 net=3561
rlabel metal2 562 -1944 562 -1944 0 net=3561
rlabel metal2 576 -1944 576 -1944 0 net=4377
rlabel metal2 621 -1944 621 -1944 0 net=7640
rlabel metal2 184 -1946 184 -1946 0 net=2909
rlabel metal2 369 -1946 369 -1946 0 net=740
rlabel metal2 583 -1946 583 -1946 0 net=4149
rlabel metal2 632 -1946 632 -1946 0 net=7515
rlabel metal2 198 -1948 198 -1948 0 net=1805
rlabel metal2 338 -1948 338 -1948 0 net=4653
rlabel metal2 660 -1948 660 -1948 0 net=5699
rlabel metal2 1017 -1948 1017 -1948 0 net=7693
rlabel metal2 198 -1950 198 -1950 0 net=1657
rlabel metal2 345 -1950 345 -1950 0 net=2987
rlabel metal2 569 -1950 569 -1950 0 net=3841
rlabel metal2 635 -1950 635 -1950 0 net=5902
rlabel metal2 989 -1950 989 -1950 0 net=7209
rlabel metal2 23 -1952 23 -1952 0 net=5393
rlabel metal2 807 -1952 807 -1952 0 net=7187
rlabel metal2 54 -1954 54 -1954 0 net=4051
rlabel metal2 635 -1954 635 -1954 0 net=5426
rlabel metal2 807 -1954 807 -1954 0 net=6667
rlabel metal2 54 -1956 54 -1956 0 net=5482
rlabel metal2 229 -1956 229 -1956 0 net=1595
rlabel metal2 352 -1956 352 -1956 0 net=3676
rlabel metal2 646 -1956 646 -1956 0 net=6688
rlabel metal2 180 -1958 180 -1958 0 net=3641
rlabel metal2 625 -1958 625 -1958 0 net=4491
rlabel metal2 117 -1960 117 -1960 0 net=7383
rlabel metal2 660 -1960 660 -1960 0 net=4959
rlabel metal2 863 -1960 863 -1960 0 net=6511
rlabel metal2 208 -1962 208 -1962 0 net=7160
rlabel metal2 149 -1964 149 -1964 0 net=7155
rlabel metal2 222 -1966 222 -1966 0 net=3028
rlabel metal2 275 -1966 275 -1966 0 net=1609
rlabel metal2 331 -1966 331 -1966 0 net=2933
rlabel metal2 359 -1966 359 -1966 0 net=7393
rlabel metal2 163 -1968 163 -1968 0 net=1867
rlabel metal2 331 -1968 331 -1968 0 net=2325
rlabel metal2 390 -1968 390 -1968 0 net=6533
rlabel metal2 163 -1970 163 -1970 0 net=2839
rlabel metal2 670 -1970 670 -1970 0 net=4493
rlabel metal2 240 -1972 240 -1972 0 net=2941
rlabel metal2 681 -1972 681 -1972 0 net=5227
rlabel metal2 751 -1972 751 -1972 0 net=6237
rlabel metal2 240 -1974 240 -1974 0 net=2949
rlabel metal2 359 -1974 359 -1974 0 net=2695
rlabel metal2 667 -1974 667 -1974 0 net=5087
rlabel metal2 688 -1974 688 -1974 0 net=6658
rlabel metal2 86 -1976 86 -1976 0 net=5543
rlabel metal2 520 -1976 520 -1976 0 net=6443
rlabel metal2 674 -1976 674 -1976 0 net=6399
rlabel metal2 61 -1978 61 -1978 0 net=3833
rlabel metal2 597 -1978 597 -1978 0 net=4249
rlabel metal2 695 -1978 695 -1978 0 net=5353
rlabel metal2 751 -1978 751 -1978 0 net=5679
rlabel metal2 233 -1980 233 -1980 0 net=4537
rlabel metal2 649 -1980 649 -1980 0 net=7599
rlabel metal2 212 -1982 212 -1982 0 net=1739
rlabel metal2 247 -1982 247 -1982 0 net=2911
rlabel metal2 758 -1982 758 -1982 0 net=5797
rlabel metal2 121 -1984 121 -1984 0 net=2515
rlabel metal2 254 -1984 254 -1984 0 net=2239
rlabel metal2 373 -1984 373 -1984 0 net=4655
rlabel metal2 653 -1984 653 -1984 0 net=4749
rlabel metal2 709 -1984 709 -1984 0 net=5385
rlabel metal2 730 -1984 730 -1984 0 net=5975
rlabel metal2 121 -1986 121 -1986 0 net=1437
rlabel metal2 303 -1986 303 -1986 0 net=1929
rlabel metal2 548 -1986 548 -1986 0 net=6617
rlabel metal2 758 -1986 758 -1986 0 net=5789
rlabel metal2 170 -1988 170 -1988 0 net=5109
rlabel metal2 170 -1990 170 -1990 0 net=1837
rlabel metal2 205 -1990 205 -1990 0 net=3743
rlabel metal2 548 -1990 548 -1990 0 net=3957
rlabel metal2 310 -1992 310 -1992 0 net=3661
rlabel metal2 639 -1992 639 -1992 0 net=4593
rlabel metal2 317 -1994 317 -1994 0 net=1426
rlabel metal2 317 -1996 317 -1996 0 net=3313
rlabel metal2 513 -1996 513 -1996 0 net=3429
rlabel metal2 590 -1996 590 -1996 0 net=4295
rlabel metal2 261 -1998 261 -1998 0 net=2413
rlabel metal2 2 -2009 2 -2009 0 net=5031
rlabel metal2 229 -2009 229 -2009 0 net=488
rlabel metal2 376 -2009 376 -2009 0 net=6488
rlabel metal2 919 -2009 919 -2009 0 net=6729
rlabel metal2 919 -2009 919 -2009 0 net=6729
rlabel metal2 926 -2009 926 -2009 0 net=6803
rlabel metal2 943 -2009 943 -2009 0 net=7210
rlabel metal2 1080 -2009 1080 -2009 0 net=6220
rlabel metal2 1104 -2009 1104 -2009 0 net=7648
rlabel metal2 1115 -2009 1115 -2009 0 net=6133
rlabel metal2 9 -2011 9 -2011 0 net=3599
rlabel metal2 30 -2011 30 -2011 0 net=1785
rlabel metal2 30 -2011 30 -2011 0 net=1785
rlabel metal2 33 -2011 33 -2011 0 net=4608
rlabel metal2 1038 -2011 1038 -2011 0 net=7517
rlabel metal2 9 -2013 9 -2013 0 net=2841
rlabel metal2 170 -2013 170 -2013 0 net=1838
rlabel metal2 275 -2013 275 -2013 0 net=1869
rlabel metal2 439 -2013 439 -2013 0 net=5808
rlabel metal2 1073 -2013 1073 -2013 0 net=7761
rlabel metal2 16 -2015 16 -2015 0 net=1986
rlabel metal2 348 -2015 348 -2015 0 net=5110
rlabel metal2 807 -2015 807 -2015 0 net=6669
rlabel metal2 947 -2015 947 -2015 0 net=6971
rlabel metal2 947 -2015 947 -2015 0 net=6971
rlabel metal2 982 -2015 982 -2015 0 net=7157
rlabel metal2 1031 -2015 1031 -2015 0 net=7425
rlabel metal2 1045 -2015 1045 -2015 0 net=7597
rlabel metal2 16 -2017 16 -2017 0 net=2967
rlabel metal2 107 -2017 107 -2017 0 net=3842
rlabel metal2 593 -2017 593 -2017 0 net=6400
rlabel metal2 996 -2017 996 -2017 0 net=7217
rlabel metal2 1059 -2017 1059 -2017 0 net=7609
rlabel metal2 51 -2019 51 -2019 0 net=5834
rlabel metal2 863 -2019 863 -2019 0 net=6239
rlabel metal2 929 -2019 929 -2019 0 net=7412
rlabel metal2 1003 -2019 1003 -2019 0 net=7315
rlabel metal2 54 -2021 54 -2021 0 net=2917
rlabel metal2 380 -2021 380 -2021 0 net=5544
rlabel metal2 464 -2021 464 -2021 0 net=4656
rlabel metal2 688 -2021 688 -2021 0 net=4250
rlabel metal2 782 -2021 782 -2021 0 net=6374
rlabel metal2 835 -2021 835 -2021 0 net=6693
rlabel metal2 940 -2021 940 -2021 0 net=6943
rlabel metal2 975 -2021 975 -2021 0 net=7141
rlabel metal2 1010 -2021 1010 -2021 0 net=7395
rlabel metal2 37 -2023 37 -2023 0 net=2569
rlabel metal2 394 -2023 394 -2023 0 net=4255
rlabel metal2 691 -2023 691 -2023 0 net=7473
rlabel metal2 37 -2025 37 -2025 0 net=5981
rlabel metal2 180 -2025 180 -2025 0 net=1740
rlabel metal2 275 -2025 275 -2025 0 net=3401
rlabel metal2 502 -2025 502 -2025 0 net=4492
rlabel metal2 954 -2025 954 -2025 0 net=7049
rlabel metal2 44 -2027 44 -2027 0 net=3135
rlabel metal2 471 -2027 471 -2027 0 net=2905
rlabel metal2 569 -2027 569 -2027 0 net=4053
rlabel metal2 716 -2027 716 -2027 0 net=6619
rlabel metal2 44 -2029 44 -2029 0 net=2517
rlabel metal2 222 -2029 222 -2029 0 net=4070
rlabel metal2 611 -2029 611 -2029 0 net=4151
rlabel metal2 58 -2031 58 -2031 0 net=99
rlabel metal2 79 -2031 79 -2031 0 net=2049
rlabel metal2 177 -2031 177 -2031 0 net=1611
rlabel metal2 324 -2031 324 -2031 0 net=3220
rlabel metal2 394 -2031 394 -2031 0 net=3755
rlabel metal2 478 -2031 478 -2031 0 net=3325
rlabel metal2 625 -2031 625 -2031 0 net=7385
rlabel metal2 58 -2033 58 -2033 0 net=4494
rlabel metal2 870 -2033 870 -2033 0 net=7015
rlabel metal2 65 -2035 65 -2035 0 net=1912
rlabel metal2 408 -2035 408 -2035 0 net=3544
rlabel metal2 579 -2035 579 -2035 0 net=5685
rlabel metal2 821 -2035 821 -2035 0 net=6003
rlabel metal2 842 -2035 842 -2035 0 net=6419
rlabel metal2 877 -2035 877 -2035 0 net=7119
rlabel metal2 65 -2037 65 -2037 0 net=2267
rlabel metal2 135 -2037 135 -2037 0 net=3260
rlabel metal2 513 -2037 513 -2037 0 net=5395
rlabel metal2 744 -2037 744 -2037 0 net=5798
rlabel metal2 842 -2037 842 -2037 0 net=6535
rlabel metal2 51 -2039 51 -2039 0 net=2183
rlabel metal2 149 -2039 149 -2039 0 net=556
rlabel metal2 534 -2039 534 -2039 0 net=3563
rlabel metal2 667 -2039 667 -2039 0 net=6445
rlabel metal2 884 -2039 884 -2039 0 net=6513
rlabel metal2 72 -2041 72 -2041 0 net=1036
rlabel metal2 110 -2041 110 -2041 0 net=1424
rlabel metal2 184 -2041 184 -2041 0 net=2910
rlabel metal2 695 -2041 695 -2041 0 net=5355
rlabel metal2 751 -2041 751 -2041 0 net=5681
rlabel metal2 891 -2041 891 -2041 0 net=7189
rlabel metal2 75 -2043 75 -2043 0 net=1123
rlabel metal2 695 -2043 695 -2043 0 net=5977
rlabel metal2 758 -2043 758 -2043 0 net=5791
rlabel metal2 79 -2045 79 -2045 0 net=2942
rlabel metal2 429 -2045 429 -2045 0 net=3033
rlabel metal2 492 -2045 492 -2045 0 net=3745
rlabel metal2 506 -2045 506 -2045 0 net=5537
rlabel metal2 761 -2045 761 -2045 0 net=7734
rlabel metal2 86 -2047 86 -2047 0 net=5741
rlabel metal2 814 -2047 814 -2047 0 net=7601
rlabel metal2 86 -2049 86 -2049 0 net=5585
rlabel metal2 765 -2049 765 -2049 0 net=7694
rlabel metal2 96 -2051 96 -2051 0 net=5700
rlabel metal2 100 -2053 100 -2053 0 net=2859
rlabel metal2 117 -2053 117 -2053 0 net=1349
rlabel metal2 184 -2053 184 -2053 0 net=1843
rlabel metal2 688 -2053 688 -2053 0 net=4543
rlabel metal2 114 -2055 114 -2055 0 net=3519
rlabel metal2 401 -2055 401 -2055 0 net=2989
rlabel metal2 443 -2055 443 -2055 0 net=4321
rlabel metal2 709 -2055 709 -2055 0 net=5387
rlabel metal2 768 -2055 768 -2055 0 net=6605
rlabel metal2 121 -2057 121 -2057 0 net=1439
rlabel metal2 226 -2057 226 -2057 0 net=3627
rlabel metal2 618 -2057 618 -2057 0 net=5089
rlabel metal2 786 -2057 786 -2057 0 net=5845
rlabel metal2 82 -2059 82 -2059 0 net=1003
rlabel metal2 128 -2059 128 -2059 0 net=2327
rlabel metal2 338 -2059 338 -2059 0 net=4654
rlabel metal2 555 -2059 555 -2059 0 net=5633
rlabel metal2 110 -2061 110 -2061 0 net=32
rlabel metal2 366 -2061 366 -2061 0 net=3959
rlabel metal2 572 -2061 572 -2061 0 net=5895
rlabel metal2 138 -2063 138 -2063 0 net=4549
rlabel metal2 138 -2065 138 -2065 0 net=6623
rlabel metal2 142 -2067 142 -2067 0 net=2097
rlabel metal2 198 -2067 198 -2067 0 net=1659
rlabel metal2 247 -2067 247 -2067 0 net=2913
rlabel metal2 443 -2067 443 -2067 0 net=4539
rlabel metal2 674 -2067 674 -2067 0 net=4751
rlabel metal2 26 -2069 26 -2069 0 net=3701
rlabel metal2 89 -2071 89 -2071 0 net=2971
rlabel metal2 247 -2071 247 -2071 0 net=1597
rlabel metal2 310 -2071 310 -2071 0 net=3663
rlabel metal2 89 -2073 89 -2073 0 net=5228
rlabel metal2 149 -2075 149 -2075 0 net=3725
rlabel metal2 254 -2075 254 -2075 0 net=2240
rlabel metal2 516 -2075 516 -2075 0 net=7095
rlabel metal2 152 -2077 152 -2077 0 net=2042
rlabel metal2 240 -2077 240 -2077 0 net=2951
rlabel metal2 282 -2077 282 -2077 0 net=2935
rlabel metal2 369 -2077 369 -2077 0 net=6123
rlabel metal2 152 -2079 152 -2079 0 net=7161
rlabel metal2 191 -2081 191 -2081 0 net=1949
rlabel metal2 289 -2081 289 -2081 0 net=1807
rlabel metal2 324 -2081 324 -2081 0 net=2833
rlabel metal2 387 -2081 387 -2081 0 net=2445
rlabel metal2 411 -2081 411 -2081 0 net=7143
rlabel metal2 240 -2083 240 -2083 0 net=3103
rlabel metal2 457 -2083 457 -2083 0 net=3269
rlabel metal2 520 -2083 520 -2083 0 net=3835
rlabel metal2 576 -2083 576 -2083 0 net=4379
rlabel metal2 737 -2083 737 -2083 0 net=6565
rlabel metal2 142 -2085 142 -2085 0 net=3633
rlabel metal2 541 -2085 541 -2085 0 net=3431
rlabel metal2 268 -2087 268 -2087 0 net=2707
rlabel metal2 541 -2087 541 -2087 0 net=3403
rlabel metal2 289 -2089 289 -2089 0 net=6976
rlabel metal2 296 -2091 296 -2091 0 net=1931
rlabel metal2 317 -2091 317 -2091 0 net=3315
rlabel metal2 411 -2091 411 -2091 0 net=4296
rlabel metal2 303 -2093 303 -2093 0 net=1913
rlabel metal2 317 -2095 317 -2095 0 net=2697
rlabel metal2 415 -2095 415 -2095 0 net=3643
rlabel metal2 639 -2095 639 -2095 0 net=7345
rlabel metal2 261 -2097 261 -2097 0 net=2415
rlabel metal2 415 -2097 415 -2097 0 net=6329
rlabel metal2 93 -2099 93 -2099 0 net=1617
rlabel metal2 331 -2099 331 -2099 0 net=1345
rlabel metal2 93 -2101 93 -2101 0 net=82
rlabel metal2 341 -2103 341 -2103 0 net=3919
rlabel metal2 548 -2103 548 -2103 0 net=4960
rlabel metal2 716 -2103 716 -2103 0 net=4665
rlabel metal2 485 -2105 485 -2105 0 net=4157
rlabel metal2 485 -2107 485 -2107 0 net=3049
rlabel metal2 653 -2109 653 -2109 0 net=4595
rlabel metal2 653 -2111 653 -2111 0 net=7391
rlabel metal2 9 -2122 9 -2122 0 net=2842
rlabel metal2 401 -2122 401 -2122 0 net=2446
rlabel metal2 432 -2122 432 -2122 0 net=3326
rlabel metal2 611 -2122 611 -2122 0 net=4152
rlabel metal2 9 -2124 9 -2124 0 net=2953
rlabel metal2 275 -2124 275 -2124 0 net=3402
rlabel metal2 436 -2124 436 -2124 0 net=1870
rlabel metal2 590 -2124 590 -2124 0 net=3664
rlabel metal2 642 -2124 642 -2124 0 net=6514
rlabel metal2 1052 -2124 1052 -2124 0 net=7392
rlabel metal2 1101 -2124 1101 -2124 0 net=6134
rlabel metal2 16 -2126 16 -2126 0 net=2969
rlabel metal2 485 -2126 485 -2126 0 net=3050
rlabel metal2 523 -2126 523 -2126 0 net=5792
rlabel metal2 821 -2126 821 -2126 0 net=6005
rlabel metal2 821 -2126 821 -2126 0 net=6005
rlabel metal2 849 -2126 849 -2126 0 net=6331
rlabel metal2 849 -2126 849 -2126 0 net=6331
rlabel metal2 873 -2126 873 -2126 0 net=6944
rlabel metal2 16 -2128 16 -2128 0 net=4939
rlabel metal2 93 -2128 93 -2128 0 net=2645
rlabel metal2 282 -2128 282 -2128 0 net=2936
rlabel metal2 359 -2128 359 -2128 0 net=2416
rlabel metal2 576 -2128 576 -2128 0 net=7050
rlabel metal2 23 -2130 23 -2130 0 net=3600
rlabel metal2 152 -2130 152 -2130 0 net=3960
rlabel metal2 373 -2130 373 -2130 0 net=3521
rlabel metal2 485 -2130 485 -2130 0 net=3405
rlabel metal2 548 -2130 548 -2130 0 net=3836
rlabel metal2 565 -2130 565 -2130 0 net=7158
rlabel metal2 23 -2132 23 -2132 0 net=3645
rlabel metal2 604 -2132 604 -2132 0 net=7316
rlabel metal2 30 -2134 30 -2134 0 net=1786
rlabel metal2 58 -2134 58 -2134 0 net=2050
rlabel metal2 173 -2134 173 -2134 0 net=2918
rlabel metal2 366 -2134 366 -2134 0 net=2571
rlabel metal2 394 -2134 394 -2134 0 net=3757
rlabel metal2 611 -2134 611 -2134 0 net=4753
rlabel metal2 730 -2134 730 -2134 0 net=5389
rlabel metal2 737 -2134 737 -2134 0 net=7120
rlabel metal2 1017 -2134 1017 -2134 0 net=7611
rlabel metal2 51 -2136 51 -2136 0 net=2185
rlabel metal2 401 -2136 401 -2136 0 net=2623
rlabel metal2 684 -2136 684 -2136 0 net=7016
rlabel metal2 982 -2136 982 -2136 0 net=7603
rlabel metal2 51 -2138 51 -2138 0 net=2211
rlabel metal2 376 -2138 376 -2138 0 net=608
rlabel metal2 415 -2138 415 -2138 0 net=2665
rlabel metal2 723 -2138 723 -2138 0 net=5357
rlabel metal2 807 -2138 807 -2138 0 net=6567
rlabel metal2 884 -2138 884 -2138 0 net=6607
rlabel metal2 884 -2138 884 -2138 0 net=6607
rlabel metal2 898 -2138 898 -2138 0 net=6241
rlabel metal2 898 -2138 898 -2138 0 net=6241
rlabel metal2 940 -2138 940 -2138 0 net=7145
rlabel metal2 961 -2138 961 -2138 0 net=7219
rlabel metal2 1038 -2138 1038 -2138 0 net=7427
rlabel metal2 58 -2140 58 -2140 0 net=3317
rlabel metal2 408 -2140 408 -2140 0 net=3747
rlabel metal2 530 -2140 530 -2140 0 net=7096
rlabel metal2 61 -2142 61 -2142 0 net=3407
rlabel metal2 548 -2142 548 -2142 0 net=4105
rlabel metal2 555 -2142 555 -2142 0 net=3432
rlabel metal2 593 -2142 593 -2142 0 net=7695
rlabel metal2 72 -2144 72 -2144 0 net=3270
rlabel metal2 534 -2144 534 -2144 0 net=3564
rlabel metal2 625 -2144 625 -2144 0 net=7142
rlabel metal2 75 -2146 75 -2146 0 net=7707
rlabel metal2 75 -2148 75 -2148 0 net=4158
rlabel metal2 691 -2148 691 -2148 0 net=5846
rlabel metal2 891 -2148 891 -2148 0 net=7191
rlabel metal2 989 -2148 989 -2148 0 net=7763
rlabel metal2 79 -2150 79 -2150 0 net=5742
rlabel metal2 814 -2150 814 -2150 0 net=6125
rlabel metal2 835 -2150 835 -2150 0 net=6695
rlabel metal2 947 -2150 947 -2150 0 net=6973
rlabel metal2 1003 -2150 1003 -2150 0 net=7519
rlabel metal2 79 -2152 79 -2152 0 net=1951
rlabel metal2 219 -2152 219 -2152 0 net=1479
rlabel metal2 443 -2152 443 -2152 0 net=4540
rlabel metal2 534 -2152 534 -2152 0 net=4323
rlabel metal2 695 -2152 695 -2152 0 net=5979
rlabel metal2 947 -2152 947 -2152 0 net=7163
rlabel metal2 86 -2154 86 -2154 0 net=2906
rlabel metal2 527 -2154 527 -2154 0 net=7235
rlabel metal2 72 -2156 72 -2156 0 net=3171
rlabel metal2 93 -2156 93 -2156 0 net=3911
rlabel metal2 226 -2156 226 -2156 0 net=3629
rlabel metal2 625 -2156 625 -2156 0 net=4597
rlabel metal2 730 -2156 730 -2156 0 net=6537
rlabel metal2 96 -2158 96 -2158 0 net=3702
rlabel metal2 653 -2158 653 -2158 0 net=4481
rlabel metal2 702 -2158 702 -2158 0 net=5683
rlabel metal2 786 -2158 786 -2158 0 net=5897
rlabel metal2 828 -2158 828 -2158 0 net=6421
rlabel metal2 100 -2160 100 -2160 0 net=2861
rlabel metal2 100 -2160 100 -2160 0 net=2861
rlabel metal2 107 -2160 107 -2160 0 net=13
rlabel metal2 317 -2160 317 -2160 0 net=2699
rlabel metal2 443 -2160 443 -2160 0 net=3137
rlabel metal2 471 -2160 471 -2160 0 net=3359
rlabel metal2 765 -2160 765 -2160 0 net=5635
rlabel metal2 779 -2160 779 -2160 0 net=5687
rlabel metal2 835 -2160 835 -2160 0 net=6447
rlabel metal2 37 -2162 37 -2162 0 net=5983
rlabel metal2 863 -2162 863 -2162 0 net=6621
rlabel metal2 44 -2164 44 -2164 0 net=2519
rlabel metal2 320 -2164 320 -2164 0 net=7299
rlabel metal2 44 -2166 44 -2166 0 net=3727
rlabel metal2 226 -2166 226 -2166 0 net=1915
rlabel metal2 324 -2166 324 -2166 0 net=2835
rlabel metal2 453 -2166 453 -2166 0 net=7767
rlabel metal2 107 -2168 107 -2168 0 net=3953
rlabel metal2 177 -2168 177 -2168 0 net=1613
rlabel metal2 303 -2168 303 -2168 0 net=2915
rlabel metal2 464 -2168 464 -2168 0 net=3035
rlabel metal2 527 -2168 527 -2168 0 net=5299
rlabel metal2 744 -2168 744 -2168 0 net=5539
rlabel metal2 905 -2168 905 -2168 0 net=7387
rlabel metal2 65 -2170 65 -2170 0 net=2268
rlabel metal2 198 -2170 198 -2170 0 net=2973
rlabel metal2 345 -2170 345 -2170 0 net=2167
rlabel metal2 555 -2170 555 -2170 0 net=4055
rlabel metal2 656 -2170 656 -2170 0 net=7598
rlabel metal2 65 -2172 65 -2172 0 net=2709
rlabel metal2 422 -2172 422 -2172 0 net=2991
rlabel metal2 597 -2172 597 -2172 0 net=6670
rlabel metal2 110 -2174 110 -2174 0 net=560
rlabel metal2 632 -2174 632 -2174 0 net=4257
rlabel metal2 660 -2174 660 -2174 0 net=4551
rlabel metal2 751 -2174 751 -2174 0 net=5587
rlabel metal2 114 -2176 114 -2176 0 net=5337
rlabel metal2 128 -2176 128 -2176 0 net=2329
rlabel metal2 138 -2176 138 -2176 0 net=7346
rlabel metal2 82 -2178 82 -2178 0 net=1395
rlabel metal2 142 -2178 142 -2178 0 net=3634
rlabel metal2 513 -2178 513 -2178 0 net=5397
rlabel metal2 117 -2180 117 -2180 0 net=4544
rlabel metal2 142 -2182 142 -2182 0 net=3105
rlabel metal2 261 -2182 261 -2182 0 net=1618
rlabel metal2 422 -2182 422 -2182 0 net=2557
rlabel metal2 149 -2184 149 -2184 0 net=2099
rlabel metal2 163 -2184 163 -2184 0 net=1351
rlabel metal2 261 -2184 261 -2184 0 net=1933
rlabel metal2 436 -2184 436 -2184 0 net=7077
rlabel metal2 121 -2186 121 -2186 0 net=3143
rlabel metal2 513 -2186 513 -2186 0 net=4673
rlabel metal2 124 -2188 124 -2188 0 net=2333
rlabel metal2 184 -2188 184 -2188 0 net=1845
rlabel metal2 268 -2188 268 -2188 0 net=1347
rlabel metal2 639 -2188 639 -2188 0 net=5889
rlabel metal2 2 -2190 2 -2190 0 net=5033
rlabel metal2 646 -2190 646 -2190 0 net=4381
rlabel metal2 688 -2190 688 -2190 0 net=6089
rlabel metal2 2 -2192 2 -2192 0 net=1307
rlabel metal2 124 -2194 124 -2194 0 net=7735
rlabel metal2 198 -2196 198 -2196 0 net=1475
rlabel metal2 667 -2196 667 -2196 0 net=7396
rlabel metal2 212 -2198 212 -2198 0 net=1511
rlabel metal2 310 -2198 310 -2198 0 net=1809
rlabel metal2 674 -2198 674 -2198 0 net=4667
rlabel metal2 758 -2198 758 -2198 0 net=6625
rlabel metal2 233 -2200 233 -2200 0 net=1660
rlabel metal2 618 -2200 618 -2200 0 net=5091
rlabel metal2 912 -2200 912 -2200 0 net=6731
rlabel metal2 205 -2202 205 -2202 0 net=1441
rlabel metal2 247 -2202 247 -2202 0 net=1599
rlabel metal2 520 -2202 520 -2202 0 net=3921
rlabel metal2 919 -2202 919 -2202 0 net=6805
rlabel metal2 205 -2204 205 -2204 0 net=3891
rlabel metal2 520 -2204 520 -2204 0 net=5035
rlabel metal2 926 -2204 926 -2204 0 net=7475
rlabel metal2 247 -2206 247 -2206 0 net=1381
rlabel metal2 9 -2217 9 -2217 0 net=2954
rlabel metal2 208 -2217 208 -2217 0 net=5034
rlabel metal2 653 -2217 653 -2217 0 net=4482
rlabel metal2 691 -2217 691 -2217 0 net=6622
rlabel metal2 870 -2217 870 -2217 0 net=7237
rlabel metal2 9 -2219 9 -2219 0 net=6559
rlabel metal2 341 -2219 341 -2219 0 net=3406
rlabel metal2 488 -2219 488 -2219 0 net=5984
rlabel metal2 856 -2219 856 -2219 0 net=6090
rlabel metal2 16 -2221 16 -2221 0 net=4940
rlabel metal2 121 -2221 121 -2221 0 net=1352
rlabel metal2 282 -2221 282 -2221 0 net=1614
rlabel metal2 348 -2221 348 -2221 0 net=2572
rlabel metal2 373 -2221 373 -2221 0 net=3361
rlabel metal2 485 -2221 485 -2221 0 net=5449
rlabel metal2 695 -2221 695 -2221 0 net=7604
rlabel metal2 30 -2223 30 -2223 0 net=2168
rlabel metal2 355 -2223 355 -2223 0 net=2700
rlabel metal2 394 -2223 394 -2223 0 net=7736
rlabel metal2 44 -2225 44 -2225 0 net=3728
rlabel metal2 387 -2225 387 -2225 0 net=2559
rlabel metal2 436 -2225 436 -2225 0 net=2863
rlabel metal2 695 -2225 695 -2225 0 net=5359
rlabel metal2 768 -2225 768 -2225 0 net=5898
rlabel metal2 856 -2225 856 -2225 0 net=7613
rlabel metal2 37 -2227 37 -2227 0 net=4121
rlabel metal2 51 -2227 51 -2227 0 net=2213
rlabel metal2 194 -2227 194 -2227 0 net=1512
rlabel metal2 215 -2227 215 -2227 0 net=3144
rlabel metal2 310 -2227 310 -2227 0 net=1601
rlabel metal2 359 -2227 359 -2227 0 net=2837
rlabel metal2 401 -2227 401 -2227 0 net=2625
rlabel metal2 439 -2227 439 -2227 0 net=7708
rlabel metal2 30 -2229 30 -2229 0 net=4177
rlabel metal2 86 -2229 86 -2229 0 net=3173
rlabel metal2 86 -2229 86 -2229 0 net=3173
rlabel metal2 93 -2229 93 -2229 0 net=3912
rlabel metal2 177 -2229 177 -2229 0 net=2916
rlabel metal2 317 -2229 317 -2229 0 net=2975
rlabel metal2 331 -2229 331 -2229 0 net=1810
rlabel metal2 359 -2229 359 -2229 0 net=5483
rlabel metal2 590 -2229 590 -2229 0 net=6448
rlabel metal2 863 -2229 863 -2229 0 net=7697
rlabel metal2 23 -2231 23 -2231 0 net=3647
rlabel metal2 331 -2231 331 -2231 0 net=2585
rlabel metal2 502 -2231 502 -2231 0 net=4273
rlabel metal2 548 -2231 548 -2231 0 net=4107
rlabel metal2 572 -2231 572 -2231 0 net=5684
rlabel metal2 723 -2231 723 -2231 0 net=6126
rlabel metal2 835 -2231 835 -2231 0 net=7221
rlabel metal2 23 -2233 23 -2233 0 net=5823
rlabel metal2 166 -2233 166 -2233 0 net=752
rlabel metal2 576 -2233 576 -2233 0 net=3631
rlabel metal2 653 -2233 653 -2233 0 net=5037
rlabel metal2 723 -2233 723 -2233 0 net=5637
rlabel metal2 779 -2233 779 -2233 0 net=5891
rlabel metal2 800 -2233 800 -2233 0 net=6733
rlabel metal2 922 -2233 922 -2233 0 net=6974
rlabel metal2 37 -2235 37 -2235 0 net=3107
rlabel metal2 156 -2235 156 -2235 0 net=2335
rlabel metal2 201 -2235 201 -2235 0 net=636
rlabel metal2 590 -2235 590 -2235 0 net=4259
rlabel metal2 667 -2235 667 -2235 0 net=6539
rlabel metal2 737 -2235 737 -2235 0 net=5689
rlabel metal2 793 -2235 793 -2235 0 net=7147
rlabel metal2 961 -2235 961 -2235 0 net=7521
rlabel metal2 2 -2237 2 -2237 0 net=1309
rlabel metal2 170 -2237 170 -2237 0 net=2647
rlabel metal2 282 -2237 282 -2237 0 net=1873
rlabel metal2 401 -2237 401 -2237 0 net=3893
rlabel metal2 506 -2237 506 -2237 0 net=4057
rlabel metal2 597 -2237 597 -2237 0 net=5093
rlabel metal2 726 -2237 726 -2237 0 net=7428
rlabel metal2 2 -2239 2 -2239 0 net=5339
rlabel metal2 121 -2239 121 -2239 0 net=3759
rlabel metal2 604 -2239 604 -2239 0 net=3922
rlabel metal2 681 -2239 681 -2239 0 net=5945
rlabel metal2 758 -2239 758 -2239 0 net=6627
rlabel metal2 814 -2239 814 -2239 0 net=6423
rlabel metal2 884 -2239 884 -2239 0 net=6609
rlabel metal2 884 -2239 884 -2239 0 net=6609
rlabel metal2 940 -2239 940 -2239 0 net=7765
rlabel metal2 79 -2241 79 -2241 0 net=1953
rlabel metal2 198 -2241 198 -2241 0 net=1477
rlabel metal2 296 -2241 296 -2241 0 net=2143
rlabel metal2 408 -2241 408 -2241 0 net=3748
rlabel metal2 513 -2241 513 -2241 0 net=4675
rlabel metal2 698 -2241 698 -2241 0 net=7388
rlabel metal2 93 -2243 93 -2243 0 net=3955
rlabel metal2 114 -2243 114 -2243 0 net=1397
rlabel metal2 135 -2243 135 -2243 0 net=2330
rlabel metal2 380 -2243 380 -2243 0 net=2187
rlabel metal2 429 -2243 429 -2243 0 net=4689
rlabel metal2 527 -2243 527 -2243 0 net=5301
rlabel metal2 583 -2243 583 -2243 0 net=5540
rlabel metal2 100 -2245 100 -2245 0 net=2862
rlabel metal2 135 -2245 135 -2245 0 net=2101
rlabel metal2 156 -2245 156 -2245 0 net=1365
rlabel metal2 205 -2245 205 -2245 0 net=1481
rlabel metal2 226 -2245 226 -2245 0 net=1916
rlabel metal2 429 -2245 429 -2245 0 net=3409
rlabel metal2 548 -2245 548 -2245 0 net=3897
rlabel metal2 604 -2245 604 -2245 0 net=4383
rlabel metal2 709 -2245 709 -2245 0 net=5589
rlabel metal2 772 -2245 772 -2245 0 net=6333
rlabel metal2 65 -2247 65 -2247 0 net=2711
rlabel metal2 212 -2247 212 -2247 0 net=1348
rlabel metal2 450 -2247 450 -2247 0 net=3523
rlabel metal2 618 -2247 618 -2247 0 net=4599
rlabel metal2 646 -2247 646 -2247 0 net=4827
rlabel metal2 716 -2247 716 -2247 0 net=6696
rlabel metal2 33 -2249 33 -2249 0 net=1849
rlabel metal2 450 -2249 450 -2249 0 net=5391
rlabel metal2 758 -2249 758 -2249 0 net=6007
rlabel metal2 828 -2249 828 -2249 0 net=7079
rlabel metal2 65 -2251 65 -2251 0 net=1879
rlabel metal2 226 -2251 226 -2251 0 net=2521
rlabel metal2 352 -2251 352 -2251 0 net=7051
rlabel metal2 821 -2251 821 -2251 0 net=7301
rlabel metal2 72 -2253 72 -2253 0 net=2023
rlabel metal2 240 -2253 240 -2253 0 net=1846
rlabel metal2 352 -2253 352 -2253 0 net=3036
rlabel metal2 467 -2253 467 -2253 0 net=2463
rlabel metal2 541 -2253 541 -2253 0 net=5980
rlabel metal2 891 -2253 891 -2253 0 net=7769
rlabel metal2 240 -2255 240 -2255 0 net=2667
rlabel metal2 457 -2255 457 -2255 0 net=2970
rlabel metal2 593 -2255 593 -2255 0 net=3391
rlabel metal2 684 -2255 684 -2255 0 net=6879
rlabel metal2 842 -2255 842 -2255 0 net=6807
rlabel metal2 968 -2255 968 -2255 0 net=5943
rlabel metal2 58 -2257 58 -2257 0 net=3319
rlabel metal2 443 -2257 443 -2257 0 net=3139
rlabel metal2 471 -2257 471 -2257 0 net=4755
rlabel metal2 849 -2257 849 -2257 0 net=6243
rlabel metal2 912 -2257 912 -2257 0 net=2209
rlabel metal2 16 -2259 16 -2259 0 net=6155
rlabel metal2 247 -2259 247 -2259 0 net=1383
rlabel metal2 247 -2259 247 -2259 0 net=1383
rlabel metal2 254 -2259 254 -2259 0 net=3735
rlabel metal2 443 -2259 443 -2259 0 net=4669
rlabel metal2 877 -2259 877 -2259 0 net=7477
rlabel metal2 261 -2261 261 -2261 0 net=1935
rlabel metal2 478 -2261 478 -2261 0 net=2993
rlabel metal2 233 -2263 233 -2263 0 net=1443
rlabel metal2 478 -2263 478 -2263 0 net=4721
rlabel metal2 534 -2263 534 -2263 0 net=4324
rlabel metal2 233 -2265 233 -2265 0 net=5329
rlabel metal2 611 -2265 611 -2265 0 net=4553
rlabel metal2 502 -2267 502 -2267 0 net=1321
rlabel metal2 660 -2267 660 -2267 0 net=5399
rlabel metal2 751 -2269 751 -2269 0 net=6569
rlabel metal2 807 -2271 807 -2271 0 net=7165
rlabel metal2 947 -2273 947 -2273 0 net=7193
rlabel metal2 464 -2275 464 -2275 0 net=5129
rlabel metal2 2 -2286 2 -2286 0 net=5340
rlabel metal2 58 -2286 58 -2286 0 net=1478
rlabel metal2 303 -2286 303 -2286 0 net=3648
rlabel metal2 481 -2286 481 -2286 0 net=7770
rlabel metal2 905 -2286 905 -2286 0 net=2210
rlabel metal2 2 -2288 2 -2288 0 net=4179
rlabel metal2 44 -2288 44 -2288 0 net=4122
rlabel metal2 58 -2288 58 -2288 0 net=2865
rlabel metal2 450 -2288 450 -2288 0 net=5392
rlabel metal2 499 -2288 499 -2288 0 net=4555
rlabel metal2 618 -2288 618 -2288 0 net=4601
rlabel metal2 618 -2288 618 -2288 0 net=4601
rlabel metal2 639 -2288 639 -2288 0 net=3632
rlabel metal2 639 -2288 639 -2288 0 net=3632
rlabel metal2 642 -2288 642 -2288 0 net=6734
rlabel metal2 877 -2288 877 -2288 0 net=7479
rlabel metal2 908 -2288 908 -2288 0 net=7194
rlabel metal2 9 -2290 9 -2290 0 net=6560
rlabel metal2 191 -2290 191 -2290 0 net=2215
rlabel metal2 226 -2290 226 -2290 0 net=2523
rlabel metal2 376 -2290 376 -2290 0 net=4828
rlabel metal2 684 -2290 684 -2290 0 net=7222
rlabel metal2 877 -2290 877 -2290 0 net=5131
rlabel metal2 12 -2292 12 -2292 0 net=1137
rlabel metal2 268 -2292 268 -2292 0 net=1850
rlabel metal2 502 -2292 502 -2292 0 net=5638
rlabel metal2 765 -2292 765 -2292 0 net=7081
rlabel metal2 884 -2292 884 -2292 0 net=6610
rlabel metal2 922 -2292 922 -2292 0 net=227
rlabel metal2 947 -2292 947 -2292 0 net=7523
rlabel metal2 16 -2294 16 -2294 0 net=6156
rlabel metal2 506 -2294 506 -2294 0 net=4059
rlabel metal2 506 -2294 506 -2294 0 net=4059
rlabel metal2 534 -2294 534 -2294 0 net=1322
rlabel metal2 569 -2294 569 -2294 0 net=4109
rlabel metal2 569 -2294 569 -2294 0 net=4109
rlabel metal2 576 -2294 576 -2294 0 net=7614
rlabel metal2 926 -2294 926 -2294 0 net=5944
rlabel metal2 16 -2296 16 -2296 0 net=5331
rlabel metal2 268 -2296 268 -2296 0 net=2144
rlabel metal2 303 -2296 303 -2296 0 net=3321
rlabel metal2 436 -2296 436 -2296 0 net=3141
rlabel metal2 464 -2296 464 -2296 0 net=3524
rlabel metal2 583 -2296 583 -2296 0 net=5400
rlabel metal2 723 -2296 723 -2296 0 net=7303
rlabel metal2 842 -2296 842 -2296 0 net=6809
rlabel metal2 23 -2298 23 -2298 0 net=5824
rlabel metal2 61 -2298 61 -2298 0 net=823
rlabel metal2 768 -2298 768 -2298 0 net=6244
rlabel metal2 856 -2298 856 -2298 0 net=1353
rlabel metal2 23 -2300 23 -2300 0 net=1875
rlabel metal2 296 -2300 296 -2300 0 net=1777
rlabel metal2 467 -2300 467 -2300 0 net=4756
rlabel metal2 520 -2300 520 -2300 0 net=4275
rlabel metal2 597 -2300 597 -2300 0 net=5095
rlabel metal2 779 -2300 779 -2300 0 net=5893
rlabel metal2 849 -2300 849 -2300 0 net=3503
rlabel metal2 30 -2302 30 -2302 0 net=3969
rlabel metal2 233 -2302 233 -2302 0 net=1445
rlabel metal2 275 -2302 275 -2302 0 net=3567
rlabel metal2 373 -2302 373 -2302 0 net=3363
rlabel metal2 562 -2302 562 -2302 0 net=6008
rlabel metal2 786 -2302 786 -2302 0 net=6629
rlabel metal2 44 -2304 44 -2304 0 net=6053
rlabel metal2 793 -2304 793 -2304 0 net=7149
rlabel metal2 47 -2306 47 -2306 0 net=319
rlabel metal2 163 -2306 163 -2306 0 net=1955
rlabel metal2 261 -2306 261 -2306 0 net=1407
rlabel metal2 310 -2306 310 -2306 0 net=1936
rlabel metal2 341 -2306 341 -2306 0 net=657
rlabel metal2 793 -2306 793 -2306 0 net=7699
rlabel metal2 65 -2308 65 -2308 0 net=1880
rlabel metal2 313 -2308 313 -2308 0 net=7099
rlabel metal2 800 -2308 800 -2308 0 net=6424
rlabel metal2 65 -2310 65 -2310 0 net=5295
rlabel metal2 107 -2310 107 -2310 0 net=3392
rlabel metal2 667 -2310 667 -2310 0 net=6541
rlabel metal2 72 -2312 72 -2312 0 net=2024
rlabel metal2 282 -2312 282 -2312 0 net=2189
rlabel metal2 415 -2312 415 -2312 0 net=5377
rlabel metal2 72 -2314 72 -2314 0 net=2131
rlabel metal2 82 -2314 82 -2314 0 net=3174
rlabel metal2 93 -2314 93 -2314 0 net=3956
rlabel metal2 107 -2314 107 -2314 0 net=51
rlabel metal2 114 -2314 114 -2314 0 net=1398
rlabel metal2 289 -2314 289 -2314 0 net=1603
rlabel metal2 355 -2314 355 -2314 0 net=3185
rlabel metal2 537 -2314 537 -2314 0 net=5693
rlabel metal2 79 -2316 79 -2316 0 net=2713
rlabel metal2 163 -2316 163 -2316 0 net=1429
rlabel metal2 355 -2316 355 -2316 0 net=5113
rlabel metal2 681 -2316 681 -2316 0 net=1811
rlabel metal2 86 -2318 86 -2318 0 net=2743
rlabel metal2 586 -2318 586 -2318 0 net=5249
rlabel metal2 93 -2320 93 -2320 0 net=707
rlabel metal2 597 -2320 597 -2320 0 net=4385
rlabel metal2 611 -2320 611 -2320 0 net=4677
rlabel metal2 100 -2322 100 -2322 0 net=2627
rlabel metal2 450 -2322 450 -2322 0 net=5947
rlabel metal2 114 -2324 114 -2324 0 net=2103
rlabel metal2 149 -2324 149 -2324 0 net=2337
rlabel metal2 198 -2324 198 -2324 0 net=1483
rlabel metal2 317 -2324 317 -2324 0 net=2976
rlabel metal2 401 -2324 401 -2324 0 net=3895
rlabel metal2 625 -2324 625 -2324 0 net=5451
rlabel metal2 54 -2326 54 -2326 0 net=6323
rlabel metal2 142 -2326 142 -2326 0 net=1311
rlabel metal2 205 -2326 205 -2326 0 net=2377
rlabel metal2 359 -2326 359 -2326 0 net=5485
rlabel metal2 128 -2328 128 -2328 0 net=2669
rlabel metal2 317 -2328 317 -2328 0 net=2995
rlabel metal2 688 -2328 688 -2328 0 net=5361
rlabel metal2 142 -2330 142 -2330 0 net=1367
rlabel metal2 177 -2330 177 -2330 0 net=1385
rlabel metal2 324 -2330 324 -2330 0 net=4671
rlabel metal2 513 -2330 513 -2330 0 net=4691
rlabel metal2 674 -2330 674 -2330 0 net=5591
rlabel metal2 37 -2332 37 -2332 0 net=3108
rlabel metal2 180 -2332 180 -2332 0 net=6453
rlabel metal2 702 -2332 702 -2332 0 net=6881
rlabel metal2 37 -2334 37 -2334 0 net=3789
rlabel metal2 121 -2334 121 -2334 0 net=3761
rlabel metal2 254 -2334 254 -2334 0 net=3737
rlabel metal2 702 -2334 702 -2334 0 net=6570
rlabel metal2 121 -2336 121 -2336 0 net=3097
rlabel metal2 359 -2336 359 -2336 0 net=2838
rlabel metal2 401 -2336 401 -2336 0 net=5038
rlabel metal2 737 -2336 737 -2336 0 net=5691
rlabel metal2 240 -2338 240 -2338 0 net=2465
rlabel metal2 737 -2338 737 -2338 0 net=7053
rlabel metal2 254 -2340 254 -2340 0 net=1399
rlabel metal2 744 -2340 744 -2340 0 net=6335
rlabel metal2 352 -2342 352 -2342 0 net=3827
rlabel metal2 772 -2342 772 -2342 0 net=7238
rlabel metal2 366 -2344 366 -2344 0 net=4499
rlabel metal2 870 -2344 870 -2344 0 net=7766
rlabel metal2 170 -2346 170 -2346 0 net=2649
rlabel metal2 380 -2346 380 -2346 0 net=6263
rlabel metal2 159 -2348 159 -2348 0 net=2019
rlabel metal2 331 -2348 331 -2348 0 net=2587
rlabel metal2 383 -2348 383 -2348 0 net=2641
rlabel metal2 422 -2348 422 -2348 0 net=3411
rlabel metal2 443 -2348 443 -2348 0 net=3899
rlabel metal2 373 -2350 373 -2350 0 net=4235
rlabel metal2 492 -2350 492 -2350 0 net=4723
rlabel metal2 387 -2352 387 -2352 0 net=2561
rlabel metal2 387 -2352 387 -2352 0 net=2561
rlabel metal2 394 -2352 394 -2352 0 net=7375
rlabel metal2 492 -2354 492 -2354 0 net=5303
rlabel metal2 548 -2356 548 -2356 0 net=4261
rlabel metal2 544 -2358 544 -2358 0 net=4643
rlabel metal2 555 -2360 555 -2360 0 net=7166
rlabel metal2 583 -2362 583 -2362 0 net=7127
rlabel metal2 16 -2373 16 -2373 0 net=5332
rlabel metal2 142 -2373 142 -2373 0 net=1369
rlabel metal2 142 -2373 142 -2373 0 net=1369
rlabel metal2 156 -2373 156 -2373 0 net=305
rlabel metal2 226 -2373 226 -2373 0 net=5250
rlabel metal2 702 -2373 702 -2373 0 net=6883
rlabel metal2 726 -2373 726 -2373 0 net=6630
rlabel metal2 884 -2373 884 -2373 0 net=6811
rlabel metal2 884 -2373 884 -2373 0 net=6811
rlabel metal2 891 -2373 891 -2373 0 net=7481
rlabel metal2 891 -2373 891 -2373 0 net=7481
rlabel metal2 926 -2373 926 -2373 0 net=3229
rlabel metal2 926 -2373 926 -2373 0 net=3229
rlabel metal2 940 -2373 940 -2373 0 net=7525
rlabel metal2 23 -2375 23 -2375 0 net=1876
rlabel metal2 240 -2375 240 -2375 0 net=2466
rlabel metal2 569 -2375 569 -2375 0 net=4111
rlabel metal2 709 -2375 709 -2375 0 net=7083
rlabel metal2 772 -2375 772 -2375 0 net=5894
rlabel metal2 30 -2377 30 -2377 0 net=3970
rlabel metal2 177 -2377 177 -2377 0 net=1387
rlabel metal2 233 -2377 233 -2377 0 net=1447
rlabel metal2 247 -2377 247 -2377 0 net=3763
rlabel metal2 376 -2377 376 -2377 0 net=5694
rlabel metal2 761 -2377 761 -2377 0 net=7150
rlabel metal2 2 -2379 2 -2379 0 net=4180
rlabel metal2 44 -2379 44 -2379 0 net=1035
rlabel metal2 72 -2379 72 -2379 0 net=2132
rlabel metal2 72 -2379 72 -2379 0 net=2132
rlabel metal2 86 -2379 86 -2379 0 net=2745
rlabel metal2 86 -2379 86 -2379 0 net=2745
rlabel metal2 93 -2379 93 -2379 0 net=625
rlabel metal2 212 -2379 212 -2379 0 net=2216
rlabel metal2 404 -2379 404 -2379 0 net=6054
rlabel metal2 828 -2379 828 -2379 0 net=5133
rlabel metal2 37 -2381 37 -2381 0 net=3791
rlabel metal2 100 -2381 100 -2381 0 net=2629
rlabel metal2 411 -2381 411 -2381 0 net=3142
rlabel metal2 457 -2381 457 -2381 0 net=4276
rlabel metal2 583 -2381 583 -2381 0 net=5115
rlabel metal2 723 -2381 723 -2381 0 net=7305
rlabel metal2 772 -2381 772 -2381 0 net=7701
rlabel metal2 51 -2383 51 -2383 0 net=5486
rlabel metal2 751 -2383 751 -2383 0 net=5692
rlabel metal2 100 -2385 100 -2385 0 net=2339
rlabel metal2 177 -2385 177 -2385 0 net=1401
rlabel metal2 261 -2385 261 -2385 0 net=1409
rlabel metal2 261 -2385 261 -2385 0 net=1409
rlabel metal2 268 -2385 268 -2385 0 net=1605
rlabel metal2 303 -2385 303 -2385 0 net=3322
rlabel metal2 460 -2385 460 -2385 0 net=4060
rlabel metal2 520 -2385 520 -2385 0 net=4263
rlabel metal2 555 -2385 555 -2385 0 net=5453
rlabel metal2 639 -2385 639 -2385 0 net=5362
rlabel metal2 723 -2385 723 -2385 0 net=3504
rlabel metal2 107 -2387 107 -2387 0 net=5948
rlabel metal2 464 -2387 464 -2387 0 net=3999
rlabel metal2 523 -2387 523 -2387 0 net=4678
rlabel metal2 618 -2387 618 -2387 0 net=4602
rlabel metal2 639 -2387 639 -2387 0 net=7377
rlabel metal2 107 -2389 107 -2389 0 net=2459
rlabel metal2 163 -2389 163 -2389 0 net=1431
rlabel metal2 310 -2389 310 -2389 0 net=4500
rlabel metal2 611 -2389 611 -2389 0 net=5593
rlabel metal2 114 -2391 114 -2391 0 net=2104
rlabel metal2 163 -2391 163 -2391 0 net=1313
rlabel metal2 205 -2391 205 -2391 0 net=2379
rlabel metal2 275 -2391 275 -2391 0 net=3568
rlabel metal2 408 -2391 408 -2391 0 net=2643
rlabel metal2 450 -2391 450 -2391 0 net=3187
rlabel metal2 481 -2391 481 -2391 0 net=5378
rlabel metal2 114 -2393 114 -2393 0 net=2021
rlabel metal2 184 -2393 184 -2393 0 net=185
rlabel metal2 233 -2393 233 -2393 0 net=2563
rlabel metal2 408 -2393 408 -2393 0 net=5096
rlabel metal2 660 -2393 660 -2393 0 net=7055
rlabel metal2 121 -2395 121 -2395 0 net=3098
rlabel metal2 275 -2395 275 -2395 0 net=3413
rlabel metal2 464 -2395 464 -2395 0 net=6542
rlabel metal2 65 -2397 65 -2397 0 net=5297
rlabel metal2 135 -2397 135 -2397 0 net=6325
rlabel metal2 310 -2397 310 -2397 0 net=3837
rlabel metal2 380 -2397 380 -2397 0 net=2589
rlabel metal2 618 -2397 618 -2397 0 net=6455
rlabel metal2 716 -2397 716 -2397 0 net=7129
rlabel metal2 170 -2399 170 -2399 0 net=1957
rlabel metal2 219 -2399 219 -2399 0 net=150
rlabel metal2 551 -2399 551 -2399 0 net=4471
rlabel metal2 674 -2399 674 -2399 0 net=7101
rlabel metal2 807 -2399 807 -2399 0 net=1813
rlabel metal2 191 -2401 191 -2401 0 net=1485
rlabel metal2 282 -2401 282 -2401 0 net=2190
rlabel metal2 471 -2401 471 -2401 0 net=5939
rlabel metal2 737 -2401 737 -2401 0 net=6337
rlabel metal2 128 -2403 128 -2403 0 net=2671
rlabel metal2 313 -2403 313 -2403 0 net=3896
rlabel metal2 744 -2403 744 -2403 0 net=1355
rlabel metal2 128 -2405 128 -2405 0 net=1779
rlabel metal2 324 -2405 324 -2405 0 net=4672
rlabel metal2 345 -2405 345 -2405 0 net=2525
rlabel metal2 527 -2405 527 -2405 0 net=3829
rlabel metal2 79 -2407 79 -2407 0 net=2714
rlabel metal2 317 -2407 317 -2407 0 net=2997
rlabel metal2 527 -2407 527 -2407 0 net=4645
rlabel metal2 58 -2409 58 -2409 0 net=2867
rlabel metal2 198 -2409 198 -2409 0 net=4853
rlabel metal2 317 -2409 317 -2409 0 net=2527
rlabel metal2 58 -2411 58 -2411 0 net=4243
rlabel metal2 324 -2411 324 -2411 0 net=3455
rlabel metal2 534 -2411 534 -2411 0 net=4386
rlabel metal2 331 -2413 331 -2413 0 net=6311
rlabel metal2 415 -2413 415 -2413 0 net=4237
rlabel metal2 499 -2413 499 -2413 0 net=4557
rlabel metal2 597 -2413 597 -2413 0 net=6265
rlabel metal2 331 -2415 331 -2415 0 net=2650
rlabel metal2 429 -2415 429 -2415 0 net=5623
rlabel metal2 653 -2415 653 -2415 0 net=4725
rlabel metal2 334 -2417 334 -2417 0 net=6937
rlabel metal2 401 -2417 401 -2417 0 net=6317
rlabel metal2 254 -2419 254 -2419 0 net=2367
rlabel metal2 338 -2419 338 -2419 0 net=3739
rlabel metal2 366 -2421 366 -2421 0 net=3365
rlabel metal2 499 -2421 499 -2421 0 net=4693
rlabel metal2 401 -2423 401 -2423 0 net=5305
rlabel metal2 513 -2423 513 -2423 0 net=3913
rlabel metal2 443 -2425 443 -2425 0 net=3901
rlabel metal2 394 -2427 394 -2427 0 net=6705
rlabel metal2 488 -2427 488 -2427 0 net=7277
rlabel metal2 65 -2438 65 -2438 0 net=4245
rlabel metal2 79 -2438 79 -2438 0 net=2868
rlabel metal2 268 -2438 268 -2438 0 net=1606
rlabel metal2 422 -2438 422 -2438 0 net=2526
rlabel metal2 471 -2438 471 -2438 0 net=5116
rlabel metal2 590 -2438 590 -2438 0 net=5624
rlabel metal2 625 -2438 625 -2438 0 net=7130
rlabel metal2 730 -2438 730 -2438 0 net=6338
rlabel metal2 754 -2438 754 -2438 0 net=1814
rlabel metal2 884 -2438 884 -2438 0 net=6813
rlabel metal2 884 -2438 884 -2438 0 net=6813
rlabel metal2 891 -2438 891 -2438 0 net=7483
rlabel metal2 891 -2438 891 -2438 0 net=7483
rlabel metal2 926 -2438 926 -2438 0 net=3230
rlabel metal2 940 -2438 940 -2438 0 net=7527
rlabel metal2 940 -2438 940 -2438 0 net=7527
rlabel metal2 93 -2440 93 -2440 0 net=3792
rlabel metal2 135 -2440 135 -2440 0 net=1371
rlabel metal2 170 -2440 170 -2440 0 net=1958
rlabel metal2 233 -2440 233 -2440 0 net=2564
rlabel metal2 401 -2440 401 -2440 0 net=5307
rlabel metal2 474 -2440 474 -2440 0 net=462
rlabel metal2 485 -2440 485 -2440 0 net=2590
rlabel metal2 625 -2440 625 -2440 0 net=7057
rlabel metal2 681 -2440 681 -2440 0 net=4727
rlabel metal2 695 -2440 695 -2440 0 net=6884
rlabel metal2 716 -2440 716 -2440 0 net=6471
rlabel metal2 730 -2440 730 -2440 0 net=7621
rlabel metal2 765 -2440 765 -2440 0 net=7307
rlabel metal2 765 -2440 765 -2440 0 net=7307
rlabel metal2 779 -2440 779 -2440 0 net=5134
rlabel metal2 100 -2442 100 -2442 0 net=2340
rlabel metal2 191 -2442 191 -2442 0 net=1486
rlabel metal2 240 -2442 240 -2442 0 net=1448
rlabel metal2 275 -2442 275 -2442 0 net=3414
rlabel metal2 334 -2442 334 -2442 0 net=290
rlabel metal2 408 -2442 408 -2442 0 net=4239
rlabel metal2 422 -2442 422 -2442 0 net=5375
rlabel metal2 502 -2442 502 -2442 0 net=3830
rlabel metal2 576 -2442 576 -2442 0 net=6318
rlabel metal2 660 -2442 660 -2442 0 net=4113
rlabel metal2 681 -2442 681 -2442 0 net=7085
rlabel metal2 100 -2444 100 -2444 0 net=5099
rlabel metal2 121 -2444 121 -2444 0 net=5298
rlabel metal2 226 -2444 226 -2444 0 net=1389
rlabel metal2 296 -2444 296 -2444 0 net=6266
rlabel metal2 604 -2444 604 -2444 0 net=5595
rlabel metal2 642 -2444 642 -2444 0 net=4472
rlabel metal2 709 -2444 709 -2444 0 net=1357
rlabel metal2 107 -2446 107 -2446 0 net=2461
rlabel metal2 128 -2446 128 -2446 0 net=1781
rlabel metal2 226 -2446 226 -2446 0 net=1411
rlabel metal2 303 -2446 303 -2446 0 net=6327
rlabel metal2 303 -2446 303 -2446 0 net=6327
rlabel metal2 310 -2446 310 -2446 0 net=3838
rlabel metal2 506 -2446 506 -2446 0 net=4000
rlabel metal2 611 -2446 611 -2446 0 net=7279
rlabel metal2 114 -2448 114 -2448 0 net=2022
rlabel metal2 254 -2448 254 -2448 0 net=2369
rlabel metal2 317 -2448 317 -2448 0 net=2528
rlabel metal2 443 -2448 443 -2448 0 net=6707
rlabel metal2 499 -2448 499 -2448 0 net=4695
rlabel metal2 513 -2448 513 -2448 0 net=3914
rlabel metal2 107 -2450 107 -2450 0 net=3357
rlabel metal2 149 -2450 149 -2450 0 net=3925
rlabel metal2 191 -2450 191 -2450 0 net=4855
rlabel metal2 222 -2450 222 -2450 0 net=4799
rlabel metal2 345 -2450 345 -2450 0 net=2999
rlabel metal2 443 -2450 443 -2450 0 net=3189
rlabel metal2 457 -2450 457 -2450 0 net=3903
rlabel metal2 513 -2450 513 -2450 0 net=4559
rlabel metal2 541 -2450 541 -2450 0 net=5941
rlabel metal2 569 -2450 569 -2450 0 net=6457
rlabel metal2 86 -2452 86 -2452 0 net=2746
rlabel metal2 460 -2452 460 -2452 0 net=4264
rlabel metal2 527 -2452 527 -2452 0 net=4646
rlabel metal2 555 -2452 555 -2452 0 net=5455
rlabel metal2 152 -2454 152 -2454 0 net=2977
rlabel metal2 282 -2454 282 -2454 0 net=2673
rlabel metal2 331 -2454 331 -2454 0 net=7649
rlabel metal2 348 -2454 348 -2454 0 net=6938
rlabel metal2 534 -2454 534 -2454 0 net=7102
rlabel metal2 163 -2456 163 -2456 0 net=1314
rlabel metal2 289 -2456 289 -2456 0 net=1432
rlabel metal2 548 -2456 548 -2456 0 net=7379
rlabel metal2 674 -2456 674 -2456 0 net=5085
rlabel metal2 163 -2458 163 -2458 0 net=3623
rlabel metal2 212 -2458 212 -2458 0 net=5559
rlabel metal2 352 -2458 352 -2458 0 net=3764
rlabel metal2 639 -2458 639 -2458 0 net=392
rlabel metal2 737 -2458 737 -2458 0 net=2303
rlabel metal2 184 -2460 184 -2460 0 net=6489
rlabel metal2 247 -2460 247 -2460 0 net=2381
rlabel metal2 324 -2460 324 -2460 0 net=3457
rlabel metal2 359 -2460 359 -2460 0 net=2630
rlabel metal2 723 -2460 723 -2460 0 net=3873
rlabel metal2 177 -2462 177 -2462 0 net=1403
rlabel metal2 338 -2462 338 -2462 0 net=3741
rlabel metal2 366 -2462 366 -2462 0 net=3367
rlabel metal2 761 -2462 761 -2462 0 net=7702
rlabel metal2 159 -2464 159 -2464 0 net=5965
rlabel metal2 299 -2464 299 -2464 0 net=1851
rlabel metal2 387 -2464 387 -2464 0 net=2644
rlabel metal2 380 -2466 380 -2466 0 net=6313
rlabel metal2 373 -2468 373 -2468 0 net=3223
rlabel metal2 394 -2468 394 -2468 0 net=1341
rlabel metal2 5 -2479 5 -2479 0 net=444
rlabel metal2 5 -2479 5 -2479 0 net=444
rlabel metal2 65 -2479 65 -2479 0 net=4246
rlabel metal2 86 -2479 86 -2479 0 net=2223
rlabel metal2 100 -2479 100 -2479 0 net=5100
rlabel metal2 114 -2479 114 -2479 0 net=2462
rlabel metal2 131 -2479 131 -2479 0 net=1372
rlabel metal2 142 -2479 142 -2479 0 net=3927
rlabel metal2 177 -2479 177 -2479 0 net=5966
rlabel metal2 198 -2479 198 -2479 0 net=2979
rlabel metal2 219 -2479 219 -2479 0 net=1783
rlabel metal2 282 -2479 282 -2479 0 net=5560
rlabel metal2 376 -2479 376 -2479 0 net=5376
rlabel metal2 432 -2479 432 -2479 0 net=3904
rlabel metal2 467 -2479 467 -2479 0 net=6708
rlabel metal2 502 -2479 502 -2479 0 net=4560
rlabel metal2 523 -2479 523 -2479 0 net=5942
rlabel metal2 576 -2479 576 -2479 0 net=5456
rlabel metal2 590 -2479 590 -2479 0 net=7058
rlabel metal2 660 -2479 660 -2479 0 net=4115
rlabel metal2 660 -2479 660 -2479 0 net=4115
rlabel metal2 667 -2479 667 -2479 0 net=7087
rlabel metal2 730 -2479 730 -2479 0 net=7622
rlabel metal2 730 -2479 730 -2479 0 net=7622
rlabel metal2 744 -2479 744 -2479 0 net=4647
rlabel metal2 758 -2479 758 -2479 0 net=7308
rlabel metal2 884 -2479 884 -2479 0 net=6814
rlabel metal2 884 -2479 884 -2479 0 net=6814
rlabel metal2 891 -2479 891 -2479 0 net=7485
rlabel metal2 891 -2479 891 -2479 0 net=7485
rlabel metal2 933 -2479 933 -2479 0 net=3975
rlabel metal2 940 -2479 940 -2479 0 net=7529
rlabel metal2 100 -2481 100 -2481 0 net=5811
rlabel metal2 138 -2481 138 -2481 0 net=173
rlabel metal2 226 -2481 226 -2481 0 net=1413
rlabel metal2 247 -2481 247 -2481 0 net=1404
rlabel metal2 338 -2481 338 -2481 0 net=1852
rlabel metal2 450 -2481 450 -2481 0 net=7380
rlabel metal2 597 -2481 597 -2481 0 net=5086
rlabel metal2 681 -2481 681 -2481 0 net=4729
rlabel metal2 758 -2481 758 -2481 0 net=6671
rlabel metal2 107 -2483 107 -2483 0 net=3358
rlabel metal2 149 -2483 149 -2483 0 net=3625
rlabel metal2 177 -2483 177 -2483 0 net=4857
rlabel metal2 205 -2483 205 -2483 0 net=6491
rlabel metal2 205 -2483 205 -2483 0 net=6491
rlabel metal2 226 -2483 226 -2483 0 net=6885
rlabel metal2 275 -2483 275 -2483 0 net=1391
rlabel metal2 352 -2483 352 -2483 0 net=3459
rlabel metal2 352 -2483 352 -2483 0 net=3459
rlabel metal2 359 -2483 359 -2483 0 net=3742
rlabel metal2 380 -2483 380 -2483 0 net=3225
rlabel metal2 380 -2483 380 -2483 0 net=3225
rlabel metal2 394 -2483 394 -2483 0 net=1343
rlabel metal2 394 -2483 394 -2483 0 net=1343
rlabel metal2 401 -2483 401 -2483 0 net=3000
rlabel metal2 443 -2483 443 -2483 0 net=3191
rlabel metal2 471 -2483 471 -2483 0 net=5308
rlabel metal2 604 -2483 604 -2483 0 net=5597
rlabel metal2 604 -2483 604 -2483 0 net=5597
rlabel metal2 611 -2483 611 -2483 0 net=7281
rlabel metal2 611 -2483 611 -2483 0 net=7281
rlabel metal2 688 -2483 688 -2483 0 net=2263
rlabel metal2 159 -2485 159 -2485 0 net=4123
rlabel metal2 233 -2485 233 -2485 0 net=5493
rlabel metal2 271 -2485 271 -2485 0 net=2551
rlabel metal2 296 -2485 296 -2485 0 net=6328
rlabel metal2 310 -2485 310 -2485 0 net=4800
rlabel metal2 401 -2485 401 -2485 0 net=30
rlabel metal2 695 -2485 695 -2485 0 net=1359
rlabel metal2 236 -2487 236 -2487 0 net=6897
rlabel metal2 359 -2487 359 -2487 0 net=4240
rlabel metal2 415 -2487 415 -2487 0 net=3369
rlabel metal2 506 -2487 506 -2487 0 net=4696
rlabel metal2 523 -2487 523 -2487 0 net=2219
rlabel metal2 709 -2487 709 -2487 0 net=6473
rlabel metal2 240 -2489 240 -2489 0 net=3753
rlabel metal2 303 -2489 303 -2489 0 net=7650
rlabel metal2 408 -2489 408 -2489 0 net=6315
rlabel metal2 520 -2489 520 -2489 0 net=6458
rlabel metal2 716 -2489 716 -2489 0 net=3875
rlabel metal2 247 -2491 247 -2491 0 net=2371
rlabel metal2 317 -2491 317 -2491 0 net=2675
rlabel metal2 723 -2491 723 -2491 0 net=2305
rlabel metal2 289 -2493 289 -2493 0 net=2383
rlabel metal2 201 -2495 201 -2495 0 net=6673
rlabel metal2 5 -2506 5 -2506 0 net=5373
rlabel metal2 86 -2506 86 -2506 0 net=2224
rlabel metal2 107 -2506 107 -2506 0 net=5812
rlabel metal2 142 -2506 142 -2506 0 net=3928
rlabel metal2 201 -2506 201 -2506 0 net=6492
rlabel metal2 219 -2506 219 -2506 0 net=3754
rlabel metal2 247 -2506 247 -2506 0 net=2372
rlabel metal2 275 -2506 275 -2506 0 net=2552
rlabel metal2 285 -2506 285 -2506 0 net=2384
rlabel metal2 331 -2506 331 -2506 0 net=2677
rlabel metal2 352 -2506 352 -2506 0 net=3460
rlabel metal2 380 -2506 380 -2506 0 net=3226
rlabel metal2 387 -2506 387 -2506 0 net=6316
rlabel metal2 450 -2506 450 -2506 0 net=3192
rlabel metal2 523 -2506 523 -2506 0 net=2220
rlabel metal2 597 -2506 597 -2506 0 net=5598
rlabel metal2 660 -2506 660 -2506 0 net=4116
rlabel metal2 667 -2506 667 -2506 0 net=7089
rlabel metal2 667 -2506 667 -2506 0 net=7089
rlabel metal2 681 -2506 681 -2506 0 net=4730
rlabel metal2 709 -2506 709 -2506 0 net=6474
rlabel metal2 716 -2506 716 -2506 0 net=3877
rlabel metal2 716 -2506 716 -2506 0 net=3877
rlabel metal2 723 -2506 723 -2506 0 net=2307
rlabel metal2 740 -2506 740 -2506 0 net=4648
rlabel metal2 887 -2506 887 -2506 0 net=7486
rlabel metal2 933 -2506 933 -2506 0 net=3976
rlabel metal2 943 -2506 943 -2506 0 net=7530
rlabel metal2 100 -2508 100 -2508 0 net=5695
rlabel metal2 114 -2508 114 -2508 0 net=1501
rlabel metal2 149 -2508 149 -2508 0 net=3626
rlabel metal2 184 -2508 184 -2508 0 net=1661
rlabel metal2 191 -2508 191 -2508 0 net=6886
rlabel metal2 229 -2508 229 -2508 0 net=1414
rlabel metal2 254 -2508 254 -2508 0 net=1784
rlabel metal2 289 -2508 289 -2508 0 net=6674
rlabel metal2 394 -2508 394 -2508 0 net=1344
rlabel metal2 404 -2508 404 -2508 0 net=671
rlabel metal2 443 -2508 443 -2508 0 net=3371
rlabel metal2 604 -2508 604 -2508 0 net=7283
rlabel metal2 688 -2508 688 -2508 0 net=2264
rlabel metal2 688 -2508 688 -2508 0 net=2264
rlabel metal2 695 -2508 695 -2508 0 net=1360
rlabel metal2 744 -2508 744 -2508 0 net=6672
rlabel metal2 156 -2510 156 -2510 0 net=976
rlabel metal2 163 -2510 163 -2510 0 net=4124
rlabel metal2 177 -2510 177 -2510 0 net=4859
rlabel metal2 212 -2510 212 -2510 0 net=2980
rlabel metal2 261 -2510 261 -2510 0 net=5494
rlabel metal2 296 -2510 296 -2510 0 net=6899
rlabel metal2 401 -2510 401 -2510 0 net=304
rlabel metal2 163 -2512 163 -2512 0 net=6661
rlabel metal2 299 -2512 299 -2512 0 net=247
rlabel metal2 310 -2514 310 -2514 0 net=1393
rlabel metal2 5 -2525 5 -2525 0 net=5374
rlabel metal2 100 -2525 100 -2525 0 net=5696
rlabel metal2 114 -2525 114 -2525 0 net=1502
rlabel metal2 163 -2525 163 -2525 0 net=6662
rlabel metal2 180 -2525 180 -2525 0 net=1662
rlabel metal2 191 -2525 191 -2525 0 net=4860
rlabel metal2 292 -2525 292 -2525 0 net=6900
rlabel metal2 303 -2525 303 -2525 0 net=1394
rlabel metal2 341 -2525 341 -2525 0 net=2678
rlabel metal2 450 -2525 450 -2525 0 net=3372
rlabel metal2 597 -2525 597 -2525 0 net=7284
rlabel metal2 663 -2525 663 -2525 0 net=7090
rlabel metal2 716 -2525 716 -2525 0 net=3878
rlabel metal2 730 -2525 730 -2525 0 net=2308
rlabel metal2 121 -2527 121 -2527 0 net=806
<< end >>
