magic
tech scmos
timestamp 1555017675 
<< pdiffusion >>
rect 1 -10 7 -4
rect 8 -10 14 -4
rect 15 -10 21 -4
rect 22 -10 28 -4
rect 29 -10 35 -4
rect 36 -10 42 -4
rect 43 -10 49 -4
rect 176 -10 179 -4
rect 183 -10 186 -4
rect 190 -10 196 -4
rect 197 -10 203 -4
rect 211 -10 217 -4
rect 218 -10 221 -4
rect 232 -10 238 -4
rect 239 -10 242 -4
rect 253 -10 259 -4
rect 260 -10 263 -4
rect 274 -10 280 -4
rect 281 -10 287 -4
rect 288 -10 291 -4
rect 295 -10 301 -4
rect 302 -10 305 -4
rect 309 -10 315 -4
rect 316 -10 322 -4
rect 337 -10 340 -4
rect 344 -10 350 -4
rect 351 -10 354 -4
rect 358 -10 364 -4
rect 365 -10 368 -4
rect 407 -10 413 -4
rect 421 -10 427 -4
rect 456 -10 462 -4
rect 463 -10 469 -4
rect 470 -10 473 -4
rect 477 -10 483 -4
rect 484 -10 487 -4
rect 533 -10 539 -4
rect 540 -10 543 -4
rect 554 -10 560 -4
rect 575 -10 581 -4
rect 582 -10 585 -4
rect 603 -10 606 -4
rect 610 -10 616 -4
rect 617 -10 623 -4
rect 729 -10 732 -4
rect 736 -10 742 -4
rect 1 -27 7 -21
rect 8 -27 14 -21
rect 15 -27 21 -21
rect 22 -27 28 -21
rect 29 -27 35 -21
rect 36 -27 42 -21
rect 43 -27 49 -21
rect 50 -27 56 -21
rect 57 -27 63 -21
rect 64 -27 70 -21
rect 78 -27 84 -21
rect 113 -27 119 -21
rect 120 -27 123 -21
rect 127 -27 133 -21
rect 155 -27 161 -21
rect 162 -27 165 -21
rect 169 -27 172 -21
rect 176 -27 182 -21
rect 183 -27 186 -21
rect 211 -27 217 -21
rect 218 -27 221 -21
rect 225 -27 228 -21
rect 239 -27 242 -21
rect 246 -27 249 -21
rect 253 -27 256 -21
rect 260 -27 266 -21
rect 267 -27 273 -21
rect 274 -27 280 -21
rect 281 -27 284 -21
rect 288 -27 291 -21
rect 295 -27 298 -21
rect 302 -27 305 -21
rect 309 -27 312 -21
rect 316 -27 319 -21
rect 330 -27 336 -21
rect 337 -27 340 -21
rect 344 -27 347 -21
rect 351 -27 354 -21
rect 358 -27 361 -21
rect 365 -27 368 -21
rect 372 -27 378 -21
rect 379 -27 385 -21
rect 407 -27 413 -21
rect 414 -27 417 -21
rect 421 -27 427 -21
rect 428 -27 431 -21
rect 435 -27 441 -21
rect 442 -27 445 -21
rect 449 -27 452 -21
rect 456 -27 459 -21
rect 463 -27 469 -21
rect 470 -27 476 -21
rect 477 -27 480 -21
rect 484 -27 487 -21
rect 491 -27 494 -21
rect 526 -27 529 -21
rect 540 -27 543 -21
rect 575 -27 581 -21
rect 582 -27 585 -21
rect 603 -27 606 -21
rect 610 -27 613 -21
rect 617 -27 620 -21
rect 687 -27 690 -21
rect 694 -27 700 -21
rect 708 -27 714 -21
rect 729 -27 732 -21
rect 1 -50 7 -44
rect 8 -50 14 -44
rect 15 -50 21 -44
rect 22 -50 28 -44
rect 29 -50 35 -44
rect 57 -50 60 -44
rect 64 -50 70 -44
rect 78 -50 81 -44
rect 106 -50 112 -44
rect 113 -50 116 -44
rect 120 -50 126 -44
rect 127 -50 133 -44
rect 134 -50 137 -44
rect 141 -50 144 -44
rect 148 -50 154 -44
rect 155 -50 158 -44
rect 162 -50 165 -44
rect 169 -50 175 -44
rect 176 -50 179 -44
rect 183 -50 186 -44
rect 190 -50 196 -44
rect 197 -50 200 -44
rect 204 -50 210 -44
rect 211 -50 214 -44
rect 218 -50 224 -44
rect 225 -50 231 -44
rect 232 -50 235 -44
rect 239 -50 242 -44
rect 246 -50 249 -44
rect 253 -50 259 -44
rect 260 -50 263 -44
rect 267 -50 270 -44
rect 274 -50 277 -44
rect 281 -50 284 -44
rect 288 -50 291 -44
rect 295 -50 298 -44
rect 302 -50 305 -44
rect 309 -50 312 -44
rect 316 -50 319 -44
rect 323 -50 326 -44
rect 330 -50 336 -44
rect 337 -50 343 -44
rect 344 -50 347 -44
rect 351 -50 354 -44
rect 358 -50 361 -44
rect 365 -50 368 -44
rect 372 -50 375 -44
rect 379 -50 382 -44
rect 386 -50 392 -44
rect 393 -50 399 -44
rect 400 -50 403 -44
rect 407 -50 410 -44
rect 421 -50 427 -44
rect 428 -50 431 -44
rect 435 -50 438 -44
rect 442 -50 448 -44
rect 449 -50 452 -44
rect 456 -50 459 -44
rect 470 -50 473 -44
rect 477 -50 480 -44
rect 484 -50 487 -44
rect 498 -50 501 -44
rect 512 -50 515 -44
rect 533 -50 539 -44
rect 540 -50 546 -44
rect 547 -50 550 -44
rect 554 -50 557 -44
rect 561 -50 564 -44
rect 568 -50 574 -44
rect 575 -50 578 -44
rect 582 -50 585 -44
rect 589 -50 595 -44
rect 596 -50 599 -44
rect 603 -50 606 -44
rect 610 -50 613 -44
rect 624 -50 627 -44
rect 631 -50 634 -44
rect 645 -50 651 -44
rect 652 -50 658 -44
rect 659 -50 662 -44
rect 687 -50 690 -44
rect 729 -50 732 -44
rect 785 -50 788 -44
rect 806 -50 809 -44
rect 813 -50 819 -44
rect 897 -50 903 -44
rect 1 -89 7 -83
rect 8 -89 14 -83
rect 15 -89 21 -83
rect 22 -89 28 -83
rect 50 -89 56 -83
rect 57 -89 60 -83
rect 64 -89 67 -83
rect 78 -89 84 -83
rect 85 -89 91 -83
rect 92 -89 95 -83
rect 99 -89 105 -83
rect 106 -89 112 -83
rect 113 -89 116 -83
rect 120 -89 126 -83
rect 127 -89 130 -83
rect 134 -89 137 -83
rect 141 -89 144 -83
rect 148 -89 151 -83
rect 155 -89 158 -83
rect 162 -89 165 -83
rect 169 -89 172 -83
rect 176 -89 182 -83
rect 183 -89 189 -83
rect 190 -89 193 -83
rect 197 -89 200 -83
rect 204 -89 210 -83
rect 211 -89 214 -83
rect 218 -89 224 -83
rect 225 -89 231 -83
rect 232 -89 235 -83
rect 239 -89 242 -83
rect 246 -89 249 -83
rect 253 -89 256 -83
rect 260 -89 263 -83
rect 267 -89 270 -83
rect 274 -89 280 -83
rect 281 -89 284 -83
rect 288 -89 291 -83
rect 295 -89 301 -83
rect 302 -89 305 -83
rect 309 -89 312 -83
rect 316 -89 319 -83
rect 323 -89 326 -83
rect 330 -89 333 -83
rect 337 -89 340 -83
rect 344 -89 347 -83
rect 351 -89 354 -83
rect 358 -89 364 -83
rect 365 -89 368 -83
rect 372 -89 375 -83
rect 379 -89 382 -83
rect 386 -89 389 -83
rect 393 -89 399 -83
rect 400 -89 403 -83
rect 407 -89 410 -83
rect 414 -89 417 -83
rect 421 -89 424 -83
rect 428 -89 431 -83
rect 435 -89 441 -83
rect 442 -89 448 -83
rect 449 -89 452 -83
rect 456 -89 462 -83
rect 463 -89 469 -83
rect 470 -89 476 -83
rect 477 -89 480 -83
rect 484 -89 487 -83
rect 491 -89 497 -83
rect 498 -89 501 -83
rect 505 -89 508 -83
rect 512 -89 515 -83
rect 519 -89 522 -83
rect 526 -89 532 -83
rect 533 -89 536 -83
rect 540 -89 543 -83
rect 547 -89 550 -83
rect 554 -89 557 -83
rect 561 -89 564 -83
rect 568 -89 571 -83
rect 575 -89 578 -83
rect 582 -89 585 -83
rect 589 -89 592 -83
rect 596 -89 599 -83
rect 603 -89 606 -83
rect 610 -89 613 -83
rect 617 -89 620 -83
rect 624 -89 627 -83
rect 631 -89 637 -83
rect 638 -89 641 -83
rect 645 -89 648 -83
rect 652 -89 655 -83
rect 659 -89 662 -83
rect 673 -89 676 -83
rect 680 -89 686 -83
rect 701 -89 704 -83
rect 729 -89 732 -83
rect 792 -89 795 -83
rect 806 -89 809 -83
rect 897 -89 900 -83
rect 974 -89 980 -83
rect 1086 -89 1089 -83
rect 1093 -89 1099 -83
rect 1 -126 7 -120
rect 8 -126 14 -120
rect 15 -126 21 -120
rect 22 -126 28 -120
rect 29 -126 32 -120
rect 36 -126 42 -120
rect 43 -126 49 -120
rect 50 -126 53 -120
rect 57 -126 60 -120
rect 64 -126 67 -120
rect 71 -126 77 -120
rect 92 -126 95 -120
rect 99 -126 102 -120
rect 106 -126 109 -120
rect 113 -126 119 -120
rect 120 -126 123 -120
rect 127 -126 130 -120
rect 134 -126 140 -120
rect 141 -126 144 -120
rect 148 -126 151 -120
rect 155 -126 158 -120
rect 162 -126 165 -120
rect 169 -126 172 -120
rect 176 -126 182 -120
rect 183 -126 189 -120
rect 190 -126 193 -120
rect 197 -126 200 -120
rect 204 -126 207 -120
rect 211 -126 214 -120
rect 218 -126 221 -120
rect 225 -126 231 -120
rect 232 -126 235 -120
rect 239 -126 245 -120
rect 246 -126 252 -120
rect 253 -126 256 -120
rect 260 -126 263 -120
rect 267 -126 270 -120
rect 274 -126 277 -120
rect 281 -126 284 -120
rect 288 -126 294 -120
rect 295 -126 301 -120
rect 302 -126 305 -120
rect 309 -126 312 -120
rect 316 -126 319 -120
rect 323 -126 329 -120
rect 330 -126 333 -120
rect 337 -126 340 -120
rect 344 -126 347 -120
rect 351 -126 357 -120
rect 358 -126 361 -120
rect 365 -126 368 -120
rect 372 -126 378 -120
rect 379 -126 385 -120
rect 386 -126 389 -120
rect 393 -126 396 -120
rect 400 -126 403 -120
rect 407 -126 413 -120
rect 414 -126 417 -120
rect 421 -126 424 -120
rect 428 -126 431 -120
rect 435 -126 438 -120
rect 442 -126 445 -120
rect 449 -126 452 -120
rect 456 -126 459 -120
rect 463 -126 469 -120
rect 470 -126 473 -120
rect 477 -126 483 -120
rect 484 -126 487 -120
rect 491 -126 494 -120
rect 498 -126 501 -120
rect 505 -126 511 -120
rect 512 -126 515 -120
rect 519 -126 522 -120
rect 526 -126 529 -120
rect 533 -126 536 -120
rect 540 -126 543 -120
rect 547 -126 553 -120
rect 554 -126 560 -120
rect 561 -126 564 -120
rect 568 -126 571 -120
rect 575 -126 578 -120
rect 582 -126 585 -120
rect 589 -126 595 -120
rect 596 -126 599 -120
rect 603 -126 606 -120
rect 610 -126 613 -120
rect 617 -126 620 -120
rect 624 -126 627 -120
rect 631 -126 634 -120
rect 638 -126 641 -120
rect 645 -126 648 -120
rect 652 -126 658 -120
rect 659 -126 662 -120
rect 666 -126 669 -120
rect 673 -126 676 -120
rect 680 -126 683 -120
rect 687 -126 690 -120
rect 694 -126 697 -120
rect 701 -126 704 -120
rect 708 -126 714 -120
rect 715 -126 718 -120
rect 722 -126 725 -120
rect 729 -126 732 -120
rect 736 -126 739 -120
rect 757 -126 763 -120
rect 764 -126 767 -120
rect 778 -126 781 -120
rect 799 -126 802 -120
rect 904 -126 907 -120
rect 974 -126 977 -120
rect 1086 -126 1089 -120
rect 1 -187 7 -181
rect 8 -187 14 -181
rect 22 -187 25 -181
rect 29 -187 32 -181
rect 36 -187 42 -181
rect 43 -187 49 -181
rect 50 -187 53 -181
rect 57 -187 60 -181
rect 64 -187 70 -181
rect 71 -187 74 -181
rect 78 -187 81 -181
rect 85 -187 91 -181
rect 92 -187 95 -181
rect 99 -187 102 -181
rect 106 -187 109 -181
rect 113 -187 116 -181
rect 120 -187 123 -181
rect 127 -187 130 -181
rect 134 -187 140 -181
rect 141 -187 144 -181
rect 148 -187 151 -181
rect 155 -187 161 -181
rect 162 -187 168 -181
rect 169 -187 172 -181
rect 176 -187 179 -181
rect 183 -187 189 -181
rect 190 -187 193 -181
rect 197 -187 203 -181
rect 204 -187 210 -181
rect 211 -187 214 -181
rect 218 -187 221 -181
rect 225 -187 228 -181
rect 232 -187 235 -181
rect 239 -187 242 -181
rect 246 -187 249 -181
rect 253 -187 256 -181
rect 260 -187 263 -181
rect 267 -187 270 -181
rect 274 -187 277 -181
rect 281 -187 284 -181
rect 288 -187 291 -181
rect 295 -187 298 -181
rect 302 -187 305 -181
rect 309 -187 312 -181
rect 316 -187 322 -181
rect 323 -187 326 -181
rect 330 -187 336 -181
rect 337 -187 343 -181
rect 344 -187 350 -181
rect 351 -187 354 -181
rect 358 -187 361 -181
rect 365 -187 368 -181
rect 372 -187 378 -181
rect 379 -187 382 -181
rect 386 -187 392 -181
rect 393 -187 396 -181
rect 400 -187 403 -181
rect 407 -187 410 -181
rect 414 -187 417 -181
rect 421 -187 427 -181
rect 428 -187 431 -181
rect 435 -187 438 -181
rect 442 -187 445 -181
rect 449 -187 452 -181
rect 456 -187 459 -181
rect 463 -187 469 -181
rect 470 -187 473 -181
rect 477 -187 480 -181
rect 484 -187 490 -181
rect 491 -187 497 -181
rect 498 -187 501 -181
rect 505 -187 508 -181
rect 512 -187 515 -181
rect 519 -187 525 -181
rect 526 -187 529 -181
rect 533 -187 539 -181
rect 540 -187 543 -181
rect 547 -187 550 -181
rect 554 -187 557 -181
rect 561 -187 564 -181
rect 568 -187 571 -181
rect 575 -187 578 -181
rect 582 -187 585 -181
rect 589 -187 592 -181
rect 596 -187 599 -181
rect 603 -187 606 -181
rect 610 -187 613 -181
rect 617 -187 620 -181
rect 624 -187 627 -181
rect 631 -187 634 -181
rect 638 -187 641 -181
rect 645 -187 648 -181
rect 652 -187 655 -181
rect 659 -187 662 -181
rect 666 -187 669 -181
rect 673 -187 676 -181
rect 680 -187 683 -181
rect 687 -187 690 -181
rect 694 -187 697 -181
rect 701 -187 704 -181
rect 708 -187 711 -181
rect 715 -187 718 -181
rect 722 -187 725 -181
rect 729 -187 732 -181
rect 736 -187 739 -181
rect 743 -187 746 -181
rect 750 -187 753 -181
rect 757 -187 760 -181
rect 764 -187 767 -181
rect 771 -187 774 -181
rect 778 -187 781 -181
rect 785 -187 788 -181
rect 792 -187 795 -181
rect 799 -187 802 -181
rect 806 -187 809 -181
rect 813 -187 819 -181
rect 820 -187 826 -181
rect 827 -187 833 -181
rect 834 -187 840 -181
rect 841 -187 847 -181
rect 848 -187 851 -181
rect 855 -187 861 -181
rect 918 -187 921 -181
rect 974 -187 977 -181
rect 1086 -187 1089 -181
rect 1 -246 7 -240
rect 8 -246 14 -240
rect 15 -246 18 -240
rect 22 -246 25 -240
rect 29 -246 32 -240
rect 36 -246 39 -240
rect 43 -246 46 -240
rect 50 -246 53 -240
rect 57 -246 63 -240
rect 64 -246 70 -240
rect 71 -246 74 -240
rect 78 -246 81 -240
rect 85 -246 91 -240
rect 92 -246 98 -240
rect 99 -246 105 -240
rect 106 -246 112 -240
rect 113 -246 119 -240
rect 120 -246 123 -240
rect 127 -246 130 -240
rect 134 -246 137 -240
rect 141 -246 144 -240
rect 148 -246 151 -240
rect 155 -246 161 -240
rect 162 -246 165 -240
rect 169 -246 175 -240
rect 176 -246 179 -240
rect 183 -246 189 -240
rect 190 -246 193 -240
rect 197 -246 203 -240
rect 204 -246 207 -240
rect 211 -246 214 -240
rect 218 -246 224 -240
rect 225 -246 231 -240
rect 232 -246 235 -240
rect 239 -246 242 -240
rect 246 -246 249 -240
rect 253 -246 256 -240
rect 260 -246 266 -240
rect 267 -246 270 -240
rect 274 -246 277 -240
rect 281 -246 287 -240
rect 288 -246 294 -240
rect 295 -246 298 -240
rect 302 -246 305 -240
rect 309 -246 312 -240
rect 316 -246 319 -240
rect 323 -246 326 -240
rect 330 -246 333 -240
rect 337 -246 340 -240
rect 344 -246 347 -240
rect 351 -246 357 -240
rect 358 -246 361 -240
rect 365 -246 368 -240
rect 372 -246 375 -240
rect 379 -246 385 -240
rect 386 -246 389 -240
rect 393 -246 396 -240
rect 400 -246 403 -240
rect 407 -246 410 -240
rect 414 -246 417 -240
rect 421 -246 424 -240
rect 428 -246 431 -240
rect 435 -246 438 -240
rect 442 -246 445 -240
rect 449 -246 452 -240
rect 456 -246 462 -240
rect 463 -246 469 -240
rect 470 -246 473 -240
rect 477 -246 483 -240
rect 484 -246 490 -240
rect 491 -246 497 -240
rect 498 -246 501 -240
rect 505 -246 508 -240
rect 512 -246 515 -240
rect 519 -246 522 -240
rect 526 -246 529 -240
rect 533 -246 536 -240
rect 540 -246 543 -240
rect 547 -246 550 -240
rect 554 -246 557 -240
rect 561 -246 564 -240
rect 568 -246 571 -240
rect 575 -246 578 -240
rect 582 -246 585 -240
rect 589 -246 595 -240
rect 596 -246 602 -240
rect 603 -246 606 -240
rect 610 -246 613 -240
rect 617 -246 620 -240
rect 624 -246 627 -240
rect 631 -246 634 -240
rect 638 -246 641 -240
rect 645 -246 651 -240
rect 652 -246 655 -240
rect 659 -246 662 -240
rect 666 -246 669 -240
rect 673 -246 676 -240
rect 680 -246 683 -240
rect 687 -246 690 -240
rect 694 -246 697 -240
rect 701 -246 704 -240
rect 708 -246 711 -240
rect 715 -246 718 -240
rect 722 -246 725 -240
rect 729 -246 732 -240
rect 736 -246 739 -240
rect 743 -246 746 -240
rect 750 -246 753 -240
rect 757 -246 760 -240
rect 764 -246 767 -240
rect 771 -246 774 -240
rect 778 -246 781 -240
rect 785 -246 788 -240
rect 792 -246 795 -240
rect 799 -246 805 -240
rect 806 -246 809 -240
rect 813 -246 816 -240
rect 820 -246 823 -240
rect 827 -246 830 -240
rect 834 -246 837 -240
rect 841 -246 844 -240
rect 848 -246 851 -240
rect 855 -246 858 -240
rect 862 -246 865 -240
rect 869 -246 872 -240
rect 876 -246 879 -240
rect 883 -246 886 -240
rect 890 -246 893 -240
rect 897 -246 900 -240
rect 904 -246 907 -240
rect 911 -246 914 -240
rect 918 -246 921 -240
rect 925 -246 928 -240
rect 932 -246 935 -240
rect 939 -246 942 -240
rect 946 -246 949 -240
rect 953 -246 959 -240
rect 974 -246 977 -240
rect 1086 -246 1089 -240
rect 1 -317 7 -311
rect 8 -317 14 -311
rect 15 -317 18 -311
rect 22 -317 25 -311
rect 29 -317 35 -311
rect 36 -317 39 -311
rect 43 -317 49 -311
rect 50 -317 56 -311
rect 57 -317 60 -311
rect 64 -317 67 -311
rect 71 -317 74 -311
rect 78 -317 84 -311
rect 85 -317 88 -311
rect 92 -317 95 -311
rect 99 -317 102 -311
rect 106 -317 112 -311
rect 113 -317 116 -311
rect 120 -317 123 -311
rect 127 -317 130 -311
rect 134 -317 137 -311
rect 141 -317 147 -311
rect 148 -317 151 -311
rect 155 -317 158 -311
rect 162 -317 168 -311
rect 169 -317 172 -311
rect 176 -317 179 -311
rect 183 -317 186 -311
rect 190 -317 196 -311
rect 197 -317 200 -311
rect 204 -317 210 -311
rect 211 -317 214 -311
rect 218 -317 221 -311
rect 225 -317 231 -311
rect 232 -317 235 -311
rect 239 -317 242 -311
rect 246 -317 249 -311
rect 253 -317 256 -311
rect 260 -317 263 -311
rect 267 -317 270 -311
rect 274 -317 277 -311
rect 281 -317 284 -311
rect 288 -317 294 -311
rect 295 -317 298 -311
rect 302 -317 305 -311
rect 309 -317 312 -311
rect 316 -317 319 -311
rect 323 -317 326 -311
rect 330 -317 333 -311
rect 337 -317 340 -311
rect 344 -317 347 -311
rect 351 -317 354 -311
rect 358 -317 361 -311
rect 365 -317 368 -311
rect 372 -317 375 -311
rect 379 -317 385 -311
rect 386 -317 392 -311
rect 393 -317 396 -311
rect 400 -317 403 -311
rect 407 -317 413 -311
rect 414 -317 420 -311
rect 421 -317 424 -311
rect 428 -317 431 -311
rect 435 -317 441 -311
rect 442 -317 445 -311
rect 449 -317 452 -311
rect 456 -317 459 -311
rect 463 -317 469 -311
rect 470 -317 476 -311
rect 477 -317 480 -311
rect 484 -317 490 -311
rect 491 -317 494 -311
rect 498 -317 501 -311
rect 505 -317 511 -311
rect 512 -317 515 -311
rect 519 -317 522 -311
rect 526 -317 529 -311
rect 533 -317 536 -311
rect 540 -317 546 -311
rect 547 -317 553 -311
rect 554 -317 557 -311
rect 561 -317 564 -311
rect 568 -317 571 -311
rect 575 -317 581 -311
rect 582 -317 588 -311
rect 589 -317 592 -311
rect 596 -317 599 -311
rect 603 -317 606 -311
rect 610 -317 613 -311
rect 617 -317 620 -311
rect 624 -317 627 -311
rect 631 -317 634 -311
rect 638 -317 641 -311
rect 645 -317 648 -311
rect 652 -317 655 -311
rect 659 -317 662 -311
rect 666 -317 669 -311
rect 673 -317 676 -311
rect 680 -317 683 -311
rect 687 -317 690 -311
rect 694 -317 697 -311
rect 701 -317 704 -311
rect 708 -317 711 -311
rect 715 -317 721 -311
rect 722 -317 725 -311
rect 729 -317 732 -311
rect 736 -317 739 -311
rect 743 -317 746 -311
rect 750 -317 753 -311
rect 757 -317 760 -311
rect 764 -317 767 -311
rect 771 -317 774 -311
rect 778 -317 781 -311
rect 785 -317 788 -311
rect 792 -317 795 -311
rect 799 -317 802 -311
rect 806 -317 809 -311
rect 813 -317 816 -311
rect 820 -317 823 -311
rect 827 -317 830 -311
rect 834 -317 837 -311
rect 841 -317 844 -311
rect 848 -317 851 -311
rect 855 -317 858 -311
rect 862 -317 865 -311
rect 869 -317 872 -311
rect 876 -317 879 -311
rect 883 -317 886 -311
rect 890 -317 893 -311
rect 897 -317 900 -311
rect 904 -317 907 -311
rect 911 -317 914 -311
rect 918 -317 921 -311
rect 925 -317 928 -311
rect 932 -317 938 -311
rect 939 -317 942 -311
rect 946 -317 952 -311
rect 953 -317 956 -311
rect 960 -317 963 -311
rect 967 -317 973 -311
rect 974 -317 977 -311
rect 981 -317 984 -311
rect 1093 -317 1096 -311
rect 1 -402 7 -396
rect 15 -402 18 -396
rect 22 -402 25 -396
rect 29 -402 35 -396
rect 36 -402 42 -396
rect 43 -402 46 -396
rect 50 -402 53 -396
rect 57 -402 60 -396
rect 64 -402 67 -396
rect 71 -402 74 -396
rect 78 -402 81 -396
rect 85 -402 88 -396
rect 92 -402 95 -396
rect 99 -402 102 -396
rect 106 -402 109 -396
rect 113 -402 119 -396
rect 120 -402 123 -396
rect 127 -402 130 -396
rect 134 -402 140 -396
rect 141 -402 147 -396
rect 148 -402 151 -396
rect 155 -402 158 -396
rect 162 -402 165 -396
rect 169 -402 175 -396
rect 176 -402 182 -396
rect 183 -402 186 -396
rect 190 -402 193 -396
rect 197 -402 200 -396
rect 204 -402 210 -396
rect 211 -402 214 -396
rect 218 -402 221 -396
rect 225 -402 228 -396
rect 232 -402 235 -396
rect 239 -402 242 -396
rect 246 -402 249 -396
rect 253 -402 256 -396
rect 260 -402 263 -396
rect 267 -402 270 -396
rect 274 -402 280 -396
rect 281 -402 284 -396
rect 288 -402 291 -396
rect 295 -402 298 -396
rect 302 -402 305 -396
rect 309 -402 312 -396
rect 316 -402 322 -396
rect 323 -402 326 -396
rect 330 -402 333 -396
rect 337 -402 343 -396
rect 344 -402 347 -396
rect 351 -402 354 -396
rect 358 -402 364 -396
rect 365 -402 368 -396
rect 372 -402 375 -396
rect 379 -402 382 -396
rect 386 -402 389 -396
rect 393 -402 396 -396
rect 400 -402 406 -396
rect 407 -402 410 -396
rect 414 -402 417 -396
rect 421 -402 427 -396
rect 428 -402 431 -396
rect 435 -402 438 -396
rect 442 -402 445 -396
rect 449 -402 455 -396
rect 456 -402 459 -396
rect 463 -402 466 -396
rect 470 -402 476 -396
rect 477 -402 480 -396
rect 484 -402 487 -396
rect 491 -402 497 -396
rect 498 -402 501 -396
rect 505 -402 511 -396
rect 512 -402 515 -396
rect 519 -402 525 -396
rect 526 -402 529 -396
rect 533 -402 536 -396
rect 540 -402 543 -396
rect 547 -402 553 -396
rect 554 -402 557 -396
rect 561 -402 567 -396
rect 568 -402 571 -396
rect 575 -402 581 -396
rect 582 -402 585 -396
rect 589 -402 592 -396
rect 596 -402 599 -396
rect 603 -402 606 -396
rect 610 -402 613 -396
rect 617 -402 620 -396
rect 624 -402 627 -396
rect 631 -402 634 -396
rect 638 -402 641 -396
rect 645 -402 648 -396
rect 652 -402 655 -396
rect 659 -402 662 -396
rect 666 -402 669 -396
rect 673 -402 676 -396
rect 680 -402 686 -396
rect 687 -402 690 -396
rect 694 -402 697 -396
rect 701 -402 704 -396
rect 708 -402 711 -396
rect 715 -402 718 -396
rect 722 -402 725 -396
rect 729 -402 732 -396
rect 736 -402 739 -396
rect 743 -402 746 -396
rect 750 -402 753 -396
rect 757 -402 760 -396
rect 764 -402 767 -396
rect 771 -402 774 -396
rect 778 -402 781 -396
rect 785 -402 788 -396
rect 792 -402 795 -396
rect 799 -402 802 -396
rect 806 -402 809 -396
rect 813 -402 816 -396
rect 820 -402 823 -396
rect 827 -402 830 -396
rect 834 -402 837 -396
rect 841 -402 844 -396
rect 848 -402 851 -396
rect 855 -402 858 -396
rect 862 -402 865 -396
rect 869 -402 872 -396
rect 876 -402 879 -396
rect 883 -402 886 -396
rect 890 -402 893 -396
rect 897 -402 903 -396
rect 904 -402 907 -396
rect 911 -402 914 -396
rect 918 -402 921 -396
rect 925 -402 928 -396
rect 932 -402 935 -396
rect 939 -402 942 -396
rect 946 -402 949 -396
rect 953 -402 956 -396
rect 960 -402 966 -396
rect 967 -402 970 -396
rect 974 -402 977 -396
rect 981 -402 984 -396
rect 988 -402 991 -396
rect 995 -402 1001 -396
rect 1002 -402 1005 -396
rect 1009 -402 1012 -396
rect 1016 -402 1019 -396
rect 1023 -402 1026 -396
rect 1030 -402 1036 -396
rect 1037 -402 1043 -396
rect 1044 -402 1050 -396
rect 1051 -402 1054 -396
rect 1065 -402 1068 -396
rect 1107 -402 1110 -396
rect 1 -471 7 -465
rect 8 -471 14 -465
rect 15 -471 18 -465
rect 22 -471 25 -465
rect 29 -471 32 -465
rect 36 -471 39 -465
rect 43 -471 46 -465
rect 50 -471 53 -465
rect 57 -471 60 -465
rect 64 -471 67 -465
rect 71 -471 74 -465
rect 78 -471 81 -465
rect 85 -471 91 -465
rect 92 -471 95 -465
rect 99 -471 102 -465
rect 106 -471 112 -465
rect 113 -471 116 -465
rect 120 -471 123 -465
rect 127 -471 130 -465
rect 134 -471 140 -465
rect 141 -471 144 -465
rect 148 -471 151 -465
rect 155 -471 158 -465
rect 162 -471 165 -465
rect 169 -471 172 -465
rect 176 -471 179 -465
rect 183 -471 186 -465
rect 190 -471 193 -465
rect 197 -471 200 -465
rect 204 -471 207 -465
rect 211 -471 217 -465
rect 218 -471 221 -465
rect 225 -471 231 -465
rect 232 -471 235 -465
rect 239 -471 242 -465
rect 246 -471 249 -465
rect 253 -471 256 -465
rect 260 -471 263 -465
rect 267 -471 270 -465
rect 274 -471 280 -465
rect 281 -471 284 -465
rect 288 -471 291 -465
rect 295 -471 298 -465
rect 302 -471 308 -465
rect 309 -471 312 -465
rect 316 -471 319 -465
rect 323 -471 326 -465
rect 330 -471 333 -465
rect 337 -471 340 -465
rect 344 -471 350 -465
rect 351 -471 354 -465
rect 358 -471 361 -465
rect 365 -471 368 -465
rect 372 -471 375 -465
rect 379 -471 382 -465
rect 386 -471 392 -465
rect 393 -471 396 -465
rect 400 -471 406 -465
rect 407 -471 413 -465
rect 414 -471 417 -465
rect 421 -471 424 -465
rect 428 -471 431 -465
rect 435 -471 438 -465
rect 442 -471 445 -465
rect 449 -471 452 -465
rect 456 -471 462 -465
rect 463 -471 466 -465
rect 470 -471 476 -465
rect 477 -471 480 -465
rect 484 -471 487 -465
rect 491 -471 494 -465
rect 498 -471 504 -465
rect 505 -471 511 -465
rect 512 -471 515 -465
rect 519 -471 525 -465
rect 526 -471 532 -465
rect 533 -471 536 -465
rect 540 -471 543 -465
rect 547 -471 550 -465
rect 554 -471 557 -465
rect 561 -471 567 -465
rect 568 -471 571 -465
rect 575 -471 578 -465
rect 582 -471 588 -465
rect 589 -471 592 -465
rect 596 -471 602 -465
rect 603 -471 606 -465
rect 610 -471 613 -465
rect 617 -471 620 -465
rect 624 -471 627 -465
rect 631 -471 637 -465
rect 638 -471 641 -465
rect 645 -471 648 -465
rect 652 -471 655 -465
rect 659 -471 665 -465
rect 666 -471 669 -465
rect 673 -471 676 -465
rect 680 -471 683 -465
rect 687 -471 690 -465
rect 694 -471 697 -465
rect 701 -471 704 -465
rect 708 -471 711 -465
rect 715 -471 718 -465
rect 722 -471 728 -465
rect 729 -471 732 -465
rect 736 -471 742 -465
rect 743 -471 746 -465
rect 750 -471 756 -465
rect 757 -471 760 -465
rect 764 -471 767 -465
rect 771 -471 774 -465
rect 778 -471 781 -465
rect 785 -471 788 -465
rect 792 -471 795 -465
rect 799 -471 802 -465
rect 806 -471 809 -465
rect 813 -471 816 -465
rect 820 -471 823 -465
rect 827 -471 830 -465
rect 834 -471 837 -465
rect 841 -471 844 -465
rect 848 -471 851 -465
rect 855 -471 858 -465
rect 862 -471 865 -465
rect 869 -471 872 -465
rect 876 -471 879 -465
rect 883 -471 886 -465
rect 890 -471 893 -465
rect 897 -471 900 -465
rect 904 -471 907 -465
rect 911 -471 914 -465
rect 918 -471 921 -465
rect 925 -471 928 -465
rect 932 -471 935 -465
rect 939 -471 942 -465
rect 946 -471 949 -465
rect 953 -471 956 -465
rect 960 -471 963 -465
rect 967 -471 970 -465
rect 974 -471 977 -465
rect 981 -471 987 -465
rect 988 -471 991 -465
rect 995 -471 998 -465
rect 1002 -471 1005 -465
rect 1009 -471 1012 -465
rect 1016 -471 1019 -465
rect 1023 -471 1026 -465
rect 1030 -471 1033 -465
rect 1037 -471 1040 -465
rect 1044 -471 1047 -465
rect 1051 -471 1054 -465
rect 1058 -471 1061 -465
rect 1065 -471 1068 -465
rect 1072 -471 1075 -465
rect 1079 -471 1082 -465
rect 1086 -471 1089 -465
rect 1093 -471 1096 -465
rect 1100 -471 1103 -465
rect 1107 -471 1110 -465
rect 1114 -471 1117 -465
rect 1121 -471 1124 -465
rect 1128 -471 1131 -465
rect 1135 -471 1141 -465
rect 1142 -471 1148 -465
rect 1149 -471 1152 -465
rect 1 -566 7 -560
rect 8 -566 11 -560
rect 15 -566 18 -560
rect 22 -566 25 -560
rect 29 -566 35 -560
rect 36 -566 39 -560
rect 43 -566 46 -560
rect 50 -566 53 -560
rect 57 -566 60 -560
rect 64 -566 67 -560
rect 71 -566 77 -560
rect 78 -566 84 -560
rect 85 -566 88 -560
rect 92 -566 95 -560
rect 99 -566 102 -560
rect 106 -566 112 -560
rect 113 -566 116 -560
rect 120 -566 123 -560
rect 127 -566 130 -560
rect 134 -566 137 -560
rect 141 -566 144 -560
rect 148 -566 154 -560
rect 155 -566 158 -560
rect 162 -566 168 -560
rect 169 -566 172 -560
rect 176 -566 179 -560
rect 183 -566 186 -560
rect 190 -566 196 -560
rect 197 -566 203 -560
rect 204 -566 207 -560
rect 211 -566 217 -560
rect 218 -566 221 -560
rect 225 -566 228 -560
rect 232 -566 235 -560
rect 239 -566 242 -560
rect 246 -566 249 -560
rect 253 -566 256 -560
rect 260 -566 263 -560
rect 267 -566 270 -560
rect 274 -566 277 -560
rect 281 -566 284 -560
rect 288 -566 291 -560
rect 295 -566 298 -560
rect 302 -566 305 -560
rect 309 -566 312 -560
rect 316 -566 322 -560
rect 323 -566 326 -560
rect 330 -566 333 -560
rect 337 -566 340 -560
rect 344 -566 347 -560
rect 351 -566 357 -560
rect 358 -566 361 -560
rect 365 -566 371 -560
rect 372 -566 375 -560
rect 379 -566 382 -560
rect 386 -566 392 -560
rect 393 -566 399 -560
rect 400 -566 403 -560
rect 407 -566 413 -560
rect 414 -566 417 -560
rect 421 -566 427 -560
rect 428 -566 431 -560
rect 435 -566 438 -560
rect 442 -566 445 -560
rect 449 -566 452 -560
rect 456 -566 459 -560
rect 463 -566 466 -560
rect 470 -566 473 -560
rect 477 -566 480 -560
rect 484 -566 487 -560
rect 491 -566 494 -560
rect 498 -566 501 -560
rect 505 -566 511 -560
rect 512 -566 515 -560
rect 519 -566 522 -560
rect 526 -566 529 -560
rect 533 -566 539 -560
rect 540 -566 543 -560
rect 547 -566 553 -560
rect 554 -566 557 -560
rect 561 -566 567 -560
rect 568 -566 574 -560
rect 575 -566 578 -560
rect 582 -566 585 -560
rect 589 -566 595 -560
rect 596 -566 602 -560
rect 603 -566 609 -560
rect 610 -566 613 -560
rect 617 -566 620 -560
rect 624 -566 630 -560
rect 631 -566 634 -560
rect 638 -566 641 -560
rect 645 -566 648 -560
rect 652 -566 655 -560
rect 659 -566 665 -560
rect 666 -566 669 -560
rect 673 -566 676 -560
rect 680 -566 683 -560
rect 687 -566 690 -560
rect 694 -566 697 -560
rect 701 -566 704 -560
rect 708 -566 714 -560
rect 715 -566 718 -560
rect 722 -566 725 -560
rect 729 -566 735 -560
rect 736 -566 739 -560
rect 743 -566 746 -560
rect 750 -566 753 -560
rect 757 -566 760 -560
rect 764 -566 767 -560
rect 771 -566 774 -560
rect 778 -566 781 -560
rect 785 -566 788 -560
rect 792 -566 795 -560
rect 799 -566 802 -560
rect 806 -566 809 -560
rect 813 -566 816 -560
rect 820 -566 823 -560
rect 827 -566 830 -560
rect 834 -566 837 -560
rect 841 -566 844 -560
rect 848 -566 851 -560
rect 855 -566 858 -560
rect 862 -566 865 -560
rect 869 -566 872 -560
rect 876 -566 879 -560
rect 883 -566 886 -560
rect 890 -566 893 -560
rect 897 -566 900 -560
rect 904 -566 907 -560
rect 911 -566 914 -560
rect 918 -566 921 -560
rect 925 -566 928 -560
rect 932 -566 935 -560
rect 939 -566 942 -560
rect 946 -566 949 -560
rect 953 -566 956 -560
rect 960 -566 963 -560
rect 967 -566 970 -560
rect 974 -566 977 -560
rect 981 -566 984 -560
rect 988 -566 991 -560
rect 995 -566 998 -560
rect 1002 -566 1005 -560
rect 1009 -566 1012 -560
rect 1016 -566 1019 -560
rect 1023 -566 1026 -560
rect 1030 -566 1033 -560
rect 1037 -566 1040 -560
rect 1044 -566 1047 -560
rect 1051 -566 1054 -560
rect 1058 -566 1061 -560
rect 1065 -566 1068 -560
rect 1072 -566 1075 -560
rect 1079 -566 1082 -560
rect 1086 -566 1089 -560
rect 1093 -566 1096 -560
rect 1100 -566 1103 -560
rect 1114 -566 1117 -560
rect 1121 -566 1124 -560
rect 1170 -566 1176 -560
rect 1177 -566 1180 -560
rect 1 -657 7 -651
rect 8 -657 11 -651
rect 15 -657 18 -651
rect 22 -657 28 -651
rect 29 -657 32 -651
rect 36 -657 39 -651
rect 43 -657 46 -651
rect 50 -657 56 -651
rect 57 -657 60 -651
rect 64 -657 70 -651
rect 71 -657 74 -651
rect 78 -657 84 -651
rect 85 -657 91 -651
rect 92 -657 95 -651
rect 99 -657 105 -651
rect 106 -657 109 -651
rect 113 -657 119 -651
rect 120 -657 123 -651
rect 127 -657 133 -651
rect 134 -657 137 -651
rect 141 -657 144 -651
rect 148 -657 151 -651
rect 155 -657 161 -651
rect 162 -657 165 -651
rect 169 -657 172 -651
rect 176 -657 179 -651
rect 183 -657 189 -651
rect 190 -657 193 -651
rect 197 -657 200 -651
rect 204 -657 210 -651
rect 211 -657 214 -651
rect 218 -657 221 -651
rect 225 -657 228 -651
rect 232 -657 238 -651
rect 239 -657 242 -651
rect 246 -657 249 -651
rect 253 -657 256 -651
rect 260 -657 263 -651
rect 267 -657 270 -651
rect 274 -657 277 -651
rect 281 -657 284 -651
rect 288 -657 291 -651
rect 295 -657 298 -651
rect 302 -657 305 -651
rect 309 -657 312 -651
rect 316 -657 319 -651
rect 323 -657 326 -651
rect 330 -657 336 -651
rect 337 -657 343 -651
rect 344 -657 350 -651
rect 351 -657 354 -651
rect 358 -657 361 -651
rect 365 -657 368 -651
rect 372 -657 375 -651
rect 379 -657 382 -651
rect 386 -657 389 -651
rect 393 -657 396 -651
rect 400 -657 403 -651
rect 407 -657 413 -651
rect 414 -657 420 -651
rect 421 -657 424 -651
rect 428 -657 431 -651
rect 435 -657 438 -651
rect 442 -657 448 -651
rect 449 -657 452 -651
rect 456 -657 459 -651
rect 463 -657 466 -651
rect 470 -657 473 -651
rect 477 -657 483 -651
rect 484 -657 487 -651
rect 491 -657 494 -651
rect 498 -657 504 -651
rect 505 -657 508 -651
rect 512 -657 518 -651
rect 519 -657 525 -651
rect 526 -657 529 -651
rect 533 -657 536 -651
rect 540 -657 543 -651
rect 547 -657 553 -651
rect 554 -657 557 -651
rect 561 -657 564 -651
rect 568 -657 571 -651
rect 575 -657 578 -651
rect 582 -657 585 -651
rect 589 -657 592 -651
rect 596 -657 599 -651
rect 603 -657 609 -651
rect 610 -657 616 -651
rect 617 -657 620 -651
rect 624 -657 627 -651
rect 631 -657 634 -651
rect 638 -657 641 -651
rect 645 -657 648 -651
rect 652 -657 658 -651
rect 659 -657 662 -651
rect 666 -657 669 -651
rect 673 -657 676 -651
rect 680 -657 683 -651
rect 687 -657 693 -651
rect 694 -657 697 -651
rect 701 -657 704 -651
rect 708 -657 711 -651
rect 715 -657 718 -651
rect 722 -657 725 -651
rect 729 -657 732 -651
rect 736 -657 739 -651
rect 743 -657 746 -651
rect 750 -657 753 -651
rect 757 -657 763 -651
rect 764 -657 767 -651
rect 771 -657 774 -651
rect 778 -657 781 -651
rect 785 -657 788 -651
rect 792 -657 795 -651
rect 799 -657 802 -651
rect 806 -657 809 -651
rect 813 -657 816 -651
rect 820 -657 823 -651
rect 827 -657 830 -651
rect 834 -657 837 -651
rect 841 -657 844 -651
rect 848 -657 851 -651
rect 855 -657 858 -651
rect 862 -657 865 -651
rect 869 -657 872 -651
rect 876 -657 879 -651
rect 883 -657 886 -651
rect 890 -657 893 -651
rect 897 -657 900 -651
rect 904 -657 907 -651
rect 911 -657 914 -651
rect 918 -657 921 -651
rect 925 -657 928 -651
rect 932 -657 938 -651
rect 939 -657 942 -651
rect 946 -657 949 -651
rect 953 -657 956 -651
rect 960 -657 963 -651
rect 967 -657 970 -651
rect 974 -657 977 -651
rect 981 -657 984 -651
rect 988 -657 991 -651
rect 995 -657 998 -651
rect 1002 -657 1005 -651
rect 1009 -657 1012 -651
rect 1016 -657 1019 -651
rect 1023 -657 1026 -651
rect 1030 -657 1033 -651
rect 1037 -657 1040 -651
rect 1044 -657 1047 -651
rect 1051 -657 1054 -651
rect 1058 -657 1061 -651
rect 1065 -657 1068 -651
rect 1072 -657 1075 -651
rect 1079 -657 1082 -651
rect 1086 -657 1089 -651
rect 1093 -657 1096 -651
rect 1100 -657 1103 -651
rect 1107 -657 1110 -651
rect 1114 -657 1117 -651
rect 1121 -657 1124 -651
rect 1128 -657 1131 -651
rect 1135 -657 1138 -651
rect 1177 -657 1180 -651
rect 8 -738 11 -732
rect 15 -738 18 -732
rect 22 -738 25 -732
rect 29 -738 35 -732
rect 36 -738 39 -732
rect 43 -738 46 -732
rect 50 -738 53 -732
rect 57 -738 60 -732
rect 64 -738 67 -732
rect 71 -738 77 -732
rect 78 -738 81 -732
rect 85 -738 88 -732
rect 92 -738 95 -732
rect 99 -738 102 -732
rect 106 -738 109 -732
rect 113 -738 116 -732
rect 120 -738 126 -732
rect 127 -738 130 -732
rect 134 -738 140 -732
rect 141 -738 144 -732
rect 148 -738 154 -732
rect 155 -738 158 -732
rect 162 -738 165 -732
rect 169 -738 172 -732
rect 176 -738 179 -732
rect 183 -738 189 -732
rect 190 -738 196 -732
rect 197 -738 200 -732
rect 204 -738 210 -732
rect 211 -738 214 -732
rect 218 -738 221 -732
rect 225 -738 228 -732
rect 232 -738 235 -732
rect 239 -738 242 -732
rect 246 -738 249 -732
rect 253 -738 256 -732
rect 260 -738 263 -732
rect 267 -738 270 -732
rect 274 -738 277 -732
rect 281 -738 284 -732
rect 288 -738 291 -732
rect 295 -738 298 -732
rect 302 -738 305 -732
rect 309 -738 315 -732
rect 316 -738 319 -732
rect 323 -738 326 -732
rect 330 -738 333 -732
rect 337 -738 343 -732
rect 344 -738 347 -732
rect 351 -738 354 -732
rect 358 -738 364 -732
rect 365 -738 368 -732
rect 372 -738 375 -732
rect 379 -738 382 -732
rect 386 -738 389 -732
rect 393 -738 399 -732
rect 400 -738 406 -732
rect 407 -738 413 -732
rect 414 -738 417 -732
rect 421 -738 427 -732
rect 428 -738 431 -732
rect 435 -738 441 -732
rect 442 -738 445 -732
rect 449 -738 452 -732
rect 456 -738 459 -732
rect 463 -738 469 -732
rect 470 -738 476 -732
rect 477 -738 480 -732
rect 484 -738 487 -732
rect 491 -738 494 -732
rect 498 -738 501 -732
rect 505 -738 508 -732
rect 512 -738 515 -732
rect 519 -738 525 -732
rect 526 -738 529 -732
rect 533 -738 536 -732
rect 540 -738 543 -732
rect 547 -738 553 -732
rect 554 -738 557 -732
rect 561 -738 564 -732
rect 568 -738 571 -732
rect 575 -738 578 -732
rect 582 -738 585 -732
rect 589 -738 592 -732
rect 596 -738 602 -732
rect 603 -738 609 -732
rect 610 -738 613 -732
rect 617 -738 620 -732
rect 624 -738 627 -732
rect 631 -738 637 -732
rect 638 -738 644 -732
rect 645 -738 648 -732
rect 652 -738 655 -732
rect 659 -738 662 -732
rect 666 -738 669 -732
rect 673 -738 676 -732
rect 680 -738 683 -732
rect 687 -738 693 -732
rect 694 -738 697 -732
rect 701 -738 704 -732
rect 708 -738 711 -732
rect 715 -738 721 -732
rect 722 -738 725 -732
rect 729 -738 732 -732
rect 736 -738 739 -732
rect 743 -738 749 -732
rect 750 -738 753 -732
rect 757 -738 760 -732
rect 764 -738 767 -732
rect 771 -738 774 -732
rect 778 -738 781 -732
rect 785 -738 788 -732
rect 792 -738 795 -732
rect 799 -738 802 -732
rect 806 -738 809 -732
rect 813 -738 816 -732
rect 820 -738 823 -732
rect 827 -738 830 -732
rect 834 -738 837 -732
rect 841 -738 844 -732
rect 848 -738 851 -732
rect 855 -738 858 -732
rect 862 -738 865 -732
rect 869 -738 872 -732
rect 876 -738 879 -732
rect 883 -738 886 -732
rect 890 -738 893 -732
rect 897 -738 900 -732
rect 904 -738 907 -732
rect 911 -738 914 -732
rect 918 -738 921 -732
rect 925 -738 928 -732
rect 932 -738 935 -732
rect 939 -738 942 -732
rect 946 -738 949 -732
rect 953 -738 956 -732
rect 960 -738 963 -732
rect 967 -738 970 -732
rect 974 -738 977 -732
rect 981 -738 984 -732
rect 988 -738 991 -732
rect 995 -738 998 -732
rect 1002 -738 1005 -732
rect 1009 -738 1012 -732
rect 1016 -738 1019 -732
rect 1023 -738 1026 -732
rect 1030 -738 1033 -732
rect 1037 -738 1040 -732
rect 1044 -738 1047 -732
rect 1051 -738 1054 -732
rect 1058 -738 1061 -732
rect 1065 -738 1068 -732
rect 1072 -738 1075 -732
rect 1079 -738 1082 -732
rect 1086 -738 1092 -732
rect 1093 -738 1096 -732
rect 1100 -738 1103 -732
rect 1107 -738 1113 -732
rect 1114 -738 1117 -732
rect 1121 -738 1124 -732
rect 1128 -738 1131 -732
rect 1135 -738 1138 -732
rect 1142 -738 1145 -732
rect 1149 -738 1152 -732
rect 1156 -738 1162 -732
rect 1163 -738 1166 -732
rect 1170 -738 1173 -732
rect 1184 -738 1187 -732
rect 1 -827 7 -821
rect 8 -827 11 -821
rect 15 -827 18 -821
rect 22 -827 25 -821
rect 29 -827 32 -821
rect 36 -827 39 -821
rect 43 -827 46 -821
rect 50 -827 53 -821
rect 57 -827 60 -821
rect 64 -827 67 -821
rect 71 -827 77 -821
rect 78 -827 81 -821
rect 85 -827 88 -821
rect 92 -827 95 -821
rect 99 -827 102 -821
rect 106 -827 109 -821
rect 113 -827 119 -821
rect 120 -827 126 -821
rect 127 -827 133 -821
rect 134 -827 140 -821
rect 141 -827 144 -821
rect 148 -827 151 -821
rect 155 -827 158 -821
rect 162 -827 168 -821
rect 169 -827 175 -821
rect 176 -827 179 -821
rect 183 -827 186 -821
rect 190 -827 193 -821
rect 197 -827 200 -821
rect 204 -827 207 -821
rect 211 -827 214 -821
rect 218 -827 221 -821
rect 225 -827 228 -821
rect 232 -827 235 -821
rect 239 -827 242 -821
rect 246 -827 249 -821
rect 253 -827 256 -821
rect 260 -827 266 -821
rect 267 -827 270 -821
rect 274 -827 277 -821
rect 281 -827 284 -821
rect 288 -827 291 -821
rect 295 -827 298 -821
rect 302 -827 305 -821
rect 309 -827 312 -821
rect 316 -827 319 -821
rect 323 -827 326 -821
rect 330 -827 333 -821
rect 337 -827 340 -821
rect 344 -827 347 -821
rect 351 -827 357 -821
rect 358 -827 364 -821
rect 365 -827 368 -821
rect 372 -827 375 -821
rect 379 -827 385 -821
rect 386 -827 389 -821
rect 393 -827 396 -821
rect 400 -827 403 -821
rect 407 -827 410 -821
rect 414 -827 417 -821
rect 421 -827 427 -821
rect 428 -827 431 -821
rect 435 -827 438 -821
rect 442 -827 445 -821
rect 449 -827 452 -821
rect 456 -827 459 -821
rect 463 -827 466 -821
rect 470 -827 473 -821
rect 477 -827 483 -821
rect 484 -827 487 -821
rect 491 -827 497 -821
rect 498 -827 504 -821
rect 505 -827 508 -821
rect 512 -827 515 -821
rect 519 -827 525 -821
rect 526 -827 529 -821
rect 533 -827 536 -821
rect 540 -827 543 -821
rect 547 -827 550 -821
rect 554 -827 560 -821
rect 561 -827 567 -821
rect 568 -827 574 -821
rect 575 -827 578 -821
rect 582 -827 585 -821
rect 589 -827 592 -821
rect 596 -827 599 -821
rect 603 -827 606 -821
rect 610 -827 613 -821
rect 617 -827 623 -821
rect 624 -827 630 -821
rect 631 -827 634 -821
rect 638 -827 644 -821
rect 645 -827 648 -821
rect 652 -827 658 -821
rect 659 -827 665 -821
rect 666 -827 669 -821
rect 673 -827 676 -821
rect 680 -827 683 -821
rect 687 -827 690 -821
rect 694 -827 700 -821
rect 701 -827 704 -821
rect 708 -827 711 -821
rect 715 -827 718 -821
rect 722 -827 728 -821
rect 729 -827 732 -821
rect 736 -827 739 -821
rect 743 -827 746 -821
rect 750 -827 753 -821
rect 757 -827 760 -821
rect 764 -827 767 -821
rect 771 -827 774 -821
rect 778 -827 784 -821
rect 785 -827 788 -821
rect 792 -827 795 -821
rect 799 -827 802 -821
rect 806 -827 809 -821
rect 813 -827 819 -821
rect 820 -827 823 -821
rect 827 -827 830 -821
rect 834 -827 837 -821
rect 841 -827 844 -821
rect 848 -827 854 -821
rect 855 -827 858 -821
rect 862 -827 865 -821
rect 869 -827 872 -821
rect 876 -827 879 -821
rect 883 -827 886 -821
rect 890 -827 893 -821
rect 897 -827 900 -821
rect 904 -827 907 -821
rect 911 -827 914 -821
rect 918 -827 921 -821
rect 925 -827 928 -821
rect 932 -827 935 -821
rect 939 -827 942 -821
rect 946 -827 949 -821
rect 953 -827 956 -821
rect 960 -827 963 -821
rect 967 -827 970 -821
rect 974 -827 977 -821
rect 981 -827 984 -821
rect 988 -827 991 -821
rect 995 -827 998 -821
rect 1002 -827 1005 -821
rect 1009 -827 1012 -821
rect 1016 -827 1019 -821
rect 1023 -827 1026 -821
rect 1030 -827 1033 -821
rect 1037 -827 1040 -821
rect 1044 -827 1047 -821
rect 1051 -827 1054 -821
rect 1058 -827 1061 -821
rect 1065 -827 1068 -821
rect 1072 -827 1075 -821
rect 1079 -827 1082 -821
rect 1086 -827 1089 -821
rect 1093 -827 1096 -821
rect 1100 -827 1103 -821
rect 1107 -827 1110 -821
rect 1114 -827 1117 -821
rect 1121 -827 1124 -821
rect 1128 -827 1131 -821
rect 1135 -827 1138 -821
rect 1142 -827 1145 -821
rect 1149 -827 1152 -821
rect 1156 -827 1159 -821
rect 1163 -827 1166 -821
rect 1170 -827 1173 -821
rect 1177 -827 1180 -821
rect 1184 -827 1187 -821
rect 1191 -827 1194 -821
rect 1198 -827 1201 -821
rect 1205 -827 1208 -821
rect 1212 -827 1215 -821
rect 1219 -827 1222 -821
rect 1 -914 7 -908
rect 8 -914 11 -908
rect 15 -914 21 -908
rect 22 -914 25 -908
rect 29 -914 35 -908
rect 36 -914 42 -908
rect 43 -914 46 -908
rect 50 -914 53 -908
rect 57 -914 60 -908
rect 64 -914 67 -908
rect 71 -914 77 -908
rect 78 -914 81 -908
rect 85 -914 88 -908
rect 92 -914 95 -908
rect 99 -914 102 -908
rect 106 -914 109 -908
rect 113 -914 119 -908
rect 120 -914 123 -908
rect 127 -914 133 -908
rect 134 -914 137 -908
rect 141 -914 144 -908
rect 148 -914 154 -908
rect 155 -914 158 -908
rect 162 -914 165 -908
rect 169 -914 172 -908
rect 176 -914 179 -908
rect 183 -914 186 -908
rect 190 -914 193 -908
rect 197 -914 200 -908
rect 204 -914 210 -908
rect 211 -914 214 -908
rect 218 -914 221 -908
rect 225 -914 228 -908
rect 232 -914 235 -908
rect 239 -914 242 -908
rect 246 -914 249 -908
rect 253 -914 256 -908
rect 260 -914 266 -908
rect 267 -914 270 -908
rect 274 -914 280 -908
rect 281 -914 284 -908
rect 288 -914 294 -908
rect 295 -914 298 -908
rect 302 -914 305 -908
rect 309 -914 315 -908
rect 316 -914 319 -908
rect 323 -914 326 -908
rect 330 -914 333 -908
rect 337 -914 340 -908
rect 344 -914 350 -908
rect 351 -914 354 -908
rect 358 -914 361 -908
rect 365 -914 368 -908
rect 372 -914 378 -908
rect 379 -914 382 -908
rect 386 -914 389 -908
rect 393 -914 396 -908
rect 400 -914 403 -908
rect 407 -914 410 -908
rect 414 -914 417 -908
rect 421 -914 427 -908
rect 428 -914 431 -908
rect 435 -914 441 -908
rect 442 -914 445 -908
rect 449 -914 452 -908
rect 456 -914 459 -908
rect 463 -914 466 -908
rect 470 -914 473 -908
rect 477 -914 483 -908
rect 484 -914 487 -908
rect 491 -914 494 -908
rect 498 -914 501 -908
rect 505 -914 508 -908
rect 512 -914 515 -908
rect 519 -914 522 -908
rect 526 -914 529 -908
rect 533 -914 536 -908
rect 540 -914 546 -908
rect 547 -914 550 -908
rect 554 -914 560 -908
rect 561 -914 564 -908
rect 568 -914 571 -908
rect 575 -914 578 -908
rect 582 -914 585 -908
rect 589 -914 592 -908
rect 596 -914 602 -908
rect 603 -914 606 -908
rect 610 -914 616 -908
rect 617 -914 623 -908
rect 624 -914 627 -908
rect 631 -914 634 -908
rect 638 -914 641 -908
rect 645 -914 648 -908
rect 652 -914 658 -908
rect 659 -914 662 -908
rect 666 -914 672 -908
rect 673 -914 679 -908
rect 680 -914 686 -908
rect 687 -914 690 -908
rect 694 -914 697 -908
rect 701 -914 704 -908
rect 708 -914 711 -908
rect 715 -914 718 -908
rect 722 -914 725 -908
rect 729 -914 732 -908
rect 736 -914 739 -908
rect 743 -914 746 -908
rect 750 -914 753 -908
rect 757 -914 760 -908
rect 764 -914 767 -908
rect 771 -914 774 -908
rect 778 -914 781 -908
rect 785 -914 788 -908
rect 792 -914 795 -908
rect 799 -914 802 -908
rect 806 -914 809 -908
rect 813 -914 816 -908
rect 820 -914 826 -908
rect 827 -914 830 -908
rect 834 -914 837 -908
rect 841 -914 844 -908
rect 848 -914 851 -908
rect 855 -914 858 -908
rect 862 -914 865 -908
rect 869 -914 872 -908
rect 876 -914 879 -908
rect 883 -914 886 -908
rect 890 -914 893 -908
rect 897 -914 903 -908
rect 904 -914 907 -908
rect 911 -914 914 -908
rect 918 -914 921 -908
rect 925 -914 928 -908
rect 932 -914 935 -908
rect 939 -914 942 -908
rect 946 -914 949 -908
rect 953 -914 956 -908
rect 960 -914 963 -908
rect 967 -914 970 -908
rect 974 -914 977 -908
rect 981 -914 984 -908
rect 988 -914 991 -908
rect 995 -914 998 -908
rect 1002 -914 1005 -908
rect 1009 -914 1012 -908
rect 1016 -914 1019 -908
rect 1023 -914 1026 -908
rect 1030 -914 1033 -908
rect 1037 -914 1040 -908
rect 1044 -914 1047 -908
rect 1051 -914 1054 -908
rect 1058 -914 1061 -908
rect 1065 -914 1068 -908
rect 1072 -914 1075 -908
rect 1079 -914 1082 -908
rect 1086 -914 1092 -908
rect 1093 -914 1096 -908
rect 1100 -914 1103 -908
rect 1107 -914 1110 -908
rect 1114 -914 1117 -908
rect 1121 -914 1124 -908
rect 1128 -914 1131 -908
rect 1163 -914 1166 -908
rect 1170 -914 1173 -908
rect 1177 -914 1180 -908
rect 1191 -914 1194 -908
rect 1 -1003 4 -997
rect 8 -1003 11 -997
rect 15 -1003 21 -997
rect 22 -1003 25 -997
rect 29 -1003 32 -997
rect 36 -1003 42 -997
rect 43 -1003 46 -997
rect 50 -1003 53 -997
rect 57 -1003 63 -997
rect 64 -1003 70 -997
rect 71 -1003 74 -997
rect 78 -1003 81 -997
rect 85 -1003 88 -997
rect 92 -1003 98 -997
rect 99 -1003 105 -997
rect 106 -1003 109 -997
rect 113 -1003 116 -997
rect 120 -1003 126 -997
rect 127 -1003 130 -997
rect 134 -1003 137 -997
rect 141 -1003 144 -997
rect 148 -1003 151 -997
rect 155 -1003 158 -997
rect 162 -1003 165 -997
rect 169 -1003 172 -997
rect 176 -1003 179 -997
rect 183 -1003 189 -997
rect 190 -1003 193 -997
rect 197 -1003 203 -997
rect 204 -1003 207 -997
rect 211 -1003 214 -997
rect 218 -1003 221 -997
rect 225 -1003 228 -997
rect 232 -1003 235 -997
rect 239 -1003 242 -997
rect 246 -1003 249 -997
rect 253 -1003 256 -997
rect 260 -1003 263 -997
rect 267 -1003 270 -997
rect 274 -1003 277 -997
rect 281 -1003 284 -997
rect 288 -1003 291 -997
rect 295 -1003 298 -997
rect 302 -1003 305 -997
rect 309 -1003 312 -997
rect 316 -1003 319 -997
rect 323 -1003 326 -997
rect 330 -1003 333 -997
rect 337 -1003 340 -997
rect 344 -1003 347 -997
rect 351 -1003 354 -997
rect 358 -1003 364 -997
rect 365 -1003 368 -997
rect 372 -1003 378 -997
rect 379 -1003 382 -997
rect 386 -1003 392 -997
rect 393 -1003 396 -997
rect 400 -1003 403 -997
rect 407 -1003 410 -997
rect 414 -1003 417 -997
rect 421 -1003 424 -997
rect 428 -1003 431 -997
rect 435 -1003 441 -997
rect 442 -1003 445 -997
rect 449 -1003 452 -997
rect 456 -1003 459 -997
rect 463 -1003 469 -997
rect 470 -1003 473 -997
rect 477 -1003 480 -997
rect 484 -1003 487 -997
rect 491 -1003 494 -997
rect 498 -1003 504 -997
rect 505 -1003 511 -997
rect 512 -1003 515 -997
rect 519 -1003 522 -997
rect 526 -1003 529 -997
rect 533 -1003 536 -997
rect 540 -1003 546 -997
rect 547 -1003 550 -997
rect 554 -1003 557 -997
rect 561 -1003 564 -997
rect 568 -1003 571 -997
rect 575 -1003 578 -997
rect 582 -1003 585 -997
rect 589 -1003 592 -997
rect 596 -1003 599 -997
rect 603 -1003 609 -997
rect 610 -1003 613 -997
rect 617 -1003 620 -997
rect 624 -1003 630 -997
rect 631 -1003 634 -997
rect 638 -1003 644 -997
rect 645 -1003 651 -997
rect 652 -1003 655 -997
rect 659 -1003 662 -997
rect 666 -1003 669 -997
rect 673 -1003 676 -997
rect 680 -1003 686 -997
rect 687 -1003 690 -997
rect 694 -1003 700 -997
rect 701 -1003 704 -997
rect 708 -1003 714 -997
rect 715 -1003 718 -997
rect 722 -1003 725 -997
rect 729 -1003 735 -997
rect 736 -1003 739 -997
rect 743 -1003 746 -997
rect 750 -1003 753 -997
rect 757 -1003 760 -997
rect 764 -1003 767 -997
rect 771 -1003 774 -997
rect 778 -1003 781 -997
rect 785 -1003 788 -997
rect 792 -1003 795 -997
rect 799 -1003 802 -997
rect 806 -1003 809 -997
rect 813 -1003 816 -997
rect 820 -1003 823 -997
rect 827 -1003 830 -997
rect 834 -1003 837 -997
rect 841 -1003 844 -997
rect 848 -1003 851 -997
rect 855 -1003 861 -997
rect 862 -1003 865 -997
rect 869 -1003 872 -997
rect 876 -1003 879 -997
rect 883 -1003 886 -997
rect 890 -1003 893 -997
rect 897 -1003 900 -997
rect 904 -1003 907 -997
rect 911 -1003 914 -997
rect 918 -1003 921 -997
rect 925 -1003 928 -997
rect 932 -1003 935 -997
rect 939 -1003 942 -997
rect 946 -1003 949 -997
rect 953 -1003 956 -997
rect 960 -1003 963 -997
rect 967 -1003 970 -997
rect 974 -1003 977 -997
rect 981 -1003 984 -997
rect 988 -1003 991 -997
rect 995 -1003 998 -997
rect 1002 -1003 1005 -997
rect 1009 -1003 1012 -997
rect 1016 -1003 1019 -997
rect 1023 -1003 1026 -997
rect 1030 -1003 1033 -997
rect 1037 -1003 1040 -997
rect 1044 -1003 1047 -997
rect 1051 -1003 1054 -997
rect 1058 -1003 1061 -997
rect 1065 -1003 1068 -997
rect 1072 -1003 1075 -997
rect 1079 -1003 1082 -997
rect 1086 -1003 1089 -997
rect 1093 -1003 1096 -997
rect 1100 -1003 1103 -997
rect 1107 -1003 1110 -997
rect 1114 -1003 1117 -997
rect 1121 -1003 1124 -997
rect 1128 -1003 1134 -997
rect 1135 -1003 1141 -997
rect 1142 -1003 1145 -997
rect 1149 -1003 1152 -997
rect 1156 -1003 1159 -997
rect 1163 -1003 1169 -997
rect 1170 -1003 1173 -997
rect 1184 -1003 1187 -997
rect 1191 -1003 1197 -997
rect 15 -1078 18 -1072
rect 22 -1078 25 -1072
rect 29 -1078 32 -1072
rect 36 -1078 39 -1072
rect 43 -1078 46 -1072
rect 50 -1078 53 -1072
rect 57 -1078 63 -1072
rect 64 -1078 70 -1072
rect 71 -1078 74 -1072
rect 78 -1078 81 -1072
rect 85 -1078 91 -1072
rect 92 -1078 98 -1072
rect 99 -1078 102 -1072
rect 106 -1078 109 -1072
rect 113 -1078 119 -1072
rect 120 -1078 123 -1072
rect 127 -1078 130 -1072
rect 134 -1078 137 -1072
rect 141 -1078 144 -1072
rect 148 -1078 154 -1072
rect 155 -1078 158 -1072
rect 162 -1078 165 -1072
rect 169 -1078 175 -1072
rect 176 -1078 179 -1072
rect 183 -1078 186 -1072
rect 190 -1078 193 -1072
rect 197 -1078 200 -1072
rect 204 -1078 210 -1072
rect 211 -1078 214 -1072
rect 218 -1078 221 -1072
rect 225 -1078 228 -1072
rect 232 -1078 235 -1072
rect 239 -1078 242 -1072
rect 246 -1078 249 -1072
rect 253 -1078 256 -1072
rect 260 -1078 266 -1072
rect 267 -1078 270 -1072
rect 274 -1078 277 -1072
rect 281 -1078 284 -1072
rect 288 -1078 291 -1072
rect 295 -1078 301 -1072
rect 302 -1078 305 -1072
rect 309 -1078 312 -1072
rect 316 -1078 322 -1072
rect 323 -1078 326 -1072
rect 330 -1078 333 -1072
rect 337 -1078 340 -1072
rect 344 -1078 347 -1072
rect 351 -1078 357 -1072
rect 358 -1078 361 -1072
rect 365 -1078 368 -1072
rect 372 -1078 375 -1072
rect 379 -1078 382 -1072
rect 386 -1078 389 -1072
rect 393 -1078 396 -1072
rect 400 -1078 403 -1072
rect 407 -1078 410 -1072
rect 414 -1078 417 -1072
rect 421 -1078 424 -1072
rect 428 -1078 431 -1072
rect 435 -1078 441 -1072
rect 442 -1078 445 -1072
rect 449 -1078 452 -1072
rect 456 -1078 459 -1072
rect 463 -1078 469 -1072
rect 470 -1078 473 -1072
rect 477 -1078 480 -1072
rect 484 -1078 487 -1072
rect 491 -1078 494 -1072
rect 498 -1078 501 -1072
rect 505 -1078 511 -1072
rect 512 -1078 515 -1072
rect 519 -1078 522 -1072
rect 526 -1078 529 -1072
rect 533 -1078 539 -1072
rect 540 -1078 543 -1072
rect 547 -1078 550 -1072
rect 554 -1078 557 -1072
rect 561 -1078 564 -1072
rect 568 -1078 574 -1072
rect 575 -1078 578 -1072
rect 582 -1078 585 -1072
rect 589 -1078 592 -1072
rect 596 -1078 602 -1072
rect 603 -1078 606 -1072
rect 610 -1078 613 -1072
rect 617 -1078 623 -1072
rect 624 -1078 627 -1072
rect 631 -1078 637 -1072
rect 638 -1078 641 -1072
rect 645 -1078 648 -1072
rect 652 -1078 655 -1072
rect 659 -1078 662 -1072
rect 666 -1078 669 -1072
rect 673 -1078 676 -1072
rect 680 -1078 683 -1072
rect 687 -1078 693 -1072
rect 694 -1078 697 -1072
rect 701 -1078 704 -1072
rect 708 -1078 711 -1072
rect 715 -1078 718 -1072
rect 722 -1078 725 -1072
rect 729 -1078 735 -1072
rect 736 -1078 739 -1072
rect 743 -1078 746 -1072
rect 750 -1078 753 -1072
rect 757 -1078 763 -1072
rect 764 -1078 767 -1072
rect 771 -1078 774 -1072
rect 778 -1078 781 -1072
rect 785 -1078 788 -1072
rect 792 -1078 795 -1072
rect 799 -1078 802 -1072
rect 806 -1078 812 -1072
rect 813 -1078 816 -1072
rect 820 -1078 823 -1072
rect 827 -1078 830 -1072
rect 834 -1078 837 -1072
rect 841 -1078 844 -1072
rect 848 -1078 851 -1072
rect 855 -1078 858 -1072
rect 862 -1078 865 -1072
rect 869 -1078 872 -1072
rect 876 -1078 879 -1072
rect 883 -1078 886 -1072
rect 890 -1078 893 -1072
rect 897 -1078 900 -1072
rect 904 -1078 907 -1072
rect 911 -1078 914 -1072
rect 918 -1078 924 -1072
rect 925 -1078 928 -1072
rect 932 -1078 935 -1072
rect 939 -1078 942 -1072
rect 946 -1078 949 -1072
rect 953 -1078 959 -1072
rect 960 -1078 963 -1072
rect 967 -1078 970 -1072
rect 974 -1078 977 -1072
rect 981 -1078 984 -1072
rect 988 -1078 991 -1072
rect 995 -1078 998 -1072
rect 1002 -1078 1005 -1072
rect 1009 -1078 1012 -1072
rect 1016 -1078 1019 -1072
rect 1023 -1078 1026 -1072
rect 1030 -1078 1036 -1072
rect 1037 -1078 1043 -1072
rect 1044 -1078 1047 -1072
rect 1051 -1078 1054 -1072
rect 1058 -1078 1064 -1072
rect 1065 -1078 1071 -1072
rect 1072 -1078 1075 -1072
rect 1079 -1078 1082 -1072
rect 1086 -1078 1089 -1072
rect 1093 -1078 1096 -1072
rect 1121 -1078 1124 -1072
rect 1184 -1078 1187 -1072
rect 22 -1161 28 -1155
rect 29 -1161 32 -1155
rect 36 -1161 39 -1155
rect 43 -1161 46 -1155
rect 50 -1161 53 -1155
rect 57 -1161 60 -1155
rect 64 -1161 67 -1155
rect 71 -1161 74 -1155
rect 78 -1161 84 -1155
rect 85 -1161 91 -1155
rect 92 -1161 95 -1155
rect 99 -1161 102 -1155
rect 106 -1161 109 -1155
rect 113 -1161 119 -1155
rect 120 -1161 123 -1155
rect 127 -1161 133 -1155
rect 134 -1161 140 -1155
rect 141 -1161 144 -1155
rect 148 -1161 151 -1155
rect 155 -1161 161 -1155
rect 162 -1161 168 -1155
rect 169 -1161 172 -1155
rect 176 -1161 179 -1155
rect 183 -1161 189 -1155
rect 190 -1161 193 -1155
rect 197 -1161 203 -1155
rect 204 -1161 207 -1155
rect 211 -1161 214 -1155
rect 218 -1161 221 -1155
rect 225 -1161 231 -1155
rect 232 -1161 235 -1155
rect 239 -1161 242 -1155
rect 246 -1161 249 -1155
rect 253 -1161 256 -1155
rect 260 -1161 263 -1155
rect 267 -1161 270 -1155
rect 274 -1161 277 -1155
rect 281 -1161 287 -1155
rect 288 -1161 291 -1155
rect 295 -1161 298 -1155
rect 302 -1161 308 -1155
rect 309 -1161 312 -1155
rect 316 -1161 319 -1155
rect 323 -1161 326 -1155
rect 330 -1161 336 -1155
rect 337 -1161 340 -1155
rect 344 -1161 347 -1155
rect 351 -1161 354 -1155
rect 358 -1161 361 -1155
rect 365 -1161 368 -1155
rect 372 -1161 375 -1155
rect 379 -1161 382 -1155
rect 386 -1161 389 -1155
rect 393 -1161 396 -1155
rect 400 -1161 403 -1155
rect 407 -1161 410 -1155
rect 414 -1161 420 -1155
rect 421 -1161 424 -1155
rect 428 -1161 431 -1155
rect 435 -1161 438 -1155
rect 442 -1161 448 -1155
rect 449 -1161 452 -1155
rect 456 -1161 459 -1155
rect 463 -1161 466 -1155
rect 470 -1161 473 -1155
rect 477 -1161 480 -1155
rect 484 -1161 487 -1155
rect 491 -1161 494 -1155
rect 498 -1161 501 -1155
rect 505 -1161 511 -1155
rect 512 -1161 515 -1155
rect 519 -1161 522 -1155
rect 526 -1161 529 -1155
rect 533 -1161 536 -1155
rect 540 -1161 543 -1155
rect 547 -1161 553 -1155
rect 554 -1161 557 -1155
rect 561 -1161 564 -1155
rect 568 -1161 571 -1155
rect 575 -1161 578 -1155
rect 582 -1161 588 -1155
rect 589 -1161 592 -1155
rect 596 -1161 599 -1155
rect 603 -1161 609 -1155
rect 610 -1161 613 -1155
rect 617 -1161 620 -1155
rect 624 -1161 630 -1155
rect 631 -1161 634 -1155
rect 638 -1161 641 -1155
rect 645 -1161 648 -1155
rect 652 -1161 658 -1155
rect 659 -1161 662 -1155
rect 666 -1161 672 -1155
rect 673 -1161 676 -1155
rect 680 -1161 683 -1155
rect 687 -1161 690 -1155
rect 694 -1161 697 -1155
rect 701 -1161 704 -1155
rect 708 -1161 711 -1155
rect 715 -1161 718 -1155
rect 722 -1161 725 -1155
rect 729 -1161 732 -1155
rect 736 -1161 739 -1155
rect 743 -1161 746 -1155
rect 750 -1161 753 -1155
rect 757 -1161 760 -1155
rect 764 -1161 767 -1155
rect 771 -1161 774 -1155
rect 778 -1161 781 -1155
rect 785 -1161 788 -1155
rect 792 -1161 795 -1155
rect 799 -1161 802 -1155
rect 806 -1161 812 -1155
rect 813 -1161 816 -1155
rect 820 -1161 823 -1155
rect 827 -1161 830 -1155
rect 834 -1161 837 -1155
rect 841 -1161 844 -1155
rect 848 -1161 854 -1155
rect 855 -1161 858 -1155
rect 862 -1161 865 -1155
rect 869 -1161 872 -1155
rect 876 -1161 879 -1155
rect 883 -1161 886 -1155
rect 890 -1161 893 -1155
rect 897 -1161 900 -1155
rect 904 -1161 907 -1155
rect 911 -1161 914 -1155
rect 918 -1161 921 -1155
rect 925 -1161 928 -1155
rect 932 -1161 938 -1155
rect 939 -1161 942 -1155
rect 946 -1161 949 -1155
rect 953 -1161 956 -1155
rect 960 -1161 963 -1155
rect 967 -1161 970 -1155
rect 974 -1161 980 -1155
rect 981 -1161 984 -1155
rect 988 -1161 991 -1155
rect 995 -1161 998 -1155
rect 1002 -1161 1008 -1155
rect 1009 -1161 1012 -1155
rect 1016 -1161 1019 -1155
rect 1023 -1161 1026 -1155
rect 1030 -1161 1033 -1155
rect 1037 -1161 1040 -1155
rect 1044 -1161 1050 -1155
rect 1058 -1161 1061 -1155
rect 1065 -1161 1068 -1155
rect 1079 -1161 1082 -1155
rect 1086 -1161 1089 -1155
rect 1107 -1161 1110 -1155
rect 1184 -1161 1190 -1155
rect 1 -1236 7 -1230
rect 8 -1236 14 -1230
rect 15 -1236 18 -1230
rect 22 -1236 28 -1230
rect 29 -1236 32 -1230
rect 36 -1236 39 -1230
rect 43 -1236 49 -1230
rect 50 -1236 53 -1230
rect 57 -1236 63 -1230
rect 64 -1236 70 -1230
rect 71 -1236 74 -1230
rect 78 -1236 81 -1230
rect 85 -1236 91 -1230
rect 92 -1236 95 -1230
rect 99 -1236 102 -1230
rect 106 -1236 109 -1230
rect 113 -1236 119 -1230
rect 120 -1236 123 -1230
rect 127 -1236 130 -1230
rect 134 -1236 137 -1230
rect 141 -1236 144 -1230
rect 148 -1236 154 -1230
rect 155 -1236 158 -1230
rect 162 -1236 165 -1230
rect 169 -1236 172 -1230
rect 176 -1236 182 -1230
rect 183 -1236 186 -1230
rect 190 -1236 193 -1230
rect 197 -1236 200 -1230
rect 204 -1236 207 -1230
rect 211 -1236 214 -1230
rect 218 -1236 221 -1230
rect 225 -1236 228 -1230
rect 232 -1236 235 -1230
rect 239 -1236 242 -1230
rect 246 -1236 249 -1230
rect 253 -1236 256 -1230
rect 260 -1236 266 -1230
rect 267 -1236 270 -1230
rect 274 -1236 277 -1230
rect 281 -1236 284 -1230
rect 288 -1236 291 -1230
rect 295 -1236 298 -1230
rect 302 -1236 305 -1230
rect 309 -1236 312 -1230
rect 316 -1236 322 -1230
rect 323 -1236 326 -1230
rect 330 -1236 333 -1230
rect 337 -1236 340 -1230
rect 344 -1236 347 -1230
rect 351 -1236 354 -1230
rect 358 -1236 361 -1230
rect 365 -1236 368 -1230
rect 372 -1236 378 -1230
rect 379 -1236 385 -1230
rect 386 -1236 392 -1230
rect 393 -1236 396 -1230
rect 400 -1236 403 -1230
rect 407 -1236 410 -1230
rect 414 -1236 417 -1230
rect 421 -1236 427 -1230
rect 428 -1236 431 -1230
rect 435 -1236 438 -1230
rect 442 -1236 448 -1230
rect 449 -1236 452 -1230
rect 456 -1236 459 -1230
rect 463 -1236 466 -1230
rect 470 -1236 473 -1230
rect 477 -1236 480 -1230
rect 484 -1236 487 -1230
rect 491 -1236 494 -1230
rect 498 -1236 501 -1230
rect 505 -1236 511 -1230
rect 512 -1236 515 -1230
rect 519 -1236 522 -1230
rect 526 -1236 529 -1230
rect 533 -1236 536 -1230
rect 540 -1236 546 -1230
rect 547 -1236 553 -1230
rect 554 -1236 557 -1230
rect 561 -1236 567 -1230
rect 568 -1236 574 -1230
rect 575 -1236 578 -1230
rect 582 -1236 585 -1230
rect 589 -1236 595 -1230
rect 596 -1236 599 -1230
rect 603 -1236 606 -1230
rect 610 -1236 613 -1230
rect 617 -1236 620 -1230
rect 624 -1236 627 -1230
rect 631 -1236 634 -1230
rect 638 -1236 644 -1230
rect 645 -1236 648 -1230
rect 652 -1236 658 -1230
rect 659 -1236 665 -1230
rect 666 -1236 669 -1230
rect 673 -1236 676 -1230
rect 680 -1236 683 -1230
rect 687 -1236 690 -1230
rect 694 -1236 697 -1230
rect 701 -1236 704 -1230
rect 708 -1236 714 -1230
rect 715 -1236 718 -1230
rect 722 -1236 728 -1230
rect 729 -1236 732 -1230
rect 736 -1236 739 -1230
rect 743 -1236 746 -1230
rect 750 -1236 753 -1230
rect 757 -1236 760 -1230
rect 764 -1236 767 -1230
rect 771 -1236 777 -1230
rect 778 -1236 781 -1230
rect 785 -1236 788 -1230
rect 792 -1236 795 -1230
rect 799 -1236 802 -1230
rect 806 -1236 809 -1230
rect 813 -1236 816 -1230
rect 820 -1236 823 -1230
rect 827 -1236 833 -1230
rect 834 -1236 837 -1230
rect 841 -1236 844 -1230
rect 848 -1236 851 -1230
rect 855 -1236 858 -1230
rect 862 -1236 865 -1230
rect 869 -1236 872 -1230
rect 876 -1236 879 -1230
rect 883 -1236 886 -1230
rect 890 -1236 893 -1230
rect 897 -1236 900 -1230
rect 904 -1236 907 -1230
rect 911 -1236 914 -1230
rect 918 -1236 921 -1230
rect 925 -1236 928 -1230
rect 932 -1236 935 -1230
rect 939 -1236 942 -1230
rect 946 -1236 949 -1230
rect 953 -1236 956 -1230
rect 960 -1236 963 -1230
rect 967 -1236 970 -1230
rect 974 -1236 977 -1230
rect 981 -1236 984 -1230
rect 988 -1236 991 -1230
rect 995 -1236 998 -1230
rect 1002 -1236 1005 -1230
rect 1009 -1236 1012 -1230
rect 1016 -1236 1019 -1230
rect 1023 -1236 1026 -1230
rect 1030 -1236 1033 -1230
rect 1037 -1236 1040 -1230
rect 1044 -1236 1047 -1230
rect 1051 -1236 1054 -1230
rect 1058 -1236 1061 -1230
rect 1065 -1236 1068 -1230
rect 1072 -1236 1075 -1230
rect 1079 -1236 1082 -1230
rect 1086 -1236 1089 -1230
rect 1093 -1236 1096 -1230
rect 1100 -1236 1103 -1230
rect 1107 -1236 1110 -1230
rect 1114 -1236 1117 -1230
rect 1121 -1236 1124 -1230
rect 1128 -1236 1131 -1230
rect 1 -1307 7 -1301
rect 8 -1307 14 -1301
rect 15 -1307 21 -1301
rect 43 -1307 46 -1301
rect 71 -1307 74 -1301
rect 78 -1307 81 -1301
rect 85 -1307 88 -1301
rect 92 -1307 98 -1301
rect 99 -1307 102 -1301
rect 106 -1307 109 -1301
rect 113 -1307 116 -1301
rect 120 -1307 123 -1301
rect 127 -1307 130 -1301
rect 134 -1307 137 -1301
rect 141 -1307 144 -1301
rect 148 -1307 154 -1301
rect 155 -1307 158 -1301
rect 162 -1307 165 -1301
rect 169 -1307 172 -1301
rect 176 -1307 179 -1301
rect 183 -1307 186 -1301
rect 190 -1307 196 -1301
rect 197 -1307 200 -1301
rect 204 -1307 207 -1301
rect 211 -1307 214 -1301
rect 218 -1307 221 -1301
rect 225 -1307 228 -1301
rect 232 -1307 235 -1301
rect 239 -1307 245 -1301
rect 246 -1307 249 -1301
rect 253 -1307 256 -1301
rect 260 -1307 263 -1301
rect 267 -1307 270 -1301
rect 274 -1307 277 -1301
rect 281 -1307 284 -1301
rect 288 -1307 291 -1301
rect 295 -1307 298 -1301
rect 302 -1307 308 -1301
rect 309 -1307 312 -1301
rect 316 -1307 319 -1301
rect 323 -1307 326 -1301
rect 330 -1307 333 -1301
rect 337 -1307 343 -1301
rect 344 -1307 347 -1301
rect 351 -1307 354 -1301
rect 358 -1307 361 -1301
rect 365 -1307 368 -1301
rect 372 -1307 375 -1301
rect 379 -1307 382 -1301
rect 386 -1307 389 -1301
rect 393 -1307 396 -1301
rect 400 -1307 406 -1301
rect 407 -1307 410 -1301
rect 414 -1307 417 -1301
rect 421 -1307 424 -1301
rect 428 -1307 431 -1301
rect 435 -1307 438 -1301
rect 442 -1307 445 -1301
rect 449 -1307 452 -1301
rect 456 -1307 459 -1301
rect 463 -1307 469 -1301
rect 470 -1307 473 -1301
rect 477 -1307 483 -1301
rect 484 -1307 487 -1301
rect 491 -1307 494 -1301
rect 498 -1307 504 -1301
rect 505 -1307 508 -1301
rect 512 -1307 515 -1301
rect 519 -1307 522 -1301
rect 526 -1307 529 -1301
rect 533 -1307 539 -1301
rect 540 -1307 543 -1301
rect 547 -1307 550 -1301
rect 554 -1307 557 -1301
rect 561 -1307 564 -1301
rect 568 -1307 574 -1301
rect 575 -1307 581 -1301
rect 582 -1307 585 -1301
rect 589 -1307 592 -1301
rect 596 -1307 602 -1301
rect 603 -1307 606 -1301
rect 610 -1307 616 -1301
rect 617 -1307 620 -1301
rect 624 -1307 627 -1301
rect 631 -1307 637 -1301
rect 638 -1307 641 -1301
rect 645 -1307 648 -1301
rect 652 -1307 658 -1301
rect 659 -1307 662 -1301
rect 666 -1307 669 -1301
rect 673 -1307 679 -1301
rect 680 -1307 683 -1301
rect 687 -1307 690 -1301
rect 694 -1307 697 -1301
rect 701 -1307 704 -1301
rect 708 -1307 711 -1301
rect 715 -1307 718 -1301
rect 722 -1307 725 -1301
rect 729 -1307 732 -1301
rect 736 -1307 739 -1301
rect 743 -1307 746 -1301
rect 750 -1307 753 -1301
rect 757 -1307 760 -1301
rect 764 -1307 767 -1301
rect 771 -1307 774 -1301
rect 778 -1307 781 -1301
rect 785 -1307 788 -1301
rect 792 -1307 798 -1301
rect 799 -1307 802 -1301
rect 806 -1307 809 -1301
rect 813 -1307 816 -1301
rect 820 -1307 823 -1301
rect 827 -1307 830 -1301
rect 834 -1307 837 -1301
rect 841 -1307 844 -1301
rect 848 -1307 851 -1301
rect 855 -1307 858 -1301
rect 862 -1307 868 -1301
rect 869 -1307 872 -1301
rect 876 -1307 879 -1301
rect 883 -1307 886 -1301
rect 890 -1307 893 -1301
rect 897 -1307 900 -1301
rect 904 -1307 907 -1301
rect 911 -1307 914 -1301
rect 918 -1307 924 -1301
rect 925 -1307 928 -1301
rect 932 -1307 935 -1301
rect 939 -1307 942 -1301
rect 946 -1307 949 -1301
rect 953 -1307 956 -1301
rect 960 -1307 963 -1301
rect 967 -1307 970 -1301
rect 974 -1307 980 -1301
rect 981 -1307 984 -1301
rect 988 -1307 991 -1301
rect 995 -1307 1001 -1301
rect 1002 -1307 1005 -1301
rect 1009 -1307 1012 -1301
rect 1016 -1307 1022 -1301
rect 1023 -1307 1029 -1301
rect 1030 -1307 1033 -1301
rect 1037 -1307 1040 -1301
rect 1044 -1307 1047 -1301
rect 1051 -1307 1054 -1301
rect 1058 -1307 1064 -1301
rect 1065 -1307 1068 -1301
rect 1079 -1307 1082 -1301
rect 1086 -1307 1089 -1301
rect 1093 -1307 1099 -1301
rect 1100 -1307 1103 -1301
rect 1 -1378 7 -1372
rect 8 -1378 14 -1372
rect 15 -1378 18 -1372
rect 22 -1378 25 -1372
rect 29 -1378 32 -1372
rect 36 -1378 39 -1372
rect 43 -1378 46 -1372
rect 50 -1378 53 -1372
rect 57 -1378 60 -1372
rect 64 -1378 70 -1372
rect 71 -1378 74 -1372
rect 78 -1378 81 -1372
rect 85 -1378 88 -1372
rect 92 -1378 98 -1372
rect 99 -1378 105 -1372
rect 106 -1378 109 -1372
rect 113 -1378 116 -1372
rect 120 -1378 123 -1372
rect 127 -1378 130 -1372
rect 134 -1378 140 -1372
rect 141 -1378 147 -1372
rect 148 -1378 151 -1372
rect 155 -1378 158 -1372
rect 162 -1378 165 -1372
rect 169 -1378 172 -1372
rect 176 -1378 182 -1372
rect 183 -1378 186 -1372
rect 190 -1378 193 -1372
rect 197 -1378 203 -1372
rect 204 -1378 207 -1372
rect 211 -1378 214 -1372
rect 218 -1378 221 -1372
rect 225 -1378 228 -1372
rect 232 -1378 238 -1372
rect 239 -1378 242 -1372
rect 246 -1378 252 -1372
rect 253 -1378 256 -1372
rect 260 -1378 263 -1372
rect 267 -1378 270 -1372
rect 274 -1378 280 -1372
rect 281 -1378 287 -1372
rect 288 -1378 291 -1372
rect 295 -1378 298 -1372
rect 302 -1378 305 -1372
rect 309 -1378 312 -1372
rect 316 -1378 319 -1372
rect 323 -1378 326 -1372
rect 330 -1378 333 -1372
rect 337 -1378 340 -1372
rect 344 -1378 350 -1372
rect 351 -1378 354 -1372
rect 358 -1378 361 -1372
rect 365 -1378 371 -1372
rect 372 -1378 375 -1372
rect 379 -1378 382 -1372
rect 386 -1378 389 -1372
rect 393 -1378 396 -1372
rect 400 -1378 403 -1372
rect 407 -1378 413 -1372
rect 414 -1378 417 -1372
rect 421 -1378 424 -1372
rect 428 -1378 431 -1372
rect 435 -1378 441 -1372
rect 442 -1378 445 -1372
rect 449 -1378 452 -1372
rect 456 -1378 459 -1372
rect 463 -1378 466 -1372
rect 470 -1378 473 -1372
rect 477 -1378 483 -1372
rect 484 -1378 487 -1372
rect 491 -1378 497 -1372
rect 498 -1378 501 -1372
rect 505 -1378 511 -1372
rect 512 -1378 515 -1372
rect 519 -1378 522 -1372
rect 526 -1378 529 -1372
rect 533 -1378 536 -1372
rect 540 -1378 546 -1372
rect 547 -1378 550 -1372
rect 554 -1378 557 -1372
rect 561 -1378 564 -1372
rect 568 -1378 574 -1372
rect 575 -1378 578 -1372
rect 582 -1378 585 -1372
rect 589 -1378 592 -1372
rect 596 -1378 599 -1372
rect 603 -1378 606 -1372
rect 610 -1378 613 -1372
rect 617 -1378 620 -1372
rect 624 -1378 630 -1372
rect 631 -1378 634 -1372
rect 638 -1378 641 -1372
rect 645 -1378 651 -1372
rect 652 -1378 658 -1372
rect 659 -1378 665 -1372
rect 666 -1378 669 -1372
rect 673 -1378 676 -1372
rect 680 -1378 683 -1372
rect 687 -1378 690 -1372
rect 694 -1378 697 -1372
rect 701 -1378 704 -1372
rect 708 -1378 711 -1372
rect 715 -1378 718 -1372
rect 722 -1378 728 -1372
rect 729 -1378 735 -1372
rect 736 -1378 739 -1372
rect 743 -1378 746 -1372
rect 750 -1378 753 -1372
rect 757 -1378 760 -1372
rect 764 -1378 767 -1372
rect 771 -1378 774 -1372
rect 778 -1378 781 -1372
rect 785 -1378 788 -1372
rect 792 -1378 795 -1372
rect 799 -1378 802 -1372
rect 806 -1378 809 -1372
rect 813 -1378 816 -1372
rect 820 -1378 823 -1372
rect 827 -1378 830 -1372
rect 834 -1378 837 -1372
rect 841 -1378 844 -1372
rect 848 -1378 851 -1372
rect 855 -1378 858 -1372
rect 862 -1378 865 -1372
rect 869 -1378 872 -1372
rect 876 -1378 879 -1372
rect 883 -1378 886 -1372
rect 890 -1378 893 -1372
rect 897 -1378 900 -1372
rect 904 -1378 907 -1372
rect 911 -1378 914 -1372
rect 918 -1378 921 -1372
rect 925 -1378 928 -1372
rect 932 -1378 935 -1372
rect 939 -1378 942 -1372
rect 946 -1378 949 -1372
rect 953 -1378 956 -1372
rect 960 -1378 963 -1372
rect 967 -1378 970 -1372
rect 974 -1378 977 -1372
rect 981 -1378 984 -1372
rect 988 -1378 991 -1372
rect 995 -1378 1001 -1372
rect 1002 -1378 1005 -1372
rect 1009 -1378 1012 -1372
rect 1016 -1378 1019 -1372
rect 1023 -1378 1029 -1372
rect 1030 -1378 1033 -1372
rect 1065 -1378 1068 -1372
rect 1 -1453 7 -1447
rect 8 -1453 11 -1447
rect 15 -1453 21 -1447
rect 22 -1453 25 -1447
rect 29 -1453 32 -1447
rect 36 -1453 42 -1447
rect 43 -1453 46 -1447
rect 50 -1453 53 -1447
rect 57 -1453 60 -1447
rect 64 -1453 70 -1447
rect 71 -1453 74 -1447
rect 78 -1453 81 -1447
rect 85 -1453 88 -1447
rect 92 -1453 95 -1447
rect 99 -1453 102 -1447
rect 106 -1453 109 -1447
rect 113 -1453 116 -1447
rect 120 -1453 123 -1447
rect 127 -1453 133 -1447
rect 134 -1453 140 -1447
rect 141 -1453 144 -1447
rect 148 -1453 151 -1447
rect 155 -1453 158 -1447
rect 162 -1453 165 -1447
rect 169 -1453 172 -1447
rect 176 -1453 179 -1447
rect 183 -1453 186 -1447
rect 190 -1453 196 -1447
rect 197 -1453 200 -1447
rect 204 -1453 210 -1447
rect 211 -1453 217 -1447
rect 218 -1453 221 -1447
rect 225 -1453 228 -1447
rect 232 -1453 235 -1447
rect 239 -1453 242 -1447
rect 246 -1453 249 -1447
rect 253 -1453 256 -1447
rect 260 -1453 263 -1447
rect 267 -1453 270 -1447
rect 274 -1453 280 -1447
rect 281 -1453 287 -1447
rect 288 -1453 291 -1447
rect 295 -1453 298 -1447
rect 302 -1453 305 -1447
rect 309 -1453 312 -1447
rect 316 -1453 322 -1447
rect 323 -1453 326 -1447
rect 330 -1453 333 -1447
rect 337 -1453 340 -1447
rect 344 -1453 347 -1447
rect 351 -1453 354 -1447
rect 358 -1453 361 -1447
rect 365 -1453 371 -1447
rect 372 -1453 378 -1447
rect 379 -1453 382 -1447
rect 386 -1453 389 -1447
rect 393 -1453 396 -1447
rect 400 -1453 403 -1447
rect 407 -1453 410 -1447
rect 414 -1453 417 -1447
rect 421 -1453 427 -1447
rect 428 -1453 431 -1447
rect 435 -1453 441 -1447
rect 442 -1453 445 -1447
rect 449 -1453 452 -1447
rect 456 -1453 462 -1447
rect 463 -1453 466 -1447
rect 470 -1453 476 -1447
rect 477 -1453 480 -1447
rect 484 -1453 490 -1447
rect 491 -1453 494 -1447
rect 498 -1453 501 -1447
rect 505 -1453 508 -1447
rect 512 -1453 515 -1447
rect 519 -1453 525 -1447
rect 526 -1453 532 -1447
rect 533 -1453 539 -1447
rect 540 -1453 543 -1447
rect 547 -1453 550 -1447
rect 554 -1453 557 -1447
rect 561 -1453 564 -1447
rect 568 -1453 571 -1447
rect 575 -1453 578 -1447
rect 582 -1453 585 -1447
rect 589 -1453 592 -1447
rect 596 -1453 599 -1447
rect 603 -1453 609 -1447
rect 610 -1453 613 -1447
rect 617 -1453 620 -1447
rect 624 -1453 627 -1447
rect 631 -1453 637 -1447
rect 638 -1453 644 -1447
rect 645 -1453 648 -1447
rect 652 -1453 655 -1447
rect 659 -1453 662 -1447
rect 666 -1453 669 -1447
rect 673 -1453 676 -1447
rect 680 -1453 683 -1447
rect 687 -1453 690 -1447
rect 694 -1453 697 -1447
rect 701 -1453 704 -1447
rect 708 -1453 711 -1447
rect 715 -1453 718 -1447
rect 722 -1453 725 -1447
rect 729 -1453 732 -1447
rect 736 -1453 739 -1447
rect 743 -1453 746 -1447
rect 750 -1453 753 -1447
rect 757 -1453 760 -1447
rect 764 -1453 770 -1447
rect 771 -1453 774 -1447
rect 778 -1453 781 -1447
rect 785 -1453 788 -1447
rect 792 -1453 798 -1447
rect 799 -1453 802 -1447
rect 806 -1453 809 -1447
rect 813 -1453 816 -1447
rect 820 -1453 826 -1447
rect 827 -1453 830 -1447
rect 834 -1453 837 -1447
rect 841 -1453 844 -1447
rect 848 -1453 851 -1447
rect 855 -1453 858 -1447
rect 862 -1453 865 -1447
rect 869 -1453 872 -1447
rect 876 -1453 879 -1447
rect 883 -1453 886 -1447
rect 890 -1453 893 -1447
rect 897 -1453 900 -1447
rect 904 -1453 907 -1447
rect 911 -1453 914 -1447
rect 918 -1453 921 -1447
rect 925 -1453 928 -1447
rect 932 -1453 935 -1447
rect 939 -1453 942 -1447
rect 946 -1453 949 -1447
rect 953 -1453 956 -1447
rect 960 -1453 963 -1447
rect 967 -1453 970 -1447
rect 974 -1453 977 -1447
rect 981 -1453 984 -1447
rect 988 -1453 991 -1447
rect 995 -1453 998 -1447
rect 1002 -1453 1005 -1447
rect 1009 -1453 1012 -1447
rect 1016 -1453 1019 -1447
rect 1023 -1453 1026 -1447
rect 1030 -1453 1033 -1447
rect 1037 -1453 1040 -1447
rect 1044 -1453 1050 -1447
rect 1051 -1453 1057 -1447
rect 1058 -1453 1061 -1447
rect 1065 -1453 1068 -1447
rect 1 -1536 4 -1530
rect 8 -1536 14 -1530
rect 15 -1536 18 -1530
rect 22 -1536 25 -1530
rect 29 -1536 32 -1530
rect 36 -1536 39 -1530
rect 43 -1536 46 -1530
rect 50 -1536 53 -1530
rect 57 -1536 60 -1530
rect 64 -1536 70 -1530
rect 71 -1536 74 -1530
rect 78 -1536 81 -1530
rect 85 -1536 88 -1530
rect 92 -1536 98 -1530
rect 99 -1536 102 -1530
rect 106 -1536 109 -1530
rect 113 -1536 119 -1530
rect 120 -1536 123 -1530
rect 127 -1536 130 -1530
rect 134 -1536 140 -1530
rect 141 -1536 144 -1530
rect 148 -1536 151 -1530
rect 155 -1536 158 -1530
rect 162 -1536 165 -1530
rect 169 -1536 172 -1530
rect 176 -1536 179 -1530
rect 183 -1536 186 -1530
rect 190 -1536 193 -1530
rect 197 -1536 203 -1530
rect 204 -1536 207 -1530
rect 211 -1536 214 -1530
rect 218 -1536 221 -1530
rect 225 -1536 228 -1530
rect 232 -1536 235 -1530
rect 239 -1536 242 -1530
rect 246 -1536 249 -1530
rect 253 -1536 256 -1530
rect 260 -1536 263 -1530
rect 267 -1536 270 -1530
rect 274 -1536 277 -1530
rect 281 -1536 284 -1530
rect 288 -1536 294 -1530
rect 295 -1536 301 -1530
rect 302 -1536 305 -1530
rect 309 -1536 312 -1530
rect 316 -1536 319 -1530
rect 323 -1536 326 -1530
rect 330 -1536 333 -1530
rect 337 -1536 340 -1530
rect 344 -1536 350 -1530
rect 351 -1536 357 -1530
rect 358 -1536 361 -1530
rect 365 -1536 368 -1530
rect 372 -1536 375 -1530
rect 379 -1536 382 -1530
rect 386 -1536 389 -1530
rect 393 -1536 396 -1530
rect 400 -1536 403 -1530
rect 407 -1536 413 -1530
rect 414 -1536 417 -1530
rect 421 -1536 424 -1530
rect 428 -1536 431 -1530
rect 435 -1536 438 -1530
rect 442 -1536 445 -1530
rect 449 -1536 452 -1530
rect 456 -1536 459 -1530
rect 463 -1536 469 -1530
rect 470 -1536 473 -1530
rect 477 -1536 480 -1530
rect 484 -1536 490 -1530
rect 491 -1536 494 -1530
rect 498 -1536 501 -1530
rect 505 -1536 511 -1530
rect 512 -1536 518 -1530
rect 519 -1536 525 -1530
rect 526 -1536 532 -1530
rect 533 -1536 539 -1530
rect 540 -1536 546 -1530
rect 547 -1536 550 -1530
rect 554 -1536 557 -1530
rect 561 -1536 567 -1530
rect 568 -1536 571 -1530
rect 575 -1536 578 -1530
rect 582 -1536 585 -1530
rect 589 -1536 595 -1530
rect 596 -1536 599 -1530
rect 603 -1536 609 -1530
rect 610 -1536 613 -1530
rect 617 -1536 623 -1530
rect 624 -1536 627 -1530
rect 631 -1536 634 -1530
rect 638 -1536 641 -1530
rect 645 -1536 648 -1530
rect 652 -1536 655 -1530
rect 659 -1536 665 -1530
rect 666 -1536 669 -1530
rect 673 -1536 676 -1530
rect 680 -1536 686 -1530
rect 687 -1536 690 -1530
rect 694 -1536 697 -1530
rect 701 -1536 704 -1530
rect 708 -1536 711 -1530
rect 715 -1536 718 -1530
rect 722 -1536 728 -1530
rect 729 -1536 732 -1530
rect 736 -1536 742 -1530
rect 743 -1536 746 -1530
rect 750 -1536 753 -1530
rect 757 -1536 760 -1530
rect 764 -1536 767 -1530
rect 771 -1536 774 -1530
rect 778 -1536 781 -1530
rect 785 -1536 788 -1530
rect 792 -1536 795 -1530
rect 799 -1536 802 -1530
rect 806 -1536 809 -1530
rect 813 -1536 816 -1530
rect 820 -1536 823 -1530
rect 827 -1536 830 -1530
rect 834 -1536 837 -1530
rect 841 -1536 847 -1530
rect 848 -1536 851 -1530
rect 855 -1536 858 -1530
rect 862 -1536 865 -1530
rect 869 -1536 872 -1530
rect 876 -1536 879 -1530
rect 883 -1536 886 -1530
rect 890 -1536 893 -1530
rect 897 -1536 900 -1530
rect 904 -1536 907 -1530
rect 911 -1536 914 -1530
rect 918 -1536 921 -1530
rect 925 -1536 928 -1530
rect 932 -1536 935 -1530
rect 939 -1536 942 -1530
rect 946 -1536 949 -1530
rect 953 -1536 956 -1530
rect 960 -1536 963 -1530
rect 967 -1536 970 -1530
rect 974 -1536 977 -1530
rect 981 -1536 984 -1530
rect 988 -1536 991 -1530
rect 995 -1536 1001 -1530
rect 1002 -1536 1005 -1530
rect 1009 -1536 1012 -1530
rect 1016 -1536 1019 -1530
rect 1044 -1536 1047 -1530
rect 1051 -1536 1054 -1530
rect 1058 -1536 1064 -1530
rect 1 -1613 7 -1607
rect 8 -1613 14 -1607
rect 22 -1613 25 -1607
rect 29 -1613 32 -1607
rect 36 -1613 39 -1607
rect 43 -1613 46 -1607
rect 50 -1613 53 -1607
rect 57 -1613 60 -1607
rect 64 -1613 70 -1607
rect 71 -1613 77 -1607
rect 78 -1613 81 -1607
rect 85 -1613 88 -1607
rect 92 -1613 95 -1607
rect 99 -1613 102 -1607
rect 106 -1613 112 -1607
rect 113 -1613 116 -1607
rect 120 -1613 123 -1607
rect 127 -1613 130 -1607
rect 134 -1613 137 -1607
rect 141 -1613 144 -1607
rect 148 -1613 154 -1607
rect 155 -1613 161 -1607
rect 162 -1613 165 -1607
rect 169 -1613 175 -1607
rect 176 -1613 179 -1607
rect 183 -1613 186 -1607
rect 190 -1613 193 -1607
rect 197 -1613 203 -1607
rect 204 -1613 207 -1607
rect 211 -1613 214 -1607
rect 218 -1613 221 -1607
rect 225 -1613 231 -1607
rect 232 -1613 235 -1607
rect 239 -1613 242 -1607
rect 246 -1613 249 -1607
rect 253 -1613 256 -1607
rect 260 -1613 263 -1607
rect 267 -1613 270 -1607
rect 274 -1613 277 -1607
rect 281 -1613 284 -1607
rect 288 -1613 291 -1607
rect 295 -1613 298 -1607
rect 302 -1613 308 -1607
rect 309 -1613 315 -1607
rect 316 -1613 319 -1607
rect 323 -1613 326 -1607
rect 330 -1613 333 -1607
rect 337 -1613 340 -1607
rect 344 -1613 347 -1607
rect 351 -1613 357 -1607
rect 358 -1613 361 -1607
rect 365 -1613 368 -1607
rect 372 -1613 378 -1607
rect 379 -1613 382 -1607
rect 386 -1613 392 -1607
rect 393 -1613 399 -1607
rect 400 -1613 403 -1607
rect 407 -1613 410 -1607
rect 414 -1613 417 -1607
rect 421 -1613 427 -1607
rect 428 -1613 431 -1607
rect 435 -1613 438 -1607
rect 442 -1613 445 -1607
rect 449 -1613 452 -1607
rect 456 -1613 459 -1607
rect 463 -1613 466 -1607
rect 470 -1613 473 -1607
rect 477 -1613 480 -1607
rect 484 -1613 487 -1607
rect 491 -1613 494 -1607
rect 498 -1613 501 -1607
rect 505 -1613 508 -1607
rect 512 -1613 515 -1607
rect 519 -1613 525 -1607
rect 526 -1613 532 -1607
rect 533 -1613 536 -1607
rect 540 -1613 543 -1607
rect 547 -1613 550 -1607
rect 554 -1613 560 -1607
rect 561 -1613 567 -1607
rect 568 -1613 574 -1607
rect 575 -1613 578 -1607
rect 582 -1613 585 -1607
rect 589 -1613 592 -1607
rect 596 -1613 599 -1607
rect 603 -1613 606 -1607
rect 610 -1613 616 -1607
rect 617 -1613 620 -1607
rect 624 -1613 630 -1607
rect 631 -1613 634 -1607
rect 638 -1613 641 -1607
rect 645 -1613 648 -1607
rect 652 -1613 655 -1607
rect 659 -1613 662 -1607
rect 666 -1613 669 -1607
rect 673 -1613 676 -1607
rect 680 -1613 686 -1607
rect 687 -1613 690 -1607
rect 694 -1613 700 -1607
rect 701 -1613 704 -1607
rect 708 -1613 711 -1607
rect 715 -1613 718 -1607
rect 722 -1613 725 -1607
rect 729 -1613 732 -1607
rect 736 -1613 739 -1607
rect 743 -1613 746 -1607
rect 750 -1613 753 -1607
rect 757 -1613 760 -1607
rect 764 -1613 767 -1607
rect 771 -1613 774 -1607
rect 778 -1613 781 -1607
rect 785 -1613 788 -1607
rect 792 -1613 795 -1607
rect 799 -1613 802 -1607
rect 806 -1613 809 -1607
rect 813 -1613 816 -1607
rect 820 -1613 823 -1607
rect 827 -1613 830 -1607
rect 834 -1613 837 -1607
rect 841 -1613 844 -1607
rect 848 -1613 851 -1607
rect 855 -1613 861 -1607
rect 862 -1613 865 -1607
rect 869 -1613 872 -1607
rect 876 -1613 879 -1607
rect 883 -1613 886 -1607
rect 890 -1613 893 -1607
rect 897 -1613 900 -1607
rect 904 -1613 907 -1607
rect 911 -1613 914 -1607
rect 918 -1613 921 -1607
rect 925 -1613 928 -1607
rect 932 -1613 938 -1607
rect 939 -1613 942 -1607
rect 946 -1613 949 -1607
rect 953 -1613 956 -1607
rect 960 -1613 963 -1607
rect 1023 -1613 1026 -1607
rect 1037 -1613 1040 -1607
rect 1044 -1613 1050 -1607
rect 1051 -1613 1057 -1607
rect 1 -1678 7 -1672
rect 8 -1678 14 -1672
rect 36 -1678 42 -1672
rect 43 -1678 49 -1672
rect 50 -1678 53 -1672
rect 64 -1678 67 -1672
rect 71 -1678 77 -1672
rect 78 -1678 84 -1672
rect 85 -1678 88 -1672
rect 92 -1678 95 -1672
rect 99 -1678 102 -1672
rect 106 -1678 109 -1672
rect 113 -1678 119 -1672
rect 120 -1678 123 -1672
rect 127 -1678 130 -1672
rect 134 -1678 137 -1672
rect 141 -1678 144 -1672
rect 148 -1678 154 -1672
rect 155 -1678 158 -1672
rect 162 -1678 165 -1672
rect 169 -1678 172 -1672
rect 176 -1678 182 -1672
rect 183 -1678 186 -1672
rect 190 -1678 193 -1672
rect 197 -1678 203 -1672
rect 204 -1678 210 -1672
rect 211 -1678 214 -1672
rect 218 -1678 221 -1672
rect 225 -1678 228 -1672
rect 232 -1678 235 -1672
rect 239 -1678 242 -1672
rect 246 -1678 249 -1672
rect 253 -1678 259 -1672
rect 260 -1678 263 -1672
rect 267 -1678 270 -1672
rect 274 -1678 277 -1672
rect 281 -1678 284 -1672
rect 288 -1678 291 -1672
rect 295 -1678 298 -1672
rect 302 -1678 308 -1672
rect 309 -1678 312 -1672
rect 316 -1678 319 -1672
rect 323 -1678 326 -1672
rect 330 -1678 336 -1672
rect 337 -1678 343 -1672
rect 344 -1678 347 -1672
rect 351 -1678 354 -1672
rect 358 -1678 361 -1672
rect 365 -1678 368 -1672
rect 372 -1678 375 -1672
rect 379 -1678 382 -1672
rect 386 -1678 389 -1672
rect 393 -1678 396 -1672
rect 400 -1678 406 -1672
rect 407 -1678 413 -1672
rect 414 -1678 417 -1672
rect 421 -1678 424 -1672
rect 428 -1678 434 -1672
rect 435 -1678 438 -1672
rect 442 -1678 445 -1672
rect 449 -1678 452 -1672
rect 456 -1678 459 -1672
rect 463 -1678 466 -1672
rect 470 -1678 473 -1672
rect 477 -1678 480 -1672
rect 484 -1678 487 -1672
rect 491 -1678 494 -1672
rect 498 -1678 501 -1672
rect 505 -1678 508 -1672
rect 512 -1678 518 -1672
rect 519 -1678 525 -1672
rect 526 -1678 529 -1672
rect 533 -1678 536 -1672
rect 540 -1678 546 -1672
rect 547 -1678 553 -1672
rect 554 -1678 557 -1672
rect 561 -1678 564 -1672
rect 568 -1678 571 -1672
rect 575 -1678 578 -1672
rect 582 -1678 585 -1672
rect 589 -1678 592 -1672
rect 596 -1678 599 -1672
rect 603 -1678 606 -1672
rect 610 -1678 613 -1672
rect 624 -1678 627 -1672
rect 631 -1678 634 -1672
rect 645 -1678 648 -1672
rect 666 -1678 669 -1672
rect 673 -1678 679 -1672
rect 680 -1678 683 -1672
rect 687 -1678 693 -1672
rect 694 -1678 697 -1672
rect 701 -1678 704 -1672
rect 708 -1678 711 -1672
rect 715 -1678 718 -1672
rect 722 -1678 725 -1672
rect 729 -1678 735 -1672
rect 736 -1678 739 -1672
rect 743 -1678 746 -1672
rect 750 -1678 753 -1672
rect 757 -1678 760 -1672
rect 764 -1678 767 -1672
rect 771 -1678 777 -1672
rect 778 -1678 784 -1672
rect 785 -1678 788 -1672
rect 792 -1678 795 -1672
rect 799 -1678 805 -1672
rect 806 -1678 809 -1672
rect 813 -1678 816 -1672
rect 820 -1678 823 -1672
rect 827 -1678 830 -1672
rect 834 -1678 840 -1672
rect 841 -1678 844 -1672
rect 848 -1678 854 -1672
rect 862 -1678 865 -1672
rect 883 -1678 886 -1672
rect 890 -1678 893 -1672
rect 904 -1678 907 -1672
rect 967 -1678 970 -1672
rect 1023 -1678 1026 -1672
rect 1 -1715 7 -1709
rect 8 -1715 14 -1709
rect 15 -1715 21 -1709
rect 22 -1715 28 -1709
rect 29 -1715 35 -1709
rect 43 -1715 46 -1709
rect 57 -1715 60 -1709
rect 92 -1715 95 -1709
rect 99 -1715 105 -1709
rect 113 -1715 119 -1709
rect 127 -1715 130 -1709
rect 141 -1715 144 -1709
rect 148 -1715 151 -1709
rect 155 -1715 158 -1709
rect 162 -1715 165 -1709
rect 169 -1715 172 -1709
rect 176 -1715 182 -1709
rect 183 -1715 189 -1709
rect 190 -1715 193 -1709
rect 197 -1715 203 -1709
rect 204 -1715 210 -1709
rect 211 -1715 217 -1709
rect 218 -1715 221 -1709
rect 225 -1715 228 -1709
rect 232 -1715 235 -1709
rect 239 -1715 242 -1709
rect 253 -1715 256 -1709
rect 260 -1715 266 -1709
rect 267 -1715 270 -1709
rect 274 -1715 280 -1709
rect 281 -1715 284 -1709
rect 288 -1715 291 -1709
rect 295 -1715 301 -1709
rect 302 -1715 305 -1709
rect 309 -1715 312 -1709
rect 316 -1715 319 -1709
rect 323 -1715 326 -1709
rect 330 -1715 333 -1709
rect 337 -1715 343 -1709
rect 344 -1715 347 -1709
rect 351 -1715 357 -1709
rect 358 -1715 361 -1709
rect 365 -1715 368 -1709
rect 372 -1715 378 -1709
rect 379 -1715 385 -1709
rect 386 -1715 389 -1709
rect 393 -1715 396 -1709
rect 400 -1715 406 -1709
rect 407 -1715 410 -1709
rect 414 -1715 417 -1709
rect 421 -1715 424 -1709
rect 428 -1715 431 -1709
rect 435 -1715 438 -1709
rect 442 -1715 445 -1709
rect 449 -1715 452 -1709
rect 456 -1715 459 -1709
rect 463 -1715 466 -1709
rect 470 -1715 476 -1709
rect 477 -1715 480 -1709
rect 484 -1715 487 -1709
rect 491 -1715 494 -1709
rect 498 -1715 504 -1709
rect 505 -1715 508 -1709
rect 512 -1715 515 -1709
rect 519 -1715 522 -1709
rect 526 -1715 529 -1709
rect 533 -1715 536 -1709
rect 540 -1715 543 -1709
rect 547 -1715 550 -1709
rect 554 -1715 557 -1709
rect 561 -1715 564 -1709
rect 568 -1715 571 -1709
rect 575 -1715 578 -1709
rect 582 -1715 585 -1709
rect 589 -1715 595 -1709
rect 596 -1715 602 -1709
rect 603 -1715 609 -1709
rect 610 -1715 616 -1709
rect 617 -1715 620 -1709
rect 638 -1715 641 -1709
rect 645 -1715 648 -1709
rect 652 -1715 655 -1709
rect 673 -1715 676 -1709
rect 680 -1715 686 -1709
rect 708 -1715 711 -1709
rect 722 -1715 725 -1709
rect 729 -1715 732 -1709
rect 736 -1715 739 -1709
rect 743 -1715 746 -1709
rect 750 -1715 753 -1709
rect 757 -1715 760 -1709
rect 764 -1715 767 -1709
rect 771 -1715 774 -1709
rect 778 -1715 781 -1709
rect 792 -1715 795 -1709
rect 799 -1715 802 -1709
rect 806 -1715 809 -1709
rect 813 -1715 819 -1709
rect 820 -1715 823 -1709
rect 827 -1715 830 -1709
rect 834 -1715 837 -1709
rect 841 -1715 847 -1709
rect 848 -1715 851 -1709
rect 855 -1715 858 -1709
rect 862 -1715 868 -1709
rect 883 -1715 886 -1709
rect 897 -1715 900 -1709
rect 967 -1715 970 -1709
rect 1023 -1715 1026 -1709
rect 1 -1748 7 -1742
rect 8 -1748 14 -1742
rect 15 -1748 21 -1742
rect 43 -1748 46 -1742
rect 57 -1748 63 -1742
rect 64 -1748 67 -1742
rect 99 -1748 102 -1742
rect 106 -1748 109 -1742
rect 113 -1748 119 -1742
rect 120 -1748 123 -1742
rect 127 -1748 133 -1742
rect 134 -1748 140 -1742
rect 141 -1748 147 -1742
rect 148 -1748 154 -1742
rect 155 -1748 161 -1742
rect 162 -1748 165 -1742
rect 169 -1748 175 -1742
rect 176 -1748 179 -1742
rect 183 -1748 186 -1742
rect 190 -1748 193 -1742
rect 204 -1748 207 -1742
rect 211 -1748 217 -1742
rect 218 -1748 224 -1742
rect 225 -1748 231 -1742
rect 232 -1748 235 -1742
rect 239 -1748 242 -1742
rect 246 -1748 249 -1742
rect 274 -1748 277 -1742
rect 295 -1748 298 -1742
rect 302 -1748 305 -1742
rect 309 -1748 312 -1742
rect 316 -1748 319 -1742
rect 323 -1748 326 -1742
rect 330 -1748 333 -1742
rect 337 -1748 340 -1742
rect 344 -1748 347 -1742
rect 351 -1748 354 -1742
rect 358 -1748 361 -1742
rect 365 -1748 371 -1742
rect 372 -1748 375 -1742
rect 379 -1748 382 -1742
rect 386 -1748 389 -1742
rect 393 -1748 396 -1742
rect 400 -1748 406 -1742
rect 407 -1748 413 -1742
rect 414 -1748 417 -1742
rect 421 -1748 424 -1742
rect 428 -1748 431 -1742
rect 435 -1748 438 -1742
rect 442 -1748 448 -1742
rect 449 -1748 452 -1742
rect 456 -1748 459 -1742
rect 463 -1748 466 -1742
rect 470 -1748 476 -1742
rect 477 -1748 480 -1742
rect 484 -1748 490 -1742
rect 491 -1748 494 -1742
rect 498 -1748 501 -1742
rect 505 -1748 511 -1742
rect 512 -1748 515 -1742
rect 519 -1748 522 -1742
rect 526 -1748 532 -1742
rect 533 -1748 536 -1742
rect 540 -1748 543 -1742
rect 547 -1748 550 -1742
rect 554 -1748 560 -1742
rect 561 -1748 567 -1742
rect 568 -1748 571 -1742
rect 575 -1748 578 -1742
rect 582 -1748 588 -1742
rect 589 -1748 592 -1742
rect 596 -1748 599 -1742
rect 645 -1748 648 -1742
rect 652 -1748 658 -1742
rect 701 -1748 704 -1742
rect 708 -1748 711 -1742
rect 715 -1748 721 -1742
rect 722 -1748 725 -1742
rect 729 -1748 732 -1742
rect 736 -1748 739 -1742
rect 743 -1748 746 -1742
rect 750 -1748 753 -1742
rect 757 -1748 760 -1742
rect 764 -1748 767 -1742
rect 771 -1748 777 -1742
rect 778 -1748 784 -1742
rect 785 -1748 788 -1742
rect 792 -1748 795 -1742
rect 799 -1748 802 -1742
rect 806 -1748 809 -1742
rect 827 -1748 830 -1742
rect 841 -1748 844 -1742
rect 855 -1748 858 -1742
rect 883 -1748 886 -1742
rect 897 -1748 900 -1742
rect 967 -1748 970 -1742
rect 974 -1748 980 -1742
rect 1023 -1748 1026 -1742
rect 1 -1775 7 -1769
rect 8 -1775 14 -1769
rect 15 -1775 21 -1769
rect 22 -1775 28 -1769
rect 29 -1775 35 -1769
rect 43 -1775 49 -1769
rect 57 -1775 60 -1769
rect 64 -1775 70 -1769
rect 71 -1775 74 -1769
rect 78 -1775 81 -1769
rect 92 -1775 95 -1769
rect 99 -1775 105 -1769
rect 106 -1775 112 -1769
rect 113 -1775 119 -1769
rect 120 -1775 126 -1769
rect 127 -1775 130 -1769
rect 134 -1775 137 -1769
rect 141 -1775 144 -1769
rect 148 -1775 154 -1769
rect 155 -1775 161 -1769
rect 169 -1775 172 -1769
rect 190 -1775 193 -1769
rect 197 -1775 203 -1769
rect 204 -1775 207 -1769
rect 211 -1775 217 -1769
rect 218 -1775 221 -1769
rect 225 -1775 231 -1769
rect 232 -1775 235 -1769
rect 239 -1775 242 -1769
rect 274 -1775 277 -1769
rect 281 -1775 284 -1769
rect 288 -1775 291 -1769
rect 295 -1775 298 -1769
rect 302 -1775 308 -1769
rect 309 -1775 312 -1769
rect 316 -1775 322 -1769
rect 323 -1775 326 -1769
rect 330 -1775 336 -1769
rect 337 -1775 340 -1769
rect 344 -1775 347 -1769
rect 351 -1775 354 -1769
rect 358 -1775 364 -1769
rect 365 -1775 371 -1769
rect 372 -1775 375 -1769
rect 379 -1775 382 -1769
rect 393 -1775 396 -1769
rect 400 -1775 403 -1769
rect 407 -1775 413 -1769
rect 414 -1775 417 -1769
rect 421 -1775 427 -1769
rect 428 -1775 434 -1769
rect 442 -1775 445 -1769
rect 449 -1775 452 -1769
rect 456 -1775 459 -1769
rect 463 -1775 466 -1769
rect 470 -1775 473 -1769
rect 477 -1775 480 -1769
rect 505 -1775 508 -1769
rect 512 -1775 515 -1769
rect 526 -1775 529 -1769
rect 561 -1775 564 -1769
rect 708 -1775 711 -1769
rect 715 -1775 721 -1769
rect 722 -1775 725 -1769
rect 729 -1775 732 -1769
rect 736 -1775 739 -1769
rect 743 -1775 749 -1769
rect 750 -1775 753 -1769
rect 757 -1775 760 -1769
rect 771 -1775 774 -1769
rect 778 -1775 784 -1769
rect 792 -1775 795 -1769
rect 813 -1775 816 -1769
rect 827 -1775 830 -1769
rect 841 -1775 847 -1769
rect 855 -1775 861 -1769
rect 876 -1775 882 -1769
rect 883 -1775 886 -1769
rect 897 -1775 900 -1769
rect 1023 -1775 1026 -1769
rect 1 -1796 7 -1790
rect 8 -1796 14 -1790
rect 15 -1796 21 -1790
rect 22 -1796 28 -1790
rect 29 -1796 35 -1790
rect 36 -1796 42 -1790
rect 43 -1796 49 -1790
rect 50 -1796 56 -1790
rect 57 -1796 63 -1790
rect 64 -1796 70 -1790
rect 71 -1796 77 -1790
rect 78 -1796 81 -1790
rect 141 -1796 144 -1790
rect 148 -1796 154 -1790
rect 155 -1796 158 -1790
rect 169 -1796 175 -1790
rect 183 -1796 189 -1790
rect 204 -1796 207 -1790
rect 225 -1796 228 -1790
rect 239 -1796 242 -1790
rect 246 -1796 252 -1790
rect 260 -1796 263 -1790
rect 281 -1796 284 -1790
rect 295 -1796 298 -1790
rect 302 -1796 308 -1790
rect 309 -1796 315 -1790
rect 316 -1796 322 -1790
rect 323 -1796 326 -1790
rect 330 -1796 333 -1790
rect 337 -1796 340 -1790
rect 344 -1796 350 -1790
rect 351 -1796 354 -1790
rect 379 -1796 382 -1790
rect 386 -1796 389 -1790
rect 407 -1796 413 -1790
rect 414 -1796 417 -1790
rect 421 -1796 424 -1790
rect 428 -1796 434 -1790
rect 435 -1796 441 -1790
rect 442 -1796 445 -1790
rect 449 -1796 452 -1790
rect 456 -1796 459 -1790
rect 470 -1796 473 -1790
rect 477 -1796 480 -1790
rect 498 -1796 504 -1790
rect 505 -1796 511 -1790
rect 512 -1796 515 -1790
rect 519 -1796 522 -1790
rect 561 -1796 567 -1790
rect 736 -1796 739 -1790
rect 743 -1796 749 -1790
rect 750 -1796 756 -1790
rect 757 -1796 760 -1790
rect 764 -1796 767 -1790
rect 771 -1796 777 -1790
rect 792 -1796 795 -1790
rect 813 -1796 819 -1790
rect 834 -1796 840 -1790
rect 897 -1796 900 -1790
rect 1023 -1796 1026 -1790
rect 1 -1811 7 -1805
rect 8 -1811 14 -1805
rect 15 -1811 21 -1805
rect 22 -1811 28 -1805
rect 29 -1811 35 -1805
rect 36 -1811 42 -1805
rect 43 -1811 49 -1805
rect 50 -1811 56 -1805
rect 57 -1811 63 -1805
rect 155 -1811 161 -1805
rect 183 -1811 189 -1805
rect 190 -1811 193 -1805
rect 204 -1811 210 -1805
rect 218 -1811 224 -1805
rect 225 -1811 228 -1805
rect 260 -1811 266 -1805
rect 267 -1811 270 -1805
rect 281 -1811 287 -1805
rect 295 -1811 298 -1805
rect 302 -1811 308 -1805
rect 323 -1811 329 -1805
rect 330 -1811 333 -1805
rect 337 -1811 343 -1805
rect 351 -1811 354 -1805
rect 358 -1811 364 -1805
rect 372 -1811 378 -1805
rect 379 -1811 385 -1805
rect 386 -1811 389 -1805
rect 421 -1811 424 -1805
rect 428 -1811 434 -1805
rect 463 -1811 469 -1805
rect 470 -1811 476 -1805
rect 477 -1811 483 -1805
rect 512 -1811 518 -1805
rect 743 -1811 749 -1805
rect 750 -1811 753 -1805
rect 792 -1811 798 -1805
rect 897 -1811 903 -1805
rect 904 -1811 907 -1805
rect 1023 -1811 1029 -1805
<< polysilicon >>
rect 177 -5 178 -3
rect 177 -11 178 -9
rect 184 -5 185 -3
rect 184 -11 185 -9
rect 194 -5 195 -3
rect 198 -5 199 -3
rect 212 -5 213 -3
rect 219 -5 220 -3
rect 219 -11 220 -9
rect 236 -5 237 -3
rect 240 -5 241 -3
rect 240 -11 241 -9
rect 254 -5 255 -3
rect 261 -5 262 -3
rect 261 -11 262 -9
rect 278 -11 279 -9
rect 285 -5 286 -3
rect 289 -5 290 -3
rect 289 -11 290 -9
rect 296 -11 297 -9
rect 303 -5 304 -3
rect 303 -11 304 -9
rect 310 -5 311 -3
rect 317 -11 318 -9
rect 338 -5 339 -3
rect 338 -11 339 -9
rect 348 -5 349 -3
rect 352 -5 353 -3
rect 352 -11 353 -9
rect 359 -5 360 -3
rect 366 -5 367 -3
rect 366 -11 367 -9
rect 408 -5 409 -3
rect 408 -11 409 -9
rect 422 -11 423 -9
rect 460 -11 461 -9
rect 467 -5 468 -3
rect 471 -5 472 -3
rect 471 -11 472 -9
rect 478 -5 479 -3
rect 485 -5 486 -3
rect 485 -11 486 -9
rect 534 -5 535 -3
rect 541 -5 542 -3
rect 541 -11 542 -9
rect 555 -11 556 -9
rect 558 -11 559 -9
rect 576 -5 577 -3
rect 583 -5 584 -3
rect 583 -11 584 -9
rect 604 -5 605 -3
rect 604 -11 605 -9
rect 611 -5 612 -3
rect 621 -11 622 -9
rect 730 -5 731 -3
rect 730 -11 731 -9
rect 740 -5 741 -3
rect 61 -28 62 -26
rect 79 -28 80 -26
rect 114 -22 115 -20
rect 121 -22 122 -20
rect 121 -28 122 -26
rect 128 -28 129 -26
rect 156 -22 157 -20
rect 163 -22 164 -20
rect 163 -28 164 -26
rect 170 -22 171 -20
rect 170 -28 171 -26
rect 180 -28 181 -26
rect 184 -22 185 -20
rect 184 -28 185 -26
rect 215 -22 216 -20
rect 219 -22 220 -20
rect 219 -28 220 -26
rect 226 -22 227 -20
rect 226 -28 227 -26
rect 240 -22 241 -20
rect 240 -28 241 -26
rect 247 -22 248 -20
rect 247 -28 248 -26
rect 254 -22 255 -20
rect 254 -28 255 -26
rect 261 -22 262 -20
rect 271 -28 272 -26
rect 278 -22 279 -20
rect 282 -22 283 -20
rect 282 -28 283 -26
rect 289 -22 290 -20
rect 289 -28 290 -26
rect 296 -22 297 -20
rect 296 -28 297 -26
rect 303 -22 304 -20
rect 303 -28 304 -26
rect 310 -22 311 -20
rect 310 -28 311 -26
rect 317 -22 318 -20
rect 317 -28 318 -26
rect 334 -22 335 -20
rect 338 -22 339 -20
rect 338 -28 339 -26
rect 345 -22 346 -20
rect 345 -28 346 -26
rect 352 -22 353 -20
rect 352 -28 353 -26
rect 359 -22 360 -20
rect 359 -28 360 -26
rect 366 -22 367 -20
rect 366 -28 367 -26
rect 373 -22 374 -20
rect 380 -28 381 -26
rect 411 -28 412 -26
rect 415 -22 416 -20
rect 415 -28 416 -26
rect 425 -22 426 -20
rect 429 -22 430 -20
rect 429 -28 430 -26
rect 436 -28 437 -26
rect 443 -22 444 -20
rect 443 -28 444 -26
rect 450 -22 451 -20
rect 450 -28 451 -26
rect 457 -22 458 -20
rect 457 -28 458 -26
rect 467 -22 468 -20
rect 474 -22 475 -20
rect 478 -22 479 -20
rect 478 -28 479 -26
rect 485 -22 486 -20
rect 485 -28 486 -26
rect 492 -22 493 -20
rect 492 -28 493 -26
rect 527 -22 528 -20
rect 527 -28 528 -26
rect 541 -22 542 -20
rect 541 -28 542 -26
rect 579 -28 580 -26
rect 583 -22 584 -20
rect 583 -28 584 -26
rect 604 -22 605 -20
rect 604 -28 605 -26
rect 611 -22 612 -20
rect 611 -28 612 -26
rect 618 -22 619 -20
rect 618 -28 619 -26
rect 688 -22 689 -20
rect 688 -28 689 -26
rect 698 -22 699 -20
rect 709 -28 710 -26
rect 712 -28 713 -26
rect 730 -22 731 -20
rect 730 -28 731 -26
rect 58 -45 59 -43
rect 58 -51 59 -49
rect 65 -51 66 -49
rect 79 -45 80 -43
rect 79 -51 80 -49
rect 107 -51 108 -49
rect 114 -45 115 -43
rect 114 -51 115 -49
rect 124 -45 125 -43
rect 121 -51 122 -49
rect 128 -45 129 -43
rect 131 -51 132 -49
rect 135 -45 136 -43
rect 135 -51 136 -49
rect 142 -45 143 -43
rect 142 -51 143 -49
rect 152 -45 153 -43
rect 156 -45 157 -43
rect 156 -51 157 -49
rect 163 -45 164 -43
rect 163 -51 164 -49
rect 170 -45 171 -43
rect 173 -45 174 -43
rect 170 -51 171 -49
rect 177 -45 178 -43
rect 177 -51 178 -49
rect 184 -45 185 -43
rect 184 -51 185 -49
rect 191 -51 192 -49
rect 198 -45 199 -43
rect 198 -51 199 -49
rect 208 -51 209 -49
rect 212 -45 213 -43
rect 212 -51 213 -49
rect 222 -51 223 -49
rect 226 -45 227 -43
rect 226 -51 227 -49
rect 229 -51 230 -49
rect 233 -45 234 -43
rect 233 -51 234 -49
rect 240 -45 241 -43
rect 240 -51 241 -49
rect 247 -45 248 -43
rect 247 -51 248 -49
rect 254 -45 255 -43
rect 257 -45 258 -43
rect 261 -45 262 -43
rect 261 -51 262 -49
rect 268 -45 269 -43
rect 268 -51 269 -49
rect 275 -45 276 -43
rect 275 -51 276 -49
rect 282 -45 283 -43
rect 282 -51 283 -49
rect 289 -45 290 -43
rect 289 -51 290 -49
rect 296 -45 297 -43
rect 296 -51 297 -49
rect 303 -45 304 -43
rect 303 -51 304 -49
rect 310 -45 311 -43
rect 310 -51 311 -49
rect 317 -45 318 -43
rect 317 -51 318 -49
rect 324 -45 325 -43
rect 324 -51 325 -49
rect 331 -45 332 -43
rect 334 -45 335 -43
rect 338 -45 339 -43
rect 345 -45 346 -43
rect 345 -51 346 -49
rect 352 -45 353 -43
rect 352 -51 353 -49
rect 359 -45 360 -43
rect 359 -51 360 -49
rect 366 -45 367 -43
rect 366 -51 367 -49
rect 373 -45 374 -43
rect 373 -51 374 -49
rect 380 -45 381 -43
rect 380 -51 381 -49
rect 387 -45 388 -43
rect 397 -45 398 -43
rect 394 -51 395 -49
rect 401 -45 402 -43
rect 401 -51 402 -49
rect 408 -45 409 -43
rect 408 -51 409 -49
rect 425 -45 426 -43
rect 422 -51 423 -49
rect 429 -45 430 -43
rect 429 -51 430 -49
rect 436 -45 437 -43
rect 436 -51 437 -49
rect 443 -51 444 -49
rect 446 -51 447 -49
rect 450 -45 451 -43
rect 450 -51 451 -49
rect 457 -45 458 -43
rect 457 -51 458 -49
rect 471 -45 472 -43
rect 471 -51 472 -49
rect 478 -45 479 -43
rect 478 -51 479 -49
rect 485 -45 486 -43
rect 485 -51 486 -49
rect 499 -45 500 -43
rect 499 -51 500 -49
rect 513 -45 514 -43
rect 513 -51 514 -49
rect 537 -45 538 -43
rect 534 -51 535 -49
rect 541 -45 542 -43
rect 548 -45 549 -43
rect 548 -51 549 -49
rect 555 -45 556 -43
rect 555 -51 556 -49
rect 562 -45 563 -43
rect 562 -51 563 -49
rect 572 -45 573 -43
rect 576 -45 577 -43
rect 576 -51 577 -49
rect 583 -45 584 -43
rect 583 -51 584 -49
rect 590 -51 591 -49
rect 597 -45 598 -43
rect 597 -51 598 -49
rect 604 -45 605 -43
rect 604 -51 605 -49
rect 611 -45 612 -43
rect 611 -51 612 -49
rect 625 -45 626 -43
rect 625 -51 626 -49
rect 632 -45 633 -43
rect 632 -51 633 -49
rect 646 -45 647 -43
rect 653 -51 654 -49
rect 660 -45 661 -43
rect 660 -51 661 -49
rect 688 -45 689 -43
rect 688 -51 689 -49
rect 730 -45 731 -43
rect 730 -51 731 -49
rect 786 -45 787 -43
rect 786 -51 787 -49
rect 807 -45 808 -43
rect 807 -51 808 -49
rect 814 -45 815 -43
rect 898 -51 899 -49
rect 54 -90 55 -88
rect 58 -84 59 -82
rect 58 -90 59 -88
rect 65 -84 66 -82
rect 65 -90 66 -88
rect 79 -84 80 -82
rect 89 -90 90 -88
rect 93 -84 94 -82
rect 93 -90 94 -88
rect 103 -84 104 -82
rect 110 -84 111 -82
rect 114 -84 115 -82
rect 114 -90 115 -88
rect 124 -90 125 -88
rect 128 -84 129 -82
rect 128 -90 129 -88
rect 135 -84 136 -82
rect 135 -90 136 -88
rect 142 -84 143 -82
rect 142 -90 143 -88
rect 149 -84 150 -82
rect 149 -90 150 -88
rect 156 -84 157 -82
rect 156 -90 157 -88
rect 163 -84 164 -82
rect 163 -90 164 -88
rect 170 -84 171 -82
rect 170 -90 171 -88
rect 180 -90 181 -88
rect 184 -84 185 -82
rect 184 -90 185 -88
rect 187 -90 188 -88
rect 191 -84 192 -82
rect 191 -90 192 -88
rect 198 -84 199 -82
rect 198 -90 199 -88
rect 205 -84 206 -82
rect 208 -84 209 -82
rect 205 -90 206 -88
rect 212 -84 213 -82
rect 212 -90 213 -88
rect 222 -90 223 -88
rect 229 -90 230 -88
rect 233 -84 234 -82
rect 233 -90 234 -88
rect 240 -84 241 -82
rect 240 -90 241 -88
rect 247 -84 248 -82
rect 247 -90 248 -88
rect 254 -84 255 -82
rect 254 -90 255 -88
rect 261 -84 262 -82
rect 261 -90 262 -88
rect 268 -84 269 -82
rect 268 -90 269 -88
rect 278 -84 279 -82
rect 282 -84 283 -82
rect 282 -90 283 -88
rect 289 -84 290 -82
rect 289 -90 290 -88
rect 299 -84 300 -82
rect 299 -90 300 -88
rect 303 -84 304 -82
rect 303 -90 304 -88
rect 310 -84 311 -82
rect 317 -84 318 -82
rect 317 -90 318 -88
rect 324 -84 325 -82
rect 324 -90 325 -88
rect 331 -84 332 -82
rect 331 -90 332 -88
rect 338 -84 339 -82
rect 338 -90 339 -88
rect 345 -84 346 -82
rect 345 -90 346 -88
rect 352 -84 353 -82
rect 352 -90 353 -88
rect 359 -90 360 -88
rect 362 -90 363 -88
rect 366 -84 367 -82
rect 366 -90 367 -88
rect 373 -84 374 -82
rect 373 -90 374 -88
rect 380 -84 381 -82
rect 380 -90 381 -88
rect 387 -84 388 -82
rect 387 -90 388 -88
rect 390 -90 391 -88
rect 394 -84 395 -82
rect 397 -90 398 -88
rect 401 -84 402 -82
rect 401 -90 402 -88
rect 408 -84 409 -82
rect 408 -90 409 -88
rect 415 -84 416 -82
rect 415 -90 416 -88
rect 422 -84 423 -82
rect 422 -90 423 -88
rect 429 -84 430 -82
rect 429 -90 430 -88
rect 439 -84 440 -82
rect 436 -90 437 -88
rect 443 -84 444 -82
rect 446 -84 447 -82
rect 450 -84 451 -82
rect 450 -90 451 -88
rect 460 -84 461 -82
rect 467 -84 468 -82
rect 474 -84 475 -82
rect 478 -84 479 -82
rect 478 -90 479 -88
rect 485 -84 486 -82
rect 485 -90 486 -88
rect 495 -84 496 -82
rect 495 -90 496 -88
rect 499 -84 500 -82
rect 499 -90 500 -88
rect 506 -84 507 -82
rect 506 -90 507 -88
rect 513 -84 514 -82
rect 513 -90 514 -88
rect 520 -84 521 -82
rect 520 -90 521 -88
rect 527 -84 528 -82
rect 534 -84 535 -82
rect 534 -90 535 -88
rect 541 -84 542 -82
rect 541 -90 542 -88
rect 548 -84 549 -82
rect 548 -90 549 -88
rect 555 -84 556 -82
rect 555 -90 556 -88
rect 562 -84 563 -82
rect 562 -90 563 -88
rect 569 -84 570 -82
rect 569 -90 570 -88
rect 576 -84 577 -82
rect 576 -90 577 -88
rect 583 -84 584 -82
rect 583 -90 584 -88
rect 590 -84 591 -82
rect 590 -90 591 -88
rect 597 -84 598 -82
rect 597 -90 598 -88
rect 604 -84 605 -82
rect 604 -90 605 -88
rect 611 -84 612 -82
rect 611 -90 612 -88
rect 618 -84 619 -82
rect 618 -90 619 -88
rect 625 -84 626 -82
rect 625 -90 626 -88
rect 632 -84 633 -82
rect 639 -84 640 -82
rect 639 -90 640 -88
rect 646 -84 647 -82
rect 646 -90 647 -88
rect 653 -84 654 -82
rect 653 -90 654 -88
rect 660 -84 661 -82
rect 660 -90 661 -88
rect 674 -84 675 -82
rect 674 -90 675 -88
rect 681 -90 682 -88
rect 702 -84 703 -82
rect 702 -90 703 -88
rect 730 -84 731 -82
rect 730 -90 731 -88
rect 793 -84 794 -82
rect 793 -90 794 -88
rect 807 -84 808 -82
rect 807 -90 808 -88
rect 898 -84 899 -82
rect 898 -90 899 -88
rect 978 -90 979 -88
rect 1087 -84 1088 -82
rect 1087 -90 1088 -88
rect 1097 -84 1098 -82
rect 30 -121 31 -119
rect 30 -127 31 -125
rect 44 -121 45 -119
rect 47 -127 48 -125
rect 51 -121 52 -119
rect 51 -127 52 -125
rect 58 -121 59 -119
rect 58 -127 59 -125
rect 65 -121 66 -119
rect 65 -127 66 -125
rect 93 -121 94 -119
rect 93 -127 94 -125
rect 100 -121 101 -119
rect 100 -127 101 -125
rect 107 -121 108 -119
rect 107 -127 108 -125
rect 114 -121 115 -119
rect 121 -121 122 -119
rect 121 -127 122 -125
rect 128 -121 129 -119
rect 128 -127 129 -125
rect 135 -127 136 -125
rect 138 -127 139 -125
rect 142 -121 143 -119
rect 142 -127 143 -125
rect 149 -121 150 -119
rect 149 -127 150 -125
rect 156 -121 157 -119
rect 156 -127 157 -125
rect 163 -121 164 -119
rect 163 -127 164 -125
rect 170 -121 171 -119
rect 170 -127 171 -125
rect 177 -121 178 -119
rect 180 -121 181 -119
rect 177 -127 178 -125
rect 187 -127 188 -125
rect 191 -121 192 -119
rect 191 -127 192 -125
rect 198 -121 199 -119
rect 198 -127 199 -125
rect 205 -121 206 -119
rect 205 -127 206 -125
rect 212 -121 213 -119
rect 212 -127 213 -125
rect 219 -121 220 -119
rect 219 -127 220 -125
rect 229 -121 230 -119
rect 229 -127 230 -125
rect 233 -121 234 -119
rect 233 -127 234 -125
rect 240 -121 241 -119
rect 243 -127 244 -125
rect 247 -127 248 -125
rect 250 -127 251 -125
rect 254 -121 255 -119
rect 254 -127 255 -125
rect 261 -121 262 -119
rect 261 -127 262 -125
rect 268 -121 269 -119
rect 268 -127 269 -125
rect 275 -121 276 -119
rect 275 -127 276 -125
rect 282 -121 283 -119
rect 282 -127 283 -125
rect 289 -121 290 -119
rect 289 -127 290 -125
rect 299 -121 300 -119
rect 303 -121 304 -119
rect 303 -127 304 -125
rect 310 -127 311 -125
rect 317 -121 318 -119
rect 317 -127 318 -125
rect 324 -121 325 -119
rect 327 -121 328 -119
rect 324 -127 325 -125
rect 331 -121 332 -119
rect 331 -127 332 -125
rect 338 -121 339 -119
rect 338 -127 339 -125
rect 345 -121 346 -119
rect 345 -127 346 -125
rect 355 -121 356 -119
rect 352 -127 353 -125
rect 359 -121 360 -119
rect 359 -127 360 -125
rect 366 -121 367 -119
rect 366 -127 367 -125
rect 373 -121 374 -119
rect 376 -127 377 -125
rect 380 -127 381 -125
rect 383 -127 384 -125
rect 387 -121 388 -119
rect 390 -121 391 -119
rect 387 -127 388 -125
rect 394 -121 395 -119
rect 394 -127 395 -125
rect 401 -121 402 -119
rect 401 -127 402 -125
rect 408 -121 409 -119
rect 411 -121 412 -119
rect 415 -121 416 -119
rect 415 -127 416 -125
rect 422 -121 423 -119
rect 422 -127 423 -125
rect 429 -121 430 -119
rect 429 -127 430 -125
rect 436 -121 437 -119
rect 436 -127 437 -125
rect 443 -121 444 -119
rect 443 -127 444 -125
rect 450 -121 451 -119
rect 450 -127 451 -125
rect 457 -121 458 -119
rect 457 -127 458 -125
rect 467 -121 468 -119
rect 464 -127 465 -125
rect 471 -121 472 -119
rect 471 -127 472 -125
rect 478 -127 479 -125
rect 481 -127 482 -125
rect 485 -121 486 -119
rect 485 -127 486 -125
rect 492 -121 493 -119
rect 492 -127 493 -125
rect 499 -121 500 -119
rect 499 -127 500 -125
rect 509 -127 510 -125
rect 513 -121 514 -119
rect 513 -127 514 -125
rect 520 -121 521 -119
rect 520 -127 521 -125
rect 527 -121 528 -119
rect 527 -127 528 -125
rect 534 -121 535 -119
rect 534 -127 535 -125
rect 541 -121 542 -119
rect 541 -127 542 -125
rect 548 -127 549 -125
rect 555 -127 556 -125
rect 562 -121 563 -119
rect 562 -127 563 -125
rect 569 -121 570 -119
rect 569 -127 570 -125
rect 576 -121 577 -119
rect 576 -127 577 -125
rect 583 -121 584 -119
rect 583 -127 584 -125
rect 593 -121 594 -119
rect 593 -127 594 -125
rect 597 -121 598 -119
rect 597 -127 598 -125
rect 604 -121 605 -119
rect 604 -127 605 -125
rect 611 -121 612 -119
rect 611 -127 612 -125
rect 618 -121 619 -119
rect 618 -127 619 -125
rect 625 -121 626 -119
rect 625 -127 626 -125
rect 632 -121 633 -119
rect 632 -127 633 -125
rect 639 -121 640 -119
rect 639 -127 640 -125
rect 646 -121 647 -119
rect 646 -127 647 -125
rect 656 -127 657 -125
rect 660 -121 661 -119
rect 660 -127 661 -125
rect 667 -121 668 -119
rect 667 -127 668 -125
rect 674 -121 675 -119
rect 674 -127 675 -125
rect 681 -121 682 -119
rect 681 -127 682 -125
rect 688 -121 689 -119
rect 688 -127 689 -125
rect 695 -121 696 -119
rect 695 -127 696 -125
rect 702 -121 703 -119
rect 702 -127 703 -125
rect 709 -127 710 -125
rect 716 -121 717 -119
rect 716 -127 717 -125
rect 723 -121 724 -119
rect 723 -127 724 -125
rect 730 -121 731 -119
rect 730 -127 731 -125
rect 737 -121 738 -119
rect 737 -127 738 -125
rect 758 -121 759 -119
rect 765 -121 766 -119
rect 765 -127 766 -125
rect 779 -121 780 -119
rect 779 -127 780 -125
rect 800 -121 801 -119
rect 800 -127 801 -125
rect 905 -121 906 -119
rect 905 -127 906 -125
rect 975 -121 976 -119
rect 975 -127 976 -125
rect 1087 -121 1088 -119
rect 1087 -127 1088 -125
rect 23 -182 24 -180
rect 23 -188 24 -186
rect 30 -182 31 -180
rect 30 -188 31 -186
rect 37 -182 38 -180
rect 44 -182 45 -180
rect 51 -182 52 -180
rect 51 -188 52 -186
rect 58 -182 59 -180
rect 58 -188 59 -186
rect 65 -188 66 -186
rect 68 -188 69 -186
rect 72 -182 73 -180
rect 72 -188 73 -186
rect 79 -182 80 -180
rect 79 -188 80 -186
rect 86 -182 87 -180
rect 93 -182 94 -180
rect 93 -188 94 -186
rect 100 -182 101 -180
rect 100 -188 101 -186
rect 107 -182 108 -180
rect 107 -188 108 -186
rect 114 -182 115 -180
rect 114 -188 115 -186
rect 121 -182 122 -180
rect 121 -188 122 -186
rect 128 -182 129 -180
rect 128 -188 129 -186
rect 138 -182 139 -180
rect 142 -182 143 -180
rect 142 -188 143 -186
rect 149 -182 150 -180
rect 149 -188 150 -186
rect 156 -182 157 -180
rect 156 -188 157 -186
rect 166 -182 167 -180
rect 170 -182 171 -180
rect 170 -188 171 -186
rect 177 -182 178 -180
rect 177 -188 178 -186
rect 184 -182 185 -180
rect 187 -188 188 -186
rect 191 -182 192 -180
rect 191 -188 192 -186
rect 198 -188 199 -186
rect 201 -188 202 -186
rect 205 -182 206 -180
rect 212 -182 213 -180
rect 212 -188 213 -186
rect 219 -182 220 -180
rect 219 -188 220 -186
rect 226 -182 227 -180
rect 226 -188 227 -186
rect 233 -182 234 -180
rect 233 -188 234 -186
rect 240 -182 241 -180
rect 240 -188 241 -186
rect 247 -182 248 -180
rect 247 -188 248 -186
rect 254 -182 255 -180
rect 254 -188 255 -186
rect 261 -182 262 -180
rect 261 -188 262 -186
rect 268 -182 269 -180
rect 268 -188 269 -186
rect 275 -182 276 -180
rect 275 -188 276 -186
rect 282 -182 283 -180
rect 282 -188 283 -186
rect 289 -182 290 -180
rect 289 -188 290 -186
rect 296 -182 297 -180
rect 296 -188 297 -186
rect 303 -182 304 -180
rect 303 -188 304 -186
rect 310 -182 311 -180
rect 310 -188 311 -186
rect 317 -182 318 -180
rect 320 -182 321 -180
rect 317 -188 318 -186
rect 324 -182 325 -180
rect 324 -188 325 -186
rect 331 -182 332 -180
rect 334 -182 335 -180
rect 338 -182 339 -180
rect 345 -182 346 -180
rect 348 -182 349 -180
rect 345 -188 346 -186
rect 348 -188 349 -186
rect 352 -182 353 -180
rect 352 -188 353 -186
rect 359 -182 360 -180
rect 359 -188 360 -186
rect 366 -182 367 -180
rect 366 -188 367 -186
rect 376 -182 377 -180
rect 373 -188 374 -186
rect 380 -182 381 -180
rect 380 -188 381 -186
rect 387 -182 388 -180
rect 390 -182 391 -180
rect 394 -182 395 -180
rect 394 -188 395 -186
rect 401 -182 402 -180
rect 401 -188 402 -186
rect 408 -182 409 -180
rect 408 -188 409 -186
rect 415 -182 416 -180
rect 415 -188 416 -186
rect 422 -182 423 -180
rect 422 -188 423 -186
rect 425 -188 426 -186
rect 429 -182 430 -180
rect 429 -188 430 -186
rect 436 -182 437 -180
rect 436 -188 437 -186
rect 443 -182 444 -180
rect 443 -188 444 -186
rect 450 -182 451 -180
rect 450 -188 451 -186
rect 457 -182 458 -180
rect 457 -188 458 -186
rect 467 -182 468 -180
rect 467 -188 468 -186
rect 471 -182 472 -180
rect 471 -188 472 -186
rect 478 -182 479 -180
rect 478 -188 479 -186
rect 488 -182 489 -180
rect 485 -188 486 -186
rect 495 -182 496 -180
rect 499 -182 500 -180
rect 499 -188 500 -186
rect 506 -182 507 -180
rect 506 -188 507 -186
rect 513 -182 514 -180
rect 513 -188 514 -186
rect 523 -182 524 -180
rect 527 -182 528 -180
rect 527 -188 528 -186
rect 537 -182 538 -180
rect 537 -188 538 -186
rect 541 -182 542 -180
rect 541 -188 542 -186
rect 548 -182 549 -180
rect 548 -188 549 -186
rect 555 -182 556 -180
rect 555 -188 556 -186
rect 562 -182 563 -180
rect 562 -188 563 -186
rect 569 -182 570 -180
rect 569 -188 570 -186
rect 576 -182 577 -180
rect 576 -188 577 -186
rect 583 -182 584 -180
rect 583 -188 584 -186
rect 590 -182 591 -180
rect 590 -188 591 -186
rect 597 -182 598 -180
rect 597 -188 598 -186
rect 604 -182 605 -180
rect 604 -188 605 -186
rect 611 -182 612 -180
rect 611 -188 612 -186
rect 618 -182 619 -180
rect 618 -188 619 -186
rect 625 -182 626 -180
rect 625 -188 626 -186
rect 632 -182 633 -180
rect 632 -188 633 -186
rect 639 -182 640 -180
rect 639 -188 640 -186
rect 646 -182 647 -180
rect 646 -188 647 -186
rect 653 -182 654 -180
rect 653 -188 654 -186
rect 660 -182 661 -180
rect 660 -188 661 -186
rect 667 -182 668 -180
rect 667 -188 668 -186
rect 674 -182 675 -180
rect 674 -188 675 -186
rect 681 -182 682 -180
rect 681 -188 682 -186
rect 688 -182 689 -180
rect 688 -188 689 -186
rect 695 -182 696 -180
rect 695 -188 696 -186
rect 702 -182 703 -180
rect 702 -188 703 -186
rect 709 -182 710 -180
rect 709 -188 710 -186
rect 716 -182 717 -180
rect 716 -188 717 -186
rect 723 -182 724 -180
rect 723 -188 724 -186
rect 730 -182 731 -180
rect 730 -188 731 -186
rect 737 -182 738 -180
rect 737 -188 738 -186
rect 744 -182 745 -180
rect 744 -188 745 -186
rect 751 -182 752 -180
rect 751 -188 752 -186
rect 758 -182 759 -180
rect 758 -188 759 -186
rect 765 -182 766 -180
rect 765 -188 766 -186
rect 772 -182 773 -180
rect 772 -188 773 -186
rect 779 -182 780 -180
rect 779 -188 780 -186
rect 786 -182 787 -180
rect 786 -188 787 -186
rect 793 -182 794 -180
rect 793 -188 794 -186
rect 800 -182 801 -180
rect 800 -188 801 -186
rect 807 -182 808 -180
rect 807 -188 808 -186
rect 814 -182 815 -180
rect 821 -188 822 -186
rect 828 -188 829 -186
rect 835 -188 836 -186
rect 845 -182 846 -180
rect 849 -182 850 -180
rect 849 -188 850 -186
rect 859 -188 860 -186
rect 919 -182 920 -180
rect 919 -188 920 -186
rect 975 -182 976 -180
rect 975 -188 976 -186
rect 1087 -182 1088 -180
rect 1087 -188 1088 -186
rect 16 -241 17 -239
rect 16 -247 17 -245
rect 23 -241 24 -239
rect 23 -247 24 -245
rect 30 -241 31 -239
rect 30 -247 31 -245
rect 37 -241 38 -239
rect 37 -247 38 -245
rect 44 -241 45 -239
rect 44 -247 45 -245
rect 51 -241 52 -239
rect 51 -247 52 -245
rect 58 -241 59 -239
rect 65 -241 66 -239
rect 68 -241 69 -239
rect 72 -241 73 -239
rect 72 -247 73 -245
rect 79 -241 80 -239
rect 79 -247 80 -245
rect 89 -247 90 -245
rect 93 -241 94 -239
rect 93 -247 94 -245
rect 100 -241 101 -239
rect 103 -241 104 -239
rect 103 -247 104 -245
rect 107 -241 108 -239
rect 107 -247 108 -245
rect 114 -241 115 -239
rect 117 -241 118 -239
rect 114 -247 115 -245
rect 117 -247 118 -245
rect 121 -241 122 -239
rect 121 -247 122 -245
rect 128 -241 129 -239
rect 128 -247 129 -245
rect 135 -241 136 -239
rect 135 -247 136 -245
rect 142 -241 143 -239
rect 142 -247 143 -245
rect 149 -241 150 -239
rect 149 -247 150 -245
rect 156 -247 157 -245
rect 159 -247 160 -245
rect 163 -241 164 -239
rect 163 -247 164 -245
rect 173 -241 174 -239
rect 170 -247 171 -245
rect 177 -241 178 -239
rect 177 -247 178 -245
rect 184 -241 185 -239
rect 187 -241 188 -239
rect 191 -241 192 -239
rect 191 -247 192 -245
rect 201 -241 202 -239
rect 205 -241 206 -239
rect 205 -247 206 -245
rect 212 -241 213 -239
rect 212 -247 213 -245
rect 219 -247 220 -245
rect 229 -241 230 -239
rect 226 -247 227 -245
rect 233 -241 234 -239
rect 233 -247 234 -245
rect 240 -241 241 -239
rect 240 -247 241 -245
rect 247 -241 248 -239
rect 247 -247 248 -245
rect 254 -241 255 -239
rect 254 -247 255 -245
rect 261 -247 262 -245
rect 264 -247 265 -245
rect 268 -241 269 -239
rect 268 -247 269 -245
rect 275 -241 276 -239
rect 275 -247 276 -245
rect 282 -241 283 -239
rect 292 -241 293 -239
rect 292 -247 293 -245
rect 296 -241 297 -239
rect 296 -247 297 -245
rect 303 -241 304 -239
rect 303 -247 304 -245
rect 310 -241 311 -239
rect 310 -247 311 -245
rect 317 -241 318 -239
rect 317 -247 318 -245
rect 324 -241 325 -239
rect 324 -247 325 -245
rect 331 -241 332 -239
rect 331 -247 332 -245
rect 338 -241 339 -239
rect 338 -247 339 -245
rect 345 -241 346 -239
rect 345 -247 346 -245
rect 352 -241 353 -239
rect 355 -241 356 -239
rect 359 -241 360 -239
rect 359 -247 360 -245
rect 366 -241 367 -239
rect 366 -247 367 -245
rect 373 -241 374 -239
rect 373 -247 374 -245
rect 380 -247 381 -245
rect 383 -247 384 -245
rect 387 -241 388 -239
rect 387 -247 388 -245
rect 394 -241 395 -239
rect 394 -247 395 -245
rect 401 -241 402 -239
rect 401 -247 402 -245
rect 408 -241 409 -239
rect 408 -247 409 -245
rect 415 -241 416 -239
rect 415 -247 416 -245
rect 422 -241 423 -239
rect 422 -247 423 -245
rect 429 -241 430 -239
rect 429 -247 430 -245
rect 436 -241 437 -239
rect 436 -247 437 -245
rect 443 -241 444 -239
rect 443 -247 444 -245
rect 450 -241 451 -239
rect 450 -247 451 -245
rect 460 -241 461 -239
rect 457 -247 458 -245
rect 464 -241 465 -239
rect 467 -241 468 -239
rect 464 -247 465 -245
rect 471 -241 472 -239
rect 471 -247 472 -245
rect 478 -241 479 -239
rect 478 -247 479 -245
rect 481 -247 482 -245
rect 485 -247 486 -245
rect 495 -241 496 -239
rect 492 -247 493 -245
rect 495 -247 496 -245
rect 499 -241 500 -239
rect 499 -247 500 -245
rect 506 -241 507 -239
rect 506 -247 507 -245
rect 513 -241 514 -239
rect 513 -247 514 -245
rect 520 -241 521 -239
rect 520 -247 521 -245
rect 527 -241 528 -239
rect 527 -247 528 -245
rect 534 -241 535 -239
rect 534 -247 535 -245
rect 541 -241 542 -239
rect 541 -247 542 -245
rect 548 -241 549 -239
rect 548 -247 549 -245
rect 555 -241 556 -239
rect 555 -247 556 -245
rect 562 -241 563 -239
rect 562 -247 563 -245
rect 569 -241 570 -239
rect 569 -247 570 -245
rect 576 -241 577 -239
rect 576 -247 577 -245
rect 583 -241 584 -239
rect 583 -247 584 -245
rect 593 -241 594 -239
rect 593 -247 594 -245
rect 597 -247 598 -245
rect 600 -247 601 -245
rect 604 -241 605 -239
rect 604 -247 605 -245
rect 611 -241 612 -239
rect 611 -247 612 -245
rect 618 -241 619 -239
rect 618 -247 619 -245
rect 625 -241 626 -239
rect 625 -247 626 -245
rect 632 -241 633 -239
rect 632 -247 633 -245
rect 639 -241 640 -239
rect 639 -247 640 -245
rect 646 -247 647 -245
rect 653 -241 654 -239
rect 653 -247 654 -245
rect 660 -241 661 -239
rect 660 -247 661 -245
rect 667 -241 668 -239
rect 667 -247 668 -245
rect 674 -241 675 -239
rect 674 -247 675 -245
rect 681 -241 682 -239
rect 681 -247 682 -245
rect 688 -241 689 -239
rect 688 -247 689 -245
rect 695 -241 696 -239
rect 695 -247 696 -245
rect 702 -241 703 -239
rect 702 -247 703 -245
rect 709 -241 710 -239
rect 709 -247 710 -245
rect 716 -241 717 -239
rect 716 -247 717 -245
rect 723 -241 724 -239
rect 723 -247 724 -245
rect 730 -241 731 -239
rect 730 -247 731 -245
rect 737 -241 738 -239
rect 737 -247 738 -245
rect 744 -241 745 -239
rect 744 -247 745 -245
rect 751 -241 752 -239
rect 751 -247 752 -245
rect 758 -241 759 -239
rect 758 -247 759 -245
rect 765 -241 766 -239
rect 765 -247 766 -245
rect 772 -241 773 -239
rect 772 -247 773 -245
rect 779 -241 780 -239
rect 779 -247 780 -245
rect 786 -241 787 -239
rect 786 -247 787 -245
rect 793 -241 794 -239
rect 793 -247 794 -245
rect 800 -241 801 -239
rect 807 -241 808 -239
rect 807 -247 808 -245
rect 814 -241 815 -239
rect 814 -247 815 -245
rect 821 -241 822 -239
rect 821 -247 822 -245
rect 828 -241 829 -239
rect 828 -247 829 -245
rect 835 -241 836 -239
rect 835 -247 836 -245
rect 842 -241 843 -239
rect 842 -247 843 -245
rect 849 -241 850 -239
rect 849 -247 850 -245
rect 856 -241 857 -239
rect 856 -247 857 -245
rect 863 -241 864 -239
rect 863 -247 864 -245
rect 870 -241 871 -239
rect 870 -247 871 -245
rect 877 -241 878 -239
rect 877 -247 878 -245
rect 884 -241 885 -239
rect 884 -247 885 -245
rect 891 -241 892 -239
rect 891 -247 892 -245
rect 898 -241 899 -239
rect 898 -247 899 -245
rect 905 -241 906 -239
rect 905 -247 906 -245
rect 912 -241 913 -239
rect 912 -247 913 -245
rect 919 -241 920 -239
rect 919 -247 920 -245
rect 926 -241 927 -239
rect 926 -247 927 -245
rect 933 -241 934 -239
rect 933 -247 934 -245
rect 940 -241 941 -239
rect 940 -247 941 -245
rect 947 -241 948 -239
rect 947 -247 948 -245
rect 954 -247 955 -245
rect 975 -241 976 -239
rect 975 -247 976 -245
rect 1087 -241 1088 -239
rect 1087 -247 1088 -245
rect 9 -318 10 -316
rect 16 -312 17 -310
rect 16 -318 17 -316
rect 23 -312 24 -310
rect 23 -318 24 -316
rect 33 -312 34 -310
rect 30 -318 31 -316
rect 37 -312 38 -310
rect 37 -318 38 -316
rect 47 -312 48 -310
rect 58 -312 59 -310
rect 58 -318 59 -316
rect 65 -312 66 -310
rect 65 -318 66 -316
rect 72 -312 73 -310
rect 72 -318 73 -316
rect 79 -312 80 -310
rect 82 -312 83 -310
rect 79 -318 80 -316
rect 86 -312 87 -310
rect 86 -318 87 -316
rect 93 -312 94 -310
rect 93 -318 94 -316
rect 100 -312 101 -310
rect 100 -318 101 -316
rect 107 -318 108 -316
rect 110 -318 111 -316
rect 114 -312 115 -310
rect 114 -318 115 -316
rect 121 -312 122 -310
rect 121 -318 122 -316
rect 128 -312 129 -310
rect 128 -318 129 -316
rect 135 -312 136 -310
rect 135 -318 136 -316
rect 145 -312 146 -310
rect 145 -318 146 -316
rect 149 -312 150 -310
rect 149 -318 150 -316
rect 156 -312 157 -310
rect 156 -318 157 -316
rect 163 -312 164 -310
rect 163 -318 164 -316
rect 170 -312 171 -310
rect 170 -318 171 -316
rect 177 -312 178 -310
rect 177 -318 178 -316
rect 184 -312 185 -310
rect 184 -318 185 -316
rect 191 -312 192 -310
rect 191 -318 192 -316
rect 198 -312 199 -310
rect 198 -318 199 -316
rect 205 -312 206 -310
rect 208 -312 209 -310
rect 208 -318 209 -316
rect 212 -312 213 -310
rect 212 -318 213 -316
rect 219 -312 220 -310
rect 219 -318 220 -316
rect 229 -312 230 -310
rect 233 -312 234 -310
rect 233 -318 234 -316
rect 240 -312 241 -310
rect 240 -318 241 -316
rect 247 -312 248 -310
rect 247 -318 248 -316
rect 254 -312 255 -310
rect 254 -318 255 -316
rect 261 -312 262 -310
rect 261 -318 262 -316
rect 268 -312 269 -310
rect 268 -318 269 -316
rect 275 -312 276 -310
rect 275 -318 276 -316
rect 282 -312 283 -310
rect 282 -318 283 -316
rect 289 -312 290 -310
rect 292 -318 293 -316
rect 296 -312 297 -310
rect 296 -318 297 -316
rect 303 -312 304 -310
rect 303 -318 304 -316
rect 310 -312 311 -310
rect 310 -318 311 -316
rect 317 -312 318 -310
rect 317 -318 318 -316
rect 324 -312 325 -310
rect 324 -318 325 -316
rect 331 -312 332 -310
rect 331 -318 332 -316
rect 338 -312 339 -310
rect 338 -318 339 -316
rect 345 -312 346 -310
rect 345 -318 346 -316
rect 352 -312 353 -310
rect 352 -318 353 -316
rect 359 -312 360 -310
rect 359 -318 360 -316
rect 366 -312 367 -310
rect 366 -318 367 -316
rect 373 -312 374 -310
rect 373 -318 374 -316
rect 380 -318 381 -316
rect 383 -318 384 -316
rect 387 -318 388 -316
rect 390 -318 391 -316
rect 394 -312 395 -310
rect 394 -318 395 -316
rect 401 -312 402 -310
rect 401 -318 402 -316
rect 411 -312 412 -310
rect 408 -318 409 -316
rect 415 -312 416 -310
rect 418 -318 419 -316
rect 422 -312 423 -310
rect 422 -318 423 -316
rect 429 -312 430 -310
rect 429 -318 430 -316
rect 439 -312 440 -310
rect 436 -318 437 -316
rect 443 -312 444 -310
rect 443 -318 444 -316
rect 450 -312 451 -310
rect 450 -318 451 -316
rect 457 -312 458 -310
rect 457 -318 458 -316
rect 464 -312 465 -310
rect 467 -318 468 -316
rect 471 -312 472 -310
rect 474 -312 475 -310
rect 474 -318 475 -316
rect 478 -312 479 -310
rect 478 -318 479 -316
rect 488 -312 489 -310
rect 485 -318 486 -316
rect 488 -318 489 -316
rect 492 -312 493 -310
rect 492 -318 493 -316
rect 499 -312 500 -310
rect 499 -318 500 -316
rect 506 -312 507 -310
rect 513 -312 514 -310
rect 513 -318 514 -316
rect 520 -312 521 -310
rect 520 -318 521 -316
rect 527 -312 528 -310
rect 527 -318 528 -316
rect 534 -312 535 -310
rect 534 -318 535 -316
rect 541 -318 542 -316
rect 544 -318 545 -316
rect 548 -312 549 -310
rect 548 -318 549 -316
rect 551 -318 552 -316
rect 555 -312 556 -310
rect 555 -318 556 -316
rect 562 -312 563 -310
rect 562 -318 563 -316
rect 569 -312 570 -310
rect 569 -318 570 -316
rect 579 -312 580 -310
rect 583 -312 584 -310
rect 586 -312 587 -310
rect 586 -318 587 -316
rect 590 -312 591 -310
rect 590 -318 591 -316
rect 597 -312 598 -310
rect 597 -318 598 -316
rect 604 -312 605 -310
rect 604 -318 605 -316
rect 611 -312 612 -310
rect 611 -318 612 -316
rect 618 -312 619 -310
rect 618 -318 619 -316
rect 625 -312 626 -310
rect 625 -318 626 -316
rect 632 -312 633 -310
rect 632 -318 633 -316
rect 639 -312 640 -310
rect 639 -318 640 -316
rect 646 -312 647 -310
rect 646 -318 647 -316
rect 653 -312 654 -310
rect 653 -318 654 -316
rect 660 -312 661 -310
rect 660 -318 661 -316
rect 667 -312 668 -310
rect 667 -318 668 -316
rect 674 -312 675 -310
rect 674 -318 675 -316
rect 681 -312 682 -310
rect 681 -318 682 -316
rect 684 -318 685 -316
rect 688 -312 689 -310
rect 688 -318 689 -316
rect 695 -312 696 -310
rect 695 -318 696 -316
rect 702 -312 703 -310
rect 702 -318 703 -316
rect 709 -312 710 -310
rect 709 -318 710 -316
rect 716 -318 717 -316
rect 719 -318 720 -316
rect 723 -312 724 -310
rect 723 -318 724 -316
rect 730 -312 731 -310
rect 730 -318 731 -316
rect 737 -312 738 -310
rect 737 -318 738 -316
rect 744 -312 745 -310
rect 744 -318 745 -316
rect 751 -312 752 -310
rect 751 -318 752 -316
rect 758 -312 759 -310
rect 758 -318 759 -316
rect 765 -312 766 -310
rect 765 -318 766 -316
rect 772 -312 773 -310
rect 772 -318 773 -316
rect 779 -312 780 -310
rect 779 -318 780 -316
rect 786 -312 787 -310
rect 786 -318 787 -316
rect 793 -312 794 -310
rect 793 -318 794 -316
rect 800 -312 801 -310
rect 800 -318 801 -316
rect 807 -312 808 -310
rect 807 -318 808 -316
rect 814 -312 815 -310
rect 814 -318 815 -316
rect 821 -312 822 -310
rect 821 -318 822 -316
rect 828 -312 829 -310
rect 828 -318 829 -316
rect 835 -312 836 -310
rect 835 -318 836 -316
rect 842 -312 843 -310
rect 842 -318 843 -316
rect 849 -312 850 -310
rect 849 -318 850 -316
rect 856 -312 857 -310
rect 856 -318 857 -316
rect 863 -312 864 -310
rect 863 -318 864 -316
rect 870 -312 871 -310
rect 870 -318 871 -316
rect 877 -312 878 -310
rect 877 -318 878 -316
rect 884 -312 885 -310
rect 884 -318 885 -316
rect 891 -312 892 -310
rect 891 -318 892 -316
rect 898 -312 899 -310
rect 898 -318 899 -316
rect 905 -312 906 -310
rect 905 -318 906 -316
rect 912 -312 913 -310
rect 912 -318 913 -316
rect 919 -312 920 -310
rect 919 -318 920 -316
rect 926 -312 927 -310
rect 926 -318 927 -316
rect 936 -312 937 -310
rect 936 -318 937 -316
rect 940 -312 941 -310
rect 940 -318 941 -316
rect 947 -318 948 -316
rect 954 -312 955 -310
rect 954 -318 955 -316
rect 961 -312 962 -310
rect 961 -318 962 -316
rect 968 -312 969 -310
rect 975 -312 976 -310
rect 975 -318 976 -316
rect 982 -312 983 -310
rect 982 -318 983 -316
rect 1094 -312 1095 -310
rect 1094 -318 1095 -316
rect 16 -397 17 -395
rect 16 -403 17 -401
rect 23 -397 24 -395
rect 23 -403 24 -401
rect 33 -397 34 -395
rect 40 -397 41 -395
rect 44 -397 45 -395
rect 44 -403 45 -401
rect 51 -397 52 -395
rect 51 -403 52 -401
rect 58 -397 59 -395
rect 58 -403 59 -401
rect 65 -397 66 -395
rect 65 -403 66 -401
rect 72 -397 73 -395
rect 72 -403 73 -401
rect 79 -397 80 -395
rect 79 -403 80 -401
rect 86 -397 87 -395
rect 86 -403 87 -401
rect 93 -397 94 -395
rect 93 -403 94 -401
rect 100 -397 101 -395
rect 100 -403 101 -401
rect 107 -397 108 -395
rect 107 -403 108 -401
rect 117 -397 118 -395
rect 114 -403 115 -401
rect 121 -397 122 -395
rect 121 -403 122 -401
rect 128 -397 129 -395
rect 128 -403 129 -401
rect 135 -397 136 -395
rect 138 -403 139 -401
rect 145 -397 146 -395
rect 142 -403 143 -401
rect 145 -403 146 -401
rect 149 -397 150 -395
rect 149 -403 150 -401
rect 156 -397 157 -395
rect 156 -403 157 -401
rect 163 -397 164 -395
rect 163 -403 164 -401
rect 170 -403 171 -401
rect 173 -403 174 -401
rect 180 -397 181 -395
rect 177 -403 178 -401
rect 180 -403 181 -401
rect 184 -397 185 -395
rect 184 -403 185 -401
rect 191 -397 192 -395
rect 191 -403 192 -401
rect 198 -397 199 -395
rect 198 -403 199 -401
rect 205 -397 206 -395
rect 208 -397 209 -395
rect 208 -403 209 -401
rect 212 -397 213 -395
rect 212 -403 213 -401
rect 219 -397 220 -395
rect 219 -403 220 -401
rect 226 -397 227 -395
rect 226 -403 227 -401
rect 233 -397 234 -395
rect 233 -403 234 -401
rect 240 -397 241 -395
rect 240 -403 241 -401
rect 247 -397 248 -395
rect 247 -403 248 -401
rect 254 -397 255 -395
rect 254 -403 255 -401
rect 261 -397 262 -395
rect 268 -397 269 -395
rect 268 -403 269 -401
rect 275 -397 276 -395
rect 278 -403 279 -401
rect 282 -397 283 -395
rect 282 -403 283 -401
rect 285 -403 286 -401
rect 289 -397 290 -395
rect 289 -403 290 -401
rect 296 -397 297 -395
rect 296 -403 297 -401
rect 303 -397 304 -395
rect 303 -403 304 -401
rect 310 -397 311 -395
rect 310 -403 311 -401
rect 317 -403 318 -401
rect 320 -403 321 -401
rect 324 -397 325 -395
rect 324 -403 325 -401
rect 331 -397 332 -395
rect 331 -403 332 -401
rect 338 -397 339 -395
rect 338 -403 339 -401
rect 341 -403 342 -401
rect 345 -397 346 -395
rect 345 -403 346 -401
rect 352 -397 353 -395
rect 352 -403 353 -401
rect 359 -397 360 -395
rect 366 -397 367 -395
rect 366 -403 367 -401
rect 373 -397 374 -395
rect 373 -403 374 -401
rect 380 -397 381 -395
rect 380 -403 381 -401
rect 387 -397 388 -395
rect 387 -403 388 -401
rect 394 -397 395 -395
rect 394 -403 395 -401
rect 401 -397 402 -395
rect 404 -397 405 -395
rect 404 -403 405 -401
rect 408 -397 409 -395
rect 408 -403 409 -401
rect 415 -397 416 -395
rect 415 -403 416 -401
rect 422 -397 423 -395
rect 425 -403 426 -401
rect 429 -397 430 -395
rect 429 -403 430 -401
rect 436 -397 437 -395
rect 436 -403 437 -401
rect 443 -397 444 -395
rect 443 -403 444 -401
rect 450 -397 451 -395
rect 453 -397 454 -395
rect 457 -397 458 -395
rect 457 -403 458 -401
rect 464 -397 465 -395
rect 464 -403 465 -401
rect 474 -397 475 -395
rect 478 -397 479 -395
rect 478 -403 479 -401
rect 485 -397 486 -395
rect 485 -403 486 -401
rect 492 -397 493 -395
rect 495 -397 496 -395
rect 492 -403 493 -401
rect 499 -397 500 -395
rect 499 -403 500 -401
rect 506 -397 507 -395
rect 513 -397 514 -395
rect 513 -403 514 -401
rect 520 -397 521 -395
rect 523 -397 524 -395
rect 520 -403 521 -401
rect 527 -397 528 -395
rect 527 -403 528 -401
rect 534 -397 535 -395
rect 534 -403 535 -401
rect 541 -397 542 -395
rect 541 -403 542 -401
rect 548 -397 549 -395
rect 551 -397 552 -395
rect 551 -403 552 -401
rect 555 -397 556 -395
rect 555 -403 556 -401
rect 562 -397 563 -395
rect 565 -397 566 -395
rect 569 -397 570 -395
rect 569 -403 570 -401
rect 579 -397 580 -395
rect 579 -403 580 -401
rect 583 -397 584 -395
rect 583 -403 584 -401
rect 590 -397 591 -395
rect 590 -403 591 -401
rect 597 -397 598 -395
rect 597 -403 598 -401
rect 604 -397 605 -395
rect 604 -403 605 -401
rect 611 -397 612 -395
rect 611 -403 612 -401
rect 618 -397 619 -395
rect 618 -403 619 -401
rect 625 -397 626 -395
rect 625 -403 626 -401
rect 632 -397 633 -395
rect 632 -403 633 -401
rect 639 -397 640 -395
rect 639 -403 640 -401
rect 646 -397 647 -395
rect 646 -403 647 -401
rect 653 -397 654 -395
rect 653 -403 654 -401
rect 660 -397 661 -395
rect 660 -403 661 -401
rect 667 -397 668 -395
rect 667 -403 668 -401
rect 674 -397 675 -395
rect 674 -403 675 -401
rect 681 -397 682 -395
rect 684 -397 685 -395
rect 681 -403 682 -401
rect 688 -397 689 -395
rect 688 -403 689 -401
rect 695 -397 696 -395
rect 695 -403 696 -401
rect 702 -397 703 -395
rect 702 -403 703 -401
rect 709 -397 710 -395
rect 709 -403 710 -401
rect 716 -397 717 -395
rect 716 -403 717 -401
rect 723 -397 724 -395
rect 723 -403 724 -401
rect 730 -397 731 -395
rect 730 -403 731 -401
rect 737 -397 738 -395
rect 737 -403 738 -401
rect 744 -397 745 -395
rect 744 -403 745 -401
rect 751 -397 752 -395
rect 751 -403 752 -401
rect 758 -397 759 -395
rect 758 -403 759 -401
rect 765 -397 766 -395
rect 765 -403 766 -401
rect 772 -397 773 -395
rect 772 -403 773 -401
rect 779 -397 780 -395
rect 779 -403 780 -401
rect 786 -397 787 -395
rect 786 -403 787 -401
rect 793 -397 794 -395
rect 793 -403 794 -401
rect 800 -397 801 -395
rect 800 -403 801 -401
rect 807 -397 808 -395
rect 807 -403 808 -401
rect 814 -397 815 -395
rect 814 -403 815 -401
rect 821 -397 822 -395
rect 821 -403 822 -401
rect 828 -397 829 -395
rect 828 -403 829 -401
rect 835 -397 836 -395
rect 835 -403 836 -401
rect 842 -397 843 -395
rect 842 -403 843 -401
rect 849 -397 850 -395
rect 849 -403 850 -401
rect 856 -397 857 -395
rect 856 -403 857 -401
rect 863 -397 864 -395
rect 863 -403 864 -401
rect 870 -397 871 -395
rect 870 -403 871 -401
rect 877 -397 878 -395
rect 877 -403 878 -401
rect 884 -397 885 -395
rect 884 -403 885 -401
rect 891 -397 892 -395
rect 891 -403 892 -401
rect 901 -397 902 -395
rect 901 -403 902 -401
rect 905 -397 906 -395
rect 905 -403 906 -401
rect 912 -397 913 -395
rect 912 -403 913 -401
rect 919 -397 920 -395
rect 919 -403 920 -401
rect 926 -397 927 -395
rect 926 -403 927 -401
rect 933 -397 934 -395
rect 933 -403 934 -401
rect 940 -397 941 -395
rect 940 -403 941 -401
rect 947 -397 948 -395
rect 947 -403 948 -401
rect 954 -397 955 -395
rect 954 -403 955 -401
rect 961 -397 962 -395
rect 964 -397 965 -395
rect 961 -403 962 -401
rect 968 -397 969 -395
rect 968 -403 969 -401
rect 975 -397 976 -395
rect 975 -403 976 -401
rect 982 -397 983 -395
rect 982 -403 983 -401
rect 989 -397 990 -395
rect 989 -403 990 -401
rect 999 -397 1000 -395
rect 996 -403 997 -401
rect 1003 -397 1004 -395
rect 1003 -403 1004 -401
rect 1010 -397 1011 -395
rect 1010 -403 1011 -401
rect 1017 -397 1018 -395
rect 1017 -403 1018 -401
rect 1024 -397 1025 -395
rect 1024 -403 1025 -401
rect 1031 -403 1032 -401
rect 1041 -403 1042 -401
rect 1048 -403 1049 -401
rect 1052 -397 1053 -395
rect 1052 -403 1053 -401
rect 1066 -397 1067 -395
rect 1066 -403 1067 -401
rect 1108 -397 1109 -395
rect 1108 -403 1109 -401
rect 12 -466 13 -464
rect 16 -466 17 -464
rect 16 -472 17 -470
rect 23 -466 24 -464
rect 23 -472 24 -470
rect 30 -466 31 -464
rect 30 -472 31 -470
rect 37 -466 38 -464
rect 37 -472 38 -470
rect 44 -466 45 -464
rect 44 -472 45 -470
rect 51 -466 52 -464
rect 51 -472 52 -470
rect 58 -466 59 -464
rect 58 -472 59 -470
rect 65 -466 66 -464
rect 65 -472 66 -470
rect 72 -466 73 -464
rect 72 -472 73 -470
rect 79 -466 80 -464
rect 79 -472 80 -470
rect 86 -466 87 -464
rect 89 -466 90 -464
rect 86 -472 87 -470
rect 93 -466 94 -464
rect 93 -472 94 -470
rect 100 -466 101 -464
rect 100 -472 101 -470
rect 110 -466 111 -464
rect 110 -472 111 -470
rect 114 -466 115 -464
rect 114 -472 115 -470
rect 121 -466 122 -464
rect 121 -472 122 -470
rect 128 -466 129 -464
rect 128 -472 129 -470
rect 135 -466 136 -464
rect 138 -472 139 -470
rect 142 -466 143 -464
rect 142 -472 143 -470
rect 149 -466 150 -464
rect 149 -472 150 -470
rect 156 -466 157 -464
rect 156 -472 157 -470
rect 163 -466 164 -464
rect 163 -472 164 -470
rect 170 -466 171 -464
rect 170 -472 171 -470
rect 177 -466 178 -464
rect 177 -472 178 -470
rect 184 -466 185 -464
rect 184 -472 185 -470
rect 191 -466 192 -464
rect 191 -472 192 -470
rect 198 -466 199 -464
rect 198 -472 199 -470
rect 205 -466 206 -464
rect 205 -472 206 -470
rect 215 -472 216 -470
rect 219 -466 220 -464
rect 219 -472 220 -470
rect 229 -466 230 -464
rect 233 -466 234 -464
rect 233 -472 234 -470
rect 240 -466 241 -464
rect 240 -472 241 -470
rect 247 -466 248 -464
rect 247 -472 248 -470
rect 254 -466 255 -464
rect 254 -472 255 -470
rect 261 -472 262 -470
rect 268 -466 269 -464
rect 268 -472 269 -470
rect 275 -466 276 -464
rect 278 -466 279 -464
rect 278 -472 279 -470
rect 282 -466 283 -464
rect 285 -466 286 -464
rect 282 -472 283 -470
rect 289 -466 290 -464
rect 289 -472 290 -470
rect 296 -466 297 -464
rect 296 -472 297 -470
rect 303 -466 304 -464
rect 306 -466 307 -464
rect 303 -472 304 -470
rect 310 -466 311 -464
rect 310 -472 311 -470
rect 317 -466 318 -464
rect 317 -472 318 -470
rect 324 -466 325 -464
rect 324 -472 325 -470
rect 331 -466 332 -464
rect 331 -472 332 -470
rect 338 -466 339 -464
rect 338 -472 339 -470
rect 345 -466 346 -464
rect 348 -472 349 -470
rect 352 -466 353 -464
rect 352 -472 353 -470
rect 359 -466 360 -464
rect 359 -472 360 -470
rect 366 -466 367 -464
rect 366 -472 367 -470
rect 373 -466 374 -464
rect 373 -472 374 -470
rect 380 -466 381 -464
rect 380 -472 381 -470
rect 390 -466 391 -464
rect 387 -472 388 -470
rect 390 -472 391 -470
rect 394 -466 395 -464
rect 394 -472 395 -470
rect 401 -466 402 -464
rect 404 -466 405 -464
rect 401 -472 402 -470
rect 404 -472 405 -470
rect 408 -466 409 -464
rect 411 -466 412 -464
rect 408 -472 409 -470
rect 415 -466 416 -464
rect 415 -472 416 -470
rect 422 -466 423 -464
rect 422 -472 423 -470
rect 429 -466 430 -464
rect 429 -472 430 -470
rect 436 -466 437 -464
rect 436 -472 437 -470
rect 443 -466 444 -464
rect 443 -472 444 -470
rect 450 -466 451 -464
rect 450 -472 451 -470
rect 457 -466 458 -464
rect 460 -472 461 -470
rect 464 -466 465 -464
rect 464 -472 465 -470
rect 471 -466 472 -464
rect 474 -466 475 -464
rect 471 -472 472 -470
rect 478 -466 479 -464
rect 478 -472 479 -470
rect 485 -466 486 -464
rect 485 -472 486 -470
rect 492 -466 493 -464
rect 492 -472 493 -470
rect 502 -466 503 -464
rect 502 -472 503 -470
rect 509 -466 510 -464
rect 509 -472 510 -470
rect 513 -466 514 -464
rect 513 -472 514 -470
rect 520 -466 521 -464
rect 523 -466 524 -464
rect 527 -466 528 -464
rect 527 -472 528 -470
rect 530 -472 531 -470
rect 534 -466 535 -464
rect 534 -472 535 -470
rect 541 -466 542 -464
rect 541 -472 542 -470
rect 548 -466 549 -464
rect 548 -472 549 -470
rect 555 -466 556 -464
rect 555 -472 556 -470
rect 562 -466 563 -464
rect 565 -466 566 -464
rect 562 -472 563 -470
rect 569 -466 570 -464
rect 569 -472 570 -470
rect 576 -466 577 -464
rect 576 -472 577 -470
rect 583 -466 584 -464
rect 586 -466 587 -464
rect 586 -472 587 -470
rect 590 -466 591 -464
rect 590 -472 591 -470
rect 597 -466 598 -464
rect 600 -466 601 -464
rect 597 -472 598 -470
rect 600 -472 601 -470
rect 604 -466 605 -464
rect 604 -472 605 -470
rect 611 -466 612 -464
rect 611 -472 612 -470
rect 618 -466 619 -464
rect 618 -472 619 -470
rect 625 -466 626 -464
rect 625 -472 626 -470
rect 635 -466 636 -464
rect 632 -472 633 -470
rect 635 -472 636 -470
rect 639 -466 640 -464
rect 639 -472 640 -470
rect 646 -466 647 -464
rect 646 -472 647 -470
rect 653 -466 654 -464
rect 653 -472 654 -470
rect 660 -466 661 -464
rect 660 -472 661 -470
rect 667 -466 668 -464
rect 667 -472 668 -470
rect 674 -466 675 -464
rect 674 -472 675 -470
rect 681 -466 682 -464
rect 681 -472 682 -470
rect 688 -466 689 -464
rect 688 -472 689 -470
rect 695 -466 696 -464
rect 695 -472 696 -470
rect 702 -466 703 -464
rect 702 -472 703 -470
rect 709 -466 710 -464
rect 709 -472 710 -470
rect 716 -466 717 -464
rect 716 -472 717 -470
rect 723 -466 724 -464
rect 723 -472 724 -470
rect 730 -466 731 -464
rect 730 -472 731 -470
rect 737 -466 738 -464
rect 740 -466 741 -464
rect 744 -466 745 -464
rect 744 -472 745 -470
rect 754 -466 755 -464
rect 754 -472 755 -470
rect 758 -466 759 -464
rect 758 -472 759 -470
rect 765 -466 766 -464
rect 765 -472 766 -470
rect 772 -466 773 -464
rect 772 -472 773 -470
rect 779 -466 780 -464
rect 779 -472 780 -470
rect 786 -466 787 -464
rect 786 -472 787 -470
rect 793 -466 794 -464
rect 793 -472 794 -470
rect 800 -466 801 -464
rect 800 -472 801 -470
rect 807 -466 808 -464
rect 807 -472 808 -470
rect 814 -466 815 -464
rect 814 -472 815 -470
rect 821 -466 822 -464
rect 821 -472 822 -470
rect 828 -466 829 -464
rect 828 -472 829 -470
rect 835 -466 836 -464
rect 835 -472 836 -470
rect 842 -466 843 -464
rect 842 -472 843 -470
rect 849 -466 850 -464
rect 849 -472 850 -470
rect 856 -466 857 -464
rect 856 -472 857 -470
rect 863 -466 864 -464
rect 863 -472 864 -470
rect 870 -466 871 -464
rect 870 -472 871 -470
rect 877 -466 878 -464
rect 877 -472 878 -470
rect 884 -466 885 -464
rect 884 -472 885 -470
rect 891 -466 892 -464
rect 891 -472 892 -470
rect 898 -466 899 -464
rect 898 -472 899 -470
rect 905 -466 906 -464
rect 905 -472 906 -470
rect 912 -466 913 -464
rect 912 -472 913 -470
rect 919 -466 920 -464
rect 919 -472 920 -470
rect 926 -466 927 -464
rect 926 -472 927 -470
rect 933 -466 934 -464
rect 933 -472 934 -470
rect 940 -466 941 -464
rect 940 -472 941 -470
rect 947 -466 948 -464
rect 947 -472 948 -470
rect 954 -466 955 -464
rect 954 -472 955 -470
rect 961 -466 962 -464
rect 961 -472 962 -470
rect 968 -466 969 -464
rect 968 -472 969 -470
rect 975 -466 976 -464
rect 975 -472 976 -470
rect 982 -466 983 -464
rect 989 -466 990 -464
rect 989 -472 990 -470
rect 996 -466 997 -464
rect 996 -472 997 -470
rect 1003 -466 1004 -464
rect 1003 -472 1004 -470
rect 1010 -466 1011 -464
rect 1010 -472 1011 -470
rect 1017 -466 1018 -464
rect 1017 -472 1018 -470
rect 1024 -466 1025 -464
rect 1024 -472 1025 -470
rect 1031 -466 1032 -464
rect 1031 -472 1032 -470
rect 1038 -466 1039 -464
rect 1038 -472 1039 -470
rect 1045 -466 1046 -464
rect 1045 -472 1046 -470
rect 1052 -466 1053 -464
rect 1052 -472 1053 -470
rect 1059 -466 1060 -464
rect 1059 -472 1060 -470
rect 1066 -466 1067 -464
rect 1066 -472 1067 -470
rect 1073 -466 1074 -464
rect 1073 -472 1074 -470
rect 1080 -466 1081 -464
rect 1080 -472 1081 -470
rect 1087 -466 1088 -464
rect 1087 -472 1088 -470
rect 1094 -466 1095 -464
rect 1094 -472 1095 -470
rect 1101 -466 1102 -464
rect 1101 -472 1102 -470
rect 1108 -466 1109 -464
rect 1108 -472 1109 -470
rect 1115 -466 1116 -464
rect 1115 -472 1116 -470
rect 1122 -466 1123 -464
rect 1122 -472 1123 -470
rect 1129 -466 1130 -464
rect 1129 -472 1130 -470
rect 1139 -466 1140 -464
rect 1139 -472 1140 -470
rect 1143 -472 1144 -470
rect 1150 -466 1151 -464
rect 1150 -472 1151 -470
rect 2 -567 3 -565
rect 9 -561 10 -559
rect 9 -567 10 -565
rect 16 -561 17 -559
rect 16 -567 17 -565
rect 23 -561 24 -559
rect 23 -567 24 -565
rect 33 -561 34 -559
rect 30 -567 31 -565
rect 33 -567 34 -565
rect 37 -561 38 -559
rect 37 -567 38 -565
rect 44 -561 45 -559
rect 44 -567 45 -565
rect 51 -561 52 -559
rect 51 -567 52 -565
rect 58 -561 59 -559
rect 58 -567 59 -565
rect 65 -561 66 -559
rect 65 -567 66 -565
rect 72 -567 73 -565
rect 75 -567 76 -565
rect 79 -567 80 -565
rect 82 -567 83 -565
rect 86 -561 87 -559
rect 86 -567 87 -565
rect 93 -561 94 -559
rect 93 -567 94 -565
rect 100 -561 101 -559
rect 100 -567 101 -565
rect 107 -561 108 -559
rect 110 -561 111 -559
rect 107 -567 108 -565
rect 114 -561 115 -559
rect 114 -567 115 -565
rect 121 -561 122 -559
rect 121 -567 122 -565
rect 128 -561 129 -559
rect 128 -567 129 -565
rect 135 -561 136 -559
rect 135 -567 136 -565
rect 142 -561 143 -559
rect 142 -567 143 -565
rect 152 -561 153 -559
rect 152 -567 153 -565
rect 156 -561 157 -559
rect 156 -567 157 -565
rect 166 -561 167 -559
rect 163 -567 164 -565
rect 166 -567 167 -565
rect 170 -561 171 -559
rect 170 -567 171 -565
rect 177 -561 178 -559
rect 177 -567 178 -565
rect 184 -561 185 -559
rect 184 -567 185 -565
rect 191 -561 192 -559
rect 194 -561 195 -559
rect 198 -561 199 -559
rect 201 -561 202 -559
rect 201 -567 202 -565
rect 205 -561 206 -559
rect 205 -567 206 -565
rect 215 -561 216 -559
rect 212 -567 213 -565
rect 219 -561 220 -559
rect 219 -567 220 -565
rect 226 -561 227 -559
rect 226 -567 227 -565
rect 233 -561 234 -559
rect 233 -567 234 -565
rect 240 -561 241 -559
rect 240 -567 241 -565
rect 247 -561 248 -559
rect 247 -567 248 -565
rect 254 -561 255 -559
rect 254 -567 255 -565
rect 261 -561 262 -559
rect 261 -567 262 -565
rect 268 -561 269 -559
rect 268 -567 269 -565
rect 275 -561 276 -559
rect 275 -567 276 -565
rect 282 -561 283 -559
rect 282 -567 283 -565
rect 289 -561 290 -559
rect 289 -567 290 -565
rect 296 -561 297 -559
rect 296 -567 297 -565
rect 303 -561 304 -559
rect 303 -567 304 -565
rect 310 -561 311 -559
rect 310 -567 311 -565
rect 317 -561 318 -559
rect 320 -561 321 -559
rect 317 -567 318 -565
rect 320 -567 321 -565
rect 324 -561 325 -559
rect 324 -567 325 -565
rect 331 -561 332 -559
rect 331 -567 332 -565
rect 338 -561 339 -559
rect 338 -567 339 -565
rect 345 -561 346 -559
rect 345 -567 346 -565
rect 355 -561 356 -559
rect 352 -567 353 -565
rect 355 -567 356 -565
rect 359 -561 360 -559
rect 359 -567 360 -565
rect 366 -567 367 -565
rect 373 -561 374 -559
rect 373 -567 374 -565
rect 380 -561 381 -559
rect 380 -567 381 -565
rect 390 -561 391 -559
rect 390 -567 391 -565
rect 397 -561 398 -559
rect 397 -567 398 -565
rect 401 -561 402 -559
rect 401 -567 402 -565
rect 408 -561 409 -559
rect 408 -567 409 -565
rect 411 -567 412 -565
rect 415 -561 416 -559
rect 415 -567 416 -565
rect 422 -561 423 -559
rect 422 -567 423 -565
rect 429 -561 430 -559
rect 429 -567 430 -565
rect 436 -561 437 -559
rect 436 -567 437 -565
rect 443 -561 444 -559
rect 443 -567 444 -565
rect 450 -561 451 -559
rect 450 -567 451 -565
rect 457 -561 458 -559
rect 457 -567 458 -565
rect 464 -561 465 -559
rect 464 -567 465 -565
rect 471 -561 472 -559
rect 471 -567 472 -565
rect 478 -561 479 -559
rect 478 -567 479 -565
rect 485 -561 486 -559
rect 485 -567 486 -565
rect 492 -561 493 -559
rect 492 -567 493 -565
rect 499 -561 500 -559
rect 499 -567 500 -565
rect 506 -561 507 -559
rect 509 -561 510 -559
rect 506 -567 507 -565
rect 509 -567 510 -565
rect 513 -561 514 -559
rect 513 -567 514 -565
rect 520 -561 521 -559
rect 520 -567 521 -565
rect 527 -561 528 -559
rect 527 -567 528 -565
rect 537 -561 538 -559
rect 537 -567 538 -565
rect 541 -561 542 -559
rect 541 -567 542 -565
rect 548 -561 549 -559
rect 551 -561 552 -559
rect 548 -567 549 -565
rect 551 -567 552 -565
rect 555 -561 556 -559
rect 555 -567 556 -565
rect 562 -561 563 -559
rect 565 -561 566 -559
rect 562 -567 563 -565
rect 569 -561 570 -559
rect 572 -561 573 -559
rect 569 -567 570 -565
rect 572 -567 573 -565
rect 576 -561 577 -559
rect 576 -567 577 -565
rect 583 -561 584 -559
rect 583 -567 584 -565
rect 593 -561 594 -559
rect 590 -567 591 -565
rect 597 -561 598 -559
rect 600 -567 601 -565
rect 604 -561 605 -559
rect 604 -567 605 -565
rect 607 -567 608 -565
rect 611 -561 612 -559
rect 611 -567 612 -565
rect 618 -561 619 -559
rect 618 -567 619 -565
rect 628 -561 629 -559
rect 628 -567 629 -565
rect 632 -561 633 -559
rect 632 -567 633 -565
rect 639 -561 640 -559
rect 639 -567 640 -565
rect 646 -561 647 -559
rect 646 -567 647 -565
rect 653 -561 654 -559
rect 653 -567 654 -565
rect 660 -561 661 -559
rect 663 -561 664 -559
rect 660 -567 661 -565
rect 663 -567 664 -565
rect 667 -561 668 -559
rect 667 -567 668 -565
rect 674 -561 675 -559
rect 674 -567 675 -565
rect 681 -561 682 -559
rect 681 -567 682 -565
rect 688 -561 689 -559
rect 688 -567 689 -565
rect 695 -561 696 -559
rect 695 -567 696 -565
rect 702 -561 703 -559
rect 702 -567 703 -565
rect 709 -561 710 -559
rect 712 -567 713 -565
rect 716 -561 717 -559
rect 716 -567 717 -565
rect 723 -561 724 -559
rect 723 -567 724 -565
rect 730 -561 731 -559
rect 733 -561 734 -559
rect 733 -567 734 -565
rect 737 -561 738 -559
rect 737 -567 738 -565
rect 744 -561 745 -559
rect 744 -567 745 -565
rect 751 -561 752 -559
rect 751 -567 752 -565
rect 758 -561 759 -559
rect 758 -567 759 -565
rect 765 -561 766 -559
rect 765 -567 766 -565
rect 772 -561 773 -559
rect 772 -567 773 -565
rect 779 -561 780 -559
rect 779 -567 780 -565
rect 786 -561 787 -559
rect 786 -567 787 -565
rect 793 -561 794 -559
rect 793 -567 794 -565
rect 800 -561 801 -559
rect 800 -567 801 -565
rect 807 -561 808 -559
rect 807 -567 808 -565
rect 814 -561 815 -559
rect 814 -567 815 -565
rect 821 -561 822 -559
rect 821 -567 822 -565
rect 828 -561 829 -559
rect 828 -567 829 -565
rect 835 -561 836 -559
rect 835 -567 836 -565
rect 842 -561 843 -559
rect 842 -567 843 -565
rect 849 -561 850 -559
rect 849 -567 850 -565
rect 856 -561 857 -559
rect 856 -567 857 -565
rect 863 -561 864 -559
rect 863 -567 864 -565
rect 870 -561 871 -559
rect 870 -567 871 -565
rect 877 -561 878 -559
rect 877 -567 878 -565
rect 884 -561 885 -559
rect 884 -567 885 -565
rect 891 -561 892 -559
rect 891 -567 892 -565
rect 898 -561 899 -559
rect 898 -567 899 -565
rect 905 -561 906 -559
rect 905 -567 906 -565
rect 912 -561 913 -559
rect 912 -567 913 -565
rect 919 -561 920 -559
rect 919 -567 920 -565
rect 926 -561 927 -559
rect 926 -567 927 -565
rect 933 -561 934 -559
rect 933 -567 934 -565
rect 940 -561 941 -559
rect 940 -567 941 -565
rect 947 -561 948 -559
rect 947 -567 948 -565
rect 954 -561 955 -559
rect 954 -567 955 -565
rect 961 -561 962 -559
rect 961 -567 962 -565
rect 968 -561 969 -559
rect 968 -567 969 -565
rect 975 -561 976 -559
rect 975 -567 976 -565
rect 982 -561 983 -559
rect 982 -567 983 -565
rect 989 -561 990 -559
rect 989 -567 990 -565
rect 996 -561 997 -559
rect 996 -567 997 -565
rect 1003 -561 1004 -559
rect 1003 -567 1004 -565
rect 1010 -561 1011 -559
rect 1010 -567 1011 -565
rect 1017 -561 1018 -559
rect 1017 -567 1018 -565
rect 1024 -561 1025 -559
rect 1024 -567 1025 -565
rect 1031 -561 1032 -559
rect 1031 -567 1032 -565
rect 1038 -561 1039 -559
rect 1038 -567 1039 -565
rect 1045 -561 1046 -559
rect 1045 -567 1046 -565
rect 1052 -561 1053 -559
rect 1052 -567 1053 -565
rect 1059 -561 1060 -559
rect 1059 -567 1060 -565
rect 1066 -561 1067 -559
rect 1066 -567 1067 -565
rect 1073 -561 1074 -559
rect 1073 -567 1074 -565
rect 1080 -561 1081 -559
rect 1080 -567 1081 -565
rect 1087 -561 1088 -559
rect 1087 -567 1088 -565
rect 1094 -561 1095 -559
rect 1094 -567 1095 -565
rect 1101 -561 1102 -559
rect 1101 -567 1102 -565
rect 1115 -561 1116 -559
rect 1115 -567 1116 -565
rect 1122 -561 1123 -559
rect 1122 -567 1123 -565
rect 1174 -561 1175 -559
rect 1178 -561 1179 -559
rect 1178 -567 1179 -565
rect 9 -652 10 -650
rect 9 -658 10 -656
rect 16 -652 17 -650
rect 16 -658 17 -656
rect 23 -652 24 -650
rect 30 -652 31 -650
rect 30 -658 31 -656
rect 37 -652 38 -650
rect 37 -658 38 -656
rect 44 -652 45 -650
rect 44 -658 45 -656
rect 54 -652 55 -650
rect 54 -658 55 -656
rect 58 -652 59 -650
rect 58 -658 59 -656
rect 68 -652 69 -650
rect 65 -658 66 -656
rect 72 -652 73 -650
rect 72 -658 73 -656
rect 79 -652 80 -650
rect 79 -658 80 -656
rect 82 -658 83 -656
rect 86 -652 87 -650
rect 89 -658 90 -656
rect 93 -652 94 -650
rect 93 -658 94 -656
rect 100 -652 101 -650
rect 103 -658 104 -656
rect 107 -652 108 -650
rect 107 -658 108 -656
rect 117 -652 118 -650
rect 117 -658 118 -656
rect 121 -652 122 -650
rect 121 -658 122 -656
rect 131 -658 132 -656
rect 135 -652 136 -650
rect 135 -658 136 -656
rect 142 -652 143 -650
rect 142 -658 143 -656
rect 149 -652 150 -650
rect 149 -658 150 -656
rect 156 -658 157 -656
rect 159 -658 160 -656
rect 163 -652 164 -650
rect 163 -658 164 -656
rect 170 -652 171 -650
rect 170 -658 171 -656
rect 177 -652 178 -650
rect 177 -658 178 -656
rect 184 -652 185 -650
rect 187 -652 188 -650
rect 184 -658 185 -656
rect 187 -658 188 -656
rect 191 -652 192 -650
rect 191 -658 192 -656
rect 198 -652 199 -650
rect 198 -658 199 -656
rect 205 -652 206 -650
rect 205 -658 206 -656
rect 212 -652 213 -650
rect 212 -658 213 -656
rect 219 -652 220 -650
rect 219 -658 220 -656
rect 226 -652 227 -650
rect 226 -658 227 -656
rect 233 -658 234 -656
rect 236 -658 237 -656
rect 240 -652 241 -650
rect 240 -658 241 -656
rect 247 -652 248 -650
rect 254 -652 255 -650
rect 254 -658 255 -656
rect 261 -652 262 -650
rect 261 -658 262 -656
rect 268 -652 269 -650
rect 268 -658 269 -656
rect 275 -652 276 -650
rect 275 -658 276 -656
rect 282 -652 283 -650
rect 282 -658 283 -656
rect 289 -652 290 -650
rect 289 -658 290 -656
rect 296 -652 297 -650
rect 296 -658 297 -656
rect 303 -652 304 -650
rect 303 -658 304 -656
rect 310 -652 311 -650
rect 310 -658 311 -656
rect 317 -652 318 -650
rect 317 -658 318 -656
rect 324 -652 325 -650
rect 324 -658 325 -656
rect 331 -652 332 -650
rect 341 -652 342 -650
rect 338 -658 339 -656
rect 345 -652 346 -650
rect 348 -652 349 -650
rect 345 -658 346 -656
rect 352 -652 353 -650
rect 352 -658 353 -656
rect 359 -652 360 -650
rect 359 -658 360 -656
rect 366 -652 367 -650
rect 366 -658 367 -656
rect 373 -652 374 -650
rect 373 -658 374 -656
rect 380 -652 381 -650
rect 380 -658 381 -656
rect 387 -652 388 -650
rect 387 -658 388 -656
rect 394 -652 395 -650
rect 394 -658 395 -656
rect 401 -652 402 -650
rect 401 -658 402 -656
rect 408 -652 409 -650
rect 408 -658 409 -656
rect 418 -652 419 -650
rect 418 -658 419 -656
rect 422 -652 423 -650
rect 422 -658 423 -656
rect 429 -652 430 -650
rect 429 -658 430 -656
rect 436 -652 437 -650
rect 436 -658 437 -656
rect 446 -652 447 -650
rect 443 -658 444 -656
rect 446 -658 447 -656
rect 450 -652 451 -650
rect 450 -658 451 -656
rect 457 -652 458 -650
rect 457 -658 458 -656
rect 464 -652 465 -650
rect 464 -658 465 -656
rect 471 -652 472 -650
rect 471 -658 472 -656
rect 481 -652 482 -650
rect 478 -658 479 -656
rect 481 -658 482 -656
rect 485 -652 486 -650
rect 485 -658 486 -656
rect 492 -652 493 -650
rect 492 -658 493 -656
rect 502 -652 503 -650
rect 499 -658 500 -656
rect 502 -658 503 -656
rect 506 -652 507 -650
rect 506 -658 507 -656
rect 513 -652 514 -650
rect 513 -658 514 -656
rect 516 -658 517 -656
rect 520 -658 521 -656
rect 523 -658 524 -656
rect 527 -652 528 -650
rect 527 -658 528 -656
rect 534 -652 535 -650
rect 534 -658 535 -656
rect 541 -652 542 -650
rect 541 -658 542 -656
rect 548 -652 549 -650
rect 551 -658 552 -656
rect 555 -652 556 -650
rect 555 -658 556 -656
rect 562 -652 563 -650
rect 562 -658 563 -656
rect 569 -652 570 -650
rect 569 -658 570 -656
rect 576 -652 577 -650
rect 576 -658 577 -656
rect 583 -652 584 -650
rect 583 -658 584 -656
rect 590 -652 591 -650
rect 590 -658 591 -656
rect 597 -652 598 -650
rect 597 -658 598 -656
rect 604 -652 605 -650
rect 607 -652 608 -650
rect 604 -658 605 -656
rect 607 -658 608 -656
rect 611 -652 612 -650
rect 614 -652 615 -650
rect 614 -658 615 -656
rect 618 -652 619 -650
rect 618 -658 619 -656
rect 625 -652 626 -650
rect 625 -658 626 -656
rect 632 -652 633 -650
rect 632 -658 633 -656
rect 639 -652 640 -650
rect 639 -658 640 -656
rect 646 -652 647 -650
rect 646 -658 647 -656
rect 653 -652 654 -650
rect 656 -652 657 -650
rect 656 -658 657 -656
rect 660 -652 661 -650
rect 660 -658 661 -656
rect 667 -652 668 -650
rect 667 -658 668 -656
rect 674 -652 675 -650
rect 674 -658 675 -656
rect 681 -652 682 -650
rect 681 -658 682 -656
rect 691 -652 692 -650
rect 688 -658 689 -656
rect 691 -658 692 -656
rect 695 -652 696 -650
rect 695 -658 696 -656
rect 702 -652 703 -650
rect 702 -658 703 -656
rect 709 -652 710 -650
rect 709 -658 710 -656
rect 716 -652 717 -650
rect 716 -658 717 -656
rect 723 -652 724 -650
rect 723 -658 724 -656
rect 730 -652 731 -650
rect 730 -658 731 -656
rect 737 -652 738 -650
rect 737 -658 738 -656
rect 744 -652 745 -650
rect 744 -658 745 -656
rect 751 -652 752 -650
rect 751 -658 752 -656
rect 758 -652 759 -650
rect 761 -652 762 -650
rect 765 -652 766 -650
rect 765 -658 766 -656
rect 772 -652 773 -650
rect 772 -658 773 -656
rect 779 -652 780 -650
rect 779 -658 780 -656
rect 786 -652 787 -650
rect 786 -658 787 -656
rect 793 -652 794 -650
rect 793 -658 794 -656
rect 800 -652 801 -650
rect 800 -658 801 -656
rect 807 -652 808 -650
rect 807 -658 808 -656
rect 814 -652 815 -650
rect 814 -658 815 -656
rect 821 -652 822 -650
rect 821 -658 822 -656
rect 828 -652 829 -650
rect 828 -658 829 -656
rect 835 -652 836 -650
rect 835 -658 836 -656
rect 842 -652 843 -650
rect 842 -658 843 -656
rect 849 -652 850 -650
rect 849 -658 850 -656
rect 856 -652 857 -650
rect 856 -658 857 -656
rect 863 -652 864 -650
rect 863 -658 864 -656
rect 870 -652 871 -650
rect 870 -658 871 -656
rect 877 -652 878 -650
rect 884 -652 885 -650
rect 884 -658 885 -656
rect 891 -652 892 -650
rect 891 -658 892 -656
rect 898 -652 899 -650
rect 898 -658 899 -656
rect 905 -652 906 -650
rect 905 -658 906 -656
rect 912 -652 913 -650
rect 912 -658 913 -656
rect 919 -652 920 -650
rect 919 -658 920 -656
rect 926 -652 927 -650
rect 926 -658 927 -656
rect 933 -658 934 -656
rect 940 -652 941 -650
rect 940 -658 941 -656
rect 947 -652 948 -650
rect 947 -658 948 -656
rect 954 -652 955 -650
rect 954 -658 955 -656
rect 961 -652 962 -650
rect 961 -658 962 -656
rect 968 -652 969 -650
rect 968 -658 969 -656
rect 975 -652 976 -650
rect 975 -658 976 -656
rect 982 -652 983 -650
rect 982 -658 983 -656
rect 989 -652 990 -650
rect 989 -658 990 -656
rect 996 -652 997 -650
rect 996 -658 997 -656
rect 1003 -652 1004 -650
rect 1003 -658 1004 -656
rect 1006 -658 1007 -656
rect 1010 -652 1011 -650
rect 1010 -658 1011 -656
rect 1017 -652 1018 -650
rect 1017 -658 1018 -656
rect 1024 -652 1025 -650
rect 1024 -658 1025 -656
rect 1031 -652 1032 -650
rect 1031 -658 1032 -656
rect 1038 -652 1039 -650
rect 1038 -658 1039 -656
rect 1041 -658 1042 -656
rect 1045 -652 1046 -650
rect 1045 -658 1046 -656
rect 1052 -652 1053 -650
rect 1052 -658 1053 -656
rect 1059 -652 1060 -650
rect 1059 -658 1060 -656
rect 1066 -652 1067 -650
rect 1066 -658 1067 -656
rect 1073 -652 1074 -650
rect 1073 -658 1074 -656
rect 1080 -652 1081 -650
rect 1080 -658 1081 -656
rect 1087 -652 1088 -650
rect 1087 -658 1088 -656
rect 1094 -652 1095 -650
rect 1094 -658 1095 -656
rect 1101 -652 1102 -650
rect 1101 -658 1102 -656
rect 1108 -652 1109 -650
rect 1108 -658 1109 -656
rect 1115 -652 1116 -650
rect 1115 -658 1116 -656
rect 1122 -652 1123 -650
rect 1122 -658 1123 -656
rect 1129 -652 1130 -650
rect 1129 -658 1130 -656
rect 1136 -652 1137 -650
rect 1136 -658 1137 -656
rect 1178 -652 1179 -650
rect 1178 -658 1179 -656
rect 9 -733 10 -731
rect 9 -739 10 -737
rect 16 -733 17 -731
rect 16 -739 17 -737
rect 23 -733 24 -731
rect 23 -739 24 -737
rect 33 -733 34 -731
rect 37 -733 38 -731
rect 37 -739 38 -737
rect 44 -733 45 -731
rect 44 -739 45 -737
rect 51 -733 52 -731
rect 51 -739 52 -737
rect 58 -733 59 -731
rect 58 -739 59 -737
rect 65 -733 66 -731
rect 65 -739 66 -737
rect 72 -733 73 -731
rect 79 -733 80 -731
rect 79 -739 80 -737
rect 86 -733 87 -731
rect 86 -739 87 -737
rect 93 -733 94 -731
rect 93 -739 94 -737
rect 100 -733 101 -731
rect 100 -739 101 -737
rect 107 -733 108 -731
rect 107 -739 108 -737
rect 114 -733 115 -731
rect 114 -739 115 -737
rect 124 -739 125 -737
rect 128 -733 129 -731
rect 128 -739 129 -737
rect 135 -733 136 -731
rect 135 -739 136 -737
rect 138 -739 139 -737
rect 142 -733 143 -731
rect 142 -739 143 -737
rect 149 -733 150 -731
rect 152 -733 153 -731
rect 156 -733 157 -731
rect 156 -739 157 -737
rect 163 -733 164 -731
rect 163 -739 164 -737
rect 170 -733 171 -731
rect 170 -739 171 -737
rect 177 -733 178 -731
rect 177 -739 178 -737
rect 184 -733 185 -731
rect 187 -739 188 -737
rect 191 -733 192 -731
rect 191 -739 192 -737
rect 198 -733 199 -731
rect 198 -739 199 -737
rect 205 -733 206 -731
rect 208 -733 209 -731
rect 212 -733 213 -731
rect 212 -739 213 -737
rect 219 -733 220 -731
rect 219 -739 220 -737
rect 226 -733 227 -731
rect 226 -739 227 -737
rect 233 -733 234 -731
rect 233 -739 234 -737
rect 240 -733 241 -731
rect 240 -739 241 -737
rect 247 -739 248 -737
rect 254 -733 255 -731
rect 254 -739 255 -737
rect 261 -733 262 -731
rect 261 -739 262 -737
rect 268 -733 269 -731
rect 268 -739 269 -737
rect 275 -733 276 -731
rect 275 -739 276 -737
rect 282 -733 283 -731
rect 282 -739 283 -737
rect 289 -733 290 -731
rect 289 -739 290 -737
rect 296 -733 297 -731
rect 296 -739 297 -737
rect 303 -733 304 -731
rect 303 -739 304 -737
rect 310 -739 311 -737
rect 317 -733 318 -731
rect 317 -739 318 -737
rect 324 -733 325 -731
rect 324 -739 325 -737
rect 331 -733 332 -731
rect 331 -739 332 -737
rect 338 -733 339 -731
rect 341 -733 342 -731
rect 338 -739 339 -737
rect 341 -739 342 -737
rect 345 -733 346 -731
rect 345 -739 346 -737
rect 352 -733 353 -731
rect 352 -739 353 -737
rect 359 -739 360 -737
rect 362 -739 363 -737
rect 366 -733 367 -731
rect 366 -739 367 -737
rect 373 -733 374 -731
rect 373 -739 374 -737
rect 380 -733 381 -731
rect 380 -739 381 -737
rect 387 -733 388 -731
rect 387 -739 388 -737
rect 394 -733 395 -731
rect 397 -733 398 -731
rect 394 -739 395 -737
rect 404 -739 405 -737
rect 411 -733 412 -731
rect 411 -739 412 -737
rect 415 -733 416 -731
rect 415 -739 416 -737
rect 425 -733 426 -731
rect 425 -739 426 -737
rect 429 -733 430 -731
rect 429 -739 430 -737
rect 439 -733 440 -731
rect 439 -739 440 -737
rect 443 -733 444 -731
rect 443 -739 444 -737
rect 450 -733 451 -731
rect 450 -739 451 -737
rect 457 -733 458 -731
rect 457 -739 458 -737
rect 464 -733 465 -731
rect 467 -733 468 -731
rect 474 -733 475 -731
rect 474 -739 475 -737
rect 478 -733 479 -731
rect 478 -739 479 -737
rect 485 -733 486 -731
rect 485 -739 486 -737
rect 492 -733 493 -731
rect 492 -739 493 -737
rect 499 -733 500 -731
rect 499 -739 500 -737
rect 506 -733 507 -731
rect 506 -739 507 -737
rect 513 -733 514 -731
rect 513 -739 514 -737
rect 523 -733 524 -731
rect 520 -739 521 -737
rect 523 -739 524 -737
rect 527 -733 528 -731
rect 527 -739 528 -737
rect 534 -733 535 -731
rect 534 -739 535 -737
rect 541 -733 542 -731
rect 541 -739 542 -737
rect 548 -733 549 -731
rect 551 -733 552 -731
rect 548 -739 549 -737
rect 555 -733 556 -731
rect 555 -739 556 -737
rect 562 -733 563 -731
rect 562 -739 563 -737
rect 569 -733 570 -731
rect 569 -739 570 -737
rect 576 -733 577 -731
rect 576 -739 577 -737
rect 583 -733 584 -731
rect 583 -739 584 -737
rect 590 -733 591 -731
rect 590 -739 591 -737
rect 597 -733 598 -731
rect 597 -739 598 -737
rect 600 -739 601 -737
rect 604 -733 605 -731
rect 604 -739 605 -737
rect 611 -733 612 -731
rect 611 -739 612 -737
rect 618 -733 619 -731
rect 618 -739 619 -737
rect 625 -733 626 -731
rect 625 -739 626 -737
rect 635 -733 636 -731
rect 632 -739 633 -737
rect 635 -739 636 -737
rect 639 -733 640 -731
rect 642 -739 643 -737
rect 646 -733 647 -731
rect 646 -739 647 -737
rect 653 -733 654 -731
rect 653 -739 654 -737
rect 660 -733 661 -731
rect 660 -739 661 -737
rect 667 -733 668 -731
rect 667 -739 668 -737
rect 674 -733 675 -731
rect 674 -739 675 -737
rect 681 -733 682 -731
rect 681 -739 682 -737
rect 688 -733 689 -731
rect 691 -733 692 -731
rect 688 -739 689 -737
rect 695 -733 696 -731
rect 695 -739 696 -737
rect 702 -733 703 -731
rect 702 -739 703 -737
rect 709 -733 710 -731
rect 709 -739 710 -737
rect 716 -733 717 -731
rect 716 -739 717 -737
rect 723 -733 724 -731
rect 723 -739 724 -737
rect 730 -733 731 -731
rect 730 -739 731 -737
rect 737 -733 738 -731
rect 737 -739 738 -737
rect 744 -733 745 -731
rect 747 -733 748 -731
rect 744 -739 745 -737
rect 747 -739 748 -737
rect 751 -733 752 -731
rect 751 -739 752 -737
rect 758 -733 759 -731
rect 758 -739 759 -737
rect 765 -733 766 -731
rect 765 -739 766 -737
rect 772 -733 773 -731
rect 772 -739 773 -737
rect 779 -733 780 -731
rect 779 -739 780 -737
rect 786 -733 787 -731
rect 786 -739 787 -737
rect 793 -733 794 -731
rect 793 -739 794 -737
rect 800 -733 801 -731
rect 800 -739 801 -737
rect 807 -733 808 -731
rect 807 -739 808 -737
rect 814 -733 815 -731
rect 814 -739 815 -737
rect 821 -733 822 -731
rect 821 -739 822 -737
rect 828 -733 829 -731
rect 828 -739 829 -737
rect 835 -733 836 -731
rect 835 -739 836 -737
rect 842 -733 843 -731
rect 842 -739 843 -737
rect 849 -733 850 -731
rect 849 -739 850 -737
rect 856 -733 857 -731
rect 856 -739 857 -737
rect 863 -733 864 -731
rect 863 -739 864 -737
rect 870 -733 871 -731
rect 870 -739 871 -737
rect 877 -739 878 -737
rect 884 -733 885 -731
rect 884 -739 885 -737
rect 891 -733 892 -731
rect 891 -739 892 -737
rect 898 -733 899 -731
rect 898 -739 899 -737
rect 905 -733 906 -731
rect 905 -739 906 -737
rect 912 -733 913 -731
rect 912 -739 913 -737
rect 919 -733 920 -731
rect 919 -739 920 -737
rect 926 -733 927 -731
rect 926 -739 927 -737
rect 933 -733 934 -731
rect 933 -739 934 -737
rect 940 -733 941 -731
rect 940 -739 941 -737
rect 947 -733 948 -731
rect 947 -739 948 -737
rect 954 -733 955 -731
rect 954 -739 955 -737
rect 961 -733 962 -731
rect 961 -739 962 -737
rect 968 -733 969 -731
rect 968 -739 969 -737
rect 975 -733 976 -731
rect 975 -739 976 -737
rect 982 -733 983 -731
rect 982 -739 983 -737
rect 989 -733 990 -731
rect 989 -739 990 -737
rect 996 -733 997 -731
rect 996 -739 997 -737
rect 1003 -733 1004 -731
rect 1006 -733 1007 -731
rect 1003 -739 1004 -737
rect 1010 -733 1011 -731
rect 1010 -739 1011 -737
rect 1017 -733 1018 -731
rect 1017 -739 1018 -737
rect 1024 -733 1025 -731
rect 1024 -739 1025 -737
rect 1031 -733 1032 -731
rect 1031 -739 1032 -737
rect 1038 -733 1039 -731
rect 1041 -733 1042 -731
rect 1038 -739 1039 -737
rect 1045 -733 1046 -731
rect 1045 -739 1046 -737
rect 1052 -733 1053 -731
rect 1052 -739 1053 -737
rect 1059 -733 1060 -731
rect 1059 -739 1060 -737
rect 1066 -733 1067 -731
rect 1066 -739 1067 -737
rect 1073 -733 1074 -731
rect 1073 -739 1074 -737
rect 1080 -733 1081 -731
rect 1080 -739 1081 -737
rect 1087 -733 1088 -731
rect 1090 -733 1091 -731
rect 1087 -739 1088 -737
rect 1090 -739 1091 -737
rect 1094 -733 1095 -731
rect 1094 -739 1095 -737
rect 1101 -733 1102 -731
rect 1101 -739 1102 -737
rect 1108 -733 1109 -731
rect 1111 -733 1112 -731
rect 1108 -739 1109 -737
rect 1115 -733 1116 -731
rect 1115 -739 1116 -737
rect 1122 -733 1123 -731
rect 1122 -739 1123 -737
rect 1129 -733 1130 -731
rect 1129 -739 1130 -737
rect 1136 -733 1137 -731
rect 1136 -739 1137 -737
rect 1143 -733 1144 -731
rect 1143 -739 1144 -737
rect 1150 -733 1151 -731
rect 1150 -739 1151 -737
rect 1157 -739 1158 -737
rect 1160 -739 1161 -737
rect 1164 -733 1165 -731
rect 1164 -739 1165 -737
rect 1171 -733 1172 -731
rect 1171 -739 1172 -737
rect 1185 -733 1186 -731
rect 1185 -739 1186 -737
rect 9 -822 10 -820
rect 9 -828 10 -826
rect 16 -822 17 -820
rect 16 -828 17 -826
rect 23 -822 24 -820
rect 23 -828 24 -826
rect 30 -822 31 -820
rect 30 -828 31 -826
rect 37 -822 38 -820
rect 37 -828 38 -826
rect 44 -822 45 -820
rect 44 -828 45 -826
rect 51 -822 52 -820
rect 51 -828 52 -826
rect 58 -822 59 -820
rect 58 -828 59 -826
rect 65 -822 66 -820
rect 65 -828 66 -826
rect 72 -828 73 -826
rect 79 -822 80 -820
rect 79 -828 80 -826
rect 86 -822 87 -820
rect 86 -828 87 -826
rect 93 -822 94 -820
rect 93 -828 94 -826
rect 100 -822 101 -820
rect 107 -822 108 -820
rect 107 -828 108 -826
rect 117 -822 118 -820
rect 114 -828 115 -826
rect 117 -828 118 -826
rect 121 -822 122 -820
rect 121 -828 122 -826
rect 124 -828 125 -826
rect 131 -822 132 -820
rect 128 -828 129 -826
rect 135 -822 136 -820
rect 138 -822 139 -820
rect 142 -822 143 -820
rect 142 -828 143 -826
rect 149 -822 150 -820
rect 149 -828 150 -826
rect 156 -822 157 -820
rect 156 -828 157 -826
rect 163 -822 164 -820
rect 163 -828 164 -826
rect 170 -822 171 -820
rect 173 -822 174 -820
rect 177 -822 178 -820
rect 177 -828 178 -826
rect 184 -822 185 -820
rect 184 -828 185 -826
rect 191 -822 192 -820
rect 191 -828 192 -826
rect 198 -822 199 -820
rect 198 -828 199 -826
rect 205 -822 206 -820
rect 205 -828 206 -826
rect 212 -822 213 -820
rect 212 -828 213 -826
rect 219 -822 220 -820
rect 219 -828 220 -826
rect 226 -822 227 -820
rect 226 -828 227 -826
rect 233 -822 234 -820
rect 233 -828 234 -826
rect 240 -822 241 -820
rect 240 -828 241 -826
rect 247 -822 248 -820
rect 247 -828 248 -826
rect 254 -822 255 -820
rect 254 -828 255 -826
rect 268 -822 269 -820
rect 268 -828 269 -826
rect 275 -822 276 -820
rect 275 -828 276 -826
rect 282 -822 283 -820
rect 282 -828 283 -826
rect 289 -822 290 -820
rect 289 -828 290 -826
rect 296 -822 297 -820
rect 296 -828 297 -826
rect 303 -822 304 -820
rect 303 -828 304 -826
rect 310 -822 311 -820
rect 310 -828 311 -826
rect 317 -822 318 -820
rect 317 -828 318 -826
rect 324 -822 325 -820
rect 324 -828 325 -826
rect 331 -822 332 -820
rect 331 -828 332 -826
rect 338 -822 339 -820
rect 338 -828 339 -826
rect 345 -822 346 -820
rect 345 -828 346 -826
rect 352 -822 353 -820
rect 352 -828 353 -826
rect 355 -828 356 -826
rect 362 -828 363 -826
rect 366 -822 367 -820
rect 366 -828 367 -826
rect 373 -822 374 -820
rect 373 -828 374 -826
rect 380 -822 381 -820
rect 383 -822 384 -820
rect 380 -828 381 -826
rect 383 -828 384 -826
rect 387 -822 388 -820
rect 387 -828 388 -826
rect 394 -822 395 -820
rect 394 -828 395 -826
rect 401 -822 402 -820
rect 401 -828 402 -826
rect 408 -822 409 -820
rect 408 -828 409 -826
rect 415 -822 416 -820
rect 415 -828 416 -826
rect 425 -822 426 -820
rect 422 -828 423 -826
rect 425 -828 426 -826
rect 429 -822 430 -820
rect 429 -828 430 -826
rect 436 -822 437 -820
rect 436 -828 437 -826
rect 443 -822 444 -820
rect 443 -828 444 -826
rect 450 -822 451 -820
rect 450 -828 451 -826
rect 457 -822 458 -820
rect 457 -828 458 -826
rect 464 -822 465 -820
rect 464 -828 465 -826
rect 471 -822 472 -820
rect 471 -828 472 -826
rect 478 -822 479 -820
rect 485 -822 486 -820
rect 485 -828 486 -826
rect 495 -822 496 -820
rect 492 -828 493 -826
rect 495 -828 496 -826
rect 499 -822 500 -820
rect 502 -822 503 -820
rect 502 -828 503 -826
rect 506 -822 507 -820
rect 506 -828 507 -826
rect 513 -822 514 -820
rect 513 -828 514 -826
rect 520 -822 521 -820
rect 523 -828 524 -826
rect 527 -822 528 -820
rect 527 -828 528 -826
rect 534 -822 535 -820
rect 534 -828 535 -826
rect 541 -822 542 -820
rect 541 -828 542 -826
rect 548 -822 549 -820
rect 548 -828 549 -826
rect 555 -822 556 -820
rect 555 -828 556 -826
rect 558 -828 559 -826
rect 562 -822 563 -820
rect 565 -822 566 -820
rect 569 -822 570 -820
rect 572 -822 573 -820
rect 569 -828 570 -826
rect 576 -822 577 -820
rect 576 -828 577 -826
rect 583 -822 584 -820
rect 583 -828 584 -826
rect 590 -822 591 -820
rect 590 -828 591 -826
rect 597 -822 598 -820
rect 597 -828 598 -826
rect 604 -822 605 -820
rect 604 -828 605 -826
rect 611 -822 612 -820
rect 611 -828 612 -826
rect 621 -822 622 -820
rect 618 -828 619 -826
rect 621 -828 622 -826
rect 625 -822 626 -820
rect 632 -822 633 -820
rect 632 -828 633 -826
rect 639 -822 640 -820
rect 642 -822 643 -820
rect 646 -822 647 -820
rect 646 -828 647 -826
rect 656 -822 657 -820
rect 656 -828 657 -826
rect 660 -822 661 -820
rect 663 -822 664 -820
rect 663 -828 664 -826
rect 667 -822 668 -820
rect 667 -828 668 -826
rect 674 -822 675 -820
rect 674 -828 675 -826
rect 681 -822 682 -820
rect 681 -828 682 -826
rect 688 -822 689 -820
rect 688 -828 689 -826
rect 695 -822 696 -820
rect 698 -822 699 -820
rect 695 -828 696 -826
rect 698 -828 699 -826
rect 702 -822 703 -820
rect 702 -828 703 -826
rect 709 -822 710 -820
rect 709 -828 710 -826
rect 716 -822 717 -820
rect 716 -828 717 -826
rect 723 -822 724 -820
rect 726 -828 727 -826
rect 730 -822 731 -820
rect 730 -828 731 -826
rect 737 -822 738 -820
rect 737 -828 738 -826
rect 744 -822 745 -820
rect 744 -828 745 -826
rect 751 -822 752 -820
rect 751 -828 752 -826
rect 758 -822 759 -820
rect 758 -828 759 -826
rect 765 -822 766 -820
rect 765 -828 766 -826
rect 772 -822 773 -820
rect 772 -828 773 -826
rect 779 -822 780 -820
rect 782 -822 783 -820
rect 786 -822 787 -820
rect 786 -828 787 -826
rect 793 -822 794 -820
rect 793 -828 794 -826
rect 800 -822 801 -820
rect 800 -828 801 -826
rect 807 -822 808 -820
rect 807 -828 808 -826
rect 817 -822 818 -820
rect 814 -828 815 -826
rect 817 -828 818 -826
rect 821 -822 822 -820
rect 821 -828 822 -826
rect 828 -822 829 -820
rect 828 -828 829 -826
rect 835 -822 836 -820
rect 835 -828 836 -826
rect 842 -822 843 -820
rect 842 -828 843 -826
rect 849 -822 850 -820
rect 852 -822 853 -820
rect 856 -822 857 -820
rect 856 -828 857 -826
rect 863 -822 864 -820
rect 863 -828 864 -826
rect 870 -822 871 -820
rect 870 -828 871 -826
rect 877 -822 878 -820
rect 877 -828 878 -826
rect 884 -822 885 -820
rect 884 -828 885 -826
rect 891 -822 892 -820
rect 891 -828 892 -826
rect 898 -822 899 -820
rect 898 -828 899 -826
rect 905 -822 906 -820
rect 905 -828 906 -826
rect 912 -822 913 -820
rect 912 -828 913 -826
rect 919 -822 920 -820
rect 919 -828 920 -826
rect 926 -822 927 -820
rect 926 -828 927 -826
rect 933 -822 934 -820
rect 933 -828 934 -826
rect 940 -822 941 -820
rect 940 -828 941 -826
rect 947 -822 948 -820
rect 947 -828 948 -826
rect 954 -822 955 -820
rect 954 -828 955 -826
rect 961 -822 962 -820
rect 961 -828 962 -826
rect 968 -822 969 -820
rect 968 -828 969 -826
rect 975 -822 976 -820
rect 975 -828 976 -826
rect 982 -822 983 -820
rect 982 -828 983 -826
rect 989 -822 990 -820
rect 989 -828 990 -826
rect 996 -822 997 -820
rect 996 -828 997 -826
rect 999 -828 1000 -826
rect 1003 -822 1004 -820
rect 1003 -828 1004 -826
rect 1010 -822 1011 -820
rect 1010 -828 1011 -826
rect 1017 -822 1018 -820
rect 1017 -828 1018 -826
rect 1024 -822 1025 -820
rect 1024 -828 1025 -826
rect 1031 -822 1032 -820
rect 1031 -828 1032 -826
rect 1038 -822 1039 -820
rect 1038 -828 1039 -826
rect 1045 -822 1046 -820
rect 1045 -828 1046 -826
rect 1052 -822 1053 -820
rect 1052 -828 1053 -826
rect 1059 -822 1060 -820
rect 1059 -828 1060 -826
rect 1066 -822 1067 -820
rect 1066 -828 1067 -826
rect 1073 -822 1074 -820
rect 1073 -828 1074 -826
rect 1080 -822 1081 -820
rect 1080 -828 1081 -826
rect 1087 -822 1088 -820
rect 1087 -828 1088 -826
rect 1094 -822 1095 -820
rect 1094 -828 1095 -826
rect 1101 -822 1102 -820
rect 1101 -828 1102 -826
rect 1108 -822 1109 -820
rect 1108 -828 1109 -826
rect 1115 -822 1116 -820
rect 1115 -828 1116 -826
rect 1122 -822 1123 -820
rect 1122 -828 1123 -826
rect 1129 -822 1130 -820
rect 1129 -828 1130 -826
rect 1136 -822 1137 -820
rect 1136 -828 1137 -826
rect 1143 -822 1144 -820
rect 1143 -828 1144 -826
rect 1150 -822 1151 -820
rect 1150 -828 1151 -826
rect 1157 -822 1158 -820
rect 1157 -828 1158 -826
rect 1164 -822 1165 -820
rect 1164 -828 1165 -826
rect 1171 -822 1172 -820
rect 1171 -828 1172 -826
rect 1178 -822 1179 -820
rect 1178 -828 1179 -826
rect 1185 -822 1186 -820
rect 1185 -828 1186 -826
rect 1192 -822 1193 -820
rect 1192 -828 1193 -826
rect 1199 -822 1200 -820
rect 1199 -828 1200 -826
rect 1206 -822 1207 -820
rect 1206 -828 1207 -826
rect 1213 -822 1214 -820
rect 1213 -828 1214 -826
rect 1220 -822 1221 -820
rect 1220 -828 1221 -826
rect 5 -909 6 -907
rect 9 -909 10 -907
rect 9 -915 10 -913
rect 19 -909 20 -907
rect 19 -915 20 -913
rect 23 -909 24 -907
rect 23 -915 24 -913
rect 33 -909 34 -907
rect 33 -915 34 -913
rect 37 -909 38 -907
rect 40 -909 41 -907
rect 37 -915 38 -913
rect 40 -915 41 -913
rect 44 -909 45 -907
rect 44 -915 45 -913
rect 51 -909 52 -907
rect 51 -915 52 -913
rect 58 -909 59 -907
rect 58 -915 59 -913
rect 65 -909 66 -907
rect 65 -915 66 -913
rect 72 -909 73 -907
rect 72 -915 73 -913
rect 79 -909 80 -907
rect 79 -915 80 -913
rect 86 -909 87 -907
rect 86 -915 87 -913
rect 93 -909 94 -907
rect 93 -915 94 -913
rect 100 -915 101 -913
rect 107 -909 108 -907
rect 107 -915 108 -913
rect 117 -909 118 -907
rect 114 -915 115 -913
rect 117 -915 118 -913
rect 121 -909 122 -907
rect 121 -915 122 -913
rect 128 -909 129 -907
rect 128 -915 129 -913
rect 135 -909 136 -907
rect 135 -915 136 -913
rect 142 -909 143 -907
rect 142 -915 143 -913
rect 149 -909 150 -907
rect 152 -915 153 -913
rect 156 -909 157 -907
rect 156 -915 157 -913
rect 163 -909 164 -907
rect 163 -915 164 -913
rect 170 -909 171 -907
rect 170 -915 171 -913
rect 177 -909 178 -907
rect 177 -915 178 -913
rect 184 -909 185 -907
rect 184 -915 185 -913
rect 191 -909 192 -907
rect 191 -915 192 -913
rect 198 -909 199 -907
rect 198 -915 199 -913
rect 205 -909 206 -907
rect 208 -915 209 -913
rect 212 -909 213 -907
rect 212 -915 213 -913
rect 219 -909 220 -907
rect 219 -915 220 -913
rect 226 -909 227 -907
rect 226 -915 227 -913
rect 233 -909 234 -907
rect 233 -915 234 -913
rect 240 -909 241 -907
rect 240 -915 241 -913
rect 247 -909 248 -907
rect 247 -915 248 -913
rect 254 -909 255 -907
rect 254 -915 255 -913
rect 264 -909 265 -907
rect 261 -915 262 -913
rect 264 -915 265 -913
rect 268 -909 269 -907
rect 268 -915 269 -913
rect 278 -909 279 -907
rect 275 -915 276 -913
rect 282 -909 283 -907
rect 282 -915 283 -913
rect 289 -909 290 -907
rect 292 -909 293 -907
rect 289 -915 290 -913
rect 296 -909 297 -907
rect 296 -915 297 -913
rect 303 -909 304 -907
rect 303 -915 304 -913
rect 310 -909 311 -907
rect 313 -909 314 -907
rect 317 -909 318 -907
rect 317 -915 318 -913
rect 324 -909 325 -907
rect 324 -915 325 -913
rect 331 -909 332 -907
rect 331 -915 332 -913
rect 338 -909 339 -907
rect 338 -915 339 -913
rect 348 -909 349 -907
rect 348 -915 349 -913
rect 352 -909 353 -907
rect 352 -915 353 -913
rect 359 -909 360 -907
rect 359 -915 360 -913
rect 366 -909 367 -907
rect 366 -915 367 -913
rect 373 -915 374 -913
rect 380 -909 381 -907
rect 380 -915 381 -913
rect 387 -909 388 -907
rect 387 -915 388 -913
rect 394 -909 395 -907
rect 394 -915 395 -913
rect 401 -909 402 -907
rect 401 -915 402 -913
rect 408 -909 409 -907
rect 408 -915 409 -913
rect 415 -909 416 -907
rect 415 -915 416 -913
rect 425 -909 426 -907
rect 422 -915 423 -913
rect 429 -909 430 -907
rect 429 -915 430 -913
rect 436 -909 437 -907
rect 436 -915 437 -913
rect 439 -915 440 -913
rect 443 -909 444 -907
rect 443 -915 444 -913
rect 450 -909 451 -907
rect 450 -915 451 -913
rect 457 -909 458 -907
rect 457 -915 458 -913
rect 464 -909 465 -907
rect 464 -915 465 -913
rect 471 -909 472 -907
rect 471 -915 472 -913
rect 478 -909 479 -907
rect 485 -909 486 -907
rect 485 -915 486 -913
rect 492 -909 493 -907
rect 492 -915 493 -913
rect 499 -909 500 -907
rect 499 -915 500 -913
rect 506 -909 507 -907
rect 506 -915 507 -913
rect 513 -909 514 -907
rect 513 -915 514 -913
rect 520 -909 521 -907
rect 520 -915 521 -913
rect 527 -909 528 -907
rect 527 -915 528 -913
rect 534 -909 535 -907
rect 534 -915 535 -913
rect 541 -909 542 -907
rect 544 -909 545 -907
rect 548 -909 549 -907
rect 548 -915 549 -913
rect 555 -909 556 -907
rect 555 -915 556 -913
rect 558 -915 559 -913
rect 562 -909 563 -907
rect 562 -915 563 -913
rect 569 -909 570 -907
rect 569 -915 570 -913
rect 576 -909 577 -907
rect 576 -915 577 -913
rect 583 -909 584 -907
rect 583 -915 584 -913
rect 590 -909 591 -907
rect 590 -915 591 -913
rect 597 -909 598 -907
rect 600 -909 601 -907
rect 597 -915 598 -913
rect 604 -909 605 -907
rect 604 -915 605 -913
rect 611 -909 612 -907
rect 614 -909 615 -907
rect 614 -915 615 -913
rect 621 -909 622 -907
rect 625 -909 626 -907
rect 625 -915 626 -913
rect 632 -909 633 -907
rect 632 -915 633 -913
rect 639 -909 640 -907
rect 639 -915 640 -913
rect 646 -909 647 -907
rect 646 -915 647 -913
rect 653 -909 654 -907
rect 656 -909 657 -907
rect 653 -915 654 -913
rect 656 -915 657 -913
rect 660 -909 661 -907
rect 660 -915 661 -913
rect 667 -909 668 -907
rect 670 -909 671 -907
rect 674 -909 675 -907
rect 677 -909 678 -907
rect 681 -909 682 -907
rect 684 -915 685 -913
rect 688 -909 689 -907
rect 688 -915 689 -913
rect 695 -909 696 -907
rect 695 -915 696 -913
rect 702 -909 703 -907
rect 702 -915 703 -913
rect 709 -909 710 -907
rect 709 -915 710 -913
rect 716 -909 717 -907
rect 716 -915 717 -913
rect 723 -909 724 -907
rect 723 -915 724 -913
rect 730 -909 731 -907
rect 730 -915 731 -913
rect 737 -909 738 -907
rect 737 -915 738 -913
rect 744 -909 745 -907
rect 744 -915 745 -913
rect 751 -909 752 -907
rect 751 -915 752 -913
rect 758 -909 759 -907
rect 758 -915 759 -913
rect 765 -909 766 -907
rect 765 -915 766 -913
rect 772 -909 773 -907
rect 772 -915 773 -913
rect 779 -909 780 -907
rect 779 -915 780 -913
rect 786 -909 787 -907
rect 786 -915 787 -913
rect 793 -909 794 -907
rect 793 -915 794 -913
rect 800 -909 801 -907
rect 800 -915 801 -913
rect 807 -909 808 -907
rect 807 -915 808 -913
rect 814 -909 815 -907
rect 814 -915 815 -913
rect 821 -915 822 -913
rect 824 -915 825 -913
rect 828 -909 829 -907
rect 828 -915 829 -913
rect 835 -909 836 -907
rect 835 -915 836 -913
rect 842 -909 843 -907
rect 842 -915 843 -913
rect 849 -909 850 -907
rect 849 -915 850 -913
rect 856 -909 857 -907
rect 856 -915 857 -913
rect 863 -909 864 -907
rect 863 -915 864 -913
rect 870 -909 871 -907
rect 870 -915 871 -913
rect 877 -909 878 -907
rect 877 -915 878 -913
rect 884 -909 885 -907
rect 884 -915 885 -913
rect 891 -909 892 -907
rect 891 -915 892 -913
rect 898 -915 899 -913
rect 901 -915 902 -913
rect 905 -909 906 -907
rect 905 -915 906 -913
rect 912 -909 913 -907
rect 912 -915 913 -913
rect 919 -909 920 -907
rect 919 -915 920 -913
rect 926 -909 927 -907
rect 926 -915 927 -913
rect 933 -909 934 -907
rect 933 -915 934 -913
rect 940 -909 941 -907
rect 940 -915 941 -913
rect 947 -909 948 -907
rect 947 -915 948 -913
rect 954 -909 955 -907
rect 954 -915 955 -913
rect 961 -909 962 -907
rect 961 -915 962 -913
rect 968 -909 969 -907
rect 968 -915 969 -913
rect 975 -909 976 -907
rect 975 -915 976 -913
rect 982 -909 983 -907
rect 982 -915 983 -913
rect 989 -909 990 -907
rect 989 -915 990 -913
rect 996 -909 997 -907
rect 999 -909 1000 -907
rect 996 -915 997 -913
rect 1003 -909 1004 -907
rect 1003 -915 1004 -913
rect 1010 -909 1011 -907
rect 1010 -915 1011 -913
rect 1017 -909 1018 -907
rect 1017 -915 1018 -913
rect 1024 -909 1025 -907
rect 1024 -915 1025 -913
rect 1031 -909 1032 -907
rect 1031 -915 1032 -913
rect 1038 -909 1039 -907
rect 1038 -915 1039 -913
rect 1045 -909 1046 -907
rect 1045 -915 1046 -913
rect 1052 -909 1053 -907
rect 1052 -915 1053 -913
rect 1059 -909 1060 -907
rect 1059 -915 1060 -913
rect 1066 -909 1067 -907
rect 1066 -915 1067 -913
rect 1073 -909 1074 -907
rect 1073 -915 1074 -913
rect 1080 -909 1081 -907
rect 1080 -915 1081 -913
rect 1087 -909 1088 -907
rect 1090 -909 1091 -907
rect 1090 -915 1091 -913
rect 1094 -909 1095 -907
rect 1094 -915 1095 -913
rect 1101 -909 1102 -907
rect 1101 -915 1102 -913
rect 1108 -909 1109 -907
rect 1108 -915 1109 -913
rect 1115 -909 1116 -907
rect 1115 -915 1116 -913
rect 1122 -909 1123 -907
rect 1122 -915 1123 -913
rect 1129 -909 1130 -907
rect 1129 -915 1130 -913
rect 1164 -909 1165 -907
rect 1164 -915 1165 -913
rect 1171 -909 1172 -907
rect 1171 -915 1172 -913
rect 1178 -909 1179 -907
rect 1178 -915 1179 -913
rect 1192 -909 1193 -907
rect 1192 -915 1193 -913
rect 2 -998 3 -996
rect 2 -1004 3 -1002
rect 9 -998 10 -996
rect 9 -1004 10 -1002
rect 16 -1004 17 -1002
rect 23 -998 24 -996
rect 23 -1004 24 -1002
rect 30 -998 31 -996
rect 30 -1004 31 -1002
rect 40 -998 41 -996
rect 40 -1004 41 -1002
rect 44 -998 45 -996
rect 44 -1004 45 -1002
rect 51 -998 52 -996
rect 51 -1004 52 -1002
rect 58 -998 59 -996
rect 61 -998 62 -996
rect 61 -1004 62 -1002
rect 65 -998 66 -996
rect 65 -1004 66 -1002
rect 72 -998 73 -996
rect 72 -1004 73 -1002
rect 79 -998 80 -996
rect 79 -1004 80 -1002
rect 86 -998 87 -996
rect 86 -1004 87 -1002
rect 93 -998 94 -996
rect 96 -998 97 -996
rect 96 -1004 97 -1002
rect 100 -998 101 -996
rect 103 -1004 104 -1002
rect 107 -998 108 -996
rect 107 -1004 108 -1002
rect 114 -998 115 -996
rect 114 -1004 115 -1002
rect 121 -998 122 -996
rect 124 -1004 125 -1002
rect 128 -998 129 -996
rect 128 -1004 129 -1002
rect 135 -998 136 -996
rect 135 -1004 136 -1002
rect 142 -998 143 -996
rect 142 -1004 143 -1002
rect 149 -998 150 -996
rect 149 -1004 150 -1002
rect 156 -998 157 -996
rect 156 -1004 157 -1002
rect 163 -998 164 -996
rect 163 -1004 164 -1002
rect 170 -998 171 -996
rect 170 -1004 171 -1002
rect 177 -998 178 -996
rect 177 -1004 178 -1002
rect 184 -998 185 -996
rect 187 -1004 188 -1002
rect 191 -998 192 -996
rect 191 -1004 192 -1002
rect 198 -998 199 -996
rect 198 -1004 199 -1002
rect 201 -1004 202 -1002
rect 205 -998 206 -996
rect 205 -1004 206 -1002
rect 212 -998 213 -996
rect 212 -1004 213 -1002
rect 219 -998 220 -996
rect 219 -1004 220 -1002
rect 226 -998 227 -996
rect 226 -1004 227 -1002
rect 233 -998 234 -996
rect 233 -1004 234 -1002
rect 240 -998 241 -996
rect 240 -1004 241 -1002
rect 247 -998 248 -996
rect 247 -1004 248 -1002
rect 254 -998 255 -996
rect 254 -1004 255 -1002
rect 261 -998 262 -996
rect 261 -1004 262 -1002
rect 268 -998 269 -996
rect 268 -1004 269 -1002
rect 275 -998 276 -996
rect 275 -1004 276 -1002
rect 282 -998 283 -996
rect 282 -1004 283 -1002
rect 289 -998 290 -996
rect 289 -1004 290 -1002
rect 296 -998 297 -996
rect 296 -1004 297 -1002
rect 303 -998 304 -996
rect 303 -1004 304 -1002
rect 310 -998 311 -996
rect 310 -1004 311 -1002
rect 317 -998 318 -996
rect 317 -1004 318 -1002
rect 324 -998 325 -996
rect 324 -1004 325 -1002
rect 331 -998 332 -996
rect 331 -1004 332 -1002
rect 338 -998 339 -996
rect 338 -1004 339 -1002
rect 345 -998 346 -996
rect 345 -1004 346 -1002
rect 352 -998 353 -996
rect 352 -1004 353 -1002
rect 362 -998 363 -996
rect 359 -1004 360 -1002
rect 362 -1004 363 -1002
rect 366 -998 367 -996
rect 366 -1004 367 -1002
rect 376 -998 377 -996
rect 373 -1004 374 -1002
rect 376 -1004 377 -1002
rect 380 -998 381 -996
rect 380 -1004 381 -1002
rect 390 -998 391 -996
rect 390 -1004 391 -1002
rect 394 -998 395 -996
rect 394 -1004 395 -1002
rect 401 -998 402 -996
rect 401 -1004 402 -1002
rect 408 -998 409 -996
rect 408 -1004 409 -1002
rect 415 -998 416 -996
rect 415 -1004 416 -1002
rect 422 -998 423 -996
rect 422 -1004 423 -1002
rect 429 -998 430 -996
rect 429 -1004 430 -1002
rect 439 -998 440 -996
rect 436 -1004 437 -1002
rect 443 -998 444 -996
rect 443 -1004 444 -1002
rect 450 -998 451 -996
rect 450 -1004 451 -1002
rect 457 -998 458 -996
rect 457 -1004 458 -1002
rect 464 -1004 465 -1002
rect 471 -998 472 -996
rect 471 -1004 472 -1002
rect 478 -998 479 -996
rect 478 -1004 479 -1002
rect 485 -998 486 -996
rect 485 -1004 486 -1002
rect 492 -998 493 -996
rect 492 -1004 493 -1002
rect 499 -998 500 -996
rect 502 -998 503 -996
rect 499 -1004 500 -1002
rect 502 -1004 503 -1002
rect 506 -1004 507 -1002
rect 509 -1004 510 -1002
rect 513 -998 514 -996
rect 513 -1004 514 -1002
rect 520 -998 521 -996
rect 520 -1004 521 -1002
rect 527 -998 528 -996
rect 527 -1004 528 -1002
rect 534 -998 535 -996
rect 534 -1004 535 -1002
rect 544 -998 545 -996
rect 541 -1004 542 -1002
rect 544 -1004 545 -1002
rect 548 -998 549 -996
rect 548 -1004 549 -1002
rect 555 -998 556 -996
rect 555 -1004 556 -1002
rect 562 -998 563 -996
rect 562 -1004 563 -1002
rect 569 -998 570 -996
rect 569 -1004 570 -1002
rect 576 -998 577 -996
rect 576 -1004 577 -1002
rect 583 -998 584 -996
rect 583 -1004 584 -1002
rect 590 -998 591 -996
rect 590 -1004 591 -1002
rect 597 -998 598 -996
rect 597 -1004 598 -1002
rect 604 -998 605 -996
rect 607 -998 608 -996
rect 607 -1004 608 -1002
rect 611 -998 612 -996
rect 611 -1004 612 -1002
rect 618 -998 619 -996
rect 618 -1004 619 -1002
rect 628 -998 629 -996
rect 632 -998 633 -996
rect 632 -1004 633 -1002
rect 639 -1004 640 -1002
rect 642 -1004 643 -1002
rect 649 -1004 650 -1002
rect 653 -998 654 -996
rect 653 -1004 654 -1002
rect 660 -998 661 -996
rect 660 -1004 661 -1002
rect 667 -998 668 -996
rect 667 -1004 668 -1002
rect 674 -998 675 -996
rect 674 -1004 675 -1002
rect 681 -998 682 -996
rect 681 -1004 682 -1002
rect 684 -1004 685 -1002
rect 688 -998 689 -996
rect 688 -1004 689 -1002
rect 695 -998 696 -996
rect 698 -1004 699 -1002
rect 702 -998 703 -996
rect 702 -1004 703 -1002
rect 709 -998 710 -996
rect 712 -998 713 -996
rect 709 -1004 710 -1002
rect 716 -998 717 -996
rect 716 -1004 717 -1002
rect 723 -998 724 -996
rect 723 -1004 724 -1002
rect 730 -998 731 -996
rect 733 -998 734 -996
rect 730 -1004 731 -1002
rect 737 -998 738 -996
rect 737 -1004 738 -1002
rect 744 -998 745 -996
rect 744 -1004 745 -1002
rect 751 -998 752 -996
rect 751 -1004 752 -1002
rect 758 -998 759 -996
rect 758 -1004 759 -1002
rect 765 -998 766 -996
rect 765 -1004 766 -1002
rect 772 -998 773 -996
rect 772 -1004 773 -1002
rect 779 -998 780 -996
rect 779 -1004 780 -1002
rect 786 -998 787 -996
rect 786 -1004 787 -1002
rect 793 -998 794 -996
rect 793 -1004 794 -1002
rect 800 -998 801 -996
rect 800 -1004 801 -1002
rect 807 -998 808 -996
rect 807 -1004 808 -1002
rect 814 -998 815 -996
rect 814 -1004 815 -1002
rect 821 -998 822 -996
rect 821 -1004 822 -1002
rect 828 -998 829 -996
rect 828 -1004 829 -1002
rect 835 -998 836 -996
rect 835 -1004 836 -1002
rect 842 -998 843 -996
rect 842 -1004 843 -1002
rect 849 -998 850 -996
rect 849 -1004 850 -1002
rect 859 -998 860 -996
rect 856 -1004 857 -1002
rect 859 -1004 860 -1002
rect 863 -998 864 -996
rect 863 -1004 864 -1002
rect 870 -998 871 -996
rect 870 -1004 871 -1002
rect 877 -998 878 -996
rect 877 -1004 878 -1002
rect 884 -998 885 -996
rect 884 -1004 885 -1002
rect 891 -998 892 -996
rect 891 -1004 892 -1002
rect 898 -998 899 -996
rect 898 -1004 899 -1002
rect 905 -998 906 -996
rect 905 -1004 906 -1002
rect 912 -998 913 -996
rect 912 -1004 913 -1002
rect 919 -998 920 -996
rect 919 -1004 920 -1002
rect 926 -998 927 -996
rect 926 -1004 927 -1002
rect 933 -998 934 -996
rect 933 -1004 934 -1002
rect 940 -998 941 -996
rect 940 -1004 941 -1002
rect 947 -998 948 -996
rect 947 -1004 948 -1002
rect 954 -998 955 -996
rect 954 -1004 955 -1002
rect 961 -998 962 -996
rect 961 -1004 962 -1002
rect 968 -998 969 -996
rect 968 -1004 969 -1002
rect 975 -998 976 -996
rect 975 -1004 976 -1002
rect 982 -998 983 -996
rect 982 -1004 983 -1002
rect 989 -998 990 -996
rect 989 -1004 990 -1002
rect 996 -998 997 -996
rect 996 -1004 997 -1002
rect 1003 -998 1004 -996
rect 1003 -1004 1004 -1002
rect 1010 -998 1011 -996
rect 1010 -1004 1011 -1002
rect 1017 -998 1018 -996
rect 1017 -1004 1018 -1002
rect 1024 -998 1025 -996
rect 1024 -1004 1025 -1002
rect 1031 -998 1032 -996
rect 1031 -1004 1032 -1002
rect 1038 -998 1039 -996
rect 1038 -1004 1039 -1002
rect 1045 -998 1046 -996
rect 1045 -1004 1046 -1002
rect 1052 -998 1053 -996
rect 1052 -1004 1053 -1002
rect 1059 -998 1060 -996
rect 1059 -1004 1060 -1002
rect 1066 -998 1067 -996
rect 1066 -1004 1067 -1002
rect 1073 -998 1074 -996
rect 1073 -1004 1074 -1002
rect 1080 -998 1081 -996
rect 1080 -1004 1081 -1002
rect 1087 -998 1088 -996
rect 1087 -1004 1088 -1002
rect 1094 -998 1095 -996
rect 1094 -1004 1095 -1002
rect 1101 -998 1102 -996
rect 1101 -1004 1102 -1002
rect 1108 -998 1109 -996
rect 1108 -1004 1109 -1002
rect 1115 -998 1116 -996
rect 1115 -1004 1116 -1002
rect 1122 -998 1123 -996
rect 1122 -1004 1123 -1002
rect 1129 -998 1130 -996
rect 1129 -1004 1130 -1002
rect 1132 -1004 1133 -1002
rect 1136 -998 1137 -996
rect 1136 -1004 1137 -1002
rect 1143 -998 1144 -996
rect 1143 -1004 1144 -1002
rect 1150 -998 1151 -996
rect 1150 -1004 1151 -1002
rect 1157 -998 1158 -996
rect 1157 -1004 1158 -1002
rect 1164 -998 1165 -996
rect 1167 -1004 1168 -1002
rect 1171 -998 1172 -996
rect 1171 -1004 1172 -1002
rect 1185 -998 1186 -996
rect 1185 -1004 1186 -1002
rect 1192 -998 1193 -996
rect 16 -1073 17 -1071
rect 16 -1079 17 -1077
rect 23 -1073 24 -1071
rect 23 -1079 24 -1077
rect 30 -1073 31 -1071
rect 30 -1079 31 -1077
rect 37 -1073 38 -1071
rect 37 -1079 38 -1077
rect 44 -1073 45 -1071
rect 44 -1079 45 -1077
rect 51 -1073 52 -1071
rect 51 -1079 52 -1077
rect 58 -1073 59 -1071
rect 61 -1073 62 -1071
rect 65 -1073 66 -1071
rect 68 -1079 69 -1077
rect 72 -1073 73 -1071
rect 72 -1079 73 -1077
rect 79 -1073 80 -1071
rect 79 -1079 80 -1077
rect 86 -1073 87 -1071
rect 89 -1073 90 -1071
rect 93 -1073 94 -1071
rect 96 -1073 97 -1071
rect 100 -1073 101 -1071
rect 100 -1079 101 -1077
rect 107 -1073 108 -1071
rect 107 -1079 108 -1077
rect 117 -1073 118 -1071
rect 121 -1073 122 -1071
rect 121 -1079 122 -1077
rect 128 -1073 129 -1071
rect 128 -1079 129 -1077
rect 135 -1073 136 -1071
rect 135 -1079 136 -1077
rect 142 -1073 143 -1071
rect 142 -1079 143 -1077
rect 152 -1073 153 -1071
rect 149 -1079 150 -1077
rect 156 -1073 157 -1071
rect 156 -1079 157 -1077
rect 163 -1073 164 -1071
rect 163 -1079 164 -1077
rect 173 -1073 174 -1071
rect 170 -1079 171 -1077
rect 177 -1073 178 -1071
rect 177 -1079 178 -1077
rect 184 -1073 185 -1071
rect 184 -1079 185 -1077
rect 191 -1073 192 -1071
rect 191 -1079 192 -1077
rect 198 -1073 199 -1071
rect 198 -1079 199 -1077
rect 205 -1073 206 -1071
rect 208 -1073 209 -1071
rect 205 -1079 206 -1077
rect 212 -1073 213 -1071
rect 212 -1079 213 -1077
rect 219 -1073 220 -1071
rect 219 -1079 220 -1077
rect 226 -1073 227 -1071
rect 226 -1079 227 -1077
rect 233 -1073 234 -1071
rect 233 -1079 234 -1077
rect 240 -1073 241 -1071
rect 240 -1079 241 -1077
rect 247 -1073 248 -1071
rect 247 -1079 248 -1077
rect 254 -1073 255 -1071
rect 254 -1079 255 -1077
rect 264 -1073 265 -1071
rect 261 -1079 262 -1077
rect 264 -1079 265 -1077
rect 268 -1073 269 -1071
rect 268 -1079 269 -1077
rect 275 -1073 276 -1071
rect 275 -1079 276 -1077
rect 282 -1073 283 -1071
rect 282 -1079 283 -1077
rect 289 -1073 290 -1071
rect 289 -1079 290 -1077
rect 296 -1079 297 -1077
rect 299 -1079 300 -1077
rect 303 -1073 304 -1071
rect 303 -1079 304 -1077
rect 310 -1073 311 -1071
rect 310 -1079 311 -1077
rect 317 -1073 318 -1071
rect 320 -1073 321 -1071
rect 317 -1079 318 -1077
rect 324 -1073 325 -1071
rect 324 -1079 325 -1077
rect 331 -1073 332 -1071
rect 331 -1079 332 -1077
rect 338 -1073 339 -1071
rect 338 -1079 339 -1077
rect 345 -1073 346 -1071
rect 345 -1079 346 -1077
rect 352 -1073 353 -1071
rect 355 -1073 356 -1071
rect 355 -1079 356 -1077
rect 359 -1073 360 -1071
rect 359 -1079 360 -1077
rect 366 -1073 367 -1071
rect 366 -1079 367 -1077
rect 373 -1073 374 -1071
rect 373 -1079 374 -1077
rect 380 -1073 381 -1071
rect 380 -1079 381 -1077
rect 387 -1073 388 -1071
rect 387 -1079 388 -1077
rect 394 -1073 395 -1071
rect 394 -1079 395 -1077
rect 401 -1073 402 -1071
rect 401 -1079 402 -1077
rect 408 -1073 409 -1071
rect 408 -1079 409 -1077
rect 415 -1073 416 -1071
rect 415 -1079 416 -1077
rect 422 -1073 423 -1071
rect 422 -1079 423 -1077
rect 429 -1073 430 -1071
rect 429 -1079 430 -1077
rect 436 -1073 437 -1071
rect 436 -1079 437 -1077
rect 443 -1073 444 -1071
rect 443 -1079 444 -1077
rect 450 -1073 451 -1071
rect 450 -1079 451 -1077
rect 457 -1073 458 -1071
rect 457 -1079 458 -1077
rect 464 -1079 465 -1077
rect 467 -1079 468 -1077
rect 471 -1073 472 -1071
rect 471 -1079 472 -1077
rect 478 -1073 479 -1071
rect 478 -1079 479 -1077
rect 485 -1073 486 -1071
rect 485 -1079 486 -1077
rect 492 -1073 493 -1071
rect 492 -1079 493 -1077
rect 499 -1073 500 -1071
rect 499 -1079 500 -1077
rect 506 -1079 507 -1077
rect 509 -1079 510 -1077
rect 513 -1073 514 -1071
rect 513 -1079 514 -1077
rect 520 -1073 521 -1071
rect 520 -1079 521 -1077
rect 527 -1073 528 -1071
rect 527 -1079 528 -1077
rect 534 -1073 535 -1071
rect 534 -1079 535 -1077
rect 537 -1079 538 -1077
rect 541 -1073 542 -1071
rect 541 -1079 542 -1077
rect 548 -1073 549 -1071
rect 548 -1079 549 -1077
rect 555 -1073 556 -1071
rect 555 -1079 556 -1077
rect 562 -1073 563 -1071
rect 562 -1079 563 -1077
rect 572 -1073 573 -1071
rect 569 -1079 570 -1077
rect 572 -1079 573 -1077
rect 576 -1073 577 -1071
rect 576 -1079 577 -1077
rect 583 -1073 584 -1071
rect 583 -1079 584 -1077
rect 590 -1073 591 -1071
rect 590 -1079 591 -1077
rect 597 -1073 598 -1071
rect 600 -1073 601 -1071
rect 600 -1079 601 -1077
rect 604 -1073 605 -1071
rect 604 -1079 605 -1077
rect 611 -1073 612 -1071
rect 611 -1079 612 -1077
rect 618 -1073 619 -1071
rect 621 -1073 622 -1071
rect 621 -1079 622 -1077
rect 625 -1073 626 -1071
rect 625 -1079 626 -1077
rect 632 -1079 633 -1077
rect 639 -1073 640 -1071
rect 639 -1079 640 -1077
rect 646 -1073 647 -1071
rect 646 -1079 647 -1077
rect 653 -1073 654 -1071
rect 653 -1079 654 -1077
rect 660 -1073 661 -1071
rect 660 -1079 661 -1077
rect 667 -1073 668 -1071
rect 667 -1079 668 -1077
rect 674 -1073 675 -1071
rect 674 -1079 675 -1077
rect 681 -1073 682 -1071
rect 681 -1079 682 -1077
rect 688 -1073 689 -1071
rect 691 -1073 692 -1071
rect 688 -1079 689 -1077
rect 695 -1073 696 -1071
rect 695 -1079 696 -1077
rect 702 -1073 703 -1071
rect 702 -1079 703 -1077
rect 709 -1073 710 -1071
rect 709 -1079 710 -1077
rect 716 -1073 717 -1071
rect 716 -1079 717 -1077
rect 723 -1073 724 -1071
rect 723 -1079 724 -1077
rect 733 -1073 734 -1071
rect 733 -1079 734 -1077
rect 737 -1073 738 -1071
rect 737 -1079 738 -1077
rect 744 -1073 745 -1071
rect 744 -1079 745 -1077
rect 751 -1073 752 -1071
rect 751 -1079 752 -1077
rect 758 -1079 759 -1077
rect 765 -1073 766 -1071
rect 765 -1079 766 -1077
rect 772 -1073 773 -1071
rect 772 -1079 773 -1077
rect 779 -1073 780 -1071
rect 779 -1079 780 -1077
rect 786 -1073 787 -1071
rect 786 -1079 787 -1077
rect 793 -1073 794 -1071
rect 793 -1079 794 -1077
rect 800 -1073 801 -1071
rect 800 -1079 801 -1077
rect 810 -1073 811 -1071
rect 810 -1079 811 -1077
rect 814 -1073 815 -1071
rect 814 -1079 815 -1077
rect 821 -1073 822 -1071
rect 821 -1079 822 -1077
rect 828 -1073 829 -1071
rect 828 -1079 829 -1077
rect 835 -1073 836 -1071
rect 835 -1079 836 -1077
rect 842 -1073 843 -1071
rect 842 -1079 843 -1077
rect 849 -1073 850 -1071
rect 849 -1079 850 -1077
rect 856 -1073 857 -1071
rect 856 -1079 857 -1077
rect 863 -1073 864 -1071
rect 863 -1079 864 -1077
rect 870 -1073 871 -1071
rect 870 -1079 871 -1077
rect 877 -1073 878 -1071
rect 877 -1079 878 -1077
rect 884 -1073 885 -1071
rect 884 -1079 885 -1077
rect 891 -1073 892 -1071
rect 891 -1079 892 -1077
rect 898 -1073 899 -1071
rect 898 -1079 899 -1077
rect 905 -1073 906 -1071
rect 905 -1079 906 -1077
rect 912 -1073 913 -1071
rect 912 -1079 913 -1077
rect 919 -1073 920 -1071
rect 919 -1079 920 -1077
rect 926 -1073 927 -1071
rect 926 -1079 927 -1077
rect 933 -1073 934 -1071
rect 933 -1079 934 -1077
rect 940 -1073 941 -1071
rect 940 -1079 941 -1077
rect 947 -1073 948 -1071
rect 947 -1079 948 -1077
rect 954 -1073 955 -1071
rect 957 -1079 958 -1077
rect 961 -1073 962 -1071
rect 961 -1079 962 -1077
rect 968 -1073 969 -1071
rect 968 -1079 969 -1077
rect 975 -1073 976 -1071
rect 975 -1079 976 -1077
rect 982 -1073 983 -1071
rect 982 -1079 983 -1077
rect 989 -1073 990 -1071
rect 989 -1079 990 -1077
rect 996 -1073 997 -1071
rect 996 -1079 997 -1077
rect 1003 -1073 1004 -1071
rect 1003 -1079 1004 -1077
rect 1010 -1073 1011 -1071
rect 1010 -1079 1011 -1077
rect 1017 -1073 1018 -1071
rect 1017 -1079 1018 -1077
rect 1024 -1073 1025 -1071
rect 1024 -1079 1025 -1077
rect 1031 -1073 1032 -1071
rect 1031 -1079 1032 -1077
rect 1038 -1073 1039 -1071
rect 1041 -1079 1042 -1077
rect 1045 -1073 1046 -1071
rect 1045 -1079 1046 -1077
rect 1052 -1073 1053 -1071
rect 1052 -1079 1053 -1077
rect 1059 -1073 1060 -1071
rect 1066 -1073 1067 -1071
rect 1069 -1073 1070 -1071
rect 1066 -1079 1067 -1077
rect 1073 -1073 1074 -1071
rect 1073 -1079 1074 -1077
rect 1080 -1073 1081 -1071
rect 1080 -1079 1081 -1077
rect 1087 -1073 1088 -1071
rect 1087 -1079 1088 -1077
rect 1094 -1073 1095 -1071
rect 1094 -1079 1095 -1077
rect 1122 -1073 1123 -1071
rect 1122 -1079 1123 -1077
rect 1185 -1073 1186 -1071
rect 1185 -1079 1186 -1077
rect 23 -1162 24 -1160
rect 30 -1156 31 -1154
rect 30 -1162 31 -1160
rect 37 -1156 38 -1154
rect 37 -1162 38 -1160
rect 44 -1156 45 -1154
rect 44 -1162 45 -1160
rect 51 -1156 52 -1154
rect 51 -1162 52 -1160
rect 58 -1156 59 -1154
rect 58 -1162 59 -1160
rect 65 -1156 66 -1154
rect 65 -1162 66 -1160
rect 72 -1156 73 -1154
rect 72 -1162 73 -1160
rect 82 -1156 83 -1154
rect 82 -1162 83 -1160
rect 89 -1162 90 -1160
rect 93 -1156 94 -1154
rect 93 -1162 94 -1160
rect 100 -1156 101 -1154
rect 100 -1162 101 -1160
rect 107 -1156 108 -1154
rect 107 -1162 108 -1160
rect 117 -1156 118 -1154
rect 114 -1162 115 -1160
rect 117 -1162 118 -1160
rect 121 -1156 122 -1154
rect 121 -1162 122 -1160
rect 128 -1156 129 -1154
rect 131 -1162 132 -1160
rect 135 -1156 136 -1154
rect 138 -1162 139 -1160
rect 142 -1156 143 -1154
rect 142 -1162 143 -1160
rect 149 -1156 150 -1154
rect 149 -1162 150 -1160
rect 156 -1156 157 -1154
rect 156 -1162 157 -1160
rect 166 -1156 167 -1154
rect 163 -1162 164 -1160
rect 166 -1162 167 -1160
rect 170 -1156 171 -1154
rect 170 -1162 171 -1160
rect 177 -1156 178 -1154
rect 177 -1162 178 -1160
rect 184 -1156 185 -1154
rect 187 -1156 188 -1154
rect 187 -1162 188 -1160
rect 191 -1156 192 -1154
rect 191 -1162 192 -1160
rect 198 -1162 199 -1160
rect 205 -1156 206 -1154
rect 205 -1162 206 -1160
rect 212 -1156 213 -1154
rect 212 -1162 213 -1160
rect 219 -1156 220 -1154
rect 219 -1162 220 -1160
rect 226 -1156 227 -1154
rect 229 -1162 230 -1160
rect 233 -1156 234 -1154
rect 233 -1162 234 -1160
rect 240 -1156 241 -1154
rect 240 -1162 241 -1160
rect 247 -1156 248 -1154
rect 247 -1162 248 -1160
rect 254 -1156 255 -1154
rect 254 -1162 255 -1160
rect 261 -1156 262 -1154
rect 261 -1162 262 -1160
rect 268 -1156 269 -1154
rect 268 -1162 269 -1160
rect 275 -1156 276 -1154
rect 275 -1162 276 -1160
rect 282 -1156 283 -1154
rect 285 -1162 286 -1160
rect 289 -1156 290 -1154
rect 289 -1162 290 -1160
rect 296 -1156 297 -1154
rect 296 -1162 297 -1160
rect 306 -1156 307 -1154
rect 306 -1162 307 -1160
rect 310 -1156 311 -1154
rect 310 -1162 311 -1160
rect 317 -1156 318 -1154
rect 317 -1162 318 -1160
rect 324 -1156 325 -1154
rect 324 -1162 325 -1160
rect 331 -1156 332 -1154
rect 338 -1156 339 -1154
rect 338 -1162 339 -1160
rect 345 -1156 346 -1154
rect 345 -1162 346 -1160
rect 352 -1156 353 -1154
rect 352 -1162 353 -1160
rect 359 -1156 360 -1154
rect 359 -1162 360 -1160
rect 366 -1156 367 -1154
rect 366 -1162 367 -1160
rect 373 -1156 374 -1154
rect 373 -1162 374 -1160
rect 380 -1156 381 -1154
rect 380 -1162 381 -1160
rect 387 -1156 388 -1154
rect 387 -1162 388 -1160
rect 394 -1156 395 -1154
rect 394 -1162 395 -1160
rect 401 -1156 402 -1154
rect 401 -1162 402 -1160
rect 408 -1156 409 -1154
rect 408 -1162 409 -1160
rect 415 -1156 416 -1154
rect 418 -1156 419 -1154
rect 415 -1162 416 -1160
rect 422 -1156 423 -1154
rect 422 -1162 423 -1160
rect 429 -1156 430 -1154
rect 429 -1162 430 -1160
rect 436 -1156 437 -1154
rect 436 -1162 437 -1160
rect 446 -1156 447 -1154
rect 446 -1162 447 -1160
rect 450 -1156 451 -1154
rect 450 -1162 451 -1160
rect 457 -1156 458 -1154
rect 457 -1162 458 -1160
rect 464 -1156 465 -1154
rect 464 -1162 465 -1160
rect 471 -1156 472 -1154
rect 471 -1162 472 -1160
rect 478 -1156 479 -1154
rect 478 -1162 479 -1160
rect 485 -1156 486 -1154
rect 485 -1162 486 -1160
rect 492 -1156 493 -1154
rect 492 -1162 493 -1160
rect 499 -1156 500 -1154
rect 499 -1162 500 -1160
rect 506 -1162 507 -1160
rect 509 -1162 510 -1160
rect 513 -1156 514 -1154
rect 513 -1162 514 -1160
rect 520 -1156 521 -1154
rect 520 -1162 521 -1160
rect 527 -1156 528 -1154
rect 527 -1162 528 -1160
rect 534 -1156 535 -1154
rect 534 -1162 535 -1160
rect 541 -1156 542 -1154
rect 541 -1162 542 -1160
rect 548 -1156 549 -1154
rect 551 -1156 552 -1154
rect 551 -1162 552 -1160
rect 555 -1156 556 -1154
rect 555 -1162 556 -1160
rect 562 -1156 563 -1154
rect 562 -1162 563 -1160
rect 569 -1156 570 -1154
rect 569 -1162 570 -1160
rect 576 -1156 577 -1154
rect 576 -1162 577 -1160
rect 583 -1156 584 -1154
rect 586 -1156 587 -1154
rect 583 -1162 584 -1160
rect 586 -1162 587 -1160
rect 590 -1156 591 -1154
rect 590 -1162 591 -1160
rect 597 -1156 598 -1154
rect 597 -1162 598 -1160
rect 607 -1156 608 -1154
rect 604 -1162 605 -1160
rect 607 -1162 608 -1160
rect 611 -1156 612 -1154
rect 611 -1162 612 -1160
rect 618 -1156 619 -1154
rect 618 -1162 619 -1160
rect 628 -1156 629 -1154
rect 625 -1162 626 -1160
rect 632 -1156 633 -1154
rect 632 -1162 633 -1160
rect 639 -1156 640 -1154
rect 639 -1162 640 -1160
rect 646 -1156 647 -1154
rect 646 -1162 647 -1160
rect 653 -1156 654 -1154
rect 656 -1162 657 -1160
rect 660 -1156 661 -1154
rect 660 -1162 661 -1160
rect 667 -1156 668 -1154
rect 670 -1156 671 -1154
rect 667 -1162 668 -1160
rect 674 -1156 675 -1154
rect 674 -1162 675 -1160
rect 681 -1156 682 -1154
rect 681 -1162 682 -1160
rect 688 -1156 689 -1154
rect 688 -1162 689 -1160
rect 695 -1156 696 -1154
rect 695 -1162 696 -1160
rect 702 -1156 703 -1154
rect 702 -1162 703 -1160
rect 709 -1156 710 -1154
rect 709 -1162 710 -1160
rect 716 -1156 717 -1154
rect 716 -1162 717 -1160
rect 723 -1156 724 -1154
rect 723 -1162 724 -1160
rect 730 -1156 731 -1154
rect 730 -1162 731 -1160
rect 737 -1156 738 -1154
rect 737 -1162 738 -1160
rect 744 -1156 745 -1154
rect 744 -1162 745 -1160
rect 751 -1156 752 -1154
rect 751 -1162 752 -1160
rect 758 -1156 759 -1154
rect 758 -1162 759 -1160
rect 765 -1156 766 -1154
rect 765 -1162 766 -1160
rect 772 -1156 773 -1154
rect 772 -1162 773 -1160
rect 779 -1156 780 -1154
rect 779 -1162 780 -1160
rect 786 -1156 787 -1154
rect 786 -1162 787 -1160
rect 793 -1156 794 -1154
rect 793 -1162 794 -1160
rect 800 -1156 801 -1154
rect 800 -1162 801 -1160
rect 807 -1156 808 -1154
rect 810 -1156 811 -1154
rect 810 -1162 811 -1160
rect 814 -1156 815 -1154
rect 814 -1162 815 -1160
rect 821 -1156 822 -1154
rect 821 -1162 822 -1160
rect 828 -1156 829 -1154
rect 828 -1162 829 -1160
rect 835 -1156 836 -1154
rect 835 -1162 836 -1160
rect 842 -1156 843 -1154
rect 842 -1162 843 -1160
rect 852 -1156 853 -1154
rect 856 -1156 857 -1154
rect 856 -1162 857 -1160
rect 863 -1156 864 -1154
rect 863 -1162 864 -1160
rect 870 -1156 871 -1154
rect 870 -1162 871 -1160
rect 877 -1156 878 -1154
rect 877 -1162 878 -1160
rect 884 -1156 885 -1154
rect 884 -1162 885 -1160
rect 891 -1156 892 -1154
rect 891 -1162 892 -1160
rect 898 -1156 899 -1154
rect 898 -1162 899 -1160
rect 905 -1156 906 -1154
rect 905 -1162 906 -1160
rect 912 -1156 913 -1154
rect 912 -1162 913 -1160
rect 919 -1156 920 -1154
rect 919 -1162 920 -1160
rect 926 -1156 927 -1154
rect 926 -1162 927 -1160
rect 933 -1156 934 -1154
rect 936 -1162 937 -1160
rect 940 -1156 941 -1154
rect 940 -1162 941 -1160
rect 947 -1156 948 -1154
rect 947 -1162 948 -1160
rect 954 -1156 955 -1154
rect 954 -1162 955 -1160
rect 961 -1156 962 -1154
rect 961 -1162 962 -1160
rect 968 -1156 969 -1154
rect 968 -1162 969 -1160
rect 978 -1156 979 -1154
rect 975 -1162 976 -1160
rect 978 -1162 979 -1160
rect 982 -1156 983 -1154
rect 982 -1162 983 -1160
rect 989 -1156 990 -1154
rect 989 -1162 990 -1160
rect 996 -1156 997 -1154
rect 996 -1162 997 -1160
rect 1003 -1156 1004 -1154
rect 1006 -1156 1007 -1154
rect 1010 -1156 1011 -1154
rect 1010 -1162 1011 -1160
rect 1017 -1156 1018 -1154
rect 1017 -1162 1018 -1160
rect 1024 -1156 1025 -1154
rect 1024 -1162 1025 -1160
rect 1031 -1156 1032 -1154
rect 1031 -1162 1032 -1160
rect 1038 -1156 1039 -1154
rect 1038 -1162 1039 -1160
rect 1048 -1156 1049 -1154
rect 1059 -1156 1060 -1154
rect 1059 -1162 1060 -1160
rect 1066 -1156 1067 -1154
rect 1066 -1162 1067 -1160
rect 1080 -1156 1081 -1154
rect 1080 -1162 1081 -1160
rect 1087 -1156 1088 -1154
rect 1087 -1162 1088 -1160
rect 1108 -1156 1109 -1154
rect 1108 -1162 1109 -1160
rect 1188 -1156 1189 -1154
rect 16 -1231 17 -1229
rect 16 -1237 17 -1235
rect 23 -1231 24 -1229
rect 26 -1231 27 -1229
rect 30 -1231 31 -1229
rect 30 -1237 31 -1235
rect 37 -1231 38 -1229
rect 37 -1237 38 -1235
rect 44 -1237 45 -1235
rect 47 -1237 48 -1235
rect 51 -1231 52 -1229
rect 51 -1237 52 -1235
rect 58 -1231 59 -1229
rect 61 -1231 62 -1229
rect 65 -1231 66 -1229
rect 68 -1237 69 -1235
rect 72 -1231 73 -1229
rect 72 -1237 73 -1235
rect 79 -1231 80 -1229
rect 79 -1237 80 -1235
rect 93 -1231 94 -1229
rect 93 -1237 94 -1235
rect 100 -1231 101 -1229
rect 100 -1237 101 -1235
rect 107 -1231 108 -1229
rect 107 -1237 108 -1235
rect 117 -1237 118 -1235
rect 121 -1231 122 -1229
rect 121 -1237 122 -1235
rect 128 -1231 129 -1229
rect 128 -1237 129 -1235
rect 135 -1231 136 -1229
rect 135 -1237 136 -1235
rect 142 -1231 143 -1229
rect 142 -1237 143 -1235
rect 152 -1231 153 -1229
rect 149 -1237 150 -1235
rect 152 -1237 153 -1235
rect 156 -1231 157 -1229
rect 156 -1237 157 -1235
rect 163 -1231 164 -1229
rect 163 -1237 164 -1235
rect 170 -1231 171 -1229
rect 170 -1237 171 -1235
rect 177 -1237 178 -1235
rect 180 -1237 181 -1235
rect 184 -1231 185 -1229
rect 184 -1237 185 -1235
rect 191 -1231 192 -1229
rect 191 -1237 192 -1235
rect 198 -1231 199 -1229
rect 198 -1237 199 -1235
rect 205 -1231 206 -1229
rect 205 -1237 206 -1235
rect 212 -1231 213 -1229
rect 212 -1237 213 -1235
rect 219 -1231 220 -1229
rect 219 -1237 220 -1235
rect 226 -1231 227 -1229
rect 226 -1237 227 -1235
rect 233 -1231 234 -1229
rect 233 -1237 234 -1235
rect 240 -1231 241 -1229
rect 240 -1237 241 -1235
rect 247 -1231 248 -1229
rect 247 -1237 248 -1235
rect 254 -1231 255 -1229
rect 254 -1237 255 -1235
rect 264 -1237 265 -1235
rect 268 -1231 269 -1229
rect 268 -1237 269 -1235
rect 275 -1231 276 -1229
rect 275 -1237 276 -1235
rect 282 -1231 283 -1229
rect 282 -1237 283 -1235
rect 289 -1231 290 -1229
rect 289 -1237 290 -1235
rect 296 -1231 297 -1229
rect 296 -1237 297 -1235
rect 303 -1231 304 -1229
rect 303 -1237 304 -1235
rect 310 -1231 311 -1229
rect 310 -1237 311 -1235
rect 317 -1231 318 -1229
rect 317 -1237 318 -1235
rect 320 -1237 321 -1235
rect 324 -1231 325 -1229
rect 324 -1237 325 -1235
rect 331 -1231 332 -1229
rect 331 -1237 332 -1235
rect 338 -1231 339 -1229
rect 338 -1237 339 -1235
rect 345 -1231 346 -1229
rect 345 -1237 346 -1235
rect 352 -1231 353 -1229
rect 352 -1237 353 -1235
rect 359 -1231 360 -1229
rect 359 -1237 360 -1235
rect 366 -1231 367 -1229
rect 366 -1237 367 -1235
rect 373 -1231 374 -1229
rect 376 -1237 377 -1235
rect 383 -1231 384 -1229
rect 380 -1237 381 -1235
rect 387 -1237 388 -1235
rect 390 -1237 391 -1235
rect 394 -1231 395 -1229
rect 394 -1237 395 -1235
rect 401 -1231 402 -1229
rect 401 -1237 402 -1235
rect 408 -1231 409 -1229
rect 408 -1237 409 -1235
rect 415 -1231 416 -1229
rect 415 -1237 416 -1235
rect 422 -1231 423 -1229
rect 422 -1237 423 -1235
rect 429 -1231 430 -1229
rect 429 -1237 430 -1235
rect 436 -1231 437 -1229
rect 436 -1237 437 -1235
rect 443 -1231 444 -1229
rect 446 -1237 447 -1235
rect 450 -1231 451 -1229
rect 450 -1237 451 -1235
rect 457 -1231 458 -1229
rect 457 -1237 458 -1235
rect 464 -1231 465 -1229
rect 464 -1237 465 -1235
rect 471 -1231 472 -1229
rect 471 -1237 472 -1235
rect 478 -1231 479 -1229
rect 478 -1237 479 -1235
rect 485 -1231 486 -1229
rect 485 -1237 486 -1235
rect 492 -1231 493 -1229
rect 492 -1237 493 -1235
rect 499 -1231 500 -1229
rect 499 -1237 500 -1235
rect 509 -1231 510 -1229
rect 506 -1237 507 -1235
rect 509 -1237 510 -1235
rect 513 -1231 514 -1229
rect 513 -1237 514 -1235
rect 520 -1231 521 -1229
rect 520 -1237 521 -1235
rect 527 -1231 528 -1229
rect 527 -1237 528 -1235
rect 534 -1231 535 -1229
rect 534 -1237 535 -1235
rect 544 -1231 545 -1229
rect 544 -1237 545 -1235
rect 548 -1231 549 -1229
rect 548 -1237 549 -1235
rect 555 -1231 556 -1229
rect 555 -1237 556 -1235
rect 562 -1231 563 -1229
rect 565 -1231 566 -1229
rect 562 -1237 563 -1235
rect 565 -1237 566 -1235
rect 569 -1231 570 -1229
rect 569 -1237 570 -1235
rect 572 -1237 573 -1235
rect 576 -1231 577 -1229
rect 576 -1237 577 -1235
rect 583 -1231 584 -1229
rect 583 -1237 584 -1235
rect 593 -1231 594 -1229
rect 590 -1237 591 -1235
rect 597 -1231 598 -1229
rect 597 -1237 598 -1235
rect 604 -1231 605 -1229
rect 604 -1237 605 -1235
rect 611 -1231 612 -1229
rect 611 -1237 612 -1235
rect 618 -1231 619 -1229
rect 618 -1237 619 -1235
rect 625 -1231 626 -1229
rect 625 -1237 626 -1235
rect 632 -1231 633 -1229
rect 632 -1237 633 -1235
rect 639 -1237 640 -1235
rect 642 -1237 643 -1235
rect 646 -1231 647 -1229
rect 646 -1237 647 -1235
rect 653 -1231 654 -1229
rect 656 -1231 657 -1229
rect 656 -1237 657 -1235
rect 660 -1237 661 -1235
rect 663 -1237 664 -1235
rect 667 -1231 668 -1229
rect 667 -1237 668 -1235
rect 674 -1231 675 -1229
rect 674 -1237 675 -1235
rect 681 -1231 682 -1229
rect 681 -1237 682 -1235
rect 688 -1231 689 -1229
rect 688 -1237 689 -1235
rect 695 -1231 696 -1229
rect 695 -1237 696 -1235
rect 702 -1231 703 -1229
rect 702 -1237 703 -1235
rect 709 -1231 710 -1229
rect 709 -1237 710 -1235
rect 716 -1231 717 -1229
rect 716 -1237 717 -1235
rect 723 -1231 724 -1229
rect 726 -1231 727 -1229
rect 723 -1237 724 -1235
rect 726 -1237 727 -1235
rect 730 -1231 731 -1229
rect 730 -1237 731 -1235
rect 737 -1231 738 -1229
rect 737 -1237 738 -1235
rect 744 -1231 745 -1229
rect 744 -1237 745 -1235
rect 751 -1231 752 -1229
rect 751 -1237 752 -1235
rect 758 -1231 759 -1229
rect 758 -1237 759 -1235
rect 765 -1231 766 -1229
rect 765 -1237 766 -1235
rect 772 -1231 773 -1229
rect 775 -1237 776 -1235
rect 779 -1231 780 -1229
rect 779 -1237 780 -1235
rect 786 -1231 787 -1229
rect 786 -1237 787 -1235
rect 793 -1231 794 -1229
rect 793 -1237 794 -1235
rect 800 -1231 801 -1229
rect 800 -1237 801 -1235
rect 807 -1231 808 -1229
rect 807 -1237 808 -1235
rect 814 -1231 815 -1229
rect 814 -1237 815 -1235
rect 821 -1231 822 -1229
rect 821 -1237 822 -1235
rect 828 -1231 829 -1229
rect 831 -1231 832 -1229
rect 828 -1237 829 -1235
rect 835 -1231 836 -1229
rect 835 -1237 836 -1235
rect 842 -1231 843 -1229
rect 842 -1237 843 -1235
rect 849 -1231 850 -1229
rect 849 -1237 850 -1235
rect 856 -1231 857 -1229
rect 856 -1237 857 -1235
rect 863 -1231 864 -1229
rect 863 -1237 864 -1235
rect 870 -1231 871 -1229
rect 870 -1237 871 -1235
rect 877 -1231 878 -1229
rect 877 -1237 878 -1235
rect 884 -1231 885 -1229
rect 884 -1237 885 -1235
rect 891 -1231 892 -1229
rect 891 -1237 892 -1235
rect 898 -1231 899 -1229
rect 898 -1237 899 -1235
rect 905 -1231 906 -1229
rect 905 -1237 906 -1235
rect 912 -1231 913 -1229
rect 912 -1237 913 -1235
rect 919 -1231 920 -1229
rect 919 -1237 920 -1235
rect 926 -1231 927 -1229
rect 926 -1237 927 -1235
rect 933 -1231 934 -1229
rect 933 -1237 934 -1235
rect 940 -1231 941 -1229
rect 940 -1237 941 -1235
rect 947 -1231 948 -1229
rect 947 -1237 948 -1235
rect 954 -1231 955 -1229
rect 954 -1237 955 -1235
rect 961 -1231 962 -1229
rect 961 -1237 962 -1235
rect 968 -1231 969 -1229
rect 968 -1237 969 -1235
rect 975 -1231 976 -1229
rect 975 -1237 976 -1235
rect 982 -1231 983 -1229
rect 982 -1237 983 -1235
rect 989 -1231 990 -1229
rect 989 -1237 990 -1235
rect 996 -1231 997 -1229
rect 996 -1237 997 -1235
rect 1003 -1231 1004 -1229
rect 1003 -1237 1004 -1235
rect 1010 -1231 1011 -1229
rect 1010 -1237 1011 -1235
rect 1017 -1231 1018 -1229
rect 1017 -1237 1018 -1235
rect 1024 -1231 1025 -1229
rect 1024 -1237 1025 -1235
rect 1031 -1231 1032 -1229
rect 1031 -1237 1032 -1235
rect 1038 -1231 1039 -1229
rect 1038 -1237 1039 -1235
rect 1045 -1231 1046 -1229
rect 1045 -1237 1046 -1235
rect 1052 -1231 1053 -1229
rect 1052 -1237 1053 -1235
rect 1059 -1231 1060 -1229
rect 1059 -1237 1060 -1235
rect 1066 -1231 1067 -1229
rect 1066 -1237 1067 -1235
rect 1073 -1231 1074 -1229
rect 1073 -1237 1074 -1235
rect 1080 -1231 1081 -1229
rect 1080 -1237 1081 -1235
rect 1087 -1231 1088 -1229
rect 1087 -1237 1088 -1235
rect 1094 -1231 1095 -1229
rect 1094 -1237 1095 -1235
rect 1101 -1231 1102 -1229
rect 1101 -1237 1102 -1235
rect 1108 -1231 1109 -1229
rect 1108 -1237 1109 -1235
rect 1115 -1231 1116 -1229
rect 1115 -1237 1116 -1235
rect 1122 -1231 1123 -1229
rect 1122 -1237 1123 -1235
rect 1129 -1231 1130 -1229
rect 1129 -1237 1130 -1235
rect 44 -1302 45 -1300
rect 44 -1308 45 -1306
rect 72 -1302 73 -1300
rect 72 -1308 73 -1306
rect 79 -1302 80 -1300
rect 79 -1308 80 -1306
rect 86 -1302 87 -1300
rect 86 -1308 87 -1306
rect 96 -1302 97 -1300
rect 93 -1308 94 -1306
rect 100 -1302 101 -1300
rect 100 -1308 101 -1306
rect 107 -1302 108 -1300
rect 107 -1308 108 -1306
rect 114 -1302 115 -1300
rect 114 -1308 115 -1306
rect 121 -1302 122 -1300
rect 121 -1308 122 -1306
rect 128 -1302 129 -1300
rect 128 -1308 129 -1306
rect 135 -1302 136 -1300
rect 135 -1308 136 -1306
rect 142 -1302 143 -1300
rect 142 -1308 143 -1306
rect 149 -1302 150 -1300
rect 149 -1308 150 -1306
rect 156 -1302 157 -1300
rect 156 -1308 157 -1306
rect 163 -1302 164 -1300
rect 163 -1308 164 -1306
rect 170 -1302 171 -1300
rect 170 -1308 171 -1306
rect 177 -1302 178 -1300
rect 177 -1308 178 -1306
rect 184 -1302 185 -1300
rect 184 -1308 185 -1306
rect 194 -1308 195 -1306
rect 198 -1302 199 -1300
rect 198 -1308 199 -1306
rect 205 -1302 206 -1300
rect 205 -1308 206 -1306
rect 212 -1302 213 -1300
rect 212 -1308 213 -1306
rect 219 -1302 220 -1300
rect 219 -1308 220 -1306
rect 226 -1302 227 -1300
rect 226 -1308 227 -1306
rect 233 -1302 234 -1300
rect 233 -1308 234 -1306
rect 240 -1302 241 -1300
rect 240 -1308 241 -1306
rect 247 -1302 248 -1300
rect 247 -1308 248 -1306
rect 254 -1302 255 -1300
rect 254 -1308 255 -1306
rect 261 -1302 262 -1300
rect 261 -1308 262 -1306
rect 268 -1302 269 -1300
rect 268 -1308 269 -1306
rect 275 -1302 276 -1300
rect 275 -1308 276 -1306
rect 282 -1302 283 -1300
rect 282 -1308 283 -1306
rect 289 -1302 290 -1300
rect 289 -1308 290 -1306
rect 296 -1302 297 -1300
rect 296 -1308 297 -1306
rect 303 -1302 304 -1300
rect 303 -1308 304 -1306
rect 306 -1308 307 -1306
rect 310 -1302 311 -1300
rect 310 -1308 311 -1306
rect 317 -1302 318 -1300
rect 317 -1308 318 -1306
rect 324 -1302 325 -1300
rect 324 -1308 325 -1306
rect 331 -1302 332 -1300
rect 331 -1308 332 -1306
rect 338 -1302 339 -1300
rect 341 -1302 342 -1300
rect 341 -1308 342 -1306
rect 345 -1302 346 -1300
rect 345 -1308 346 -1306
rect 352 -1302 353 -1300
rect 352 -1308 353 -1306
rect 359 -1302 360 -1300
rect 359 -1308 360 -1306
rect 366 -1302 367 -1300
rect 366 -1308 367 -1306
rect 373 -1302 374 -1300
rect 373 -1308 374 -1306
rect 380 -1302 381 -1300
rect 380 -1308 381 -1306
rect 387 -1302 388 -1300
rect 387 -1308 388 -1306
rect 394 -1302 395 -1300
rect 394 -1308 395 -1306
rect 401 -1302 402 -1300
rect 404 -1302 405 -1300
rect 404 -1308 405 -1306
rect 408 -1302 409 -1300
rect 408 -1308 409 -1306
rect 415 -1302 416 -1300
rect 415 -1308 416 -1306
rect 422 -1302 423 -1300
rect 422 -1308 423 -1306
rect 429 -1302 430 -1300
rect 429 -1308 430 -1306
rect 436 -1302 437 -1300
rect 436 -1308 437 -1306
rect 443 -1302 444 -1300
rect 443 -1308 444 -1306
rect 450 -1302 451 -1300
rect 450 -1308 451 -1306
rect 457 -1302 458 -1300
rect 457 -1308 458 -1306
rect 464 -1302 465 -1300
rect 467 -1302 468 -1300
rect 464 -1308 465 -1306
rect 467 -1308 468 -1306
rect 471 -1302 472 -1300
rect 471 -1308 472 -1306
rect 478 -1302 479 -1300
rect 481 -1302 482 -1300
rect 478 -1308 479 -1306
rect 481 -1308 482 -1306
rect 485 -1302 486 -1300
rect 485 -1308 486 -1306
rect 492 -1302 493 -1300
rect 492 -1308 493 -1306
rect 499 -1302 500 -1300
rect 502 -1302 503 -1300
rect 506 -1302 507 -1300
rect 506 -1308 507 -1306
rect 513 -1302 514 -1300
rect 513 -1308 514 -1306
rect 520 -1302 521 -1300
rect 520 -1308 521 -1306
rect 527 -1302 528 -1300
rect 527 -1308 528 -1306
rect 534 -1308 535 -1306
rect 537 -1308 538 -1306
rect 541 -1302 542 -1300
rect 541 -1308 542 -1306
rect 548 -1302 549 -1300
rect 548 -1308 549 -1306
rect 555 -1302 556 -1300
rect 555 -1308 556 -1306
rect 562 -1302 563 -1300
rect 562 -1308 563 -1306
rect 572 -1302 573 -1300
rect 569 -1308 570 -1306
rect 572 -1308 573 -1306
rect 579 -1302 580 -1300
rect 576 -1308 577 -1306
rect 583 -1302 584 -1300
rect 583 -1308 584 -1306
rect 590 -1302 591 -1300
rect 590 -1308 591 -1306
rect 597 -1308 598 -1306
rect 600 -1308 601 -1306
rect 604 -1302 605 -1300
rect 604 -1308 605 -1306
rect 611 -1302 612 -1300
rect 614 -1308 615 -1306
rect 618 -1302 619 -1300
rect 618 -1308 619 -1306
rect 625 -1302 626 -1300
rect 625 -1308 626 -1306
rect 635 -1308 636 -1306
rect 639 -1302 640 -1300
rect 639 -1308 640 -1306
rect 646 -1302 647 -1300
rect 646 -1308 647 -1306
rect 656 -1302 657 -1300
rect 660 -1302 661 -1300
rect 660 -1308 661 -1306
rect 667 -1302 668 -1300
rect 667 -1308 668 -1306
rect 674 -1302 675 -1300
rect 677 -1302 678 -1300
rect 674 -1308 675 -1306
rect 677 -1308 678 -1306
rect 681 -1302 682 -1300
rect 681 -1308 682 -1306
rect 688 -1302 689 -1300
rect 688 -1308 689 -1306
rect 695 -1302 696 -1300
rect 695 -1308 696 -1306
rect 702 -1302 703 -1300
rect 702 -1308 703 -1306
rect 709 -1302 710 -1300
rect 709 -1308 710 -1306
rect 716 -1302 717 -1300
rect 716 -1308 717 -1306
rect 723 -1302 724 -1300
rect 723 -1308 724 -1306
rect 730 -1302 731 -1300
rect 730 -1308 731 -1306
rect 737 -1302 738 -1300
rect 737 -1308 738 -1306
rect 744 -1302 745 -1300
rect 744 -1308 745 -1306
rect 751 -1302 752 -1300
rect 751 -1308 752 -1306
rect 758 -1302 759 -1300
rect 758 -1308 759 -1306
rect 765 -1302 766 -1300
rect 765 -1308 766 -1306
rect 772 -1302 773 -1300
rect 772 -1308 773 -1306
rect 779 -1302 780 -1300
rect 779 -1308 780 -1306
rect 786 -1302 787 -1300
rect 786 -1308 787 -1306
rect 793 -1302 794 -1300
rect 796 -1302 797 -1300
rect 793 -1308 794 -1306
rect 796 -1308 797 -1306
rect 800 -1302 801 -1300
rect 800 -1308 801 -1306
rect 807 -1302 808 -1300
rect 807 -1308 808 -1306
rect 814 -1302 815 -1300
rect 814 -1308 815 -1306
rect 821 -1302 822 -1300
rect 821 -1308 822 -1306
rect 828 -1302 829 -1300
rect 828 -1308 829 -1306
rect 835 -1302 836 -1300
rect 835 -1308 836 -1306
rect 842 -1302 843 -1300
rect 842 -1308 843 -1306
rect 849 -1302 850 -1300
rect 849 -1308 850 -1306
rect 856 -1302 857 -1300
rect 856 -1308 857 -1306
rect 866 -1302 867 -1300
rect 863 -1308 864 -1306
rect 870 -1302 871 -1300
rect 870 -1308 871 -1306
rect 877 -1302 878 -1300
rect 877 -1308 878 -1306
rect 884 -1302 885 -1300
rect 884 -1308 885 -1306
rect 891 -1302 892 -1300
rect 891 -1308 892 -1306
rect 898 -1302 899 -1300
rect 898 -1308 899 -1306
rect 905 -1302 906 -1300
rect 905 -1308 906 -1306
rect 912 -1302 913 -1300
rect 912 -1308 913 -1306
rect 922 -1308 923 -1306
rect 926 -1302 927 -1300
rect 926 -1308 927 -1306
rect 933 -1302 934 -1300
rect 933 -1308 934 -1306
rect 940 -1302 941 -1300
rect 940 -1308 941 -1306
rect 947 -1302 948 -1300
rect 947 -1308 948 -1306
rect 954 -1302 955 -1300
rect 954 -1308 955 -1306
rect 961 -1302 962 -1300
rect 961 -1308 962 -1306
rect 968 -1302 969 -1300
rect 968 -1308 969 -1306
rect 978 -1302 979 -1300
rect 975 -1308 976 -1306
rect 982 -1302 983 -1300
rect 982 -1308 983 -1306
rect 989 -1302 990 -1300
rect 989 -1308 990 -1306
rect 999 -1302 1000 -1300
rect 1003 -1302 1004 -1300
rect 1003 -1308 1004 -1306
rect 1010 -1302 1011 -1300
rect 1010 -1308 1011 -1306
rect 1017 -1302 1018 -1300
rect 1017 -1308 1018 -1306
rect 1020 -1308 1021 -1306
rect 1024 -1302 1025 -1300
rect 1027 -1302 1028 -1300
rect 1031 -1302 1032 -1300
rect 1031 -1308 1032 -1306
rect 1038 -1302 1039 -1300
rect 1038 -1308 1039 -1306
rect 1045 -1302 1046 -1300
rect 1045 -1308 1046 -1306
rect 1052 -1302 1053 -1300
rect 1052 -1308 1053 -1306
rect 1059 -1302 1060 -1300
rect 1062 -1302 1063 -1300
rect 1059 -1308 1060 -1306
rect 1066 -1302 1067 -1300
rect 1066 -1308 1067 -1306
rect 1080 -1302 1081 -1300
rect 1080 -1308 1081 -1306
rect 1087 -1302 1088 -1300
rect 1087 -1308 1088 -1306
rect 1097 -1302 1098 -1300
rect 1097 -1308 1098 -1306
rect 1101 -1302 1102 -1300
rect 1101 -1308 1102 -1306
rect 2 -1379 3 -1377
rect 9 -1373 10 -1371
rect 16 -1373 17 -1371
rect 16 -1379 17 -1377
rect 23 -1373 24 -1371
rect 23 -1379 24 -1377
rect 30 -1373 31 -1371
rect 30 -1379 31 -1377
rect 37 -1373 38 -1371
rect 37 -1379 38 -1377
rect 44 -1373 45 -1371
rect 44 -1379 45 -1377
rect 51 -1373 52 -1371
rect 51 -1379 52 -1377
rect 58 -1373 59 -1371
rect 58 -1379 59 -1377
rect 65 -1373 66 -1371
rect 68 -1373 69 -1371
rect 72 -1373 73 -1371
rect 72 -1379 73 -1377
rect 79 -1373 80 -1371
rect 79 -1379 80 -1377
rect 86 -1373 87 -1371
rect 86 -1379 87 -1377
rect 93 -1373 94 -1371
rect 93 -1379 94 -1377
rect 100 -1373 101 -1371
rect 107 -1373 108 -1371
rect 107 -1379 108 -1377
rect 114 -1373 115 -1371
rect 114 -1379 115 -1377
rect 121 -1373 122 -1371
rect 121 -1379 122 -1377
rect 128 -1373 129 -1371
rect 128 -1379 129 -1377
rect 135 -1373 136 -1371
rect 138 -1379 139 -1377
rect 142 -1373 143 -1371
rect 142 -1379 143 -1377
rect 149 -1373 150 -1371
rect 149 -1379 150 -1377
rect 156 -1373 157 -1371
rect 156 -1379 157 -1377
rect 163 -1373 164 -1371
rect 163 -1379 164 -1377
rect 170 -1373 171 -1371
rect 170 -1379 171 -1377
rect 177 -1373 178 -1371
rect 180 -1373 181 -1371
rect 184 -1373 185 -1371
rect 184 -1379 185 -1377
rect 191 -1373 192 -1371
rect 191 -1379 192 -1377
rect 198 -1373 199 -1371
rect 201 -1373 202 -1371
rect 201 -1379 202 -1377
rect 205 -1373 206 -1371
rect 205 -1379 206 -1377
rect 212 -1373 213 -1371
rect 212 -1379 213 -1377
rect 219 -1373 220 -1371
rect 219 -1379 220 -1377
rect 226 -1373 227 -1371
rect 226 -1379 227 -1377
rect 233 -1373 234 -1371
rect 233 -1379 234 -1377
rect 240 -1373 241 -1371
rect 240 -1379 241 -1377
rect 247 -1379 248 -1377
rect 250 -1379 251 -1377
rect 254 -1373 255 -1371
rect 254 -1379 255 -1377
rect 261 -1373 262 -1371
rect 261 -1379 262 -1377
rect 268 -1373 269 -1371
rect 268 -1379 269 -1377
rect 275 -1373 276 -1371
rect 278 -1373 279 -1371
rect 275 -1379 276 -1377
rect 285 -1373 286 -1371
rect 285 -1379 286 -1377
rect 289 -1373 290 -1371
rect 289 -1379 290 -1377
rect 296 -1373 297 -1371
rect 296 -1379 297 -1377
rect 303 -1373 304 -1371
rect 303 -1379 304 -1377
rect 310 -1373 311 -1371
rect 310 -1379 311 -1377
rect 317 -1373 318 -1371
rect 317 -1379 318 -1377
rect 324 -1373 325 -1371
rect 324 -1379 325 -1377
rect 331 -1373 332 -1371
rect 331 -1379 332 -1377
rect 338 -1373 339 -1371
rect 338 -1379 339 -1377
rect 345 -1373 346 -1371
rect 348 -1373 349 -1371
rect 345 -1379 346 -1377
rect 348 -1379 349 -1377
rect 352 -1373 353 -1371
rect 352 -1379 353 -1377
rect 359 -1373 360 -1371
rect 359 -1379 360 -1377
rect 366 -1373 367 -1371
rect 369 -1373 370 -1371
rect 366 -1379 367 -1377
rect 369 -1379 370 -1377
rect 373 -1373 374 -1371
rect 373 -1379 374 -1377
rect 380 -1373 381 -1371
rect 380 -1379 381 -1377
rect 387 -1373 388 -1371
rect 387 -1379 388 -1377
rect 394 -1373 395 -1371
rect 394 -1379 395 -1377
rect 401 -1373 402 -1371
rect 401 -1379 402 -1377
rect 408 -1373 409 -1371
rect 411 -1373 412 -1371
rect 408 -1379 409 -1377
rect 415 -1373 416 -1371
rect 415 -1379 416 -1377
rect 422 -1373 423 -1371
rect 422 -1379 423 -1377
rect 429 -1373 430 -1371
rect 429 -1379 430 -1377
rect 436 -1373 437 -1371
rect 439 -1373 440 -1371
rect 436 -1379 437 -1377
rect 443 -1373 444 -1371
rect 443 -1379 444 -1377
rect 450 -1373 451 -1371
rect 450 -1379 451 -1377
rect 457 -1373 458 -1371
rect 457 -1379 458 -1377
rect 464 -1373 465 -1371
rect 464 -1379 465 -1377
rect 471 -1373 472 -1371
rect 471 -1379 472 -1377
rect 478 -1373 479 -1371
rect 481 -1373 482 -1371
rect 485 -1373 486 -1371
rect 485 -1379 486 -1377
rect 492 -1379 493 -1377
rect 495 -1379 496 -1377
rect 499 -1373 500 -1371
rect 499 -1379 500 -1377
rect 506 -1373 507 -1371
rect 509 -1379 510 -1377
rect 513 -1373 514 -1371
rect 513 -1379 514 -1377
rect 520 -1373 521 -1371
rect 520 -1379 521 -1377
rect 527 -1373 528 -1371
rect 527 -1379 528 -1377
rect 534 -1373 535 -1371
rect 534 -1379 535 -1377
rect 541 -1373 542 -1371
rect 544 -1373 545 -1371
rect 541 -1379 542 -1377
rect 544 -1379 545 -1377
rect 548 -1373 549 -1371
rect 548 -1379 549 -1377
rect 555 -1373 556 -1371
rect 555 -1379 556 -1377
rect 562 -1373 563 -1371
rect 562 -1379 563 -1377
rect 569 -1373 570 -1371
rect 572 -1373 573 -1371
rect 569 -1379 570 -1377
rect 576 -1373 577 -1371
rect 576 -1379 577 -1377
rect 583 -1373 584 -1371
rect 583 -1379 584 -1377
rect 590 -1373 591 -1371
rect 590 -1379 591 -1377
rect 597 -1373 598 -1371
rect 597 -1379 598 -1377
rect 604 -1373 605 -1371
rect 604 -1379 605 -1377
rect 611 -1373 612 -1371
rect 611 -1379 612 -1377
rect 618 -1373 619 -1371
rect 618 -1379 619 -1377
rect 625 -1373 626 -1371
rect 628 -1373 629 -1371
rect 628 -1379 629 -1377
rect 632 -1373 633 -1371
rect 632 -1379 633 -1377
rect 639 -1373 640 -1371
rect 639 -1379 640 -1377
rect 646 -1373 647 -1371
rect 646 -1379 647 -1377
rect 653 -1373 654 -1371
rect 653 -1379 654 -1377
rect 656 -1379 657 -1377
rect 660 -1373 661 -1371
rect 663 -1379 664 -1377
rect 667 -1373 668 -1371
rect 667 -1379 668 -1377
rect 674 -1373 675 -1371
rect 674 -1379 675 -1377
rect 681 -1373 682 -1371
rect 681 -1379 682 -1377
rect 688 -1373 689 -1371
rect 688 -1379 689 -1377
rect 695 -1373 696 -1371
rect 695 -1379 696 -1377
rect 702 -1373 703 -1371
rect 702 -1379 703 -1377
rect 709 -1373 710 -1371
rect 709 -1379 710 -1377
rect 716 -1373 717 -1371
rect 716 -1379 717 -1377
rect 723 -1373 724 -1371
rect 726 -1373 727 -1371
rect 723 -1379 724 -1377
rect 726 -1379 727 -1377
rect 730 -1373 731 -1371
rect 733 -1373 734 -1371
rect 737 -1373 738 -1371
rect 737 -1379 738 -1377
rect 744 -1373 745 -1371
rect 744 -1379 745 -1377
rect 751 -1373 752 -1371
rect 751 -1379 752 -1377
rect 758 -1373 759 -1371
rect 758 -1379 759 -1377
rect 765 -1373 766 -1371
rect 765 -1379 766 -1377
rect 772 -1373 773 -1371
rect 772 -1379 773 -1377
rect 779 -1373 780 -1371
rect 779 -1379 780 -1377
rect 786 -1373 787 -1371
rect 786 -1379 787 -1377
rect 793 -1373 794 -1371
rect 793 -1379 794 -1377
rect 800 -1373 801 -1371
rect 800 -1379 801 -1377
rect 807 -1373 808 -1371
rect 807 -1379 808 -1377
rect 814 -1373 815 -1371
rect 814 -1379 815 -1377
rect 821 -1373 822 -1371
rect 821 -1379 822 -1377
rect 828 -1373 829 -1371
rect 828 -1379 829 -1377
rect 835 -1373 836 -1371
rect 835 -1379 836 -1377
rect 842 -1373 843 -1371
rect 842 -1379 843 -1377
rect 849 -1373 850 -1371
rect 849 -1379 850 -1377
rect 856 -1373 857 -1371
rect 856 -1379 857 -1377
rect 863 -1373 864 -1371
rect 863 -1379 864 -1377
rect 870 -1373 871 -1371
rect 870 -1379 871 -1377
rect 877 -1373 878 -1371
rect 877 -1379 878 -1377
rect 884 -1373 885 -1371
rect 884 -1379 885 -1377
rect 891 -1373 892 -1371
rect 891 -1379 892 -1377
rect 898 -1373 899 -1371
rect 898 -1379 899 -1377
rect 905 -1373 906 -1371
rect 905 -1379 906 -1377
rect 912 -1373 913 -1371
rect 912 -1379 913 -1377
rect 919 -1373 920 -1371
rect 919 -1379 920 -1377
rect 926 -1373 927 -1371
rect 926 -1379 927 -1377
rect 933 -1373 934 -1371
rect 933 -1379 934 -1377
rect 940 -1373 941 -1371
rect 940 -1379 941 -1377
rect 947 -1373 948 -1371
rect 947 -1379 948 -1377
rect 954 -1373 955 -1371
rect 954 -1379 955 -1377
rect 961 -1373 962 -1371
rect 961 -1379 962 -1377
rect 968 -1373 969 -1371
rect 968 -1379 969 -1377
rect 975 -1373 976 -1371
rect 975 -1379 976 -1377
rect 982 -1373 983 -1371
rect 982 -1379 983 -1377
rect 989 -1373 990 -1371
rect 989 -1379 990 -1377
rect 996 -1373 997 -1371
rect 999 -1373 1000 -1371
rect 996 -1379 997 -1377
rect 1003 -1373 1004 -1371
rect 1003 -1379 1004 -1377
rect 1010 -1373 1011 -1371
rect 1010 -1379 1011 -1377
rect 1017 -1373 1018 -1371
rect 1017 -1379 1018 -1377
rect 1024 -1373 1025 -1371
rect 1031 -1373 1032 -1371
rect 1031 -1379 1032 -1377
rect 1066 -1373 1067 -1371
rect 1066 -1379 1067 -1377
rect 5 -1448 6 -1446
rect 9 -1448 10 -1446
rect 9 -1454 10 -1452
rect 19 -1454 20 -1452
rect 23 -1448 24 -1446
rect 23 -1454 24 -1452
rect 30 -1448 31 -1446
rect 30 -1454 31 -1452
rect 37 -1454 38 -1452
rect 40 -1454 41 -1452
rect 44 -1448 45 -1446
rect 44 -1454 45 -1452
rect 51 -1448 52 -1446
rect 51 -1454 52 -1452
rect 58 -1448 59 -1446
rect 58 -1454 59 -1452
rect 68 -1454 69 -1452
rect 72 -1448 73 -1446
rect 72 -1454 73 -1452
rect 79 -1448 80 -1446
rect 79 -1454 80 -1452
rect 86 -1448 87 -1446
rect 86 -1454 87 -1452
rect 93 -1448 94 -1446
rect 93 -1454 94 -1452
rect 100 -1448 101 -1446
rect 100 -1454 101 -1452
rect 107 -1448 108 -1446
rect 107 -1454 108 -1452
rect 114 -1448 115 -1446
rect 114 -1454 115 -1452
rect 121 -1448 122 -1446
rect 121 -1454 122 -1452
rect 128 -1448 129 -1446
rect 128 -1454 129 -1452
rect 135 -1448 136 -1446
rect 135 -1454 136 -1452
rect 138 -1454 139 -1452
rect 142 -1448 143 -1446
rect 142 -1454 143 -1452
rect 149 -1448 150 -1446
rect 149 -1454 150 -1452
rect 156 -1448 157 -1446
rect 156 -1454 157 -1452
rect 163 -1448 164 -1446
rect 163 -1454 164 -1452
rect 170 -1448 171 -1446
rect 170 -1454 171 -1452
rect 177 -1448 178 -1446
rect 177 -1454 178 -1452
rect 184 -1448 185 -1446
rect 184 -1454 185 -1452
rect 191 -1454 192 -1452
rect 194 -1454 195 -1452
rect 198 -1448 199 -1446
rect 198 -1454 199 -1452
rect 205 -1448 206 -1446
rect 208 -1448 209 -1446
rect 215 -1454 216 -1452
rect 219 -1448 220 -1446
rect 219 -1454 220 -1452
rect 226 -1448 227 -1446
rect 226 -1454 227 -1452
rect 233 -1448 234 -1446
rect 233 -1454 234 -1452
rect 240 -1448 241 -1446
rect 240 -1454 241 -1452
rect 247 -1448 248 -1446
rect 247 -1454 248 -1452
rect 254 -1448 255 -1446
rect 254 -1454 255 -1452
rect 261 -1448 262 -1446
rect 261 -1454 262 -1452
rect 268 -1448 269 -1446
rect 268 -1454 269 -1452
rect 275 -1454 276 -1452
rect 278 -1454 279 -1452
rect 285 -1454 286 -1452
rect 289 -1448 290 -1446
rect 289 -1454 290 -1452
rect 296 -1448 297 -1446
rect 296 -1454 297 -1452
rect 303 -1448 304 -1446
rect 303 -1454 304 -1452
rect 310 -1448 311 -1446
rect 310 -1454 311 -1452
rect 324 -1448 325 -1446
rect 324 -1454 325 -1452
rect 331 -1448 332 -1446
rect 331 -1454 332 -1452
rect 338 -1448 339 -1446
rect 338 -1454 339 -1452
rect 345 -1448 346 -1446
rect 345 -1454 346 -1452
rect 352 -1448 353 -1446
rect 352 -1454 353 -1452
rect 359 -1448 360 -1446
rect 359 -1454 360 -1452
rect 366 -1448 367 -1446
rect 369 -1448 370 -1446
rect 366 -1454 367 -1452
rect 373 -1448 374 -1446
rect 376 -1448 377 -1446
rect 373 -1454 374 -1452
rect 376 -1454 377 -1452
rect 380 -1448 381 -1446
rect 380 -1454 381 -1452
rect 387 -1448 388 -1446
rect 387 -1454 388 -1452
rect 394 -1448 395 -1446
rect 394 -1454 395 -1452
rect 401 -1448 402 -1446
rect 401 -1454 402 -1452
rect 408 -1448 409 -1446
rect 408 -1454 409 -1452
rect 415 -1448 416 -1446
rect 415 -1454 416 -1452
rect 422 -1448 423 -1446
rect 422 -1454 423 -1452
rect 425 -1454 426 -1452
rect 429 -1448 430 -1446
rect 429 -1454 430 -1452
rect 436 -1448 437 -1446
rect 439 -1448 440 -1446
rect 436 -1454 437 -1452
rect 443 -1448 444 -1446
rect 443 -1454 444 -1452
rect 450 -1448 451 -1446
rect 450 -1454 451 -1452
rect 460 -1448 461 -1446
rect 457 -1454 458 -1452
rect 460 -1454 461 -1452
rect 464 -1448 465 -1446
rect 464 -1454 465 -1452
rect 474 -1448 475 -1446
rect 471 -1454 472 -1452
rect 474 -1454 475 -1452
rect 478 -1448 479 -1446
rect 478 -1454 479 -1452
rect 485 -1448 486 -1446
rect 488 -1448 489 -1446
rect 488 -1454 489 -1452
rect 492 -1448 493 -1446
rect 492 -1454 493 -1452
rect 499 -1448 500 -1446
rect 499 -1454 500 -1452
rect 506 -1448 507 -1446
rect 506 -1454 507 -1452
rect 513 -1448 514 -1446
rect 513 -1454 514 -1452
rect 520 -1448 521 -1446
rect 523 -1448 524 -1446
rect 520 -1454 521 -1452
rect 527 -1448 528 -1446
rect 530 -1448 531 -1446
rect 527 -1454 528 -1452
rect 534 -1448 535 -1446
rect 537 -1448 538 -1446
rect 537 -1454 538 -1452
rect 541 -1448 542 -1446
rect 541 -1454 542 -1452
rect 548 -1448 549 -1446
rect 548 -1454 549 -1452
rect 555 -1448 556 -1446
rect 555 -1454 556 -1452
rect 562 -1448 563 -1446
rect 562 -1454 563 -1452
rect 569 -1448 570 -1446
rect 569 -1454 570 -1452
rect 576 -1448 577 -1446
rect 576 -1454 577 -1452
rect 583 -1448 584 -1446
rect 583 -1454 584 -1452
rect 590 -1448 591 -1446
rect 590 -1454 591 -1452
rect 597 -1448 598 -1446
rect 597 -1454 598 -1452
rect 607 -1454 608 -1452
rect 611 -1448 612 -1446
rect 611 -1454 612 -1452
rect 618 -1448 619 -1446
rect 618 -1454 619 -1452
rect 625 -1448 626 -1446
rect 625 -1454 626 -1452
rect 635 -1454 636 -1452
rect 639 -1448 640 -1446
rect 639 -1454 640 -1452
rect 642 -1454 643 -1452
rect 646 -1448 647 -1446
rect 646 -1454 647 -1452
rect 653 -1448 654 -1446
rect 653 -1454 654 -1452
rect 660 -1448 661 -1446
rect 660 -1454 661 -1452
rect 667 -1448 668 -1446
rect 667 -1454 668 -1452
rect 674 -1448 675 -1446
rect 674 -1454 675 -1452
rect 681 -1448 682 -1446
rect 681 -1454 682 -1452
rect 688 -1448 689 -1446
rect 688 -1454 689 -1452
rect 695 -1448 696 -1446
rect 695 -1454 696 -1452
rect 702 -1448 703 -1446
rect 702 -1454 703 -1452
rect 709 -1448 710 -1446
rect 709 -1454 710 -1452
rect 716 -1448 717 -1446
rect 723 -1448 724 -1446
rect 723 -1454 724 -1452
rect 730 -1448 731 -1446
rect 730 -1454 731 -1452
rect 737 -1448 738 -1446
rect 737 -1454 738 -1452
rect 744 -1448 745 -1446
rect 744 -1454 745 -1452
rect 747 -1454 748 -1452
rect 751 -1448 752 -1446
rect 751 -1454 752 -1452
rect 758 -1448 759 -1446
rect 758 -1454 759 -1452
rect 765 -1454 766 -1452
rect 768 -1454 769 -1452
rect 772 -1448 773 -1446
rect 772 -1454 773 -1452
rect 779 -1448 780 -1446
rect 779 -1454 780 -1452
rect 786 -1448 787 -1446
rect 786 -1454 787 -1452
rect 793 -1448 794 -1446
rect 796 -1448 797 -1446
rect 793 -1454 794 -1452
rect 796 -1454 797 -1452
rect 800 -1448 801 -1446
rect 800 -1454 801 -1452
rect 807 -1448 808 -1446
rect 807 -1454 808 -1452
rect 814 -1448 815 -1446
rect 814 -1454 815 -1452
rect 821 -1448 822 -1446
rect 824 -1454 825 -1452
rect 828 -1448 829 -1446
rect 828 -1454 829 -1452
rect 835 -1448 836 -1446
rect 835 -1454 836 -1452
rect 842 -1448 843 -1446
rect 842 -1454 843 -1452
rect 849 -1448 850 -1446
rect 849 -1454 850 -1452
rect 856 -1448 857 -1446
rect 856 -1454 857 -1452
rect 863 -1448 864 -1446
rect 863 -1454 864 -1452
rect 870 -1448 871 -1446
rect 870 -1454 871 -1452
rect 877 -1448 878 -1446
rect 877 -1454 878 -1452
rect 884 -1448 885 -1446
rect 884 -1454 885 -1452
rect 891 -1448 892 -1446
rect 891 -1454 892 -1452
rect 898 -1448 899 -1446
rect 898 -1454 899 -1452
rect 905 -1448 906 -1446
rect 905 -1454 906 -1452
rect 912 -1448 913 -1446
rect 912 -1454 913 -1452
rect 919 -1448 920 -1446
rect 919 -1454 920 -1452
rect 926 -1448 927 -1446
rect 926 -1454 927 -1452
rect 933 -1448 934 -1446
rect 933 -1454 934 -1452
rect 940 -1448 941 -1446
rect 940 -1454 941 -1452
rect 947 -1448 948 -1446
rect 947 -1454 948 -1452
rect 954 -1448 955 -1446
rect 954 -1454 955 -1452
rect 961 -1448 962 -1446
rect 961 -1454 962 -1452
rect 968 -1448 969 -1446
rect 968 -1454 969 -1452
rect 975 -1448 976 -1446
rect 975 -1454 976 -1452
rect 982 -1448 983 -1446
rect 982 -1454 983 -1452
rect 989 -1448 990 -1446
rect 989 -1454 990 -1452
rect 996 -1448 997 -1446
rect 996 -1454 997 -1452
rect 1003 -1448 1004 -1446
rect 1003 -1454 1004 -1452
rect 1010 -1448 1011 -1446
rect 1010 -1454 1011 -1452
rect 1017 -1448 1018 -1446
rect 1017 -1454 1018 -1452
rect 1024 -1448 1025 -1446
rect 1024 -1454 1025 -1452
rect 1031 -1448 1032 -1446
rect 1031 -1454 1032 -1452
rect 1038 -1448 1039 -1446
rect 1038 -1454 1039 -1452
rect 1045 -1448 1046 -1446
rect 1048 -1448 1049 -1446
rect 1048 -1454 1049 -1452
rect 1052 -1448 1053 -1446
rect 1055 -1448 1056 -1446
rect 1059 -1448 1060 -1446
rect 1059 -1454 1060 -1452
rect 1066 -1448 1067 -1446
rect 1066 -1454 1067 -1452
rect 2 -1531 3 -1529
rect 2 -1537 3 -1535
rect 16 -1531 17 -1529
rect 16 -1537 17 -1535
rect 23 -1531 24 -1529
rect 23 -1537 24 -1535
rect 30 -1531 31 -1529
rect 30 -1537 31 -1535
rect 37 -1531 38 -1529
rect 37 -1537 38 -1535
rect 44 -1531 45 -1529
rect 44 -1537 45 -1535
rect 51 -1531 52 -1529
rect 51 -1537 52 -1535
rect 58 -1531 59 -1529
rect 58 -1537 59 -1535
rect 68 -1531 69 -1529
rect 68 -1537 69 -1535
rect 72 -1531 73 -1529
rect 72 -1537 73 -1535
rect 79 -1531 80 -1529
rect 79 -1537 80 -1535
rect 86 -1531 87 -1529
rect 86 -1537 87 -1535
rect 93 -1531 94 -1529
rect 96 -1531 97 -1529
rect 100 -1531 101 -1529
rect 100 -1537 101 -1535
rect 107 -1531 108 -1529
rect 107 -1537 108 -1535
rect 114 -1531 115 -1529
rect 114 -1537 115 -1535
rect 117 -1537 118 -1535
rect 121 -1531 122 -1529
rect 121 -1537 122 -1535
rect 128 -1531 129 -1529
rect 128 -1537 129 -1535
rect 135 -1531 136 -1529
rect 135 -1537 136 -1535
rect 142 -1531 143 -1529
rect 142 -1537 143 -1535
rect 149 -1531 150 -1529
rect 149 -1537 150 -1535
rect 156 -1531 157 -1529
rect 156 -1537 157 -1535
rect 163 -1531 164 -1529
rect 163 -1537 164 -1535
rect 170 -1531 171 -1529
rect 170 -1537 171 -1535
rect 177 -1531 178 -1529
rect 177 -1537 178 -1535
rect 184 -1531 185 -1529
rect 184 -1537 185 -1535
rect 191 -1531 192 -1529
rect 191 -1537 192 -1535
rect 198 -1531 199 -1529
rect 201 -1537 202 -1535
rect 205 -1531 206 -1529
rect 205 -1537 206 -1535
rect 212 -1531 213 -1529
rect 212 -1537 213 -1535
rect 219 -1531 220 -1529
rect 219 -1537 220 -1535
rect 226 -1531 227 -1529
rect 226 -1537 227 -1535
rect 233 -1531 234 -1529
rect 233 -1537 234 -1535
rect 240 -1531 241 -1529
rect 240 -1537 241 -1535
rect 247 -1531 248 -1529
rect 247 -1537 248 -1535
rect 254 -1531 255 -1529
rect 254 -1537 255 -1535
rect 261 -1531 262 -1529
rect 261 -1537 262 -1535
rect 268 -1531 269 -1529
rect 268 -1537 269 -1535
rect 275 -1531 276 -1529
rect 275 -1537 276 -1535
rect 282 -1531 283 -1529
rect 282 -1537 283 -1535
rect 289 -1531 290 -1529
rect 289 -1537 290 -1535
rect 296 -1531 297 -1529
rect 296 -1537 297 -1535
rect 303 -1531 304 -1529
rect 303 -1537 304 -1535
rect 310 -1531 311 -1529
rect 310 -1537 311 -1535
rect 317 -1531 318 -1529
rect 317 -1537 318 -1535
rect 324 -1531 325 -1529
rect 324 -1537 325 -1535
rect 331 -1531 332 -1529
rect 331 -1537 332 -1535
rect 338 -1531 339 -1529
rect 338 -1537 339 -1535
rect 348 -1531 349 -1529
rect 352 -1531 353 -1529
rect 355 -1537 356 -1535
rect 359 -1531 360 -1529
rect 359 -1537 360 -1535
rect 366 -1531 367 -1529
rect 366 -1537 367 -1535
rect 373 -1531 374 -1529
rect 373 -1537 374 -1535
rect 380 -1531 381 -1529
rect 380 -1537 381 -1535
rect 387 -1531 388 -1529
rect 387 -1537 388 -1535
rect 394 -1531 395 -1529
rect 394 -1537 395 -1535
rect 401 -1531 402 -1529
rect 401 -1537 402 -1535
rect 408 -1531 409 -1529
rect 408 -1537 409 -1535
rect 411 -1537 412 -1535
rect 415 -1531 416 -1529
rect 415 -1537 416 -1535
rect 422 -1531 423 -1529
rect 422 -1537 423 -1535
rect 429 -1531 430 -1529
rect 429 -1537 430 -1535
rect 436 -1531 437 -1529
rect 436 -1537 437 -1535
rect 443 -1531 444 -1529
rect 443 -1537 444 -1535
rect 450 -1531 451 -1529
rect 450 -1537 451 -1535
rect 457 -1531 458 -1529
rect 457 -1537 458 -1535
rect 464 -1531 465 -1529
rect 471 -1531 472 -1529
rect 471 -1537 472 -1535
rect 478 -1531 479 -1529
rect 478 -1537 479 -1535
rect 488 -1531 489 -1529
rect 488 -1537 489 -1535
rect 492 -1531 493 -1529
rect 492 -1537 493 -1535
rect 499 -1531 500 -1529
rect 499 -1537 500 -1535
rect 506 -1531 507 -1529
rect 509 -1531 510 -1529
rect 509 -1537 510 -1535
rect 516 -1531 517 -1529
rect 513 -1537 514 -1535
rect 520 -1531 521 -1529
rect 523 -1531 524 -1529
rect 520 -1537 521 -1535
rect 527 -1537 528 -1535
rect 534 -1531 535 -1529
rect 537 -1531 538 -1529
rect 537 -1537 538 -1535
rect 541 -1531 542 -1529
rect 544 -1531 545 -1529
rect 548 -1531 549 -1529
rect 548 -1537 549 -1535
rect 555 -1531 556 -1529
rect 555 -1537 556 -1535
rect 565 -1531 566 -1529
rect 565 -1537 566 -1535
rect 569 -1531 570 -1529
rect 569 -1537 570 -1535
rect 576 -1531 577 -1529
rect 576 -1537 577 -1535
rect 583 -1531 584 -1529
rect 583 -1537 584 -1535
rect 590 -1531 591 -1529
rect 593 -1531 594 -1529
rect 590 -1537 591 -1535
rect 597 -1531 598 -1529
rect 597 -1537 598 -1535
rect 604 -1531 605 -1529
rect 611 -1531 612 -1529
rect 611 -1537 612 -1535
rect 618 -1537 619 -1535
rect 625 -1531 626 -1529
rect 625 -1537 626 -1535
rect 632 -1531 633 -1529
rect 632 -1537 633 -1535
rect 639 -1531 640 -1529
rect 639 -1537 640 -1535
rect 646 -1531 647 -1529
rect 646 -1537 647 -1535
rect 653 -1531 654 -1529
rect 653 -1537 654 -1535
rect 660 -1531 661 -1529
rect 660 -1537 661 -1535
rect 663 -1537 664 -1535
rect 667 -1531 668 -1529
rect 667 -1537 668 -1535
rect 674 -1531 675 -1529
rect 674 -1537 675 -1535
rect 681 -1531 682 -1529
rect 684 -1531 685 -1529
rect 684 -1537 685 -1535
rect 688 -1531 689 -1529
rect 688 -1537 689 -1535
rect 695 -1531 696 -1529
rect 695 -1537 696 -1535
rect 702 -1531 703 -1529
rect 702 -1537 703 -1535
rect 709 -1531 710 -1529
rect 709 -1537 710 -1535
rect 716 -1537 717 -1535
rect 723 -1531 724 -1529
rect 726 -1531 727 -1529
rect 726 -1537 727 -1535
rect 730 -1531 731 -1529
rect 730 -1537 731 -1535
rect 740 -1531 741 -1529
rect 737 -1537 738 -1535
rect 740 -1537 741 -1535
rect 744 -1531 745 -1529
rect 747 -1531 748 -1529
rect 744 -1537 745 -1535
rect 751 -1531 752 -1529
rect 751 -1537 752 -1535
rect 758 -1531 759 -1529
rect 758 -1537 759 -1535
rect 765 -1531 766 -1529
rect 765 -1537 766 -1535
rect 772 -1531 773 -1529
rect 772 -1537 773 -1535
rect 779 -1531 780 -1529
rect 779 -1537 780 -1535
rect 786 -1531 787 -1529
rect 786 -1537 787 -1535
rect 793 -1531 794 -1529
rect 793 -1537 794 -1535
rect 800 -1531 801 -1529
rect 800 -1537 801 -1535
rect 807 -1531 808 -1529
rect 807 -1537 808 -1535
rect 814 -1531 815 -1529
rect 814 -1537 815 -1535
rect 821 -1531 822 -1529
rect 821 -1537 822 -1535
rect 828 -1531 829 -1529
rect 828 -1537 829 -1535
rect 835 -1531 836 -1529
rect 835 -1537 836 -1535
rect 842 -1531 843 -1529
rect 845 -1531 846 -1529
rect 849 -1531 850 -1529
rect 849 -1537 850 -1535
rect 856 -1531 857 -1529
rect 856 -1537 857 -1535
rect 863 -1531 864 -1529
rect 863 -1537 864 -1535
rect 870 -1531 871 -1529
rect 870 -1537 871 -1535
rect 877 -1531 878 -1529
rect 877 -1537 878 -1535
rect 884 -1531 885 -1529
rect 884 -1537 885 -1535
rect 891 -1531 892 -1529
rect 891 -1537 892 -1535
rect 898 -1531 899 -1529
rect 898 -1537 899 -1535
rect 905 -1531 906 -1529
rect 905 -1537 906 -1535
rect 912 -1531 913 -1529
rect 912 -1537 913 -1535
rect 919 -1531 920 -1529
rect 919 -1537 920 -1535
rect 926 -1531 927 -1529
rect 926 -1537 927 -1535
rect 933 -1531 934 -1529
rect 933 -1537 934 -1535
rect 940 -1531 941 -1529
rect 940 -1537 941 -1535
rect 947 -1531 948 -1529
rect 947 -1537 948 -1535
rect 954 -1531 955 -1529
rect 954 -1537 955 -1535
rect 961 -1531 962 -1529
rect 961 -1537 962 -1535
rect 968 -1531 969 -1529
rect 968 -1537 969 -1535
rect 975 -1531 976 -1529
rect 975 -1537 976 -1535
rect 982 -1531 983 -1529
rect 982 -1537 983 -1535
rect 989 -1531 990 -1529
rect 989 -1537 990 -1535
rect 996 -1531 997 -1529
rect 999 -1531 1000 -1529
rect 996 -1537 997 -1535
rect 1003 -1531 1004 -1529
rect 1003 -1537 1004 -1535
rect 1010 -1531 1011 -1529
rect 1010 -1537 1011 -1535
rect 1017 -1531 1018 -1529
rect 1017 -1537 1018 -1535
rect 1045 -1531 1046 -1529
rect 1045 -1537 1046 -1535
rect 1052 -1531 1053 -1529
rect 1052 -1537 1053 -1535
rect 1059 -1531 1060 -1529
rect 23 -1608 24 -1606
rect 23 -1614 24 -1612
rect 30 -1608 31 -1606
rect 30 -1614 31 -1612
rect 37 -1608 38 -1606
rect 37 -1614 38 -1612
rect 44 -1608 45 -1606
rect 44 -1614 45 -1612
rect 51 -1608 52 -1606
rect 51 -1614 52 -1612
rect 58 -1608 59 -1606
rect 58 -1614 59 -1612
rect 68 -1608 69 -1606
rect 68 -1614 69 -1612
rect 72 -1608 73 -1606
rect 79 -1608 80 -1606
rect 79 -1614 80 -1612
rect 86 -1608 87 -1606
rect 86 -1614 87 -1612
rect 93 -1608 94 -1606
rect 93 -1614 94 -1612
rect 100 -1608 101 -1606
rect 100 -1614 101 -1612
rect 107 -1608 108 -1606
rect 107 -1614 108 -1612
rect 110 -1614 111 -1612
rect 114 -1608 115 -1606
rect 114 -1614 115 -1612
rect 121 -1608 122 -1606
rect 121 -1614 122 -1612
rect 128 -1608 129 -1606
rect 128 -1614 129 -1612
rect 135 -1608 136 -1606
rect 135 -1614 136 -1612
rect 142 -1608 143 -1606
rect 142 -1614 143 -1612
rect 152 -1608 153 -1606
rect 152 -1614 153 -1612
rect 156 -1608 157 -1606
rect 156 -1614 157 -1612
rect 159 -1614 160 -1612
rect 163 -1608 164 -1606
rect 163 -1614 164 -1612
rect 173 -1608 174 -1606
rect 170 -1614 171 -1612
rect 177 -1608 178 -1606
rect 177 -1614 178 -1612
rect 184 -1608 185 -1606
rect 184 -1614 185 -1612
rect 191 -1608 192 -1606
rect 191 -1614 192 -1612
rect 198 -1614 199 -1612
rect 201 -1614 202 -1612
rect 205 -1608 206 -1606
rect 205 -1614 206 -1612
rect 212 -1608 213 -1606
rect 212 -1614 213 -1612
rect 219 -1608 220 -1606
rect 219 -1614 220 -1612
rect 226 -1614 227 -1612
rect 229 -1614 230 -1612
rect 233 -1608 234 -1606
rect 233 -1614 234 -1612
rect 240 -1608 241 -1606
rect 240 -1614 241 -1612
rect 247 -1608 248 -1606
rect 247 -1614 248 -1612
rect 254 -1608 255 -1606
rect 254 -1614 255 -1612
rect 261 -1608 262 -1606
rect 261 -1614 262 -1612
rect 268 -1608 269 -1606
rect 268 -1614 269 -1612
rect 275 -1608 276 -1606
rect 275 -1614 276 -1612
rect 282 -1608 283 -1606
rect 282 -1614 283 -1612
rect 289 -1608 290 -1606
rect 289 -1614 290 -1612
rect 296 -1608 297 -1606
rect 296 -1614 297 -1612
rect 306 -1608 307 -1606
rect 303 -1614 304 -1612
rect 306 -1614 307 -1612
rect 313 -1608 314 -1606
rect 310 -1614 311 -1612
rect 313 -1614 314 -1612
rect 317 -1608 318 -1606
rect 317 -1614 318 -1612
rect 324 -1608 325 -1606
rect 324 -1614 325 -1612
rect 331 -1608 332 -1606
rect 331 -1614 332 -1612
rect 338 -1608 339 -1606
rect 338 -1614 339 -1612
rect 345 -1608 346 -1606
rect 345 -1614 346 -1612
rect 355 -1608 356 -1606
rect 352 -1614 353 -1612
rect 355 -1614 356 -1612
rect 359 -1608 360 -1606
rect 359 -1614 360 -1612
rect 366 -1608 367 -1606
rect 366 -1614 367 -1612
rect 373 -1608 374 -1606
rect 373 -1614 374 -1612
rect 376 -1614 377 -1612
rect 380 -1608 381 -1606
rect 380 -1614 381 -1612
rect 387 -1608 388 -1606
rect 390 -1614 391 -1612
rect 394 -1608 395 -1606
rect 394 -1614 395 -1612
rect 401 -1608 402 -1606
rect 401 -1614 402 -1612
rect 408 -1608 409 -1606
rect 408 -1614 409 -1612
rect 415 -1608 416 -1606
rect 415 -1614 416 -1612
rect 425 -1608 426 -1606
rect 422 -1614 423 -1612
rect 425 -1614 426 -1612
rect 429 -1608 430 -1606
rect 429 -1614 430 -1612
rect 436 -1608 437 -1606
rect 436 -1614 437 -1612
rect 443 -1608 444 -1606
rect 443 -1614 444 -1612
rect 450 -1608 451 -1606
rect 450 -1614 451 -1612
rect 457 -1608 458 -1606
rect 457 -1614 458 -1612
rect 464 -1608 465 -1606
rect 464 -1614 465 -1612
rect 471 -1608 472 -1606
rect 471 -1614 472 -1612
rect 478 -1608 479 -1606
rect 478 -1614 479 -1612
rect 485 -1608 486 -1606
rect 485 -1614 486 -1612
rect 492 -1608 493 -1606
rect 492 -1614 493 -1612
rect 499 -1608 500 -1606
rect 499 -1614 500 -1612
rect 506 -1608 507 -1606
rect 506 -1614 507 -1612
rect 513 -1608 514 -1606
rect 513 -1614 514 -1612
rect 523 -1614 524 -1612
rect 530 -1608 531 -1606
rect 530 -1614 531 -1612
rect 534 -1608 535 -1606
rect 534 -1614 535 -1612
rect 541 -1608 542 -1606
rect 541 -1614 542 -1612
rect 548 -1608 549 -1606
rect 548 -1614 549 -1612
rect 555 -1608 556 -1606
rect 558 -1608 559 -1606
rect 555 -1614 556 -1612
rect 562 -1608 563 -1606
rect 565 -1608 566 -1606
rect 562 -1614 563 -1612
rect 565 -1614 566 -1612
rect 572 -1608 573 -1606
rect 569 -1614 570 -1612
rect 576 -1608 577 -1606
rect 576 -1614 577 -1612
rect 583 -1608 584 -1606
rect 583 -1614 584 -1612
rect 590 -1608 591 -1606
rect 590 -1614 591 -1612
rect 597 -1608 598 -1606
rect 597 -1614 598 -1612
rect 604 -1608 605 -1606
rect 604 -1614 605 -1612
rect 614 -1614 615 -1612
rect 618 -1608 619 -1606
rect 618 -1614 619 -1612
rect 628 -1608 629 -1606
rect 632 -1608 633 -1606
rect 632 -1614 633 -1612
rect 639 -1608 640 -1606
rect 639 -1614 640 -1612
rect 646 -1608 647 -1606
rect 646 -1614 647 -1612
rect 653 -1608 654 -1606
rect 653 -1614 654 -1612
rect 660 -1608 661 -1606
rect 660 -1614 661 -1612
rect 667 -1608 668 -1606
rect 667 -1614 668 -1612
rect 674 -1608 675 -1606
rect 674 -1614 675 -1612
rect 681 -1614 682 -1612
rect 684 -1614 685 -1612
rect 688 -1608 689 -1606
rect 688 -1614 689 -1612
rect 695 -1608 696 -1606
rect 695 -1614 696 -1612
rect 702 -1608 703 -1606
rect 702 -1614 703 -1612
rect 709 -1608 710 -1606
rect 709 -1614 710 -1612
rect 716 -1608 717 -1606
rect 716 -1614 717 -1612
rect 723 -1608 724 -1606
rect 723 -1614 724 -1612
rect 730 -1608 731 -1606
rect 730 -1614 731 -1612
rect 737 -1608 738 -1606
rect 737 -1614 738 -1612
rect 744 -1608 745 -1606
rect 744 -1614 745 -1612
rect 751 -1608 752 -1606
rect 751 -1614 752 -1612
rect 758 -1608 759 -1606
rect 758 -1614 759 -1612
rect 765 -1608 766 -1606
rect 765 -1614 766 -1612
rect 772 -1608 773 -1606
rect 772 -1614 773 -1612
rect 779 -1608 780 -1606
rect 779 -1614 780 -1612
rect 786 -1608 787 -1606
rect 786 -1614 787 -1612
rect 793 -1608 794 -1606
rect 793 -1614 794 -1612
rect 800 -1608 801 -1606
rect 800 -1614 801 -1612
rect 807 -1608 808 -1606
rect 807 -1614 808 -1612
rect 814 -1608 815 -1606
rect 814 -1614 815 -1612
rect 821 -1608 822 -1606
rect 821 -1614 822 -1612
rect 828 -1608 829 -1606
rect 828 -1614 829 -1612
rect 835 -1608 836 -1606
rect 835 -1614 836 -1612
rect 842 -1608 843 -1606
rect 842 -1614 843 -1612
rect 849 -1608 850 -1606
rect 849 -1614 850 -1612
rect 856 -1608 857 -1606
rect 859 -1614 860 -1612
rect 863 -1608 864 -1606
rect 863 -1614 864 -1612
rect 870 -1608 871 -1606
rect 870 -1614 871 -1612
rect 877 -1608 878 -1606
rect 877 -1614 878 -1612
rect 884 -1608 885 -1606
rect 884 -1614 885 -1612
rect 891 -1608 892 -1606
rect 891 -1614 892 -1612
rect 898 -1608 899 -1606
rect 898 -1614 899 -1612
rect 905 -1608 906 -1606
rect 905 -1614 906 -1612
rect 912 -1608 913 -1606
rect 912 -1614 913 -1612
rect 919 -1608 920 -1606
rect 919 -1614 920 -1612
rect 926 -1608 927 -1606
rect 926 -1614 927 -1612
rect 936 -1608 937 -1606
rect 936 -1614 937 -1612
rect 940 -1608 941 -1606
rect 940 -1614 941 -1612
rect 947 -1608 948 -1606
rect 947 -1614 948 -1612
rect 954 -1608 955 -1606
rect 954 -1614 955 -1612
rect 961 -1608 962 -1606
rect 961 -1614 962 -1612
rect 1024 -1608 1025 -1606
rect 1024 -1614 1025 -1612
rect 1038 -1608 1039 -1606
rect 1038 -1614 1039 -1612
rect 1045 -1614 1046 -1612
rect 1052 -1608 1053 -1606
rect 37 -1673 38 -1671
rect 40 -1673 41 -1671
rect 44 -1673 45 -1671
rect 47 -1679 48 -1677
rect 51 -1673 52 -1671
rect 51 -1679 52 -1677
rect 65 -1673 66 -1671
rect 65 -1679 66 -1677
rect 72 -1673 73 -1671
rect 75 -1679 76 -1677
rect 79 -1673 80 -1671
rect 86 -1673 87 -1671
rect 86 -1679 87 -1677
rect 93 -1673 94 -1671
rect 93 -1679 94 -1677
rect 100 -1673 101 -1671
rect 100 -1679 101 -1677
rect 107 -1673 108 -1671
rect 107 -1679 108 -1677
rect 114 -1673 115 -1671
rect 117 -1679 118 -1677
rect 121 -1673 122 -1671
rect 121 -1679 122 -1677
rect 128 -1673 129 -1671
rect 128 -1679 129 -1677
rect 135 -1673 136 -1671
rect 135 -1679 136 -1677
rect 142 -1673 143 -1671
rect 142 -1679 143 -1677
rect 149 -1673 150 -1671
rect 152 -1673 153 -1671
rect 156 -1673 157 -1671
rect 156 -1679 157 -1677
rect 163 -1673 164 -1671
rect 163 -1679 164 -1677
rect 170 -1673 171 -1671
rect 170 -1679 171 -1677
rect 177 -1679 178 -1677
rect 180 -1679 181 -1677
rect 184 -1673 185 -1671
rect 184 -1679 185 -1677
rect 191 -1673 192 -1671
rect 191 -1679 192 -1677
rect 198 -1679 199 -1677
rect 201 -1679 202 -1677
rect 205 -1673 206 -1671
rect 208 -1673 209 -1671
rect 212 -1673 213 -1671
rect 212 -1679 213 -1677
rect 219 -1673 220 -1671
rect 219 -1679 220 -1677
rect 226 -1673 227 -1671
rect 226 -1679 227 -1677
rect 233 -1673 234 -1671
rect 233 -1679 234 -1677
rect 240 -1673 241 -1671
rect 240 -1679 241 -1677
rect 247 -1673 248 -1671
rect 247 -1679 248 -1677
rect 257 -1673 258 -1671
rect 261 -1673 262 -1671
rect 261 -1679 262 -1677
rect 268 -1673 269 -1671
rect 268 -1679 269 -1677
rect 275 -1673 276 -1671
rect 275 -1679 276 -1677
rect 282 -1673 283 -1671
rect 282 -1679 283 -1677
rect 289 -1673 290 -1671
rect 289 -1679 290 -1677
rect 296 -1673 297 -1671
rect 303 -1673 304 -1671
rect 306 -1673 307 -1671
rect 306 -1679 307 -1677
rect 310 -1673 311 -1671
rect 310 -1679 311 -1677
rect 317 -1673 318 -1671
rect 317 -1679 318 -1677
rect 324 -1673 325 -1671
rect 324 -1679 325 -1677
rect 331 -1673 332 -1671
rect 334 -1673 335 -1671
rect 331 -1679 332 -1677
rect 334 -1679 335 -1677
rect 341 -1679 342 -1677
rect 345 -1673 346 -1671
rect 345 -1679 346 -1677
rect 352 -1673 353 -1671
rect 352 -1679 353 -1677
rect 359 -1673 360 -1671
rect 359 -1679 360 -1677
rect 366 -1673 367 -1671
rect 366 -1679 367 -1677
rect 373 -1673 374 -1671
rect 373 -1679 374 -1677
rect 380 -1673 381 -1671
rect 380 -1679 381 -1677
rect 387 -1673 388 -1671
rect 387 -1679 388 -1677
rect 394 -1673 395 -1671
rect 394 -1679 395 -1677
rect 401 -1673 402 -1671
rect 404 -1673 405 -1671
rect 401 -1679 402 -1677
rect 411 -1673 412 -1671
rect 408 -1679 409 -1677
rect 415 -1673 416 -1671
rect 415 -1679 416 -1677
rect 422 -1673 423 -1671
rect 422 -1679 423 -1677
rect 425 -1679 426 -1677
rect 429 -1673 430 -1671
rect 432 -1673 433 -1671
rect 432 -1679 433 -1677
rect 436 -1673 437 -1671
rect 436 -1679 437 -1677
rect 443 -1673 444 -1671
rect 443 -1679 444 -1677
rect 450 -1673 451 -1671
rect 450 -1679 451 -1677
rect 457 -1673 458 -1671
rect 457 -1679 458 -1677
rect 464 -1673 465 -1671
rect 464 -1679 465 -1677
rect 471 -1673 472 -1671
rect 471 -1679 472 -1677
rect 478 -1673 479 -1671
rect 478 -1679 479 -1677
rect 485 -1673 486 -1671
rect 485 -1679 486 -1677
rect 492 -1673 493 -1671
rect 492 -1679 493 -1677
rect 499 -1673 500 -1671
rect 499 -1679 500 -1677
rect 506 -1673 507 -1671
rect 506 -1679 507 -1677
rect 513 -1673 514 -1671
rect 516 -1673 517 -1671
rect 520 -1673 521 -1671
rect 523 -1673 524 -1671
rect 520 -1679 521 -1677
rect 523 -1679 524 -1677
rect 527 -1673 528 -1671
rect 527 -1679 528 -1677
rect 534 -1673 535 -1671
rect 534 -1679 535 -1677
rect 541 -1673 542 -1671
rect 544 -1673 545 -1671
rect 551 -1673 552 -1671
rect 548 -1679 549 -1677
rect 555 -1673 556 -1671
rect 555 -1679 556 -1677
rect 562 -1673 563 -1671
rect 562 -1679 563 -1677
rect 569 -1673 570 -1671
rect 569 -1679 570 -1677
rect 576 -1673 577 -1671
rect 576 -1679 577 -1677
rect 583 -1673 584 -1671
rect 583 -1679 584 -1677
rect 590 -1673 591 -1671
rect 590 -1679 591 -1677
rect 597 -1673 598 -1671
rect 597 -1679 598 -1677
rect 604 -1673 605 -1671
rect 604 -1679 605 -1677
rect 611 -1673 612 -1671
rect 611 -1679 612 -1677
rect 625 -1673 626 -1671
rect 625 -1679 626 -1677
rect 632 -1673 633 -1671
rect 632 -1679 633 -1677
rect 646 -1673 647 -1671
rect 646 -1679 647 -1677
rect 667 -1673 668 -1671
rect 667 -1679 668 -1677
rect 677 -1679 678 -1677
rect 681 -1673 682 -1671
rect 681 -1679 682 -1677
rect 688 -1673 689 -1671
rect 688 -1679 689 -1677
rect 691 -1679 692 -1677
rect 695 -1673 696 -1671
rect 695 -1679 696 -1677
rect 702 -1673 703 -1671
rect 702 -1679 703 -1677
rect 709 -1673 710 -1671
rect 709 -1679 710 -1677
rect 716 -1673 717 -1671
rect 716 -1679 717 -1677
rect 723 -1673 724 -1671
rect 723 -1679 724 -1677
rect 733 -1673 734 -1671
rect 737 -1673 738 -1671
rect 737 -1679 738 -1677
rect 744 -1673 745 -1671
rect 744 -1679 745 -1677
rect 751 -1673 752 -1671
rect 751 -1679 752 -1677
rect 758 -1673 759 -1671
rect 758 -1679 759 -1677
rect 765 -1673 766 -1671
rect 765 -1679 766 -1677
rect 775 -1673 776 -1671
rect 779 -1673 780 -1671
rect 782 -1679 783 -1677
rect 786 -1673 787 -1671
rect 786 -1679 787 -1677
rect 793 -1673 794 -1671
rect 793 -1679 794 -1677
rect 800 -1673 801 -1671
rect 803 -1673 804 -1671
rect 807 -1673 808 -1671
rect 807 -1679 808 -1677
rect 814 -1673 815 -1671
rect 814 -1679 815 -1677
rect 821 -1673 822 -1671
rect 821 -1679 822 -1677
rect 828 -1673 829 -1671
rect 828 -1679 829 -1677
rect 835 -1673 836 -1671
rect 838 -1673 839 -1671
rect 842 -1673 843 -1671
rect 842 -1679 843 -1677
rect 849 -1679 850 -1677
rect 852 -1679 853 -1677
rect 863 -1673 864 -1671
rect 863 -1679 864 -1677
rect 884 -1673 885 -1671
rect 884 -1679 885 -1677
rect 891 -1673 892 -1671
rect 891 -1679 892 -1677
rect 905 -1673 906 -1671
rect 905 -1679 906 -1677
rect 968 -1673 969 -1671
rect 968 -1679 969 -1677
rect 1024 -1673 1025 -1671
rect 1024 -1679 1025 -1677
rect 44 -1710 45 -1708
rect 44 -1716 45 -1714
rect 58 -1710 59 -1708
rect 58 -1716 59 -1714
rect 93 -1710 94 -1708
rect 93 -1716 94 -1714
rect 103 -1710 104 -1708
rect 100 -1716 101 -1714
rect 103 -1716 104 -1714
rect 114 -1710 115 -1708
rect 117 -1716 118 -1714
rect 128 -1710 129 -1708
rect 128 -1716 129 -1714
rect 142 -1710 143 -1708
rect 142 -1716 143 -1714
rect 149 -1710 150 -1708
rect 149 -1716 150 -1714
rect 156 -1710 157 -1708
rect 156 -1716 157 -1714
rect 163 -1710 164 -1708
rect 163 -1716 164 -1714
rect 170 -1710 171 -1708
rect 170 -1716 171 -1714
rect 177 -1710 178 -1708
rect 180 -1710 181 -1708
rect 184 -1716 185 -1714
rect 191 -1710 192 -1708
rect 191 -1716 192 -1714
rect 201 -1710 202 -1708
rect 208 -1710 209 -1708
rect 215 -1710 216 -1708
rect 212 -1716 213 -1714
rect 215 -1716 216 -1714
rect 219 -1710 220 -1708
rect 219 -1716 220 -1714
rect 226 -1710 227 -1708
rect 226 -1716 227 -1714
rect 233 -1710 234 -1708
rect 233 -1716 234 -1714
rect 240 -1710 241 -1708
rect 240 -1716 241 -1714
rect 254 -1710 255 -1708
rect 254 -1716 255 -1714
rect 264 -1710 265 -1708
rect 261 -1716 262 -1714
rect 268 -1710 269 -1708
rect 268 -1716 269 -1714
rect 275 -1710 276 -1708
rect 278 -1716 279 -1714
rect 282 -1710 283 -1708
rect 282 -1716 283 -1714
rect 289 -1710 290 -1708
rect 289 -1716 290 -1714
rect 296 -1716 297 -1714
rect 299 -1716 300 -1714
rect 303 -1710 304 -1708
rect 303 -1716 304 -1714
rect 310 -1710 311 -1708
rect 310 -1716 311 -1714
rect 317 -1710 318 -1708
rect 317 -1716 318 -1714
rect 324 -1710 325 -1708
rect 324 -1716 325 -1714
rect 331 -1710 332 -1708
rect 331 -1716 332 -1714
rect 341 -1710 342 -1708
rect 338 -1716 339 -1714
rect 345 -1710 346 -1708
rect 345 -1716 346 -1714
rect 355 -1710 356 -1708
rect 352 -1716 353 -1714
rect 359 -1710 360 -1708
rect 359 -1716 360 -1714
rect 366 -1710 367 -1708
rect 366 -1716 367 -1714
rect 373 -1710 374 -1708
rect 376 -1710 377 -1708
rect 373 -1716 374 -1714
rect 383 -1710 384 -1708
rect 383 -1716 384 -1714
rect 387 -1710 388 -1708
rect 394 -1710 395 -1708
rect 394 -1716 395 -1714
rect 404 -1710 405 -1708
rect 401 -1716 402 -1714
rect 408 -1710 409 -1708
rect 408 -1716 409 -1714
rect 415 -1710 416 -1708
rect 415 -1716 416 -1714
rect 422 -1710 423 -1708
rect 425 -1710 426 -1708
rect 422 -1716 423 -1714
rect 429 -1710 430 -1708
rect 429 -1716 430 -1714
rect 436 -1710 437 -1708
rect 436 -1716 437 -1714
rect 443 -1710 444 -1708
rect 443 -1716 444 -1714
rect 450 -1710 451 -1708
rect 450 -1716 451 -1714
rect 457 -1710 458 -1708
rect 457 -1716 458 -1714
rect 464 -1710 465 -1708
rect 464 -1716 465 -1714
rect 474 -1710 475 -1708
rect 471 -1716 472 -1714
rect 478 -1710 479 -1708
rect 478 -1716 479 -1714
rect 485 -1710 486 -1708
rect 485 -1716 486 -1714
rect 492 -1710 493 -1708
rect 492 -1716 493 -1714
rect 499 -1716 500 -1714
rect 506 -1710 507 -1708
rect 506 -1716 507 -1714
rect 513 -1710 514 -1708
rect 513 -1716 514 -1714
rect 520 -1710 521 -1708
rect 520 -1716 521 -1714
rect 527 -1710 528 -1708
rect 527 -1716 528 -1714
rect 534 -1710 535 -1708
rect 534 -1716 535 -1714
rect 541 -1710 542 -1708
rect 541 -1716 542 -1714
rect 548 -1710 549 -1708
rect 548 -1716 549 -1714
rect 555 -1710 556 -1708
rect 555 -1716 556 -1714
rect 562 -1710 563 -1708
rect 562 -1716 563 -1714
rect 569 -1710 570 -1708
rect 569 -1716 570 -1714
rect 576 -1710 577 -1708
rect 576 -1716 577 -1714
rect 583 -1710 584 -1708
rect 583 -1716 584 -1714
rect 590 -1710 591 -1708
rect 593 -1710 594 -1708
rect 593 -1716 594 -1714
rect 597 -1716 598 -1714
rect 604 -1710 605 -1708
rect 604 -1716 605 -1714
rect 611 -1710 612 -1708
rect 611 -1716 612 -1714
rect 618 -1710 619 -1708
rect 618 -1716 619 -1714
rect 639 -1710 640 -1708
rect 639 -1716 640 -1714
rect 646 -1710 647 -1708
rect 646 -1716 647 -1714
rect 653 -1710 654 -1708
rect 653 -1716 654 -1714
rect 674 -1710 675 -1708
rect 674 -1716 675 -1714
rect 681 -1716 682 -1714
rect 709 -1710 710 -1708
rect 709 -1716 710 -1714
rect 723 -1710 724 -1708
rect 723 -1716 724 -1714
rect 730 -1710 731 -1708
rect 730 -1716 731 -1714
rect 737 -1710 738 -1708
rect 737 -1716 738 -1714
rect 744 -1710 745 -1708
rect 744 -1716 745 -1714
rect 751 -1710 752 -1708
rect 751 -1716 752 -1714
rect 758 -1710 759 -1708
rect 758 -1716 759 -1714
rect 765 -1710 766 -1708
rect 765 -1716 766 -1714
rect 772 -1710 773 -1708
rect 772 -1716 773 -1714
rect 779 -1710 780 -1708
rect 779 -1716 780 -1714
rect 793 -1710 794 -1708
rect 793 -1716 794 -1714
rect 796 -1716 797 -1714
rect 800 -1710 801 -1708
rect 800 -1716 801 -1714
rect 807 -1710 808 -1708
rect 807 -1716 808 -1714
rect 817 -1710 818 -1708
rect 821 -1710 822 -1708
rect 821 -1716 822 -1714
rect 828 -1710 829 -1708
rect 828 -1716 829 -1714
rect 835 -1710 836 -1708
rect 835 -1716 836 -1714
rect 845 -1716 846 -1714
rect 849 -1710 850 -1708
rect 849 -1716 850 -1714
rect 856 -1710 857 -1708
rect 856 -1716 857 -1714
rect 863 -1710 864 -1708
rect 866 -1710 867 -1708
rect 866 -1716 867 -1714
rect 884 -1710 885 -1708
rect 884 -1716 885 -1714
rect 898 -1710 899 -1708
rect 898 -1716 899 -1714
rect 968 -1710 969 -1708
rect 968 -1716 969 -1714
rect 1024 -1710 1025 -1708
rect 1024 -1716 1025 -1714
rect 44 -1743 45 -1741
rect 44 -1749 45 -1747
rect 61 -1749 62 -1747
rect 65 -1743 66 -1741
rect 65 -1749 66 -1747
rect 100 -1743 101 -1741
rect 100 -1749 101 -1747
rect 107 -1743 108 -1741
rect 107 -1749 108 -1747
rect 114 -1743 115 -1741
rect 121 -1743 122 -1741
rect 121 -1749 122 -1747
rect 128 -1749 129 -1747
rect 131 -1749 132 -1747
rect 135 -1749 136 -1747
rect 138 -1749 139 -1747
rect 142 -1743 143 -1741
rect 145 -1743 146 -1741
rect 142 -1749 143 -1747
rect 145 -1749 146 -1747
rect 152 -1743 153 -1741
rect 156 -1743 157 -1741
rect 156 -1749 157 -1747
rect 159 -1749 160 -1747
rect 163 -1743 164 -1741
rect 163 -1749 164 -1747
rect 170 -1749 171 -1747
rect 173 -1749 174 -1747
rect 177 -1743 178 -1741
rect 177 -1749 178 -1747
rect 184 -1743 185 -1741
rect 184 -1749 185 -1747
rect 191 -1743 192 -1741
rect 191 -1749 192 -1747
rect 205 -1743 206 -1741
rect 205 -1749 206 -1747
rect 212 -1743 213 -1741
rect 219 -1749 220 -1747
rect 226 -1743 227 -1741
rect 233 -1743 234 -1741
rect 233 -1749 234 -1747
rect 240 -1743 241 -1741
rect 240 -1749 241 -1747
rect 247 -1743 248 -1741
rect 247 -1749 248 -1747
rect 275 -1743 276 -1741
rect 275 -1749 276 -1747
rect 296 -1743 297 -1741
rect 296 -1749 297 -1747
rect 303 -1743 304 -1741
rect 303 -1749 304 -1747
rect 310 -1743 311 -1741
rect 310 -1749 311 -1747
rect 317 -1743 318 -1741
rect 317 -1749 318 -1747
rect 324 -1743 325 -1741
rect 324 -1749 325 -1747
rect 331 -1743 332 -1741
rect 331 -1749 332 -1747
rect 338 -1743 339 -1741
rect 338 -1749 339 -1747
rect 345 -1743 346 -1741
rect 345 -1749 346 -1747
rect 352 -1743 353 -1741
rect 352 -1749 353 -1747
rect 359 -1743 360 -1741
rect 359 -1749 360 -1747
rect 366 -1743 367 -1741
rect 369 -1743 370 -1741
rect 366 -1749 367 -1747
rect 373 -1743 374 -1741
rect 373 -1749 374 -1747
rect 380 -1743 381 -1741
rect 380 -1749 381 -1747
rect 387 -1749 388 -1747
rect 394 -1743 395 -1741
rect 394 -1749 395 -1747
rect 404 -1749 405 -1747
rect 411 -1743 412 -1741
rect 411 -1749 412 -1747
rect 415 -1743 416 -1741
rect 415 -1749 416 -1747
rect 422 -1743 423 -1741
rect 422 -1749 423 -1747
rect 429 -1743 430 -1741
rect 429 -1749 430 -1747
rect 436 -1743 437 -1741
rect 436 -1749 437 -1747
rect 446 -1743 447 -1741
rect 450 -1743 451 -1741
rect 450 -1749 451 -1747
rect 457 -1743 458 -1741
rect 457 -1749 458 -1747
rect 464 -1743 465 -1741
rect 464 -1749 465 -1747
rect 471 -1749 472 -1747
rect 478 -1743 479 -1741
rect 478 -1749 479 -1747
rect 485 -1743 486 -1741
rect 488 -1749 489 -1747
rect 492 -1743 493 -1741
rect 492 -1749 493 -1747
rect 499 -1743 500 -1741
rect 499 -1749 500 -1747
rect 506 -1749 507 -1747
rect 509 -1749 510 -1747
rect 513 -1743 514 -1741
rect 513 -1749 514 -1747
rect 520 -1743 521 -1741
rect 520 -1749 521 -1747
rect 530 -1749 531 -1747
rect 534 -1743 535 -1741
rect 534 -1749 535 -1747
rect 541 -1743 542 -1741
rect 541 -1749 542 -1747
rect 548 -1743 549 -1741
rect 548 -1749 549 -1747
rect 555 -1743 556 -1741
rect 555 -1749 556 -1747
rect 562 -1749 563 -1747
rect 569 -1743 570 -1741
rect 569 -1749 570 -1747
rect 576 -1743 577 -1741
rect 576 -1749 577 -1747
rect 586 -1749 587 -1747
rect 590 -1743 591 -1741
rect 590 -1749 591 -1747
rect 597 -1743 598 -1741
rect 597 -1749 598 -1747
rect 646 -1743 647 -1741
rect 646 -1749 647 -1747
rect 656 -1743 657 -1741
rect 656 -1749 657 -1747
rect 702 -1743 703 -1741
rect 702 -1749 703 -1747
rect 709 -1743 710 -1741
rect 709 -1749 710 -1747
rect 716 -1749 717 -1747
rect 723 -1743 724 -1741
rect 723 -1749 724 -1747
rect 730 -1743 731 -1741
rect 730 -1749 731 -1747
rect 737 -1743 738 -1741
rect 737 -1749 738 -1747
rect 744 -1743 745 -1741
rect 744 -1749 745 -1747
rect 751 -1743 752 -1741
rect 751 -1749 752 -1747
rect 758 -1743 759 -1741
rect 758 -1749 759 -1747
rect 765 -1743 766 -1741
rect 765 -1749 766 -1747
rect 772 -1749 773 -1747
rect 782 -1743 783 -1741
rect 779 -1749 780 -1747
rect 782 -1749 783 -1747
rect 786 -1743 787 -1741
rect 786 -1749 787 -1747
rect 793 -1743 794 -1741
rect 796 -1743 797 -1741
rect 793 -1749 794 -1747
rect 800 -1743 801 -1741
rect 800 -1749 801 -1747
rect 807 -1743 808 -1741
rect 807 -1749 808 -1747
rect 828 -1743 829 -1741
rect 828 -1749 829 -1747
rect 842 -1743 843 -1741
rect 842 -1749 843 -1747
rect 856 -1743 857 -1741
rect 856 -1749 857 -1747
rect 884 -1743 885 -1741
rect 884 -1749 885 -1747
rect 898 -1743 899 -1741
rect 898 -1749 899 -1747
rect 968 -1743 969 -1741
rect 968 -1749 969 -1747
rect 975 -1749 976 -1747
rect 1024 -1743 1025 -1741
rect 1024 -1749 1025 -1747
rect 47 -1770 48 -1768
rect 58 -1770 59 -1768
rect 58 -1776 59 -1774
rect 65 -1770 66 -1768
rect 65 -1776 66 -1774
rect 72 -1770 73 -1768
rect 72 -1776 73 -1774
rect 79 -1770 80 -1768
rect 79 -1776 80 -1774
rect 93 -1770 94 -1768
rect 93 -1776 94 -1774
rect 100 -1770 101 -1768
rect 110 -1776 111 -1774
rect 117 -1770 118 -1768
rect 117 -1776 118 -1774
rect 121 -1770 122 -1768
rect 128 -1770 129 -1768
rect 128 -1776 129 -1774
rect 135 -1770 136 -1768
rect 135 -1776 136 -1774
rect 142 -1770 143 -1768
rect 142 -1776 143 -1774
rect 152 -1776 153 -1774
rect 156 -1770 157 -1768
rect 170 -1770 171 -1768
rect 170 -1776 171 -1774
rect 191 -1770 192 -1768
rect 191 -1776 192 -1774
rect 198 -1776 199 -1774
rect 205 -1770 206 -1768
rect 205 -1776 206 -1774
rect 212 -1770 213 -1768
rect 219 -1770 220 -1768
rect 219 -1776 220 -1774
rect 229 -1770 230 -1768
rect 226 -1776 227 -1774
rect 233 -1770 234 -1768
rect 233 -1776 234 -1774
rect 240 -1770 241 -1768
rect 240 -1776 241 -1774
rect 275 -1770 276 -1768
rect 275 -1776 276 -1774
rect 282 -1770 283 -1768
rect 282 -1776 283 -1774
rect 289 -1770 290 -1768
rect 289 -1776 290 -1774
rect 296 -1770 297 -1768
rect 296 -1776 297 -1774
rect 306 -1776 307 -1774
rect 310 -1770 311 -1768
rect 310 -1776 311 -1774
rect 317 -1770 318 -1768
rect 324 -1770 325 -1768
rect 324 -1776 325 -1774
rect 331 -1776 332 -1774
rect 338 -1770 339 -1768
rect 338 -1776 339 -1774
rect 345 -1770 346 -1768
rect 345 -1776 346 -1774
rect 352 -1770 353 -1768
rect 352 -1776 353 -1774
rect 359 -1770 360 -1768
rect 362 -1776 363 -1774
rect 369 -1770 370 -1768
rect 373 -1770 374 -1768
rect 373 -1776 374 -1774
rect 380 -1770 381 -1768
rect 380 -1776 381 -1774
rect 394 -1770 395 -1768
rect 394 -1776 395 -1774
rect 401 -1770 402 -1768
rect 401 -1776 402 -1774
rect 411 -1776 412 -1774
rect 415 -1770 416 -1768
rect 415 -1776 416 -1774
rect 422 -1770 423 -1768
rect 429 -1770 430 -1768
rect 443 -1770 444 -1768
rect 443 -1776 444 -1774
rect 450 -1770 451 -1768
rect 450 -1776 451 -1774
rect 457 -1770 458 -1768
rect 457 -1776 458 -1774
rect 464 -1770 465 -1768
rect 464 -1776 465 -1774
rect 471 -1770 472 -1768
rect 471 -1776 472 -1774
rect 478 -1770 479 -1768
rect 478 -1776 479 -1774
rect 506 -1770 507 -1768
rect 506 -1776 507 -1774
rect 513 -1770 514 -1768
rect 513 -1776 514 -1774
rect 527 -1770 528 -1768
rect 527 -1776 528 -1774
rect 562 -1770 563 -1768
rect 562 -1776 563 -1774
rect 709 -1770 710 -1768
rect 709 -1776 710 -1774
rect 716 -1776 717 -1774
rect 723 -1770 724 -1768
rect 723 -1776 724 -1774
rect 730 -1770 731 -1768
rect 730 -1776 731 -1774
rect 737 -1770 738 -1768
rect 737 -1776 738 -1774
rect 747 -1776 748 -1774
rect 751 -1770 752 -1768
rect 751 -1776 752 -1774
rect 758 -1770 759 -1768
rect 758 -1776 759 -1774
rect 772 -1770 773 -1768
rect 772 -1776 773 -1774
rect 779 -1776 780 -1774
rect 793 -1770 794 -1768
rect 793 -1776 794 -1774
rect 814 -1770 815 -1768
rect 814 -1776 815 -1774
rect 828 -1770 829 -1768
rect 828 -1776 829 -1774
rect 845 -1770 846 -1768
rect 856 -1770 857 -1768
rect 880 -1776 881 -1774
rect 884 -1770 885 -1768
rect 884 -1776 885 -1774
rect 898 -1770 899 -1768
rect 898 -1776 899 -1774
rect 1024 -1770 1025 -1768
rect 1024 -1776 1025 -1774
rect 68 -1797 69 -1795
rect 75 -1791 76 -1789
rect 79 -1791 80 -1789
rect 79 -1797 80 -1795
rect 142 -1791 143 -1789
rect 142 -1797 143 -1795
rect 152 -1791 153 -1789
rect 149 -1797 150 -1795
rect 156 -1791 157 -1789
rect 156 -1797 157 -1795
rect 173 -1791 174 -1789
rect 184 -1797 185 -1795
rect 205 -1791 206 -1789
rect 205 -1797 206 -1795
rect 226 -1791 227 -1789
rect 226 -1797 227 -1795
rect 240 -1791 241 -1789
rect 240 -1797 241 -1795
rect 247 -1791 248 -1789
rect 247 -1797 248 -1795
rect 261 -1791 262 -1789
rect 261 -1797 262 -1795
rect 282 -1791 283 -1789
rect 282 -1797 283 -1795
rect 296 -1791 297 -1789
rect 296 -1797 297 -1795
rect 303 -1791 304 -1789
rect 306 -1791 307 -1789
rect 313 -1791 314 -1789
rect 320 -1791 321 -1789
rect 324 -1791 325 -1789
rect 324 -1797 325 -1795
rect 331 -1791 332 -1789
rect 331 -1797 332 -1795
rect 338 -1791 339 -1789
rect 338 -1797 339 -1795
rect 345 -1797 346 -1795
rect 352 -1791 353 -1789
rect 352 -1797 353 -1795
rect 380 -1791 381 -1789
rect 380 -1797 381 -1795
rect 387 -1791 388 -1789
rect 387 -1797 388 -1795
rect 411 -1791 412 -1789
rect 415 -1791 416 -1789
rect 415 -1797 416 -1795
rect 422 -1791 423 -1789
rect 422 -1797 423 -1795
rect 429 -1797 430 -1795
rect 432 -1797 433 -1795
rect 439 -1797 440 -1795
rect 443 -1791 444 -1789
rect 443 -1797 444 -1795
rect 450 -1791 451 -1789
rect 450 -1797 451 -1795
rect 457 -1791 458 -1789
rect 457 -1797 458 -1795
rect 471 -1791 472 -1789
rect 471 -1797 472 -1795
rect 478 -1791 479 -1789
rect 478 -1797 479 -1795
rect 502 -1791 503 -1789
rect 506 -1797 507 -1795
rect 513 -1791 514 -1789
rect 513 -1797 514 -1795
rect 520 -1791 521 -1789
rect 520 -1797 521 -1795
rect 565 -1791 566 -1789
rect 737 -1791 738 -1789
rect 737 -1797 738 -1795
rect 744 -1797 745 -1795
rect 754 -1797 755 -1795
rect 758 -1791 759 -1789
rect 758 -1797 759 -1795
rect 765 -1791 766 -1789
rect 765 -1797 766 -1795
rect 772 -1791 773 -1789
rect 793 -1791 794 -1789
rect 793 -1797 794 -1795
rect 814 -1791 815 -1789
rect 838 -1791 839 -1789
rect 898 -1791 899 -1789
rect 898 -1797 899 -1795
rect 1024 -1791 1025 -1789
rect 1024 -1797 1025 -1795
rect 159 -1806 160 -1804
rect 187 -1812 188 -1810
rect 191 -1806 192 -1804
rect 191 -1812 192 -1810
rect 208 -1806 209 -1804
rect 222 -1812 223 -1810
rect 226 -1806 227 -1804
rect 226 -1812 227 -1810
rect 264 -1812 265 -1810
rect 268 -1806 269 -1804
rect 268 -1812 269 -1810
rect 282 -1806 283 -1804
rect 296 -1806 297 -1804
rect 296 -1812 297 -1810
rect 306 -1812 307 -1810
rect 324 -1812 325 -1810
rect 331 -1806 332 -1804
rect 331 -1812 332 -1810
rect 341 -1806 342 -1804
rect 352 -1806 353 -1804
rect 352 -1812 353 -1810
rect 359 -1812 360 -1810
rect 376 -1812 377 -1810
rect 383 -1806 384 -1804
rect 387 -1806 388 -1804
rect 387 -1812 388 -1810
rect 422 -1806 423 -1804
rect 422 -1812 423 -1810
rect 429 -1812 430 -1810
rect 464 -1806 465 -1804
rect 471 -1806 472 -1804
rect 481 -1806 482 -1804
rect 516 -1806 517 -1804
rect 747 -1812 748 -1810
rect 751 -1806 752 -1804
rect 751 -1812 752 -1810
rect 796 -1806 797 -1804
rect 901 -1812 902 -1810
rect 905 -1806 906 -1804
rect 905 -1812 906 -1810
rect 1027 -1806 1028 -1804
<< metal1 >>
rect 177 0 199 1
rect 212 0 220 1
rect 236 0 241 1
rect 254 0 262 1
rect 285 0 290 1
rect 303 0 311 1
rect 338 0 349 1
rect 352 0 360 1
rect 366 0 409 1
rect 467 0 472 1
rect 478 0 486 1
rect 534 0 542 1
rect 576 0 584 1
rect 604 0 612 1
rect 730 0 741 1
rect 184 -2 195 -1
rect 114 -13 122 -12
rect 156 -13 164 -12
rect 170 -13 178 -12
rect 219 -13 227 -12
rect 240 -13 255 -12
rect 278 -13 283 -12
rect 303 -13 311 -12
rect 345 -13 367 -12
rect 408 -13 444 -12
rect 450 -13 461 -12
rect 474 -13 479 -12
rect 485 -13 493 -12
rect 527 -13 559 -12
rect 604 -13 612 -12
rect 618 -13 622 -12
rect 688 -13 699 -12
rect 215 -15 220 -14
rect 247 -15 262 -14
rect 289 -15 304 -14
rect 352 -15 360 -14
rect 366 -15 374 -14
rect 415 -15 423 -14
rect 425 -15 430 -14
rect 457 -15 468 -14
rect 471 -15 486 -14
rect 555 -15 605 -14
rect 240 -17 262 -16
rect 278 -17 290 -16
rect 338 -17 353 -16
rect 334 -19 339 -18
rect 58 -30 62 -29
rect 114 -30 125 -29
rect 142 -30 171 -29
rect 184 -30 199 -29
rect 212 -30 220 -29
rect 226 -30 262 -29
rect 268 -30 297 -29
rect 317 -30 325 -29
rect 334 -30 346 -29
rect 352 -30 374 -29
rect 387 -30 402 -29
rect 408 -30 412 -29
rect 415 -30 426 -29
rect 429 -30 433 -29
rect 443 -30 472 -29
rect 492 -30 500 -29
rect 513 -30 538 -29
rect 541 -30 549 -29
rect 576 -30 580 -29
rect 583 -30 598 -29
rect 604 -30 633 -29
rect 646 -30 661 -29
rect 709 -30 787 -29
rect 807 -30 815 -29
rect 121 -32 136 -31
rect 152 -32 157 -31
rect 163 -32 174 -31
rect 177 -32 227 -31
rect 233 -32 241 -31
rect 254 -32 297 -31
rect 345 -32 367 -31
rect 429 -32 437 -31
rect 527 -32 556 -31
rect 572 -32 584 -31
rect 604 -32 612 -31
rect 625 -32 713 -31
rect 163 -34 171 -33
rect 180 -34 185 -33
rect 240 -34 283 -33
rect 352 -34 398 -33
rect 432 -34 437 -33
rect 541 -34 563 -33
rect 611 -34 619 -33
rect 247 -36 255 -35
rect 257 -36 276 -35
rect 282 -36 311 -35
rect 359 -36 367 -35
rect 247 -38 272 -37
rect 303 -38 311 -37
rect 338 -38 360 -37
rect 303 -40 332 -39
rect 317 -42 339 -41
rect 93 -53 104 -52
rect 107 -53 150 -52
rect 170 -53 185 -52
rect 226 -53 279 -52
rect 310 -53 332 -52
rect 338 -53 402 -52
rect 415 -53 461 -52
rect 478 -53 507 -52
rect 513 -53 521 -52
rect 534 -53 619 -52
rect 660 -53 675 -52
rect 688 -53 703 -52
rect 793 -53 808 -52
rect 1087 -53 1098 -52
rect 110 -55 206 -54
rect 229 -55 297 -54
rect 373 -55 388 -54
rect 429 -55 444 -54
rect 485 -55 514 -54
rect 541 -55 584 -54
rect 653 -55 661 -54
rect 786 -55 808 -54
rect 121 -57 136 -56
rect 170 -57 192 -56
rect 233 -57 255 -56
rect 289 -57 311 -56
rect 373 -57 468 -56
rect 474 -57 486 -56
rect 499 -57 535 -56
rect 555 -57 647 -56
rect 128 -59 178 -58
rect 184 -59 276 -58
rect 289 -59 300 -58
rect 380 -59 402 -58
rect 422 -59 444 -58
rect 471 -59 500 -58
rect 527 -59 556 -58
rect 569 -59 626 -58
rect 632 -59 654 -58
rect 135 -61 157 -60
rect 191 -61 209 -60
rect 233 -61 262 -60
rect 380 -61 409 -60
rect 422 -61 451 -60
rect 495 -61 626 -60
rect 632 -61 640 -60
rect 156 -63 199 -62
rect 208 -63 213 -62
rect 247 -63 262 -62
rect 408 -63 458 -62
rect 576 -63 584 -62
rect 198 -65 283 -64
rect 429 -65 447 -64
rect 576 -65 605 -64
rect 212 -67 304 -66
rect 436 -67 451 -66
rect 597 -67 605 -66
rect 222 -69 248 -68
rect 268 -69 304 -68
rect 439 -69 479 -68
rect 590 -69 598 -68
rect 268 -71 360 -70
rect 562 -71 591 -70
rect 282 -73 318 -72
rect 548 -73 563 -72
rect 317 -75 353 -74
rect 446 -75 549 -74
rect 324 -77 353 -76
rect 324 -79 395 -78
rect 131 -81 395 -80
rect 30 -92 45 -91
rect 51 -92 66 -91
rect 89 -92 94 -91
rect 100 -92 157 -91
rect 219 -92 269 -91
rect 275 -92 290 -91
rect 299 -92 353 -91
rect 366 -92 395 -91
rect 397 -92 412 -91
rect 429 -92 496 -91
rect 527 -92 556 -91
rect 597 -92 633 -91
rect 646 -92 689 -91
rect 730 -92 738 -91
rect 758 -92 780 -91
rect 800 -92 808 -91
rect 898 -92 906 -91
rect 975 -92 979 -91
rect 54 -94 66 -93
rect 93 -94 143 -93
rect 149 -94 188 -93
rect 261 -94 269 -93
rect 282 -94 290 -93
rect 303 -94 307 -93
rect 338 -94 367 -93
rect 387 -94 391 -93
rect 401 -94 430 -93
rect 450 -94 472 -93
rect 478 -94 493 -93
rect 541 -94 598 -93
rect 604 -94 668 -93
rect 674 -94 717 -93
rect 765 -94 794 -93
rect 107 -96 416 -95
rect 450 -96 640 -95
rect 681 -96 724 -95
rect 121 -98 185 -97
rect 240 -98 262 -97
rect 282 -98 318 -97
rect 327 -98 339 -97
rect 373 -98 416 -97
rect 457 -98 486 -97
rect 534 -98 640 -97
rect 702 -98 731 -97
rect 124 -100 178 -99
rect 240 -100 248 -99
rect 303 -100 311 -99
rect 317 -100 325 -99
rect 380 -100 402 -99
rect 408 -100 444 -99
rect 467 -100 486 -99
rect 499 -100 535 -99
rect 541 -100 570 -99
rect 590 -100 647 -99
rect 660 -100 703 -99
rect 128 -102 181 -101
rect 324 -102 437 -101
rect 520 -102 570 -101
rect 593 -102 682 -101
rect 128 -104 346 -103
rect 355 -104 521 -103
rect 562 -104 605 -103
rect 611 -104 661 -103
rect 135 -106 181 -105
rect 212 -106 346 -105
rect 362 -106 500 -105
rect 506 -106 563 -105
rect 618 -106 675 -105
rect 142 -108 199 -107
rect 212 -108 234 -107
rect 373 -108 437 -107
rect 548 -108 612 -107
rect 625 -108 696 -107
rect 149 -110 206 -109
rect 233 -110 255 -109
rect 387 -110 423 -109
rect 513 -110 626 -109
rect 156 -112 164 -111
rect 198 -112 230 -111
rect 390 -112 423 -111
rect 576 -112 619 -111
rect 163 -114 171 -113
rect 205 -114 360 -113
rect 408 -114 514 -113
rect 576 -114 654 -113
rect 170 -116 192 -115
rect 229 -116 255 -115
rect 299 -116 360 -115
rect 191 -118 223 -117
rect 23 -129 45 -128
rect 47 -129 66 -128
rect 79 -129 87 -128
rect 121 -129 185 -128
rect 219 -129 325 -128
rect 338 -129 409 -128
rect 457 -129 465 -128
rect 495 -129 507 -128
rect 541 -129 594 -128
rect 656 -129 759 -128
rect 779 -129 850 -128
rect 905 -129 920 -128
rect 30 -131 38 -130
rect 121 -131 206 -130
rect 219 -131 283 -130
rect 296 -131 304 -130
rect 324 -131 339 -130
rect 345 -131 353 -130
rect 380 -131 430 -130
rect 443 -131 458 -130
rect 509 -131 542 -130
rect 555 -131 696 -130
rect 737 -131 752 -130
rect 30 -133 52 -132
rect 149 -133 377 -132
rect 394 -133 430 -132
rect 471 -133 556 -132
rect 583 -133 654 -132
rect 667 -133 787 -132
rect 51 -135 59 -134
rect 149 -135 482 -134
rect 513 -135 584 -134
rect 590 -135 689 -134
rect 695 -135 766 -134
rect 156 -137 167 -136
rect 170 -137 381 -136
rect 394 -137 416 -136
rect 450 -137 472 -136
rect 520 -137 780 -136
rect 58 -139 157 -138
rect 170 -139 188 -138
rect 198 -139 377 -138
rect 401 -139 416 -138
rect 450 -139 549 -138
rect 604 -139 668 -138
rect 674 -139 794 -138
rect 142 -141 402 -140
rect 499 -141 549 -140
rect 562 -141 675 -140
rect 681 -141 808 -140
rect 135 -143 500 -142
rect 527 -143 563 -142
rect 604 -143 724 -142
rect 744 -143 801 -142
rect 142 -145 164 -144
rect 205 -145 213 -144
rect 226 -145 349 -144
rect 492 -145 528 -144
rect 569 -145 724 -144
rect 730 -145 801 -144
rect 212 -147 276 -146
rect 282 -147 391 -146
rect 569 -147 703 -146
rect 709 -147 738 -146
rect 229 -149 360 -148
rect 618 -149 682 -148
rect 702 -149 846 -148
rect 233 -151 353 -150
rect 359 -151 367 -150
rect 534 -151 619 -150
rect 625 -151 731 -150
rect 233 -153 248 -152
rect 250 -153 255 -152
rect 275 -153 468 -152
rect 597 -153 626 -152
rect 632 -153 689 -152
rect 240 -155 318 -154
rect 334 -155 514 -154
rect 597 -155 717 -154
rect 72 -157 318 -156
rect 345 -157 423 -156
rect 478 -157 633 -156
rect 639 -157 766 -156
rect 243 -159 321 -158
rect 366 -159 384 -158
rect 422 -159 773 -158
rect 247 -161 262 -160
rect 303 -161 332 -160
rect 436 -161 640 -160
rect 646 -161 710 -160
rect 254 -163 290 -162
rect 331 -163 444 -162
rect 478 -163 815 -162
rect 107 -165 290 -164
rect 387 -165 437 -164
rect 611 -165 647 -164
rect 660 -165 717 -164
rect 107 -167 129 -166
rect 261 -167 269 -166
rect 387 -167 486 -166
rect 537 -167 661 -166
rect 128 -169 139 -168
rect 268 -169 311 -168
rect 576 -169 612 -168
rect 100 -171 311 -170
rect 523 -171 577 -170
rect 93 -173 101 -172
rect 114 -173 139 -172
rect 93 -175 178 -174
rect 177 -177 192 -176
rect 191 -179 489 -178
rect 16 -190 304 -189
rect 317 -190 577 -189
rect 758 -190 871 -189
rect 919 -190 948 -189
rect 30 -192 66 -191
rect 68 -192 104 -191
rect 117 -192 199 -191
rect 201 -192 234 -191
rect 240 -192 332 -191
rect 338 -192 437 -191
rect 460 -192 731 -191
rect 765 -192 815 -191
rect 821 -192 920 -191
rect 23 -194 69 -193
rect 72 -194 202 -193
rect 205 -194 353 -193
rect 355 -194 437 -193
rect 485 -194 885 -193
rect 23 -196 101 -195
rect 163 -196 178 -195
rect 184 -196 213 -195
rect 233 -196 269 -195
rect 292 -196 388 -195
rect 422 -196 556 -195
rect 660 -196 731 -195
rect 744 -196 766 -195
rect 772 -196 878 -195
rect 30 -198 115 -197
rect 142 -198 213 -197
rect 261 -198 269 -197
rect 296 -198 318 -197
rect 345 -198 906 -197
rect 37 -200 248 -199
rect 303 -200 374 -199
rect 380 -200 556 -199
rect 674 -200 759 -199
rect 786 -200 857 -199
rect 859 -200 934 -199
rect 44 -202 283 -201
rect 352 -202 640 -201
rect 702 -202 745 -201
rect 751 -202 787 -201
rect 793 -202 864 -201
rect 72 -204 157 -203
rect 170 -204 178 -203
rect 187 -204 297 -203
rect 373 -204 395 -203
rect 408 -204 423 -203
rect 495 -204 521 -203
rect 527 -204 675 -203
rect 681 -204 752 -203
rect 800 -204 892 -203
rect 79 -206 241 -205
rect 247 -206 276 -205
rect 408 -206 538 -205
rect 541 -206 577 -205
rect 604 -206 640 -205
rect 681 -206 689 -205
rect 709 -206 773 -205
rect 800 -206 843 -205
rect 79 -208 349 -207
rect 450 -208 528 -207
rect 534 -208 591 -207
rect 625 -208 689 -207
rect 737 -208 794 -207
rect 807 -208 941 -207
rect 107 -210 395 -209
rect 429 -210 451 -209
rect 478 -210 542 -209
rect 548 -210 626 -209
rect 646 -210 710 -209
rect 716 -210 808 -209
rect 821 -210 850 -209
rect 58 -212 549 -211
rect 583 -212 605 -211
rect 667 -212 738 -211
rect 779 -212 850 -211
rect 51 -214 59 -213
rect 107 -214 136 -213
rect 142 -214 150 -213
rect 187 -214 584 -213
rect 695 -214 717 -213
rect 723 -214 780 -213
rect 828 -214 927 -213
rect 51 -216 66 -215
rect 114 -216 129 -215
rect 149 -216 220 -215
rect 254 -216 283 -215
rect 324 -216 430 -215
rect 464 -216 829 -215
rect 835 -216 899 -215
rect 121 -218 129 -217
rect 191 -218 255 -217
rect 275 -218 619 -217
rect 632 -218 696 -217
rect 93 -220 192 -219
rect 310 -220 325 -219
rect 345 -220 479 -219
rect 499 -220 661 -219
rect 93 -222 913 -221
rect 121 -224 230 -223
rect 467 -224 668 -223
rect 173 -226 311 -225
rect 366 -226 468 -225
rect 471 -226 500 -225
rect 513 -226 703 -225
rect 289 -228 367 -227
rect 457 -228 472 -227
rect 506 -228 514 -227
rect 593 -228 836 -227
rect 443 -230 507 -229
rect 597 -230 633 -229
rect 653 -230 724 -229
rect 415 -232 444 -231
rect 611 -232 619 -231
rect 401 -234 416 -233
rect 425 -234 654 -233
rect 100 -236 402 -235
rect 569 -236 612 -235
rect 226 -238 570 -237
rect 30 -249 160 -248
rect 170 -249 213 -248
rect 233 -249 293 -248
rect 352 -249 507 -248
rect 579 -249 773 -248
rect 877 -249 962 -248
rect 975 -249 983 -248
rect 1087 -249 1095 -248
rect 33 -251 486 -250
rect 488 -251 780 -250
rect 877 -251 934 -250
rect 947 -251 976 -250
rect 37 -253 199 -252
rect 208 -253 556 -252
rect 586 -253 829 -252
rect 37 -255 90 -254
rect 93 -255 248 -254
rect 254 -255 283 -254
rect 380 -255 395 -254
rect 436 -255 507 -254
rect 527 -255 556 -254
rect 593 -255 654 -254
rect 758 -255 773 -254
rect 779 -255 794 -254
rect 828 -255 885 -254
rect 44 -257 290 -256
rect 383 -257 591 -256
rect 600 -257 710 -256
rect 765 -257 801 -256
rect 884 -257 892 -256
rect 47 -259 87 -258
rect 93 -259 304 -258
rect 394 -259 514 -258
rect 520 -259 528 -258
rect 597 -259 766 -258
rect 891 -259 955 -258
rect 58 -261 192 -260
rect 205 -261 255 -260
rect 275 -261 482 -260
rect 495 -261 675 -260
rect 702 -261 955 -260
rect 23 -263 192 -262
rect 233 -263 458 -262
rect 464 -263 647 -262
rect 653 -263 731 -262
rect 23 -265 52 -264
rect 65 -265 440 -264
rect 478 -265 836 -264
rect 79 -267 213 -266
rect 338 -267 458 -266
rect 499 -267 514 -266
rect 562 -267 598 -266
rect 604 -267 675 -266
rect 695 -267 731 -266
rect 79 -269 794 -268
rect 82 -271 101 -270
rect 103 -271 129 -270
rect 135 -271 248 -270
rect 331 -271 339 -270
rect 373 -271 521 -270
rect 541 -271 563 -270
rect 583 -271 605 -270
rect 618 -271 647 -270
rect 695 -271 738 -270
rect 107 -273 570 -272
rect 576 -273 619 -272
rect 667 -273 738 -272
rect 117 -275 332 -274
rect 359 -275 374 -274
rect 411 -275 759 -274
rect 128 -277 325 -276
rect 359 -277 416 -276
rect 450 -277 479 -276
rect 583 -277 682 -276
rect 702 -277 724 -276
rect 135 -279 262 -278
rect 317 -279 325 -278
rect 415 -279 836 -278
rect 142 -281 276 -280
rect 422 -281 451 -280
rect 471 -281 500 -280
rect 639 -281 668 -280
rect 681 -281 689 -280
rect 709 -281 850 -280
rect 114 -283 689 -282
rect 723 -283 752 -282
rect 849 -283 927 -282
rect 114 -285 164 -284
rect 170 -285 297 -284
rect 422 -285 430 -284
rect 471 -285 815 -284
rect 912 -285 927 -284
rect 145 -287 304 -286
rect 429 -287 444 -286
rect 474 -287 570 -286
rect 625 -287 640 -286
rect 744 -287 752 -286
rect 912 -287 941 -286
rect 156 -289 549 -288
rect 625 -289 661 -288
rect 716 -289 745 -288
rect 821 -289 941 -288
rect 156 -291 206 -290
rect 219 -291 297 -290
rect 401 -291 444 -290
rect 492 -291 815 -290
rect 163 -293 549 -292
rect 632 -293 661 -292
rect 786 -293 822 -292
rect 177 -295 185 -294
rect 219 -295 241 -294
rect 264 -295 318 -294
rect 366 -295 402 -294
rect 492 -295 871 -294
rect 16 -297 178 -296
rect 226 -297 241 -296
rect 310 -297 367 -296
rect 611 -297 633 -296
rect 786 -297 808 -296
rect 870 -297 920 -296
rect 16 -299 465 -298
rect 807 -299 857 -298
rect 863 -299 920 -298
rect 72 -301 311 -300
rect 408 -301 612 -300
rect 842 -301 857 -300
rect 863 -301 899 -300
rect 72 -303 346 -302
rect 842 -303 969 -302
rect 149 -305 346 -304
rect 898 -305 937 -304
rect 149 -307 388 -306
rect 229 -309 262 -308
rect 9 -320 146 -319
rect 205 -320 209 -319
rect 226 -320 269 -319
rect 296 -320 409 -319
rect 436 -320 927 -319
rect 933 -320 983 -319
rect 999 -320 1067 -319
rect 1094 -320 1109 -319
rect 16 -322 475 -321
rect 523 -322 654 -321
rect 681 -322 685 -321
rect 716 -322 906 -321
rect 947 -322 969 -321
rect 16 -324 136 -323
rect 208 -324 293 -323
rect 317 -324 465 -323
rect 527 -324 545 -323
rect 548 -324 962 -323
rect 964 -324 1053 -323
rect 23 -326 118 -325
rect 121 -326 297 -325
rect 331 -326 468 -325
rect 541 -326 955 -325
rect 23 -328 304 -327
rect 345 -328 384 -327
rect 390 -328 521 -327
rect 534 -328 542 -327
rect 548 -328 920 -327
rect 37 -330 52 -329
rect 58 -330 419 -329
rect 443 -330 584 -329
rect 632 -330 654 -329
rect 681 -330 885 -329
rect 898 -330 983 -329
rect 40 -332 59 -331
rect 65 -332 164 -331
rect 212 -332 437 -331
rect 443 -332 489 -331
rect 499 -332 535 -331
rect 579 -332 906 -331
rect 44 -334 146 -333
rect 212 -334 486 -333
rect 618 -334 633 -333
rect 716 -334 815 -333
rect 821 -334 927 -333
rect 65 -336 108 -335
rect 121 -336 325 -335
rect 338 -336 346 -335
rect 352 -336 356 -335
rect 359 -336 416 -335
rect 422 -336 500 -335
rect 786 -336 885 -335
rect 901 -336 976 -335
rect 30 -338 423 -337
rect 453 -338 773 -337
rect 807 -338 822 -337
rect 828 -338 976 -337
rect 93 -340 290 -339
rect 352 -340 395 -339
rect 401 -340 409 -339
rect 457 -340 528 -339
rect 702 -340 773 -339
rect 835 -340 1011 -339
rect 93 -342 181 -341
rect 191 -342 619 -341
rect 639 -342 703 -341
rect 744 -342 787 -341
rect 842 -342 948 -341
rect 100 -344 108 -343
rect 135 -344 164 -343
rect 254 -344 269 -343
rect 275 -344 304 -343
rect 359 -344 479 -343
rect 506 -344 829 -343
rect 849 -344 1018 -343
rect 79 -346 479 -345
rect 590 -346 640 -345
rect 723 -346 850 -345
rect 863 -346 990 -345
rect 79 -348 171 -347
rect 219 -348 255 -347
rect 261 -348 332 -347
rect 380 -348 920 -347
rect 72 -350 381 -349
rect 394 -350 472 -349
rect 474 -350 724 -349
rect 751 -350 808 -349
rect 870 -350 1004 -349
rect 72 -352 87 -351
rect 100 -352 111 -351
rect 149 -352 486 -351
rect 569 -352 591 -351
rect 684 -352 745 -351
rect 758 -352 864 -351
rect 870 -352 913 -351
rect 86 -354 367 -353
rect 401 -354 815 -353
rect 877 -354 1025 -353
rect 149 -356 248 -355
rect 275 -356 451 -355
rect 555 -356 570 -355
rect 586 -356 759 -355
rect 765 -356 878 -355
rect 891 -356 913 -355
rect 191 -358 451 -357
rect 513 -358 556 -357
rect 730 -358 766 -357
rect 793 -358 892 -357
rect 198 -360 262 -359
rect 282 -360 325 -359
rect 366 -360 552 -359
rect 688 -360 794 -359
rect 800 -360 843 -359
rect 114 -362 283 -361
rect 404 -362 836 -361
rect 128 -364 199 -363
rect 219 -364 566 -363
rect 611 -364 689 -363
rect 695 -364 801 -363
rect 33 -366 129 -365
rect 240 -366 248 -365
rect 429 -366 458 -365
rect 492 -366 514 -365
rect 611 -366 675 -365
rect 719 -366 731 -365
rect 737 -366 752 -365
rect 240 -368 937 -367
rect 429 -370 521 -369
rect 625 -370 696 -369
rect 737 -370 941 -369
rect 492 -372 955 -371
rect 495 -374 552 -373
rect 597 -374 626 -373
rect 660 -374 675 -373
rect 856 -374 941 -373
rect 562 -376 598 -375
rect 646 -376 661 -375
rect 779 -376 857 -375
rect 338 -378 647 -377
rect 779 -378 962 -377
rect 562 -380 710 -379
rect 667 -382 710 -381
rect 604 -384 668 -383
rect 387 -386 605 -385
rect 373 -388 388 -387
rect 310 -390 374 -389
rect 233 -392 311 -391
rect 177 -394 234 -393
rect 16 -405 139 -404
rect 142 -405 150 -404
rect 180 -405 199 -404
rect 233 -405 276 -404
rect 282 -405 286 -404
rect 306 -405 325 -404
rect 331 -405 405 -404
rect 422 -405 755 -404
rect 800 -405 1046 -404
rect 1066 -405 1140 -404
rect 16 -407 52 -406
rect 58 -407 199 -406
rect 233 -407 566 -406
rect 576 -407 591 -406
rect 600 -407 871 -406
rect 877 -407 1102 -406
rect 1108 -407 1151 -406
rect 23 -409 391 -408
rect 401 -409 794 -408
rect 800 -409 808 -408
rect 863 -409 1116 -408
rect 23 -411 115 -410
rect 142 -411 174 -410
rect 191 -411 206 -410
rect 247 -411 251 -410
rect 254 -411 321 -410
rect 331 -411 486 -410
rect 502 -411 997 -410
rect 1003 -411 1088 -410
rect 37 -413 213 -412
rect 247 -413 262 -412
rect 268 -413 279 -412
rect 282 -413 290 -412
rect 296 -413 325 -412
rect 338 -413 430 -412
rect 436 -413 493 -412
rect 509 -413 696 -412
rect 740 -413 1081 -412
rect 51 -415 111 -414
rect 128 -415 192 -414
rect 219 -415 297 -414
rect 317 -415 451 -414
rect 478 -415 493 -414
rect 523 -415 899 -414
rect 919 -415 997 -414
rect 1010 -415 1109 -414
rect 58 -417 80 -416
rect 107 -417 115 -416
rect 128 -417 157 -416
rect 219 -417 304 -416
rect 317 -417 381 -416
rect 425 -417 1067 -416
rect 65 -419 90 -418
rect 145 -419 209 -418
rect 240 -419 339 -418
rect 341 -419 346 -418
rect 359 -419 416 -418
rect 429 -419 552 -418
rect 586 -419 717 -418
rect 730 -419 920 -418
rect 947 -419 1039 -418
rect 1041 -419 1053 -418
rect 44 -421 948 -420
rect 954 -421 1053 -420
rect 44 -423 279 -422
rect 285 -423 290 -422
rect 345 -423 500 -422
rect 548 -423 1032 -422
rect 65 -425 353 -424
rect 366 -425 437 -424
rect 485 -425 528 -424
rect 590 -425 598 -424
rect 646 -425 955 -424
rect 975 -425 1095 -424
rect 72 -427 136 -426
rect 156 -427 412 -426
rect 478 -427 598 -426
rect 639 -427 647 -426
rect 660 -427 696 -426
rect 709 -427 717 -426
rect 744 -427 878 -426
rect 905 -427 1011 -426
rect 1017 -427 1123 -426
rect 30 -429 661 -428
rect 674 -429 710 -428
rect 744 -429 759 -428
rect 772 -429 1004 -428
rect 1024 -429 1130 -428
rect 72 -431 87 -430
rect 93 -431 353 -430
rect 380 -431 902 -430
rect 926 -431 1025 -430
rect 12 -433 87 -432
rect 93 -433 122 -432
rect 240 -433 636 -432
rect 653 -433 675 -432
rect 688 -433 731 -432
rect 765 -433 773 -432
rect 793 -433 850 -432
rect 870 -433 913 -432
rect 926 -433 990 -432
rect 79 -435 514 -434
rect 527 -435 563 -434
rect 569 -435 766 -434
rect 779 -435 990 -434
rect 121 -437 164 -436
rect 254 -437 395 -436
rect 408 -437 416 -436
rect 457 -437 514 -436
rect 534 -437 570 -436
rect 625 -437 640 -436
rect 653 -437 738 -436
rect 807 -437 822 -436
rect 835 -437 976 -436
rect 982 -437 1074 -436
rect 149 -439 458 -438
rect 471 -439 780 -438
rect 814 -439 906 -438
rect 940 -439 1032 -438
rect 163 -441 178 -440
rect 268 -441 444 -440
rect 520 -441 822 -440
rect 835 -441 885 -440
rect 940 -441 962 -440
rect 982 -441 1060 -440
rect 170 -443 815 -442
rect 842 -443 864 -442
rect 884 -443 969 -442
rect 170 -445 227 -444
rect 303 -445 843 -444
rect 856 -445 969 -444
rect 177 -447 311 -446
rect 387 -447 395 -446
rect 408 -447 1018 -446
rect 310 -449 580 -448
rect 604 -449 626 -448
rect 681 -449 913 -448
rect 933 -449 962 -448
rect 443 -451 465 -450
rect 474 -451 857 -450
rect 891 -451 934 -450
rect 464 -453 738 -452
rect 828 -453 892 -452
rect 520 -455 668 -454
rect 681 -455 1049 -454
rect 534 -457 542 -456
rect 604 -457 619 -456
rect 632 -457 668 -456
rect 688 -457 703 -456
rect 723 -457 759 -456
rect 786 -457 829 -456
rect 229 -459 542 -458
rect 583 -459 619 -458
rect 723 -459 850 -458
rect 366 -461 584 -460
rect 751 -461 787 -460
rect 404 -463 703 -462
rect 9 -474 311 -473
rect 324 -474 346 -473
rect 348 -474 636 -473
rect 660 -474 969 -473
rect 975 -474 1144 -473
rect 1174 -474 1179 -473
rect 16 -476 111 -475
rect 135 -476 143 -475
rect 156 -476 531 -475
rect 537 -476 1046 -475
rect 16 -478 101 -477
rect 107 -478 255 -477
rect 261 -478 279 -477
rect 296 -478 311 -477
rect 397 -478 521 -477
rect 527 -478 990 -477
rect 1045 -478 1060 -477
rect 37 -480 304 -479
rect 401 -480 514 -479
rect 527 -480 535 -479
rect 562 -480 1123 -479
rect 37 -482 202 -481
rect 205 -482 227 -481
rect 240 -482 297 -481
rect 352 -482 402 -481
rect 436 -482 601 -481
rect 632 -482 1130 -481
rect 23 -484 206 -483
rect 219 -484 391 -483
rect 415 -484 437 -483
rect 450 -484 664 -483
rect 695 -484 738 -483
rect 751 -484 857 -483
rect 870 -484 969 -483
rect 975 -484 997 -483
rect 1059 -484 1109 -483
rect 1122 -484 1140 -483
rect 23 -486 31 -485
rect 72 -486 276 -485
rect 289 -486 304 -485
rect 380 -486 514 -485
rect 565 -486 1095 -485
rect 58 -488 381 -487
rect 415 -488 479 -487
rect 506 -488 731 -487
rect 733 -488 1102 -487
rect 58 -490 374 -489
rect 450 -490 486 -489
rect 583 -490 591 -489
rect 593 -490 1116 -489
rect 79 -492 500 -491
rect 586 -492 1004 -491
rect 1010 -492 1102 -491
rect 1115 -492 1151 -491
rect 86 -494 948 -493
rect 961 -494 983 -493
rect 989 -494 1025 -493
rect 86 -496 115 -495
rect 142 -496 367 -495
rect 457 -496 843 -495
rect 961 -496 1018 -495
rect 93 -498 157 -497
rect 166 -498 1067 -497
rect 93 -500 122 -499
rect 170 -500 220 -499
rect 240 -500 248 -499
rect 261 -500 430 -499
rect 460 -500 941 -499
rect 996 -500 1039 -499
rect 100 -502 129 -501
rect 149 -502 171 -501
rect 177 -502 255 -501
rect 289 -502 321 -501
rect 331 -502 374 -501
rect 429 -502 510 -501
rect 611 -502 857 -501
rect 884 -502 1067 -501
rect 44 -504 332 -503
rect 443 -504 510 -503
rect 548 -504 612 -503
rect 632 -504 654 -503
rect 660 -504 941 -503
rect 1003 -504 1053 -503
rect 44 -506 318 -505
rect 387 -506 1053 -505
rect 110 -508 178 -507
rect 191 -508 325 -507
rect 471 -508 570 -507
rect 604 -508 654 -507
rect 723 -508 906 -507
rect 1010 -508 1032 -507
rect 33 -510 605 -509
rect 730 -510 1025 -509
rect 1031 -510 1081 -509
rect 114 -512 395 -511
rect 478 -512 493 -511
rect 502 -512 724 -511
rect 754 -512 815 -511
rect 828 -512 843 -511
rect 849 -512 885 -511
rect 898 -512 906 -511
rect 1017 -512 1074 -511
rect 1080 -512 1088 -511
rect 128 -514 409 -513
rect 485 -514 573 -513
rect 597 -514 1088 -513
rect 152 -516 570 -515
rect 597 -516 878 -515
rect 926 -516 1074 -515
rect 163 -518 472 -517
rect 492 -518 629 -517
rect 765 -518 1095 -517
rect 191 -520 696 -519
rect 779 -520 829 -519
rect 835 -520 948 -519
rect 247 -522 405 -521
rect 422 -522 836 -521
rect 877 -522 913 -521
rect 121 -524 423 -523
rect 551 -524 927 -523
rect 268 -526 444 -525
rect 688 -526 766 -525
rect 786 -526 815 -525
rect 821 -526 899 -525
rect 268 -528 283 -527
rect 317 -528 360 -527
rect 667 -528 689 -527
rect 716 -528 780 -527
rect 793 -528 850 -527
rect 891 -528 913 -527
rect 138 -530 360 -529
rect 639 -530 668 -529
rect 681 -530 717 -529
rect 744 -530 787 -529
rect 800 -530 822 -529
rect 863 -530 892 -529
rect 233 -532 283 -531
rect 355 -532 794 -531
rect 807 -532 1039 -531
rect 51 -534 234 -533
rect 408 -534 801 -533
rect 863 -534 955 -533
rect 51 -536 339 -535
rect 548 -536 682 -535
rect 744 -536 759 -535
rect 772 -536 808 -535
rect 933 -536 955 -535
rect 338 -538 391 -537
rect 625 -538 640 -537
rect 702 -538 773 -537
rect 919 -538 934 -537
rect 562 -540 920 -539
rect 674 -542 703 -541
rect 709 -542 759 -541
rect 646 -544 675 -543
rect 709 -544 871 -543
rect 618 -546 647 -545
rect 576 -548 619 -547
rect 65 -550 577 -549
rect 65 -552 199 -551
rect 198 -554 465 -553
rect 215 -556 465 -555
rect 194 -558 216 -557
rect 2 -569 510 -568
rect 534 -569 542 -568
rect 548 -569 871 -568
rect 1059 -569 1109 -568
rect 9 -571 73 -570
rect 82 -571 710 -570
rect 712 -571 899 -570
rect 1087 -571 1130 -570
rect 9 -573 381 -572
rect 408 -573 836 -572
rect 842 -573 899 -572
rect 1024 -573 1088 -572
rect 1101 -573 1137 -572
rect 16 -575 871 -574
rect 975 -575 1025 -574
rect 16 -577 87 -576
rect 121 -577 563 -576
rect 569 -577 1039 -576
rect 23 -579 542 -578
rect 548 -579 1060 -578
rect 23 -581 419 -580
rect 443 -581 573 -580
rect 600 -581 885 -580
rect 919 -581 1039 -580
rect 30 -583 80 -582
rect 86 -583 297 -582
rect 338 -583 388 -582
rect 464 -583 692 -582
rect 733 -583 745 -582
rect 751 -583 920 -582
rect 968 -583 976 -582
rect 30 -585 262 -584
rect 268 -585 353 -584
rect 380 -585 493 -584
rect 506 -585 1102 -584
rect 33 -587 412 -586
rect 471 -587 598 -586
rect 604 -587 1067 -586
rect 37 -589 188 -588
rect 191 -589 227 -588
rect 254 -589 503 -588
rect 513 -589 563 -588
rect 604 -589 962 -588
rect 1003 -589 1067 -588
rect 37 -591 101 -590
rect 107 -591 262 -590
rect 275 -591 356 -590
rect 436 -591 472 -590
rect 478 -591 514 -590
rect 551 -591 857 -590
rect 877 -591 962 -590
rect 44 -593 465 -592
rect 555 -593 570 -592
rect 625 -593 682 -592
rect 688 -593 745 -592
rect 751 -593 759 -592
rect 761 -593 1011 -592
rect 44 -595 94 -594
rect 107 -595 118 -594
rect 121 -595 202 -594
rect 205 -595 398 -594
rect 415 -595 437 -594
rect 555 -595 640 -594
rect 656 -595 1081 -594
rect 54 -597 801 -596
rect 807 -597 878 -596
rect 926 -597 969 -596
rect 982 -597 1011 -596
rect 1017 -597 1081 -596
rect 65 -599 507 -598
rect 611 -599 640 -598
rect 660 -599 1074 -598
rect 68 -601 458 -600
rect 628 -601 731 -600
rect 765 -601 857 -600
rect 926 -601 948 -600
rect 954 -601 1004 -600
rect 1045 -601 1074 -600
rect 72 -603 374 -602
rect 450 -603 458 -602
rect 632 -603 682 -602
rect 723 -603 808 -602
rect 821 -603 843 -602
rect 849 -603 955 -602
rect 989 -603 1046 -602
rect 79 -605 836 -604
rect 905 -605 948 -604
rect 989 -605 1053 -604
rect 75 -607 906 -606
rect 933 -607 983 -606
rect 996 -607 1053 -606
rect 93 -609 608 -608
rect 611 -609 633 -608
rect 646 -609 661 -608
rect 765 -609 780 -608
rect 793 -609 885 -608
rect 940 -609 1018 -608
rect 114 -611 451 -610
rect 485 -611 647 -610
rect 674 -611 780 -610
rect 800 -611 1095 -610
rect 128 -613 447 -612
rect 537 -613 724 -612
rect 772 -613 822 -612
rect 863 -613 997 -612
rect 1031 -613 1095 -612
rect 149 -615 409 -614
rect 663 -615 1032 -614
rect 152 -617 297 -616
rect 331 -617 353 -616
rect 373 -617 482 -616
rect 667 -617 675 -616
rect 695 -617 794 -616
rect 814 -617 850 -616
rect 166 -619 913 -618
rect 170 -621 199 -620
rect 212 -621 367 -620
rect 390 -621 864 -620
rect 891 -621 913 -620
rect 51 -623 367 -622
rect 583 -623 668 -622
rect 695 -623 759 -622
rect 828 -623 892 -622
rect 170 -625 248 -624
rect 289 -625 486 -624
rect 583 -625 619 -624
rect 716 -625 773 -624
rect 786 -625 829 -624
rect 177 -627 227 -626
rect 233 -627 255 -626
rect 289 -627 608 -626
rect 653 -627 717 -626
rect 737 -627 815 -626
rect 100 -629 738 -628
rect 177 -631 185 -630
rect 212 -631 318 -630
rect 341 -631 941 -630
rect 142 -633 318 -632
rect 345 -633 395 -632
rect 422 -633 654 -632
rect 58 -635 346 -634
rect 348 -635 493 -634
rect 576 -635 619 -634
rect 58 -637 241 -636
rect 247 -637 283 -636
rect 359 -637 787 -636
rect 135 -639 241 -638
rect 282 -639 321 -638
rect 359 -639 402 -638
rect 422 -639 615 -638
rect 135 -641 164 -640
rect 184 -641 269 -640
rect 401 -641 430 -640
rect 527 -641 577 -640
rect 142 -643 591 -642
rect 163 -645 206 -644
rect 219 -645 276 -644
rect 324 -645 430 -644
rect 499 -645 528 -644
rect 156 -647 220 -646
rect 310 -647 325 -646
rect 520 -647 591 -646
rect 310 -649 332 -648
rect 16 -660 129 -659
rect 149 -660 234 -659
rect 254 -660 416 -659
rect 425 -660 608 -659
rect 611 -660 633 -659
rect 691 -660 976 -659
rect 1003 -660 1007 -659
rect 1038 -660 1042 -659
rect 1059 -660 1151 -659
rect 1178 -660 1186 -659
rect 16 -662 185 -661
rect 187 -662 237 -661
rect 254 -662 269 -661
rect 324 -662 339 -661
rect 408 -662 794 -661
rect 807 -662 811 -661
rect 933 -662 1018 -661
rect 1038 -662 1116 -661
rect 23 -664 423 -663
rect 439 -664 636 -663
rect 747 -664 780 -663
rect 807 -664 815 -663
rect 933 -664 948 -663
rect 975 -664 1025 -663
rect 1045 -664 1060 -663
rect 1087 -664 1116 -663
rect 30 -666 479 -665
rect 481 -666 920 -665
rect 947 -666 983 -665
rect 996 -666 1018 -665
rect 1087 -666 1130 -665
rect 37 -668 132 -667
rect 142 -668 339 -667
rect 345 -668 479 -667
rect 513 -668 661 -667
rect 695 -668 780 -667
rect 814 -668 878 -667
rect 898 -668 920 -667
rect 968 -668 997 -667
rect 1003 -668 1053 -667
rect 1090 -668 1172 -667
rect 37 -670 122 -669
rect 142 -670 192 -669
rect 205 -670 398 -669
rect 443 -670 1025 -669
rect 1031 -670 1053 -669
rect 1101 -670 1130 -669
rect 44 -672 118 -671
rect 159 -672 598 -671
rect 604 -672 990 -671
rect 1010 -672 1046 -671
rect 1080 -672 1102 -671
rect 1108 -672 1144 -671
rect 44 -674 199 -673
rect 208 -674 213 -673
rect 233 -674 262 -673
rect 268 -674 692 -673
rect 758 -674 773 -673
rect 842 -674 899 -673
rect 940 -674 969 -673
rect 1073 -674 1081 -673
rect 1108 -674 1137 -673
rect 51 -676 192 -675
rect 198 -676 304 -675
rect 324 -676 374 -675
rect 380 -676 514 -675
rect 523 -676 1165 -675
rect 54 -678 66 -677
rect 72 -678 447 -677
rect 464 -678 475 -677
rect 502 -678 843 -677
rect 940 -678 955 -677
rect 961 -678 990 -677
rect 1073 -678 1095 -677
rect 1122 -678 1137 -677
rect 58 -680 262 -679
rect 303 -680 451 -679
rect 464 -680 710 -679
rect 905 -680 955 -679
rect 58 -682 353 -681
rect 366 -682 444 -681
rect 450 -682 472 -681
rect 516 -682 1123 -681
rect 65 -684 524 -683
rect 551 -684 857 -683
rect 884 -684 906 -683
rect 912 -684 962 -683
rect 72 -686 213 -685
rect 317 -686 353 -685
rect 366 -686 521 -685
rect 551 -686 584 -685
rect 597 -686 836 -685
rect 891 -686 913 -685
rect 79 -688 97 -687
rect 100 -688 220 -687
rect 310 -688 318 -687
rect 345 -688 437 -687
rect 499 -688 885 -687
rect 79 -690 108 -689
rect 114 -690 136 -689
rect 152 -690 374 -689
rect 380 -690 419 -689
rect 485 -690 500 -689
rect 569 -690 584 -689
rect 604 -690 864 -689
rect 870 -690 892 -689
rect 82 -692 549 -691
rect 576 -692 654 -691
rect 660 -692 717 -691
rect 765 -692 864 -691
rect 86 -694 150 -693
rect 156 -694 1011 -693
rect 89 -696 206 -695
rect 219 -696 276 -695
rect 506 -696 577 -695
rect 614 -696 927 -695
rect 93 -698 108 -697
rect 135 -698 836 -697
rect 93 -700 164 -699
rect 184 -700 332 -699
rect 506 -700 801 -699
rect 821 -700 857 -699
rect 103 -702 556 -701
rect 646 -702 710 -701
rect 716 -702 794 -701
rect 800 -702 829 -701
rect 156 -704 171 -703
rect 240 -704 486 -703
rect 534 -704 570 -703
rect 646 -704 682 -703
rect 688 -704 696 -703
rect 702 -704 773 -703
rect 163 -706 248 -705
rect 275 -706 283 -705
rect 467 -706 822 -705
rect 170 -708 360 -707
rect 527 -708 535 -707
rect 541 -708 556 -707
rect 667 -708 682 -707
rect 688 -708 983 -707
rect 1041 -708 1095 -707
rect 240 -710 297 -709
rect 429 -710 542 -709
rect 639 -710 668 -709
rect 730 -710 927 -709
rect 282 -712 395 -711
rect 401 -712 430 -711
rect 527 -712 619 -711
rect 639 -712 703 -711
rect 730 -712 787 -711
rect 33 -714 395 -713
rect 411 -714 787 -713
rect 289 -716 297 -715
rect 562 -716 619 -715
rect 744 -716 766 -715
rect 289 -718 493 -717
rect 562 -718 591 -717
rect 744 -718 871 -717
rect 341 -720 591 -719
rect 751 -720 829 -719
rect 492 -722 724 -721
rect 625 -724 752 -723
rect 625 -726 1112 -725
rect 674 -728 724 -727
rect 656 -730 675 -729
rect 9 -741 139 -740
rect 149 -741 584 -740
rect 600 -741 941 -740
rect 1038 -741 1088 -740
rect 1108 -741 1137 -740
rect 1143 -741 1193 -740
rect 9 -743 80 -742
rect 86 -743 132 -742
rect 163 -743 363 -742
rect 373 -743 384 -742
rect 404 -743 500 -742
rect 502 -743 528 -742
rect 583 -743 748 -742
rect 782 -743 1004 -742
rect 1031 -743 1039 -742
rect 1052 -743 1109 -742
rect 1122 -743 1179 -742
rect 1185 -743 1214 -742
rect 16 -745 339 -744
rect 359 -745 1053 -744
rect 1059 -745 1123 -744
rect 1129 -745 1186 -744
rect 16 -747 367 -746
rect 373 -747 388 -746
rect 408 -747 626 -746
rect 639 -747 818 -746
rect 821 -747 853 -746
rect 884 -747 1004 -746
rect 1059 -747 1091 -746
rect 1101 -747 1144 -746
rect 1150 -747 1161 -746
rect 1164 -747 1200 -746
rect 23 -749 402 -748
rect 411 -749 416 -748
rect 439 -749 472 -748
rect 495 -749 948 -748
rect 968 -749 1032 -748
rect 1080 -749 1137 -748
rect 1171 -749 1221 -748
rect 23 -751 346 -750
rect 387 -751 570 -750
rect 572 -751 1165 -750
rect 30 -753 171 -752
rect 173 -753 206 -752
rect 212 -753 426 -752
rect 464 -753 479 -752
rect 513 -753 636 -752
rect 642 -753 864 -752
rect 926 -753 941 -752
rect 947 -753 955 -752
rect 989 -753 1081 -752
rect 1115 -753 1151 -752
rect 37 -755 125 -754
rect 177 -755 185 -754
rect 187 -755 542 -754
rect 625 -755 878 -754
rect 954 -755 1158 -754
rect 37 -757 118 -756
rect 156 -757 178 -756
rect 191 -757 255 -756
rect 331 -757 437 -756
rect 485 -757 514 -756
rect 520 -757 969 -756
rect 982 -757 990 -756
rect 996 -757 1088 -756
rect 58 -759 346 -758
rect 366 -759 521 -758
rect 523 -759 661 -758
rect 663 -759 1130 -758
rect 58 -761 94 -760
rect 100 -761 213 -760
rect 338 -761 598 -760
rect 604 -761 1158 -760
rect 65 -763 332 -762
rect 380 -763 661 -762
rect 688 -763 899 -762
rect 933 -763 983 -762
rect 996 -763 1025 -762
rect 1073 -763 1172 -762
rect 44 -765 381 -764
rect 394 -765 885 -764
rect 1010 -765 1116 -764
rect 44 -767 269 -766
rect 341 -767 1025 -766
rect 1073 -767 1095 -766
rect 65 -769 507 -768
rect 527 -769 535 -768
rect 541 -769 556 -768
rect 565 -769 934 -768
rect 1017 -769 1095 -768
rect 79 -771 426 -770
rect 499 -771 535 -770
rect 569 -771 1011 -770
rect 1017 -771 1067 -770
rect 86 -773 318 -772
rect 394 -773 430 -772
rect 506 -773 577 -772
rect 590 -773 605 -772
rect 688 -773 696 -772
rect 698 -773 1102 -772
rect 93 -775 241 -774
rect 268 -775 311 -774
rect 317 -775 353 -774
rect 415 -775 643 -774
rect 716 -775 857 -774
rect 870 -775 878 -774
rect 100 -777 136 -776
rect 138 -777 157 -776
rect 163 -777 255 -776
rect 429 -777 892 -776
rect 114 -779 122 -778
rect 135 -779 290 -778
rect 457 -779 577 -778
rect 590 -779 619 -778
rect 744 -779 976 -778
rect 170 -781 241 -780
rect 247 -781 311 -780
rect 443 -781 458 -780
rect 485 -781 696 -780
rect 786 -781 899 -780
rect 191 -783 297 -782
rect 443 -783 451 -782
rect 492 -783 717 -782
rect 786 -783 808 -782
rect 842 -783 927 -782
rect 226 -785 248 -784
rect 289 -785 353 -784
rect 548 -785 745 -784
rect 779 -785 808 -784
rect 835 -785 843 -784
rect 849 -785 864 -784
rect 891 -785 906 -784
rect 128 -787 227 -786
rect 296 -787 612 -786
rect 656 -787 976 -786
rect 303 -789 451 -788
rect 548 -789 563 -788
rect 597 -789 752 -788
rect 779 -789 871 -788
rect 198 -791 304 -790
rect 555 -791 1067 -790
rect 107 -793 199 -792
rect 562 -793 731 -792
rect 751 -793 829 -792
rect 849 -793 1207 -792
rect 107 -795 220 -794
rect 474 -795 829 -794
rect 856 -795 920 -794
rect 219 -797 654 -796
rect 793 -797 822 -796
rect 912 -797 920 -796
rect 611 -799 668 -798
rect 772 -799 794 -798
rect 800 -799 906 -798
rect 912 -799 962 -798
rect 478 -801 773 -800
rect 814 -801 836 -800
rect 632 -803 962 -802
rect 632 -805 682 -804
rect 758 -805 801 -804
rect 51 -807 682 -806
rect 51 -809 283 -808
rect 621 -809 759 -808
rect 233 -811 283 -810
rect 667 -811 710 -810
rect 233 -813 276 -812
rect 646 -813 710 -812
rect 261 -815 276 -814
rect 646 -815 675 -814
rect 674 -817 724 -816
rect 723 -819 731 -818
rect 19 -830 314 -829
rect 355 -830 1004 -829
rect 30 -832 118 -831
rect 121 -832 1102 -831
rect 33 -834 171 -833
rect 198 -834 500 -833
rect 523 -834 591 -833
rect 618 -834 906 -833
rect 996 -834 1000 -833
rect 1003 -834 1039 -833
rect 44 -836 570 -835
rect 590 -836 633 -835
rect 639 -836 703 -835
rect 726 -836 1067 -835
rect 44 -838 290 -837
rect 359 -838 384 -837
rect 387 -838 479 -837
rect 485 -838 521 -837
rect 555 -838 612 -837
rect 656 -838 731 -837
rect 758 -838 850 -837
rect 905 -838 990 -837
rect 996 -838 1011 -837
rect 1017 -838 1067 -837
rect 37 -840 388 -839
rect 394 -840 496 -839
rect 558 -840 633 -839
rect 656 -840 1081 -839
rect 51 -842 265 -841
rect 296 -842 556 -841
rect 562 -842 605 -841
rect 611 -842 1095 -841
rect 51 -844 192 -843
rect 198 -844 234 -843
rect 296 -844 325 -843
rect 362 -844 458 -843
rect 464 -844 622 -843
rect 660 -844 668 -843
rect 695 -844 1088 -843
rect 1094 -844 1179 -843
rect 16 -846 192 -845
rect 205 -846 605 -845
rect 621 -846 766 -845
rect 779 -846 829 -845
rect 968 -846 1039 -845
rect 1073 -846 1088 -845
rect 1178 -846 1221 -845
rect 58 -848 62 -847
rect 86 -848 353 -847
rect 380 -848 1102 -847
rect 58 -850 241 -849
rect 289 -850 829 -849
rect 968 -850 983 -849
rect 989 -850 1130 -849
rect 86 -852 682 -851
rect 695 -852 717 -851
rect 730 -852 801 -851
rect 814 -852 1193 -851
rect 5 -854 815 -853
rect 982 -854 1116 -853
rect 1129 -854 1186 -853
rect 1192 -854 1214 -853
rect 93 -856 241 -855
rect 292 -856 801 -855
rect 1017 -856 1060 -855
rect 1073 -856 1137 -855
rect 93 -858 101 -857
rect 114 -858 1032 -857
rect 1059 -858 1123 -857
rect 117 -860 381 -859
rect 422 -860 507 -859
rect 569 -860 584 -859
rect 663 -860 668 -859
rect 681 -860 885 -859
rect 999 -860 1011 -859
rect 1024 -860 1116 -859
rect 1122 -860 1172 -859
rect 121 -862 615 -861
rect 698 -862 1165 -861
rect 1171 -862 1207 -861
rect 124 -864 227 -863
rect 324 -864 332 -863
rect 352 -864 437 -863
rect 450 -864 458 -863
rect 464 -864 503 -863
rect 506 -864 577 -863
rect 583 -864 689 -863
rect 702 -864 745 -863
rect 751 -864 766 -863
rect 863 -864 885 -863
rect 1024 -864 1109 -863
rect 1164 -864 1200 -863
rect 135 -866 346 -865
rect 425 -866 626 -865
rect 674 -866 689 -865
rect 716 -866 773 -865
rect 863 -866 892 -865
rect 1031 -866 1046 -865
rect 1080 -866 1151 -865
rect 23 -868 426 -867
rect 429 -868 745 -867
rect 751 -868 794 -867
rect 856 -868 892 -867
rect 1045 -868 1144 -867
rect 23 -870 220 -869
rect 226 -870 279 -869
rect 317 -870 332 -869
rect 429 -870 444 -869
rect 471 -870 724 -869
rect 758 -870 808 -869
rect 835 -870 857 -869
rect 870 -870 1109 -869
rect 107 -872 318 -871
rect 436 -872 598 -871
rect 600 -872 794 -871
rect 807 -872 843 -871
rect 870 -872 962 -871
rect 65 -874 598 -873
rect 674 -874 1053 -873
rect 65 -876 535 -875
rect 576 -876 647 -875
rect 677 -876 836 -875
rect 842 -876 878 -875
rect 898 -876 1053 -875
rect 79 -878 108 -877
rect 149 -878 444 -877
rect 471 -878 671 -877
rect 772 -878 822 -877
rect 877 -878 920 -877
rect 37 -880 80 -879
rect 163 -880 1158 -879
rect 156 -882 164 -881
rect 177 -882 234 -881
rect 485 -882 514 -881
rect 534 -882 549 -881
rect 646 -882 710 -881
rect 817 -882 962 -881
rect 142 -884 178 -883
rect 205 -884 248 -883
rect 415 -884 549 -883
rect 709 -884 738 -883
rect 128 -886 143 -885
rect 149 -886 248 -885
rect 348 -886 416 -885
rect 513 -886 528 -885
rect 544 -886 920 -885
rect 9 -888 129 -887
rect 156 -888 493 -887
rect 527 -888 654 -887
rect 737 -888 934 -887
rect 9 -890 255 -889
rect 366 -890 493 -889
rect 933 -890 941 -889
rect 212 -892 395 -891
rect 926 -892 941 -891
rect 212 -894 409 -893
rect 926 -894 955 -893
rect 219 -896 283 -895
rect 366 -896 374 -895
rect 912 -896 955 -895
rect 40 -898 283 -897
rect 912 -898 1091 -897
rect 254 -900 339 -899
rect 268 -902 409 -901
rect 268 -904 276 -903
rect 310 -904 339 -903
rect 310 -906 451 -905
rect 2 -917 87 -916
rect 96 -917 486 -916
rect 502 -917 514 -916
rect 548 -917 682 -916
rect 684 -917 1116 -916
rect 1136 -917 1179 -916
rect 19 -919 815 -918
rect 824 -919 1088 -918
rect 1101 -919 1116 -918
rect 1150 -919 1165 -918
rect 30 -921 171 -920
rect 205 -921 577 -920
rect 597 -921 871 -920
rect 898 -921 1123 -920
rect 1157 -921 1172 -920
rect 33 -923 500 -922
rect 506 -923 514 -922
rect 548 -923 563 -922
rect 597 -923 829 -922
rect 1108 -923 1172 -922
rect 37 -925 605 -924
rect 618 -925 703 -924
rect 716 -925 1144 -924
rect 1164 -925 1193 -924
rect 40 -927 325 -926
rect 345 -927 493 -926
rect 499 -927 899 -926
rect 1066 -927 1109 -926
rect 1122 -927 1130 -926
rect 1185 -927 1193 -926
rect 9 -929 325 -928
rect 348 -929 409 -928
rect 415 -929 493 -928
rect 555 -929 1102 -928
rect 40 -931 577 -930
rect 628 -931 710 -930
rect 716 -931 731 -930
rect 737 -931 829 -930
rect 1052 -931 1130 -930
rect 44 -933 612 -932
rect 656 -933 990 -932
rect 1052 -933 1081 -932
rect 44 -935 101 -934
rect 117 -935 391 -934
rect 408 -935 559 -934
rect 562 -935 570 -934
rect 667 -935 696 -934
rect 702 -935 773 -934
rect 975 -935 1081 -934
rect 51 -937 115 -936
rect 142 -937 153 -936
rect 170 -937 209 -936
rect 219 -937 437 -936
rect 439 -937 633 -936
rect 674 -937 731 -936
rect 737 -937 787 -936
rect 975 -937 1018 -936
rect 51 -939 62 -938
rect 65 -939 556 -938
rect 632 -939 647 -938
rect 695 -939 871 -938
rect 989 -939 1032 -938
rect 58 -941 115 -940
rect 142 -941 265 -940
rect 268 -941 290 -940
rect 303 -941 311 -940
rect 331 -941 416 -940
rect 439 -941 860 -940
rect 996 -941 1032 -940
rect 58 -943 108 -942
rect 149 -943 234 -942
rect 247 -943 290 -942
rect 303 -943 734 -942
rect 772 -943 864 -942
rect 961 -943 997 -942
rect 1017 -943 1074 -942
rect 72 -945 713 -944
rect 786 -945 801 -944
rect 961 -945 1011 -944
rect 1038 -945 1074 -944
rect 79 -947 108 -946
rect 191 -947 220 -946
rect 233 -947 377 -946
rect 380 -947 654 -946
rect 709 -947 983 -946
rect 1010 -947 1095 -946
rect 79 -949 129 -948
rect 156 -949 192 -948
rect 212 -949 248 -948
rect 261 -949 332 -948
rect 362 -949 815 -948
rect 982 -949 1091 -948
rect 86 -951 94 -950
rect 121 -951 129 -950
rect 156 -951 199 -950
rect 240 -951 262 -950
rect 268 -951 367 -950
rect 373 -951 724 -950
rect 800 -951 857 -950
rect 1059 -951 1095 -950
rect 9 -953 122 -952
rect 177 -953 213 -952
rect 240 -953 255 -952
rect 275 -953 297 -952
rect 352 -953 367 -952
rect 380 -953 388 -952
rect 471 -953 570 -952
rect 607 -953 1039 -952
rect 23 -955 255 -954
rect 275 -955 283 -954
rect 296 -955 318 -954
rect 471 -955 584 -954
rect 625 -955 864 -954
rect 1024 -955 1060 -954
rect 23 -957 101 -956
rect 135 -957 353 -956
rect 478 -957 521 -956
rect 583 -957 661 -956
rect 723 -957 780 -956
rect 821 -957 1025 -956
rect 72 -959 199 -958
rect 317 -959 451 -958
rect 485 -959 528 -958
rect 544 -959 661 -958
rect 744 -959 780 -958
rect 821 -959 906 -958
rect 93 -961 1067 -960
rect 135 -963 615 -962
rect 653 -963 689 -962
rect 744 -963 794 -962
rect 905 -963 955 -962
rect 177 -965 185 -964
rect 359 -965 521 -964
rect 527 -965 535 -964
rect 688 -965 752 -964
rect 793 -965 808 -964
rect 954 -965 969 -964
rect 184 -967 283 -966
rect 443 -967 535 -966
rect 751 -967 850 -966
rect 968 -967 1046 -966
rect 422 -969 1046 -968
rect 422 -971 465 -970
rect 807 -971 878 -970
rect 429 -973 444 -972
rect 450 -973 591 -972
rect 849 -973 892 -972
rect 429 -975 458 -974
rect 590 -975 836 -974
rect 877 -975 920 -974
rect 457 -977 640 -976
rect 765 -977 892 -976
rect 758 -979 766 -978
rect 835 -979 948 -978
rect 65 -981 759 -980
rect 884 -981 920 -980
rect 933 -981 948 -980
rect 842 -983 934 -982
rect 842 -985 902 -984
rect 884 -987 927 -986
rect 926 -989 941 -988
rect 940 -991 1004 -990
rect 912 -993 1004 -992
rect 604 -995 913 -994
rect 9 -1006 94 -1005
rect 100 -1006 108 -1005
rect 121 -1006 339 -1005
rect 359 -1006 423 -1005
rect 464 -1006 514 -1005
rect 541 -1006 766 -1005
rect 810 -1006 955 -1005
rect 1129 -1006 1158 -1005
rect 37 -1008 66 -1007
rect 89 -1008 864 -1007
rect 884 -1008 888 -1007
rect 954 -1008 1116 -1007
rect 1136 -1008 1151 -1007
rect 40 -1010 545 -1009
rect 569 -1010 608 -1009
rect 625 -1010 724 -1009
rect 730 -1010 1095 -1009
rect 44 -1012 199 -1011
rect 208 -1012 213 -1011
rect 219 -1012 356 -1011
rect 362 -1012 1039 -1011
rect 1094 -1012 1172 -1011
rect 16 -1014 45 -1013
rect 58 -1014 73 -1013
rect 107 -1014 395 -1013
rect 401 -1014 514 -1013
rect 527 -1014 542 -1013
rect 597 -1014 643 -1013
rect 646 -1014 675 -1013
rect 681 -1014 706 -1013
rect 723 -1014 836 -1013
rect 856 -1014 1081 -1013
rect 16 -1016 104 -1015
rect 124 -1016 360 -1015
rect 457 -1016 528 -1015
rect 600 -1016 794 -1015
rect 856 -1016 878 -1015
rect 884 -1016 906 -1015
rect 1024 -1016 1039 -1015
rect 1069 -1016 1081 -1015
rect 30 -1018 220 -1017
rect 254 -1018 388 -1017
rect 443 -1018 458 -1017
rect 499 -1018 983 -1017
rect 996 -1018 1025 -1017
rect 30 -1020 143 -1019
rect 184 -1020 283 -1019
rect 289 -1020 321 -1019
rect 338 -1020 381 -1019
rect 429 -1020 444 -1019
rect 499 -1020 584 -1019
rect 604 -1020 692 -1019
rect 695 -1020 738 -1019
rect 751 -1020 766 -1019
rect 786 -1020 836 -1019
rect 859 -1020 1109 -1019
rect 61 -1022 549 -1021
rect 632 -1022 675 -1021
rect 681 -1022 689 -1021
rect 698 -1022 794 -1021
rect 863 -1022 899 -1021
rect 905 -1022 969 -1021
rect 982 -1022 1011 -1021
rect 65 -1024 409 -1023
rect 429 -1024 486 -1023
rect 502 -1024 1102 -1023
rect 72 -1026 276 -1025
rect 289 -1026 297 -1025
rect 317 -1026 423 -1025
rect 471 -1026 584 -1025
rect 639 -1026 1088 -1025
rect 79 -1028 283 -1027
rect 317 -1028 598 -1027
rect 639 -1028 654 -1027
rect 660 -1028 738 -1027
rect 751 -1028 822 -1027
rect 968 -1028 990 -1027
rect 996 -1028 1018 -1027
rect 1087 -1028 1123 -1027
rect 79 -1030 150 -1029
rect 187 -1030 780 -1029
rect 786 -1030 920 -1029
rect 989 -1030 1067 -1029
rect 1122 -1030 1168 -1029
rect 96 -1032 395 -1031
rect 408 -1032 416 -1031
rect 485 -1032 563 -1031
rect 649 -1032 892 -1031
rect 919 -1032 1074 -1031
rect 86 -1034 97 -1033
rect 114 -1034 143 -1033
rect 191 -1034 199 -1033
rect 205 -1034 472 -1033
rect 509 -1034 535 -1033
rect 653 -1034 703 -1033
rect 716 -1034 878 -1033
rect 891 -1034 913 -1033
rect 1010 -1034 1133 -1033
rect 2 -1036 206 -1035
rect 212 -1036 241 -1035
rect 268 -1036 374 -1035
rect 376 -1036 899 -1035
rect 912 -1036 927 -1035
rect 1017 -1036 1053 -1035
rect 170 -1038 269 -1037
rect 331 -1038 549 -1037
rect 572 -1038 927 -1037
rect 177 -1040 192 -1039
rect 226 -1040 276 -1039
rect 303 -1040 332 -1039
rect 373 -1040 479 -1039
rect 506 -1040 703 -1039
rect 716 -1040 773 -1039
rect 779 -1040 808 -1039
rect 821 -1040 871 -1039
rect 86 -1042 227 -1041
rect 233 -1042 255 -1041
rect 303 -1042 311 -1041
rect 380 -1042 437 -1041
rect 450 -1042 563 -1041
rect 660 -1042 668 -1041
rect 684 -1042 1060 -1041
rect 117 -1044 234 -1043
rect 240 -1044 265 -1043
rect 401 -1044 437 -1043
rect 450 -1044 612 -1043
rect 667 -1044 710 -1043
rect 733 -1044 1032 -1043
rect 1059 -1044 1074 -1043
rect 152 -1046 311 -1045
rect 415 -1046 622 -1045
rect 688 -1046 815 -1045
rect 842 -1046 871 -1045
rect 1031 -1046 1053 -1045
rect 156 -1048 178 -1047
rect 390 -1048 843 -1047
rect 156 -1050 164 -1049
rect 478 -1050 493 -1049
rect 534 -1050 934 -1049
rect 135 -1052 164 -1051
rect 201 -1052 934 -1051
rect 135 -1054 325 -1053
rect 345 -1054 493 -1053
rect 576 -1054 612 -1053
rect 709 -1054 745 -1053
rect 772 -1054 801 -1053
rect 814 -1054 850 -1053
rect 247 -1056 325 -1055
rect 345 -1056 353 -1055
rect 576 -1056 619 -1055
rect 744 -1056 829 -1055
rect 849 -1056 1046 -1055
rect 247 -1058 262 -1057
rect 352 -1058 591 -1057
rect 618 -1058 948 -1057
rect 520 -1060 591 -1059
rect 758 -1060 829 -1059
rect 887 -1060 1067 -1059
rect 173 -1062 521 -1061
rect 800 -1062 1144 -1061
rect 940 -1064 948 -1063
rect 940 -1066 962 -1065
rect 961 -1068 976 -1067
rect 61 -1070 976 -1069
rect 16 -1081 188 -1080
rect 219 -1081 447 -1080
rect 471 -1081 619 -1080
rect 632 -1081 696 -1080
rect 852 -1081 878 -1080
rect 884 -1081 888 -1080
rect 954 -1081 962 -1080
rect 978 -1081 1018 -1080
rect 1031 -1081 1039 -1080
rect 1041 -1081 1053 -1080
rect 1108 -1081 1123 -1080
rect 1185 -1081 1189 -1080
rect 23 -1083 150 -1082
rect 170 -1083 591 -1082
rect 600 -1083 731 -1082
rect 877 -1083 927 -1082
rect 940 -1083 962 -1082
rect 1006 -1083 1095 -1082
rect 30 -1085 265 -1084
rect 268 -1085 307 -1084
rect 355 -1085 598 -1084
rect 607 -1085 752 -1084
rect 884 -1085 899 -1084
rect 940 -1085 948 -1084
rect 1017 -1085 1025 -1084
rect 1045 -1085 1060 -1084
rect 30 -1087 45 -1086
rect 58 -1087 167 -1086
rect 170 -1087 178 -1086
rect 191 -1087 220 -1086
rect 247 -1087 269 -1086
rect 275 -1087 507 -1086
rect 509 -1087 850 -1086
rect 891 -1087 899 -1086
rect 947 -1087 1004 -1086
rect 1010 -1087 1025 -1086
rect 1048 -1087 1088 -1086
rect 37 -1089 300 -1088
rect 387 -1089 468 -1088
rect 485 -1089 629 -1088
rect 667 -1089 752 -1088
rect 887 -1089 892 -1088
rect 989 -1089 1011 -1088
rect 1080 -1089 1088 -1088
rect 37 -1091 129 -1090
rect 149 -1091 157 -1090
rect 177 -1091 213 -1090
rect 296 -1091 612 -1090
rect 621 -1091 633 -1090
rect 667 -1091 843 -1090
rect 982 -1091 990 -1090
rect 1073 -1091 1081 -1090
rect 44 -1093 451 -1092
rect 551 -1093 577 -1092
rect 586 -1093 927 -1092
rect 968 -1093 983 -1092
rect 65 -1095 69 -1094
rect 72 -1095 465 -1094
rect 499 -1095 577 -1094
rect 590 -1095 738 -1094
rect 842 -1095 871 -1094
rect 968 -1095 976 -1094
rect 72 -1097 83 -1096
rect 93 -1097 101 -1096
rect 121 -1097 353 -1096
rect 366 -1097 465 -1096
rect 499 -1097 556 -1096
rect 572 -1097 584 -1096
rect 604 -1097 612 -1096
rect 670 -1097 1032 -1096
rect 79 -1099 129 -1098
rect 156 -1099 535 -1098
rect 583 -1099 654 -1098
rect 681 -1099 696 -1098
rect 702 -1099 871 -1098
rect 100 -1101 118 -1100
rect 121 -1101 185 -1100
rect 191 -1101 325 -1100
rect 359 -1101 703 -1100
rect 709 -1101 738 -1100
rect 184 -1103 419 -1102
rect 422 -1103 472 -1102
rect 534 -1103 734 -1102
rect 212 -1105 332 -1104
rect 373 -1105 556 -1104
rect 646 -1105 710 -1104
rect 226 -1107 367 -1106
rect 387 -1107 514 -1106
rect 646 -1107 920 -1106
rect 226 -1109 248 -1108
rect 282 -1109 325 -1108
rect 338 -1109 374 -1108
rect 422 -1109 570 -1108
rect 688 -1109 724 -1108
rect 919 -1109 934 -1108
rect 240 -1111 360 -1110
rect 436 -1111 479 -1110
rect 513 -1111 528 -1110
rect 562 -1111 570 -1110
rect 688 -1111 801 -1110
rect 933 -1111 1067 -1110
rect 240 -1113 538 -1112
rect 723 -1113 829 -1112
rect 1003 -1113 1067 -1112
rect 275 -1115 283 -1114
rect 289 -1115 297 -1114
rect 317 -1115 682 -1114
rect 800 -1115 815 -1114
rect 821 -1115 829 -1114
rect 233 -1117 290 -1116
rect 303 -1117 318 -1116
rect 331 -1117 437 -1116
rect 443 -1117 486 -1116
rect 492 -1117 563 -1116
rect 744 -1117 822 -1116
rect 163 -1119 234 -1118
rect 338 -1119 416 -1118
rect 429 -1119 493 -1118
rect 527 -1119 542 -1118
rect 744 -1119 864 -1118
rect 401 -1121 430 -1120
rect 450 -1121 458 -1120
rect 478 -1121 808 -1120
rect 814 -1121 836 -1120
rect 205 -1123 458 -1122
rect 541 -1123 626 -1122
rect 653 -1123 836 -1122
rect 198 -1125 206 -1124
rect 261 -1125 402 -1124
rect 408 -1125 416 -1124
rect 793 -1125 864 -1124
rect 261 -1127 311 -1126
rect 779 -1127 794 -1126
rect 310 -1129 811 -1128
rect 772 -1131 780 -1130
rect 810 -1131 906 -1130
rect 758 -1133 773 -1132
rect 786 -1133 906 -1132
rect 716 -1135 787 -1134
rect 520 -1137 717 -1136
rect 758 -1137 766 -1136
rect 520 -1139 958 -1138
rect 548 -1141 766 -1140
rect 394 -1143 549 -1142
rect 380 -1145 395 -1144
rect 107 -1147 381 -1146
rect 107 -1149 143 -1148
rect 135 -1151 143 -1150
rect 135 -1153 409 -1152
rect 16 -1164 122 -1163
rect 149 -1164 164 -1163
rect 170 -1164 199 -1163
rect 226 -1164 269 -1163
rect 285 -1164 318 -1163
rect 331 -1164 353 -1163
rect 446 -1164 934 -1163
rect 975 -1164 1039 -1163
rect 1066 -1164 1123 -1163
rect 23 -1166 27 -1165
rect 30 -1166 157 -1165
rect 163 -1166 248 -1165
rect 254 -1166 668 -1165
rect 695 -1166 808 -1165
rect 828 -1166 937 -1165
rect 961 -1166 976 -1165
rect 989 -1166 1067 -1165
rect 1080 -1166 1130 -1165
rect 30 -1168 500 -1167
rect 506 -1168 556 -1167
rect 562 -1168 605 -1167
rect 618 -1168 657 -1167
rect 667 -1168 689 -1167
rect 695 -1168 766 -1167
rect 831 -1168 878 -1167
rect 884 -1168 962 -1167
rect 996 -1168 1004 -1167
rect 1010 -1168 1039 -1167
rect 1087 -1168 1116 -1167
rect 37 -1170 139 -1169
rect 152 -1170 479 -1169
rect 499 -1170 510 -1169
rect 544 -1170 885 -1169
rect 919 -1170 997 -1169
rect 1024 -1170 1053 -1169
rect 1101 -1170 1109 -1169
rect 37 -1172 727 -1171
rect 730 -1172 1081 -1171
rect 44 -1174 115 -1173
rect 117 -1174 122 -1173
rect 170 -1174 276 -1173
rect 352 -1174 594 -1173
rect 607 -1174 878 -1173
rect 926 -1174 1074 -1173
rect 58 -1176 157 -1175
rect 177 -1176 199 -1175
rect 229 -1176 360 -1175
rect 443 -1176 1011 -1175
rect 1031 -1176 1088 -1175
rect 51 -1178 59 -1177
rect 72 -1178 129 -1177
rect 184 -1178 346 -1177
rect 359 -1178 381 -1177
rect 478 -1178 486 -1177
rect 562 -1178 822 -1177
rect 842 -1178 920 -1177
rect 954 -1178 990 -1177
rect 1017 -1178 1032 -1177
rect 1059 -1178 1109 -1177
rect 65 -1180 73 -1179
rect 79 -1180 584 -1179
rect 586 -1180 724 -1179
rect 730 -1180 794 -1179
rect 814 -1180 843 -1179
rect 849 -1180 892 -1179
rect 940 -1180 1018 -1179
rect 51 -1182 66 -1181
rect 82 -1182 339 -1181
rect 429 -1182 584 -1181
rect 590 -1182 605 -1181
rect 625 -1182 1046 -1181
rect 89 -1184 136 -1183
rect 187 -1184 815 -1183
rect 863 -1184 979 -1183
rect 107 -1186 346 -1185
rect 429 -1186 647 -1185
rect 653 -1186 717 -1185
rect 765 -1186 857 -1185
rect 870 -1186 927 -1185
rect 968 -1186 1060 -1185
rect 61 -1188 969 -1187
rect 107 -1190 384 -1189
rect 450 -1190 486 -1189
rect 565 -1190 871 -1189
rect 891 -1190 913 -1189
rect 233 -1192 304 -1191
rect 306 -1192 339 -1191
rect 401 -1192 451 -1191
rect 569 -1192 619 -1191
rect 625 -1192 640 -1191
rect 646 -1192 675 -1191
rect 688 -1192 759 -1191
rect 772 -1192 1025 -1191
rect 131 -1194 759 -1193
rect 772 -1194 1095 -1193
rect 233 -1196 549 -1195
rect 555 -1196 570 -1195
rect 611 -1196 864 -1195
rect 898 -1196 941 -1195
rect 240 -1198 248 -1197
rect 254 -1198 811 -1197
rect 898 -1198 948 -1197
rect 240 -1200 290 -1199
rect 317 -1200 717 -1199
rect 744 -1200 913 -1199
rect 261 -1202 283 -1201
rect 289 -1202 297 -1201
rect 394 -1202 402 -1201
rect 597 -1202 745 -1201
rect 779 -1202 822 -1201
rect 166 -1204 395 -1203
rect 408 -1204 780 -1203
rect 786 -1204 794 -1203
rect 800 -1204 857 -1203
rect 212 -1206 297 -1205
rect 408 -1206 458 -1205
rect 509 -1206 801 -1205
rect 191 -1208 213 -1207
rect 268 -1208 311 -1207
rect 457 -1208 472 -1207
rect 534 -1208 598 -1207
rect 611 -1208 657 -1207
rect 674 -1208 738 -1207
rect 751 -1208 787 -1207
rect 191 -1210 521 -1209
rect 527 -1210 535 -1209
rect 660 -1210 738 -1209
rect 751 -1210 836 -1209
rect 275 -1212 374 -1211
rect 464 -1212 472 -1211
rect 513 -1212 521 -1211
rect 527 -1212 552 -1211
rect 681 -1212 948 -1211
rect 23 -1214 465 -1213
rect 541 -1214 836 -1213
rect 310 -1216 325 -1215
rect 436 -1216 514 -1215
rect 681 -1216 710 -1215
rect 324 -1218 388 -1217
rect 436 -1218 493 -1217
rect 632 -1218 710 -1217
rect 492 -1220 724 -1219
rect 576 -1222 633 -1221
rect 702 -1222 955 -1221
rect 366 -1224 577 -1223
rect 366 -1226 374 -1225
rect 415 -1226 703 -1225
rect 415 -1228 829 -1227
rect 30 -1239 566 -1238
rect 569 -1239 727 -1238
rect 772 -1239 822 -1238
rect 828 -1239 1018 -1238
rect 47 -1241 178 -1240
rect 180 -1241 465 -1240
rect 481 -1241 864 -1240
rect 866 -1241 906 -1240
rect 999 -1241 1032 -1240
rect 68 -1243 73 -1242
rect 86 -1243 164 -1242
rect 177 -1243 206 -1242
rect 212 -1243 391 -1242
rect 394 -1243 776 -1242
rect 807 -1243 1032 -1242
rect 72 -1245 388 -1244
rect 394 -1245 468 -1244
rect 509 -1245 535 -1244
rect 541 -1245 580 -1244
rect 590 -1245 1060 -1244
rect 93 -1247 97 -1246
rect 114 -1247 129 -1246
rect 149 -1247 563 -1246
rect 590 -1247 619 -1246
rect 642 -1247 836 -1246
rect 905 -1247 1053 -1246
rect 1059 -1247 1116 -1246
rect 16 -1249 150 -1248
rect 163 -1249 290 -1248
rect 324 -1249 381 -1248
rect 387 -1249 409 -1248
rect 443 -1249 479 -1248
rect 544 -1249 948 -1248
rect 1017 -1249 1074 -1248
rect 117 -1251 213 -1250
rect 233 -1251 503 -1250
rect 548 -1251 1025 -1250
rect 1052 -1251 1098 -1250
rect 128 -1253 199 -1252
rect 205 -1253 255 -1252
rect 264 -1253 353 -1252
rect 373 -1253 556 -1252
rect 618 -1253 640 -1252
rect 656 -1253 962 -1252
rect 184 -1255 262 -1254
rect 289 -1255 297 -1254
rect 324 -1255 423 -1254
rect 478 -1255 605 -1254
rect 639 -1255 668 -1254
rect 677 -1255 731 -1254
rect 796 -1255 948 -1254
rect 961 -1255 1088 -1254
rect 184 -1257 227 -1256
rect 233 -1257 311 -1256
rect 341 -1257 584 -1256
rect 604 -1257 647 -1256
rect 656 -1257 738 -1256
rect 807 -1257 878 -1256
rect 1087 -1257 1123 -1256
rect 156 -1259 227 -1258
rect 240 -1259 447 -1258
rect 506 -1259 556 -1258
rect 572 -1259 738 -1258
rect 821 -1259 1063 -1258
rect 152 -1261 157 -1260
rect 191 -1261 321 -1260
rect 345 -1261 381 -1260
rect 404 -1261 430 -1260
rect 506 -1261 528 -1260
rect 548 -1261 598 -1260
rect 646 -1261 675 -1260
rect 709 -1261 997 -1260
rect 198 -1263 241 -1262
rect 254 -1263 269 -1262
rect 282 -1263 346 -1262
rect 352 -1263 577 -1262
rect 583 -1263 675 -1262
rect 709 -1263 815 -1262
rect 828 -1263 913 -1262
rect 121 -1265 283 -1264
rect 296 -1265 304 -1264
rect 310 -1265 633 -1264
rect 660 -1265 671 -1264
rect 723 -1265 1067 -1264
rect 107 -1267 122 -1266
rect 268 -1267 276 -1266
rect 317 -1267 573 -1266
rect 660 -1267 682 -1266
rect 723 -1267 759 -1266
rect 814 -1267 979 -1266
rect 1066 -1267 1109 -1266
rect 79 -1269 276 -1268
rect 366 -1269 528 -1268
rect 663 -1269 794 -1268
rect 835 -1269 850 -1268
rect 877 -1269 941 -1268
rect 79 -1271 136 -1270
rect 247 -1271 318 -1270
rect 376 -1271 472 -1270
rect 667 -1271 703 -1270
rect 730 -1271 780 -1270
rect 793 -1271 899 -1270
rect 912 -1271 1046 -1270
rect 37 -1273 136 -1272
rect 247 -1273 360 -1272
rect 408 -1273 451 -1272
rect 464 -1273 899 -1272
rect 940 -1273 1039 -1272
rect 1045 -1273 1095 -1272
rect 107 -1275 171 -1274
rect 359 -1275 493 -1274
rect 670 -1275 682 -1274
rect 702 -1275 717 -1274
rect 751 -1275 759 -1274
rect 779 -1275 885 -1274
rect 142 -1277 171 -1276
rect 338 -1277 493 -1276
rect 695 -1277 717 -1276
rect 751 -1277 766 -1276
rect 849 -1277 920 -1276
rect 142 -1279 332 -1278
rect 338 -1279 367 -1278
rect 415 -1279 472 -1278
rect 695 -1279 745 -1278
rect 765 -1279 955 -1278
rect 303 -1281 332 -1280
rect 401 -1281 416 -1280
rect 429 -1281 458 -1280
rect 688 -1281 745 -1280
rect 856 -1281 1039 -1280
rect 44 -1283 402 -1282
rect 436 -1283 458 -1282
rect 688 -1283 787 -1282
rect 856 -1283 934 -1282
rect 954 -1283 983 -1282
rect 44 -1285 52 -1284
rect 436 -1285 521 -1284
rect 786 -1285 843 -1284
rect 884 -1285 1028 -1284
rect 450 -1287 486 -1286
rect 520 -1287 612 -1286
rect 842 -1287 927 -1286
rect 933 -1287 1004 -1286
rect 485 -1289 514 -1288
rect 562 -1289 612 -1288
rect 891 -1289 983 -1288
rect 1003 -1289 1011 -1288
rect 499 -1291 514 -1290
rect 800 -1291 1011 -1290
rect 422 -1293 500 -1292
rect 800 -1293 871 -1292
rect 891 -1293 990 -1292
rect 870 -1295 969 -1294
rect 989 -1295 1081 -1294
rect 926 -1297 1025 -1296
rect 1080 -1297 1130 -1296
rect 968 -1299 976 -1298
rect 9 -1310 31 -1309
rect 37 -1310 115 -1309
rect 135 -1310 370 -1309
rect 408 -1310 482 -1309
rect 499 -1310 514 -1309
rect 534 -1310 591 -1309
rect 611 -1310 626 -1309
rect 628 -1310 920 -1309
rect 922 -1310 969 -1309
rect 975 -1310 983 -1309
rect 996 -1310 1004 -1309
rect 1020 -1310 1067 -1309
rect 1097 -1310 1102 -1309
rect 16 -1312 73 -1311
rect 93 -1312 101 -1311
rect 114 -1312 202 -1311
rect 212 -1312 339 -1311
rect 380 -1312 591 -1311
rect 614 -1312 752 -1311
rect 793 -1312 1011 -1311
rect 1059 -1312 1088 -1311
rect 23 -1314 241 -1313
rect 261 -1314 349 -1313
rect 380 -1314 423 -1313
rect 429 -1314 465 -1313
rect 471 -1314 514 -1313
rect 527 -1314 752 -1313
rect 793 -1314 1032 -1313
rect 1066 -1314 1081 -1313
rect 51 -1316 248 -1315
rect 268 -1316 304 -1315
rect 310 -1316 598 -1315
rect 625 -1316 703 -1315
rect 726 -1316 1025 -1315
rect 1031 -1316 1053 -1315
rect 58 -1318 538 -1317
rect 555 -1318 570 -1317
rect 576 -1318 601 -1317
rect 653 -1318 745 -1317
rect 863 -1318 941 -1317
rect 961 -1318 1011 -1317
rect 68 -1320 307 -1319
rect 408 -1320 486 -1319
rect 492 -1320 535 -1319
rect 541 -1320 556 -1319
rect 597 -1320 605 -1319
rect 677 -1320 703 -1319
rect 709 -1320 745 -1319
rect 821 -1320 864 -1319
rect 905 -1320 969 -1319
rect 999 -1320 1046 -1319
rect 72 -1322 545 -1321
rect 569 -1322 605 -1321
rect 681 -1322 710 -1321
rect 733 -1322 766 -1321
rect 870 -1322 906 -1321
rect 912 -1322 976 -1321
rect 93 -1324 482 -1323
rect 506 -1324 633 -1323
rect 737 -1324 741 -1323
rect 758 -1324 822 -1323
rect 870 -1324 885 -1323
rect 891 -1324 913 -1323
rect 933 -1324 962 -1323
rect 100 -1326 353 -1325
rect 411 -1326 682 -1325
rect 723 -1326 759 -1325
rect 765 -1326 787 -1325
rect 877 -1326 885 -1325
rect 891 -1326 1018 -1325
rect 128 -1328 262 -1327
rect 268 -1328 297 -1327
rect 345 -1328 353 -1327
rect 422 -1328 444 -1327
rect 471 -1328 521 -1327
rect 527 -1328 584 -1327
rect 660 -1328 1018 -1327
rect 86 -1330 297 -1329
rect 345 -1330 983 -1329
rect 86 -1332 276 -1331
rect 285 -1332 486 -1331
rect 506 -1332 1004 -1331
rect 128 -1334 360 -1333
rect 366 -1334 444 -1333
rect 520 -1334 675 -1333
rect 716 -1334 787 -1333
rect 856 -1334 878 -1333
rect 933 -1334 948 -1333
rect 79 -1336 360 -1335
rect 366 -1336 402 -1335
rect 429 -1336 451 -1335
rect 572 -1336 675 -1335
rect 688 -1336 717 -1335
rect 723 -1336 850 -1335
rect 856 -1336 1039 -1335
rect 79 -1338 185 -1337
rect 191 -1338 206 -1337
rect 212 -1338 279 -1337
rect 415 -1338 451 -1337
rect 572 -1338 731 -1337
rect 737 -1338 773 -1337
rect 835 -1338 850 -1337
rect 926 -1338 948 -1337
rect 170 -1340 241 -1339
rect 254 -1340 304 -1339
rect 310 -1340 731 -1339
rect 740 -1340 773 -1339
rect 926 -1340 955 -1339
rect 163 -1342 171 -1341
rect 177 -1342 206 -1341
rect 254 -1342 479 -1341
rect 583 -1342 619 -1341
rect 646 -1342 689 -1341
rect 954 -1342 990 -1341
rect 107 -1344 164 -1343
rect 177 -1344 416 -1343
rect 436 -1344 465 -1343
rect 478 -1344 549 -1343
rect 618 -1344 640 -1343
rect 646 -1344 941 -1343
rect 107 -1346 136 -1345
rect 180 -1346 227 -1345
rect 275 -1346 563 -1345
rect 660 -1346 780 -1345
rect 898 -1346 990 -1345
rect 65 -1348 563 -1347
rect 779 -1348 801 -1347
rect 184 -1350 199 -1349
rect 226 -1350 234 -1349
rect 394 -1350 899 -1349
rect 194 -1352 220 -1351
rect 233 -1352 318 -1351
rect 373 -1352 395 -1351
rect 436 -1352 458 -1351
rect 467 -1352 640 -1351
rect 800 -1352 808 -1351
rect 121 -1354 220 -1353
rect 341 -1354 458 -1353
rect 548 -1354 797 -1353
rect 807 -1354 815 -1353
rect 121 -1356 150 -1355
rect 198 -1356 325 -1355
rect 373 -1356 542 -1355
rect 814 -1356 829 -1355
rect 142 -1358 318 -1357
rect 439 -1358 577 -1357
rect 828 -1358 843 -1357
rect 142 -1360 836 -1359
rect 149 -1362 157 -1361
rect 282 -1362 325 -1361
rect 635 -1362 843 -1361
rect 156 -1364 388 -1363
rect 331 -1366 388 -1365
rect 289 -1368 332 -1367
rect 289 -1370 405 -1369
rect 2 -1381 6 -1380
rect 9 -1381 115 -1380
rect 142 -1381 241 -1380
rect 250 -1381 269 -1380
rect 369 -1381 675 -1380
rect 702 -1381 731 -1380
rect 996 -1381 1060 -1380
rect 30 -1383 34 -1382
rect 72 -1383 276 -1382
rect 369 -1383 521 -1382
rect 530 -1383 787 -1382
rect 947 -1383 997 -1382
rect 1003 -1383 1025 -1382
rect 1031 -1383 1039 -1382
rect 1045 -1383 1067 -1382
rect 30 -1385 45 -1384
rect 72 -1385 202 -1384
rect 208 -1385 591 -1384
rect 618 -1385 626 -1384
rect 632 -1385 675 -1384
rect 681 -1385 948 -1384
rect 975 -1385 1004 -1384
rect 1010 -1385 1032 -1384
rect 1055 -1385 1067 -1384
rect 33 -1387 45 -1386
rect 79 -1387 269 -1386
rect 380 -1387 437 -1386
rect 443 -1387 479 -1386
rect 488 -1387 507 -1386
rect 509 -1387 563 -1386
rect 646 -1387 759 -1386
rect 786 -1387 815 -1386
rect 940 -1387 976 -1386
rect 982 -1387 1011 -1386
rect 79 -1389 122 -1388
rect 128 -1389 437 -1388
rect 457 -1389 493 -1388
rect 499 -1389 545 -1388
rect 555 -1389 619 -1388
rect 653 -1389 990 -1388
rect 86 -1391 475 -1390
rect 513 -1391 563 -1390
rect 569 -1391 941 -1390
rect 961 -1391 990 -1390
rect 86 -1393 346 -1392
rect 366 -1393 654 -1392
rect 660 -1393 794 -1392
rect 912 -1393 962 -1392
rect 100 -1395 108 -1394
rect 114 -1395 157 -1394
rect 177 -1395 192 -1394
rect 198 -1395 248 -1394
rect 261 -1395 286 -1394
rect 289 -1395 983 -1394
rect 93 -1397 290 -1396
rect 380 -1397 402 -1396
rect 408 -1397 493 -1396
rect 534 -1397 591 -1396
rect 604 -1397 647 -1396
rect 667 -1397 682 -1396
rect 702 -1397 773 -1396
rect 793 -1397 815 -1396
rect 912 -1397 927 -1396
rect 16 -1399 94 -1398
rect 121 -1399 524 -1398
rect 537 -1399 822 -1398
rect 842 -1399 927 -1398
rect 128 -1401 899 -1400
rect 142 -1403 171 -1402
rect 212 -1403 402 -1402
rect 408 -1403 657 -1402
rect 667 -1403 752 -1402
rect 772 -1403 801 -1402
rect 821 -1403 920 -1402
rect 58 -1405 171 -1404
rect 219 -1405 262 -1404
rect 345 -1405 535 -1404
rect 541 -1405 969 -1404
rect 156 -1407 549 -1406
rect 569 -1407 724 -1406
rect 726 -1407 934 -1406
rect 135 -1409 549 -1408
rect 663 -1409 969 -1408
rect 205 -1411 220 -1410
rect 226 -1411 377 -1410
rect 415 -1411 444 -1410
rect 450 -1411 500 -1410
rect 541 -1411 745 -1410
rect 751 -1411 766 -1410
rect 828 -1411 843 -1410
rect 891 -1411 899 -1410
rect 905 -1411 920 -1410
rect 107 -1413 206 -1412
rect 226 -1413 255 -1412
rect 366 -1413 934 -1412
rect 233 -1415 1053 -1414
rect 51 -1417 234 -1416
rect 240 -1417 339 -1416
rect 415 -1417 423 -1416
rect 439 -1417 556 -1416
rect 597 -1417 745 -1416
rect 796 -1417 906 -1416
rect 51 -1419 388 -1418
rect 450 -1419 808 -1418
rect 828 -1419 885 -1418
rect 58 -1421 423 -1420
rect 471 -1421 514 -1420
rect 520 -1421 598 -1420
rect 695 -1421 724 -1420
rect 779 -1421 808 -1420
rect 877 -1421 885 -1420
rect 247 -1423 304 -1422
rect 310 -1423 339 -1422
rect 387 -1423 528 -1422
rect 688 -1423 696 -1422
rect 709 -1423 801 -1422
rect 870 -1423 878 -1422
rect 254 -1425 486 -1424
rect 527 -1425 836 -1424
rect 863 -1425 871 -1424
rect 138 -1427 864 -1426
rect 303 -1429 318 -1428
rect 348 -1429 836 -1428
rect 310 -1431 332 -1430
rect 464 -1431 486 -1430
rect 628 -1431 710 -1430
rect 716 -1431 759 -1430
rect 779 -1431 857 -1430
rect 331 -1433 353 -1432
rect 359 -1433 465 -1432
rect 576 -1433 857 -1432
rect 23 -1435 353 -1434
rect 460 -1435 717 -1434
rect 23 -1437 164 -1436
rect 324 -1437 360 -1436
rect 576 -1437 584 -1436
rect 639 -1437 689 -1436
rect 163 -1439 185 -1438
rect 296 -1439 325 -1438
rect 583 -1439 1049 -1438
rect 37 -1441 185 -1440
rect 296 -1441 374 -1440
rect 639 -1441 1018 -1440
rect 373 -1443 892 -1442
rect 954 -1443 1018 -1442
rect 495 -1445 955 -1444
rect 2 -1456 38 -1455
rect 68 -1456 395 -1455
rect 422 -1456 815 -1455
rect 824 -1456 1025 -1455
rect 1045 -1456 1060 -1455
rect 9 -1458 129 -1457
rect 142 -1458 286 -1457
rect 310 -1458 318 -1457
rect 348 -1458 444 -1457
rect 457 -1458 983 -1457
rect 999 -1458 1039 -1457
rect 1048 -1458 1053 -1457
rect 1059 -1458 1067 -1457
rect 19 -1460 59 -1459
rect 72 -1460 139 -1459
rect 142 -1460 178 -1459
rect 184 -1460 311 -1459
rect 352 -1460 461 -1459
rect 506 -1460 538 -1459
rect 593 -1460 846 -1459
rect 982 -1460 1032 -1459
rect 23 -1462 353 -1461
rect 387 -1462 475 -1461
rect 509 -1462 619 -1461
rect 625 -1462 629 -1461
rect 632 -1462 682 -1461
rect 684 -1462 934 -1461
rect 23 -1464 426 -1463
rect 436 -1464 969 -1463
rect 30 -1466 41 -1465
rect 72 -1466 563 -1465
rect 604 -1466 612 -1465
rect 625 -1466 717 -1465
rect 744 -1466 748 -1465
rect 765 -1466 864 -1465
rect 37 -1468 45 -1467
rect 93 -1468 423 -1467
rect 436 -1468 465 -1467
rect 520 -1468 759 -1467
rect 765 -1468 871 -1467
rect 44 -1470 409 -1469
rect 443 -1470 570 -1469
rect 607 -1470 948 -1469
rect 58 -1472 409 -1471
rect 450 -1472 538 -1471
rect 611 -1472 675 -1471
rect 681 -1472 927 -1471
rect 93 -1474 178 -1473
rect 191 -1474 479 -1473
rect 520 -1474 941 -1473
rect 96 -1476 759 -1475
rect 768 -1476 829 -1475
rect 856 -1476 871 -1475
rect 926 -1476 976 -1475
rect 128 -1478 304 -1477
rect 345 -1478 451 -1477
rect 464 -1478 514 -1477
rect 534 -1478 549 -1477
rect 635 -1478 661 -1477
rect 667 -1478 675 -1477
rect 709 -1478 948 -1477
rect 975 -1478 997 -1477
rect 163 -1480 185 -1479
rect 191 -1480 241 -1479
rect 247 -1480 377 -1479
rect 387 -1480 654 -1479
rect 660 -1480 668 -1479
rect 709 -1480 738 -1479
rect 744 -1480 780 -1479
rect 793 -1480 962 -1479
rect 163 -1482 199 -1481
rect 215 -1482 570 -1481
rect 639 -1482 703 -1481
rect 772 -1482 780 -1481
rect 793 -1482 843 -1481
rect 856 -1482 899 -1481
rect 170 -1484 206 -1483
rect 226 -1484 248 -1483
rect 268 -1484 276 -1483
rect 282 -1484 325 -1483
rect 373 -1484 941 -1483
rect 107 -1486 227 -1485
rect 233 -1486 325 -1485
rect 373 -1486 489 -1485
rect 544 -1486 962 -1485
rect 107 -1488 528 -1487
rect 548 -1488 577 -1487
rect 639 -1488 696 -1487
rect 702 -1488 727 -1487
rect 772 -1488 808 -1487
rect 814 -1488 885 -1487
rect 898 -1488 920 -1487
rect 68 -1490 885 -1489
rect 114 -1492 269 -1491
rect 275 -1492 360 -1491
rect 394 -1492 556 -1491
rect 642 -1492 864 -1491
rect 79 -1494 115 -1493
rect 121 -1494 171 -1493
rect 194 -1494 213 -1493
rect 233 -1494 332 -1493
rect 359 -1494 402 -1493
rect 478 -1494 598 -1493
rect 653 -1494 689 -1493
rect 695 -1494 741 -1493
rect 796 -1494 829 -1493
rect 842 -1494 1018 -1493
rect 51 -1496 122 -1495
rect 240 -1496 524 -1495
rect 541 -1496 577 -1495
rect 590 -1496 598 -1495
rect 807 -1496 878 -1495
rect 989 -1496 1018 -1495
rect 51 -1498 255 -1497
rect 296 -1498 402 -1497
rect 492 -1498 920 -1497
rect 79 -1500 157 -1499
rect 254 -1500 584 -1499
rect 590 -1500 836 -1499
rect 877 -1500 1004 -1499
rect 86 -1502 157 -1501
rect 278 -1502 493 -1501
rect 506 -1502 836 -1501
rect 905 -1502 990 -1501
rect 86 -1504 136 -1503
rect 296 -1504 458 -1503
rect 516 -1504 689 -1503
rect 747 -1504 1004 -1503
rect 16 -1506 136 -1505
rect 303 -1506 381 -1505
rect 541 -1506 934 -1505
rect 331 -1508 489 -1507
rect 555 -1508 566 -1507
rect 583 -1508 647 -1507
rect 821 -1508 997 -1507
rect 338 -1510 381 -1509
rect 646 -1510 731 -1509
rect 905 -1510 913 -1509
rect 338 -1512 367 -1511
rect 499 -1512 731 -1511
rect 912 -1512 955 -1511
rect 198 -1514 500 -1513
rect 954 -1514 1011 -1513
rect 366 -1516 724 -1515
rect 800 -1516 1011 -1515
rect 723 -1518 969 -1517
rect 800 -1520 850 -1519
rect 849 -1522 892 -1521
rect 471 -1524 892 -1523
rect 289 -1526 472 -1525
rect 30 -1528 290 -1527
rect 23 -1539 136 -1538
rect 152 -1539 962 -1538
rect 1017 -1539 1025 -1538
rect 1038 -1539 1046 -1538
rect 2 -1541 24 -1540
rect 30 -1541 426 -1540
rect 488 -1541 738 -1540
rect 740 -1541 983 -1540
rect 30 -1543 304 -1542
rect 306 -1543 507 -1542
rect 520 -1543 920 -1542
rect 961 -1543 997 -1542
rect 68 -1545 87 -1544
rect 93 -1545 416 -1544
rect 527 -1545 549 -1544
rect 558 -1545 976 -1544
rect 68 -1547 759 -1546
rect 842 -1547 885 -1546
rect 86 -1549 101 -1548
rect 135 -1549 262 -1548
rect 289 -1549 668 -1548
rect 723 -1549 815 -1548
rect 877 -1549 920 -1548
rect 100 -1551 227 -1550
rect 247 -1551 262 -1550
rect 296 -1551 360 -1550
rect 366 -1551 629 -1550
rect 663 -1551 829 -1550
rect 884 -1551 1004 -1550
rect 128 -1553 290 -1552
rect 373 -1553 486 -1552
rect 499 -1553 549 -1552
rect 565 -1553 948 -1552
rect 72 -1555 500 -1554
rect 534 -1555 556 -1554
rect 583 -1555 668 -1554
rect 684 -1555 878 -1554
rect 947 -1555 1011 -1554
rect 16 -1557 73 -1556
rect 121 -1557 129 -1556
rect 156 -1557 314 -1556
rect 359 -1557 566 -1556
rect 583 -1557 696 -1556
rect 726 -1557 899 -1556
rect 121 -1559 276 -1558
rect 366 -1559 556 -1558
rect 590 -1559 829 -1558
rect 898 -1559 934 -1558
rect 44 -1561 276 -1560
rect 373 -1561 538 -1560
rect 541 -1561 612 -1560
rect 618 -1561 654 -1560
rect 737 -1561 822 -1560
rect 44 -1563 143 -1562
rect 156 -1563 339 -1562
rect 355 -1563 654 -1562
rect 758 -1563 801 -1562
rect 814 -1563 864 -1562
rect 107 -1565 339 -1564
rect 380 -1565 416 -1564
rect 590 -1565 640 -1564
rect 800 -1565 808 -1564
rect 821 -1565 850 -1564
rect 863 -1565 913 -1564
rect 142 -1567 150 -1566
rect 170 -1567 696 -1566
rect 807 -1567 871 -1566
rect 912 -1567 990 -1566
rect 177 -1569 381 -1568
rect 387 -1569 514 -1568
rect 576 -1569 640 -1568
rect 660 -1569 850 -1568
rect 870 -1569 927 -1568
rect 177 -1571 192 -1570
rect 201 -1571 311 -1570
rect 401 -1571 465 -1570
rect 478 -1571 514 -1570
rect 562 -1571 927 -1570
rect 191 -1573 206 -1572
rect 212 -1573 297 -1572
rect 394 -1573 479 -1572
rect 576 -1573 633 -1572
rect 660 -1573 689 -1572
rect 205 -1575 234 -1574
rect 240 -1575 356 -1574
rect 401 -1575 430 -1574
rect 569 -1575 633 -1574
rect 688 -1575 710 -1574
rect 163 -1577 234 -1576
rect 240 -1577 423 -1576
rect 429 -1577 458 -1576
rect 604 -1577 626 -1576
rect 709 -1577 745 -1576
rect 58 -1579 164 -1578
rect 212 -1579 220 -1578
rect 247 -1579 283 -1578
rect 345 -1579 395 -1578
rect 408 -1579 703 -1578
rect 744 -1579 780 -1578
rect 58 -1581 174 -1580
rect 408 -1581 444 -1580
rect 450 -1581 458 -1580
rect 597 -1581 780 -1580
rect 51 -1583 451 -1582
rect 618 -1583 675 -1582
rect 702 -1583 941 -1582
rect 51 -1585 573 -1584
rect 716 -1585 941 -1584
rect 114 -1587 220 -1586
rect 387 -1587 598 -1586
rect 716 -1587 752 -1586
rect 107 -1589 115 -1588
rect 117 -1589 283 -1588
rect 411 -1589 731 -1588
rect 751 -1589 787 -1588
rect 443 -1591 531 -1590
rect 730 -1591 773 -1590
rect 786 -1591 857 -1590
rect 492 -1593 675 -1592
rect 765 -1593 773 -1592
rect 856 -1593 937 -1592
rect 331 -1595 493 -1594
rect 765 -1595 794 -1594
rect 317 -1597 332 -1596
rect 793 -1597 836 -1596
rect 268 -1599 318 -1598
rect 835 -1599 892 -1598
rect 254 -1601 269 -1600
rect 891 -1601 955 -1600
rect 254 -1603 510 -1602
rect 905 -1603 955 -1602
rect 905 -1605 969 -1604
rect 30 -1616 356 -1615
rect 366 -1616 528 -1615
rect 530 -1616 780 -1615
rect 926 -1616 937 -1615
rect 954 -1616 969 -1615
rect 1038 -1616 1046 -1615
rect 58 -1618 304 -1617
rect 310 -1618 472 -1617
rect 523 -1618 668 -1617
rect 681 -1618 738 -1617
rect 775 -1618 850 -1617
rect 65 -1620 111 -1619
rect 121 -1620 307 -1619
rect 310 -1620 353 -1619
rect 366 -1620 402 -1619
rect 425 -1620 472 -1619
rect 544 -1620 794 -1619
rect 68 -1622 241 -1621
rect 257 -1622 325 -1621
rect 352 -1622 409 -1621
rect 429 -1622 517 -1621
rect 551 -1622 640 -1621
rect 646 -1622 668 -1621
rect 681 -1622 685 -1621
rect 695 -1622 920 -1621
rect 72 -1624 412 -1623
rect 562 -1624 839 -1623
rect 79 -1626 402 -1625
rect 562 -1626 703 -1625
rect 723 -1626 738 -1625
rect 751 -1626 794 -1625
rect 79 -1628 230 -1627
rect 268 -1628 423 -1627
rect 565 -1628 619 -1627
rect 688 -1628 752 -1627
rect 779 -1628 822 -1627
rect 107 -1630 514 -1629
rect 569 -1630 815 -1629
rect 93 -1632 108 -1631
rect 121 -1632 160 -1631
rect 163 -1632 241 -1631
rect 268 -1632 405 -1631
rect 513 -1632 860 -1631
rect 93 -1634 255 -1633
rect 282 -1634 524 -1633
rect 569 -1634 633 -1633
rect 688 -1634 871 -1633
rect 128 -1636 164 -1635
rect 198 -1636 346 -1635
rect 376 -1636 381 -1635
rect 387 -1636 444 -1635
rect 576 -1636 633 -1635
rect 695 -1636 804 -1635
rect 814 -1636 941 -1635
rect 114 -1638 129 -1637
rect 149 -1638 171 -1637
rect 208 -1638 423 -1637
rect 443 -1638 465 -1637
rect 478 -1638 577 -1637
rect 590 -1638 626 -1637
rect 702 -1638 766 -1637
rect 86 -1640 115 -1639
rect 152 -1640 248 -1639
rect 275 -1640 283 -1639
rect 296 -1640 433 -1639
rect 478 -1640 500 -1639
rect 590 -1640 661 -1639
rect 709 -1640 766 -1639
rect 86 -1642 206 -1641
rect 212 -1642 227 -1641
rect 247 -1642 290 -1641
rect 296 -1642 332 -1641
rect 359 -1642 381 -1641
rect 390 -1642 493 -1641
rect 499 -1642 521 -1641
rect 604 -1642 647 -1641
rect 709 -1642 745 -1641
rect 758 -1642 822 -1641
rect 44 -1644 206 -1643
rect 212 -1644 220 -1643
rect 226 -1644 234 -1643
rect 289 -1644 437 -1643
rect 485 -1644 493 -1643
rect 583 -1644 605 -1643
rect 611 -1644 654 -1643
rect 716 -1644 724 -1643
rect 730 -1644 759 -1643
rect 23 -1646 45 -1645
rect 135 -1646 234 -1645
rect 317 -1646 346 -1645
rect 373 -1646 465 -1645
rect 485 -1646 507 -1645
rect 541 -1646 584 -1645
rect 614 -1646 843 -1645
rect 135 -1648 153 -1647
rect 156 -1648 899 -1647
rect 100 -1650 157 -1649
rect 170 -1650 202 -1649
rect 306 -1650 374 -1649
rect 394 -1650 829 -1649
rect 842 -1650 878 -1649
rect 51 -1652 101 -1651
rect 177 -1652 220 -1651
rect 317 -1652 556 -1651
rect 716 -1652 836 -1651
rect 40 -1654 52 -1653
rect 184 -1654 276 -1653
rect 324 -1654 542 -1653
rect 555 -1654 675 -1653
rect 733 -1654 885 -1653
rect 184 -1656 192 -1655
rect 331 -1656 416 -1655
rect 436 -1656 458 -1655
rect 506 -1656 549 -1655
rect 744 -1656 808 -1655
rect 884 -1656 948 -1655
rect 191 -1658 335 -1657
rect 338 -1658 360 -1657
rect 394 -1658 451 -1657
rect 786 -1658 829 -1657
rect 303 -1660 458 -1659
rect 772 -1660 787 -1659
rect 800 -1660 836 -1659
rect 313 -1662 416 -1661
rect 429 -1662 451 -1661
rect 800 -1662 962 -1661
rect 807 -1664 864 -1663
rect 863 -1666 892 -1665
rect 891 -1668 906 -1667
rect 905 -1670 913 -1669
rect 44 -1681 52 -1680
rect 65 -1681 104 -1680
rect 107 -1681 255 -1680
rect 264 -1681 325 -1680
rect 383 -1681 388 -1680
rect 408 -1681 500 -1680
rect 513 -1681 524 -1680
rect 541 -1681 570 -1680
rect 593 -1681 598 -1680
rect 611 -1681 619 -1680
rect 625 -1681 640 -1680
rect 646 -1681 689 -1680
rect 723 -1681 731 -1680
rect 758 -1681 773 -1680
rect 779 -1681 853 -1680
rect 856 -1681 864 -1680
rect 898 -1681 906 -1680
rect 47 -1683 59 -1682
rect 86 -1683 307 -1682
rect 310 -1683 377 -1682
rect 380 -1683 388 -1682
rect 422 -1683 426 -1682
rect 429 -1683 444 -1682
rect 450 -1683 475 -1682
rect 520 -1683 591 -1682
rect 604 -1683 612 -1682
rect 632 -1683 647 -1682
rect 653 -1683 696 -1682
rect 709 -1683 724 -1682
rect 737 -1683 759 -1682
rect 782 -1683 808 -1682
rect 817 -1683 885 -1682
rect 93 -1685 202 -1684
rect 212 -1685 335 -1684
rect 373 -1685 409 -1684
rect 422 -1685 437 -1684
rect 450 -1685 486 -1684
rect 569 -1685 692 -1684
rect 709 -1685 717 -1684
rect 737 -1685 745 -1684
rect 786 -1685 850 -1684
rect 884 -1685 892 -1684
rect 75 -1687 94 -1686
rect 100 -1687 181 -1686
rect 201 -1687 227 -1686
rect 240 -1687 244 -1686
rect 282 -1687 304 -1686
rect 310 -1687 346 -1686
rect 373 -1687 465 -1686
rect 576 -1687 605 -1686
rect 667 -1687 675 -1686
rect 677 -1687 682 -1686
rect 744 -1687 752 -1686
rect 793 -1687 801 -1686
rect 807 -1687 843 -1686
rect 849 -1687 867 -1686
rect 114 -1689 150 -1688
rect 156 -1689 199 -1688
rect 219 -1689 227 -1688
rect 240 -1689 276 -1688
rect 324 -1689 342 -1688
rect 345 -1689 353 -1688
rect 401 -1689 521 -1688
rect 527 -1689 577 -1688
rect 702 -1689 752 -1688
rect 765 -1689 794 -1688
rect 821 -1689 836 -1688
rect 117 -1691 122 -1690
rect 128 -1691 181 -1690
rect 184 -1691 220 -1690
rect 247 -1691 342 -1690
rect 404 -1691 444 -1690
rect 464 -1691 535 -1690
rect 765 -1691 815 -1690
rect 821 -1691 864 -1690
rect 128 -1693 136 -1692
rect 156 -1693 178 -1692
rect 268 -1693 283 -1692
rect 415 -1693 486 -1692
rect 527 -1693 556 -1692
rect 163 -1695 209 -1694
rect 261 -1695 269 -1694
rect 275 -1695 290 -1694
rect 394 -1695 416 -1694
rect 436 -1695 479 -1694
rect 163 -1697 192 -1696
rect 289 -1697 318 -1696
rect 394 -1697 433 -1696
rect 457 -1697 535 -1696
rect 177 -1699 356 -1698
rect 457 -1699 549 -1698
rect 191 -1701 216 -1700
rect 317 -1701 332 -1700
rect 471 -1701 556 -1700
rect 296 -1703 332 -1702
rect 478 -1703 507 -1702
rect 548 -1703 563 -1702
rect 492 -1705 507 -1704
rect 562 -1705 584 -1704
rect 425 -1707 493 -1706
rect 583 -1707 591 -1706
rect 58 -1718 66 -1717
rect 93 -1718 118 -1717
rect 121 -1718 129 -1717
rect 142 -1718 153 -1717
rect 156 -1718 185 -1717
rect 212 -1718 241 -1717
rect 268 -1718 276 -1717
rect 289 -1718 402 -1717
rect 411 -1718 521 -1717
rect 562 -1718 591 -1717
rect 593 -1718 783 -1717
rect 793 -1718 797 -1717
rect 828 -1718 867 -1717
rect 103 -1720 146 -1719
rect 149 -1720 178 -1719
rect 205 -1720 213 -1719
rect 215 -1720 279 -1719
rect 299 -1720 570 -1719
rect 583 -1720 598 -1719
rect 604 -1720 654 -1719
rect 674 -1720 682 -1719
rect 702 -1720 710 -1719
rect 730 -1720 734 -1719
rect 772 -1720 787 -1719
rect 793 -1720 808 -1719
rect 821 -1720 829 -1719
rect 835 -1720 843 -1719
rect 845 -1720 857 -1719
rect 107 -1722 115 -1721
rect 142 -1722 157 -1721
rect 163 -1722 185 -1721
rect 219 -1722 262 -1721
rect 324 -1722 370 -1721
rect 380 -1722 409 -1721
rect 422 -1722 447 -1721
rect 464 -1722 500 -1721
rect 597 -1722 619 -1721
rect 639 -1722 657 -1721
rect 709 -1722 780 -1721
rect 849 -1722 857 -1721
rect 163 -1724 171 -1723
rect 226 -1724 241 -1723
rect 296 -1724 325 -1723
rect 338 -1724 346 -1723
rect 352 -1724 612 -1723
rect 730 -1724 738 -1723
rect 233 -1726 248 -1725
rect 282 -1726 297 -1725
rect 338 -1726 374 -1725
rect 422 -1726 430 -1725
rect 464 -1726 479 -1725
rect 492 -1726 521 -1725
rect 737 -1726 745 -1725
rect 226 -1728 234 -1727
rect 331 -1728 374 -1727
rect 429 -1728 458 -1727
rect 471 -1728 577 -1727
rect 744 -1728 766 -1727
rect 317 -1730 332 -1729
rect 345 -1730 360 -1729
rect 366 -1730 377 -1729
rect 457 -1730 549 -1729
rect 555 -1730 577 -1729
rect 758 -1730 766 -1729
rect 254 -1732 318 -1731
rect 352 -1732 384 -1731
rect 478 -1732 507 -1731
rect 534 -1732 549 -1731
rect 555 -1732 570 -1731
rect 751 -1732 759 -1731
rect 359 -1734 416 -1733
rect 485 -1734 493 -1733
rect 499 -1734 528 -1733
rect 366 -1736 395 -1735
rect 415 -1736 451 -1735
rect 513 -1736 535 -1735
rect 387 -1738 395 -1737
rect 436 -1738 451 -1737
rect 485 -1738 514 -1737
rect 436 -1740 444 -1739
rect 796 -1740 808 -1739
rect 44 -1751 48 -1750
rect 58 -1751 62 -1750
rect 65 -1751 73 -1750
rect 93 -1751 118 -1750
rect 121 -1751 136 -1750
rect 159 -1751 178 -1750
rect 184 -1751 213 -1750
rect 219 -1751 248 -1750
rect 282 -1751 304 -1750
rect 352 -1751 370 -1750
rect 373 -1751 402 -1750
rect 443 -1751 458 -1750
rect 464 -1751 472 -1750
rect 488 -1751 577 -1750
rect 586 -1751 591 -1750
rect 646 -1751 657 -1750
rect 716 -1751 731 -1750
rect 765 -1751 783 -1750
rect 807 -1751 815 -1750
rect 842 -1751 846 -1750
rect 968 -1751 976 -1750
rect 65 -1753 80 -1752
rect 107 -1753 122 -1752
rect 128 -1753 146 -1752
rect 163 -1753 174 -1752
rect 219 -1753 234 -1752
rect 289 -1753 311 -1752
rect 317 -1753 353 -1752
rect 366 -1753 374 -1752
rect 387 -1753 405 -1752
rect 450 -1753 465 -1752
rect 471 -1753 493 -1752
rect 499 -1753 510 -1752
rect 527 -1753 542 -1752
rect 548 -1753 556 -1752
rect 562 -1753 598 -1752
rect 709 -1753 731 -1752
rect 772 -1753 787 -1752
rect 128 -1755 132 -1754
rect 135 -1755 143 -1754
rect 233 -1755 241 -1754
rect 296 -1755 318 -1754
rect 429 -1755 451 -1754
rect 457 -1755 521 -1754
rect 530 -1755 535 -1754
rect 562 -1755 570 -1754
rect 702 -1755 710 -1754
rect 758 -1755 773 -1754
rect 779 -1755 794 -1754
rect 138 -1757 143 -1756
rect 229 -1757 241 -1756
rect 296 -1757 332 -1756
rect 429 -1757 437 -1756
rect 751 -1757 759 -1756
rect 793 -1757 801 -1756
rect 310 -1759 339 -1758
rect 737 -1759 752 -1758
rect 324 -1761 339 -1760
rect 737 -1761 745 -1760
rect 324 -1763 346 -1762
rect 345 -1765 360 -1764
rect 359 -1767 412 -1766
rect 58 -1778 66 -1777
rect 75 -1778 80 -1777
rect 93 -1778 111 -1777
rect 117 -1778 129 -1777
rect 135 -1778 153 -1777
rect 170 -1778 174 -1777
rect 191 -1778 199 -1777
rect 219 -1778 227 -1777
rect 247 -1778 262 -1777
rect 282 -1778 321 -1777
rect 331 -1778 346 -1777
rect 380 -1778 388 -1777
rect 394 -1778 412 -1777
rect 502 -1778 507 -1777
rect 520 -1778 528 -1777
rect 562 -1778 566 -1777
rect 709 -1778 717 -1777
rect 723 -1778 748 -1777
rect 751 -1778 766 -1777
rect 772 -1778 780 -1777
rect 828 -1778 839 -1777
rect 880 -1778 885 -1777
rect 72 -1780 80 -1779
rect 152 -1780 157 -1779
rect 226 -1780 234 -1779
rect 275 -1780 283 -1779
rect 289 -1780 307 -1779
rect 324 -1780 332 -1779
rect 373 -1780 381 -1779
rect 401 -1780 423 -1779
rect 730 -1780 773 -1779
rect 296 -1782 314 -1781
rect 411 -1782 458 -1781
rect 296 -1784 304 -1783
rect 306 -1784 363 -1783
rect 450 -1784 458 -1783
rect 310 -1786 325 -1785
rect 450 -1786 472 -1785
rect 464 -1788 472 -1787
rect 68 -1799 80 -1798
rect 142 -1799 150 -1798
rect 156 -1799 160 -1798
rect 184 -1799 192 -1798
rect 205 -1799 209 -1798
rect 240 -1799 248 -1798
rect 261 -1799 269 -1798
rect 324 -1799 342 -1798
rect 380 -1799 384 -1798
rect 422 -1799 430 -1798
rect 432 -1799 444 -1798
rect 457 -1799 465 -1798
rect 471 -1799 482 -1798
rect 506 -1799 514 -1798
rect 516 -1799 521 -1798
rect 737 -1799 752 -1798
rect 754 -1799 766 -1798
rect 793 -1799 797 -1798
rect 898 -1799 906 -1798
rect 1024 -1799 1028 -1798
rect 331 -1801 346 -1800
rect 415 -1801 423 -1800
rect 439 -1801 451 -1800
rect 471 -1801 479 -1800
rect 744 -1801 759 -1800
rect 331 -1803 339 -1802
rect 187 -1814 192 -1813
rect 222 -1814 227 -1813
rect 264 -1814 269 -1813
rect 296 -1814 307 -1813
rect 324 -1814 332 -1813
rect 352 -1814 360 -1813
rect 376 -1814 388 -1813
rect 422 -1814 430 -1813
rect 747 -1814 752 -1813
rect 901 -1814 906 -1813
<< m2contact >>
rect 177 0 178 1
rect 198 0 199 1
rect 212 0 213 1
rect 219 0 220 1
rect 236 0 237 1
rect 240 0 241 1
rect 254 0 255 1
rect 261 0 262 1
rect 285 0 286 1
rect 289 0 290 1
rect 303 0 304 1
rect 310 0 311 1
rect 338 0 339 1
rect 348 0 349 1
rect 352 0 353 1
rect 359 0 360 1
rect 366 0 367 1
rect 408 0 409 1
rect 467 0 468 1
rect 471 0 472 1
rect 478 0 479 1
rect 485 0 486 1
rect 534 0 535 1
rect 541 0 542 1
rect 576 0 577 1
rect 583 0 584 1
rect 604 0 605 1
rect 611 0 612 1
rect 730 0 731 1
rect 740 0 741 1
rect 184 -2 185 -1
rect 194 -2 195 -1
rect 114 -13 115 -12
rect 121 -13 122 -12
rect 156 -13 157 -12
rect 163 -13 164 -12
rect 170 -13 171 -12
rect 177 -13 178 -12
rect 219 -13 220 -12
rect 226 -13 227 -12
rect 240 -13 241 -12
rect 254 -13 255 -12
rect 278 -13 279 -12
rect 282 -13 283 -12
rect 303 -13 304 -12
rect 310 -13 311 -12
rect 345 -13 346 -12
rect 366 -13 367 -12
rect 408 -13 409 -12
rect 443 -13 444 -12
rect 450 -13 451 -12
rect 460 -13 461 -12
rect 474 -13 475 -12
rect 478 -13 479 -12
rect 485 -13 486 -12
rect 492 -13 493 -12
rect 527 -13 528 -12
rect 558 -13 559 -12
rect 604 -13 605 -12
rect 611 -13 612 -12
rect 618 -13 619 -12
rect 621 -13 622 -12
rect 688 -13 689 -12
rect 698 -13 699 -12
rect 215 -15 216 -14
rect 219 -15 220 -14
rect 247 -15 248 -14
rect 261 -15 262 -14
rect 289 -15 290 -14
rect 303 -15 304 -14
rect 352 -15 353 -14
rect 359 -15 360 -14
rect 366 -15 367 -14
rect 373 -15 374 -14
rect 415 -15 416 -14
rect 422 -15 423 -14
rect 425 -15 426 -14
rect 429 -15 430 -14
rect 457 -15 458 -14
rect 467 -15 468 -14
rect 471 -15 472 -14
rect 485 -15 486 -14
rect 555 -15 556 -14
rect 604 -15 605 -14
rect 240 -17 241 -16
rect 261 -17 262 -16
rect 278 -17 279 -16
rect 289 -17 290 -16
rect 338 -17 339 -16
rect 352 -17 353 -16
rect 334 -19 335 -18
rect 338 -19 339 -18
rect 58 -30 59 -29
rect 61 -30 62 -29
rect 114 -30 115 -29
rect 124 -30 125 -29
rect 142 -30 143 -29
rect 170 -30 171 -29
rect 184 -30 185 -29
rect 198 -30 199 -29
rect 212 -30 213 -29
rect 219 -30 220 -29
rect 226 -30 227 -29
rect 261 -30 262 -29
rect 268 -30 269 -29
rect 296 -30 297 -29
rect 317 -30 318 -29
rect 324 -30 325 -29
rect 334 -30 335 -29
rect 345 -30 346 -29
rect 352 -30 353 -29
rect 373 -30 374 -29
rect 387 -30 388 -29
rect 401 -30 402 -29
rect 408 -30 409 -29
rect 411 -30 412 -29
rect 415 -30 416 -29
rect 425 -30 426 -29
rect 429 -30 430 -29
rect 432 -30 433 -29
rect 443 -30 444 -29
rect 471 -30 472 -29
rect 492 -30 493 -29
rect 499 -30 500 -29
rect 513 -30 514 -29
rect 537 -30 538 -29
rect 541 -30 542 -29
rect 548 -30 549 -29
rect 576 -30 577 -29
rect 579 -30 580 -29
rect 583 -30 584 -29
rect 597 -30 598 -29
rect 604 -30 605 -29
rect 632 -30 633 -29
rect 646 -30 647 -29
rect 660 -30 661 -29
rect 709 -30 710 -29
rect 786 -30 787 -29
rect 807 -30 808 -29
rect 814 -30 815 -29
rect 121 -32 122 -31
rect 135 -32 136 -31
rect 152 -32 153 -31
rect 156 -32 157 -31
rect 163 -32 164 -31
rect 173 -32 174 -31
rect 177 -32 178 -31
rect 226 -32 227 -31
rect 233 -32 234 -31
rect 240 -32 241 -31
rect 254 -32 255 -31
rect 296 -32 297 -31
rect 345 -32 346 -31
rect 366 -32 367 -31
rect 429 -32 430 -31
rect 436 -32 437 -31
rect 527 -32 528 -31
rect 555 -32 556 -31
rect 572 -32 573 -31
rect 583 -32 584 -31
rect 604 -32 605 -31
rect 611 -32 612 -31
rect 625 -32 626 -31
rect 712 -32 713 -31
rect 163 -34 164 -33
rect 170 -34 171 -33
rect 180 -34 181 -33
rect 184 -34 185 -33
rect 240 -34 241 -33
rect 282 -34 283 -33
rect 352 -34 353 -33
rect 397 -34 398 -33
rect 432 -34 433 -33
rect 436 -34 437 -33
rect 541 -34 542 -33
rect 562 -34 563 -33
rect 611 -34 612 -33
rect 618 -34 619 -33
rect 247 -36 248 -35
rect 254 -36 255 -35
rect 257 -36 258 -35
rect 275 -36 276 -35
rect 282 -36 283 -35
rect 310 -36 311 -35
rect 359 -36 360 -35
rect 366 -36 367 -35
rect 247 -38 248 -37
rect 271 -38 272 -37
rect 303 -38 304 -37
rect 310 -38 311 -37
rect 338 -38 339 -37
rect 359 -38 360 -37
rect 303 -40 304 -39
rect 331 -40 332 -39
rect 317 -42 318 -41
rect 338 -42 339 -41
rect 93 -53 94 -52
rect 103 -53 104 -52
rect 107 -53 108 -52
rect 149 -53 150 -52
rect 170 -53 171 -52
rect 184 -53 185 -52
rect 226 -53 227 -52
rect 278 -53 279 -52
rect 310 -53 311 -52
rect 331 -53 332 -52
rect 338 -53 339 -52
rect 401 -53 402 -52
rect 415 -53 416 -52
rect 460 -53 461 -52
rect 478 -53 479 -52
rect 506 -53 507 -52
rect 513 -53 514 -52
rect 520 -53 521 -52
rect 534 -53 535 -52
rect 618 -53 619 -52
rect 660 -53 661 -52
rect 674 -53 675 -52
rect 688 -53 689 -52
rect 702 -53 703 -52
rect 793 -53 794 -52
rect 807 -53 808 -52
rect 1087 -53 1088 -52
rect 1097 -53 1098 -52
rect 110 -55 111 -54
rect 205 -55 206 -54
rect 229 -55 230 -54
rect 296 -55 297 -54
rect 373 -55 374 -54
rect 387 -55 388 -54
rect 429 -55 430 -54
rect 443 -55 444 -54
rect 485 -55 486 -54
rect 513 -55 514 -54
rect 541 -55 542 -54
rect 583 -55 584 -54
rect 653 -55 654 -54
rect 660 -55 661 -54
rect 786 -55 787 -54
rect 807 -55 808 -54
rect 121 -57 122 -56
rect 135 -57 136 -56
rect 170 -57 171 -56
rect 191 -57 192 -56
rect 233 -57 234 -56
rect 254 -57 255 -56
rect 289 -57 290 -56
rect 310 -57 311 -56
rect 373 -57 374 -56
rect 467 -57 468 -56
rect 474 -57 475 -56
rect 485 -57 486 -56
rect 499 -57 500 -56
rect 534 -57 535 -56
rect 555 -57 556 -56
rect 646 -57 647 -56
rect 128 -59 129 -58
rect 177 -59 178 -58
rect 184 -59 185 -58
rect 275 -59 276 -58
rect 289 -59 290 -58
rect 299 -59 300 -58
rect 380 -59 381 -58
rect 401 -59 402 -58
rect 422 -59 423 -58
rect 443 -59 444 -58
rect 471 -59 472 -58
rect 499 -59 500 -58
rect 527 -59 528 -58
rect 555 -59 556 -58
rect 569 -59 570 -58
rect 625 -59 626 -58
rect 632 -59 633 -58
rect 653 -59 654 -58
rect 135 -61 136 -60
rect 156 -61 157 -60
rect 191 -61 192 -60
rect 208 -61 209 -60
rect 233 -61 234 -60
rect 261 -61 262 -60
rect 380 -61 381 -60
rect 408 -61 409 -60
rect 422 -61 423 -60
rect 450 -61 451 -60
rect 495 -61 496 -60
rect 625 -61 626 -60
rect 632 -61 633 -60
rect 639 -61 640 -60
rect 156 -63 157 -62
rect 198 -63 199 -62
rect 208 -63 209 -62
rect 212 -63 213 -62
rect 247 -63 248 -62
rect 261 -63 262 -62
rect 408 -63 409 -62
rect 457 -63 458 -62
rect 576 -63 577 -62
rect 583 -63 584 -62
rect 198 -65 199 -64
rect 282 -65 283 -64
rect 429 -65 430 -64
rect 446 -65 447 -64
rect 576 -65 577 -64
rect 604 -65 605 -64
rect 212 -67 213 -66
rect 303 -67 304 -66
rect 436 -67 437 -66
rect 450 -67 451 -66
rect 597 -67 598 -66
rect 604 -67 605 -66
rect 222 -69 223 -68
rect 247 -69 248 -68
rect 268 -69 269 -68
rect 303 -69 304 -68
rect 439 -69 440 -68
rect 478 -69 479 -68
rect 590 -69 591 -68
rect 597 -69 598 -68
rect 268 -71 269 -70
rect 359 -71 360 -70
rect 562 -71 563 -70
rect 590 -71 591 -70
rect 282 -73 283 -72
rect 317 -73 318 -72
rect 548 -73 549 -72
rect 562 -73 563 -72
rect 317 -75 318 -74
rect 352 -75 353 -74
rect 446 -75 447 -74
rect 548 -75 549 -74
rect 324 -77 325 -76
rect 352 -77 353 -76
rect 324 -79 325 -78
rect 394 -79 395 -78
rect 131 -81 132 -80
rect 394 -81 395 -80
rect 30 -92 31 -91
rect 44 -92 45 -91
rect 51 -92 52 -91
rect 65 -92 66 -91
rect 89 -92 90 -91
rect 93 -92 94 -91
rect 100 -92 101 -91
rect 156 -92 157 -91
rect 219 -92 220 -91
rect 268 -92 269 -91
rect 275 -92 276 -91
rect 289 -92 290 -91
rect 299 -92 300 -91
rect 352 -92 353 -91
rect 366 -92 367 -91
rect 394 -92 395 -91
rect 397 -92 398 -91
rect 411 -92 412 -91
rect 429 -92 430 -91
rect 495 -92 496 -91
rect 527 -92 528 -91
rect 555 -92 556 -91
rect 597 -92 598 -91
rect 632 -92 633 -91
rect 646 -92 647 -91
rect 688 -92 689 -91
rect 730 -92 731 -91
rect 737 -92 738 -91
rect 758 -92 759 -91
rect 779 -92 780 -91
rect 800 -92 801 -91
rect 807 -92 808 -91
rect 898 -92 899 -91
rect 905 -92 906 -91
rect 975 -92 976 -91
rect 978 -92 979 -91
rect 54 -94 55 -93
rect 65 -94 66 -93
rect 93 -94 94 -93
rect 142 -94 143 -93
rect 149 -94 150 -93
rect 187 -94 188 -93
rect 261 -94 262 -93
rect 268 -94 269 -93
rect 282 -94 283 -93
rect 289 -94 290 -93
rect 303 -94 304 -93
rect 306 -94 307 -93
rect 338 -94 339 -93
rect 366 -94 367 -93
rect 387 -94 388 -93
rect 390 -94 391 -93
rect 401 -94 402 -93
rect 429 -94 430 -93
rect 450 -94 451 -93
rect 471 -94 472 -93
rect 478 -94 479 -93
rect 492 -94 493 -93
rect 541 -94 542 -93
rect 597 -94 598 -93
rect 604 -94 605 -93
rect 667 -94 668 -93
rect 674 -94 675 -93
rect 716 -94 717 -93
rect 765 -94 766 -93
rect 793 -94 794 -93
rect 107 -96 108 -95
rect 415 -96 416 -95
rect 450 -96 451 -95
rect 639 -96 640 -95
rect 681 -96 682 -95
rect 723 -96 724 -95
rect 121 -98 122 -97
rect 184 -98 185 -97
rect 240 -98 241 -97
rect 261 -98 262 -97
rect 282 -98 283 -97
rect 317 -98 318 -97
rect 327 -98 328 -97
rect 338 -98 339 -97
rect 373 -98 374 -97
rect 415 -98 416 -97
rect 457 -98 458 -97
rect 485 -98 486 -97
rect 534 -98 535 -97
rect 639 -98 640 -97
rect 702 -98 703 -97
rect 730 -98 731 -97
rect 124 -100 125 -99
rect 177 -100 178 -99
rect 240 -100 241 -99
rect 247 -100 248 -99
rect 303 -100 304 -99
rect 310 -100 311 -99
rect 317 -100 318 -99
rect 324 -100 325 -99
rect 380 -100 381 -99
rect 401 -100 402 -99
rect 408 -100 409 -99
rect 443 -100 444 -99
rect 467 -100 468 -99
rect 485 -100 486 -99
rect 499 -100 500 -99
rect 534 -100 535 -99
rect 541 -100 542 -99
rect 569 -100 570 -99
rect 590 -100 591 -99
rect 646 -100 647 -99
rect 660 -100 661 -99
rect 702 -100 703 -99
rect 128 -102 129 -101
rect 180 -102 181 -101
rect 324 -102 325 -101
rect 436 -102 437 -101
rect 520 -102 521 -101
rect 569 -102 570 -101
rect 593 -102 594 -101
rect 681 -102 682 -101
rect 128 -104 129 -103
rect 345 -104 346 -103
rect 355 -104 356 -103
rect 520 -104 521 -103
rect 562 -104 563 -103
rect 604 -104 605 -103
rect 611 -104 612 -103
rect 660 -104 661 -103
rect 135 -106 136 -105
rect 180 -106 181 -105
rect 212 -106 213 -105
rect 345 -106 346 -105
rect 362 -106 363 -105
rect 499 -106 500 -105
rect 506 -106 507 -105
rect 562 -106 563 -105
rect 618 -106 619 -105
rect 674 -106 675 -105
rect 142 -108 143 -107
rect 198 -108 199 -107
rect 212 -108 213 -107
rect 233 -108 234 -107
rect 373 -108 374 -107
rect 436 -108 437 -107
rect 548 -108 549 -107
rect 611 -108 612 -107
rect 625 -108 626 -107
rect 695 -108 696 -107
rect 149 -110 150 -109
rect 205 -110 206 -109
rect 233 -110 234 -109
rect 254 -110 255 -109
rect 387 -110 388 -109
rect 422 -110 423 -109
rect 513 -110 514 -109
rect 625 -110 626 -109
rect 156 -112 157 -111
rect 163 -112 164 -111
rect 198 -112 199 -111
rect 229 -112 230 -111
rect 390 -112 391 -111
rect 422 -112 423 -111
rect 576 -112 577 -111
rect 618 -112 619 -111
rect 163 -114 164 -113
rect 170 -114 171 -113
rect 205 -114 206 -113
rect 359 -114 360 -113
rect 408 -114 409 -113
rect 513 -114 514 -113
rect 576 -114 577 -113
rect 653 -114 654 -113
rect 170 -116 171 -115
rect 191 -116 192 -115
rect 229 -116 230 -115
rect 254 -116 255 -115
rect 299 -116 300 -115
rect 359 -116 360 -115
rect 191 -118 192 -117
rect 222 -118 223 -117
rect 23 -129 24 -128
rect 44 -129 45 -128
rect 47 -129 48 -128
rect 65 -129 66 -128
rect 79 -129 80 -128
rect 86 -129 87 -128
rect 121 -129 122 -128
rect 184 -129 185 -128
rect 219 -129 220 -128
rect 324 -129 325 -128
rect 338 -129 339 -128
rect 408 -129 409 -128
rect 457 -129 458 -128
rect 464 -129 465 -128
rect 495 -129 496 -128
rect 506 -129 507 -128
rect 541 -129 542 -128
rect 593 -129 594 -128
rect 656 -129 657 -128
rect 758 -129 759 -128
rect 779 -129 780 -128
rect 849 -129 850 -128
rect 905 -129 906 -128
rect 919 -129 920 -128
rect 30 -131 31 -130
rect 37 -131 38 -130
rect 121 -131 122 -130
rect 205 -131 206 -130
rect 219 -131 220 -130
rect 282 -131 283 -130
rect 296 -131 297 -130
rect 303 -131 304 -130
rect 324 -131 325 -130
rect 338 -131 339 -130
rect 345 -131 346 -130
rect 352 -131 353 -130
rect 380 -131 381 -130
rect 429 -131 430 -130
rect 443 -131 444 -130
rect 457 -131 458 -130
rect 509 -131 510 -130
rect 541 -131 542 -130
rect 555 -131 556 -130
rect 695 -131 696 -130
rect 737 -131 738 -130
rect 751 -131 752 -130
rect 30 -133 31 -132
rect 51 -133 52 -132
rect 149 -133 150 -132
rect 376 -133 377 -132
rect 394 -133 395 -132
rect 429 -133 430 -132
rect 471 -133 472 -132
rect 555 -133 556 -132
rect 583 -133 584 -132
rect 653 -133 654 -132
rect 667 -133 668 -132
rect 786 -133 787 -132
rect 51 -135 52 -134
rect 58 -135 59 -134
rect 149 -135 150 -134
rect 481 -135 482 -134
rect 513 -135 514 -134
rect 583 -135 584 -134
rect 590 -135 591 -134
rect 688 -135 689 -134
rect 695 -135 696 -134
rect 765 -135 766 -134
rect 156 -137 157 -136
rect 166 -137 167 -136
rect 170 -137 171 -136
rect 380 -137 381 -136
rect 394 -137 395 -136
rect 415 -137 416 -136
rect 450 -137 451 -136
rect 471 -137 472 -136
rect 520 -137 521 -136
rect 779 -137 780 -136
rect 58 -139 59 -138
rect 156 -139 157 -138
rect 170 -139 171 -138
rect 187 -139 188 -138
rect 198 -139 199 -138
rect 376 -139 377 -138
rect 401 -139 402 -138
rect 415 -139 416 -138
rect 450 -139 451 -138
rect 548 -139 549 -138
rect 604 -139 605 -138
rect 667 -139 668 -138
rect 674 -139 675 -138
rect 793 -139 794 -138
rect 142 -141 143 -140
rect 401 -141 402 -140
rect 499 -141 500 -140
rect 548 -141 549 -140
rect 562 -141 563 -140
rect 674 -141 675 -140
rect 681 -141 682 -140
rect 807 -141 808 -140
rect 135 -143 136 -142
rect 499 -143 500 -142
rect 527 -143 528 -142
rect 562 -143 563 -142
rect 604 -143 605 -142
rect 723 -143 724 -142
rect 744 -143 745 -142
rect 800 -143 801 -142
rect 142 -145 143 -144
rect 163 -145 164 -144
rect 205 -145 206 -144
rect 212 -145 213 -144
rect 226 -145 227 -144
rect 348 -145 349 -144
rect 492 -145 493 -144
rect 527 -145 528 -144
rect 569 -145 570 -144
rect 723 -145 724 -144
rect 730 -145 731 -144
rect 800 -145 801 -144
rect 212 -147 213 -146
rect 275 -147 276 -146
rect 282 -147 283 -146
rect 390 -147 391 -146
rect 569 -147 570 -146
rect 702 -147 703 -146
rect 709 -147 710 -146
rect 737 -147 738 -146
rect 229 -149 230 -148
rect 359 -149 360 -148
rect 618 -149 619 -148
rect 681 -149 682 -148
rect 702 -149 703 -148
rect 845 -149 846 -148
rect 233 -151 234 -150
rect 352 -151 353 -150
rect 359 -151 360 -150
rect 366 -151 367 -150
rect 534 -151 535 -150
rect 618 -151 619 -150
rect 625 -151 626 -150
rect 730 -151 731 -150
rect 233 -153 234 -152
rect 247 -153 248 -152
rect 250 -153 251 -152
rect 254 -153 255 -152
rect 275 -153 276 -152
rect 467 -153 468 -152
rect 597 -153 598 -152
rect 625 -153 626 -152
rect 632 -153 633 -152
rect 688 -153 689 -152
rect 240 -155 241 -154
rect 317 -155 318 -154
rect 334 -155 335 -154
rect 513 -155 514 -154
rect 597 -155 598 -154
rect 716 -155 717 -154
rect 72 -157 73 -156
rect 317 -157 318 -156
rect 345 -157 346 -156
rect 422 -157 423 -156
rect 478 -157 479 -156
rect 632 -157 633 -156
rect 639 -157 640 -156
rect 765 -157 766 -156
rect 243 -159 244 -158
rect 320 -159 321 -158
rect 366 -159 367 -158
rect 383 -159 384 -158
rect 422 -159 423 -158
rect 772 -159 773 -158
rect 247 -161 248 -160
rect 261 -161 262 -160
rect 303 -161 304 -160
rect 331 -161 332 -160
rect 436 -161 437 -160
rect 639 -161 640 -160
rect 646 -161 647 -160
rect 709 -161 710 -160
rect 254 -163 255 -162
rect 289 -163 290 -162
rect 331 -163 332 -162
rect 443 -163 444 -162
rect 478 -163 479 -162
rect 814 -163 815 -162
rect 107 -165 108 -164
rect 289 -165 290 -164
rect 387 -165 388 -164
rect 436 -165 437 -164
rect 611 -165 612 -164
rect 646 -165 647 -164
rect 660 -165 661 -164
rect 716 -165 717 -164
rect 107 -167 108 -166
rect 128 -167 129 -166
rect 261 -167 262 -166
rect 268 -167 269 -166
rect 387 -167 388 -166
rect 485 -167 486 -166
rect 537 -167 538 -166
rect 660 -167 661 -166
rect 128 -169 129 -168
rect 138 -169 139 -168
rect 268 -169 269 -168
rect 310 -169 311 -168
rect 576 -169 577 -168
rect 611 -169 612 -168
rect 100 -171 101 -170
rect 310 -171 311 -170
rect 523 -171 524 -170
rect 576 -171 577 -170
rect 93 -173 94 -172
rect 100 -173 101 -172
rect 114 -173 115 -172
rect 138 -173 139 -172
rect 93 -175 94 -174
rect 177 -175 178 -174
rect 177 -177 178 -176
rect 191 -177 192 -176
rect 191 -179 192 -178
rect 488 -179 489 -178
rect 16 -190 17 -189
rect 303 -190 304 -189
rect 317 -190 318 -189
rect 576 -190 577 -189
rect 758 -190 759 -189
rect 870 -190 871 -189
rect 919 -190 920 -189
rect 947 -190 948 -189
rect 30 -192 31 -191
rect 65 -192 66 -191
rect 68 -192 69 -191
rect 103 -192 104 -191
rect 117 -192 118 -191
rect 198 -192 199 -191
rect 201 -192 202 -191
rect 233 -192 234 -191
rect 240 -192 241 -191
rect 331 -192 332 -191
rect 338 -192 339 -191
rect 436 -192 437 -191
rect 460 -192 461 -191
rect 730 -192 731 -191
rect 765 -192 766 -191
rect 814 -192 815 -191
rect 821 -192 822 -191
rect 919 -192 920 -191
rect 23 -194 24 -193
rect 68 -194 69 -193
rect 72 -194 73 -193
rect 201 -194 202 -193
rect 205 -194 206 -193
rect 352 -194 353 -193
rect 355 -194 356 -193
rect 436 -194 437 -193
rect 485 -194 486 -193
rect 884 -194 885 -193
rect 23 -196 24 -195
rect 100 -196 101 -195
rect 163 -196 164 -195
rect 177 -196 178 -195
rect 184 -196 185 -195
rect 212 -196 213 -195
rect 233 -196 234 -195
rect 268 -196 269 -195
rect 292 -196 293 -195
rect 387 -196 388 -195
rect 422 -196 423 -195
rect 555 -196 556 -195
rect 660 -196 661 -195
rect 730 -196 731 -195
rect 744 -196 745 -195
rect 765 -196 766 -195
rect 772 -196 773 -195
rect 877 -196 878 -195
rect 30 -198 31 -197
rect 114 -198 115 -197
rect 142 -198 143 -197
rect 212 -198 213 -197
rect 261 -198 262 -197
rect 268 -198 269 -197
rect 296 -198 297 -197
rect 317 -198 318 -197
rect 345 -198 346 -197
rect 905 -198 906 -197
rect 37 -200 38 -199
rect 247 -200 248 -199
rect 303 -200 304 -199
rect 373 -200 374 -199
rect 380 -200 381 -199
rect 555 -200 556 -199
rect 674 -200 675 -199
rect 758 -200 759 -199
rect 786 -200 787 -199
rect 856 -200 857 -199
rect 859 -200 860 -199
rect 933 -200 934 -199
rect 44 -202 45 -201
rect 282 -202 283 -201
rect 352 -202 353 -201
rect 639 -202 640 -201
rect 702 -202 703 -201
rect 744 -202 745 -201
rect 751 -202 752 -201
rect 786 -202 787 -201
rect 793 -202 794 -201
rect 863 -202 864 -201
rect 72 -204 73 -203
rect 156 -204 157 -203
rect 170 -204 171 -203
rect 177 -204 178 -203
rect 187 -204 188 -203
rect 296 -204 297 -203
rect 373 -204 374 -203
rect 394 -204 395 -203
rect 408 -204 409 -203
rect 422 -204 423 -203
rect 495 -204 496 -203
rect 520 -204 521 -203
rect 527 -204 528 -203
rect 674 -204 675 -203
rect 681 -204 682 -203
rect 751 -204 752 -203
rect 800 -204 801 -203
rect 891 -204 892 -203
rect 79 -206 80 -205
rect 240 -206 241 -205
rect 247 -206 248 -205
rect 275 -206 276 -205
rect 408 -206 409 -205
rect 537 -206 538 -205
rect 541 -206 542 -205
rect 576 -206 577 -205
rect 604 -206 605 -205
rect 639 -206 640 -205
rect 681 -206 682 -205
rect 688 -206 689 -205
rect 709 -206 710 -205
rect 772 -206 773 -205
rect 800 -206 801 -205
rect 842 -206 843 -205
rect 79 -208 80 -207
rect 348 -208 349 -207
rect 450 -208 451 -207
rect 527 -208 528 -207
rect 534 -208 535 -207
rect 590 -208 591 -207
rect 625 -208 626 -207
rect 688 -208 689 -207
rect 737 -208 738 -207
rect 793 -208 794 -207
rect 807 -208 808 -207
rect 940 -208 941 -207
rect 107 -210 108 -209
rect 394 -210 395 -209
rect 429 -210 430 -209
rect 450 -210 451 -209
rect 478 -210 479 -209
rect 541 -210 542 -209
rect 548 -210 549 -209
rect 625 -210 626 -209
rect 646 -210 647 -209
rect 709 -210 710 -209
rect 716 -210 717 -209
rect 807 -210 808 -209
rect 821 -210 822 -209
rect 849 -210 850 -209
rect 58 -212 59 -211
rect 548 -212 549 -211
rect 583 -212 584 -211
rect 604 -212 605 -211
rect 667 -212 668 -211
rect 737 -212 738 -211
rect 779 -212 780 -211
rect 849 -212 850 -211
rect 51 -214 52 -213
rect 58 -214 59 -213
rect 107 -214 108 -213
rect 135 -214 136 -213
rect 142 -214 143 -213
rect 149 -214 150 -213
rect 187 -214 188 -213
rect 583 -214 584 -213
rect 695 -214 696 -213
rect 716 -214 717 -213
rect 723 -214 724 -213
rect 779 -214 780 -213
rect 828 -214 829 -213
rect 926 -214 927 -213
rect 51 -216 52 -215
rect 65 -216 66 -215
rect 114 -216 115 -215
rect 128 -216 129 -215
rect 149 -216 150 -215
rect 219 -216 220 -215
rect 254 -216 255 -215
rect 282 -216 283 -215
rect 324 -216 325 -215
rect 429 -216 430 -215
rect 464 -216 465 -215
rect 828 -216 829 -215
rect 835 -216 836 -215
rect 898 -216 899 -215
rect 121 -218 122 -217
rect 128 -218 129 -217
rect 191 -218 192 -217
rect 254 -218 255 -217
rect 275 -218 276 -217
rect 618 -218 619 -217
rect 632 -218 633 -217
rect 695 -218 696 -217
rect 93 -220 94 -219
rect 191 -220 192 -219
rect 310 -220 311 -219
rect 324 -220 325 -219
rect 345 -220 346 -219
rect 478 -220 479 -219
rect 499 -220 500 -219
rect 660 -220 661 -219
rect 93 -222 94 -221
rect 912 -222 913 -221
rect 121 -224 122 -223
rect 229 -224 230 -223
rect 467 -224 468 -223
rect 667 -224 668 -223
rect 173 -226 174 -225
rect 310 -226 311 -225
rect 366 -226 367 -225
rect 467 -226 468 -225
rect 471 -226 472 -225
rect 499 -226 500 -225
rect 513 -226 514 -225
rect 702 -226 703 -225
rect 289 -228 290 -227
rect 366 -228 367 -227
rect 457 -228 458 -227
rect 471 -228 472 -227
rect 506 -228 507 -227
rect 513 -228 514 -227
rect 593 -228 594 -227
rect 835 -228 836 -227
rect 443 -230 444 -229
rect 506 -230 507 -229
rect 597 -230 598 -229
rect 632 -230 633 -229
rect 653 -230 654 -229
rect 723 -230 724 -229
rect 415 -232 416 -231
rect 443 -232 444 -231
rect 611 -232 612 -231
rect 618 -232 619 -231
rect 401 -234 402 -233
rect 415 -234 416 -233
rect 425 -234 426 -233
rect 653 -234 654 -233
rect 100 -236 101 -235
rect 401 -236 402 -235
rect 569 -236 570 -235
rect 611 -236 612 -235
rect 226 -238 227 -237
rect 569 -238 570 -237
rect 30 -249 31 -248
rect 159 -249 160 -248
rect 170 -249 171 -248
rect 212 -249 213 -248
rect 233 -249 234 -248
rect 292 -249 293 -248
rect 352 -249 353 -248
rect 506 -249 507 -248
rect 579 -249 580 -248
rect 772 -249 773 -248
rect 877 -249 878 -248
rect 961 -249 962 -248
rect 975 -249 976 -248
rect 982 -249 983 -248
rect 1087 -249 1088 -248
rect 1094 -249 1095 -248
rect 33 -251 34 -250
rect 485 -251 486 -250
rect 488 -251 489 -250
rect 779 -251 780 -250
rect 877 -251 878 -250
rect 933 -251 934 -250
rect 947 -251 948 -250
rect 975 -251 976 -250
rect 37 -253 38 -252
rect 198 -253 199 -252
rect 208 -253 209 -252
rect 555 -253 556 -252
rect 586 -253 587 -252
rect 828 -253 829 -252
rect 37 -255 38 -254
rect 89 -255 90 -254
rect 93 -255 94 -254
rect 247 -255 248 -254
rect 254 -255 255 -254
rect 282 -255 283 -254
rect 380 -255 381 -254
rect 394 -255 395 -254
rect 436 -255 437 -254
rect 506 -255 507 -254
rect 527 -255 528 -254
rect 555 -255 556 -254
rect 593 -255 594 -254
rect 653 -255 654 -254
rect 758 -255 759 -254
rect 772 -255 773 -254
rect 779 -255 780 -254
rect 793 -255 794 -254
rect 828 -255 829 -254
rect 884 -255 885 -254
rect 44 -257 45 -256
rect 289 -257 290 -256
rect 383 -257 384 -256
rect 590 -257 591 -256
rect 600 -257 601 -256
rect 709 -257 710 -256
rect 765 -257 766 -256
rect 800 -257 801 -256
rect 884 -257 885 -256
rect 891 -257 892 -256
rect 47 -259 48 -258
rect 86 -259 87 -258
rect 93 -259 94 -258
rect 303 -259 304 -258
rect 394 -259 395 -258
rect 513 -259 514 -258
rect 520 -259 521 -258
rect 527 -259 528 -258
rect 597 -259 598 -258
rect 765 -259 766 -258
rect 891 -259 892 -258
rect 954 -259 955 -258
rect 58 -261 59 -260
rect 191 -261 192 -260
rect 205 -261 206 -260
rect 254 -261 255 -260
rect 275 -261 276 -260
rect 481 -261 482 -260
rect 495 -261 496 -260
rect 674 -261 675 -260
rect 702 -261 703 -260
rect 954 -261 955 -260
rect 23 -263 24 -262
rect 191 -263 192 -262
rect 233 -263 234 -262
rect 457 -263 458 -262
rect 464 -263 465 -262
rect 646 -263 647 -262
rect 653 -263 654 -262
rect 730 -263 731 -262
rect 23 -265 24 -264
rect 51 -265 52 -264
rect 65 -265 66 -264
rect 439 -265 440 -264
rect 478 -265 479 -264
rect 835 -265 836 -264
rect 79 -267 80 -266
rect 212 -267 213 -266
rect 338 -267 339 -266
rect 457 -267 458 -266
rect 499 -267 500 -266
rect 513 -267 514 -266
rect 562 -267 563 -266
rect 597 -267 598 -266
rect 604 -267 605 -266
rect 674 -267 675 -266
rect 695 -267 696 -266
rect 730 -267 731 -266
rect 79 -269 80 -268
rect 793 -269 794 -268
rect 82 -271 83 -270
rect 100 -271 101 -270
rect 103 -271 104 -270
rect 128 -271 129 -270
rect 135 -271 136 -270
rect 247 -271 248 -270
rect 331 -271 332 -270
rect 338 -271 339 -270
rect 373 -271 374 -270
rect 520 -271 521 -270
rect 541 -271 542 -270
rect 562 -271 563 -270
rect 583 -271 584 -270
rect 604 -271 605 -270
rect 618 -271 619 -270
rect 646 -271 647 -270
rect 695 -271 696 -270
rect 737 -271 738 -270
rect 107 -273 108 -272
rect 569 -273 570 -272
rect 576 -273 577 -272
rect 618 -273 619 -272
rect 667 -273 668 -272
rect 737 -273 738 -272
rect 117 -275 118 -274
rect 331 -275 332 -274
rect 359 -275 360 -274
rect 373 -275 374 -274
rect 411 -275 412 -274
rect 758 -275 759 -274
rect 128 -277 129 -276
rect 324 -277 325 -276
rect 359 -277 360 -276
rect 415 -277 416 -276
rect 450 -277 451 -276
rect 478 -277 479 -276
rect 583 -277 584 -276
rect 681 -277 682 -276
rect 702 -277 703 -276
rect 723 -277 724 -276
rect 135 -279 136 -278
rect 261 -279 262 -278
rect 317 -279 318 -278
rect 324 -279 325 -278
rect 415 -279 416 -278
rect 835 -279 836 -278
rect 142 -281 143 -280
rect 275 -281 276 -280
rect 422 -281 423 -280
rect 450 -281 451 -280
rect 471 -281 472 -280
rect 499 -281 500 -280
rect 639 -281 640 -280
rect 667 -281 668 -280
rect 681 -281 682 -280
rect 688 -281 689 -280
rect 709 -281 710 -280
rect 849 -281 850 -280
rect 114 -283 115 -282
rect 688 -283 689 -282
rect 723 -283 724 -282
rect 751 -283 752 -282
rect 849 -283 850 -282
rect 926 -283 927 -282
rect 114 -285 115 -284
rect 163 -285 164 -284
rect 170 -285 171 -284
rect 296 -285 297 -284
rect 422 -285 423 -284
rect 429 -285 430 -284
rect 471 -285 472 -284
rect 814 -285 815 -284
rect 912 -285 913 -284
rect 926 -285 927 -284
rect 145 -287 146 -286
rect 303 -287 304 -286
rect 429 -287 430 -286
rect 443 -287 444 -286
rect 474 -287 475 -286
rect 569 -287 570 -286
rect 625 -287 626 -286
rect 639 -287 640 -286
rect 744 -287 745 -286
rect 751 -287 752 -286
rect 912 -287 913 -286
rect 940 -287 941 -286
rect 156 -289 157 -288
rect 548 -289 549 -288
rect 625 -289 626 -288
rect 660 -289 661 -288
rect 716 -289 717 -288
rect 744 -289 745 -288
rect 821 -289 822 -288
rect 940 -289 941 -288
rect 156 -291 157 -290
rect 205 -291 206 -290
rect 219 -291 220 -290
rect 296 -291 297 -290
rect 401 -291 402 -290
rect 443 -291 444 -290
rect 492 -291 493 -290
rect 814 -291 815 -290
rect 163 -293 164 -292
rect 548 -293 549 -292
rect 632 -293 633 -292
rect 660 -293 661 -292
rect 786 -293 787 -292
rect 821 -293 822 -292
rect 177 -295 178 -294
rect 184 -295 185 -294
rect 219 -295 220 -294
rect 240 -295 241 -294
rect 264 -295 265 -294
rect 317 -295 318 -294
rect 366 -295 367 -294
rect 401 -295 402 -294
rect 492 -295 493 -294
rect 870 -295 871 -294
rect 16 -297 17 -296
rect 177 -297 178 -296
rect 226 -297 227 -296
rect 240 -297 241 -296
rect 310 -297 311 -296
rect 366 -297 367 -296
rect 611 -297 612 -296
rect 632 -297 633 -296
rect 786 -297 787 -296
rect 807 -297 808 -296
rect 870 -297 871 -296
rect 919 -297 920 -296
rect 16 -299 17 -298
rect 464 -299 465 -298
rect 807 -299 808 -298
rect 856 -299 857 -298
rect 863 -299 864 -298
rect 919 -299 920 -298
rect 72 -301 73 -300
rect 310 -301 311 -300
rect 408 -301 409 -300
rect 611 -301 612 -300
rect 842 -301 843 -300
rect 856 -301 857 -300
rect 863 -301 864 -300
rect 898 -301 899 -300
rect 72 -303 73 -302
rect 345 -303 346 -302
rect 842 -303 843 -302
rect 968 -303 969 -302
rect 149 -305 150 -304
rect 345 -305 346 -304
rect 898 -305 899 -304
rect 936 -305 937 -304
rect 149 -307 150 -306
rect 387 -307 388 -306
rect 229 -309 230 -308
rect 261 -309 262 -308
rect 9 -320 10 -319
rect 145 -320 146 -319
rect 205 -320 206 -319
rect 208 -320 209 -319
rect 226 -320 227 -319
rect 268 -320 269 -319
rect 296 -320 297 -319
rect 408 -320 409 -319
rect 436 -320 437 -319
rect 926 -320 927 -319
rect 933 -320 934 -319
rect 982 -320 983 -319
rect 999 -320 1000 -319
rect 1066 -320 1067 -319
rect 1094 -320 1095 -319
rect 1108 -320 1109 -319
rect 16 -322 17 -321
rect 474 -322 475 -321
rect 523 -322 524 -321
rect 653 -322 654 -321
rect 681 -322 682 -321
rect 684 -322 685 -321
rect 716 -322 717 -321
rect 905 -322 906 -321
rect 947 -322 948 -321
rect 968 -322 969 -321
rect 16 -324 17 -323
rect 135 -324 136 -323
rect 208 -324 209 -323
rect 292 -324 293 -323
rect 317 -324 318 -323
rect 464 -324 465 -323
rect 527 -324 528 -323
rect 544 -324 545 -323
rect 548 -324 549 -323
rect 961 -324 962 -323
rect 964 -324 965 -323
rect 1052 -324 1053 -323
rect 23 -326 24 -325
rect 117 -326 118 -325
rect 121 -326 122 -325
rect 296 -326 297 -325
rect 331 -326 332 -325
rect 467 -326 468 -325
rect 541 -326 542 -325
rect 954 -326 955 -325
rect 23 -328 24 -327
rect 303 -328 304 -327
rect 345 -328 346 -327
rect 383 -328 384 -327
rect 390 -328 391 -327
rect 520 -328 521 -327
rect 534 -328 535 -327
rect 541 -328 542 -327
rect 548 -328 549 -327
rect 919 -328 920 -327
rect 37 -330 38 -329
rect 51 -330 52 -329
rect 58 -330 59 -329
rect 418 -330 419 -329
rect 443 -330 444 -329
rect 583 -330 584 -329
rect 632 -330 633 -329
rect 653 -330 654 -329
rect 681 -330 682 -329
rect 884 -330 885 -329
rect 898 -330 899 -329
rect 982 -330 983 -329
rect 40 -332 41 -331
rect 58 -332 59 -331
rect 65 -332 66 -331
rect 163 -332 164 -331
rect 212 -332 213 -331
rect 436 -332 437 -331
rect 443 -332 444 -331
rect 488 -332 489 -331
rect 499 -332 500 -331
rect 534 -332 535 -331
rect 579 -332 580 -331
rect 905 -332 906 -331
rect 44 -334 45 -333
rect 145 -334 146 -333
rect 212 -334 213 -333
rect 485 -334 486 -333
rect 618 -334 619 -333
rect 632 -334 633 -333
rect 716 -334 717 -333
rect 814 -334 815 -333
rect 821 -334 822 -333
rect 926 -334 927 -333
rect 65 -336 66 -335
rect 107 -336 108 -335
rect 121 -336 122 -335
rect 324 -336 325 -335
rect 338 -336 339 -335
rect 345 -336 346 -335
rect 352 -336 353 -335
rect 355 -336 356 -335
rect 359 -336 360 -335
rect 415 -336 416 -335
rect 422 -336 423 -335
rect 499 -336 500 -335
rect 786 -336 787 -335
rect 884 -336 885 -335
rect 901 -336 902 -335
rect 975 -336 976 -335
rect 30 -338 31 -337
rect 422 -338 423 -337
rect 453 -338 454 -337
rect 772 -338 773 -337
rect 807 -338 808 -337
rect 821 -338 822 -337
rect 828 -338 829 -337
rect 975 -338 976 -337
rect 93 -340 94 -339
rect 289 -340 290 -339
rect 352 -340 353 -339
rect 394 -340 395 -339
rect 401 -340 402 -339
rect 408 -340 409 -339
rect 457 -340 458 -339
rect 527 -340 528 -339
rect 702 -340 703 -339
rect 772 -340 773 -339
rect 835 -340 836 -339
rect 1010 -340 1011 -339
rect 93 -342 94 -341
rect 180 -342 181 -341
rect 191 -342 192 -341
rect 618 -342 619 -341
rect 639 -342 640 -341
rect 702 -342 703 -341
rect 744 -342 745 -341
rect 786 -342 787 -341
rect 842 -342 843 -341
rect 947 -342 948 -341
rect 100 -344 101 -343
rect 107 -344 108 -343
rect 135 -344 136 -343
rect 163 -344 164 -343
rect 254 -344 255 -343
rect 268 -344 269 -343
rect 275 -344 276 -343
rect 303 -344 304 -343
rect 359 -344 360 -343
rect 478 -344 479 -343
rect 506 -344 507 -343
rect 828 -344 829 -343
rect 849 -344 850 -343
rect 1017 -344 1018 -343
rect 79 -346 80 -345
rect 478 -346 479 -345
rect 590 -346 591 -345
rect 639 -346 640 -345
rect 723 -346 724 -345
rect 849 -346 850 -345
rect 863 -346 864 -345
rect 989 -346 990 -345
rect 79 -348 80 -347
rect 170 -348 171 -347
rect 219 -348 220 -347
rect 254 -348 255 -347
rect 261 -348 262 -347
rect 331 -348 332 -347
rect 380 -348 381 -347
rect 919 -348 920 -347
rect 72 -350 73 -349
rect 380 -350 381 -349
rect 394 -350 395 -349
rect 471 -350 472 -349
rect 474 -350 475 -349
rect 723 -350 724 -349
rect 751 -350 752 -349
rect 807 -350 808 -349
rect 870 -350 871 -349
rect 1003 -350 1004 -349
rect 72 -352 73 -351
rect 86 -352 87 -351
rect 100 -352 101 -351
rect 110 -352 111 -351
rect 149 -352 150 -351
rect 485 -352 486 -351
rect 569 -352 570 -351
rect 590 -352 591 -351
rect 684 -352 685 -351
rect 744 -352 745 -351
rect 758 -352 759 -351
rect 863 -352 864 -351
rect 870 -352 871 -351
rect 912 -352 913 -351
rect 86 -354 87 -353
rect 366 -354 367 -353
rect 401 -354 402 -353
rect 814 -354 815 -353
rect 877 -354 878 -353
rect 1024 -354 1025 -353
rect 149 -356 150 -355
rect 247 -356 248 -355
rect 275 -356 276 -355
rect 450 -356 451 -355
rect 555 -356 556 -355
rect 569 -356 570 -355
rect 586 -356 587 -355
rect 758 -356 759 -355
rect 765 -356 766 -355
rect 877 -356 878 -355
rect 891 -356 892 -355
rect 912 -356 913 -355
rect 191 -358 192 -357
rect 450 -358 451 -357
rect 513 -358 514 -357
rect 555 -358 556 -357
rect 730 -358 731 -357
rect 765 -358 766 -357
rect 793 -358 794 -357
rect 891 -358 892 -357
rect 198 -360 199 -359
rect 261 -360 262 -359
rect 282 -360 283 -359
rect 324 -360 325 -359
rect 366 -360 367 -359
rect 551 -360 552 -359
rect 688 -360 689 -359
rect 793 -360 794 -359
rect 800 -360 801 -359
rect 842 -360 843 -359
rect 114 -362 115 -361
rect 282 -362 283 -361
rect 404 -362 405 -361
rect 835 -362 836 -361
rect 128 -364 129 -363
rect 198 -364 199 -363
rect 219 -364 220 -363
rect 565 -364 566 -363
rect 611 -364 612 -363
rect 688 -364 689 -363
rect 695 -364 696 -363
rect 800 -364 801 -363
rect 33 -366 34 -365
rect 128 -366 129 -365
rect 240 -366 241 -365
rect 247 -366 248 -365
rect 429 -366 430 -365
rect 457 -366 458 -365
rect 492 -366 493 -365
rect 513 -366 514 -365
rect 611 -366 612 -365
rect 674 -366 675 -365
rect 719 -366 720 -365
rect 730 -366 731 -365
rect 737 -366 738 -365
rect 751 -366 752 -365
rect 240 -368 241 -367
rect 936 -368 937 -367
rect 429 -370 430 -369
rect 520 -370 521 -369
rect 625 -370 626 -369
rect 695 -370 696 -369
rect 737 -370 738 -369
rect 940 -370 941 -369
rect 492 -372 493 -371
rect 954 -372 955 -371
rect 495 -374 496 -373
rect 551 -374 552 -373
rect 597 -374 598 -373
rect 625 -374 626 -373
rect 660 -374 661 -373
rect 674 -374 675 -373
rect 856 -374 857 -373
rect 940 -374 941 -373
rect 562 -376 563 -375
rect 597 -376 598 -375
rect 646 -376 647 -375
rect 660 -376 661 -375
rect 779 -376 780 -375
rect 856 -376 857 -375
rect 338 -378 339 -377
rect 646 -378 647 -377
rect 779 -378 780 -377
rect 961 -378 962 -377
rect 562 -380 563 -379
rect 709 -380 710 -379
rect 667 -382 668 -381
rect 709 -382 710 -381
rect 604 -384 605 -383
rect 667 -384 668 -383
rect 387 -386 388 -385
rect 604 -386 605 -385
rect 373 -388 374 -387
rect 387 -388 388 -387
rect 310 -390 311 -389
rect 373 -390 374 -389
rect 233 -392 234 -391
rect 310 -392 311 -391
rect 177 -394 178 -393
rect 233 -394 234 -393
rect 16 -405 17 -404
rect 138 -405 139 -404
rect 142 -405 143 -404
rect 149 -405 150 -404
rect 180 -405 181 -404
rect 198 -405 199 -404
rect 233 -405 234 -404
rect 275 -405 276 -404
rect 282 -405 283 -404
rect 285 -405 286 -404
rect 306 -405 307 -404
rect 324 -405 325 -404
rect 331 -405 332 -404
rect 404 -405 405 -404
rect 422 -405 423 -404
rect 754 -405 755 -404
rect 800 -405 801 -404
rect 1045 -405 1046 -404
rect 1066 -405 1067 -404
rect 1139 -405 1140 -404
rect 16 -407 17 -406
rect 51 -407 52 -406
rect 58 -407 59 -406
rect 198 -407 199 -406
rect 233 -407 234 -406
rect 565 -407 566 -406
rect 576 -407 577 -406
rect 590 -407 591 -406
rect 600 -407 601 -406
rect 870 -407 871 -406
rect 877 -407 878 -406
rect 1101 -407 1102 -406
rect 1108 -407 1109 -406
rect 1150 -407 1151 -406
rect 23 -409 24 -408
rect 390 -409 391 -408
rect 401 -409 402 -408
rect 793 -409 794 -408
rect 800 -409 801 -408
rect 807 -409 808 -408
rect 863 -409 864 -408
rect 1115 -409 1116 -408
rect 23 -411 24 -410
rect 114 -411 115 -410
rect 142 -411 143 -410
rect 173 -411 174 -410
rect 191 -411 192 -410
rect 205 -411 206 -410
rect 247 -411 248 -410
rect 250 -411 251 -410
rect 254 -411 255 -410
rect 320 -411 321 -410
rect 331 -411 332 -410
rect 485 -411 486 -410
rect 502 -411 503 -410
rect 996 -411 997 -410
rect 1003 -411 1004 -410
rect 1087 -411 1088 -410
rect 37 -413 38 -412
rect 212 -413 213 -412
rect 247 -413 248 -412
rect 261 -413 262 -412
rect 268 -413 269 -412
rect 278 -413 279 -412
rect 282 -413 283 -412
rect 289 -413 290 -412
rect 296 -413 297 -412
rect 324 -413 325 -412
rect 338 -413 339 -412
rect 429 -413 430 -412
rect 436 -413 437 -412
rect 492 -413 493 -412
rect 509 -413 510 -412
rect 695 -413 696 -412
rect 740 -413 741 -412
rect 1080 -413 1081 -412
rect 51 -415 52 -414
rect 110 -415 111 -414
rect 128 -415 129 -414
rect 191 -415 192 -414
rect 219 -415 220 -414
rect 296 -415 297 -414
rect 317 -415 318 -414
rect 450 -415 451 -414
rect 478 -415 479 -414
rect 492 -415 493 -414
rect 523 -415 524 -414
rect 898 -415 899 -414
rect 919 -415 920 -414
rect 996 -415 997 -414
rect 1010 -415 1011 -414
rect 1108 -415 1109 -414
rect 58 -417 59 -416
rect 79 -417 80 -416
rect 107 -417 108 -416
rect 114 -417 115 -416
rect 128 -417 129 -416
rect 156 -417 157 -416
rect 219 -417 220 -416
rect 303 -417 304 -416
rect 317 -417 318 -416
rect 380 -417 381 -416
rect 425 -417 426 -416
rect 1066 -417 1067 -416
rect 65 -419 66 -418
rect 89 -419 90 -418
rect 145 -419 146 -418
rect 208 -419 209 -418
rect 240 -419 241 -418
rect 338 -419 339 -418
rect 341 -419 342 -418
rect 345 -419 346 -418
rect 359 -419 360 -418
rect 415 -419 416 -418
rect 429 -419 430 -418
rect 551 -419 552 -418
rect 586 -419 587 -418
rect 716 -419 717 -418
rect 730 -419 731 -418
rect 919 -419 920 -418
rect 947 -419 948 -418
rect 1038 -419 1039 -418
rect 1041 -419 1042 -418
rect 1052 -419 1053 -418
rect 44 -421 45 -420
rect 947 -421 948 -420
rect 954 -421 955 -420
rect 1052 -421 1053 -420
rect 44 -423 45 -422
rect 278 -423 279 -422
rect 285 -423 286 -422
rect 289 -423 290 -422
rect 345 -423 346 -422
rect 499 -423 500 -422
rect 548 -423 549 -422
rect 1031 -423 1032 -422
rect 65 -425 66 -424
rect 352 -425 353 -424
rect 366 -425 367 -424
rect 436 -425 437 -424
rect 485 -425 486 -424
rect 527 -425 528 -424
rect 590 -425 591 -424
rect 597 -425 598 -424
rect 646 -425 647 -424
rect 954 -425 955 -424
rect 975 -425 976 -424
rect 1094 -425 1095 -424
rect 72 -427 73 -426
rect 135 -427 136 -426
rect 156 -427 157 -426
rect 411 -427 412 -426
rect 478 -427 479 -426
rect 597 -427 598 -426
rect 639 -427 640 -426
rect 646 -427 647 -426
rect 660 -427 661 -426
rect 695 -427 696 -426
rect 709 -427 710 -426
rect 716 -427 717 -426
rect 744 -427 745 -426
rect 877 -427 878 -426
rect 905 -427 906 -426
rect 1010 -427 1011 -426
rect 1017 -427 1018 -426
rect 1122 -427 1123 -426
rect 30 -429 31 -428
rect 660 -429 661 -428
rect 674 -429 675 -428
rect 709 -429 710 -428
rect 744 -429 745 -428
rect 758 -429 759 -428
rect 772 -429 773 -428
rect 1003 -429 1004 -428
rect 1024 -429 1025 -428
rect 1129 -429 1130 -428
rect 72 -431 73 -430
rect 86 -431 87 -430
rect 93 -431 94 -430
rect 352 -431 353 -430
rect 380 -431 381 -430
rect 901 -431 902 -430
rect 926 -431 927 -430
rect 1024 -431 1025 -430
rect 12 -433 13 -432
rect 86 -433 87 -432
rect 93 -433 94 -432
rect 121 -433 122 -432
rect 240 -433 241 -432
rect 635 -433 636 -432
rect 653 -433 654 -432
rect 674 -433 675 -432
rect 688 -433 689 -432
rect 730 -433 731 -432
rect 765 -433 766 -432
rect 772 -433 773 -432
rect 793 -433 794 -432
rect 849 -433 850 -432
rect 870 -433 871 -432
rect 912 -433 913 -432
rect 926 -433 927 -432
rect 989 -433 990 -432
rect 79 -435 80 -434
rect 513 -435 514 -434
rect 527 -435 528 -434
rect 562 -435 563 -434
rect 569 -435 570 -434
rect 765 -435 766 -434
rect 779 -435 780 -434
rect 989 -435 990 -434
rect 121 -437 122 -436
rect 163 -437 164 -436
rect 254 -437 255 -436
rect 394 -437 395 -436
rect 408 -437 409 -436
rect 415 -437 416 -436
rect 457 -437 458 -436
rect 513 -437 514 -436
rect 534 -437 535 -436
rect 569 -437 570 -436
rect 625 -437 626 -436
rect 639 -437 640 -436
rect 653 -437 654 -436
rect 737 -437 738 -436
rect 807 -437 808 -436
rect 821 -437 822 -436
rect 835 -437 836 -436
rect 975 -437 976 -436
rect 982 -437 983 -436
rect 1073 -437 1074 -436
rect 149 -439 150 -438
rect 457 -439 458 -438
rect 471 -439 472 -438
rect 779 -439 780 -438
rect 814 -439 815 -438
rect 905 -439 906 -438
rect 940 -439 941 -438
rect 1031 -439 1032 -438
rect 163 -441 164 -440
rect 177 -441 178 -440
rect 268 -441 269 -440
rect 443 -441 444 -440
rect 520 -441 521 -440
rect 821 -441 822 -440
rect 835 -441 836 -440
rect 884 -441 885 -440
rect 940 -441 941 -440
rect 961 -441 962 -440
rect 982 -441 983 -440
rect 1059 -441 1060 -440
rect 170 -443 171 -442
rect 814 -443 815 -442
rect 842 -443 843 -442
rect 863 -443 864 -442
rect 884 -443 885 -442
rect 968 -443 969 -442
rect 170 -445 171 -444
rect 226 -445 227 -444
rect 303 -445 304 -444
rect 842 -445 843 -444
rect 856 -445 857 -444
rect 968 -445 969 -444
rect 177 -447 178 -446
rect 310 -447 311 -446
rect 387 -447 388 -446
rect 394 -447 395 -446
rect 408 -447 409 -446
rect 1017 -447 1018 -446
rect 310 -449 311 -448
rect 579 -449 580 -448
rect 604 -449 605 -448
rect 625 -449 626 -448
rect 681 -449 682 -448
rect 912 -449 913 -448
rect 933 -449 934 -448
rect 961 -449 962 -448
rect 443 -451 444 -450
rect 464 -451 465 -450
rect 474 -451 475 -450
rect 856 -451 857 -450
rect 891 -451 892 -450
rect 933 -451 934 -450
rect 464 -453 465 -452
rect 737 -453 738 -452
rect 828 -453 829 -452
rect 891 -453 892 -452
rect 520 -455 521 -454
rect 667 -455 668 -454
rect 681 -455 682 -454
rect 1048 -455 1049 -454
rect 534 -457 535 -456
rect 541 -457 542 -456
rect 604 -457 605 -456
rect 618 -457 619 -456
rect 632 -457 633 -456
rect 667 -457 668 -456
rect 688 -457 689 -456
rect 702 -457 703 -456
rect 723 -457 724 -456
rect 758 -457 759 -456
rect 786 -457 787 -456
rect 828 -457 829 -456
rect 229 -459 230 -458
rect 541 -459 542 -458
rect 583 -459 584 -458
rect 618 -459 619 -458
rect 723 -459 724 -458
rect 849 -459 850 -458
rect 366 -461 367 -460
rect 583 -461 584 -460
rect 751 -461 752 -460
rect 786 -461 787 -460
rect 404 -463 405 -462
rect 702 -463 703 -462
rect 9 -474 10 -473
rect 310 -474 311 -473
rect 324 -474 325 -473
rect 345 -474 346 -473
rect 348 -474 349 -473
rect 635 -474 636 -473
rect 660 -474 661 -473
rect 968 -474 969 -473
rect 975 -474 976 -473
rect 1143 -474 1144 -473
rect 1174 -474 1175 -473
rect 1178 -474 1179 -473
rect 16 -476 17 -475
rect 110 -476 111 -475
rect 135 -476 136 -475
rect 142 -476 143 -475
rect 156 -476 157 -475
rect 530 -476 531 -475
rect 537 -476 538 -475
rect 1045 -476 1046 -475
rect 16 -478 17 -477
rect 100 -478 101 -477
rect 107 -478 108 -477
rect 254 -478 255 -477
rect 261 -478 262 -477
rect 278 -478 279 -477
rect 296 -478 297 -477
rect 310 -478 311 -477
rect 397 -478 398 -477
rect 520 -478 521 -477
rect 527 -478 528 -477
rect 989 -478 990 -477
rect 1045 -478 1046 -477
rect 1059 -478 1060 -477
rect 37 -480 38 -479
rect 303 -480 304 -479
rect 401 -480 402 -479
rect 513 -480 514 -479
rect 527 -480 528 -479
rect 534 -480 535 -479
rect 562 -480 563 -479
rect 1122 -480 1123 -479
rect 37 -482 38 -481
rect 201 -482 202 -481
rect 205 -482 206 -481
rect 226 -482 227 -481
rect 240 -482 241 -481
rect 296 -482 297 -481
rect 352 -482 353 -481
rect 401 -482 402 -481
rect 436 -482 437 -481
rect 600 -482 601 -481
rect 632 -482 633 -481
rect 1129 -482 1130 -481
rect 23 -484 24 -483
rect 205 -484 206 -483
rect 219 -484 220 -483
rect 390 -484 391 -483
rect 415 -484 416 -483
rect 436 -484 437 -483
rect 450 -484 451 -483
rect 663 -484 664 -483
rect 695 -484 696 -483
rect 737 -484 738 -483
rect 751 -484 752 -483
rect 856 -484 857 -483
rect 870 -484 871 -483
rect 968 -484 969 -483
rect 975 -484 976 -483
rect 996 -484 997 -483
rect 1059 -484 1060 -483
rect 1108 -484 1109 -483
rect 1122 -484 1123 -483
rect 1139 -484 1140 -483
rect 23 -486 24 -485
rect 30 -486 31 -485
rect 72 -486 73 -485
rect 275 -486 276 -485
rect 289 -486 290 -485
rect 303 -486 304 -485
rect 380 -486 381 -485
rect 513 -486 514 -485
rect 565 -486 566 -485
rect 1094 -486 1095 -485
rect 58 -488 59 -487
rect 380 -488 381 -487
rect 415 -488 416 -487
rect 478 -488 479 -487
rect 506 -488 507 -487
rect 730 -488 731 -487
rect 733 -488 734 -487
rect 1101 -488 1102 -487
rect 58 -490 59 -489
rect 373 -490 374 -489
rect 450 -490 451 -489
rect 485 -490 486 -489
rect 583 -490 584 -489
rect 590 -490 591 -489
rect 593 -490 594 -489
rect 1115 -490 1116 -489
rect 79 -492 80 -491
rect 499 -492 500 -491
rect 586 -492 587 -491
rect 1003 -492 1004 -491
rect 1010 -492 1011 -491
rect 1101 -492 1102 -491
rect 1115 -492 1116 -491
rect 1150 -492 1151 -491
rect 86 -494 87 -493
rect 947 -494 948 -493
rect 961 -494 962 -493
rect 982 -494 983 -493
rect 989 -494 990 -493
rect 1024 -494 1025 -493
rect 86 -496 87 -495
rect 114 -496 115 -495
rect 142 -496 143 -495
rect 366 -496 367 -495
rect 457 -496 458 -495
rect 842 -496 843 -495
rect 961 -496 962 -495
rect 1017 -496 1018 -495
rect 93 -498 94 -497
rect 156 -498 157 -497
rect 166 -498 167 -497
rect 1066 -498 1067 -497
rect 93 -500 94 -499
rect 121 -500 122 -499
rect 170 -500 171 -499
rect 219 -500 220 -499
rect 240 -500 241 -499
rect 247 -500 248 -499
rect 261 -500 262 -499
rect 429 -500 430 -499
rect 460 -500 461 -499
rect 940 -500 941 -499
rect 996 -500 997 -499
rect 1038 -500 1039 -499
rect 100 -502 101 -501
rect 128 -502 129 -501
rect 149 -502 150 -501
rect 170 -502 171 -501
rect 177 -502 178 -501
rect 254 -502 255 -501
rect 289 -502 290 -501
rect 320 -502 321 -501
rect 331 -502 332 -501
rect 373 -502 374 -501
rect 429 -502 430 -501
rect 509 -502 510 -501
rect 611 -502 612 -501
rect 856 -502 857 -501
rect 884 -502 885 -501
rect 1066 -502 1067 -501
rect 44 -504 45 -503
rect 331 -504 332 -503
rect 443 -504 444 -503
rect 509 -504 510 -503
rect 548 -504 549 -503
rect 611 -504 612 -503
rect 632 -504 633 -503
rect 653 -504 654 -503
rect 660 -504 661 -503
rect 940 -504 941 -503
rect 1003 -504 1004 -503
rect 1052 -504 1053 -503
rect 44 -506 45 -505
rect 317 -506 318 -505
rect 387 -506 388 -505
rect 1052 -506 1053 -505
rect 110 -508 111 -507
rect 177 -508 178 -507
rect 191 -508 192 -507
rect 324 -508 325 -507
rect 471 -508 472 -507
rect 569 -508 570 -507
rect 604 -508 605 -507
rect 653 -508 654 -507
rect 723 -508 724 -507
rect 905 -508 906 -507
rect 1010 -508 1011 -507
rect 1031 -508 1032 -507
rect 33 -510 34 -509
rect 604 -510 605 -509
rect 730 -510 731 -509
rect 1024 -510 1025 -509
rect 1031 -510 1032 -509
rect 1080 -510 1081 -509
rect 114 -512 115 -511
rect 394 -512 395 -511
rect 478 -512 479 -511
rect 492 -512 493 -511
rect 502 -512 503 -511
rect 723 -512 724 -511
rect 754 -512 755 -511
rect 814 -512 815 -511
rect 828 -512 829 -511
rect 842 -512 843 -511
rect 849 -512 850 -511
rect 884 -512 885 -511
rect 898 -512 899 -511
rect 905 -512 906 -511
rect 1017 -512 1018 -511
rect 1073 -512 1074 -511
rect 1080 -512 1081 -511
rect 1087 -512 1088 -511
rect 128 -514 129 -513
rect 408 -514 409 -513
rect 485 -514 486 -513
rect 572 -514 573 -513
rect 597 -514 598 -513
rect 1087 -514 1088 -513
rect 152 -516 153 -515
rect 569 -516 570 -515
rect 597 -516 598 -515
rect 877 -516 878 -515
rect 926 -516 927 -515
rect 1073 -516 1074 -515
rect 163 -518 164 -517
rect 471 -518 472 -517
rect 492 -518 493 -517
rect 628 -518 629 -517
rect 765 -518 766 -517
rect 1094 -518 1095 -517
rect 191 -520 192 -519
rect 695 -520 696 -519
rect 779 -520 780 -519
rect 828 -520 829 -519
rect 835 -520 836 -519
rect 947 -520 948 -519
rect 247 -522 248 -521
rect 404 -522 405 -521
rect 422 -522 423 -521
rect 835 -522 836 -521
rect 877 -522 878 -521
rect 912 -522 913 -521
rect 121 -524 122 -523
rect 422 -524 423 -523
rect 551 -524 552 -523
rect 926 -524 927 -523
rect 268 -526 269 -525
rect 443 -526 444 -525
rect 688 -526 689 -525
rect 765 -526 766 -525
rect 786 -526 787 -525
rect 814 -526 815 -525
rect 821 -526 822 -525
rect 898 -526 899 -525
rect 268 -528 269 -527
rect 282 -528 283 -527
rect 317 -528 318 -527
rect 359 -528 360 -527
rect 667 -528 668 -527
rect 688 -528 689 -527
rect 716 -528 717 -527
rect 779 -528 780 -527
rect 793 -528 794 -527
rect 849 -528 850 -527
rect 891 -528 892 -527
rect 912 -528 913 -527
rect 138 -530 139 -529
rect 359 -530 360 -529
rect 639 -530 640 -529
rect 667 -530 668 -529
rect 681 -530 682 -529
rect 716 -530 717 -529
rect 744 -530 745 -529
rect 786 -530 787 -529
rect 800 -530 801 -529
rect 821 -530 822 -529
rect 863 -530 864 -529
rect 891 -530 892 -529
rect 233 -532 234 -531
rect 282 -532 283 -531
rect 355 -532 356 -531
rect 793 -532 794 -531
rect 807 -532 808 -531
rect 1038 -532 1039 -531
rect 51 -534 52 -533
rect 233 -534 234 -533
rect 408 -534 409 -533
rect 800 -534 801 -533
rect 863 -534 864 -533
rect 954 -534 955 -533
rect 51 -536 52 -535
rect 338 -536 339 -535
rect 548 -536 549 -535
rect 681 -536 682 -535
rect 744 -536 745 -535
rect 758 -536 759 -535
rect 772 -536 773 -535
rect 807 -536 808 -535
rect 933 -536 934 -535
rect 954 -536 955 -535
rect 338 -538 339 -537
rect 390 -538 391 -537
rect 625 -538 626 -537
rect 639 -538 640 -537
rect 702 -538 703 -537
rect 772 -538 773 -537
rect 919 -538 920 -537
rect 933 -538 934 -537
rect 562 -540 563 -539
rect 919 -540 920 -539
rect 674 -542 675 -541
rect 702 -542 703 -541
rect 709 -542 710 -541
rect 758 -542 759 -541
rect 646 -544 647 -543
rect 674 -544 675 -543
rect 709 -544 710 -543
rect 870 -544 871 -543
rect 618 -546 619 -545
rect 646 -546 647 -545
rect 576 -548 577 -547
rect 618 -548 619 -547
rect 65 -550 66 -549
rect 576 -550 577 -549
rect 65 -552 66 -551
rect 198 -552 199 -551
rect 198 -554 199 -553
rect 464 -554 465 -553
rect 215 -556 216 -555
rect 464 -556 465 -555
rect 194 -558 195 -557
rect 215 -558 216 -557
rect 2 -569 3 -568
rect 509 -569 510 -568
rect 534 -569 535 -568
rect 541 -569 542 -568
rect 548 -569 549 -568
rect 870 -569 871 -568
rect 1059 -569 1060 -568
rect 1108 -569 1109 -568
rect 9 -571 10 -570
rect 72 -571 73 -570
rect 82 -571 83 -570
rect 709 -571 710 -570
rect 712 -571 713 -570
rect 898 -571 899 -570
rect 1087 -571 1088 -570
rect 1129 -571 1130 -570
rect 9 -573 10 -572
rect 380 -573 381 -572
rect 408 -573 409 -572
rect 835 -573 836 -572
rect 842 -573 843 -572
rect 898 -573 899 -572
rect 1024 -573 1025 -572
rect 1087 -573 1088 -572
rect 1101 -573 1102 -572
rect 1136 -573 1137 -572
rect 16 -575 17 -574
rect 870 -575 871 -574
rect 975 -575 976 -574
rect 1024 -575 1025 -574
rect 16 -577 17 -576
rect 86 -577 87 -576
rect 121 -577 122 -576
rect 562 -577 563 -576
rect 569 -577 570 -576
rect 1038 -577 1039 -576
rect 23 -579 24 -578
rect 541 -579 542 -578
rect 548 -579 549 -578
rect 1059 -579 1060 -578
rect 23 -581 24 -580
rect 418 -581 419 -580
rect 443 -581 444 -580
rect 572 -581 573 -580
rect 600 -581 601 -580
rect 884 -581 885 -580
rect 919 -581 920 -580
rect 1038 -581 1039 -580
rect 30 -583 31 -582
rect 79 -583 80 -582
rect 86 -583 87 -582
rect 296 -583 297 -582
rect 338 -583 339 -582
rect 387 -583 388 -582
rect 464 -583 465 -582
rect 691 -583 692 -582
rect 733 -583 734 -582
rect 744 -583 745 -582
rect 751 -583 752 -582
rect 919 -583 920 -582
rect 968 -583 969 -582
rect 975 -583 976 -582
rect 30 -585 31 -584
rect 261 -585 262 -584
rect 268 -585 269 -584
rect 352 -585 353 -584
rect 380 -585 381 -584
rect 492 -585 493 -584
rect 506 -585 507 -584
rect 1101 -585 1102 -584
rect 33 -587 34 -586
rect 411 -587 412 -586
rect 471 -587 472 -586
rect 597 -587 598 -586
rect 604 -587 605 -586
rect 1066 -587 1067 -586
rect 37 -589 38 -588
rect 187 -589 188 -588
rect 191 -589 192 -588
rect 226 -589 227 -588
rect 254 -589 255 -588
rect 502 -589 503 -588
rect 513 -589 514 -588
rect 562 -589 563 -588
rect 604 -589 605 -588
rect 961 -589 962 -588
rect 1003 -589 1004 -588
rect 1066 -589 1067 -588
rect 37 -591 38 -590
rect 100 -591 101 -590
rect 107 -591 108 -590
rect 261 -591 262 -590
rect 275 -591 276 -590
rect 355 -591 356 -590
rect 436 -591 437 -590
rect 471 -591 472 -590
rect 478 -591 479 -590
rect 513 -591 514 -590
rect 551 -591 552 -590
rect 856 -591 857 -590
rect 877 -591 878 -590
rect 961 -591 962 -590
rect 44 -593 45 -592
rect 464 -593 465 -592
rect 555 -593 556 -592
rect 569 -593 570 -592
rect 625 -593 626 -592
rect 681 -593 682 -592
rect 688 -593 689 -592
rect 744 -593 745 -592
rect 751 -593 752 -592
rect 758 -593 759 -592
rect 761 -593 762 -592
rect 1010 -593 1011 -592
rect 44 -595 45 -594
rect 93 -595 94 -594
rect 107 -595 108 -594
rect 117 -595 118 -594
rect 121 -595 122 -594
rect 201 -595 202 -594
rect 205 -595 206 -594
rect 397 -595 398 -594
rect 415 -595 416 -594
rect 436 -595 437 -594
rect 555 -595 556 -594
rect 639 -595 640 -594
rect 656 -595 657 -594
rect 1080 -595 1081 -594
rect 54 -597 55 -596
rect 800 -597 801 -596
rect 807 -597 808 -596
rect 877 -597 878 -596
rect 926 -597 927 -596
rect 968 -597 969 -596
rect 982 -597 983 -596
rect 1010 -597 1011 -596
rect 1017 -597 1018 -596
rect 1080 -597 1081 -596
rect 65 -599 66 -598
rect 506 -599 507 -598
rect 611 -599 612 -598
rect 639 -599 640 -598
rect 660 -599 661 -598
rect 1073 -599 1074 -598
rect 68 -601 69 -600
rect 457 -601 458 -600
rect 628 -601 629 -600
rect 730 -601 731 -600
rect 765 -601 766 -600
rect 856 -601 857 -600
rect 926 -601 927 -600
rect 947 -601 948 -600
rect 954 -601 955 -600
rect 1003 -601 1004 -600
rect 1045 -601 1046 -600
rect 1073 -601 1074 -600
rect 72 -603 73 -602
rect 373 -603 374 -602
rect 450 -603 451 -602
rect 457 -603 458 -602
rect 632 -603 633 -602
rect 681 -603 682 -602
rect 723 -603 724 -602
rect 807 -603 808 -602
rect 821 -603 822 -602
rect 842 -603 843 -602
rect 849 -603 850 -602
rect 954 -603 955 -602
rect 989 -603 990 -602
rect 1045 -603 1046 -602
rect 79 -605 80 -604
rect 835 -605 836 -604
rect 905 -605 906 -604
rect 947 -605 948 -604
rect 989 -605 990 -604
rect 1052 -605 1053 -604
rect 75 -607 76 -606
rect 905 -607 906 -606
rect 933 -607 934 -606
rect 982 -607 983 -606
rect 996 -607 997 -606
rect 1052 -607 1053 -606
rect 93 -609 94 -608
rect 607 -609 608 -608
rect 611 -609 612 -608
rect 632 -609 633 -608
rect 646 -609 647 -608
rect 660 -609 661 -608
rect 765 -609 766 -608
rect 779 -609 780 -608
rect 793 -609 794 -608
rect 884 -609 885 -608
rect 940 -609 941 -608
rect 1017 -609 1018 -608
rect 114 -611 115 -610
rect 450 -611 451 -610
rect 485 -611 486 -610
rect 646 -611 647 -610
rect 674 -611 675 -610
rect 779 -611 780 -610
rect 800 -611 801 -610
rect 1094 -611 1095 -610
rect 128 -613 129 -612
rect 446 -613 447 -612
rect 537 -613 538 -612
rect 723 -613 724 -612
rect 772 -613 773 -612
rect 821 -613 822 -612
rect 863 -613 864 -612
rect 996 -613 997 -612
rect 1031 -613 1032 -612
rect 1094 -613 1095 -612
rect 149 -615 150 -614
rect 408 -615 409 -614
rect 663 -615 664 -614
rect 1031 -615 1032 -614
rect 152 -617 153 -616
rect 296 -617 297 -616
rect 331 -617 332 -616
rect 352 -617 353 -616
rect 373 -617 374 -616
rect 481 -617 482 -616
rect 667 -617 668 -616
rect 674 -617 675 -616
rect 695 -617 696 -616
rect 793 -617 794 -616
rect 814 -617 815 -616
rect 849 -617 850 -616
rect 166 -619 167 -618
rect 912 -619 913 -618
rect 170 -621 171 -620
rect 198 -621 199 -620
rect 212 -621 213 -620
rect 366 -621 367 -620
rect 390 -621 391 -620
rect 863 -621 864 -620
rect 891 -621 892 -620
rect 912 -621 913 -620
rect 51 -623 52 -622
rect 366 -623 367 -622
rect 583 -623 584 -622
rect 667 -623 668 -622
rect 695 -623 696 -622
rect 758 -623 759 -622
rect 828 -623 829 -622
rect 891 -623 892 -622
rect 170 -625 171 -624
rect 247 -625 248 -624
rect 289 -625 290 -624
rect 485 -625 486 -624
rect 583 -625 584 -624
rect 618 -625 619 -624
rect 716 -625 717 -624
rect 772 -625 773 -624
rect 786 -625 787 -624
rect 828 -625 829 -624
rect 177 -627 178 -626
rect 226 -627 227 -626
rect 233 -627 234 -626
rect 254 -627 255 -626
rect 289 -627 290 -626
rect 607 -627 608 -626
rect 653 -627 654 -626
rect 716 -627 717 -626
rect 737 -627 738 -626
rect 814 -627 815 -626
rect 100 -629 101 -628
rect 737 -629 738 -628
rect 177 -631 178 -630
rect 184 -631 185 -630
rect 212 -631 213 -630
rect 317 -631 318 -630
rect 341 -631 342 -630
rect 940 -631 941 -630
rect 142 -633 143 -632
rect 317 -633 318 -632
rect 345 -633 346 -632
rect 394 -633 395 -632
rect 422 -633 423 -632
rect 653 -633 654 -632
rect 58 -635 59 -634
rect 345 -635 346 -634
rect 348 -635 349 -634
rect 492 -635 493 -634
rect 576 -635 577 -634
rect 618 -635 619 -634
rect 58 -637 59 -636
rect 240 -637 241 -636
rect 247 -637 248 -636
rect 282 -637 283 -636
rect 359 -637 360 -636
rect 786 -637 787 -636
rect 135 -639 136 -638
rect 240 -639 241 -638
rect 282 -639 283 -638
rect 320 -639 321 -638
rect 359 -639 360 -638
rect 401 -639 402 -638
rect 422 -639 423 -638
rect 614 -639 615 -638
rect 135 -641 136 -640
rect 163 -641 164 -640
rect 184 -641 185 -640
rect 268 -641 269 -640
rect 401 -641 402 -640
rect 429 -641 430 -640
rect 527 -641 528 -640
rect 576 -641 577 -640
rect 142 -643 143 -642
rect 590 -643 591 -642
rect 163 -645 164 -644
rect 205 -645 206 -644
rect 219 -645 220 -644
rect 275 -645 276 -644
rect 324 -645 325 -644
rect 429 -645 430 -644
rect 499 -645 500 -644
rect 527 -645 528 -644
rect 156 -647 157 -646
rect 219 -647 220 -646
rect 310 -647 311 -646
rect 324 -647 325 -646
rect 520 -647 521 -646
rect 590 -647 591 -646
rect 310 -649 311 -648
rect 331 -649 332 -648
rect 16 -660 17 -659
rect 128 -660 129 -659
rect 149 -660 150 -659
rect 233 -660 234 -659
rect 254 -660 255 -659
rect 415 -660 416 -659
rect 425 -660 426 -659
rect 607 -660 608 -659
rect 611 -660 612 -659
rect 632 -660 633 -659
rect 691 -660 692 -659
rect 975 -660 976 -659
rect 1003 -660 1004 -659
rect 1006 -660 1007 -659
rect 1038 -660 1039 -659
rect 1041 -660 1042 -659
rect 1059 -660 1060 -659
rect 1150 -660 1151 -659
rect 1178 -660 1179 -659
rect 1185 -660 1186 -659
rect 16 -662 17 -661
rect 184 -662 185 -661
rect 187 -662 188 -661
rect 236 -662 237 -661
rect 254 -662 255 -661
rect 268 -662 269 -661
rect 324 -662 325 -661
rect 338 -662 339 -661
rect 408 -662 409 -661
rect 793 -662 794 -661
rect 807 -662 808 -661
rect 810 -662 811 -661
rect 933 -662 934 -661
rect 1017 -662 1018 -661
rect 1038 -662 1039 -661
rect 1115 -662 1116 -661
rect 23 -664 24 -663
rect 422 -664 423 -663
rect 439 -664 440 -663
rect 635 -664 636 -663
rect 747 -664 748 -663
rect 779 -664 780 -663
rect 807 -664 808 -663
rect 814 -664 815 -663
rect 933 -664 934 -663
rect 947 -664 948 -663
rect 975 -664 976 -663
rect 1024 -664 1025 -663
rect 1045 -664 1046 -663
rect 1059 -664 1060 -663
rect 1087 -664 1088 -663
rect 1115 -664 1116 -663
rect 30 -666 31 -665
rect 478 -666 479 -665
rect 481 -666 482 -665
rect 919 -666 920 -665
rect 947 -666 948 -665
rect 982 -666 983 -665
rect 996 -666 997 -665
rect 1017 -666 1018 -665
rect 1087 -666 1088 -665
rect 1129 -666 1130 -665
rect 37 -668 38 -667
rect 131 -668 132 -667
rect 142 -668 143 -667
rect 338 -668 339 -667
rect 345 -668 346 -667
rect 478 -668 479 -667
rect 513 -668 514 -667
rect 660 -668 661 -667
rect 695 -668 696 -667
rect 779 -668 780 -667
rect 814 -668 815 -667
rect 877 -668 878 -667
rect 898 -668 899 -667
rect 919 -668 920 -667
rect 968 -668 969 -667
rect 996 -668 997 -667
rect 1003 -668 1004 -667
rect 1052 -668 1053 -667
rect 1090 -668 1091 -667
rect 1171 -668 1172 -667
rect 37 -670 38 -669
rect 121 -670 122 -669
rect 142 -670 143 -669
rect 191 -670 192 -669
rect 205 -670 206 -669
rect 397 -670 398 -669
rect 443 -670 444 -669
rect 1024 -670 1025 -669
rect 1031 -670 1032 -669
rect 1052 -670 1053 -669
rect 1101 -670 1102 -669
rect 1129 -670 1130 -669
rect 44 -672 45 -671
rect 117 -672 118 -671
rect 159 -672 160 -671
rect 597 -672 598 -671
rect 604 -672 605 -671
rect 989 -672 990 -671
rect 1010 -672 1011 -671
rect 1045 -672 1046 -671
rect 1080 -672 1081 -671
rect 1101 -672 1102 -671
rect 1108 -672 1109 -671
rect 1143 -672 1144 -671
rect 44 -674 45 -673
rect 198 -674 199 -673
rect 208 -674 209 -673
rect 212 -674 213 -673
rect 233 -674 234 -673
rect 261 -674 262 -673
rect 268 -674 269 -673
rect 691 -674 692 -673
rect 758 -674 759 -673
rect 772 -674 773 -673
rect 842 -674 843 -673
rect 898 -674 899 -673
rect 940 -674 941 -673
rect 968 -674 969 -673
rect 1073 -674 1074 -673
rect 1080 -674 1081 -673
rect 1108 -674 1109 -673
rect 1136 -674 1137 -673
rect 51 -676 52 -675
rect 191 -676 192 -675
rect 198 -676 199 -675
rect 303 -676 304 -675
rect 324 -676 325 -675
rect 373 -676 374 -675
rect 380 -676 381 -675
rect 513 -676 514 -675
rect 523 -676 524 -675
rect 1164 -676 1165 -675
rect 54 -678 55 -677
rect 65 -678 66 -677
rect 72 -678 73 -677
rect 446 -678 447 -677
rect 464 -678 465 -677
rect 474 -678 475 -677
rect 502 -678 503 -677
rect 842 -678 843 -677
rect 940 -678 941 -677
rect 954 -678 955 -677
rect 961 -678 962 -677
rect 989 -678 990 -677
rect 1073 -678 1074 -677
rect 1094 -678 1095 -677
rect 1122 -678 1123 -677
rect 1136 -678 1137 -677
rect 58 -680 59 -679
rect 261 -680 262 -679
rect 303 -680 304 -679
rect 450 -680 451 -679
rect 464 -680 465 -679
rect 709 -680 710 -679
rect 905 -680 906 -679
rect 954 -680 955 -679
rect 58 -682 59 -681
rect 352 -682 353 -681
rect 366 -682 367 -681
rect 443 -682 444 -681
rect 450 -682 451 -681
rect 471 -682 472 -681
rect 516 -682 517 -681
rect 1122 -682 1123 -681
rect 65 -684 66 -683
rect 523 -684 524 -683
rect 551 -684 552 -683
rect 856 -684 857 -683
rect 884 -684 885 -683
rect 905 -684 906 -683
rect 912 -684 913 -683
rect 961 -684 962 -683
rect 72 -686 73 -685
rect 212 -686 213 -685
rect 317 -686 318 -685
rect 352 -686 353 -685
rect 366 -686 367 -685
rect 520 -686 521 -685
rect 551 -686 552 -685
rect 583 -686 584 -685
rect 597 -686 598 -685
rect 835 -686 836 -685
rect 891 -686 892 -685
rect 912 -686 913 -685
rect 79 -688 80 -687
rect 96 -688 97 -687
rect 100 -688 101 -687
rect 219 -688 220 -687
rect 310 -688 311 -687
rect 317 -688 318 -687
rect 345 -688 346 -687
rect 436 -688 437 -687
rect 499 -688 500 -687
rect 884 -688 885 -687
rect 79 -690 80 -689
rect 107 -690 108 -689
rect 114 -690 115 -689
rect 135 -690 136 -689
rect 152 -690 153 -689
rect 373 -690 374 -689
rect 380 -690 381 -689
rect 418 -690 419 -689
rect 485 -690 486 -689
rect 499 -690 500 -689
rect 569 -690 570 -689
rect 583 -690 584 -689
rect 604 -690 605 -689
rect 863 -690 864 -689
rect 870 -690 871 -689
rect 891 -690 892 -689
rect 82 -692 83 -691
rect 548 -692 549 -691
rect 576 -692 577 -691
rect 653 -692 654 -691
rect 660 -692 661 -691
rect 716 -692 717 -691
rect 765 -692 766 -691
rect 863 -692 864 -691
rect 86 -694 87 -693
rect 149 -694 150 -693
rect 156 -694 157 -693
rect 1010 -694 1011 -693
rect 89 -696 90 -695
rect 205 -696 206 -695
rect 219 -696 220 -695
rect 275 -696 276 -695
rect 506 -696 507 -695
rect 576 -696 577 -695
rect 614 -696 615 -695
rect 926 -696 927 -695
rect 93 -698 94 -697
rect 107 -698 108 -697
rect 135 -698 136 -697
rect 835 -698 836 -697
rect 93 -700 94 -699
rect 163 -700 164 -699
rect 184 -700 185 -699
rect 331 -700 332 -699
rect 506 -700 507 -699
rect 800 -700 801 -699
rect 821 -700 822 -699
rect 856 -700 857 -699
rect 103 -702 104 -701
rect 555 -702 556 -701
rect 646 -702 647 -701
rect 709 -702 710 -701
rect 716 -702 717 -701
rect 793 -702 794 -701
rect 800 -702 801 -701
rect 828 -702 829 -701
rect 156 -704 157 -703
rect 170 -704 171 -703
rect 240 -704 241 -703
rect 485 -704 486 -703
rect 534 -704 535 -703
rect 569 -704 570 -703
rect 646 -704 647 -703
rect 681 -704 682 -703
rect 688 -704 689 -703
rect 695 -704 696 -703
rect 702 -704 703 -703
rect 772 -704 773 -703
rect 163 -706 164 -705
rect 247 -706 248 -705
rect 275 -706 276 -705
rect 282 -706 283 -705
rect 467 -706 468 -705
rect 821 -706 822 -705
rect 170 -708 171 -707
rect 359 -708 360 -707
rect 527 -708 528 -707
rect 534 -708 535 -707
rect 541 -708 542 -707
rect 555 -708 556 -707
rect 667 -708 668 -707
rect 681 -708 682 -707
rect 688 -708 689 -707
rect 982 -708 983 -707
rect 1041 -708 1042 -707
rect 1094 -708 1095 -707
rect 240 -710 241 -709
rect 296 -710 297 -709
rect 429 -710 430 -709
rect 541 -710 542 -709
rect 639 -710 640 -709
rect 667 -710 668 -709
rect 730 -710 731 -709
rect 926 -710 927 -709
rect 282 -712 283 -711
rect 394 -712 395 -711
rect 401 -712 402 -711
rect 429 -712 430 -711
rect 527 -712 528 -711
rect 618 -712 619 -711
rect 639 -712 640 -711
rect 702 -712 703 -711
rect 730 -712 731 -711
rect 786 -712 787 -711
rect 33 -714 34 -713
rect 394 -714 395 -713
rect 411 -714 412 -713
rect 786 -714 787 -713
rect 289 -716 290 -715
rect 296 -716 297 -715
rect 562 -716 563 -715
rect 618 -716 619 -715
rect 744 -716 745 -715
rect 765 -716 766 -715
rect 289 -718 290 -717
rect 492 -718 493 -717
rect 562 -718 563 -717
rect 590 -718 591 -717
rect 744 -718 745 -717
rect 870 -718 871 -717
rect 341 -720 342 -719
rect 590 -720 591 -719
rect 751 -720 752 -719
rect 828 -720 829 -719
rect 492 -722 493 -721
rect 723 -722 724 -721
rect 625 -724 626 -723
rect 751 -724 752 -723
rect 625 -726 626 -725
rect 1111 -726 1112 -725
rect 674 -728 675 -727
rect 723 -728 724 -727
rect 656 -730 657 -729
rect 674 -730 675 -729
rect 9 -741 10 -740
rect 138 -741 139 -740
rect 149 -741 150 -740
rect 583 -741 584 -740
rect 600 -741 601 -740
rect 940 -741 941 -740
rect 1038 -741 1039 -740
rect 1087 -741 1088 -740
rect 1108 -741 1109 -740
rect 1136 -741 1137 -740
rect 1143 -741 1144 -740
rect 1192 -741 1193 -740
rect 9 -743 10 -742
rect 79 -743 80 -742
rect 86 -743 87 -742
rect 131 -743 132 -742
rect 163 -743 164 -742
rect 362 -743 363 -742
rect 373 -743 374 -742
rect 383 -743 384 -742
rect 404 -743 405 -742
rect 499 -743 500 -742
rect 502 -743 503 -742
rect 527 -743 528 -742
rect 583 -743 584 -742
rect 747 -743 748 -742
rect 782 -743 783 -742
rect 1003 -743 1004 -742
rect 1031 -743 1032 -742
rect 1038 -743 1039 -742
rect 1052 -743 1053 -742
rect 1108 -743 1109 -742
rect 1122 -743 1123 -742
rect 1178 -743 1179 -742
rect 1185 -743 1186 -742
rect 1213 -743 1214 -742
rect 16 -745 17 -744
rect 338 -745 339 -744
rect 359 -745 360 -744
rect 1052 -745 1053 -744
rect 1059 -745 1060 -744
rect 1122 -745 1123 -744
rect 1129 -745 1130 -744
rect 1185 -745 1186 -744
rect 16 -747 17 -746
rect 366 -747 367 -746
rect 373 -747 374 -746
rect 387 -747 388 -746
rect 408 -747 409 -746
rect 625 -747 626 -746
rect 639 -747 640 -746
rect 817 -747 818 -746
rect 821 -747 822 -746
rect 852 -747 853 -746
rect 884 -747 885 -746
rect 1003 -747 1004 -746
rect 1059 -747 1060 -746
rect 1090 -747 1091 -746
rect 1101 -747 1102 -746
rect 1143 -747 1144 -746
rect 1150 -747 1151 -746
rect 1160 -747 1161 -746
rect 1164 -747 1165 -746
rect 1199 -747 1200 -746
rect 23 -749 24 -748
rect 401 -749 402 -748
rect 411 -749 412 -748
rect 415 -749 416 -748
rect 439 -749 440 -748
rect 471 -749 472 -748
rect 495 -749 496 -748
rect 947 -749 948 -748
rect 968 -749 969 -748
rect 1031 -749 1032 -748
rect 1080 -749 1081 -748
rect 1136 -749 1137 -748
rect 1171 -749 1172 -748
rect 1220 -749 1221 -748
rect 23 -751 24 -750
rect 345 -751 346 -750
rect 387 -751 388 -750
rect 569 -751 570 -750
rect 572 -751 573 -750
rect 1164 -751 1165 -750
rect 30 -753 31 -752
rect 170 -753 171 -752
rect 173 -753 174 -752
rect 205 -753 206 -752
rect 212 -753 213 -752
rect 425 -753 426 -752
rect 464 -753 465 -752
rect 478 -753 479 -752
rect 513 -753 514 -752
rect 635 -753 636 -752
rect 642 -753 643 -752
rect 863 -753 864 -752
rect 926 -753 927 -752
rect 940 -753 941 -752
rect 947 -753 948 -752
rect 954 -753 955 -752
rect 989 -753 990 -752
rect 1080 -753 1081 -752
rect 1115 -753 1116 -752
rect 1150 -753 1151 -752
rect 37 -755 38 -754
rect 124 -755 125 -754
rect 177 -755 178 -754
rect 184 -755 185 -754
rect 187 -755 188 -754
rect 541 -755 542 -754
rect 625 -755 626 -754
rect 877 -755 878 -754
rect 954 -755 955 -754
rect 1157 -755 1158 -754
rect 37 -757 38 -756
rect 117 -757 118 -756
rect 156 -757 157 -756
rect 177 -757 178 -756
rect 191 -757 192 -756
rect 254 -757 255 -756
rect 331 -757 332 -756
rect 436 -757 437 -756
rect 485 -757 486 -756
rect 513 -757 514 -756
rect 520 -757 521 -756
rect 968 -757 969 -756
rect 982 -757 983 -756
rect 989 -757 990 -756
rect 996 -757 997 -756
rect 1087 -757 1088 -756
rect 58 -759 59 -758
rect 345 -759 346 -758
rect 366 -759 367 -758
rect 520 -759 521 -758
rect 523 -759 524 -758
rect 660 -759 661 -758
rect 663 -759 664 -758
rect 1129 -759 1130 -758
rect 58 -761 59 -760
rect 93 -761 94 -760
rect 100 -761 101 -760
rect 212 -761 213 -760
rect 338 -761 339 -760
rect 597 -761 598 -760
rect 604 -761 605 -760
rect 1157 -761 1158 -760
rect 65 -763 66 -762
rect 331 -763 332 -762
rect 380 -763 381 -762
rect 660 -763 661 -762
rect 688 -763 689 -762
rect 898 -763 899 -762
rect 933 -763 934 -762
rect 982 -763 983 -762
rect 996 -763 997 -762
rect 1024 -763 1025 -762
rect 1073 -763 1074 -762
rect 1171 -763 1172 -762
rect 44 -765 45 -764
rect 380 -765 381 -764
rect 394 -765 395 -764
rect 884 -765 885 -764
rect 1010 -765 1011 -764
rect 1115 -765 1116 -764
rect 44 -767 45 -766
rect 268 -767 269 -766
rect 341 -767 342 -766
rect 1024 -767 1025 -766
rect 1073 -767 1074 -766
rect 1094 -767 1095 -766
rect 65 -769 66 -768
rect 506 -769 507 -768
rect 527 -769 528 -768
rect 534 -769 535 -768
rect 541 -769 542 -768
rect 555 -769 556 -768
rect 565 -769 566 -768
rect 933 -769 934 -768
rect 1017 -769 1018 -768
rect 1094 -769 1095 -768
rect 79 -771 80 -770
rect 425 -771 426 -770
rect 499 -771 500 -770
rect 534 -771 535 -770
rect 569 -771 570 -770
rect 1010 -771 1011 -770
rect 1017 -771 1018 -770
rect 1066 -771 1067 -770
rect 86 -773 87 -772
rect 317 -773 318 -772
rect 394 -773 395 -772
rect 429 -773 430 -772
rect 506 -773 507 -772
rect 576 -773 577 -772
rect 590 -773 591 -772
rect 604 -773 605 -772
rect 688 -773 689 -772
rect 695 -773 696 -772
rect 698 -773 699 -772
rect 1101 -773 1102 -772
rect 93 -775 94 -774
rect 240 -775 241 -774
rect 268 -775 269 -774
rect 310 -775 311 -774
rect 317 -775 318 -774
rect 352 -775 353 -774
rect 415 -775 416 -774
rect 642 -775 643 -774
rect 716 -775 717 -774
rect 856 -775 857 -774
rect 870 -775 871 -774
rect 877 -775 878 -774
rect 100 -777 101 -776
rect 135 -777 136 -776
rect 138 -777 139 -776
rect 156 -777 157 -776
rect 163 -777 164 -776
rect 254 -777 255 -776
rect 429 -777 430 -776
rect 891 -777 892 -776
rect 114 -779 115 -778
rect 121 -779 122 -778
rect 135 -779 136 -778
rect 289 -779 290 -778
rect 457 -779 458 -778
rect 576 -779 577 -778
rect 590 -779 591 -778
rect 618 -779 619 -778
rect 744 -779 745 -778
rect 975 -779 976 -778
rect 170 -781 171 -780
rect 240 -781 241 -780
rect 247 -781 248 -780
rect 310 -781 311 -780
rect 443 -781 444 -780
rect 457 -781 458 -780
rect 485 -781 486 -780
rect 695 -781 696 -780
rect 786 -781 787 -780
rect 898 -781 899 -780
rect 191 -783 192 -782
rect 296 -783 297 -782
rect 443 -783 444 -782
rect 450 -783 451 -782
rect 492 -783 493 -782
rect 716 -783 717 -782
rect 786 -783 787 -782
rect 807 -783 808 -782
rect 842 -783 843 -782
rect 926 -783 927 -782
rect 226 -785 227 -784
rect 247 -785 248 -784
rect 289 -785 290 -784
rect 352 -785 353 -784
rect 548 -785 549 -784
rect 744 -785 745 -784
rect 779 -785 780 -784
rect 807 -785 808 -784
rect 835 -785 836 -784
rect 842 -785 843 -784
rect 849 -785 850 -784
rect 863 -785 864 -784
rect 891 -785 892 -784
rect 905 -785 906 -784
rect 128 -787 129 -786
rect 226 -787 227 -786
rect 296 -787 297 -786
rect 611 -787 612 -786
rect 656 -787 657 -786
rect 975 -787 976 -786
rect 303 -789 304 -788
rect 450 -789 451 -788
rect 548 -789 549 -788
rect 562 -789 563 -788
rect 597 -789 598 -788
rect 751 -789 752 -788
rect 779 -789 780 -788
rect 870 -789 871 -788
rect 198 -791 199 -790
rect 303 -791 304 -790
rect 555 -791 556 -790
rect 1066 -791 1067 -790
rect 107 -793 108 -792
rect 198 -793 199 -792
rect 562 -793 563 -792
rect 730 -793 731 -792
rect 751 -793 752 -792
rect 828 -793 829 -792
rect 849 -793 850 -792
rect 1206 -793 1207 -792
rect 107 -795 108 -794
rect 219 -795 220 -794
rect 474 -795 475 -794
rect 828 -795 829 -794
rect 856 -795 857 -794
rect 919 -795 920 -794
rect 219 -797 220 -796
rect 653 -797 654 -796
rect 793 -797 794 -796
rect 821 -797 822 -796
rect 912 -797 913 -796
rect 919 -797 920 -796
rect 611 -799 612 -798
rect 667 -799 668 -798
rect 772 -799 773 -798
rect 793 -799 794 -798
rect 800 -799 801 -798
rect 905 -799 906 -798
rect 912 -799 913 -798
rect 961 -799 962 -798
rect 478 -801 479 -800
rect 772 -801 773 -800
rect 814 -801 815 -800
rect 835 -801 836 -800
rect 632 -803 633 -802
rect 961 -803 962 -802
rect 632 -805 633 -804
rect 681 -805 682 -804
rect 758 -805 759 -804
rect 800 -805 801 -804
rect 51 -807 52 -806
rect 681 -807 682 -806
rect 51 -809 52 -808
rect 282 -809 283 -808
rect 621 -809 622 -808
rect 758 -809 759 -808
rect 233 -811 234 -810
rect 282 -811 283 -810
rect 667 -811 668 -810
rect 709 -811 710 -810
rect 233 -813 234 -812
rect 275 -813 276 -812
rect 646 -813 647 -812
rect 709 -813 710 -812
rect 261 -815 262 -814
rect 275 -815 276 -814
rect 646 -815 647 -814
rect 674 -815 675 -814
rect 674 -817 675 -816
rect 723 -817 724 -816
rect 723 -819 724 -818
rect 730 -819 731 -818
rect 19 -830 20 -829
rect 313 -830 314 -829
rect 355 -830 356 -829
rect 1003 -830 1004 -829
rect 30 -832 31 -831
rect 117 -832 118 -831
rect 121 -832 122 -831
rect 1101 -832 1102 -831
rect 33 -834 34 -833
rect 170 -834 171 -833
rect 198 -834 199 -833
rect 499 -834 500 -833
rect 523 -834 524 -833
rect 590 -834 591 -833
rect 618 -834 619 -833
rect 905 -834 906 -833
rect 996 -834 997 -833
rect 999 -834 1000 -833
rect 1003 -834 1004 -833
rect 1038 -834 1039 -833
rect 44 -836 45 -835
rect 569 -836 570 -835
rect 590 -836 591 -835
rect 632 -836 633 -835
rect 639 -836 640 -835
rect 702 -836 703 -835
rect 726 -836 727 -835
rect 1066 -836 1067 -835
rect 44 -838 45 -837
rect 289 -838 290 -837
rect 359 -838 360 -837
rect 383 -838 384 -837
rect 387 -838 388 -837
rect 478 -838 479 -837
rect 485 -838 486 -837
rect 520 -838 521 -837
rect 555 -838 556 -837
rect 611 -838 612 -837
rect 656 -838 657 -837
rect 730 -838 731 -837
rect 758 -838 759 -837
rect 849 -838 850 -837
rect 905 -838 906 -837
rect 989 -838 990 -837
rect 996 -838 997 -837
rect 1010 -838 1011 -837
rect 1017 -838 1018 -837
rect 1066 -838 1067 -837
rect 37 -840 38 -839
rect 387 -840 388 -839
rect 394 -840 395 -839
rect 495 -840 496 -839
rect 558 -840 559 -839
rect 632 -840 633 -839
rect 656 -840 657 -839
rect 1080 -840 1081 -839
rect 51 -842 52 -841
rect 264 -842 265 -841
rect 296 -842 297 -841
rect 555 -842 556 -841
rect 562 -842 563 -841
rect 604 -842 605 -841
rect 611 -842 612 -841
rect 1094 -842 1095 -841
rect 51 -844 52 -843
rect 191 -844 192 -843
rect 198 -844 199 -843
rect 233 -844 234 -843
rect 296 -844 297 -843
rect 324 -844 325 -843
rect 362 -844 363 -843
rect 457 -844 458 -843
rect 464 -844 465 -843
rect 621 -844 622 -843
rect 660 -844 661 -843
rect 667 -844 668 -843
rect 695 -844 696 -843
rect 1087 -844 1088 -843
rect 1094 -844 1095 -843
rect 1178 -844 1179 -843
rect 16 -846 17 -845
rect 191 -846 192 -845
rect 205 -846 206 -845
rect 604 -846 605 -845
rect 621 -846 622 -845
rect 765 -846 766 -845
rect 779 -846 780 -845
rect 828 -846 829 -845
rect 968 -846 969 -845
rect 1038 -846 1039 -845
rect 1073 -846 1074 -845
rect 1087 -846 1088 -845
rect 1178 -846 1179 -845
rect 1220 -846 1221 -845
rect 58 -848 59 -847
rect 61 -848 62 -847
rect 86 -848 87 -847
rect 352 -848 353 -847
rect 380 -848 381 -847
rect 1101 -848 1102 -847
rect 58 -850 59 -849
rect 240 -850 241 -849
rect 289 -850 290 -849
rect 828 -850 829 -849
rect 968 -850 969 -849
rect 982 -850 983 -849
rect 989 -850 990 -849
rect 1129 -850 1130 -849
rect 86 -852 87 -851
rect 681 -852 682 -851
rect 695 -852 696 -851
rect 716 -852 717 -851
rect 730 -852 731 -851
rect 800 -852 801 -851
rect 814 -852 815 -851
rect 1192 -852 1193 -851
rect 5 -854 6 -853
rect 814 -854 815 -853
rect 982 -854 983 -853
rect 1115 -854 1116 -853
rect 1129 -854 1130 -853
rect 1185 -854 1186 -853
rect 1192 -854 1193 -853
rect 1213 -854 1214 -853
rect 93 -856 94 -855
rect 240 -856 241 -855
rect 292 -856 293 -855
rect 800 -856 801 -855
rect 1017 -856 1018 -855
rect 1059 -856 1060 -855
rect 1073 -856 1074 -855
rect 1136 -856 1137 -855
rect 93 -858 94 -857
rect 100 -858 101 -857
rect 114 -858 115 -857
rect 1031 -858 1032 -857
rect 1059 -858 1060 -857
rect 1122 -858 1123 -857
rect 117 -860 118 -859
rect 380 -860 381 -859
rect 422 -860 423 -859
rect 506 -860 507 -859
rect 569 -860 570 -859
rect 583 -860 584 -859
rect 663 -860 664 -859
rect 667 -860 668 -859
rect 681 -860 682 -859
rect 884 -860 885 -859
rect 999 -860 1000 -859
rect 1010 -860 1011 -859
rect 1024 -860 1025 -859
rect 1115 -860 1116 -859
rect 1122 -860 1123 -859
rect 1171 -860 1172 -859
rect 121 -862 122 -861
rect 614 -862 615 -861
rect 698 -862 699 -861
rect 1164 -862 1165 -861
rect 1171 -862 1172 -861
rect 1206 -862 1207 -861
rect 124 -864 125 -863
rect 226 -864 227 -863
rect 324 -864 325 -863
rect 331 -864 332 -863
rect 352 -864 353 -863
rect 436 -864 437 -863
rect 450 -864 451 -863
rect 457 -864 458 -863
rect 464 -864 465 -863
rect 502 -864 503 -863
rect 506 -864 507 -863
rect 576 -864 577 -863
rect 583 -864 584 -863
rect 688 -864 689 -863
rect 702 -864 703 -863
rect 744 -864 745 -863
rect 751 -864 752 -863
rect 765 -864 766 -863
rect 863 -864 864 -863
rect 884 -864 885 -863
rect 1024 -864 1025 -863
rect 1108 -864 1109 -863
rect 1164 -864 1165 -863
rect 1199 -864 1200 -863
rect 135 -866 136 -865
rect 345 -866 346 -865
rect 425 -866 426 -865
rect 625 -866 626 -865
rect 674 -866 675 -865
rect 688 -866 689 -865
rect 716 -866 717 -865
rect 772 -866 773 -865
rect 863 -866 864 -865
rect 891 -866 892 -865
rect 1031 -866 1032 -865
rect 1045 -866 1046 -865
rect 1080 -866 1081 -865
rect 1150 -866 1151 -865
rect 23 -868 24 -867
rect 425 -868 426 -867
rect 429 -868 430 -867
rect 744 -868 745 -867
rect 751 -868 752 -867
rect 793 -868 794 -867
rect 856 -868 857 -867
rect 891 -868 892 -867
rect 1045 -868 1046 -867
rect 1143 -868 1144 -867
rect 23 -870 24 -869
rect 219 -870 220 -869
rect 226 -870 227 -869
rect 278 -870 279 -869
rect 317 -870 318 -869
rect 331 -870 332 -869
rect 429 -870 430 -869
rect 443 -870 444 -869
rect 471 -870 472 -869
rect 723 -870 724 -869
rect 758 -870 759 -869
rect 807 -870 808 -869
rect 835 -870 836 -869
rect 856 -870 857 -869
rect 870 -870 871 -869
rect 1108 -870 1109 -869
rect 107 -872 108 -871
rect 317 -872 318 -871
rect 436 -872 437 -871
rect 597 -872 598 -871
rect 600 -872 601 -871
rect 793 -872 794 -871
rect 807 -872 808 -871
rect 842 -872 843 -871
rect 870 -872 871 -871
rect 961 -872 962 -871
rect 65 -874 66 -873
rect 597 -874 598 -873
rect 674 -874 675 -873
rect 1052 -874 1053 -873
rect 65 -876 66 -875
rect 534 -876 535 -875
rect 576 -876 577 -875
rect 646 -876 647 -875
rect 677 -876 678 -875
rect 835 -876 836 -875
rect 842 -876 843 -875
rect 877 -876 878 -875
rect 898 -876 899 -875
rect 1052 -876 1053 -875
rect 79 -878 80 -877
rect 107 -878 108 -877
rect 149 -878 150 -877
rect 443 -878 444 -877
rect 471 -878 472 -877
rect 670 -878 671 -877
rect 772 -878 773 -877
rect 821 -878 822 -877
rect 877 -878 878 -877
rect 919 -878 920 -877
rect 37 -880 38 -879
rect 79 -880 80 -879
rect 163 -880 164 -879
rect 1157 -880 1158 -879
rect 156 -882 157 -881
rect 163 -882 164 -881
rect 177 -882 178 -881
rect 233 -882 234 -881
rect 485 -882 486 -881
rect 513 -882 514 -881
rect 534 -882 535 -881
rect 548 -882 549 -881
rect 646 -882 647 -881
rect 709 -882 710 -881
rect 817 -882 818 -881
rect 961 -882 962 -881
rect 142 -884 143 -883
rect 177 -884 178 -883
rect 205 -884 206 -883
rect 247 -884 248 -883
rect 415 -884 416 -883
rect 548 -884 549 -883
rect 709 -884 710 -883
rect 737 -884 738 -883
rect 128 -886 129 -885
rect 142 -886 143 -885
rect 149 -886 150 -885
rect 247 -886 248 -885
rect 348 -886 349 -885
rect 415 -886 416 -885
rect 513 -886 514 -885
rect 527 -886 528 -885
rect 544 -886 545 -885
rect 919 -886 920 -885
rect 9 -888 10 -887
rect 128 -888 129 -887
rect 156 -888 157 -887
rect 492 -888 493 -887
rect 527 -888 528 -887
rect 653 -888 654 -887
rect 737 -888 738 -887
rect 933 -888 934 -887
rect 9 -890 10 -889
rect 254 -890 255 -889
rect 366 -890 367 -889
rect 492 -890 493 -889
rect 933 -890 934 -889
rect 940 -890 941 -889
rect 212 -892 213 -891
rect 394 -892 395 -891
rect 926 -892 927 -891
rect 940 -892 941 -891
rect 212 -894 213 -893
rect 408 -894 409 -893
rect 926 -894 927 -893
rect 954 -894 955 -893
rect 219 -896 220 -895
rect 282 -896 283 -895
rect 366 -896 367 -895
rect 373 -896 374 -895
rect 912 -896 913 -895
rect 954 -896 955 -895
rect 40 -898 41 -897
rect 282 -898 283 -897
rect 912 -898 913 -897
rect 1090 -898 1091 -897
rect 254 -900 255 -899
rect 338 -900 339 -899
rect 268 -902 269 -901
rect 408 -902 409 -901
rect 268 -904 269 -903
rect 275 -904 276 -903
rect 310 -904 311 -903
rect 338 -904 339 -903
rect 310 -906 311 -905
rect 450 -906 451 -905
rect 2 -917 3 -916
rect 86 -917 87 -916
rect 96 -917 97 -916
rect 485 -917 486 -916
rect 502 -917 503 -916
rect 513 -917 514 -916
rect 548 -917 549 -916
rect 681 -917 682 -916
rect 684 -917 685 -916
rect 1115 -917 1116 -916
rect 1136 -917 1137 -916
rect 1178 -917 1179 -916
rect 19 -919 20 -918
rect 814 -919 815 -918
rect 824 -919 825 -918
rect 1087 -919 1088 -918
rect 1101 -919 1102 -918
rect 1115 -919 1116 -918
rect 1150 -919 1151 -918
rect 1164 -919 1165 -918
rect 30 -921 31 -920
rect 170 -921 171 -920
rect 205 -921 206 -920
rect 576 -921 577 -920
rect 597 -921 598 -920
rect 870 -921 871 -920
rect 898 -921 899 -920
rect 1122 -921 1123 -920
rect 1157 -921 1158 -920
rect 1171 -921 1172 -920
rect 33 -923 34 -922
rect 499 -923 500 -922
rect 506 -923 507 -922
rect 513 -923 514 -922
rect 548 -923 549 -922
rect 562 -923 563 -922
rect 597 -923 598 -922
rect 828 -923 829 -922
rect 1108 -923 1109 -922
rect 1171 -923 1172 -922
rect 37 -925 38 -924
rect 604 -925 605 -924
rect 618 -925 619 -924
rect 702 -925 703 -924
rect 716 -925 717 -924
rect 1143 -925 1144 -924
rect 1164 -925 1165 -924
rect 1192 -925 1193 -924
rect 40 -927 41 -926
rect 324 -927 325 -926
rect 345 -927 346 -926
rect 492 -927 493 -926
rect 499 -927 500 -926
rect 898 -927 899 -926
rect 1066 -927 1067 -926
rect 1108 -927 1109 -926
rect 1122 -927 1123 -926
rect 1129 -927 1130 -926
rect 1185 -927 1186 -926
rect 1192 -927 1193 -926
rect 9 -929 10 -928
rect 324 -929 325 -928
rect 348 -929 349 -928
rect 408 -929 409 -928
rect 415 -929 416 -928
rect 492 -929 493 -928
rect 555 -929 556 -928
rect 1101 -929 1102 -928
rect 40 -931 41 -930
rect 576 -931 577 -930
rect 628 -931 629 -930
rect 709 -931 710 -930
rect 716 -931 717 -930
rect 730 -931 731 -930
rect 737 -931 738 -930
rect 828 -931 829 -930
rect 1052 -931 1053 -930
rect 1129 -931 1130 -930
rect 44 -933 45 -932
rect 611 -933 612 -932
rect 656 -933 657 -932
rect 989 -933 990 -932
rect 1052 -933 1053 -932
rect 1080 -933 1081 -932
rect 44 -935 45 -934
rect 100 -935 101 -934
rect 117 -935 118 -934
rect 390 -935 391 -934
rect 408 -935 409 -934
rect 558 -935 559 -934
rect 562 -935 563 -934
rect 569 -935 570 -934
rect 667 -935 668 -934
rect 695 -935 696 -934
rect 702 -935 703 -934
rect 772 -935 773 -934
rect 975 -935 976 -934
rect 1080 -935 1081 -934
rect 51 -937 52 -936
rect 114 -937 115 -936
rect 142 -937 143 -936
rect 152 -937 153 -936
rect 170 -937 171 -936
rect 208 -937 209 -936
rect 219 -937 220 -936
rect 436 -937 437 -936
rect 439 -937 440 -936
rect 632 -937 633 -936
rect 674 -937 675 -936
rect 730 -937 731 -936
rect 737 -937 738 -936
rect 786 -937 787 -936
rect 975 -937 976 -936
rect 1017 -937 1018 -936
rect 51 -939 52 -938
rect 61 -939 62 -938
rect 65 -939 66 -938
rect 555 -939 556 -938
rect 632 -939 633 -938
rect 646 -939 647 -938
rect 695 -939 696 -938
rect 870 -939 871 -938
rect 989 -939 990 -938
rect 1031 -939 1032 -938
rect 58 -941 59 -940
rect 114 -941 115 -940
rect 142 -941 143 -940
rect 264 -941 265 -940
rect 268 -941 269 -940
rect 289 -941 290 -940
rect 303 -941 304 -940
rect 310 -941 311 -940
rect 331 -941 332 -940
rect 415 -941 416 -940
rect 439 -941 440 -940
rect 859 -941 860 -940
rect 996 -941 997 -940
rect 1031 -941 1032 -940
rect 58 -943 59 -942
rect 107 -943 108 -942
rect 149 -943 150 -942
rect 233 -943 234 -942
rect 247 -943 248 -942
rect 289 -943 290 -942
rect 303 -943 304 -942
rect 733 -943 734 -942
rect 772 -943 773 -942
rect 863 -943 864 -942
rect 961 -943 962 -942
rect 996 -943 997 -942
rect 1017 -943 1018 -942
rect 1073 -943 1074 -942
rect 72 -945 73 -944
rect 712 -945 713 -944
rect 786 -945 787 -944
rect 800 -945 801 -944
rect 961 -945 962 -944
rect 1010 -945 1011 -944
rect 1038 -945 1039 -944
rect 1073 -945 1074 -944
rect 79 -947 80 -946
rect 107 -947 108 -946
rect 191 -947 192 -946
rect 219 -947 220 -946
rect 233 -947 234 -946
rect 376 -947 377 -946
rect 380 -947 381 -946
rect 653 -947 654 -946
rect 709 -947 710 -946
rect 982 -947 983 -946
rect 1010 -947 1011 -946
rect 1094 -947 1095 -946
rect 79 -949 80 -948
rect 128 -949 129 -948
rect 156 -949 157 -948
rect 191 -949 192 -948
rect 212 -949 213 -948
rect 247 -949 248 -948
rect 261 -949 262 -948
rect 331 -949 332 -948
rect 362 -949 363 -948
rect 814 -949 815 -948
rect 982 -949 983 -948
rect 1090 -949 1091 -948
rect 86 -951 87 -950
rect 93 -951 94 -950
rect 121 -951 122 -950
rect 128 -951 129 -950
rect 156 -951 157 -950
rect 198 -951 199 -950
rect 240 -951 241 -950
rect 261 -951 262 -950
rect 268 -951 269 -950
rect 366 -951 367 -950
rect 373 -951 374 -950
rect 723 -951 724 -950
rect 800 -951 801 -950
rect 856 -951 857 -950
rect 1059 -951 1060 -950
rect 1094 -951 1095 -950
rect 9 -953 10 -952
rect 121 -953 122 -952
rect 177 -953 178 -952
rect 212 -953 213 -952
rect 240 -953 241 -952
rect 254 -953 255 -952
rect 275 -953 276 -952
rect 296 -953 297 -952
rect 352 -953 353 -952
rect 366 -953 367 -952
rect 380 -953 381 -952
rect 387 -953 388 -952
rect 471 -953 472 -952
rect 569 -953 570 -952
rect 607 -953 608 -952
rect 1038 -953 1039 -952
rect 23 -955 24 -954
rect 254 -955 255 -954
rect 275 -955 276 -954
rect 282 -955 283 -954
rect 296 -955 297 -954
rect 317 -955 318 -954
rect 471 -955 472 -954
rect 583 -955 584 -954
rect 625 -955 626 -954
rect 863 -955 864 -954
rect 1024 -955 1025 -954
rect 1059 -955 1060 -954
rect 23 -957 24 -956
rect 100 -957 101 -956
rect 135 -957 136 -956
rect 352 -957 353 -956
rect 478 -957 479 -956
rect 520 -957 521 -956
rect 583 -957 584 -956
rect 660 -957 661 -956
rect 723 -957 724 -956
rect 779 -957 780 -956
rect 821 -957 822 -956
rect 1024 -957 1025 -956
rect 72 -959 73 -958
rect 198 -959 199 -958
rect 317 -959 318 -958
rect 450 -959 451 -958
rect 485 -959 486 -958
rect 527 -959 528 -958
rect 544 -959 545 -958
rect 660 -959 661 -958
rect 744 -959 745 -958
rect 779 -959 780 -958
rect 821 -959 822 -958
rect 905 -959 906 -958
rect 93 -961 94 -960
rect 1066 -961 1067 -960
rect 135 -963 136 -962
rect 614 -963 615 -962
rect 653 -963 654 -962
rect 688 -963 689 -962
rect 744 -963 745 -962
rect 793 -963 794 -962
rect 905 -963 906 -962
rect 954 -963 955 -962
rect 177 -965 178 -964
rect 184 -965 185 -964
rect 359 -965 360 -964
rect 520 -965 521 -964
rect 527 -965 528 -964
rect 534 -965 535 -964
rect 688 -965 689 -964
rect 751 -965 752 -964
rect 793 -965 794 -964
rect 807 -965 808 -964
rect 954 -965 955 -964
rect 968 -965 969 -964
rect 184 -967 185 -966
rect 282 -967 283 -966
rect 443 -967 444 -966
rect 534 -967 535 -966
rect 751 -967 752 -966
rect 849 -967 850 -966
rect 968 -967 969 -966
rect 1045 -967 1046 -966
rect 422 -969 423 -968
rect 1045 -969 1046 -968
rect 422 -971 423 -970
rect 464 -971 465 -970
rect 807 -971 808 -970
rect 877 -971 878 -970
rect 429 -973 430 -972
rect 443 -973 444 -972
rect 450 -973 451 -972
rect 590 -973 591 -972
rect 849 -973 850 -972
rect 891 -973 892 -972
rect 429 -975 430 -974
rect 457 -975 458 -974
rect 590 -975 591 -974
rect 835 -975 836 -974
rect 877 -975 878 -974
rect 919 -975 920 -974
rect 457 -977 458 -976
rect 639 -977 640 -976
rect 765 -977 766 -976
rect 891 -977 892 -976
rect 758 -979 759 -978
rect 765 -979 766 -978
rect 835 -979 836 -978
rect 947 -979 948 -978
rect 65 -981 66 -980
rect 758 -981 759 -980
rect 884 -981 885 -980
rect 919 -981 920 -980
rect 933 -981 934 -980
rect 947 -981 948 -980
rect 842 -983 843 -982
rect 933 -983 934 -982
rect 842 -985 843 -984
rect 901 -985 902 -984
rect 884 -987 885 -986
rect 926 -987 927 -986
rect 926 -989 927 -988
rect 940 -989 941 -988
rect 940 -991 941 -990
rect 1003 -991 1004 -990
rect 912 -993 913 -992
rect 1003 -993 1004 -992
rect 604 -995 605 -994
rect 912 -995 913 -994
rect 9 -1006 10 -1005
rect 93 -1006 94 -1005
rect 100 -1006 101 -1005
rect 107 -1006 108 -1005
rect 121 -1006 122 -1005
rect 338 -1006 339 -1005
rect 359 -1006 360 -1005
rect 422 -1006 423 -1005
rect 464 -1006 465 -1005
rect 513 -1006 514 -1005
rect 541 -1006 542 -1005
rect 765 -1006 766 -1005
rect 810 -1006 811 -1005
rect 954 -1006 955 -1005
rect 1129 -1006 1130 -1005
rect 1157 -1006 1158 -1005
rect 37 -1008 38 -1007
rect 65 -1008 66 -1007
rect 89 -1008 90 -1007
rect 863 -1008 864 -1007
rect 884 -1008 885 -1007
rect 887 -1008 888 -1007
rect 954 -1008 955 -1007
rect 1115 -1008 1116 -1007
rect 1136 -1008 1137 -1007
rect 1150 -1008 1151 -1007
rect 40 -1010 41 -1009
rect 544 -1010 545 -1009
rect 569 -1010 570 -1009
rect 607 -1010 608 -1009
rect 625 -1010 626 -1009
rect 723 -1010 724 -1009
rect 730 -1010 731 -1009
rect 1094 -1010 1095 -1009
rect 44 -1012 45 -1011
rect 198 -1012 199 -1011
rect 208 -1012 209 -1011
rect 212 -1012 213 -1011
rect 219 -1012 220 -1011
rect 355 -1012 356 -1011
rect 362 -1012 363 -1011
rect 1038 -1012 1039 -1011
rect 1094 -1012 1095 -1011
rect 1171 -1012 1172 -1011
rect 16 -1014 17 -1013
rect 44 -1014 45 -1013
rect 58 -1014 59 -1013
rect 72 -1014 73 -1013
rect 107 -1014 108 -1013
rect 394 -1014 395 -1013
rect 401 -1014 402 -1013
rect 513 -1014 514 -1013
rect 527 -1014 528 -1013
rect 541 -1014 542 -1013
rect 597 -1014 598 -1013
rect 642 -1014 643 -1013
rect 646 -1014 647 -1013
rect 674 -1014 675 -1013
rect 681 -1014 682 -1013
rect 705 -1014 706 -1013
rect 723 -1014 724 -1013
rect 835 -1014 836 -1013
rect 856 -1014 857 -1013
rect 1080 -1014 1081 -1013
rect 16 -1016 17 -1015
rect 103 -1016 104 -1015
rect 124 -1016 125 -1015
rect 359 -1016 360 -1015
rect 457 -1016 458 -1015
rect 527 -1016 528 -1015
rect 600 -1016 601 -1015
rect 793 -1016 794 -1015
rect 856 -1016 857 -1015
rect 877 -1016 878 -1015
rect 884 -1016 885 -1015
rect 905 -1016 906 -1015
rect 1024 -1016 1025 -1015
rect 1038 -1016 1039 -1015
rect 1069 -1016 1070 -1015
rect 1080 -1016 1081 -1015
rect 30 -1018 31 -1017
rect 219 -1018 220 -1017
rect 254 -1018 255 -1017
rect 387 -1018 388 -1017
rect 443 -1018 444 -1017
rect 457 -1018 458 -1017
rect 499 -1018 500 -1017
rect 982 -1018 983 -1017
rect 996 -1018 997 -1017
rect 1024 -1018 1025 -1017
rect 30 -1020 31 -1019
rect 142 -1020 143 -1019
rect 184 -1020 185 -1019
rect 282 -1020 283 -1019
rect 289 -1020 290 -1019
rect 320 -1020 321 -1019
rect 338 -1020 339 -1019
rect 380 -1020 381 -1019
rect 429 -1020 430 -1019
rect 443 -1020 444 -1019
rect 499 -1020 500 -1019
rect 583 -1020 584 -1019
rect 604 -1020 605 -1019
rect 691 -1020 692 -1019
rect 695 -1020 696 -1019
rect 737 -1020 738 -1019
rect 751 -1020 752 -1019
rect 765 -1020 766 -1019
rect 786 -1020 787 -1019
rect 835 -1020 836 -1019
rect 859 -1020 860 -1019
rect 1108 -1020 1109 -1019
rect 61 -1022 62 -1021
rect 548 -1022 549 -1021
rect 632 -1022 633 -1021
rect 674 -1022 675 -1021
rect 681 -1022 682 -1021
rect 688 -1022 689 -1021
rect 698 -1022 699 -1021
rect 793 -1022 794 -1021
rect 863 -1022 864 -1021
rect 898 -1022 899 -1021
rect 905 -1022 906 -1021
rect 968 -1022 969 -1021
rect 982 -1022 983 -1021
rect 1010 -1022 1011 -1021
rect 65 -1024 66 -1023
rect 408 -1024 409 -1023
rect 429 -1024 430 -1023
rect 485 -1024 486 -1023
rect 502 -1024 503 -1023
rect 1101 -1024 1102 -1023
rect 72 -1026 73 -1025
rect 275 -1026 276 -1025
rect 289 -1026 290 -1025
rect 296 -1026 297 -1025
rect 317 -1026 318 -1025
rect 422 -1026 423 -1025
rect 471 -1026 472 -1025
rect 583 -1026 584 -1025
rect 639 -1026 640 -1025
rect 1087 -1026 1088 -1025
rect 79 -1028 80 -1027
rect 282 -1028 283 -1027
rect 317 -1028 318 -1027
rect 597 -1028 598 -1027
rect 639 -1028 640 -1027
rect 653 -1028 654 -1027
rect 660 -1028 661 -1027
rect 737 -1028 738 -1027
rect 751 -1028 752 -1027
rect 821 -1028 822 -1027
rect 968 -1028 969 -1027
rect 989 -1028 990 -1027
rect 996 -1028 997 -1027
rect 1017 -1028 1018 -1027
rect 1087 -1028 1088 -1027
rect 1122 -1028 1123 -1027
rect 79 -1030 80 -1029
rect 149 -1030 150 -1029
rect 187 -1030 188 -1029
rect 779 -1030 780 -1029
rect 786 -1030 787 -1029
rect 919 -1030 920 -1029
rect 989 -1030 990 -1029
rect 1066 -1030 1067 -1029
rect 1122 -1030 1123 -1029
rect 1167 -1030 1168 -1029
rect 96 -1032 97 -1031
rect 394 -1032 395 -1031
rect 408 -1032 409 -1031
rect 415 -1032 416 -1031
rect 485 -1032 486 -1031
rect 562 -1032 563 -1031
rect 649 -1032 650 -1031
rect 891 -1032 892 -1031
rect 919 -1032 920 -1031
rect 1073 -1032 1074 -1031
rect 86 -1034 87 -1033
rect 96 -1034 97 -1033
rect 114 -1034 115 -1033
rect 142 -1034 143 -1033
rect 191 -1034 192 -1033
rect 198 -1034 199 -1033
rect 205 -1034 206 -1033
rect 471 -1034 472 -1033
rect 509 -1034 510 -1033
rect 534 -1034 535 -1033
rect 653 -1034 654 -1033
rect 702 -1034 703 -1033
rect 716 -1034 717 -1033
rect 877 -1034 878 -1033
rect 891 -1034 892 -1033
rect 912 -1034 913 -1033
rect 1010 -1034 1011 -1033
rect 1132 -1034 1133 -1033
rect 2 -1036 3 -1035
rect 205 -1036 206 -1035
rect 212 -1036 213 -1035
rect 240 -1036 241 -1035
rect 268 -1036 269 -1035
rect 373 -1036 374 -1035
rect 376 -1036 377 -1035
rect 898 -1036 899 -1035
rect 912 -1036 913 -1035
rect 926 -1036 927 -1035
rect 1017 -1036 1018 -1035
rect 1052 -1036 1053 -1035
rect 170 -1038 171 -1037
rect 268 -1038 269 -1037
rect 331 -1038 332 -1037
rect 548 -1038 549 -1037
rect 572 -1038 573 -1037
rect 926 -1038 927 -1037
rect 177 -1040 178 -1039
rect 191 -1040 192 -1039
rect 226 -1040 227 -1039
rect 275 -1040 276 -1039
rect 303 -1040 304 -1039
rect 331 -1040 332 -1039
rect 373 -1040 374 -1039
rect 478 -1040 479 -1039
rect 506 -1040 507 -1039
rect 702 -1040 703 -1039
rect 716 -1040 717 -1039
rect 772 -1040 773 -1039
rect 779 -1040 780 -1039
rect 807 -1040 808 -1039
rect 821 -1040 822 -1039
rect 870 -1040 871 -1039
rect 86 -1042 87 -1041
rect 226 -1042 227 -1041
rect 233 -1042 234 -1041
rect 254 -1042 255 -1041
rect 303 -1042 304 -1041
rect 310 -1042 311 -1041
rect 380 -1042 381 -1041
rect 436 -1042 437 -1041
rect 450 -1042 451 -1041
rect 562 -1042 563 -1041
rect 660 -1042 661 -1041
rect 667 -1042 668 -1041
rect 684 -1042 685 -1041
rect 1059 -1042 1060 -1041
rect 117 -1044 118 -1043
rect 233 -1044 234 -1043
rect 240 -1044 241 -1043
rect 264 -1044 265 -1043
rect 401 -1044 402 -1043
rect 436 -1044 437 -1043
rect 450 -1044 451 -1043
rect 611 -1044 612 -1043
rect 667 -1044 668 -1043
rect 709 -1044 710 -1043
rect 733 -1044 734 -1043
rect 1031 -1044 1032 -1043
rect 1059 -1044 1060 -1043
rect 1073 -1044 1074 -1043
rect 152 -1046 153 -1045
rect 310 -1046 311 -1045
rect 415 -1046 416 -1045
rect 621 -1046 622 -1045
rect 688 -1046 689 -1045
rect 814 -1046 815 -1045
rect 842 -1046 843 -1045
rect 870 -1046 871 -1045
rect 1031 -1046 1032 -1045
rect 1052 -1046 1053 -1045
rect 156 -1048 157 -1047
rect 177 -1048 178 -1047
rect 390 -1048 391 -1047
rect 842 -1048 843 -1047
rect 156 -1050 157 -1049
rect 163 -1050 164 -1049
rect 478 -1050 479 -1049
rect 492 -1050 493 -1049
rect 534 -1050 535 -1049
rect 933 -1050 934 -1049
rect 135 -1052 136 -1051
rect 163 -1052 164 -1051
rect 201 -1052 202 -1051
rect 933 -1052 934 -1051
rect 135 -1054 136 -1053
rect 324 -1054 325 -1053
rect 345 -1054 346 -1053
rect 492 -1054 493 -1053
rect 576 -1054 577 -1053
rect 611 -1054 612 -1053
rect 709 -1054 710 -1053
rect 744 -1054 745 -1053
rect 772 -1054 773 -1053
rect 800 -1054 801 -1053
rect 814 -1054 815 -1053
rect 849 -1054 850 -1053
rect 247 -1056 248 -1055
rect 324 -1056 325 -1055
rect 345 -1056 346 -1055
rect 352 -1056 353 -1055
rect 576 -1056 577 -1055
rect 618 -1056 619 -1055
rect 744 -1056 745 -1055
rect 828 -1056 829 -1055
rect 849 -1056 850 -1055
rect 1045 -1056 1046 -1055
rect 247 -1058 248 -1057
rect 261 -1058 262 -1057
rect 352 -1058 353 -1057
rect 590 -1058 591 -1057
rect 618 -1058 619 -1057
rect 947 -1058 948 -1057
rect 520 -1060 521 -1059
rect 590 -1060 591 -1059
rect 758 -1060 759 -1059
rect 828 -1060 829 -1059
rect 887 -1060 888 -1059
rect 1066 -1060 1067 -1059
rect 173 -1062 174 -1061
rect 520 -1062 521 -1061
rect 800 -1062 801 -1061
rect 1143 -1062 1144 -1061
rect 940 -1064 941 -1063
rect 947 -1064 948 -1063
rect 940 -1066 941 -1065
rect 961 -1066 962 -1065
rect 961 -1068 962 -1067
rect 975 -1068 976 -1067
rect 61 -1070 62 -1069
rect 975 -1070 976 -1069
rect 16 -1081 17 -1080
rect 187 -1081 188 -1080
rect 219 -1081 220 -1080
rect 446 -1081 447 -1080
rect 471 -1081 472 -1080
rect 618 -1081 619 -1080
rect 632 -1081 633 -1080
rect 695 -1081 696 -1080
rect 852 -1081 853 -1080
rect 877 -1081 878 -1080
rect 884 -1081 885 -1080
rect 887 -1081 888 -1080
rect 954 -1081 955 -1080
rect 961 -1081 962 -1080
rect 978 -1081 979 -1080
rect 1017 -1081 1018 -1080
rect 1031 -1081 1032 -1080
rect 1038 -1081 1039 -1080
rect 1041 -1081 1042 -1080
rect 1052 -1081 1053 -1080
rect 1108 -1081 1109 -1080
rect 1122 -1081 1123 -1080
rect 1185 -1081 1186 -1080
rect 1188 -1081 1189 -1080
rect 23 -1083 24 -1082
rect 149 -1083 150 -1082
rect 170 -1083 171 -1082
rect 590 -1083 591 -1082
rect 600 -1083 601 -1082
rect 730 -1083 731 -1082
rect 877 -1083 878 -1082
rect 926 -1083 927 -1082
rect 940 -1083 941 -1082
rect 961 -1083 962 -1082
rect 1006 -1083 1007 -1082
rect 1094 -1083 1095 -1082
rect 30 -1085 31 -1084
rect 264 -1085 265 -1084
rect 268 -1085 269 -1084
rect 306 -1085 307 -1084
rect 355 -1085 356 -1084
rect 597 -1085 598 -1084
rect 607 -1085 608 -1084
rect 751 -1085 752 -1084
rect 884 -1085 885 -1084
rect 898 -1085 899 -1084
rect 940 -1085 941 -1084
rect 947 -1085 948 -1084
rect 1017 -1085 1018 -1084
rect 1024 -1085 1025 -1084
rect 1045 -1085 1046 -1084
rect 1059 -1085 1060 -1084
rect 30 -1087 31 -1086
rect 44 -1087 45 -1086
rect 58 -1087 59 -1086
rect 166 -1087 167 -1086
rect 170 -1087 171 -1086
rect 177 -1087 178 -1086
rect 191 -1087 192 -1086
rect 219 -1087 220 -1086
rect 247 -1087 248 -1086
rect 268 -1087 269 -1086
rect 275 -1087 276 -1086
rect 506 -1087 507 -1086
rect 509 -1087 510 -1086
rect 849 -1087 850 -1086
rect 891 -1087 892 -1086
rect 898 -1087 899 -1086
rect 947 -1087 948 -1086
rect 1003 -1087 1004 -1086
rect 1010 -1087 1011 -1086
rect 1024 -1087 1025 -1086
rect 1048 -1087 1049 -1086
rect 1087 -1087 1088 -1086
rect 37 -1089 38 -1088
rect 299 -1089 300 -1088
rect 387 -1089 388 -1088
rect 467 -1089 468 -1088
rect 485 -1089 486 -1088
rect 628 -1089 629 -1088
rect 667 -1089 668 -1088
rect 751 -1089 752 -1088
rect 887 -1089 888 -1088
rect 891 -1089 892 -1088
rect 989 -1089 990 -1088
rect 1010 -1089 1011 -1088
rect 1080 -1089 1081 -1088
rect 1087 -1089 1088 -1088
rect 37 -1091 38 -1090
rect 128 -1091 129 -1090
rect 149 -1091 150 -1090
rect 156 -1091 157 -1090
rect 177 -1091 178 -1090
rect 212 -1091 213 -1090
rect 296 -1091 297 -1090
rect 611 -1091 612 -1090
rect 621 -1091 622 -1090
rect 632 -1091 633 -1090
rect 667 -1091 668 -1090
rect 842 -1091 843 -1090
rect 982 -1091 983 -1090
rect 989 -1091 990 -1090
rect 1073 -1091 1074 -1090
rect 1080 -1091 1081 -1090
rect 44 -1093 45 -1092
rect 450 -1093 451 -1092
rect 551 -1093 552 -1092
rect 576 -1093 577 -1092
rect 586 -1093 587 -1092
rect 926 -1093 927 -1092
rect 968 -1093 969 -1092
rect 982 -1093 983 -1092
rect 65 -1095 66 -1094
rect 68 -1095 69 -1094
rect 72 -1095 73 -1094
rect 464 -1095 465 -1094
rect 499 -1095 500 -1094
rect 576 -1095 577 -1094
rect 590 -1095 591 -1094
rect 737 -1095 738 -1094
rect 842 -1095 843 -1094
rect 870 -1095 871 -1094
rect 968 -1095 969 -1094
rect 975 -1095 976 -1094
rect 72 -1097 73 -1096
rect 82 -1097 83 -1096
rect 93 -1097 94 -1096
rect 100 -1097 101 -1096
rect 121 -1097 122 -1096
rect 352 -1097 353 -1096
rect 366 -1097 367 -1096
rect 464 -1097 465 -1096
rect 499 -1097 500 -1096
rect 555 -1097 556 -1096
rect 572 -1097 573 -1096
rect 583 -1097 584 -1096
rect 604 -1097 605 -1096
rect 611 -1097 612 -1096
rect 670 -1097 671 -1096
rect 1031 -1097 1032 -1096
rect 79 -1099 80 -1098
rect 128 -1099 129 -1098
rect 156 -1099 157 -1098
rect 534 -1099 535 -1098
rect 583 -1099 584 -1098
rect 653 -1099 654 -1098
rect 681 -1099 682 -1098
rect 695 -1099 696 -1098
rect 702 -1099 703 -1098
rect 870 -1099 871 -1098
rect 100 -1101 101 -1100
rect 117 -1101 118 -1100
rect 121 -1101 122 -1100
rect 184 -1101 185 -1100
rect 191 -1101 192 -1100
rect 324 -1101 325 -1100
rect 359 -1101 360 -1100
rect 702 -1101 703 -1100
rect 709 -1101 710 -1100
rect 737 -1101 738 -1100
rect 184 -1103 185 -1102
rect 418 -1103 419 -1102
rect 422 -1103 423 -1102
rect 471 -1103 472 -1102
rect 534 -1103 535 -1102
rect 733 -1103 734 -1102
rect 212 -1105 213 -1104
rect 331 -1105 332 -1104
rect 373 -1105 374 -1104
rect 555 -1105 556 -1104
rect 646 -1105 647 -1104
rect 709 -1105 710 -1104
rect 226 -1107 227 -1106
rect 366 -1107 367 -1106
rect 387 -1107 388 -1106
rect 513 -1107 514 -1106
rect 646 -1107 647 -1106
rect 919 -1107 920 -1106
rect 226 -1109 227 -1108
rect 247 -1109 248 -1108
rect 282 -1109 283 -1108
rect 324 -1109 325 -1108
rect 338 -1109 339 -1108
rect 373 -1109 374 -1108
rect 422 -1109 423 -1108
rect 569 -1109 570 -1108
rect 688 -1109 689 -1108
rect 723 -1109 724 -1108
rect 919 -1109 920 -1108
rect 933 -1109 934 -1108
rect 240 -1111 241 -1110
rect 359 -1111 360 -1110
rect 436 -1111 437 -1110
rect 478 -1111 479 -1110
rect 513 -1111 514 -1110
rect 527 -1111 528 -1110
rect 562 -1111 563 -1110
rect 569 -1111 570 -1110
rect 688 -1111 689 -1110
rect 800 -1111 801 -1110
rect 933 -1111 934 -1110
rect 1066 -1111 1067 -1110
rect 240 -1113 241 -1112
rect 537 -1113 538 -1112
rect 723 -1113 724 -1112
rect 828 -1113 829 -1112
rect 1003 -1113 1004 -1112
rect 1066 -1113 1067 -1112
rect 275 -1115 276 -1114
rect 282 -1115 283 -1114
rect 289 -1115 290 -1114
rect 296 -1115 297 -1114
rect 317 -1115 318 -1114
rect 681 -1115 682 -1114
rect 800 -1115 801 -1114
rect 814 -1115 815 -1114
rect 821 -1115 822 -1114
rect 828 -1115 829 -1114
rect 233 -1117 234 -1116
rect 289 -1117 290 -1116
rect 303 -1117 304 -1116
rect 317 -1117 318 -1116
rect 331 -1117 332 -1116
rect 436 -1117 437 -1116
rect 443 -1117 444 -1116
rect 485 -1117 486 -1116
rect 492 -1117 493 -1116
rect 562 -1117 563 -1116
rect 744 -1117 745 -1116
rect 821 -1117 822 -1116
rect 163 -1119 164 -1118
rect 233 -1119 234 -1118
rect 338 -1119 339 -1118
rect 415 -1119 416 -1118
rect 429 -1119 430 -1118
rect 492 -1119 493 -1118
rect 527 -1119 528 -1118
rect 541 -1119 542 -1118
rect 744 -1119 745 -1118
rect 863 -1119 864 -1118
rect 401 -1121 402 -1120
rect 429 -1121 430 -1120
rect 450 -1121 451 -1120
rect 457 -1121 458 -1120
rect 478 -1121 479 -1120
rect 807 -1121 808 -1120
rect 814 -1121 815 -1120
rect 835 -1121 836 -1120
rect 205 -1123 206 -1122
rect 457 -1123 458 -1122
rect 541 -1123 542 -1122
rect 625 -1123 626 -1122
rect 653 -1123 654 -1122
rect 835 -1123 836 -1122
rect 198 -1125 199 -1124
rect 205 -1125 206 -1124
rect 261 -1125 262 -1124
rect 401 -1125 402 -1124
rect 408 -1125 409 -1124
rect 415 -1125 416 -1124
rect 793 -1125 794 -1124
rect 863 -1125 864 -1124
rect 261 -1127 262 -1126
rect 310 -1127 311 -1126
rect 779 -1127 780 -1126
rect 793 -1127 794 -1126
rect 310 -1129 311 -1128
rect 810 -1129 811 -1128
rect 772 -1131 773 -1130
rect 779 -1131 780 -1130
rect 810 -1131 811 -1130
rect 905 -1131 906 -1130
rect 758 -1133 759 -1132
rect 772 -1133 773 -1132
rect 786 -1133 787 -1132
rect 905 -1133 906 -1132
rect 716 -1135 717 -1134
rect 786 -1135 787 -1134
rect 520 -1137 521 -1136
rect 716 -1137 717 -1136
rect 758 -1137 759 -1136
rect 765 -1137 766 -1136
rect 520 -1139 521 -1138
rect 957 -1139 958 -1138
rect 548 -1141 549 -1140
rect 765 -1141 766 -1140
rect 394 -1143 395 -1142
rect 548 -1143 549 -1142
rect 380 -1145 381 -1144
rect 394 -1145 395 -1144
rect 107 -1147 108 -1146
rect 380 -1147 381 -1146
rect 107 -1149 108 -1148
rect 142 -1149 143 -1148
rect 135 -1151 136 -1150
rect 142 -1151 143 -1150
rect 135 -1153 136 -1152
rect 408 -1153 409 -1152
rect 16 -1164 17 -1163
rect 121 -1164 122 -1163
rect 149 -1164 150 -1163
rect 163 -1164 164 -1163
rect 170 -1164 171 -1163
rect 198 -1164 199 -1163
rect 226 -1164 227 -1163
rect 268 -1164 269 -1163
rect 285 -1164 286 -1163
rect 317 -1164 318 -1163
rect 331 -1164 332 -1163
rect 352 -1164 353 -1163
rect 446 -1164 447 -1163
rect 933 -1164 934 -1163
rect 975 -1164 976 -1163
rect 1038 -1164 1039 -1163
rect 1066 -1164 1067 -1163
rect 1122 -1164 1123 -1163
rect 23 -1166 24 -1165
rect 26 -1166 27 -1165
rect 30 -1166 31 -1165
rect 156 -1166 157 -1165
rect 163 -1166 164 -1165
rect 247 -1166 248 -1165
rect 254 -1166 255 -1165
rect 667 -1166 668 -1165
rect 695 -1166 696 -1165
rect 807 -1166 808 -1165
rect 828 -1166 829 -1165
rect 936 -1166 937 -1165
rect 961 -1166 962 -1165
rect 975 -1166 976 -1165
rect 989 -1166 990 -1165
rect 1066 -1166 1067 -1165
rect 1080 -1166 1081 -1165
rect 1129 -1166 1130 -1165
rect 30 -1168 31 -1167
rect 499 -1168 500 -1167
rect 506 -1168 507 -1167
rect 555 -1168 556 -1167
rect 562 -1168 563 -1167
rect 604 -1168 605 -1167
rect 618 -1168 619 -1167
rect 656 -1168 657 -1167
rect 667 -1168 668 -1167
rect 688 -1168 689 -1167
rect 695 -1168 696 -1167
rect 765 -1168 766 -1167
rect 831 -1168 832 -1167
rect 877 -1168 878 -1167
rect 884 -1168 885 -1167
rect 961 -1168 962 -1167
rect 996 -1168 997 -1167
rect 1003 -1168 1004 -1167
rect 1010 -1168 1011 -1167
rect 1038 -1168 1039 -1167
rect 1087 -1168 1088 -1167
rect 1115 -1168 1116 -1167
rect 37 -1170 38 -1169
rect 138 -1170 139 -1169
rect 152 -1170 153 -1169
rect 478 -1170 479 -1169
rect 499 -1170 500 -1169
rect 509 -1170 510 -1169
rect 544 -1170 545 -1169
rect 884 -1170 885 -1169
rect 919 -1170 920 -1169
rect 996 -1170 997 -1169
rect 1024 -1170 1025 -1169
rect 1052 -1170 1053 -1169
rect 1101 -1170 1102 -1169
rect 1108 -1170 1109 -1169
rect 37 -1172 38 -1171
rect 726 -1172 727 -1171
rect 730 -1172 731 -1171
rect 1080 -1172 1081 -1171
rect 44 -1174 45 -1173
rect 114 -1174 115 -1173
rect 117 -1174 118 -1173
rect 121 -1174 122 -1173
rect 170 -1174 171 -1173
rect 275 -1174 276 -1173
rect 352 -1174 353 -1173
rect 593 -1174 594 -1173
rect 607 -1174 608 -1173
rect 877 -1174 878 -1173
rect 926 -1174 927 -1173
rect 1073 -1174 1074 -1173
rect 58 -1176 59 -1175
rect 156 -1176 157 -1175
rect 177 -1176 178 -1175
rect 198 -1176 199 -1175
rect 229 -1176 230 -1175
rect 359 -1176 360 -1175
rect 443 -1176 444 -1175
rect 1010 -1176 1011 -1175
rect 1031 -1176 1032 -1175
rect 1087 -1176 1088 -1175
rect 51 -1178 52 -1177
rect 58 -1178 59 -1177
rect 72 -1178 73 -1177
rect 128 -1178 129 -1177
rect 184 -1178 185 -1177
rect 345 -1178 346 -1177
rect 359 -1178 360 -1177
rect 380 -1178 381 -1177
rect 478 -1178 479 -1177
rect 485 -1178 486 -1177
rect 562 -1178 563 -1177
rect 821 -1178 822 -1177
rect 842 -1178 843 -1177
rect 919 -1178 920 -1177
rect 954 -1178 955 -1177
rect 989 -1178 990 -1177
rect 1017 -1178 1018 -1177
rect 1031 -1178 1032 -1177
rect 1059 -1178 1060 -1177
rect 1108 -1178 1109 -1177
rect 65 -1180 66 -1179
rect 72 -1180 73 -1179
rect 79 -1180 80 -1179
rect 583 -1180 584 -1179
rect 586 -1180 587 -1179
rect 723 -1180 724 -1179
rect 730 -1180 731 -1179
rect 793 -1180 794 -1179
rect 814 -1180 815 -1179
rect 842 -1180 843 -1179
rect 849 -1180 850 -1179
rect 891 -1180 892 -1179
rect 940 -1180 941 -1179
rect 1017 -1180 1018 -1179
rect 51 -1182 52 -1181
rect 65 -1182 66 -1181
rect 82 -1182 83 -1181
rect 338 -1182 339 -1181
rect 429 -1182 430 -1181
rect 583 -1182 584 -1181
rect 590 -1182 591 -1181
rect 604 -1182 605 -1181
rect 625 -1182 626 -1181
rect 1045 -1182 1046 -1181
rect 89 -1184 90 -1183
rect 135 -1184 136 -1183
rect 187 -1184 188 -1183
rect 814 -1184 815 -1183
rect 863 -1184 864 -1183
rect 978 -1184 979 -1183
rect 107 -1186 108 -1185
rect 345 -1186 346 -1185
rect 429 -1186 430 -1185
rect 646 -1186 647 -1185
rect 653 -1186 654 -1185
rect 716 -1186 717 -1185
rect 765 -1186 766 -1185
rect 856 -1186 857 -1185
rect 870 -1186 871 -1185
rect 926 -1186 927 -1185
rect 968 -1186 969 -1185
rect 1059 -1186 1060 -1185
rect 61 -1188 62 -1187
rect 968 -1188 969 -1187
rect 107 -1190 108 -1189
rect 383 -1190 384 -1189
rect 450 -1190 451 -1189
rect 485 -1190 486 -1189
rect 565 -1190 566 -1189
rect 870 -1190 871 -1189
rect 891 -1190 892 -1189
rect 912 -1190 913 -1189
rect 233 -1192 234 -1191
rect 303 -1192 304 -1191
rect 306 -1192 307 -1191
rect 338 -1192 339 -1191
rect 401 -1192 402 -1191
rect 450 -1192 451 -1191
rect 569 -1192 570 -1191
rect 618 -1192 619 -1191
rect 625 -1192 626 -1191
rect 639 -1192 640 -1191
rect 646 -1192 647 -1191
rect 674 -1192 675 -1191
rect 688 -1192 689 -1191
rect 758 -1192 759 -1191
rect 772 -1192 773 -1191
rect 1024 -1192 1025 -1191
rect 131 -1194 132 -1193
rect 758 -1194 759 -1193
rect 772 -1194 773 -1193
rect 1094 -1194 1095 -1193
rect 233 -1196 234 -1195
rect 548 -1196 549 -1195
rect 555 -1196 556 -1195
rect 569 -1196 570 -1195
rect 611 -1196 612 -1195
rect 863 -1196 864 -1195
rect 898 -1196 899 -1195
rect 940 -1196 941 -1195
rect 240 -1198 241 -1197
rect 247 -1198 248 -1197
rect 254 -1198 255 -1197
rect 810 -1198 811 -1197
rect 898 -1198 899 -1197
rect 947 -1198 948 -1197
rect 240 -1200 241 -1199
rect 289 -1200 290 -1199
rect 317 -1200 318 -1199
rect 716 -1200 717 -1199
rect 744 -1200 745 -1199
rect 912 -1200 913 -1199
rect 261 -1202 262 -1201
rect 282 -1202 283 -1201
rect 289 -1202 290 -1201
rect 296 -1202 297 -1201
rect 394 -1202 395 -1201
rect 401 -1202 402 -1201
rect 597 -1202 598 -1201
rect 744 -1202 745 -1201
rect 779 -1202 780 -1201
rect 821 -1202 822 -1201
rect 166 -1204 167 -1203
rect 394 -1204 395 -1203
rect 408 -1204 409 -1203
rect 779 -1204 780 -1203
rect 786 -1204 787 -1203
rect 793 -1204 794 -1203
rect 800 -1204 801 -1203
rect 856 -1204 857 -1203
rect 212 -1206 213 -1205
rect 296 -1206 297 -1205
rect 408 -1206 409 -1205
rect 457 -1206 458 -1205
rect 509 -1206 510 -1205
rect 800 -1206 801 -1205
rect 191 -1208 192 -1207
rect 212 -1208 213 -1207
rect 268 -1208 269 -1207
rect 310 -1208 311 -1207
rect 457 -1208 458 -1207
rect 471 -1208 472 -1207
rect 534 -1208 535 -1207
rect 597 -1208 598 -1207
rect 611 -1208 612 -1207
rect 656 -1208 657 -1207
rect 674 -1208 675 -1207
rect 737 -1208 738 -1207
rect 751 -1208 752 -1207
rect 786 -1208 787 -1207
rect 191 -1210 192 -1209
rect 520 -1210 521 -1209
rect 527 -1210 528 -1209
rect 534 -1210 535 -1209
rect 660 -1210 661 -1209
rect 737 -1210 738 -1209
rect 751 -1210 752 -1209
rect 835 -1210 836 -1209
rect 275 -1212 276 -1211
rect 373 -1212 374 -1211
rect 464 -1212 465 -1211
rect 471 -1212 472 -1211
rect 513 -1212 514 -1211
rect 520 -1212 521 -1211
rect 527 -1212 528 -1211
rect 551 -1212 552 -1211
rect 681 -1212 682 -1211
rect 947 -1212 948 -1211
rect 23 -1214 24 -1213
rect 464 -1214 465 -1213
rect 541 -1214 542 -1213
rect 835 -1214 836 -1213
rect 310 -1216 311 -1215
rect 324 -1216 325 -1215
rect 436 -1216 437 -1215
rect 513 -1216 514 -1215
rect 681 -1216 682 -1215
rect 709 -1216 710 -1215
rect 324 -1218 325 -1217
rect 387 -1218 388 -1217
rect 436 -1218 437 -1217
rect 492 -1218 493 -1217
rect 632 -1218 633 -1217
rect 709 -1218 710 -1217
rect 492 -1220 493 -1219
rect 723 -1220 724 -1219
rect 576 -1222 577 -1221
rect 632 -1222 633 -1221
rect 702 -1222 703 -1221
rect 954 -1222 955 -1221
rect 366 -1224 367 -1223
rect 576 -1224 577 -1223
rect 366 -1226 367 -1225
rect 373 -1226 374 -1225
rect 415 -1226 416 -1225
rect 702 -1226 703 -1225
rect 415 -1228 416 -1227
rect 828 -1228 829 -1227
rect 30 -1239 31 -1238
rect 565 -1239 566 -1238
rect 569 -1239 570 -1238
rect 726 -1239 727 -1238
rect 772 -1239 773 -1238
rect 821 -1239 822 -1238
rect 828 -1239 829 -1238
rect 1017 -1239 1018 -1238
rect 47 -1241 48 -1240
rect 177 -1241 178 -1240
rect 180 -1241 181 -1240
rect 464 -1241 465 -1240
rect 481 -1241 482 -1240
rect 863 -1241 864 -1240
rect 866 -1241 867 -1240
rect 905 -1241 906 -1240
rect 999 -1241 1000 -1240
rect 1031 -1241 1032 -1240
rect 68 -1243 69 -1242
rect 72 -1243 73 -1242
rect 86 -1243 87 -1242
rect 163 -1243 164 -1242
rect 177 -1243 178 -1242
rect 205 -1243 206 -1242
rect 212 -1243 213 -1242
rect 390 -1243 391 -1242
rect 394 -1243 395 -1242
rect 775 -1243 776 -1242
rect 807 -1243 808 -1242
rect 1031 -1243 1032 -1242
rect 72 -1245 73 -1244
rect 387 -1245 388 -1244
rect 394 -1245 395 -1244
rect 467 -1245 468 -1244
rect 509 -1245 510 -1244
rect 534 -1245 535 -1244
rect 541 -1245 542 -1244
rect 579 -1245 580 -1244
rect 590 -1245 591 -1244
rect 1059 -1245 1060 -1244
rect 93 -1247 94 -1246
rect 96 -1247 97 -1246
rect 114 -1247 115 -1246
rect 128 -1247 129 -1246
rect 149 -1247 150 -1246
rect 562 -1247 563 -1246
rect 590 -1247 591 -1246
rect 618 -1247 619 -1246
rect 642 -1247 643 -1246
rect 835 -1247 836 -1246
rect 905 -1247 906 -1246
rect 1052 -1247 1053 -1246
rect 1059 -1247 1060 -1246
rect 1115 -1247 1116 -1246
rect 16 -1249 17 -1248
rect 149 -1249 150 -1248
rect 163 -1249 164 -1248
rect 289 -1249 290 -1248
rect 324 -1249 325 -1248
rect 380 -1249 381 -1248
rect 387 -1249 388 -1248
rect 408 -1249 409 -1248
rect 443 -1249 444 -1248
rect 478 -1249 479 -1248
rect 544 -1249 545 -1248
rect 947 -1249 948 -1248
rect 1017 -1249 1018 -1248
rect 1073 -1249 1074 -1248
rect 117 -1251 118 -1250
rect 212 -1251 213 -1250
rect 233 -1251 234 -1250
rect 502 -1251 503 -1250
rect 548 -1251 549 -1250
rect 1024 -1251 1025 -1250
rect 1052 -1251 1053 -1250
rect 1097 -1251 1098 -1250
rect 128 -1253 129 -1252
rect 198 -1253 199 -1252
rect 205 -1253 206 -1252
rect 254 -1253 255 -1252
rect 264 -1253 265 -1252
rect 352 -1253 353 -1252
rect 373 -1253 374 -1252
rect 555 -1253 556 -1252
rect 618 -1253 619 -1252
rect 639 -1253 640 -1252
rect 656 -1253 657 -1252
rect 961 -1253 962 -1252
rect 184 -1255 185 -1254
rect 261 -1255 262 -1254
rect 289 -1255 290 -1254
rect 296 -1255 297 -1254
rect 324 -1255 325 -1254
rect 422 -1255 423 -1254
rect 478 -1255 479 -1254
rect 604 -1255 605 -1254
rect 639 -1255 640 -1254
rect 667 -1255 668 -1254
rect 677 -1255 678 -1254
rect 730 -1255 731 -1254
rect 796 -1255 797 -1254
rect 947 -1255 948 -1254
rect 961 -1255 962 -1254
rect 1087 -1255 1088 -1254
rect 184 -1257 185 -1256
rect 226 -1257 227 -1256
rect 233 -1257 234 -1256
rect 310 -1257 311 -1256
rect 341 -1257 342 -1256
rect 583 -1257 584 -1256
rect 604 -1257 605 -1256
rect 646 -1257 647 -1256
rect 656 -1257 657 -1256
rect 737 -1257 738 -1256
rect 807 -1257 808 -1256
rect 877 -1257 878 -1256
rect 1087 -1257 1088 -1256
rect 1122 -1257 1123 -1256
rect 156 -1259 157 -1258
rect 226 -1259 227 -1258
rect 240 -1259 241 -1258
rect 446 -1259 447 -1258
rect 506 -1259 507 -1258
rect 555 -1259 556 -1258
rect 572 -1259 573 -1258
rect 737 -1259 738 -1258
rect 821 -1259 822 -1258
rect 1062 -1259 1063 -1258
rect 152 -1261 153 -1260
rect 156 -1261 157 -1260
rect 191 -1261 192 -1260
rect 320 -1261 321 -1260
rect 345 -1261 346 -1260
rect 380 -1261 381 -1260
rect 404 -1261 405 -1260
rect 429 -1261 430 -1260
rect 506 -1261 507 -1260
rect 527 -1261 528 -1260
rect 548 -1261 549 -1260
rect 597 -1261 598 -1260
rect 646 -1261 647 -1260
rect 674 -1261 675 -1260
rect 709 -1261 710 -1260
rect 996 -1261 997 -1260
rect 198 -1263 199 -1262
rect 240 -1263 241 -1262
rect 254 -1263 255 -1262
rect 268 -1263 269 -1262
rect 282 -1263 283 -1262
rect 345 -1263 346 -1262
rect 352 -1263 353 -1262
rect 576 -1263 577 -1262
rect 583 -1263 584 -1262
rect 674 -1263 675 -1262
rect 709 -1263 710 -1262
rect 814 -1263 815 -1262
rect 828 -1263 829 -1262
rect 912 -1263 913 -1262
rect 121 -1265 122 -1264
rect 282 -1265 283 -1264
rect 296 -1265 297 -1264
rect 303 -1265 304 -1264
rect 310 -1265 311 -1264
rect 632 -1265 633 -1264
rect 660 -1265 661 -1264
rect 670 -1265 671 -1264
rect 723 -1265 724 -1264
rect 1066 -1265 1067 -1264
rect 107 -1267 108 -1266
rect 121 -1267 122 -1266
rect 268 -1267 269 -1266
rect 275 -1267 276 -1266
rect 317 -1267 318 -1266
rect 572 -1267 573 -1266
rect 660 -1267 661 -1266
rect 681 -1267 682 -1266
rect 723 -1267 724 -1266
rect 758 -1267 759 -1266
rect 814 -1267 815 -1266
rect 978 -1267 979 -1266
rect 1066 -1267 1067 -1266
rect 1108 -1267 1109 -1266
rect 79 -1269 80 -1268
rect 275 -1269 276 -1268
rect 366 -1269 367 -1268
rect 527 -1269 528 -1268
rect 663 -1269 664 -1268
rect 793 -1269 794 -1268
rect 835 -1269 836 -1268
rect 849 -1269 850 -1268
rect 877 -1269 878 -1268
rect 940 -1269 941 -1268
rect 79 -1271 80 -1270
rect 135 -1271 136 -1270
rect 247 -1271 248 -1270
rect 317 -1271 318 -1270
rect 376 -1271 377 -1270
rect 471 -1271 472 -1270
rect 667 -1271 668 -1270
rect 702 -1271 703 -1270
rect 730 -1271 731 -1270
rect 779 -1271 780 -1270
rect 793 -1271 794 -1270
rect 898 -1271 899 -1270
rect 912 -1271 913 -1270
rect 1045 -1271 1046 -1270
rect 37 -1273 38 -1272
rect 135 -1273 136 -1272
rect 247 -1273 248 -1272
rect 359 -1273 360 -1272
rect 408 -1273 409 -1272
rect 450 -1273 451 -1272
rect 464 -1273 465 -1272
rect 898 -1273 899 -1272
rect 940 -1273 941 -1272
rect 1038 -1273 1039 -1272
rect 1045 -1273 1046 -1272
rect 1094 -1273 1095 -1272
rect 107 -1275 108 -1274
rect 170 -1275 171 -1274
rect 359 -1275 360 -1274
rect 492 -1275 493 -1274
rect 670 -1275 671 -1274
rect 681 -1275 682 -1274
rect 702 -1275 703 -1274
rect 716 -1275 717 -1274
rect 751 -1275 752 -1274
rect 758 -1275 759 -1274
rect 779 -1275 780 -1274
rect 884 -1275 885 -1274
rect 142 -1277 143 -1276
rect 170 -1277 171 -1276
rect 338 -1277 339 -1276
rect 492 -1277 493 -1276
rect 695 -1277 696 -1276
rect 716 -1277 717 -1276
rect 751 -1277 752 -1276
rect 765 -1277 766 -1276
rect 849 -1277 850 -1276
rect 919 -1277 920 -1276
rect 142 -1279 143 -1278
rect 331 -1279 332 -1278
rect 338 -1279 339 -1278
rect 366 -1279 367 -1278
rect 415 -1279 416 -1278
rect 471 -1279 472 -1278
rect 695 -1279 696 -1278
rect 744 -1279 745 -1278
rect 765 -1279 766 -1278
rect 954 -1279 955 -1278
rect 303 -1281 304 -1280
rect 331 -1281 332 -1280
rect 401 -1281 402 -1280
rect 415 -1281 416 -1280
rect 429 -1281 430 -1280
rect 457 -1281 458 -1280
rect 688 -1281 689 -1280
rect 744 -1281 745 -1280
rect 856 -1281 857 -1280
rect 1038 -1281 1039 -1280
rect 44 -1283 45 -1282
rect 401 -1283 402 -1282
rect 436 -1283 437 -1282
rect 457 -1283 458 -1282
rect 688 -1283 689 -1282
rect 786 -1283 787 -1282
rect 856 -1283 857 -1282
rect 933 -1283 934 -1282
rect 954 -1283 955 -1282
rect 982 -1283 983 -1282
rect 44 -1285 45 -1284
rect 51 -1285 52 -1284
rect 436 -1285 437 -1284
rect 520 -1285 521 -1284
rect 786 -1285 787 -1284
rect 842 -1285 843 -1284
rect 884 -1285 885 -1284
rect 1027 -1285 1028 -1284
rect 450 -1287 451 -1286
rect 485 -1287 486 -1286
rect 520 -1287 521 -1286
rect 611 -1287 612 -1286
rect 842 -1287 843 -1286
rect 926 -1287 927 -1286
rect 933 -1287 934 -1286
rect 1003 -1287 1004 -1286
rect 485 -1289 486 -1288
rect 513 -1289 514 -1288
rect 562 -1289 563 -1288
rect 611 -1289 612 -1288
rect 891 -1289 892 -1288
rect 982 -1289 983 -1288
rect 1003 -1289 1004 -1288
rect 1010 -1289 1011 -1288
rect 499 -1291 500 -1290
rect 513 -1291 514 -1290
rect 800 -1291 801 -1290
rect 1010 -1291 1011 -1290
rect 422 -1293 423 -1292
rect 499 -1293 500 -1292
rect 800 -1293 801 -1292
rect 870 -1293 871 -1292
rect 891 -1293 892 -1292
rect 989 -1293 990 -1292
rect 870 -1295 871 -1294
rect 968 -1295 969 -1294
rect 989 -1295 990 -1294
rect 1080 -1295 1081 -1294
rect 926 -1297 927 -1296
rect 1024 -1297 1025 -1296
rect 1080 -1297 1081 -1296
rect 1129 -1297 1130 -1296
rect 968 -1299 969 -1298
rect 975 -1299 976 -1298
rect 9 -1310 10 -1309
rect 30 -1310 31 -1309
rect 37 -1310 38 -1309
rect 114 -1310 115 -1309
rect 135 -1310 136 -1309
rect 369 -1310 370 -1309
rect 408 -1310 409 -1309
rect 481 -1310 482 -1309
rect 499 -1310 500 -1309
rect 513 -1310 514 -1309
rect 534 -1310 535 -1309
rect 590 -1310 591 -1309
rect 611 -1310 612 -1309
rect 625 -1310 626 -1309
rect 628 -1310 629 -1309
rect 919 -1310 920 -1309
rect 922 -1310 923 -1309
rect 968 -1310 969 -1309
rect 975 -1310 976 -1309
rect 982 -1310 983 -1309
rect 996 -1310 997 -1309
rect 1003 -1310 1004 -1309
rect 1020 -1310 1021 -1309
rect 1066 -1310 1067 -1309
rect 1097 -1310 1098 -1309
rect 1101 -1310 1102 -1309
rect 16 -1312 17 -1311
rect 72 -1312 73 -1311
rect 93 -1312 94 -1311
rect 100 -1312 101 -1311
rect 114 -1312 115 -1311
rect 201 -1312 202 -1311
rect 212 -1312 213 -1311
rect 338 -1312 339 -1311
rect 380 -1312 381 -1311
rect 590 -1312 591 -1311
rect 614 -1312 615 -1311
rect 751 -1312 752 -1311
rect 793 -1312 794 -1311
rect 1010 -1312 1011 -1311
rect 1059 -1312 1060 -1311
rect 1087 -1312 1088 -1311
rect 23 -1314 24 -1313
rect 240 -1314 241 -1313
rect 261 -1314 262 -1313
rect 348 -1314 349 -1313
rect 380 -1314 381 -1313
rect 422 -1314 423 -1313
rect 429 -1314 430 -1313
rect 464 -1314 465 -1313
rect 471 -1314 472 -1313
rect 513 -1314 514 -1313
rect 527 -1314 528 -1313
rect 751 -1314 752 -1313
rect 793 -1314 794 -1313
rect 1031 -1314 1032 -1313
rect 1066 -1314 1067 -1313
rect 1080 -1314 1081 -1313
rect 51 -1316 52 -1315
rect 247 -1316 248 -1315
rect 268 -1316 269 -1315
rect 303 -1316 304 -1315
rect 310 -1316 311 -1315
rect 597 -1316 598 -1315
rect 625 -1316 626 -1315
rect 702 -1316 703 -1315
rect 726 -1316 727 -1315
rect 1024 -1316 1025 -1315
rect 1031 -1316 1032 -1315
rect 1052 -1316 1053 -1315
rect 58 -1318 59 -1317
rect 537 -1318 538 -1317
rect 555 -1318 556 -1317
rect 569 -1318 570 -1317
rect 576 -1318 577 -1317
rect 600 -1318 601 -1317
rect 653 -1318 654 -1317
rect 744 -1318 745 -1317
rect 863 -1318 864 -1317
rect 940 -1318 941 -1317
rect 961 -1318 962 -1317
rect 1010 -1318 1011 -1317
rect 68 -1320 69 -1319
rect 306 -1320 307 -1319
rect 408 -1320 409 -1319
rect 485 -1320 486 -1319
rect 492 -1320 493 -1319
rect 534 -1320 535 -1319
rect 541 -1320 542 -1319
rect 555 -1320 556 -1319
rect 597 -1320 598 -1319
rect 604 -1320 605 -1319
rect 677 -1320 678 -1319
rect 702 -1320 703 -1319
rect 709 -1320 710 -1319
rect 744 -1320 745 -1319
rect 821 -1320 822 -1319
rect 863 -1320 864 -1319
rect 905 -1320 906 -1319
rect 968 -1320 969 -1319
rect 999 -1320 1000 -1319
rect 1045 -1320 1046 -1319
rect 72 -1322 73 -1321
rect 544 -1322 545 -1321
rect 569 -1322 570 -1321
rect 604 -1322 605 -1321
rect 681 -1322 682 -1321
rect 709 -1322 710 -1321
rect 733 -1322 734 -1321
rect 765 -1322 766 -1321
rect 870 -1322 871 -1321
rect 905 -1322 906 -1321
rect 912 -1322 913 -1321
rect 975 -1322 976 -1321
rect 93 -1324 94 -1323
rect 481 -1324 482 -1323
rect 506 -1324 507 -1323
rect 632 -1324 633 -1323
rect 737 -1324 738 -1323
rect 740 -1324 741 -1323
rect 758 -1324 759 -1323
rect 821 -1324 822 -1323
rect 870 -1324 871 -1323
rect 884 -1324 885 -1323
rect 891 -1324 892 -1323
rect 912 -1324 913 -1323
rect 933 -1324 934 -1323
rect 961 -1324 962 -1323
rect 100 -1326 101 -1325
rect 352 -1326 353 -1325
rect 411 -1326 412 -1325
rect 681 -1326 682 -1325
rect 723 -1326 724 -1325
rect 758 -1326 759 -1325
rect 765 -1326 766 -1325
rect 786 -1326 787 -1325
rect 877 -1326 878 -1325
rect 884 -1326 885 -1325
rect 891 -1326 892 -1325
rect 1017 -1326 1018 -1325
rect 128 -1328 129 -1327
rect 261 -1328 262 -1327
rect 268 -1328 269 -1327
rect 296 -1328 297 -1327
rect 345 -1328 346 -1327
rect 352 -1328 353 -1327
rect 422 -1328 423 -1327
rect 443 -1328 444 -1327
rect 471 -1328 472 -1327
rect 520 -1328 521 -1327
rect 527 -1328 528 -1327
rect 583 -1328 584 -1327
rect 660 -1328 661 -1327
rect 1017 -1328 1018 -1327
rect 86 -1330 87 -1329
rect 296 -1330 297 -1329
rect 345 -1330 346 -1329
rect 982 -1330 983 -1329
rect 86 -1332 87 -1331
rect 275 -1332 276 -1331
rect 285 -1332 286 -1331
rect 485 -1332 486 -1331
rect 506 -1332 507 -1331
rect 1003 -1332 1004 -1331
rect 128 -1334 129 -1333
rect 359 -1334 360 -1333
rect 366 -1334 367 -1333
rect 443 -1334 444 -1333
rect 520 -1334 521 -1333
rect 674 -1334 675 -1333
rect 716 -1334 717 -1333
rect 786 -1334 787 -1333
rect 856 -1334 857 -1333
rect 877 -1334 878 -1333
rect 933 -1334 934 -1333
rect 947 -1334 948 -1333
rect 79 -1336 80 -1335
rect 359 -1336 360 -1335
rect 366 -1336 367 -1335
rect 401 -1336 402 -1335
rect 429 -1336 430 -1335
rect 450 -1336 451 -1335
rect 572 -1336 573 -1335
rect 674 -1336 675 -1335
rect 688 -1336 689 -1335
rect 716 -1336 717 -1335
rect 723 -1336 724 -1335
rect 849 -1336 850 -1335
rect 856 -1336 857 -1335
rect 1038 -1336 1039 -1335
rect 79 -1338 80 -1337
rect 184 -1338 185 -1337
rect 191 -1338 192 -1337
rect 205 -1338 206 -1337
rect 212 -1338 213 -1337
rect 278 -1338 279 -1337
rect 415 -1338 416 -1337
rect 450 -1338 451 -1337
rect 572 -1338 573 -1337
rect 730 -1338 731 -1337
rect 737 -1338 738 -1337
rect 772 -1338 773 -1337
rect 835 -1338 836 -1337
rect 849 -1338 850 -1337
rect 926 -1338 927 -1337
rect 947 -1338 948 -1337
rect 170 -1340 171 -1339
rect 240 -1340 241 -1339
rect 254 -1340 255 -1339
rect 303 -1340 304 -1339
rect 310 -1340 311 -1339
rect 730 -1340 731 -1339
rect 740 -1340 741 -1339
rect 772 -1340 773 -1339
rect 926 -1340 927 -1339
rect 954 -1340 955 -1339
rect 163 -1342 164 -1341
rect 170 -1342 171 -1341
rect 177 -1342 178 -1341
rect 205 -1342 206 -1341
rect 254 -1342 255 -1341
rect 478 -1342 479 -1341
rect 583 -1342 584 -1341
rect 618 -1342 619 -1341
rect 646 -1342 647 -1341
rect 688 -1342 689 -1341
rect 954 -1342 955 -1341
rect 989 -1342 990 -1341
rect 107 -1344 108 -1343
rect 163 -1344 164 -1343
rect 177 -1344 178 -1343
rect 415 -1344 416 -1343
rect 436 -1344 437 -1343
rect 464 -1344 465 -1343
rect 478 -1344 479 -1343
rect 548 -1344 549 -1343
rect 618 -1344 619 -1343
rect 639 -1344 640 -1343
rect 646 -1344 647 -1343
rect 940 -1344 941 -1343
rect 107 -1346 108 -1345
rect 135 -1346 136 -1345
rect 180 -1346 181 -1345
rect 226 -1346 227 -1345
rect 275 -1346 276 -1345
rect 562 -1346 563 -1345
rect 660 -1346 661 -1345
rect 779 -1346 780 -1345
rect 898 -1346 899 -1345
rect 989 -1346 990 -1345
rect 65 -1348 66 -1347
rect 562 -1348 563 -1347
rect 779 -1348 780 -1347
rect 800 -1348 801 -1347
rect 184 -1350 185 -1349
rect 198 -1350 199 -1349
rect 226 -1350 227 -1349
rect 233 -1350 234 -1349
rect 394 -1350 395 -1349
rect 898 -1350 899 -1349
rect 194 -1352 195 -1351
rect 219 -1352 220 -1351
rect 233 -1352 234 -1351
rect 317 -1352 318 -1351
rect 373 -1352 374 -1351
rect 394 -1352 395 -1351
rect 436 -1352 437 -1351
rect 457 -1352 458 -1351
rect 467 -1352 468 -1351
rect 639 -1352 640 -1351
rect 800 -1352 801 -1351
rect 807 -1352 808 -1351
rect 121 -1354 122 -1353
rect 219 -1354 220 -1353
rect 341 -1354 342 -1353
rect 457 -1354 458 -1353
rect 548 -1354 549 -1353
rect 796 -1354 797 -1353
rect 807 -1354 808 -1353
rect 814 -1354 815 -1353
rect 121 -1356 122 -1355
rect 149 -1356 150 -1355
rect 198 -1356 199 -1355
rect 324 -1356 325 -1355
rect 373 -1356 374 -1355
rect 541 -1356 542 -1355
rect 814 -1356 815 -1355
rect 828 -1356 829 -1355
rect 142 -1358 143 -1357
rect 317 -1358 318 -1357
rect 439 -1358 440 -1357
rect 576 -1358 577 -1357
rect 828 -1358 829 -1357
rect 842 -1358 843 -1357
rect 142 -1360 143 -1359
rect 835 -1360 836 -1359
rect 149 -1362 150 -1361
rect 156 -1362 157 -1361
rect 282 -1362 283 -1361
rect 324 -1362 325 -1361
rect 635 -1362 636 -1361
rect 842 -1362 843 -1361
rect 156 -1364 157 -1363
rect 387 -1364 388 -1363
rect 331 -1366 332 -1365
rect 387 -1366 388 -1365
rect 289 -1368 290 -1367
rect 331 -1368 332 -1367
rect 289 -1370 290 -1369
rect 404 -1370 405 -1369
rect 2 -1381 3 -1380
rect 5 -1381 6 -1380
rect 9 -1381 10 -1380
rect 114 -1381 115 -1380
rect 142 -1381 143 -1380
rect 240 -1381 241 -1380
rect 250 -1381 251 -1380
rect 268 -1381 269 -1380
rect 369 -1381 370 -1380
rect 674 -1381 675 -1380
rect 702 -1381 703 -1380
rect 730 -1381 731 -1380
rect 996 -1381 997 -1380
rect 1059 -1381 1060 -1380
rect 30 -1383 31 -1382
rect 33 -1383 34 -1382
rect 72 -1383 73 -1382
rect 275 -1383 276 -1382
rect 369 -1383 370 -1382
rect 520 -1383 521 -1382
rect 530 -1383 531 -1382
rect 786 -1383 787 -1382
rect 947 -1383 948 -1382
rect 996 -1383 997 -1382
rect 1003 -1383 1004 -1382
rect 1024 -1383 1025 -1382
rect 1031 -1383 1032 -1382
rect 1038 -1383 1039 -1382
rect 1045 -1383 1046 -1382
rect 1066 -1383 1067 -1382
rect 30 -1385 31 -1384
rect 44 -1385 45 -1384
rect 72 -1385 73 -1384
rect 201 -1385 202 -1384
rect 208 -1385 209 -1384
rect 590 -1385 591 -1384
rect 618 -1385 619 -1384
rect 625 -1385 626 -1384
rect 632 -1385 633 -1384
rect 674 -1385 675 -1384
rect 681 -1385 682 -1384
rect 947 -1385 948 -1384
rect 975 -1385 976 -1384
rect 1003 -1385 1004 -1384
rect 1010 -1385 1011 -1384
rect 1031 -1385 1032 -1384
rect 1055 -1385 1056 -1384
rect 1066 -1385 1067 -1384
rect 33 -1387 34 -1386
rect 44 -1387 45 -1386
rect 79 -1387 80 -1386
rect 268 -1387 269 -1386
rect 380 -1387 381 -1386
rect 436 -1387 437 -1386
rect 443 -1387 444 -1386
rect 478 -1387 479 -1386
rect 488 -1387 489 -1386
rect 506 -1387 507 -1386
rect 509 -1387 510 -1386
rect 562 -1387 563 -1386
rect 646 -1387 647 -1386
rect 758 -1387 759 -1386
rect 786 -1387 787 -1386
rect 814 -1387 815 -1386
rect 940 -1387 941 -1386
rect 975 -1387 976 -1386
rect 982 -1387 983 -1386
rect 1010 -1387 1011 -1386
rect 79 -1389 80 -1388
rect 121 -1389 122 -1388
rect 128 -1389 129 -1388
rect 436 -1389 437 -1388
rect 457 -1389 458 -1388
rect 492 -1389 493 -1388
rect 499 -1389 500 -1388
rect 544 -1389 545 -1388
rect 555 -1389 556 -1388
rect 618 -1389 619 -1388
rect 653 -1389 654 -1388
rect 989 -1389 990 -1388
rect 86 -1391 87 -1390
rect 474 -1391 475 -1390
rect 513 -1391 514 -1390
rect 562 -1391 563 -1390
rect 569 -1391 570 -1390
rect 940 -1391 941 -1390
rect 961 -1391 962 -1390
rect 989 -1391 990 -1390
rect 86 -1393 87 -1392
rect 345 -1393 346 -1392
rect 366 -1393 367 -1392
rect 653 -1393 654 -1392
rect 660 -1393 661 -1392
rect 793 -1393 794 -1392
rect 912 -1393 913 -1392
rect 961 -1393 962 -1392
rect 100 -1395 101 -1394
rect 107 -1395 108 -1394
rect 114 -1395 115 -1394
rect 156 -1395 157 -1394
rect 177 -1395 178 -1394
rect 191 -1395 192 -1394
rect 198 -1395 199 -1394
rect 247 -1395 248 -1394
rect 261 -1395 262 -1394
rect 285 -1395 286 -1394
rect 289 -1395 290 -1394
rect 982 -1395 983 -1394
rect 93 -1397 94 -1396
rect 289 -1397 290 -1396
rect 380 -1397 381 -1396
rect 401 -1397 402 -1396
rect 408 -1397 409 -1396
rect 492 -1397 493 -1396
rect 534 -1397 535 -1396
rect 590 -1397 591 -1396
rect 604 -1397 605 -1396
rect 646 -1397 647 -1396
rect 667 -1397 668 -1396
rect 681 -1397 682 -1396
rect 702 -1397 703 -1396
rect 772 -1397 773 -1396
rect 793 -1397 794 -1396
rect 814 -1397 815 -1396
rect 912 -1397 913 -1396
rect 926 -1397 927 -1396
rect 16 -1399 17 -1398
rect 93 -1399 94 -1398
rect 121 -1399 122 -1398
rect 523 -1399 524 -1398
rect 537 -1399 538 -1398
rect 821 -1399 822 -1398
rect 842 -1399 843 -1398
rect 926 -1399 927 -1398
rect 128 -1401 129 -1400
rect 898 -1401 899 -1400
rect 142 -1403 143 -1402
rect 170 -1403 171 -1402
rect 212 -1403 213 -1402
rect 401 -1403 402 -1402
rect 408 -1403 409 -1402
rect 656 -1403 657 -1402
rect 667 -1403 668 -1402
rect 751 -1403 752 -1402
rect 772 -1403 773 -1402
rect 800 -1403 801 -1402
rect 821 -1403 822 -1402
rect 919 -1403 920 -1402
rect 58 -1405 59 -1404
rect 170 -1405 171 -1404
rect 219 -1405 220 -1404
rect 261 -1405 262 -1404
rect 345 -1405 346 -1404
rect 534 -1405 535 -1404
rect 541 -1405 542 -1404
rect 968 -1405 969 -1404
rect 156 -1407 157 -1406
rect 548 -1407 549 -1406
rect 569 -1407 570 -1406
rect 723 -1407 724 -1406
rect 726 -1407 727 -1406
rect 933 -1407 934 -1406
rect 135 -1409 136 -1408
rect 548 -1409 549 -1408
rect 663 -1409 664 -1408
rect 968 -1409 969 -1408
rect 205 -1411 206 -1410
rect 219 -1411 220 -1410
rect 226 -1411 227 -1410
rect 376 -1411 377 -1410
rect 415 -1411 416 -1410
rect 443 -1411 444 -1410
rect 450 -1411 451 -1410
rect 499 -1411 500 -1410
rect 541 -1411 542 -1410
rect 744 -1411 745 -1410
rect 751 -1411 752 -1410
rect 765 -1411 766 -1410
rect 828 -1411 829 -1410
rect 842 -1411 843 -1410
rect 891 -1411 892 -1410
rect 898 -1411 899 -1410
rect 905 -1411 906 -1410
rect 919 -1411 920 -1410
rect 107 -1413 108 -1412
rect 205 -1413 206 -1412
rect 226 -1413 227 -1412
rect 254 -1413 255 -1412
rect 366 -1413 367 -1412
rect 933 -1413 934 -1412
rect 233 -1415 234 -1414
rect 1052 -1415 1053 -1414
rect 51 -1417 52 -1416
rect 233 -1417 234 -1416
rect 240 -1417 241 -1416
rect 338 -1417 339 -1416
rect 415 -1417 416 -1416
rect 422 -1417 423 -1416
rect 439 -1417 440 -1416
rect 555 -1417 556 -1416
rect 597 -1417 598 -1416
rect 744 -1417 745 -1416
rect 796 -1417 797 -1416
rect 905 -1417 906 -1416
rect 51 -1419 52 -1418
rect 387 -1419 388 -1418
rect 450 -1419 451 -1418
rect 807 -1419 808 -1418
rect 828 -1419 829 -1418
rect 884 -1419 885 -1418
rect 58 -1421 59 -1420
rect 422 -1421 423 -1420
rect 471 -1421 472 -1420
rect 513 -1421 514 -1420
rect 520 -1421 521 -1420
rect 597 -1421 598 -1420
rect 695 -1421 696 -1420
rect 723 -1421 724 -1420
rect 779 -1421 780 -1420
rect 807 -1421 808 -1420
rect 877 -1421 878 -1420
rect 884 -1421 885 -1420
rect 247 -1423 248 -1422
rect 303 -1423 304 -1422
rect 310 -1423 311 -1422
rect 338 -1423 339 -1422
rect 387 -1423 388 -1422
rect 527 -1423 528 -1422
rect 688 -1423 689 -1422
rect 695 -1423 696 -1422
rect 709 -1423 710 -1422
rect 800 -1423 801 -1422
rect 870 -1423 871 -1422
rect 877 -1423 878 -1422
rect 254 -1425 255 -1424
rect 485 -1425 486 -1424
rect 527 -1425 528 -1424
rect 835 -1425 836 -1424
rect 863 -1425 864 -1424
rect 870 -1425 871 -1424
rect 138 -1427 139 -1426
rect 863 -1427 864 -1426
rect 303 -1429 304 -1428
rect 317 -1429 318 -1428
rect 348 -1429 349 -1428
rect 835 -1429 836 -1428
rect 310 -1431 311 -1430
rect 331 -1431 332 -1430
rect 464 -1431 465 -1430
rect 485 -1431 486 -1430
rect 628 -1431 629 -1430
rect 709 -1431 710 -1430
rect 716 -1431 717 -1430
rect 758 -1431 759 -1430
rect 779 -1431 780 -1430
rect 856 -1431 857 -1430
rect 331 -1433 332 -1432
rect 352 -1433 353 -1432
rect 359 -1433 360 -1432
rect 464 -1433 465 -1432
rect 576 -1433 577 -1432
rect 856 -1433 857 -1432
rect 23 -1435 24 -1434
rect 352 -1435 353 -1434
rect 460 -1435 461 -1434
rect 716 -1435 717 -1434
rect 23 -1437 24 -1436
rect 163 -1437 164 -1436
rect 324 -1437 325 -1436
rect 359 -1437 360 -1436
rect 576 -1437 577 -1436
rect 583 -1437 584 -1436
rect 639 -1437 640 -1436
rect 688 -1437 689 -1436
rect 163 -1439 164 -1438
rect 184 -1439 185 -1438
rect 296 -1439 297 -1438
rect 324 -1439 325 -1438
rect 583 -1439 584 -1438
rect 1048 -1439 1049 -1438
rect 37 -1441 38 -1440
rect 184 -1441 185 -1440
rect 296 -1441 297 -1440
rect 373 -1441 374 -1440
rect 639 -1441 640 -1440
rect 1017 -1441 1018 -1440
rect 373 -1443 374 -1442
rect 891 -1443 892 -1442
rect 954 -1443 955 -1442
rect 1017 -1443 1018 -1442
rect 495 -1445 496 -1444
rect 954 -1445 955 -1444
rect 2 -1456 3 -1455
rect 37 -1456 38 -1455
rect 68 -1456 69 -1455
rect 394 -1456 395 -1455
rect 422 -1456 423 -1455
rect 814 -1456 815 -1455
rect 824 -1456 825 -1455
rect 1024 -1456 1025 -1455
rect 1045 -1456 1046 -1455
rect 1059 -1456 1060 -1455
rect 9 -1458 10 -1457
rect 128 -1458 129 -1457
rect 142 -1458 143 -1457
rect 285 -1458 286 -1457
rect 310 -1458 311 -1457
rect 317 -1458 318 -1457
rect 348 -1458 349 -1457
rect 443 -1458 444 -1457
rect 457 -1458 458 -1457
rect 982 -1458 983 -1457
rect 999 -1458 1000 -1457
rect 1038 -1458 1039 -1457
rect 1048 -1458 1049 -1457
rect 1052 -1458 1053 -1457
rect 1059 -1458 1060 -1457
rect 1066 -1458 1067 -1457
rect 19 -1460 20 -1459
rect 58 -1460 59 -1459
rect 72 -1460 73 -1459
rect 138 -1460 139 -1459
rect 142 -1460 143 -1459
rect 177 -1460 178 -1459
rect 184 -1460 185 -1459
rect 310 -1460 311 -1459
rect 352 -1460 353 -1459
rect 460 -1460 461 -1459
rect 506 -1460 507 -1459
rect 537 -1460 538 -1459
rect 593 -1460 594 -1459
rect 845 -1460 846 -1459
rect 982 -1460 983 -1459
rect 1031 -1460 1032 -1459
rect 23 -1462 24 -1461
rect 352 -1462 353 -1461
rect 387 -1462 388 -1461
rect 474 -1462 475 -1461
rect 509 -1462 510 -1461
rect 618 -1462 619 -1461
rect 625 -1462 626 -1461
rect 628 -1462 629 -1461
rect 632 -1462 633 -1461
rect 681 -1462 682 -1461
rect 684 -1462 685 -1461
rect 933 -1462 934 -1461
rect 23 -1464 24 -1463
rect 425 -1464 426 -1463
rect 436 -1464 437 -1463
rect 968 -1464 969 -1463
rect 30 -1466 31 -1465
rect 40 -1466 41 -1465
rect 72 -1466 73 -1465
rect 562 -1466 563 -1465
rect 604 -1466 605 -1465
rect 611 -1466 612 -1465
rect 625 -1466 626 -1465
rect 716 -1466 717 -1465
rect 744 -1466 745 -1465
rect 747 -1466 748 -1465
rect 765 -1466 766 -1465
rect 863 -1466 864 -1465
rect 37 -1468 38 -1467
rect 44 -1468 45 -1467
rect 93 -1468 94 -1467
rect 422 -1468 423 -1467
rect 436 -1468 437 -1467
rect 464 -1468 465 -1467
rect 520 -1468 521 -1467
rect 758 -1468 759 -1467
rect 765 -1468 766 -1467
rect 870 -1468 871 -1467
rect 44 -1470 45 -1469
rect 408 -1470 409 -1469
rect 443 -1470 444 -1469
rect 569 -1470 570 -1469
rect 607 -1470 608 -1469
rect 947 -1470 948 -1469
rect 58 -1472 59 -1471
rect 408 -1472 409 -1471
rect 450 -1472 451 -1471
rect 537 -1472 538 -1471
rect 611 -1472 612 -1471
rect 674 -1472 675 -1471
rect 681 -1472 682 -1471
rect 926 -1472 927 -1471
rect 93 -1474 94 -1473
rect 177 -1474 178 -1473
rect 191 -1474 192 -1473
rect 478 -1474 479 -1473
rect 520 -1474 521 -1473
rect 940 -1474 941 -1473
rect 96 -1476 97 -1475
rect 758 -1476 759 -1475
rect 768 -1476 769 -1475
rect 828 -1476 829 -1475
rect 856 -1476 857 -1475
rect 870 -1476 871 -1475
rect 926 -1476 927 -1475
rect 975 -1476 976 -1475
rect 128 -1478 129 -1477
rect 303 -1478 304 -1477
rect 345 -1478 346 -1477
rect 450 -1478 451 -1477
rect 464 -1478 465 -1477
rect 513 -1478 514 -1477
rect 534 -1478 535 -1477
rect 548 -1478 549 -1477
rect 635 -1478 636 -1477
rect 660 -1478 661 -1477
rect 667 -1478 668 -1477
rect 674 -1478 675 -1477
rect 709 -1478 710 -1477
rect 947 -1478 948 -1477
rect 975 -1478 976 -1477
rect 996 -1478 997 -1477
rect 163 -1480 164 -1479
rect 184 -1480 185 -1479
rect 191 -1480 192 -1479
rect 240 -1480 241 -1479
rect 247 -1480 248 -1479
rect 376 -1480 377 -1479
rect 387 -1480 388 -1479
rect 653 -1480 654 -1479
rect 660 -1480 661 -1479
rect 667 -1480 668 -1479
rect 709 -1480 710 -1479
rect 737 -1480 738 -1479
rect 744 -1480 745 -1479
rect 779 -1480 780 -1479
rect 793 -1480 794 -1479
rect 961 -1480 962 -1479
rect 163 -1482 164 -1481
rect 198 -1482 199 -1481
rect 215 -1482 216 -1481
rect 569 -1482 570 -1481
rect 639 -1482 640 -1481
rect 702 -1482 703 -1481
rect 772 -1482 773 -1481
rect 779 -1482 780 -1481
rect 793 -1482 794 -1481
rect 842 -1482 843 -1481
rect 856 -1482 857 -1481
rect 898 -1482 899 -1481
rect 170 -1484 171 -1483
rect 205 -1484 206 -1483
rect 226 -1484 227 -1483
rect 247 -1484 248 -1483
rect 268 -1484 269 -1483
rect 275 -1484 276 -1483
rect 282 -1484 283 -1483
rect 324 -1484 325 -1483
rect 373 -1484 374 -1483
rect 940 -1484 941 -1483
rect 107 -1486 108 -1485
rect 226 -1486 227 -1485
rect 233 -1486 234 -1485
rect 324 -1486 325 -1485
rect 373 -1486 374 -1485
rect 488 -1486 489 -1485
rect 544 -1486 545 -1485
rect 961 -1486 962 -1485
rect 107 -1488 108 -1487
rect 527 -1488 528 -1487
rect 548 -1488 549 -1487
rect 576 -1488 577 -1487
rect 639 -1488 640 -1487
rect 695 -1488 696 -1487
rect 702 -1488 703 -1487
rect 726 -1488 727 -1487
rect 772 -1488 773 -1487
rect 807 -1488 808 -1487
rect 814 -1488 815 -1487
rect 884 -1488 885 -1487
rect 898 -1488 899 -1487
rect 919 -1488 920 -1487
rect 68 -1490 69 -1489
rect 884 -1490 885 -1489
rect 114 -1492 115 -1491
rect 268 -1492 269 -1491
rect 275 -1492 276 -1491
rect 359 -1492 360 -1491
rect 394 -1492 395 -1491
rect 555 -1492 556 -1491
rect 642 -1492 643 -1491
rect 863 -1492 864 -1491
rect 79 -1494 80 -1493
rect 114 -1494 115 -1493
rect 121 -1494 122 -1493
rect 170 -1494 171 -1493
rect 194 -1494 195 -1493
rect 212 -1494 213 -1493
rect 233 -1494 234 -1493
rect 331 -1494 332 -1493
rect 359 -1494 360 -1493
rect 401 -1494 402 -1493
rect 478 -1494 479 -1493
rect 597 -1494 598 -1493
rect 653 -1494 654 -1493
rect 688 -1494 689 -1493
rect 695 -1494 696 -1493
rect 740 -1494 741 -1493
rect 796 -1494 797 -1493
rect 828 -1494 829 -1493
rect 842 -1494 843 -1493
rect 1017 -1494 1018 -1493
rect 51 -1496 52 -1495
rect 121 -1496 122 -1495
rect 240 -1496 241 -1495
rect 523 -1496 524 -1495
rect 541 -1496 542 -1495
rect 576 -1496 577 -1495
rect 590 -1496 591 -1495
rect 597 -1496 598 -1495
rect 807 -1496 808 -1495
rect 877 -1496 878 -1495
rect 989 -1496 990 -1495
rect 1017 -1496 1018 -1495
rect 51 -1498 52 -1497
rect 254 -1498 255 -1497
rect 296 -1498 297 -1497
rect 401 -1498 402 -1497
rect 492 -1498 493 -1497
rect 919 -1498 920 -1497
rect 79 -1500 80 -1499
rect 156 -1500 157 -1499
rect 254 -1500 255 -1499
rect 583 -1500 584 -1499
rect 590 -1500 591 -1499
rect 835 -1500 836 -1499
rect 877 -1500 878 -1499
rect 1003 -1500 1004 -1499
rect 86 -1502 87 -1501
rect 156 -1502 157 -1501
rect 278 -1502 279 -1501
rect 492 -1502 493 -1501
rect 506 -1502 507 -1501
rect 835 -1502 836 -1501
rect 905 -1502 906 -1501
rect 989 -1502 990 -1501
rect 86 -1504 87 -1503
rect 135 -1504 136 -1503
rect 296 -1504 297 -1503
rect 457 -1504 458 -1503
rect 516 -1504 517 -1503
rect 688 -1504 689 -1503
rect 747 -1504 748 -1503
rect 1003 -1504 1004 -1503
rect 16 -1506 17 -1505
rect 135 -1506 136 -1505
rect 303 -1506 304 -1505
rect 380 -1506 381 -1505
rect 541 -1506 542 -1505
rect 933 -1506 934 -1505
rect 331 -1508 332 -1507
rect 488 -1508 489 -1507
rect 555 -1508 556 -1507
rect 565 -1508 566 -1507
rect 583 -1508 584 -1507
rect 646 -1508 647 -1507
rect 821 -1508 822 -1507
rect 996 -1508 997 -1507
rect 338 -1510 339 -1509
rect 380 -1510 381 -1509
rect 646 -1510 647 -1509
rect 730 -1510 731 -1509
rect 905 -1510 906 -1509
rect 912 -1510 913 -1509
rect 338 -1512 339 -1511
rect 366 -1512 367 -1511
rect 499 -1512 500 -1511
rect 730 -1512 731 -1511
rect 912 -1512 913 -1511
rect 954 -1512 955 -1511
rect 198 -1514 199 -1513
rect 499 -1514 500 -1513
rect 954 -1514 955 -1513
rect 1010 -1514 1011 -1513
rect 366 -1516 367 -1515
rect 723 -1516 724 -1515
rect 800 -1516 801 -1515
rect 1010 -1516 1011 -1515
rect 723 -1518 724 -1517
rect 968 -1518 969 -1517
rect 800 -1520 801 -1519
rect 849 -1520 850 -1519
rect 849 -1522 850 -1521
rect 891 -1522 892 -1521
rect 471 -1524 472 -1523
rect 891 -1524 892 -1523
rect 289 -1526 290 -1525
rect 471 -1526 472 -1525
rect 30 -1528 31 -1527
rect 289 -1528 290 -1527
rect 23 -1539 24 -1538
rect 135 -1539 136 -1538
rect 152 -1539 153 -1538
rect 961 -1539 962 -1538
rect 1017 -1539 1018 -1538
rect 1024 -1539 1025 -1538
rect 1038 -1539 1039 -1538
rect 1045 -1539 1046 -1538
rect 2 -1541 3 -1540
rect 23 -1541 24 -1540
rect 30 -1541 31 -1540
rect 425 -1541 426 -1540
rect 488 -1541 489 -1540
rect 737 -1541 738 -1540
rect 740 -1541 741 -1540
rect 982 -1541 983 -1540
rect 30 -1543 31 -1542
rect 303 -1543 304 -1542
rect 306 -1543 307 -1542
rect 506 -1543 507 -1542
rect 520 -1543 521 -1542
rect 919 -1543 920 -1542
rect 961 -1543 962 -1542
rect 996 -1543 997 -1542
rect 68 -1545 69 -1544
rect 86 -1545 87 -1544
rect 93 -1545 94 -1544
rect 415 -1545 416 -1544
rect 527 -1545 528 -1544
rect 548 -1545 549 -1544
rect 558 -1545 559 -1544
rect 975 -1545 976 -1544
rect 68 -1547 69 -1546
rect 758 -1547 759 -1546
rect 842 -1547 843 -1546
rect 884 -1547 885 -1546
rect 86 -1549 87 -1548
rect 100 -1549 101 -1548
rect 135 -1549 136 -1548
rect 261 -1549 262 -1548
rect 289 -1549 290 -1548
rect 667 -1549 668 -1548
rect 723 -1549 724 -1548
rect 814 -1549 815 -1548
rect 877 -1549 878 -1548
rect 919 -1549 920 -1548
rect 100 -1551 101 -1550
rect 226 -1551 227 -1550
rect 247 -1551 248 -1550
rect 261 -1551 262 -1550
rect 296 -1551 297 -1550
rect 359 -1551 360 -1550
rect 366 -1551 367 -1550
rect 628 -1551 629 -1550
rect 663 -1551 664 -1550
rect 828 -1551 829 -1550
rect 884 -1551 885 -1550
rect 1003 -1551 1004 -1550
rect 128 -1553 129 -1552
rect 289 -1553 290 -1552
rect 373 -1553 374 -1552
rect 485 -1553 486 -1552
rect 499 -1553 500 -1552
rect 548 -1553 549 -1552
rect 565 -1553 566 -1552
rect 947 -1553 948 -1552
rect 72 -1555 73 -1554
rect 499 -1555 500 -1554
rect 534 -1555 535 -1554
rect 555 -1555 556 -1554
rect 583 -1555 584 -1554
rect 667 -1555 668 -1554
rect 684 -1555 685 -1554
rect 877 -1555 878 -1554
rect 947 -1555 948 -1554
rect 1010 -1555 1011 -1554
rect 16 -1557 17 -1556
rect 72 -1557 73 -1556
rect 121 -1557 122 -1556
rect 128 -1557 129 -1556
rect 156 -1557 157 -1556
rect 313 -1557 314 -1556
rect 359 -1557 360 -1556
rect 565 -1557 566 -1556
rect 583 -1557 584 -1556
rect 695 -1557 696 -1556
rect 726 -1557 727 -1556
rect 898 -1557 899 -1556
rect 121 -1559 122 -1558
rect 275 -1559 276 -1558
rect 366 -1559 367 -1558
rect 555 -1559 556 -1558
rect 590 -1559 591 -1558
rect 828 -1559 829 -1558
rect 898 -1559 899 -1558
rect 933 -1559 934 -1558
rect 44 -1561 45 -1560
rect 275 -1561 276 -1560
rect 373 -1561 374 -1560
rect 537 -1561 538 -1560
rect 541 -1561 542 -1560
rect 611 -1561 612 -1560
rect 618 -1561 619 -1560
rect 653 -1561 654 -1560
rect 737 -1561 738 -1560
rect 821 -1561 822 -1560
rect 44 -1563 45 -1562
rect 142 -1563 143 -1562
rect 156 -1563 157 -1562
rect 338 -1563 339 -1562
rect 355 -1563 356 -1562
rect 653 -1563 654 -1562
rect 758 -1563 759 -1562
rect 800 -1563 801 -1562
rect 814 -1563 815 -1562
rect 863 -1563 864 -1562
rect 107 -1565 108 -1564
rect 338 -1565 339 -1564
rect 380 -1565 381 -1564
rect 415 -1565 416 -1564
rect 590 -1565 591 -1564
rect 639 -1565 640 -1564
rect 800 -1565 801 -1564
rect 807 -1565 808 -1564
rect 821 -1565 822 -1564
rect 849 -1565 850 -1564
rect 863 -1565 864 -1564
rect 912 -1565 913 -1564
rect 142 -1567 143 -1566
rect 149 -1567 150 -1566
rect 170 -1567 171 -1566
rect 695 -1567 696 -1566
rect 807 -1567 808 -1566
rect 870 -1567 871 -1566
rect 912 -1567 913 -1566
rect 989 -1567 990 -1566
rect 177 -1569 178 -1568
rect 380 -1569 381 -1568
rect 387 -1569 388 -1568
rect 513 -1569 514 -1568
rect 576 -1569 577 -1568
rect 639 -1569 640 -1568
rect 660 -1569 661 -1568
rect 849 -1569 850 -1568
rect 870 -1569 871 -1568
rect 926 -1569 927 -1568
rect 177 -1571 178 -1570
rect 191 -1571 192 -1570
rect 201 -1571 202 -1570
rect 310 -1571 311 -1570
rect 401 -1571 402 -1570
rect 464 -1571 465 -1570
rect 478 -1571 479 -1570
rect 513 -1571 514 -1570
rect 562 -1571 563 -1570
rect 926 -1571 927 -1570
rect 191 -1573 192 -1572
rect 205 -1573 206 -1572
rect 212 -1573 213 -1572
rect 296 -1573 297 -1572
rect 394 -1573 395 -1572
rect 478 -1573 479 -1572
rect 576 -1573 577 -1572
rect 632 -1573 633 -1572
rect 660 -1573 661 -1572
rect 688 -1573 689 -1572
rect 205 -1575 206 -1574
rect 233 -1575 234 -1574
rect 240 -1575 241 -1574
rect 355 -1575 356 -1574
rect 401 -1575 402 -1574
rect 429 -1575 430 -1574
rect 569 -1575 570 -1574
rect 632 -1575 633 -1574
rect 688 -1575 689 -1574
rect 709 -1575 710 -1574
rect 163 -1577 164 -1576
rect 233 -1577 234 -1576
rect 240 -1577 241 -1576
rect 422 -1577 423 -1576
rect 429 -1577 430 -1576
rect 457 -1577 458 -1576
rect 604 -1577 605 -1576
rect 625 -1577 626 -1576
rect 709 -1577 710 -1576
rect 744 -1577 745 -1576
rect 58 -1579 59 -1578
rect 163 -1579 164 -1578
rect 212 -1579 213 -1578
rect 219 -1579 220 -1578
rect 247 -1579 248 -1578
rect 282 -1579 283 -1578
rect 345 -1579 346 -1578
rect 394 -1579 395 -1578
rect 408 -1579 409 -1578
rect 702 -1579 703 -1578
rect 744 -1579 745 -1578
rect 779 -1579 780 -1578
rect 58 -1581 59 -1580
rect 173 -1581 174 -1580
rect 408 -1581 409 -1580
rect 443 -1581 444 -1580
rect 450 -1581 451 -1580
rect 457 -1581 458 -1580
rect 597 -1581 598 -1580
rect 779 -1581 780 -1580
rect 51 -1583 52 -1582
rect 450 -1583 451 -1582
rect 618 -1583 619 -1582
rect 674 -1583 675 -1582
rect 702 -1583 703 -1582
rect 940 -1583 941 -1582
rect 51 -1585 52 -1584
rect 572 -1585 573 -1584
rect 716 -1585 717 -1584
rect 940 -1585 941 -1584
rect 114 -1587 115 -1586
rect 219 -1587 220 -1586
rect 387 -1587 388 -1586
rect 597 -1587 598 -1586
rect 716 -1587 717 -1586
rect 751 -1587 752 -1586
rect 107 -1589 108 -1588
rect 114 -1589 115 -1588
rect 117 -1589 118 -1588
rect 282 -1589 283 -1588
rect 411 -1589 412 -1588
rect 730 -1589 731 -1588
rect 751 -1589 752 -1588
rect 786 -1589 787 -1588
rect 443 -1591 444 -1590
rect 530 -1591 531 -1590
rect 730 -1591 731 -1590
rect 772 -1591 773 -1590
rect 786 -1591 787 -1590
rect 856 -1591 857 -1590
rect 492 -1593 493 -1592
rect 674 -1593 675 -1592
rect 765 -1593 766 -1592
rect 772 -1593 773 -1592
rect 856 -1593 857 -1592
rect 936 -1593 937 -1592
rect 331 -1595 332 -1594
rect 492 -1595 493 -1594
rect 765 -1595 766 -1594
rect 793 -1595 794 -1594
rect 317 -1597 318 -1596
rect 331 -1597 332 -1596
rect 793 -1597 794 -1596
rect 835 -1597 836 -1596
rect 268 -1599 269 -1598
rect 317 -1599 318 -1598
rect 835 -1599 836 -1598
rect 891 -1599 892 -1598
rect 254 -1601 255 -1600
rect 268 -1601 269 -1600
rect 891 -1601 892 -1600
rect 954 -1601 955 -1600
rect 254 -1603 255 -1602
rect 509 -1603 510 -1602
rect 905 -1603 906 -1602
rect 954 -1603 955 -1602
rect 905 -1605 906 -1604
rect 968 -1605 969 -1604
rect 30 -1616 31 -1615
rect 355 -1616 356 -1615
rect 366 -1616 367 -1615
rect 527 -1616 528 -1615
rect 530 -1616 531 -1615
rect 779 -1616 780 -1615
rect 926 -1616 927 -1615
rect 936 -1616 937 -1615
rect 954 -1616 955 -1615
rect 968 -1616 969 -1615
rect 1038 -1616 1039 -1615
rect 1045 -1616 1046 -1615
rect 58 -1618 59 -1617
rect 303 -1618 304 -1617
rect 310 -1618 311 -1617
rect 471 -1618 472 -1617
rect 523 -1618 524 -1617
rect 667 -1618 668 -1617
rect 681 -1618 682 -1617
rect 737 -1618 738 -1617
rect 775 -1618 776 -1617
rect 849 -1618 850 -1617
rect 65 -1620 66 -1619
rect 110 -1620 111 -1619
rect 121 -1620 122 -1619
rect 306 -1620 307 -1619
rect 310 -1620 311 -1619
rect 352 -1620 353 -1619
rect 366 -1620 367 -1619
rect 401 -1620 402 -1619
rect 425 -1620 426 -1619
rect 471 -1620 472 -1619
rect 544 -1620 545 -1619
rect 793 -1620 794 -1619
rect 68 -1622 69 -1621
rect 240 -1622 241 -1621
rect 257 -1622 258 -1621
rect 324 -1622 325 -1621
rect 352 -1622 353 -1621
rect 408 -1622 409 -1621
rect 429 -1622 430 -1621
rect 516 -1622 517 -1621
rect 551 -1622 552 -1621
rect 639 -1622 640 -1621
rect 646 -1622 647 -1621
rect 667 -1622 668 -1621
rect 681 -1622 682 -1621
rect 684 -1622 685 -1621
rect 695 -1622 696 -1621
rect 919 -1622 920 -1621
rect 72 -1624 73 -1623
rect 411 -1624 412 -1623
rect 562 -1624 563 -1623
rect 838 -1624 839 -1623
rect 79 -1626 80 -1625
rect 401 -1626 402 -1625
rect 562 -1626 563 -1625
rect 702 -1626 703 -1625
rect 723 -1626 724 -1625
rect 737 -1626 738 -1625
rect 751 -1626 752 -1625
rect 793 -1626 794 -1625
rect 79 -1628 80 -1627
rect 229 -1628 230 -1627
rect 268 -1628 269 -1627
rect 422 -1628 423 -1627
rect 565 -1628 566 -1627
rect 618 -1628 619 -1627
rect 688 -1628 689 -1627
rect 751 -1628 752 -1627
rect 779 -1628 780 -1627
rect 821 -1628 822 -1627
rect 107 -1630 108 -1629
rect 513 -1630 514 -1629
rect 569 -1630 570 -1629
rect 814 -1630 815 -1629
rect 93 -1632 94 -1631
rect 107 -1632 108 -1631
rect 121 -1632 122 -1631
rect 159 -1632 160 -1631
rect 163 -1632 164 -1631
rect 240 -1632 241 -1631
rect 268 -1632 269 -1631
rect 404 -1632 405 -1631
rect 513 -1632 514 -1631
rect 859 -1632 860 -1631
rect 93 -1634 94 -1633
rect 254 -1634 255 -1633
rect 282 -1634 283 -1633
rect 523 -1634 524 -1633
rect 569 -1634 570 -1633
rect 632 -1634 633 -1633
rect 688 -1634 689 -1633
rect 870 -1634 871 -1633
rect 128 -1636 129 -1635
rect 163 -1636 164 -1635
rect 198 -1636 199 -1635
rect 345 -1636 346 -1635
rect 376 -1636 377 -1635
rect 380 -1636 381 -1635
rect 387 -1636 388 -1635
rect 443 -1636 444 -1635
rect 576 -1636 577 -1635
rect 632 -1636 633 -1635
rect 695 -1636 696 -1635
rect 803 -1636 804 -1635
rect 814 -1636 815 -1635
rect 940 -1636 941 -1635
rect 114 -1638 115 -1637
rect 128 -1638 129 -1637
rect 149 -1638 150 -1637
rect 170 -1638 171 -1637
rect 208 -1638 209 -1637
rect 422 -1638 423 -1637
rect 443 -1638 444 -1637
rect 464 -1638 465 -1637
rect 478 -1638 479 -1637
rect 576 -1638 577 -1637
rect 590 -1638 591 -1637
rect 625 -1638 626 -1637
rect 702 -1638 703 -1637
rect 765 -1638 766 -1637
rect 86 -1640 87 -1639
rect 114 -1640 115 -1639
rect 152 -1640 153 -1639
rect 247 -1640 248 -1639
rect 275 -1640 276 -1639
rect 282 -1640 283 -1639
rect 296 -1640 297 -1639
rect 432 -1640 433 -1639
rect 478 -1640 479 -1639
rect 499 -1640 500 -1639
rect 590 -1640 591 -1639
rect 660 -1640 661 -1639
rect 709 -1640 710 -1639
rect 765 -1640 766 -1639
rect 86 -1642 87 -1641
rect 205 -1642 206 -1641
rect 212 -1642 213 -1641
rect 226 -1642 227 -1641
rect 247 -1642 248 -1641
rect 289 -1642 290 -1641
rect 296 -1642 297 -1641
rect 331 -1642 332 -1641
rect 359 -1642 360 -1641
rect 380 -1642 381 -1641
rect 390 -1642 391 -1641
rect 492 -1642 493 -1641
rect 499 -1642 500 -1641
rect 520 -1642 521 -1641
rect 604 -1642 605 -1641
rect 646 -1642 647 -1641
rect 709 -1642 710 -1641
rect 744 -1642 745 -1641
rect 758 -1642 759 -1641
rect 821 -1642 822 -1641
rect 44 -1644 45 -1643
rect 205 -1644 206 -1643
rect 212 -1644 213 -1643
rect 219 -1644 220 -1643
rect 226 -1644 227 -1643
rect 233 -1644 234 -1643
rect 289 -1644 290 -1643
rect 436 -1644 437 -1643
rect 485 -1644 486 -1643
rect 492 -1644 493 -1643
rect 583 -1644 584 -1643
rect 604 -1644 605 -1643
rect 611 -1644 612 -1643
rect 653 -1644 654 -1643
rect 716 -1644 717 -1643
rect 723 -1644 724 -1643
rect 730 -1644 731 -1643
rect 758 -1644 759 -1643
rect 23 -1646 24 -1645
rect 44 -1646 45 -1645
rect 135 -1646 136 -1645
rect 233 -1646 234 -1645
rect 317 -1646 318 -1645
rect 345 -1646 346 -1645
rect 373 -1646 374 -1645
rect 464 -1646 465 -1645
rect 485 -1646 486 -1645
rect 506 -1646 507 -1645
rect 541 -1646 542 -1645
rect 583 -1646 584 -1645
rect 614 -1646 615 -1645
rect 842 -1646 843 -1645
rect 135 -1648 136 -1647
rect 152 -1648 153 -1647
rect 156 -1648 157 -1647
rect 898 -1648 899 -1647
rect 100 -1650 101 -1649
rect 156 -1650 157 -1649
rect 170 -1650 171 -1649
rect 201 -1650 202 -1649
rect 306 -1650 307 -1649
rect 373 -1650 374 -1649
rect 394 -1650 395 -1649
rect 828 -1650 829 -1649
rect 842 -1650 843 -1649
rect 877 -1650 878 -1649
rect 51 -1652 52 -1651
rect 100 -1652 101 -1651
rect 177 -1652 178 -1651
rect 219 -1652 220 -1651
rect 317 -1652 318 -1651
rect 555 -1652 556 -1651
rect 716 -1652 717 -1651
rect 835 -1652 836 -1651
rect 40 -1654 41 -1653
rect 51 -1654 52 -1653
rect 184 -1654 185 -1653
rect 275 -1654 276 -1653
rect 324 -1654 325 -1653
rect 541 -1654 542 -1653
rect 555 -1654 556 -1653
rect 674 -1654 675 -1653
rect 733 -1654 734 -1653
rect 884 -1654 885 -1653
rect 184 -1656 185 -1655
rect 191 -1656 192 -1655
rect 331 -1656 332 -1655
rect 415 -1656 416 -1655
rect 436 -1656 437 -1655
rect 457 -1656 458 -1655
rect 506 -1656 507 -1655
rect 548 -1656 549 -1655
rect 744 -1656 745 -1655
rect 807 -1656 808 -1655
rect 884 -1656 885 -1655
rect 947 -1656 948 -1655
rect 191 -1658 192 -1657
rect 334 -1658 335 -1657
rect 338 -1658 339 -1657
rect 359 -1658 360 -1657
rect 394 -1658 395 -1657
rect 450 -1658 451 -1657
rect 786 -1658 787 -1657
rect 828 -1658 829 -1657
rect 303 -1660 304 -1659
rect 457 -1660 458 -1659
rect 772 -1660 773 -1659
rect 786 -1660 787 -1659
rect 800 -1660 801 -1659
rect 835 -1660 836 -1659
rect 313 -1662 314 -1661
rect 415 -1662 416 -1661
rect 429 -1662 430 -1661
rect 450 -1662 451 -1661
rect 800 -1662 801 -1661
rect 961 -1662 962 -1661
rect 807 -1664 808 -1663
rect 863 -1664 864 -1663
rect 863 -1666 864 -1665
rect 891 -1666 892 -1665
rect 891 -1668 892 -1667
rect 905 -1668 906 -1667
rect 905 -1670 906 -1669
rect 912 -1670 913 -1669
rect 44 -1681 45 -1680
rect 51 -1681 52 -1680
rect 65 -1681 66 -1680
rect 103 -1681 104 -1680
rect 107 -1681 108 -1680
rect 254 -1681 255 -1680
rect 264 -1681 265 -1680
rect 324 -1681 325 -1680
rect 383 -1681 384 -1680
rect 387 -1681 388 -1680
rect 408 -1681 409 -1680
rect 499 -1681 500 -1680
rect 513 -1681 514 -1680
rect 523 -1681 524 -1680
rect 541 -1681 542 -1680
rect 569 -1681 570 -1680
rect 593 -1681 594 -1680
rect 597 -1681 598 -1680
rect 611 -1681 612 -1680
rect 618 -1681 619 -1680
rect 625 -1681 626 -1680
rect 639 -1681 640 -1680
rect 646 -1681 647 -1680
rect 688 -1681 689 -1680
rect 723 -1681 724 -1680
rect 730 -1681 731 -1680
rect 758 -1681 759 -1680
rect 772 -1681 773 -1680
rect 779 -1681 780 -1680
rect 852 -1681 853 -1680
rect 856 -1681 857 -1680
rect 863 -1681 864 -1680
rect 898 -1681 899 -1680
rect 905 -1681 906 -1680
rect 47 -1683 48 -1682
rect 58 -1683 59 -1682
rect 86 -1683 87 -1682
rect 306 -1683 307 -1682
rect 310 -1683 311 -1682
rect 376 -1683 377 -1682
rect 380 -1683 381 -1682
rect 387 -1683 388 -1682
rect 422 -1683 423 -1682
rect 425 -1683 426 -1682
rect 429 -1683 430 -1682
rect 443 -1683 444 -1682
rect 450 -1683 451 -1682
rect 474 -1683 475 -1682
rect 520 -1683 521 -1682
rect 590 -1683 591 -1682
rect 604 -1683 605 -1682
rect 611 -1683 612 -1682
rect 632 -1683 633 -1682
rect 646 -1683 647 -1682
rect 653 -1683 654 -1682
rect 695 -1683 696 -1682
rect 709 -1683 710 -1682
rect 723 -1683 724 -1682
rect 737 -1683 738 -1682
rect 758 -1683 759 -1682
rect 782 -1683 783 -1682
rect 807 -1683 808 -1682
rect 817 -1683 818 -1682
rect 884 -1683 885 -1682
rect 93 -1685 94 -1684
rect 201 -1685 202 -1684
rect 212 -1685 213 -1684
rect 334 -1685 335 -1684
rect 373 -1685 374 -1684
rect 408 -1685 409 -1684
rect 422 -1685 423 -1684
rect 436 -1685 437 -1684
rect 450 -1685 451 -1684
rect 485 -1685 486 -1684
rect 569 -1685 570 -1684
rect 691 -1685 692 -1684
rect 709 -1685 710 -1684
rect 716 -1685 717 -1684
rect 737 -1685 738 -1684
rect 744 -1685 745 -1684
rect 786 -1685 787 -1684
rect 849 -1685 850 -1684
rect 884 -1685 885 -1684
rect 891 -1685 892 -1684
rect 75 -1687 76 -1686
rect 93 -1687 94 -1686
rect 100 -1687 101 -1686
rect 180 -1687 181 -1686
rect 201 -1687 202 -1686
rect 226 -1687 227 -1686
rect 240 -1687 241 -1686
rect 243 -1687 244 -1686
rect 282 -1687 283 -1686
rect 303 -1687 304 -1686
rect 310 -1687 311 -1686
rect 345 -1687 346 -1686
rect 373 -1687 374 -1686
rect 464 -1687 465 -1686
rect 576 -1687 577 -1686
rect 604 -1687 605 -1686
rect 667 -1687 668 -1686
rect 674 -1687 675 -1686
rect 677 -1687 678 -1686
rect 681 -1687 682 -1686
rect 744 -1687 745 -1686
rect 751 -1687 752 -1686
rect 793 -1687 794 -1686
rect 800 -1687 801 -1686
rect 807 -1687 808 -1686
rect 842 -1687 843 -1686
rect 849 -1687 850 -1686
rect 866 -1687 867 -1686
rect 114 -1689 115 -1688
rect 149 -1689 150 -1688
rect 156 -1689 157 -1688
rect 198 -1689 199 -1688
rect 219 -1689 220 -1688
rect 226 -1689 227 -1688
rect 240 -1689 241 -1688
rect 275 -1689 276 -1688
rect 324 -1689 325 -1688
rect 341 -1689 342 -1688
rect 345 -1689 346 -1688
rect 352 -1689 353 -1688
rect 401 -1689 402 -1688
rect 520 -1689 521 -1688
rect 527 -1689 528 -1688
rect 576 -1689 577 -1688
rect 702 -1689 703 -1688
rect 751 -1689 752 -1688
rect 765 -1689 766 -1688
rect 793 -1689 794 -1688
rect 821 -1689 822 -1688
rect 835 -1689 836 -1688
rect 117 -1691 118 -1690
rect 121 -1691 122 -1690
rect 128 -1691 129 -1690
rect 180 -1691 181 -1690
rect 184 -1691 185 -1690
rect 219 -1691 220 -1690
rect 247 -1691 248 -1690
rect 341 -1691 342 -1690
rect 404 -1691 405 -1690
rect 443 -1691 444 -1690
rect 464 -1691 465 -1690
rect 534 -1691 535 -1690
rect 765 -1691 766 -1690
rect 814 -1691 815 -1690
rect 821 -1691 822 -1690
rect 863 -1691 864 -1690
rect 128 -1693 129 -1692
rect 135 -1693 136 -1692
rect 156 -1693 157 -1692
rect 177 -1693 178 -1692
rect 268 -1693 269 -1692
rect 282 -1693 283 -1692
rect 415 -1693 416 -1692
rect 485 -1693 486 -1692
rect 527 -1693 528 -1692
rect 555 -1693 556 -1692
rect 163 -1695 164 -1694
rect 208 -1695 209 -1694
rect 261 -1695 262 -1694
rect 268 -1695 269 -1694
rect 275 -1695 276 -1694
rect 289 -1695 290 -1694
rect 394 -1695 395 -1694
rect 415 -1695 416 -1694
rect 436 -1695 437 -1694
rect 478 -1695 479 -1694
rect 163 -1697 164 -1696
rect 191 -1697 192 -1696
rect 289 -1697 290 -1696
rect 317 -1697 318 -1696
rect 394 -1697 395 -1696
rect 432 -1697 433 -1696
rect 457 -1697 458 -1696
rect 534 -1697 535 -1696
rect 177 -1699 178 -1698
rect 355 -1699 356 -1698
rect 457 -1699 458 -1698
rect 548 -1699 549 -1698
rect 191 -1701 192 -1700
rect 215 -1701 216 -1700
rect 317 -1701 318 -1700
rect 331 -1701 332 -1700
rect 471 -1701 472 -1700
rect 555 -1701 556 -1700
rect 296 -1703 297 -1702
rect 331 -1703 332 -1702
rect 478 -1703 479 -1702
rect 506 -1703 507 -1702
rect 548 -1703 549 -1702
rect 562 -1703 563 -1702
rect 492 -1705 493 -1704
rect 506 -1705 507 -1704
rect 562 -1705 563 -1704
rect 583 -1705 584 -1704
rect 425 -1707 426 -1706
rect 492 -1707 493 -1706
rect 583 -1707 584 -1706
rect 590 -1707 591 -1706
rect 58 -1718 59 -1717
rect 65 -1718 66 -1717
rect 93 -1718 94 -1717
rect 117 -1718 118 -1717
rect 121 -1718 122 -1717
rect 128 -1718 129 -1717
rect 142 -1718 143 -1717
rect 152 -1718 153 -1717
rect 156 -1718 157 -1717
rect 184 -1718 185 -1717
rect 212 -1718 213 -1717
rect 240 -1718 241 -1717
rect 268 -1718 269 -1717
rect 275 -1718 276 -1717
rect 289 -1718 290 -1717
rect 401 -1718 402 -1717
rect 411 -1718 412 -1717
rect 520 -1718 521 -1717
rect 562 -1718 563 -1717
rect 590 -1718 591 -1717
rect 593 -1718 594 -1717
rect 782 -1718 783 -1717
rect 793 -1718 794 -1717
rect 796 -1718 797 -1717
rect 828 -1718 829 -1717
rect 866 -1718 867 -1717
rect 103 -1720 104 -1719
rect 145 -1720 146 -1719
rect 149 -1720 150 -1719
rect 177 -1720 178 -1719
rect 205 -1720 206 -1719
rect 212 -1720 213 -1719
rect 215 -1720 216 -1719
rect 278 -1720 279 -1719
rect 299 -1720 300 -1719
rect 569 -1720 570 -1719
rect 583 -1720 584 -1719
rect 597 -1720 598 -1719
rect 604 -1720 605 -1719
rect 653 -1720 654 -1719
rect 674 -1720 675 -1719
rect 681 -1720 682 -1719
rect 702 -1720 703 -1719
rect 709 -1720 710 -1719
rect 730 -1720 731 -1719
rect 733 -1720 734 -1719
rect 772 -1720 773 -1719
rect 786 -1720 787 -1719
rect 793 -1720 794 -1719
rect 807 -1720 808 -1719
rect 821 -1720 822 -1719
rect 828 -1720 829 -1719
rect 835 -1720 836 -1719
rect 842 -1720 843 -1719
rect 845 -1720 846 -1719
rect 856 -1720 857 -1719
rect 107 -1722 108 -1721
rect 114 -1722 115 -1721
rect 142 -1722 143 -1721
rect 156 -1722 157 -1721
rect 163 -1722 164 -1721
rect 184 -1722 185 -1721
rect 219 -1722 220 -1721
rect 261 -1722 262 -1721
rect 324 -1722 325 -1721
rect 369 -1722 370 -1721
rect 380 -1722 381 -1721
rect 408 -1722 409 -1721
rect 422 -1722 423 -1721
rect 446 -1722 447 -1721
rect 464 -1722 465 -1721
rect 499 -1722 500 -1721
rect 597 -1722 598 -1721
rect 618 -1722 619 -1721
rect 639 -1722 640 -1721
rect 656 -1722 657 -1721
rect 709 -1722 710 -1721
rect 779 -1722 780 -1721
rect 849 -1722 850 -1721
rect 856 -1722 857 -1721
rect 163 -1724 164 -1723
rect 170 -1724 171 -1723
rect 226 -1724 227 -1723
rect 240 -1724 241 -1723
rect 296 -1724 297 -1723
rect 324 -1724 325 -1723
rect 338 -1724 339 -1723
rect 345 -1724 346 -1723
rect 352 -1724 353 -1723
rect 611 -1724 612 -1723
rect 730 -1724 731 -1723
rect 737 -1724 738 -1723
rect 233 -1726 234 -1725
rect 247 -1726 248 -1725
rect 282 -1726 283 -1725
rect 296 -1726 297 -1725
rect 338 -1726 339 -1725
rect 373 -1726 374 -1725
rect 422 -1726 423 -1725
rect 429 -1726 430 -1725
rect 464 -1726 465 -1725
rect 478 -1726 479 -1725
rect 492 -1726 493 -1725
rect 520 -1726 521 -1725
rect 737 -1726 738 -1725
rect 744 -1726 745 -1725
rect 226 -1728 227 -1727
rect 233 -1728 234 -1727
rect 331 -1728 332 -1727
rect 373 -1728 374 -1727
rect 429 -1728 430 -1727
rect 457 -1728 458 -1727
rect 471 -1728 472 -1727
rect 576 -1728 577 -1727
rect 744 -1728 745 -1727
rect 765 -1728 766 -1727
rect 317 -1730 318 -1729
rect 331 -1730 332 -1729
rect 345 -1730 346 -1729
rect 359 -1730 360 -1729
rect 366 -1730 367 -1729
rect 376 -1730 377 -1729
rect 457 -1730 458 -1729
rect 548 -1730 549 -1729
rect 555 -1730 556 -1729
rect 576 -1730 577 -1729
rect 758 -1730 759 -1729
rect 765 -1730 766 -1729
rect 254 -1732 255 -1731
rect 317 -1732 318 -1731
rect 352 -1732 353 -1731
rect 383 -1732 384 -1731
rect 478 -1732 479 -1731
rect 506 -1732 507 -1731
rect 534 -1732 535 -1731
rect 548 -1732 549 -1731
rect 555 -1732 556 -1731
rect 569 -1732 570 -1731
rect 751 -1732 752 -1731
rect 758 -1732 759 -1731
rect 359 -1734 360 -1733
rect 415 -1734 416 -1733
rect 485 -1734 486 -1733
rect 492 -1734 493 -1733
rect 499 -1734 500 -1733
rect 527 -1734 528 -1733
rect 366 -1736 367 -1735
rect 394 -1736 395 -1735
rect 415 -1736 416 -1735
rect 450 -1736 451 -1735
rect 513 -1736 514 -1735
rect 534 -1736 535 -1735
rect 387 -1738 388 -1737
rect 394 -1738 395 -1737
rect 436 -1738 437 -1737
rect 450 -1738 451 -1737
rect 485 -1738 486 -1737
rect 513 -1738 514 -1737
rect 436 -1740 437 -1739
rect 443 -1740 444 -1739
rect 796 -1740 797 -1739
rect 807 -1740 808 -1739
rect 44 -1751 45 -1750
rect 47 -1751 48 -1750
rect 58 -1751 59 -1750
rect 61 -1751 62 -1750
rect 65 -1751 66 -1750
rect 72 -1751 73 -1750
rect 93 -1751 94 -1750
rect 117 -1751 118 -1750
rect 121 -1751 122 -1750
rect 135 -1751 136 -1750
rect 159 -1751 160 -1750
rect 177 -1751 178 -1750
rect 184 -1751 185 -1750
rect 212 -1751 213 -1750
rect 219 -1751 220 -1750
rect 247 -1751 248 -1750
rect 282 -1751 283 -1750
rect 303 -1751 304 -1750
rect 352 -1751 353 -1750
rect 369 -1751 370 -1750
rect 373 -1751 374 -1750
rect 401 -1751 402 -1750
rect 443 -1751 444 -1750
rect 457 -1751 458 -1750
rect 464 -1751 465 -1750
rect 471 -1751 472 -1750
rect 488 -1751 489 -1750
rect 576 -1751 577 -1750
rect 586 -1751 587 -1750
rect 590 -1751 591 -1750
rect 646 -1751 647 -1750
rect 656 -1751 657 -1750
rect 716 -1751 717 -1750
rect 730 -1751 731 -1750
rect 765 -1751 766 -1750
rect 782 -1751 783 -1750
rect 807 -1751 808 -1750
rect 814 -1751 815 -1750
rect 842 -1751 843 -1750
rect 845 -1751 846 -1750
rect 968 -1751 969 -1750
rect 975 -1751 976 -1750
rect 65 -1753 66 -1752
rect 79 -1753 80 -1752
rect 107 -1753 108 -1752
rect 121 -1753 122 -1752
rect 128 -1753 129 -1752
rect 145 -1753 146 -1752
rect 163 -1753 164 -1752
rect 173 -1753 174 -1752
rect 219 -1753 220 -1752
rect 233 -1753 234 -1752
rect 289 -1753 290 -1752
rect 310 -1753 311 -1752
rect 317 -1753 318 -1752
rect 352 -1753 353 -1752
rect 366 -1753 367 -1752
rect 373 -1753 374 -1752
rect 387 -1753 388 -1752
rect 404 -1753 405 -1752
rect 450 -1753 451 -1752
rect 464 -1753 465 -1752
rect 471 -1753 472 -1752
rect 492 -1753 493 -1752
rect 499 -1753 500 -1752
rect 509 -1753 510 -1752
rect 527 -1753 528 -1752
rect 541 -1753 542 -1752
rect 548 -1753 549 -1752
rect 555 -1753 556 -1752
rect 562 -1753 563 -1752
rect 597 -1753 598 -1752
rect 709 -1753 710 -1752
rect 730 -1753 731 -1752
rect 772 -1753 773 -1752
rect 786 -1753 787 -1752
rect 128 -1755 129 -1754
rect 131 -1755 132 -1754
rect 135 -1755 136 -1754
rect 142 -1755 143 -1754
rect 233 -1755 234 -1754
rect 240 -1755 241 -1754
rect 296 -1755 297 -1754
rect 317 -1755 318 -1754
rect 429 -1755 430 -1754
rect 450 -1755 451 -1754
rect 457 -1755 458 -1754
rect 520 -1755 521 -1754
rect 530 -1755 531 -1754
rect 534 -1755 535 -1754
rect 562 -1755 563 -1754
rect 569 -1755 570 -1754
rect 702 -1755 703 -1754
rect 709 -1755 710 -1754
rect 758 -1755 759 -1754
rect 772 -1755 773 -1754
rect 779 -1755 780 -1754
rect 793 -1755 794 -1754
rect 138 -1757 139 -1756
rect 142 -1757 143 -1756
rect 229 -1757 230 -1756
rect 240 -1757 241 -1756
rect 296 -1757 297 -1756
rect 331 -1757 332 -1756
rect 429 -1757 430 -1756
rect 436 -1757 437 -1756
rect 751 -1757 752 -1756
rect 758 -1757 759 -1756
rect 793 -1757 794 -1756
rect 800 -1757 801 -1756
rect 310 -1759 311 -1758
rect 338 -1759 339 -1758
rect 737 -1759 738 -1758
rect 751 -1759 752 -1758
rect 324 -1761 325 -1760
rect 338 -1761 339 -1760
rect 737 -1761 738 -1760
rect 744 -1761 745 -1760
rect 324 -1763 325 -1762
rect 345 -1763 346 -1762
rect 345 -1765 346 -1764
rect 359 -1765 360 -1764
rect 359 -1767 360 -1766
rect 411 -1767 412 -1766
rect 58 -1778 59 -1777
rect 65 -1778 66 -1777
rect 75 -1778 76 -1777
rect 79 -1778 80 -1777
rect 93 -1778 94 -1777
rect 110 -1778 111 -1777
rect 117 -1778 118 -1777
rect 128 -1778 129 -1777
rect 135 -1778 136 -1777
rect 152 -1778 153 -1777
rect 170 -1778 171 -1777
rect 173 -1778 174 -1777
rect 191 -1778 192 -1777
rect 198 -1778 199 -1777
rect 219 -1778 220 -1777
rect 226 -1778 227 -1777
rect 247 -1778 248 -1777
rect 261 -1778 262 -1777
rect 282 -1778 283 -1777
rect 320 -1778 321 -1777
rect 331 -1778 332 -1777
rect 345 -1778 346 -1777
rect 380 -1778 381 -1777
rect 387 -1778 388 -1777
rect 394 -1778 395 -1777
rect 411 -1778 412 -1777
rect 502 -1778 503 -1777
rect 506 -1778 507 -1777
rect 520 -1778 521 -1777
rect 527 -1778 528 -1777
rect 562 -1778 563 -1777
rect 565 -1778 566 -1777
rect 709 -1778 710 -1777
rect 716 -1778 717 -1777
rect 723 -1778 724 -1777
rect 747 -1778 748 -1777
rect 751 -1778 752 -1777
rect 765 -1778 766 -1777
rect 772 -1778 773 -1777
rect 779 -1778 780 -1777
rect 828 -1778 829 -1777
rect 838 -1778 839 -1777
rect 880 -1778 881 -1777
rect 884 -1778 885 -1777
rect 72 -1780 73 -1779
rect 79 -1780 80 -1779
rect 152 -1780 153 -1779
rect 156 -1780 157 -1779
rect 226 -1780 227 -1779
rect 233 -1780 234 -1779
rect 275 -1780 276 -1779
rect 282 -1780 283 -1779
rect 289 -1780 290 -1779
rect 306 -1780 307 -1779
rect 324 -1780 325 -1779
rect 331 -1780 332 -1779
rect 373 -1780 374 -1779
rect 380 -1780 381 -1779
rect 401 -1780 402 -1779
rect 422 -1780 423 -1779
rect 730 -1780 731 -1779
rect 772 -1780 773 -1779
rect 296 -1782 297 -1781
rect 313 -1782 314 -1781
rect 411 -1782 412 -1781
rect 457 -1782 458 -1781
rect 296 -1784 297 -1783
rect 303 -1784 304 -1783
rect 306 -1784 307 -1783
rect 362 -1784 363 -1783
rect 450 -1784 451 -1783
rect 457 -1784 458 -1783
rect 310 -1786 311 -1785
rect 324 -1786 325 -1785
rect 450 -1786 451 -1785
rect 471 -1786 472 -1785
rect 464 -1788 465 -1787
rect 471 -1788 472 -1787
rect 68 -1799 69 -1798
rect 79 -1799 80 -1798
rect 142 -1799 143 -1798
rect 149 -1799 150 -1798
rect 156 -1799 157 -1798
rect 159 -1799 160 -1798
rect 184 -1799 185 -1798
rect 191 -1799 192 -1798
rect 205 -1799 206 -1798
rect 208 -1799 209 -1798
rect 240 -1799 241 -1798
rect 247 -1799 248 -1798
rect 261 -1799 262 -1798
rect 268 -1799 269 -1798
rect 324 -1799 325 -1798
rect 341 -1799 342 -1798
rect 380 -1799 381 -1798
rect 383 -1799 384 -1798
rect 422 -1799 423 -1798
rect 429 -1799 430 -1798
rect 432 -1799 433 -1798
rect 443 -1799 444 -1798
rect 457 -1799 458 -1798
rect 464 -1799 465 -1798
rect 471 -1799 472 -1798
rect 481 -1799 482 -1798
rect 506 -1799 507 -1798
rect 513 -1799 514 -1798
rect 516 -1799 517 -1798
rect 520 -1799 521 -1798
rect 737 -1799 738 -1798
rect 751 -1799 752 -1798
rect 754 -1799 755 -1798
rect 765 -1799 766 -1798
rect 793 -1799 794 -1798
rect 796 -1799 797 -1798
rect 898 -1799 899 -1798
rect 905 -1799 906 -1798
rect 1024 -1799 1025 -1798
rect 1027 -1799 1028 -1798
rect 331 -1801 332 -1800
rect 345 -1801 346 -1800
rect 415 -1801 416 -1800
rect 422 -1801 423 -1800
rect 439 -1801 440 -1800
rect 450 -1801 451 -1800
rect 471 -1801 472 -1800
rect 478 -1801 479 -1800
rect 744 -1801 745 -1800
rect 758 -1801 759 -1800
rect 331 -1803 332 -1802
rect 338 -1803 339 -1802
rect 187 -1814 188 -1813
rect 191 -1814 192 -1813
rect 222 -1814 223 -1813
rect 226 -1814 227 -1813
rect 264 -1814 265 -1813
rect 268 -1814 269 -1813
rect 296 -1814 297 -1813
rect 306 -1814 307 -1813
rect 324 -1814 325 -1813
rect 331 -1814 332 -1813
rect 352 -1814 353 -1813
rect 359 -1814 360 -1813
rect 376 -1814 377 -1813
rect 387 -1814 388 -1813
rect 422 -1814 423 -1813
rect 429 -1814 430 -1813
rect 747 -1814 748 -1813
rect 751 -1814 752 -1813
rect 901 -1814 902 -1813
rect 905 -1814 906 -1813
<< metal2 >>
rect 177 -3 178 1
rect 198 -3 199 1
rect 212 -3 213 1
rect 219 -3 220 1
rect 236 -3 237 1
rect 240 -3 241 1
rect 254 -3 255 1
rect 261 -3 262 1
rect 285 -3 286 1
rect 289 -3 290 1
rect 303 -3 304 1
rect 310 -3 311 1
rect 338 -3 339 1
rect 348 -3 349 1
rect 352 -3 353 1
rect 359 -3 360 1
rect 366 -3 367 1
rect 408 -3 409 1
rect 467 -3 468 1
rect 471 -3 472 1
rect 478 -3 479 1
rect 485 -3 486 1
rect 534 -3 535 1
rect 541 -3 542 1
rect 576 -3 577 1
rect 583 -3 584 1
rect 604 -3 605 1
rect 611 -3 612 1
rect 730 -3 731 1
rect 740 -3 741 1
rect 184 -3 185 -1
rect 194 -3 195 -1
rect 114 -20 115 -12
rect 121 -20 122 -12
rect 156 -20 157 -12
rect 163 -20 164 -12
rect 170 -20 171 -12
rect 177 -13 178 -11
rect 184 -13 185 -11
rect 184 -20 185 -12
rect 184 -13 185 -11
rect 184 -20 185 -12
rect 219 -13 220 -11
rect 226 -20 227 -12
rect 240 -13 241 -11
rect 254 -20 255 -12
rect 278 -13 279 -11
rect 282 -20 283 -12
rect 296 -13 297 -11
rect 296 -20 297 -12
rect 296 -13 297 -11
rect 296 -20 297 -12
rect 303 -13 304 -11
rect 310 -20 311 -12
rect 317 -13 318 -11
rect 317 -20 318 -12
rect 317 -13 318 -11
rect 317 -20 318 -12
rect 345 -20 346 -12
rect 366 -13 367 -11
rect 408 -13 409 -11
rect 443 -20 444 -12
rect 450 -20 451 -12
rect 460 -13 461 -11
rect 474 -20 475 -12
rect 478 -20 479 -12
rect 485 -13 486 -11
rect 492 -20 493 -12
rect 527 -20 528 -12
rect 558 -13 559 -11
rect 583 -13 584 -11
rect 583 -20 584 -12
rect 583 -13 584 -11
rect 583 -20 584 -12
rect 604 -13 605 -11
rect 611 -20 612 -12
rect 618 -20 619 -12
rect 621 -13 622 -11
rect 688 -20 689 -12
rect 698 -20 699 -12
rect 730 -13 731 -11
rect 730 -20 731 -12
rect 730 -13 731 -11
rect 730 -20 731 -12
rect 215 -20 216 -14
rect 219 -20 220 -14
rect 247 -20 248 -14
rect 261 -15 262 -11
rect 289 -15 290 -11
rect 303 -20 304 -14
rect 352 -15 353 -11
rect 359 -20 360 -14
rect 366 -20 367 -14
rect 373 -20 374 -14
rect 415 -20 416 -14
rect 422 -15 423 -11
rect 425 -20 426 -14
rect 429 -20 430 -14
rect 457 -20 458 -14
rect 467 -20 468 -14
rect 471 -15 472 -11
rect 485 -20 486 -14
rect 541 -15 542 -11
rect 541 -20 542 -14
rect 541 -15 542 -11
rect 541 -20 542 -14
rect 555 -15 556 -11
rect 604 -20 605 -14
rect 240 -20 241 -16
rect 261 -20 262 -16
rect 278 -20 279 -16
rect 289 -20 290 -16
rect 338 -17 339 -11
rect 352 -20 353 -16
rect 334 -20 335 -18
rect 338 -20 339 -18
rect 58 -43 59 -29
rect 61 -30 62 -28
rect 79 -30 80 -28
rect 79 -43 80 -29
rect 79 -30 80 -28
rect 79 -43 80 -29
rect 114 -43 115 -29
rect 124 -43 125 -29
rect 128 -30 129 -28
rect 128 -43 129 -29
rect 128 -30 129 -28
rect 128 -43 129 -29
rect 142 -43 143 -29
rect 170 -30 171 -28
rect 184 -30 185 -28
rect 198 -43 199 -29
rect 212 -43 213 -29
rect 219 -30 220 -28
rect 226 -30 227 -28
rect 261 -43 262 -29
rect 268 -43 269 -29
rect 296 -30 297 -28
rect 317 -30 318 -28
rect 324 -43 325 -29
rect 334 -43 335 -29
rect 345 -30 346 -28
rect 352 -30 353 -28
rect 373 -43 374 -29
rect 380 -30 381 -28
rect 380 -43 381 -29
rect 380 -30 381 -28
rect 380 -43 381 -29
rect 387 -43 388 -29
rect 401 -43 402 -29
rect 408 -43 409 -29
rect 411 -30 412 -28
rect 415 -30 416 -28
rect 425 -43 426 -29
rect 429 -30 430 -28
rect 432 -34 433 -29
rect 443 -30 444 -28
rect 471 -43 472 -29
rect 478 -30 479 -28
rect 478 -43 479 -29
rect 478 -30 479 -28
rect 478 -43 479 -29
rect 485 -30 486 -28
rect 485 -43 486 -29
rect 485 -30 486 -28
rect 485 -43 486 -29
rect 492 -30 493 -28
rect 499 -43 500 -29
rect 513 -43 514 -29
rect 537 -43 538 -29
rect 541 -30 542 -28
rect 548 -43 549 -29
rect 576 -43 577 -29
rect 579 -30 580 -28
rect 583 -30 584 -28
rect 597 -43 598 -29
rect 604 -30 605 -28
rect 632 -43 633 -29
rect 646 -43 647 -29
rect 660 -43 661 -29
rect 688 -30 689 -28
rect 688 -43 689 -29
rect 688 -30 689 -28
rect 688 -43 689 -29
rect 709 -30 710 -28
rect 786 -43 787 -29
rect 807 -43 808 -29
rect 814 -43 815 -29
rect 121 -32 122 -28
rect 135 -43 136 -31
rect 152 -43 153 -31
rect 156 -43 157 -31
rect 163 -32 164 -28
rect 173 -43 174 -31
rect 177 -43 178 -31
rect 226 -43 227 -31
rect 233 -43 234 -31
rect 240 -32 241 -28
rect 254 -32 255 -28
rect 296 -43 297 -31
rect 345 -43 346 -31
rect 366 -32 367 -28
rect 429 -43 430 -31
rect 436 -32 437 -28
rect 450 -32 451 -28
rect 450 -43 451 -31
rect 450 -32 451 -28
rect 450 -43 451 -31
rect 457 -32 458 -28
rect 457 -43 458 -31
rect 457 -32 458 -28
rect 457 -43 458 -31
rect 527 -32 528 -28
rect 555 -43 556 -31
rect 572 -43 573 -31
rect 583 -43 584 -31
rect 604 -43 605 -31
rect 611 -32 612 -28
rect 625 -43 626 -31
rect 712 -32 713 -28
rect 730 -32 731 -28
rect 730 -43 731 -31
rect 730 -32 731 -28
rect 730 -43 731 -31
rect 163 -43 164 -33
rect 170 -43 171 -33
rect 180 -34 181 -28
rect 184 -43 185 -33
rect 240 -43 241 -33
rect 282 -34 283 -28
rect 289 -34 290 -28
rect 289 -43 290 -33
rect 289 -34 290 -28
rect 289 -43 290 -33
rect 352 -43 353 -33
rect 397 -43 398 -33
rect 436 -43 437 -33
rect 541 -43 542 -33
rect 562 -43 563 -33
rect 611 -43 612 -33
rect 618 -34 619 -28
rect 247 -36 248 -28
rect 254 -43 255 -35
rect 257 -43 258 -35
rect 275 -43 276 -35
rect 282 -43 283 -35
rect 310 -36 311 -28
rect 359 -36 360 -28
rect 366 -43 367 -35
rect 247 -43 248 -37
rect 271 -38 272 -28
rect 303 -38 304 -28
rect 310 -43 311 -37
rect 338 -38 339 -28
rect 359 -43 360 -37
rect 303 -43 304 -39
rect 331 -43 332 -39
rect 317 -43 318 -41
rect 338 -43 339 -41
rect 58 -53 59 -51
rect 58 -82 59 -52
rect 58 -53 59 -51
rect 58 -82 59 -52
rect 65 -53 66 -51
rect 65 -82 66 -52
rect 65 -53 66 -51
rect 65 -82 66 -52
rect 79 -53 80 -51
rect 79 -82 80 -52
rect 79 -53 80 -51
rect 79 -82 80 -52
rect 93 -82 94 -52
rect 103 -82 104 -52
rect 107 -53 108 -51
rect 149 -82 150 -52
rect 163 -53 164 -51
rect 163 -82 164 -52
rect 163 -53 164 -51
rect 163 -82 164 -52
rect 170 -53 171 -51
rect 184 -53 185 -51
rect 226 -53 227 -51
rect 278 -82 279 -52
rect 310 -53 311 -51
rect 331 -82 332 -52
rect 338 -82 339 -52
rect 401 -53 402 -51
rect 415 -82 416 -52
rect 460 -82 461 -52
rect 478 -53 479 -51
rect 506 -82 507 -52
rect 513 -53 514 -51
rect 520 -82 521 -52
rect 534 -53 535 -51
rect 618 -82 619 -52
rect 660 -53 661 -51
rect 674 -82 675 -52
rect 688 -53 689 -51
rect 702 -82 703 -52
rect 730 -53 731 -51
rect 730 -82 731 -52
rect 730 -53 731 -51
rect 730 -82 731 -52
rect 793 -82 794 -52
rect 807 -53 808 -51
rect 898 -53 899 -51
rect 898 -82 899 -52
rect 898 -53 899 -51
rect 898 -82 899 -52
rect 1087 -82 1088 -52
rect 1097 -82 1098 -52
rect 110 -82 111 -54
rect 205 -82 206 -54
rect 229 -55 230 -51
rect 296 -55 297 -51
rect 345 -55 346 -51
rect 345 -82 346 -54
rect 345 -55 346 -51
rect 345 -82 346 -54
rect 366 -55 367 -51
rect 366 -82 367 -54
rect 366 -55 367 -51
rect 366 -82 367 -54
rect 373 -55 374 -51
rect 387 -82 388 -54
rect 429 -55 430 -51
rect 443 -55 444 -51
rect 485 -55 486 -51
rect 513 -82 514 -54
rect 541 -82 542 -54
rect 583 -55 584 -51
rect 611 -55 612 -51
rect 611 -82 612 -54
rect 611 -55 612 -51
rect 611 -82 612 -54
rect 653 -55 654 -51
rect 660 -82 661 -54
rect 786 -55 787 -51
rect 807 -82 808 -54
rect 114 -57 115 -51
rect 114 -82 115 -56
rect 114 -57 115 -51
rect 114 -82 115 -56
rect 121 -57 122 -51
rect 135 -57 136 -51
rect 142 -57 143 -51
rect 142 -82 143 -56
rect 142 -57 143 -51
rect 142 -82 143 -56
rect 170 -82 171 -56
rect 191 -57 192 -51
rect 233 -57 234 -51
rect 254 -82 255 -56
rect 289 -57 290 -51
rect 310 -82 311 -56
rect 373 -82 374 -56
rect 467 -82 468 -56
rect 474 -82 475 -56
rect 485 -82 486 -56
rect 499 -57 500 -51
rect 534 -82 535 -56
rect 555 -57 556 -51
rect 646 -82 647 -56
rect 128 -82 129 -58
rect 177 -59 178 -51
rect 184 -82 185 -58
rect 275 -59 276 -51
rect 289 -82 290 -58
rect 299 -82 300 -58
rect 380 -59 381 -51
rect 401 -82 402 -58
rect 422 -59 423 -51
rect 443 -82 444 -58
rect 471 -59 472 -51
rect 499 -82 500 -58
rect 527 -82 528 -58
rect 555 -82 556 -58
rect 569 -82 570 -58
rect 625 -59 626 -51
rect 632 -59 633 -51
rect 653 -82 654 -58
rect 135 -82 136 -60
rect 156 -61 157 -51
rect 191 -82 192 -60
rect 208 -61 209 -51
rect 233 -82 234 -60
rect 261 -61 262 -51
rect 380 -82 381 -60
rect 408 -61 409 -51
rect 422 -82 423 -60
rect 450 -61 451 -51
rect 495 -82 496 -60
rect 625 -82 626 -60
rect 632 -82 633 -60
rect 639 -82 640 -60
rect 156 -82 157 -62
rect 198 -63 199 -51
rect 208 -82 209 -62
rect 212 -63 213 -51
rect 240 -63 241 -51
rect 240 -82 241 -62
rect 240 -63 241 -51
rect 240 -82 241 -62
rect 247 -63 248 -51
rect 261 -82 262 -62
rect 408 -82 409 -62
rect 457 -63 458 -51
rect 576 -63 577 -51
rect 583 -82 584 -62
rect 198 -82 199 -64
rect 282 -65 283 -51
rect 429 -82 430 -64
rect 446 -65 447 -51
rect 576 -82 577 -64
rect 604 -65 605 -51
rect 212 -82 213 -66
rect 303 -67 304 -51
rect 436 -67 437 -51
rect 450 -82 451 -66
rect 597 -67 598 -51
rect 604 -82 605 -66
rect 222 -69 223 -51
rect 247 -82 248 -68
rect 268 -69 269 -51
rect 303 -82 304 -68
rect 439 -82 440 -68
rect 478 -82 479 -68
rect 590 -69 591 -51
rect 597 -82 598 -68
rect 268 -82 269 -70
rect 359 -71 360 -51
rect 562 -71 563 -51
rect 590 -82 591 -70
rect 282 -82 283 -72
rect 317 -73 318 -51
rect 548 -73 549 -51
rect 562 -82 563 -72
rect 317 -82 318 -74
rect 352 -75 353 -51
rect 446 -82 447 -74
rect 548 -82 549 -74
rect 324 -77 325 -51
rect 352 -82 353 -76
rect 324 -82 325 -78
rect 394 -79 395 -51
rect 131 -81 132 -51
rect 394 -82 395 -80
rect 30 -119 31 -91
rect 44 -119 45 -91
rect 51 -119 52 -91
rect 65 -92 66 -90
rect 89 -92 90 -90
rect 93 -92 94 -90
rect 100 -119 101 -91
rect 156 -92 157 -90
rect 219 -119 220 -91
rect 268 -92 269 -90
rect 275 -119 276 -91
rect 289 -92 290 -90
rect 299 -92 300 -90
rect 352 -92 353 -90
rect 366 -92 367 -90
rect 394 -119 395 -91
rect 397 -92 398 -90
rect 411 -119 412 -91
rect 429 -92 430 -90
rect 495 -92 496 -90
rect 527 -119 528 -91
rect 555 -92 556 -90
rect 583 -92 584 -90
rect 583 -119 584 -91
rect 583 -92 584 -90
rect 583 -119 584 -91
rect 597 -92 598 -90
rect 632 -119 633 -91
rect 646 -92 647 -90
rect 688 -119 689 -91
rect 730 -92 731 -90
rect 737 -119 738 -91
rect 758 -119 759 -91
rect 779 -119 780 -91
rect 800 -119 801 -91
rect 807 -92 808 -90
rect 898 -92 899 -90
rect 905 -119 906 -91
rect 975 -119 976 -91
rect 978 -92 979 -90
rect 1087 -92 1088 -90
rect 1087 -119 1088 -91
rect 1087 -92 1088 -90
rect 1087 -119 1088 -91
rect 54 -94 55 -90
rect 65 -119 66 -93
rect 93 -119 94 -93
rect 142 -94 143 -90
rect 149 -94 150 -90
rect 187 -94 188 -90
rect 261 -94 262 -90
rect 268 -119 269 -93
rect 282 -94 283 -90
rect 289 -119 290 -93
rect 303 -94 304 -90
rect 306 -112 307 -93
rect 331 -94 332 -90
rect 331 -119 332 -93
rect 331 -94 332 -90
rect 331 -119 332 -93
rect 338 -94 339 -90
rect 366 -119 367 -93
rect 387 -94 388 -90
rect 390 -94 391 -90
rect 401 -94 402 -90
rect 429 -119 430 -93
rect 450 -94 451 -90
rect 471 -119 472 -93
rect 478 -94 479 -90
rect 492 -119 493 -93
rect 541 -94 542 -90
rect 597 -119 598 -93
rect 604 -94 605 -90
rect 667 -119 668 -93
rect 674 -94 675 -90
rect 716 -119 717 -93
rect 765 -119 766 -93
rect 793 -94 794 -90
rect 58 -96 59 -90
rect 58 -119 59 -95
rect 58 -96 59 -90
rect 58 -119 59 -95
rect 107 -119 108 -95
rect 415 -96 416 -90
rect 450 -119 451 -95
rect 639 -96 640 -90
rect 681 -96 682 -90
rect 723 -119 724 -95
rect 114 -98 115 -90
rect 114 -119 115 -97
rect 114 -98 115 -90
rect 114 -119 115 -97
rect 121 -119 122 -97
rect 184 -98 185 -90
rect 240 -98 241 -90
rect 261 -119 262 -97
rect 282 -119 283 -97
rect 317 -98 318 -90
rect 327 -119 328 -97
rect 338 -119 339 -97
rect 373 -98 374 -90
rect 415 -119 416 -97
rect 457 -119 458 -97
rect 485 -98 486 -90
rect 534 -98 535 -90
rect 639 -119 640 -97
rect 702 -98 703 -90
rect 730 -119 731 -97
rect 124 -100 125 -90
rect 177 -119 178 -99
rect 240 -119 241 -99
rect 247 -100 248 -90
rect 303 -119 304 -99
rect 317 -119 318 -99
rect 324 -100 325 -90
rect 380 -100 381 -90
rect 401 -119 402 -99
rect 408 -100 409 -90
rect 443 -119 444 -99
rect 467 -119 468 -99
rect 485 -119 486 -99
rect 499 -100 500 -90
rect 534 -119 535 -99
rect 541 -119 542 -99
rect 569 -100 570 -90
rect 590 -100 591 -90
rect 646 -119 647 -99
rect 660 -100 661 -90
rect 702 -119 703 -99
rect 128 -102 129 -90
rect 180 -102 181 -90
rect 324 -119 325 -101
rect 436 -102 437 -90
rect 520 -102 521 -90
rect 569 -119 570 -101
rect 593 -119 594 -101
rect 681 -119 682 -101
rect 128 -119 129 -103
rect 345 -104 346 -90
rect 355 -119 356 -103
rect 520 -119 521 -103
rect 562 -104 563 -90
rect 604 -119 605 -103
rect 611 -104 612 -90
rect 660 -119 661 -103
rect 135 -106 136 -90
rect 180 -119 181 -105
rect 212 -106 213 -90
rect 345 -119 346 -105
rect 362 -106 363 -90
rect 499 -119 500 -105
rect 506 -106 507 -90
rect 562 -119 563 -105
rect 618 -106 619 -90
rect 674 -119 675 -105
rect 142 -119 143 -107
rect 198 -108 199 -90
rect 212 -119 213 -107
rect 233 -108 234 -90
rect 373 -119 374 -107
rect 436 -119 437 -107
rect 548 -108 549 -90
rect 611 -119 612 -107
rect 625 -108 626 -90
rect 695 -119 696 -107
rect 149 -119 150 -109
rect 205 -110 206 -90
rect 233 -119 234 -109
rect 254 -110 255 -90
rect 387 -119 388 -109
rect 422 -110 423 -90
rect 513 -110 514 -90
rect 625 -119 626 -109
rect 156 -119 157 -111
rect 163 -112 164 -90
rect 198 -119 199 -111
rect 229 -112 230 -90
rect 390 -119 391 -111
rect 422 -119 423 -111
rect 576 -112 577 -90
rect 618 -119 619 -111
rect 163 -119 164 -113
rect 170 -114 171 -90
rect 205 -119 206 -113
rect 359 -114 360 -90
rect 408 -119 409 -113
rect 513 -119 514 -113
rect 576 -119 577 -113
rect 653 -114 654 -90
rect 170 -119 171 -115
rect 191 -116 192 -90
rect 229 -119 230 -115
rect 254 -119 255 -115
rect 299 -119 300 -115
rect 359 -119 360 -115
rect 191 -119 192 -117
rect 222 -118 223 -90
rect 23 -180 24 -128
rect 44 -180 45 -128
rect 47 -129 48 -127
rect 65 -129 66 -127
rect 79 -180 80 -128
rect 86 -180 87 -128
rect 121 -129 122 -127
rect 184 -180 185 -128
rect 219 -129 220 -127
rect 324 -129 325 -127
rect 338 -129 339 -127
rect 408 -180 409 -128
rect 457 -129 458 -127
rect 464 -129 465 -127
rect 495 -180 496 -128
rect 506 -180 507 -128
rect 541 -129 542 -127
rect 593 -129 594 -127
rect 656 -129 657 -127
rect 758 -180 759 -128
rect 779 -129 780 -127
rect 849 -180 850 -128
rect 905 -129 906 -127
rect 919 -180 920 -128
rect 975 -129 976 -127
rect 975 -180 976 -128
rect 975 -129 976 -127
rect 975 -180 976 -128
rect 1087 -129 1088 -127
rect 1087 -180 1088 -128
rect 1087 -129 1088 -127
rect 1087 -180 1088 -128
rect 30 -131 31 -127
rect 37 -180 38 -130
rect 121 -180 122 -130
rect 205 -131 206 -127
rect 219 -180 220 -130
rect 282 -131 283 -127
rect 296 -180 297 -130
rect 303 -131 304 -127
rect 324 -180 325 -130
rect 338 -180 339 -130
rect 345 -131 346 -127
rect 352 -131 353 -127
rect 380 -131 381 -127
rect 429 -131 430 -127
rect 443 -131 444 -127
rect 457 -180 458 -130
rect 509 -131 510 -127
rect 541 -180 542 -130
rect 555 -131 556 -127
rect 695 -131 696 -127
rect 737 -131 738 -127
rect 751 -180 752 -130
rect 30 -180 31 -132
rect 51 -133 52 -127
rect 149 -133 150 -127
rect 376 -133 377 -127
rect 394 -133 395 -127
rect 429 -180 430 -132
rect 471 -133 472 -127
rect 555 -180 556 -132
rect 583 -133 584 -127
rect 653 -180 654 -132
rect 667 -133 668 -127
rect 786 -180 787 -132
rect 51 -180 52 -134
rect 58 -135 59 -127
rect 149 -180 150 -134
rect 481 -135 482 -127
rect 513 -135 514 -127
rect 583 -180 584 -134
rect 590 -180 591 -134
rect 688 -135 689 -127
rect 695 -180 696 -134
rect 765 -135 766 -127
rect 156 -137 157 -127
rect 166 -180 167 -136
rect 170 -137 171 -127
rect 380 -180 381 -136
rect 394 -180 395 -136
rect 415 -137 416 -127
rect 450 -137 451 -127
rect 471 -180 472 -136
rect 520 -137 521 -127
rect 779 -180 780 -136
rect 58 -180 59 -138
rect 156 -180 157 -138
rect 170 -180 171 -138
rect 187 -139 188 -127
rect 198 -139 199 -127
rect 376 -180 377 -138
rect 401 -139 402 -127
rect 415 -180 416 -138
rect 450 -180 451 -138
rect 548 -139 549 -127
rect 604 -139 605 -127
rect 667 -180 668 -138
rect 674 -139 675 -127
rect 793 -180 794 -138
rect 142 -141 143 -127
rect 401 -180 402 -140
rect 499 -141 500 -127
rect 548 -180 549 -140
rect 562 -141 563 -127
rect 674 -180 675 -140
rect 681 -141 682 -127
rect 807 -180 808 -140
rect 135 -143 136 -127
rect 499 -180 500 -142
rect 527 -143 528 -127
rect 562 -180 563 -142
rect 604 -180 605 -142
rect 723 -143 724 -127
rect 744 -180 745 -142
rect 800 -143 801 -127
rect 142 -180 143 -144
rect 163 -145 164 -127
rect 205 -180 206 -144
rect 212 -145 213 -127
rect 226 -180 227 -144
rect 348 -180 349 -144
rect 492 -145 493 -127
rect 527 -180 528 -144
rect 569 -145 570 -127
rect 723 -180 724 -144
rect 730 -145 731 -127
rect 800 -180 801 -144
rect 212 -180 213 -146
rect 275 -147 276 -127
rect 282 -180 283 -146
rect 390 -180 391 -146
rect 569 -180 570 -146
rect 702 -147 703 -127
rect 709 -147 710 -127
rect 737 -180 738 -146
rect 229 -149 230 -127
rect 359 -149 360 -127
rect 618 -149 619 -127
rect 681 -180 682 -148
rect 702 -180 703 -148
rect 845 -180 846 -148
rect 233 -151 234 -127
rect 352 -180 353 -150
rect 359 -180 360 -150
rect 366 -151 367 -127
rect 534 -151 535 -127
rect 618 -180 619 -150
rect 625 -151 626 -127
rect 730 -180 731 -150
rect 233 -180 234 -152
rect 247 -153 248 -127
rect 250 -153 251 -127
rect 254 -153 255 -127
rect 275 -180 276 -152
rect 467 -180 468 -152
rect 597 -153 598 -127
rect 625 -180 626 -152
rect 632 -153 633 -127
rect 688 -180 689 -152
rect 240 -180 241 -154
rect 317 -155 318 -127
rect 334 -180 335 -154
rect 513 -180 514 -154
rect 597 -180 598 -154
rect 716 -155 717 -127
rect 72 -180 73 -156
rect 317 -180 318 -156
rect 345 -180 346 -156
rect 422 -157 423 -127
rect 478 -157 479 -127
rect 632 -180 633 -156
rect 639 -157 640 -127
rect 765 -180 766 -156
rect 243 -159 244 -127
rect 320 -180 321 -158
rect 366 -180 367 -158
rect 383 -159 384 -127
rect 422 -180 423 -158
rect 772 -180 773 -158
rect 247 -180 248 -160
rect 261 -161 262 -127
rect 303 -180 304 -160
rect 331 -161 332 -127
rect 436 -161 437 -127
rect 639 -180 640 -160
rect 646 -161 647 -127
rect 709 -180 710 -160
rect 254 -180 255 -162
rect 289 -163 290 -127
rect 331 -180 332 -162
rect 443 -180 444 -162
rect 478 -180 479 -162
rect 814 -180 815 -162
rect 107 -165 108 -127
rect 289 -180 290 -164
rect 387 -165 388 -127
rect 436 -180 437 -164
rect 611 -165 612 -127
rect 646 -180 647 -164
rect 660 -165 661 -127
rect 716 -180 717 -164
rect 107 -180 108 -166
rect 128 -167 129 -127
rect 261 -180 262 -166
rect 268 -167 269 -127
rect 387 -180 388 -166
rect 485 -167 486 -127
rect 537 -180 538 -166
rect 660 -180 661 -166
rect 128 -180 129 -168
rect 138 -169 139 -127
rect 268 -180 269 -168
rect 310 -169 311 -127
rect 576 -169 577 -127
rect 611 -180 612 -168
rect 100 -171 101 -127
rect 310 -180 311 -170
rect 523 -180 524 -170
rect 576 -180 577 -170
rect 93 -173 94 -127
rect 100 -180 101 -172
rect 114 -180 115 -172
rect 138 -180 139 -172
rect 93 -180 94 -174
rect 177 -175 178 -127
rect 177 -180 178 -176
rect 191 -177 192 -127
rect 191 -180 192 -178
rect 488 -180 489 -178
rect 16 -239 17 -189
rect 303 -190 304 -188
rect 317 -190 318 -188
rect 576 -190 577 -188
rect 758 -190 759 -188
rect 870 -239 871 -189
rect 919 -190 920 -188
rect 947 -239 948 -189
rect 975 -190 976 -188
rect 975 -239 976 -189
rect 975 -190 976 -188
rect 975 -239 976 -189
rect 1087 -190 1088 -188
rect 1087 -239 1088 -189
rect 1087 -190 1088 -188
rect 1087 -239 1088 -189
rect 30 -192 31 -188
rect 65 -192 66 -188
rect 68 -192 69 -188
rect 103 -239 104 -191
rect 117 -239 118 -191
rect 198 -192 199 -188
rect 201 -192 202 -188
rect 233 -192 234 -188
rect 240 -192 241 -188
rect 331 -239 332 -191
rect 338 -239 339 -191
rect 436 -192 437 -188
rect 460 -239 461 -191
rect 730 -192 731 -188
rect 765 -192 766 -188
rect 814 -239 815 -191
rect 821 -192 822 -188
rect 919 -239 920 -191
rect 23 -194 24 -188
rect 68 -239 69 -193
rect 72 -194 73 -188
rect 201 -239 202 -193
rect 205 -239 206 -193
rect 352 -194 353 -188
rect 355 -239 356 -193
rect 436 -239 437 -193
rect 485 -194 486 -188
rect 884 -239 885 -193
rect 23 -239 24 -195
rect 100 -196 101 -188
rect 163 -239 164 -195
rect 177 -196 178 -188
rect 184 -239 185 -195
rect 212 -196 213 -188
rect 233 -239 234 -195
rect 268 -196 269 -188
rect 292 -239 293 -195
rect 387 -239 388 -195
rect 422 -196 423 -188
rect 555 -196 556 -188
rect 562 -196 563 -188
rect 562 -239 563 -195
rect 562 -196 563 -188
rect 562 -239 563 -195
rect 660 -196 661 -188
rect 730 -239 731 -195
rect 744 -196 745 -188
rect 765 -239 766 -195
rect 772 -196 773 -188
rect 877 -239 878 -195
rect 30 -239 31 -197
rect 114 -198 115 -188
rect 142 -198 143 -188
rect 212 -239 213 -197
rect 261 -198 262 -188
rect 268 -239 269 -197
rect 296 -198 297 -188
rect 317 -239 318 -197
rect 345 -198 346 -188
rect 905 -239 906 -197
rect 37 -239 38 -199
rect 247 -200 248 -188
rect 303 -239 304 -199
rect 373 -200 374 -188
rect 380 -200 381 -188
rect 555 -239 556 -199
rect 674 -200 675 -188
rect 758 -239 759 -199
rect 786 -200 787 -188
rect 856 -239 857 -199
rect 859 -200 860 -188
rect 933 -239 934 -199
rect 44 -239 45 -201
rect 282 -202 283 -188
rect 352 -239 353 -201
rect 639 -202 640 -188
rect 702 -202 703 -188
rect 744 -239 745 -201
rect 751 -202 752 -188
rect 786 -239 787 -201
rect 793 -202 794 -188
rect 863 -239 864 -201
rect 72 -239 73 -203
rect 156 -204 157 -188
rect 170 -204 171 -188
rect 177 -239 178 -203
rect 187 -204 188 -188
rect 296 -239 297 -203
rect 359 -204 360 -188
rect 359 -239 360 -203
rect 359 -204 360 -188
rect 359 -239 360 -203
rect 373 -239 374 -203
rect 394 -204 395 -188
rect 408 -204 409 -188
rect 422 -239 423 -203
rect 495 -239 496 -203
rect 520 -239 521 -203
rect 527 -204 528 -188
rect 674 -239 675 -203
rect 681 -204 682 -188
rect 751 -239 752 -203
rect 800 -204 801 -188
rect 891 -239 892 -203
rect 79 -206 80 -188
rect 240 -239 241 -205
rect 247 -239 248 -205
rect 275 -206 276 -188
rect 408 -239 409 -205
rect 537 -206 538 -188
rect 541 -206 542 -188
rect 576 -239 577 -205
rect 604 -206 605 -188
rect 639 -239 640 -205
rect 681 -239 682 -205
rect 688 -206 689 -188
rect 709 -206 710 -188
rect 772 -239 773 -205
rect 800 -239 801 -205
rect 842 -239 843 -205
rect 79 -239 80 -207
rect 348 -208 349 -188
rect 450 -208 451 -188
rect 527 -239 528 -207
rect 534 -239 535 -207
rect 590 -208 591 -188
rect 625 -208 626 -188
rect 688 -239 689 -207
rect 737 -208 738 -188
rect 793 -239 794 -207
rect 807 -208 808 -188
rect 940 -239 941 -207
rect 107 -210 108 -188
rect 394 -239 395 -209
rect 429 -210 430 -188
rect 450 -239 451 -209
rect 478 -210 479 -188
rect 541 -239 542 -209
rect 548 -210 549 -188
rect 625 -239 626 -209
rect 646 -210 647 -188
rect 709 -239 710 -209
rect 716 -210 717 -188
rect 807 -239 808 -209
rect 821 -239 822 -209
rect 849 -210 850 -188
rect 58 -212 59 -188
rect 548 -239 549 -211
rect 583 -212 584 -188
rect 604 -239 605 -211
rect 667 -212 668 -188
rect 737 -239 738 -211
rect 779 -212 780 -188
rect 849 -239 850 -211
rect 51 -214 52 -188
rect 58 -239 59 -213
rect 107 -239 108 -213
rect 135 -239 136 -213
rect 142 -239 143 -213
rect 149 -214 150 -188
rect 187 -239 188 -213
rect 583 -239 584 -213
rect 695 -214 696 -188
rect 716 -239 717 -213
rect 723 -214 724 -188
rect 779 -239 780 -213
rect 828 -214 829 -188
rect 926 -239 927 -213
rect 51 -239 52 -215
rect 65 -239 66 -215
rect 114 -239 115 -215
rect 128 -216 129 -188
rect 149 -239 150 -215
rect 219 -216 220 -188
rect 254 -216 255 -188
rect 282 -239 283 -215
rect 324 -216 325 -188
rect 429 -239 430 -215
rect 464 -239 465 -215
rect 828 -239 829 -215
rect 835 -216 836 -188
rect 898 -239 899 -215
rect 121 -218 122 -188
rect 128 -239 129 -217
rect 191 -218 192 -188
rect 254 -239 255 -217
rect 275 -239 276 -217
rect 618 -218 619 -188
rect 632 -218 633 -188
rect 695 -239 696 -217
rect 93 -220 94 -188
rect 191 -239 192 -219
rect 310 -220 311 -188
rect 324 -239 325 -219
rect 345 -239 346 -219
rect 478 -239 479 -219
rect 499 -220 500 -188
rect 660 -239 661 -219
rect 93 -239 94 -221
rect 912 -239 913 -221
rect 121 -239 122 -223
rect 229 -239 230 -223
rect 467 -224 468 -188
rect 667 -239 668 -223
rect 173 -239 174 -225
rect 310 -239 311 -225
rect 366 -226 367 -188
rect 467 -239 468 -225
rect 471 -226 472 -188
rect 499 -239 500 -225
rect 513 -226 514 -188
rect 702 -239 703 -225
rect 289 -228 290 -188
rect 366 -239 367 -227
rect 457 -228 458 -188
rect 471 -239 472 -227
rect 506 -228 507 -188
rect 513 -239 514 -227
rect 593 -239 594 -227
rect 835 -239 836 -227
rect 443 -230 444 -188
rect 506 -239 507 -229
rect 597 -230 598 -188
rect 632 -239 633 -229
rect 653 -230 654 -188
rect 723 -239 724 -229
rect 415 -232 416 -188
rect 443 -239 444 -231
rect 611 -232 612 -188
rect 618 -239 619 -231
rect 401 -234 402 -188
rect 415 -239 416 -233
rect 425 -234 426 -188
rect 653 -239 654 -233
rect 100 -239 101 -235
rect 401 -239 402 -235
rect 569 -236 570 -188
rect 611 -239 612 -235
rect 226 -238 227 -188
rect 569 -239 570 -237
rect 30 -249 31 -247
rect 159 -249 160 -247
rect 170 -249 171 -247
rect 212 -249 213 -247
rect 233 -249 234 -247
rect 292 -249 293 -247
rect 352 -310 353 -248
rect 506 -249 507 -247
rect 534 -249 535 -247
rect 534 -310 535 -248
rect 534 -249 535 -247
rect 534 -310 535 -248
rect 579 -310 580 -248
rect 772 -249 773 -247
rect 877 -249 878 -247
rect 961 -310 962 -248
rect 975 -249 976 -247
rect 982 -310 983 -248
rect 1087 -249 1088 -247
rect 1094 -310 1095 -248
rect 33 -310 34 -250
rect 485 -251 486 -247
rect 488 -310 489 -250
rect 779 -251 780 -247
rect 877 -310 878 -250
rect 933 -251 934 -247
rect 947 -251 948 -247
rect 975 -310 976 -250
rect 37 -253 38 -247
rect 198 -310 199 -252
rect 208 -310 209 -252
rect 555 -253 556 -247
rect 586 -310 587 -252
rect 828 -253 829 -247
rect 905 -253 906 -247
rect 905 -310 906 -252
rect 905 -253 906 -247
rect 905 -310 906 -252
rect 37 -310 38 -254
rect 89 -255 90 -247
rect 93 -255 94 -247
rect 247 -255 248 -247
rect 254 -255 255 -247
rect 282 -310 283 -254
rect 380 -255 381 -247
rect 394 -255 395 -247
rect 436 -255 437 -247
rect 506 -310 507 -254
rect 527 -255 528 -247
rect 555 -310 556 -254
rect 593 -255 594 -247
rect 653 -255 654 -247
rect 758 -255 759 -247
rect 772 -310 773 -254
rect 779 -310 780 -254
rect 793 -255 794 -247
rect 828 -310 829 -254
rect 884 -255 885 -247
rect 44 -257 45 -247
rect 289 -310 290 -256
rect 383 -257 384 -247
rect 590 -310 591 -256
rect 600 -257 601 -247
rect 709 -257 710 -247
rect 765 -257 766 -247
rect 800 -310 801 -256
rect 884 -310 885 -256
rect 891 -257 892 -247
rect 47 -310 48 -258
rect 86 -310 87 -258
rect 93 -310 94 -258
rect 303 -259 304 -247
rect 394 -310 395 -258
rect 513 -259 514 -247
rect 520 -259 521 -247
rect 527 -310 528 -258
rect 597 -259 598 -247
rect 765 -310 766 -258
rect 891 -310 892 -258
rect 954 -259 955 -247
rect 58 -310 59 -260
rect 191 -261 192 -247
rect 205 -261 206 -247
rect 254 -310 255 -260
rect 268 -261 269 -247
rect 268 -310 269 -260
rect 268 -261 269 -247
rect 268 -310 269 -260
rect 275 -261 276 -247
rect 481 -261 482 -247
rect 495 -261 496 -247
rect 674 -261 675 -247
rect 702 -261 703 -247
rect 954 -310 955 -260
rect 23 -263 24 -247
rect 191 -310 192 -262
rect 233 -310 234 -262
rect 457 -263 458 -247
rect 464 -263 465 -247
rect 646 -263 647 -247
rect 653 -310 654 -262
rect 730 -263 731 -247
rect 23 -310 24 -264
rect 51 -265 52 -247
rect 65 -310 66 -264
rect 439 -310 440 -264
rect 478 -265 479 -247
rect 835 -265 836 -247
rect 79 -267 80 -247
rect 212 -310 213 -266
rect 338 -267 339 -247
rect 457 -310 458 -266
rect 499 -267 500 -247
rect 513 -310 514 -266
rect 562 -267 563 -247
rect 597 -310 598 -266
rect 604 -267 605 -247
rect 674 -310 675 -266
rect 695 -267 696 -247
rect 730 -310 731 -266
rect 79 -310 80 -268
rect 793 -310 794 -268
rect 82 -310 83 -270
rect 100 -310 101 -270
rect 103 -271 104 -247
rect 128 -271 129 -247
rect 135 -271 136 -247
rect 247 -310 248 -270
rect 331 -271 332 -247
rect 338 -310 339 -270
rect 373 -271 374 -247
rect 520 -310 521 -270
rect 541 -271 542 -247
rect 562 -310 563 -270
rect 583 -271 584 -247
rect 604 -310 605 -270
rect 618 -271 619 -247
rect 646 -310 647 -270
rect 695 -310 696 -270
rect 737 -271 738 -247
rect 107 -273 108 -247
rect 569 -273 570 -247
rect 576 -273 577 -247
rect 618 -310 619 -272
rect 667 -273 668 -247
rect 737 -310 738 -272
rect 117 -275 118 -247
rect 331 -310 332 -274
rect 359 -275 360 -247
rect 373 -310 374 -274
rect 411 -310 412 -274
rect 758 -310 759 -274
rect 121 -277 122 -247
rect 121 -310 122 -276
rect 121 -277 122 -247
rect 121 -310 122 -276
rect 128 -310 129 -276
rect 324 -277 325 -247
rect 359 -310 360 -276
rect 415 -277 416 -247
rect 450 -277 451 -247
rect 478 -310 479 -276
rect 583 -310 584 -276
rect 681 -277 682 -247
rect 702 -310 703 -276
rect 723 -277 724 -247
rect 135 -310 136 -278
rect 261 -279 262 -247
rect 317 -279 318 -247
rect 324 -310 325 -278
rect 415 -310 416 -278
rect 835 -310 836 -278
rect 142 -281 143 -247
rect 275 -310 276 -280
rect 422 -281 423 -247
rect 450 -310 451 -280
rect 471 -281 472 -247
rect 499 -310 500 -280
rect 639 -281 640 -247
rect 667 -310 668 -280
rect 681 -310 682 -280
rect 688 -281 689 -247
rect 709 -310 710 -280
rect 849 -281 850 -247
rect 114 -283 115 -247
rect 688 -310 689 -282
rect 723 -310 724 -282
rect 751 -283 752 -247
rect 849 -310 850 -282
rect 926 -283 927 -247
rect 114 -310 115 -284
rect 163 -285 164 -247
rect 170 -310 171 -284
rect 296 -285 297 -247
rect 422 -310 423 -284
rect 429 -285 430 -247
rect 471 -310 472 -284
rect 814 -285 815 -247
rect 912 -285 913 -247
rect 926 -310 927 -284
rect 145 -310 146 -286
rect 303 -310 304 -286
rect 429 -310 430 -286
rect 443 -287 444 -247
rect 474 -310 475 -286
rect 569 -310 570 -286
rect 625 -287 626 -247
rect 639 -310 640 -286
rect 744 -287 745 -247
rect 751 -310 752 -286
rect 912 -310 913 -286
rect 940 -287 941 -247
rect 156 -289 157 -247
rect 548 -289 549 -247
rect 625 -310 626 -288
rect 660 -289 661 -247
rect 716 -289 717 -247
rect 744 -310 745 -288
rect 821 -289 822 -247
rect 940 -310 941 -288
rect 156 -310 157 -290
rect 205 -310 206 -290
rect 219 -291 220 -247
rect 296 -310 297 -290
rect 401 -291 402 -247
rect 443 -310 444 -290
rect 492 -291 493 -247
rect 814 -310 815 -290
rect 163 -310 164 -292
rect 548 -310 549 -292
rect 632 -293 633 -247
rect 660 -310 661 -292
rect 786 -293 787 -247
rect 821 -310 822 -292
rect 177 -295 178 -247
rect 184 -310 185 -294
rect 219 -310 220 -294
rect 240 -295 241 -247
rect 264 -295 265 -247
rect 317 -310 318 -294
rect 366 -295 367 -247
rect 401 -310 402 -294
rect 492 -310 493 -294
rect 870 -295 871 -247
rect 16 -297 17 -247
rect 177 -310 178 -296
rect 226 -297 227 -247
rect 240 -310 241 -296
rect 310 -297 311 -247
rect 366 -310 367 -296
rect 611 -297 612 -247
rect 632 -310 633 -296
rect 786 -310 787 -296
rect 807 -297 808 -247
rect 870 -310 871 -296
rect 919 -297 920 -247
rect 16 -310 17 -298
rect 464 -310 465 -298
rect 807 -310 808 -298
rect 856 -299 857 -247
rect 863 -299 864 -247
rect 919 -310 920 -298
rect 72 -301 73 -247
rect 310 -310 311 -300
rect 408 -301 409 -247
rect 611 -310 612 -300
rect 842 -301 843 -247
rect 856 -310 857 -300
rect 863 -310 864 -300
rect 898 -301 899 -247
rect 72 -310 73 -302
rect 345 -303 346 -247
rect 842 -310 843 -302
rect 968 -310 969 -302
rect 149 -305 150 -247
rect 345 -310 346 -304
rect 898 -310 899 -304
rect 936 -310 937 -304
rect 149 -310 150 -306
rect 387 -307 388 -247
rect 229 -310 230 -308
rect 261 -310 262 -308
rect 9 -320 10 -318
rect 145 -320 146 -318
rect 156 -320 157 -318
rect 156 -395 157 -319
rect 156 -320 157 -318
rect 156 -395 157 -319
rect 184 -320 185 -318
rect 184 -395 185 -319
rect 184 -320 185 -318
rect 184 -395 185 -319
rect 205 -395 206 -319
rect 208 -320 209 -318
rect 226 -395 227 -319
rect 268 -320 269 -318
rect 296 -320 297 -318
rect 408 -320 409 -318
rect 436 -320 437 -318
rect 926 -320 927 -318
rect 933 -395 934 -319
rect 982 -320 983 -318
rect 999 -395 1000 -319
rect 1066 -395 1067 -319
rect 1094 -320 1095 -318
rect 1108 -395 1109 -319
rect 16 -322 17 -318
rect 474 -322 475 -318
rect 523 -395 524 -321
rect 653 -322 654 -318
rect 681 -322 682 -318
rect 684 -322 685 -318
rect 716 -322 717 -318
rect 905 -322 906 -318
rect 947 -322 948 -318
rect 968 -395 969 -321
rect 16 -395 17 -323
rect 135 -324 136 -318
rect 208 -395 209 -323
rect 292 -324 293 -318
rect 317 -324 318 -318
rect 464 -395 465 -323
rect 527 -324 528 -318
rect 544 -324 545 -318
rect 548 -324 549 -318
rect 961 -324 962 -318
rect 964 -395 965 -323
rect 1052 -395 1053 -323
rect 23 -326 24 -318
rect 117 -395 118 -325
rect 121 -326 122 -318
rect 296 -395 297 -325
rect 331 -326 332 -318
rect 467 -326 468 -318
rect 541 -326 542 -318
rect 954 -326 955 -318
rect 23 -395 24 -327
rect 303 -328 304 -318
rect 345 -328 346 -318
rect 383 -328 384 -318
rect 390 -328 391 -318
rect 520 -328 521 -318
rect 534 -328 535 -318
rect 541 -395 542 -327
rect 548 -395 549 -327
rect 919 -328 920 -318
rect 37 -330 38 -318
rect 51 -395 52 -329
rect 58 -330 59 -318
rect 418 -330 419 -318
rect 443 -330 444 -318
rect 583 -395 584 -329
rect 632 -330 633 -318
rect 653 -395 654 -329
rect 681 -395 682 -329
rect 884 -330 885 -318
rect 898 -330 899 -318
rect 982 -395 983 -329
rect 40 -395 41 -331
rect 58 -395 59 -331
rect 65 -332 66 -318
rect 163 -332 164 -318
rect 212 -332 213 -318
rect 436 -395 437 -331
rect 443 -395 444 -331
rect 488 -332 489 -318
rect 499 -332 500 -318
rect 534 -395 535 -331
rect 579 -395 580 -331
rect 905 -395 906 -331
rect 44 -395 45 -333
rect 145 -395 146 -333
rect 212 -395 213 -333
rect 485 -334 486 -318
rect 618 -334 619 -318
rect 632 -395 633 -333
rect 716 -395 717 -333
rect 814 -334 815 -318
rect 821 -334 822 -318
rect 926 -395 927 -333
rect 65 -395 66 -335
rect 107 -336 108 -318
rect 121 -395 122 -335
rect 324 -336 325 -318
rect 338 -336 339 -318
rect 345 -395 346 -335
rect 352 -336 353 -318
rect 355 -352 356 -335
rect 359 -336 360 -318
rect 415 -395 416 -335
rect 422 -336 423 -318
rect 499 -395 500 -335
rect 786 -336 787 -318
rect 884 -395 885 -335
rect 901 -395 902 -335
rect 975 -336 976 -318
rect 30 -338 31 -318
rect 422 -395 423 -337
rect 453 -395 454 -337
rect 772 -338 773 -318
rect 807 -338 808 -318
rect 821 -395 822 -337
rect 828 -338 829 -318
rect 975 -395 976 -337
rect 93 -340 94 -318
rect 289 -395 290 -339
rect 352 -395 353 -339
rect 394 -340 395 -318
rect 401 -340 402 -318
rect 408 -395 409 -339
rect 457 -340 458 -318
rect 527 -395 528 -339
rect 702 -340 703 -318
rect 772 -395 773 -339
rect 835 -340 836 -318
rect 1010 -395 1011 -339
rect 93 -395 94 -341
rect 180 -395 181 -341
rect 191 -342 192 -318
rect 618 -395 619 -341
rect 639 -342 640 -318
rect 702 -395 703 -341
rect 744 -342 745 -318
rect 786 -395 787 -341
rect 842 -342 843 -318
rect 947 -395 948 -341
rect 100 -344 101 -318
rect 107 -395 108 -343
rect 135 -395 136 -343
rect 163 -395 164 -343
rect 254 -344 255 -318
rect 268 -395 269 -343
rect 275 -344 276 -318
rect 303 -395 304 -343
rect 359 -395 360 -343
rect 478 -344 479 -318
rect 506 -395 507 -343
rect 828 -395 829 -343
rect 849 -344 850 -318
rect 1017 -395 1018 -343
rect 79 -346 80 -318
rect 478 -395 479 -345
rect 590 -346 591 -318
rect 639 -395 640 -345
rect 723 -346 724 -318
rect 849 -395 850 -345
rect 863 -346 864 -318
rect 989 -395 990 -345
rect 79 -395 80 -347
rect 170 -348 171 -318
rect 219 -348 220 -318
rect 254 -395 255 -347
rect 261 -348 262 -318
rect 331 -395 332 -347
rect 380 -348 381 -318
rect 919 -395 920 -347
rect 72 -350 73 -318
rect 380 -395 381 -349
rect 394 -395 395 -349
rect 474 -395 475 -349
rect 723 -395 724 -349
rect 751 -350 752 -318
rect 807 -395 808 -349
rect 870 -350 871 -318
rect 1003 -395 1004 -349
rect 72 -395 73 -351
rect 86 -352 87 -318
rect 100 -395 101 -351
rect 110 -352 111 -318
rect 149 -352 150 -318
rect 485 -395 486 -351
rect 569 -352 570 -318
rect 590 -395 591 -351
rect 684 -395 685 -351
rect 744 -395 745 -351
rect 758 -352 759 -318
rect 863 -395 864 -351
rect 870 -395 871 -351
rect 912 -352 913 -318
rect 86 -395 87 -353
rect 366 -354 367 -318
rect 401 -395 402 -353
rect 814 -395 815 -353
rect 877 -354 878 -318
rect 1024 -395 1025 -353
rect 149 -395 150 -355
rect 247 -356 248 -318
rect 275 -395 276 -355
rect 450 -356 451 -318
rect 555 -356 556 -318
rect 569 -395 570 -355
rect 586 -356 587 -318
rect 758 -395 759 -355
rect 765 -356 766 -318
rect 877 -395 878 -355
rect 891 -356 892 -318
rect 912 -395 913 -355
rect 191 -395 192 -357
rect 450 -395 451 -357
rect 513 -358 514 -318
rect 555 -395 556 -357
rect 730 -358 731 -318
rect 765 -395 766 -357
rect 793 -358 794 -318
rect 891 -395 892 -357
rect 198 -360 199 -318
rect 261 -395 262 -359
rect 282 -360 283 -318
rect 324 -395 325 -359
rect 366 -395 367 -359
rect 551 -360 552 -318
rect 688 -360 689 -318
rect 793 -395 794 -359
rect 800 -360 801 -318
rect 842 -395 843 -359
rect 114 -362 115 -318
rect 282 -395 283 -361
rect 404 -395 405 -361
rect 835 -395 836 -361
rect 128 -364 129 -318
rect 198 -395 199 -363
rect 219 -395 220 -363
rect 565 -395 566 -363
rect 611 -364 612 -318
rect 688 -395 689 -363
rect 695 -364 696 -318
rect 800 -395 801 -363
rect 33 -395 34 -365
rect 128 -395 129 -365
rect 240 -366 241 -318
rect 247 -395 248 -365
rect 429 -366 430 -318
rect 457 -395 458 -365
rect 492 -366 493 -318
rect 513 -395 514 -365
rect 611 -395 612 -365
rect 674 -366 675 -318
rect 719 -366 720 -318
rect 730 -395 731 -365
rect 737 -366 738 -318
rect 751 -395 752 -365
rect 240 -395 241 -367
rect 936 -368 937 -318
rect 429 -395 430 -369
rect 520 -395 521 -369
rect 625 -370 626 -318
rect 695 -395 696 -369
rect 737 -395 738 -369
rect 940 -370 941 -318
rect 492 -395 493 -371
rect 954 -395 955 -371
rect 495 -395 496 -373
rect 551 -395 552 -373
rect 597 -374 598 -318
rect 625 -395 626 -373
rect 660 -374 661 -318
rect 674 -395 675 -373
rect 856 -374 857 -318
rect 940 -395 941 -373
rect 562 -376 563 -318
rect 597 -395 598 -375
rect 646 -376 647 -318
rect 660 -395 661 -375
rect 779 -376 780 -318
rect 856 -395 857 -375
rect 338 -395 339 -377
rect 646 -395 647 -377
rect 779 -395 780 -377
rect 961 -395 962 -377
rect 562 -395 563 -379
rect 709 -380 710 -318
rect 667 -382 668 -318
rect 709 -395 710 -381
rect 604 -384 605 -318
rect 667 -395 668 -383
rect 387 -386 388 -318
rect 604 -395 605 -385
rect 373 -388 374 -318
rect 387 -395 388 -387
rect 310 -390 311 -318
rect 373 -395 374 -389
rect 233 -392 234 -318
rect 310 -395 311 -391
rect 177 -394 178 -318
rect 233 -395 234 -393
rect 16 -405 17 -403
rect 138 -405 139 -403
rect 142 -405 143 -403
rect 149 -405 150 -403
rect 180 -405 181 -403
rect 198 -405 199 -403
rect 233 -405 234 -403
rect 275 -464 276 -404
rect 282 -405 283 -403
rect 285 -405 286 -403
rect 306 -464 307 -404
rect 324 -405 325 -403
rect 331 -405 332 -403
rect 404 -405 405 -403
rect 422 -464 423 -404
rect 754 -464 755 -404
rect 800 -405 801 -403
rect 1045 -464 1046 -404
rect 1066 -405 1067 -403
rect 1139 -464 1140 -404
rect 16 -464 17 -406
rect 51 -407 52 -403
rect 58 -407 59 -403
rect 198 -464 199 -406
rect 233 -464 234 -406
rect 565 -464 566 -406
rect 576 -464 577 -406
rect 590 -407 591 -403
rect 600 -464 601 -406
rect 870 -407 871 -403
rect 877 -407 878 -403
rect 1101 -464 1102 -406
rect 1108 -407 1109 -403
rect 1150 -464 1151 -406
rect 23 -409 24 -403
rect 390 -464 391 -408
rect 401 -464 402 -408
rect 793 -409 794 -403
rect 800 -464 801 -408
rect 807 -409 808 -403
rect 863 -409 864 -403
rect 1115 -464 1116 -408
rect 23 -464 24 -410
rect 114 -411 115 -403
rect 142 -464 143 -410
rect 173 -411 174 -403
rect 184 -411 185 -403
rect 184 -464 185 -410
rect 184 -411 185 -403
rect 184 -464 185 -410
rect 191 -411 192 -403
rect 205 -464 206 -410
rect 247 -411 248 -403
rect 250 -423 251 -410
rect 254 -411 255 -403
rect 320 -411 321 -403
rect 331 -464 332 -410
rect 485 -411 486 -403
rect 502 -464 503 -410
rect 996 -411 997 -403
rect 1003 -411 1004 -403
rect 1087 -464 1088 -410
rect 37 -464 38 -412
rect 212 -413 213 -403
rect 247 -464 248 -412
rect 268 -413 269 -403
rect 278 -413 279 -403
rect 282 -464 283 -412
rect 289 -413 290 -403
rect 296 -413 297 -403
rect 324 -464 325 -412
rect 338 -413 339 -403
rect 429 -413 430 -403
rect 436 -413 437 -403
rect 492 -413 493 -403
rect 509 -464 510 -412
rect 695 -413 696 -403
rect 740 -464 741 -412
rect 1080 -464 1081 -412
rect 51 -464 52 -414
rect 110 -464 111 -414
rect 128 -415 129 -403
rect 191 -464 192 -414
rect 219 -415 220 -403
rect 296 -464 297 -414
rect 317 -415 318 -403
rect 450 -464 451 -414
rect 478 -415 479 -403
rect 492 -464 493 -414
rect 523 -464 524 -414
rect 898 -464 899 -414
rect 919 -415 920 -403
rect 996 -464 997 -414
rect 1010 -415 1011 -403
rect 1108 -464 1109 -414
rect 58 -464 59 -416
rect 79 -417 80 -403
rect 100 -417 101 -403
rect 100 -464 101 -416
rect 100 -417 101 -403
rect 100 -464 101 -416
rect 107 -417 108 -403
rect 114 -464 115 -416
rect 128 -464 129 -416
rect 156 -417 157 -403
rect 219 -464 220 -416
rect 303 -417 304 -403
rect 317 -464 318 -416
rect 380 -417 381 -403
rect 425 -417 426 -403
rect 1066 -464 1067 -416
rect 65 -419 66 -403
rect 89 -464 90 -418
rect 145 -419 146 -403
rect 208 -419 209 -403
rect 240 -419 241 -403
rect 338 -464 339 -418
rect 341 -419 342 -403
rect 345 -419 346 -403
rect 359 -464 360 -418
rect 415 -419 416 -403
rect 429 -464 430 -418
rect 551 -419 552 -403
rect 555 -419 556 -403
rect 555 -464 556 -418
rect 555 -419 556 -403
rect 555 -464 556 -418
rect 586 -464 587 -418
rect 716 -419 717 -403
rect 730 -419 731 -403
rect 919 -464 920 -418
rect 947 -419 948 -403
rect 1038 -464 1039 -418
rect 1041 -419 1042 -403
rect 1052 -419 1053 -403
rect 44 -421 45 -403
rect 947 -464 948 -420
rect 954 -421 955 -403
rect 1052 -464 1053 -420
rect 44 -464 45 -422
rect 278 -464 279 -422
rect 285 -464 286 -422
rect 289 -464 290 -422
rect 345 -464 346 -422
rect 499 -423 500 -403
rect 548 -464 549 -422
rect 1031 -423 1032 -403
rect 65 -464 66 -424
rect 352 -425 353 -403
rect 366 -425 367 -403
rect 436 -464 437 -424
rect 485 -464 486 -424
rect 527 -425 528 -403
rect 590 -464 591 -424
rect 597 -425 598 -403
rect 611 -425 612 -403
rect 611 -464 612 -424
rect 611 -425 612 -403
rect 611 -464 612 -424
rect 646 -425 647 -403
rect 954 -464 955 -424
rect 975 -425 976 -403
rect 1094 -464 1095 -424
rect 72 -427 73 -403
rect 135 -464 136 -426
rect 156 -464 157 -426
rect 411 -464 412 -426
rect 478 -464 479 -426
rect 597 -464 598 -426
rect 639 -427 640 -403
rect 646 -464 647 -426
rect 660 -427 661 -403
rect 695 -464 696 -426
rect 709 -427 710 -403
rect 716 -464 717 -426
rect 744 -427 745 -403
rect 877 -464 878 -426
rect 905 -427 906 -403
rect 1010 -464 1011 -426
rect 1017 -427 1018 -403
rect 1122 -464 1123 -426
rect 30 -464 31 -428
rect 660 -464 661 -428
rect 674 -429 675 -403
rect 709 -464 710 -428
rect 744 -464 745 -428
rect 758 -429 759 -403
rect 772 -429 773 -403
rect 1003 -464 1004 -428
rect 1024 -429 1025 -403
rect 1129 -464 1130 -428
rect 72 -464 73 -430
rect 86 -431 87 -403
rect 93 -431 94 -403
rect 352 -464 353 -430
rect 373 -431 374 -403
rect 373 -464 374 -430
rect 373 -431 374 -403
rect 373 -464 374 -430
rect 380 -464 381 -430
rect 901 -431 902 -403
rect 926 -431 927 -403
rect 1024 -464 1025 -430
rect 12 -464 13 -432
rect 86 -464 87 -432
rect 93 -464 94 -432
rect 121 -433 122 -403
rect 240 -464 241 -432
rect 635 -464 636 -432
rect 653 -433 654 -403
rect 674 -464 675 -432
rect 688 -433 689 -403
rect 730 -464 731 -432
rect 765 -433 766 -403
rect 772 -464 773 -432
rect 793 -464 794 -432
rect 849 -433 850 -403
rect 870 -464 871 -432
rect 912 -433 913 -403
rect 926 -464 927 -432
rect 989 -433 990 -403
rect 79 -464 80 -434
rect 513 -435 514 -403
rect 527 -464 528 -434
rect 562 -464 563 -434
rect 569 -435 570 -403
rect 765 -464 766 -434
rect 779 -435 780 -403
rect 989 -464 990 -434
rect 121 -464 122 -436
rect 163 -437 164 -403
rect 254 -464 255 -436
rect 394 -437 395 -403
rect 408 -437 409 -403
rect 415 -464 416 -436
rect 457 -437 458 -403
rect 513 -464 514 -436
rect 534 -437 535 -403
rect 569 -464 570 -436
rect 625 -437 626 -403
rect 639 -464 640 -436
rect 653 -464 654 -436
rect 737 -437 738 -403
rect 807 -464 808 -436
rect 821 -437 822 -403
rect 835 -437 836 -403
rect 975 -464 976 -436
rect 982 -437 983 -403
rect 1073 -464 1074 -436
rect 149 -464 150 -438
rect 457 -464 458 -438
rect 471 -464 472 -438
rect 779 -464 780 -438
rect 814 -439 815 -403
rect 905 -464 906 -438
rect 940 -439 941 -403
rect 1031 -464 1032 -438
rect 163 -464 164 -440
rect 177 -441 178 -403
rect 268 -464 269 -440
rect 443 -441 444 -403
rect 520 -441 521 -403
rect 821 -464 822 -440
rect 835 -464 836 -440
rect 884 -441 885 -403
rect 940 -464 941 -440
rect 961 -441 962 -403
rect 982 -464 983 -440
rect 1059 -464 1060 -440
rect 170 -443 171 -403
rect 814 -464 815 -442
rect 842 -443 843 -403
rect 863 -464 864 -442
rect 884 -464 885 -442
rect 968 -443 969 -403
rect 170 -464 171 -444
rect 226 -445 227 -403
rect 303 -464 304 -444
rect 842 -464 843 -444
rect 856 -445 857 -403
rect 968 -464 969 -444
rect 177 -464 178 -446
rect 310 -447 311 -403
rect 387 -447 388 -403
rect 394 -464 395 -446
rect 408 -464 409 -446
rect 1017 -464 1018 -446
rect 310 -464 311 -448
rect 579 -449 580 -403
rect 604 -449 605 -403
rect 625 -464 626 -448
rect 681 -449 682 -403
rect 912 -464 913 -448
rect 933 -449 934 -403
rect 961 -464 962 -448
rect 443 -464 444 -450
rect 464 -451 465 -403
rect 474 -464 475 -450
rect 856 -464 857 -450
rect 891 -451 892 -403
rect 933 -464 934 -450
rect 464 -464 465 -452
rect 737 -464 738 -452
rect 828 -453 829 -403
rect 891 -464 892 -452
rect 520 -464 521 -454
rect 667 -455 668 -403
rect 681 -464 682 -454
rect 1048 -455 1049 -403
rect 534 -464 535 -456
rect 541 -457 542 -403
rect 604 -464 605 -456
rect 618 -457 619 -403
rect 632 -457 633 -403
rect 667 -464 668 -456
rect 688 -464 689 -456
rect 702 -457 703 -403
rect 723 -457 724 -403
rect 758 -464 759 -456
rect 786 -457 787 -403
rect 828 -464 829 -456
rect 229 -464 230 -458
rect 541 -464 542 -458
rect 583 -459 584 -403
rect 618 -464 619 -458
rect 723 -464 724 -458
rect 849 -464 850 -458
rect 366 -464 367 -460
rect 583 -464 584 -460
rect 751 -461 752 -403
rect 786 -464 787 -460
rect 404 -464 405 -462
rect 702 -464 703 -462
rect 9 -559 10 -473
rect 310 -474 311 -472
rect 324 -474 325 -472
rect 345 -559 346 -473
rect 348 -474 349 -472
rect 635 -474 636 -472
rect 660 -474 661 -472
rect 968 -474 969 -472
rect 975 -474 976 -472
rect 1143 -474 1144 -472
rect 1174 -559 1175 -473
rect 1178 -559 1179 -473
rect 16 -476 17 -472
rect 110 -476 111 -472
rect 135 -559 136 -475
rect 142 -476 143 -472
rect 156 -476 157 -472
rect 530 -476 531 -472
rect 537 -559 538 -475
rect 1045 -476 1046 -472
rect 16 -559 17 -477
rect 100 -478 101 -472
rect 107 -559 108 -477
rect 254 -478 255 -472
rect 261 -478 262 -472
rect 278 -478 279 -472
rect 296 -478 297 -472
rect 310 -559 311 -477
rect 397 -559 398 -477
rect 520 -559 521 -477
rect 527 -478 528 -472
rect 989 -478 990 -472
rect 1045 -559 1046 -477
rect 1059 -478 1060 -472
rect 37 -480 38 -472
rect 303 -480 304 -472
rect 401 -480 402 -472
rect 513 -480 514 -472
rect 527 -559 528 -479
rect 534 -480 535 -472
rect 541 -480 542 -472
rect 541 -559 542 -479
rect 541 -480 542 -472
rect 541 -559 542 -479
rect 555 -480 556 -472
rect 555 -559 556 -479
rect 555 -480 556 -472
rect 555 -559 556 -479
rect 562 -480 563 -472
rect 1122 -480 1123 -472
rect 37 -559 38 -481
rect 201 -559 202 -481
rect 205 -482 206 -472
rect 226 -559 227 -481
rect 240 -482 241 -472
rect 296 -559 297 -481
rect 352 -482 353 -472
rect 401 -559 402 -481
rect 436 -482 437 -472
rect 600 -482 601 -472
rect 632 -482 633 -472
rect 1129 -482 1130 -472
rect 23 -484 24 -472
rect 205 -559 206 -483
rect 219 -484 220 -472
rect 390 -484 391 -472
rect 415 -484 416 -472
rect 436 -559 437 -483
rect 450 -484 451 -472
rect 663 -559 664 -483
rect 695 -484 696 -472
rect 737 -559 738 -483
rect 751 -559 752 -483
rect 856 -484 857 -472
rect 870 -484 871 -472
rect 968 -559 969 -483
rect 975 -559 976 -483
rect 996 -484 997 -472
rect 1059 -559 1060 -483
rect 1108 -484 1109 -472
rect 1122 -559 1123 -483
rect 1139 -484 1140 -472
rect 23 -559 24 -485
rect 30 -486 31 -472
rect 72 -486 73 -472
rect 275 -559 276 -485
rect 289 -486 290 -472
rect 303 -559 304 -485
rect 380 -486 381 -472
rect 513 -559 514 -485
rect 565 -559 566 -485
rect 1094 -486 1095 -472
rect 58 -488 59 -472
rect 380 -559 381 -487
rect 415 -559 416 -487
rect 478 -488 479 -472
rect 506 -559 507 -487
rect 730 -488 731 -472
rect 733 -559 734 -487
rect 1101 -488 1102 -472
rect 58 -559 59 -489
rect 373 -490 374 -472
rect 450 -559 451 -489
rect 485 -490 486 -472
rect 583 -559 584 -489
rect 590 -490 591 -472
rect 593 -559 594 -489
rect 1115 -490 1116 -472
rect 79 -492 80 -472
rect 499 -559 500 -491
rect 586 -492 587 -472
rect 1003 -492 1004 -472
rect 1010 -492 1011 -472
rect 1101 -559 1102 -491
rect 1115 -559 1116 -491
rect 1150 -492 1151 -472
rect 86 -494 87 -472
rect 947 -494 948 -472
rect 961 -494 962 -472
rect 982 -559 983 -493
rect 989 -559 990 -493
rect 1024 -494 1025 -472
rect 86 -559 87 -495
rect 114 -496 115 -472
rect 142 -559 143 -495
rect 366 -496 367 -472
rect 457 -559 458 -495
rect 842 -496 843 -472
rect 961 -559 962 -495
rect 1017 -496 1018 -472
rect 93 -498 94 -472
rect 156 -559 157 -497
rect 166 -559 167 -497
rect 1066 -498 1067 -472
rect 93 -559 94 -499
rect 121 -500 122 -472
rect 170 -500 171 -472
rect 219 -559 220 -499
rect 240 -559 241 -499
rect 247 -500 248 -472
rect 261 -559 262 -499
rect 429 -500 430 -472
rect 460 -500 461 -472
rect 940 -500 941 -472
rect 996 -559 997 -499
rect 1038 -500 1039 -472
rect 100 -559 101 -501
rect 128 -502 129 -472
rect 149 -502 150 -472
rect 170 -559 171 -501
rect 177 -502 178 -472
rect 254 -559 255 -501
rect 289 -559 290 -501
rect 320 -559 321 -501
rect 331 -502 332 -472
rect 373 -559 374 -501
rect 429 -559 430 -501
rect 509 -502 510 -472
rect 611 -502 612 -472
rect 856 -559 857 -501
rect 884 -502 885 -472
rect 1066 -559 1067 -501
rect 44 -504 45 -472
rect 331 -559 332 -503
rect 443 -504 444 -472
rect 509 -559 510 -503
rect 548 -504 549 -472
rect 611 -559 612 -503
rect 632 -559 633 -503
rect 653 -504 654 -472
rect 660 -559 661 -503
rect 940 -559 941 -503
rect 1003 -559 1004 -503
rect 1052 -504 1053 -472
rect 44 -559 45 -505
rect 317 -506 318 -472
rect 387 -506 388 -472
rect 1052 -559 1053 -505
rect 110 -559 111 -507
rect 177 -559 178 -507
rect 184 -508 185 -472
rect 184 -559 185 -507
rect 184 -508 185 -472
rect 184 -559 185 -507
rect 191 -508 192 -472
rect 324 -559 325 -507
rect 471 -508 472 -472
rect 569 -508 570 -472
rect 604 -508 605 -472
rect 653 -559 654 -507
rect 723 -508 724 -472
rect 905 -508 906 -472
rect 1010 -559 1011 -507
rect 1031 -508 1032 -472
rect 33 -559 34 -509
rect 604 -559 605 -509
rect 730 -559 731 -509
rect 1024 -559 1025 -509
rect 1031 -559 1032 -509
rect 1080 -510 1081 -472
rect 114 -559 115 -511
rect 394 -512 395 -472
rect 478 -559 479 -511
rect 492 -512 493 -472
rect 502 -512 503 -472
rect 723 -559 724 -511
rect 754 -512 755 -472
rect 814 -512 815 -472
rect 828 -512 829 -472
rect 842 -559 843 -511
rect 849 -512 850 -472
rect 884 -559 885 -511
rect 898 -512 899 -472
rect 905 -559 906 -511
rect 1017 -559 1018 -511
rect 1073 -512 1074 -472
rect 1080 -559 1081 -511
rect 1087 -512 1088 -472
rect 128 -559 129 -513
rect 408 -514 409 -472
rect 485 -559 486 -513
rect 572 -559 573 -513
rect 597 -514 598 -472
rect 1087 -559 1088 -513
rect 152 -559 153 -515
rect 569 -559 570 -515
rect 597 -559 598 -515
rect 877 -516 878 -472
rect 926 -516 927 -472
rect 1073 -559 1074 -515
rect 163 -518 164 -472
rect 471 -559 472 -517
rect 492 -559 493 -517
rect 628 -559 629 -517
rect 765 -518 766 -472
rect 1094 -559 1095 -517
rect 191 -559 192 -519
rect 695 -559 696 -519
rect 779 -520 780 -472
rect 828 -559 829 -519
rect 835 -520 836 -472
rect 947 -559 948 -519
rect 247 -559 248 -521
rect 404 -522 405 -472
rect 422 -522 423 -472
rect 835 -559 836 -521
rect 877 -559 878 -521
rect 912 -522 913 -472
rect 121 -559 122 -523
rect 422 -559 423 -523
rect 551 -559 552 -523
rect 926 -559 927 -523
rect 268 -526 269 -472
rect 443 -559 444 -525
rect 688 -526 689 -472
rect 765 -559 766 -525
rect 786 -526 787 -472
rect 814 -559 815 -525
rect 821 -526 822 -472
rect 898 -559 899 -525
rect 268 -559 269 -527
rect 282 -528 283 -472
rect 317 -559 318 -527
rect 359 -528 360 -472
rect 667 -528 668 -472
rect 688 -559 689 -527
rect 716 -528 717 -472
rect 779 -559 780 -527
rect 793 -528 794 -472
rect 849 -559 850 -527
rect 891 -528 892 -472
rect 912 -559 913 -527
rect 138 -530 139 -472
rect 359 -559 360 -529
rect 639 -530 640 -472
rect 667 -559 668 -529
rect 681 -530 682 -472
rect 716 -559 717 -529
rect 744 -530 745 -472
rect 786 -559 787 -529
rect 800 -530 801 -472
rect 821 -559 822 -529
rect 863 -530 864 -472
rect 891 -559 892 -529
rect 233 -532 234 -472
rect 282 -559 283 -531
rect 355 -559 356 -531
rect 793 -559 794 -531
rect 807 -532 808 -472
rect 1038 -559 1039 -531
rect 51 -534 52 -472
rect 233 -559 234 -533
rect 408 -559 409 -533
rect 800 -559 801 -533
rect 863 -559 864 -533
rect 954 -534 955 -472
rect 51 -559 52 -535
rect 338 -536 339 -472
rect 548 -559 549 -535
rect 681 -559 682 -535
rect 744 -559 745 -535
rect 758 -536 759 -472
rect 772 -536 773 -472
rect 807 -559 808 -535
rect 933 -536 934 -472
rect 954 -559 955 -535
rect 338 -559 339 -537
rect 390 -559 391 -537
rect 625 -538 626 -472
rect 639 -559 640 -537
rect 702 -538 703 -472
rect 772 -559 773 -537
rect 919 -538 920 -472
rect 933 -559 934 -537
rect 562 -559 563 -539
rect 919 -559 920 -539
rect 674 -542 675 -472
rect 702 -559 703 -541
rect 709 -542 710 -472
rect 758 -559 759 -541
rect 646 -544 647 -472
rect 674 -559 675 -543
rect 709 -559 710 -543
rect 870 -559 871 -543
rect 618 -546 619 -472
rect 646 -559 647 -545
rect 576 -548 577 -472
rect 618 -559 619 -547
rect 65 -550 66 -472
rect 576 -559 577 -549
rect 65 -559 66 -551
rect 198 -552 199 -472
rect 198 -559 199 -553
rect 464 -554 465 -472
rect 215 -556 216 -472
rect 464 -559 465 -555
rect 194 -559 195 -557
rect 215 -559 216 -557
rect 2 -569 3 -567
rect 509 -569 510 -567
rect 534 -650 535 -568
rect 541 -569 542 -567
rect 548 -569 549 -567
rect 870 -569 871 -567
rect 1059 -569 1060 -567
rect 1108 -650 1109 -568
rect 1115 -569 1116 -567
rect 1115 -650 1116 -568
rect 1115 -569 1116 -567
rect 1115 -650 1116 -568
rect 1122 -569 1123 -567
rect 1122 -650 1123 -568
rect 1122 -569 1123 -567
rect 1122 -650 1123 -568
rect 1178 -569 1179 -567
rect 1178 -650 1179 -568
rect 1178 -569 1179 -567
rect 1178 -650 1179 -568
rect 9 -571 10 -567
rect 72 -571 73 -567
rect 82 -571 83 -567
rect 709 -650 710 -570
rect 712 -571 713 -567
rect 898 -571 899 -567
rect 1087 -571 1088 -567
rect 1129 -650 1130 -570
rect 9 -650 10 -572
rect 380 -573 381 -567
rect 408 -573 409 -567
rect 835 -573 836 -567
rect 842 -573 843 -567
rect 898 -650 899 -572
rect 1024 -573 1025 -567
rect 1087 -650 1088 -572
rect 1101 -573 1102 -567
rect 1136 -650 1137 -572
rect 16 -575 17 -567
rect 870 -650 871 -574
rect 975 -575 976 -567
rect 1024 -650 1025 -574
rect 16 -650 17 -576
rect 86 -577 87 -567
rect 121 -577 122 -567
rect 562 -577 563 -567
rect 569 -577 570 -567
rect 1038 -577 1039 -567
rect 23 -579 24 -567
rect 541 -650 542 -578
rect 548 -650 549 -578
rect 1059 -650 1060 -578
rect 23 -650 24 -580
rect 418 -650 419 -580
rect 443 -581 444 -567
rect 572 -581 573 -567
rect 600 -581 601 -567
rect 884 -581 885 -567
rect 919 -581 920 -567
rect 1038 -650 1039 -580
rect 30 -583 31 -567
rect 79 -583 80 -567
rect 86 -650 87 -582
rect 296 -583 297 -567
rect 303 -583 304 -567
rect 303 -650 304 -582
rect 303 -583 304 -567
rect 303 -650 304 -582
rect 338 -583 339 -567
rect 387 -650 388 -582
rect 464 -583 465 -567
rect 691 -650 692 -582
rect 702 -583 703 -567
rect 702 -650 703 -582
rect 702 -583 703 -567
rect 702 -650 703 -582
rect 733 -583 734 -567
rect 744 -583 745 -567
rect 751 -583 752 -567
rect 919 -650 920 -582
rect 968 -583 969 -567
rect 975 -650 976 -582
rect 30 -650 31 -584
rect 261 -585 262 -567
rect 268 -585 269 -567
rect 352 -585 353 -567
rect 380 -650 381 -584
rect 492 -585 493 -567
rect 506 -585 507 -567
rect 1101 -650 1102 -584
rect 33 -587 34 -567
rect 411 -587 412 -567
rect 471 -587 472 -567
rect 597 -650 598 -586
rect 604 -587 605 -567
rect 1066 -587 1067 -567
rect 37 -589 38 -567
rect 187 -650 188 -588
rect 191 -650 192 -588
rect 226 -589 227 -567
rect 254 -589 255 -567
rect 502 -650 503 -588
rect 513 -589 514 -567
rect 562 -650 563 -588
rect 604 -650 605 -588
rect 961 -589 962 -567
rect 1003 -589 1004 -567
rect 1066 -650 1067 -588
rect 37 -650 38 -590
rect 100 -591 101 -567
rect 107 -591 108 -567
rect 261 -650 262 -590
rect 275 -591 276 -567
rect 355 -591 356 -567
rect 436 -591 437 -567
rect 471 -650 472 -590
rect 478 -591 479 -567
rect 513 -650 514 -590
rect 551 -591 552 -567
rect 856 -591 857 -567
rect 877 -591 878 -567
rect 961 -650 962 -590
rect 44 -593 45 -567
rect 464 -650 465 -592
rect 555 -593 556 -567
rect 569 -650 570 -592
rect 625 -650 626 -592
rect 681 -593 682 -567
rect 688 -593 689 -567
rect 744 -650 745 -592
rect 751 -650 752 -592
rect 758 -593 759 -567
rect 761 -650 762 -592
rect 1010 -593 1011 -567
rect 44 -650 45 -594
rect 93 -595 94 -567
rect 107 -650 108 -594
rect 117 -650 118 -594
rect 121 -650 122 -594
rect 201 -595 202 -567
rect 205 -595 206 -567
rect 397 -595 398 -567
rect 415 -595 416 -567
rect 436 -650 437 -594
rect 555 -650 556 -594
rect 639 -595 640 -567
rect 656 -650 657 -594
rect 1080 -595 1081 -567
rect 54 -650 55 -596
rect 800 -597 801 -567
rect 807 -597 808 -567
rect 877 -650 878 -596
rect 926 -597 927 -567
rect 968 -650 969 -596
rect 982 -597 983 -567
rect 1010 -650 1011 -596
rect 1017 -597 1018 -567
rect 1080 -650 1081 -596
rect 65 -599 66 -567
rect 506 -650 507 -598
rect 611 -599 612 -567
rect 639 -650 640 -598
rect 660 -599 661 -567
rect 1073 -599 1074 -567
rect 68 -650 69 -600
rect 457 -601 458 -567
rect 628 -601 629 -567
rect 730 -650 731 -600
rect 765 -601 766 -567
rect 856 -650 857 -600
rect 926 -650 927 -600
rect 947 -601 948 -567
rect 954 -601 955 -567
rect 1003 -650 1004 -600
rect 1045 -601 1046 -567
rect 1073 -650 1074 -600
rect 72 -650 73 -602
rect 373 -603 374 -567
rect 450 -603 451 -567
rect 457 -650 458 -602
rect 632 -603 633 -567
rect 681 -650 682 -602
rect 723 -603 724 -567
rect 807 -650 808 -602
rect 821 -603 822 -567
rect 842 -650 843 -602
rect 849 -603 850 -567
rect 954 -650 955 -602
rect 989 -603 990 -567
rect 1045 -650 1046 -602
rect 79 -650 80 -604
rect 835 -650 836 -604
rect 905 -605 906 -567
rect 947 -650 948 -604
rect 989 -650 990 -604
rect 1052 -605 1053 -567
rect 75 -607 76 -567
rect 905 -650 906 -606
rect 933 -607 934 -567
rect 982 -650 983 -606
rect 996 -607 997 -567
rect 1052 -650 1053 -606
rect 93 -650 94 -608
rect 607 -609 608 -567
rect 611 -650 612 -608
rect 632 -650 633 -608
rect 646 -609 647 -567
rect 660 -650 661 -608
rect 765 -650 766 -608
rect 779 -609 780 -567
rect 793 -609 794 -567
rect 884 -650 885 -608
rect 940 -609 941 -567
rect 1017 -650 1018 -608
rect 114 -611 115 -567
rect 450 -650 451 -610
rect 485 -611 486 -567
rect 646 -650 647 -610
rect 674 -611 675 -567
rect 779 -650 780 -610
rect 800 -650 801 -610
rect 1094 -611 1095 -567
rect 128 -613 129 -567
rect 446 -650 447 -612
rect 537 -613 538 -567
rect 723 -650 724 -612
rect 772 -613 773 -567
rect 821 -650 822 -612
rect 863 -613 864 -567
rect 996 -650 997 -612
rect 1031 -613 1032 -567
rect 1094 -650 1095 -612
rect 149 -650 150 -614
rect 408 -650 409 -614
rect 663 -615 664 -567
rect 1031 -650 1032 -614
rect 152 -617 153 -567
rect 296 -650 297 -616
rect 331 -617 332 -567
rect 352 -650 353 -616
rect 373 -650 374 -616
rect 481 -650 482 -616
rect 667 -617 668 -567
rect 674 -650 675 -616
rect 695 -617 696 -567
rect 793 -650 794 -616
rect 814 -617 815 -567
rect 849 -650 850 -616
rect 166 -619 167 -567
rect 912 -619 913 -567
rect 170 -621 171 -567
rect 198 -650 199 -620
rect 212 -621 213 -567
rect 366 -621 367 -567
rect 390 -621 391 -567
rect 863 -650 864 -620
rect 891 -621 892 -567
rect 912 -650 913 -620
rect 51 -623 52 -567
rect 366 -650 367 -622
rect 583 -623 584 -567
rect 667 -650 668 -622
rect 695 -650 696 -622
rect 758 -650 759 -622
rect 828 -623 829 -567
rect 891 -650 892 -622
rect 170 -650 171 -624
rect 247 -625 248 -567
rect 289 -625 290 -567
rect 485 -650 486 -624
rect 583 -650 584 -624
rect 618 -625 619 -567
rect 716 -625 717 -567
rect 772 -650 773 -624
rect 786 -625 787 -567
rect 828 -650 829 -624
rect 177 -627 178 -567
rect 226 -650 227 -626
rect 233 -627 234 -567
rect 254 -650 255 -626
rect 289 -650 290 -626
rect 607 -650 608 -626
rect 653 -627 654 -567
rect 716 -650 717 -626
rect 737 -627 738 -567
rect 814 -650 815 -626
rect 100 -650 101 -628
rect 737 -650 738 -628
rect 177 -650 178 -630
rect 184 -631 185 -567
rect 212 -650 213 -630
rect 317 -631 318 -567
rect 341 -650 342 -630
rect 940 -650 941 -630
rect 142 -633 143 -567
rect 317 -650 318 -632
rect 345 -633 346 -567
rect 394 -650 395 -632
rect 422 -633 423 -567
rect 653 -650 654 -632
rect 58 -635 59 -567
rect 345 -650 346 -634
rect 348 -650 349 -634
rect 492 -650 493 -634
rect 576 -635 577 -567
rect 618 -650 619 -634
rect 58 -650 59 -636
rect 240 -637 241 -567
rect 247 -650 248 -636
rect 282 -637 283 -567
rect 359 -637 360 -567
rect 786 -650 787 -636
rect 135 -639 136 -567
rect 240 -650 241 -638
rect 282 -650 283 -638
rect 320 -639 321 -567
rect 359 -650 360 -638
rect 401 -639 402 -567
rect 422 -650 423 -638
rect 614 -650 615 -638
rect 135 -650 136 -640
rect 163 -641 164 -567
rect 184 -650 185 -640
rect 268 -650 269 -640
rect 401 -650 402 -640
rect 429 -641 430 -567
rect 527 -641 528 -567
rect 576 -650 577 -640
rect 142 -650 143 -642
rect 590 -643 591 -567
rect 163 -650 164 -644
rect 205 -650 206 -644
rect 219 -645 220 -567
rect 275 -650 276 -644
rect 324 -645 325 -567
rect 429 -650 430 -644
rect 499 -645 500 -567
rect 527 -650 528 -644
rect 156 -647 157 -567
rect 219 -650 220 -646
rect 310 -647 311 -567
rect 324 -650 325 -646
rect 520 -647 521 -567
rect 590 -650 591 -646
rect 310 -650 311 -648
rect 331 -650 332 -648
rect 9 -660 10 -658
rect 9 -731 10 -659
rect 9 -660 10 -658
rect 9 -731 10 -659
rect 16 -660 17 -658
rect 128 -731 129 -659
rect 149 -660 150 -658
rect 233 -660 234 -658
rect 254 -660 255 -658
rect 415 -731 416 -659
rect 425 -731 426 -659
rect 607 -660 608 -658
rect 611 -731 612 -659
rect 632 -660 633 -658
rect 691 -660 692 -658
rect 975 -660 976 -658
rect 1003 -660 1004 -658
rect 1006 -660 1007 -658
rect 1038 -660 1039 -658
rect 1041 -660 1042 -658
rect 1059 -660 1060 -658
rect 1150 -731 1151 -659
rect 1178 -660 1179 -658
rect 1185 -731 1186 -659
rect 16 -731 17 -661
rect 184 -662 185 -658
rect 187 -662 188 -658
rect 236 -662 237 -658
rect 254 -731 255 -661
rect 268 -662 269 -658
rect 324 -662 325 -658
rect 338 -662 339 -658
rect 387 -662 388 -658
rect 387 -731 388 -661
rect 387 -662 388 -658
rect 387 -731 388 -661
rect 408 -662 409 -658
rect 793 -662 794 -658
rect 807 -662 808 -658
rect 810 -708 811 -661
rect 849 -662 850 -658
rect 849 -731 850 -661
rect 849 -662 850 -658
rect 849 -731 850 -661
rect 933 -662 934 -658
rect 1017 -662 1018 -658
rect 1038 -731 1039 -661
rect 1115 -662 1116 -658
rect 23 -731 24 -663
rect 422 -664 423 -658
rect 439 -731 440 -663
rect 635 -731 636 -663
rect 737 -664 738 -658
rect 737 -731 738 -663
rect 737 -664 738 -658
rect 737 -731 738 -663
rect 747 -731 748 -663
rect 779 -664 780 -658
rect 807 -731 808 -663
rect 814 -664 815 -658
rect 933 -731 934 -663
rect 947 -664 948 -658
rect 975 -731 976 -663
rect 1024 -664 1025 -658
rect 1045 -664 1046 -658
rect 1059 -731 1060 -663
rect 1066 -664 1067 -658
rect 1066 -731 1067 -663
rect 1066 -664 1067 -658
rect 1066 -731 1067 -663
rect 1087 -664 1088 -658
rect 1115 -731 1116 -663
rect 30 -666 31 -658
rect 478 -666 479 -658
rect 481 -666 482 -658
rect 919 -666 920 -658
rect 947 -731 948 -665
rect 982 -666 983 -658
rect 996 -666 997 -658
rect 1017 -731 1018 -665
rect 1087 -731 1088 -665
rect 1129 -666 1130 -658
rect 37 -668 38 -658
rect 131 -668 132 -658
rect 142 -668 143 -658
rect 338 -731 339 -667
rect 345 -668 346 -658
rect 478 -731 479 -667
rect 513 -668 514 -658
rect 660 -668 661 -658
rect 695 -668 696 -658
rect 779 -731 780 -667
rect 814 -731 815 -667
rect 898 -668 899 -658
rect 919 -731 920 -667
rect 968 -668 969 -658
rect 996 -731 997 -667
rect 1003 -731 1004 -667
rect 1052 -668 1053 -658
rect 1090 -731 1091 -667
rect 1171 -731 1172 -667
rect 37 -731 38 -669
rect 121 -670 122 -658
rect 142 -731 143 -669
rect 191 -670 192 -658
rect 205 -670 206 -658
rect 397 -731 398 -669
rect 443 -670 444 -658
rect 1024 -731 1025 -669
rect 1031 -670 1032 -658
rect 1052 -731 1053 -669
rect 1101 -670 1102 -658
rect 1129 -731 1130 -669
rect 44 -672 45 -658
rect 117 -672 118 -658
rect 159 -672 160 -658
rect 597 -672 598 -658
rect 604 -672 605 -658
rect 989 -672 990 -658
rect 1010 -672 1011 -658
rect 1045 -731 1046 -671
rect 1080 -672 1081 -658
rect 1101 -731 1102 -671
rect 1108 -672 1109 -658
rect 1143 -731 1144 -671
rect 44 -731 45 -673
rect 198 -674 199 -658
rect 208 -731 209 -673
rect 212 -674 213 -658
rect 226 -674 227 -658
rect 226 -731 227 -673
rect 226 -674 227 -658
rect 226 -731 227 -673
rect 233 -731 234 -673
rect 261 -674 262 -658
rect 268 -731 269 -673
rect 691 -731 692 -673
rect 758 -731 759 -673
rect 772 -674 773 -658
rect 842 -674 843 -658
rect 898 -731 899 -673
rect 940 -674 941 -658
rect 968 -731 969 -673
rect 1073 -674 1074 -658
rect 1080 -731 1081 -673
rect 1108 -731 1109 -673
rect 1136 -674 1137 -658
rect 51 -731 52 -675
rect 191 -731 192 -675
rect 198 -731 199 -675
rect 303 -676 304 -658
rect 324 -731 325 -675
rect 373 -676 374 -658
rect 380 -676 381 -658
rect 513 -731 514 -675
rect 523 -676 524 -658
rect 1164 -731 1165 -675
rect 54 -678 55 -658
rect 65 -678 66 -658
rect 72 -678 73 -658
rect 446 -678 447 -658
rect 457 -678 458 -658
rect 457 -731 458 -677
rect 457 -678 458 -658
rect 457 -731 458 -677
rect 464 -678 465 -658
rect 474 -731 475 -677
rect 502 -678 503 -658
rect 842 -731 843 -677
rect 940 -731 941 -677
rect 954 -678 955 -658
rect 961 -678 962 -658
rect 989 -731 990 -677
rect 1073 -731 1074 -677
rect 1094 -678 1095 -658
rect 1122 -678 1123 -658
rect 1136 -731 1137 -677
rect 58 -680 59 -658
rect 261 -731 262 -679
rect 303 -731 304 -679
rect 450 -680 451 -658
rect 464 -731 465 -679
rect 709 -680 710 -658
rect 905 -680 906 -658
rect 954 -731 955 -679
rect 58 -731 59 -681
rect 352 -682 353 -658
rect 366 -682 367 -658
rect 443 -731 444 -681
rect 450 -731 451 -681
rect 471 -682 472 -658
rect 516 -682 517 -658
rect 1122 -731 1123 -681
rect 65 -731 66 -683
rect 523 -731 524 -683
rect 551 -684 552 -658
rect 856 -684 857 -658
rect 884 -684 885 -658
rect 905 -731 906 -683
rect 912 -684 913 -658
rect 961 -731 962 -683
rect 72 -731 73 -685
rect 212 -731 213 -685
rect 317 -686 318 -658
rect 352 -731 353 -685
rect 366 -731 367 -685
rect 520 -686 521 -658
rect 551 -731 552 -685
rect 583 -686 584 -658
rect 597 -731 598 -685
rect 835 -686 836 -658
rect 891 -686 892 -658
rect 912 -731 913 -685
rect 79 -688 80 -658
rect 96 -708 97 -687
rect 100 -731 101 -687
rect 219 -688 220 -658
rect 310 -688 311 -658
rect 317 -731 318 -687
rect 345 -731 346 -687
rect 436 -688 437 -658
rect 499 -688 500 -658
rect 884 -731 885 -687
rect 79 -731 80 -689
rect 107 -690 108 -658
rect 114 -731 115 -689
rect 135 -690 136 -658
rect 152 -731 153 -689
rect 373 -731 374 -689
rect 380 -731 381 -689
rect 418 -690 419 -658
rect 485 -690 486 -658
rect 499 -731 500 -689
rect 569 -690 570 -658
rect 583 -731 584 -689
rect 604 -731 605 -689
rect 863 -690 864 -658
rect 870 -690 871 -658
rect 891 -731 892 -689
rect 82 -692 83 -658
rect 548 -731 549 -691
rect 576 -692 577 -658
rect 653 -731 654 -691
rect 660 -731 661 -691
rect 716 -692 717 -658
rect 765 -692 766 -658
rect 863 -731 864 -691
rect 86 -731 87 -693
rect 149 -731 150 -693
rect 156 -694 157 -658
rect 1010 -731 1011 -693
rect 89 -696 90 -658
rect 205 -731 206 -695
rect 219 -731 220 -695
rect 275 -696 276 -658
rect 506 -696 507 -658
rect 576 -731 577 -695
rect 614 -696 615 -658
rect 926 -696 927 -658
rect 93 -698 94 -658
rect 107 -731 108 -697
rect 135 -731 136 -697
rect 835 -731 836 -697
rect 93 -731 94 -699
rect 163 -700 164 -658
rect 177 -700 178 -658
rect 177 -731 178 -699
rect 177 -700 178 -658
rect 177 -731 178 -699
rect 184 -731 185 -699
rect 331 -731 332 -699
rect 506 -731 507 -699
rect 800 -700 801 -658
rect 821 -700 822 -658
rect 856 -731 857 -699
rect 103 -702 104 -658
rect 555 -702 556 -658
rect 646 -702 647 -658
rect 709 -731 710 -701
rect 716 -731 717 -701
rect 793 -731 794 -701
rect 800 -731 801 -701
rect 828 -702 829 -658
rect 156 -731 157 -703
rect 170 -704 171 -658
rect 240 -704 241 -658
rect 485 -731 486 -703
rect 534 -704 535 -658
rect 569 -731 570 -703
rect 646 -731 647 -703
rect 681 -704 682 -658
rect 688 -704 689 -658
rect 695 -731 696 -703
rect 702 -704 703 -658
rect 772 -731 773 -703
rect 163 -731 164 -705
rect 275 -731 276 -705
rect 282 -706 283 -658
rect 467 -731 468 -705
rect 821 -731 822 -705
rect 170 -731 171 -707
rect 359 -708 360 -658
rect 527 -708 528 -658
rect 534 -731 535 -707
rect 541 -708 542 -658
rect 555 -731 556 -707
rect 667 -708 668 -658
rect 681 -731 682 -707
rect 688 -731 689 -707
rect 982 -731 983 -707
rect 1041 -731 1042 -707
rect 1094 -731 1095 -707
rect 240 -731 241 -709
rect 296 -710 297 -658
rect 429 -710 430 -658
rect 541 -731 542 -709
rect 639 -710 640 -658
rect 667 -731 668 -709
rect 730 -710 731 -658
rect 926 -731 927 -709
rect 282 -731 283 -711
rect 394 -712 395 -658
rect 401 -712 402 -658
rect 429 -731 430 -711
rect 527 -731 528 -711
rect 618 -712 619 -658
rect 639 -731 640 -711
rect 702 -731 703 -711
rect 730 -731 731 -711
rect 786 -712 787 -658
rect 33 -731 34 -713
rect 394 -731 395 -713
rect 411 -731 412 -713
rect 786 -731 787 -713
rect 289 -716 290 -658
rect 296 -731 297 -715
rect 562 -716 563 -658
rect 618 -731 619 -715
rect 744 -716 745 -658
rect 765 -731 766 -715
rect 289 -731 290 -717
rect 492 -718 493 -658
rect 562 -731 563 -717
rect 590 -718 591 -658
rect 744 -731 745 -717
rect 870 -731 871 -717
rect 341 -731 342 -719
rect 590 -731 591 -719
rect 751 -720 752 -658
rect 828 -731 829 -719
rect 492 -731 493 -721
rect 723 -722 724 -658
rect 625 -724 626 -658
rect 751 -731 752 -723
rect 625 -731 626 -725
rect 1111 -731 1112 -725
rect 674 -728 675 -658
rect 723 -731 724 -727
rect 656 -730 657 -658
rect 674 -731 675 -729
rect 9 -741 10 -739
rect 138 -741 139 -739
rect 142 -741 143 -739
rect 142 -820 143 -740
rect 142 -741 143 -739
rect 142 -820 143 -740
rect 149 -820 150 -740
rect 583 -741 584 -739
rect 600 -741 601 -739
rect 940 -741 941 -739
rect 1038 -741 1039 -739
rect 1087 -741 1088 -739
rect 1108 -741 1109 -739
rect 1136 -741 1137 -739
rect 1143 -741 1144 -739
rect 1192 -820 1193 -740
rect 9 -820 10 -742
rect 79 -743 80 -739
rect 86 -743 87 -739
rect 131 -820 132 -742
rect 163 -743 164 -739
rect 362 -743 363 -739
rect 373 -743 374 -739
rect 383 -820 384 -742
rect 404 -743 405 -739
rect 499 -743 500 -739
rect 502 -820 503 -742
rect 527 -743 528 -739
rect 583 -820 584 -742
rect 747 -743 748 -739
rect 765 -743 766 -739
rect 765 -820 766 -742
rect 765 -743 766 -739
rect 765 -820 766 -742
rect 782 -820 783 -742
rect 1003 -743 1004 -739
rect 1031 -743 1032 -739
rect 1038 -820 1039 -742
rect 1045 -743 1046 -739
rect 1045 -820 1046 -742
rect 1045 -743 1046 -739
rect 1045 -820 1046 -742
rect 1052 -743 1053 -739
rect 1108 -820 1109 -742
rect 1122 -743 1123 -739
rect 1178 -820 1179 -742
rect 1185 -743 1186 -739
rect 1213 -820 1214 -742
rect 16 -745 17 -739
rect 338 -745 339 -739
rect 359 -745 360 -739
rect 1052 -820 1053 -744
rect 1059 -745 1060 -739
rect 1122 -820 1123 -744
rect 1129 -745 1130 -739
rect 1185 -820 1186 -744
rect 16 -820 17 -746
rect 366 -747 367 -739
rect 373 -820 374 -746
rect 387 -747 388 -739
rect 408 -820 409 -746
rect 625 -747 626 -739
rect 639 -820 640 -746
rect 817 -820 818 -746
rect 821 -747 822 -739
rect 852 -820 853 -746
rect 884 -747 885 -739
rect 1003 -820 1004 -746
rect 1059 -820 1060 -746
rect 1090 -747 1091 -739
rect 1101 -747 1102 -739
rect 1143 -820 1144 -746
rect 1150 -747 1151 -739
rect 1160 -747 1161 -739
rect 1164 -747 1165 -739
rect 1199 -820 1200 -746
rect 23 -749 24 -739
rect 401 -820 402 -748
rect 411 -749 412 -739
rect 415 -749 416 -739
rect 439 -749 440 -739
rect 471 -820 472 -748
rect 495 -820 496 -748
rect 947 -749 948 -739
rect 968 -749 969 -739
rect 1031 -820 1032 -748
rect 1080 -749 1081 -739
rect 1136 -820 1137 -748
rect 1171 -749 1172 -739
rect 1220 -820 1221 -748
rect 23 -820 24 -750
rect 345 -751 346 -739
rect 387 -820 388 -750
rect 569 -751 570 -739
rect 572 -820 573 -750
rect 1164 -820 1165 -750
rect 30 -820 31 -752
rect 170 -753 171 -739
rect 173 -820 174 -752
rect 205 -820 206 -752
rect 212 -753 213 -739
rect 425 -753 426 -739
rect 464 -820 465 -752
rect 478 -753 479 -739
rect 513 -753 514 -739
rect 635 -753 636 -739
rect 642 -753 643 -739
rect 863 -753 864 -739
rect 926 -753 927 -739
rect 940 -820 941 -752
rect 947 -820 948 -752
rect 954 -753 955 -739
rect 989 -753 990 -739
rect 1080 -820 1081 -752
rect 1115 -753 1116 -739
rect 1150 -820 1151 -752
rect 37 -755 38 -739
rect 124 -755 125 -739
rect 177 -755 178 -739
rect 184 -820 185 -754
rect 187 -755 188 -739
rect 541 -755 542 -739
rect 625 -820 626 -754
rect 877 -755 878 -739
rect 954 -820 955 -754
rect 1157 -755 1158 -739
rect 37 -820 38 -756
rect 117 -820 118 -756
rect 156 -757 157 -739
rect 177 -820 178 -756
rect 191 -757 192 -739
rect 254 -757 255 -739
rect 324 -757 325 -739
rect 324 -820 325 -756
rect 324 -757 325 -739
rect 324 -820 325 -756
rect 331 -757 332 -739
rect 436 -820 437 -756
rect 485 -757 486 -739
rect 513 -820 514 -756
rect 520 -757 521 -739
rect 968 -820 969 -756
rect 982 -757 983 -739
rect 989 -820 990 -756
rect 996 -757 997 -739
rect 1087 -820 1088 -756
rect 58 -759 59 -739
rect 345 -820 346 -758
rect 366 -820 367 -758
rect 520 -820 521 -758
rect 523 -759 524 -739
rect 660 -759 661 -739
rect 663 -820 664 -758
rect 1129 -820 1130 -758
rect 58 -820 59 -760
rect 93 -761 94 -739
rect 100 -761 101 -739
rect 212 -820 213 -760
rect 338 -820 339 -760
rect 597 -761 598 -739
rect 604 -761 605 -739
rect 1157 -820 1158 -760
rect 65 -763 66 -739
rect 331 -820 332 -762
rect 380 -763 381 -739
rect 660 -820 661 -762
rect 688 -763 689 -739
rect 898 -763 899 -739
rect 933 -763 934 -739
rect 982 -820 983 -762
rect 996 -820 997 -762
rect 1024 -763 1025 -739
rect 1073 -763 1074 -739
rect 1171 -820 1172 -762
rect 44 -765 45 -739
rect 380 -820 381 -764
rect 394 -765 395 -739
rect 884 -820 885 -764
rect 1010 -765 1011 -739
rect 1115 -820 1116 -764
rect 44 -820 45 -766
rect 268 -767 269 -739
rect 341 -767 342 -739
rect 1024 -820 1025 -766
rect 1073 -820 1074 -766
rect 1094 -767 1095 -739
rect 65 -820 66 -768
rect 506 -769 507 -739
rect 527 -820 528 -768
rect 534 -769 535 -739
rect 541 -820 542 -768
rect 555 -769 556 -739
rect 565 -820 566 -768
rect 933 -820 934 -768
rect 1017 -769 1018 -739
rect 1094 -820 1095 -768
rect 79 -820 80 -770
rect 425 -820 426 -770
rect 499 -820 500 -770
rect 534 -820 535 -770
rect 569 -820 570 -770
rect 1010 -820 1011 -770
rect 1017 -820 1018 -770
rect 1066 -771 1067 -739
rect 86 -820 87 -772
rect 317 -773 318 -739
rect 394 -820 395 -772
rect 429 -773 430 -739
rect 506 -820 507 -772
rect 576 -773 577 -739
rect 590 -773 591 -739
rect 604 -820 605 -772
rect 688 -820 689 -772
rect 695 -773 696 -739
rect 698 -820 699 -772
rect 1101 -820 1102 -772
rect 93 -820 94 -774
rect 240 -775 241 -739
rect 268 -820 269 -774
rect 310 -775 311 -739
rect 317 -820 318 -774
rect 352 -775 353 -739
rect 415 -820 416 -774
rect 642 -820 643 -774
rect 702 -775 703 -739
rect 702 -820 703 -774
rect 702 -775 703 -739
rect 702 -820 703 -774
rect 716 -775 717 -739
rect 856 -775 857 -739
rect 870 -775 871 -739
rect 877 -820 878 -774
rect 100 -820 101 -776
rect 135 -777 136 -739
rect 138 -820 139 -776
rect 156 -820 157 -776
rect 163 -820 164 -776
rect 254 -820 255 -776
rect 429 -820 430 -776
rect 891 -777 892 -739
rect 114 -779 115 -739
rect 121 -820 122 -778
rect 135 -820 136 -778
rect 289 -779 290 -739
rect 457 -779 458 -739
rect 576 -820 577 -778
rect 590 -820 591 -778
rect 618 -779 619 -739
rect 737 -779 738 -739
rect 737 -820 738 -778
rect 737 -779 738 -739
rect 737 -820 738 -778
rect 744 -779 745 -739
rect 975 -779 976 -739
rect 170 -820 171 -780
rect 240 -820 241 -780
rect 247 -781 248 -739
rect 310 -820 311 -780
rect 443 -781 444 -739
rect 457 -820 458 -780
rect 485 -820 486 -780
rect 695 -820 696 -780
rect 786 -781 787 -739
rect 898 -820 899 -780
rect 191 -820 192 -782
rect 296 -783 297 -739
rect 443 -820 444 -782
rect 450 -783 451 -739
rect 492 -783 493 -739
rect 716 -820 717 -782
rect 786 -820 787 -782
rect 807 -783 808 -739
rect 842 -783 843 -739
rect 926 -820 927 -782
rect 226 -785 227 -739
rect 247 -820 248 -784
rect 289 -820 290 -784
rect 352 -820 353 -784
rect 548 -785 549 -739
rect 744 -820 745 -784
rect 779 -785 780 -739
rect 807 -820 808 -784
rect 835 -785 836 -739
rect 842 -820 843 -784
rect 849 -785 850 -739
rect 863 -820 864 -784
rect 891 -820 892 -784
rect 905 -785 906 -739
rect 128 -787 129 -739
rect 226 -820 227 -786
rect 296 -820 297 -786
rect 611 -787 612 -739
rect 656 -820 657 -786
rect 975 -820 976 -786
rect 303 -789 304 -739
rect 450 -820 451 -788
rect 548 -820 549 -788
rect 562 -789 563 -739
rect 597 -820 598 -788
rect 751 -789 752 -739
rect 779 -820 780 -788
rect 870 -820 871 -788
rect 198 -791 199 -739
rect 303 -820 304 -790
rect 555 -820 556 -790
rect 1066 -820 1067 -790
rect 107 -793 108 -739
rect 198 -820 199 -792
rect 562 -820 563 -792
rect 730 -793 731 -739
rect 751 -820 752 -792
rect 828 -793 829 -739
rect 849 -820 850 -792
rect 1206 -820 1207 -792
rect 107 -820 108 -794
rect 219 -795 220 -739
rect 474 -795 475 -739
rect 828 -820 829 -794
rect 856 -820 857 -794
rect 919 -795 920 -739
rect 219 -820 220 -796
rect 653 -797 654 -739
rect 793 -797 794 -739
rect 821 -820 822 -796
rect 912 -797 913 -739
rect 919 -820 920 -796
rect 611 -820 612 -798
rect 667 -799 668 -739
rect 772 -799 773 -739
rect 793 -820 794 -798
rect 800 -799 801 -739
rect 905 -820 906 -798
rect 912 -820 913 -798
rect 961 -799 962 -739
rect 478 -820 479 -800
rect 772 -820 773 -800
rect 814 -801 815 -739
rect 835 -820 836 -800
rect 632 -803 633 -739
rect 961 -820 962 -802
rect 632 -820 633 -804
rect 681 -805 682 -739
rect 758 -805 759 -739
rect 800 -820 801 -804
rect 51 -807 52 -739
rect 681 -820 682 -806
rect 51 -820 52 -808
rect 282 -809 283 -739
rect 621 -820 622 -808
rect 758 -820 759 -808
rect 233 -811 234 -739
rect 282 -820 283 -810
rect 667 -820 668 -810
rect 709 -811 710 -739
rect 233 -820 234 -812
rect 275 -813 276 -739
rect 646 -813 647 -739
rect 709 -820 710 -812
rect 261 -815 262 -739
rect 275 -820 276 -814
rect 646 -820 647 -814
rect 674 -815 675 -739
rect 674 -820 675 -816
rect 723 -817 724 -739
rect 723 -820 724 -818
rect 730 -820 731 -818
rect 19 -907 20 -829
rect 313 -907 314 -829
rect 355 -830 356 -828
rect 1003 -830 1004 -828
rect 30 -832 31 -828
rect 117 -832 118 -828
rect 121 -832 122 -828
rect 1101 -832 1102 -828
rect 33 -907 34 -833
rect 170 -907 171 -833
rect 184 -834 185 -828
rect 184 -907 185 -833
rect 184 -834 185 -828
rect 184 -907 185 -833
rect 198 -834 199 -828
rect 499 -907 500 -833
rect 523 -834 524 -828
rect 590 -834 591 -828
rect 618 -834 619 -828
rect 905 -834 906 -828
rect 947 -834 948 -828
rect 947 -907 948 -833
rect 947 -834 948 -828
rect 947 -907 948 -833
rect 975 -834 976 -828
rect 975 -907 976 -833
rect 975 -834 976 -828
rect 975 -907 976 -833
rect 996 -834 997 -828
rect 999 -834 1000 -828
rect 1003 -907 1004 -833
rect 1038 -834 1039 -828
rect 44 -836 45 -828
rect 569 -836 570 -828
rect 590 -907 591 -835
rect 632 -836 633 -828
rect 639 -907 640 -835
rect 702 -836 703 -828
rect 726 -836 727 -828
rect 1066 -836 1067 -828
rect 44 -907 45 -837
rect 289 -838 290 -828
rect 303 -838 304 -828
rect 303 -907 304 -837
rect 303 -838 304 -828
rect 303 -907 304 -837
rect 359 -907 360 -837
rect 383 -838 384 -828
rect 387 -838 388 -828
rect 478 -907 479 -837
rect 485 -838 486 -828
rect 520 -907 521 -837
rect 541 -838 542 -828
rect 541 -907 542 -837
rect 541 -838 542 -828
rect 541 -907 542 -837
rect 555 -838 556 -828
rect 611 -838 612 -828
rect 656 -838 657 -828
rect 730 -838 731 -828
rect 758 -838 759 -828
rect 849 -907 850 -837
rect 905 -907 906 -837
rect 989 -838 990 -828
rect 996 -907 997 -837
rect 1010 -838 1011 -828
rect 1017 -838 1018 -828
rect 1066 -907 1067 -837
rect 37 -840 38 -828
rect 387 -907 388 -839
rect 394 -840 395 -828
rect 495 -840 496 -828
rect 558 -840 559 -828
rect 632 -907 633 -839
rect 656 -907 657 -839
rect 1080 -840 1081 -828
rect 51 -842 52 -828
rect 264 -907 265 -841
rect 296 -842 297 -828
rect 555 -907 556 -841
rect 562 -907 563 -841
rect 604 -842 605 -828
rect 611 -907 612 -841
rect 1094 -842 1095 -828
rect 51 -907 52 -843
rect 191 -844 192 -828
rect 198 -907 199 -843
rect 233 -844 234 -828
rect 296 -907 297 -843
rect 324 -844 325 -828
rect 362 -844 363 -828
rect 457 -844 458 -828
rect 464 -844 465 -828
rect 621 -844 622 -828
rect 660 -907 661 -843
rect 667 -844 668 -828
rect 695 -844 696 -828
rect 1087 -844 1088 -828
rect 1094 -907 1095 -843
rect 1178 -844 1179 -828
rect 16 -846 17 -828
rect 191 -907 192 -845
rect 205 -846 206 -828
rect 604 -907 605 -845
rect 621 -907 622 -845
rect 765 -846 766 -828
rect 779 -907 780 -845
rect 828 -846 829 -828
rect 968 -846 969 -828
rect 1038 -907 1039 -845
rect 1073 -846 1074 -828
rect 1087 -907 1088 -845
rect 1178 -907 1179 -845
rect 1220 -846 1221 -828
rect 58 -848 59 -828
rect 61 -860 62 -847
rect 72 -848 73 -828
rect 72 -907 73 -847
rect 72 -848 73 -828
rect 72 -907 73 -847
rect 86 -848 87 -828
rect 352 -848 353 -828
rect 380 -848 381 -828
rect 1101 -907 1102 -847
rect 58 -907 59 -849
rect 240 -850 241 -828
rect 289 -907 290 -849
rect 828 -907 829 -849
rect 968 -907 969 -849
rect 982 -850 983 -828
rect 989 -907 990 -849
rect 1129 -850 1130 -828
rect 86 -907 87 -851
rect 681 -852 682 -828
rect 695 -907 696 -851
rect 716 -852 717 -828
rect 730 -907 731 -851
rect 800 -852 801 -828
rect 814 -852 815 -828
rect 1192 -852 1193 -828
rect 5 -907 6 -853
rect 814 -907 815 -853
rect 982 -907 983 -853
rect 1115 -854 1116 -828
rect 1129 -907 1130 -853
rect 1185 -854 1186 -828
rect 1192 -907 1193 -853
rect 1213 -854 1214 -828
rect 93 -856 94 -828
rect 240 -907 241 -855
rect 292 -907 293 -855
rect 800 -907 801 -855
rect 1017 -907 1018 -855
rect 1059 -856 1060 -828
rect 1073 -907 1074 -855
rect 1136 -856 1137 -828
rect 93 -907 94 -857
rect 114 -858 115 -828
rect 1031 -858 1032 -828
rect 1059 -907 1060 -857
rect 1122 -858 1123 -828
rect 117 -907 118 -859
rect 380 -907 381 -859
rect 401 -860 402 -828
rect 401 -907 402 -859
rect 401 -860 402 -828
rect 401 -907 402 -859
rect 422 -860 423 -828
rect 506 -860 507 -828
rect 569 -907 570 -859
rect 583 -860 584 -828
rect 663 -860 664 -828
rect 667 -907 668 -859
rect 681 -907 682 -859
rect 884 -860 885 -828
rect 999 -907 1000 -859
rect 1010 -907 1011 -859
rect 1024 -860 1025 -828
rect 1115 -907 1116 -859
rect 1122 -907 1123 -859
rect 1171 -860 1172 -828
rect 121 -907 122 -861
rect 614 -907 615 -861
rect 698 -862 699 -828
rect 1164 -862 1165 -828
rect 1171 -907 1172 -861
rect 1206 -862 1207 -828
rect 124 -864 125 -828
rect 226 -864 227 -828
rect 324 -907 325 -863
rect 331 -864 332 -828
rect 352 -907 353 -863
rect 436 -864 437 -828
rect 450 -864 451 -828
rect 457 -907 458 -863
rect 464 -907 465 -863
rect 502 -864 503 -828
rect 506 -907 507 -863
rect 576 -864 577 -828
rect 583 -907 584 -863
rect 688 -864 689 -828
rect 702 -907 703 -863
rect 744 -864 745 -828
rect 751 -864 752 -828
rect 765 -907 766 -863
rect 786 -864 787 -828
rect 786 -907 787 -863
rect 786 -864 787 -828
rect 786 -907 787 -863
rect 863 -864 864 -828
rect 884 -907 885 -863
rect 1024 -907 1025 -863
rect 1108 -864 1109 -828
rect 1164 -907 1165 -863
rect 1199 -864 1200 -828
rect 135 -907 136 -865
rect 345 -866 346 -828
rect 425 -866 426 -828
rect 625 -907 626 -865
rect 674 -866 675 -828
rect 688 -907 689 -865
rect 716 -907 717 -865
rect 772 -866 773 -828
rect 863 -907 864 -865
rect 891 -866 892 -828
rect 1031 -907 1032 -865
rect 1045 -866 1046 -828
rect 1080 -907 1081 -865
rect 1150 -866 1151 -828
rect 23 -868 24 -828
rect 425 -907 426 -867
rect 429 -868 430 -828
rect 744 -907 745 -867
rect 751 -907 752 -867
rect 793 -868 794 -828
rect 856 -868 857 -828
rect 891 -907 892 -867
rect 1045 -907 1046 -867
rect 1143 -868 1144 -828
rect 23 -907 24 -869
rect 219 -870 220 -828
rect 226 -907 227 -869
rect 278 -907 279 -869
rect 317 -870 318 -828
rect 331 -907 332 -869
rect 429 -907 430 -869
rect 443 -870 444 -828
rect 471 -870 472 -828
rect 723 -907 724 -869
rect 758 -907 759 -869
rect 807 -870 808 -828
rect 835 -870 836 -828
rect 856 -907 857 -869
rect 870 -870 871 -828
rect 1108 -907 1109 -869
rect 107 -872 108 -828
rect 317 -907 318 -871
rect 436 -907 437 -871
rect 597 -872 598 -828
rect 600 -907 601 -871
rect 793 -907 794 -871
rect 807 -907 808 -871
rect 842 -872 843 -828
rect 870 -907 871 -871
rect 961 -872 962 -828
rect 65 -874 66 -828
rect 597 -907 598 -873
rect 674 -907 675 -873
rect 1052 -874 1053 -828
rect 65 -907 66 -875
rect 534 -876 535 -828
rect 576 -907 577 -875
rect 646 -876 647 -828
rect 677 -907 678 -875
rect 835 -907 836 -875
rect 842 -907 843 -875
rect 877 -876 878 -828
rect 898 -876 899 -828
rect 1052 -907 1053 -875
rect 79 -878 80 -828
rect 107 -907 108 -877
rect 149 -878 150 -828
rect 443 -907 444 -877
rect 471 -907 472 -877
rect 670 -907 671 -877
rect 772 -907 773 -877
rect 821 -878 822 -828
rect 877 -907 878 -877
rect 919 -878 920 -828
rect 37 -907 38 -879
rect 79 -907 80 -879
rect 163 -880 164 -828
rect 1157 -880 1158 -828
rect 156 -882 157 -828
rect 163 -907 164 -881
rect 177 -882 178 -828
rect 233 -907 234 -881
rect 485 -907 486 -881
rect 513 -882 514 -828
rect 534 -907 535 -881
rect 548 -882 549 -828
rect 646 -907 647 -881
rect 709 -882 710 -828
rect 817 -882 818 -828
rect 961 -907 962 -881
rect 142 -884 143 -828
rect 177 -907 178 -883
rect 205 -907 206 -883
rect 247 -884 248 -828
rect 415 -884 416 -828
rect 548 -907 549 -883
rect 709 -907 710 -883
rect 737 -884 738 -828
rect 128 -886 129 -828
rect 142 -907 143 -885
rect 149 -907 150 -885
rect 247 -907 248 -885
rect 348 -907 349 -885
rect 415 -907 416 -885
rect 513 -907 514 -885
rect 527 -886 528 -828
rect 544 -907 545 -885
rect 919 -907 920 -885
rect 9 -888 10 -828
rect 128 -907 129 -887
rect 156 -907 157 -887
rect 492 -888 493 -828
rect 527 -907 528 -887
rect 653 -907 654 -887
rect 737 -907 738 -887
rect 933 -888 934 -828
rect 9 -907 10 -889
rect 254 -890 255 -828
rect 366 -890 367 -828
rect 492 -907 493 -889
rect 933 -907 934 -889
rect 940 -890 941 -828
rect 212 -892 213 -828
rect 394 -907 395 -891
rect 926 -892 927 -828
rect 940 -907 941 -891
rect 212 -907 213 -893
rect 408 -894 409 -828
rect 926 -907 927 -893
rect 954 -894 955 -828
rect 219 -907 220 -895
rect 282 -896 283 -828
rect 366 -907 367 -895
rect 373 -896 374 -828
rect 912 -896 913 -828
rect 954 -907 955 -895
rect 40 -907 41 -897
rect 282 -907 283 -897
rect 912 -907 913 -897
rect 1090 -907 1091 -897
rect 254 -907 255 -899
rect 338 -900 339 -828
rect 268 -902 269 -828
rect 408 -907 409 -901
rect 268 -907 269 -903
rect 275 -904 276 -828
rect 310 -904 311 -828
rect 338 -907 339 -903
rect 310 -907 311 -905
rect 450 -907 451 -905
rect 2 -996 3 -916
rect 86 -917 87 -915
rect 96 -996 97 -916
rect 485 -917 486 -915
rect 502 -996 503 -916
rect 513 -917 514 -915
rect 548 -917 549 -915
rect 681 -996 682 -916
rect 684 -917 685 -915
rect 1115 -917 1116 -915
rect 1136 -996 1137 -916
rect 1178 -917 1179 -915
rect 19 -919 20 -915
rect 814 -919 815 -915
rect 824 -919 825 -915
rect 1087 -996 1088 -918
rect 1101 -919 1102 -915
rect 1115 -996 1116 -918
rect 1150 -996 1151 -918
rect 1164 -919 1165 -915
rect 30 -996 31 -920
rect 170 -921 171 -915
rect 205 -996 206 -920
rect 576 -921 577 -915
rect 597 -921 598 -915
rect 870 -921 871 -915
rect 898 -921 899 -915
rect 1122 -921 1123 -915
rect 1157 -996 1158 -920
rect 1171 -921 1172 -915
rect 33 -923 34 -915
rect 499 -923 500 -915
rect 506 -923 507 -915
rect 513 -996 514 -922
rect 548 -996 549 -922
rect 562 -923 563 -915
rect 597 -996 598 -922
rect 828 -923 829 -915
rect 1108 -923 1109 -915
rect 1171 -996 1172 -922
rect 37 -925 38 -915
rect 604 -925 605 -915
rect 618 -996 619 -924
rect 702 -925 703 -915
rect 716 -925 717 -915
rect 1143 -996 1144 -924
rect 1164 -996 1165 -924
rect 1192 -925 1193 -915
rect 40 -927 41 -915
rect 324 -927 325 -915
rect 338 -927 339 -915
rect 338 -996 339 -926
rect 338 -927 339 -915
rect 338 -996 339 -926
rect 345 -996 346 -926
rect 492 -927 493 -915
rect 499 -996 500 -926
rect 898 -996 899 -926
rect 1066 -927 1067 -915
rect 1108 -996 1109 -926
rect 1122 -996 1123 -926
rect 1129 -927 1130 -915
rect 1185 -996 1186 -926
rect 1192 -996 1193 -926
rect 9 -929 10 -915
rect 324 -996 325 -928
rect 348 -929 349 -915
rect 408 -929 409 -915
rect 415 -929 416 -915
rect 492 -996 493 -928
rect 555 -929 556 -915
rect 1101 -996 1102 -928
rect 40 -996 41 -930
rect 576 -996 577 -930
rect 628 -996 629 -930
rect 709 -931 710 -915
rect 716 -996 717 -930
rect 730 -931 731 -915
rect 737 -931 738 -915
rect 828 -996 829 -930
rect 1052 -931 1053 -915
rect 1129 -996 1130 -930
rect 44 -933 45 -915
rect 611 -996 612 -932
rect 656 -933 657 -915
rect 989 -933 990 -915
rect 1052 -996 1053 -932
rect 1080 -933 1081 -915
rect 44 -996 45 -934
rect 100 -935 101 -915
rect 117 -935 118 -915
rect 390 -996 391 -934
rect 394 -935 395 -915
rect 394 -996 395 -934
rect 394 -935 395 -915
rect 394 -996 395 -934
rect 401 -935 402 -915
rect 401 -996 402 -934
rect 401 -935 402 -915
rect 401 -996 402 -934
rect 408 -996 409 -934
rect 558 -935 559 -915
rect 562 -996 563 -934
rect 569 -935 570 -915
rect 667 -996 668 -934
rect 695 -935 696 -915
rect 702 -996 703 -934
rect 772 -935 773 -915
rect 975 -935 976 -915
rect 1080 -996 1081 -934
rect 51 -937 52 -915
rect 114 -937 115 -915
rect 142 -937 143 -915
rect 152 -937 153 -915
rect 163 -937 164 -915
rect 163 -996 164 -936
rect 163 -937 164 -915
rect 163 -996 164 -936
rect 170 -996 171 -936
rect 208 -937 209 -915
rect 219 -937 220 -915
rect 436 -937 437 -915
rect 439 -937 440 -915
rect 632 -937 633 -915
rect 674 -996 675 -936
rect 730 -996 731 -936
rect 737 -996 738 -936
rect 786 -937 787 -915
rect 975 -996 976 -936
rect 1017 -937 1018 -915
rect 51 -996 52 -938
rect 61 -996 62 -938
rect 65 -939 66 -915
rect 555 -996 556 -938
rect 632 -996 633 -938
rect 646 -939 647 -915
rect 695 -996 696 -938
rect 870 -996 871 -938
rect 989 -996 990 -938
rect 1031 -939 1032 -915
rect 58 -941 59 -915
rect 114 -996 115 -940
rect 142 -996 143 -940
rect 264 -941 265 -915
rect 268 -941 269 -915
rect 289 -941 290 -915
rect 303 -941 304 -915
rect 310 -996 311 -940
rect 331 -941 332 -915
rect 415 -996 416 -940
rect 439 -996 440 -940
rect 859 -996 860 -940
rect 996 -941 997 -915
rect 1031 -996 1032 -940
rect 58 -996 59 -942
rect 107 -943 108 -915
rect 149 -996 150 -942
rect 233 -943 234 -915
rect 247 -943 248 -915
rect 289 -996 290 -942
rect 303 -996 304 -942
rect 733 -996 734 -942
rect 772 -996 773 -942
rect 863 -943 864 -915
rect 961 -943 962 -915
rect 996 -996 997 -942
rect 1017 -996 1018 -942
rect 1073 -943 1074 -915
rect 72 -945 73 -915
rect 712 -996 713 -944
rect 786 -996 787 -944
rect 800 -945 801 -915
rect 961 -996 962 -944
rect 1010 -945 1011 -915
rect 1038 -945 1039 -915
rect 1073 -996 1074 -944
rect 79 -947 80 -915
rect 107 -996 108 -946
rect 191 -947 192 -915
rect 219 -996 220 -946
rect 226 -947 227 -915
rect 226 -996 227 -946
rect 226 -947 227 -915
rect 226 -996 227 -946
rect 233 -996 234 -946
rect 376 -996 377 -946
rect 380 -947 381 -915
rect 653 -947 654 -915
rect 709 -996 710 -946
rect 982 -947 983 -915
rect 1010 -996 1011 -946
rect 1094 -947 1095 -915
rect 79 -996 80 -948
rect 128 -949 129 -915
rect 156 -949 157 -915
rect 191 -996 192 -948
rect 212 -949 213 -915
rect 247 -996 248 -948
rect 261 -949 262 -915
rect 331 -996 332 -948
rect 362 -996 363 -948
rect 814 -996 815 -948
rect 982 -996 983 -948
rect 1090 -949 1091 -915
rect 86 -996 87 -950
rect 93 -951 94 -915
rect 121 -951 122 -915
rect 128 -996 129 -950
rect 156 -996 157 -950
rect 198 -951 199 -915
rect 240 -951 241 -915
rect 261 -996 262 -950
rect 268 -996 269 -950
rect 366 -951 367 -915
rect 373 -951 374 -915
rect 723 -951 724 -915
rect 800 -996 801 -950
rect 856 -951 857 -915
rect 1059 -951 1060 -915
rect 1094 -996 1095 -950
rect 9 -996 10 -952
rect 121 -996 122 -952
rect 177 -953 178 -915
rect 212 -996 213 -952
rect 240 -996 241 -952
rect 254 -953 255 -915
rect 275 -953 276 -915
rect 296 -953 297 -915
rect 352 -953 353 -915
rect 366 -996 367 -952
rect 380 -996 381 -952
rect 387 -953 388 -915
rect 471 -953 472 -915
rect 569 -996 570 -952
rect 607 -996 608 -952
rect 1038 -996 1039 -952
rect 23 -955 24 -915
rect 254 -996 255 -954
rect 275 -996 276 -954
rect 282 -955 283 -915
rect 296 -996 297 -954
rect 317 -955 318 -915
rect 471 -996 472 -954
rect 583 -955 584 -915
rect 625 -955 626 -915
rect 863 -996 864 -954
rect 1024 -955 1025 -915
rect 1059 -996 1060 -954
rect 23 -996 24 -956
rect 100 -996 101 -956
rect 135 -957 136 -915
rect 352 -996 353 -956
rect 478 -996 479 -956
rect 520 -957 521 -915
rect 583 -996 584 -956
rect 660 -957 661 -915
rect 723 -996 724 -956
rect 779 -957 780 -915
rect 821 -957 822 -915
rect 1024 -996 1025 -956
rect 72 -996 73 -958
rect 198 -996 199 -958
rect 317 -996 318 -958
rect 450 -959 451 -915
rect 485 -996 486 -958
rect 527 -959 528 -915
rect 544 -996 545 -958
rect 660 -996 661 -958
rect 744 -959 745 -915
rect 779 -996 780 -958
rect 821 -996 822 -958
rect 905 -959 906 -915
rect 93 -996 94 -960
rect 1066 -996 1067 -960
rect 135 -996 136 -962
rect 614 -963 615 -915
rect 653 -996 654 -962
rect 688 -963 689 -915
rect 744 -996 745 -962
rect 793 -963 794 -915
rect 905 -996 906 -962
rect 954 -963 955 -915
rect 177 -996 178 -964
rect 184 -965 185 -915
rect 359 -965 360 -915
rect 520 -996 521 -964
rect 527 -996 528 -964
rect 534 -965 535 -915
rect 688 -996 689 -964
rect 751 -965 752 -915
rect 793 -996 794 -964
rect 807 -965 808 -915
rect 954 -996 955 -964
rect 968 -965 969 -915
rect 184 -996 185 -966
rect 282 -996 283 -966
rect 443 -967 444 -915
rect 534 -996 535 -966
rect 751 -996 752 -966
rect 849 -967 850 -915
rect 968 -996 969 -966
rect 1045 -967 1046 -915
rect 422 -969 423 -915
rect 1045 -996 1046 -968
rect 422 -996 423 -970
rect 464 -971 465 -915
rect 807 -996 808 -970
rect 877 -971 878 -915
rect 429 -973 430 -915
rect 443 -996 444 -972
rect 450 -996 451 -972
rect 590 -973 591 -915
rect 849 -996 850 -972
rect 891 -973 892 -915
rect 429 -996 430 -974
rect 457 -975 458 -915
rect 590 -996 591 -974
rect 835 -975 836 -915
rect 877 -996 878 -974
rect 919 -975 920 -915
rect 457 -996 458 -976
rect 639 -977 640 -915
rect 765 -977 766 -915
rect 891 -996 892 -976
rect 758 -979 759 -915
rect 765 -996 766 -978
rect 835 -996 836 -978
rect 947 -979 948 -915
rect 65 -996 66 -980
rect 758 -996 759 -980
rect 884 -981 885 -915
rect 919 -996 920 -980
rect 933 -981 934 -915
rect 947 -996 948 -980
rect 842 -983 843 -915
rect 933 -996 934 -982
rect 842 -996 843 -984
rect 901 -985 902 -915
rect 884 -996 885 -986
rect 926 -987 927 -915
rect 926 -996 927 -988
rect 940 -989 941 -915
rect 940 -996 941 -990
rect 1003 -991 1004 -915
rect 912 -993 913 -915
rect 1003 -996 1004 -992
rect 604 -996 605 -994
rect 912 -996 913 -994
rect 9 -1006 10 -1004
rect 93 -1071 94 -1005
rect 100 -1071 101 -1005
rect 107 -1006 108 -1004
rect 121 -1071 122 -1005
rect 338 -1006 339 -1004
rect 359 -1006 360 -1004
rect 422 -1006 423 -1004
rect 464 -1006 465 -1004
rect 513 -1006 514 -1004
rect 541 -1006 542 -1004
rect 765 -1006 766 -1004
rect 810 -1071 811 -1005
rect 954 -1006 955 -1004
rect 1003 -1006 1004 -1004
rect 1003 -1071 1004 -1005
rect 1003 -1006 1004 -1004
rect 1003 -1071 1004 -1005
rect 1129 -1006 1130 -1004
rect 1157 -1006 1158 -1004
rect 1185 -1006 1186 -1004
rect 1185 -1071 1186 -1005
rect 1185 -1006 1186 -1004
rect 1185 -1071 1186 -1005
rect 23 -1008 24 -1004
rect 23 -1071 24 -1007
rect 23 -1008 24 -1004
rect 23 -1071 24 -1007
rect 37 -1071 38 -1007
rect 65 -1008 66 -1004
rect 89 -1071 90 -1007
rect 863 -1008 864 -1004
rect 884 -1008 885 -1004
rect 887 -1060 888 -1007
rect 954 -1071 955 -1007
rect 1115 -1008 1116 -1004
rect 1136 -1008 1137 -1004
rect 1150 -1008 1151 -1004
rect 40 -1010 41 -1004
rect 544 -1010 545 -1004
rect 555 -1010 556 -1004
rect 555 -1071 556 -1009
rect 555 -1010 556 -1004
rect 555 -1071 556 -1009
rect 569 -1010 570 -1004
rect 607 -1010 608 -1004
rect 625 -1071 626 -1009
rect 723 -1010 724 -1004
rect 730 -1010 731 -1004
rect 1094 -1010 1095 -1004
rect 44 -1012 45 -1004
rect 198 -1012 199 -1004
rect 208 -1071 209 -1011
rect 212 -1012 213 -1004
rect 219 -1012 220 -1004
rect 355 -1071 356 -1011
rect 362 -1012 363 -1004
rect 1038 -1012 1039 -1004
rect 1094 -1071 1095 -1011
rect 1171 -1012 1172 -1004
rect 16 -1014 17 -1004
rect 44 -1071 45 -1013
rect 51 -1014 52 -1004
rect 51 -1071 52 -1013
rect 51 -1014 52 -1004
rect 51 -1071 52 -1013
rect 58 -1071 59 -1013
rect 72 -1014 73 -1004
rect 107 -1071 108 -1013
rect 394 -1014 395 -1004
rect 401 -1014 402 -1004
rect 513 -1071 514 -1013
rect 527 -1014 528 -1004
rect 541 -1071 542 -1013
rect 597 -1014 598 -1004
rect 642 -1014 643 -1004
rect 646 -1071 647 -1013
rect 674 -1014 675 -1004
rect 681 -1014 682 -1004
rect 705 -1060 706 -1013
rect 723 -1071 724 -1013
rect 835 -1014 836 -1004
rect 856 -1014 857 -1004
rect 1080 -1014 1081 -1004
rect 16 -1071 17 -1015
rect 103 -1016 104 -1004
rect 124 -1016 125 -1004
rect 359 -1071 360 -1015
rect 366 -1016 367 -1004
rect 366 -1071 367 -1015
rect 366 -1016 367 -1004
rect 366 -1071 367 -1015
rect 457 -1016 458 -1004
rect 527 -1071 528 -1015
rect 600 -1071 601 -1015
rect 793 -1016 794 -1004
rect 856 -1071 857 -1015
rect 877 -1016 878 -1004
rect 884 -1071 885 -1015
rect 905 -1016 906 -1004
rect 1024 -1016 1025 -1004
rect 1038 -1071 1039 -1015
rect 1069 -1071 1070 -1015
rect 1080 -1071 1081 -1015
rect 30 -1018 31 -1004
rect 219 -1071 220 -1017
rect 254 -1018 255 -1004
rect 387 -1071 388 -1017
rect 443 -1018 444 -1004
rect 457 -1071 458 -1017
rect 499 -1018 500 -1004
rect 982 -1018 983 -1004
rect 996 -1018 997 -1004
rect 1024 -1071 1025 -1017
rect 30 -1071 31 -1019
rect 142 -1020 143 -1004
rect 184 -1071 185 -1019
rect 282 -1020 283 -1004
rect 289 -1020 290 -1004
rect 320 -1071 321 -1019
rect 338 -1071 339 -1019
rect 380 -1020 381 -1004
rect 429 -1020 430 -1004
rect 443 -1071 444 -1019
rect 499 -1071 500 -1019
rect 583 -1020 584 -1004
rect 604 -1071 605 -1019
rect 691 -1071 692 -1019
rect 695 -1071 696 -1019
rect 737 -1020 738 -1004
rect 751 -1020 752 -1004
rect 765 -1071 766 -1019
rect 786 -1020 787 -1004
rect 835 -1071 836 -1019
rect 859 -1020 860 -1004
rect 1108 -1020 1109 -1004
rect 61 -1022 62 -1004
rect 548 -1022 549 -1004
rect 632 -1022 633 -1004
rect 674 -1071 675 -1021
rect 681 -1071 682 -1021
rect 688 -1022 689 -1004
rect 698 -1022 699 -1004
rect 793 -1071 794 -1021
rect 863 -1071 864 -1021
rect 898 -1022 899 -1004
rect 905 -1071 906 -1021
rect 968 -1022 969 -1004
rect 982 -1071 983 -1021
rect 1010 -1022 1011 -1004
rect 65 -1071 66 -1023
rect 408 -1024 409 -1004
rect 429 -1071 430 -1023
rect 485 -1024 486 -1004
rect 502 -1024 503 -1004
rect 1101 -1024 1102 -1004
rect 72 -1071 73 -1025
rect 275 -1026 276 -1004
rect 289 -1071 290 -1025
rect 296 -1026 297 -1004
rect 317 -1026 318 -1004
rect 422 -1071 423 -1025
rect 471 -1026 472 -1004
rect 583 -1071 584 -1025
rect 639 -1026 640 -1004
rect 1087 -1026 1088 -1004
rect 79 -1028 80 -1004
rect 282 -1071 283 -1027
rect 317 -1071 318 -1027
rect 597 -1071 598 -1027
rect 639 -1071 640 -1027
rect 653 -1028 654 -1004
rect 660 -1028 661 -1004
rect 737 -1071 738 -1027
rect 751 -1071 752 -1027
rect 821 -1028 822 -1004
rect 968 -1071 969 -1027
rect 989 -1028 990 -1004
rect 996 -1071 997 -1027
rect 1017 -1028 1018 -1004
rect 1087 -1071 1088 -1027
rect 1122 -1028 1123 -1004
rect 79 -1071 80 -1029
rect 149 -1030 150 -1004
rect 187 -1030 188 -1004
rect 779 -1030 780 -1004
rect 786 -1071 787 -1029
rect 919 -1030 920 -1004
rect 989 -1071 990 -1029
rect 1066 -1030 1067 -1004
rect 1122 -1071 1123 -1029
rect 1167 -1030 1168 -1004
rect 96 -1032 97 -1004
rect 394 -1071 395 -1031
rect 408 -1071 409 -1031
rect 415 -1032 416 -1004
rect 485 -1071 486 -1031
rect 562 -1032 563 -1004
rect 649 -1032 650 -1004
rect 891 -1032 892 -1004
rect 919 -1071 920 -1031
rect 1073 -1032 1074 -1004
rect 86 -1034 87 -1004
rect 96 -1071 97 -1033
rect 114 -1034 115 -1004
rect 142 -1071 143 -1033
rect 191 -1034 192 -1004
rect 198 -1071 199 -1033
rect 205 -1034 206 -1004
rect 471 -1071 472 -1033
rect 509 -1034 510 -1004
rect 534 -1034 535 -1004
rect 653 -1071 654 -1033
rect 702 -1034 703 -1004
rect 716 -1034 717 -1004
rect 877 -1071 878 -1033
rect 891 -1071 892 -1033
rect 912 -1034 913 -1004
rect 1010 -1071 1011 -1033
rect 1132 -1034 1133 -1004
rect 2 -1036 3 -1004
rect 205 -1071 206 -1035
rect 212 -1071 213 -1035
rect 240 -1036 241 -1004
rect 268 -1036 269 -1004
rect 373 -1036 374 -1004
rect 376 -1036 377 -1004
rect 898 -1071 899 -1035
rect 912 -1071 913 -1035
rect 926 -1036 927 -1004
rect 1017 -1071 1018 -1035
rect 1052 -1036 1053 -1004
rect 128 -1038 129 -1004
rect 128 -1071 129 -1037
rect 128 -1038 129 -1004
rect 128 -1071 129 -1037
rect 170 -1038 171 -1004
rect 268 -1071 269 -1037
rect 331 -1038 332 -1004
rect 548 -1071 549 -1037
rect 572 -1071 573 -1037
rect 926 -1071 927 -1037
rect 177 -1040 178 -1004
rect 191 -1071 192 -1039
rect 226 -1040 227 -1004
rect 275 -1071 276 -1039
rect 303 -1040 304 -1004
rect 331 -1071 332 -1039
rect 373 -1071 374 -1039
rect 478 -1040 479 -1004
rect 506 -1040 507 -1004
rect 702 -1071 703 -1039
rect 716 -1071 717 -1039
rect 772 -1040 773 -1004
rect 779 -1071 780 -1039
rect 807 -1040 808 -1004
rect 821 -1071 822 -1039
rect 870 -1040 871 -1004
rect 86 -1071 87 -1041
rect 226 -1071 227 -1041
rect 233 -1042 234 -1004
rect 254 -1071 255 -1041
rect 303 -1071 304 -1041
rect 310 -1042 311 -1004
rect 380 -1071 381 -1041
rect 436 -1042 437 -1004
rect 450 -1042 451 -1004
rect 562 -1071 563 -1041
rect 660 -1071 661 -1041
rect 667 -1042 668 -1004
rect 684 -1042 685 -1004
rect 1059 -1042 1060 -1004
rect 117 -1071 118 -1043
rect 233 -1071 234 -1043
rect 240 -1071 241 -1043
rect 264 -1071 265 -1043
rect 401 -1071 402 -1043
rect 436 -1071 437 -1043
rect 450 -1071 451 -1043
rect 611 -1044 612 -1004
rect 667 -1071 668 -1043
rect 709 -1044 710 -1004
rect 733 -1071 734 -1043
rect 1031 -1044 1032 -1004
rect 1059 -1071 1060 -1043
rect 1073 -1071 1074 -1043
rect 152 -1071 153 -1045
rect 310 -1071 311 -1045
rect 415 -1071 416 -1045
rect 621 -1071 622 -1045
rect 688 -1071 689 -1045
rect 814 -1046 815 -1004
rect 842 -1046 843 -1004
rect 870 -1071 871 -1045
rect 1031 -1071 1032 -1045
rect 1052 -1071 1053 -1045
rect 156 -1048 157 -1004
rect 177 -1071 178 -1047
rect 390 -1048 391 -1004
rect 842 -1071 843 -1047
rect 156 -1071 157 -1049
rect 163 -1050 164 -1004
rect 478 -1071 479 -1049
rect 492 -1050 493 -1004
rect 534 -1071 535 -1049
rect 933 -1050 934 -1004
rect 135 -1052 136 -1004
rect 163 -1071 164 -1051
rect 201 -1052 202 -1004
rect 933 -1071 934 -1051
rect 135 -1071 136 -1053
rect 324 -1054 325 -1004
rect 345 -1054 346 -1004
rect 492 -1071 493 -1053
rect 576 -1054 577 -1004
rect 611 -1071 612 -1053
rect 709 -1071 710 -1053
rect 744 -1054 745 -1004
rect 772 -1071 773 -1053
rect 800 -1054 801 -1004
rect 814 -1071 815 -1053
rect 849 -1054 850 -1004
rect 247 -1056 248 -1004
rect 324 -1071 325 -1055
rect 345 -1071 346 -1055
rect 352 -1056 353 -1004
rect 576 -1071 577 -1055
rect 618 -1056 619 -1004
rect 744 -1071 745 -1055
rect 828 -1056 829 -1004
rect 849 -1071 850 -1055
rect 1045 -1056 1046 -1004
rect 247 -1071 248 -1057
rect 261 -1058 262 -1004
rect 352 -1071 353 -1057
rect 590 -1058 591 -1004
rect 618 -1071 619 -1057
rect 947 -1058 948 -1004
rect 520 -1060 521 -1004
rect 590 -1071 591 -1059
rect 758 -1060 759 -1004
rect 828 -1071 829 -1059
rect 1066 -1071 1067 -1059
rect 173 -1071 174 -1061
rect 520 -1071 521 -1061
rect 800 -1071 801 -1061
rect 1143 -1062 1144 -1004
rect 940 -1064 941 -1004
rect 947 -1071 948 -1063
rect 940 -1071 941 -1065
rect 961 -1066 962 -1004
rect 961 -1071 962 -1067
rect 975 -1068 976 -1004
rect 61 -1071 62 -1069
rect 975 -1071 976 -1069
rect 16 -1081 17 -1079
rect 187 -1154 188 -1080
rect 219 -1081 220 -1079
rect 446 -1154 447 -1080
rect 471 -1081 472 -1079
rect 618 -1154 619 -1080
rect 632 -1081 633 -1079
rect 695 -1081 696 -1079
rect 852 -1154 853 -1080
rect 877 -1081 878 -1079
rect 884 -1081 885 -1079
rect 887 -1089 888 -1080
rect 912 -1081 913 -1079
rect 912 -1154 913 -1080
rect 912 -1081 913 -1079
rect 912 -1154 913 -1080
rect 954 -1154 955 -1080
rect 961 -1081 962 -1079
rect 978 -1154 979 -1080
rect 1017 -1081 1018 -1079
rect 1031 -1081 1032 -1079
rect 1038 -1154 1039 -1080
rect 1041 -1081 1042 -1079
rect 1052 -1081 1053 -1079
rect 1108 -1154 1109 -1080
rect 1122 -1081 1123 -1079
rect 1185 -1081 1186 -1079
rect 1188 -1154 1189 -1080
rect 23 -1083 24 -1079
rect 149 -1083 150 -1079
rect 170 -1083 171 -1079
rect 590 -1083 591 -1079
rect 600 -1083 601 -1079
rect 730 -1154 731 -1082
rect 856 -1083 857 -1079
rect 856 -1154 857 -1082
rect 856 -1083 857 -1079
rect 856 -1154 857 -1082
rect 877 -1154 878 -1082
rect 926 -1083 927 -1079
rect 940 -1083 941 -1079
rect 961 -1154 962 -1082
rect 996 -1083 997 -1079
rect 996 -1154 997 -1082
rect 996 -1083 997 -1079
rect 996 -1154 997 -1082
rect 1006 -1154 1007 -1082
rect 1094 -1083 1095 -1079
rect 30 -1085 31 -1079
rect 264 -1085 265 -1079
rect 268 -1085 269 -1079
rect 306 -1154 307 -1084
rect 345 -1085 346 -1079
rect 345 -1154 346 -1084
rect 345 -1085 346 -1079
rect 345 -1154 346 -1084
rect 355 -1085 356 -1079
rect 597 -1154 598 -1084
rect 607 -1154 608 -1084
rect 751 -1085 752 -1079
rect 884 -1154 885 -1084
rect 898 -1085 899 -1079
rect 940 -1154 941 -1084
rect 947 -1085 948 -1079
rect 1017 -1154 1018 -1084
rect 1024 -1085 1025 -1079
rect 1045 -1085 1046 -1079
rect 1059 -1154 1060 -1084
rect 30 -1154 31 -1086
rect 44 -1087 45 -1079
rect 51 -1087 52 -1079
rect 51 -1154 52 -1086
rect 51 -1087 52 -1079
rect 51 -1154 52 -1086
rect 58 -1154 59 -1086
rect 166 -1154 167 -1086
rect 170 -1154 171 -1086
rect 177 -1087 178 -1079
rect 191 -1087 192 -1079
rect 219 -1154 220 -1086
rect 247 -1087 248 -1079
rect 268 -1154 269 -1086
rect 275 -1087 276 -1079
rect 506 -1087 507 -1079
rect 509 -1087 510 -1079
rect 849 -1087 850 -1079
rect 891 -1087 892 -1079
rect 898 -1154 899 -1086
rect 947 -1154 948 -1086
rect 1003 -1087 1004 -1079
rect 1010 -1087 1011 -1079
rect 1024 -1154 1025 -1086
rect 1048 -1154 1049 -1086
rect 1087 -1087 1088 -1079
rect 37 -1089 38 -1079
rect 299 -1089 300 -1079
rect 387 -1089 388 -1079
rect 467 -1089 468 -1079
rect 485 -1089 486 -1079
rect 628 -1154 629 -1088
rect 639 -1089 640 -1079
rect 639 -1154 640 -1088
rect 639 -1089 640 -1079
rect 639 -1154 640 -1088
rect 660 -1089 661 -1079
rect 660 -1154 661 -1088
rect 660 -1089 661 -1079
rect 660 -1154 661 -1088
rect 667 -1089 668 -1079
rect 751 -1154 752 -1088
rect 891 -1154 892 -1088
rect 989 -1089 990 -1079
rect 1010 -1154 1011 -1088
rect 1080 -1089 1081 -1079
rect 1087 -1154 1088 -1088
rect 37 -1154 38 -1090
rect 128 -1091 129 -1079
rect 149 -1154 150 -1090
rect 156 -1091 157 -1079
rect 177 -1154 178 -1090
rect 212 -1091 213 -1079
rect 254 -1091 255 -1079
rect 254 -1154 255 -1090
rect 254 -1091 255 -1079
rect 254 -1154 255 -1090
rect 296 -1091 297 -1079
rect 611 -1091 612 -1079
rect 621 -1091 622 -1079
rect 632 -1154 633 -1090
rect 667 -1154 668 -1090
rect 842 -1091 843 -1079
rect 982 -1091 983 -1079
rect 989 -1154 990 -1090
rect 1073 -1091 1074 -1079
rect 1080 -1154 1081 -1090
rect 44 -1154 45 -1092
rect 450 -1093 451 -1079
rect 551 -1154 552 -1092
rect 576 -1093 577 -1079
rect 586 -1154 587 -1092
rect 926 -1154 927 -1092
rect 968 -1093 969 -1079
rect 982 -1154 983 -1092
rect 65 -1154 66 -1094
rect 68 -1095 69 -1079
rect 72 -1095 73 -1079
rect 464 -1095 465 -1079
rect 499 -1095 500 -1079
rect 576 -1154 577 -1094
rect 590 -1154 591 -1094
rect 737 -1095 738 -1079
rect 842 -1154 843 -1094
rect 870 -1095 871 -1079
rect 968 -1154 969 -1094
rect 975 -1095 976 -1079
rect 72 -1154 73 -1096
rect 82 -1154 83 -1096
rect 93 -1154 94 -1096
rect 100 -1097 101 -1079
rect 121 -1097 122 -1079
rect 352 -1154 353 -1096
rect 366 -1097 367 -1079
rect 464 -1154 465 -1096
rect 499 -1154 500 -1096
rect 555 -1097 556 -1079
rect 572 -1097 573 -1079
rect 583 -1097 584 -1079
rect 604 -1097 605 -1079
rect 611 -1154 612 -1096
rect 670 -1154 671 -1096
rect 1031 -1154 1032 -1096
rect 79 -1099 80 -1079
rect 128 -1154 129 -1098
rect 156 -1154 157 -1098
rect 534 -1099 535 -1079
rect 583 -1154 584 -1098
rect 653 -1099 654 -1079
rect 674 -1099 675 -1079
rect 674 -1154 675 -1098
rect 674 -1099 675 -1079
rect 674 -1154 675 -1098
rect 681 -1099 682 -1079
rect 695 -1154 696 -1098
rect 702 -1099 703 -1079
rect 870 -1154 871 -1098
rect 100 -1154 101 -1100
rect 117 -1154 118 -1100
rect 121 -1154 122 -1100
rect 184 -1101 185 -1079
rect 191 -1154 192 -1100
rect 324 -1101 325 -1079
rect 359 -1101 360 -1079
rect 702 -1154 703 -1100
rect 709 -1101 710 -1079
rect 737 -1154 738 -1100
rect 184 -1154 185 -1102
rect 418 -1154 419 -1102
rect 422 -1103 423 -1079
rect 471 -1154 472 -1102
rect 534 -1154 535 -1102
rect 733 -1103 734 -1079
rect 212 -1154 213 -1104
rect 331 -1105 332 -1079
rect 373 -1105 374 -1079
rect 555 -1154 556 -1104
rect 646 -1105 647 -1079
rect 709 -1154 710 -1104
rect 226 -1107 227 -1079
rect 366 -1154 367 -1106
rect 387 -1154 388 -1106
rect 513 -1107 514 -1079
rect 646 -1154 647 -1106
rect 919 -1107 920 -1079
rect 226 -1154 227 -1108
rect 247 -1154 248 -1108
rect 282 -1109 283 -1079
rect 324 -1154 325 -1108
rect 338 -1109 339 -1079
rect 373 -1154 374 -1108
rect 422 -1154 423 -1108
rect 569 -1109 570 -1079
rect 688 -1109 689 -1079
rect 723 -1109 724 -1079
rect 919 -1154 920 -1108
rect 933 -1109 934 -1079
rect 240 -1111 241 -1079
rect 359 -1154 360 -1110
rect 436 -1111 437 -1079
rect 478 -1111 479 -1079
rect 513 -1154 514 -1110
rect 527 -1111 528 -1079
rect 562 -1111 563 -1079
rect 569 -1154 570 -1110
rect 688 -1154 689 -1110
rect 800 -1111 801 -1079
rect 933 -1154 934 -1110
rect 1066 -1111 1067 -1079
rect 240 -1154 241 -1112
rect 537 -1113 538 -1079
rect 723 -1154 724 -1112
rect 828 -1113 829 -1079
rect 1003 -1154 1004 -1112
rect 1066 -1154 1067 -1112
rect 275 -1154 276 -1114
rect 282 -1154 283 -1114
rect 289 -1115 290 -1079
rect 296 -1154 297 -1114
rect 317 -1115 318 -1079
rect 681 -1154 682 -1114
rect 800 -1154 801 -1114
rect 814 -1115 815 -1079
rect 821 -1115 822 -1079
rect 828 -1154 829 -1114
rect 233 -1117 234 -1079
rect 289 -1154 290 -1116
rect 303 -1117 304 -1079
rect 317 -1154 318 -1116
rect 331 -1154 332 -1116
rect 436 -1154 437 -1116
rect 443 -1117 444 -1079
rect 485 -1154 486 -1116
rect 492 -1117 493 -1079
rect 562 -1154 563 -1116
rect 744 -1117 745 -1079
rect 821 -1154 822 -1116
rect 163 -1119 164 -1079
rect 233 -1154 234 -1118
rect 338 -1154 339 -1118
rect 415 -1119 416 -1079
rect 429 -1119 430 -1079
rect 492 -1154 493 -1118
rect 527 -1154 528 -1118
rect 541 -1119 542 -1079
rect 744 -1154 745 -1118
rect 863 -1119 864 -1079
rect 401 -1121 402 -1079
rect 429 -1154 430 -1120
rect 450 -1154 451 -1120
rect 457 -1121 458 -1079
rect 478 -1154 479 -1120
rect 807 -1154 808 -1120
rect 814 -1154 815 -1120
rect 835 -1121 836 -1079
rect 205 -1123 206 -1079
rect 457 -1154 458 -1122
rect 541 -1154 542 -1122
rect 625 -1123 626 -1079
rect 653 -1154 654 -1122
rect 835 -1154 836 -1122
rect 198 -1125 199 -1079
rect 205 -1154 206 -1124
rect 261 -1125 262 -1079
rect 401 -1154 402 -1124
rect 408 -1125 409 -1079
rect 415 -1154 416 -1124
rect 793 -1125 794 -1079
rect 863 -1154 864 -1124
rect 261 -1154 262 -1126
rect 310 -1127 311 -1079
rect 779 -1127 780 -1079
rect 793 -1154 794 -1126
rect 310 -1154 311 -1128
rect 810 -1129 811 -1079
rect 772 -1131 773 -1079
rect 779 -1154 780 -1130
rect 810 -1154 811 -1130
rect 905 -1131 906 -1079
rect 758 -1133 759 -1079
rect 772 -1154 773 -1132
rect 786 -1133 787 -1079
rect 905 -1154 906 -1132
rect 716 -1135 717 -1079
rect 786 -1154 787 -1134
rect 520 -1137 521 -1079
rect 716 -1154 717 -1136
rect 758 -1154 759 -1136
rect 765 -1137 766 -1079
rect 520 -1154 521 -1138
rect 957 -1139 958 -1079
rect 548 -1141 549 -1079
rect 765 -1154 766 -1140
rect 394 -1143 395 -1079
rect 548 -1154 549 -1142
rect 380 -1145 381 -1079
rect 394 -1154 395 -1144
rect 107 -1147 108 -1079
rect 380 -1154 381 -1146
rect 107 -1154 108 -1148
rect 142 -1149 143 -1079
rect 135 -1151 136 -1079
rect 142 -1154 143 -1150
rect 135 -1154 136 -1152
rect 408 -1154 409 -1152
rect 16 -1229 17 -1163
rect 121 -1164 122 -1162
rect 142 -1164 143 -1162
rect 142 -1229 143 -1163
rect 142 -1164 143 -1162
rect 142 -1229 143 -1163
rect 149 -1164 150 -1162
rect 163 -1164 164 -1162
rect 170 -1164 171 -1162
rect 198 -1164 199 -1162
rect 205 -1164 206 -1162
rect 205 -1229 206 -1163
rect 205 -1164 206 -1162
rect 205 -1229 206 -1163
rect 219 -1164 220 -1162
rect 219 -1229 220 -1163
rect 219 -1164 220 -1162
rect 219 -1229 220 -1163
rect 226 -1229 227 -1163
rect 268 -1164 269 -1162
rect 285 -1164 286 -1162
rect 317 -1164 318 -1162
rect 331 -1229 332 -1163
rect 352 -1164 353 -1162
rect 422 -1164 423 -1162
rect 422 -1229 423 -1163
rect 422 -1164 423 -1162
rect 422 -1229 423 -1163
rect 446 -1164 447 -1162
rect 933 -1229 934 -1163
rect 975 -1164 976 -1162
rect 1038 -1164 1039 -1162
rect 1066 -1164 1067 -1162
rect 1122 -1229 1123 -1163
rect 23 -1166 24 -1162
rect 26 -1229 27 -1165
rect 30 -1166 31 -1162
rect 156 -1166 157 -1162
rect 163 -1229 164 -1165
rect 247 -1166 248 -1162
rect 254 -1166 255 -1162
rect 667 -1166 668 -1162
rect 695 -1166 696 -1162
rect 807 -1229 808 -1165
rect 828 -1166 829 -1162
rect 936 -1166 937 -1162
rect 961 -1166 962 -1162
rect 975 -1229 976 -1165
rect 982 -1166 983 -1162
rect 982 -1229 983 -1165
rect 982 -1166 983 -1162
rect 982 -1229 983 -1165
rect 989 -1166 990 -1162
rect 1066 -1229 1067 -1165
rect 1080 -1166 1081 -1162
rect 1129 -1229 1130 -1165
rect 30 -1229 31 -1167
rect 499 -1168 500 -1162
rect 506 -1168 507 -1162
rect 555 -1168 556 -1162
rect 562 -1168 563 -1162
rect 604 -1168 605 -1162
rect 618 -1168 619 -1162
rect 656 -1168 657 -1162
rect 667 -1229 668 -1167
rect 688 -1168 689 -1162
rect 695 -1229 696 -1167
rect 765 -1168 766 -1162
rect 831 -1229 832 -1167
rect 877 -1168 878 -1162
rect 884 -1168 885 -1162
rect 961 -1229 962 -1167
rect 996 -1168 997 -1162
rect 1003 -1229 1004 -1167
rect 1010 -1168 1011 -1162
rect 1038 -1229 1039 -1167
rect 1087 -1168 1088 -1162
rect 1115 -1229 1116 -1167
rect 37 -1170 38 -1162
rect 138 -1170 139 -1162
rect 152 -1229 153 -1169
rect 478 -1170 479 -1162
rect 499 -1229 500 -1169
rect 509 -1170 510 -1162
rect 544 -1229 545 -1169
rect 884 -1229 885 -1169
rect 905 -1170 906 -1162
rect 905 -1229 906 -1169
rect 905 -1170 906 -1162
rect 905 -1229 906 -1169
rect 919 -1170 920 -1162
rect 996 -1229 997 -1169
rect 1024 -1170 1025 -1162
rect 1052 -1229 1053 -1169
rect 1101 -1229 1102 -1169
rect 1108 -1170 1109 -1162
rect 37 -1229 38 -1171
rect 726 -1229 727 -1171
rect 730 -1172 731 -1162
rect 1080 -1229 1081 -1171
rect 44 -1174 45 -1162
rect 114 -1174 115 -1162
rect 117 -1174 118 -1162
rect 121 -1229 122 -1173
rect 170 -1229 171 -1173
rect 275 -1174 276 -1162
rect 352 -1229 353 -1173
rect 593 -1229 594 -1173
rect 607 -1174 608 -1162
rect 877 -1229 878 -1173
rect 926 -1174 927 -1162
rect 1073 -1229 1074 -1173
rect 58 -1176 59 -1162
rect 156 -1229 157 -1175
rect 177 -1176 178 -1162
rect 198 -1229 199 -1175
rect 229 -1176 230 -1162
rect 359 -1176 360 -1162
rect 443 -1229 444 -1175
rect 1010 -1229 1011 -1175
rect 1031 -1176 1032 -1162
rect 1087 -1229 1088 -1175
rect 51 -1178 52 -1162
rect 58 -1229 59 -1177
rect 72 -1178 73 -1162
rect 128 -1229 129 -1177
rect 184 -1229 185 -1177
rect 345 -1178 346 -1162
rect 359 -1229 360 -1177
rect 380 -1178 381 -1162
rect 478 -1229 479 -1177
rect 485 -1178 486 -1162
rect 562 -1229 563 -1177
rect 821 -1178 822 -1162
rect 842 -1178 843 -1162
rect 919 -1229 920 -1177
rect 954 -1178 955 -1162
rect 989 -1229 990 -1177
rect 1017 -1178 1018 -1162
rect 1031 -1229 1032 -1177
rect 1059 -1178 1060 -1162
rect 1108 -1229 1109 -1177
rect 65 -1180 66 -1162
rect 72 -1229 73 -1179
rect 79 -1229 80 -1179
rect 583 -1180 584 -1162
rect 586 -1180 587 -1162
rect 723 -1180 724 -1162
rect 730 -1229 731 -1179
rect 793 -1180 794 -1162
rect 814 -1180 815 -1162
rect 842 -1229 843 -1179
rect 849 -1229 850 -1179
rect 891 -1180 892 -1162
rect 940 -1180 941 -1162
rect 1017 -1229 1018 -1179
rect 51 -1229 52 -1181
rect 65 -1229 66 -1181
rect 82 -1182 83 -1162
rect 338 -1182 339 -1162
rect 429 -1182 430 -1162
rect 583 -1229 584 -1181
rect 590 -1182 591 -1162
rect 604 -1229 605 -1181
rect 625 -1182 626 -1162
rect 1045 -1229 1046 -1181
rect 89 -1184 90 -1162
rect 135 -1229 136 -1183
rect 187 -1184 188 -1162
rect 814 -1229 815 -1183
rect 863 -1184 864 -1162
rect 978 -1184 979 -1162
rect 93 -1186 94 -1162
rect 93 -1229 94 -1185
rect 93 -1186 94 -1162
rect 93 -1229 94 -1185
rect 100 -1186 101 -1162
rect 100 -1229 101 -1185
rect 100 -1186 101 -1162
rect 100 -1229 101 -1185
rect 107 -1186 108 -1162
rect 345 -1229 346 -1185
rect 429 -1229 430 -1185
rect 646 -1186 647 -1162
rect 653 -1229 654 -1185
rect 716 -1186 717 -1162
rect 765 -1229 766 -1185
rect 856 -1186 857 -1162
rect 870 -1186 871 -1162
rect 926 -1229 927 -1185
rect 968 -1186 969 -1162
rect 1059 -1229 1060 -1185
rect 61 -1229 62 -1187
rect 968 -1229 969 -1187
rect 107 -1229 108 -1189
rect 383 -1229 384 -1189
rect 450 -1190 451 -1162
rect 485 -1229 486 -1189
rect 565 -1229 566 -1189
rect 870 -1229 871 -1189
rect 891 -1229 892 -1189
rect 912 -1190 913 -1162
rect 233 -1192 234 -1162
rect 303 -1229 304 -1191
rect 306 -1192 307 -1162
rect 338 -1229 339 -1191
rect 401 -1192 402 -1162
rect 450 -1229 451 -1191
rect 569 -1192 570 -1162
rect 618 -1229 619 -1191
rect 625 -1229 626 -1191
rect 639 -1192 640 -1162
rect 646 -1229 647 -1191
rect 674 -1192 675 -1162
rect 688 -1229 689 -1191
rect 758 -1192 759 -1162
rect 772 -1192 773 -1162
rect 1024 -1229 1025 -1191
rect 131 -1194 132 -1162
rect 758 -1229 759 -1193
rect 772 -1229 773 -1193
rect 1094 -1229 1095 -1193
rect 233 -1229 234 -1195
rect 548 -1229 549 -1195
rect 555 -1229 556 -1195
rect 569 -1229 570 -1195
rect 611 -1196 612 -1162
rect 863 -1229 864 -1195
rect 898 -1196 899 -1162
rect 940 -1229 941 -1195
rect 240 -1198 241 -1162
rect 247 -1229 248 -1197
rect 254 -1229 255 -1197
rect 810 -1198 811 -1162
rect 898 -1229 899 -1197
rect 947 -1198 948 -1162
rect 240 -1229 241 -1199
rect 289 -1200 290 -1162
rect 317 -1229 318 -1199
rect 716 -1229 717 -1199
rect 744 -1200 745 -1162
rect 912 -1229 913 -1199
rect 261 -1202 262 -1162
rect 282 -1229 283 -1201
rect 289 -1229 290 -1201
rect 296 -1202 297 -1162
rect 394 -1202 395 -1162
rect 401 -1229 402 -1201
rect 597 -1202 598 -1162
rect 744 -1229 745 -1201
rect 779 -1202 780 -1162
rect 821 -1229 822 -1201
rect 166 -1204 167 -1162
rect 394 -1229 395 -1203
rect 408 -1204 409 -1162
rect 779 -1229 780 -1203
rect 786 -1204 787 -1162
rect 793 -1229 794 -1203
rect 800 -1204 801 -1162
rect 856 -1229 857 -1203
rect 212 -1206 213 -1162
rect 296 -1229 297 -1205
rect 408 -1229 409 -1205
rect 457 -1206 458 -1162
rect 509 -1229 510 -1205
rect 800 -1229 801 -1205
rect 191 -1208 192 -1162
rect 212 -1229 213 -1207
rect 268 -1229 269 -1207
rect 310 -1208 311 -1162
rect 457 -1229 458 -1207
rect 471 -1208 472 -1162
rect 534 -1208 535 -1162
rect 597 -1229 598 -1207
rect 611 -1229 612 -1207
rect 656 -1229 657 -1207
rect 674 -1229 675 -1207
rect 737 -1208 738 -1162
rect 751 -1208 752 -1162
rect 786 -1229 787 -1207
rect 191 -1229 192 -1209
rect 520 -1210 521 -1162
rect 527 -1210 528 -1162
rect 534 -1229 535 -1209
rect 660 -1210 661 -1162
rect 737 -1229 738 -1209
rect 751 -1229 752 -1209
rect 835 -1210 836 -1162
rect 275 -1229 276 -1211
rect 373 -1212 374 -1162
rect 464 -1212 465 -1162
rect 471 -1229 472 -1211
rect 513 -1212 514 -1162
rect 520 -1229 521 -1211
rect 527 -1229 528 -1211
rect 551 -1212 552 -1162
rect 681 -1212 682 -1162
rect 947 -1229 948 -1211
rect 23 -1229 24 -1213
rect 464 -1229 465 -1213
rect 541 -1214 542 -1162
rect 835 -1229 836 -1213
rect 310 -1229 311 -1215
rect 324 -1216 325 -1162
rect 436 -1216 437 -1162
rect 513 -1229 514 -1215
rect 681 -1229 682 -1215
rect 709 -1216 710 -1162
rect 324 -1229 325 -1217
rect 387 -1218 388 -1162
rect 436 -1229 437 -1217
rect 492 -1218 493 -1162
rect 632 -1218 633 -1162
rect 709 -1229 710 -1217
rect 492 -1229 493 -1219
rect 723 -1229 724 -1219
rect 576 -1222 577 -1162
rect 632 -1229 633 -1221
rect 702 -1222 703 -1162
rect 954 -1229 955 -1221
rect 366 -1224 367 -1162
rect 576 -1229 577 -1223
rect 366 -1229 367 -1225
rect 373 -1229 374 -1225
rect 415 -1226 416 -1162
rect 702 -1229 703 -1225
rect 415 -1229 416 -1227
rect 828 -1229 829 -1227
rect 30 -1239 31 -1237
rect 565 -1239 566 -1237
rect 569 -1239 570 -1237
rect 726 -1239 727 -1237
rect 772 -1300 773 -1238
rect 821 -1239 822 -1237
rect 828 -1239 829 -1237
rect 1017 -1239 1018 -1237
rect 1101 -1239 1102 -1237
rect 1101 -1300 1102 -1238
rect 1101 -1239 1102 -1237
rect 1101 -1300 1102 -1238
rect 47 -1241 48 -1237
rect 177 -1241 178 -1237
rect 180 -1241 181 -1237
rect 464 -1241 465 -1237
rect 481 -1300 482 -1240
rect 863 -1241 864 -1237
rect 866 -1300 867 -1240
rect 905 -1241 906 -1237
rect 999 -1300 1000 -1240
rect 1031 -1241 1032 -1237
rect 68 -1243 69 -1237
rect 72 -1243 73 -1237
rect 86 -1300 87 -1242
rect 163 -1243 164 -1237
rect 177 -1300 178 -1242
rect 205 -1243 206 -1237
rect 212 -1243 213 -1237
rect 390 -1243 391 -1237
rect 394 -1243 395 -1237
rect 775 -1243 776 -1237
rect 807 -1243 808 -1237
rect 1031 -1300 1032 -1242
rect 72 -1300 73 -1244
rect 387 -1245 388 -1237
rect 394 -1300 395 -1244
rect 467 -1300 468 -1244
rect 509 -1245 510 -1237
rect 534 -1245 535 -1237
rect 541 -1300 542 -1244
rect 579 -1300 580 -1244
rect 590 -1245 591 -1237
rect 1059 -1245 1060 -1237
rect 93 -1247 94 -1237
rect 96 -1300 97 -1246
rect 100 -1247 101 -1237
rect 100 -1300 101 -1246
rect 100 -1247 101 -1237
rect 100 -1300 101 -1246
rect 114 -1300 115 -1246
rect 128 -1247 129 -1237
rect 149 -1247 150 -1237
rect 562 -1247 563 -1237
rect 590 -1300 591 -1246
rect 618 -1247 619 -1237
rect 625 -1247 626 -1237
rect 625 -1300 626 -1246
rect 625 -1247 626 -1237
rect 625 -1300 626 -1246
rect 642 -1247 643 -1237
rect 835 -1247 836 -1237
rect 905 -1300 906 -1246
rect 1052 -1247 1053 -1237
rect 1059 -1300 1060 -1246
rect 1115 -1247 1116 -1237
rect 16 -1249 17 -1237
rect 149 -1300 150 -1248
rect 163 -1300 164 -1248
rect 289 -1249 290 -1237
rect 324 -1249 325 -1237
rect 380 -1249 381 -1237
rect 387 -1300 388 -1248
rect 408 -1249 409 -1237
rect 443 -1300 444 -1248
rect 478 -1249 479 -1237
rect 544 -1249 545 -1237
rect 947 -1249 948 -1237
rect 1017 -1300 1018 -1248
rect 1073 -1249 1074 -1237
rect 117 -1251 118 -1237
rect 212 -1300 213 -1250
rect 219 -1251 220 -1237
rect 219 -1300 220 -1250
rect 219 -1251 220 -1237
rect 219 -1300 220 -1250
rect 233 -1251 234 -1237
rect 502 -1300 503 -1250
rect 548 -1251 549 -1237
rect 1024 -1251 1025 -1237
rect 1052 -1300 1053 -1250
rect 1097 -1300 1098 -1250
rect 128 -1300 129 -1252
rect 198 -1253 199 -1237
rect 205 -1300 206 -1252
rect 254 -1253 255 -1237
rect 264 -1253 265 -1237
rect 352 -1253 353 -1237
rect 373 -1300 374 -1252
rect 555 -1253 556 -1237
rect 618 -1300 619 -1252
rect 639 -1253 640 -1237
rect 656 -1253 657 -1237
rect 961 -1253 962 -1237
rect 184 -1255 185 -1237
rect 261 -1300 262 -1254
rect 289 -1300 290 -1254
rect 296 -1255 297 -1237
rect 324 -1300 325 -1254
rect 422 -1255 423 -1237
rect 478 -1300 479 -1254
rect 604 -1255 605 -1237
rect 639 -1300 640 -1254
rect 667 -1255 668 -1237
rect 677 -1300 678 -1254
rect 730 -1255 731 -1237
rect 796 -1300 797 -1254
rect 947 -1300 948 -1254
rect 961 -1300 962 -1254
rect 1087 -1255 1088 -1237
rect 184 -1300 185 -1256
rect 226 -1257 227 -1237
rect 233 -1300 234 -1256
rect 310 -1257 311 -1237
rect 341 -1300 342 -1256
rect 583 -1257 584 -1237
rect 604 -1300 605 -1256
rect 646 -1257 647 -1237
rect 656 -1300 657 -1256
rect 737 -1257 738 -1237
rect 807 -1300 808 -1256
rect 877 -1257 878 -1237
rect 1087 -1300 1088 -1256
rect 1122 -1257 1123 -1237
rect 156 -1259 157 -1237
rect 226 -1300 227 -1258
rect 240 -1259 241 -1237
rect 446 -1259 447 -1237
rect 506 -1259 507 -1237
rect 555 -1300 556 -1258
rect 572 -1259 573 -1237
rect 737 -1300 738 -1258
rect 821 -1300 822 -1258
rect 1062 -1300 1063 -1258
rect 152 -1261 153 -1237
rect 156 -1300 157 -1260
rect 191 -1261 192 -1237
rect 320 -1261 321 -1237
rect 345 -1261 346 -1237
rect 380 -1300 381 -1260
rect 404 -1300 405 -1260
rect 429 -1261 430 -1237
rect 506 -1300 507 -1260
rect 527 -1261 528 -1237
rect 548 -1300 549 -1260
rect 597 -1261 598 -1237
rect 646 -1300 647 -1260
rect 674 -1261 675 -1237
rect 709 -1261 710 -1237
rect 996 -1261 997 -1237
rect 198 -1300 199 -1262
rect 240 -1300 241 -1262
rect 254 -1300 255 -1262
rect 268 -1263 269 -1237
rect 282 -1263 283 -1237
rect 345 -1300 346 -1262
rect 352 -1300 353 -1262
rect 576 -1263 577 -1237
rect 583 -1300 584 -1262
rect 674 -1300 675 -1262
rect 709 -1300 710 -1262
rect 814 -1263 815 -1237
rect 828 -1300 829 -1262
rect 912 -1263 913 -1237
rect 121 -1265 122 -1237
rect 282 -1300 283 -1264
rect 296 -1300 297 -1264
rect 303 -1265 304 -1237
rect 310 -1300 311 -1264
rect 632 -1265 633 -1237
rect 660 -1265 661 -1237
rect 670 -1275 671 -1264
rect 723 -1265 724 -1237
rect 1066 -1265 1067 -1237
rect 107 -1267 108 -1237
rect 121 -1300 122 -1266
rect 268 -1300 269 -1266
rect 275 -1267 276 -1237
rect 317 -1267 318 -1237
rect 572 -1300 573 -1266
rect 660 -1300 661 -1266
rect 681 -1267 682 -1237
rect 723 -1300 724 -1266
rect 758 -1267 759 -1237
rect 814 -1300 815 -1266
rect 978 -1300 979 -1266
rect 1066 -1300 1067 -1266
rect 1108 -1267 1109 -1237
rect 79 -1269 80 -1237
rect 275 -1300 276 -1268
rect 366 -1269 367 -1237
rect 527 -1300 528 -1268
rect 663 -1269 664 -1237
rect 793 -1269 794 -1237
rect 835 -1300 836 -1268
rect 849 -1269 850 -1237
rect 877 -1300 878 -1268
rect 940 -1269 941 -1237
rect 79 -1300 80 -1270
rect 135 -1271 136 -1237
rect 247 -1271 248 -1237
rect 317 -1300 318 -1270
rect 376 -1271 377 -1237
rect 471 -1271 472 -1237
rect 667 -1300 668 -1270
rect 702 -1271 703 -1237
rect 730 -1300 731 -1270
rect 779 -1271 780 -1237
rect 793 -1300 794 -1270
rect 898 -1271 899 -1237
rect 912 -1300 913 -1270
rect 1045 -1271 1046 -1237
rect 37 -1273 38 -1237
rect 135 -1300 136 -1272
rect 247 -1300 248 -1272
rect 359 -1273 360 -1237
rect 408 -1300 409 -1272
rect 450 -1273 451 -1237
rect 464 -1300 465 -1272
rect 898 -1300 899 -1272
rect 940 -1300 941 -1272
rect 1038 -1273 1039 -1237
rect 1045 -1300 1046 -1272
rect 1094 -1273 1095 -1237
rect 107 -1300 108 -1274
rect 170 -1275 171 -1237
rect 359 -1300 360 -1274
rect 492 -1275 493 -1237
rect 681 -1300 682 -1274
rect 702 -1300 703 -1274
rect 716 -1275 717 -1237
rect 751 -1275 752 -1237
rect 758 -1300 759 -1274
rect 779 -1300 780 -1274
rect 884 -1275 885 -1237
rect 142 -1277 143 -1237
rect 170 -1300 171 -1276
rect 338 -1277 339 -1237
rect 492 -1300 493 -1276
rect 695 -1277 696 -1237
rect 716 -1300 717 -1276
rect 751 -1300 752 -1276
rect 765 -1277 766 -1237
rect 849 -1300 850 -1276
rect 919 -1277 920 -1237
rect 142 -1300 143 -1278
rect 331 -1279 332 -1237
rect 338 -1300 339 -1278
rect 366 -1300 367 -1278
rect 415 -1279 416 -1237
rect 471 -1300 472 -1278
rect 695 -1300 696 -1278
rect 744 -1279 745 -1237
rect 765 -1300 766 -1278
rect 954 -1279 955 -1237
rect 303 -1300 304 -1280
rect 331 -1300 332 -1280
rect 401 -1281 402 -1237
rect 415 -1300 416 -1280
rect 429 -1300 430 -1280
rect 457 -1281 458 -1237
rect 688 -1281 689 -1237
rect 744 -1300 745 -1280
rect 856 -1281 857 -1237
rect 1038 -1300 1039 -1280
rect 44 -1283 45 -1237
rect 401 -1300 402 -1282
rect 436 -1283 437 -1237
rect 457 -1300 458 -1282
rect 688 -1300 689 -1282
rect 786 -1283 787 -1237
rect 856 -1300 857 -1282
rect 933 -1283 934 -1237
rect 954 -1300 955 -1282
rect 982 -1283 983 -1237
rect 44 -1300 45 -1284
rect 51 -1285 52 -1237
rect 436 -1300 437 -1284
rect 520 -1285 521 -1237
rect 786 -1300 787 -1284
rect 842 -1285 843 -1237
rect 884 -1300 885 -1284
rect 1027 -1300 1028 -1284
rect 450 -1300 451 -1286
rect 485 -1287 486 -1237
rect 520 -1300 521 -1286
rect 611 -1287 612 -1237
rect 842 -1300 843 -1286
rect 926 -1287 927 -1237
rect 933 -1300 934 -1286
rect 1003 -1287 1004 -1237
rect 485 -1300 486 -1288
rect 513 -1289 514 -1237
rect 562 -1300 563 -1288
rect 611 -1300 612 -1288
rect 891 -1289 892 -1237
rect 982 -1300 983 -1288
rect 1003 -1300 1004 -1288
rect 1010 -1289 1011 -1237
rect 499 -1291 500 -1237
rect 513 -1300 514 -1290
rect 800 -1291 801 -1237
rect 1010 -1300 1011 -1290
rect 422 -1300 423 -1292
rect 499 -1300 500 -1292
rect 800 -1300 801 -1292
rect 870 -1293 871 -1237
rect 891 -1300 892 -1292
rect 989 -1293 990 -1237
rect 870 -1300 871 -1294
rect 968 -1295 969 -1237
rect 989 -1300 990 -1294
rect 1080 -1295 1081 -1237
rect 926 -1300 927 -1296
rect 1024 -1300 1025 -1296
rect 1080 -1300 1081 -1296
rect 1129 -1297 1130 -1237
rect 968 -1300 969 -1298
rect 975 -1299 976 -1237
rect 9 -1371 10 -1309
rect 30 -1371 31 -1309
rect 37 -1371 38 -1309
rect 114 -1310 115 -1308
rect 135 -1310 136 -1308
rect 369 -1371 370 -1309
rect 408 -1310 409 -1308
rect 481 -1310 482 -1308
rect 499 -1371 500 -1309
rect 513 -1310 514 -1308
rect 534 -1310 535 -1308
rect 590 -1310 591 -1308
rect 611 -1371 612 -1309
rect 625 -1310 626 -1308
rect 628 -1371 629 -1309
rect 919 -1371 920 -1309
rect 922 -1310 923 -1308
rect 968 -1310 969 -1308
rect 975 -1310 976 -1308
rect 982 -1310 983 -1308
rect 996 -1371 997 -1309
rect 1003 -1310 1004 -1308
rect 1020 -1310 1021 -1308
rect 1066 -1310 1067 -1308
rect 1097 -1310 1098 -1308
rect 1101 -1310 1102 -1308
rect 16 -1371 17 -1311
rect 72 -1312 73 -1308
rect 93 -1312 94 -1308
rect 100 -1312 101 -1308
rect 114 -1371 115 -1311
rect 201 -1371 202 -1311
rect 212 -1312 213 -1308
rect 338 -1371 339 -1311
rect 380 -1312 381 -1308
rect 590 -1371 591 -1311
rect 614 -1312 615 -1308
rect 751 -1312 752 -1308
rect 793 -1312 794 -1308
rect 1010 -1312 1011 -1308
rect 1059 -1312 1060 -1308
rect 1087 -1312 1088 -1308
rect 23 -1371 24 -1313
rect 240 -1314 241 -1308
rect 261 -1314 262 -1308
rect 348 -1371 349 -1313
rect 380 -1371 381 -1313
rect 422 -1314 423 -1308
rect 429 -1314 430 -1308
rect 464 -1314 465 -1308
rect 471 -1314 472 -1308
rect 513 -1371 514 -1313
rect 527 -1314 528 -1308
rect 751 -1371 752 -1313
rect 793 -1371 794 -1313
rect 1031 -1314 1032 -1308
rect 1066 -1371 1067 -1313
rect 1080 -1314 1081 -1308
rect 44 -1316 45 -1308
rect 44 -1371 45 -1315
rect 44 -1316 45 -1308
rect 44 -1371 45 -1315
rect 51 -1371 52 -1315
rect 247 -1316 248 -1308
rect 268 -1316 269 -1308
rect 303 -1316 304 -1308
rect 310 -1316 311 -1308
rect 597 -1316 598 -1308
rect 625 -1371 626 -1315
rect 702 -1316 703 -1308
rect 726 -1371 727 -1315
rect 1024 -1371 1025 -1315
rect 1031 -1371 1032 -1315
rect 1052 -1316 1053 -1308
rect 58 -1371 59 -1317
rect 537 -1318 538 -1308
rect 555 -1318 556 -1308
rect 569 -1318 570 -1308
rect 576 -1318 577 -1308
rect 600 -1318 601 -1308
rect 653 -1371 654 -1317
rect 744 -1318 745 -1308
rect 863 -1318 864 -1308
rect 940 -1318 941 -1308
rect 961 -1318 962 -1308
rect 1010 -1371 1011 -1317
rect 68 -1371 69 -1319
rect 306 -1320 307 -1308
rect 408 -1371 409 -1319
rect 485 -1320 486 -1308
rect 492 -1320 493 -1308
rect 534 -1371 535 -1319
rect 541 -1320 542 -1308
rect 555 -1371 556 -1319
rect 597 -1371 598 -1319
rect 604 -1320 605 -1308
rect 667 -1320 668 -1308
rect 667 -1371 668 -1319
rect 667 -1320 668 -1308
rect 667 -1371 668 -1319
rect 677 -1320 678 -1308
rect 702 -1371 703 -1319
rect 709 -1320 710 -1308
rect 744 -1371 745 -1319
rect 821 -1320 822 -1308
rect 863 -1371 864 -1319
rect 905 -1320 906 -1308
rect 968 -1371 969 -1319
rect 999 -1371 1000 -1319
rect 1045 -1320 1046 -1308
rect 72 -1371 73 -1321
rect 544 -1371 545 -1321
rect 569 -1371 570 -1321
rect 604 -1371 605 -1321
rect 681 -1322 682 -1308
rect 709 -1371 710 -1321
rect 733 -1371 734 -1321
rect 765 -1322 766 -1308
rect 870 -1322 871 -1308
rect 905 -1371 906 -1321
rect 912 -1322 913 -1308
rect 975 -1371 976 -1321
rect 93 -1371 94 -1323
rect 481 -1371 482 -1323
rect 506 -1324 507 -1308
rect 632 -1371 633 -1323
rect 695 -1324 696 -1308
rect 695 -1371 696 -1323
rect 695 -1324 696 -1308
rect 695 -1371 696 -1323
rect 737 -1324 738 -1308
rect 740 -1340 741 -1323
rect 758 -1324 759 -1308
rect 821 -1371 822 -1323
rect 870 -1371 871 -1323
rect 884 -1324 885 -1308
rect 891 -1324 892 -1308
rect 912 -1371 913 -1323
rect 933 -1324 934 -1308
rect 961 -1371 962 -1323
rect 100 -1371 101 -1325
rect 352 -1326 353 -1308
rect 411 -1371 412 -1325
rect 681 -1371 682 -1325
rect 723 -1326 724 -1308
rect 758 -1371 759 -1325
rect 765 -1371 766 -1325
rect 786 -1326 787 -1308
rect 877 -1326 878 -1308
rect 884 -1371 885 -1325
rect 891 -1371 892 -1325
rect 1017 -1326 1018 -1308
rect 128 -1328 129 -1308
rect 261 -1371 262 -1327
rect 268 -1371 269 -1327
rect 296 -1328 297 -1308
rect 345 -1328 346 -1308
rect 352 -1371 353 -1327
rect 422 -1371 423 -1327
rect 443 -1328 444 -1308
rect 471 -1371 472 -1327
rect 520 -1328 521 -1308
rect 527 -1371 528 -1327
rect 583 -1328 584 -1308
rect 660 -1328 661 -1308
rect 1017 -1371 1018 -1327
rect 86 -1330 87 -1308
rect 296 -1371 297 -1329
rect 345 -1371 346 -1329
rect 982 -1371 983 -1329
rect 86 -1371 87 -1331
rect 275 -1332 276 -1308
rect 285 -1371 286 -1331
rect 485 -1371 486 -1331
rect 506 -1371 507 -1331
rect 1003 -1371 1004 -1331
rect 128 -1371 129 -1333
rect 359 -1334 360 -1308
rect 366 -1334 367 -1308
rect 443 -1371 444 -1333
rect 520 -1371 521 -1333
rect 674 -1334 675 -1308
rect 716 -1334 717 -1308
rect 786 -1371 787 -1333
rect 856 -1334 857 -1308
rect 877 -1371 878 -1333
rect 933 -1371 934 -1333
rect 947 -1334 948 -1308
rect 79 -1336 80 -1308
rect 359 -1371 360 -1335
rect 366 -1371 367 -1335
rect 401 -1371 402 -1335
rect 429 -1371 430 -1335
rect 450 -1336 451 -1308
rect 572 -1336 573 -1308
rect 674 -1371 675 -1335
rect 688 -1336 689 -1308
rect 716 -1371 717 -1335
rect 723 -1371 724 -1335
rect 849 -1336 850 -1308
rect 856 -1371 857 -1335
rect 1038 -1336 1039 -1308
rect 79 -1371 80 -1337
rect 184 -1338 185 -1308
rect 191 -1371 192 -1337
rect 205 -1338 206 -1308
rect 212 -1371 213 -1337
rect 278 -1371 279 -1337
rect 415 -1338 416 -1308
rect 450 -1371 451 -1337
rect 572 -1371 573 -1337
rect 730 -1338 731 -1308
rect 737 -1371 738 -1337
rect 772 -1338 773 -1308
rect 835 -1338 836 -1308
rect 849 -1371 850 -1337
rect 926 -1338 927 -1308
rect 947 -1371 948 -1337
rect 170 -1340 171 -1308
rect 240 -1371 241 -1339
rect 254 -1340 255 -1308
rect 303 -1371 304 -1339
rect 310 -1371 311 -1339
rect 730 -1371 731 -1339
rect 772 -1371 773 -1339
rect 926 -1371 927 -1339
rect 954 -1340 955 -1308
rect 163 -1342 164 -1308
rect 170 -1371 171 -1341
rect 177 -1342 178 -1308
rect 205 -1371 206 -1341
rect 254 -1371 255 -1341
rect 478 -1342 479 -1308
rect 583 -1371 584 -1341
rect 618 -1342 619 -1308
rect 646 -1342 647 -1308
rect 688 -1371 689 -1341
rect 954 -1371 955 -1341
rect 989 -1342 990 -1308
rect 107 -1344 108 -1308
rect 163 -1371 164 -1343
rect 177 -1371 178 -1343
rect 415 -1371 416 -1343
rect 436 -1344 437 -1308
rect 464 -1371 465 -1343
rect 478 -1371 479 -1343
rect 548 -1344 549 -1308
rect 618 -1371 619 -1343
rect 639 -1344 640 -1308
rect 646 -1371 647 -1343
rect 940 -1371 941 -1343
rect 107 -1371 108 -1345
rect 135 -1371 136 -1345
rect 180 -1371 181 -1345
rect 226 -1346 227 -1308
rect 275 -1371 276 -1345
rect 562 -1346 563 -1308
rect 660 -1371 661 -1345
rect 779 -1346 780 -1308
rect 898 -1346 899 -1308
rect 989 -1371 990 -1345
rect 65 -1371 66 -1347
rect 562 -1371 563 -1347
rect 779 -1371 780 -1347
rect 800 -1348 801 -1308
rect 184 -1371 185 -1349
rect 198 -1350 199 -1308
rect 226 -1371 227 -1349
rect 233 -1350 234 -1308
rect 394 -1350 395 -1308
rect 898 -1371 899 -1349
rect 194 -1352 195 -1308
rect 219 -1352 220 -1308
rect 233 -1371 234 -1351
rect 317 -1352 318 -1308
rect 373 -1352 374 -1308
rect 394 -1371 395 -1351
rect 436 -1371 437 -1351
rect 457 -1352 458 -1308
rect 467 -1352 468 -1308
rect 639 -1371 640 -1351
rect 800 -1371 801 -1351
rect 807 -1352 808 -1308
rect 121 -1354 122 -1308
rect 219 -1371 220 -1353
rect 341 -1354 342 -1308
rect 457 -1371 458 -1353
rect 548 -1371 549 -1353
rect 796 -1354 797 -1308
rect 807 -1371 808 -1353
rect 814 -1354 815 -1308
rect 121 -1371 122 -1355
rect 149 -1356 150 -1308
rect 198 -1371 199 -1355
rect 324 -1356 325 -1308
rect 373 -1371 374 -1355
rect 541 -1371 542 -1355
rect 814 -1371 815 -1355
rect 828 -1356 829 -1308
rect 142 -1358 143 -1308
rect 317 -1371 318 -1357
rect 439 -1371 440 -1357
rect 576 -1371 577 -1357
rect 828 -1371 829 -1357
rect 842 -1358 843 -1308
rect 142 -1371 143 -1359
rect 835 -1371 836 -1359
rect 149 -1371 150 -1361
rect 156 -1362 157 -1308
rect 282 -1362 283 -1308
rect 324 -1371 325 -1361
rect 635 -1362 636 -1308
rect 842 -1371 843 -1361
rect 156 -1371 157 -1363
rect 387 -1364 388 -1308
rect 331 -1366 332 -1308
rect 387 -1371 388 -1365
rect 289 -1368 290 -1308
rect 331 -1371 332 -1367
rect 289 -1371 290 -1369
rect 404 -1370 405 -1308
rect 2 -1381 3 -1379
rect 5 -1446 6 -1380
rect 9 -1446 10 -1380
rect 114 -1381 115 -1379
rect 142 -1381 143 -1379
rect 240 -1381 241 -1379
rect 250 -1381 251 -1379
rect 268 -1381 269 -1379
rect 369 -1381 370 -1379
rect 674 -1381 675 -1379
rect 702 -1381 703 -1379
rect 730 -1446 731 -1380
rect 737 -1381 738 -1379
rect 737 -1446 738 -1380
rect 737 -1381 738 -1379
rect 737 -1446 738 -1380
rect 849 -1381 850 -1379
rect 849 -1446 850 -1380
rect 849 -1381 850 -1379
rect 849 -1446 850 -1380
rect 996 -1381 997 -1379
rect 1059 -1446 1060 -1380
rect 30 -1383 31 -1379
rect 33 -1387 34 -1382
rect 72 -1383 73 -1379
rect 275 -1383 276 -1379
rect 369 -1446 370 -1382
rect 520 -1383 521 -1379
rect 530 -1446 531 -1382
rect 786 -1383 787 -1379
rect 947 -1383 948 -1379
rect 996 -1446 997 -1382
rect 1003 -1383 1004 -1379
rect 1024 -1446 1025 -1382
rect 1031 -1383 1032 -1379
rect 1038 -1446 1039 -1382
rect 1045 -1446 1046 -1382
rect 1066 -1383 1067 -1379
rect 30 -1446 31 -1384
rect 44 -1385 45 -1379
rect 72 -1446 73 -1384
rect 201 -1385 202 -1379
rect 208 -1446 209 -1384
rect 590 -1385 591 -1379
rect 611 -1385 612 -1379
rect 611 -1446 612 -1384
rect 611 -1385 612 -1379
rect 611 -1446 612 -1384
rect 618 -1385 619 -1379
rect 625 -1446 626 -1384
rect 632 -1385 633 -1379
rect 674 -1446 675 -1384
rect 681 -1385 682 -1379
rect 947 -1446 948 -1384
rect 975 -1385 976 -1379
rect 1003 -1446 1004 -1384
rect 1010 -1385 1011 -1379
rect 1031 -1446 1032 -1384
rect 1055 -1446 1056 -1384
rect 1066 -1446 1067 -1384
rect 44 -1446 45 -1386
rect 79 -1387 80 -1379
rect 268 -1446 269 -1386
rect 380 -1387 381 -1379
rect 436 -1387 437 -1379
rect 443 -1387 444 -1379
rect 478 -1446 479 -1386
rect 488 -1446 489 -1386
rect 506 -1446 507 -1386
rect 509 -1387 510 -1379
rect 562 -1387 563 -1379
rect 646 -1387 647 -1379
rect 758 -1387 759 -1379
rect 786 -1446 787 -1386
rect 814 -1387 815 -1379
rect 940 -1387 941 -1379
rect 975 -1446 976 -1386
rect 982 -1387 983 -1379
rect 1010 -1446 1011 -1386
rect 79 -1446 80 -1388
rect 121 -1389 122 -1379
rect 128 -1389 129 -1379
rect 436 -1446 437 -1388
rect 457 -1389 458 -1379
rect 492 -1389 493 -1379
rect 499 -1389 500 -1379
rect 544 -1389 545 -1379
rect 555 -1389 556 -1379
rect 618 -1446 619 -1388
rect 653 -1389 654 -1379
rect 989 -1389 990 -1379
rect 86 -1391 87 -1379
rect 474 -1446 475 -1390
rect 513 -1391 514 -1379
rect 562 -1446 563 -1390
rect 569 -1391 570 -1379
rect 940 -1446 941 -1390
rect 961 -1391 962 -1379
rect 989 -1446 990 -1390
rect 86 -1446 87 -1392
rect 345 -1393 346 -1379
rect 366 -1393 367 -1379
rect 653 -1446 654 -1392
rect 660 -1446 661 -1392
rect 793 -1393 794 -1379
rect 912 -1393 913 -1379
rect 961 -1446 962 -1392
rect 100 -1446 101 -1394
rect 107 -1395 108 -1379
rect 114 -1446 115 -1394
rect 156 -1395 157 -1379
rect 177 -1446 178 -1394
rect 191 -1395 192 -1379
rect 198 -1446 199 -1394
rect 247 -1395 248 -1379
rect 261 -1395 262 -1379
rect 285 -1395 286 -1379
rect 289 -1395 290 -1379
rect 982 -1446 983 -1394
rect 93 -1397 94 -1379
rect 289 -1446 290 -1396
rect 380 -1446 381 -1396
rect 401 -1397 402 -1379
rect 408 -1397 409 -1379
rect 492 -1446 493 -1396
rect 534 -1397 535 -1379
rect 590 -1446 591 -1396
rect 604 -1397 605 -1379
rect 646 -1446 647 -1396
rect 667 -1397 668 -1379
rect 681 -1446 682 -1396
rect 702 -1446 703 -1396
rect 772 -1397 773 -1379
rect 793 -1446 794 -1396
rect 814 -1446 815 -1396
rect 912 -1446 913 -1396
rect 926 -1397 927 -1379
rect 16 -1399 17 -1379
rect 93 -1446 94 -1398
rect 121 -1446 122 -1398
rect 523 -1446 524 -1398
rect 537 -1446 538 -1398
rect 821 -1399 822 -1379
rect 842 -1399 843 -1379
rect 926 -1446 927 -1398
rect 128 -1446 129 -1400
rect 898 -1401 899 -1379
rect 142 -1446 143 -1402
rect 170 -1403 171 -1379
rect 212 -1403 213 -1379
rect 401 -1446 402 -1402
rect 408 -1446 409 -1402
rect 656 -1403 657 -1379
rect 667 -1446 668 -1402
rect 751 -1403 752 -1379
rect 772 -1446 773 -1402
rect 800 -1403 801 -1379
rect 821 -1446 822 -1402
rect 919 -1403 920 -1379
rect 58 -1405 59 -1379
rect 170 -1446 171 -1404
rect 219 -1405 220 -1379
rect 261 -1446 262 -1404
rect 345 -1446 346 -1404
rect 534 -1446 535 -1404
rect 541 -1405 542 -1379
rect 968 -1405 969 -1379
rect 149 -1407 150 -1379
rect 149 -1446 150 -1406
rect 149 -1407 150 -1379
rect 149 -1446 150 -1406
rect 156 -1446 157 -1406
rect 548 -1407 549 -1379
rect 569 -1446 570 -1406
rect 723 -1407 724 -1379
rect 726 -1407 727 -1379
rect 933 -1407 934 -1379
rect 135 -1446 136 -1408
rect 548 -1446 549 -1408
rect 663 -1409 664 -1379
rect 968 -1446 969 -1408
rect 205 -1411 206 -1379
rect 219 -1446 220 -1410
rect 226 -1411 227 -1379
rect 376 -1446 377 -1410
rect 394 -1411 395 -1379
rect 394 -1446 395 -1410
rect 394 -1411 395 -1379
rect 394 -1446 395 -1410
rect 415 -1411 416 -1379
rect 443 -1446 444 -1410
rect 450 -1411 451 -1379
rect 499 -1446 500 -1410
rect 541 -1446 542 -1410
rect 744 -1411 745 -1379
rect 751 -1446 752 -1410
rect 765 -1411 766 -1379
rect 828 -1411 829 -1379
rect 842 -1446 843 -1410
rect 891 -1411 892 -1379
rect 898 -1446 899 -1410
rect 905 -1411 906 -1379
rect 919 -1446 920 -1410
rect 107 -1446 108 -1412
rect 205 -1446 206 -1412
rect 226 -1446 227 -1412
rect 254 -1413 255 -1379
rect 366 -1446 367 -1412
rect 933 -1446 934 -1412
rect 233 -1415 234 -1379
rect 1052 -1446 1053 -1414
rect 51 -1417 52 -1379
rect 233 -1446 234 -1416
rect 240 -1446 241 -1416
rect 338 -1417 339 -1379
rect 415 -1446 416 -1416
rect 422 -1417 423 -1379
rect 429 -1417 430 -1379
rect 429 -1446 430 -1416
rect 429 -1417 430 -1379
rect 429 -1446 430 -1416
rect 439 -1446 440 -1416
rect 555 -1446 556 -1416
rect 597 -1417 598 -1379
rect 744 -1446 745 -1416
rect 796 -1446 797 -1416
rect 905 -1446 906 -1416
rect 51 -1446 52 -1418
rect 387 -1419 388 -1379
rect 450 -1446 451 -1418
rect 807 -1419 808 -1379
rect 828 -1446 829 -1418
rect 884 -1419 885 -1379
rect 58 -1446 59 -1420
rect 422 -1446 423 -1420
rect 471 -1421 472 -1379
rect 513 -1446 514 -1420
rect 520 -1446 521 -1420
rect 597 -1446 598 -1420
rect 695 -1421 696 -1379
rect 723 -1446 724 -1420
rect 779 -1421 780 -1379
rect 807 -1446 808 -1420
rect 877 -1421 878 -1379
rect 884 -1446 885 -1420
rect 247 -1446 248 -1422
rect 303 -1423 304 -1379
rect 310 -1423 311 -1379
rect 338 -1446 339 -1422
rect 387 -1446 388 -1422
rect 527 -1423 528 -1379
rect 688 -1423 689 -1379
rect 695 -1446 696 -1422
rect 709 -1423 710 -1379
rect 800 -1446 801 -1422
rect 870 -1423 871 -1379
rect 877 -1446 878 -1422
rect 254 -1446 255 -1424
rect 485 -1425 486 -1379
rect 527 -1446 528 -1424
rect 835 -1425 836 -1379
rect 863 -1425 864 -1379
rect 870 -1446 871 -1424
rect 138 -1427 139 -1379
rect 863 -1446 864 -1426
rect 303 -1446 304 -1428
rect 317 -1429 318 -1379
rect 348 -1429 349 -1379
rect 835 -1446 836 -1428
rect 310 -1446 311 -1430
rect 331 -1431 332 -1379
rect 464 -1431 465 -1379
rect 485 -1446 486 -1430
rect 628 -1431 629 -1379
rect 709 -1446 710 -1430
rect 716 -1431 717 -1379
rect 758 -1446 759 -1430
rect 779 -1446 780 -1430
rect 856 -1431 857 -1379
rect 331 -1446 332 -1432
rect 352 -1433 353 -1379
rect 359 -1433 360 -1379
rect 464 -1446 465 -1432
rect 576 -1433 577 -1379
rect 856 -1446 857 -1432
rect 23 -1435 24 -1379
rect 352 -1446 353 -1434
rect 460 -1446 461 -1434
rect 716 -1446 717 -1434
rect 23 -1446 24 -1436
rect 163 -1437 164 -1379
rect 324 -1437 325 -1379
rect 359 -1446 360 -1436
rect 576 -1446 577 -1436
rect 583 -1437 584 -1379
rect 639 -1437 640 -1379
rect 688 -1446 689 -1436
rect 163 -1446 164 -1438
rect 184 -1439 185 -1379
rect 296 -1439 297 -1379
rect 324 -1446 325 -1438
rect 583 -1446 584 -1438
rect 1048 -1446 1049 -1438
rect 37 -1441 38 -1379
rect 184 -1446 185 -1440
rect 296 -1446 297 -1440
rect 373 -1441 374 -1379
rect 639 -1446 640 -1440
rect 1017 -1441 1018 -1379
rect 373 -1446 374 -1442
rect 891 -1446 892 -1442
rect 954 -1443 955 -1379
rect 1017 -1446 1018 -1442
rect 495 -1445 496 -1379
rect 954 -1446 955 -1444
rect 2 -1529 3 -1455
rect 37 -1456 38 -1454
rect 68 -1456 69 -1454
rect 394 -1456 395 -1454
rect 415 -1456 416 -1454
rect 415 -1529 416 -1455
rect 415 -1456 416 -1454
rect 415 -1529 416 -1455
rect 422 -1456 423 -1454
rect 814 -1456 815 -1454
rect 824 -1456 825 -1454
rect 1024 -1456 1025 -1454
rect 1045 -1529 1046 -1455
rect 1059 -1456 1060 -1454
rect 9 -1458 10 -1454
rect 128 -1458 129 -1454
rect 142 -1458 143 -1454
rect 285 -1458 286 -1454
rect 310 -1458 311 -1454
rect 317 -1529 318 -1457
rect 348 -1529 349 -1457
rect 443 -1458 444 -1454
rect 457 -1458 458 -1454
rect 982 -1458 983 -1454
rect 999 -1529 1000 -1457
rect 1038 -1458 1039 -1454
rect 1048 -1458 1049 -1454
rect 1052 -1529 1053 -1457
rect 1059 -1529 1060 -1457
rect 1066 -1458 1067 -1454
rect 19 -1460 20 -1454
rect 58 -1460 59 -1454
rect 72 -1460 73 -1454
rect 138 -1460 139 -1454
rect 142 -1529 143 -1459
rect 177 -1460 178 -1454
rect 184 -1460 185 -1454
rect 310 -1529 311 -1459
rect 352 -1460 353 -1454
rect 460 -1460 461 -1454
rect 506 -1460 507 -1454
rect 537 -1460 538 -1454
rect 593 -1529 594 -1459
rect 845 -1529 846 -1459
rect 982 -1529 983 -1459
rect 1031 -1460 1032 -1454
rect 23 -1462 24 -1454
rect 352 -1529 353 -1461
rect 387 -1462 388 -1454
rect 474 -1462 475 -1454
rect 509 -1529 510 -1461
rect 618 -1462 619 -1454
rect 625 -1462 626 -1454
rect 628 -1504 629 -1461
rect 632 -1529 633 -1461
rect 681 -1462 682 -1454
rect 684 -1529 685 -1461
rect 933 -1462 934 -1454
rect 23 -1529 24 -1463
rect 425 -1464 426 -1454
rect 429 -1464 430 -1454
rect 429 -1529 430 -1463
rect 429 -1464 430 -1454
rect 429 -1529 430 -1463
rect 436 -1464 437 -1454
rect 968 -1464 969 -1454
rect 30 -1466 31 -1454
rect 40 -1466 41 -1454
rect 72 -1529 73 -1465
rect 562 -1466 563 -1454
rect 604 -1529 605 -1465
rect 611 -1466 612 -1454
rect 625 -1529 626 -1465
rect 744 -1466 745 -1454
rect 747 -1466 748 -1454
rect 751 -1466 752 -1454
rect 751 -1529 752 -1465
rect 751 -1466 752 -1454
rect 751 -1529 752 -1465
rect 765 -1466 766 -1454
rect 863 -1466 864 -1454
rect 37 -1529 38 -1467
rect 44 -1468 45 -1454
rect 93 -1468 94 -1454
rect 422 -1529 423 -1467
rect 436 -1529 437 -1467
rect 464 -1468 465 -1454
rect 520 -1468 521 -1454
rect 758 -1468 759 -1454
rect 765 -1529 766 -1467
rect 870 -1468 871 -1454
rect 44 -1529 45 -1469
rect 408 -1470 409 -1454
rect 443 -1529 444 -1469
rect 569 -1470 570 -1454
rect 607 -1470 608 -1454
rect 947 -1470 948 -1454
rect 58 -1529 59 -1471
rect 408 -1529 409 -1471
rect 450 -1472 451 -1454
rect 537 -1529 538 -1471
rect 611 -1529 612 -1471
rect 674 -1472 675 -1454
rect 681 -1529 682 -1471
rect 926 -1472 927 -1454
rect 93 -1529 94 -1473
rect 177 -1529 178 -1473
rect 191 -1474 192 -1454
rect 478 -1474 479 -1454
rect 520 -1529 521 -1473
rect 940 -1474 941 -1454
rect 96 -1529 97 -1475
rect 758 -1529 759 -1475
rect 768 -1476 769 -1454
rect 828 -1476 829 -1454
rect 856 -1476 857 -1454
rect 870 -1529 871 -1475
rect 926 -1529 927 -1475
rect 975 -1476 976 -1454
rect 100 -1478 101 -1454
rect 100 -1529 101 -1477
rect 100 -1478 101 -1454
rect 100 -1529 101 -1477
rect 128 -1529 129 -1477
rect 303 -1478 304 -1454
rect 345 -1478 346 -1454
rect 450 -1529 451 -1477
rect 464 -1529 465 -1477
rect 513 -1478 514 -1454
rect 534 -1529 535 -1477
rect 548 -1478 549 -1454
rect 635 -1478 636 -1454
rect 660 -1478 661 -1454
rect 667 -1478 668 -1454
rect 674 -1529 675 -1477
rect 709 -1478 710 -1454
rect 947 -1529 948 -1477
rect 975 -1529 976 -1477
rect 996 -1478 997 -1454
rect 149 -1480 150 -1454
rect 149 -1529 150 -1479
rect 149 -1480 150 -1454
rect 149 -1529 150 -1479
rect 163 -1480 164 -1454
rect 184 -1529 185 -1479
rect 191 -1529 192 -1479
rect 240 -1480 241 -1454
rect 247 -1480 248 -1454
rect 376 -1480 377 -1454
rect 387 -1529 388 -1479
rect 653 -1480 654 -1454
rect 660 -1529 661 -1479
rect 667 -1529 668 -1479
rect 709 -1529 710 -1479
rect 737 -1480 738 -1454
rect 744 -1529 745 -1479
rect 779 -1480 780 -1454
rect 786 -1480 787 -1454
rect 786 -1529 787 -1479
rect 786 -1480 787 -1454
rect 786 -1529 787 -1479
rect 793 -1480 794 -1454
rect 961 -1480 962 -1454
rect 163 -1529 164 -1481
rect 198 -1482 199 -1454
rect 215 -1482 216 -1454
rect 569 -1529 570 -1481
rect 639 -1482 640 -1454
rect 702 -1482 703 -1454
rect 772 -1482 773 -1454
rect 779 -1529 780 -1481
rect 793 -1529 794 -1481
rect 842 -1482 843 -1454
rect 856 -1529 857 -1481
rect 898 -1482 899 -1454
rect 170 -1484 171 -1454
rect 205 -1529 206 -1483
rect 219 -1484 220 -1454
rect 219 -1529 220 -1483
rect 219 -1484 220 -1454
rect 219 -1529 220 -1483
rect 226 -1484 227 -1454
rect 247 -1529 248 -1483
rect 261 -1484 262 -1454
rect 261 -1529 262 -1483
rect 261 -1484 262 -1454
rect 261 -1529 262 -1483
rect 268 -1484 269 -1454
rect 275 -1484 276 -1454
rect 282 -1529 283 -1483
rect 324 -1484 325 -1454
rect 373 -1484 374 -1454
rect 940 -1529 941 -1483
rect 107 -1486 108 -1454
rect 226 -1529 227 -1485
rect 233 -1486 234 -1454
rect 324 -1529 325 -1485
rect 373 -1529 374 -1485
rect 488 -1486 489 -1454
rect 544 -1529 545 -1485
rect 961 -1529 962 -1485
rect 107 -1529 108 -1487
rect 527 -1488 528 -1454
rect 548 -1529 549 -1487
rect 576 -1488 577 -1454
rect 639 -1529 640 -1487
rect 695 -1488 696 -1454
rect 702 -1529 703 -1487
rect 726 -1529 727 -1487
rect 772 -1529 773 -1487
rect 807 -1488 808 -1454
rect 814 -1529 815 -1487
rect 884 -1488 885 -1454
rect 898 -1529 899 -1487
rect 919 -1488 920 -1454
rect 68 -1529 69 -1489
rect 884 -1529 885 -1489
rect 114 -1492 115 -1454
rect 268 -1529 269 -1491
rect 275 -1529 276 -1491
rect 359 -1492 360 -1454
rect 394 -1529 395 -1491
rect 555 -1492 556 -1454
rect 642 -1492 643 -1454
rect 863 -1529 864 -1491
rect 79 -1494 80 -1454
rect 114 -1529 115 -1493
rect 121 -1494 122 -1454
rect 170 -1529 171 -1493
rect 194 -1494 195 -1454
rect 212 -1529 213 -1493
rect 233 -1529 234 -1493
rect 331 -1494 332 -1454
rect 359 -1529 360 -1493
rect 401 -1494 402 -1454
rect 478 -1529 479 -1493
rect 597 -1494 598 -1454
rect 653 -1529 654 -1493
rect 688 -1494 689 -1454
rect 695 -1529 696 -1493
rect 740 -1529 741 -1493
rect 796 -1494 797 -1454
rect 828 -1529 829 -1493
rect 842 -1529 843 -1493
rect 1017 -1494 1018 -1454
rect 51 -1496 52 -1454
rect 121 -1529 122 -1495
rect 240 -1529 241 -1495
rect 523 -1529 524 -1495
rect 541 -1496 542 -1454
rect 576 -1529 577 -1495
rect 590 -1496 591 -1454
rect 597 -1529 598 -1495
rect 807 -1529 808 -1495
rect 877 -1496 878 -1454
rect 989 -1496 990 -1454
rect 1017 -1529 1018 -1495
rect 51 -1529 52 -1497
rect 254 -1498 255 -1454
rect 296 -1498 297 -1454
rect 401 -1529 402 -1497
rect 492 -1498 493 -1454
rect 919 -1529 920 -1497
rect 79 -1529 80 -1499
rect 156 -1500 157 -1454
rect 254 -1529 255 -1499
rect 583 -1500 584 -1454
rect 590 -1529 591 -1499
rect 835 -1500 836 -1454
rect 877 -1529 878 -1499
rect 1003 -1500 1004 -1454
rect 86 -1502 87 -1454
rect 156 -1529 157 -1501
rect 278 -1502 279 -1454
rect 492 -1529 493 -1501
rect 506 -1529 507 -1501
rect 835 -1529 836 -1501
rect 905 -1502 906 -1454
rect 989 -1529 990 -1501
rect 86 -1529 87 -1503
rect 135 -1504 136 -1454
rect 296 -1529 297 -1503
rect 457 -1529 458 -1503
rect 516 -1529 517 -1503
rect 688 -1529 689 -1503
rect 747 -1529 748 -1503
rect 1003 -1529 1004 -1503
rect 16 -1529 17 -1505
rect 135 -1529 136 -1505
rect 303 -1529 304 -1505
rect 380 -1506 381 -1454
rect 541 -1529 542 -1505
rect 933 -1529 934 -1505
rect 331 -1529 332 -1507
rect 488 -1529 489 -1507
rect 555 -1529 556 -1507
rect 565 -1529 566 -1507
rect 583 -1529 584 -1507
rect 646 -1508 647 -1454
rect 821 -1529 822 -1507
rect 996 -1529 997 -1507
rect 338 -1510 339 -1454
rect 380 -1529 381 -1509
rect 646 -1529 647 -1509
rect 730 -1510 731 -1454
rect 905 -1529 906 -1509
rect 912 -1510 913 -1454
rect 338 -1529 339 -1511
rect 366 -1512 367 -1454
rect 499 -1512 500 -1454
rect 730 -1529 731 -1511
rect 912 -1529 913 -1511
rect 954 -1512 955 -1454
rect 198 -1529 199 -1513
rect 499 -1529 500 -1513
rect 954 -1529 955 -1513
rect 1010 -1514 1011 -1454
rect 366 -1529 367 -1515
rect 723 -1516 724 -1454
rect 800 -1516 801 -1454
rect 1010 -1529 1011 -1515
rect 723 -1529 724 -1517
rect 968 -1529 969 -1517
rect 800 -1529 801 -1519
rect 849 -1520 850 -1454
rect 849 -1529 850 -1521
rect 891 -1522 892 -1454
rect 471 -1524 472 -1454
rect 891 -1529 892 -1523
rect 289 -1526 290 -1454
rect 471 -1529 472 -1525
rect 30 -1529 31 -1527
rect 289 -1529 290 -1527
rect 23 -1539 24 -1537
rect 135 -1539 136 -1537
rect 152 -1606 153 -1538
rect 961 -1539 962 -1537
rect 1017 -1539 1018 -1537
rect 1024 -1606 1025 -1538
rect 1038 -1606 1039 -1538
rect 1045 -1539 1046 -1537
rect 1052 -1539 1053 -1537
rect 1052 -1606 1053 -1538
rect 1052 -1539 1053 -1537
rect 1052 -1606 1053 -1538
rect 2 -1541 3 -1537
rect 23 -1606 24 -1540
rect 30 -1541 31 -1537
rect 425 -1606 426 -1540
rect 436 -1541 437 -1537
rect 436 -1606 437 -1540
rect 436 -1541 437 -1537
rect 436 -1606 437 -1540
rect 471 -1541 472 -1537
rect 471 -1606 472 -1540
rect 471 -1541 472 -1537
rect 471 -1606 472 -1540
rect 488 -1541 489 -1537
rect 737 -1541 738 -1537
rect 740 -1541 741 -1537
rect 982 -1541 983 -1537
rect 30 -1606 31 -1542
rect 303 -1543 304 -1537
rect 306 -1606 307 -1542
rect 506 -1606 507 -1542
rect 520 -1543 521 -1537
rect 919 -1543 920 -1537
rect 961 -1606 962 -1542
rect 996 -1543 997 -1537
rect 37 -1545 38 -1537
rect 37 -1606 38 -1544
rect 37 -1545 38 -1537
rect 37 -1606 38 -1544
rect 68 -1545 69 -1537
rect 86 -1545 87 -1537
rect 93 -1606 94 -1544
rect 415 -1545 416 -1537
rect 527 -1545 528 -1537
rect 548 -1545 549 -1537
rect 558 -1606 559 -1544
rect 975 -1545 976 -1537
rect 68 -1606 69 -1546
rect 758 -1547 759 -1537
rect 842 -1606 843 -1546
rect 884 -1547 885 -1537
rect 79 -1549 80 -1537
rect 79 -1606 80 -1548
rect 79 -1549 80 -1537
rect 79 -1606 80 -1548
rect 86 -1606 87 -1548
rect 100 -1549 101 -1537
rect 135 -1606 136 -1548
rect 261 -1549 262 -1537
rect 289 -1549 290 -1537
rect 667 -1549 668 -1537
rect 723 -1606 724 -1548
rect 814 -1549 815 -1537
rect 877 -1549 878 -1537
rect 919 -1606 920 -1548
rect 100 -1606 101 -1550
rect 226 -1551 227 -1537
rect 247 -1551 248 -1537
rect 261 -1606 262 -1550
rect 296 -1551 297 -1537
rect 359 -1551 360 -1537
rect 366 -1551 367 -1537
rect 628 -1606 629 -1550
rect 646 -1551 647 -1537
rect 646 -1606 647 -1550
rect 646 -1551 647 -1537
rect 646 -1606 647 -1550
rect 663 -1551 664 -1537
rect 828 -1551 829 -1537
rect 884 -1606 885 -1550
rect 1003 -1551 1004 -1537
rect 128 -1553 129 -1537
rect 289 -1606 290 -1552
rect 324 -1553 325 -1537
rect 324 -1606 325 -1552
rect 324 -1553 325 -1537
rect 324 -1606 325 -1552
rect 373 -1553 374 -1537
rect 485 -1606 486 -1552
rect 499 -1553 500 -1537
rect 548 -1606 549 -1552
rect 565 -1553 566 -1537
rect 947 -1553 948 -1537
rect 72 -1555 73 -1537
rect 499 -1606 500 -1554
rect 534 -1606 535 -1554
rect 555 -1555 556 -1537
rect 583 -1555 584 -1537
rect 667 -1606 668 -1554
rect 684 -1555 685 -1537
rect 877 -1606 878 -1554
rect 947 -1606 948 -1554
rect 1010 -1555 1011 -1537
rect 16 -1557 17 -1537
rect 72 -1606 73 -1556
rect 121 -1557 122 -1537
rect 128 -1606 129 -1556
rect 156 -1557 157 -1537
rect 313 -1606 314 -1556
rect 359 -1606 360 -1556
rect 565 -1606 566 -1556
rect 583 -1606 584 -1556
rect 695 -1557 696 -1537
rect 726 -1557 727 -1537
rect 898 -1557 899 -1537
rect 121 -1606 122 -1558
rect 275 -1559 276 -1537
rect 366 -1606 367 -1558
rect 555 -1606 556 -1558
rect 590 -1559 591 -1537
rect 828 -1606 829 -1558
rect 898 -1606 899 -1558
rect 933 -1559 934 -1537
rect 44 -1561 45 -1537
rect 275 -1606 276 -1560
rect 373 -1606 374 -1560
rect 537 -1561 538 -1537
rect 541 -1606 542 -1560
rect 611 -1561 612 -1537
rect 618 -1561 619 -1537
rect 653 -1561 654 -1537
rect 737 -1606 738 -1560
rect 821 -1561 822 -1537
rect 44 -1606 45 -1562
rect 142 -1563 143 -1537
rect 156 -1606 157 -1562
rect 338 -1563 339 -1537
rect 355 -1563 356 -1537
rect 653 -1606 654 -1562
rect 758 -1606 759 -1562
rect 800 -1563 801 -1537
rect 814 -1606 815 -1562
rect 863 -1563 864 -1537
rect 107 -1565 108 -1537
rect 338 -1606 339 -1564
rect 380 -1565 381 -1537
rect 415 -1606 416 -1564
rect 590 -1606 591 -1564
rect 639 -1565 640 -1537
rect 800 -1606 801 -1564
rect 807 -1565 808 -1537
rect 821 -1606 822 -1564
rect 849 -1565 850 -1537
rect 863 -1606 864 -1564
rect 912 -1565 913 -1537
rect 142 -1606 143 -1566
rect 149 -1567 150 -1537
rect 170 -1567 171 -1537
rect 695 -1606 696 -1566
rect 807 -1606 808 -1566
rect 870 -1567 871 -1537
rect 912 -1606 913 -1566
rect 989 -1567 990 -1537
rect 177 -1569 178 -1537
rect 380 -1606 381 -1568
rect 387 -1569 388 -1537
rect 513 -1569 514 -1537
rect 576 -1569 577 -1537
rect 639 -1606 640 -1568
rect 660 -1569 661 -1537
rect 849 -1606 850 -1568
rect 870 -1606 871 -1568
rect 926 -1569 927 -1537
rect 177 -1606 178 -1570
rect 191 -1571 192 -1537
rect 201 -1571 202 -1537
rect 310 -1571 311 -1537
rect 401 -1571 402 -1537
rect 464 -1606 465 -1570
rect 478 -1571 479 -1537
rect 513 -1606 514 -1570
rect 562 -1606 563 -1570
rect 926 -1606 927 -1570
rect 184 -1573 185 -1537
rect 184 -1606 185 -1572
rect 184 -1573 185 -1537
rect 184 -1606 185 -1572
rect 191 -1606 192 -1572
rect 205 -1573 206 -1537
rect 212 -1573 213 -1537
rect 296 -1606 297 -1572
rect 394 -1573 395 -1537
rect 478 -1606 479 -1572
rect 576 -1606 577 -1572
rect 632 -1573 633 -1537
rect 660 -1606 661 -1572
rect 688 -1573 689 -1537
rect 205 -1606 206 -1574
rect 233 -1575 234 -1537
rect 240 -1575 241 -1537
rect 355 -1606 356 -1574
rect 401 -1606 402 -1574
rect 429 -1575 430 -1537
rect 569 -1575 570 -1537
rect 632 -1606 633 -1574
rect 688 -1606 689 -1574
rect 709 -1575 710 -1537
rect 163 -1577 164 -1537
rect 233 -1606 234 -1576
rect 240 -1606 241 -1576
rect 422 -1577 423 -1537
rect 429 -1606 430 -1576
rect 457 -1577 458 -1537
rect 604 -1606 605 -1576
rect 625 -1577 626 -1537
rect 709 -1606 710 -1576
rect 744 -1577 745 -1537
rect 58 -1579 59 -1537
rect 163 -1606 164 -1578
rect 212 -1606 213 -1578
rect 219 -1579 220 -1537
rect 247 -1606 248 -1578
rect 282 -1579 283 -1537
rect 345 -1606 346 -1578
rect 394 -1606 395 -1578
rect 408 -1579 409 -1537
rect 702 -1579 703 -1537
rect 744 -1606 745 -1578
rect 779 -1579 780 -1537
rect 58 -1606 59 -1580
rect 173 -1606 174 -1580
rect 408 -1606 409 -1580
rect 443 -1581 444 -1537
rect 450 -1581 451 -1537
rect 457 -1606 458 -1580
rect 597 -1581 598 -1537
rect 779 -1606 780 -1580
rect 51 -1583 52 -1537
rect 450 -1606 451 -1582
rect 618 -1606 619 -1582
rect 674 -1583 675 -1537
rect 702 -1606 703 -1582
rect 940 -1583 941 -1537
rect 51 -1606 52 -1584
rect 572 -1606 573 -1584
rect 716 -1585 717 -1537
rect 940 -1606 941 -1584
rect 114 -1587 115 -1537
rect 219 -1606 220 -1586
rect 387 -1606 388 -1586
rect 597 -1606 598 -1586
rect 716 -1606 717 -1586
rect 751 -1587 752 -1537
rect 107 -1606 108 -1588
rect 114 -1606 115 -1588
rect 117 -1589 118 -1537
rect 282 -1606 283 -1588
rect 411 -1589 412 -1537
rect 730 -1589 731 -1537
rect 751 -1606 752 -1588
rect 786 -1589 787 -1537
rect 443 -1606 444 -1590
rect 530 -1606 531 -1590
rect 730 -1606 731 -1590
rect 772 -1591 773 -1537
rect 786 -1606 787 -1590
rect 856 -1591 857 -1537
rect 492 -1593 493 -1537
rect 674 -1606 675 -1592
rect 765 -1593 766 -1537
rect 772 -1606 773 -1592
rect 856 -1606 857 -1592
rect 936 -1606 937 -1592
rect 331 -1595 332 -1537
rect 492 -1606 493 -1594
rect 765 -1606 766 -1594
rect 793 -1595 794 -1537
rect 317 -1597 318 -1537
rect 331 -1606 332 -1596
rect 793 -1606 794 -1596
rect 835 -1597 836 -1537
rect 268 -1599 269 -1537
rect 317 -1606 318 -1598
rect 835 -1606 836 -1598
rect 891 -1599 892 -1537
rect 254 -1601 255 -1537
rect 268 -1606 269 -1600
rect 891 -1606 892 -1600
rect 954 -1601 955 -1537
rect 254 -1606 255 -1602
rect 509 -1603 510 -1537
rect 905 -1603 906 -1537
rect 954 -1606 955 -1602
rect 905 -1606 906 -1604
rect 968 -1605 969 -1537
rect 30 -1616 31 -1614
rect 355 -1616 356 -1614
rect 366 -1616 367 -1614
rect 527 -1671 528 -1615
rect 530 -1616 531 -1614
rect 779 -1616 780 -1614
rect 926 -1616 927 -1614
rect 936 -1616 937 -1614
rect 954 -1616 955 -1614
rect 968 -1671 969 -1615
rect 1024 -1616 1025 -1614
rect 1024 -1671 1025 -1615
rect 1024 -1616 1025 -1614
rect 1024 -1671 1025 -1615
rect 1038 -1616 1039 -1614
rect 1045 -1616 1046 -1614
rect 37 -1618 38 -1614
rect 37 -1671 38 -1617
rect 37 -1618 38 -1614
rect 37 -1671 38 -1617
rect 58 -1618 59 -1614
rect 303 -1618 304 -1614
rect 310 -1618 311 -1614
rect 471 -1618 472 -1614
rect 523 -1618 524 -1614
rect 667 -1618 668 -1614
rect 681 -1618 682 -1614
rect 737 -1618 738 -1614
rect 775 -1671 776 -1617
rect 849 -1618 850 -1614
rect 65 -1671 66 -1619
rect 110 -1620 111 -1614
rect 121 -1620 122 -1614
rect 306 -1620 307 -1614
rect 310 -1671 311 -1619
rect 352 -1620 353 -1614
rect 366 -1671 367 -1619
rect 401 -1620 402 -1614
rect 425 -1620 426 -1614
rect 471 -1671 472 -1619
rect 534 -1620 535 -1614
rect 534 -1671 535 -1619
rect 534 -1620 535 -1614
rect 534 -1671 535 -1619
rect 544 -1671 545 -1619
rect 793 -1620 794 -1614
rect 68 -1622 69 -1614
rect 240 -1622 241 -1614
rect 257 -1671 258 -1621
rect 324 -1622 325 -1614
rect 352 -1671 353 -1621
rect 408 -1622 409 -1614
rect 429 -1622 430 -1614
rect 516 -1671 517 -1621
rect 551 -1671 552 -1621
rect 639 -1622 640 -1614
rect 646 -1622 647 -1614
rect 667 -1671 668 -1621
rect 681 -1671 682 -1621
rect 684 -1622 685 -1614
rect 695 -1622 696 -1614
rect 919 -1622 920 -1614
rect 72 -1671 73 -1623
rect 411 -1671 412 -1623
rect 562 -1624 563 -1614
rect 838 -1671 839 -1623
rect 79 -1626 80 -1614
rect 401 -1671 402 -1625
rect 562 -1671 563 -1625
rect 702 -1626 703 -1614
rect 723 -1626 724 -1614
rect 737 -1671 738 -1625
rect 751 -1626 752 -1614
rect 793 -1671 794 -1625
rect 79 -1671 80 -1627
rect 229 -1628 230 -1614
rect 261 -1628 262 -1614
rect 261 -1671 262 -1627
rect 261 -1628 262 -1614
rect 261 -1671 262 -1627
rect 268 -1628 269 -1614
rect 422 -1628 423 -1614
rect 565 -1628 566 -1614
rect 618 -1628 619 -1614
rect 688 -1628 689 -1614
rect 751 -1671 752 -1627
rect 779 -1671 780 -1627
rect 821 -1628 822 -1614
rect 107 -1630 108 -1614
rect 513 -1630 514 -1614
rect 569 -1630 570 -1614
rect 814 -1630 815 -1614
rect 93 -1632 94 -1614
rect 107 -1671 108 -1631
rect 121 -1671 122 -1631
rect 159 -1632 160 -1614
rect 163 -1632 164 -1614
rect 240 -1671 241 -1631
rect 268 -1671 269 -1631
rect 404 -1671 405 -1631
rect 513 -1671 514 -1631
rect 859 -1632 860 -1614
rect 93 -1671 94 -1633
rect 254 -1634 255 -1614
rect 282 -1634 283 -1614
rect 523 -1671 524 -1633
rect 569 -1671 570 -1633
rect 632 -1634 633 -1614
rect 688 -1671 689 -1633
rect 870 -1634 871 -1614
rect 128 -1636 129 -1614
rect 163 -1671 164 -1635
rect 198 -1636 199 -1614
rect 345 -1636 346 -1614
rect 376 -1636 377 -1614
rect 380 -1636 381 -1614
rect 387 -1671 388 -1635
rect 443 -1636 444 -1614
rect 576 -1636 577 -1614
rect 632 -1671 633 -1635
rect 695 -1671 696 -1635
rect 803 -1671 804 -1635
rect 814 -1671 815 -1635
rect 940 -1636 941 -1614
rect 114 -1638 115 -1614
rect 128 -1671 129 -1637
rect 142 -1638 143 -1614
rect 142 -1671 143 -1637
rect 142 -1638 143 -1614
rect 142 -1671 143 -1637
rect 149 -1671 150 -1637
rect 170 -1638 171 -1614
rect 208 -1671 209 -1637
rect 422 -1671 423 -1637
rect 443 -1671 444 -1637
rect 464 -1638 465 -1614
rect 478 -1638 479 -1614
rect 576 -1671 577 -1637
rect 590 -1638 591 -1614
rect 625 -1671 626 -1637
rect 702 -1671 703 -1637
rect 765 -1638 766 -1614
rect 86 -1640 87 -1614
rect 114 -1671 115 -1639
rect 152 -1640 153 -1614
rect 247 -1640 248 -1614
rect 275 -1640 276 -1614
rect 282 -1671 283 -1639
rect 296 -1640 297 -1614
rect 432 -1671 433 -1639
rect 478 -1671 479 -1639
rect 499 -1640 500 -1614
rect 590 -1671 591 -1639
rect 660 -1640 661 -1614
rect 709 -1640 710 -1614
rect 765 -1671 766 -1639
rect 86 -1671 87 -1641
rect 205 -1642 206 -1614
rect 212 -1642 213 -1614
rect 226 -1642 227 -1614
rect 247 -1671 248 -1641
rect 289 -1642 290 -1614
rect 296 -1671 297 -1641
rect 331 -1642 332 -1614
rect 359 -1642 360 -1614
rect 380 -1671 381 -1641
rect 390 -1642 391 -1614
rect 492 -1642 493 -1614
rect 499 -1671 500 -1641
rect 520 -1671 521 -1641
rect 597 -1642 598 -1614
rect 597 -1671 598 -1641
rect 597 -1642 598 -1614
rect 597 -1671 598 -1641
rect 604 -1642 605 -1614
rect 646 -1671 647 -1641
rect 709 -1671 710 -1641
rect 744 -1642 745 -1614
rect 758 -1642 759 -1614
rect 821 -1671 822 -1641
rect 44 -1644 45 -1614
rect 205 -1671 206 -1643
rect 212 -1671 213 -1643
rect 219 -1644 220 -1614
rect 226 -1671 227 -1643
rect 233 -1644 234 -1614
rect 289 -1671 290 -1643
rect 436 -1644 437 -1614
rect 485 -1644 486 -1614
rect 492 -1671 493 -1643
rect 583 -1644 584 -1614
rect 604 -1671 605 -1643
rect 611 -1671 612 -1643
rect 653 -1644 654 -1614
rect 716 -1644 717 -1614
rect 723 -1671 724 -1643
rect 730 -1644 731 -1614
rect 758 -1671 759 -1643
rect 23 -1646 24 -1614
rect 44 -1671 45 -1645
rect 135 -1646 136 -1614
rect 233 -1671 234 -1645
rect 317 -1646 318 -1614
rect 345 -1671 346 -1645
rect 373 -1646 374 -1614
rect 464 -1671 465 -1645
rect 485 -1671 486 -1645
rect 506 -1646 507 -1614
rect 541 -1646 542 -1614
rect 583 -1671 584 -1645
rect 614 -1646 615 -1614
rect 842 -1646 843 -1614
rect 135 -1671 136 -1647
rect 152 -1671 153 -1647
rect 156 -1648 157 -1614
rect 898 -1648 899 -1614
rect 100 -1650 101 -1614
rect 156 -1671 157 -1649
rect 170 -1671 171 -1649
rect 201 -1650 202 -1614
rect 306 -1671 307 -1649
rect 373 -1671 374 -1649
rect 394 -1650 395 -1614
rect 828 -1650 829 -1614
rect 842 -1671 843 -1649
rect 877 -1650 878 -1614
rect 51 -1652 52 -1614
rect 100 -1671 101 -1651
rect 177 -1652 178 -1614
rect 219 -1671 220 -1651
rect 317 -1671 318 -1651
rect 555 -1652 556 -1614
rect 716 -1671 717 -1651
rect 835 -1652 836 -1614
rect 40 -1671 41 -1653
rect 51 -1671 52 -1653
rect 184 -1654 185 -1614
rect 275 -1671 276 -1653
rect 324 -1671 325 -1653
rect 541 -1671 542 -1653
rect 555 -1671 556 -1653
rect 674 -1654 675 -1614
rect 733 -1671 734 -1653
rect 884 -1654 885 -1614
rect 184 -1671 185 -1655
rect 191 -1656 192 -1614
rect 331 -1671 332 -1655
rect 415 -1656 416 -1614
rect 436 -1671 437 -1655
rect 457 -1656 458 -1614
rect 506 -1671 507 -1655
rect 548 -1656 549 -1614
rect 744 -1671 745 -1655
rect 807 -1656 808 -1614
rect 884 -1671 885 -1655
rect 947 -1656 948 -1614
rect 191 -1671 192 -1657
rect 334 -1671 335 -1657
rect 338 -1658 339 -1614
rect 359 -1671 360 -1657
rect 394 -1671 395 -1657
rect 450 -1658 451 -1614
rect 786 -1658 787 -1614
rect 828 -1671 829 -1657
rect 303 -1671 304 -1659
rect 457 -1671 458 -1659
rect 772 -1660 773 -1614
rect 786 -1671 787 -1659
rect 800 -1660 801 -1614
rect 835 -1671 836 -1659
rect 313 -1662 314 -1614
rect 415 -1671 416 -1661
rect 429 -1671 430 -1661
rect 450 -1671 451 -1661
rect 800 -1671 801 -1661
rect 961 -1662 962 -1614
rect 807 -1671 808 -1663
rect 863 -1664 864 -1614
rect 863 -1671 864 -1665
rect 891 -1666 892 -1614
rect 891 -1671 892 -1667
rect 905 -1668 906 -1614
rect 905 -1671 906 -1669
rect 912 -1670 913 -1614
rect 44 -1708 45 -1680
rect 51 -1681 52 -1679
rect 65 -1681 66 -1679
rect 103 -1708 104 -1680
rect 107 -1681 108 -1679
rect 254 -1708 255 -1680
rect 264 -1708 265 -1680
rect 324 -1681 325 -1679
rect 359 -1681 360 -1679
rect 359 -1708 360 -1680
rect 359 -1681 360 -1679
rect 359 -1708 360 -1680
rect 366 -1681 367 -1679
rect 366 -1708 367 -1680
rect 366 -1681 367 -1679
rect 366 -1708 367 -1680
rect 383 -1708 384 -1680
rect 387 -1681 388 -1679
rect 408 -1681 409 -1679
rect 499 -1681 500 -1679
rect 513 -1708 514 -1680
rect 523 -1681 524 -1679
rect 541 -1708 542 -1680
rect 569 -1681 570 -1679
rect 593 -1708 594 -1680
rect 597 -1681 598 -1679
rect 611 -1681 612 -1679
rect 618 -1708 619 -1680
rect 625 -1681 626 -1679
rect 639 -1708 640 -1680
rect 646 -1681 647 -1679
rect 688 -1681 689 -1679
rect 723 -1681 724 -1679
rect 730 -1708 731 -1680
rect 758 -1681 759 -1679
rect 772 -1708 773 -1680
rect 779 -1708 780 -1680
rect 852 -1681 853 -1679
rect 856 -1708 857 -1680
rect 863 -1681 864 -1679
rect 898 -1708 899 -1680
rect 905 -1681 906 -1679
rect 968 -1681 969 -1679
rect 968 -1708 969 -1680
rect 968 -1681 969 -1679
rect 968 -1708 969 -1680
rect 1024 -1681 1025 -1679
rect 1024 -1708 1025 -1680
rect 1024 -1681 1025 -1679
rect 1024 -1708 1025 -1680
rect 47 -1683 48 -1679
rect 58 -1708 59 -1682
rect 86 -1683 87 -1679
rect 306 -1683 307 -1679
rect 310 -1683 311 -1679
rect 376 -1708 377 -1682
rect 380 -1683 381 -1679
rect 387 -1708 388 -1682
rect 422 -1683 423 -1679
rect 425 -1683 426 -1679
rect 429 -1708 430 -1682
rect 443 -1683 444 -1679
rect 450 -1683 451 -1679
rect 474 -1708 475 -1682
rect 520 -1683 521 -1679
rect 590 -1683 591 -1679
rect 604 -1683 605 -1679
rect 611 -1708 612 -1682
rect 632 -1683 633 -1679
rect 646 -1708 647 -1682
rect 653 -1708 654 -1682
rect 695 -1683 696 -1679
rect 709 -1683 710 -1679
rect 723 -1708 724 -1682
rect 737 -1683 738 -1679
rect 758 -1708 759 -1682
rect 782 -1683 783 -1679
rect 807 -1683 808 -1679
rect 817 -1708 818 -1682
rect 884 -1683 885 -1679
rect 93 -1685 94 -1679
rect 201 -1685 202 -1679
rect 212 -1685 213 -1679
rect 334 -1685 335 -1679
rect 373 -1685 374 -1679
rect 408 -1708 409 -1684
rect 422 -1708 423 -1684
rect 436 -1685 437 -1679
rect 450 -1708 451 -1684
rect 485 -1685 486 -1679
rect 569 -1708 570 -1684
rect 691 -1685 692 -1679
rect 709 -1708 710 -1684
rect 716 -1685 717 -1679
rect 737 -1708 738 -1684
rect 744 -1685 745 -1679
rect 786 -1685 787 -1679
rect 849 -1685 850 -1679
rect 884 -1708 885 -1684
rect 891 -1685 892 -1679
rect 75 -1687 76 -1679
rect 93 -1708 94 -1686
rect 100 -1687 101 -1679
rect 180 -1687 181 -1679
rect 201 -1708 202 -1686
rect 226 -1687 227 -1679
rect 233 -1687 234 -1679
rect 233 -1708 234 -1686
rect 233 -1687 234 -1679
rect 233 -1708 234 -1686
rect 240 -1687 241 -1679
rect 243 -1707 244 -1686
rect 282 -1687 283 -1679
rect 303 -1708 304 -1686
rect 310 -1708 311 -1686
rect 345 -1687 346 -1679
rect 373 -1708 374 -1686
rect 464 -1687 465 -1679
rect 576 -1687 577 -1679
rect 604 -1708 605 -1686
rect 667 -1687 668 -1679
rect 674 -1708 675 -1686
rect 677 -1687 678 -1679
rect 681 -1687 682 -1679
rect 744 -1708 745 -1686
rect 751 -1687 752 -1679
rect 793 -1687 794 -1679
rect 800 -1708 801 -1686
rect 807 -1708 808 -1686
rect 842 -1687 843 -1679
rect 849 -1708 850 -1686
rect 866 -1708 867 -1686
rect 114 -1708 115 -1688
rect 149 -1708 150 -1688
rect 156 -1689 157 -1679
rect 198 -1689 199 -1679
rect 219 -1689 220 -1679
rect 226 -1708 227 -1688
rect 240 -1708 241 -1688
rect 275 -1689 276 -1679
rect 324 -1708 325 -1688
rect 341 -1689 342 -1679
rect 345 -1708 346 -1688
rect 352 -1689 353 -1679
rect 401 -1689 402 -1679
rect 520 -1708 521 -1688
rect 527 -1689 528 -1679
rect 576 -1708 577 -1688
rect 702 -1689 703 -1679
rect 751 -1708 752 -1688
rect 765 -1689 766 -1679
rect 793 -1708 794 -1688
rect 821 -1689 822 -1679
rect 835 -1708 836 -1688
rect 117 -1691 118 -1679
rect 121 -1691 122 -1679
rect 128 -1691 129 -1679
rect 180 -1708 181 -1690
rect 184 -1691 185 -1679
rect 219 -1708 220 -1690
rect 247 -1691 248 -1679
rect 341 -1708 342 -1690
rect 404 -1708 405 -1690
rect 443 -1708 444 -1690
rect 464 -1708 465 -1690
rect 534 -1691 535 -1679
rect 765 -1708 766 -1690
rect 814 -1691 815 -1679
rect 821 -1708 822 -1690
rect 863 -1708 864 -1690
rect 128 -1708 129 -1692
rect 135 -1693 136 -1679
rect 142 -1693 143 -1679
rect 142 -1708 143 -1692
rect 142 -1693 143 -1679
rect 142 -1708 143 -1692
rect 156 -1708 157 -1692
rect 177 -1693 178 -1679
rect 268 -1693 269 -1679
rect 282 -1708 283 -1692
rect 415 -1693 416 -1679
rect 485 -1708 486 -1692
rect 527 -1708 528 -1692
rect 555 -1693 556 -1679
rect 828 -1693 829 -1679
rect 828 -1708 829 -1692
rect 828 -1693 829 -1679
rect 828 -1708 829 -1692
rect 163 -1695 164 -1679
rect 208 -1708 209 -1694
rect 261 -1695 262 -1679
rect 268 -1708 269 -1694
rect 275 -1708 276 -1694
rect 289 -1695 290 -1679
rect 394 -1695 395 -1679
rect 415 -1708 416 -1694
rect 436 -1708 437 -1694
rect 478 -1695 479 -1679
rect 163 -1708 164 -1696
rect 191 -1697 192 -1679
rect 289 -1708 290 -1696
rect 317 -1697 318 -1679
rect 394 -1708 395 -1696
rect 432 -1697 433 -1679
rect 457 -1697 458 -1679
rect 534 -1708 535 -1696
rect 170 -1699 171 -1679
rect 170 -1708 171 -1698
rect 170 -1699 171 -1679
rect 170 -1708 171 -1698
rect 177 -1708 178 -1698
rect 355 -1708 356 -1698
rect 457 -1708 458 -1698
rect 548 -1699 549 -1679
rect 191 -1708 192 -1700
rect 215 -1708 216 -1700
rect 317 -1708 318 -1700
rect 331 -1701 332 -1679
rect 471 -1701 472 -1679
rect 555 -1708 556 -1700
rect 331 -1708 332 -1702
rect 478 -1708 479 -1702
rect 506 -1703 507 -1679
rect 548 -1708 549 -1702
rect 562 -1703 563 -1679
rect 492 -1705 493 -1679
rect 506 -1708 507 -1704
rect 562 -1708 563 -1704
rect 583 -1705 584 -1679
rect 425 -1708 426 -1706
rect 492 -1708 493 -1706
rect 583 -1708 584 -1706
rect 590 -1708 591 -1706
rect 44 -1718 45 -1716
rect 44 -1741 45 -1717
rect 44 -1718 45 -1716
rect 44 -1741 45 -1717
rect 58 -1718 59 -1716
rect 65 -1741 66 -1717
rect 93 -1718 94 -1716
rect 117 -1718 118 -1716
rect 121 -1741 122 -1717
rect 128 -1718 129 -1716
rect 142 -1718 143 -1716
rect 152 -1741 153 -1717
rect 156 -1718 157 -1716
rect 184 -1718 185 -1716
rect 191 -1718 192 -1716
rect 191 -1741 192 -1717
rect 191 -1718 192 -1716
rect 191 -1741 192 -1717
rect 212 -1718 213 -1716
rect 240 -1718 241 -1716
rect 268 -1718 269 -1716
rect 275 -1741 276 -1717
rect 289 -1718 290 -1716
rect 401 -1718 402 -1716
rect 411 -1741 412 -1717
rect 520 -1718 521 -1716
rect 541 -1718 542 -1716
rect 541 -1741 542 -1717
rect 541 -1718 542 -1716
rect 541 -1741 542 -1717
rect 562 -1718 563 -1716
rect 590 -1741 591 -1717
rect 593 -1718 594 -1716
rect 782 -1741 783 -1717
rect 793 -1718 794 -1716
rect 796 -1718 797 -1716
rect 800 -1718 801 -1716
rect 800 -1741 801 -1717
rect 800 -1718 801 -1716
rect 800 -1741 801 -1717
rect 828 -1718 829 -1716
rect 866 -1718 867 -1716
rect 884 -1718 885 -1716
rect 884 -1741 885 -1717
rect 884 -1718 885 -1716
rect 884 -1741 885 -1717
rect 898 -1718 899 -1716
rect 898 -1741 899 -1717
rect 898 -1718 899 -1716
rect 898 -1741 899 -1717
rect 968 -1718 969 -1716
rect 968 -1741 969 -1717
rect 968 -1718 969 -1716
rect 968 -1741 969 -1717
rect 1024 -1718 1025 -1716
rect 1024 -1741 1025 -1717
rect 1024 -1718 1025 -1716
rect 1024 -1741 1025 -1717
rect 100 -1720 101 -1716
rect 100 -1741 101 -1719
rect 100 -1720 101 -1716
rect 100 -1741 101 -1719
rect 103 -1720 104 -1716
rect 145 -1741 146 -1719
rect 149 -1720 150 -1716
rect 177 -1741 178 -1719
rect 205 -1741 206 -1719
rect 212 -1741 213 -1719
rect 215 -1720 216 -1716
rect 278 -1720 279 -1716
rect 299 -1720 300 -1716
rect 569 -1720 570 -1716
rect 583 -1720 584 -1716
rect 597 -1720 598 -1716
rect 604 -1720 605 -1716
rect 653 -1720 654 -1716
rect 674 -1720 675 -1716
rect 681 -1720 682 -1716
rect 702 -1741 703 -1719
rect 709 -1720 710 -1716
rect 723 -1720 724 -1716
rect 723 -1741 724 -1719
rect 723 -1720 724 -1716
rect 723 -1741 724 -1719
rect 730 -1720 731 -1716
rect 733 -1740 734 -1719
rect 772 -1720 773 -1716
rect 786 -1741 787 -1719
rect 793 -1741 794 -1719
rect 807 -1720 808 -1716
rect 821 -1720 822 -1716
rect 828 -1741 829 -1719
rect 835 -1720 836 -1716
rect 842 -1741 843 -1719
rect 845 -1720 846 -1716
rect 856 -1720 857 -1716
rect 107 -1741 108 -1721
rect 114 -1741 115 -1721
rect 142 -1741 143 -1721
rect 156 -1741 157 -1721
rect 163 -1722 164 -1716
rect 184 -1741 185 -1721
rect 219 -1722 220 -1716
rect 261 -1722 262 -1716
rect 303 -1722 304 -1716
rect 303 -1741 304 -1721
rect 303 -1722 304 -1716
rect 303 -1741 304 -1721
rect 310 -1722 311 -1716
rect 310 -1741 311 -1721
rect 310 -1722 311 -1716
rect 310 -1741 311 -1721
rect 324 -1722 325 -1716
rect 369 -1741 370 -1721
rect 380 -1741 381 -1721
rect 408 -1722 409 -1716
rect 422 -1722 423 -1716
rect 446 -1741 447 -1721
rect 464 -1722 465 -1716
rect 499 -1722 500 -1716
rect 597 -1741 598 -1721
rect 618 -1722 619 -1716
rect 639 -1722 640 -1716
rect 656 -1741 657 -1721
rect 709 -1741 710 -1721
rect 779 -1722 780 -1716
rect 849 -1722 850 -1716
rect 856 -1741 857 -1721
rect 163 -1741 164 -1723
rect 170 -1724 171 -1716
rect 226 -1724 227 -1716
rect 240 -1741 241 -1723
rect 296 -1724 297 -1716
rect 324 -1741 325 -1723
rect 338 -1724 339 -1716
rect 345 -1724 346 -1716
rect 352 -1724 353 -1716
rect 611 -1724 612 -1716
rect 646 -1724 647 -1716
rect 646 -1741 647 -1723
rect 646 -1724 647 -1716
rect 646 -1741 647 -1723
rect 730 -1741 731 -1723
rect 737 -1724 738 -1716
rect 233 -1726 234 -1716
rect 247 -1741 248 -1725
rect 282 -1726 283 -1716
rect 296 -1741 297 -1725
rect 338 -1741 339 -1725
rect 373 -1726 374 -1716
rect 422 -1741 423 -1725
rect 429 -1726 430 -1716
rect 464 -1741 465 -1725
rect 478 -1726 479 -1716
rect 492 -1726 493 -1716
rect 520 -1741 521 -1725
rect 737 -1741 738 -1725
rect 744 -1726 745 -1716
rect 226 -1741 227 -1727
rect 233 -1741 234 -1727
rect 331 -1728 332 -1716
rect 373 -1741 374 -1727
rect 429 -1741 430 -1727
rect 457 -1728 458 -1716
rect 471 -1728 472 -1716
rect 576 -1728 577 -1716
rect 744 -1741 745 -1727
rect 765 -1728 766 -1716
rect 317 -1730 318 -1716
rect 331 -1741 332 -1729
rect 345 -1741 346 -1729
rect 359 -1730 360 -1716
rect 366 -1730 367 -1716
rect 376 -1740 377 -1729
rect 457 -1741 458 -1729
rect 548 -1730 549 -1716
rect 555 -1730 556 -1716
rect 576 -1741 577 -1729
rect 758 -1730 759 -1716
rect 765 -1741 766 -1729
rect 254 -1732 255 -1716
rect 317 -1741 318 -1731
rect 352 -1741 353 -1731
rect 383 -1732 384 -1716
rect 478 -1741 479 -1731
rect 506 -1732 507 -1716
rect 534 -1732 535 -1716
rect 548 -1741 549 -1731
rect 555 -1741 556 -1731
rect 569 -1741 570 -1731
rect 751 -1732 752 -1716
rect 758 -1741 759 -1731
rect 359 -1741 360 -1733
rect 415 -1734 416 -1716
rect 485 -1734 486 -1716
rect 492 -1741 493 -1733
rect 499 -1741 500 -1733
rect 527 -1734 528 -1716
rect 366 -1741 367 -1735
rect 394 -1736 395 -1716
rect 415 -1741 416 -1735
rect 450 -1736 451 -1716
rect 513 -1736 514 -1716
rect 534 -1741 535 -1735
rect 394 -1741 395 -1737
rect 436 -1738 437 -1716
rect 450 -1741 451 -1737
rect 485 -1741 486 -1737
rect 513 -1741 514 -1737
rect 436 -1741 437 -1739
rect 443 -1740 444 -1716
rect 796 -1741 797 -1739
rect 807 -1741 808 -1739
rect 44 -1751 45 -1749
rect 47 -1768 48 -1750
rect 58 -1768 59 -1750
rect 61 -1751 62 -1749
rect 65 -1751 66 -1749
rect 72 -1768 73 -1750
rect 93 -1768 94 -1750
rect 117 -1768 118 -1750
rect 121 -1751 122 -1749
rect 135 -1751 136 -1749
rect 156 -1751 157 -1749
rect 156 -1768 157 -1750
rect 156 -1751 157 -1749
rect 156 -1768 157 -1750
rect 159 -1751 160 -1749
rect 177 -1751 178 -1749
rect 184 -1751 185 -1749
rect 212 -1768 213 -1750
rect 219 -1751 220 -1749
rect 247 -1751 248 -1749
rect 275 -1751 276 -1749
rect 275 -1768 276 -1750
rect 275 -1751 276 -1749
rect 275 -1768 276 -1750
rect 282 -1768 283 -1750
rect 303 -1751 304 -1749
rect 352 -1751 353 -1749
rect 369 -1768 370 -1750
rect 373 -1751 374 -1749
rect 401 -1768 402 -1750
rect 415 -1751 416 -1749
rect 415 -1768 416 -1750
rect 415 -1751 416 -1749
rect 415 -1768 416 -1750
rect 422 -1751 423 -1749
rect 422 -1768 423 -1750
rect 422 -1751 423 -1749
rect 422 -1768 423 -1750
rect 443 -1768 444 -1750
rect 457 -1751 458 -1749
rect 464 -1751 465 -1749
rect 471 -1751 472 -1749
rect 478 -1751 479 -1749
rect 478 -1768 479 -1750
rect 478 -1751 479 -1749
rect 478 -1768 479 -1750
rect 488 -1751 489 -1749
rect 576 -1751 577 -1749
rect 586 -1751 587 -1749
rect 590 -1751 591 -1749
rect 646 -1751 647 -1749
rect 656 -1751 657 -1749
rect 716 -1751 717 -1749
rect 730 -1751 731 -1749
rect 765 -1751 766 -1749
rect 782 -1751 783 -1749
rect 807 -1751 808 -1749
rect 814 -1768 815 -1750
rect 828 -1751 829 -1749
rect 828 -1768 829 -1750
rect 828 -1751 829 -1749
rect 828 -1768 829 -1750
rect 842 -1751 843 -1749
rect 845 -1768 846 -1750
rect 856 -1751 857 -1749
rect 856 -1768 857 -1750
rect 856 -1751 857 -1749
rect 856 -1768 857 -1750
rect 884 -1751 885 -1749
rect 884 -1768 885 -1750
rect 884 -1751 885 -1749
rect 884 -1768 885 -1750
rect 898 -1751 899 -1749
rect 898 -1768 899 -1750
rect 898 -1751 899 -1749
rect 898 -1768 899 -1750
rect 968 -1751 969 -1749
rect 975 -1751 976 -1749
rect 1024 -1751 1025 -1749
rect 1024 -1768 1025 -1750
rect 1024 -1751 1025 -1749
rect 1024 -1768 1025 -1750
rect 65 -1768 66 -1752
rect 79 -1768 80 -1752
rect 100 -1753 101 -1749
rect 100 -1768 101 -1752
rect 100 -1753 101 -1749
rect 100 -1768 101 -1752
rect 107 -1753 108 -1749
rect 121 -1768 122 -1752
rect 128 -1753 129 -1749
rect 145 -1753 146 -1749
rect 163 -1753 164 -1749
rect 173 -1753 174 -1749
rect 191 -1753 192 -1749
rect 191 -1768 192 -1752
rect 191 -1753 192 -1749
rect 191 -1768 192 -1752
rect 205 -1753 206 -1749
rect 205 -1768 206 -1752
rect 205 -1753 206 -1749
rect 205 -1768 206 -1752
rect 219 -1768 220 -1752
rect 233 -1753 234 -1749
rect 289 -1768 290 -1752
rect 310 -1753 311 -1749
rect 317 -1753 318 -1749
rect 352 -1768 353 -1752
rect 366 -1753 367 -1749
rect 373 -1768 374 -1752
rect 380 -1753 381 -1749
rect 380 -1768 381 -1752
rect 380 -1753 381 -1749
rect 380 -1768 381 -1752
rect 387 -1753 388 -1749
rect 404 -1753 405 -1749
rect 450 -1753 451 -1749
rect 464 -1768 465 -1752
rect 471 -1768 472 -1752
rect 492 -1753 493 -1749
rect 499 -1753 500 -1749
rect 509 -1753 510 -1749
rect 513 -1753 514 -1749
rect 513 -1768 514 -1752
rect 513 -1753 514 -1749
rect 513 -1768 514 -1752
rect 527 -1768 528 -1752
rect 541 -1753 542 -1749
rect 548 -1753 549 -1749
rect 555 -1753 556 -1749
rect 562 -1753 563 -1749
rect 597 -1753 598 -1749
rect 709 -1753 710 -1749
rect 730 -1768 731 -1752
rect 772 -1753 773 -1749
rect 786 -1753 787 -1749
rect 128 -1768 129 -1754
rect 131 -1755 132 -1749
rect 135 -1768 136 -1754
rect 142 -1755 143 -1749
rect 170 -1755 171 -1749
rect 170 -1768 171 -1754
rect 170 -1755 171 -1749
rect 170 -1768 171 -1754
rect 233 -1768 234 -1754
rect 240 -1755 241 -1749
rect 296 -1755 297 -1749
rect 317 -1768 318 -1754
rect 394 -1755 395 -1749
rect 394 -1768 395 -1754
rect 394 -1755 395 -1749
rect 394 -1768 395 -1754
rect 429 -1755 430 -1749
rect 450 -1768 451 -1754
rect 457 -1768 458 -1754
rect 520 -1755 521 -1749
rect 530 -1755 531 -1749
rect 534 -1755 535 -1749
rect 562 -1768 563 -1754
rect 569 -1755 570 -1749
rect 702 -1755 703 -1749
rect 709 -1768 710 -1754
rect 723 -1755 724 -1749
rect 723 -1768 724 -1754
rect 723 -1755 724 -1749
rect 723 -1768 724 -1754
rect 758 -1755 759 -1749
rect 772 -1768 773 -1754
rect 779 -1755 780 -1749
rect 793 -1755 794 -1749
rect 138 -1757 139 -1749
rect 142 -1768 143 -1756
rect 229 -1768 230 -1756
rect 240 -1768 241 -1756
rect 296 -1768 297 -1756
rect 331 -1757 332 -1749
rect 429 -1768 430 -1756
rect 436 -1757 437 -1749
rect 506 -1757 507 -1749
rect 506 -1768 507 -1756
rect 506 -1757 507 -1749
rect 506 -1768 507 -1756
rect 751 -1757 752 -1749
rect 758 -1768 759 -1756
rect 793 -1768 794 -1756
rect 800 -1757 801 -1749
rect 310 -1768 311 -1758
rect 338 -1759 339 -1749
rect 737 -1759 738 -1749
rect 751 -1768 752 -1758
rect 324 -1761 325 -1749
rect 338 -1768 339 -1760
rect 737 -1768 738 -1760
rect 744 -1761 745 -1749
rect 324 -1768 325 -1762
rect 345 -1763 346 -1749
rect 345 -1768 346 -1764
rect 359 -1765 360 -1749
rect 359 -1768 360 -1766
rect 411 -1767 412 -1749
rect 58 -1778 59 -1776
rect 65 -1778 66 -1776
rect 75 -1789 76 -1777
rect 79 -1778 80 -1776
rect 93 -1778 94 -1776
rect 110 -1778 111 -1776
rect 117 -1778 118 -1776
rect 128 -1778 129 -1776
rect 135 -1778 136 -1776
rect 152 -1778 153 -1776
rect 170 -1778 171 -1776
rect 173 -1789 174 -1777
rect 191 -1778 192 -1776
rect 198 -1778 199 -1776
rect 205 -1778 206 -1776
rect 205 -1789 206 -1777
rect 205 -1778 206 -1776
rect 205 -1789 206 -1777
rect 219 -1778 220 -1776
rect 226 -1778 227 -1776
rect 240 -1778 241 -1776
rect 240 -1789 241 -1777
rect 240 -1778 241 -1776
rect 240 -1789 241 -1777
rect 247 -1789 248 -1777
rect 261 -1789 262 -1777
rect 282 -1778 283 -1776
rect 320 -1789 321 -1777
rect 331 -1778 332 -1776
rect 345 -1778 346 -1776
rect 352 -1778 353 -1776
rect 352 -1789 353 -1777
rect 352 -1778 353 -1776
rect 352 -1789 353 -1777
rect 380 -1778 381 -1776
rect 387 -1789 388 -1777
rect 394 -1778 395 -1776
rect 411 -1778 412 -1776
rect 415 -1778 416 -1776
rect 415 -1789 416 -1777
rect 415 -1778 416 -1776
rect 415 -1789 416 -1777
rect 443 -1778 444 -1776
rect 443 -1789 444 -1777
rect 443 -1778 444 -1776
rect 443 -1789 444 -1777
rect 478 -1778 479 -1776
rect 478 -1789 479 -1777
rect 478 -1778 479 -1776
rect 478 -1789 479 -1777
rect 502 -1789 503 -1777
rect 506 -1778 507 -1776
rect 513 -1778 514 -1776
rect 513 -1789 514 -1777
rect 513 -1778 514 -1776
rect 513 -1789 514 -1777
rect 520 -1789 521 -1777
rect 527 -1778 528 -1776
rect 562 -1778 563 -1776
rect 565 -1789 566 -1777
rect 709 -1778 710 -1776
rect 716 -1778 717 -1776
rect 723 -1778 724 -1776
rect 747 -1778 748 -1776
rect 751 -1778 752 -1776
rect 765 -1789 766 -1777
rect 772 -1778 773 -1776
rect 779 -1778 780 -1776
rect 793 -1778 794 -1776
rect 793 -1789 794 -1777
rect 793 -1778 794 -1776
rect 793 -1789 794 -1777
rect 814 -1778 815 -1776
rect 814 -1789 815 -1777
rect 814 -1778 815 -1776
rect 814 -1789 815 -1777
rect 828 -1778 829 -1776
rect 838 -1789 839 -1777
rect 880 -1778 881 -1776
rect 884 -1778 885 -1776
rect 898 -1778 899 -1776
rect 898 -1789 899 -1777
rect 898 -1778 899 -1776
rect 898 -1789 899 -1777
rect 1024 -1778 1025 -1776
rect 1024 -1789 1025 -1777
rect 1024 -1778 1025 -1776
rect 1024 -1789 1025 -1777
rect 72 -1780 73 -1776
rect 79 -1789 80 -1779
rect 142 -1780 143 -1776
rect 142 -1789 143 -1779
rect 142 -1780 143 -1776
rect 142 -1789 143 -1779
rect 152 -1789 153 -1779
rect 156 -1789 157 -1779
rect 226 -1789 227 -1779
rect 233 -1780 234 -1776
rect 275 -1780 276 -1776
rect 282 -1789 283 -1779
rect 289 -1780 290 -1776
rect 306 -1780 307 -1776
rect 324 -1780 325 -1776
rect 331 -1789 332 -1779
rect 338 -1780 339 -1776
rect 338 -1789 339 -1779
rect 338 -1780 339 -1776
rect 338 -1789 339 -1779
rect 373 -1780 374 -1776
rect 380 -1789 381 -1779
rect 401 -1780 402 -1776
rect 422 -1789 423 -1779
rect 730 -1780 731 -1776
rect 772 -1789 773 -1779
rect 296 -1782 297 -1776
rect 313 -1789 314 -1781
rect 411 -1789 412 -1781
rect 457 -1782 458 -1776
rect 737 -1782 738 -1776
rect 737 -1789 738 -1781
rect 737 -1782 738 -1776
rect 737 -1789 738 -1781
rect 758 -1782 759 -1776
rect 758 -1789 759 -1781
rect 758 -1782 759 -1776
rect 758 -1789 759 -1781
rect 296 -1789 297 -1783
rect 303 -1789 304 -1783
rect 306 -1789 307 -1783
rect 362 -1784 363 -1776
rect 450 -1784 451 -1776
rect 457 -1789 458 -1783
rect 310 -1786 311 -1776
rect 324 -1789 325 -1785
rect 450 -1789 451 -1785
rect 471 -1786 472 -1776
rect 464 -1788 465 -1776
rect 471 -1789 472 -1787
rect 68 -1799 69 -1797
rect 79 -1799 80 -1797
rect 142 -1799 143 -1797
rect 149 -1799 150 -1797
rect 156 -1799 157 -1797
rect 159 -1804 160 -1798
rect 184 -1799 185 -1797
rect 191 -1804 192 -1798
rect 205 -1799 206 -1797
rect 208 -1804 209 -1798
rect 226 -1799 227 -1797
rect 226 -1804 227 -1798
rect 226 -1799 227 -1797
rect 226 -1804 227 -1798
rect 240 -1799 241 -1797
rect 247 -1799 248 -1797
rect 261 -1799 262 -1797
rect 268 -1804 269 -1798
rect 282 -1799 283 -1797
rect 282 -1804 283 -1798
rect 282 -1799 283 -1797
rect 282 -1804 283 -1798
rect 296 -1799 297 -1797
rect 296 -1804 297 -1798
rect 296 -1799 297 -1797
rect 296 -1804 297 -1798
rect 324 -1799 325 -1797
rect 341 -1804 342 -1798
rect 352 -1799 353 -1797
rect 352 -1804 353 -1798
rect 352 -1799 353 -1797
rect 352 -1804 353 -1798
rect 380 -1799 381 -1797
rect 383 -1804 384 -1798
rect 387 -1799 388 -1797
rect 387 -1804 388 -1798
rect 387 -1799 388 -1797
rect 387 -1804 388 -1798
rect 422 -1799 423 -1797
rect 429 -1799 430 -1797
rect 432 -1799 433 -1797
rect 443 -1799 444 -1797
rect 457 -1799 458 -1797
rect 464 -1804 465 -1798
rect 471 -1799 472 -1797
rect 481 -1804 482 -1798
rect 506 -1799 507 -1797
rect 513 -1799 514 -1797
rect 516 -1804 517 -1798
rect 520 -1799 521 -1797
rect 737 -1799 738 -1797
rect 751 -1804 752 -1798
rect 754 -1799 755 -1797
rect 765 -1799 766 -1797
rect 793 -1799 794 -1797
rect 796 -1804 797 -1798
rect 898 -1799 899 -1797
rect 905 -1804 906 -1798
rect 1024 -1799 1025 -1797
rect 1027 -1804 1028 -1798
rect 331 -1801 332 -1797
rect 345 -1801 346 -1797
rect 415 -1801 416 -1797
rect 422 -1804 423 -1800
rect 439 -1801 440 -1797
rect 450 -1801 451 -1797
rect 471 -1804 472 -1800
rect 478 -1801 479 -1797
rect 744 -1801 745 -1797
rect 758 -1801 759 -1797
rect 331 -1804 332 -1802
rect 338 -1803 339 -1797
rect 187 -1814 188 -1812
rect 191 -1814 192 -1812
rect 222 -1814 223 -1812
rect 226 -1814 227 -1812
rect 264 -1814 265 -1812
rect 268 -1814 269 -1812
rect 296 -1814 297 -1812
rect 306 -1814 307 -1812
rect 324 -1814 325 -1812
rect 331 -1814 332 -1812
rect 352 -1814 353 -1812
rect 359 -1814 360 -1812
rect 376 -1814 377 -1812
rect 387 -1814 388 -1812
rect 422 -1814 423 -1812
rect 429 -1814 430 -1812
rect 747 -1814 748 -1812
rect 751 -1814 752 -1812
rect 901 -1814 902 -1812
rect 905 -1814 906 -1812
<< labels >>
rlabel pdiffusion 3 -8 3 -8 0 cellNo=73
rlabel pdiffusion 10 -8 10 -8 0 cellNo=281
rlabel pdiffusion 17 -8 17 -8 0 cellNo=262
rlabel pdiffusion 24 -8 24 -8 0 cellNo=342
rlabel pdiffusion 31 -8 31 -8 0 cellNo=409
rlabel pdiffusion 38 -8 38 -8 0 cellNo=561
rlabel pdiffusion 45 -8 45 -8 0 cellNo=695
rlabel pdiffusion 178 -8 178 -8 0 feedthrough
rlabel pdiffusion 185 -8 185 -8 0 feedthrough
rlabel pdiffusion 192 -8 192 -8 0 cellNo=24
rlabel pdiffusion 199 -8 199 -8 0 cellNo=130
rlabel pdiffusion 213 -8 213 -8 0 cellNo=80
rlabel pdiffusion 220 -8 220 -8 0 feedthrough
rlabel pdiffusion 234 -8 234 -8 0 cellNo=252
rlabel pdiffusion 241 -8 241 -8 0 feedthrough
rlabel pdiffusion 255 -8 255 -8 0 cellNo=642
rlabel pdiffusion 262 -8 262 -8 0 feedthrough
rlabel pdiffusion 276 -8 276 -8 0 cellNo=5
rlabel pdiffusion 283 -8 283 -8 0 cellNo=249
rlabel pdiffusion 290 -8 290 -8 0 feedthrough
rlabel pdiffusion 297 -8 297 -8 0 cellNo=394
rlabel pdiffusion 304 -8 304 -8 0 feedthrough
rlabel pdiffusion 311 -8 311 -8 0 cellNo=26
rlabel pdiffusion 318 -8 318 -8 0 cellNo=79
rlabel pdiffusion 339 -8 339 -8 0 feedthrough
rlabel pdiffusion 346 -8 346 -8 0 cellNo=131
rlabel pdiffusion 353 -8 353 -8 0 feedthrough
rlabel pdiffusion 360 -8 360 -8 0 cellNo=311
rlabel pdiffusion 367 -8 367 -8 0 feedthrough
rlabel pdiffusion 409 -8 409 -8 0 cellNo=866
rlabel pdiffusion 423 -8 423 -8 0 cellNo=17
rlabel pdiffusion 458 -8 458 -8 0 cellNo=625
rlabel pdiffusion 465 -8 465 -8 0 cellNo=21
rlabel pdiffusion 472 -8 472 -8 0 feedthrough
rlabel pdiffusion 479 -8 479 -8 0 cellNo=3
rlabel pdiffusion 486 -8 486 -8 0 feedthrough
rlabel pdiffusion 535 -8 535 -8 0 cellNo=213
rlabel pdiffusion 542 -8 542 -8 0 feedthrough
rlabel pdiffusion 556 -8 556 -8 0 cellNo=826
rlabel pdiffusion 577 -8 577 -8 0 cellNo=731
rlabel pdiffusion 584 -8 584 -8 0 feedthrough
rlabel pdiffusion 605 -8 605 -8 0 feedthrough
rlabel pdiffusion 612 -8 612 -8 0 cellNo=433
rlabel pdiffusion 619 -8 619 -8 0 cellNo=802
rlabel pdiffusion 731 -8 731 -8 0 feedthrough
rlabel pdiffusion 738 -8 738 -8 0 cellNo=483
rlabel pdiffusion 3 -25 3 -25 0 cellNo=35
rlabel pdiffusion 10 -25 10 -25 0 cellNo=322
rlabel pdiffusion 17 -25 17 -25 0 cellNo=365
rlabel pdiffusion 24 -25 24 -25 0 cellNo=40
rlabel pdiffusion 31 -25 31 -25 0 cellNo=47
rlabel pdiffusion 38 -25 38 -25 0 cellNo=60
rlabel pdiffusion 45 -25 45 -25 0 cellNo=293
rlabel pdiffusion 52 -25 52 -25 0 cellNo=347
rlabel pdiffusion 59 -25 59 -25 0 cellNo=42
rlabel pdiffusion 66 -25 66 -25 0 cellNo=559
rlabel pdiffusion 80 -25 80 -25 0 cellNo=46
rlabel pdiffusion 115 -25 115 -25 0 cellNo=431
rlabel pdiffusion 122 -25 122 -25 0 feedthrough
rlabel pdiffusion 129 -25 129 -25 0 cellNo=324
rlabel pdiffusion 157 -25 157 -25 0 cellNo=297
rlabel pdiffusion 164 -25 164 -25 0 feedthrough
rlabel pdiffusion 171 -25 171 -25 0 feedthrough
rlabel pdiffusion 178 -25 178 -25 0 cellNo=615
rlabel pdiffusion 185 -25 185 -25 0 feedthrough
rlabel pdiffusion 213 -25 213 -25 0 cellNo=747
rlabel pdiffusion 220 -25 220 -25 0 feedthrough
rlabel pdiffusion 227 -25 227 -25 0 feedthrough
rlabel pdiffusion 241 -25 241 -25 0 feedthrough
rlabel pdiffusion 248 -25 248 -25 0 feedthrough
rlabel pdiffusion 255 -25 255 -25 0 feedthrough
rlabel pdiffusion 262 -25 262 -25 0 cellNo=52
rlabel pdiffusion 269 -25 269 -25 0 cellNo=59
rlabel pdiffusion 276 -25 276 -25 0 cellNo=554
rlabel pdiffusion 283 -25 283 -25 0 feedthrough
rlabel pdiffusion 290 -25 290 -25 0 feedthrough
rlabel pdiffusion 297 -25 297 -25 0 feedthrough
rlabel pdiffusion 304 -25 304 -25 0 feedthrough
rlabel pdiffusion 311 -25 311 -25 0 feedthrough
rlabel pdiffusion 318 -25 318 -25 0 feedthrough
rlabel pdiffusion 332 -25 332 -25 0 cellNo=36
rlabel pdiffusion 339 -25 339 -25 0 feedthrough
rlabel pdiffusion 346 -25 346 -25 0 feedthrough
rlabel pdiffusion 353 -25 353 -25 0 feedthrough
rlabel pdiffusion 360 -25 360 -25 0 feedthrough
rlabel pdiffusion 367 -25 367 -25 0 feedthrough
rlabel pdiffusion 374 -25 374 -25 0 cellNo=135
rlabel pdiffusion 381 -25 381 -25 0 cellNo=502
rlabel pdiffusion 409 -25 409 -25 0 cellNo=45
rlabel pdiffusion 416 -25 416 -25 0 feedthrough
rlabel pdiffusion 423 -25 423 -25 0 cellNo=459
rlabel pdiffusion 430 -25 430 -25 0 feedthrough
rlabel pdiffusion 437 -25 437 -25 0 cellNo=53
rlabel pdiffusion 444 -25 444 -25 0 feedthrough
rlabel pdiffusion 451 -25 451 -25 0 feedthrough
rlabel pdiffusion 458 -25 458 -25 0 feedthrough
rlabel pdiffusion 465 -25 465 -25 0 cellNo=37
rlabel pdiffusion 472 -25 472 -25 0 cellNo=34
rlabel pdiffusion 479 -25 479 -25 0 feedthrough
rlabel pdiffusion 486 -25 486 -25 0 feedthrough
rlabel pdiffusion 493 -25 493 -25 0 feedthrough
rlabel pdiffusion 528 -25 528 -25 0 feedthrough
rlabel pdiffusion 542 -25 542 -25 0 feedthrough
rlabel pdiffusion 577 -25 577 -25 0 cellNo=221
rlabel pdiffusion 584 -25 584 -25 0 feedthrough
rlabel pdiffusion 605 -25 605 -25 0 feedthrough
rlabel pdiffusion 612 -25 612 -25 0 feedthrough
rlabel pdiffusion 619 -25 619 -25 0 feedthrough
rlabel pdiffusion 689 -25 689 -25 0 feedthrough
rlabel pdiffusion 696 -25 696 -25 0 cellNo=505
rlabel pdiffusion 710 -25 710 -25 0 cellNo=865
rlabel pdiffusion 731 -25 731 -25 0 feedthrough
rlabel pdiffusion 3 -48 3 -48 0 cellNo=68
rlabel pdiffusion 10 -48 10 -48 0 cellNo=474
rlabel pdiffusion 17 -48 17 -48 0 cellNo=536
rlabel pdiffusion 24 -48 24 -48 0 cellNo=556
rlabel pdiffusion 31 -48 31 -48 0 cellNo=671
rlabel pdiffusion 59 -48 59 -48 0 feedthrough
rlabel pdiffusion 66 -48 66 -48 0 cellNo=384
rlabel pdiffusion 80 -48 80 -48 0 feedthrough
rlabel pdiffusion 108 -48 108 -48 0 cellNo=257
rlabel pdiffusion 115 -48 115 -48 0 feedthrough
rlabel pdiffusion 122 -48 122 -48 0 cellNo=774
rlabel pdiffusion 129 -48 129 -48 0 cellNo=11
rlabel pdiffusion 136 -48 136 -48 0 feedthrough
rlabel pdiffusion 143 -48 143 -48 0 feedthrough
rlabel pdiffusion 150 -48 150 -48 0 cellNo=255
rlabel pdiffusion 157 -48 157 -48 0 feedthrough
rlabel pdiffusion 164 -48 164 -48 0 feedthrough
rlabel pdiffusion 171 -48 171 -48 0 cellNo=571
rlabel pdiffusion 178 -48 178 -48 0 feedthrough
rlabel pdiffusion 185 -48 185 -48 0 feedthrough
rlabel pdiffusion 192 -48 192 -48 0 cellNo=644
rlabel pdiffusion 199 -48 199 -48 0 feedthrough
rlabel pdiffusion 206 -48 206 -48 0 cellNo=282
rlabel pdiffusion 213 -48 213 -48 0 feedthrough
rlabel pdiffusion 220 -48 220 -48 0 cellNo=87
rlabel pdiffusion 227 -48 227 -48 0 cellNo=744
rlabel pdiffusion 234 -48 234 -48 0 feedthrough
rlabel pdiffusion 241 -48 241 -48 0 feedthrough
rlabel pdiffusion 248 -48 248 -48 0 feedthrough
rlabel pdiffusion 255 -48 255 -48 0 cellNo=376
rlabel pdiffusion 262 -48 262 -48 0 feedthrough
rlabel pdiffusion 269 -48 269 -48 0 feedthrough
rlabel pdiffusion 276 -48 276 -48 0 feedthrough
rlabel pdiffusion 283 -48 283 -48 0 feedthrough
rlabel pdiffusion 290 -48 290 -48 0 feedthrough
rlabel pdiffusion 297 -48 297 -48 0 feedthrough
rlabel pdiffusion 304 -48 304 -48 0 feedthrough
rlabel pdiffusion 311 -48 311 -48 0 feedthrough
rlabel pdiffusion 318 -48 318 -48 0 feedthrough
rlabel pdiffusion 325 -48 325 -48 0 feedthrough
rlabel pdiffusion 332 -48 332 -48 0 cellNo=356
rlabel pdiffusion 339 -48 339 -48 0 cellNo=90
rlabel pdiffusion 346 -48 346 -48 0 feedthrough
rlabel pdiffusion 353 -48 353 -48 0 feedthrough
rlabel pdiffusion 360 -48 360 -48 0 feedthrough
rlabel pdiffusion 367 -48 367 -48 0 feedthrough
rlabel pdiffusion 374 -48 374 -48 0 feedthrough
rlabel pdiffusion 381 -48 381 -48 0 feedthrough
rlabel pdiffusion 388 -48 388 -48 0 cellNo=61
rlabel pdiffusion 395 -48 395 -48 0 cellNo=800
rlabel pdiffusion 402 -48 402 -48 0 feedthrough
rlabel pdiffusion 409 -48 409 -48 0 feedthrough
rlabel pdiffusion 423 -48 423 -48 0 cellNo=66
rlabel pdiffusion 430 -48 430 -48 0 feedthrough
rlabel pdiffusion 437 -48 437 -48 0 feedthrough
rlabel pdiffusion 444 -48 444 -48 0 cellNo=128
rlabel pdiffusion 451 -48 451 -48 0 feedthrough
rlabel pdiffusion 458 -48 458 -48 0 feedthrough
rlabel pdiffusion 472 -48 472 -48 0 feedthrough
rlabel pdiffusion 479 -48 479 -48 0 feedthrough
rlabel pdiffusion 486 -48 486 -48 0 feedthrough
rlabel pdiffusion 500 -48 500 -48 0 feedthrough
rlabel pdiffusion 514 -48 514 -48 0 feedthrough
rlabel pdiffusion 535 -48 535 -48 0 cellNo=454
rlabel pdiffusion 542 -48 542 -48 0 cellNo=235
rlabel pdiffusion 549 -48 549 -48 0 feedthrough
rlabel pdiffusion 556 -48 556 -48 0 feedthrough
rlabel pdiffusion 563 -48 563 -48 0 feedthrough
rlabel pdiffusion 570 -48 570 -48 0 cellNo=82
rlabel pdiffusion 577 -48 577 -48 0 feedthrough
rlabel pdiffusion 584 -48 584 -48 0 feedthrough
rlabel pdiffusion 591 -48 591 -48 0 cellNo=250
rlabel pdiffusion 598 -48 598 -48 0 feedthrough
rlabel pdiffusion 605 -48 605 -48 0 feedthrough
rlabel pdiffusion 612 -48 612 -48 0 feedthrough
rlabel pdiffusion 626 -48 626 -48 0 feedthrough
rlabel pdiffusion 633 -48 633 -48 0 feedthrough
rlabel pdiffusion 647 -48 647 -48 0 cellNo=265
rlabel pdiffusion 654 -48 654 -48 0 cellNo=607
rlabel pdiffusion 661 -48 661 -48 0 feedthrough
rlabel pdiffusion 689 -48 689 -48 0 feedthrough
rlabel pdiffusion 731 -48 731 -48 0 feedthrough
rlabel pdiffusion 787 -48 787 -48 0 feedthrough
rlabel pdiffusion 808 -48 808 -48 0 feedthrough
rlabel pdiffusion 815 -48 815 -48 0 cellNo=398
rlabel pdiffusion 899 -48 899 -48 0 cellNo=64
rlabel pdiffusion 3 -87 3 -87 0 cellNo=91
rlabel pdiffusion 10 -87 10 -87 0 cellNo=228
rlabel pdiffusion 17 -87 17 -87 0 cellNo=683
rlabel pdiffusion 24 -87 24 -87 0 cellNo=438
rlabel pdiffusion 52 -87 52 -87 0 cellNo=97
rlabel pdiffusion 59 -87 59 -87 0 feedthrough
rlabel pdiffusion 66 -87 66 -87 0 feedthrough
rlabel pdiffusion 80 -87 80 -87 0 cellNo=490
rlabel pdiffusion 87 -87 87 -87 0 cellNo=116
rlabel pdiffusion 94 -87 94 -87 0 feedthrough
rlabel pdiffusion 101 -87 101 -87 0 cellNo=94
rlabel pdiffusion 108 -87 108 -87 0 cellNo=413
rlabel pdiffusion 115 -87 115 -87 0 feedthrough
rlabel pdiffusion 122 -87 122 -87 0 cellNo=238
rlabel pdiffusion 129 -87 129 -87 0 feedthrough
rlabel pdiffusion 136 -87 136 -87 0 feedthrough
rlabel pdiffusion 143 -87 143 -87 0 feedthrough
rlabel pdiffusion 150 -87 150 -87 0 feedthrough
rlabel pdiffusion 157 -87 157 -87 0 feedthrough
rlabel pdiffusion 164 -87 164 -87 0 feedthrough
rlabel pdiffusion 171 -87 171 -87 0 feedthrough
rlabel pdiffusion 178 -87 178 -87 0 cellNo=503
rlabel pdiffusion 185 -87 185 -87 0 cellNo=646
rlabel pdiffusion 192 -87 192 -87 0 feedthrough
rlabel pdiffusion 199 -87 199 -87 0 feedthrough
rlabel pdiffusion 206 -87 206 -87 0 cellNo=31
rlabel pdiffusion 213 -87 213 -87 0 feedthrough
rlabel pdiffusion 220 -87 220 -87 0 cellNo=117
rlabel pdiffusion 227 -87 227 -87 0 cellNo=640
rlabel pdiffusion 234 -87 234 -87 0 feedthrough
rlabel pdiffusion 241 -87 241 -87 0 feedthrough
rlabel pdiffusion 248 -87 248 -87 0 feedthrough
rlabel pdiffusion 255 -87 255 -87 0 feedthrough
rlabel pdiffusion 262 -87 262 -87 0 feedthrough
rlabel pdiffusion 269 -87 269 -87 0 feedthrough
rlabel pdiffusion 276 -87 276 -87 0 cellNo=417
rlabel pdiffusion 283 -87 283 -87 0 feedthrough
rlabel pdiffusion 290 -87 290 -87 0 feedthrough
rlabel pdiffusion 297 -87 297 -87 0 cellNo=443
rlabel pdiffusion 304 -87 304 -87 0 feedthrough
rlabel pdiffusion 311 -87 311 -87 0 feedthrough
rlabel pdiffusion 318 -87 318 -87 0 feedthrough
rlabel pdiffusion 325 -87 325 -87 0 feedthrough
rlabel pdiffusion 332 -87 332 -87 0 feedthrough
rlabel pdiffusion 339 -87 339 -87 0 feedthrough
rlabel pdiffusion 346 -87 346 -87 0 feedthrough
rlabel pdiffusion 353 -87 353 -87 0 feedthrough
rlabel pdiffusion 360 -87 360 -87 0 cellNo=543
rlabel pdiffusion 367 -87 367 -87 0 feedthrough
rlabel pdiffusion 374 -87 374 -87 0 feedthrough
rlabel pdiffusion 381 -87 381 -87 0 feedthrough
rlabel pdiffusion 388 -87 388 -87 0 feedthrough
rlabel pdiffusion 395 -87 395 -87 0 cellNo=57
rlabel pdiffusion 402 -87 402 -87 0 feedthrough
rlabel pdiffusion 409 -87 409 -87 0 feedthrough
rlabel pdiffusion 416 -87 416 -87 0 feedthrough
rlabel pdiffusion 423 -87 423 -87 0 feedthrough
rlabel pdiffusion 430 -87 430 -87 0 feedthrough
rlabel pdiffusion 437 -87 437 -87 0 cellNo=218
rlabel pdiffusion 444 -87 444 -87 0 cellNo=225
rlabel pdiffusion 451 -87 451 -87 0 feedthrough
rlabel pdiffusion 458 -87 458 -87 0 cellNo=174
rlabel pdiffusion 465 -87 465 -87 0 cellNo=803
rlabel pdiffusion 472 -87 472 -87 0 cellNo=81
rlabel pdiffusion 479 -87 479 -87 0 feedthrough
rlabel pdiffusion 486 -87 486 -87 0 feedthrough
rlabel pdiffusion 493 -87 493 -87 0 cellNo=407
rlabel pdiffusion 500 -87 500 -87 0 feedthrough
rlabel pdiffusion 507 -87 507 -87 0 feedthrough
rlabel pdiffusion 514 -87 514 -87 0 feedthrough
rlabel pdiffusion 521 -87 521 -87 0 feedthrough
rlabel pdiffusion 528 -87 528 -87 0 cellNo=118
rlabel pdiffusion 535 -87 535 -87 0 feedthrough
rlabel pdiffusion 542 -87 542 -87 0 feedthrough
rlabel pdiffusion 549 -87 549 -87 0 feedthrough
rlabel pdiffusion 556 -87 556 -87 0 feedthrough
rlabel pdiffusion 563 -87 563 -87 0 feedthrough
rlabel pdiffusion 570 -87 570 -87 0 feedthrough
rlabel pdiffusion 577 -87 577 -87 0 feedthrough
rlabel pdiffusion 584 -87 584 -87 0 feedthrough
rlabel pdiffusion 591 -87 591 -87 0 feedthrough
rlabel pdiffusion 598 -87 598 -87 0 feedthrough
rlabel pdiffusion 605 -87 605 -87 0 feedthrough
rlabel pdiffusion 612 -87 612 -87 0 feedthrough
rlabel pdiffusion 619 -87 619 -87 0 feedthrough
rlabel pdiffusion 626 -87 626 -87 0 feedthrough
rlabel pdiffusion 633 -87 633 -87 0 cellNo=378
rlabel pdiffusion 640 -87 640 -87 0 feedthrough
rlabel pdiffusion 647 -87 647 -87 0 feedthrough
rlabel pdiffusion 654 -87 654 -87 0 feedthrough
rlabel pdiffusion 661 -87 661 -87 0 feedthrough
rlabel pdiffusion 675 -87 675 -87 0 feedthrough
rlabel pdiffusion 682 -87 682 -87 0 cellNo=277
rlabel pdiffusion 703 -87 703 -87 0 feedthrough
rlabel pdiffusion 731 -87 731 -87 0 feedthrough
rlabel pdiffusion 794 -87 794 -87 0 feedthrough
rlabel pdiffusion 808 -87 808 -87 0 feedthrough
rlabel pdiffusion 899 -87 899 -87 0 feedthrough
rlabel pdiffusion 976 -87 976 -87 0 cellNo=108
rlabel pdiffusion 1088 -87 1088 -87 0 feedthrough
rlabel pdiffusion 1095 -87 1095 -87 0 cellNo=368
rlabel pdiffusion 3 -124 3 -124 0 cellNo=121
rlabel pdiffusion 10 -124 10 -124 0 cellNo=195
rlabel pdiffusion 17 -124 17 -124 0 cellNo=148
rlabel pdiffusion 24 -124 24 -124 0 cellNo=233
rlabel pdiffusion 31 -124 31 -124 0 feedthrough
rlabel pdiffusion 38 -124 38 -124 0 cellNo=335
rlabel pdiffusion 45 -124 45 -124 0 cellNo=20
rlabel pdiffusion 52 -124 52 -124 0 feedthrough
rlabel pdiffusion 59 -124 59 -124 0 feedthrough
rlabel pdiffusion 66 -124 66 -124 0 feedthrough
rlabel pdiffusion 73 -124 73 -124 0 cellNo=441
rlabel pdiffusion 94 -124 94 -124 0 feedthrough
rlabel pdiffusion 101 -124 101 -124 0 feedthrough
rlabel pdiffusion 108 -124 108 -124 0 feedthrough
rlabel pdiffusion 115 -124 115 -124 0 cellNo=566
rlabel pdiffusion 122 -124 122 -124 0 feedthrough
rlabel pdiffusion 129 -124 129 -124 0 feedthrough
rlabel pdiffusion 136 -124 136 -124 0 cellNo=768
rlabel pdiffusion 143 -124 143 -124 0 feedthrough
rlabel pdiffusion 150 -124 150 -124 0 feedthrough
rlabel pdiffusion 157 -124 157 -124 0 feedthrough
rlabel pdiffusion 164 -124 164 -124 0 feedthrough
rlabel pdiffusion 171 -124 171 -124 0 feedthrough
rlabel pdiffusion 178 -124 178 -124 0 cellNo=689
rlabel pdiffusion 185 -124 185 -124 0 cellNo=243
rlabel pdiffusion 192 -124 192 -124 0 feedthrough
rlabel pdiffusion 199 -124 199 -124 0 feedthrough
rlabel pdiffusion 206 -124 206 -124 0 feedthrough
rlabel pdiffusion 213 -124 213 -124 0 feedthrough
rlabel pdiffusion 220 -124 220 -124 0 feedthrough
rlabel pdiffusion 227 -124 227 -124 0 cellNo=793
rlabel pdiffusion 234 -124 234 -124 0 feedthrough
rlabel pdiffusion 241 -124 241 -124 0 cellNo=146
rlabel pdiffusion 248 -124 248 -124 0 cellNo=196
rlabel pdiffusion 255 -124 255 -124 0 feedthrough
rlabel pdiffusion 262 -124 262 -124 0 feedthrough
rlabel pdiffusion 269 -124 269 -124 0 feedthrough
rlabel pdiffusion 276 -124 276 -124 0 feedthrough
rlabel pdiffusion 283 -124 283 -124 0 feedthrough
rlabel pdiffusion 290 -124 290 -124 0 cellNo=712
rlabel pdiffusion 297 -124 297 -124 0 cellNo=534
rlabel pdiffusion 304 -124 304 -124 0 feedthrough
rlabel pdiffusion 311 -124 311 -124 0 feedthrough
rlabel pdiffusion 318 -124 318 -124 0 feedthrough
rlabel pdiffusion 325 -124 325 -124 0 cellNo=654
rlabel pdiffusion 332 -124 332 -124 0 feedthrough
rlabel pdiffusion 339 -124 339 -124 0 feedthrough
rlabel pdiffusion 346 -124 346 -124 0 feedthrough
rlabel pdiffusion 353 -124 353 -124 0 cellNo=404
rlabel pdiffusion 360 -124 360 -124 0 feedthrough
rlabel pdiffusion 367 -124 367 -124 0 feedthrough
rlabel pdiffusion 374 -124 374 -124 0 cellNo=343
rlabel pdiffusion 381 -124 381 -124 0 cellNo=44
rlabel pdiffusion 388 -124 388 -124 0 feedthrough
rlabel pdiffusion 395 -124 395 -124 0 feedthrough
rlabel pdiffusion 402 -124 402 -124 0 feedthrough
rlabel pdiffusion 409 -124 409 -124 0 cellNo=564
rlabel pdiffusion 416 -124 416 -124 0 feedthrough
rlabel pdiffusion 423 -124 423 -124 0 feedthrough
rlabel pdiffusion 430 -124 430 -124 0 feedthrough
rlabel pdiffusion 437 -124 437 -124 0 feedthrough
rlabel pdiffusion 444 -124 444 -124 0 feedthrough
rlabel pdiffusion 451 -124 451 -124 0 feedthrough
rlabel pdiffusion 458 -124 458 -124 0 feedthrough
rlabel pdiffusion 465 -124 465 -124 0 cellNo=718
rlabel pdiffusion 472 -124 472 -124 0 feedthrough
rlabel pdiffusion 479 -124 479 -124 0 cellNo=807
rlabel pdiffusion 486 -124 486 -124 0 feedthrough
rlabel pdiffusion 493 -124 493 -124 0 feedthrough
rlabel pdiffusion 500 -124 500 -124 0 feedthrough
rlabel pdiffusion 507 -124 507 -124 0 cellNo=198
rlabel pdiffusion 514 -124 514 -124 0 feedthrough
rlabel pdiffusion 521 -124 521 -124 0 feedthrough
rlabel pdiffusion 528 -124 528 -124 0 feedthrough
rlabel pdiffusion 535 -124 535 -124 0 feedthrough
rlabel pdiffusion 542 -124 542 -124 0 feedthrough
rlabel pdiffusion 549 -124 549 -124 0 cellNo=680
rlabel pdiffusion 556 -124 556 -124 0 cellNo=229
rlabel pdiffusion 563 -124 563 -124 0 feedthrough
rlabel pdiffusion 570 -124 570 -124 0 feedthrough
rlabel pdiffusion 577 -124 577 -124 0 feedthrough
rlabel pdiffusion 584 -124 584 -124 0 feedthrough
rlabel pdiffusion 591 -124 591 -124 0 cellNo=748
rlabel pdiffusion 598 -124 598 -124 0 feedthrough
rlabel pdiffusion 605 -124 605 -124 0 feedthrough
rlabel pdiffusion 612 -124 612 -124 0 feedthrough
rlabel pdiffusion 619 -124 619 -124 0 feedthrough
rlabel pdiffusion 626 -124 626 -124 0 feedthrough
rlabel pdiffusion 633 -124 633 -124 0 feedthrough
rlabel pdiffusion 640 -124 640 -124 0 feedthrough
rlabel pdiffusion 647 -124 647 -124 0 feedthrough
rlabel pdiffusion 654 -124 654 -124 0 cellNo=613
rlabel pdiffusion 661 -124 661 -124 0 feedthrough
rlabel pdiffusion 668 -124 668 -124 0 feedthrough
rlabel pdiffusion 675 -124 675 -124 0 feedthrough
rlabel pdiffusion 682 -124 682 -124 0 feedthrough
rlabel pdiffusion 689 -124 689 -124 0 feedthrough
rlabel pdiffusion 696 -124 696 -124 0 feedthrough
rlabel pdiffusion 703 -124 703 -124 0 feedthrough
rlabel pdiffusion 710 -124 710 -124 0 cellNo=524
rlabel pdiffusion 717 -124 717 -124 0 feedthrough
rlabel pdiffusion 724 -124 724 -124 0 feedthrough
rlabel pdiffusion 731 -124 731 -124 0 feedthrough
rlabel pdiffusion 738 -124 738 -124 0 feedthrough
rlabel pdiffusion 759 -124 759 -124 0 cellNo=528
rlabel pdiffusion 766 -124 766 -124 0 feedthrough
rlabel pdiffusion 780 -124 780 -124 0 feedthrough
rlabel pdiffusion 801 -124 801 -124 0 feedthrough
rlabel pdiffusion 906 -124 906 -124 0 feedthrough
rlabel pdiffusion 976 -124 976 -124 0 feedthrough
rlabel pdiffusion 1088 -124 1088 -124 0 feedthrough
rlabel pdiffusion 3 -185 3 -185 0 cellNo=267
rlabel pdiffusion 10 -185 10 -185 0 cellNo=827
rlabel pdiffusion 24 -185 24 -185 0 feedthrough
rlabel pdiffusion 31 -185 31 -185 0 feedthrough
rlabel pdiffusion 38 -185 38 -185 0 cellNo=332
rlabel pdiffusion 45 -185 45 -185 0 cellNo=251
rlabel pdiffusion 52 -185 52 -185 0 feedthrough
rlabel pdiffusion 59 -185 59 -185 0 feedthrough
rlabel pdiffusion 66 -185 66 -185 0 cellNo=596
rlabel pdiffusion 73 -185 73 -185 0 feedthrough
rlabel pdiffusion 80 -185 80 -185 0 feedthrough
rlabel pdiffusion 87 -185 87 -185 0 cellNo=176
rlabel pdiffusion 94 -185 94 -185 0 feedthrough
rlabel pdiffusion 101 -185 101 -185 0 feedthrough
rlabel pdiffusion 108 -185 108 -185 0 feedthrough
rlabel pdiffusion 115 -185 115 -185 0 feedthrough
rlabel pdiffusion 122 -185 122 -185 0 feedthrough
rlabel pdiffusion 129 -185 129 -185 0 feedthrough
rlabel pdiffusion 136 -185 136 -185 0 cellNo=258
rlabel pdiffusion 143 -185 143 -185 0 feedthrough
rlabel pdiffusion 150 -185 150 -185 0 feedthrough
rlabel pdiffusion 157 -185 157 -185 0 cellNo=620
rlabel pdiffusion 164 -185 164 -185 0 cellNo=179
rlabel pdiffusion 171 -185 171 -185 0 feedthrough
rlabel pdiffusion 178 -185 178 -185 0 feedthrough
rlabel pdiffusion 185 -185 185 -185 0 cellNo=635
rlabel pdiffusion 192 -185 192 -185 0 feedthrough
rlabel pdiffusion 199 -185 199 -185 0 cellNo=457
rlabel pdiffusion 206 -185 206 -185 0 cellNo=339
rlabel pdiffusion 213 -185 213 -185 0 feedthrough
rlabel pdiffusion 220 -185 220 -185 0 feedthrough
rlabel pdiffusion 227 -185 227 -185 0 feedthrough
rlabel pdiffusion 234 -185 234 -185 0 feedthrough
rlabel pdiffusion 241 -185 241 -185 0 feedthrough
rlabel pdiffusion 248 -185 248 -185 0 feedthrough
rlabel pdiffusion 255 -185 255 -185 0 feedthrough
rlabel pdiffusion 262 -185 262 -185 0 feedthrough
rlabel pdiffusion 269 -185 269 -185 0 feedthrough
rlabel pdiffusion 276 -185 276 -185 0 feedthrough
rlabel pdiffusion 283 -185 283 -185 0 feedthrough
rlabel pdiffusion 290 -185 290 -185 0 feedthrough
rlabel pdiffusion 297 -185 297 -185 0 feedthrough
rlabel pdiffusion 304 -185 304 -185 0 feedthrough
rlabel pdiffusion 311 -185 311 -185 0 feedthrough
rlabel pdiffusion 318 -185 318 -185 0 cellNo=180
rlabel pdiffusion 325 -185 325 -185 0 feedthrough
rlabel pdiffusion 332 -185 332 -185 0 cellNo=653
rlabel pdiffusion 339 -185 339 -185 0 cellNo=711
rlabel pdiffusion 346 -185 346 -185 0 cellNo=745
rlabel pdiffusion 353 -185 353 -185 0 feedthrough
rlabel pdiffusion 360 -185 360 -185 0 feedthrough
rlabel pdiffusion 367 -185 367 -185 0 feedthrough
rlabel pdiffusion 374 -185 374 -185 0 cellNo=519
rlabel pdiffusion 381 -185 381 -185 0 feedthrough
rlabel pdiffusion 388 -185 388 -185 0 cellNo=129
rlabel pdiffusion 395 -185 395 -185 0 feedthrough
rlabel pdiffusion 402 -185 402 -185 0 feedthrough
rlabel pdiffusion 409 -185 409 -185 0 feedthrough
rlabel pdiffusion 416 -185 416 -185 0 feedthrough
rlabel pdiffusion 423 -185 423 -185 0 cellNo=491
rlabel pdiffusion 430 -185 430 -185 0 feedthrough
rlabel pdiffusion 437 -185 437 -185 0 feedthrough
rlabel pdiffusion 444 -185 444 -185 0 feedthrough
rlabel pdiffusion 451 -185 451 -185 0 feedthrough
rlabel pdiffusion 458 -185 458 -185 0 feedthrough
rlabel pdiffusion 465 -185 465 -185 0 cellNo=190
rlabel pdiffusion 472 -185 472 -185 0 feedthrough
rlabel pdiffusion 479 -185 479 -185 0 feedthrough
rlabel pdiffusion 486 -185 486 -185 0 cellNo=790
rlabel pdiffusion 493 -185 493 -185 0 cellNo=448
rlabel pdiffusion 500 -185 500 -185 0 feedthrough
rlabel pdiffusion 507 -185 507 -185 0 feedthrough
rlabel pdiffusion 514 -185 514 -185 0 feedthrough
rlabel pdiffusion 521 -185 521 -185 0 cellNo=285
rlabel pdiffusion 528 -185 528 -185 0 feedthrough
rlabel pdiffusion 535 -185 535 -185 0 cellNo=352
rlabel pdiffusion 542 -185 542 -185 0 feedthrough
rlabel pdiffusion 549 -185 549 -185 0 feedthrough
rlabel pdiffusion 556 -185 556 -185 0 feedthrough
rlabel pdiffusion 563 -185 563 -185 0 feedthrough
rlabel pdiffusion 570 -185 570 -185 0 feedthrough
rlabel pdiffusion 577 -185 577 -185 0 feedthrough
rlabel pdiffusion 584 -185 584 -185 0 feedthrough
rlabel pdiffusion 591 -185 591 -185 0 feedthrough
rlabel pdiffusion 598 -185 598 -185 0 feedthrough
rlabel pdiffusion 605 -185 605 -185 0 feedthrough
rlabel pdiffusion 612 -185 612 -185 0 feedthrough
rlabel pdiffusion 619 -185 619 -185 0 feedthrough
rlabel pdiffusion 626 -185 626 -185 0 feedthrough
rlabel pdiffusion 633 -185 633 -185 0 feedthrough
rlabel pdiffusion 640 -185 640 -185 0 feedthrough
rlabel pdiffusion 647 -185 647 -185 0 feedthrough
rlabel pdiffusion 654 -185 654 -185 0 feedthrough
rlabel pdiffusion 661 -185 661 -185 0 feedthrough
rlabel pdiffusion 668 -185 668 -185 0 feedthrough
rlabel pdiffusion 675 -185 675 -185 0 feedthrough
rlabel pdiffusion 682 -185 682 -185 0 feedthrough
rlabel pdiffusion 689 -185 689 -185 0 feedthrough
rlabel pdiffusion 696 -185 696 -185 0 feedthrough
rlabel pdiffusion 703 -185 703 -185 0 feedthrough
rlabel pdiffusion 710 -185 710 -185 0 feedthrough
rlabel pdiffusion 717 -185 717 -185 0 feedthrough
rlabel pdiffusion 724 -185 724 -185 0 feedthrough
rlabel pdiffusion 731 -185 731 -185 0 feedthrough
rlabel pdiffusion 738 -185 738 -185 0 feedthrough
rlabel pdiffusion 745 -185 745 -185 0 feedthrough
rlabel pdiffusion 752 -185 752 -185 0 feedthrough
rlabel pdiffusion 759 -185 759 -185 0 feedthrough
rlabel pdiffusion 766 -185 766 -185 0 feedthrough
rlabel pdiffusion 773 -185 773 -185 0 feedthrough
rlabel pdiffusion 780 -185 780 -185 0 feedthrough
rlabel pdiffusion 787 -185 787 -185 0 feedthrough
rlabel pdiffusion 794 -185 794 -185 0 feedthrough
rlabel pdiffusion 801 -185 801 -185 0 feedthrough
rlabel pdiffusion 808 -185 808 -185 0 feedthrough
rlabel pdiffusion 815 -185 815 -185 0 cellNo=216
rlabel pdiffusion 822 -185 822 -185 0 cellNo=369
rlabel pdiffusion 829 -185 829 -185 0 cellNo=439
rlabel pdiffusion 836 -185 836 -185 0 cellNo=501
rlabel pdiffusion 843 -185 843 -185 0 cellNo=527
rlabel pdiffusion 850 -185 850 -185 0 feedthrough
rlabel pdiffusion 857 -185 857 -185 0 cellNo=575
rlabel pdiffusion 920 -185 920 -185 0 feedthrough
rlabel pdiffusion 976 -185 976 -185 0 feedthrough
rlabel pdiffusion 1088 -185 1088 -185 0 feedthrough
rlabel pdiffusion 3 -244 3 -244 0 cellNo=109
rlabel pdiffusion 10 -244 10 -244 0 cellNo=795
rlabel pdiffusion 17 -244 17 -244 0 feedthrough
rlabel pdiffusion 24 -244 24 -244 0 feedthrough
rlabel pdiffusion 31 -244 31 -244 0 feedthrough
rlabel pdiffusion 38 -244 38 -244 0 feedthrough
rlabel pdiffusion 45 -244 45 -244 0 feedthrough
rlabel pdiffusion 52 -244 52 -244 0 feedthrough
rlabel pdiffusion 59 -244 59 -244 0 cellNo=161
rlabel pdiffusion 66 -244 66 -244 0 cellNo=220
rlabel pdiffusion 73 -244 73 -244 0 feedthrough
rlabel pdiffusion 80 -244 80 -244 0 feedthrough
rlabel pdiffusion 87 -244 87 -244 0 cellNo=562
rlabel pdiffusion 94 -244 94 -244 0 cellNo=759
rlabel pdiffusion 101 -244 101 -244 0 cellNo=55
rlabel pdiffusion 108 -244 108 -244 0 cellNo=535
rlabel pdiffusion 115 -244 115 -244 0 cellNo=240
rlabel pdiffusion 122 -244 122 -244 0 feedthrough
rlabel pdiffusion 129 -244 129 -244 0 feedthrough
rlabel pdiffusion 136 -244 136 -244 0 feedthrough
rlabel pdiffusion 143 -244 143 -244 0 feedthrough
rlabel pdiffusion 150 -244 150 -244 0 feedthrough
rlabel pdiffusion 157 -244 157 -244 0 cellNo=623
rlabel pdiffusion 164 -244 164 -244 0 feedthrough
rlabel pdiffusion 171 -244 171 -244 0 cellNo=142
rlabel pdiffusion 178 -244 178 -244 0 feedthrough
rlabel pdiffusion 185 -244 185 -244 0 cellNo=860
rlabel pdiffusion 192 -244 192 -244 0 feedthrough
rlabel pdiffusion 199 -244 199 -244 0 cellNo=338
rlabel pdiffusion 206 -244 206 -244 0 feedthrough
rlabel pdiffusion 213 -244 213 -244 0 feedthrough
rlabel pdiffusion 220 -244 220 -244 0 cellNo=296
rlabel pdiffusion 227 -244 227 -244 0 cellNo=787
rlabel pdiffusion 234 -244 234 -244 0 feedthrough
rlabel pdiffusion 241 -244 241 -244 0 feedthrough
rlabel pdiffusion 248 -244 248 -244 0 feedthrough
rlabel pdiffusion 255 -244 255 -244 0 feedthrough
rlabel pdiffusion 262 -244 262 -244 0 cellNo=738
rlabel pdiffusion 269 -244 269 -244 0 feedthrough
rlabel pdiffusion 276 -244 276 -244 0 feedthrough
rlabel pdiffusion 283 -244 283 -244 0 cellNo=597
rlabel pdiffusion 290 -244 290 -244 0 cellNo=643
rlabel pdiffusion 297 -244 297 -244 0 feedthrough
rlabel pdiffusion 304 -244 304 -244 0 feedthrough
rlabel pdiffusion 311 -244 311 -244 0 feedthrough
rlabel pdiffusion 318 -244 318 -244 0 feedthrough
rlabel pdiffusion 325 -244 325 -244 0 feedthrough
rlabel pdiffusion 332 -244 332 -244 0 feedthrough
rlabel pdiffusion 339 -244 339 -244 0 feedthrough
rlabel pdiffusion 346 -244 346 -244 0 feedthrough
rlabel pdiffusion 353 -244 353 -244 0 cellNo=215
rlabel pdiffusion 360 -244 360 -244 0 feedthrough
rlabel pdiffusion 367 -244 367 -244 0 feedthrough
rlabel pdiffusion 374 -244 374 -244 0 feedthrough
rlabel pdiffusion 381 -244 381 -244 0 cellNo=395
rlabel pdiffusion 388 -244 388 -244 0 feedthrough
rlabel pdiffusion 395 -244 395 -244 0 feedthrough
rlabel pdiffusion 402 -244 402 -244 0 feedthrough
rlabel pdiffusion 409 -244 409 -244 0 feedthrough
rlabel pdiffusion 416 -244 416 -244 0 feedthrough
rlabel pdiffusion 423 -244 423 -244 0 feedthrough
rlabel pdiffusion 430 -244 430 -244 0 feedthrough
rlabel pdiffusion 437 -244 437 -244 0 feedthrough
rlabel pdiffusion 444 -244 444 -244 0 feedthrough
rlabel pdiffusion 451 -244 451 -244 0 feedthrough
rlabel pdiffusion 458 -244 458 -244 0 cellNo=320
rlabel pdiffusion 465 -244 465 -244 0 cellNo=152
rlabel pdiffusion 472 -244 472 -244 0 feedthrough
rlabel pdiffusion 479 -244 479 -244 0 cellNo=856
rlabel pdiffusion 486 -244 486 -244 0 cellNo=230
rlabel pdiffusion 493 -244 493 -244 0 cellNo=85
rlabel pdiffusion 500 -244 500 -244 0 feedthrough
rlabel pdiffusion 507 -244 507 -244 0 feedthrough
rlabel pdiffusion 514 -244 514 -244 0 feedthrough
rlabel pdiffusion 521 -244 521 -244 0 feedthrough
rlabel pdiffusion 528 -244 528 -244 0 feedthrough
rlabel pdiffusion 535 -244 535 -244 0 feedthrough
rlabel pdiffusion 542 -244 542 -244 0 feedthrough
rlabel pdiffusion 549 -244 549 -244 0 feedthrough
rlabel pdiffusion 556 -244 556 -244 0 feedthrough
rlabel pdiffusion 563 -244 563 -244 0 feedthrough
rlabel pdiffusion 570 -244 570 -244 0 feedthrough
rlabel pdiffusion 577 -244 577 -244 0 feedthrough
rlabel pdiffusion 584 -244 584 -244 0 feedthrough
rlabel pdiffusion 591 -244 591 -244 0 cellNo=56
rlabel pdiffusion 598 -244 598 -244 0 cellNo=419
rlabel pdiffusion 605 -244 605 -244 0 feedthrough
rlabel pdiffusion 612 -244 612 -244 0 feedthrough
rlabel pdiffusion 619 -244 619 -244 0 feedthrough
rlabel pdiffusion 626 -244 626 -244 0 feedthrough
rlabel pdiffusion 633 -244 633 -244 0 feedthrough
rlabel pdiffusion 640 -244 640 -244 0 feedthrough
rlabel pdiffusion 647 -244 647 -244 0 cellNo=760
rlabel pdiffusion 654 -244 654 -244 0 feedthrough
rlabel pdiffusion 661 -244 661 -244 0 feedthrough
rlabel pdiffusion 668 -244 668 -244 0 feedthrough
rlabel pdiffusion 675 -244 675 -244 0 feedthrough
rlabel pdiffusion 682 -244 682 -244 0 feedthrough
rlabel pdiffusion 689 -244 689 -244 0 feedthrough
rlabel pdiffusion 696 -244 696 -244 0 feedthrough
rlabel pdiffusion 703 -244 703 -244 0 feedthrough
rlabel pdiffusion 710 -244 710 -244 0 feedthrough
rlabel pdiffusion 717 -244 717 -244 0 feedthrough
rlabel pdiffusion 724 -244 724 -244 0 feedthrough
rlabel pdiffusion 731 -244 731 -244 0 feedthrough
rlabel pdiffusion 738 -244 738 -244 0 feedthrough
rlabel pdiffusion 745 -244 745 -244 0 feedthrough
rlabel pdiffusion 752 -244 752 -244 0 feedthrough
rlabel pdiffusion 759 -244 759 -244 0 feedthrough
rlabel pdiffusion 766 -244 766 -244 0 feedthrough
rlabel pdiffusion 773 -244 773 -244 0 feedthrough
rlabel pdiffusion 780 -244 780 -244 0 feedthrough
rlabel pdiffusion 787 -244 787 -244 0 feedthrough
rlabel pdiffusion 794 -244 794 -244 0 feedthrough
rlabel pdiffusion 801 -244 801 -244 0 cellNo=736
rlabel pdiffusion 808 -244 808 -244 0 feedthrough
rlabel pdiffusion 815 -244 815 -244 0 feedthrough
rlabel pdiffusion 822 -244 822 -244 0 feedthrough
rlabel pdiffusion 829 -244 829 -244 0 feedthrough
rlabel pdiffusion 836 -244 836 -244 0 feedthrough
rlabel pdiffusion 843 -244 843 -244 0 feedthrough
rlabel pdiffusion 850 -244 850 -244 0 feedthrough
rlabel pdiffusion 857 -244 857 -244 0 feedthrough
rlabel pdiffusion 864 -244 864 -244 0 feedthrough
rlabel pdiffusion 871 -244 871 -244 0 feedthrough
rlabel pdiffusion 878 -244 878 -244 0 feedthrough
rlabel pdiffusion 885 -244 885 -244 0 feedthrough
rlabel pdiffusion 892 -244 892 -244 0 feedthrough
rlabel pdiffusion 899 -244 899 -244 0 feedthrough
rlabel pdiffusion 906 -244 906 -244 0 feedthrough
rlabel pdiffusion 913 -244 913 -244 0 feedthrough
rlabel pdiffusion 920 -244 920 -244 0 feedthrough
rlabel pdiffusion 927 -244 927 -244 0 feedthrough
rlabel pdiffusion 934 -244 934 -244 0 feedthrough
rlabel pdiffusion 941 -244 941 -244 0 feedthrough
rlabel pdiffusion 948 -244 948 -244 0 feedthrough
rlabel pdiffusion 955 -244 955 -244 0 cellNo=725
rlabel pdiffusion 976 -244 976 -244 0 feedthrough
rlabel pdiffusion 1088 -244 1088 -244 0 feedthrough
rlabel pdiffusion 3 -315 3 -315 0 cellNo=401
rlabel pdiffusion 10 -315 10 -315 0 cellNo=306
rlabel pdiffusion 17 -315 17 -315 0 feedthrough
rlabel pdiffusion 24 -315 24 -315 0 feedthrough
rlabel pdiffusion 31 -315 31 -315 0 cellNo=705
rlabel pdiffusion 38 -315 38 -315 0 feedthrough
rlabel pdiffusion 45 -315 45 -315 0 cellNo=304
rlabel pdiffusion 52 -315 52 -315 0 cellNo=473
rlabel pdiffusion 59 -315 59 -315 0 feedthrough
rlabel pdiffusion 66 -315 66 -315 0 feedthrough
rlabel pdiffusion 73 -315 73 -315 0 feedthrough
rlabel pdiffusion 80 -315 80 -315 0 cellNo=776
rlabel pdiffusion 87 -315 87 -315 0 feedthrough
rlabel pdiffusion 94 -315 94 -315 0 feedthrough
rlabel pdiffusion 101 -315 101 -315 0 feedthrough
rlabel pdiffusion 108 -315 108 -315 0 cellNo=274
rlabel pdiffusion 115 -315 115 -315 0 feedthrough
rlabel pdiffusion 122 -315 122 -315 0 feedthrough
rlabel pdiffusion 129 -315 129 -315 0 feedthrough
rlabel pdiffusion 136 -315 136 -315 0 feedthrough
rlabel pdiffusion 143 -315 143 -315 0 cellNo=728
rlabel pdiffusion 150 -315 150 -315 0 feedthrough
rlabel pdiffusion 157 -315 157 -315 0 feedthrough
rlabel pdiffusion 164 -315 164 -315 0 cellNo=254
rlabel pdiffusion 171 -315 171 -315 0 feedthrough
rlabel pdiffusion 178 -315 178 -315 0 feedthrough
rlabel pdiffusion 185 -315 185 -315 0 feedthrough
rlabel pdiffusion 192 -315 192 -315 0 cellNo=602
rlabel pdiffusion 199 -315 199 -315 0 feedthrough
rlabel pdiffusion 206 -315 206 -315 0 cellNo=170
rlabel pdiffusion 213 -315 213 -315 0 feedthrough
rlabel pdiffusion 220 -315 220 -315 0 feedthrough
rlabel pdiffusion 227 -315 227 -315 0 cellNo=266
rlabel pdiffusion 234 -315 234 -315 0 feedthrough
rlabel pdiffusion 241 -315 241 -315 0 feedthrough
rlabel pdiffusion 248 -315 248 -315 0 feedthrough
rlabel pdiffusion 255 -315 255 -315 0 feedthrough
rlabel pdiffusion 262 -315 262 -315 0 feedthrough
rlabel pdiffusion 269 -315 269 -315 0 feedthrough
rlabel pdiffusion 276 -315 276 -315 0 feedthrough
rlabel pdiffusion 283 -315 283 -315 0 feedthrough
rlabel pdiffusion 290 -315 290 -315 0 cellNo=150
rlabel pdiffusion 297 -315 297 -315 0 feedthrough
rlabel pdiffusion 304 -315 304 -315 0 feedthrough
rlabel pdiffusion 311 -315 311 -315 0 feedthrough
rlabel pdiffusion 318 -315 318 -315 0 feedthrough
rlabel pdiffusion 325 -315 325 -315 0 feedthrough
rlabel pdiffusion 332 -315 332 -315 0 feedthrough
rlabel pdiffusion 339 -315 339 -315 0 feedthrough
rlabel pdiffusion 346 -315 346 -315 0 feedthrough
rlabel pdiffusion 353 -315 353 -315 0 feedthrough
rlabel pdiffusion 360 -315 360 -315 0 feedthrough
rlabel pdiffusion 367 -315 367 -315 0 feedthrough
rlabel pdiffusion 374 -315 374 -315 0 feedthrough
rlabel pdiffusion 381 -315 381 -315 0 cellNo=525
rlabel pdiffusion 388 -315 388 -315 0 cellNo=102
rlabel pdiffusion 395 -315 395 -315 0 feedthrough
rlabel pdiffusion 402 -315 402 -315 0 feedthrough
rlabel pdiffusion 409 -315 409 -315 0 cellNo=248
rlabel pdiffusion 416 -315 416 -315 0 cellNo=539
rlabel pdiffusion 423 -315 423 -315 0 feedthrough
rlabel pdiffusion 430 -315 430 -315 0 feedthrough
rlabel pdiffusion 437 -315 437 -315 0 cellNo=734
rlabel pdiffusion 444 -315 444 -315 0 feedthrough
rlabel pdiffusion 451 -315 451 -315 0 feedthrough
rlabel pdiffusion 458 -315 458 -315 0 feedthrough
rlabel pdiffusion 465 -315 465 -315 0 cellNo=406
rlabel pdiffusion 472 -315 472 -315 0 cellNo=520
rlabel pdiffusion 479 -315 479 -315 0 feedthrough
rlabel pdiffusion 486 -315 486 -315 0 cellNo=194
rlabel pdiffusion 493 -315 493 -315 0 feedthrough
rlabel pdiffusion 500 -315 500 -315 0 feedthrough
rlabel pdiffusion 507 -315 507 -315 0 cellNo=606
rlabel pdiffusion 514 -315 514 -315 0 feedthrough
rlabel pdiffusion 521 -315 521 -315 0 feedthrough
rlabel pdiffusion 528 -315 528 -315 0 feedthrough
rlabel pdiffusion 535 -315 535 -315 0 feedthrough
rlabel pdiffusion 542 -315 542 -315 0 cellNo=43
rlabel pdiffusion 549 -315 549 -315 0 cellNo=98
rlabel pdiffusion 556 -315 556 -315 0 feedthrough
rlabel pdiffusion 563 -315 563 -315 0 feedthrough
rlabel pdiffusion 570 -315 570 -315 0 feedthrough
rlabel pdiffusion 577 -315 577 -315 0 cellNo=508
rlabel pdiffusion 584 -315 584 -315 0 cellNo=279
rlabel pdiffusion 591 -315 591 -315 0 feedthrough
rlabel pdiffusion 598 -315 598 -315 0 feedthrough
rlabel pdiffusion 605 -315 605 -315 0 feedthrough
rlabel pdiffusion 612 -315 612 -315 0 feedthrough
rlabel pdiffusion 619 -315 619 -315 0 feedthrough
rlabel pdiffusion 626 -315 626 -315 0 feedthrough
rlabel pdiffusion 633 -315 633 -315 0 feedthrough
rlabel pdiffusion 640 -315 640 -315 0 feedthrough
rlabel pdiffusion 647 -315 647 -315 0 feedthrough
rlabel pdiffusion 654 -315 654 -315 0 feedthrough
rlabel pdiffusion 661 -315 661 -315 0 feedthrough
rlabel pdiffusion 668 -315 668 -315 0 feedthrough
rlabel pdiffusion 675 -315 675 -315 0 feedthrough
rlabel pdiffusion 682 -315 682 -315 0 feedthrough
rlabel pdiffusion 689 -315 689 -315 0 feedthrough
rlabel pdiffusion 696 -315 696 -315 0 feedthrough
rlabel pdiffusion 703 -315 703 -315 0 feedthrough
rlabel pdiffusion 710 -315 710 -315 0 feedthrough
rlabel pdiffusion 717 -315 717 -315 0 cellNo=288
rlabel pdiffusion 724 -315 724 -315 0 feedthrough
rlabel pdiffusion 731 -315 731 -315 0 feedthrough
rlabel pdiffusion 738 -315 738 -315 0 feedthrough
rlabel pdiffusion 745 -315 745 -315 0 feedthrough
rlabel pdiffusion 752 -315 752 -315 0 feedthrough
rlabel pdiffusion 759 -315 759 -315 0 feedthrough
rlabel pdiffusion 766 -315 766 -315 0 feedthrough
rlabel pdiffusion 773 -315 773 -315 0 feedthrough
rlabel pdiffusion 780 -315 780 -315 0 feedthrough
rlabel pdiffusion 787 -315 787 -315 0 feedthrough
rlabel pdiffusion 794 -315 794 -315 0 feedthrough
rlabel pdiffusion 801 -315 801 -315 0 feedthrough
rlabel pdiffusion 808 -315 808 -315 0 feedthrough
rlabel pdiffusion 815 -315 815 -315 0 feedthrough
rlabel pdiffusion 822 -315 822 -315 0 feedthrough
rlabel pdiffusion 829 -315 829 -315 0 feedthrough
rlabel pdiffusion 836 -315 836 -315 0 feedthrough
rlabel pdiffusion 843 -315 843 -315 0 feedthrough
rlabel pdiffusion 850 -315 850 -315 0 feedthrough
rlabel pdiffusion 857 -315 857 -315 0 feedthrough
rlabel pdiffusion 864 -315 864 -315 0 feedthrough
rlabel pdiffusion 871 -315 871 -315 0 feedthrough
rlabel pdiffusion 878 -315 878 -315 0 feedthrough
rlabel pdiffusion 885 -315 885 -315 0 feedthrough
rlabel pdiffusion 892 -315 892 -315 0 feedthrough
rlabel pdiffusion 899 -315 899 -315 0 feedthrough
rlabel pdiffusion 906 -315 906 -315 0 feedthrough
rlabel pdiffusion 913 -315 913 -315 0 feedthrough
rlabel pdiffusion 920 -315 920 -315 0 feedthrough
rlabel pdiffusion 927 -315 927 -315 0 feedthrough
rlabel pdiffusion 934 -315 934 -315 0 cellNo=859
rlabel pdiffusion 941 -315 941 -315 0 feedthrough
rlabel pdiffusion 948 -315 948 -315 0 cellNo=211
rlabel pdiffusion 955 -315 955 -315 0 feedthrough
rlabel pdiffusion 962 -315 962 -315 0 feedthrough
rlabel pdiffusion 969 -315 969 -315 0 cellNo=302
rlabel pdiffusion 976 -315 976 -315 0 feedthrough
rlabel pdiffusion 983 -315 983 -315 0 feedthrough
rlabel pdiffusion 1095 -315 1095 -315 0 feedthrough
rlabel pdiffusion 3 -400 3 -400 0 cellNo=49
rlabel pdiffusion 17 -400 17 -400 0 feedthrough
rlabel pdiffusion 24 -400 24 -400 0 feedthrough
rlabel pdiffusion 31 -400 31 -400 0 cellNo=504
rlabel pdiffusion 38 -400 38 -400 0 cellNo=241
rlabel pdiffusion 45 -400 45 -400 0 feedthrough
rlabel pdiffusion 52 -400 52 -400 0 feedthrough
rlabel pdiffusion 59 -400 59 -400 0 feedthrough
rlabel pdiffusion 66 -400 66 -400 0 feedthrough
rlabel pdiffusion 73 -400 73 -400 0 feedthrough
rlabel pdiffusion 80 -400 80 -400 0 feedthrough
rlabel pdiffusion 87 -400 87 -400 0 feedthrough
rlabel pdiffusion 94 -400 94 -400 0 feedthrough
rlabel pdiffusion 101 -400 101 -400 0 feedthrough
rlabel pdiffusion 108 -400 108 -400 0 feedthrough
rlabel pdiffusion 115 -400 115 -400 0 cellNo=106
rlabel pdiffusion 122 -400 122 -400 0 feedthrough
rlabel pdiffusion 129 -400 129 -400 0 feedthrough
rlabel pdiffusion 136 -400 136 -400 0 cellNo=163
rlabel pdiffusion 143 -400 143 -400 0 cellNo=658
rlabel pdiffusion 150 -400 150 -400 0 feedthrough
rlabel pdiffusion 157 -400 157 -400 0 feedthrough
rlabel pdiffusion 164 -400 164 -400 0 feedthrough
rlabel pdiffusion 171 -400 171 -400 0 cellNo=7
rlabel pdiffusion 178 -400 178 -400 0 cellNo=788
rlabel pdiffusion 185 -400 185 -400 0 feedthrough
rlabel pdiffusion 192 -400 192 -400 0 feedthrough
rlabel pdiffusion 199 -400 199 -400 0 feedthrough
rlabel pdiffusion 206 -400 206 -400 0 cellNo=794
rlabel pdiffusion 213 -400 213 -400 0 feedthrough
rlabel pdiffusion 220 -400 220 -400 0 feedthrough
rlabel pdiffusion 227 -400 227 -400 0 feedthrough
rlabel pdiffusion 234 -400 234 -400 0 feedthrough
rlabel pdiffusion 241 -400 241 -400 0 feedthrough
rlabel pdiffusion 248 -400 248 -400 0 feedthrough
rlabel pdiffusion 255 -400 255 -400 0 feedthrough
rlabel pdiffusion 262 -400 262 -400 0 feedthrough
rlabel pdiffusion 269 -400 269 -400 0 feedthrough
rlabel pdiffusion 276 -400 276 -400 0 cellNo=601
rlabel pdiffusion 283 -400 283 -400 0 feedthrough
rlabel pdiffusion 290 -400 290 -400 0 feedthrough
rlabel pdiffusion 297 -400 297 -400 0 feedthrough
rlabel pdiffusion 304 -400 304 -400 0 feedthrough
rlabel pdiffusion 311 -400 311 -400 0 feedthrough
rlabel pdiffusion 318 -400 318 -400 0 cellNo=813
rlabel pdiffusion 325 -400 325 -400 0 feedthrough
rlabel pdiffusion 332 -400 332 -400 0 feedthrough
rlabel pdiffusion 339 -400 339 -400 0 cellNo=8
rlabel pdiffusion 346 -400 346 -400 0 feedthrough
rlabel pdiffusion 353 -400 353 -400 0 feedthrough
rlabel pdiffusion 360 -400 360 -400 0 cellNo=208
rlabel pdiffusion 367 -400 367 -400 0 feedthrough
rlabel pdiffusion 374 -400 374 -400 0 feedthrough
rlabel pdiffusion 381 -400 381 -400 0 feedthrough
rlabel pdiffusion 388 -400 388 -400 0 feedthrough
rlabel pdiffusion 395 -400 395 -400 0 feedthrough
rlabel pdiffusion 402 -400 402 -400 0 cellNo=317
rlabel pdiffusion 409 -400 409 -400 0 feedthrough
rlabel pdiffusion 416 -400 416 -400 0 feedthrough
rlabel pdiffusion 423 -400 423 -400 0 cellNo=560
rlabel pdiffusion 430 -400 430 -400 0 feedthrough
rlabel pdiffusion 437 -400 437 -400 0 feedthrough
rlabel pdiffusion 444 -400 444 -400 0 feedthrough
rlabel pdiffusion 451 -400 451 -400 0 cellNo=13
rlabel pdiffusion 458 -400 458 -400 0 feedthrough
rlabel pdiffusion 465 -400 465 -400 0 feedthrough
rlabel pdiffusion 472 -400 472 -400 0 cellNo=766
rlabel pdiffusion 479 -400 479 -400 0 feedthrough
rlabel pdiffusion 486 -400 486 -400 0 feedthrough
rlabel pdiffusion 493 -400 493 -400 0 cellNo=23
rlabel pdiffusion 500 -400 500 -400 0 feedthrough
rlabel pdiffusion 507 -400 507 -400 0 cellNo=551
rlabel pdiffusion 514 -400 514 -400 0 feedthrough
rlabel pdiffusion 521 -400 521 -400 0 cellNo=552
rlabel pdiffusion 528 -400 528 -400 0 feedthrough
rlabel pdiffusion 535 -400 535 -400 0 feedthrough
rlabel pdiffusion 542 -400 542 -400 0 feedthrough
rlabel pdiffusion 549 -400 549 -400 0 cellNo=698
rlabel pdiffusion 556 -400 556 -400 0 feedthrough
rlabel pdiffusion 563 -400 563 -400 0 cellNo=214
rlabel pdiffusion 570 -400 570 -400 0 feedthrough
rlabel pdiffusion 577 -400 577 -400 0 cellNo=421
rlabel pdiffusion 584 -400 584 -400 0 feedthrough
rlabel pdiffusion 591 -400 591 -400 0 feedthrough
rlabel pdiffusion 598 -400 598 -400 0 feedthrough
rlabel pdiffusion 605 -400 605 -400 0 feedthrough
rlabel pdiffusion 612 -400 612 -400 0 feedthrough
rlabel pdiffusion 619 -400 619 -400 0 feedthrough
rlabel pdiffusion 626 -400 626 -400 0 feedthrough
rlabel pdiffusion 633 -400 633 -400 0 feedthrough
rlabel pdiffusion 640 -400 640 -400 0 feedthrough
rlabel pdiffusion 647 -400 647 -400 0 feedthrough
rlabel pdiffusion 654 -400 654 -400 0 feedthrough
rlabel pdiffusion 661 -400 661 -400 0 feedthrough
rlabel pdiffusion 668 -400 668 -400 0 feedthrough
rlabel pdiffusion 675 -400 675 -400 0 feedthrough
rlabel pdiffusion 682 -400 682 -400 0 cellNo=175
rlabel pdiffusion 689 -400 689 -400 0 feedthrough
rlabel pdiffusion 696 -400 696 -400 0 feedthrough
rlabel pdiffusion 703 -400 703 -400 0 feedthrough
rlabel pdiffusion 710 -400 710 -400 0 feedthrough
rlabel pdiffusion 717 -400 717 -400 0 feedthrough
rlabel pdiffusion 724 -400 724 -400 0 feedthrough
rlabel pdiffusion 731 -400 731 -400 0 feedthrough
rlabel pdiffusion 738 -400 738 -400 0 feedthrough
rlabel pdiffusion 745 -400 745 -400 0 feedthrough
rlabel pdiffusion 752 -400 752 -400 0 feedthrough
rlabel pdiffusion 759 -400 759 -400 0 feedthrough
rlabel pdiffusion 766 -400 766 -400 0 feedthrough
rlabel pdiffusion 773 -400 773 -400 0 feedthrough
rlabel pdiffusion 780 -400 780 -400 0 feedthrough
rlabel pdiffusion 787 -400 787 -400 0 feedthrough
rlabel pdiffusion 794 -400 794 -400 0 feedthrough
rlabel pdiffusion 801 -400 801 -400 0 feedthrough
rlabel pdiffusion 808 -400 808 -400 0 feedthrough
rlabel pdiffusion 815 -400 815 -400 0 feedthrough
rlabel pdiffusion 822 -400 822 -400 0 feedthrough
rlabel pdiffusion 829 -400 829 -400 0 feedthrough
rlabel pdiffusion 836 -400 836 -400 0 feedthrough
rlabel pdiffusion 843 -400 843 -400 0 feedthrough
rlabel pdiffusion 850 -400 850 -400 0 feedthrough
rlabel pdiffusion 857 -400 857 -400 0 feedthrough
rlabel pdiffusion 864 -400 864 -400 0 feedthrough
rlabel pdiffusion 871 -400 871 -400 0 feedthrough
rlabel pdiffusion 878 -400 878 -400 0 feedthrough
rlabel pdiffusion 885 -400 885 -400 0 feedthrough
rlabel pdiffusion 892 -400 892 -400 0 feedthrough
rlabel pdiffusion 899 -400 899 -400 0 cellNo=69
rlabel pdiffusion 906 -400 906 -400 0 feedthrough
rlabel pdiffusion 913 -400 913 -400 0 feedthrough
rlabel pdiffusion 920 -400 920 -400 0 feedthrough
rlabel pdiffusion 927 -400 927 -400 0 feedthrough
rlabel pdiffusion 934 -400 934 -400 0 feedthrough
rlabel pdiffusion 941 -400 941 -400 0 feedthrough
rlabel pdiffusion 948 -400 948 -400 0 feedthrough
rlabel pdiffusion 955 -400 955 -400 0 feedthrough
rlabel pdiffusion 962 -400 962 -400 0 cellNo=572
rlabel pdiffusion 969 -400 969 -400 0 feedthrough
rlabel pdiffusion 976 -400 976 -400 0 feedthrough
rlabel pdiffusion 983 -400 983 -400 0 feedthrough
rlabel pdiffusion 990 -400 990 -400 0 feedthrough
rlabel pdiffusion 997 -400 997 -400 0 cellNo=428
rlabel pdiffusion 1004 -400 1004 -400 0 feedthrough
rlabel pdiffusion 1011 -400 1011 -400 0 feedthrough
rlabel pdiffusion 1018 -400 1018 -400 0 feedthrough
rlabel pdiffusion 1025 -400 1025 -400 0 feedthrough
rlabel pdiffusion 1032 -400 1032 -400 0 cellNo=244
rlabel pdiffusion 1039 -400 1039 -400 0 cellNo=608
rlabel pdiffusion 1046 -400 1046 -400 0 cellNo=702
rlabel pdiffusion 1053 -400 1053 -400 0 feedthrough
rlabel pdiffusion 1067 -400 1067 -400 0 feedthrough
rlabel pdiffusion 1109 -400 1109 -400 0 feedthrough
rlabel pdiffusion 3 -469 3 -469 0 cellNo=416
rlabel pdiffusion 10 -469 10 -469 0 cellNo=271
rlabel pdiffusion 17 -469 17 -469 0 feedthrough
rlabel pdiffusion 24 -469 24 -469 0 feedthrough
rlabel pdiffusion 31 -469 31 -469 0 feedthrough
rlabel pdiffusion 38 -469 38 -469 0 feedthrough
rlabel pdiffusion 45 -469 45 -469 0 feedthrough
rlabel pdiffusion 52 -469 52 -469 0 feedthrough
rlabel pdiffusion 59 -469 59 -469 0 feedthrough
rlabel pdiffusion 66 -469 66 -469 0 feedthrough
rlabel pdiffusion 73 -469 73 -469 0 feedthrough
rlabel pdiffusion 80 -469 80 -469 0 feedthrough
rlabel pdiffusion 87 -469 87 -469 0 cellNo=412
rlabel pdiffusion 94 -469 94 -469 0 feedthrough
rlabel pdiffusion 101 -469 101 -469 0 feedthrough
rlabel pdiffusion 108 -469 108 -469 0 cellNo=168
rlabel pdiffusion 115 -469 115 -469 0 feedthrough
rlabel pdiffusion 122 -469 122 -469 0 feedthrough
rlabel pdiffusion 129 -469 129 -469 0 feedthrough
rlabel pdiffusion 136 -469 136 -469 0 cellNo=426
rlabel pdiffusion 143 -469 143 -469 0 feedthrough
rlabel pdiffusion 150 -469 150 -469 0 feedthrough
rlabel pdiffusion 157 -469 157 -469 0 feedthrough
rlabel pdiffusion 164 -469 164 -469 0 feedthrough
rlabel pdiffusion 171 -469 171 -469 0 feedthrough
rlabel pdiffusion 178 -469 178 -469 0 feedthrough
rlabel pdiffusion 185 -469 185 -469 0 feedthrough
rlabel pdiffusion 192 -469 192 -469 0 feedthrough
rlabel pdiffusion 199 -469 199 -469 0 feedthrough
rlabel pdiffusion 206 -469 206 -469 0 feedthrough
rlabel pdiffusion 213 -469 213 -469 0 cellNo=169
rlabel pdiffusion 220 -469 220 -469 0 feedthrough
rlabel pdiffusion 227 -469 227 -469 0 cellNo=350
rlabel pdiffusion 234 -469 234 -469 0 feedthrough
rlabel pdiffusion 241 -469 241 -469 0 feedthrough
rlabel pdiffusion 248 -469 248 -469 0 feedthrough
rlabel pdiffusion 255 -469 255 -469 0 feedthrough
rlabel pdiffusion 262 -469 262 -469 0 feedthrough
rlabel pdiffusion 269 -469 269 -469 0 feedthrough
rlabel pdiffusion 276 -469 276 -469 0 cellNo=291
rlabel pdiffusion 283 -469 283 -469 0 feedthrough
rlabel pdiffusion 290 -469 290 -469 0 feedthrough
rlabel pdiffusion 297 -469 297 -469 0 feedthrough
rlabel pdiffusion 304 -469 304 -469 0 cellNo=529
rlabel pdiffusion 311 -469 311 -469 0 feedthrough
rlabel pdiffusion 318 -469 318 -469 0 feedthrough
rlabel pdiffusion 325 -469 325 -469 0 feedthrough
rlabel pdiffusion 332 -469 332 -469 0 feedthrough
rlabel pdiffusion 339 -469 339 -469 0 feedthrough
rlabel pdiffusion 346 -469 346 -469 0 cellNo=178
rlabel pdiffusion 353 -469 353 -469 0 feedthrough
rlabel pdiffusion 360 -469 360 -469 0 feedthrough
rlabel pdiffusion 367 -469 367 -469 0 feedthrough
rlabel pdiffusion 374 -469 374 -469 0 feedthrough
rlabel pdiffusion 381 -469 381 -469 0 feedthrough
rlabel pdiffusion 388 -469 388 -469 0 cellNo=688
rlabel pdiffusion 395 -469 395 -469 0 feedthrough
rlabel pdiffusion 402 -469 402 -469 0 cellNo=645
rlabel pdiffusion 409 -469 409 -469 0 cellNo=355
rlabel pdiffusion 416 -469 416 -469 0 feedthrough
rlabel pdiffusion 423 -469 423 -469 0 feedthrough
rlabel pdiffusion 430 -469 430 -469 0 feedthrough
rlabel pdiffusion 437 -469 437 -469 0 feedthrough
rlabel pdiffusion 444 -469 444 -469 0 feedthrough
rlabel pdiffusion 451 -469 451 -469 0 feedthrough
rlabel pdiffusion 458 -469 458 -469 0 cellNo=755
rlabel pdiffusion 465 -469 465 -469 0 feedthrough
rlabel pdiffusion 472 -469 472 -469 0 cellNo=604
rlabel pdiffusion 479 -469 479 -469 0 feedthrough
rlabel pdiffusion 486 -469 486 -469 0 feedthrough
rlabel pdiffusion 493 -469 493 -469 0 feedthrough
rlabel pdiffusion 500 -469 500 -469 0 cellNo=708
rlabel pdiffusion 507 -469 507 -469 0 cellNo=639
rlabel pdiffusion 514 -469 514 -469 0 feedthrough
rlabel pdiffusion 521 -469 521 -469 0 cellNo=587
rlabel pdiffusion 528 -469 528 -469 0 cellNo=603
rlabel pdiffusion 535 -469 535 -469 0 feedthrough
rlabel pdiffusion 542 -469 542 -469 0 feedthrough
rlabel pdiffusion 549 -469 549 -469 0 feedthrough
rlabel pdiffusion 556 -469 556 -469 0 feedthrough
rlabel pdiffusion 563 -469 563 -469 0 cellNo=309
rlabel pdiffusion 570 -469 570 -469 0 feedthrough
rlabel pdiffusion 577 -469 577 -469 0 feedthrough
rlabel pdiffusion 584 -469 584 -469 0 cellNo=388
rlabel pdiffusion 591 -469 591 -469 0 feedthrough
rlabel pdiffusion 598 -469 598 -469 0 cellNo=307
rlabel pdiffusion 605 -469 605 -469 0 feedthrough
rlabel pdiffusion 612 -469 612 -469 0 feedthrough
rlabel pdiffusion 619 -469 619 -469 0 feedthrough
rlabel pdiffusion 626 -469 626 -469 0 feedthrough
rlabel pdiffusion 633 -469 633 -469 0 cellNo=207
rlabel pdiffusion 640 -469 640 -469 0 feedthrough
rlabel pdiffusion 647 -469 647 -469 0 feedthrough
rlabel pdiffusion 654 -469 654 -469 0 feedthrough
rlabel pdiffusion 661 -469 661 -469 0 cellNo=122
rlabel pdiffusion 668 -469 668 -469 0 feedthrough
rlabel pdiffusion 675 -469 675 -469 0 feedthrough
rlabel pdiffusion 682 -469 682 -469 0 feedthrough
rlabel pdiffusion 689 -469 689 -469 0 feedthrough
rlabel pdiffusion 696 -469 696 -469 0 feedthrough
rlabel pdiffusion 703 -469 703 -469 0 feedthrough
rlabel pdiffusion 710 -469 710 -469 0 feedthrough
rlabel pdiffusion 717 -469 717 -469 0 feedthrough
rlabel pdiffusion 724 -469 724 -469 0 cellNo=449
rlabel pdiffusion 731 -469 731 -469 0 feedthrough
rlabel pdiffusion 738 -469 738 -469 0 cellNo=887
rlabel pdiffusion 745 -469 745 -469 0 feedthrough
rlabel pdiffusion 752 -469 752 -469 0 cellNo=472
rlabel pdiffusion 759 -469 759 -469 0 feedthrough
rlabel pdiffusion 766 -469 766 -469 0 feedthrough
rlabel pdiffusion 773 -469 773 -469 0 feedthrough
rlabel pdiffusion 780 -469 780 -469 0 feedthrough
rlabel pdiffusion 787 -469 787 -469 0 feedthrough
rlabel pdiffusion 794 -469 794 -469 0 feedthrough
rlabel pdiffusion 801 -469 801 -469 0 feedthrough
rlabel pdiffusion 808 -469 808 -469 0 feedthrough
rlabel pdiffusion 815 -469 815 -469 0 feedthrough
rlabel pdiffusion 822 -469 822 -469 0 feedthrough
rlabel pdiffusion 829 -469 829 -469 0 feedthrough
rlabel pdiffusion 836 -469 836 -469 0 feedthrough
rlabel pdiffusion 843 -469 843 -469 0 feedthrough
rlabel pdiffusion 850 -469 850 -469 0 feedthrough
rlabel pdiffusion 857 -469 857 -469 0 feedthrough
rlabel pdiffusion 864 -469 864 -469 0 feedthrough
rlabel pdiffusion 871 -469 871 -469 0 feedthrough
rlabel pdiffusion 878 -469 878 -469 0 feedthrough
rlabel pdiffusion 885 -469 885 -469 0 feedthrough
rlabel pdiffusion 892 -469 892 -469 0 feedthrough
rlabel pdiffusion 899 -469 899 -469 0 feedthrough
rlabel pdiffusion 906 -469 906 -469 0 feedthrough
rlabel pdiffusion 913 -469 913 -469 0 feedthrough
rlabel pdiffusion 920 -469 920 -469 0 feedthrough
rlabel pdiffusion 927 -469 927 -469 0 feedthrough
rlabel pdiffusion 934 -469 934 -469 0 feedthrough
rlabel pdiffusion 941 -469 941 -469 0 feedthrough
rlabel pdiffusion 948 -469 948 -469 0 feedthrough
rlabel pdiffusion 955 -469 955 -469 0 feedthrough
rlabel pdiffusion 962 -469 962 -469 0 feedthrough
rlabel pdiffusion 969 -469 969 -469 0 feedthrough
rlabel pdiffusion 976 -469 976 -469 0 feedthrough
rlabel pdiffusion 983 -469 983 -469 0 cellNo=798
rlabel pdiffusion 990 -469 990 -469 0 feedthrough
rlabel pdiffusion 997 -469 997 -469 0 feedthrough
rlabel pdiffusion 1004 -469 1004 -469 0 feedthrough
rlabel pdiffusion 1011 -469 1011 -469 0 feedthrough
rlabel pdiffusion 1018 -469 1018 -469 0 feedthrough
rlabel pdiffusion 1025 -469 1025 -469 0 feedthrough
rlabel pdiffusion 1032 -469 1032 -469 0 feedthrough
rlabel pdiffusion 1039 -469 1039 -469 0 feedthrough
rlabel pdiffusion 1046 -469 1046 -469 0 feedthrough
rlabel pdiffusion 1053 -469 1053 -469 0 feedthrough
rlabel pdiffusion 1060 -469 1060 -469 0 feedthrough
rlabel pdiffusion 1067 -469 1067 -469 0 feedthrough
rlabel pdiffusion 1074 -469 1074 -469 0 feedthrough
rlabel pdiffusion 1081 -469 1081 -469 0 feedthrough
rlabel pdiffusion 1088 -469 1088 -469 0 feedthrough
rlabel pdiffusion 1095 -469 1095 -469 0 feedthrough
rlabel pdiffusion 1102 -469 1102 -469 0 feedthrough
rlabel pdiffusion 1109 -469 1109 -469 0 feedthrough
rlabel pdiffusion 1116 -469 1116 -469 0 feedthrough
rlabel pdiffusion 1123 -469 1123 -469 0 feedthrough
rlabel pdiffusion 1130 -469 1130 -469 0 feedthrough
rlabel pdiffusion 1137 -469 1137 -469 0 cellNo=189
rlabel pdiffusion 1144 -469 1144 -469 0 cellNo=300
rlabel pdiffusion 1151 -469 1151 -469 0 feedthrough
rlabel pdiffusion 3 -564 3 -564 0 cellNo=403
rlabel pdiffusion 10 -564 10 -564 0 feedthrough
rlabel pdiffusion 17 -564 17 -564 0 feedthrough
rlabel pdiffusion 24 -564 24 -564 0 feedthrough
rlabel pdiffusion 31 -564 31 -564 0 cellNo=874
rlabel pdiffusion 38 -564 38 -564 0 feedthrough
rlabel pdiffusion 45 -564 45 -564 0 feedthrough
rlabel pdiffusion 52 -564 52 -564 0 feedthrough
rlabel pdiffusion 59 -564 59 -564 0 feedthrough
rlabel pdiffusion 66 -564 66 -564 0 feedthrough
rlabel pdiffusion 73 -564 73 -564 0 cellNo=78
rlabel pdiffusion 80 -564 80 -564 0 cellNo=649
rlabel pdiffusion 87 -564 87 -564 0 feedthrough
rlabel pdiffusion 94 -564 94 -564 0 feedthrough
rlabel pdiffusion 101 -564 101 -564 0 feedthrough
rlabel pdiffusion 108 -564 108 -564 0 cellNo=828
rlabel pdiffusion 115 -564 115 -564 0 feedthrough
rlabel pdiffusion 122 -564 122 -564 0 feedthrough
rlabel pdiffusion 129 -564 129 -564 0 feedthrough
rlabel pdiffusion 136 -564 136 -564 0 feedthrough
rlabel pdiffusion 143 -564 143 -564 0 feedthrough
rlabel pdiffusion 150 -564 150 -564 0 cellNo=353
rlabel pdiffusion 157 -564 157 -564 0 feedthrough
rlabel pdiffusion 164 -564 164 -564 0 cellNo=270
rlabel pdiffusion 171 -564 171 -564 0 feedthrough
rlabel pdiffusion 178 -564 178 -564 0 feedthrough
rlabel pdiffusion 185 -564 185 -564 0 feedthrough
rlabel pdiffusion 192 -564 192 -564 0 cellNo=881
rlabel pdiffusion 199 -564 199 -564 0 cellNo=661
rlabel pdiffusion 206 -564 206 -564 0 feedthrough
rlabel pdiffusion 213 -564 213 -564 0 cellNo=159
rlabel pdiffusion 220 -564 220 -564 0 feedthrough
rlabel pdiffusion 227 -564 227 -564 0 feedthrough
rlabel pdiffusion 234 -564 234 -564 0 feedthrough
rlabel pdiffusion 241 -564 241 -564 0 feedthrough
rlabel pdiffusion 248 -564 248 -564 0 feedthrough
rlabel pdiffusion 255 -564 255 -564 0 feedthrough
rlabel pdiffusion 262 -564 262 -564 0 feedthrough
rlabel pdiffusion 269 -564 269 -564 0 feedthrough
rlabel pdiffusion 276 -564 276 -564 0 feedthrough
rlabel pdiffusion 283 -564 283 -564 0 feedthrough
rlabel pdiffusion 290 -564 290 -564 0 feedthrough
rlabel pdiffusion 297 -564 297 -564 0 feedthrough
rlabel pdiffusion 304 -564 304 -564 0 feedthrough
rlabel pdiffusion 311 -564 311 -564 0 feedthrough
rlabel pdiffusion 318 -564 318 -564 0 cellNo=783
rlabel pdiffusion 325 -564 325 -564 0 feedthrough
rlabel pdiffusion 332 -564 332 -564 0 feedthrough
rlabel pdiffusion 339 -564 339 -564 0 feedthrough
rlabel pdiffusion 346 -564 346 -564 0 feedthrough
rlabel pdiffusion 353 -564 353 -564 0 cellNo=119
rlabel pdiffusion 360 -564 360 -564 0 feedthrough
rlabel pdiffusion 367 -564 367 -564 0 cellNo=796
rlabel pdiffusion 374 -564 374 -564 0 feedthrough
rlabel pdiffusion 381 -564 381 -564 0 feedthrough
rlabel pdiffusion 388 -564 388 -564 0 cellNo=636
rlabel pdiffusion 395 -564 395 -564 0 cellNo=287
rlabel pdiffusion 402 -564 402 -564 0 feedthrough
rlabel pdiffusion 409 -564 409 -564 0 cellNo=193
rlabel pdiffusion 416 -564 416 -564 0 feedthrough
rlabel pdiffusion 423 -564 423 -564 0 cellNo=678
rlabel pdiffusion 430 -564 430 -564 0 feedthrough
rlabel pdiffusion 437 -564 437 -564 0 feedthrough
rlabel pdiffusion 444 -564 444 -564 0 feedthrough
rlabel pdiffusion 451 -564 451 -564 0 feedthrough
rlabel pdiffusion 458 -564 458 -564 0 feedthrough
rlabel pdiffusion 465 -564 465 -564 0 feedthrough
rlabel pdiffusion 472 -564 472 -564 0 feedthrough
rlabel pdiffusion 479 -564 479 -564 0 feedthrough
rlabel pdiffusion 486 -564 486 -564 0 feedthrough
rlabel pdiffusion 493 -564 493 -564 0 feedthrough
rlabel pdiffusion 500 -564 500 -564 0 feedthrough
rlabel pdiffusion 507 -564 507 -564 0 cellNo=383
rlabel pdiffusion 514 -564 514 -564 0 feedthrough
rlabel pdiffusion 521 -564 521 -564 0 feedthrough
rlabel pdiffusion 528 -564 528 -564 0 feedthrough
rlabel pdiffusion 535 -564 535 -564 0 cellNo=400
rlabel pdiffusion 542 -564 542 -564 0 feedthrough
rlabel pdiffusion 549 -564 549 -564 0 cellNo=754
rlabel pdiffusion 556 -564 556 -564 0 feedthrough
rlabel pdiffusion 563 -564 563 -564 0 cellNo=107
rlabel pdiffusion 570 -564 570 -564 0 cellNo=188
rlabel pdiffusion 577 -564 577 -564 0 feedthrough
rlabel pdiffusion 584 -564 584 -564 0 feedthrough
rlabel pdiffusion 591 -564 591 -564 0 cellNo=120
rlabel pdiffusion 598 -564 598 -564 0 cellNo=348
rlabel pdiffusion 605 -564 605 -564 0 cellNo=199
rlabel pdiffusion 612 -564 612 -564 0 feedthrough
rlabel pdiffusion 619 -564 619 -564 0 feedthrough
rlabel pdiffusion 626 -564 626 -564 0 cellNo=436
rlabel pdiffusion 633 -564 633 -564 0 feedthrough
rlabel pdiffusion 640 -564 640 -564 0 feedthrough
rlabel pdiffusion 647 -564 647 -564 0 feedthrough
rlabel pdiffusion 654 -564 654 -564 0 feedthrough
rlabel pdiffusion 661 -564 661 -564 0 cellNo=70
rlabel pdiffusion 668 -564 668 -564 0 feedthrough
rlabel pdiffusion 675 -564 675 -564 0 feedthrough
rlabel pdiffusion 682 -564 682 -564 0 feedthrough
rlabel pdiffusion 689 -564 689 -564 0 feedthrough
rlabel pdiffusion 696 -564 696 -564 0 feedthrough
rlabel pdiffusion 703 -564 703 -564 0 feedthrough
rlabel pdiffusion 710 -564 710 -564 0 cellNo=160
rlabel pdiffusion 717 -564 717 -564 0 feedthrough
rlabel pdiffusion 724 -564 724 -564 0 feedthrough
rlabel pdiffusion 731 -564 731 -564 0 cellNo=93
rlabel pdiffusion 738 -564 738 -564 0 feedthrough
rlabel pdiffusion 745 -564 745 -564 0 feedthrough
rlabel pdiffusion 752 -564 752 -564 0 feedthrough
rlabel pdiffusion 759 -564 759 -564 0 feedthrough
rlabel pdiffusion 766 -564 766 -564 0 feedthrough
rlabel pdiffusion 773 -564 773 -564 0 feedthrough
rlabel pdiffusion 780 -564 780 -564 0 feedthrough
rlabel pdiffusion 787 -564 787 -564 0 feedthrough
rlabel pdiffusion 794 -564 794 -564 0 feedthrough
rlabel pdiffusion 801 -564 801 -564 0 feedthrough
rlabel pdiffusion 808 -564 808 -564 0 feedthrough
rlabel pdiffusion 815 -564 815 -564 0 feedthrough
rlabel pdiffusion 822 -564 822 -564 0 feedthrough
rlabel pdiffusion 829 -564 829 -564 0 feedthrough
rlabel pdiffusion 836 -564 836 -564 0 feedthrough
rlabel pdiffusion 843 -564 843 -564 0 feedthrough
rlabel pdiffusion 850 -564 850 -564 0 feedthrough
rlabel pdiffusion 857 -564 857 -564 0 feedthrough
rlabel pdiffusion 864 -564 864 -564 0 feedthrough
rlabel pdiffusion 871 -564 871 -564 0 feedthrough
rlabel pdiffusion 878 -564 878 -564 0 feedthrough
rlabel pdiffusion 885 -564 885 -564 0 feedthrough
rlabel pdiffusion 892 -564 892 -564 0 feedthrough
rlabel pdiffusion 899 -564 899 -564 0 feedthrough
rlabel pdiffusion 906 -564 906 -564 0 feedthrough
rlabel pdiffusion 913 -564 913 -564 0 feedthrough
rlabel pdiffusion 920 -564 920 -564 0 feedthrough
rlabel pdiffusion 927 -564 927 -564 0 feedthrough
rlabel pdiffusion 934 -564 934 -564 0 feedthrough
rlabel pdiffusion 941 -564 941 -564 0 feedthrough
rlabel pdiffusion 948 -564 948 -564 0 feedthrough
rlabel pdiffusion 955 -564 955 -564 0 feedthrough
rlabel pdiffusion 962 -564 962 -564 0 feedthrough
rlabel pdiffusion 969 -564 969 -564 0 feedthrough
rlabel pdiffusion 976 -564 976 -564 0 feedthrough
rlabel pdiffusion 983 -564 983 -564 0 feedthrough
rlabel pdiffusion 990 -564 990 -564 0 feedthrough
rlabel pdiffusion 997 -564 997 -564 0 feedthrough
rlabel pdiffusion 1004 -564 1004 -564 0 feedthrough
rlabel pdiffusion 1011 -564 1011 -564 0 feedthrough
rlabel pdiffusion 1018 -564 1018 -564 0 feedthrough
rlabel pdiffusion 1025 -564 1025 -564 0 feedthrough
rlabel pdiffusion 1032 -564 1032 -564 0 feedthrough
rlabel pdiffusion 1039 -564 1039 -564 0 feedthrough
rlabel pdiffusion 1046 -564 1046 -564 0 feedthrough
rlabel pdiffusion 1053 -564 1053 -564 0 feedthrough
rlabel pdiffusion 1060 -564 1060 -564 0 feedthrough
rlabel pdiffusion 1067 -564 1067 -564 0 feedthrough
rlabel pdiffusion 1074 -564 1074 -564 0 feedthrough
rlabel pdiffusion 1081 -564 1081 -564 0 feedthrough
rlabel pdiffusion 1088 -564 1088 -564 0 feedthrough
rlabel pdiffusion 1095 -564 1095 -564 0 feedthrough
rlabel pdiffusion 1102 -564 1102 -564 0 feedthrough
rlabel pdiffusion 1116 -564 1116 -564 0 feedthrough
rlabel pdiffusion 1123 -564 1123 -564 0 feedthrough
rlabel pdiffusion 1172 -564 1172 -564 0 cellNo=177
rlabel pdiffusion 1179 -564 1179 -564 0 feedthrough
rlabel pdiffusion 3 -655 3 -655 0 cellNo=430
rlabel pdiffusion 10 -655 10 -655 0 feedthrough
rlabel pdiffusion 17 -655 17 -655 0 feedthrough
rlabel pdiffusion 24 -655 24 -655 0 cellNo=648
rlabel pdiffusion 31 -655 31 -655 0 feedthrough
rlabel pdiffusion 38 -655 38 -655 0 feedthrough
rlabel pdiffusion 45 -655 45 -655 0 feedthrough
rlabel pdiffusion 52 -655 52 -655 0 cellNo=523
rlabel pdiffusion 59 -655 59 -655 0 feedthrough
rlabel pdiffusion 66 -655 66 -655 0 cellNo=729
rlabel pdiffusion 73 -655 73 -655 0 feedthrough
rlabel pdiffusion 80 -655 80 -655 0 cellNo=714
rlabel pdiffusion 87 -655 87 -655 0 cellNo=619
rlabel pdiffusion 94 -655 94 -655 0 feedthrough
rlabel pdiffusion 101 -655 101 -655 0 cellNo=480
rlabel pdiffusion 108 -655 108 -655 0 feedthrough
rlabel pdiffusion 115 -655 115 -655 0 cellNo=303
rlabel pdiffusion 122 -655 122 -655 0 feedthrough
rlabel pdiffusion 129 -655 129 -655 0 cellNo=201
rlabel pdiffusion 136 -655 136 -655 0 feedthrough
rlabel pdiffusion 143 -655 143 -655 0 feedthrough
rlabel pdiffusion 150 -655 150 -655 0 feedthrough
rlabel pdiffusion 157 -655 157 -655 0 cellNo=153
rlabel pdiffusion 164 -655 164 -655 0 feedthrough
rlabel pdiffusion 171 -655 171 -655 0 feedthrough
rlabel pdiffusion 178 -655 178 -655 0 feedthrough
rlabel pdiffusion 185 -655 185 -655 0 cellNo=836
rlabel pdiffusion 192 -655 192 -655 0 feedthrough
rlabel pdiffusion 199 -655 199 -655 0 feedthrough
rlabel pdiffusion 206 -655 206 -655 0 cellNo=749
rlabel pdiffusion 213 -655 213 -655 0 feedthrough
rlabel pdiffusion 220 -655 220 -655 0 feedthrough
rlabel pdiffusion 227 -655 227 -655 0 feedthrough
rlabel pdiffusion 234 -655 234 -655 0 cellNo=629
rlabel pdiffusion 241 -655 241 -655 0 feedthrough
rlabel pdiffusion 248 -655 248 -655 0 feedthrough
rlabel pdiffusion 255 -655 255 -655 0 feedthrough
rlabel pdiffusion 262 -655 262 -655 0 feedthrough
rlabel pdiffusion 269 -655 269 -655 0 feedthrough
rlabel pdiffusion 276 -655 276 -655 0 feedthrough
rlabel pdiffusion 283 -655 283 -655 0 feedthrough
rlabel pdiffusion 290 -655 290 -655 0 feedthrough
rlabel pdiffusion 297 -655 297 -655 0 feedthrough
rlabel pdiffusion 304 -655 304 -655 0 feedthrough
rlabel pdiffusion 311 -655 311 -655 0 feedthrough
rlabel pdiffusion 318 -655 318 -655 0 feedthrough
rlabel pdiffusion 325 -655 325 -655 0 feedthrough
rlabel pdiffusion 332 -655 332 -655 0 cellNo=364
rlabel pdiffusion 339 -655 339 -655 0 cellNo=387
rlabel pdiffusion 346 -655 346 -655 0 cellNo=115
rlabel pdiffusion 353 -655 353 -655 0 feedthrough
rlabel pdiffusion 360 -655 360 -655 0 feedthrough
rlabel pdiffusion 367 -655 367 -655 0 feedthrough
rlabel pdiffusion 374 -655 374 -655 0 feedthrough
rlabel pdiffusion 381 -655 381 -655 0 feedthrough
rlabel pdiffusion 388 -655 388 -655 0 feedthrough
rlabel pdiffusion 395 -655 395 -655 0 feedthrough
rlabel pdiffusion 402 -655 402 -655 0 feedthrough
rlabel pdiffusion 409 -655 409 -655 0 cellNo=732
rlabel pdiffusion 416 -655 416 -655 0 cellNo=326
rlabel pdiffusion 423 -655 423 -655 0 feedthrough
rlabel pdiffusion 430 -655 430 -655 0 feedthrough
rlabel pdiffusion 437 -655 437 -655 0 feedthrough
rlabel pdiffusion 444 -655 444 -655 0 cellNo=344
rlabel pdiffusion 451 -655 451 -655 0 feedthrough
rlabel pdiffusion 458 -655 458 -655 0 feedthrough
rlabel pdiffusion 465 -655 465 -655 0 feedthrough
rlabel pdiffusion 472 -655 472 -655 0 feedthrough
rlabel pdiffusion 479 -655 479 -655 0 cellNo=666
rlabel pdiffusion 486 -655 486 -655 0 feedthrough
rlabel pdiffusion 493 -655 493 -655 0 feedthrough
rlabel pdiffusion 500 -655 500 -655 0 cellNo=777
rlabel pdiffusion 507 -655 507 -655 0 feedthrough
rlabel pdiffusion 514 -655 514 -655 0 cellNo=83
rlabel pdiffusion 521 -655 521 -655 0 cellNo=456
rlabel pdiffusion 528 -655 528 -655 0 feedthrough
rlabel pdiffusion 535 -655 535 -655 0 feedthrough
rlabel pdiffusion 542 -655 542 -655 0 feedthrough
rlabel pdiffusion 549 -655 549 -655 0 cellNo=319
rlabel pdiffusion 556 -655 556 -655 0 feedthrough
rlabel pdiffusion 563 -655 563 -655 0 feedthrough
rlabel pdiffusion 570 -655 570 -655 0 feedthrough
rlabel pdiffusion 577 -655 577 -655 0 feedthrough
rlabel pdiffusion 584 -655 584 -655 0 feedthrough
rlabel pdiffusion 591 -655 591 -655 0 feedthrough
rlabel pdiffusion 598 -655 598 -655 0 feedthrough
rlabel pdiffusion 605 -655 605 -655 0 cellNo=206
rlabel pdiffusion 612 -655 612 -655 0 cellNo=789
rlabel pdiffusion 619 -655 619 -655 0 feedthrough
rlabel pdiffusion 626 -655 626 -655 0 feedthrough
rlabel pdiffusion 633 -655 633 -655 0 feedthrough
rlabel pdiffusion 640 -655 640 -655 0 feedthrough
rlabel pdiffusion 647 -655 647 -655 0 feedthrough
rlabel pdiffusion 654 -655 654 -655 0 cellNo=434
rlabel pdiffusion 661 -655 661 -655 0 feedthrough
rlabel pdiffusion 668 -655 668 -655 0 feedthrough
rlabel pdiffusion 675 -655 675 -655 0 feedthrough
rlabel pdiffusion 682 -655 682 -655 0 feedthrough
rlabel pdiffusion 689 -655 689 -655 0 cellNo=299
rlabel pdiffusion 696 -655 696 -655 0 feedthrough
rlabel pdiffusion 703 -655 703 -655 0 feedthrough
rlabel pdiffusion 710 -655 710 -655 0 feedthrough
rlabel pdiffusion 717 -655 717 -655 0 feedthrough
rlabel pdiffusion 724 -655 724 -655 0 feedthrough
rlabel pdiffusion 731 -655 731 -655 0 feedthrough
rlabel pdiffusion 738 -655 738 -655 0 feedthrough
rlabel pdiffusion 745 -655 745 -655 0 feedthrough
rlabel pdiffusion 752 -655 752 -655 0 feedthrough
rlabel pdiffusion 759 -655 759 -655 0 cellNo=405
rlabel pdiffusion 766 -655 766 -655 0 feedthrough
rlabel pdiffusion 773 -655 773 -655 0 feedthrough
rlabel pdiffusion 780 -655 780 -655 0 feedthrough
rlabel pdiffusion 787 -655 787 -655 0 feedthrough
rlabel pdiffusion 794 -655 794 -655 0 feedthrough
rlabel pdiffusion 801 -655 801 -655 0 feedthrough
rlabel pdiffusion 808 -655 808 -655 0 feedthrough
rlabel pdiffusion 815 -655 815 -655 0 feedthrough
rlabel pdiffusion 822 -655 822 -655 0 feedthrough
rlabel pdiffusion 829 -655 829 -655 0 feedthrough
rlabel pdiffusion 836 -655 836 -655 0 feedthrough
rlabel pdiffusion 843 -655 843 -655 0 feedthrough
rlabel pdiffusion 850 -655 850 -655 0 feedthrough
rlabel pdiffusion 857 -655 857 -655 0 feedthrough
rlabel pdiffusion 864 -655 864 -655 0 feedthrough
rlabel pdiffusion 871 -655 871 -655 0 feedthrough
rlabel pdiffusion 878 -655 878 -655 0 feedthrough
rlabel pdiffusion 885 -655 885 -655 0 feedthrough
rlabel pdiffusion 892 -655 892 -655 0 feedthrough
rlabel pdiffusion 899 -655 899 -655 0 feedthrough
rlabel pdiffusion 906 -655 906 -655 0 feedthrough
rlabel pdiffusion 913 -655 913 -655 0 feedthrough
rlabel pdiffusion 920 -655 920 -655 0 feedthrough
rlabel pdiffusion 927 -655 927 -655 0 feedthrough
rlabel pdiffusion 934 -655 934 -655 0 cellNo=616
rlabel pdiffusion 941 -655 941 -655 0 feedthrough
rlabel pdiffusion 948 -655 948 -655 0 feedthrough
rlabel pdiffusion 955 -655 955 -655 0 feedthrough
rlabel pdiffusion 962 -655 962 -655 0 feedthrough
rlabel pdiffusion 969 -655 969 -655 0 feedthrough
rlabel pdiffusion 976 -655 976 -655 0 feedthrough
rlabel pdiffusion 983 -655 983 -655 0 feedthrough
rlabel pdiffusion 990 -655 990 -655 0 feedthrough
rlabel pdiffusion 997 -655 997 -655 0 feedthrough
rlabel pdiffusion 1004 -655 1004 -655 0 feedthrough
rlabel pdiffusion 1011 -655 1011 -655 0 feedthrough
rlabel pdiffusion 1018 -655 1018 -655 0 feedthrough
rlabel pdiffusion 1025 -655 1025 -655 0 feedthrough
rlabel pdiffusion 1032 -655 1032 -655 0 feedthrough
rlabel pdiffusion 1039 -655 1039 -655 0 feedthrough
rlabel pdiffusion 1046 -655 1046 -655 0 feedthrough
rlabel pdiffusion 1053 -655 1053 -655 0 feedthrough
rlabel pdiffusion 1060 -655 1060 -655 0 feedthrough
rlabel pdiffusion 1067 -655 1067 -655 0 feedthrough
rlabel pdiffusion 1074 -655 1074 -655 0 feedthrough
rlabel pdiffusion 1081 -655 1081 -655 0 feedthrough
rlabel pdiffusion 1088 -655 1088 -655 0 feedthrough
rlabel pdiffusion 1095 -655 1095 -655 0 feedthrough
rlabel pdiffusion 1102 -655 1102 -655 0 feedthrough
rlabel pdiffusion 1109 -655 1109 -655 0 feedthrough
rlabel pdiffusion 1116 -655 1116 -655 0 feedthrough
rlabel pdiffusion 1123 -655 1123 -655 0 feedthrough
rlabel pdiffusion 1130 -655 1130 -655 0 feedthrough
rlabel pdiffusion 1137 -655 1137 -655 0 feedthrough
rlabel pdiffusion 1179 -655 1179 -655 0 feedthrough
rlabel pdiffusion 10 -736 10 -736 0 feedthrough
rlabel pdiffusion 17 -736 17 -736 0 feedthrough
rlabel pdiffusion 24 -736 24 -736 0 feedthrough
rlabel pdiffusion 31 -736 31 -736 0 cellNo=362
rlabel pdiffusion 38 -736 38 -736 0 feedthrough
rlabel pdiffusion 45 -736 45 -736 0 feedthrough
rlabel pdiffusion 52 -736 52 -736 0 feedthrough
rlabel pdiffusion 59 -736 59 -736 0 feedthrough
rlabel pdiffusion 66 -736 66 -736 0 feedthrough
rlabel pdiffusion 73 -736 73 -736 0 cellNo=791
rlabel pdiffusion 80 -736 80 -736 0 feedthrough
rlabel pdiffusion 87 -736 87 -736 0 feedthrough
rlabel pdiffusion 94 -736 94 -736 0 feedthrough
rlabel pdiffusion 101 -736 101 -736 0 feedthrough
rlabel pdiffusion 108 -736 108 -736 0 feedthrough
rlabel pdiffusion 115 -736 115 -736 0 feedthrough
rlabel pdiffusion 122 -736 122 -736 0 cellNo=553
rlabel pdiffusion 129 -736 129 -736 0 feedthrough
rlabel pdiffusion 136 -736 136 -736 0 cellNo=726
rlabel pdiffusion 143 -736 143 -736 0 feedthrough
rlabel pdiffusion 150 -736 150 -736 0 cellNo=622
rlabel pdiffusion 157 -736 157 -736 0 feedthrough
rlabel pdiffusion 164 -736 164 -736 0 feedthrough
rlabel pdiffusion 171 -736 171 -736 0 feedthrough
rlabel pdiffusion 178 -736 178 -736 0 feedthrough
rlabel pdiffusion 185 -736 185 -736 0 cellNo=410
rlabel pdiffusion 192 -736 192 -736 0 cellNo=488
rlabel pdiffusion 199 -736 199 -736 0 feedthrough
rlabel pdiffusion 206 -736 206 -736 0 cellNo=14
rlabel pdiffusion 213 -736 213 -736 0 feedthrough
rlabel pdiffusion 220 -736 220 -736 0 feedthrough
rlabel pdiffusion 227 -736 227 -736 0 feedthrough
rlabel pdiffusion 234 -736 234 -736 0 feedthrough
rlabel pdiffusion 241 -736 241 -736 0 feedthrough
rlabel pdiffusion 248 -736 248 -736 0 feedthrough
rlabel pdiffusion 255 -736 255 -736 0 feedthrough
rlabel pdiffusion 262 -736 262 -736 0 feedthrough
rlabel pdiffusion 269 -736 269 -736 0 feedthrough
rlabel pdiffusion 276 -736 276 -736 0 feedthrough
rlabel pdiffusion 283 -736 283 -736 0 feedthrough
rlabel pdiffusion 290 -736 290 -736 0 feedthrough
rlabel pdiffusion 297 -736 297 -736 0 feedthrough
rlabel pdiffusion 304 -736 304 -736 0 feedthrough
rlabel pdiffusion 311 -736 311 -736 0 cellNo=390
rlabel pdiffusion 318 -736 318 -736 0 feedthrough
rlabel pdiffusion 325 -736 325 -736 0 feedthrough
rlabel pdiffusion 332 -736 332 -736 0 feedthrough
rlabel pdiffusion 339 -736 339 -736 0 cellNo=264
rlabel pdiffusion 346 -736 346 -736 0 feedthrough
rlabel pdiffusion 353 -736 353 -736 0 feedthrough
rlabel pdiffusion 360 -736 360 -736 0 cellNo=2
rlabel pdiffusion 367 -736 367 -736 0 feedthrough
rlabel pdiffusion 374 -736 374 -736 0 feedthrough
rlabel pdiffusion 381 -736 381 -736 0 feedthrough
rlabel pdiffusion 388 -736 388 -736 0 feedthrough
rlabel pdiffusion 395 -736 395 -736 0 cellNo=101
rlabel pdiffusion 402 -736 402 -736 0 cellNo=209
rlabel pdiffusion 409 -736 409 -736 0 cellNo=6
rlabel pdiffusion 416 -736 416 -736 0 feedthrough
rlabel pdiffusion 423 -736 423 -736 0 cellNo=38
rlabel pdiffusion 430 -736 430 -736 0 feedthrough
rlabel pdiffusion 437 -736 437 -736 0 cellNo=382
rlabel pdiffusion 444 -736 444 -736 0 feedthrough
rlabel pdiffusion 451 -736 451 -736 0 feedthrough
rlabel pdiffusion 458 -736 458 -736 0 feedthrough
rlabel pdiffusion 465 -736 465 -736 0 cellNo=435
rlabel pdiffusion 472 -736 472 -736 0 cellNo=806
rlabel pdiffusion 479 -736 479 -736 0 feedthrough
rlabel pdiffusion 486 -736 486 -736 0 feedthrough
rlabel pdiffusion 493 -736 493 -736 0 feedthrough
rlabel pdiffusion 500 -736 500 -736 0 feedthrough
rlabel pdiffusion 507 -736 507 -736 0 feedthrough
rlabel pdiffusion 514 -736 514 -736 0 feedthrough
rlabel pdiffusion 521 -736 521 -736 0 cellNo=289
rlabel pdiffusion 528 -736 528 -736 0 feedthrough
rlabel pdiffusion 535 -736 535 -736 0 feedthrough
rlabel pdiffusion 542 -736 542 -736 0 feedthrough
rlabel pdiffusion 549 -736 549 -736 0 cellNo=310
rlabel pdiffusion 556 -736 556 -736 0 feedthrough
rlabel pdiffusion 563 -736 563 -736 0 feedthrough
rlabel pdiffusion 570 -736 570 -736 0 feedthrough
rlabel pdiffusion 577 -736 577 -736 0 feedthrough
rlabel pdiffusion 584 -736 584 -736 0 feedthrough
rlabel pdiffusion 591 -736 591 -736 0 feedthrough
rlabel pdiffusion 598 -736 598 -736 0 cellNo=15
rlabel pdiffusion 605 -736 605 -736 0 cellNo=854
rlabel pdiffusion 612 -736 612 -736 0 feedthrough
rlabel pdiffusion 619 -736 619 -736 0 feedthrough
rlabel pdiffusion 626 -736 626 -736 0 feedthrough
rlabel pdiffusion 633 -736 633 -736 0 cellNo=314
rlabel pdiffusion 640 -736 640 -736 0 cellNo=145
rlabel pdiffusion 647 -736 647 -736 0 feedthrough
rlabel pdiffusion 654 -736 654 -736 0 feedthrough
rlabel pdiffusion 661 -736 661 -736 0 feedthrough
rlabel pdiffusion 668 -736 668 -736 0 feedthrough
rlabel pdiffusion 675 -736 675 -736 0 feedthrough
rlabel pdiffusion 682 -736 682 -736 0 feedthrough
rlabel pdiffusion 689 -736 689 -736 0 cellNo=234
rlabel pdiffusion 696 -736 696 -736 0 feedthrough
rlabel pdiffusion 703 -736 703 -736 0 feedthrough
rlabel pdiffusion 710 -736 710 -736 0 feedthrough
rlabel pdiffusion 717 -736 717 -736 0 cellNo=363
rlabel pdiffusion 724 -736 724 -736 0 feedthrough
rlabel pdiffusion 731 -736 731 -736 0 feedthrough
rlabel pdiffusion 738 -736 738 -736 0 feedthrough
rlabel pdiffusion 745 -736 745 -736 0 cellNo=484
rlabel pdiffusion 752 -736 752 -736 0 feedthrough
rlabel pdiffusion 759 -736 759 -736 0 feedthrough
rlabel pdiffusion 766 -736 766 -736 0 feedthrough
rlabel pdiffusion 773 -736 773 -736 0 feedthrough
rlabel pdiffusion 780 -736 780 -736 0 feedthrough
rlabel pdiffusion 787 -736 787 -736 0 feedthrough
rlabel pdiffusion 794 -736 794 -736 0 feedthrough
rlabel pdiffusion 801 -736 801 -736 0 feedthrough
rlabel pdiffusion 808 -736 808 -736 0 feedthrough
rlabel pdiffusion 815 -736 815 -736 0 feedthrough
rlabel pdiffusion 822 -736 822 -736 0 feedthrough
rlabel pdiffusion 829 -736 829 -736 0 feedthrough
rlabel pdiffusion 836 -736 836 -736 0 feedthrough
rlabel pdiffusion 843 -736 843 -736 0 feedthrough
rlabel pdiffusion 850 -736 850 -736 0 feedthrough
rlabel pdiffusion 857 -736 857 -736 0 feedthrough
rlabel pdiffusion 864 -736 864 -736 0 feedthrough
rlabel pdiffusion 871 -736 871 -736 0 feedthrough
rlabel pdiffusion 878 -736 878 -736 0 feedthrough
rlabel pdiffusion 885 -736 885 -736 0 feedthrough
rlabel pdiffusion 892 -736 892 -736 0 feedthrough
rlabel pdiffusion 899 -736 899 -736 0 feedthrough
rlabel pdiffusion 906 -736 906 -736 0 feedthrough
rlabel pdiffusion 913 -736 913 -736 0 feedthrough
rlabel pdiffusion 920 -736 920 -736 0 feedthrough
rlabel pdiffusion 927 -736 927 -736 0 feedthrough
rlabel pdiffusion 934 -736 934 -736 0 feedthrough
rlabel pdiffusion 941 -736 941 -736 0 feedthrough
rlabel pdiffusion 948 -736 948 -736 0 feedthrough
rlabel pdiffusion 955 -736 955 -736 0 feedthrough
rlabel pdiffusion 962 -736 962 -736 0 feedthrough
rlabel pdiffusion 969 -736 969 -736 0 feedthrough
rlabel pdiffusion 976 -736 976 -736 0 feedthrough
rlabel pdiffusion 983 -736 983 -736 0 feedthrough
rlabel pdiffusion 990 -736 990 -736 0 feedthrough
rlabel pdiffusion 997 -736 997 -736 0 feedthrough
rlabel pdiffusion 1004 -736 1004 -736 0 feedthrough
rlabel pdiffusion 1011 -736 1011 -736 0 feedthrough
rlabel pdiffusion 1018 -736 1018 -736 0 feedthrough
rlabel pdiffusion 1025 -736 1025 -736 0 feedthrough
rlabel pdiffusion 1032 -736 1032 -736 0 feedthrough
rlabel pdiffusion 1039 -736 1039 -736 0 feedthrough
rlabel pdiffusion 1046 -736 1046 -736 0 feedthrough
rlabel pdiffusion 1053 -736 1053 -736 0 feedthrough
rlabel pdiffusion 1060 -736 1060 -736 0 feedthrough
rlabel pdiffusion 1067 -736 1067 -736 0 feedthrough
rlabel pdiffusion 1074 -736 1074 -736 0 feedthrough
rlabel pdiffusion 1081 -736 1081 -736 0 feedthrough
rlabel pdiffusion 1088 -736 1088 -736 0 cellNo=124
rlabel pdiffusion 1095 -736 1095 -736 0 feedthrough
rlabel pdiffusion 1102 -736 1102 -736 0 feedthrough
rlabel pdiffusion 1109 -736 1109 -736 0 cellNo=461
rlabel pdiffusion 1116 -736 1116 -736 0 feedthrough
rlabel pdiffusion 1123 -736 1123 -736 0 feedthrough
rlabel pdiffusion 1130 -736 1130 -736 0 feedthrough
rlabel pdiffusion 1137 -736 1137 -736 0 feedthrough
rlabel pdiffusion 1144 -736 1144 -736 0 feedthrough
rlabel pdiffusion 1151 -736 1151 -736 0 feedthrough
rlabel pdiffusion 1158 -736 1158 -736 0 cellNo=158
rlabel pdiffusion 1165 -736 1165 -736 0 feedthrough
rlabel pdiffusion 1172 -736 1172 -736 0 feedthrough
rlabel pdiffusion 1186 -736 1186 -736 0 feedthrough
rlabel pdiffusion 3 -825 3 -825 0 cellNo=156
rlabel pdiffusion 10 -825 10 -825 0 feedthrough
rlabel pdiffusion 17 -825 17 -825 0 feedthrough
rlabel pdiffusion 24 -825 24 -825 0 feedthrough
rlabel pdiffusion 31 -825 31 -825 0 feedthrough
rlabel pdiffusion 38 -825 38 -825 0 feedthrough
rlabel pdiffusion 45 -825 45 -825 0 feedthrough
rlabel pdiffusion 52 -825 52 -825 0 feedthrough
rlabel pdiffusion 59 -825 59 -825 0 feedthrough
rlabel pdiffusion 66 -825 66 -825 0 feedthrough
rlabel pdiffusion 73 -825 73 -825 0 cellNo=546
rlabel pdiffusion 80 -825 80 -825 0 feedthrough
rlabel pdiffusion 87 -825 87 -825 0 feedthrough
rlabel pdiffusion 94 -825 94 -825 0 feedthrough
rlabel pdiffusion 101 -825 101 -825 0 feedthrough
rlabel pdiffusion 108 -825 108 -825 0 feedthrough
rlabel pdiffusion 115 -825 115 -825 0 cellNo=612
rlabel pdiffusion 122 -825 122 -825 0 cellNo=893
rlabel pdiffusion 129 -825 129 -825 0 cellNo=181
rlabel pdiffusion 136 -825 136 -825 0 cellNo=268
rlabel pdiffusion 143 -825 143 -825 0 feedthrough
rlabel pdiffusion 150 -825 150 -825 0 feedthrough
rlabel pdiffusion 157 -825 157 -825 0 feedthrough
rlabel pdiffusion 164 -825 164 -825 0 cellNo=396
rlabel pdiffusion 171 -825 171 -825 0 cellNo=872
rlabel pdiffusion 178 -825 178 -825 0 feedthrough
rlabel pdiffusion 185 -825 185 -825 0 feedthrough
rlabel pdiffusion 192 -825 192 -825 0 feedthrough
rlabel pdiffusion 199 -825 199 -825 0 feedthrough
rlabel pdiffusion 206 -825 206 -825 0 feedthrough
rlabel pdiffusion 213 -825 213 -825 0 feedthrough
rlabel pdiffusion 220 -825 220 -825 0 feedthrough
rlabel pdiffusion 227 -825 227 -825 0 feedthrough
rlabel pdiffusion 234 -825 234 -825 0 feedthrough
rlabel pdiffusion 241 -825 241 -825 0 feedthrough
rlabel pdiffusion 248 -825 248 -825 0 feedthrough
rlabel pdiffusion 255 -825 255 -825 0 feedthrough
rlabel pdiffusion 262 -825 262 -825 0 cellNo=408
rlabel pdiffusion 269 -825 269 -825 0 feedthrough
rlabel pdiffusion 276 -825 276 -825 0 feedthrough
rlabel pdiffusion 283 -825 283 -825 0 feedthrough
rlabel pdiffusion 290 -825 290 -825 0 feedthrough
rlabel pdiffusion 297 -825 297 -825 0 feedthrough
rlabel pdiffusion 304 -825 304 -825 0 feedthrough
rlabel pdiffusion 311 -825 311 -825 0 feedthrough
rlabel pdiffusion 318 -825 318 -825 0 feedthrough
rlabel pdiffusion 325 -825 325 -825 0 feedthrough
rlabel pdiffusion 332 -825 332 -825 0 feedthrough
rlabel pdiffusion 339 -825 339 -825 0 feedthrough
rlabel pdiffusion 346 -825 346 -825 0 feedthrough
rlabel pdiffusion 353 -825 353 -825 0 cellNo=337
rlabel pdiffusion 360 -825 360 -825 0 cellNo=358
rlabel pdiffusion 367 -825 367 -825 0 feedthrough
rlabel pdiffusion 374 -825 374 -825 0 feedthrough
rlabel pdiffusion 381 -825 381 -825 0 cellNo=100
rlabel pdiffusion 388 -825 388 -825 0 feedthrough
rlabel pdiffusion 395 -825 395 -825 0 feedthrough
rlabel pdiffusion 402 -825 402 -825 0 feedthrough
rlabel pdiffusion 409 -825 409 -825 0 feedthrough
rlabel pdiffusion 416 -825 416 -825 0 feedthrough
rlabel pdiffusion 423 -825 423 -825 0 cellNo=391
rlabel pdiffusion 430 -825 430 -825 0 feedthrough
rlabel pdiffusion 437 -825 437 -825 0 feedthrough
rlabel pdiffusion 444 -825 444 -825 0 feedthrough
rlabel pdiffusion 451 -825 451 -825 0 feedthrough
rlabel pdiffusion 458 -825 458 -825 0 feedthrough
rlabel pdiffusion 465 -825 465 -825 0 feedthrough
rlabel pdiffusion 472 -825 472 -825 0 feedthrough
rlabel pdiffusion 479 -825 479 -825 0 cellNo=392
rlabel pdiffusion 486 -825 486 -825 0 feedthrough
rlabel pdiffusion 493 -825 493 -825 0 cellNo=4
rlabel pdiffusion 500 -825 500 -825 0 cellNo=65
rlabel pdiffusion 507 -825 507 -825 0 feedthrough
rlabel pdiffusion 514 -825 514 -825 0 feedthrough
rlabel pdiffusion 521 -825 521 -825 0 cellNo=848
rlabel pdiffusion 528 -825 528 -825 0 feedthrough
rlabel pdiffusion 535 -825 535 -825 0 feedthrough
rlabel pdiffusion 542 -825 542 -825 0 feedthrough
rlabel pdiffusion 549 -825 549 -825 0 feedthrough
rlabel pdiffusion 556 -825 556 -825 0 cellNo=149
rlabel pdiffusion 563 -825 563 -825 0 cellNo=136
rlabel pdiffusion 570 -825 570 -825 0 cellNo=851
rlabel pdiffusion 577 -825 577 -825 0 feedthrough
rlabel pdiffusion 584 -825 584 -825 0 feedthrough
rlabel pdiffusion 591 -825 591 -825 0 feedthrough
rlabel pdiffusion 598 -825 598 -825 0 feedthrough
rlabel pdiffusion 605 -825 605 -825 0 feedthrough
rlabel pdiffusion 612 -825 612 -825 0 feedthrough
rlabel pdiffusion 619 -825 619 -825 0 cellNo=450
rlabel pdiffusion 626 -825 626 -825 0 cellNo=420
rlabel pdiffusion 633 -825 633 -825 0 feedthrough
rlabel pdiffusion 640 -825 640 -825 0 cellNo=393
rlabel pdiffusion 647 -825 647 -825 0 feedthrough
rlabel pdiffusion 654 -825 654 -825 0 cellNo=263
rlabel pdiffusion 661 -825 661 -825 0 cellNo=735
rlabel pdiffusion 668 -825 668 -825 0 feedthrough
rlabel pdiffusion 675 -825 675 -825 0 feedthrough
rlabel pdiffusion 682 -825 682 -825 0 feedthrough
rlabel pdiffusion 689 -825 689 -825 0 feedthrough
rlabel pdiffusion 696 -825 696 -825 0 cellNo=204
rlabel pdiffusion 703 -825 703 -825 0 feedthrough
rlabel pdiffusion 710 -825 710 -825 0 feedthrough
rlabel pdiffusion 717 -825 717 -825 0 feedthrough
rlabel pdiffusion 724 -825 724 -825 0 cellNo=650
rlabel pdiffusion 731 -825 731 -825 0 feedthrough
rlabel pdiffusion 738 -825 738 -825 0 feedthrough
rlabel pdiffusion 745 -825 745 -825 0 feedthrough
rlabel pdiffusion 752 -825 752 -825 0 feedthrough
rlabel pdiffusion 759 -825 759 -825 0 feedthrough
rlabel pdiffusion 766 -825 766 -825 0 feedthrough
rlabel pdiffusion 773 -825 773 -825 0 feedthrough
rlabel pdiffusion 780 -825 780 -825 0 cellNo=496
rlabel pdiffusion 787 -825 787 -825 0 feedthrough
rlabel pdiffusion 794 -825 794 -825 0 feedthrough
rlabel pdiffusion 801 -825 801 -825 0 feedthrough
rlabel pdiffusion 808 -825 808 -825 0 feedthrough
rlabel pdiffusion 815 -825 815 -825 0 cellNo=286
rlabel pdiffusion 822 -825 822 -825 0 feedthrough
rlabel pdiffusion 829 -825 829 -825 0 feedthrough
rlabel pdiffusion 836 -825 836 -825 0 feedthrough
rlabel pdiffusion 843 -825 843 -825 0 feedthrough
rlabel pdiffusion 850 -825 850 -825 0 cellNo=717
rlabel pdiffusion 857 -825 857 -825 0 feedthrough
rlabel pdiffusion 864 -825 864 -825 0 feedthrough
rlabel pdiffusion 871 -825 871 -825 0 feedthrough
rlabel pdiffusion 878 -825 878 -825 0 feedthrough
rlabel pdiffusion 885 -825 885 -825 0 feedthrough
rlabel pdiffusion 892 -825 892 -825 0 feedthrough
rlabel pdiffusion 899 -825 899 -825 0 feedthrough
rlabel pdiffusion 906 -825 906 -825 0 feedthrough
rlabel pdiffusion 913 -825 913 -825 0 feedthrough
rlabel pdiffusion 920 -825 920 -825 0 feedthrough
rlabel pdiffusion 927 -825 927 -825 0 feedthrough
rlabel pdiffusion 934 -825 934 -825 0 feedthrough
rlabel pdiffusion 941 -825 941 -825 0 feedthrough
rlabel pdiffusion 948 -825 948 -825 0 feedthrough
rlabel pdiffusion 955 -825 955 -825 0 feedthrough
rlabel pdiffusion 962 -825 962 -825 0 feedthrough
rlabel pdiffusion 969 -825 969 -825 0 feedthrough
rlabel pdiffusion 976 -825 976 -825 0 feedthrough
rlabel pdiffusion 983 -825 983 -825 0 feedthrough
rlabel pdiffusion 990 -825 990 -825 0 feedthrough
rlabel pdiffusion 997 -825 997 -825 0 feedthrough
rlabel pdiffusion 1004 -825 1004 -825 0 feedthrough
rlabel pdiffusion 1011 -825 1011 -825 0 feedthrough
rlabel pdiffusion 1018 -825 1018 -825 0 feedthrough
rlabel pdiffusion 1025 -825 1025 -825 0 feedthrough
rlabel pdiffusion 1032 -825 1032 -825 0 feedthrough
rlabel pdiffusion 1039 -825 1039 -825 0 feedthrough
rlabel pdiffusion 1046 -825 1046 -825 0 feedthrough
rlabel pdiffusion 1053 -825 1053 -825 0 feedthrough
rlabel pdiffusion 1060 -825 1060 -825 0 feedthrough
rlabel pdiffusion 1067 -825 1067 -825 0 feedthrough
rlabel pdiffusion 1074 -825 1074 -825 0 feedthrough
rlabel pdiffusion 1081 -825 1081 -825 0 feedthrough
rlabel pdiffusion 1088 -825 1088 -825 0 feedthrough
rlabel pdiffusion 1095 -825 1095 -825 0 feedthrough
rlabel pdiffusion 1102 -825 1102 -825 0 feedthrough
rlabel pdiffusion 1109 -825 1109 -825 0 feedthrough
rlabel pdiffusion 1116 -825 1116 -825 0 feedthrough
rlabel pdiffusion 1123 -825 1123 -825 0 feedthrough
rlabel pdiffusion 1130 -825 1130 -825 0 feedthrough
rlabel pdiffusion 1137 -825 1137 -825 0 feedthrough
rlabel pdiffusion 1144 -825 1144 -825 0 feedthrough
rlabel pdiffusion 1151 -825 1151 -825 0 feedthrough
rlabel pdiffusion 1158 -825 1158 -825 0 feedthrough
rlabel pdiffusion 1165 -825 1165 -825 0 feedthrough
rlabel pdiffusion 1172 -825 1172 -825 0 feedthrough
rlabel pdiffusion 1179 -825 1179 -825 0 feedthrough
rlabel pdiffusion 1186 -825 1186 -825 0 feedthrough
rlabel pdiffusion 1193 -825 1193 -825 0 feedthrough
rlabel pdiffusion 1200 -825 1200 -825 0 feedthrough
rlabel pdiffusion 1207 -825 1207 -825 0 feedthrough
rlabel pdiffusion 1214 -825 1214 -825 0 feedthrough
rlabel pdiffusion 1221 -825 1221 -825 0 feedthrough
rlabel pdiffusion 3 -912 3 -912 0 cellNo=103
rlabel pdiffusion 10 -912 10 -912 0 feedthrough
rlabel pdiffusion 17 -912 17 -912 0 cellNo=487
rlabel pdiffusion 24 -912 24 -912 0 feedthrough
rlabel pdiffusion 31 -912 31 -912 0 cellNo=723
rlabel pdiffusion 38 -912 38 -912 0 cellNo=50
rlabel pdiffusion 45 -912 45 -912 0 feedthrough
rlabel pdiffusion 52 -912 52 -912 0 feedthrough
rlabel pdiffusion 59 -912 59 -912 0 feedthrough
rlabel pdiffusion 66 -912 66 -912 0 feedthrough
rlabel pdiffusion 73 -912 73 -912 0 cellNo=567
rlabel pdiffusion 80 -912 80 -912 0 feedthrough
rlabel pdiffusion 87 -912 87 -912 0 feedthrough
rlabel pdiffusion 94 -912 94 -912 0 feedthrough
rlabel pdiffusion 101 -912 101 -912 0 feedthrough
rlabel pdiffusion 108 -912 108 -912 0 feedthrough
rlabel pdiffusion 115 -912 115 -912 0 cellNo=701
rlabel pdiffusion 122 -912 122 -912 0 feedthrough
rlabel pdiffusion 129 -912 129 -912 0 cellNo=586
rlabel pdiffusion 136 -912 136 -912 0 feedthrough
rlabel pdiffusion 143 -912 143 -912 0 feedthrough
rlabel pdiffusion 150 -912 150 -912 0 cellNo=565
rlabel pdiffusion 157 -912 157 -912 0 feedthrough
rlabel pdiffusion 164 -912 164 -912 0 feedthrough
rlabel pdiffusion 171 -912 171 -912 0 feedthrough
rlabel pdiffusion 178 -912 178 -912 0 feedthrough
rlabel pdiffusion 185 -912 185 -912 0 feedthrough
rlabel pdiffusion 192 -912 192 -912 0 feedthrough
rlabel pdiffusion 199 -912 199 -912 0 feedthrough
rlabel pdiffusion 206 -912 206 -912 0 cellNo=739
rlabel pdiffusion 213 -912 213 -912 0 feedthrough
rlabel pdiffusion 220 -912 220 -912 0 feedthrough
rlabel pdiffusion 227 -912 227 -912 0 feedthrough
rlabel pdiffusion 234 -912 234 -912 0 feedthrough
rlabel pdiffusion 241 -912 241 -912 0 feedthrough
rlabel pdiffusion 248 -912 248 -912 0 feedthrough
rlabel pdiffusion 255 -912 255 -912 0 feedthrough
rlabel pdiffusion 262 -912 262 -912 0 cellNo=414
rlabel pdiffusion 269 -912 269 -912 0 feedthrough
rlabel pdiffusion 276 -912 276 -912 0 cellNo=336
rlabel pdiffusion 283 -912 283 -912 0 feedthrough
rlabel pdiffusion 290 -912 290 -912 0 cellNo=570
rlabel pdiffusion 297 -912 297 -912 0 feedthrough
rlabel pdiffusion 304 -912 304 -912 0 feedthrough
rlabel pdiffusion 311 -912 311 -912 0 cellNo=664
rlabel pdiffusion 318 -912 318 -912 0 feedthrough
rlabel pdiffusion 325 -912 325 -912 0 feedthrough
rlabel pdiffusion 332 -912 332 -912 0 feedthrough
rlabel pdiffusion 339 -912 339 -912 0 feedthrough
rlabel pdiffusion 346 -912 346 -912 0 cellNo=699
rlabel pdiffusion 353 -912 353 -912 0 feedthrough
rlabel pdiffusion 360 -912 360 -912 0 feedthrough
rlabel pdiffusion 367 -912 367 -912 0 feedthrough
rlabel pdiffusion 374 -912 374 -912 0 cellNo=518
rlabel pdiffusion 381 -912 381 -912 0 feedthrough
rlabel pdiffusion 388 -912 388 -912 0 feedthrough
rlabel pdiffusion 395 -912 395 -912 0 feedthrough
rlabel pdiffusion 402 -912 402 -912 0 feedthrough
rlabel pdiffusion 409 -912 409 -912 0 feedthrough
rlabel pdiffusion 416 -912 416 -912 0 feedthrough
rlabel pdiffusion 423 -912 423 -912 0 cellNo=656
rlabel pdiffusion 430 -912 430 -912 0 feedthrough
rlabel pdiffusion 437 -912 437 -912 0 cellNo=367
rlabel pdiffusion 444 -912 444 -912 0 feedthrough
rlabel pdiffusion 451 -912 451 -912 0 feedthrough
rlabel pdiffusion 458 -912 458 -912 0 feedthrough
rlabel pdiffusion 465 -912 465 -912 0 feedthrough
rlabel pdiffusion 472 -912 472 -912 0 feedthrough
rlabel pdiffusion 479 -912 479 -912 0 cellNo=191
rlabel pdiffusion 486 -912 486 -912 0 feedthrough
rlabel pdiffusion 493 -912 493 -912 0 feedthrough
rlabel pdiffusion 500 -912 500 -912 0 feedthrough
rlabel pdiffusion 507 -912 507 -912 0 feedthrough
rlabel pdiffusion 514 -912 514 -912 0 feedthrough
rlabel pdiffusion 521 -912 521 -912 0 feedthrough
rlabel pdiffusion 528 -912 528 -912 0 feedthrough
rlabel pdiffusion 535 -912 535 -912 0 feedthrough
rlabel pdiffusion 542 -912 542 -912 0 cellNo=32
rlabel pdiffusion 549 -912 549 -912 0 feedthrough
rlabel pdiffusion 556 -912 556 -912 0 cellNo=883
rlabel pdiffusion 563 -912 563 -912 0 feedthrough
rlabel pdiffusion 570 -912 570 -912 0 feedthrough
rlabel pdiffusion 577 -912 577 -912 0 feedthrough
rlabel pdiffusion 584 -912 584 -912 0 feedthrough
rlabel pdiffusion 591 -912 591 -912 0 feedthrough
rlabel pdiffusion 598 -912 598 -912 0 cellNo=162
rlabel pdiffusion 605 -912 605 -912 0 feedthrough
rlabel pdiffusion 612 -912 612 -912 0 cellNo=537
rlabel pdiffusion 619 -912 619 -912 0 cellNo=516
rlabel pdiffusion 626 -912 626 -912 0 feedthrough
rlabel pdiffusion 633 -912 633 -912 0 feedthrough
rlabel pdiffusion 640 -912 640 -912 0 feedthrough
rlabel pdiffusion 647 -912 647 -912 0 feedthrough
rlabel pdiffusion 654 -912 654 -912 0 cellNo=704
rlabel pdiffusion 661 -912 661 -912 0 feedthrough
rlabel pdiffusion 668 -912 668 -912 0 cellNo=74
rlabel pdiffusion 675 -912 675 -912 0 cellNo=269
rlabel pdiffusion 682 -912 682 -912 0 cellNo=549
rlabel pdiffusion 689 -912 689 -912 0 feedthrough
rlabel pdiffusion 696 -912 696 -912 0 feedthrough
rlabel pdiffusion 703 -912 703 -912 0 feedthrough
rlabel pdiffusion 710 -912 710 -912 0 feedthrough
rlabel pdiffusion 717 -912 717 -912 0 feedthrough
rlabel pdiffusion 724 -912 724 -912 0 feedthrough
rlabel pdiffusion 731 -912 731 -912 0 feedthrough
rlabel pdiffusion 738 -912 738 -912 0 feedthrough
rlabel pdiffusion 745 -912 745 -912 0 feedthrough
rlabel pdiffusion 752 -912 752 -912 0 feedthrough
rlabel pdiffusion 759 -912 759 -912 0 feedthrough
rlabel pdiffusion 766 -912 766 -912 0 feedthrough
rlabel pdiffusion 773 -912 773 -912 0 feedthrough
rlabel pdiffusion 780 -912 780 -912 0 feedthrough
rlabel pdiffusion 787 -912 787 -912 0 feedthrough
rlabel pdiffusion 794 -912 794 -912 0 feedthrough
rlabel pdiffusion 801 -912 801 -912 0 feedthrough
rlabel pdiffusion 808 -912 808 -912 0 feedthrough
rlabel pdiffusion 815 -912 815 -912 0 feedthrough
rlabel pdiffusion 822 -912 822 -912 0 cellNo=327
rlabel pdiffusion 829 -912 829 -912 0 feedthrough
rlabel pdiffusion 836 -912 836 -912 0 feedthrough
rlabel pdiffusion 843 -912 843 -912 0 feedthrough
rlabel pdiffusion 850 -912 850 -912 0 feedthrough
rlabel pdiffusion 857 -912 857 -912 0 feedthrough
rlabel pdiffusion 864 -912 864 -912 0 feedthrough
rlabel pdiffusion 871 -912 871 -912 0 feedthrough
rlabel pdiffusion 878 -912 878 -912 0 feedthrough
rlabel pdiffusion 885 -912 885 -912 0 feedthrough
rlabel pdiffusion 892 -912 892 -912 0 feedthrough
rlabel pdiffusion 899 -912 899 -912 0 cellNo=453
rlabel pdiffusion 906 -912 906 -912 0 feedthrough
rlabel pdiffusion 913 -912 913 -912 0 feedthrough
rlabel pdiffusion 920 -912 920 -912 0 feedthrough
rlabel pdiffusion 927 -912 927 -912 0 feedthrough
rlabel pdiffusion 934 -912 934 -912 0 feedthrough
rlabel pdiffusion 941 -912 941 -912 0 feedthrough
rlabel pdiffusion 948 -912 948 -912 0 feedthrough
rlabel pdiffusion 955 -912 955 -912 0 feedthrough
rlabel pdiffusion 962 -912 962 -912 0 feedthrough
rlabel pdiffusion 969 -912 969 -912 0 feedthrough
rlabel pdiffusion 976 -912 976 -912 0 feedthrough
rlabel pdiffusion 983 -912 983 -912 0 feedthrough
rlabel pdiffusion 990 -912 990 -912 0 feedthrough
rlabel pdiffusion 997 -912 997 -912 0 feedthrough
rlabel pdiffusion 1004 -912 1004 -912 0 feedthrough
rlabel pdiffusion 1011 -912 1011 -912 0 feedthrough
rlabel pdiffusion 1018 -912 1018 -912 0 feedthrough
rlabel pdiffusion 1025 -912 1025 -912 0 feedthrough
rlabel pdiffusion 1032 -912 1032 -912 0 feedthrough
rlabel pdiffusion 1039 -912 1039 -912 0 feedthrough
rlabel pdiffusion 1046 -912 1046 -912 0 feedthrough
rlabel pdiffusion 1053 -912 1053 -912 0 feedthrough
rlabel pdiffusion 1060 -912 1060 -912 0 feedthrough
rlabel pdiffusion 1067 -912 1067 -912 0 feedthrough
rlabel pdiffusion 1074 -912 1074 -912 0 feedthrough
rlabel pdiffusion 1081 -912 1081 -912 0 feedthrough
rlabel pdiffusion 1088 -912 1088 -912 0 cellNo=280
rlabel pdiffusion 1095 -912 1095 -912 0 feedthrough
rlabel pdiffusion 1102 -912 1102 -912 0 feedthrough
rlabel pdiffusion 1109 -912 1109 -912 0 feedthrough
rlabel pdiffusion 1116 -912 1116 -912 0 feedthrough
rlabel pdiffusion 1123 -912 1123 -912 0 feedthrough
rlabel pdiffusion 1130 -912 1130 -912 0 feedthrough
rlabel pdiffusion 1165 -912 1165 -912 0 feedthrough
rlabel pdiffusion 1172 -912 1172 -912 0 feedthrough
rlabel pdiffusion 1179 -912 1179 -912 0 feedthrough
rlabel pdiffusion 1193 -912 1193 -912 0 feedthrough
rlabel pdiffusion 3 -1001 3 -1001 0 feedthrough
rlabel pdiffusion 10 -1001 10 -1001 0 feedthrough
rlabel pdiffusion 17 -1001 17 -1001 0 cellNo=157
rlabel pdiffusion 24 -1001 24 -1001 0 feedthrough
rlabel pdiffusion 31 -1001 31 -1001 0 feedthrough
rlabel pdiffusion 38 -1001 38 -1001 0 cellNo=822
rlabel pdiffusion 45 -1001 45 -1001 0 feedthrough
rlabel pdiffusion 52 -1001 52 -1001 0 feedthrough
rlabel pdiffusion 59 -1001 59 -1001 0 cellNo=740
rlabel pdiffusion 66 -1001 66 -1001 0 cellNo=651
rlabel pdiffusion 73 -1001 73 -1001 0 feedthrough
rlabel pdiffusion 80 -1001 80 -1001 0 feedthrough
rlabel pdiffusion 87 -1001 87 -1001 0 feedthrough
rlabel pdiffusion 94 -1001 94 -1001 0 cellNo=75
rlabel pdiffusion 101 -1001 101 -1001 0 cellNo=440
rlabel pdiffusion 108 -1001 108 -1001 0 feedthrough
rlabel pdiffusion 115 -1001 115 -1001 0 feedthrough
rlabel pdiffusion 122 -1001 122 -1001 0 cellNo=39
rlabel pdiffusion 129 -1001 129 -1001 0 feedthrough
rlabel pdiffusion 136 -1001 136 -1001 0 feedthrough
rlabel pdiffusion 143 -1001 143 -1001 0 feedthrough
rlabel pdiffusion 150 -1001 150 -1001 0 feedthrough
rlabel pdiffusion 157 -1001 157 -1001 0 feedthrough
rlabel pdiffusion 164 -1001 164 -1001 0 feedthrough
rlabel pdiffusion 171 -1001 171 -1001 0 feedthrough
rlabel pdiffusion 178 -1001 178 -1001 0 feedthrough
rlabel pdiffusion 185 -1001 185 -1001 0 cellNo=896
rlabel pdiffusion 192 -1001 192 -1001 0 feedthrough
rlabel pdiffusion 199 -1001 199 -1001 0 cellNo=27
rlabel pdiffusion 206 -1001 206 -1001 0 feedthrough
rlabel pdiffusion 213 -1001 213 -1001 0 feedthrough
rlabel pdiffusion 220 -1001 220 -1001 0 feedthrough
rlabel pdiffusion 227 -1001 227 -1001 0 feedthrough
rlabel pdiffusion 234 -1001 234 -1001 0 feedthrough
rlabel pdiffusion 241 -1001 241 -1001 0 feedthrough
rlabel pdiffusion 248 -1001 248 -1001 0 feedthrough
rlabel pdiffusion 255 -1001 255 -1001 0 feedthrough
rlabel pdiffusion 262 -1001 262 -1001 0 feedthrough
rlabel pdiffusion 269 -1001 269 -1001 0 feedthrough
rlabel pdiffusion 276 -1001 276 -1001 0 feedthrough
rlabel pdiffusion 283 -1001 283 -1001 0 feedthrough
rlabel pdiffusion 290 -1001 290 -1001 0 feedthrough
rlabel pdiffusion 297 -1001 297 -1001 0 feedthrough
rlabel pdiffusion 304 -1001 304 -1001 0 feedthrough
rlabel pdiffusion 311 -1001 311 -1001 0 feedthrough
rlabel pdiffusion 318 -1001 318 -1001 0 feedthrough
rlabel pdiffusion 325 -1001 325 -1001 0 feedthrough
rlabel pdiffusion 332 -1001 332 -1001 0 feedthrough
rlabel pdiffusion 339 -1001 339 -1001 0 feedthrough
rlabel pdiffusion 346 -1001 346 -1001 0 feedthrough
rlabel pdiffusion 353 -1001 353 -1001 0 feedthrough
rlabel pdiffusion 360 -1001 360 -1001 0 cellNo=114
rlabel pdiffusion 367 -1001 367 -1001 0 feedthrough
rlabel pdiffusion 374 -1001 374 -1001 0 cellNo=499
rlabel pdiffusion 381 -1001 381 -1001 0 feedthrough
rlabel pdiffusion 388 -1001 388 -1001 0 cellNo=41
rlabel pdiffusion 395 -1001 395 -1001 0 feedthrough
rlabel pdiffusion 402 -1001 402 -1001 0 feedthrough
rlabel pdiffusion 409 -1001 409 -1001 0 feedthrough
rlabel pdiffusion 416 -1001 416 -1001 0 feedthrough
rlabel pdiffusion 423 -1001 423 -1001 0 feedthrough
rlabel pdiffusion 430 -1001 430 -1001 0 feedthrough
rlabel pdiffusion 437 -1001 437 -1001 0 cellNo=742
rlabel pdiffusion 444 -1001 444 -1001 0 feedthrough
rlabel pdiffusion 451 -1001 451 -1001 0 feedthrough
rlabel pdiffusion 458 -1001 458 -1001 0 feedthrough
rlabel pdiffusion 465 -1001 465 -1001 0 cellNo=478
rlabel pdiffusion 472 -1001 472 -1001 0 feedthrough
rlabel pdiffusion 479 -1001 479 -1001 0 feedthrough
rlabel pdiffusion 486 -1001 486 -1001 0 feedthrough
rlabel pdiffusion 493 -1001 493 -1001 0 feedthrough
rlabel pdiffusion 500 -1001 500 -1001 0 cellNo=462
rlabel pdiffusion 507 -1001 507 -1001 0 cellNo=371
rlabel pdiffusion 514 -1001 514 -1001 0 feedthrough
rlabel pdiffusion 521 -1001 521 -1001 0 feedthrough
rlabel pdiffusion 528 -1001 528 -1001 0 feedthrough
rlabel pdiffusion 535 -1001 535 -1001 0 feedthrough
rlabel pdiffusion 542 -1001 542 -1001 0 cellNo=223
rlabel pdiffusion 549 -1001 549 -1001 0 feedthrough
rlabel pdiffusion 556 -1001 556 -1001 0 feedthrough
rlabel pdiffusion 563 -1001 563 -1001 0 feedthrough
rlabel pdiffusion 570 -1001 570 -1001 0 feedthrough
rlabel pdiffusion 577 -1001 577 -1001 0 feedthrough
rlabel pdiffusion 584 -1001 584 -1001 0 feedthrough
rlabel pdiffusion 591 -1001 591 -1001 0 feedthrough
rlabel pdiffusion 598 -1001 598 -1001 0 feedthrough
rlabel pdiffusion 605 -1001 605 -1001 0 cellNo=665
rlabel pdiffusion 612 -1001 612 -1001 0 feedthrough
rlabel pdiffusion 619 -1001 619 -1001 0 feedthrough
rlabel pdiffusion 626 -1001 626 -1001 0 cellNo=222
rlabel pdiffusion 633 -1001 633 -1001 0 feedthrough
rlabel pdiffusion 640 -1001 640 -1001 0 cellNo=133
rlabel pdiffusion 647 -1001 647 -1001 0 cellNo=359
rlabel pdiffusion 654 -1001 654 -1001 0 feedthrough
rlabel pdiffusion 661 -1001 661 -1001 0 feedthrough
rlabel pdiffusion 668 -1001 668 -1001 0 feedthrough
rlabel pdiffusion 675 -1001 675 -1001 0 feedthrough
rlabel pdiffusion 682 -1001 682 -1001 0 cellNo=126
rlabel pdiffusion 689 -1001 689 -1001 0 feedthrough
rlabel pdiffusion 696 -1001 696 -1001 0 cellNo=321
rlabel pdiffusion 703 -1001 703 -1001 0 feedthrough
rlabel pdiffusion 710 -1001 710 -1001 0 cellNo=323
rlabel pdiffusion 717 -1001 717 -1001 0 feedthrough
rlabel pdiffusion 724 -1001 724 -1001 0 feedthrough
rlabel pdiffusion 731 -1001 731 -1001 0 cellNo=125
rlabel pdiffusion 738 -1001 738 -1001 0 feedthrough
rlabel pdiffusion 745 -1001 745 -1001 0 feedthrough
rlabel pdiffusion 752 -1001 752 -1001 0 feedthrough
rlabel pdiffusion 759 -1001 759 -1001 0 feedthrough
rlabel pdiffusion 766 -1001 766 -1001 0 feedthrough
rlabel pdiffusion 773 -1001 773 -1001 0 feedthrough
rlabel pdiffusion 780 -1001 780 -1001 0 feedthrough
rlabel pdiffusion 787 -1001 787 -1001 0 feedthrough
rlabel pdiffusion 794 -1001 794 -1001 0 feedthrough
rlabel pdiffusion 801 -1001 801 -1001 0 feedthrough
rlabel pdiffusion 808 -1001 808 -1001 0 feedthrough
rlabel pdiffusion 815 -1001 815 -1001 0 feedthrough
rlabel pdiffusion 822 -1001 822 -1001 0 feedthrough
rlabel pdiffusion 829 -1001 829 -1001 0 feedthrough
rlabel pdiffusion 836 -1001 836 -1001 0 feedthrough
rlabel pdiffusion 843 -1001 843 -1001 0 feedthrough
rlabel pdiffusion 850 -1001 850 -1001 0 feedthrough
rlabel pdiffusion 857 -1001 857 -1001 0 cellNo=672
rlabel pdiffusion 864 -1001 864 -1001 0 feedthrough
rlabel pdiffusion 871 -1001 871 -1001 0 feedthrough
rlabel pdiffusion 878 -1001 878 -1001 0 feedthrough
rlabel pdiffusion 885 -1001 885 -1001 0 feedthrough
rlabel pdiffusion 892 -1001 892 -1001 0 feedthrough
rlabel pdiffusion 899 -1001 899 -1001 0 feedthrough
rlabel pdiffusion 906 -1001 906 -1001 0 feedthrough
rlabel pdiffusion 913 -1001 913 -1001 0 feedthrough
rlabel pdiffusion 920 -1001 920 -1001 0 feedthrough
rlabel pdiffusion 927 -1001 927 -1001 0 feedthrough
rlabel pdiffusion 934 -1001 934 -1001 0 feedthrough
rlabel pdiffusion 941 -1001 941 -1001 0 feedthrough
rlabel pdiffusion 948 -1001 948 -1001 0 feedthrough
rlabel pdiffusion 955 -1001 955 -1001 0 feedthrough
rlabel pdiffusion 962 -1001 962 -1001 0 feedthrough
rlabel pdiffusion 969 -1001 969 -1001 0 feedthrough
rlabel pdiffusion 976 -1001 976 -1001 0 feedthrough
rlabel pdiffusion 983 -1001 983 -1001 0 feedthrough
rlabel pdiffusion 990 -1001 990 -1001 0 feedthrough
rlabel pdiffusion 997 -1001 997 -1001 0 feedthrough
rlabel pdiffusion 1004 -1001 1004 -1001 0 feedthrough
rlabel pdiffusion 1011 -1001 1011 -1001 0 feedthrough
rlabel pdiffusion 1018 -1001 1018 -1001 0 feedthrough
rlabel pdiffusion 1025 -1001 1025 -1001 0 feedthrough
rlabel pdiffusion 1032 -1001 1032 -1001 0 feedthrough
rlabel pdiffusion 1039 -1001 1039 -1001 0 feedthrough
rlabel pdiffusion 1046 -1001 1046 -1001 0 feedthrough
rlabel pdiffusion 1053 -1001 1053 -1001 0 feedthrough
rlabel pdiffusion 1060 -1001 1060 -1001 0 feedthrough
rlabel pdiffusion 1067 -1001 1067 -1001 0 feedthrough
rlabel pdiffusion 1074 -1001 1074 -1001 0 feedthrough
rlabel pdiffusion 1081 -1001 1081 -1001 0 feedthrough
rlabel pdiffusion 1088 -1001 1088 -1001 0 feedthrough
rlabel pdiffusion 1095 -1001 1095 -1001 0 feedthrough
rlabel pdiffusion 1102 -1001 1102 -1001 0 feedthrough
rlabel pdiffusion 1109 -1001 1109 -1001 0 feedthrough
rlabel pdiffusion 1116 -1001 1116 -1001 0 feedthrough
rlabel pdiffusion 1123 -1001 1123 -1001 0 feedthrough
rlabel pdiffusion 1130 -1001 1130 -1001 0 cellNo=256
rlabel pdiffusion 1137 -1001 1137 -1001 0 cellNo=682
rlabel pdiffusion 1144 -1001 1144 -1001 0 feedthrough
rlabel pdiffusion 1151 -1001 1151 -1001 0 feedthrough
rlabel pdiffusion 1158 -1001 1158 -1001 0 feedthrough
rlabel pdiffusion 1165 -1001 1165 -1001 0 cellNo=224
rlabel pdiffusion 1172 -1001 1172 -1001 0 feedthrough
rlabel pdiffusion 1186 -1001 1186 -1001 0 feedthrough
rlabel pdiffusion 1193 -1001 1193 -1001 0 cellNo=237
rlabel pdiffusion 17 -1076 17 -1076 0 feedthrough
rlabel pdiffusion 24 -1076 24 -1076 0 feedthrough
rlabel pdiffusion 31 -1076 31 -1076 0 feedthrough
rlabel pdiffusion 38 -1076 38 -1076 0 feedthrough
rlabel pdiffusion 45 -1076 45 -1076 0 feedthrough
rlabel pdiffusion 52 -1076 52 -1076 0 feedthrough
rlabel pdiffusion 59 -1076 59 -1076 0 cellNo=62
rlabel pdiffusion 66 -1076 66 -1076 0 cellNo=18
rlabel pdiffusion 73 -1076 73 -1076 0 feedthrough
rlabel pdiffusion 80 -1076 80 -1076 0 feedthrough
rlabel pdiffusion 87 -1076 87 -1076 0 cellNo=226
rlabel pdiffusion 94 -1076 94 -1076 0 cellNo=137
rlabel pdiffusion 101 -1076 101 -1076 0 feedthrough
rlabel pdiffusion 108 -1076 108 -1076 0 feedthrough
rlabel pdiffusion 115 -1076 115 -1076 0 cellNo=432
rlabel pdiffusion 122 -1076 122 -1076 0 feedthrough
rlabel pdiffusion 129 -1076 129 -1076 0 feedthrough
rlabel pdiffusion 136 -1076 136 -1076 0 feedthrough
rlabel pdiffusion 143 -1076 143 -1076 0 feedthrough
rlabel pdiffusion 150 -1076 150 -1076 0 cellNo=86
rlabel pdiffusion 157 -1076 157 -1076 0 feedthrough
rlabel pdiffusion 164 -1076 164 -1076 0 feedthrough
rlabel pdiffusion 171 -1076 171 -1076 0 cellNo=331
rlabel pdiffusion 178 -1076 178 -1076 0 feedthrough
rlabel pdiffusion 185 -1076 185 -1076 0 feedthrough
rlabel pdiffusion 192 -1076 192 -1076 0 feedthrough
rlabel pdiffusion 199 -1076 199 -1076 0 feedthrough
rlabel pdiffusion 206 -1076 206 -1076 0 cellNo=84
rlabel pdiffusion 213 -1076 213 -1076 0 feedthrough
rlabel pdiffusion 220 -1076 220 -1076 0 feedthrough
rlabel pdiffusion 227 -1076 227 -1076 0 feedthrough
rlabel pdiffusion 234 -1076 234 -1076 0 feedthrough
rlabel pdiffusion 241 -1076 241 -1076 0 feedthrough
rlabel pdiffusion 248 -1076 248 -1076 0 feedthrough
rlabel pdiffusion 255 -1076 255 -1076 0 feedthrough
rlabel pdiffusion 262 -1076 262 -1076 0 cellNo=687
rlabel pdiffusion 269 -1076 269 -1076 0 feedthrough
rlabel pdiffusion 276 -1076 276 -1076 0 feedthrough
rlabel pdiffusion 283 -1076 283 -1076 0 feedthrough
rlabel pdiffusion 290 -1076 290 -1076 0 feedthrough
rlabel pdiffusion 297 -1076 297 -1076 0 cellNo=515
rlabel pdiffusion 304 -1076 304 -1076 0 feedthrough
rlabel pdiffusion 311 -1076 311 -1076 0 feedthrough
rlabel pdiffusion 318 -1076 318 -1076 0 cellNo=313
rlabel pdiffusion 325 -1076 325 -1076 0 feedthrough
rlabel pdiffusion 332 -1076 332 -1076 0 feedthrough
rlabel pdiffusion 339 -1076 339 -1076 0 feedthrough
rlabel pdiffusion 346 -1076 346 -1076 0 feedthrough
rlabel pdiffusion 353 -1076 353 -1076 0 cellNo=600
rlabel pdiffusion 360 -1076 360 -1076 0 feedthrough
rlabel pdiffusion 367 -1076 367 -1076 0 feedthrough
rlabel pdiffusion 374 -1076 374 -1076 0 feedthrough
rlabel pdiffusion 381 -1076 381 -1076 0 feedthrough
rlabel pdiffusion 388 -1076 388 -1076 0 feedthrough
rlabel pdiffusion 395 -1076 395 -1076 0 feedthrough
rlabel pdiffusion 402 -1076 402 -1076 0 feedthrough
rlabel pdiffusion 409 -1076 409 -1076 0 feedthrough
rlabel pdiffusion 416 -1076 416 -1076 0 feedthrough
rlabel pdiffusion 423 -1076 423 -1076 0 feedthrough
rlabel pdiffusion 430 -1076 430 -1076 0 feedthrough
rlabel pdiffusion 437 -1076 437 -1076 0 cellNo=301
rlabel pdiffusion 444 -1076 444 -1076 0 feedthrough
rlabel pdiffusion 451 -1076 451 -1076 0 feedthrough
rlabel pdiffusion 458 -1076 458 -1076 0 feedthrough
rlabel pdiffusion 465 -1076 465 -1076 0 cellNo=674
rlabel pdiffusion 472 -1076 472 -1076 0 feedthrough
rlabel pdiffusion 479 -1076 479 -1076 0 feedthrough
rlabel pdiffusion 486 -1076 486 -1076 0 feedthrough
rlabel pdiffusion 493 -1076 493 -1076 0 feedthrough
rlabel pdiffusion 500 -1076 500 -1076 0 feedthrough
rlabel pdiffusion 507 -1076 507 -1076 0 cellNo=374
rlabel pdiffusion 514 -1076 514 -1076 0 feedthrough
rlabel pdiffusion 521 -1076 521 -1076 0 feedthrough
rlabel pdiffusion 528 -1076 528 -1076 0 feedthrough
rlabel pdiffusion 535 -1076 535 -1076 0 cellNo=573
rlabel pdiffusion 542 -1076 542 -1076 0 feedthrough
rlabel pdiffusion 549 -1076 549 -1076 0 feedthrough
rlabel pdiffusion 556 -1076 556 -1076 0 feedthrough
rlabel pdiffusion 563 -1076 563 -1076 0 feedthrough
rlabel pdiffusion 570 -1076 570 -1076 0 cellNo=166
rlabel pdiffusion 577 -1076 577 -1076 0 feedthrough
rlabel pdiffusion 584 -1076 584 -1076 0 feedthrough
rlabel pdiffusion 591 -1076 591 -1076 0 feedthrough
rlabel pdiffusion 598 -1076 598 -1076 0 cellNo=574
rlabel pdiffusion 605 -1076 605 -1076 0 feedthrough
rlabel pdiffusion 612 -1076 612 -1076 0 feedthrough
rlabel pdiffusion 619 -1076 619 -1076 0 cellNo=890
rlabel pdiffusion 626 -1076 626 -1076 0 feedthrough
rlabel pdiffusion 633 -1076 633 -1076 0 cellNo=510
rlabel pdiffusion 640 -1076 640 -1076 0 feedthrough
rlabel pdiffusion 647 -1076 647 -1076 0 feedthrough
rlabel pdiffusion 654 -1076 654 -1076 0 feedthrough
rlabel pdiffusion 661 -1076 661 -1076 0 feedthrough
rlabel pdiffusion 668 -1076 668 -1076 0 feedthrough
rlabel pdiffusion 675 -1076 675 -1076 0 feedthrough
rlabel pdiffusion 682 -1076 682 -1076 0 feedthrough
rlabel pdiffusion 689 -1076 689 -1076 0 cellNo=514
rlabel pdiffusion 696 -1076 696 -1076 0 feedthrough
rlabel pdiffusion 703 -1076 703 -1076 0 feedthrough
rlabel pdiffusion 710 -1076 710 -1076 0 feedthrough
rlabel pdiffusion 717 -1076 717 -1076 0 feedthrough
rlabel pdiffusion 724 -1076 724 -1076 0 feedthrough
rlabel pdiffusion 731 -1076 731 -1076 0 cellNo=273
rlabel pdiffusion 738 -1076 738 -1076 0 feedthrough
rlabel pdiffusion 745 -1076 745 -1076 0 feedthrough
rlabel pdiffusion 752 -1076 752 -1076 0 feedthrough
rlabel pdiffusion 759 -1076 759 -1076 0 cellNo=247
rlabel pdiffusion 766 -1076 766 -1076 0 feedthrough
rlabel pdiffusion 773 -1076 773 -1076 0 feedthrough
rlabel pdiffusion 780 -1076 780 -1076 0 feedthrough
rlabel pdiffusion 787 -1076 787 -1076 0 feedthrough
rlabel pdiffusion 794 -1076 794 -1076 0 feedthrough
rlabel pdiffusion 801 -1076 801 -1076 0 feedthrough
rlabel pdiffusion 808 -1076 808 -1076 0 cellNo=676
rlabel pdiffusion 815 -1076 815 -1076 0 feedthrough
rlabel pdiffusion 822 -1076 822 -1076 0 feedthrough
rlabel pdiffusion 829 -1076 829 -1076 0 feedthrough
rlabel pdiffusion 836 -1076 836 -1076 0 feedthrough
rlabel pdiffusion 843 -1076 843 -1076 0 feedthrough
rlabel pdiffusion 850 -1076 850 -1076 0 feedthrough
rlabel pdiffusion 857 -1076 857 -1076 0 feedthrough
rlabel pdiffusion 864 -1076 864 -1076 0 feedthrough
rlabel pdiffusion 871 -1076 871 -1076 0 feedthrough
rlabel pdiffusion 878 -1076 878 -1076 0 feedthrough
rlabel pdiffusion 885 -1076 885 -1076 0 feedthrough
rlabel pdiffusion 892 -1076 892 -1076 0 feedthrough
rlabel pdiffusion 899 -1076 899 -1076 0 feedthrough
rlabel pdiffusion 906 -1076 906 -1076 0 feedthrough
rlabel pdiffusion 913 -1076 913 -1076 0 feedthrough
rlabel pdiffusion 920 -1076 920 -1076 0 cellNo=340
rlabel pdiffusion 927 -1076 927 -1076 0 feedthrough
rlabel pdiffusion 934 -1076 934 -1076 0 feedthrough
rlabel pdiffusion 941 -1076 941 -1076 0 feedthrough
rlabel pdiffusion 948 -1076 948 -1076 0 feedthrough
rlabel pdiffusion 955 -1076 955 -1076 0 cellNo=139
rlabel pdiffusion 962 -1076 962 -1076 0 feedthrough
rlabel pdiffusion 969 -1076 969 -1076 0 feedthrough
rlabel pdiffusion 976 -1076 976 -1076 0 feedthrough
rlabel pdiffusion 983 -1076 983 -1076 0 feedthrough
rlabel pdiffusion 990 -1076 990 -1076 0 feedthrough
rlabel pdiffusion 997 -1076 997 -1076 0 feedthrough
rlabel pdiffusion 1004 -1076 1004 -1076 0 feedthrough
rlabel pdiffusion 1011 -1076 1011 -1076 0 feedthrough
rlabel pdiffusion 1018 -1076 1018 -1076 0 feedthrough
rlabel pdiffusion 1025 -1076 1025 -1076 0 feedthrough
rlabel pdiffusion 1032 -1076 1032 -1076 0 cellNo=63
rlabel pdiffusion 1039 -1076 1039 -1076 0 cellNo=784
rlabel pdiffusion 1046 -1076 1046 -1076 0 feedthrough
rlabel pdiffusion 1053 -1076 1053 -1076 0 feedthrough
rlabel pdiffusion 1060 -1076 1060 -1076 0 cellNo=447
rlabel pdiffusion 1067 -1076 1067 -1076 0 cellNo=71
rlabel pdiffusion 1074 -1076 1074 -1076 0 feedthrough
rlabel pdiffusion 1081 -1076 1081 -1076 0 feedthrough
rlabel pdiffusion 1088 -1076 1088 -1076 0 feedthrough
rlabel pdiffusion 1095 -1076 1095 -1076 0 feedthrough
rlabel pdiffusion 1123 -1076 1123 -1076 0 feedthrough
rlabel pdiffusion 1186 -1076 1186 -1076 0 feedthrough
rlabel pdiffusion 24 -1159 24 -1159 0 cellNo=51
rlabel pdiffusion 31 -1159 31 -1159 0 feedthrough
rlabel pdiffusion 38 -1159 38 -1159 0 feedthrough
rlabel pdiffusion 45 -1159 45 -1159 0 feedthrough
rlabel pdiffusion 52 -1159 52 -1159 0 feedthrough
rlabel pdiffusion 59 -1159 59 -1159 0 feedthrough
rlabel pdiffusion 66 -1159 66 -1159 0 feedthrough
rlabel pdiffusion 73 -1159 73 -1159 0 feedthrough
rlabel pdiffusion 80 -1159 80 -1159 0 cellNo=681
rlabel pdiffusion 87 -1159 87 -1159 0 cellNo=377
rlabel pdiffusion 94 -1159 94 -1159 0 feedthrough
rlabel pdiffusion 101 -1159 101 -1159 0 feedthrough
rlabel pdiffusion 108 -1159 108 -1159 0 feedthrough
rlabel pdiffusion 115 -1159 115 -1159 0 cellNo=823
rlabel pdiffusion 122 -1159 122 -1159 0 feedthrough
rlabel pdiffusion 129 -1159 129 -1159 0 cellNo=239
rlabel pdiffusion 136 -1159 136 -1159 0 cellNo=16
rlabel pdiffusion 143 -1159 143 -1159 0 feedthrough
rlabel pdiffusion 150 -1159 150 -1159 0 feedthrough
rlabel pdiffusion 157 -1159 157 -1159 0 cellNo=513
rlabel pdiffusion 164 -1159 164 -1159 0 cellNo=855
rlabel pdiffusion 171 -1159 171 -1159 0 feedthrough
rlabel pdiffusion 178 -1159 178 -1159 0 feedthrough
rlabel pdiffusion 185 -1159 185 -1159 0 cellNo=481
rlabel pdiffusion 192 -1159 192 -1159 0 feedthrough
rlabel pdiffusion 199 -1159 199 -1159 0 cellNo=538
rlabel pdiffusion 206 -1159 206 -1159 0 feedthrough
rlabel pdiffusion 213 -1159 213 -1159 0 feedthrough
rlabel pdiffusion 220 -1159 220 -1159 0 feedthrough
rlabel pdiffusion 227 -1159 227 -1159 0 cellNo=492
rlabel pdiffusion 234 -1159 234 -1159 0 feedthrough
rlabel pdiffusion 241 -1159 241 -1159 0 feedthrough
rlabel pdiffusion 248 -1159 248 -1159 0 feedthrough
rlabel pdiffusion 255 -1159 255 -1159 0 feedthrough
rlabel pdiffusion 262 -1159 262 -1159 0 feedthrough
rlabel pdiffusion 269 -1159 269 -1159 0 feedthrough
rlabel pdiffusion 276 -1159 276 -1159 0 feedthrough
rlabel pdiffusion 283 -1159 283 -1159 0 cellNo=511
rlabel pdiffusion 290 -1159 290 -1159 0 feedthrough
rlabel pdiffusion 297 -1159 297 -1159 0 feedthrough
rlabel pdiffusion 304 -1159 304 -1159 0 cellNo=879
rlabel pdiffusion 311 -1159 311 -1159 0 feedthrough
rlabel pdiffusion 318 -1159 318 -1159 0 feedthrough
rlabel pdiffusion 325 -1159 325 -1159 0 feedthrough
rlabel pdiffusion 332 -1159 332 -1159 0 cellNo=592
rlabel pdiffusion 339 -1159 339 -1159 0 feedthrough
rlabel pdiffusion 346 -1159 346 -1159 0 feedthrough
rlabel pdiffusion 353 -1159 353 -1159 0 feedthrough
rlabel pdiffusion 360 -1159 360 -1159 0 feedthrough
rlabel pdiffusion 367 -1159 367 -1159 0 feedthrough
rlabel pdiffusion 374 -1159 374 -1159 0 feedthrough
rlabel pdiffusion 381 -1159 381 -1159 0 feedthrough
rlabel pdiffusion 388 -1159 388 -1159 0 feedthrough
rlabel pdiffusion 395 -1159 395 -1159 0 feedthrough
rlabel pdiffusion 402 -1159 402 -1159 0 feedthrough
rlabel pdiffusion 409 -1159 409 -1159 0 feedthrough
rlabel pdiffusion 416 -1159 416 -1159 0 cellNo=22
rlabel pdiffusion 423 -1159 423 -1159 0 feedthrough
rlabel pdiffusion 430 -1159 430 -1159 0 feedthrough
rlabel pdiffusion 437 -1159 437 -1159 0 feedthrough
rlabel pdiffusion 444 -1159 444 -1159 0 cellNo=19
rlabel pdiffusion 451 -1159 451 -1159 0 feedthrough
rlabel pdiffusion 458 -1159 458 -1159 0 feedthrough
rlabel pdiffusion 465 -1159 465 -1159 0 feedthrough
rlabel pdiffusion 472 -1159 472 -1159 0 feedthrough
rlabel pdiffusion 479 -1159 479 -1159 0 feedthrough
rlabel pdiffusion 486 -1159 486 -1159 0 feedthrough
rlabel pdiffusion 493 -1159 493 -1159 0 feedthrough
rlabel pdiffusion 500 -1159 500 -1159 0 feedthrough
rlabel pdiffusion 507 -1159 507 -1159 0 cellNo=557
rlabel pdiffusion 514 -1159 514 -1159 0 feedthrough
rlabel pdiffusion 521 -1159 521 -1159 0 feedthrough
rlabel pdiffusion 528 -1159 528 -1159 0 feedthrough
rlabel pdiffusion 535 -1159 535 -1159 0 feedthrough
rlabel pdiffusion 542 -1159 542 -1159 0 feedthrough
rlabel pdiffusion 549 -1159 549 -1159 0 cellNo=242
rlabel pdiffusion 556 -1159 556 -1159 0 feedthrough
rlabel pdiffusion 563 -1159 563 -1159 0 feedthrough
rlabel pdiffusion 570 -1159 570 -1159 0 feedthrough
rlabel pdiffusion 577 -1159 577 -1159 0 feedthrough
rlabel pdiffusion 584 -1159 584 -1159 0 cellNo=746
rlabel pdiffusion 591 -1159 591 -1159 0 feedthrough
rlabel pdiffusion 598 -1159 598 -1159 0 feedthrough
rlabel pdiffusion 605 -1159 605 -1159 0 cellNo=555
rlabel pdiffusion 612 -1159 612 -1159 0 feedthrough
rlabel pdiffusion 619 -1159 619 -1159 0 feedthrough
rlabel pdiffusion 626 -1159 626 -1159 0 cellNo=231
rlabel pdiffusion 633 -1159 633 -1159 0 feedthrough
rlabel pdiffusion 640 -1159 640 -1159 0 feedthrough
rlabel pdiffusion 647 -1159 647 -1159 0 feedthrough
rlabel pdiffusion 654 -1159 654 -1159 0 cellNo=852
rlabel pdiffusion 661 -1159 661 -1159 0 feedthrough
rlabel pdiffusion 668 -1159 668 -1159 0 cellNo=679
rlabel pdiffusion 675 -1159 675 -1159 0 feedthrough
rlabel pdiffusion 682 -1159 682 -1159 0 feedthrough
rlabel pdiffusion 689 -1159 689 -1159 0 feedthrough
rlabel pdiffusion 696 -1159 696 -1159 0 feedthrough
rlabel pdiffusion 703 -1159 703 -1159 0 feedthrough
rlabel pdiffusion 710 -1159 710 -1159 0 feedthrough
rlabel pdiffusion 717 -1159 717 -1159 0 feedthrough
rlabel pdiffusion 724 -1159 724 -1159 0 feedthrough
rlabel pdiffusion 731 -1159 731 -1159 0 feedthrough
rlabel pdiffusion 738 -1159 738 -1159 0 feedthrough
rlabel pdiffusion 745 -1159 745 -1159 0 feedthrough
rlabel pdiffusion 752 -1159 752 -1159 0 feedthrough
rlabel pdiffusion 759 -1159 759 -1159 0 feedthrough
rlabel pdiffusion 766 -1159 766 -1159 0 feedthrough
rlabel pdiffusion 773 -1159 773 -1159 0 feedthrough
rlabel pdiffusion 780 -1159 780 -1159 0 feedthrough
rlabel pdiffusion 787 -1159 787 -1159 0 feedthrough
rlabel pdiffusion 794 -1159 794 -1159 0 feedthrough
rlabel pdiffusion 801 -1159 801 -1159 0 feedthrough
rlabel pdiffusion 808 -1159 808 -1159 0 cellNo=253
rlabel pdiffusion 815 -1159 815 -1159 0 feedthrough
rlabel pdiffusion 822 -1159 822 -1159 0 feedthrough
rlabel pdiffusion 829 -1159 829 -1159 0 feedthrough
rlabel pdiffusion 836 -1159 836 -1159 0 feedthrough
rlabel pdiffusion 843 -1159 843 -1159 0 feedthrough
rlabel pdiffusion 850 -1159 850 -1159 0 cellNo=821
rlabel pdiffusion 857 -1159 857 -1159 0 feedthrough
rlabel pdiffusion 864 -1159 864 -1159 0 feedthrough
rlabel pdiffusion 871 -1159 871 -1159 0 feedthrough
rlabel pdiffusion 878 -1159 878 -1159 0 feedthrough
rlabel pdiffusion 885 -1159 885 -1159 0 feedthrough
rlabel pdiffusion 892 -1159 892 -1159 0 feedthrough
rlabel pdiffusion 899 -1159 899 -1159 0 feedthrough
rlabel pdiffusion 906 -1159 906 -1159 0 feedthrough
rlabel pdiffusion 913 -1159 913 -1159 0 feedthrough
rlabel pdiffusion 920 -1159 920 -1159 0 feedthrough
rlabel pdiffusion 927 -1159 927 -1159 0 feedthrough
rlabel pdiffusion 934 -1159 934 -1159 0 cellNo=628
rlabel pdiffusion 941 -1159 941 -1159 0 feedthrough
rlabel pdiffusion 948 -1159 948 -1159 0 feedthrough
rlabel pdiffusion 955 -1159 955 -1159 0 feedthrough
rlabel pdiffusion 962 -1159 962 -1159 0 feedthrough
rlabel pdiffusion 969 -1159 969 -1159 0 feedthrough
rlabel pdiffusion 976 -1159 976 -1159 0 cellNo=876
rlabel pdiffusion 983 -1159 983 -1159 0 feedthrough
rlabel pdiffusion 990 -1159 990 -1159 0 feedthrough
rlabel pdiffusion 997 -1159 997 -1159 0 feedthrough
rlabel pdiffusion 1004 -1159 1004 -1159 0 cellNo=631
rlabel pdiffusion 1011 -1159 1011 -1159 0 feedthrough
rlabel pdiffusion 1018 -1159 1018 -1159 0 feedthrough
rlabel pdiffusion 1025 -1159 1025 -1159 0 feedthrough
rlabel pdiffusion 1032 -1159 1032 -1159 0 feedthrough
rlabel pdiffusion 1039 -1159 1039 -1159 0 feedthrough
rlabel pdiffusion 1046 -1159 1046 -1159 0 cellNo=341
rlabel pdiffusion 1060 -1159 1060 -1159 0 feedthrough
rlabel pdiffusion 1067 -1159 1067 -1159 0 feedthrough
rlabel pdiffusion 1081 -1159 1081 -1159 0 feedthrough
rlabel pdiffusion 1088 -1159 1088 -1159 0 feedthrough
rlabel pdiffusion 1109 -1159 1109 -1159 0 feedthrough
rlabel pdiffusion 1186 -1159 1186 -1159 0 cellNo=710
rlabel pdiffusion 3 -1234 3 -1234 0 cellNo=541
rlabel pdiffusion 10 -1234 10 -1234 0 cellNo=542
rlabel pdiffusion 17 -1234 17 -1234 0 feedthrough
rlabel pdiffusion 24 -1234 24 -1234 0 cellNo=634
rlabel pdiffusion 31 -1234 31 -1234 0 feedthrough
rlabel pdiffusion 38 -1234 38 -1234 0 feedthrough
rlabel pdiffusion 45 -1234 45 -1234 0 cellNo=33
rlabel pdiffusion 52 -1234 52 -1234 0 feedthrough
rlabel pdiffusion 59 -1234 59 -1234 0 cellNo=333
rlabel pdiffusion 66 -1234 66 -1234 0 cellNo=605
rlabel pdiffusion 73 -1234 73 -1234 0 feedthrough
rlabel pdiffusion 80 -1234 80 -1234 0 feedthrough
rlabel pdiffusion 87 -1234 87 -1234 0 cellNo=670
rlabel pdiffusion 94 -1234 94 -1234 0 feedthrough
rlabel pdiffusion 101 -1234 101 -1234 0 feedthrough
rlabel pdiffusion 108 -1234 108 -1234 0 feedthrough
rlabel pdiffusion 115 -1234 115 -1234 0 cellNo=290
rlabel pdiffusion 122 -1234 122 -1234 0 feedthrough
rlabel pdiffusion 129 -1234 129 -1234 0 feedthrough
rlabel pdiffusion 136 -1234 136 -1234 0 feedthrough
rlabel pdiffusion 143 -1234 143 -1234 0 feedthrough
rlabel pdiffusion 150 -1234 150 -1234 0 cellNo=522
rlabel pdiffusion 157 -1234 157 -1234 0 feedthrough
rlabel pdiffusion 164 -1234 164 -1234 0 feedthrough
rlabel pdiffusion 171 -1234 171 -1234 0 feedthrough
rlabel pdiffusion 178 -1234 178 -1234 0 cellNo=30
rlabel pdiffusion 185 -1234 185 -1234 0 feedthrough
rlabel pdiffusion 192 -1234 192 -1234 0 feedthrough
rlabel pdiffusion 199 -1234 199 -1234 0 feedthrough
rlabel pdiffusion 206 -1234 206 -1234 0 feedthrough
rlabel pdiffusion 213 -1234 213 -1234 0 feedthrough
rlabel pdiffusion 220 -1234 220 -1234 0 feedthrough
rlabel pdiffusion 227 -1234 227 -1234 0 feedthrough
rlabel pdiffusion 234 -1234 234 -1234 0 feedthrough
rlabel pdiffusion 241 -1234 241 -1234 0 feedthrough
rlabel pdiffusion 248 -1234 248 -1234 0 feedthrough
rlabel pdiffusion 255 -1234 255 -1234 0 feedthrough
rlabel pdiffusion 262 -1234 262 -1234 0 cellNo=545
rlabel pdiffusion 269 -1234 269 -1234 0 feedthrough
rlabel pdiffusion 276 -1234 276 -1234 0 feedthrough
rlabel pdiffusion 283 -1234 283 -1234 0 feedthrough
rlabel pdiffusion 290 -1234 290 -1234 0 feedthrough
rlabel pdiffusion 297 -1234 297 -1234 0 feedthrough
rlabel pdiffusion 304 -1234 304 -1234 0 feedthrough
rlabel pdiffusion 311 -1234 311 -1234 0 feedthrough
rlabel pdiffusion 318 -1234 318 -1234 0 cellNo=427
rlabel pdiffusion 325 -1234 325 -1234 0 feedthrough
rlabel pdiffusion 332 -1234 332 -1234 0 feedthrough
rlabel pdiffusion 339 -1234 339 -1234 0 feedthrough
rlabel pdiffusion 346 -1234 346 -1234 0 feedthrough
rlabel pdiffusion 353 -1234 353 -1234 0 feedthrough
rlabel pdiffusion 360 -1234 360 -1234 0 feedthrough
rlabel pdiffusion 367 -1234 367 -1234 0 feedthrough
rlabel pdiffusion 374 -1234 374 -1234 0 cellNo=582
rlabel pdiffusion 381 -1234 381 -1234 0 cellNo=25
rlabel pdiffusion 388 -1234 388 -1234 0 cellNo=182
rlabel pdiffusion 395 -1234 395 -1234 0 feedthrough
rlabel pdiffusion 402 -1234 402 -1234 0 feedthrough
rlabel pdiffusion 409 -1234 409 -1234 0 feedthrough
rlabel pdiffusion 416 -1234 416 -1234 0 feedthrough
rlabel pdiffusion 423 -1234 423 -1234 0 cellNo=444
rlabel pdiffusion 430 -1234 430 -1234 0 feedthrough
rlabel pdiffusion 437 -1234 437 -1234 0 feedthrough
rlabel pdiffusion 444 -1234 444 -1234 0 cellNo=834
rlabel pdiffusion 451 -1234 451 -1234 0 feedthrough
rlabel pdiffusion 458 -1234 458 -1234 0 feedthrough
rlabel pdiffusion 465 -1234 465 -1234 0 feedthrough
rlabel pdiffusion 472 -1234 472 -1234 0 feedthrough
rlabel pdiffusion 479 -1234 479 -1234 0 feedthrough
rlabel pdiffusion 486 -1234 486 -1234 0 feedthrough
rlabel pdiffusion 493 -1234 493 -1234 0 feedthrough
rlabel pdiffusion 500 -1234 500 -1234 0 feedthrough
rlabel pdiffusion 507 -1234 507 -1234 0 cellNo=721
rlabel pdiffusion 514 -1234 514 -1234 0 feedthrough
rlabel pdiffusion 521 -1234 521 -1234 0 feedthrough
rlabel pdiffusion 528 -1234 528 -1234 0 feedthrough
rlabel pdiffusion 535 -1234 535 -1234 0 feedthrough
rlabel pdiffusion 542 -1234 542 -1234 0 cellNo=92
rlabel pdiffusion 549 -1234 549 -1234 0 cellNo=423
rlabel pdiffusion 556 -1234 556 -1234 0 feedthrough
rlabel pdiffusion 563 -1234 563 -1234 0 cellNo=110
rlabel pdiffusion 570 -1234 570 -1234 0 cellNo=471
rlabel pdiffusion 577 -1234 577 -1234 0 feedthrough
rlabel pdiffusion 584 -1234 584 -1234 0 feedthrough
rlabel pdiffusion 591 -1234 591 -1234 0 cellNo=112
rlabel pdiffusion 598 -1234 598 -1234 0 feedthrough
rlabel pdiffusion 605 -1234 605 -1234 0 feedthrough
rlabel pdiffusion 612 -1234 612 -1234 0 feedthrough
rlabel pdiffusion 619 -1234 619 -1234 0 feedthrough
rlabel pdiffusion 626 -1234 626 -1234 0 feedthrough
rlabel pdiffusion 633 -1234 633 -1234 0 feedthrough
rlabel pdiffusion 640 -1234 640 -1234 0 cellNo=375
rlabel pdiffusion 647 -1234 647 -1234 0 feedthrough
rlabel pdiffusion 654 -1234 654 -1234 0 cellNo=618
rlabel pdiffusion 661 -1234 661 -1234 0 cellNo=641
rlabel pdiffusion 668 -1234 668 -1234 0 feedthrough
rlabel pdiffusion 675 -1234 675 -1234 0 feedthrough
rlabel pdiffusion 682 -1234 682 -1234 0 feedthrough
rlabel pdiffusion 689 -1234 689 -1234 0 feedthrough
rlabel pdiffusion 696 -1234 696 -1234 0 feedthrough
rlabel pdiffusion 703 -1234 703 -1234 0 feedthrough
rlabel pdiffusion 710 -1234 710 -1234 0 cellNo=463
rlabel pdiffusion 717 -1234 717 -1234 0 feedthrough
rlabel pdiffusion 724 -1234 724 -1234 0 cellNo=173
rlabel pdiffusion 731 -1234 731 -1234 0 feedthrough
rlabel pdiffusion 738 -1234 738 -1234 0 feedthrough
rlabel pdiffusion 745 -1234 745 -1234 0 feedthrough
rlabel pdiffusion 752 -1234 752 -1234 0 feedthrough
rlabel pdiffusion 759 -1234 759 -1234 0 feedthrough
rlabel pdiffusion 766 -1234 766 -1234 0 feedthrough
rlabel pdiffusion 773 -1234 773 -1234 0 cellNo=446
rlabel pdiffusion 780 -1234 780 -1234 0 feedthrough
rlabel pdiffusion 787 -1234 787 -1234 0 feedthrough
rlabel pdiffusion 794 -1234 794 -1234 0 feedthrough
rlabel pdiffusion 801 -1234 801 -1234 0 feedthrough
rlabel pdiffusion 808 -1234 808 -1234 0 feedthrough
rlabel pdiffusion 815 -1234 815 -1234 0 feedthrough
rlabel pdiffusion 822 -1234 822 -1234 0 feedthrough
rlabel pdiffusion 829 -1234 829 -1234 0 cellNo=111
rlabel pdiffusion 836 -1234 836 -1234 0 feedthrough
rlabel pdiffusion 843 -1234 843 -1234 0 feedthrough
rlabel pdiffusion 850 -1234 850 -1234 0 feedthrough
rlabel pdiffusion 857 -1234 857 -1234 0 feedthrough
rlabel pdiffusion 864 -1234 864 -1234 0 feedthrough
rlabel pdiffusion 871 -1234 871 -1234 0 feedthrough
rlabel pdiffusion 878 -1234 878 -1234 0 feedthrough
rlabel pdiffusion 885 -1234 885 -1234 0 feedthrough
rlabel pdiffusion 892 -1234 892 -1234 0 feedthrough
rlabel pdiffusion 899 -1234 899 -1234 0 feedthrough
rlabel pdiffusion 906 -1234 906 -1234 0 feedthrough
rlabel pdiffusion 913 -1234 913 -1234 0 feedthrough
rlabel pdiffusion 920 -1234 920 -1234 0 feedthrough
rlabel pdiffusion 927 -1234 927 -1234 0 feedthrough
rlabel pdiffusion 934 -1234 934 -1234 0 feedthrough
rlabel pdiffusion 941 -1234 941 -1234 0 feedthrough
rlabel pdiffusion 948 -1234 948 -1234 0 feedthrough
rlabel pdiffusion 955 -1234 955 -1234 0 feedthrough
rlabel pdiffusion 962 -1234 962 -1234 0 feedthrough
rlabel pdiffusion 969 -1234 969 -1234 0 feedthrough
rlabel pdiffusion 976 -1234 976 -1234 0 feedthrough
rlabel pdiffusion 983 -1234 983 -1234 0 feedthrough
rlabel pdiffusion 990 -1234 990 -1234 0 feedthrough
rlabel pdiffusion 997 -1234 997 -1234 0 feedthrough
rlabel pdiffusion 1004 -1234 1004 -1234 0 feedthrough
rlabel pdiffusion 1011 -1234 1011 -1234 0 feedthrough
rlabel pdiffusion 1018 -1234 1018 -1234 0 feedthrough
rlabel pdiffusion 1025 -1234 1025 -1234 0 feedthrough
rlabel pdiffusion 1032 -1234 1032 -1234 0 feedthrough
rlabel pdiffusion 1039 -1234 1039 -1234 0 feedthrough
rlabel pdiffusion 1046 -1234 1046 -1234 0 feedthrough
rlabel pdiffusion 1053 -1234 1053 -1234 0 feedthrough
rlabel pdiffusion 1060 -1234 1060 -1234 0 feedthrough
rlabel pdiffusion 1067 -1234 1067 -1234 0 feedthrough
rlabel pdiffusion 1074 -1234 1074 -1234 0 feedthrough
rlabel pdiffusion 1081 -1234 1081 -1234 0 feedthrough
rlabel pdiffusion 1088 -1234 1088 -1234 0 feedthrough
rlabel pdiffusion 1095 -1234 1095 -1234 0 feedthrough
rlabel pdiffusion 1102 -1234 1102 -1234 0 feedthrough
rlabel pdiffusion 1109 -1234 1109 -1234 0 feedthrough
rlabel pdiffusion 1116 -1234 1116 -1234 0 feedthrough
rlabel pdiffusion 1123 -1234 1123 -1234 0 feedthrough
rlabel pdiffusion 1130 -1234 1130 -1234 0 feedthrough
rlabel pdiffusion 3 -1305 3 -1305 0 cellNo=28
rlabel pdiffusion 10 -1305 10 -1305 0 cellNo=657
rlabel pdiffusion 17 -1305 17 -1305 0 cellNo=354
rlabel pdiffusion 45 -1305 45 -1305 0 feedthrough
rlabel pdiffusion 73 -1305 73 -1305 0 feedthrough
rlabel pdiffusion 80 -1305 80 -1305 0 feedthrough
rlabel pdiffusion 87 -1305 87 -1305 0 feedthrough
rlabel pdiffusion 94 -1305 94 -1305 0 cellNo=379
rlabel pdiffusion 101 -1305 101 -1305 0 feedthrough
rlabel pdiffusion 108 -1305 108 -1305 0 feedthrough
rlabel pdiffusion 115 -1305 115 -1305 0 feedthrough
rlabel pdiffusion 122 -1305 122 -1305 0 feedthrough
rlabel pdiffusion 129 -1305 129 -1305 0 feedthrough
rlabel pdiffusion 136 -1305 136 -1305 0 feedthrough
rlabel pdiffusion 143 -1305 143 -1305 0 feedthrough
rlabel pdiffusion 150 -1305 150 -1305 0 cellNo=486
rlabel pdiffusion 157 -1305 157 -1305 0 feedthrough
rlabel pdiffusion 164 -1305 164 -1305 0 feedthrough
rlabel pdiffusion 171 -1305 171 -1305 0 feedthrough
rlabel pdiffusion 178 -1305 178 -1305 0 feedthrough
rlabel pdiffusion 185 -1305 185 -1305 0 feedthrough
rlabel pdiffusion 192 -1305 192 -1305 0 cellNo=294
rlabel pdiffusion 199 -1305 199 -1305 0 feedthrough
rlabel pdiffusion 206 -1305 206 -1305 0 feedthrough
rlabel pdiffusion 213 -1305 213 -1305 0 feedthrough
rlabel pdiffusion 220 -1305 220 -1305 0 feedthrough
rlabel pdiffusion 227 -1305 227 -1305 0 feedthrough
rlabel pdiffusion 234 -1305 234 -1305 0 feedthrough
rlabel pdiffusion 241 -1305 241 -1305 0 cellNo=611
rlabel pdiffusion 248 -1305 248 -1305 0 feedthrough
rlabel pdiffusion 255 -1305 255 -1305 0 feedthrough
rlabel pdiffusion 262 -1305 262 -1305 0 feedthrough
rlabel pdiffusion 269 -1305 269 -1305 0 feedthrough
rlabel pdiffusion 276 -1305 276 -1305 0 feedthrough
rlabel pdiffusion 283 -1305 283 -1305 0 feedthrough
rlabel pdiffusion 290 -1305 290 -1305 0 feedthrough
rlabel pdiffusion 297 -1305 297 -1305 0 feedthrough
rlabel pdiffusion 304 -1305 304 -1305 0 cellNo=506
rlabel pdiffusion 311 -1305 311 -1305 0 feedthrough
rlabel pdiffusion 318 -1305 318 -1305 0 feedthrough
rlabel pdiffusion 325 -1305 325 -1305 0 feedthrough
rlabel pdiffusion 332 -1305 332 -1305 0 feedthrough
rlabel pdiffusion 339 -1305 339 -1305 0 cellNo=563
rlabel pdiffusion 346 -1305 346 -1305 0 feedthrough
rlabel pdiffusion 353 -1305 353 -1305 0 feedthrough
rlabel pdiffusion 360 -1305 360 -1305 0 feedthrough
rlabel pdiffusion 367 -1305 367 -1305 0 feedthrough
rlabel pdiffusion 374 -1305 374 -1305 0 feedthrough
rlabel pdiffusion 381 -1305 381 -1305 0 feedthrough
rlabel pdiffusion 388 -1305 388 -1305 0 feedthrough
rlabel pdiffusion 395 -1305 395 -1305 0 feedthrough
rlabel pdiffusion 402 -1305 402 -1305 0 cellNo=165
rlabel pdiffusion 409 -1305 409 -1305 0 feedthrough
rlabel pdiffusion 416 -1305 416 -1305 0 feedthrough
rlabel pdiffusion 423 -1305 423 -1305 0 feedthrough
rlabel pdiffusion 430 -1305 430 -1305 0 feedthrough
rlabel pdiffusion 437 -1305 437 -1305 0 feedthrough
rlabel pdiffusion 444 -1305 444 -1305 0 feedthrough
rlabel pdiffusion 451 -1305 451 -1305 0 feedthrough
rlabel pdiffusion 458 -1305 458 -1305 0 feedthrough
rlabel pdiffusion 465 -1305 465 -1305 0 cellNo=445
rlabel pdiffusion 472 -1305 472 -1305 0 feedthrough
rlabel pdiffusion 479 -1305 479 -1305 0 cellNo=95
rlabel pdiffusion 486 -1305 486 -1305 0 feedthrough
rlabel pdiffusion 493 -1305 493 -1305 0 feedthrough
rlabel pdiffusion 500 -1305 500 -1305 0 cellNo=442
rlabel pdiffusion 507 -1305 507 -1305 0 feedthrough
rlabel pdiffusion 514 -1305 514 -1305 0 feedthrough
rlabel pdiffusion 521 -1305 521 -1305 0 feedthrough
rlabel pdiffusion 528 -1305 528 -1305 0 feedthrough
rlabel pdiffusion 535 -1305 535 -1305 0 cellNo=151
rlabel pdiffusion 542 -1305 542 -1305 0 feedthrough
rlabel pdiffusion 549 -1305 549 -1305 0 feedthrough
rlabel pdiffusion 556 -1305 556 -1305 0 feedthrough
rlabel pdiffusion 563 -1305 563 -1305 0 feedthrough
rlabel pdiffusion 570 -1305 570 -1305 0 cellNo=686
rlabel pdiffusion 577 -1305 577 -1305 0 cellNo=781
rlabel pdiffusion 584 -1305 584 -1305 0 feedthrough
rlabel pdiffusion 591 -1305 591 -1305 0 feedthrough
rlabel pdiffusion 598 -1305 598 -1305 0 cellNo=104
rlabel pdiffusion 605 -1305 605 -1305 0 feedthrough
rlabel pdiffusion 612 -1305 612 -1305 0 cellNo=799
rlabel pdiffusion 619 -1305 619 -1305 0 feedthrough
rlabel pdiffusion 626 -1305 626 -1305 0 feedthrough
rlabel pdiffusion 633 -1305 633 -1305 0 cellNo=569
rlabel pdiffusion 640 -1305 640 -1305 0 feedthrough
rlabel pdiffusion 647 -1305 647 -1305 0 feedthrough
rlabel pdiffusion 654 -1305 654 -1305 0 cellNo=578
rlabel pdiffusion 661 -1305 661 -1305 0 feedthrough
rlabel pdiffusion 668 -1305 668 -1305 0 feedthrough
rlabel pdiffusion 675 -1305 675 -1305 0 cellNo=610
rlabel pdiffusion 682 -1305 682 -1305 0 feedthrough
rlabel pdiffusion 689 -1305 689 -1305 0 feedthrough
rlabel pdiffusion 696 -1305 696 -1305 0 feedthrough
rlabel pdiffusion 703 -1305 703 -1305 0 feedthrough
rlabel pdiffusion 710 -1305 710 -1305 0 feedthrough
rlabel pdiffusion 717 -1305 717 -1305 0 feedthrough
rlabel pdiffusion 724 -1305 724 -1305 0 feedthrough
rlabel pdiffusion 731 -1305 731 -1305 0 feedthrough
rlabel pdiffusion 738 -1305 738 -1305 0 feedthrough
rlabel pdiffusion 745 -1305 745 -1305 0 feedthrough
rlabel pdiffusion 752 -1305 752 -1305 0 feedthrough
rlabel pdiffusion 759 -1305 759 -1305 0 feedthrough
rlabel pdiffusion 766 -1305 766 -1305 0 feedthrough
rlabel pdiffusion 773 -1305 773 -1305 0 feedthrough
rlabel pdiffusion 780 -1305 780 -1305 0 feedthrough
rlabel pdiffusion 787 -1305 787 -1305 0 feedthrough
rlabel pdiffusion 794 -1305 794 -1305 0 cellNo=815
rlabel pdiffusion 801 -1305 801 -1305 0 feedthrough
rlabel pdiffusion 808 -1305 808 -1305 0 feedthrough
rlabel pdiffusion 815 -1305 815 -1305 0 feedthrough
rlabel pdiffusion 822 -1305 822 -1305 0 feedthrough
rlabel pdiffusion 829 -1305 829 -1305 0 feedthrough
rlabel pdiffusion 836 -1305 836 -1305 0 feedthrough
rlabel pdiffusion 843 -1305 843 -1305 0 feedthrough
rlabel pdiffusion 850 -1305 850 -1305 0 feedthrough
rlabel pdiffusion 857 -1305 857 -1305 0 feedthrough
rlabel pdiffusion 864 -1305 864 -1305 0 cellNo=197
rlabel pdiffusion 871 -1305 871 -1305 0 feedthrough
rlabel pdiffusion 878 -1305 878 -1305 0 feedthrough
rlabel pdiffusion 885 -1305 885 -1305 0 feedthrough
rlabel pdiffusion 892 -1305 892 -1305 0 feedthrough
rlabel pdiffusion 899 -1305 899 -1305 0 feedthrough
rlabel pdiffusion 906 -1305 906 -1305 0 feedthrough
rlabel pdiffusion 913 -1305 913 -1305 0 feedthrough
rlabel pdiffusion 920 -1305 920 -1305 0 cellNo=785
rlabel pdiffusion 927 -1305 927 -1305 0 feedthrough
rlabel pdiffusion 934 -1305 934 -1305 0 feedthrough
rlabel pdiffusion 941 -1305 941 -1305 0 feedthrough
rlabel pdiffusion 948 -1305 948 -1305 0 feedthrough
rlabel pdiffusion 955 -1305 955 -1305 0 feedthrough
rlabel pdiffusion 962 -1305 962 -1305 0 feedthrough
rlabel pdiffusion 969 -1305 969 -1305 0 feedthrough
rlabel pdiffusion 976 -1305 976 -1305 0 cellNo=334
rlabel pdiffusion 983 -1305 983 -1305 0 feedthrough
rlabel pdiffusion 990 -1305 990 -1305 0 feedthrough
rlabel pdiffusion 997 -1305 997 -1305 0 cellNo=312
rlabel pdiffusion 1004 -1305 1004 -1305 0 feedthrough
rlabel pdiffusion 1011 -1305 1011 -1305 0 feedthrough
rlabel pdiffusion 1018 -1305 1018 -1305 0 cellNo=385
rlabel pdiffusion 1025 -1305 1025 -1305 0 cellNo=141
rlabel pdiffusion 1032 -1305 1032 -1305 0 feedthrough
rlabel pdiffusion 1039 -1305 1039 -1305 0 feedthrough
rlabel pdiffusion 1046 -1305 1046 -1305 0 feedthrough
rlabel pdiffusion 1053 -1305 1053 -1305 0 feedthrough
rlabel pdiffusion 1060 -1305 1060 -1305 0 cellNo=716
rlabel pdiffusion 1067 -1305 1067 -1305 0 feedthrough
rlabel pdiffusion 1081 -1305 1081 -1305 0 feedthrough
rlabel pdiffusion 1088 -1305 1088 -1305 0 feedthrough
rlabel pdiffusion 1095 -1305 1095 -1305 0 cellNo=144
rlabel pdiffusion 1102 -1305 1102 -1305 0 feedthrough
rlabel pdiffusion 3 -1376 3 -1376 0 cellNo=512
rlabel pdiffusion 10 -1376 10 -1376 0 cellNo=771
rlabel pdiffusion 17 -1376 17 -1376 0 feedthrough
rlabel pdiffusion 24 -1376 24 -1376 0 feedthrough
rlabel pdiffusion 31 -1376 31 -1376 0 feedthrough
rlabel pdiffusion 38 -1376 38 -1376 0 feedthrough
rlabel pdiffusion 45 -1376 45 -1376 0 feedthrough
rlabel pdiffusion 52 -1376 52 -1376 0 feedthrough
rlabel pdiffusion 59 -1376 59 -1376 0 feedthrough
rlabel pdiffusion 66 -1376 66 -1376 0 cellNo=389
rlabel pdiffusion 73 -1376 73 -1376 0 feedthrough
rlabel pdiffusion 80 -1376 80 -1376 0 feedthrough
rlabel pdiffusion 87 -1376 87 -1376 0 feedthrough
rlabel pdiffusion 94 -1376 94 -1376 0 cellNo=232
rlabel pdiffusion 101 -1376 101 -1376 0 cellNo=792
rlabel pdiffusion 108 -1376 108 -1376 0 feedthrough
rlabel pdiffusion 115 -1376 115 -1376 0 feedthrough
rlabel pdiffusion 122 -1376 122 -1376 0 feedthrough
rlabel pdiffusion 129 -1376 129 -1376 0 feedthrough
rlabel pdiffusion 136 -1376 136 -1376 0 cellNo=425
rlabel pdiffusion 143 -1376 143 -1376 0 cellNo=507
rlabel pdiffusion 150 -1376 150 -1376 0 feedthrough
rlabel pdiffusion 157 -1376 157 -1376 0 feedthrough
rlabel pdiffusion 164 -1376 164 -1376 0 feedthrough
rlabel pdiffusion 171 -1376 171 -1376 0 feedthrough
rlabel pdiffusion 178 -1376 178 -1376 0 cellNo=132
rlabel pdiffusion 185 -1376 185 -1376 0 feedthrough
rlabel pdiffusion 192 -1376 192 -1376 0 feedthrough
rlabel pdiffusion 199 -1376 199 -1376 0 cellNo=767
rlabel pdiffusion 206 -1376 206 -1376 0 feedthrough
rlabel pdiffusion 213 -1376 213 -1376 0 feedthrough
rlabel pdiffusion 220 -1376 220 -1376 0 feedthrough
rlabel pdiffusion 227 -1376 227 -1376 0 feedthrough
rlabel pdiffusion 234 -1376 234 -1376 0 cellNo=737
rlabel pdiffusion 241 -1376 241 -1376 0 feedthrough
rlabel pdiffusion 248 -1376 248 -1376 0 cellNo=617
rlabel pdiffusion 255 -1376 255 -1376 0 feedthrough
rlabel pdiffusion 262 -1376 262 -1376 0 feedthrough
rlabel pdiffusion 269 -1376 269 -1376 0 feedthrough
rlabel pdiffusion 276 -1376 276 -1376 0 cellNo=498
rlabel pdiffusion 283 -1376 283 -1376 0 cellNo=315
rlabel pdiffusion 290 -1376 290 -1376 0 feedthrough
rlabel pdiffusion 297 -1376 297 -1376 0 feedthrough
rlabel pdiffusion 304 -1376 304 -1376 0 feedthrough
rlabel pdiffusion 311 -1376 311 -1376 0 feedthrough
rlabel pdiffusion 318 -1376 318 -1376 0 feedthrough
rlabel pdiffusion 325 -1376 325 -1376 0 feedthrough
rlabel pdiffusion 332 -1376 332 -1376 0 feedthrough
rlabel pdiffusion 339 -1376 339 -1376 0 feedthrough
rlabel pdiffusion 346 -1376 346 -1376 0 cellNo=113
rlabel pdiffusion 353 -1376 353 -1376 0 feedthrough
rlabel pdiffusion 360 -1376 360 -1376 0 feedthrough
rlabel pdiffusion 367 -1376 367 -1376 0 cellNo=411
rlabel pdiffusion 374 -1376 374 -1376 0 feedthrough
rlabel pdiffusion 381 -1376 381 -1376 0 feedthrough
rlabel pdiffusion 388 -1376 388 -1376 0 feedthrough
rlabel pdiffusion 395 -1376 395 -1376 0 feedthrough
rlabel pdiffusion 402 -1376 402 -1376 0 feedthrough
rlabel pdiffusion 409 -1376 409 -1376 0 cellNo=598
rlabel pdiffusion 416 -1376 416 -1376 0 feedthrough
rlabel pdiffusion 423 -1376 423 -1376 0 feedthrough
rlabel pdiffusion 430 -1376 430 -1376 0 feedthrough
rlabel pdiffusion 437 -1376 437 -1376 0 cellNo=530
rlabel pdiffusion 444 -1376 444 -1376 0 feedthrough
rlabel pdiffusion 451 -1376 451 -1376 0 feedthrough
rlabel pdiffusion 458 -1376 458 -1376 0 feedthrough
rlabel pdiffusion 465 -1376 465 -1376 0 feedthrough
rlabel pdiffusion 472 -1376 472 -1376 0 feedthrough
rlabel pdiffusion 479 -1376 479 -1376 0 cellNo=164
rlabel pdiffusion 486 -1376 486 -1376 0 feedthrough
rlabel pdiffusion 493 -1376 493 -1376 0 cellNo=558
rlabel pdiffusion 500 -1376 500 -1376 0 feedthrough
rlabel pdiffusion 507 -1376 507 -1376 0 cellNo=843
rlabel pdiffusion 514 -1376 514 -1376 0 feedthrough
rlabel pdiffusion 521 -1376 521 -1376 0 feedthrough
rlabel pdiffusion 528 -1376 528 -1376 0 feedthrough
rlabel pdiffusion 535 -1376 535 -1376 0 feedthrough
rlabel pdiffusion 542 -1376 542 -1376 0 cellNo=361
rlabel pdiffusion 549 -1376 549 -1376 0 feedthrough
rlabel pdiffusion 556 -1376 556 -1376 0 feedthrough
rlabel pdiffusion 563 -1376 563 -1376 0 feedthrough
rlabel pdiffusion 570 -1376 570 -1376 0 cellNo=185
rlabel pdiffusion 577 -1376 577 -1376 0 feedthrough
rlabel pdiffusion 584 -1376 584 -1376 0 feedthrough
rlabel pdiffusion 591 -1376 591 -1376 0 feedthrough
rlabel pdiffusion 598 -1376 598 -1376 0 feedthrough
rlabel pdiffusion 605 -1376 605 -1376 0 feedthrough
rlabel pdiffusion 612 -1376 612 -1376 0 feedthrough
rlabel pdiffusion 619 -1376 619 -1376 0 feedthrough
rlabel pdiffusion 626 -1376 626 -1376 0 cellNo=272
rlabel pdiffusion 633 -1376 633 -1376 0 feedthrough
rlabel pdiffusion 640 -1376 640 -1376 0 feedthrough
rlabel pdiffusion 647 -1376 647 -1376 0 cellNo=495
rlabel pdiffusion 654 -1376 654 -1376 0 cellNo=186
rlabel pdiffusion 661 -1376 661 -1376 0 cellNo=58
rlabel pdiffusion 668 -1376 668 -1376 0 feedthrough
rlabel pdiffusion 675 -1376 675 -1376 0 feedthrough
rlabel pdiffusion 682 -1376 682 -1376 0 feedthrough
rlabel pdiffusion 689 -1376 689 -1376 0 feedthrough
rlabel pdiffusion 696 -1376 696 -1376 0 feedthrough
rlabel pdiffusion 703 -1376 703 -1376 0 feedthrough
rlabel pdiffusion 710 -1376 710 -1376 0 feedthrough
rlabel pdiffusion 717 -1376 717 -1376 0 feedthrough
rlabel pdiffusion 724 -1376 724 -1376 0 cellNo=532
rlabel pdiffusion 731 -1376 731 -1376 0 cellNo=48
rlabel pdiffusion 738 -1376 738 -1376 0 feedthrough
rlabel pdiffusion 745 -1376 745 -1376 0 feedthrough
rlabel pdiffusion 752 -1376 752 -1376 0 feedthrough
rlabel pdiffusion 759 -1376 759 -1376 0 feedthrough
rlabel pdiffusion 766 -1376 766 -1376 0 feedthrough
rlabel pdiffusion 773 -1376 773 -1376 0 feedthrough
rlabel pdiffusion 780 -1376 780 -1376 0 feedthrough
rlabel pdiffusion 787 -1376 787 -1376 0 feedthrough
rlabel pdiffusion 794 -1376 794 -1376 0 feedthrough
rlabel pdiffusion 801 -1376 801 -1376 0 feedthrough
rlabel pdiffusion 808 -1376 808 -1376 0 feedthrough
rlabel pdiffusion 815 -1376 815 -1376 0 feedthrough
rlabel pdiffusion 822 -1376 822 -1376 0 feedthrough
rlabel pdiffusion 829 -1376 829 -1376 0 feedthrough
rlabel pdiffusion 836 -1376 836 -1376 0 feedthrough
rlabel pdiffusion 843 -1376 843 -1376 0 feedthrough
rlabel pdiffusion 850 -1376 850 -1376 0 feedthrough
rlabel pdiffusion 857 -1376 857 -1376 0 feedthrough
rlabel pdiffusion 864 -1376 864 -1376 0 feedthrough
rlabel pdiffusion 871 -1376 871 -1376 0 feedthrough
rlabel pdiffusion 878 -1376 878 -1376 0 feedthrough
rlabel pdiffusion 885 -1376 885 -1376 0 feedthrough
rlabel pdiffusion 892 -1376 892 -1376 0 feedthrough
rlabel pdiffusion 899 -1376 899 -1376 0 feedthrough
rlabel pdiffusion 906 -1376 906 -1376 0 feedthrough
rlabel pdiffusion 913 -1376 913 -1376 0 feedthrough
rlabel pdiffusion 920 -1376 920 -1376 0 feedthrough
rlabel pdiffusion 927 -1376 927 -1376 0 feedthrough
rlabel pdiffusion 934 -1376 934 -1376 0 feedthrough
rlabel pdiffusion 941 -1376 941 -1376 0 feedthrough
rlabel pdiffusion 948 -1376 948 -1376 0 feedthrough
rlabel pdiffusion 955 -1376 955 -1376 0 feedthrough
rlabel pdiffusion 962 -1376 962 -1376 0 feedthrough
rlabel pdiffusion 969 -1376 969 -1376 0 feedthrough
rlabel pdiffusion 976 -1376 976 -1376 0 feedthrough
rlabel pdiffusion 983 -1376 983 -1376 0 feedthrough
rlabel pdiffusion 990 -1376 990 -1376 0 feedthrough
rlabel pdiffusion 997 -1376 997 -1376 0 cellNo=630
rlabel pdiffusion 1004 -1376 1004 -1376 0 feedthrough
rlabel pdiffusion 1011 -1376 1011 -1376 0 feedthrough
rlabel pdiffusion 1018 -1376 1018 -1376 0 feedthrough
rlabel pdiffusion 1025 -1376 1025 -1376 0 cellNo=521
rlabel pdiffusion 1032 -1376 1032 -1376 0 feedthrough
rlabel pdiffusion 1067 -1376 1067 -1376 0 feedthrough
rlabel pdiffusion 3 -1451 3 -1451 0 cellNo=797
rlabel pdiffusion 10 -1451 10 -1451 0 feedthrough
rlabel pdiffusion 17 -1451 17 -1451 0 cellNo=380
rlabel pdiffusion 24 -1451 24 -1451 0 feedthrough
rlabel pdiffusion 31 -1451 31 -1451 0 feedthrough
rlabel pdiffusion 38 -1451 38 -1451 0 cellNo=259
rlabel pdiffusion 45 -1451 45 -1451 0 feedthrough
rlabel pdiffusion 52 -1451 52 -1451 0 feedthrough
rlabel pdiffusion 59 -1451 59 -1451 0 feedthrough
rlabel pdiffusion 66 -1451 66 -1451 0 cellNo=684
rlabel pdiffusion 73 -1451 73 -1451 0 feedthrough
rlabel pdiffusion 80 -1451 80 -1451 0 feedthrough
rlabel pdiffusion 87 -1451 87 -1451 0 feedthrough
rlabel pdiffusion 94 -1451 94 -1451 0 feedthrough
rlabel pdiffusion 101 -1451 101 -1451 0 feedthrough
rlabel pdiffusion 108 -1451 108 -1451 0 feedthrough
rlabel pdiffusion 115 -1451 115 -1451 0 feedthrough
rlabel pdiffusion 122 -1451 122 -1451 0 feedthrough
rlabel pdiffusion 129 -1451 129 -1451 0 cellNo=236
rlabel pdiffusion 136 -1451 136 -1451 0 cellNo=154
rlabel pdiffusion 143 -1451 143 -1451 0 feedthrough
rlabel pdiffusion 150 -1451 150 -1451 0 feedthrough
rlabel pdiffusion 157 -1451 157 -1451 0 feedthrough
rlabel pdiffusion 164 -1451 164 -1451 0 feedthrough
rlabel pdiffusion 171 -1451 171 -1451 0 feedthrough
rlabel pdiffusion 178 -1451 178 -1451 0 feedthrough
rlabel pdiffusion 185 -1451 185 -1451 0 feedthrough
rlabel pdiffusion 192 -1451 192 -1451 0 cellNo=54
rlabel pdiffusion 199 -1451 199 -1451 0 feedthrough
rlabel pdiffusion 206 -1451 206 -1451 0 cellNo=585
rlabel pdiffusion 213 -1451 213 -1451 0 cellNo=660
rlabel pdiffusion 220 -1451 220 -1451 0 feedthrough
rlabel pdiffusion 227 -1451 227 -1451 0 feedthrough
rlabel pdiffusion 234 -1451 234 -1451 0 feedthrough
rlabel pdiffusion 241 -1451 241 -1451 0 feedthrough
rlabel pdiffusion 248 -1451 248 -1451 0 feedthrough
rlabel pdiffusion 255 -1451 255 -1451 0 feedthrough
rlabel pdiffusion 262 -1451 262 -1451 0 feedthrough
rlabel pdiffusion 269 -1451 269 -1451 0 feedthrough
rlabel pdiffusion 276 -1451 276 -1451 0 cellNo=172
rlabel pdiffusion 283 -1451 283 -1451 0 cellNo=509
rlabel pdiffusion 290 -1451 290 -1451 0 feedthrough
rlabel pdiffusion 297 -1451 297 -1451 0 feedthrough
rlabel pdiffusion 304 -1451 304 -1451 0 feedthrough
rlabel pdiffusion 311 -1451 311 -1451 0 feedthrough
rlabel pdiffusion 318 -1451 318 -1451 0 cellNo=470
rlabel pdiffusion 325 -1451 325 -1451 0 feedthrough
rlabel pdiffusion 332 -1451 332 -1451 0 feedthrough
rlabel pdiffusion 339 -1451 339 -1451 0 feedthrough
rlabel pdiffusion 346 -1451 346 -1451 0 feedthrough
rlabel pdiffusion 353 -1451 353 -1451 0 feedthrough
rlabel pdiffusion 360 -1451 360 -1451 0 feedthrough
rlabel pdiffusion 367 -1451 367 -1451 0 cellNo=370
rlabel pdiffusion 374 -1451 374 -1451 0 cellNo=210
rlabel pdiffusion 381 -1451 381 -1451 0 feedthrough
rlabel pdiffusion 388 -1451 388 -1451 0 feedthrough
rlabel pdiffusion 395 -1451 395 -1451 0 feedthrough
rlabel pdiffusion 402 -1451 402 -1451 0 feedthrough
rlabel pdiffusion 409 -1451 409 -1451 0 feedthrough
rlabel pdiffusion 416 -1451 416 -1451 0 feedthrough
rlabel pdiffusion 423 -1451 423 -1451 0 cellNo=632
rlabel pdiffusion 430 -1451 430 -1451 0 feedthrough
rlabel pdiffusion 437 -1451 437 -1451 0 cellNo=500
rlabel pdiffusion 444 -1451 444 -1451 0 feedthrough
rlabel pdiffusion 451 -1451 451 -1451 0 feedthrough
rlabel pdiffusion 458 -1451 458 -1451 0 cellNo=873
rlabel pdiffusion 465 -1451 465 -1451 0 feedthrough
rlabel pdiffusion 472 -1451 472 -1451 0 cellNo=589
rlabel pdiffusion 479 -1451 479 -1451 0 feedthrough
rlabel pdiffusion 486 -1451 486 -1451 0 cellNo=627
rlabel pdiffusion 493 -1451 493 -1451 0 feedthrough
rlabel pdiffusion 500 -1451 500 -1451 0 feedthrough
rlabel pdiffusion 507 -1451 507 -1451 0 feedthrough
rlabel pdiffusion 514 -1451 514 -1451 0 feedthrough
rlabel pdiffusion 521 -1451 521 -1451 0 cellNo=184
rlabel pdiffusion 528 -1451 528 -1451 0 cellNo=614
rlabel pdiffusion 535 -1451 535 -1451 0 cellNo=260
rlabel pdiffusion 542 -1451 542 -1451 0 feedthrough
rlabel pdiffusion 549 -1451 549 -1451 0 feedthrough
rlabel pdiffusion 556 -1451 556 -1451 0 feedthrough
rlabel pdiffusion 563 -1451 563 -1451 0 feedthrough
rlabel pdiffusion 570 -1451 570 -1451 0 feedthrough
rlabel pdiffusion 577 -1451 577 -1451 0 feedthrough
rlabel pdiffusion 584 -1451 584 -1451 0 feedthrough
rlabel pdiffusion 591 -1451 591 -1451 0 feedthrough
rlabel pdiffusion 598 -1451 598 -1451 0 feedthrough
rlabel pdiffusion 605 -1451 605 -1451 0 cellNo=217
rlabel pdiffusion 612 -1451 612 -1451 0 feedthrough
rlabel pdiffusion 619 -1451 619 -1451 0 feedthrough
rlabel pdiffusion 626 -1451 626 -1451 0 feedthrough
rlabel pdiffusion 633 -1451 633 -1451 0 cellNo=659
rlabel pdiffusion 640 -1451 640 -1451 0 cellNo=846
rlabel pdiffusion 647 -1451 647 -1451 0 feedthrough
rlabel pdiffusion 654 -1451 654 -1451 0 feedthrough
rlabel pdiffusion 661 -1451 661 -1451 0 feedthrough
rlabel pdiffusion 668 -1451 668 -1451 0 feedthrough
rlabel pdiffusion 675 -1451 675 -1451 0 feedthrough
rlabel pdiffusion 682 -1451 682 -1451 0 feedthrough
rlabel pdiffusion 689 -1451 689 -1451 0 feedthrough
rlabel pdiffusion 696 -1451 696 -1451 0 feedthrough
rlabel pdiffusion 703 -1451 703 -1451 0 feedthrough
rlabel pdiffusion 710 -1451 710 -1451 0 feedthrough
rlabel pdiffusion 717 -1451 717 -1451 0 feedthrough
rlabel pdiffusion 724 -1451 724 -1451 0 feedthrough
rlabel pdiffusion 731 -1451 731 -1451 0 feedthrough
rlabel pdiffusion 738 -1451 738 -1451 0 feedthrough
rlabel pdiffusion 745 -1451 745 -1451 0 feedthrough
rlabel pdiffusion 752 -1451 752 -1451 0 feedthrough
rlabel pdiffusion 759 -1451 759 -1451 0 feedthrough
rlabel pdiffusion 766 -1451 766 -1451 0 cellNo=633
rlabel pdiffusion 773 -1451 773 -1451 0 feedthrough
rlabel pdiffusion 780 -1451 780 -1451 0 feedthrough
rlabel pdiffusion 787 -1451 787 -1451 0 feedthrough
rlabel pdiffusion 794 -1451 794 -1451 0 cellNo=67
rlabel pdiffusion 801 -1451 801 -1451 0 feedthrough
rlabel pdiffusion 808 -1451 808 -1451 0 feedthrough
rlabel pdiffusion 815 -1451 815 -1451 0 feedthrough
rlabel pdiffusion 822 -1451 822 -1451 0 cellNo=402
rlabel pdiffusion 829 -1451 829 -1451 0 feedthrough
rlabel pdiffusion 836 -1451 836 -1451 0 feedthrough
rlabel pdiffusion 843 -1451 843 -1451 0 feedthrough
rlabel pdiffusion 850 -1451 850 -1451 0 feedthrough
rlabel pdiffusion 857 -1451 857 -1451 0 feedthrough
rlabel pdiffusion 864 -1451 864 -1451 0 feedthrough
rlabel pdiffusion 871 -1451 871 -1451 0 feedthrough
rlabel pdiffusion 878 -1451 878 -1451 0 feedthrough
rlabel pdiffusion 885 -1451 885 -1451 0 feedthrough
rlabel pdiffusion 892 -1451 892 -1451 0 feedthrough
rlabel pdiffusion 899 -1451 899 -1451 0 feedthrough
rlabel pdiffusion 906 -1451 906 -1451 0 feedthrough
rlabel pdiffusion 913 -1451 913 -1451 0 feedthrough
rlabel pdiffusion 920 -1451 920 -1451 0 feedthrough
rlabel pdiffusion 927 -1451 927 -1451 0 feedthrough
rlabel pdiffusion 934 -1451 934 -1451 0 feedthrough
rlabel pdiffusion 941 -1451 941 -1451 0 feedthrough
rlabel pdiffusion 948 -1451 948 -1451 0 feedthrough
rlabel pdiffusion 955 -1451 955 -1451 0 feedthrough
rlabel pdiffusion 962 -1451 962 -1451 0 feedthrough
rlabel pdiffusion 969 -1451 969 -1451 0 feedthrough
rlabel pdiffusion 976 -1451 976 -1451 0 feedthrough
rlabel pdiffusion 983 -1451 983 -1451 0 feedthrough
rlabel pdiffusion 990 -1451 990 -1451 0 feedthrough
rlabel pdiffusion 997 -1451 997 -1451 0 feedthrough
rlabel pdiffusion 1004 -1451 1004 -1451 0 feedthrough
rlabel pdiffusion 1011 -1451 1011 -1451 0 feedthrough
rlabel pdiffusion 1018 -1451 1018 -1451 0 feedthrough
rlabel pdiffusion 1025 -1451 1025 -1451 0 feedthrough
rlabel pdiffusion 1032 -1451 1032 -1451 0 feedthrough
rlabel pdiffusion 1039 -1451 1039 -1451 0 feedthrough
rlabel pdiffusion 1046 -1451 1046 -1451 0 cellNo=841
rlabel pdiffusion 1053 -1451 1053 -1451 0 cellNo=579
rlabel pdiffusion 1060 -1451 1060 -1451 0 feedthrough
rlabel pdiffusion 1067 -1451 1067 -1451 0 feedthrough
rlabel pdiffusion 3 -1534 3 -1534 0 feedthrough
rlabel pdiffusion 10 -1534 10 -1534 0 cellNo=399
rlabel pdiffusion 17 -1534 17 -1534 0 feedthrough
rlabel pdiffusion 24 -1534 24 -1534 0 feedthrough
rlabel pdiffusion 31 -1534 31 -1534 0 feedthrough
rlabel pdiffusion 38 -1534 38 -1534 0 feedthrough
rlabel pdiffusion 45 -1534 45 -1534 0 feedthrough
rlabel pdiffusion 52 -1534 52 -1534 0 feedthrough
rlabel pdiffusion 59 -1534 59 -1534 0 feedthrough
rlabel pdiffusion 66 -1534 66 -1534 0 cellNo=183
rlabel pdiffusion 73 -1534 73 -1534 0 feedthrough
rlabel pdiffusion 80 -1534 80 -1534 0 feedthrough
rlabel pdiffusion 87 -1534 87 -1534 0 feedthrough
rlabel pdiffusion 94 -1534 94 -1534 0 cellNo=882
rlabel pdiffusion 101 -1534 101 -1534 0 feedthrough
rlabel pdiffusion 108 -1534 108 -1534 0 feedthrough
rlabel pdiffusion 115 -1534 115 -1534 0 cellNo=138
rlabel pdiffusion 122 -1534 122 -1534 0 feedthrough
rlabel pdiffusion 129 -1534 129 -1534 0 feedthrough
rlabel pdiffusion 136 -1534 136 -1534 0 cellNo=591
rlabel pdiffusion 143 -1534 143 -1534 0 feedthrough
rlabel pdiffusion 150 -1534 150 -1534 0 feedthrough
rlabel pdiffusion 157 -1534 157 -1534 0 feedthrough
rlabel pdiffusion 164 -1534 164 -1534 0 feedthrough
rlabel pdiffusion 171 -1534 171 -1534 0 feedthrough
rlabel pdiffusion 178 -1534 178 -1534 0 feedthrough
rlabel pdiffusion 185 -1534 185 -1534 0 feedthrough
rlabel pdiffusion 192 -1534 192 -1534 0 feedthrough
rlabel pdiffusion 199 -1534 199 -1534 0 cellNo=155
rlabel pdiffusion 206 -1534 206 -1534 0 feedthrough
rlabel pdiffusion 213 -1534 213 -1534 0 feedthrough
rlabel pdiffusion 220 -1534 220 -1534 0 feedthrough
rlabel pdiffusion 227 -1534 227 -1534 0 feedthrough
rlabel pdiffusion 234 -1534 234 -1534 0 feedthrough
rlabel pdiffusion 241 -1534 241 -1534 0 feedthrough
rlabel pdiffusion 248 -1534 248 -1534 0 feedthrough
rlabel pdiffusion 255 -1534 255 -1534 0 feedthrough
rlabel pdiffusion 262 -1534 262 -1534 0 feedthrough
rlabel pdiffusion 269 -1534 269 -1534 0 feedthrough
rlabel pdiffusion 276 -1534 276 -1534 0 feedthrough
rlabel pdiffusion 283 -1534 283 -1534 0 feedthrough
rlabel pdiffusion 290 -1534 290 -1534 0 cellNo=140
rlabel pdiffusion 297 -1534 297 -1534 0 cellNo=805
rlabel pdiffusion 304 -1534 304 -1534 0 feedthrough
rlabel pdiffusion 311 -1534 311 -1534 0 feedthrough
rlabel pdiffusion 318 -1534 318 -1534 0 feedthrough
rlabel pdiffusion 325 -1534 325 -1534 0 feedthrough
rlabel pdiffusion 332 -1534 332 -1534 0 feedthrough
rlabel pdiffusion 339 -1534 339 -1534 0 feedthrough
rlabel pdiffusion 346 -1534 346 -1534 0 cellNo=804
rlabel pdiffusion 353 -1534 353 -1534 0 cellNo=782
rlabel pdiffusion 360 -1534 360 -1534 0 feedthrough
rlabel pdiffusion 367 -1534 367 -1534 0 feedthrough
rlabel pdiffusion 374 -1534 374 -1534 0 feedthrough
rlabel pdiffusion 381 -1534 381 -1534 0 feedthrough
rlabel pdiffusion 388 -1534 388 -1534 0 feedthrough
rlabel pdiffusion 395 -1534 395 -1534 0 feedthrough
rlabel pdiffusion 402 -1534 402 -1534 0 feedthrough
rlabel pdiffusion 409 -1534 409 -1534 0 cellNo=864
rlabel pdiffusion 416 -1534 416 -1534 0 feedthrough
rlabel pdiffusion 423 -1534 423 -1534 0 feedthrough
rlabel pdiffusion 430 -1534 430 -1534 0 feedthrough
rlabel pdiffusion 437 -1534 437 -1534 0 feedthrough
rlabel pdiffusion 444 -1534 444 -1534 0 feedthrough
rlabel pdiffusion 451 -1534 451 -1534 0 feedthrough
rlabel pdiffusion 458 -1534 458 -1534 0 feedthrough
rlabel pdiffusion 465 -1534 465 -1534 0 cellNo=690
rlabel pdiffusion 472 -1534 472 -1534 0 feedthrough
rlabel pdiffusion 479 -1534 479 -1534 0 feedthrough
rlabel pdiffusion 486 -1534 486 -1534 0 cellNo=1
rlabel pdiffusion 493 -1534 493 -1534 0 feedthrough
rlabel pdiffusion 500 -1534 500 -1534 0 feedthrough
rlabel pdiffusion 507 -1534 507 -1534 0 cellNo=722
rlabel pdiffusion 514 -1534 514 -1534 0 cellNo=824
rlabel pdiffusion 521 -1534 521 -1534 0 cellNo=437
rlabel pdiffusion 528 -1534 528 -1534 0 cellNo=464
rlabel pdiffusion 535 -1534 535 -1534 0 cellNo=203
rlabel pdiffusion 542 -1534 542 -1534 0 cellNo=476
rlabel pdiffusion 549 -1534 549 -1534 0 feedthrough
rlabel pdiffusion 556 -1534 556 -1534 0 feedthrough
rlabel pdiffusion 563 -1534 563 -1534 0 cellNo=261
rlabel pdiffusion 570 -1534 570 -1534 0 feedthrough
rlabel pdiffusion 577 -1534 577 -1534 0 feedthrough
rlabel pdiffusion 584 -1534 584 -1534 0 feedthrough
rlabel pdiffusion 591 -1534 591 -1534 0 cellNo=526
rlabel pdiffusion 598 -1534 598 -1534 0 feedthrough
rlabel pdiffusion 605 -1534 605 -1534 0 cellNo=652
rlabel pdiffusion 612 -1534 612 -1534 0 feedthrough
rlabel pdiffusion 619 -1534 619 -1534 0 cellNo=397
rlabel pdiffusion 626 -1534 626 -1534 0 feedthrough
rlabel pdiffusion 633 -1534 633 -1534 0 feedthrough
rlabel pdiffusion 640 -1534 640 -1534 0 feedthrough
rlabel pdiffusion 647 -1534 647 -1534 0 feedthrough
rlabel pdiffusion 654 -1534 654 -1534 0 feedthrough
rlabel pdiffusion 661 -1534 661 -1534 0 cellNo=547
rlabel pdiffusion 668 -1534 668 -1534 0 feedthrough
rlabel pdiffusion 675 -1534 675 -1534 0 feedthrough
rlabel pdiffusion 682 -1534 682 -1534 0 cellNo=325
rlabel pdiffusion 689 -1534 689 -1534 0 feedthrough
rlabel pdiffusion 696 -1534 696 -1534 0 feedthrough
rlabel pdiffusion 703 -1534 703 -1534 0 feedthrough
rlabel pdiffusion 710 -1534 710 -1534 0 feedthrough
rlabel pdiffusion 717 -1534 717 -1534 0 feedthrough
rlabel pdiffusion 724 -1534 724 -1534 0 cellNo=677
rlabel pdiffusion 731 -1534 731 -1534 0 feedthrough
rlabel pdiffusion 738 -1534 738 -1534 0 cellNo=778
rlabel pdiffusion 745 -1534 745 -1534 0 feedthrough
rlabel pdiffusion 752 -1534 752 -1534 0 feedthrough
rlabel pdiffusion 759 -1534 759 -1534 0 feedthrough
rlabel pdiffusion 766 -1534 766 -1534 0 feedthrough
rlabel pdiffusion 773 -1534 773 -1534 0 feedthrough
rlabel pdiffusion 780 -1534 780 -1534 0 feedthrough
rlabel pdiffusion 787 -1534 787 -1534 0 feedthrough
rlabel pdiffusion 794 -1534 794 -1534 0 feedthrough
rlabel pdiffusion 801 -1534 801 -1534 0 feedthrough
rlabel pdiffusion 808 -1534 808 -1534 0 feedthrough
rlabel pdiffusion 815 -1534 815 -1534 0 feedthrough
rlabel pdiffusion 822 -1534 822 -1534 0 feedthrough
rlabel pdiffusion 829 -1534 829 -1534 0 feedthrough
rlabel pdiffusion 836 -1534 836 -1534 0 feedthrough
rlabel pdiffusion 843 -1534 843 -1534 0 cellNo=316
rlabel pdiffusion 850 -1534 850 -1534 0 feedthrough
rlabel pdiffusion 857 -1534 857 -1534 0 feedthrough
rlabel pdiffusion 864 -1534 864 -1534 0 feedthrough
rlabel pdiffusion 871 -1534 871 -1534 0 feedthrough
rlabel pdiffusion 878 -1534 878 -1534 0 feedthrough
rlabel pdiffusion 885 -1534 885 -1534 0 feedthrough
rlabel pdiffusion 892 -1534 892 -1534 0 feedthrough
rlabel pdiffusion 899 -1534 899 -1534 0 feedthrough
rlabel pdiffusion 906 -1534 906 -1534 0 feedthrough
rlabel pdiffusion 913 -1534 913 -1534 0 feedthrough
rlabel pdiffusion 920 -1534 920 -1534 0 feedthrough
rlabel pdiffusion 927 -1534 927 -1534 0 feedthrough
rlabel pdiffusion 934 -1534 934 -1534 0 feedthrough
rlabel pdiffusion 941 -1534 941 -1534 0 feedthrough
rlabel pdiffusion 948 -1534 948 -1534 0 feedthrough
rlabel pdiffusion 955 -1534 955 -1534 0 feedthrough
rlabel pdiffusion 962 -1534 962 -1534 0 feedthrough
rlabel pdiffusion 969 -1534 969 -1534 0 feedthrough
rlabel pdiffusion 976 -1534 976 -1534 0 feedthrough
rlabel pdiffusion 983 -1534 983 -1534 0 feedthrough
rlabel pdiffusion 990 -1534 990 -1534 0 feedthrough
rlabel pdiffusion 997 -1534 997 -1534 0 cellNo=147
rlabel pdiffusion 1004 -1534 1004 -1534 0 feedthrough
rlabel pdiffusion 1011 -1534 1011 -1534 0 feedthrough
rlabel pdiffusion 1018 -1534 1018 -1534 0 feedthrough
rlabel pdiffusion 1046 -1534 1046 -1534 0 feedthrough
rlabel pdiffusion 1053 -1534 1053 -1534 0 feedthrough
rlabel pdiffusion 1060 -1534 1060 -1534 0 cellNo=638
rlabel pdiffusion 3 -1611 3 -1611 0 cellNo=167
rlabel pdiffusion 10 -1611 10 -1611 0 cellNo=424
rlabel pdiffusion 24 -1611 24 -1611 0 feedthrough
rlabel pdiffusion 31 -1611 31 -1611 0 feedthrough
rlabel pdiffusion 38 -1611 38 -1611 0 feedthrough
rlabel pdiffusion 45 -1611 45 -1611 0 feedthrough
rlabel pdiffusion 52 -1611 52 -1611 0 feedthrough
rlabel pdiffusion 59 -1611 59 -1611 0 feedthrough
rlabel pdiffusion 66 -1611 66 -1611 0 cellNo=576
rlabel pdiffusion 73 -1611 73 -1611 0 cellNo=692
rlabel pdiffusion 80 -1611 80 -1611 0 feedthrough
rlabel pdiffusion 87 -1611 87 -1611 0 feedthrough
rlabel pdiffusion 94 -1611 94 -1611 0 feedthrough
rlabel pdiffusion 101 -1611 101 -1611 0 feedthrough
rlabel pdiffusion 108 -1611 108 -1611 0 cellNo=10
rlabel pdiffusion 115 -1611 115 -1611 0 feedthrough
rlabel pdiffusion 122 -1611 122 -1611 0 feedthrough
rlabel pdiffusion 129 -1611 129 -1611 0 feedthrough
rlabel pdiffusion 136 -1611 136 -1611 0 feedthrough
rlabel pdiffusion 143 -1611 143 -1611 0 feedthrough
rlabel pdiffusion 150 -1611 150 -1611 0 cellNo=765
rlabel pdiffusion 157 -1611 157 -1611 0 cellNo=809
rlabel pdiffusion 164 -1611 164 -1611 0 feedthrough
rlabel pdiffusion 171 -1611 171 -1611 0 cellNo=675
rlabel pdiffusion 178 -1611 178 -1611 0 feedthrough
rlabel pdiffusion 185 -1611 185 -1611 0 feedthrough
rlabel pdiffusion 192 -1611 192 -1611 0 feedthrough
rlabel pdiffusion 199 -1611 199 -1611 0 cellNo=884
rlabel pdiffusion 206 -1611 206 -1611 0 feedthrough
rlabel pdiffusion 213 -1611 213 -1611 0 feedthrough
rlabel pdiffusion 220 -1611 220 -1611 0 feedthrough
rlabel pdiffusion 227 -1611 227 -1611 0 cellNo=637
rlabel pdiffusion 234 -1611 234 -1611 0 feedthrough
rlabel pdiffusion 241 -1611 241 -1611 0 feedthrough
rlabel pdiffusion 248 -1611 248 -1611 0 feedthrough
rlabel pdiffusion 255 -1611 255 -1611 0 feedthrough
rlabel pdiffusion 262 -1611 262 -1611 0 feedthrough
rlabel pdiffusion 269 -1611 269 -1611 0 feedthrough
rlabel pdiffusion 276 -1611 276 -1611 0 feedthrough
rlabel pdiffusion 283 -1611 283 -1611 0 feedthrough
rlabel pdiffusion 290 -1611 290 -1611 0 feedthrough
rlabel pdiffusion 297 -1611 297 -1611 0 feedthrough
rlabel pdiffusion 304 -1611 304 -1611 0 cellNo=386
rlabel pdiffusion 311 -1611 311 -1611 0 cellNo=849
rlabel pdiffusion 318 -1611 318 -1611 0 feedthrough
rlabel pdiffusion 325 -1611 325 -1611 0 feedthrough
rlabel pdiffusion 332 -1611 332 -1611 0 feedthrough
rlabel pdiffusion 339 -1611 339 -1611 0 feedthrough
rlabel pdiffusion 346 -1611 346 -1611 0 feedthrough
rlabel pdiffusion 353 -1611 353 -1611 0 cellNo=655
rlabel pdiffusion 360 -1611 360 -1611 0 feedthrough
rlabel pdiffusion 367 -1611 367 -1611 0 feedthrough
rlabel pdiffusion 374 -1611 374 -1611 0 cellNo=667
rlabel pdiffusion 381 -1611 381 -1611 0 feedthrough
rlabel pdiffusion 388 -1611 388 -1611 0 cellNo=694
rlabel pdiffusion 395 -1611 395 -1611 0 cellNo=88
rlabel pdiffusion 402 -1611 402 -1611 0 feedthrough
rlabel pdiffusion 409 -1611 409 -1611 0 feedthrough
rlabel pdiffusion 416 -1611 416 -1611 0 feedthrough
rlabel pdiffusion 423 -1611 423 -1611 0 cellNo=540
rlabel pdiffusion 430 -1611 430 -1611 0 feedthrough
rlabel pdiffusion 437 -1611 437 -1611 0 feedthrough
rlabel pdiffusion 444 -1611 444 -1611 0 feedthrough
rlabel pdiffusion 451 -1611 451 -1611 0 feedthrough
rlabel pdiffusion 458 -1611 458 -1611 0 feedthrough
rlabel pdiffusion 465 -1611 465 -1611 0 feedthrough
rlabel pdiffusion 472 -1611 472 -1611 0 feedthrough
rlabel pdiffusion 479 -1611 479 -1611 0 feedthrough
rlabel pdiffusion 486 -1611 486 -1611 0 feedthrough
rlabel pdiffusion 493 -1611 493 -1611 0 feedthrough
rlabel pdiffusion 500 -1611 500 -1611 0 feedthrough
rlabel pdiffusion 507 -1611 507 -1611 0 feedthrough
rlabel pdiffusion 514 -1611 514 -1611 0 feedthrough
rlabel pdiffusion 521 -1611 521 -1611 0 cellNo=719
rlabel pdiffusion 528 -1611 528 -1611 0 cellNo=89
rlabel pdiffusion 535 -1611 535 -1611 0 feedthrough
rlabel pdiffusion 542 -1611 542 -1611 0 feedthrough
rlabel pdiffusion 549 -1611 549 -1611 0 feedthrough
rlabel pdiffusion 556 -1611 556 -1611 0 cellNo=466
rlabel pdiffusion 563 -1611 563 -1611 0 cellNo=123
rlabel pdiffusion 570 -1611 570 -1611 0 cellNo=715
rlabel pdiffusion 577 -1611 577 -1611 0 feedthrough
rlabel pdiffusion 584 -1611 584 -1611 0 feedthrough
rlabel pdiffusion 591 -1611 591 -1611 0 feedthrough
rlabel pdiffusion 598 -1611 598 -1611 0 feedthrough
rlabel pdiffusion 605 -1611 605 -1611 0 feedthrough
rlabel pdiffusion 612 -1611 612 -1611 0 cellNo=452
rlabel pdiffusion 619 -1611 619 -1611 0 feedthrough
rlabel pdiffusion 626 -1611 626 -1611 0 cellNo=691
rlabel pdiffusion 633 -1611 633 -1611 0 feedthrough
rlabel pdiffusion 640 -1611 640 -1611 0 feedthrough
rlabel pdiffusion 647 -1611 647 -1611 0 feedthrough
rlabel pdiffusion 654 -1611 654 -1611 0 feedthrough
rlabel pdiffusion 661 -1611 661 -1611 0 feedthrough
rlabel pdiffusion 668 -1611 668 -1611 0 feedthrough
rlabel pdiffusion 675 -1611 675 -1611 0 feedthrough
rlabel pdiffusion 682 -1611 682 -1611 0 cellNo=12
rlabel pdiffusion 689 -1611 689 -1611 0 feedthrough
rlabel pdiffusion 696 -1611 696 -1611 0 cellNo=594
rlabel pdiffusion 703 -1611 703 -1611 0 feedthrough
rlabel pdiffusion 710 -1611 710 -1611 0 feedthrough
rlabel pdiffusion 717 -1611 717 -1611 0 feedthrough
rlabel pdiffusion 724 -1611 724 -1611 0 feedthrough
rlabel pdiffusion 731 -1611 731 -1611 0 feedthrough
rlabel pdiffusion 738 -1611 738 -1611 0 feedthrough
rlabel pdiffusion 745 -1611 745 -1611 0 feedthrough
rlabel pdiffusion 752 -1611 752 -1611 0 feedthrough
rlabel pdiffusion 759 -1611 759 -1611 0 feedthrough
rlabel pdiffusion 766 -1611 766 -1611 0 feedthrough
rlabel pdiffusion 773 -1611 773 -1611 0 feedthrough
rlabel pdiffusion 780 -1611 780 -1611 0 feedthrough
rlabel pdiffusion 787 -1611 787 -1611 0 feedthrough
rlabel pdiffusion 794 -1611 794 -1611 0 feedthrough
rlabel pdiffusion 801 -1611 801 -1611 0 feedthrough
rlabel pdiffusion 808 -1611 808 -1611 0 feedthrough
rlabel pdiffusion 815 -1611 815 -1611 0 feedthrough
rlabel pdiffusion 822 -1611 822 -1611 0 feedthrough
rlabel pdiffusion 829 -1611 829 -1611 0 feedthrough
rlabel pdiffusion 836 -1611 836 -1611 0 feedthrough
rlabel pdiffusion 843 -1611 843 -1611 0 feedthrough
rlabel pdiffusion 850 -1611 850 -1611 0 feedthrough
rlabel pdiffusion 857 -1611 857 -1611 0 cellNo=283
rlabel pdiffusion 864 -1611 864 -1611 0 feedthrough
rlabel pdiffusion 871 -1611 871 -1611 0 feedthrough
rlabel pdiffusion 878 -1611 878 -1611 0 feedthrough
rlabel pdiffusion 885 -1611 885 -1611 0 feedthrough
rlabel pdiffusion 892 -1611 892 -1611 0 feedthrough
rlabel pdiffusion 899 -1611 899 -1611 0 feedthrough
rlabel pdiffusion 906 -1611 906 -1611 0 feedthrough
rlabel pdiffusion 913 -1611 913 -1611 0 feedthrough
rlabel pdiffusion 920 -1611 920 -1611 0 feedthrough
rlabel pdiffusion 927 -1611 927 -1611 0 feedthrough
rlabel pdiffusion 934 -1611 934 -1611 0 cellNo=77
rlabel pdiffusion 941 -1611 941 -1611 0 feedthrough
rlabel pdiffusion 948 -1611 948 -1611 0 feedthrough
rlabel pdiffusion 955 -1611 955 -1611 0 feedthrough
rlabel pdiffusion 962 -1611 962 -1611 0 feedthrough
rlabel pdiffusion 1025 -1611 1025 -1611 0 feedthrough
rlabel pdiffusion 1039 -1611 1039 -1611 0 feedthrough
rlabel pdiffusion 1046 -1611 1046 -1611 0 cellNo=720
rlabel pdiffusion 1053 -1611 1053 -1611 0 cellNo=105
rlabel pdiffusion 3 -1676 3 -1676 0 cellNo=469
rlabel pdiffusion 10 -1676 10 -1676 0 cellNo=673
rlabel pdiffusion 38 -1676 38 -1676 0 cellNo=733
rlabel pdiffusion 45 -1676 45 -1676 0 cellNo=127
rlabel pdiffusion 52 -1676 52 -1676 0 feedthrough
rlabel pdiffusion 66 -1676 66 -1676 0 feedthrough
rlabel pdiffusion 73 -1676 73 -1676 0 cellNo=599
rlabel pdiffusion 80 -1676 80 -1676 0 cellNo=750
rlabel pdiffusion 87 -1676 87 -1676 0 feedthrough
rlabel pdiffusion 94 -1676 94 -1676 0 feedthrough
rlabel pdiffusion 101 -1676 101 -1676 0 feedthrough
rlabel pdiffusion 108 -1676 108 -1676 0 feedthrough
rlabel pdiffusion 115 -1676 115 -1676 0 cellNo=187
rlabel pdiffusion 122 -1676 122 -1676 0 feedthrough
rlabel pdiffusion 129 -1676 129 -1676 0 feedthrough
rlabel pdiffusion 136 -1676 136 -1676 0 feedthrough
rlabel pdiffusion 143 -1676 143 -1676 0 feedthrough
rlabel pdiffusion 150 -1676 150 -1676 0 cellNo=829
rlabel pdiffusion 157 -1676 157 -1676 0 feedthrough
rlabel pdiffusion 164 -1676 164 -1676 0 feedthrough
rlabel pdiffusion 171 -1676 171 -1676 0 feedthrough
rlabel pdiffusion 178 -1676 178 -1676 0 cellNo=663
rlabel pdiffusion 185 -1676 185 -1676 0 feedthrough
rlabel pdiffusion 192 -1676 192 -1676 0 feedthrough
rlabel pdiffusion 199 -1676 199 -1676 0 cellNo=533
rlabel pdiffusion 206 -1676 206 -1676 0 cellNo=847
rlabel pdiffusion 213 -1676 213 -1676 0 feedthrough
rlabel pdiffusion 220 -1676 220 -1676 0 feedthrough
rlabel pdiffusion 227 -1676 227 -1676 0 feedthrough
rlabel pdiffusion 234 -1676 234 -1676 0 feedthrough
rlabel pdiffusion 241 -1676 241 -1676 0 feedthrough
rlabel pdiffusion 248 -1676 248 -1676 0 feedthrough
rlabel pdiffusion 255 -1676 255 -1676 0 cellNo=724
rlabel pdiffusion 262 -1676 262 -1676 0 feedthrough
rlabel pdiffusion 269 -1676 269 -1676 0 feedthrough
rlabel pdiffusion 276 -1676 276 -1676 0 feedthrough
rlabel pdiffusion 283 -1676 283 -1676 0 feedthrough
rlabel pdiffusion 290 -1676 290 -1676 0 feedthrough
rlabel pdiffusion 297 -1676 297 -1676 0 feedthrough
rlabel pdiffusion 304 -1676 304 -1676 0 cellNo=9
rlabel pdiffusion 311 -1676 311 -1676 0 feedthrough
rlabel pdiffusion 318 -1676 318 -1676 0 feedthrough
rlabel pdiffusion 325 -1676 325 -1676 0 feedthrough
rlabel pdiffusion 332 -1676 332 -1676 0 cellNo=621
rlabel pdiffusion 339 -1676 339 -1676 0 cellNo=298
rlabel pdiffusion 346 -1676 346 -1676 0 feedthrough
rlabel pdiffusion 353 -1676 353 -1676 0 feedthrough
rlabel pdiffusion 360 -1676 360 -1676 0 feedthrough
rlabel pdiffusion 367 -1676 367 -1676 0 feedthrough
rlabel pdiffusion 374 -1676 374 -1676 0 feedthrough
rlabel pdiffusion 381 -1676 381 -1676 0 feedthrough
rlabel pdiffusion 388 -1676 388 -1676 0 feedthrough
rlabel pdiffusion 395 -1676 395 -1676 0 feedthrough
rlabel pdiffusion 402 -1676 402 -1676 0 cellNo=171
rlabel pdiffusion 409 -1676 409 -1676 0 cellNo=489
rlabel pdiffusion 416 -1676 416 -1676 0 feedthrough
rlabel pdiffusion 423 -1676 423 -1676 0 feedthrough
rlabel pdiffusion 430 -1676 430 -1676 0 cellNo=465
rlabel pdiffusion 437 -1676 437 -1676 0 feedthrough
rlabel pdiffusion 444 -1676 444 -1676 0 feedthrough
rlabel pdiffusion 451 -1676 451 -1676 0 feedthrough
rlabel pdiffusion 458 -1676 458 -1676 0 feedthrough
rlabel pdiffusion 465 -1676 465 -1676 0 feedthrough
rlabel pdiffusion 472 -1676 472 -1676 0 feedthrough
rlabel pdiffusion 479 -1676 479 -1676 0 feedthrough
rlabel pdiffusion 486 -1676 486 -1676 0 feedthrough
rlabel pdiffusion 493 -1676 493 -1676 0 feedthrough
rlabel pdiffusion 500 -1676 500 -1676 0 feedthrough
rlabel pdiffusion 507 -1676 507 -1676 0 feedthrough
rlabel pdiffusion 514 -1676 514 -1676 0 cellNo=497
rlabel pdiffusion 521 -1676 521 -1676 0 cellNo=899
rlabel pdiffusion 528 -1676 528 -1676 0 feedthrough
rlabel pdiffusion 535 -1676 535 -1676 0 feedthrough
rlabel pdiffusion 542 -1676 542 -1676 0 cellNo=897
rlabel pdiffusion 549 -1676 549 -1676 0 cellNo=246
rlabel pdiffusion 556 -1676 556 -1676 0 feedthrough
rlabel pdiffusion 563 -1676 563 -1676 0 feedthrough
rlabel pdiffusion 570 -1676 570 -1676 0 feedthrough
rlabel pdiffusion 577 -1676 577 -1676 0 feedthrough
rlabel pdiffusion 584 -1676 584 -1676 0 feedthrough
rlabel pdiffusion 591 -1676 591 -1676 0 feedthrough
rlabel pdiffusion 598 -1676 598 -1676 0 feedthrough
rlabel pdiffusion 605 -1676 605 -1676 0 feedthrough
rlabel pdiffusion 612 -1676 612 -1676 0 feedthrough
rlabel pdiffusion 626 -1676 626 -1676 0 feedthrough
rlabel pdiffusion 633 -1676 633 -1676 0 feedthrough
rlabel pdiffusion 647 -1676 647 -1676 0 feedthrough
rlabel pdiffusion 668 -1676 668 -1676 0 feedthrough
rlabel pdiffusion 675 -1676 675 -1676 0 cellNo=808
rlabel pdiffusion 682 -1676 682 -1676 0 feedthrough
rlabel pdiffusion 689 -1676 689 -1676 0 cellNo=706
rlabel pdiffusion 696 -1676 696 -1676 0 feedthrough
rlabel pdiffusion 703 -1676 703 -1676 0 feedthrough
rlabel pdiffusion 710 -1676 710 -1676 0 feedthrough
rlabel pdiffusion 717 -1676 717 -1676 0 feedthrough
rlabel pdiffusion 724 -1676 724 -1676 0 feedthrough
rlabel pdiffusion 731 -1676 731 -1676 0 cellNo=458
rlabel pdiffusion 738 -1676 738 -1676 0 feedthrough
rlabel pdiffusion 745 -1676 745 -1676 0 feedthrough
rlabel pdiffusion 752 -1676 752 -1676 0 feedthrough
rlabel pdiffusion 759 -1676 759 -1676 0 feedthrough
rlabel pdiffusion 766 -1676 766 -1676 0 feedthrough
rlabel pdiffusion 773 -1676 773 -1676 0 cellNo=143
rlabel pdiffusion 780 -1676 780 -1676 0 cellNo=583
rlabel pdiffusion 787 -1676 787 -1676 0 feedthrough
rlabel pdiffusion 794 -1676 794 -1676 0 feedthrough
rlabel pdiffusion 801 -1676 801 -1676 0 cellNo=205
rlabel pdiffusion 808 -1676 808 -1676 0 feedthrough
rlabel pdiffusion 815 -1676 815 -1676 0 feedthrough
rlabel pdiffusion 822 -1676 822 -1676 0 feedthrough
rlabel pdiffusion 829 -1676 829 -1676 0 feedthrough
rlabel pdiffusion 836 -1676 836 -1676 0 cellNo=360
rlabel pdiffusion 843 -1676 843 -1676 0 feedthrough
rlabel pdiffusion 850 -1676 850 -1676 0 cellNo=862
rlabel pdiffusion 864 -1676 864 -1676 0 feedthrough
rlabel pdiffusion 885 -1676 885 -1676 0 feedthrough
rlabel pdiffusion 892 -1676 892 -1676 0 feedthrough
rlabel pdiffusion 906 -1676 906 -1676 0 feedthrough
rlabel pdiffusion 969 -1676 969 -1676 0 feedthrough
rlabel pdiffusion 1025 -1676 1025 -1676 0 feedthrough
rlabel pdiffusion 3 -1713 3 -1713 0 cellNo=99
rlabel pdiffusion 10 -1713 10 -1713 0 cellNo=278
rlabel pdiffusion 17 -1713 17 -1713 0 cellNo=366
rlabel pdiffusion 24 -1713 24 -1713 0 cellNo=662
rlabel pdiffusion 31 -1713 31 -1713 0 cellNo=780
rlabel pdiffusion 45 -1713 45 -1713 0 feedthrough
rlabel pdiffusion 59 -1713 59 -1713 0 feedthrough
rlabel pdiffusion 94 -1713 94 -1713 0 feedthrough
rlabel pdiffusion 101 -1713 101 -1713 0 cellNo=741
rlabel pdiffusion 115 -1713 115 -1713 0 cellNo=550
rlabel pdiffusion 129 -1713 129 -1713 0 feedthrough
rlabel pdiffusion 143 -1713 143 -1713 0 feedthrough
rlabel pdiffusion 150 -1713 150 -1713 0 feedthrough
rlabel pdiffusion 157 -1713 157 -1713 0 feedthrough
rlabel pdiffusion 164 -1713 164 -1713 0 feedthrough
rlabel pdiffusion 171 -1713 171 -1713 0 feedthrough
rlabel pdiffusion 178 -1713 178 -1713 0 cellNo=743
rlabel pdiffusion 185 -1713 185 -1713 0 cellNo=451
rlabel pdiffusion 192 -1713 192 -1713 0 feedthrough
rlabel pdiffusion 199 -1713 199 -1713 0 cellNo=727
rlabel pdiffusion 206 -1713 206 -1713 0 cellNo=762
rlabel pdiffusion 213 -1713 213 -1713 0 cellNo=482
rlabel pdiffusion 220 -1713 220 -1713 0 feedthrough
rlabel pdiffusion 227 -1713 227 -1713 0 feedthrough
rlabel pdiffusion 234 -1713 234 -1713 0 feedthrough
rlabel pdiffusion 241 -1713 241 -1713 0 feedthrough
rlabel pdiffusion 255 -1713 255 -1713 0 feedthrough
rlabel pdiffusion 262 -1713 262 -1713 0 cellNo=840
rlabel pdiffusion 269 -1713 269 -1713 0 feedthrough
rlabel pdiffusion 276 -1713 276 -1713 0 cellNo=329
rlabel pdiffusion 283 -1713 283 -1713 0 feedthrough
rlabel pdiffusion 290 -1713 290 -1713 0 feedthrough
rlabel pdiffusion 297 -1713 297 -1713 0 cellNo=877
rlabel pdiffusion 304 -1713 304 -1713 0 feedthrough
rlabel pdiffusion 311 -1713 311 -1713 0 feedthrough
rlabel pdiffusion 318 -1713 318 -1713 0 feedthrough
rlabel pdiffusion 325 -1713 325 -1713 0 feedthrough
rlabel pdiffusion 332 -1713 332 -1713 0 feedthrough
rlabel pdiffusion 339 -1713 339 -1713 0 cellNo=853
rlabel pdiffusion 346 -1713 346 -1713 0 feedthrough
rlabel pdiffusion 353 -1713 353 -1713 0 cellNo=779
rlabel pdiffusion 360 -1713 360 -1713 0 feedthrough
rlabel pdiffusion 367 -1713 367 -1713 0 feedthrough
rlabel pdiffusion 374 -1713 374 -1713 0 cellNo=422
rlabel pdiffusion 381 -1713 381 -1713 0 cellNo=531
rlabel pdiffusion 388 -1713 388 -1713 0 feedthrough
rlabel pdiffusion 395 -1713 395 -1713 0 feedthrough
rlabel pdiffusion 402 -1713 402 -1713 0 cellNo=839
rlabel pdiffusion 409 -1713 409 -1713 0 feedthrough
rlabel pdiffusion 416 -1713 416 -1713 0 feedthrough
rlabel pdiffusion 423 -1713 423 -1713 0 feedthrough
rlabel pdiffusion 430 -1713 430 -1713 0 feedthrough
rlabel pdiffusion 437 -1713 437 -1713 0 feedthrough
rlabel pdiffusion 444 -1713 444 -1713 0 feedthrough
rlabel pdiffusion 451 -1713 451 -1713 0 feedthrough
rlabel pdiffusion 458 -1713 458 -1713 0 feedthrough
rlabel pdiffusion 465 -1713 465 -1713 0 feedthrough
rlabel pdiffusion 472 -1713 472 -1713 0 cellNo=76
rlabel pdiffusion 479 -1713 479 -1713 0 feedthrough
rlabel pdiffusion 486 -1713 486 -1713 0 feedthrough
rlabel pdiffusion 493 -1713 493 -1713 0 feedthrough
rlabel pdiffusion 500 -1713 500 -1713 0 cellNo=769
rlabel pdiffusion 507 -1713 507 -1713 0 feedthrough
rlabel pdiffusion 514 -1713 514 -1713 0 feedthrough
rlabel pdiffusion 521 -1713 521 -1713 0 feedthrough
rlabel pdiffusion 528 -1713 528 -1713 0 feedthrough
rlabel pdiffusion 535 -1713 535 -1713 0 feedthrough
rlabel pdiffusion 542 -1713 542 -1713 0 feedthrough
rlabel pdiffusion 549 -1713 549 -1713 0 feedthrough
rlabel pdiffusion 556 -1713 556 -1713 0 feedthrough
rlabel pdiffusion 563 -1713 563 -1713 0 feedthrough
rlabel pdiffusion 570 -1713 570 -1713 0 feedthrough
rlabel pdiffusion 577 -1713 577 -1713 0 feedthrough
rlabel pdiffusion 584 -1713 584 -1713 0 feedthrough
rlabel pdiffusion 591 -1713 591 -1713 0 cellNo=192
rlabel pdiffusion 598 -1713 598 -1713 0 cellNo=349
rlabel pdiffusion 605 -1713 605 -1713 0 cellNo=816
rlabel pdiffusion 612 -1713 612 -1713 0 cellNo=626
rlabel pdiffusion 619 -1713 619 -1713 0 feedthrough
rlabel pdiffusion 640 -1713 640 -1713 0 feedthrough
rlabel pdiffusion 647 -1713 647 -1713 0 feedthrough
rlabel pdiffusion 654 -1713 654 -1713 0 feedthrough
rlabel pdiffusion 675 -1713 675 -1713 0 feedthrough
rlabel pdiffusion 682 -1713 682 -1713 0 cellNo=685
rlabel pdiffusion 710 -1713 710 -1713 0 feedthrough
rlabel pdiffusion 724 -1713 724 -1713 0 feedthrough
rlabel pdiffusion 731 -1713 731 -1713 0 feedthrough
rlabel pdiffusion 738 -1713 738 -1713 0 feedthrough
rlabel pdiffusion 745 -1713 745 -1713 0 feedthrough
rlabel pdiffusion 752 -1713 752 -1713 0 feedthrough
rlabel pdiffusion 759 -1713 759 -1713 0 feedthrough
rlabel pdiffusion 766 -1713 766 -1713 0 feedthrough
rlabel pdiffusion 773 -1713 773 -1713 0 feedthrough
rlabel pdiffusion 780 -1713 780 -1713 0 feedthrough
rlabel pdiffusion 794 -1713 794 -1713 0 feedthrough
rlabel pdiffusion 801 -1713 801 -1713 0 feedthrough
rlabel pdiffusion 808 -1713 808 -1713 0 feedthrough
rlabel pdiffusion 815 -1713 815 -1713 0 cellNo=751
rlabel pdiffusion 822 -1713 822 -1713 0 feedthrough
rlabel pdiffusion 829 -1713 829 -1713 0 feedthrough
rlabel pdiffusion 836 -1713 836 -1713 0 feedthrough
rlabel pdiffusion 843 -1713 843 -1713 0 cellNo=753
rlabel pdiffusion 850 -1713 850 -1713 0 feedthrough
rlabel pdiffusion 857 -1713 857 -1713 0 feedthrough
rlabel pdiffusion 864 -1713 864 -1713 0 cellNo=134
rlabel pdiffusion 885 -1713 885 -1713 0 feedthrough
rlabel pdiffusion 899 -1713 899 -1713 0 feedthrough
rlabel pdiffusion 969 -1713 969 -1713 0 feedthrough
rlabel pdiffusion 1025 -1713 1025 -1713 0 feedthrough
rlabel pdiffusion 3 -1746 3 -1746 0 cellNo=345
rlabel pdiffusion 10 -1746 10 -1746 0 cellNo=581
rlabel pdiffusion 17 -1746 17 -1746 0 cellNo=479
rlabel pdiffusion 45 -1746 45 -1746 0 feedthrough
rlabel pdiffusion 59 -1746 59 -1746 0 cellNo=693
rlabel pdiffusion 66 -1746 66 -1746 0 feedthrough
rlabel pdiffusion 101 -1746 101 -1746 0 feedthrough
rlabel pdiffusion 108 -1746 108 -1746 0 feedthrough
rlabel pdiffusion 115 -1746 115 -1746 0 cellNo=429
rlabel pdiffusion 122 -1746 122 -1746 0 feedthrough
rlabel pdiffusion 129 -1746 129 -1746 0 cellNo=200
rlabel pdiffusion 136 -1746 136 -1746 0 cellNo=330
rlabel pdiffusion 143 -1746 143 -1746 0 cellNo=584
rlabel pdiffusion 150 -1746 150 -1746 0 cellNo=328
rlabel pdiffusion 157 -1746 157 -1746 0 cellNo=814
rlabel pdiffusion 164 -1746 164 -1746 0 feedthrough
rlabel pdiffusion 171 -1746 171 -1746 0 cellNo=752
rlabel pdiffusion 178 -1746 178 -1746 0 feedthrough
rlabel pdiffusion 185 -1746 185 -1746 0 feedthrough
rlabel pdiffusion 192 -1746 192 -1746 0 feedthrough
rlabel pdiffusion 206 -1746 206 -1746 0 feedthrough
rlabel pdiffusion 213 -1746 213 -1746 0 cellNo=758
rlabel pdiffusion 220 -1746 220 -1746 0 cellNo=772
rlabel pdiffusion 227 -1746 227 -1746 0 cellNo=761
rlabel pdiffusion 234 -1746 234 -1746 0 feedthrough
rlabel pdiffusion 241 -1746 241 -1746 0 feedthrough
rlabel pdiffusion 248 -1746 248 -1746 0 feedthrough
rlabel pdiffusion 276 -1746 276 -1746 0 feedthrough
rlabel pdiffusion 297 -1746 297 -1746 0 feedthrough
rlabel pdiffusion 304 -1746 304 -1746 0 feedthrough
rlabel pdiffusion 311 -1746 311 -1746 0 feedthrough
rlabel pdiffusion 318 -1746 318 -1746 0 feedthrough
rlabel pdiffusion 325 -1746 325 -1746 0 feedthrough
rlabel pdiffusion 332 -1746 332 -1746 0 feedthrough
rlabel pdiffusion 339 -1746 339 -1746 0 feedthrough
rlabel pdiffusion 346 -1746 346 -1746 0 feedthrough
rlabel pdiffusion 353 -1746 353 -1746 0 feedthrough
rlabel pdiffusion 360 -1746 360 -1746 0 feedthrough
rlabel pdiffusion 367 -1746 367 -1746 0 cellNo=227
rlabel pdiffusion 374 -1746 374 -1746 0 feedthrough
rlabel pdiffusion 381 -1746 381 -1746 0 feedthrough
rlabel pdiffusion 388 -1746 388 -1746 0 feedthrough
rlabel pdiffusion 395 -1746 395 -1746 0 feedthrough
rlabel pdiffusion 402 -1746 402 -1746 0 cellNo=775
rlabel pdiffusion 409 -1746 409 -1746 0 cellNo=869
rlabel pdiffusion 416 -1746 416 -1746 0 feedthrough
rlabel pdiffusion 423 -1746 423 -1746 0 feedthrough
rlabel pdiffusion 430 -1746 430 -1746 0 feedthrough
rlabel pdiffusion 437 -1746 437 -1746 0 feedthrough
rlabel pdiffusion 444 -1746 444 -1746 0 cellNo=845
rlabel pdiffusion 451 -1746 451 -1746 0 feedthrough
rlabel pdiffusion 458 -1746 458 -1746 0 feedthrough
rlabel pdiffusion 465 -1746 465 -1746 0 feedthrough
rlabel pdiffusion 472 -1746 472 -1746 0 cellNo=707
rlabel pdiffusion 479 -1746 479 -1746 0 feedthrough
rlabel pdiffusion 486 -1746 486 -1746 0 cellNo=590
rlabel pdiffusion 493 -1746 493 -1746 0 feedthrough
rlabel pdiffusion 500 -1746 500 -1746 0 feedthrough
rlabel pdiffusion 507 -1746 507 -1746 0 cellNo=212
rlabel pdiffusion 514 -1746 514 -1746 0 feedthrough
rlabel pdiffusion 521 -1746 521 -1746 0 feedthrough
rlabel pdiffusion 528 -1746 528 -1746 0 cellNo=668
rlabel pdiffusion 535 -1746 535 -1746 0 feedthrough
rlabel pdiffusion 542 -1746 542 -1746 0 feedthrough
rlabel pdiffusion 549 -1746 549 -1746 0 feedthrough
rlabel pdiffusion 556 -1746 556 -1746 0 cellNo=844
rlabel pdiffusion 563 -1746 563 -1746 0 cellNo=544
rlabel pdiffusion 570 -1746 570 -1746 0 feedthrough
rlabel pdiffusion 577 -1746 577 -1746 0 feedthrough
rlabel pdiffusion 584 -1746 584 -1746 0 cellNo=832
rlabel pdiffusion 591 -1746 591 -1746 0 feedthrough
rlabel pdiffusion 598 -1746 598 -1746 0 feedthrough
rlabel pdiffusion 647 -1746 647 -1746 0 feedthrough
rlabel pdiffusion 654 -1746 654 -1746 0 cellNo=810
rlabel pdiffusion 703 -1746 703 -1746 0 feedthrough
rlabel pdiffusion 710 -1746 710 -1746 0 feedthrough
rlabel pdiffusion 717 -1746 717 -1746 0 cellNo=276
rlabel pdiffusion 724 -1746 724 -1746 0 feedthrough
rlabel pdiffusion 731 -1746 731 -1746 0 feedthrough
rlabel pdiffusion 738 -1746 738 -1746 0 feedthrough
rlabel pdiffusion 745 -1746 745 -1746 0 feedthrough
rlabel pdiffusion 752 -1746 752 -1746 0 feedthrough
rlabel pdiffusion 759 -1746 759 -1746 0 feedthrough
rlabel pdiffusion 766 -1746 766 -1746 0 feedthrough
rlabel pdiffusion 773 -1746 773 -1746 0 cellNo=757
rlabel pdiffusion 780 -1746 780 -1746 0 cellNo=713
rlabel pdiffusion 787 -1746 787 -1746 0 feedthrough
rlabel pdiffusion 794 -1746 794 -1746 0 feedthrough
rlabel pdiffusion 801 -1746 801 -1746 0 feedthrough
rlabel pdiffusion 808 -1746 808 -1746 0 feedthrough
rlabel pdiffusion 829 -1746 829 -1746 0 feedthrough
rlabel pdiffusion 843 -1746 843 -1746 0 feedthrough
rlabel pdiffusion 857 -1746 857 -1746 0 feedthrough
rlabel pdiffusion 885 -1746 885 -1746 0 feedthrough
rlabel pdiffusion 899 -1746 899 -1746 0 feedthrough
rlabel pdiffusion 969 -1746 969 -1746 0 feedthrough
rlabel pdiffusion 976 -1746 976 -1746 0 cellNo=831
rlabel pdiffusion 1025 -1746 1025 -1746 0 feedthrough
rlabel pdiffusion 3 -1773 3 -1773 0 cellNo=818
rlabel pdiffusion 10 -1773 10 -1773 0 cellNo=830
rlabel pdiffusion 17 -1773 17 -1773 0 cellNo=838
rlabel pdiffusion 24 -1773 24 -1773 0 cellNo=820
rlabel pdiffusion 31 -1773 31 -1773 0 cellNo=825
rlabel pdiffusion 45 -1773 45 -1773 0 cellNo=812
rlabel pdiffusion 59 -1773 59 -1773 0 feedthrough
rlabel pdiffusion 66 -1773 66 -1773 0 cellNo=875
rlabel pdiffusion 73 -1773 73 -1773 0 feedthrough
rlabel pdiffusion 80 -1773 80 -1773 0 feedthrough
rlabel pdiffusion 94 -1773 94 -1773 0 feedthrough
rlabel pdiffusion 101 -1773 101 -1773 0 cellNo=455
rlabel pdiffusion 108 -1773 108 -1773 0 cellNo=835
rlabel pdiffusion 115 -1773 115 -1773 0 cellNo=867
rlabel pdiffusion 122 -1773 122 -1773 0 cellNo=786
rlabel pdiffusion 129 -1773 129 -1773 0 feedthrough
rlabel pdiffusion 136 -1773 136 -1773 0 feedthrough
rlabel pdiffusion 143 -1773 143 -1773 0 feedthrough
rlabel pdiffusion 150 -1773 150 -1773 0 cellNo=817
rlabel pdiffusion 157 -1773 157 -1773 0 cellNo=295
rlabel pdiffusion 171 -1773 171 -1773 0 feedthrough
rlabel pdiffusion 192 -1773 192 -1773 0 feedthrough
rlabel pdiffusion 199 -1773 199 -1773 0 cellNo=493
rlabel pdiffusion 206 -1773 206 -1773 0 feedthrough
rlabel pdiffusion 213 -1773 213 -1773 0 cellNo=819
rlabel pdiffusion 220 -1773 220 -1773 0 feedthrough
rlabel pdiffusion 227 -1773 227 -1773 0 cellNo=357
rlabel pdiffusion 234 -1773 234 -1773 0 feedthrough
rlabel pdiffusion 241 -1773 241 -1773 0 feedthrough
rlabel pdiffusion 276 -1773 276 -1773 0 feedthrough
rlabel pdiffusion 283 -1773 283 -1773 0 feedthrough
rlabel pdiffusion 290 -1773 290 -1773 0 feedthrough
rlabel pdiffusion 297 -1773 297 -1773 0 feedthrough
rlabel pdiffusion 304 -1773 304 -1773 0 cellNo=811
rlabel pdiffusion 311 -1773 311 -1773 0 feedthrough
rlabel pdiffusion 318 -1773 318 -1773 0 cellNo=373
rlabel pdiffusion 325 -1773 325 -1773 0 feedthrough
rlabel pdiffusion 332 -1773 332 -1773 0 cellNo=837
rlabel pdiffusion 339 -1773 339 -1773 0 feedthrough
rlabel pdiffusion 346 -1773 346 -1773 0 feedthrough
rlabel pdiffusion 353 -1773 353 -1773 0 feedthrough
rlabel pdiffusion 360 -1773 360 -1773 0 cellNo=96
rlabel pdiffusion 367 -1773 367 -1773 0 cellNo=346
rlabel pdiffusion 374 -1773 374 -1773 0 feedthrough
rlabel pdiffusion 381 -1773 381 -1773 0 feedthrough
rlabel pdiffusion 395 -1773 395 -1773 0 feedthrough
rlabel pdiffusion 402 -1773 402 -1773 0 feedthrough
rlabel pdiffusion 409 -1773 409 -1773 0 cellNo=593
rlabel pdiffusion 416 -1773 416 -1773 0 feedthrough
rlabel pdiffusion 423 -1773 423 -1773 0 cellNo=275
rlabel pdiffusion 430 -1773 430 -1773 0 cellNo=568
rlabel pdiffusion 444 -1773 444 -1773 0 feedthrough
rlabel pdiffusion 451 -1773 451 -1773 0 feedthrough
rlabel pdiffusion 458 -1773 458 -1773 0 feedthrough
rlabel pdiffusion 465 -1773 465 -1773 0 feedthrough
rlabel pdiffusion 472 -1773 472 -1773 0 feedthrough
rlabel pdiffusion 479 -1773 479 -1773 0 feedthrough
rlabel pdiffusion 507 -1773 507 -1773 0 feedthrough
rlabel pdiffusion 514 -1773 514 -1773 0 feedthrough
rlabel pdiffusion 528 -1773 528 -1773 0 feedthrough
rlabel pdiffusion 563 -1773 563 -1773 0 feedthrough
rlabel pdiffusion 710 -1773 710 -1773 0 feedthrough
rlabel pdiffusion 717 -1773 717 -1773 0 cellNo=647
rlabel pdiffusion 724 -1773 724 -1773 0 feedthrough
rlabel pdiffusion 731 -1773 731 -1773 0 feedthrough
rlabel pdiffusion 738 -1773 738 -1773 0 feedthrough
rlabel pdiffusion 745 -1773 745 -1773 0 cellNo=460
rlabel pdiffusion 752 -1773 752 -1773 0 feedthrough
rlabel pdiffusion 759 -1773 759 -1773 0 feedthrough
rlabel pdiffusion 773 -1773 773 -1773 0 feedthrough
rlabel pdiffusion 780 -1773 780 -1773 0 cellNo=709
rlabel pdiffusion 794 -1773 794 -1773 0 feedthrough
rlabel pdiffusion 815 -1773 815 -1773 0 feedthrough
rlabel pdiffusion 829 -1773 829 -1773 0 feedthrough
rlabel pdiffusion 843 -1773 843 -1773 0 cellNo=700
rlabel pdiffusion 857 -1773 857 -1773 0 cellNo=833
rlabel pdiffusion 878 -1773 878 -1773 0 cellNo=548
rlabel pdiffusion 885 -1773 885 -1773 0 feedthrough
rlabel pdiffusion 899 -1773 899 -1773 0 feedthrough
rlabel pdiffusion 1025 -1773 1025 -1773 0 feedthrough
rlabel pdiffusion 3 -1794 3 -1794 0 cellNo=219
rlabel pdiffusion 10 -1794 10 -1794 0 cellNo=381
rlabel pdiffusion 17 -1794 17 -1794 0 cellNo=696
rlabel pdiffusion 24 -1794 24 -1794 0 cellNo=245
rlabel pdiffusion 31 -1794 31 -1794 0 cellNo=756
rlabel pdiffusion 38 -1794 38 -1794 0 cellNo=730
rlabel pdiffusion 45 -1794 45 -1794 0 cellNo=475
rlabel pdiffusion 52 -1794 52 -1794 0 cellNo=372
rlabel pdiffusion 59 -1794 59 -1794 0 cellNo=857
rlabel pdiffusion 66 -1794 66 -1794 0 cellNo=850
rlabel pdiffusion 73 -1794 73 -1794 0 cellNo=842
rlabel pdiffusion 80 -1794 80 -1794 0 feedthrough
rlabel pdiffusion 143 -1794 143 -1794 0 feedthrough
rlabel pdiffusion 150 -1794 150 -1794 0 cellNo=763
rlabel pdiffusion 157 -1794 157 -1794 0 feedthrough
rlabel pdiffusion 171 -1794 171 -1794 0 cellNo=858
rlabel pdiffusion 185 -1794 185 -1794 0 cellNo=870
rlabel pdiffusion 206 -1794 206 -1794 0 feedthrough
rlabel pdiffusion 227 -1794 227 -1794 0 feedthrough
rlabel pdiffusion 241 -1794 241 -1794 0 feedthrough
rlabel pdiffusion 248 -1794 248 -1794 0 cellNo=477
rlabel pdiffusion 262 -1794 262 -1794 0 feedthrough
rlabel pdiffusion 283 -1794 283 -1794 0 feedthrough
rlabel pdiffusion 297 -1794 297 -1794 0 feedthrough
rlabel pdiffusion 304 -1794 304 -1794 0 cellNo=29
rlabel pdiffusion 311 -1794 311 -1794 0 cellNo=72
rlabel pdiffusion 318 -1794 318 -1794 0 cellNo=624
rlabel pdiffusion 325 -1794 325 -1794 0 feedthrough
rlabel pdiffusion 332 -1794 332 -1794 0 feedthrough
rlabel pdiffusion 339 -1794 339 -1794 0 feedthrough
rlabel pdiffusion 346 -1794 346 -1794 0 cellNo=468
rlabel pdiffusion 353 -1794 353 -1794 0 feedthrough
rlabel pdiffusion 381 -1794 381 -1794 0 feedthrough
rlabel pdiffusion 388 -1794 388 -1794 0 feedthrough
rlabel pdiffusion 409 -1794 409 -1794 0 cellNo=318
rlabel pdiffusion 416 -1794 416 -1794 0 feedthrough
rlabel pdiffusion 423 -1794 423 -1794 0 feedthrough
rlabel pdiffusion 430 -1794 430 -1794 0 cellNo=863
rlabel pdiffusion 437 -1794 437 -1794 0 cellNo=202
rlabel pdiffusion 444 -1794 444 -1794 0 feedthrough
rlabel pdiffusion 451 -1794 451 -1794 0 feedthrough
rlabel pdiffusion 458 -1794 458 -1794 0 feedthrough
rlabel pdiffusion 472 -1794 472 -1794 0 feedthrough
rlabel pdiffusion 479 -1794 479 -1794 0 feedthrough
rlabel pdiffusion 500 -1794 500 -1794 0 cellNo=861
rlabel pdiffusion 507 -1794 507 -1794 0 cellNo=773
rlabel pdiffusion 514 -1794 514 -1794 0 feedthrough
rlabel pdiffusion 521 -1794 521 -1794 0 feedthrough
rlabel pdiffusion 563 -1794 563 -1794 0 cellNo=305
rlabel pdiffusion 738 -1794 738 -1794 0 feedthrough
rlabel pdiffusion 745 -1794 745 -1794 0 cellNo=467
rlabel pdiffusion 752 -1794 752 -1794 0 cellNo=580
rlabel pdiffusion 759 -1794 759 -1794 0 feedthrough
rlabel pdiffusion 766 -1794 766 -1794 0 feedthrough
rlabel pdiffusion 773 -1794 773 -1794 0 cellNo=415
rlabel pdiffusion 794 -1794 794 -1794 0 feedthrough
rlabel pdiffusion 815 -1794 815 -1794 0 cellNo=868
rlabel pdiffusion 836 -1794 836 -1794 0 cellNo=485
rlabel pdiffusion 899 -1794 899 -1794 0 feedthrough
rlabel pdiffusion 1025 -1794 1025 -1794 0 feedthrough
rlabel pdiffusion 3 -1809 3 -1809 0 cellNo=292
rlabel pdiffusion 10 -1809 10 -1809 0 cellNo=871
rlabel pdiffusion 17 -1809 17 -1809 0 cellNo=895
rlabel pdiffusion 24 -1809 24 -1809 0 cellNo=801
rlabel pdiffusion 31 -1809 31 -1809 0 cellNo=764
rlabel pdiffusion 38 -1809 38 -1809 0 cellNo=517
rlabel pdiffusion 45 -1809 45 -1809 0 cellNo=588
rlabel pdiffusion 52 -1809 52 -1809 0 cellNo=595
rlabel pdiffusion 59 -1809 59 -1809 0 cellNo=889
rlabel pdiffusion 157 -1809 157 -1809 0 cellNo=886
rlabel pdiffusion 185 -1809 185 -1809 0 cellNo=878
rlabel pdiffusion 192 -1809 192 -1809 0 feedthrough
rlabel pdiffusion 206 -1809 206 -1809 0 cellNo=284
rlabel pdiffusion 220 -1809 220 -1809 0 cellNo=494
rlabel pdiffusion 227 -1809 227 -1809 0 feedthrough
rlabel pdiffusion 262 -1809 262 -1809 0 cellNo=900
rlabel pdiffusion 269 -1809 269 -1809 0 feedthrough
rlabel pdiffusion 283 -1809 283 -1809 0 cellNo=418
rlabel pdiffusion 297 -1809 297 -1809 0 feedthrough
rlabel pdiffusion 304 -1809 304 -1809 0 cellNo=770
rlabel pdiffusion 325 -1809 325 -1809 0 cellNo=703
rlabel pdiffusion 332 -1809 332 -1809 0 feedthrough
rlabel pdiffusion 339 -1809 339 -1809 0 cellNo=609
rlabel pdiffusion 353 -1809 353 -1809 0 feedthrough
rlabel pdiffusion 360 -1809 360 -1809 0 cellNo=697
rlabel pdiffusion 374 -1809 374 -1809 0 cellNo=351
rlabel pdiffusion 381 -1809 381 -1809 0 cellNo=892
rlabel pdiffusion 388 -1809 388 -1809 0 feedthrough
rlabel pdiffusion 423 -1809 423 -1809 0 feedthrough
rlabel pdiffusion 430 -1809 430 -1809 0 cellNo=308
rlabel pdiffusion 465 -1809 465 -1809 0 cellNo=894
rlabel pdiffusion 472 -1809 472 -1809 0 cellNo=669
rlabel pdiffusion 479 -1809 479 -1809 0 cellNo=888
rlabel pdiffusion 514 -1809 514 -1809 0 cellNo=880
rlabel pdiffusion 745 -1809 745 -1809 0 cellNo=577
rlabel pdiffusion 752 -1809 752 -1809 0 feedthrough
rlabel pdiffusion 794 -1809 794 -1809 0 cellNo=891
rlabel pdiffusion 899 -1809 899 -1809 0 cellNo=898
rlabel pdiffusion 906 -1809 906 -1809 0 feedthrough
rlabel pdiffusion 1025 -1809 1025 -1809 0 cellNo=885
rlabel polysilicon 177 -4 177 -4 0 1
rlabel polysilicon 177 -10 177 -10 0 3
rlabel polysilicon 184 -4 184 -4 0 1
rlabel polysilicon 184 -10 184 -10 0 3
rlabel polysilicon 194 -4 194 -4 0 2
rlabel polysilicon 198 -4 198 -4 0 1
rlabel polysilicon 212 -4 212 -4 0 1
rlabel polysilicon 219 -4 219 -4 0 1
rlabel polysilicon 219 -10 219 -10 0 3
rlabel polysilicon 236 -4 236 -4 0 2
rlabel polysilicon 240 -4 240 -4 0 1
rlabel polysilicon 240 -10 240 -10 0 3
rlabel polysilicon 254 -4 254 -4 0 1
rlabel polysilicon 261 -4 261 -4 0 1
rlabel polysilicon 261 -10 261 -10 0 3
rlabel polysilicon 278 -10 278 -10 0 4
rlabel polysilicon 285 -4 285 -4 0 2
rlabel polysilicon 289 -4 289 -4 0 1
rlabel polysilicon 289 -10 289 -10 0 3
rlabel polysilicon 296 -10 296 -10 0 3
rlabel polysilicon 303 -4 303 -4 0 1
rlabel polysilicon 303 -10 303 -10 0 3
rlabel polysilicon 310 -4 310 -4 0 1
rlabel polysilicon 317 -10 317 -10 0 3
rlabel polysilicon 338 -4 338 -4 0 1
rlabel polysilicon 338 -10 338 -10 0 3
rlabel polysilicon 348 -4 348 -4 0 2
rlabel polysilicon 352 -4 352 -4 0 1
rlabel polysilicon 352 -10 352 -10 0 3
rlabel polysilicon 359 -4 359 -4 0 1
rlabel polysilicon 366 -4 366 -4 0 1
rlabel polysilicon 366 -10 366 -10 0 3
rlabel polysilicon 408 -4 408 -4 0 1
rlabel polysilicon 408 -10 408 -10 0 3
rlabel polysilicon 422 -10 422 -10 0 3
rlabel polysilicon 460 -10 460 -10 0 4
rlabel polysilicon 467 -4 467 -4 0 2
rlabel polysilicon 471 -4 471 -4 0 1
rlabel polysilicon 471 -10 471 -10 0 3
rlabel polysilicon 478 -4 478 -4 0 1
rlabel polysilicon 485 -4 485 -4 0 1
rlabel polysilicon 485 -10 485 -10 0 3
rlabel polysilicon 534 -4 534 -4 0 1
rlabel polysilicon 541 -4 541 -4 0 1
rlabel polysilicon 541 -10 541 -10 0 3
rlabel polysilicon 555 -10 555 -10 0 3
rlabel polysilicon 558 -10 558 -10 0 4
rlabel polysilicon 576 -4 576 -4 0 1
rlabel polysilicon 583 -4 583 -4 0 1
rlabel polysilicon 583 -10 583 -10 0 3
rlabel polysilicon 604 -4 604 -4 0 1
rlabel polysilicon 604 -10 604 -10 0 3
rlabel polysilicon 611 -4 611 -4 0 1
rlabel polysilicon 621 -10 621 -10 0 4
rlabel polysilicon 730 -4 730 -4 0 1
rlabel polysilicon 730 -10 730 -10 0 3
rlabel polysilicon 740 -4 740 -4 0 2
rlabel polysilicon 61 -27 61 -27 0 4
rlabel polysilicon 79 -27 79 -27 0 3
rlabel polysilicon 114 -21 114 -21 0 1
rlabel polysilicon 121 -21 121 -21 0 1
rlabel polysilicon 121 -27 121 -27 0 3
rlabel polysilicon 128 -27 128 -27 0 3
rlabel polysilicon 156 -21 156 -21 0 1
rlabel polysilicon 163 -21 163 -21 0 1
rlabel polysilicon 163 -27 163 -27 0 3
rlabel polysilicon 170 -21 170 -21 0 1
rlabel polysilicon 170 -27 170 -27 0 3
rlabel polysilicon 180 -27 180 -27 0 4
rlabel polysilicon 184 -21 184 -21 0 1
rlabel polysilicon 184 -27 184 -27 0 3
rlabel polysilicon 215 -21 215 -21 0 2
rlabel polysilicon 219 -21 219 -21 0 1
rlabel polysilicon 219 -27 219 -27 0 3
rlabel polysilicon 226 -21 226 -21 0 1
rlabel polysilicon 226 -27 226 -27 0 3
rlabel polysilicon 240 -21 240 -21 0 1
rlabel polysilicon 240 -27 240 -27 0 3
rlabel polysilicon 247 -21 247 -21 0 1
rlabel polysilicon 247 -27 247 -27 0 3
rlabel polysilicon 254 -21 254 -21 0 1
rlabel polysilicon 254 -27 254 -27 0 3
rlabel polysilicon 261 -21 261 -21 0 1
rlabel polysilicon 271 -27 271 -27 0 4
rlabel polysilicon 278 -21 278 -21 0 2
rlabel polysilicon 282 -21 282 -21 0 1
rlabel polysilicon 282 -27 282 -27 0 3
rlabel polysilicon 289 -21 289 -21 0 1
rlabel polysilicon 289 -27 289 -27 0 3
rlabel polysilicon 296 -21 296 -21 0 1
rlabel polysilicon 296 -27 296 -27 0 3
rlabel polysilicon 303 -21 303 -21 0 1
rlabel polysilicon 303 -27 303 -27 0 3
rlabel polysilicon 310 -21 310 -21 0 1
rlabel polysilicon 310 -27 310 -27 0 3
rlabel polysilicon 317 -21 317 -21 0 1
rlabel polysilicon 317 -27 317 -27 0 3
rlabel polysilicon 334 -21 334 -21 0 2
rlabel polysilicon 338 -21 338 -21 0 1
rlabel polysilicon 338 -27 338 -27 0 3
rlabel polysilicon 345 -21 345 -21 0 1
rlabel polysilicon 345 -27 345 -27 0 3
rlabel polysilicon 352 -21 352 -21 0 1
rlabel polysilicon 352 -27 352 -27 0 3
rlabel polysilicon 359 -21 359 -21 0 1
rlabel polysilicon 359 -27 359 -27 0 3
rlabel polysilicon 366 -21 366 -21 0 1
rlabel polysilicon 366 -27 366 -27 0 3
rlabel polysilicon 373 -21 373 -21 0 1
rlabel polysilicon 380 -27 380 -27 0 3
rlabel polysilicon 411 -27 411 -27 0 4
rlabel polysilicon 415 -21 415 -21 0 1
rlabel polysilicon 415 -27 415 -27 0 3
rlabel polysilicon 425 -21 425 -21 0 2
rlabel polysilicon 429 -21 429 -21 0 1
rlabel polysilicon 429 -27 429 -27 0 3
rlabel polysilicon 436 -27 436 -27 0 3
rlabel polysilicon 443 -21 443 -21 0 1
rlabel polysilicon 443 -27 443 -27 0 3
rlabel polysilicon 450 -21 450 -21 0 1
rlabel polysilicon 450 -27 450 -27 0 3
rlabel polysilicon 457 -21 457 -21 0 1
rlabel polysilicon 457 -27 457 -27 0 3
rlabel polysilicon 467 -21 467 -21 0 2
rlabel polysilicon 474 -21 474 -21 0 2
rlabel polysilicon 478 -21 478 -21 0 1
rlabel polysilicon 478 -27 478 -27 0 3
rlabel polysilicon 485 -21 485 -21 0 1
rlabel polysilicon 485 -27 485 -27 0 3
rlabel polysilicon 492 -21 492 -21 0 1
rlabel polysilicon 492 -27 492 -27 0 3
rlabel polysilicon 527 -21 527 -21 0 1
rlabel polysilicon 527 -27 527 -27 0 3
rlabel polysilicon 541 -21 541 -21 0 1
rlabel polysilicon 541 -27 541 -27 0 3
rlabel polysilicon 579 -27 579 -27 0 4
rlabel polysilicon 583 -21 583 -21 0 1
rlabel polysilicon 583 -27 583 -27 0 3
rlabel polysilicon 604 -21 604 -21 0 1
rlabel polysilicon 604 -27 604 -27 0 3
rlabel polysilicon 611 -21 611 -21 0 1
rlabel polysilicon 611 -27 611 -27 0 3
rlabel polysilicon 618 -21 618 -21 0 1
rlabel polysilicon 618 -27 618 -27 0 3
rlabel polysilicon 688 -21 688 -21 0 1
rlabel polysilicon 688 -27 688 -27 0 3
rlabel polysilicon 698 -21 698 -21 0 2
rlabel polysilicon 709 -27 709 -27 0 3
rlabel polysilicon 712 -27 712 -27 0 4
rlabel polysilicon 730 -21 730 -21 0 1
rlabel polysilicon 730 -27 730 -27 0 3
rlabel polysilicon 58 -44 58 -44 0 1
rlabel polysilicon 58 -50 58 -50 0 3
rlabel polysilicon 65 -50 65 -50 0 3
rlabel polysilicon 79 -44 79 -44 0 1
rlabel polysilicon 79 -50 79 -50 0 3
rlabel polysilicon 107 -50 107 -50 0 3
rlabel polysilicon 114 -44 114 -44 0 1
rlabel polysilicon 114 -50 114 -50 0 3
rlabel polysilicon 124 -44 124 -44 0 2
rlabel polysilicon 121 -50 121 -50 0 3
rlabel polysilicon 128 -44 128 -44 0 1
rlabel polysilicon 131 -50 131 -50 0 4
rlabel polysilicon 135 -44 135 -44 0 1
rlabel polysilicon 135 -50 135 -50 0 3
rlabel polysilicon 142 -44 142 -44 0 1
rlabel polysilicon 142 -50 142 -50 0 3
rlabel polysilicon 152 -44 152 -44 0 2
rlabel polysilicon 156 -44 156 -44 0 1
rlabel polysilicon 156 -50 156 -50 0 3
rlabel polysilicon 163 -44 163 -44 0 1
rlabel polysilicon 163 -50 163 -50 0 3
rlabel polysilicon 170 -44 170 -44 0 1
rlabel polysilicon 173 -44 173 -44 0 2
rlabel polysilicon 170 -50 170 -50 0 3
rlabel polysilicon 177 -44 177 -44 0 1
rlabel polysilicon 177 -50 177 -50 0 3
rlabel polysilicon 184 -44 184 -44 0 1
rlabel polysilicon 184 -50 184 -50 0 3
rlabel polysilicon 191 -50 191 -50 0 3
rlabel polysilicon 198 -44 198 -44 0 1
rlabel polysilicon 198 -50 198 -50 0 3
rlabel polysilicon 208 -50 208 -50 0 4
rlabel polysilicon 212 -44 212 -44 0 1
rlabel polysilicon 212 -50 212 -50 0 3
rlabel polysilicon 222 -50 222 -50 0 4
rlabel polysilicon 226 -44 226 -44 0 1
rlabel polysilicon 226 -50 226 -50 0 3
rlabel polysilicon 229 -50 229 -50 0 4
rlabel polysilicon 233 -44 233 -44 0 1
rlabel polysilicon 233 -50 233 -50 0 3
rlabel polysilicon 240 -44 240 -44 0 1
rlabel polysilicon 240 -50 240 -50 0 3
rlabel polysilicon 247 -44 247 -44 0 1
rlabel polysilicon 247 -50 247 -50 0 3
rlabel polysilicon 254 -44 254 -44 0 1
rlabel polysilicon 257 -44 257 -44 0 2
rlabel polysilicon 261 -44 261 -44 0 1
rlabel polysilicon 261 -50 261 -50 0 3
rlabel polysilicon 268 -44 268 -44 0 1
rlabel polysilicon 268 -50 268 -50 0 3
rlabel polysilicon 275 -44 275 -44 0 1
rlabel polysilicon 275 -50 275 -50 0 3
rlabel polysilicon 282 -44 282 -44 0 1
rlabel polysilicon 282 -50 282 -50 0 3
rlabel polysilicon 289 -44 289 -44 0 1
rlabel polysilicon 289 -50 289 -50 0 3
rlabel polysilicon 296 -44 296 -44 0 1
rlabel polysilicon 296 -50 296 -50 0 3
rlabel polysilicon 303 -44 303 -44 0 1
rlabel polysilicon 303 -50 303 -50 0 3
rlabel polysilicon 310 -44 310 -44 0 1
rlabel polysilicon 310 -50 310 -50 0 3
rlabel polysilicon 317 -44 317 -44 0 1
rlabel polysilicon 317 -50 317 -50 0 3
rlabel polysilicon 324 -44 324 -44 0 1
rlabel polysilicon 324 -50 324 -50 0 3
rlabel polysilicon 331 -44 331 -44 0 1
rlabel polysilicon 334 -44 334 -44 0 2
rlabel polysilicon 338 -44 338 -44 0 1
rlabel polysilicon 345 -44 345 -44 0 1
rlabel polysilicon 345 -50 345 -50 0 3
rlabel polysilicon 352 -44 352 -44 0 1
rlabel polysilicon 352 -50 352 -50 0 3
rlabel polysilicon 359 -44 359 -44 0 1
rlabel polysilicon 359 -50 359 -50 0 3
rlabel polysilicon 366 -44 366 -44 0 1
rlabel polysilicon 366 -50 366 -50 0 3
rlabel polysilicon 373 -44 373 -44 0 1
rlabel polysilicon 373 -50 373 -50 0 3
rlabel polysilicon 380 -44 380 -44 0 1
rlabel polysilicon 380 -50 380 -50 0 3
rlabel polysilicon 387 -44 387 -44 0 1
rlabel polysilicon 397 -44 397 -44 0 2
rlabel polysilicon 394 -50 394 -50 0 3
rlabel polysilicon 401 -44 401 -44 0 1
rlabel polysilicon 401 -50 401 -50 0 3
rlabel polysilicon 408 -44 408 -44 0 1
rlabel polysilicon 408 -50 408 -50 0 3
rlabel polysilicon 425 -44 425 -44 0 2
rlabel polysilicon 422 -50 422 -50 0 3
rlabel polysilicon 429 -44 429 -44 0 1
rlabel polysilicon 429 -50 429 -50 0 3
rlabel polysilicon 436 -44 436 -44 0 1
rlabel polysilicon 436 -50 436 -50 0 3
rlabel polysilicon 443 -50 443 -50 0 3
rlabel polysilicon 446 -50 446 -50 0 4
rlabel polysilicon 450 -44 450 -44 0 1
rlabel polysilicon 450 -50 450 -50 0 3
rlabel polysilicon 457 -44 457 -44 0 1
rlabel polysilicon 457 -50 457 -50 0 3
rlabel polysilicon 471 -44 471 -44 0 1
rlabel polysilicon 471 -50 471 -50 0 3
rlabel polysilicon 478 -44 478 -44 0 1
rlabel polysilicon 478 -50 478 -50 0 3
rlabel polysilicon 485 -44 485 -44 0 1
rlabel polysilicon 485 -50 485 -50 0 3
rlabel polysilicon 499 -44 499 -44 0 1
rlabel polysilicon 499 -50 499 -50 0 3
rlabel polysilicon 513 -44 513 -44 0 1
rlabel polysilicon 513 -50 513 -50 0 3
rlabel polysilicon 537 -44 537 -44 0 2
rlabel polysilicon 534 -50 534 -50 0 3
rlabel polysilicon 541 -44 541 -44 0 1
rlabel polysilicon 548 -44 548 -44 0 1
rlabel polysilicon 548 -50 548 -50 0 3
rlabel polysilicon 555 -44 555 -44 0 1
rlabel polysilicon 555 -50 555 -50 0 3
rlabel polysilicon 562 -44 562 -44 0 1
rlabel polysilicon 562 -50 562 -50 0 3
rlabel polysilicon 572 -44 572 -44 0 2
rlabel polysilicon 576 -44 576 -44 0 1
rlabel polysilicon 576 -50 576 -50 0 3
rlabel polysilicon 583 -44 583 -44 0 1
rlabel polysilicon 583 -50 583 -50 0 3
rlabel polysilicon 590 -50 590 -50 0 3
rlabel polysilicon 597 -44 597 -44 0 1
rlabel polysilicon 597 -50 597 -50 0 3
rlabel polysilicon 604 -44 604 -44 0 1
rlabel polysilicon 604 -50 604 -50 0 3
rlabel polysilicon 611 -44 611 -44 0 1
rlabel polysilicon 611 -50 611 -50 0 3
rlabel polysilicon 625 -44 625 -44 0 1
rlabel polysilicon 625 -50 625 -50 0 3
rlabel polysilicon 632 -44 632 -44 0 1
rlabel polysilicon 632 -50 632 -50 0 3
rlabel polysilicon 646 -44 646 -44 0 1
rlabel polysilicon 653 -50 653 -50 0 3
rlabel polysilicon 660 -44 660 -44 0 1
rlabel polysilicon 660 -50 660 -50 0 3
rlabel polysilicon 688 -44 688 -44 0 1
rlabel polysilicon 688 -50 688 -50 0 3
rlabel polysilicon 730 -44 730 -44 0 1
rlabel polysilicon 730 -50 730 -50 0 3
rlabel polysilicon 786 -44 786 -44 0 1
rlabel polysilicon 786 -50 786 -50 0 3
rlabel polysilicon 807 -44 807 -44 0 1
rlabel polysilicon 807 -50 807 -50 0 3
rlabel polysilicon 814 -44 814 -44 0 1
rlabel polysilicon 898 -50 898 -50 0 3
rlabel polysilicon 54 -89 54 -89 0 4
rlabel polysilicon 58 -83 58 -83 0 1
rlabel polysilicon 58 -89 58 -89 0 3
rlabel polysilicon 65 -83 65 -83 0 1
rlabel polysilicon 65 -89 65 -89 0 3
rlabel polysilicon 79 -83 79 -83 0 1
rlabel polysilicon 89 -89 89 -89 0 4
rlabel polysilicon 93 -83 93 -83 0 1
rlabel polysilicon 93 -89 93 -89 0 3
rlabel polysilicon 103 -83 103 -83 0 2
rlabel polysilicon 110 -83 110 -83 0 2
rlabel polysilicon 114 -83 114 -83 0 1
rlabel polysilicon 114 -89 114 -89 0 3
rlabel polysilicon 124 -89 124 -89 0 4
rlabel polysilicon 128 -83 128 -83 0 1
rlabel polysilicon 128 -89 128 -89 0 3
rlabel polysilicon 135 -83 135 -83 0 1
rlabel polysilicon 135 -89 135 -89 0 3
rlabel polysilicon 142 -83 142 -83 0 1
rlabel polysilicon 142 -89 142 -89 0 3
rlabel polysilicon 149 -83 149 -83 0 1
rlabel polysilicon 149 -89 149 -89 0 3
rlabel polysilicon 156 -83 156 -83 0 1
rlabel polysilicon 156 -89 156 -89 0 3
rlabel polysilicon 163 -83 163 -83 0 1
rlabel polysilicon 163 -89 163 -89 0 3
rlabel polysilicon 170 -83 170 -83 0 1
rlabel polysilicon 170 -89 170 -89 0 3
rlabel polysilicon 180 -89 180 -89 0 4
rlabel polysilicon 184 -83 184 -83 0 1
rlabel polysilicon 184 -89 184 -89 0 3
rlabel polysilicon 187 -89 187 -89 0 4
rlabel polysilicon 191 -83 191 -83 0 1
rlabel polysilicon 191 -89 191 -89 0 3
rlabel polysilicon 198 -83 198 -83 0 1
rlabel polysilicon 198 -89 198 -89 0 3
rlabel polysilicon 205 -83 205 -83 0 1
rlabel polysilicon 208 -83 208 -83 0 2
rlabel polysilicon 205 -89 205 -89 0 3
rlabel polysilicon 212 -83 212 -83 0 1
rlabel polysilicon 212 -89 212 -89 0 3
rlabel polysilicon 222 -89 222 -89 0 4
rlabel polysilicon 229 -89 229 -89 0 4
rlabel polysilicon 233 -83 233 -83 0 1
rlabel polysilicon 233 -89 233 -89 0 3
rlabel polysilicon 240 -83 240 -83 0 1
rlabel polysilicon 240 -89 240 -89 0 3
rlabel polysilicon 247 -83 247 -83 0 1
rlabel polysilicon 247 -89 247 -89 0 3
rlabel polysilicon 254 -83 254 -83 0 1
rlabel polysilicon 254 -89 254 -89 0 3
rlabel polysilicon 261 -83 261 -83 0 1
rlabel polysilicon 261 -89 261 -89 0 3
rlabel polysilicon 268 -83 268 -83 0 1
rlabel polysilicon 268 -89 268 -89 0 3
rlabel polysilicon 278 -83 278 -83 0 2
rlabel polysilicon 282 -83 282 -83 0 1
rlabel polysilicon 282 -89 282 -89 0 3
rlabel polysilicon 289 -83 289 -83 0 1
rlabel polysilicon 289 -89 289 -89 0 3
rlabel polysilicon 299 -83 299 -83 0 2
rlabel polysilicon 299 -89 299 -89 0 4
rlabel polysilicon 303 -83 303 -83 0 1
rlabel polysilicon 303 -89 303 -89 0 3
rlabel polysilicon 310 -83 310 -83 0 1
rlabel polysilicon 317 -83 317 -83 0 1
rlabel polysilicon 317 -89 317 -89 0 3
rlabel polysilicon 324 -83 324 -83 0 1
rlabel polysilicon 324 -89 324 -89 0 3
rlabel polysilicon 331 -83 331 -83 0 1
rlabel polysilicon 331 -89 331 -89 0 3
rlabel polysilicon 338 -83 338 -83 0 1
rlabel polysilicon 338 -89 338 -89 0 3
rlabel polysilicon 345 -83 345 -83 0 1
rlabel polysilicon 345 -89 345 -89 0 3
rlabel polysilicon 352 -83 352 -83 0 1
rlabel polysilicon 352 -89 352 -89 0 3
rlabel polysilicon 359 -89 359 -89 0 3
rlabel polysilicon 362 -89 362 -89 0 4
rlabel polysilicon 366 -83 366 -83 0 1
rlabel polysilicon 366 -89 366 -89 0 3
rlabel polysilicon 373 -83 373 -83 0 1
rlabel polysilicon 373 -89 373 -89 0 3
rlabel polysilicon 380 -83 380 -83 0 1
rlabel polysilicon 380 -89 380 -89 0 3
rlabel polysilicon 387 -83 387 -83 0 1
rlabel polysilicon 387 -89 387 -89 0 3
rlabel polysilicon 390 -89 390 -89 0 4
rlabel polysilicon 394 -83 394 -83 0 1
rlabel polysilicon 397 -89 397 -89 0 4
rlabel polysilicon 401 -83 401 -83 0 1
rlabel polysilicon 401 -89 401 -89 0 3
rlabel polysilicon 408 -83 408 -83 0 1
rlabel polysilicon 408 -89 408 -89 0 3
rlabel polysilicon 415 -83 415 -83 0 1
rlabel polysilicon 415 -89 415 -89 0 3
rlabel polysilicon 422 -83 422 -83 0 1
rlabel polysilicon 422 -89 422 -89 0 3
rlabel polysilicon 429 -83 429 -83 0 1
rlabel polysilicon 429 -89 429 -89 0 3
rlabel polysilicon 439 -83 439 -83 0 2
rlabel polysilicon 436 -89 436 -89 0 3
rlabel polysilicon 443 -83 443 -83 0 1
rlabel polysilicon 446 -83 446 -83 0 2
rlabel polysilicon 450 -83 450 -83 0 1
rlabel polysilicon 450 -89 450 -89 0 3
rlabel polysilicon 460 -83 460 -83 0 2
rlabel polysilicon 467 -83 467 -83 0 2
rlabel polysilicon 474 -83 474 -83 0 2
rlabel polysilicon 478 -83 478 -83 0 1
rlabel polysilicon 478 -89 478 -89 0 3
rlabel polysilicon 485 -83 485 -83 0 1
rlabel polysilicon 485 -89 485 -89 0 3
rlabel polysilicon 495 -83 495 -83 0 2
rlabel polysilicon 495 -89 495 -89 0 4
rlabel polysilicon 499 -83 499 -83 0 1
rlabel polysilicon 499 -89 499 -89 0 3
rlabel polysilicon 506 -83 506 -83 0 1
rlabel polysilicon 506 -89 506 -89 0 3
rlabel polysilicon 513 -83 513 -83 0 1
rlabel polysilicon 513 -89 513 -89 0 3
rlabel polysilicon 520 -83 520 -83 0 1
rlabel polysilicon 520 -89 520 -89 0 3
rlabel polysilicon 527 -83 527 -83 0 1
rlabel polysilicon 534 -83 534 -83 0 1
rlabel polysilicon 534 -89 534 -89 0 3
rlabel polysilicon 541 -83 541 -83 0 1
rlabel polysilicon 541 -89 541 -89 0 3
rlabel polysilicon 548 -83 548 -83 0 1
rlabel polysilicon 548 -89 548 -89 0 3
rlabel polysilicon 555 -83 555 -83 0 1
rlabel polysilicon 555 -89 555 -89 0 3
rlabel polysilicon 562 -83 562 -83 0 1
rlabel polysilicon 562 -89 562 -89 0 3
rlabel polysilicon 569 -83 569 -83 0 1
rlabel polysilicon 569 -89 569 -89 0 3
rlabel polysilicon 576 -83 576 -83 0 1
rlabel polysilicon 576 -89 576 -89 0 3
rlabel polysilicon 583 -83 583 -83 0 1
rlabel polysilicon 583 -89 583 -89 0 3
rlabel polysilicon 590 -83 590 -83 0 1
rlabel polysilicon 590 -89 590 -89 0 3
rlabel polysilicon 597 -83 597 -83 0 1
rlabel polysilicon 597 -89 597 -89 0 3
rlabel polysilicon 604 -83 604 -83 0 1
rlabel polysilicon 604 -89 604 -89 0 3
rlabel polysilicon 611 -83 611 -83 0 1
rlabel polysilicon 611 -89 611 -89 0 3
rlabel polysilicon 618 -83 618 -83 0 1
rlabel polysilicon 618 -89 618 -89 0 3
rlabel polysilicon 625 -83 625 -83 0 1
rlabel polysilicon 625 -89 625 -89 0 3
rlabel polysilicon 632 -83 632 -83 0 1
rlabel polysilicon 639 -83 639 -83 0 1
rlabel polysilicon 639 -89 639 -89 0 3
rlabel polysilicon 646 -83 646 -83 0 1
rlabel polysilicon 646 -89 646 -89 0 3
rlabel polysilicon 653 -83 653 -83 0 1
rlabel polysilicon 653 -89 653 -89 0 3
rlabel polysilicon 660 -83 660 -83 0 1
rlabel polysilicon 660 -89 660 -89 0 3
rlabel polysilicon 674 -83 674 -83 0 1
rlabel polysilicon 674 -89 674 -89 0 3
rlabel polysilicon 681 -89 681 -89 0 3
rlabel polysilicon 702 -83 702 -83 0 1
rlabel polysilicon 702 -89 702 -89 0 3
rlabel polysilicon 730 -83 730 -83 0 1
rlabel polysilicon 730 -89 730 -89 0 3
rlabel polysilicon 793 -83 793 -83 0 1
rlabel polysilicon 793 -89 793 -89 0 3
rlabel polysilicon 807 -83 807 -83 0 1
rlabel polysilicon 807 -89 807 -89 0 3
rlabel polysilicon 898 -83 898 -83 0 1
rlabel polysilicon 898 -89 898 -89 0 3
rlabel polysilicon 978 -89 978 -89 0 4
rlabel polysilicon 1087 -83 1087 -83 0 1
rlabel polysilicon 1087 -89 1087 -89 0 3
rlabel polysilicon 1097 -83 1097 -83 0 2
rlabel polysilicon 30 -120 30 -120 0 1
rlabel polysilicon 30 -126 30 -126 0 3
rlabel polysilicon 44 -120 44 -120 0 1
rlabel polysilicon 47 -126 47 -126 0 4
rlabel polysilicon 51 -120 51 -120 0 1
rlabel polysilicon 51 -126 51 -126 0 3
rlabel polysilicon 58 -120 58 -120 0 1
rlabel polysilicon 58 -126 58 -126 0 3
rlabel polysilicon 65 -120 65 -120 0 1
rlabel polysilicon 65 -126 65 -126 0 3
rlabel polysilicon 93 -120 93 -120 0 1
rlabel polysilicon 93 -126 93 -126 0 3
rlabel polysilicon 100 -120 100 -120 0 1
rlabel polysilicon 100 -126 100 -126 0 3
rlabel polysilicon 107 -120 107 -120 0 1
rlabel polysilicon 107 -126 107 -126 0 3
rlabel polysilicon 114 -120 114 -120 0 1
rlabel polysilicon 121 -120 121 -120 0 1
rlabel polysilicon 121 -126 121 -126 0 3
rlabel polysilicon 128 -120 128 -120 0 1
rlabel polysilicon 128 -126 128 -126 0 3
rlabel polysilicon 135 -126 135 -126 0 3
rlabel polysilicon 138 -126 138 -126 0 4
rlabel polysilicon 142 -120 142 -120 0 1
rlabel polysilicon 142 -126 142 -126 0 3
rlabel polysilicon 149 -120 149 -120 0 1
rlabel polysilicon 149 -126 149 -126 0 3
rlabel polysilicon 156 -120 156 -120 0 1
rlabel polysilicon 156 -126 156 -126 0 3
rlabel polysilicon 163 -120 163 -120 0 1
rlabel polysilicon 163 -126 163 -126 0 3
rlabel polysilicon 170 -120 170 -120 0 1
rlabel polysilicon 170 -126 170 -126 0 3
rlabel polysilicon 177 -120 177 -120 0 1
rlabel polysilicon 180 -120 180 -120 0 2
rlabel polysilicon 177 -126 177 -126 0 3
rlabel polysilicon 187 -126 187 -126 0 4
rlabel polysilicon 191 -120 191 -120 0 1
rlabel polysilicon 191 -126 191 -126 0 3
rlabel polysilicon 198 -120 198 -120 0 1
rlabel polysilicon 198 -126 198 -126 0 3
rlabel polysilicon 205 -120 205 -120 0 1
rlabel polysilicon 205 -126 205 -126 0 3
rlabel polysilicon 212 -120 212 -120 0 1
rlabel polysilicon 212 -126 212 -126 0 3
rlabel polysilicon 219 -120 219 -120 0 1
rlabel polysilicon 219 -126 219 -126 0 3
rlabel polysilicon 229 -120 229 -120 0 2
rlabel polysilicon 229 -126 229 -126 0 4
rlabel polysilicon 233 -120 233 -120 0 1
rlabel polysilicon 233 -126 233 -126 0 3
rlabel polysilicon 240 -120 240 -120 0 1
rlabel polysilicon 243 -126 243 -126 0 4
rlabel polysilicon 247 -126 247 -126 0 3
rlabel polysilicon 250 -126 250 -126 0 4
rlabel polysilicon 254 -120 254 -120 0 1
rlabel polysilicon 254 -126 254 -126 0 3
rlabel polysilicon 261 -120 261 -120 0 1
rlabel polysilicon 261 -126 261 -126 0 3
rlabel polysilicon 268 -120 268 -120 0 1
rlabel polysilicon 268 -126 268 -126 0 3
rlabel polysilicon 275 -120 275 -120 0 1
rlabel polysilicon 275 -126 275 -126 0 3
rlabel polysilicon 282 -120 282 -120 0 1
rlabel polysilicon 282 -126 282 -126 0 3
rlabel polysilicon 289 -120 289 -120 0 1
rlabel polysilicon 289 -126 289 -126 0 3
rlabel polysilicon 299 -120 299 -120 0 2
rlabel polysilicon 303 -120 303 -120 0 1
rlabel polysilicon 303 -126 303 -126 0 3
rlabel polysilicon 310 -126 310 -126 0 3
rlabel polysilicon 317 -120 317 -120 0 1
rlabel polysilicon 317 -126 317 -126 0 3
rlabel polysilicon 324 -120 324 -120 0 1
rlabel polysilicon 327 -120 327 -120 0 2
rlabel polysilicon 324 -126 324 -126 0 3
rlabel polysilicon 331 -120 331 -120 0 1
rlabel polysilicon 331 -126 331 -126 0 3
rlabel polysilicon 338 -120 338 -120 0 1
rlabel polysilicon 338 -126 338 -126 0 3
rlabel polysilicon 345 -120 345 -120 0 1
rlabel polysilicon 345 -126 345 -126 0 3
rlabel polysilicon 355 -120 355 -120 0 2
rlabel polysilicon 352 -126 352 -126 0 3
rlabel polysilicon 359 -120 359 -120 0 1
rlabel polysilicon 359 -126 359 -126 0 3
rlabel polysilicon 366 -120 366 -120 0 1
rlabel polysilicon 366 -126 366 -126 0 3
rlabel polysilicon 373 -120 373 -120 0 1
rlabel polysilicon 376 -126 376 -126 0 4
rlabel polysilicon 380 -126 380 -126 0 3
rlabel polysilicon 383 -126 383 -126 0 4
rlabel polysilicon 387 -120 387 -120 0 1
rlabel polysilicon 390 -120 390 -120 0 2
rlabel polysilicon 387 -126 387 -126 0 3
rlabel polysilicon 394 -120 394 -120 0 1
rlabel polysilicon 394 -126 394 -126 0 3
rlabel polysilicon 401 -120 401 -120 0 1
rlabel polysilicon 401 -126 401 -126 0 3
rlabel polysilicon 408 -120 408 -120 0 1
rlabel polysilicon 411 -120 411 -120 0 2
rlabel polysilicon 415 -120 415 -120 0 1
rlabel polysilicon 415 -126 415 -126 0 3
rlabel polysilicon 422 -120 422 -120 0 1
rlabel polysilicon 422 -126 422 -126 0 3
rlabel polysilicon 429 -120 429 -120 0 1
rlabel polysilicon 429 -126 429 -126 0 3
rlabel polysilicon 436 -120 436 -120 0 1
rlabel polysilicon 436 -126 436 -126 0 3
rlabel polysilicon 443 -120 443 -120 0 1
rlabel polysilicon 443 -126 443 -126 0 3
rlabel polysilicon 450 -120 450 -120 0 1
rlabel polysilicon 450 -126 450 -126 0 3
rlabel polysilicon 457 -120 457 -120 0 1
rlabel polysilicon 457 -126 457 -126 0 3
rlabel polysilicon 467 -120 467 -120 0 2
rlabel polysilicon 464 -126 464 -126 0 3
rlabel polysilicon 471 -120 471 -120 0 1
rlabel polysilicon 471 -126 471 -126 0 3
rlabel polysilicon 478 -126 478 -126 0 3
rlabel polysilicon 481 -126 481 -126 0 4
rlabel polysilicon 485 -120 485 -120 0 1
rlabel polysilicon 485 -126 485 -126 0 3
rlabel polysilicon 492 -120 492 -120 0 1
rlabel polysilicon 492 -126 492 -126 0 3
rlabel polysilicon 499 -120 499 -120 0 1
rlabel polysilicon 499 -126 499 -126 0 3
rlabel polysilicon 509 -126 509 -126 0 4
rlabel polysilicon 513 -120 513 -120 0 1
rlabel polysilicon 513 -126 513 -126 0 3
rlabel polysilicon 520 -120 520 -120 0 1
rlabel polysilicon 520 -126 520 -126 0 3
rlabel polysilicon 527 -120 527 -120 0 1
rlabel polysilicon 527 -126 527 -126 0 3
rlabel polysilicon 534 -120 534 -120 0 1
rlabel polysilicon 534 -126 534 -126 0 3
rlabel polysilicon 541 -120 541 -120 0 1
rlabel polysilicon 541 -126 541 -126 0 3
rlabel polysilicon 548 -126 548 -126 0 3
rlabel polysilicon 555 -126 555 -126 0 3
rlabel polysilicon 562 -120 562 -120 0 1
rlabel polysilicon 562 -126 562 -126 0 3
rlabel polysilicon 569 -120 569 -120 0 1
rlabel polysilicon 569 -126 569 -126 0 3
rlabel polysilicon 576 -120 576 -120 0 1
rlabel polysilicon 576 -126 576 -126 0 3
rlabel polysilicon 583 -120 583 -120 0 1
rlabel polysilicon 583 -126 583 -126 0 3
rlabel polysilicon 593 -120 593 -120 0 2
rlabel polysilicon 593 -126 593 -126 0 4
rlabel polysilicon 597 -120 597 -120 0 1
rlabel polysilicon 597 -126 597 -126 0 3
rlabel polysilicon 604 -120 604 -120 0 1
rlabel polysilicon 604 -126 604 -126 0 3
rlabel polysilicon 611 -120 611 -120 0 1
rlabel polysilicon 611 -126 611 -126 0 3
rlabel polysilicon 618 -120 618 -120 0 1
rlabel polysilicon 618 -126 618 -126 0 3
rlabel polysilicon 625 -120 625 -120 0 1
rlabel polysilicon 625 -126 625 -126 0 3
rlabel polysilicon 632 -120 632 -120 0 1
rlabel polysilicon 632 -126 632 -126 0 3
rlabel polysilicon 639 -120 639 -120 0 1
rlabel polysilicon 639 -126 639 -126 0 3
rlabel polysilicon 646 -120 646 -120 0 1
rlabel polysilicon 646 -126 646 -126 0 3
rlabel polysilicon 656 -126 656 -126 0 4
rlabel polysilicon 660 -120 660 -120 0 1
rlabel polysilicon 660 -126 660 -126 0 3
rlabel polysilicon 667 -120 667 -120 0 1
rlabel polysilicon 667 -126 667 -126 0 3
rlabel polysilicon 674 -120 674 -120 0 1
rlabel polysilicon 674 -126 674 -126 0 3
rlabel polysilicon 681 -120 681 -120 0 1
rlabel polysilicon 681 -126 681 -126 0 3
rlabel polysilicon 688 -120 688 -120 0 1
rlabel polysilicon 688 -126 688 -126 0 3
rlabel polysilicon 695 -120 695 -120 0 1
rlabel polysilicon 695 -126 695 -126 0 3
rlabel polysilicon 702 -120 702 -120 0 1
rlabel polysilicon 702 -126 702 -126 0 3
rlabel polysilicon 709 -126 709 -126 0 3
rlabel polysilicon 716 -120 716 -120 0 1
rlabel polysilicon 716 -126 716 -126 0 3
rlabel polysilicon 723 -120 723 -120 0 1
rlabel polysilicon 723 -126 723 -126 0 3
rlabel polysilicon 730 -120 730 -120 0 1
rlabel polysilicon 730 -126 730 -126 0 3
rlabel polysilicon 737 -120 737 -120 0 1
rlabel polysilicon 737 -126 737 -126 0 3
rlabel polysilicon 758 -120 758 -120 0 1
rlabel polysilicon 765 -120 765 -120 0 1
rlabel polysilicon 765 -126 765 -126 0 3
rlabel polysilicon 779 -120 779 -120 0 1
rlabel polysilicon 779 -126 779 -126 0 3
rlabel polysilicon 800 -120 800 -120 0 1
rlabel polysilicon 800 -126 800 -126 0 3
rlabel polysilicon 905 -120 905 -120 0 1
rlabel polysilicon 905 -126 905 -126 0 3
rlabel polysilicon 975 -120 975 -120 0 1
rlabel polysilicon 975 -126 975 -126 0 3
rlabel polysilicon 1087 -120 1087 -120 0 1
rlabel polysilicon 1087 -126 1087 -126 0 3
rlabel polysilicon 23 -181 23 -181 0 1
rlabel polysilicon 23 -187 23 -187 0 3
rlabel polysilicon 30 -181 30 -181 0 1
rlabel polysilicon 30 -187 30 -187 0 3
rlabel polysilicon 37 -181 37 -181 0 1
rlabel polysilicon 44 -181 44 -181 0 1
rlabel polysilicon 51 -181 51 -181 0 1
rlabel polysilicon 51 -187 51 -187 0 3
rlabel polysilicon 58 -181 58 -181 0 1
rlabel polysilicon 58 -187 58 -187 0 3
rlabel polysilicon 65 -187 65 -187 0 3
rlabel polysilicon 68 -187 68 -187 0 4
rlabel polysilicon 72 -181 72 -181 0 1
rlabel polysilicon 72 -187 72 -187 0 3
rlabel polysilicon 79 -181 79 -181 0 1
rlabel polysilicon 79 -187 79 -187 0 3
rlabel polysilicon 86 -181 86 -181 0 1
rlabel polysilicon 93 -181 93 -181 0 1
rlabel polysilicon 93 -187 93 -187 0 3
rlabel polysilicon 100 -181 100 -181 0 1
rlabel polysilicon 100 -187 100 -187 0 3
rlabel polysilicon 107 -181 107 -181 0 1
rlabel polysilicon 107 -187 107 -187 0 3
rlabel polysilicon 114 -181 114 -181 0 1
rlabel polysilicon 114 -187 114 -187 0 3
rlabel polysilicon 121 -181 121 -181 0 1
rlabel polysilicon 121 -187 121 -187 0 3
rlabel polysilicon 128 -181 128 -181 0 1
rlabel polysilicon 128 -187 128 -187 0 3
rlabel polysilicon 138 -181 138 -181 0 2
rlabel polysilicon 142 -181 142 -181 0 1
rlabel polysilicon 142 -187 142 -187 0 3
rlabel polysilicon 149 -181 149 -181 0 1
rlabel polysilicon 149 -187 149 -187 0 3
rlabel polysilicon 156 -181 156 -181 0 1
rlabel polysilicon 156 -187 156 -187 0 3
rlabel polysilicon 166 -181 166 -181 0 2
rlabel polysilicon 170 -181 170 -181 0 1
rlabel polysilicon 170 -187 170 -187 0 3
rlabel polysilicon 177 -181 177 -181 0 1
rlabel polysilicon 177 -187 177 -187 0 3
rlabel polysilicon 184 -181 184 -181 0 1
rlabel polysilicon 187 -187 187 -187 0 4
rlabel polysilicon 191 -181 191 -181 0 1
rlabel polysilicon 191 -187 191 -187 0 3
rlabel polysilicon 198 -187 198 -187 0 3
rlabel polysilicon 201 -187 201 -187 0 4
rlabel polysilicon 205 -181 205 -181 0 1
rlabel polysilicon 212 -181 212 -181 0 1
rlabel polysilicon 212 -187 212 -187 0 3
rlabel polysilicon 219 -181 219 -181 0 1
rlabel polysilicon 219 -187 219 -187 0 3
rlabel polysilicon 226 -181 226 -181 0 1
rlabel polysilicon 226 -187 226 -187 0 3
rlabel polysilicon 233 -181 233 -181 0 1
rlabel polysilicon 233 -187 233 -187 0 3
rlabel polysilicon 240 -181 240 -181 0 1
rlabel polysilicon 240 -187 240 -187 0 3
rlabel polysilicon 247 -181 247 -181 0 1
rlabel polysilicon 247 -187 247 -187 0 3
rlabel polysilicon 254 -181 254 -181 0 1
rlabel polysilicon 254 -187 254 -187 0 3
rlabel polysilicon 261 -181 261 -181 0 1
rlabel polysilicon 261 -187 261 -187 0 3
rlabel polysilicon 268 -181 268 -181 0 1
rlabel polysilicon 268 -187 268 -187 0 3
rlabel polysilicon 275 -181 275 -181 0 1
rlabel polysilicon 275 -187 275 -187 0 3
rlabel polysilicon 282 -181 282 -181 0 1
rlabel polysilicon 282 -187 282 -187 0 3
rlabel polysilicon 289 -181 289 -181 0 1
rlabel polysilicon 289 -187 289 -187 0 3
rlabel polysilicon 296 -181 296 -181 0 1
rlabel polysilicon 296 -187 296 -187 0 3
rlabel polysilicon 303 -181 303 -181 0 1
rlabel polysilicon 303 -187 303 -187 0 3
rlabel polysilicon 310 -181 310 -181 0 1
rlabel polysilicon 310 -187 310 -187 0 3
rlabel polysilicon 317 -181 317 -181 0 1
rlabel polysilicon 320 -181 320 -181 0 2
rlabel polysilicon 317 -187 317 -187 0 3
rlabel polysilicon 324 -181 324 -181 0 1
rlabel polysilicon 324 -187 324 -187 0 3
rlabel polysilicon 331 -181 331 -181 0 1
rlabel polysilicon 334 -181 334 -181 0 2
rlabel polysilicon 338 -181 338 -181 0 1
rlabel polysilicon 345 -181 345 -181 0 1
rlabel polysilicon 348 -181 348 -181 0 2
rlabel polysilicon 345 -187 345 -187 0 3
rlabel polysilicon 348 -187 348 -187 0 4
rlabel polysilicon 352 -181 352 -181 0 1
rlabel polysilicon 352 -187 352 -187 0 3
rlabel polysilicon 359 -181 359 -181 0 1
rlabel polysilicon 359 -187 359 -187 0 3
rlabel polysilicon 366 -181 366 -181 0 1
rlabel polysilicon 366 -187 366 -187 0 3
rlabel polysilicon 376 -181 376 -181 0 2
rlabel polysilicon 373 -187 373 -187 0 3
rlabel polysilicon 380 -181 380 -181 0 1
rlabel polysilicon 380 -187 380 -187 0 3
rlabel polysilicon 387 -181 387 -181 0 1
rlabel polysilicon 390 -181 390 -181 0 2
rlabel polysilicon 394 -181 394 -181 0 1
rlabel polysilicon 394 -187 394 -187 0 3
rlabel polysilicon 401 -181 401 -181 0 1
rlabel polysilicon 401 -187 401 -187 0 3
rlabel polysilicon 408 -181 408 -181 0 1
rlabel polysilicon 408 -187 408 -187 0 3
rlabel polysilicon 415 -181 415 -181 0 1
rlabel polysilicon 415 -187 415 -187 0 3
rlabel polysilicon 422 -181 422 -181 0 1
rlabel polysilicon 422 -187 422 -187 0 3
rlabel polysilicon 425 -187 425 -187 0 4
rlabel polysilicon 429 -181 429 -181 0 1
rlabel polysilicon 429 -187 429 -187 0 3
rlabel polysilicon 436 -181 436 -181 0 1
rlabel polysilicon 436 -187 436 -187 0 3
rlabel polysilicon 443 -181 443 -181 0 1
rlabel polysilicon 443 -187 443 -187 0 3
rlabel polysilicon 450 -181 450 -181 0 1
rlabel polysilicon 450 -187 450 -187 0 3
rlabel polysilicon 457 -181 457 -181 0 1
rlabel polysilicon 457 -187 457 -187 0 3
rlabel polysilicon 467 -181 467 -181 0 2
rlabel polysilicon 467 -187 467 -187 0 4
rlabel polysilicon 471 -181 471 -181 0 1
rlabel polysilicon 471 -187 471 -187 0 3
rlabel polysilicon 478 -181 478 -181 0 1
rlabel polysilicon 478 -187 478 -187 0 3
rlabel polysilicon 488 -181 488 -181 0 2
rlabel polysilicon 485 -187 485 -187 0 3
rlabel polysilicon 495 -181 495 -181 0 2
rlabel polysilicon 499 -181 499 -181 0 1
rlabel polysilicon 499 -187 499 -187 0 3
rlabel polysilicon 506 -181 506 -181 0 1
rlabel polysilicon 506 -187 506 -187 0 3
rlabel polysilicon 513 -181 513 -181 0 1
rlabel polysilicon 513 -187 513 -187 0 3
rlabel polysilicon 523 -181 523 -181 0 2
rlabel polysilicon 527 -181 527 -181 0 1
rlabel polysilicon 527 -187 527 -187 0 3
rlabel polysilicon 537 -181 537 -181 0 2
rlabel polysilicon 537 -187 537 -187 0 4
rlabel polysilicon 541 -181 541 -181 0 1
rlabel polysilicon 541 -187 541 -187 0 3
rlabel polysilicon 548 -181 548 -181 0 1
rlabel polysilicon 548 -187 548 -187 0 3
rlabel polysilicon 555 -181 555 -181 0 1
rlabel polysilicon 555 -187 555 -187 0 3
rlabel polysilicon 562 -181 562 -181 0 1
rlabel polysilicon 562 -187 562 -187 0 3
rlabel polysilicon 569 -181 569 -181 0 1
rlabel polysilicon 569 -187 569 -187 0 3
rlabel polysilicon 576 -181 576 -181 0 1
rlabel polysilicon 576 -187 576 -187 0 3
rlabel polysilicon 583 -181 583 -181 0 1
rlabel polysilicon 583 -187 583 -187 0 3
rlabel polysilicon 590 -181 590 -181 0 1
rlabel polysilicon 590 -187 590 -187 0 3
rlabel polysilicon 597 -181 597 -181 0 1
rlabel polysilicon 597 -187 597 -187 0 3
rlabel polysilicon 604 -181 604 -181 0 1
rlabel polysilicon 604 -187 604 -187 0 3
rlabel polysilicon 611 -181 611 -181 0 1
rlabel polysilicon 611 -187 611 -187 0 3
rlabel polysilicon 618 -181 618 -181 0 1
rlabel polysilicon 618 -187 618 -187 0 3
rlabel polysilicon 625 -181 625 -181 0 1
rlabel polysilicon 625 -187 625 -187 0 3
rlabel polysilicon 632 -181 632 -181 0 1
rlabel polysilicon 632 -187 632 -187 0 3
rlabel polysilicon 639 -181 639 -181 0 1
rlabel polysilicon 639 -187 639 -187 0 3
rlabel polysilicon 646 -181 646 -181 0 1
rlabel polysilicon 646 -187 646 -187 0 3
rlabel polysilicon 653 -181 653 -181 0 1
rlabel polysilicon 653 -187 653 -187 0 3
rlabel polysilicon 660 -181 660 -181 0 1
rlabel polysilicon 660 -187 660 -187 0 3
rlabel polysilicon 667 -181 667 -181 0 1
rlabel polysilicon 667 -187 667 -187 0 3
rlabel polysilicon 674 -181 674 -181 0 1
rlabel polysilicon 674 -187 674 -187 0 3
rlabel polysilicon 681 -181 681 -181 0 1
rlabel polysilicon 681 -187 681 -187 0 3
rlabel polysilicon 688 -181 688 -181 0 1
rlabel polysilicon 688 -187 688 -187 0 3
rlabel polysilicon 695 -181 695 -181 0 1
rlabel polysilicon 695 -187 695 -187 0 3
rlabel polysilicon 702 -181 702 -181 0 1
rlabel polysilicon 702 -187 702 -187 0 3
rlabel polysilicon 709 -181 709 -181 0 1
rlabel polysilicon 709 -187 709 -187 0 3
rlabel polysilicon 716 -181 716 -181 0 1
rlabel polysilicon 716 -187 716 -187 0 3
rlabel polysilicon 723 -181 723 -181 0 1
rlabel polysilicon 723 -187 723 -187 0 3
rlabel polysilicon 730 -181 730 -181 0 1
rlabel polysilicon 730 -187 730 -187 0 3
rlabel polysilicon 737 -181 737 -181 0 1
rlabel polysilicon 737 -187 737 -187 0 3
rlabel polysilicon 744 -181 744 -181 0 1
rlabel polysilicon 744 -187 744 -187 0 3
rlabel polysilicon 751 -181 751 -181 0 1
rlabel polysilicon 751 -187 751 -187 0 3
rlabel polysilicon 758 -181 758 -181 0 1
rlabel polysilicon 758 -187 758 -187 0 3
rlabel polysilicon 765 -181 765 -181 0 1
rlabel polysilicon 765 -187 765 -187 0 3
rlabel polysilicon 772 -181 772 -181 0 1
rlabel polysilicon 772 -187 772 -187 0 3
rlabel polysilicon 779 -181 779 -181 0 1
rlabel polysilicon 779 -187 779 -187 0 3
rlabel polysilicon 786 -181 786 -181 0 1
rlabel polysilicon 786 -187 786 -187 0 3
rlabel polysilicon 793 -181 793 -181 0 1
rlabel polysilicon 793 -187 793 -187 0 3
rlabel polysilicon 800 -181 800 -181 0 1
rlabel polysilicon 800 -187 800 -187 0 3
rlabel polysilicon 807 -181 807 -181 0 1
rlabel polysilicon 807 -187 807 -187 0 3
rlabel polysilicon 814 -181 814 -181 0 1
rlabel polysilicon 821 -187 821 -187 0 3
rlabel polysilicon 828 -187 828 -187 0 3
rlabel polysilicon 835 -187 835 -187 0 3
rlabel polysilicon 845 -181 845 -181 0 2
rlabel polysilicon 849 -181 849 -181 0 1
rlabel polysilicon 849 -187 849 -187 0 3
rlabel polysilicon 859 -187 859 -187 0 4
rlabel polysilicon 919 -181 919 -181 0 1
rlabel polysilicon 919 -187 919 -187 0 3
rlabel polysilicon 975 -181 975 -181 0 1
rlabel polysilicon 975 -187 975 -187 0 3
rlabel polysilicon 1087 -181 1087 -181 0 1
rlabel polysilicon 1087 -187 1087 -187 0 3
rlabel polysilicon 16 -240 16 -240 0 1
rlabel polysilicon 16 -246 16 -246 0 3
rlabel polysilicon 23 -240 23 -240 0 1
rlabel polysilicon 23 -246 23 -246 0 3
rlabel polysilicon 30 -240 30 -240 0 1
rlabel polysilicon 30 -246 30 -246 0 3
rlabel polysilicon 37 -240 37 -240 0 1
rlabel polysilicon 37 -246 37 -246 0 3
rlabel polysilicon 44 -240 44 -240 0 1
rlabel polysilicon 44 -246 44 -246 0 3
rlabel polysilicon 51 -240 51 -240 0 1
rlabel polysilicon 51 -246 51 -246 0 3
rlabel polysilicon 58 -240 58 -240 0 1
rlabel polysilicon 65 -240 65 -240 0 1
rlabel polysilicon 68 -240 68 -240 0 2
rlabel polysilicon 72 -240 72 -240 0 1
rlabel polysilicon 72 -246 72 -246 0 3
rlabel polysilicon 79 -240 79 -240 0 1
rlabel polysilicon 79 -246 79 -246 0 3
rlabel polysilicon 89 -246 89 -246 0 4
rlabel polysilicon 93 -240 93 -240 0 1
rlabel polysilicon 93 -246 93 -246 0 3
rlabel polysilicon 100 -240 100 -240 0 1
rlabel polysilicon 103 -240 103 -240 0 2
rlabel polysilicon 103 -246 103 -246 0 4
rlabel polysilicon 107 -240 107 -240 0 1
rlabel polysilicon 107 -246 107 -246 0 3
rlabel polysilicon 114 -240 114 -240 0 1
rlabel polysilicon 117 -240 117 -240 0 2
rlabel polysilicon 114 -246 114 -246 0 3
rlabel polysilicon 117 -246 117 -246 0 4
rlabel polysilicon 121 -240 121 -240 0 1
rlabel polysilicon 121 -246 121 -246 0 3
rlabel polysilicon 128 -240 128 -240 0 1
rlabel polysilicon 128 -246 128 -246 0 3
rlabel polysilicon 135 -240 135 -240 0 1
rlabel polysilicon 135 -246 135 -246 0 3
rlabel polysilicon 142 -240 142 -240 0 1
rlabel polysilicon 142 -246 142 -246 0 3
rlabel polysilicon 149 -240 149 -240 0 1
rlabel polysilicon 149 -246 149 -246 0 3
rlabel polysilicon 156 -246 156 -246 0 3
rlabel polysilicon 159 -246 159 -246 0 4
rlabel polysilicon 163 -240 163 -240 0 1
rlabel polysilicon 163 -246 163 -246 0 3
rlabel polysilicon 173 -240 173 -240 0 2
rlabel polysilicon 170 -246 170 -246 0 3
rlabel polysilicon 177 -240 177 -240 0 1
rlabel polysilicon 177 -246 177 -246 0 3
rlabel polysilicon 184 -240 184 -240 0 1
rlabel polysilicon 187 -240 187 -240 0 2
rlabel polysilicon 191 -240 191 -240 0 1
rlabel polysilicon 191 -246 191 -246 0 3
rlabel polysilicon 201 -240 201 -240 0 2
rlabel polysilicon 205 -240 205 -240 0 1
rlabel polysilicon 205 -246 205 -246 0 3
rlabel polysilicon 212 -240 212 -240 0 1
rlabel polysilicon 212 -246 212 -246 0 3
rlabel polysilicon 219 -246 219 -246 0 3
rlabel polysilicon 229 -240 229 -240 0 2
rlabel polysilicon 226 -246 226 -246 0 3
rlabel polysilicon 233 -240 233 -240 0 1
rlabel polysilicon 233 -246 233 -246 0 3
rlabel polysilicon 240 -240 240 -240 0 1
rlabel polysilicon 240 -246 240 -246 0 3
rlabel polysilicon 247 -240 247 -240 0 1
rlabel polysilicon 247 -246 247 -246 0 3
rlabel polysilicon 254 -240 254 -240 0 1
rlabel polysilicon 254 -246 254 -246 0 3
rlabel polysilicon 261 -246 261 -246 0 3
rlabel polysilicon 264 -246 264 -246 0 4
rlabel polysilicon 268 -240 268 -240 0 1
rlabel polysilicon 268 -246 268 -246 0 3
rlabel polysilicon 275 -240 275 -240 0 1
rlabel polysilicon 275 -246 275 -246 0 3
rlabel polysilicon 282 -240 282 -240 0 1
rlabel polysilicon 292 -240 292 -240 0 2
rlabel polysilicon 292 -246 292 -246 0 4
rlabel polysilicon 296 -240 296 -240 0 1
rlabel polysilicon 296 -246 296 -246 0 3
rlabel polysilicon 303 -240 303 -240 0 1
rlabel polysilicon 303 -246 303 -246 0 3
rlabel polysilicon 310 -240 310 -240 0 1
rlabel polysilicon 310 -246 310 -246 0 3
rlabel polysilicon 317 -240 317 -240 0 1
rlabel polysilicon 317 -246 317 -246 0 3
rlabel polysilicon 324 -240 324 -240 0 1
rlabel polysilicon 324 -246 324 -246 0 3
rlabel polysilicon 331 -240 331 -240 0 1
rlabel polysilicon 331 -246 331 -246 0 3
rlabel polysilicon 338 -240 338 -240 0 1
rlabel polysilicon 338 -246 338 -246 0 3
rlabel polysilicon 345 -240 345 -240 0 1
rlabel polysilicon 345 -246 345 -246 0 3
rlabel polysilicon 352 -240 352 -240 0 1
rlabel polysilicon 355 -240 355 -240 0 2
rlabel polysilicon 359 -240 359 -240 0 1
rlabel polysilicon 359 -246 359 -246 0 3
rlabel polysilicon 366 -240 366 -240 0 1
rlabel polysilicon 366 -246 366 -246 0 3
rlabel polysilicon 373 -240 373 -240 0 1
rlabel polysilicon 373 -246 373 -246 0 3
rlabel polysilicon 380 -246 380 -246 0 3
rlabel polysilicon 383 -246 383 -246 0 4
rlabel polysilicon 387 -240 387 -240 0 1
rlabel polysilicon 387 -246 387 -246 0 3
rlabel polysilicon 394 -240 394 -240 0 1
rlabel polysilicon 394 -246 394 -246 0 3
rlabel polysilicon 401 -240 401 -240 0 1
rlabel polysilicon 401 -246 401 -246 0 3
rlabel polysilicon 408 -240 408 -240 0 1
rlabel polysilicon 408 -246 408 -246 0 3
rlabel polysilicon 415 -240 415 -240 0 1
rlabel polysilicon 415 -246 415 -246 0 3
rlabel polysilicon 422 -240 422 -240 0 1
rlabel polysilicon 422 -246 422 -246 0 3
rlabel polysilicon 429 -240 429 -240 0 1
rlabel polysilicon 429 -246 429 -246 0 3
rlabel polysilicon 436 -240 436 -240 0 1
rlabel polysilicon 436 -246 436 -246 0 3
rlabel polysilicon 443 -240 443 -240 0 1
rlabel polysilicon 443 -246 443 -246 0 3
rlabel polysilicon 450 -240 450 -240 0 1
rlabel polysilicon 450 -246 450 -246 0 3
rlabel polysilicon 460 -240 460 -240 0 2
rlabel polysilicon 457 -246 457 -246 0 3
rlabel polysilicon 464 -240 464 -240 0 1
rlabel polysilicon 467 -240 467 -240 0 2
rlabel polysilicon 464 -246 464 -246 0 3
rlabel polysilicon 471 -240 471 -240 0 1
rlabel polysilicon 471 -246 471 -246 0 3
rlabel polysilicon 478 -240 478 -240 0 1
rlabel polysilicon 478 -246 478 -246 0 3
rlabel polysilicon 481 -246 481 -246 0 4
rlabel polysilicon 485 -246 485 -246 0 3
rlabel polysilicon 495 -240 495 -240 0 2
rlabel polysilicon 492 -246 492 -246 0 3
rlabel polysilicon 495 -246 495 -246 0 4
rlabel polysilicon 499 -240 499 -240 0 1
rlabel polysilicon 499 -246 499 -246 0 3
rlabel polysilicon 506 -240 506 -240 0 1
rlabel polysilicon 506 -246 506 -246 0 3
rlabel polysilicon 513 -240 513 -240 0 1
rlabel polysilicon 513 -246 513 -246 0 3
rlabel polysilicon 520 -240 520 -240 0 1
rlabel polysilicon 520 -246 520 -246 0 3
rlabel polysilicon 527 -240 527 -240 0 1
rlabel polysilicon 527 -246 527 -246 0 3
rlabel polysilicon 534 -240 534 -240 0 1
rlabel polysilicon 534 -246 534 -246 0 3
rlabel polysilicon 541 -240 541 -240 0 1
rlabel polysilicon 541 -246 541 -246 0 3
rlabel polysilicon 548 -240 548 -240 0 1
rlabel polysilicon 548 -246 548 -246 0 3
rlabel polysilicon 555 -240 555 -240 0 1
rlabel polysilicon 555 -246 555 -246 0 3
rlabel polysilicon 562 -240 562 -240 0 1
rlabel polysilicon 562 -246 562 -246 0 3
rlabel polysilicon 569 -240 569 -240 0 1
rlabel polysilicon 569 -246 569 -246 0 3
rlabel polysilicon 576 -240 576 -240 0 1
rlabel polysilicon 576 -246 576 -246 0 3
rlabel polysilicon 583 -240 583 -240 0 1
rlabel polysilicon 583 -246 583 -246 0 3
rlabel polysilicon 593 -240 593 -240 0 2
rlabel polysilicon 593 -246 593 -246 0 4
rlabel polysilicon 597 -246 597 -246 0 3
rlabel polysilicon 600 -246 600 -246 0 4
rlabel polysilicon 604 -240 604 -240 0 1
rlabel polysilicon 604 -246 604 -246 0 3
rlabel polysilicon 611 -240 611 -240 0 1
rlabel polysilicon 611 -246 611 -246 0 3
rlabel polysilicon 618 -240 618 -240 0 1
rlabel polysilicon 618 -246 618 -246 0 3
rlabel polysilicon 625 -240 625 -240 0 1
rlabel polysilicon 625 -246 625 -246 0 3
rlabel polysilicon 632 -240 632 -240 0 1
rlabel polysilicon 632 -246 632 -246 0 3
rlabel polysilicon 639 -240 639 -240 0 1
rlabel polysilicon 639 -246 639 -246 0 3
rlabel polysilicon 646 -246 646 -246 0 3
rlabel polysilicon 653 -240 653 -240 0 1
rlabel polysilicon 653 -246 653 -246 0 3
rlabel polysilicon 660 -240 660 -240 0 1
rlabel polysilicon 660 -246 660 -246 0 3
rlabel polysilicon 667 -240 667 -240 0 1
rlabel polysilicon 667 -246 667 -246 0 3
rlabel polysilicon 674 -240 674 -240 0 1
rlabel polysilicon 674 -246 674 -246 0 3
rlabel polysilicon 681 -240 681 -240 0 1
rlabel polysilicon 681 -246 681 -246 0 3
rlabel polysilicon 688 -240 688 -240 0 1
rlabel polysilicon 688 -246 688 -246 0 3
rlabel polysilicon 695 -240 695 -240 0 1
rlabel polysilicon 695 -246 695 -246 0 3
rlabel polysilicon 702 -240 702 -240 0 1
rlabel polysilicon 702 -246 702 -246 0 3
rlabel polysilicon 709 -240 709 -240 0 1
rlabel polysilicon 709 -246 709 -246 0 3
rlabel polysilicon 716 -240 716 -240 0 1
rlabel polysilicon 716 -246 716 -246 0 3
rlabel polysilicon 723 -240 723 -240 0 1
rlabel polysilicon 723 -246 723 -246 0 3
rlabel polysilicon 730 -240 730 -240 0 1
rlabel polysilicon 730 -246 730 -246 0 3
rlabel polysilicon 737 -240 737 -240 0 1
rlabel polysilicon 737 -246 737 -246 0 3
rlabel polysilicon 744 -240 744 -240 0 1
rlabel polysilicon 744 -246 744 -246 0 3
rlabel polysilicon 751 -240 751 -240 0 1
rlabel polysilicon 751 -246 751 -246 0 3
rlabel polysilicon 758 -240 758 -240 0 1
rlabel polysilicon 758 -246 758 -246 0 3
rlabel polysilicon 765 -240 765 -240 0 1
rlabel polysilicon 765 -246 765 -246 0 3
rlabel polysilicon 772 -240 772 -240 0 1
rlabel polysilicon 772 -246 772 -246 0 3
rlabel polysilicon 779 -240 779 -240 0 1
rlabel polysilicon 779 -246 779 -246 0 3
rlabel polysilicon 786 -240 786 -240 0 1
rlabel polysilicon 786 -246 786 -246 0 3
rlabel polysilicon 793 -240 793 -240 0 1
rlabel polysilicon 793 -246 793 -246 0 3
rlabel polysilicon 800 -240 800 -240 0 1
rlabel polysilicon 807 -240 807 -240 0 1
rlabel polysilicon 807 -246 807 -246 0 3
rlabel polysilicon 814 -240 814 -240 0 1
rlabel polysilicon 814 -246 814 -246 0 3
rlabel polysilicon 821 -240 821 -240 0 1
rlabel polysilicon 821 -246 821 -246 0 3
rlabel polysilicon 828 -240 828 -240 0 1
rlabel polysilicon 828 -246 828 -246 0 3
rlabel polysilicon 835 -240 835 -240 0 1
rlabel polysilicon 835 -246 835 -246 0 3
rlabel polysilicon 842 -240 842 -240 0 1
rlabel polysilicon 842 -246 842 -246 0 3
rlabel polysilicon 849 -240 849 -240 0 1
rlabel polysilicon 849 -246 849 -246 0 3
rlabel polysilicon 856 -240 856 -240 0 1
rlabel polysilicon 856 -246 856 -246 0 3
rlabel polysilicon 863 -240 863 -240 0 1
rlabel polysilicon 863 -246 863 -246 0 3
rlabel polysilicon 870 -240 870 -240 0 1
rlabel polysilicon 870 -246 870 -246 0 3
rlabel polysilicon 877 -240 877 -240 0 1
rlabel polysilicon 877 -246 877 -246 0 3
rlabel polysilicon 884 -240 884 -240 0 1
rlabel polysilicon 884 -246 884 -246 0 3
rlabel polysilicon 891 -240 891 -240 0 1
rlabel polysilicon 891 -246 891 -246 0 3
rlabel polysilicon 898 -240 898 -240 0 1
rlabel polysilicon 898 -246 898 -246 0 3
rlabel polysilicon 905 -240 905 -240 0 1
rlabel polysilicon 905 -246 905 -246 0 3
rlabel polysilicon 912 -240 912 -240 0 1
rlabel polysilicon 912 -246 912 -246 0 3
rlabel polysilicon 919 -240 919 -240 0 1
rlabel polysilicon 919 -246 919 -246 0 3
rlabel polysilicon 926 -240 926 -240 0 1
rlabel polysilicon 926 -246 926 -246 0 3
rlabel polysilicon 933 -240 933 -240 0 1
rlabel polysilicon 933 -246 933 -246 0 3
rlabel polysilicon 940 -240 940 -240 0 1
rlabel polysilicon 940 -246 940 -246 0 3
rlabel polysilicon 947 -240 947 -240 0 1
rlabel polysilicon 947 -246 947 -246 0 3
rlabel polysilicon 954 -246 954 -246 0 3
rlabel polysilicon 975 -240 975 -240 0 1
rlabel polysilicon 975 -246 975 -246 0 3
rlabel polysilicon 1087 -240 1087 -240 0 1
rlabel polysilicon 1087 -246 1087 -246 0 3
rlabel polysilicon 9 -317 9 -317 0 3
rlabel polysilicon 16 -311 16 -311 0 1
rlabel polysilicon 16 -317 16 -317 0 3
rlabel polysilicon 23 -311 23 -311 0 1
rlabel polysilicon 23 -317 23 -317 0 3
rlabel polysilicon 33 -311 33 -311 0 2
rlabel polysilicon 30 -317 30 -317 0 3
rlabel polysilicon 37 -311 37 -311 0 1
rlabel polysilicon 37 -317 37 -317 0 3
rlabel polysilicon 47 -311 47 -311 0 2
rlabel polysilicon 58 -311 58 -311 0 1
rlabel polysilicon 58 -317 58 -317 0 3
rlabel polysilicon 65 -311 65 -311 0 1
rlabel polysilicon 65 -317 65 -317 0 3
rlabel polysilicon 72 -311 72 -311 0 1
rlabel polysilicon 72 -317 72 -317 0 3
rlabel polysilicon 79 -311 79 -311 0 1
rlabel polysilicon 82 -311 82 -311 0 2
rlabel polysilicon 79 -317 79 -317 0 3
rlabel polysilicon 86 -311 86 -311 0 1
rlabel polysilicon 86 -317 86 -317 0 3
rlabel polysilicon 93 -311 93 -311 0 1
rlabel polysilicon 93 -317 93 -317 0 3
rlabel polysilicon 100 -311 100 -311 0 1
rlabel polysilicon 100 -317 100 -317 0 3
rlabel polysilicon 107 -317 107 -317 0 3
rlabel polysilicon 110 -317 110 -317 0 4
rlabel polysilicon 114 -311 114 -311 0 1
rlabel polysilicon 114 -317 114 -317 0 3
rlabel polysilicon 121 -311 121 -311 0 1
rlabel polysilicon 121 -317 121 -317 0 3
rlabel polysilicon 128 -311 128 -311 0 1
rlabel polysilicon 128 -317 128 -317 0 3
rlabel polysilicon 135 -311 135 -311 0 1
rlabel polysilicon 135 -317 135 -317 0 3
rlabel polysilicon 145 -311 145 -311 0 2
rlabel polysilicon 145 -317 145 -317 0 4
rlabel polysilicon 149 -311 149 -311 0 1
rlabel polysilicon 149 -317 149 -317 0 3
rlabel polysilicon 156 -311 156 -311 0 1
rlabel polysilicon 156 -317 156 -317 0 3
rlabel polysilicon 163 -311 163 -311 0 1
rlabel polysilicon 163 -317 163 -317 0 3
rlabel polysilicon 170 -311 170 -311 0 1
rlabel polysilicon 170 -317 170 -317 0 3
rlabel polysilicon 177 -311 177 -311 0 1
rlabel polysilicon 177 -317 177 -317 0 3
rlabel polysilicon 184 -311 184 -311 0 1
rlabel polysilicon 184 -317 184 -317 0 3
rlabel polysilicon 191 -311 191 -311 0 1
rlabel polysilicon 191 -317 191 -317 0 3
rlabel polysilicon 198 -311 198 -311 0 1
rlabel polysilicon 198 -317 198 -317 0 3
rlabel polysilicon 205 -311 205 -311 0 1
rlabel polysilicon 208 -311 208 -311 0 2
rlabel polysilicon 208 -317 208 -317 0 4
rlabel polysilicon 212 -311 212 -311 0 1
rlabel polysilicon 212 -317 212 -317 0 3
rlabel polysilicon 219 -311 219 -311 0 1
rlabel polysilicon 219 -317 219 -317 0 3
rlabel polysilicon 229 -311 229 -311 0 2
rlabel polysilicon 233 -311 233 -311 0 1
rlabel polysilicon 233 -317 233 -317 0 3
rlabel polysilicon 240 -311 240 -311 0 1
rlabel polysilicon 240 -317 240 -317 0 3
rlabel polysilicon 247 -311 247 -311 0 1
rlabel polysilicon 247 -317 247 -317 0 3
rlabel polysilicon 254 -311 254 -311 0 1
rlabel polysilicon 254 -317 254 -317 0 3
rlabel polysilicon 261 -311 261 -311 0 1
rlabel polysilicon 261 -317 261 -317 0 3
rlabel polysilicon 268 -311 268 -311 0 1
rlabel polysilicon 268 -317 268 -317 0 3
rlabel polysilicon 275 -311 275 -311 0 1
rlabel polysilicon 275 -317 275 -317 0 3
rlabel polysilicon 282 -311 282 -311 0 1
rlabel polysilicon 282 -317 282 -317 0 3
rlabel polysilicon 289 -311 289 -311 0 1
rlabel polysilicon 292 -317 292 -317 0 4
rlabel polysilicon 296 -311 296 -311 0 1
rlabel polysilicon 296 -317 296 -317 0 3
rlabel polysilicon 303 -311 303 -311 0 1
rlabel polysilicon 303 -317 303 -317 0 3
rlabel polysilicon 310 -311 310 -311 0 1
rlabel polysilicon 310 -317 310 -317 0 3
rlabel polysilicon 317 -311 317 -311 0 1
rlabel polysilicon 317 -317 317 -317 0 3
rlabel polysilicon 324 -311 324 -311 0 1
rlabel polysilicon 324 -317 324 -317 0 3
rlabel polysilicon 331 -311 331 -311 0 1
rlabel polysilicon 331 -317 331 -317 0 3
rlabel polysilicon 338 -311 338 -311 0 1
rlabel polysilicon 338 -317 338 -317 0 3
rlabel polysilicon 345 -311 345 -311 0 1
rlabel polysilicon 345 -317 345 -317 0 3
rlabel polysilicon 352 -311 352 -311 0 1
rlabel polysilicon 352 -317 352 -317 0 3
rlabel polysilicon 359 -311 359 -311 0 1
rlabel polysilicon 359 -317 359 -317 0 3
rlabel polysilicon 366 -311 366 -311 0 1
rlabel polysilicon 366 -317 366 -317 0 3
rlabel polysilicon 373 -311 373 -311 0 1
rlabel polysilicon 373 -317 373 -317 0 3
rlabel polysilicon 380 -317 380 -317 0 3
rlabel polysilicon 383 -317 383 -317 0 4
rlabel polysilicon 387 -317 387 -317 0 3
rlabel polysilicon 390 -317 390 -317 0 4
rlabel polysilicon 394 -311 394 -311 0 1
rlabel polysilicon 394 -317 394 -317 0 3
rlabel polysilicon 401 -311 401 -311 0 1
rlabel polysilicon 401 -317 401 -317 0 3
rlabel polysilicon 411 -311 411 -311 0 2
rlabel polysilicon 408 -317 408 -317 0 3
rlabel polysilicon 415 -311 415 -311 0 1
rlabel polysilicon 418 -317 418 -317 0 4
rlabel polysilicon 422 -311 422 -311 0 1
rlabel polysilicon 422 -317 422 -317 0 3
rlabel polysilicon 429 -311 429 -311 0 1
rlabel polysilicon 429 -317 429 -317 0 3
rlabel polysilicon 439 -311 439 -311 0 2
rlabel polysilicon 436 -317 436 -317 0 3
rlabel polysilicon 443 -311 443 -311 0 1
rlabel polysilicon 443 -317 443 -317 0 3
rlabel polysilicon 450 -311 450 -311 0 1
rlabel polysilicon 450 -317 450 -317 0 3
rlabel polysilicon 457 -311 457 -311 0 1
rlabel polysilicon 457 -317 457 -317 0 3
rlabel polysilicon 464 -311 464 -311 0 1
rlabel polysilicon 467 -317 467 -317 0 4
rlabel polysilicon 471 -311 471 -311 0 1
rlabel polysilicon 474 -311 474 -311 0 2
rlabel polysilicon 474 -317 474 -317 0 4
rlabel polysilicon 478 -311 478 -311 0 1
rlabel polysilicon 478 -317 478 -317 0 3
rlabel polysilicon 488 -311 488 -311 0 2
rlabel polysilicon 485 -317 485 -317 0 3
rlabel polysilicon 488 -317 488 -317 0 4
rlabel polysilicon 492 -311 492 -311 0 1
rlabel polysilicon 492 -317 492 -317 0 3
rlabel polysilicon 499 -311 499 -311 0 1
rlabel polysilicon 499 -317 499 -317 0 3
rlabel polysilicon 506 -311 506 -311 0 1
rlabel polysilicon 513 -311 513 -311 0 1
rlabel polysilicon 513 -317 513 -317 0 3
rlabel polysilicon 520 -311 520 -311 0 1
rlabel polysilicon 520 -317 520 -317 0 3
rlabel polysilicon 527 -311 527 -311 0 1
rlabel polysilicon 527 -317 527 -317 0 3
rlabel polysilicon 534 -311 534 -311 0 1
rlabel polysilicon 534 -317 534 -317 0 3
rlabel polysilicon 541 -317 541 -317 0 3
rlabel polysilicon 544 -317 544 -317 0 4
rlabel polysilicon 548 -311 548 -311 0 1
rlabel polysilicon 548 -317 548 -317 0 3
rlabel polysilicon 551 -317 551 -317 0 4
rlabel polysilicon 555 -311 555 -311 0 1
rlabel polysilicon 555 -317 555 -317 0 3
rlabel polysilicon 562 -311 562 -311 0 1
rlabel polysilicon 562 -317 562 -317 0 3
rlabel polysilicon 569 -311 569 -311 0 1
rlabel polysilicon 569 -317 569 -317 0 3
rlabel polysilicon 579 -311 579 -311 0 2
rlabel polysilicon 583 -311 583 -311 0 1
rlabel polysilicon 586 -311 586 -311 0 2
rlabel polysilicon 586 -317 586 -317 0 4
rlabel polysilicon 590 -311 590 -311 0 1
rlabel polysilicon 590 -317 590 -317 0 3
rlabel polysilicon 597 -311 597 -311 0 1
rlabel polysilicon 597 -317 597 -317 0 3
rlabel polysilicon 604 -311 604 -311 0 1
rlabel polysilicon 604 -317 604 -317 0 3
rlabel polysilicon 611 -311 611 -311 0 1
rlabel polysilicon 611 -317 611 -317 0 3
rlabel polysilicon 618 -311 618 -311 0 1
rlabel polysilicon 618 -317 618 -317 0 3
rlabel polysilicon 625 -311 625 -311 0 1
rlabel polysilicon 625 -317 625 -317 0 3
rlabel polysilicon 632 -311 632 -311 0 1
rlabel polysilicon 632 -317 632 -317 0 3
rlabel polysilicon 639 -311 639 -311 0 1
rlabel polysilicon 639 -317 639 -317 0 3
rlabel polysilicon 646 -311 646 -311 0 1
rlabel polysilicon 646 -317 646 -317 0 3
rlabel polysilicon 653 -311 653 -311 0 1
rlabel polysilicon 653 -317 653 -317 0 3
rlabel polysilicon 660 -311 660 -311 0 1
rlabel polysilicon 660 -317 660 -317 0 3
rlabel polysilicon 667 -311 667 -311 0 1
rlabel polysilicon 667 -317 667 -317 0 3
rlabel polysilicon 674 -311 674 -311 0 1
rlabel polysilicon 674 -317 674 -317 0 3
rlabel polysilicon 681 -311 681 -311 0 1
rlabel polysilicon 681 -317 681 -317 0 3
rlabel polysilicon 684 -317 684 -317 0 4
rlabel polysilicon 688 -311 688 -311 0 1
rlabel polysilicon 688 -317 688 -317 0 3
rlabel polysilicon 695 -311 695 -311 0 1
rlabel polysilicon 695 -317 695 -317 0 3
rlabel polysilicon 702 -311 702 -311 0 1
rlabel polysilicon 702 -317 702 -317 0 3
rlabel polysilicon 709 -311 709 -311 0 1
rlabel polysilicon 709 -317 709 -317 0 3
rlabel polysilicon 716 -317 716 -317 0 3
rlabel polysilicon 719 -317 719 -317 0 4
rlabel polysilicon 723 -311 723 -311 0 1
rlabel polysilicon 723 -317 723 -317 0 3
rlabel polysilicon 730 -311 730 -311 0 1
rlabel polysilicon 730 -317 730 -317 0 3
rlabel polysilicon 737 -311 737 -311 0 1
rlabel polysilicon 737 -317 737 -317 0 3
rlabel polysilicon 744 -311 744 -311 0 1
rlabel polysilicon 744 -317 744 -317 0 3
rlabel polysilicon 751 -311 751 -311 0 1
rlabel polysilicon 751 -317 751 -317 0 3
rlabel polysilicon 758 -311 758 -311 0 1
rlabel polysilicon 758 -317 758 -317 0 3
rlabel polysilicon 765 -311 765 -311 0 1
rlabel polysilicon 765 -317 765 -317 0 3
rlabel polysilicon 772 -311 772 -311 0 1
rlabel polysilicon 772 -317 772 -317 0 3
rlabel polysilicon 779 -311 779 -311 0 1
rlabel polysilicon 779 -317 779 -317 0 3
rlabel polysilicon 786 -311 786 -311 0 1
rlabel polysilicon 786 -317 786 -317 0 3
rlabel polysilicon 793 -311 793 -311 0 1
rlabel polysilicon 793 -317 793 -317 0 3
rlabel polysilicon 800 -311 800 -311 0 1
rlabel polysilicon 800 -317 800 -317 0 3
rlabel polysilicon 807 -311 807 -311 0 1
rlabel polysilicon 807 -317 807 -317 0 3
rlabel polysilicon 814 -311 814 -311 0 1
rlabel polysilicon 814 -317 814 -317 0 3
rlabel polysilicon 821 -311 821 -311 0 1
rlabel polysilicon 821 -317 821 -317 0 3
rlabel polysilicon 828 -311 828 -311 0 1
rlabel polysilicon 828 -317 828 -317 0 3
rlabel polysilicon 835 -311 835 -311 0 1
rlabel polysilicon 835 -317 835 -317 0 3
rlabel polysilicon 842 -311 842 -311 0 1
rlabel polysilicon 842 -317 842 -317 0 3
rlabel polysilicon 849 -311 849 -311 0 1
rlabel polysilicon 849 -317 849 -317 0 3
rlabel polysilicon 856 -311 856 -311 0 1
rlabel polysilicon 856 -317 856 -317 0 3
rlabel polysilicon 863 -311 863 -311 0 1
rlabel polysilicon 863 -317 863 -317 0 3
rlabel polysilicon 870 -311 870 -311 0 1
rlabel polysilicon 870 -317 870 -317 0 3
rlabel polysilicon 877 -311 877 -311 0 1
rlabel polysilicon 877 -317 877 -317 0 3
rlabel polysilicon 884 -311 884 -311 0 1
rlabel polysilicon 884 -317 884 -317 0 3
rlabel polysilicon 891 -311 891 -311 0 1
rlabel polysilicon 891 -317 891 -317 0 3
rlabel polysilicon 898 -311 898 -311 0 1
rlabel polysilicon 898 -317 898 -317 0 3
rlabel polysilicon 905 -311 905 -311 0 1
rlabel polysilicon 905 -317 905 -317 0 3
rlabel polysilicon 912 -311 912 -311 0 1
rlabel polysilicon 912 -317 912 -317 0 3
rlabel polysilicon 919 -311 919 -311 0 1
rlabel polysilicon 919 -317 919 -317 0 3
rlabel polysilicon 926 -311 926 -311 0 1
rlabel polysilicon 926 -317 926 -317 0 3
rlabel polysilicon 936 -311 936 -311 0 2
rlabel polysilicon 936 -317 936 -317 0 4
rlabel polysilicon 940 -311 940 -311 0 1
rlabel polysilicon 940 -317 940 -317 0 3
rlabel polysilicon 947 -317 947 -317 0 3
rlabel polysilicon 954 -311 954 -311 0 1
rlabel polysilicon 954 -317 954 -317 0 3
rlabel polysilicon 961 -311 961 -311 0 1
rlabel polysilicon 961 -317 961 -317 0 3
rlabel polysilicon 968 -311 968 -311 0 1
rlabel polysilicon 975 -311 975 -311 0 1
rlabel polysilicon 975 -317 975 -317 0 3
rlabel polysilicon 982 -311 982 -311 0 1
rlabel polysilicon 982 -317 982 -317 0 3
rlabel polysilicon 1094 -311 1094 -311 0 1
rlabel polysilicon 1094 -317 1094 -317 0 3
rlabel polysilicon 16 -396 16 -396 0 1
rlabel polysilicon 16 -402 16 -402 0 3
rlabel polysilicon 23 -396 23 -396 0 1
rlabel polysilicon 23 -402 23 -402 0 3
rlabel polysilicon 33 -396 33 -396 0 2
rlabel polysilicon 40 -396 40 -396 0 2
rlabel polysilicon 44 -396 44 -396 0 1
rlabel polysilicon 44 -402 44 -402 0 3
rlabel polysilicon 51 -396 51 -396 0 1
rlabel polysilicon 51 -402 51 -402 0 3
rlabel polysilicon 58 -396 58 -396 0 1
rlabel polysilicon 58 -402 58 -402 0 3
rlabel polysilicon 65 -396 65 -396 0 1
rlabel polysilicon 65 -402 65 -402 0 3
rlabel polysilicon 72 -396 72 -396 0 1
rlabel polysilicon 72 -402 72 -402 0 3
rlabel polysilicon 79 -396 79 -396 0 1
rlabel polysilicon 79 -402 79 -402 0 3
rlabel polysilicon 86 -396 86 -396 0 1
rlabel polysilicon 86 -402 86 -402 0 3
rlabel polysilicon 93 -396 93 -396 0 1
rlabel polysilicon 93 -402 93 -402 0 3
rlabel polysilicon 100 -396 100 -396 0 1
rlabel polysilicon 100 -402 100 -402 0 3
rlabel polysilicon 107 -396 107 -396 0 1
rlabel polysilicon 107 -402 107 -402 0 3
rlabel polysilicon 117 -396 117 -396 0 2
rlabel polysilicon 114 -402 114 -402 0 3
rlabel polysilicon 121 -396 121 -396 0 1
rlabel polysilicon 121 -402 121 -402 0 3
rlabel polysilicon 128 -396 128 -396 0 1
rlabel polysilicon 128 -402 128 -402 0 3
rlabel polysilicon 135 -396 135 -396 0 1
rlabel polysilicon 138 -402 138 -402 0 4
rlabel polysilicon 145 -396 145 -396 0 2
rlabel polysilicon 142 -402 142 -402 0 3
rlabel polysilicon 145 -402 145 -402 0 4
rlabel polysilicon 149 -396 149 -396 0 1
rlabel polysilicon 149 -402 149 -402 0 3
rlabel polysilicon 156 -396 156 -396 0 1
rlabel polysilicon 156 -402 156 -402 0 3
rlabel polysilicon 163 -396 163 -396 0 1
rlabel polysilicon 163 -402 163 -402 0 3
rlabel polysilicon 170 -402 170 -402 0 3
rlabel polysilicon 173 -402 173 -402 0 4
rlabel polysilicon 180 -396 180 -396 0 2
rlabel polysilicon 177 -402 177 -402 0 3
rlabel polysilicon 180 -402 180 -402 0 4
rlabel polysilicon 184 -396 184 -396 0 1
rlabel polysilicon 184 -402 184 -402 0 3
rlabel polysilicon 191 -396 191 -396 0 1
rlabel polysilicon 191 -402 191 -402 0 3
rlabel polysilicon 198 -396 198 -396 0 1
rlabel polysilicon 198 -402 198 -402 0 3
rlabel polysilicon 205 -396 205 -396 0 1
rlabel polysilicon 208 -396 208 -396 0 2
rlabel polysilicon 208 -402 208 -402 0 4
rlabel polysilicon 212 -396 212 -396 0 1
rlabel polysilicon 212 -402 212 -402 0 3
rlabel polysilicon 219 -396 219 -396 0 1
rlabel polysilicon 219 -402 219 -402 0 3
rlabel polysilicon 226 -396 226 -396 0 1
rlabel polysilicon 226 -402 226 -402 0 3
rlabel polysilicon 233 -396 233 -396 0 1
rlabel polysilicon 233 -402 233 -402 0 3
rlabel polysilicon 240 -396 240 -396 0 1
rlabel polysilicon 240 -402 240 -402 0 3
rlabel polysilicon 247 -396 247 -396 0 1
rlabel polysilicon 247 -402 247 -402 0 3
rlabel polysilicon 254 -396 254 -396 0 1
rlabel polysilicon 254 -402 254 -402 0 3
rlabel polysilicon 261 -396 261 -396 0 1
rlabel polysilicon 268 -396 268 -396 0 1
rlabel polysilicon 268 -402 268 -402 0 3
rlabel polysilicon 275 -396 275 -396 0 1
rlabel polysilicon 278 -402 278 -402 0 4
rlabel polysilicon 282 -396 282 -396 0 1
rlabel polysilicon 282 -402 282 -402 0 3
rlabel polysilicon 285 -402 285 -402 0 4
rlabel polysilicon 289 -396 289 -396 0 1
rlabel polysilicon 289 -402 289 -402 0 3
rlabel polysilicon 296 -396 296 -396 0 1
rlabel polysilicon 296 -402 296 -402 0 3
rlabel polysilicon 303 -396 303 -396 0 1
rlabel polysilicon 303 -402 303 -402 0 3
rlabel polysilicon 310 -396 310 -396 0 1
rlabel polysilicon 310 -402 310 -402 0 3
rlabel polysilicon 317 -402 317 -402 0 3
rlabel polysilicon 320 -402 320 -402 0 4
rlabel polysilicon 324 -396 324 -396 0 1
rlabel polysilicon 324 -402 324 -402 0 3
rlabel polysilicon 331 -396 331 -396 0 1
rlabel polysilicon 331 -402 331 -402 0 3
rlabel polysilicon 338 -396 338 -396 0 1
rlabel polysilicon 338 -402 338 -402 0 3
rlabel polysilicon 341 -402 341 -402 0 4
rlabel polysilicon 345 -396 345 -396 0 1
rlabel polysilicon 345 -402 345 -402 0 3
rlabel polysilicon 352 -396 352 -396 0 1
rlabel polysilicon 352 -402 352 -402 0 3
rlabel polysilicon 359 -396 359 -396 0 1
rlabel polysilicon 366 -396 366 -396 0 1
rlabel polysilicon 366 -402 366 -402 0 3
rlabel polysilicon 373 -396 373 -396 0 1
rlabel polysilicon 373 -402 373 -402 0 3
rlabel polysilicon 380 -396 380 -396 0 1
rlabel polysilicon 380 -402 380 -402 0 3
rlabel polysilicon 387 -396 387 -396 0 1
rlabel polysilicon 387 -402 387 -402 0 3
rlabel polysilicon 394 -396 394 -396 0 1
rlabel polysilicon 394 -402 394 -402 0 3
rlabel polysilicon 401 -396 401 -396 0 1
rlabel polysilicon 404 -396 404 -396 0 2
rlabel polysilicon 404 -402 404 -402 0 4
rlabel polysilicon 408 -396 408 -396 0 1
rlabel polysilicon 408 -402 408 -402 0 3
rlabel polysilicon 415 -396 415 -396 0 1
rlabel polysilicon 415 -402 415 -402 0 3
rlabel polysilicon 422 -396 422 -396 0 1
rlabel polysilicon 425 -402 425 -402 0 4
rlabel polysilicon 429 -396 429 -396 0 1
rlabel polysilicon 429 -402 429 -402 0 3
rlabel polysilicon 436 -396 436 -396 0 1
rlabel polysilicon 436 -402 436 -402 0 3
rlabel polysilicon 443 -396 443 -396 0 1
rlabel polysilicon 443 -402 443 -402 0 3
rlabel polysilicon 450 -396 450 -396 0 1
rlabel polysilicon 453 -396 453 -396 0 2
rlabel polysilicon 457 -396 457 -396 0 1
rlabel polysilicon 457 -402 457 -402 0 3
rlabel polysilicon 464 -396 464 -396 0 1
rlabel polysilicon 464 -402 464 -402 0 3
rlabel polysilicon 474 -396 474 -396 0 2
rlabel polysilicon 478 -396 478 -396 0 1
rlabel polysilicon 478 -402 478 -402 0 3
rlabel polysilicon 485 -396 485 -396 0 1
rlabel polysilicon 485 -402 485 -402 0 3
rlabel polysilicon 492 -396 492 -396 0 1
rlabel polysilicon 495 -396 495 -396 0 2
rlabel polysilicon 492 -402 492 -402 0 3
rlabel polysilicon 499 -396 499 -396 0 1
rlabel polysilicon 499 -402 499 -402 0 3
rlabel polysilicon 506 -396 506 -396 0 1
rlabel polysilicon 513 -396 513 -396 0 1
rlabel polysilicon 513 -402 513 -402 0 3
rlabel polysilicon 520 -396 520 -396 0 1
rlabel polysilicon 523 -396 523 -396 0 2
rlabel polysilicon 520 -402 520 -402 0 3
rlabel polysilicon 527 -396 527 -396 0 1
rlabel polysilicon 527 -402 527 -402 0 3
rlabel polysilicon 534 -396 534 -396 0 1
rlabel polysilicon 534 -402 534 -402 0 3
rlabel polysilicon 541 -396 541 -396 0 1
rlabel polysilicon 541 -402 541 -402 0 3
rlabel polysilicon 548 -396 548 -396 0 1
rlabel polysilicon 551 -396 551 -396 0 2
rlabel polysilicon 551 -402 551 -402 0 4
rlabel polysilicon 555 -396 555 -396 0 1
rlabel polysilicon 555 -402 555 -402 0 3
rlabel polysilicon 562 -396 562 -396 0 1
rlabel polysilicon 565 -396 565 -396 0 2
rlabel polysilicon 569 -396 569 -396 0 1
rlabel polysilicon 569 -402 569 -402 0 3
rlabel polysilicon 579 -396 579 -396 0 2
rlabel polysilicon 579 -402 579 -402 0 4
rlabel polysilicon 583 -396 583 -396 0 1
rlabel polysilicon 583 -402 583 -402 0 3
rlabel polysilicon 590 -396 590 -396 0 1
rlabel polysilicon 590 -402 590 -402 0 3
rlabel polysilicon 597 -396 597 -396 0 1
rlabel polysilicon 597 -402 597 -402 0 3
rlabel polysilicon 604 -396 604 -396 0 1
rlabel polysilicon 604 -402 604 -402 0 3
rlabel polysilicon 611 -396 611 -396 0 1
rlabel polysilicon 611 -402 611 -402 0 3
rlabel polysilicon 618 -396 618 -396 0 1
rlabel polysilicon 618 -402 618 -402 0 3
rlabel polysilicon 625 -396 625 -396 0 1
rlabel polysilicon 625 -402 625 -402 0 3
rlabel polysilicon 632 -396 632 -396 0 1
rlabel polysilicon 632 -402 632 -402 0 3
rlabel polysilicon 639 -396 639 -396 0 1
rlabel polysilicon 639 -402 639 -402 0 3
rlabel polysilicon 646 -396 646 -396 0 1
rlabel polysilicon 646 -402 646 -402 0 3
rlabel polysilicon 653 -396 653 -396 0 1
rlabel polysilicon 653 -402 653 -402 0 3
rlabel polysilicon 660 -396 660 -396 0 1
rlabel polysilicon 660 -402 660 -402 0 3
rlabel polysilicon 667 -396 667 -396 0 1
rlabel polysilicon 667 -402 667 -402 0 3
rlabel polysilicon 674 -396 674 -396 0 1
rlabel polysilicon 674 -402 674 -402 0 3
rlabel polysilicon 681 -396 681 -396 0 1
rlabel polysilicon 684 -396 684 -396 0 2
rlabel polysilicon 681 -402 681 -402 0 3
rlabel polysilicon 688 -396 688 -396 0 1
rlabel polysilicon 688 -402 688 -402 0 3
rlabel polysilicon 695 -396 695 -396 0 1
rlabel polysilicon 695 -402 695 -402 0 3
rlabel polysilicon 702 -396 702 -396 0 1
rlabel polysilicon 702 -402 702 -402 0 3
rlabel polysilicon 709 -396 709 -396 0 1
rlabel polysilicon 709 -402 709 -402 0 3
rlabel polysilicon 716 -396 716 -396 0 1
rlabel polysilicon 716 -402 716 -402 0 3
rlabel polysilicon 723 -396 723 -396 0 1
rlabel polysilicon 723 -402 723 -402 0 3
rlabel polysilicon 730 -396 730 -396 0 1
rlabel polysilicon 730 -402 730 -402 0 3
rlabel polysilicon 737 -396 737 -396 0 1
rlabel polysilicon 737 -402 737 -402 0 3
rlabel polysilicon 744 -396 744 -396 0 1
rlabel polysilicon 744 -402 744 -402 0 3
rlabel polysilicon 751 -396 751 -396 0 1
rlabel polysilicon 751 -402 751 -402 0 3
rlabel polysilicon 758 -396 758 -396 0 1
rlabel polysilicon 758 -402 758 -402 0 3
rlabel polysilicon 765 -396 765 -396 0 1
rlabel polysilicon 765 -402 765 -402 0 3
rlabel polysilicon 772 -396 772 -396 0 1
rlabel polysilicon 772 -402 772 -402 0 3
rlabel polysilicon 779 -396 779 -396 0 1
rlabel polysilicon 779 -402 779 -402 0 3
rlabel polysilicon 786 -396 786 -396 0 1
rlabel polysilicon 786 -402 786 -402 0 3
rlabel polysilicon 793 -396 793 -396 0 1
rlabel polysilicon 793 -402 793 -402 0 3
rlabel polysilicon 800 -396 800 -396 0 1
rlabel polysilicon 800 -402 800 -402 0 3
rlabel polysilicon 807 -396 807 -396 0 1
rlabel polysilicon 807 -402 807 -402 0 3
rlabel polysilicon 814 -396 814 -396 0 1
rlabel polysilicon 814 -402 814 -402 0 3
rlabel polysilicon 821 -396 821 -396 0 1
rlabel polysilicon 821 -402 821 -402 0 3
rlabel polysilicon 828 -396 828 -396 0 1
rlabel polysilicon 828 -402 828 -402 0 3
rlabel polysilicon 835 -396 835 -396 0 1
rlabel polysilicon 835 -402 835 -402 0 3
rlabel polysilicon 842 -396 842 -396 0 1
rlabel polysilicon 842 -402 842 -402 0 3
rlabel polysilicon 849 -396 849 -396 0 1
rlabel polysilicon 849 -402 849 -402 0 3
rlabel polysilicon 856 -396 856 -396 0 1
rlabel polysilicon 856 -402 856 -402 0 3
rlabel polysilicon 863 -396 863 -396 0 1
rlabel polysilicon 863 -402 863 -402 0 3
rlabel polysilicon 870 -396 870 -396 0 1
rlabel polysilicon 870 -402 870 -402 0 3
rlabel polysilicon 877 -396 877 -396 0 1
rlabel polysilicon 877 -402 877 -402 0 3
rlabel polysilicon 884 -396 884 -396 0 1
rlabel polysilicon 884 -402 884 -402 0 3
rlabel polysilicon 891 -396 891 -396 0 1
rlabel polysilicon 891 -402 891 -402 0 3
rlabel polysilicon 901 -396 901 -396 0 2
rlabel polysilicon 901 -402 901 -402 0 4
rlabel polysilicon 905 -396 905 -396 0 1
rlabel polysilicon 905 -402 905 -402 0 3
rlabel polysilicon 912 -396 912 -396 0 1
rlabel polysilicon 912 -402 912 -402 0 3
rlabel polysilicon 919 -396 919 -396 0 1
rlabel polysilicon 919 -402 919 -402 0 3
rlabel polysilicon 926 -396 926 -396 0 1
rlabel polysilicon 926 -402 926 -402 0 3
rlabel polysilicon 933 -396 933 -396 0 1
rlabel polysilicon 933 -402 933 -402 0 3
rlabel polysilicon 940 -396 940 -396 0 1
rlabel polysilicon 940 -402 940 -402 0 3
rlabel polysilicon 947 -396 947 -396 0 1
rlabel polysilicon 947 -402 947 -402 0 3
rlabel polysilicon 954 -396 954 -396 0 1
rlabel polysilicon 954 -402 954 -402 0 3
rlabel polysilicon 961 -396 961 -396 0 1
rlabel polysilicon 964 -396 964 -396 0 2
rlabel polysilicon 961 -402 961 -402 0 3
rlabel polysilicon 968 -396 968 -396 0 1
rlabel polysilicon 968 -402 968 -402 0 3
rlabel polysilicon 975 -396 975 -396 0 1
rlabel polysilicon 975 -402 975 -402 0 3
rlabel polysilicon 982 -396 982 -396 0 1
rlabel polysilicon 982 -402 982 -402 0 3
rlabel polysilicon 989 -396 989 -396 0 1
rlabel polysilicon 989 -402 989 -402 0 3
rlabel polysilicon 999 -396 999 -396 0 2
rlabel polysilicon 996 -402 996 -402 0 3
rlabel polysilicon 1003 -396 1003 -396 0 1
rlabel polysilicon 1003 -402 1003 -402 0 3
rlabel polysilicon 1010 -396 1010 -396 0 1
rlabel polysilicon 1010 -402 1010 -402 0 3
rlabel polysilicon 1017 -396 1017 -396 0 1
rlabel polysilicon 1017 -402 1017 -402 0 3
rlabel polysilicon 1024 -396 1024 -396 0 1
rlabel polysilicon 1024 -402 1024 -402 0 3
rlabel polysilicon 1031 -402 1031 -402 0 3
rlabel polysilicon 1041 -402 1041 -402 0 4
rlabel polysilicon 1048 -402 1048 -402 0 4
rlabel polysilicon 1052 -396 1052 -396 0 1
rlabel polysilicon 1052 -402 1052 -402 0 3
rlabel polysilicon 1066 -396 1066 -396 0 1
rlabel polysilicon 1066 -402 1066 -402 0 3
rlabel polysilicon 1108 -396 1108 -396 0 1
rlabel polysilicon 1108 -402 1108 -402 0 3
rlabel polysilicon 12 -465 12 -465 0 2
rlabel polysilicon 16 -465 16 -465 0 1
rlabel polysilicon 16 -471 16 -471 0 3
rlabel polysilicon 23 -465 23 -465 0 1
rlabel polysilicon 23 -471 23 -471 0 3
rlabel polysilicon 30 -465 30 -465 0 1
rlabel polysilicon 30 -471 30 -471 0 3
rlabel polysilicon 37 -465 37 -465 0 1
rlabel polysilicon 37 -471 37 -471 0 3
rlabel polysilicon 44 -465 44 -465 0 1
rlabel polysilicon 44 -471 44 -471 0 3
rlabel polysilicon 51 -465 51 -465 0 1
rlabel polysilicon 51 -471 51 -471 0 3
rlabel polysilicon 58 -465 58 -465 0 1
rlabel polysilicon 58 -471 58 -471 0 3
rlabel polysilicon 65 -465 65 -465 0 1
rlabel polysilicon 65 -471 65 -471 0 3
rlabel polysilicon 72 -465 72 -465 0 1
rlabel polysilicon 72 -471 72 -471 0 3
rlabel polysilicon 79 -465 79 -465 0 1
rlabel polysilicon 79 -471 79 -471 0 3
rlabel polysilicon 86 -465 86 -465 0 1
rlabel polysilicon 89 -465 89 -465 0 2
rlabel polysilicon 86 -471 86 -471 0 3
rlabel polysilicon 93 -465 93 -465 0 1
rlabel polysilicon 93 -471 93 -471 0 3
rlabel polysilicon 100 -465 100 -465 0 1
rlabel polysilicon 100 -471 100 -471 0 3
rlabel polysilicon 110 -465 110 -465 0 2
rlabel polysilicon 110 -471 110 -471 0 4
rlabel polysilicon 114 -465 114 -465 0 1
rlabel polysilicon 114 -471 114 -471 0 3
rlabel polysilicon 121 -465 121 -465 0 1
rlabel polysilicon 121 -471 121 -471 0 3
rlabel polysilicon 128 -465 128 -465 0 1
rlabel polysilicon 128 -471 128 -471 0 3
rlabel polysilicon 135 -465 135 -465 0 1
rlabel polysilicon 138 -471 138 -471 0 4
rlabel polysilicon 142 -465 142 -465 0 1
rlabel polysilicon 142 -471 142 -471 0 3
rlabel polysilicon 149 -465 149 -465 0 1
rlabel polysilicon 149 -471 149 -471 0 3
rlabel polysilicon 156 -465 156 -465 0 1
rlabel polysilicon 156 -471 156 -471 0 3
rlabel polysilicon 163 -465 163 -465 0 1
rlabel polysilicon 163 -471 163 -471 0 3
rlabel polysilicon 170 -465 170 -465 0 1
rlabel polysilicon 170 -471 170 -471 0 3
rlabel polysilicon 177 -465 177 -465 0 1
rlabel polysilicon 177 -471 177 -471 0 3
rlabel polysilicon 184 -465 184 -465 0 1
rlabel polysilicon 184 -471 184 -471 0 3
rlabel polysilicon 191 -465 191 -465 0 1
rlabel polysilicon 191 -471 191 -471 0 3
rlabel polysilicon 198 -465 198 -465 0 1
rlabel polysilicon 198 -471 198 -471 0 3
rlabel polysilicon 205 -465 205 -465 0 1
rlabel polysilicon 205 -471 205 -471 0 3
rlabel polysilicon 215 -471 215 -471 0 4
rlabel polysilicon 219 -465 219 -465 0 1
rlabel polysilicon 219 -471 219 -471 0 3
rlabel polysilicon 229 -465 229 -465 0 2
rlabel polysilicon 233 -465 233 -465 0 1
rlabel polysilicon 233 -471 233 -471 0 3
rlabel polysilicon 240 -465 240 -465 0 1
rlabel polysilicon 240 -471 240 -471 0 3
rlabel polysilicon 247 -465 247 -465 0 1
rlabel polysilicon 247 -471 247 -471 0 3
rlabel polysilicon 254 -465 254 -465 0 1
rlabel polysilicon 254 -471 254 -471 0 3
rlabel polysilicon 261 -471 261 -471 0 3
rlabel polysilicon 268 -465 268 -465 0 1
rlabel polysilicon 268 -471 268 -471 0 3
rlabel polysilicon 275 -465 275 -465 0 1
rlabel polysilicon 278 -465 278 -465 0 2
rlabel polysilicon 278 -471 278 -471 0 4
rlabel polysilicon 282 -465 282 -465 0 1
rlabel polysilicon 285 -465 285 -465 0 2
rlabel polysilicon 282 -471 282 -471 0 3
rlabel polysilicon 289 -465 289 -465 0 1
rlabel polysilicon 289 -471 289 -471 0 3
rlabel polysilicon 296 -465 296 -465 0 1
rlabel polysilicon 296 -471 296 -471 0 3
rlabel polysilicon 303 -465 303 -465 0 1
rlabel polysilicon 306 -465 306 -465 0 2
rlabel polysilicon 303 -471 303 -471 0 3
rlabel polysilicon 310 -465 310 -465 0 1
rlabel polysilicon 310 -471 310 -471 0 3
rlabel polysilicon 317 -465 317 -465 0 1
rlabel polysilicon 317 -471 317 -471 0 3
rlabel polysilicon 324 -465 324 -465 0 1
rlabel polysilicon 324 -471 324 -471 0 3
rlabel polysilicon 331 -465 331 -465 0 1
rlabel polysilicon 331 -471 331 -471 0 3
rlabel polysilicon 338 -465 338 -465 0 1
rlabel polysilicon 338 -471 338 -471 0 3
rlabel polysilicon 345 -465 345 -465 0 1
rlabel polysilicon 348 -471 348 -471 0 4
rlabel polysilicon 352 -465 352 -465 0 1
rlabel polysilicon 352 -471 352 -471 0 3
rlabel polysilicon 359 -465 359 -465 0 1
rlabel polysilicon 359 -471 359 -471 0 3
rlabel polysilicon 366 -465 366 -465 0 1
rlabel polysilicon 366 -471 366 -471 0 3
rlabel polysilicon 373 -465 373 -465 0 1
rlabel polysilicon 373 -471 373 -471 0 3
rlabel polysilicon 380 -465 380 -465 0 1
rlabel polysilicon 380 -471 380 -471 0 3
rlabel polysilicon 390 -465 390 -465 0 2
rlabel polysilicon 387 -471 387 -471 0 3
rlabel polysilicon 390 -471 390 -471 0 4
rlabel polysilicon 394 -465 394 -465 0 1
rlabel polysilicon 394 -471 394 -471 0 3
rlabel polysilicon 401 -465 401 -465 0 1
rlabel polysilicon 404 -465 404 -465 0 2
rlabel polysilicon 401 -471 401 -471 0 3
rlabel polysilicon 404 -471 404 -471 0 4
rlabel polysilicon 408 -465 408 -465 0 1
rlabel polysilicon 411 -465 411 -465 0 2
rlabel polysilicon 408 -471 408 -471 0 3
rlabel polysilicon 415 -465 415 -465 0 1
rlabel polysilicon 415 -471 415 -471 0 3
rlabel polysilicon 422 -465 422 -465 0 1
rlabel polysilicon 422 -471 422 -471 0 3
rlabel polysilicon 429 -465 429 -465 0 1
rlabel polysilicon 429 -471 429 -471 0 3
rlabel polysilicon 436 -465 436 -465 0 1
rlabel polysilicon 436 -471 436 -471 0 3
rlabel polysilicon 443 -465 443 -465 0 1
rlabel polysilicon 443 -471 443 -471 0 3
rlabel polysilicon 450 -465 450 -465 0 1
rlabel polysilicon 450 -471 450 -471 0 3
rlabel polysilicon 457 -465 457 -465 0 1
rlabel polysilicon 460 -471 460 -471 0 4
rlabel polysilicon 464 -465 464 -465 0 1
rlabel polysilicon 464 -471 464 -471 0 3
rlabel polysilicon 471 -465 471 -465 0 1
rlabel polysilicon 474 -465 474 -465 0 2
rlabel polysilicon 471 -471 471 -471 0 3
rlabel polysilicon 478 -465 478 -465 0 1
rlabel polysilicon 478 -471 478 -471 0 3
rlabel polysilicon 485 -465 485 -465 0 1
rlabel polysilicon 485 -471 485 -471 0 3
rlabel polysilicon 492 -465 492 -465 0 1
rlabel polysilicon 492 -471 492 -471 0 3
rlabel polysilicon 502 -465 502 -465 0 2
rlabel polysilicon 502 -471 502 -471 0 4
rlabel polysilicon 509 -465 509 -465 0 2
rlabel polysilicon 509 -471 509 -471 0 4
rlabel polysilicon 513 -465 513 -465 0 1
rlabel polysilicon 513 -471 513 -471 0 3
rlabel polysilicon 520 -465 520 -465 0 1
rlabel polysilicon 523 -465 523 -465 0 2
rlabel polysilicon 527 -465 527 -465 0 1
rlabel polysilicon 527 -471 527 -471 0 3
rlabel polysilicon 530 -471 530 -471 0 4
rlabel polysilicon 534 -465 534 -465 0 1
rlabel polysilicon 534 -471 534 -471 0 3
rlabel polysilicon 541 -465 541 -465 0 1
rlabel polysilicon 541 -471 541 -471 0 3
rlabel polysilicon 548 -465 548 -465 0 1
rlabel polysilicon 548 -471 548 -471 0 3
rlabel polysilicon 555 -465 555 -465 0 1
rlabel polysilicon 555 -471 555 -471 0 3
rlabel polysilicon 562 -465 562 -465 0 1
rlabel polysilicon 565 -465 565 -465 0 2
rlabel polysilicon 562 -471 562 -471 0 3
rlabel polysilicon 569 -465 569 -465 0 1
rlabel polysilicon 569 -471 569 -471 0 3
rlabel polysilicon 576 -465 576 -465 0 1
rlabel polysilicon 576 -471 576 -471 0 3
rlabel polysilicon 583 -465 583 -465 0 1
rlabel polysilicon 586 -465 586 -465 0 2
rlabel polysilicon 586 -471 586 -471 0 4
rlabel polysilicon 590 -465 590 -465 0 1
rlabel polysilicon 590 -471 590 -471 0 3
rlabel polysilicon 597 -465 597 -465 0 1
rlabel polysilicon 600 -465 600 -465 0 2
rlabel polysilicon 597 -471 597 -471 0 3
rlabel polysilicon 600 -471 600 -471 0 4
rlabel polysilicon 604 -465 604 -465 0 1
rlabel polysilicon 604 -471 604 -471 0 3
rlabel polysilicon 611 -465 611 -465 0 1
rlabel polysilicon 611 -471 611 -471 0 3
rlabel polysilicon 618 -465 618 -465 0 1
rlabel polysilicon 618 -471 618 -471 0 3
rlabel polysilicon 625 -465 625 -465 0 1
rlabel polysilicon 625 -471 625 -471 0 3
rlabel polysilicon 635 -465 635 -465 0 2
rlabel polysilicon 632 -471 632 -471 0 3
rlabel polysilicon 635 -471 635 -471 0 4
rlabel polysilicon 639 -465 639 -465 0 1
rlabel polysilicon 639 -471 639 -471 0 3
rlabel polysilicon 646 -465 646 -465 0 1
rlabel polysilicon 646 -471 646 -471 0 3
rlabel polysilicon 653 -465 653 -465 0 1
rlabel polysilicon 653 -471 653 -471 0 3
rlabel polysilicon 660 -465 660 -465 0 1
rlabel polysilicon 660 -471 660 -471 0 3
rlabel polysilicon 667 -465 667 -465 0 1
rlabel polysilicon 667 -471 667 -471 0 3
rlabel polysilicon 674 -465 674 -465 0 1
rlabel polysilicon 674 -471 674 -471 0 3
rlabel polysilicon 681 -465 681 -465 0 1
rlabel polysilicon 681 -471 681 -471 0 3
rlabel polysilicon 688 -465 688 -465 0 1
rlabel polysilicon 688 -471 688 -471 0 3
rlabel polysilicon 695 -465 695 -465 0 1
rlabel polysilicon 695 -471 695 -471 0 3
rlabel polysilicon 702 -465 702 -465 0 1
rlabel polysilicon 702 -471 702 -471 0 3
rlabel polysilicon 709 -465 709 -465 0 1
rlabel polysilicon 709 -471 709 -471 0 3
rlabel polysilicon 716 -465 716 -465 0 1
rlabel polysilicon 716 -471 716 -471 0 3
rlabel polysilicon 723 -465 723 -465 0 1
rlabel polysilicon 723 -471 723 -471 0 3
rlabel polysilicon 730 -465 730 -465 0 1
rlabel polysilicon 730 -471 730 -471 0 3
rlabel polysilicon 737 -465 737 -465 0 1
rlabel polysilicon 740 -465 740 -465 0 2
rlabel polysilicon 744 -465 744 -465 0 1
rlabel polysilicon 744 -471 744 -471 0 3
rlabel polysilicon 754 -465 754 -465 0 2
rlabel polysilicon 754 -471 754 -471 0 4
rlabel polysilicon 758 -465 758 -465 0 1
rlabel polysilicon 758 -471 758 -471 0 3
rlabel polysilicon 765 -465 765 -465 0 1
rlabel polysilicon 765 -471 765 -471 0 3
rlabel polysilicon 772 -465 772 -465 0 1
rlabel polysilicon 772 -471 772 -471 0 3
rlabel polysilicon 779 -465 779 -465 0 1
rlabel polysilicon 779 -471 779 -471 0 3
rlabel polysilicon 786 -465 786 -465 0 1
rlabel polysilicon 786 -471 786 -471 0 3
rlabel polysilicon 793 -465 793 -465 0 1
rlabel polysilicon 793 -471 793 -471 0 3
rlabel polysilicon 800 -465 800 -465 0 1
rlabel polysilicon 800 -471 800 -471 0 3
rlabel polysilicon 807 -465 807 -465 0 1
rlabel polysilicon 807 -471 807 -471 0 3
rlabel polysilicon 814 -465 814 -465 0 1
rlabel polysilicon 814 -471 814 -471 0 3
rlabel polysilicon 821 -465 821 -465 0 1
rlabel polysilicon 821 -471 821 -471 0 3
rlabel polysilicon 828 -465 828 -465 0 1
rlabel polysilicon 828 -471 828 -471 0 3
rlabel polysilicon 835 -465 835 -465 0 1
rlabel polysilicon 835 -471 835 -471 0 3
rlabel polysilicon 842 -465 842 -465 0 1
rlabel polysilicon 842 -471 842 -471 0 3
rlabel polysilicon 849 -465 849 -465 0 1
rlabel polysilicon 849 -471 849 -471 0 3
rlabel polysilicon 856 -465 856 -465 0 1
rlabel polysilicon 856 -471 856 -471 0 3
rlabel polysilicon 863 -465 863 -465 0 1
rlabel polysilicon 863 -471 863 -471 0 3
rlabel polysilicon 870 -465 870 -465 0 1
rlabel polysilicon 870 -471 870 -471 0 3
rlabel polysilicon 877 -465 877 -465 0 1
rlabel polysilicon 877 -471 877 -471 0 3
rlabel polysilicon 884 -465 884 -465 0 1
rlabel polysilicon 884 -471 884 -471 0 3
rlabel polysilicon 891 -465 891 -465 0 1
rlabel polysilicon 891 -471 891 -471 0 3
rlabel polysilicon 898 -465 898 -465 0 1
rlabel polysilicon 898 -471 898 -471 0 3
rlabel polysilicon 905 -465 905 -465 0 1
rlabel polysilicon 905 -471 905 -471 0 3
rlabel polysilicon 912 -465 912 -465 0 1
rlabel polysilicon 912 -471 912 -471 0 3
rlabel polysilicon 919 -465 919 -465 0 1
rlabel polysilicon 919 -471 919 -471 0 3
rlabel polysilicon 926 -465 926 -465 0 1
rlabel polysilicon 926 -471 926 -471 0 3
rlabel polysilicon 933 -465 933 -465 0 1
rlabel polysilicon 933 -471 933 -471 0 3
rlabel polysilicon 940 -465 940 -465 0 1
rlabel polysilicon 940 -471 940 -471 0 3
rlabel polysilicon 947 -465 947 -465 0 1
rlabel polysilicon 947 -471 947 -471 0 3
rlabel polysilicon 954 -465 954 -465 0 1
rlabel polysilicon 954 -471 954 -471 0 3
rlabel polysilicon 961 -465 961 -465 0 1
rlabel polysilicon 961 -471 961 -471 0 3
rlabel polysilicon 968 -465 968 -465 0 1
rlabel polysilicon 968 -471 968 -471 0 3
rlabel polysilicon 975 -465 975 -465 0 1
rlabel polysilicon 975 -471 975 -471 0 3
rlabel polysilicon 982 -465 982 -465 0 1
rlabel polysilicon 989 -465 989 -465 0 1
rlabel polysilicon 989 -471 989 -471 0 3
rlabel polysilicon 996 -465 996 -465 0 1
rlabel polysilicon 996 -471 996 -471 0 3
rlabel polysilicon 1003 -465 1003 -465 0 1
rlabel polysilicon 1003 -471 1003 -471 0 3
rlabel polysilicon 1010 -465 1010 -465 0 1
rlabel polysilicon 1010 -471 1010 -471 0 3
rlabel polysilicon 1017 -465 1017 -465 0 1
rlabel polysilicon 1017 -471 1017 -471 0 3
rlabel polysilicon 1024 -465 1024 -465 0 1
rlabel polysilicon 1024 -471 1024 -471 0 3
rlabel polysilicon 1031 -465 1031 -465 0 1
rlabel polysilicon 1031 -471 1031 -471 0 3
rlabel polysilicon 1038 -465 1038 -465 0 1
rlabel polysilicon 1038 -471 1038 -471 0 3
rlabel polysilicon 1045 -465 1045 -465 0 1
rlabel polysilicon 1045 -471 1045 -471 0 3
rlabel polysilicon 1052 -465 1052 -465 0 1
rlabel polysilicon 1052 -471 1052 -471 0 3
rlabel polysilicon 1059 -465 1059 -465 0 1
rlabel polysilicon 1059 -471 1059 -471 0 3
rlabel polysilicon 1066 -465 1066 -465 0 1
rlabel polysilicon 1066 -471 1066 -471 0 3
rlabel polysilicon 1073 -465 1073 -465 0 1
rlabel polysilicon 1073 -471 1073 -471 0 3
rlabel polysilicon 1080 -465 1080 -465 0 1
rlabel polysilicon 1080 -471 1080 -471 0 3
rlabel polysilicon 1087 -465 1087 -465 0 1
rlabel polysilicon 1087 -471 1087 -471 0 3
rlabel polysilicon 1094 -465 1094 -465 0 1
rlabel polysilicon 1094 -471 1094 -471 0 3
rlabel polysilicon 1101 -465 1101 -465 0 1
rlabel polysilicon 1101 -471 1101 -471 0 3
rlabel polysilicon 1108 -465 1108 -465 0 1
rlabel polysilicon 1108 -471 1108 -471 0 3
rlabel polysilicon 1115 -465 1115 -465 0 1
rlabel polysilicon 1115 -471 1115 -471 0 3
rlabel polysilicon 1122 -465 1122 -465 0 1
rlabel polysilicon 1122 -471 1122 -471 0 3
rlabel polysilicon 1129 -465 1129 -465 0 1
rlabel polysilicon 1129 -471 1129 -471 0 3
rlabel polysilicon 1139 -465 1139 -465 0 2
rlabel polysilicon 1139 -471 1139 -471 0 4
rlabel polysilicon 1143 -471 1143 -471 0 3
rlabel polysilicon 1150 -465 1150 -465 0 1
rlabel polysilicon 1150 -471 1150 -471 0 3
rlabel polysilicon 2 -566 2 -566 0 3
rlabel polysilicon 9 -560 9 -560 0 1
rlabel polysilicon 9 -566 9 -566 0 3
rlabel polysilicon 16 -560 16 -560 0 1
rlabel polysilicon 16 -566 16 -566 0 3
rlabel polysilicon 23 -560 23 -560 0 1
rlabel polysilicon 23 -566 23 -566 0 3
rlabel polysilicon 33 -560 33 -560 0 2
rlabel polysilicon 30 -566 30 -566 0 3
rlabel polysilicon 33 -566 33 -566 0 4
rlabel polysilicon 37 -560 37 -560 0 1
rlabel polysilicon 37 -566 37 -566 0 3
rlabel polysilicon 44 -560 44 -560 0 1
rlabel polysilicon 44 -566 44 -566 0 3
rlabel polysilicon 51 -560 51 -560 0 1
rlabel polysilicon 51 -566 51 -566 0 3
rlabel polysilicon 58 -560 58 -560 0 1
rlabel polysilicon 58 -566 58 -566 0 3
rlabel polysilicon 65 -560 65 -560 0 1
rlabel polysilicon 65 -566 65 -566 0 3
rlabel polysilicon 72 -566 72 -566 0 3
rlabel polysilicon 75 -566 75 -566 0 4
rlabel polysilicon 79 -566 79 -566 0 3
rlabel polysilicon 82 -566 82 -566 0 4
rlabel polysilicon 86 -560 86 -560 0 1
rlabel polysilicon 86 -566 86 -566 0 3
rlabel polysilicon 93 -560 93 -560 0 1
rlabel polysilicon 93 -566 93 -566 0 3
rlabel polysilicon 100 -560 100 -560 0 1
rlabel polysilicon 100 -566 100 -566 0 3
rlabel polysilicon 107 -560 107 -560 0 1
rlabel polysilicon 110 -560 110 -560 0 2
rlabel polysilicon 107 -566 107 -566 0 3
rlabel polysilicon 114 -560 114 -560 0 1
rlabel polysilicon 114 -566 114 -566 0 3
rlabel polysilicon 121 -560 121 -560 0 1
rlabel polysilicon 121 -566 121 -566 0 3
rlabel polysilicon 128 -560 128 -560 0 1
rlabel polysilicon 128 -566 128 -566 0 3
rlabel polysilicon 135 -560 135 -560 0 1
rlabel polysilicon 135 -566 135 -566 0 3
rlabel polysilicon 142 -560 142 -560 0 1
rlabel polysilicon 142 -566 142 -566 0 3
rlabel polysilicon 152 -560 152 -560 0 2
rlabel polysilicon 152 -566 152 -566 0 4
rlabel polysilicon 156 -560 156 -560 0 1
rlabel polysilicon 156 -566 156 -566 0 3
rlabel polysilicon 166 -560 166 -560 0 2
rlabel polysilicon 163 -566 163 -566 0 3
rlabel polysilicon 166 -566 166 -566 0 4
rlabel polysilicon 170 -560 170 -560 0 1
rlabel polysilicon 170 -566 170 -566 0 3
rlabel polysilicon 177 -560 177 -560 0 1
rlabel polysilicon 177 -566 177 -566 0 3
rlabel polysilicon 184 -560 184 -560 0 1
rlabel polysilicon 184 -566 184 -566 0 3
rlabel polysilicon 191 -560 191 -560 0 1
rlabel polysilicon 194 -560 194 -560 0 2
rlabel polysilicon 198 -560 198 -560 0 1
rlabel polysilicon 201 -560 201 -560 0 2
rlabel polysilicon 201 -566 201 -566 0 4
rlabel polysilicon 205 -560 205 -560 0 1
rlabel polysilicon 205 -566 205 -566 0 3
rlabel polysilicon 215 -560 215 -560 0 2
rlabel polysilicon 212 -566 212 -566 0 3
rlabel polysilicon 219 -560 219 -560 0 1
rlabel polysilicon 219 -566 219 -566 0 3
rlabel polysilicon 226 -560 226 -560 0 1
rlabel polysilicon 226 -566 226 -566 0 3
rlabel polysilicon 233 -560 233 -560 0 1
rlabel polysilicon 233 -566 233 -566 0 3
rlabel polysilicon 240 -560 240 -560 0 1
rlabel polysilicon 240 -566 240 -566 0 3
rlabel polysilicon 247 -560 247 -560 0 1
rlabel polysilicon 247 -566 247 -566 0 3
rlabel polysilicon 254 -560 254 -560 0 1
rlabel polysilicon 254 -566 254 -566 0 3
rlabel polysilicon 261 -560 261 -560 0 1
rlabel polysilicon 261 -566 261 -566 0 3
rlabel polysilicon 268 -560 268 -560 0 1
rlabel polysilicon 268 -566 268 -566 0 3
rlabel polysilicon 275 -560 275 -560 0 1
rlabel polysilicon 275 -566 275 -566 0 3
rlabel polysilicon 282 -560 282 -560 0 1
rlabel polysilicon 282 -566 282 -566 0 3
rlabel polysilicon 289 -560 289 -560 0 1
rlabel polysilicon 289 -566 289 -566 0 3
rlabel polysilicon 296 -560 296 -560 0 1
rlabel polysilicon 296 -566 296 -566 0 3
rlabel polysilicon 303 -560 303 -560 0 1
rlabel polysilicon 303 -566 303 -566 0 3
rlabel polysilicon 310 -560 310 -560 0 1
rlabel polysilicon 310 -566 310 -566 0 3
rlabel polysilicon 317 -560 317 -560 0 1
rlabel polysilicon 320 -560 320 -560 0 2
rlabel polysilicon 317 -566 317 -566 0 3
rlabel polysilicon 320 -566 320 -566 0 4
rlabel polysilicon 324 -560 324 -560 0 1
rlabel polysilicon 324 -566 324 -566 0 3
rlabel polysilicon 331 -560 331 -560 0 1
rlabel polysilicon 331 -566 331 -566 0 3
rlabel polysilicon 338 -560 338 -560 0 1
rlabel polysilicon 338 -566 338 -566 0 3
rlabel polysilicon 345 -560 345 -560 0 1
rlabel polysilicon 345 -566 345 -566 0 3
rlabel polysilicon 355 -560 355 -560 0 2
rlabel polysilicon 352 -566 352 -566 0 3
rlabel polysilicon 355 -566 355 -566 0 4
rlabel polysilicon 359 -560 359 -560 0 1
rlabel polysilicon 359 -566 359 -566 0 3
rlabel polysilicon 366 -566 366 -566 0 3
rlabel polysilicon 373 -560 373 -560 0 1
rlabel polysilicon 373 -566 373 -566 0 3
rlabel polysilicon 380 -560 380 -560 0 1
rlabel polysilicon 380 -566 380 -566 0 3
rlabel polysilicon 390 -560 390 -560 0 2
rlabel polysilicon 390 -566 390 -566 0 4
rlabel polysilicon 397 -560 397 -560 0 2
rlabel polysilicon 397 -566 397 -566 0 4
rlabel polysilicon 401 -560 401 -560 0 1
rlabel polysilicon 401 -566 401 -566 0 3
rlabel polysilicon 408 -560 408 -560 0 1
rlabel polysilicon 408 -566 408 -566 0 3
rlabel polysilicon 411 -566 411 -566 0 4
rlabel polysilicon 415 -560 415 -560 0 1
rlabel polysilicon 415 -566 415 -566 0 3
rlabel polysilicon 422 -560 422 -560 0 1
rlabel polysilicon 422 -566 422 -566 0 3
rlabel polysilicon 429 -560 429 -560 0 1
rlabel polysilicon 429 -566 429 -566 0 3
rlabel polysilicon 436 -560 436 -560 0 1
rlabel polysilicon 436 -566 436 -566 0 3
rlabel polysilicon 443 -560 443 -560 0 1
rlabel polysilicon 443 -566 443 -566 0 3
rlabel polysilicon 450 -560 450 -560 0 1
rlabel polysilicon 450 -566 450 -566 0 3
rlabel polysilicon 457 -560 457 -560 0 1
rlabel polysilicon 457 -566 457 -566 0 3
rlabel polysilicon 464 -560 464 -560 0 1
rlabel polysilicon 464 -566 464 -566 0 3
rlabel polysilicon 471 -560 471 -560 0 1
rlabel polysilicon 471 -566 471 -566 0 3
rlabel polysilicon 478 -560 478 -560 0 1
rlabel polysilicon 478 -566 478 -566 0 3
rlabel polysilicon 485 -560 485 -560 0 1
rlabel polysilicon 485 -566 485 -566 0 3
rlabel polysilicon 492 -560 492 -560 0 1
rlabel polysilicon 492 -566 492 -566 0 3
rlabel polysilicon 499 -560 499 -560 0 1
rlabel polysilicon 499 -566 499 -566 0 3
rlabel polysilicon 506 -560 506 -560 0 1
rlabel polysilicon 509 -560 509 -560 0 2
rlabel polysilicon 506 -566 506 -566 0 3
rlabel polysilicon 509 -566 509 -566 0 4
rlabel polysilicon 513 -560 513 -560 0 1
rlabel polysilicon 513 -566 513 -566 0 3
rlabel polysilicon 520 -560 520 -560 0 1
rlabel polysilicon 520 -566 520 -566 0 3
rlabel polysilicon 527 -560 527 -560 0 1
rlabel polysilicon 527 -566 527 -566 0 3
rlabel polysilicon 537 -560 537 -560 0 2
rlabel polysilicon 537 -566 537 -566 0 4
rlabel polysilicon 541 -560 541 -560 0 1
rlabel polysilicon 541 -566 541 -566 0 3
rlabel polysilicon 548 -560 548 -560 0 1
rlabel polysilicon 551 -560 551 -560 0 2
rlabel polysilicon 548 -566 548 -566 0 3
rlabel polysilicon 551 -566 551 -566 0 4
rlabel polysilicon 555 -560 555 -560 0 1
rlabel polysilicon 555 -566 555 -566 0 3
rlabel polysilicon 562 -560 562 -560 0 1
rlabel polysilicon 565 -560 565 -560 0 2
rlabel polysilicon 562 -566 562 -566 0 3
rlabel polysilicon 569 -560 569 -560 0 1
rlabel polysilicon 572 -560 572 -560 0 2
rlabel polysilicon 569 -566 569 -566 0 3
rlabel polysilicon 572 -566 572 -566 0 4
rlabel polysilicon 576 -560 576 -560 0 1
rlabel polysilicon 576 -566 576 -566 0 3
rlabel polysilicon 583 -560 583 -560 0 1
rlabel polysilicon 583 -566 583 -566 0 3
rlabel polysilicon 593 -560 593 -560 0 2
rlabel polysilicon 590 -566 590 -566 0 3
rlabel polysilicon 597 -560 597 -560 0 1
rlabel polysilicon 600 -566 600 -566 0 4
rlabel polysilicon 604 -560 604 -560 0 1
rlabel polysilicon 604 -566 604 -566 0 3
rlabel polysilicon 607 -566 607 -566 0 4
rlabel polysilicon 611 -560 611 -560 0 1
rlabel polysilicon 611 -566 611 -566 0 3
rlabel polysilicon 618 -560 618 -560 0 1
rlabel polysilicon 618 -566 618 -566 0 3
rlabel polysilicon 628 -560 628 -560 0 2
rlabel polysilicon 628 -566 628 -566 0 4
rlabel polysilicon 632 -560 632 -560 0 1
rlabel polysilicon 632 -566 632 -566 0 3
rlabel polysilicon 639 -560 639 -560 0 1
rlabel polysilicon 639 -566 639 -566 0 3
rlabel polysilicon 646 -560 646 -560 0 1
rlabel polysilicon 646 -566 646 -566 0 3
rlabel polysilicon 653 -560 653 -560 0 1
rlabel polysilicon 653 -566 653 -566 0 3
rlabel polysilicon 660 -560 660 -560 0 1
rlabel polysilicon 663 -560 663 -560 0 2
rlabel polysilicon 660 -566 660 -566 0 3
rlabel polysilicon 663 -566 663 -566 0 4
rlabel polysilicon 667 -560 667 -560 0 1
rlabel polysilicon 667 -566 667 -566 0 3
rlabel polysilicon 674 -560 674 -560 0 1
rlabel polysilicon 674 -566 674 -566 0 3
rlabel polysilicon 681 -560 681 -560 0 1
rlabel polysilicon 681 -566 681 -566 0 3
rlabel polysilicon 688 -560 688 -560 0 1
rlabel polysilicon 688 -566 688 -566 0 3
rlabel polysilicon 695 -560 695 -560 0 1
rlabel polysilicon 695 -566 695 -566 0 3
rlabel polysilicon 702 -560 702 -560 0 1
rlabel polysilicon 702 -566 702 -566 0 3
rlabel polysilicon 709 -560 709 -560 0 1
rlabel polysilicon 712 -566 712 -566 0 4
rlabel polysilicon 716 -560 716 -560 0 1
rlabel polysilicon 716 -566 716 -566 0 3
rlabel polysilicon 723 -560 723 -560 0 1
rlabel polysilicon 723 -566 723 -566 0 3
rlabel polysilicon 730 -560 730 -560 0 1
rlabel polysilicon 733 -560 733 -560 0 2
rlabel polysilicon 733 -566 733 -566 0 4
rlabel polysilicon 737 -560 737 -560 0 1
rlabel polysilicon 737 -566 737 -566 0 3
rlabel polysilicon 744 -560 744 -560 0 1
rlabel polysilicon 744 -566 744 -566 0 3
rlabel polysilicon 751 -560 751 -560 0 1
rlabel polysilicon 751 -566 751 -566 0 3
rlabel polysilicon 758 -560 758 -560 0 1
rlabel polysilicon 758 -566 758 -566 0 3
rlabel polysilicon 765 -560 765 -560 0 1
rlabel polysilicon 765 -566 765 -566 0 3
rlabel polysilicon 772 -560 772 -560 0 1
rlabel polysilicon 772 -566 772 -566 0 3
rlabel polysilicon 779 -560 779 -560 0 1
rlabel polysilicon 779 -566 779 -566 0 3
rlabel polysilicon 786 -560 786 -560 0 1
rlabel polysilicon 786 -566 786 -566 0 3
rlabel polysilicon 793 -560 793 -560 0 1
rlabel polysilicon 793 -566 793 -566 0 3
rlabel polysilicon 800 -560 800 -560 0 1
rlabel polysilicon 800 -566 800 -566 0 3
rlabel polysilicon 807 -560 807 -560 0 1
rlabel polysilicon 807 -566 807 -566 0 3
rlabel polysilicon 814 -560 814 -560 0 1
rlabel polysilicon 814 -566 814 -566 0 3
rlabel polysilicon 821 -560 821 -560 0 1
rlabel polysilicon 821 -566 821 -566 0 3
rlabel polysilicon 828 -560 828 -560 0 1
rlabel polysilicon 828 -566 828 -566 0 3
rlabel polysilicon 835 -560 835 -560 0 1
rlabel polysilicon 835 -566 835 -566 0 3
rlabel polysilicon 842 -560 842 -560 0 1
rlabel polysilicon 842 -566 842 -566 0 3
rlabel polysilicon 849 -560 849 -560 0 1
rlabel polysilicon 849 -566 849 -566 0 3
rlabel polysilicon 856 -560 856 -560 0 1
rlabel polysilicon 856 -566 856 -566 0 3
rlabel polysilicon 863 -560 863 -560 0 1
rlabel polysilicon 863 -566 863 -566 0 3
rlabel polysilicon 870 -560 870 -560 0 1
rlabel polysilicon 870 -566 870 -566 0 3
rlabel polysilicon 877 -560 877 -560 0 1
rlabel polysilicon 877 -566 877 -566 0 3
rlabel polysilicon 884 -560 884 -560 0 1
rlabel polysilicon 884 -566 884 -566 0 3
rlabel polysilicon 891 -560 891 -560 0 1
rlabel polysilicon 891 -566 891 -566 0 3
rlabel polysilicon 898 -560 898 -560 0 1
rlabel polysilicon 898 -566 898 -566 0 3
rlabel polysilicon 905 -560 905 -560 0 1
rlabel polysilicon 905 -566 905 -566 0 3
rlabel polysilicon 912 -560 912 -560 0 1
rlabel polysilicon 912 -566 912 -566 0 3
rlabel polysilicon 919 -560 919 -560 0 1
rlabel polysilicon 919 -566 919 -566 0 3
rlabel polysilicon 926 -560 926 -560 0 1
rlabel polysilicon 926 -566 926 -566 0 3
rlabel polysilicon 933 -560 933 -560 0 1
rlabel polysilicon 933 -566 933 -566 0 3
rlabel polysilicon 940 -560 940 -560 0 1
rlabel polysilicon 940 -566 940 -566 0 3
rlabel polysilicon 947 -560 947 -560 0 1
rlabel polysilicon 947 -566 947 -566 0 3
rlabel polysilicon 954 -560 954 -560 0 1
rlabel polysilicon 954 -566 954 -566 0 3
rlabel polysilicon 961 -560 961 -560 0 1
rlabel polysilicon 961 -566 961 -566 0 3
rlabel polysilicon 968 -560 968 -560 0 1
rlabel polysilicon 968 -566 968 -566 0 3
rlabel polysilicon 975 -560 975 -560 0 1
rlabel polysilicon 975 -566 975 -566 0 3
rlabel polysilicon 982 -560 982 -560 0 1
rlabel polysilicon 982 -566 982 -566 0 3
rlabel polysilicon 989 -560 989 -560 0 1
rlabel polysilicon 989 -566 989 -566 0 3
rlabel polysilicon 996 -560 996 -560 0 1
rlabel polysilicon 996 -566 996 -566 0 3
rlabel polysilicon 1003 -560 1003 -560 0 1
rlabel polysilicon 1003 -566 1003 -566 0 3
rlabel polysilicon 1010 -560 1010 -560 0 1
rlabel polysilicon 1010 -566 1010 -566 0 3
rlabel polysilicon 1017 -560 1017 -560 0 1
rlabel polysilicon 1017 -566 1017 -566 0 3
rlabel polysilicon 1024 -560 1024 -560 0 1
rlabel polysilicon 1024 -566 1024 -566 0 3
rlabel polysilicon 1031 -560 1031 -560 0 1
rlabel polysilicon 1031 -566 1031 -566 0 3
rlabel polysilicon 1038 -560 1038 -560 0 1
rlabel polysilicon 1038 -566 1038 -566 0 3
rlabel polysilicon 1045 -560 1045 -560 0 1
rlabel polysilicon 1045 -566 1045 -566 0 3
rlabel polysilicon 1052 -560 1052 -560 0 1
rlabel polysilicon 1052 -566 1052 -566 0 3
rlabel polysilicon 1059 -560 1059 -560 0 1
rlabel polysilicon 1059 -566 1059 -566 0 3
rlabel polysilicon 1066 -560 1066 -560 0 1
rlabel polysilicon 1066 -566 1066 -566 0 3
rlabel polysilicon 1073 -560 1073 -560 0 1
rlabel polysilicon 1073 -566 1073 -566 0 3
rlabel polysilicon 1080 -560 1080 -560 0 1
rlabel polysilicon 1080 -566 1080 -566 0 3
rlabel polysilicon 1087 -560 1087 -560 0 1
rlabel polysilicon 1087 -566 1087 -566 0 3
rlabel polysilicon 1094 -560 1094 -560 0 1
rlabel polysilicon 1094 -566 1094 -566 0 3
rlabel polysilicon 1101 -560 1101 -560 0 1
rlabel polysilicon 1101 -566 1101 -566 0 3
rlabel polysilicon 1115 -560 1115 -560 0 1
rlabel polysilicon 1115 -566 1115 -566 0 3
rlabel polysilicon 1122 -560 1122 -560 0 1
rlabel polysilicon 1122 -566 1122 -566 0 3
rlabel polysilicon 1174 -560 1174 -560 0 2
rlabel polysilicon 1178 -560 1178 -560 0 1
rlabel polysilicon 1178 -566 1178 -566 0 3
rlabel polysilicon 9 -651 9 -651 0 1
rlabel polysilicon 9 -657 9 -657 0 3
rlabel polysilicon 16 -651 16 -651 0 1
rlabel polysilicon 16 -657 16 -657 0 3
rlabel polysilicon 23 -651 23 -651 0 1
rlabel polysilicon 30 -651 30 -651 0 1
rlabel polysilicon 30 -657 30 -657 0 3
rlabel polysilicon 37 -651 37 -651 0 1
rlabel polysilicon 37 -657 37 -657 0 3
rlabel polysilicon 44 -651 44 -651 0 1
rlabel polysilicon 44 -657 44 -657 0 3
rlabel polysilicon 54 -651 54 -651 0 2
rlabel polysilicon 54 -657 54 -657 0 4
rlabel polysilicon 58 -651 58 -651 0 1
rlabel polysilicon 58 -657 58 -657 0 3
rlabel polysilicon 68 -651 68 -651 0 2
rlabel polysilicon 65 -657 65 -657 0 3
rlabel polysilicon 72 -651 72 -651 0 1
rlabel polysilicon 72 -657 72 -657 0 3
rlabel polysilicon 79 -651 79 -651 0 1
rlabel polysilicon 79 -657 79 -657 0 3
rlabel polysilicon 82 -657 82 -657 0 4
rlabel polysilicon 86 -651 86 -651 0 1
rlabel polysilicon 89 -657 89 -657 0 4
rlabel polysilicon 93 -651 93 -651 0 1
rlabel polysilicon 93 -657 93 -657 0 3
rlabel polysilicon 100 -651 100 -651 0 1
rlabel polysilicon 103 -657 103 -657 0 4
rlabel polysilicon 107 -651 107 -651 0 1
rlabel polysilicon 107 -657 107 -657 0 3
rlabel polysilicon 117 -651 117 -651 0 2
rlabel polysilicon 117 -657 117 -657 0 4
rlabel polysilicon 121 -651 121 -651 0 1
rlabel polysilicon 121 -657 121 -657 0 3
rlabel polysilicon 131 -657 131 -657 0 4
rlabel polysilicon 135 -651 135 -651 0 1
rlabel polysilicon 135 -657 135 -657 0 3
rlabel polysilicon 142 -651 142 -651 0 1
rlabel polysilicon 142 -657 142 -657 0 3
rlabel polysilicon 149 -651 149 -651 0 1
rlabel polysilicon 149 -657 149 -657 0 3
rlabel polysilicon 156 -657 156 -657 0 3
rlabel polysilicon 159 -657 159 -657 0 4
rlabel polysilicon 163 -651 163 -651 0 1
rlabel polysilicon 163 -657 163 -657 0 3
rlabel polysilicon 170 -651 170 -651 0 1
rlabel polysilicon 170 -657 170 -657 0 3
rlabel polysilicon 177 -651 177 -651 0 1
rlabel polysilicon 177 -657 177 -657 0 3
rlabel polysilicon 184 -651 184 -651 0 1
rlabel polysilicon 187 -651 187 -651 0 2
rlabel polysilicon 184 -657 184 -657 0 3
rlabel polysilicon 187 -657 187 -657 0 4
rlabel polysilicon 191 -651 191 -651 0 1
rlabel polysilicon 191 -657 191 -657 0 3
rlabel polysilicon 198 -651 198 -651 0 1
rlabel polysilicon 198 -657 198 -657 0 3
rlabel polysilicon 205 -651 205 -651 0 1
rlabel polysilicon 205 -657 205 -657 0 3
rlabel polysilicon 212 -651 212 -651 0 1
rlabel polysilicon 212 -657 212 -657 0 3
rlabel polysilicon 219 -651 219 -651 0 1
rlabel polysilicon 219 -657 219 -657 0 3
rlabel polysilicon 226 -651 226 -651 0 1
rlabel polysilicon 226 -657 226 -657 0 3
rlabel polysilicon 233 -657 233 -657 0 3
rlabel polysilicon 236 -657 236 -657 0 4
rlabel polysilicon 240 -651 240 -651 0 1
rlabel polysilicon 240 -657 240 -657 0 3
rlabel polysilicon 247 -651 247 -651 0 1
rlabel polysilicon 254 -651 254 -651 0 1
rlabel polysilicon 254 -657 254 -657 0 3
rlabel polysilicon 261 -651 261 -651 0 1
rlabel polysilicon 261 -657 261 -657 0 3
rlabel polysilicon 268 -651 268 -651 0 1
rlabel polysilicon 268 -657 268 -657 0 3
rlabel polysilicon 275 -651 275 -651 0 1
rlabel polysilicon 275 -657 275 -657 0 3
rlabel polysilicon 282 -651 282 -651 0 1
rlabel polysilicon 282 -657 282 -657 0 3
rlabel polysilicon 289 -651 289 -651 0 1
rlabel polysilicon 289 -657 289 -657 0 3
rlabel polysilicon 296 -651 296 -651 0 1
rlabel polysilicon 296 -657 296 -657 0 3
rlabel polysilicon 303 -651 303 -651 0 1
rlabel polysilicon 303 -657 303 -657 0 3
rlabel polysilicon 310 -651 310 -651 0 1
rlabel polysilicon 310 -657 310 -657 0 3
rlabel polysilicon 317 -651 317 -651 0 1
rlabel polysilicon 317 -657 317 -657 0 3
rlabel polysilicon 324 -651 324 -651 0 1
rlabel polysilicon 324 -657 324 -657 0 3
rlabel polysilicon 331 -651 331 -651 0 1
rlabel polysilicon 341 -651 341 -651 0 2
rlabel polysilicon 338 -657 338 -657 0 3
rlabel polysilicon 345 -651 345 -651 0 1
rlabel polysilicon 348 -651 348 -651 0 2
rlabel polysilicon 345 -657 345 -657 0 3
rlabel polysilicon 352 -651 352 -651 0 1
rlabel polysilicon 352 -657 352 -657 0 3
rlabel polysilicon 359 -651 359 -651 0 1
rlabel polysilicon 359 -657 359 -657 0 3
rlabel polysilicon 366 -651 366 -651 0 1
rlabel polysilicon 366 -657 366 -657 0 3
rlabel polysilicon 373 -651 373 -651 0 1
rlabel polysilicon 373 -657 373 -657 0 3
rlabel polysilicon 380 -651 380 -651 0 1
rlabel polysilicon 380 -657 380 -657 0 3
rlabel polysilicon 387 -651 387 -651 0 1
rlabel polysilicon 387 -657 387 -657 0 3
rlabel polysilicon 394 -651 394 -651 0 1
rlabel polysilicon 394 -657 394 -657 0 3
rlabel polysilicon 401 -651 401 -651 0 1
rlabel polysilicon 401 -657 401 -657 0 3
rlabel polysilicon 408 -651 408 -651 0 1
rlabel polysilicon 408 -657 408 -657 0 3
rlabel polysilicon 418 -651 418 -651 0 2
rlabel polysilicon 418 -657 418 -657 0 4
rlabel polysilicon 422 -651 422 -651 0 1
rlabel polysilicon 422 -657 422 -657 0 3
rlabel polysilicon 429 -651 429 -651 0 1
rlabel polysilicon 429 -657 429 -657 0 3
rlabel polysilicon 436 -651 436 -651 0 1
rlabel polysilicon 436 -657 436 -657 0 3
rlabel polysilicon 446 -651 446 -651 0 2
rlabel polysilicon 443 -657 443 -657 0 3
rlabel polysilicon 446 -657 446 -657 0 4
rlabel polysilicon 450 -651 450 -651 0 1
rlabel polysilicon 450 -657 450 -657 0 3
rlabel polysilicon 457 -651 457 -651 0 1
rlabel polysilicon 457 -657 457 -657 0 3
rlabel polysilicon 464 -651 464 -651 0 1
rlabel polysilicon 464 -657 464 -657 0 3
rlabel polysilicon 471 -651 471 -651 0 1
rlabel polysilicon 471 -657 471 -657 0 3
rlabel polysilicon 481 -651 481 -651 0 2
rlabel polysilicon 478 -657 478 -657 0 3
rlabel polysilicon 481 -657 481 -657 0 4
rlabel polysilicon 485 -651 485 -651 0 1
rlabel polysilicon 485 -657 485 -657 0 3
rlabel polysilicon 492 -651 492 -651 0 1
rlabel polysilicon 492 -657 492 -657 0 3
rlabel polysilicon 502 -651 502 -651 0 2
rlabel polysilicon 499 -657 499 -657 0 3
rlabel polysilicon 502 -657 502 -657 0 4
rlabel polysilicon 506 -651 506 -651 0 1
rlabel polysilicon 506 -657 506 -657 0 3
rlabel polysilicon 513 -651 513 -651 0 1
rlabel polysilicon 513 -657 513 -657 0 3
rlabel polysilicon 516 -657 516 -657 0 4
rlabel polysilicon 520 -657 520 -657 0 3
rlabel polysilicon 523 -657 523 -657 0 4
rlabel polysilicon 527 -651 527 -651 0 1
rlabel polysilicon 527 -657 527 -657 0 3
rlabel polysilicon 534 -651 534 -651 0 1
rlabel polysilicon 534 -657 534 -657 0 3
rlabel polysilicon 541 -651 541 -651 0 1
rlabel polysilicon 541 -657 541 -657 0 3
rlabel polysilicon 548 -651 548 -651 0 1
rlabel polysilicon 551 -657 551 -657 0 4
rlabel polysilicon 555 -651 555 -651 0 1
rlabel polysilicon 555 -657 555 -657 0 3
rlabel polysilicon 562 -651 562 -651 0 1
rlabel polysilicon 562 -657 562 -657 0 3
rlabel polysilicon 569 -651 569 -651 0 1
rlabel polysilicon 569 -657 569 -657 0 3
rlabel polysilicon 576 -651 576 -651 0 1
rlabel polysilicon 576 -657 576 -657 0 3
rlabel polysilicon 583 -651 583 -651 0 1
rlabel polysilicon 583 -657 583 -657 0 3
rlabel polysilicon 590 -651 590 -651 0 1
rlabel polysilicon 590 -657 590 -657 0 3
rlabel polysilicon 597 -651 597 -651 0 1
rlabel polysilicon 597 -657 597 -657 0 3
rlabel polysilicon 604 -651 604 -651 0 1
rlabel polysilicon 607 -651 607 -651 0 2
rlabel polysilicon 604 -657 604 -657 0 3
rlabel polysilicon 607 -657 607 -657 0 4
rlabel polysilicon 611 -651 611 -651 0 1
rlabel polysilicon 614 -651 614 -651 0 2
rlabel polysilicon 614 -657 614 -657 0 4
rlabel polysilicon 618 -651 618 -651 0 1
rlabel polysilicon 618 -657 618 -657 0 3
rlabel polysilicon 625 -651 625 -651 0 1
rlabel polysilicon 625 -657 625 -657 0 3
rlabel polysilicon 632 -651 632 -651 0 1
rlabel polysilicon 632 -657 632 -657 0 3
rlabel polysilicon 639 -651 639 -651 0 1
rlabel polysilicon 639 -657 639 -657 0 3
rlabel polysilicon 646 -651 646 -651 0 1
rlabel polysilicon 646 -657 646 -657 0 3
rlabel polysilicon 653 -651 653 -651 0 1
rlabel polysilicon 656 -651 656 -651 0 2
rlabel polysilicon 656 -657 656 -657 0 4
rlabel polysilicon 660 -651 660 -651 0 1
rlabel polysilicon 660 -657 660 -657 0 3
rlabel polysilicon 667 -651 667 -651 0 1
rlabel polysilicon 667 -657 667 -657 0 3
rlabel polysilicon 674 -651 674 -651 0 1
rlabel polysilicon 674 -657 674 -657 0 3
rlabel polysilicon 681 -651 681 -651 0 1
rlabel polysilicon 681 -657 681 -657 0 3
rlabel polysilicon 691 -651 691 -651 0 2
rlabel polysilicon 688 -657 688 -657 0 3
rlabel polysilicon 691 -657 691 -657 0 4
rlabel polysilicon 695 -651 695 -651 0 1
rlabel polysilicon 695 -657 695 -657 0 3
rlabel polysilicon 702 -651 702 -651 0 1
rlabel polysilicon 702 -657 702 -657 0 3
rlabel polysilicon 709 -651 709 -651 0 1
rlabel polysilicon 709 -657 709 -657 0 3
rlabel polysilicon 716 -651 716 -651 0 1
rlabel polysilicon 716 -657 716 -657 0 3
rlabel polysilicon 723 -651 723 -651 0 1
rlabel polysilicon 723 -657 723 -657 0 3
rlabel polysilicon 730 -651 730 -651 0 1
rlabel polysilicon 730 -657 730 -657 0 3
rlabel polysilicon 737 -651 737 -651 0 1
rlabel polysilicon 737 -657 737 -657 0 3
rlabel polysilicon 744 -651 744 -651 0 1
rlabel polysilicon 744 -657 744 -657 0 3
rlabel polysilicon 751 -651 751 -651 0 1
rlabel polysilicon 751 -657 751 -657 0 3
rlabel polysilicon 758 -651 758 -651 0 1
rlabel polysilicon 761 -651 761 -651 0 2
rlabel polysilicon 765 -651 765 -651 0 1
rlabel polysilicon 765 -657 765 -657 0 3
rlabel polysilicon 772 -651 772 -651 0 1
rlabel polysilicon 772 -657 772 -657 0 3
rlabel polysilicon 779 -651 779 -651 0 1
rlabel polysilicon 779 -657 779 -657 0 3
rlabel polysilicon 786 -651 786 -651 0 1
rlabel polysilicon 786 -657 786 -657 0 3
rlabel polysilicon 793 -651 793 -651 0 1
rlabel polysilicon 793 -657 793 -657 0 3
rlabel polysilicon 800 -651 800 -651 0 1
rlabel polysilicon 800 -657 800 -657 0 3
rlabel polysilicon 807 -651 807 -651 0 1
rlabel polysilicon 807 -657 807 -657 0 3
rlabel polysilicon 814 -651 814 -651 0 1
rlabel polysilicon 814 -657 814 -657 0 3
rlabel polysilicon 821 -651 821 -651 0 1
rlabel polysilicon 821 -657 821 -657 0 3
rlabel polysilicon 828 -651 828 -651 0 1
rlabel polysilicon 828 -657 828 -657 0 3
rlabel polysilicon 835 -651 835 -651 0 1
rlabel polysilicon 835 -657 835 -657 0 3
rlabel polysilicon 842 -651 842 -651 0 1
rlabel polysilicon 842 -657 842 -657 0 3
rlabel polysilicon 849 -651 849 -651 0 1
rlabel polysilicon 849 -657 849 -657 0 3
rlabel polysilicon 856 -651 856 -651 0 1
rlabel polysilicon 856 -657 856 -657 0 3
rlabel polysilicon 863 -651 863 -651 0 1
rlabel polysilicon 863 -657 863 -657 0 3
rlabel polysilicon 870 -651 870 -651 0 1
rlabel polysilicon 870 -657 870 -657 0 3
rlabel polysilicon 877 -651 877 -651 0 1
rlabel polysilicon 884 -651 884 -651 0 1
rlabel polysilicon 884 -657 884 -657 0 3
rlabel polysilicon 891 -651 891 -651 0 1
rlabel polysilicon 891 -657 891 -657 0 3
rlabel polysilicon 898 -651 898 -651 0 1
rlabel polysilicon 898 -657 898 -657 0 3
rlabel polysilicon 905 -651 905 -651 0 1
rlabel polysilicon 905 -657 905 -657 0 3
rlabel polysilicon 912 -651 912 -651 0 1
rlabel polysilicon 912 -657 912 -657 0 3
rlabel polysilicon 919 -651 919 -651 0 1
rlabel polysilicon 919 -657 919 -657 0 3
rlabel polysilicon 926 -651 926 -651 0 1
rlabel polysilicon 926 -657 926 -657 0 3
rlabel polysilicon 933 -657 933 -657 0 3
rlabel polysilicon 940 -651 940 -651 0 1
rlabel polysilicon 940 -657 940 -657 0 3
rlabel polysilicon 947 -651 947 -651 0 1
rlabel polysilicon 947 -657 947 -657 0 3
rlabel polysilicon 954 -651 954 -651 0 1
rlabel polysilicon 954 -657 954 -657 0 3
rlabel polysilicon 961 -651 961 -651 0 1
rlabel polysilicon 961 -657 961 -657 0 3
rlabel polysilicon 968 -651 968 -651 0 1
rlabel polysilicon 968 -657 968 -657 0 3
rlabel polysilicon 975 -651 975 -651 0 1
rlabel polysilicon 975 -657 975 -657 0 3
rlabel polysilicon 982 -651 982 -651 0 1
rlabel polysilicon 982 -657 982 -657 0 3
rlabel polysilicon 989 -651 989 -651 0 1
rlabel polysilicon 989 -657 989 -657 0 3
rlabel polysilicon 996 -651 996 -651 0 1
rlabel polysilicon 996 -657 996 -657 0 3
rlabel polysilicon 1003 -651 1003 -651 0 1
rlabel polysilicon 1003 -657 1003 -657 0 3
rlabel polysilicon 1006 -657 1006 -657 0 4
rlabel polysilicon 1010 -651 1010 -651 0 1
rlabel polysilicon 1010 -657 1010 -657 0 3
rlabel polysilicon 1017 -651 1017 -651 0 1
rlabel polysilicon 1017 -657 1017 -657 0 3
rlabel polysilicon 1024 -651 1024 -651 0 1
rlabel polysilicon 1024 -657 1024 -657 0 3
rlabel polysilicon 1031 -651 1031 -651 0 1
rlabel polysilicon 1031 -657 1031 -657 0 3
rlabel polysilicon 1038 -651 1038 -651 0 1
rlabel polysilicon 1038 -657 1038 -657 0 3
rlabel polysilicon 1041 -657 1041 -657 0 4
rlabel polysilicon 1045 -651 1045 -651 0 1
rlabel polysilicon 1045 -657 1045 -657 0 3
rlabel polysilicon 1052 -651 1052 -651 0 1
rlabel polysilicon 1052 -657 1052 -657 0 3
rlabel polysilicon 1059 -651 1059 -651 0 1
rlabel polysilicon 1059 -657 1059 -657 0 3
rlabel polysilicon 1066 -651 1066 -651 0 1
rlabel polysilicon 1066 -657 1066 -657 0 3
rlabel polysilicon 1073 -651 1073 -651 0 1
rlabel polysilicon 1073 -657 1073 -657 0 3
rlabel polysilicon 1080 -651 1080 -651 0 1
rlabel polysilicon 1080 -657 1080 -657 0 3
rlabel polysilicon 1087 -651 1087 -651 0 1
rlabel polysilicon 1087 -657 1087 -657 0 3
rlabel polysilicon 1094 -651 1094 -651 0 1
rlabel polysilicon 1094 -657 1094 -657 0 3
rlabel polysilicon 1101 -651 1101 -651 0 1
rlabel polysilicon 1101 -657 1101 -657 0 3
rlabel polysilicon 1108 -651 1108 -651 0 1
rlabel polysilicon 1108 -657 1108 -657 0 3
rlabel polysilicon 1115 -651 1115 -651 0 1
rlabel polysilicon 1115 -657 1115 -657 0 3
rlabel polysilicon 1122 -651 1122 -651 0 1
rlabel polysilicon 1122 -657 1122 -657 0 3
rlabel polysilicon 1129 -651 1129 -651 0 1
rlabel polysilicon 1129 -657 1129 -657 0 3
rlabel polysilicon 1136 -651 1136 -651 0 1
rlabel polysilicon 1136 -657 1136 -657 0 3
rlabel polysilicon 1178 -651 1178 -651 0 1
rlabel polysilicon 1178 -657 1178 -657 0 3
rlabel polysilicon 9 -732 9 -732 0 1
rlabel polysilicon 9 -738 9 -738 0 3
rlabel polysilicon 16 -732 16 -732 0 1
rlabel polysilicon 16 -738 16 -738 0 3
rlabel polysilicon 23 -732 23 -732 0 1
rlabel polysilicon 23 -738 23 -738 0 3
rlabel polysilicon 33 -732 33 -732 0 2
rlabel polysilicon 37 -732 37 -732 0 1
rlabel polysilicon 37 -738 37 -738 0 3
rlabel polysilicon 44 -732 44 -732 0 1
rlabel polysilicon 44 -738 44 -738 0 3
rlabel polysilicon 51 -732 51 -732 0 1
rlabel polysilicon 51 -738 51 -738 0 3
rlabel polysilicon 58 -732 58 -732 0 1
rlabel polysilicon 58 -738 58 -738 0 3
rlabel polysilicon 65 -732 65 -732 0 1
rlabel polysilicon 65 -738 65 -738 0 3
rlabel polysilicon 72 -732 72 -732 0 1
rlabel polysilicon 79 -732 79 -732 0 1
rlabel polysilicon 79 -738 79 -738 0 3
rlabel polysilicon 86 -732 86 -732 0 1
rlabel polysilicon 86 -738 86 -738 0 3
rlabel polysilicon 93 -732 93 -732 0 1
rlabel polysilicon 93 -738 93 -738 0 3
rlabel polysilicon 100 -732 100 -732 0 1
rlabel polysilicon 100 -738 100 -738 0 3
rlabel polysilicon 107 -732 107 -732 0 1
rlabel polysilicon 107 -738 107 -738 0 3
rlabel polysilicon 114 -732 114 -732 0 1
rlabel polysilicon 114 -738 114 -738 0 3
rlabel polysilicon 124 -738 124 -738 0 4
rlabel polysilicon 128 -732 128 -732 0 1
rlabel polysilicon 128 -738 128 -738 0 3
rlabel polysilicon 135 -732 135 -732 0 1
rlabel polysilicon 135 -738 135 -738 0 3
rlabel polysilicon 138 -738 138 -738 0 4
rlabel polysilicon 142 -732 142 -732 0 1
rlabel polysilicon 142 -738 142 -738 0 3
rlabel polysilicon 149 -732 149 -732 0 1
rlabel polysilicon 152 -732 152 -732 0 2
rlabel polysilicon 156 -732 156 -732 0 1
rlabel polysilicon 156 -738 156 -738 0 3
rlabel polysilicon 163 -732 163 -732 0 1
rlabel polysilicon 163 -738 163 -738 0 3
rlabel polysilicon 170 -732 170 -732 0 1
rlabel polysilicon 170 -738 170 -738 0 3
rlabel polysilicon 177 -732 177 -732 0 1
rlabel polysilicon 177 -738 177 -738 0 3
rlabel polysilicon 184 -732 184 -732 0 1
rlabel polysilicon 187 -738 187 -738 0 4
rlabel polysilicon 191 -732 191 -732 0 1
rlabel polysilicon 191 -738 191 -738 0 3
rlabel polysilicon 198 -732 198 -732 0 1
rlabel polysilicon 198 -738 198 -738 0 3
rlabel polysilicon 205 -732 205 -732 0 1
rlabel polysilicon 208 -732 208 -732 0 2
rlabel polysilicon 212 -732 212 -732 0 1
rlabel polysilicon 212 -738 212 -738 0 3
rlabel polysilicon 219 -732 219 -732 0 1
rlabel polysilicon 219 -738 219 -738 0 3
rlabel polysilicon 226 -732 226 -732 0 1
rlabel polysilicon 226 -738 226 -738 0 3
rlabel polysilicon 233 -732 233 -732 0 1
rlabel polysilicon 233 -738 233 -738 0 3
rlabel polysilicon 240 -732 240 -732 0 1
rlabel polysilicon 240 -738 240 -738 0 3
rlabel polysilicon 247 -738 247 -738 0 3
rlabel polysilicon 254 -732 254 -732 0 1
rlabel polysilicon 254 -738 254 -738 0 3
rlabel polysilicon 261 -732 261 -732 0 1
rlabel polysilicon 261 -738 261 -738 0 3
rlabel polysilicon 268 -732 268 -732 0 1
rlabel polysilicon 268 -738 268 -738 0 3
rlabel polysilicon 275 -732 275 -732 0 1
rlabel polysilicon 275 -738 275 -738 0 3
rlabel polysilicon 282 -732 282 -732 0 1
rlabel polysilicon 282 -738 282 -738 0 3
rlabel polysilicon 289 -732 289 -732 0 1
rlabel polysilicon 289 -738 289 -738 0 3
rlabel polysilicon 296 -732 296 -732 0 1
rlabel polysilicon 296 -738 296 -738 0 3
rlabel polysilicon 303 -732 303 -732 0 1
rlabel polysilicon 303 -738 303 -738 0 3
rlabel polysilicon 310 -738 310 -738 0 3
rlabel polysilicon 317 -732 317 -732 0 1
rlabel polysilicon 317 -738 317 -738 0 3
rlabel polysilicon 324 -732 324 -732 0 1
rlabel polysilicon 324 -738 324 -738 0 3
rlabel polysilicon 331 -732 331 -732 0 1
rlabel polysilicon 331 -738 331 -738 0 3
rlabel polysilicon 338 -732 338 -732 0 1
rlabel polysilicon 341 -732 341 -732 0 2
rlabel polysilicon 338 -738 338 -738 0 3
rlabel polysilicon 341 -738 341 -738 0 4
rlabel polysilicon 345 -732 345 -732 0 1
rlabel polysilicon 345 -738 345 -738 0 3
rlabel polysilicon 352 -732 352 -732 0 1
rlabel polysilicon 352 -738 352 -738 0 3
rlabel polysilicon 359 -738 359 -738 0 3
rlabel polysilicon 362 -738 362 -738 0 4
rlabel polysilicon 366 -732 366 -732 0 1
rlabel polysilicon 366 -738 366 -738 0 3
rlabel polysilicon 373 -732 373 -732 0 1
rlabel polysilicon 373 -738 373 -738 0 3
rlabel polysilicon 380 -732 380 -732 0 1
rlabel polysilicon 380 -738 380 -738 0 3
rlabel polysilicon 387 -732 387 -732 0 1
rlabel polysilicon 387 -738 387 -738 0 3
rlabel polysilicon 394 -732 394 -732 0 1
rlabel polysilicon 397 -732 397 -732 0 2
rlabel polysilicon 394 -738 394 -738 0 3
rlabel polysilicon 404 -738 404 -738 0 4
rlabel polysilicon 411 -732 411 -732 0 2
rlabel polysilicon 411 -738 411 -738 0 4
rlabel polysilicon 415 -732 415 -732 0 1
rlabel polysilicon 415 -738 415 -738 0 3
rlabel polysilicon 425 -732 425 -732 0 2
rlabel polysilicon 425 -738 425 -738 0 4
rlabel polysilicon 429 -732 429 -732 0 1
rlabel polysilicon 429 -738 429 -738 0 3
rlabel polysilicon 439 -732 439 -732 0 2
rlabel polysilicon 439 -738 439 -738 0 4
rlabel polysilicon 443 -732 443 -732 0 1
rlabel polysilicon 443 -738 443 -738 0 3
rlabel polysilicon 450 -732 450 -732 0 1
rlabel polysilicon 450 -738 450 -738 0 3
rlabel polysilicon 457 -732 457 -732 0 1
rlabel polysilicon 457 -738 457 -738 0 3
rlabel polysilicon 464 -732 464 -732 0 1
rlabel polysilicon 467 -732 467 -732 0 2
rlabel polysilicon 474 -732 474 -732 0 2
rlabel polysilicon 474 -738 474 -738 0 4
rlabel polysilicon 478 -732 478 -732 0 1
rlabel polysilicon 478 -738 478 -738 0 3
rlabel polysilicon 485 -732 485 -732 0 1
rlabel polysilicon 485 -738 485 -738 0 3
rlabel polysilicon 492 -732 492 -732 0 1
rlabel polysilicon 492 -738 492 -738 0 3
rlabel polysilicon 499 -732 499 -732 0 1
rlabel polysilicon 499 -738 499 -738 0 3
rlabel polysilicon 506 -732 506 -732 0 1
rlabel polysilicon 506 -738 506 -738 0 3
rlabel polysilicon 513 -732 513 -732 0 1
rlabel polysilicon 513 -738 513 -738 0 3
rlabel polysilicon 523 -732 523 -732 0 2
rlabel polysilicon 520 -738 520 -738 0 3
rlabel polysilicon 523 -738 523 -738 0 4
rlabel polysilicon 527 -732 527 -732 0 1
rlabel polysilicon 527 -738 527 -738 0 3
rlabel polysilicon 534 -732 534 -732 0 1
rlabel polysilicon 534 -738 534 -738 0 3
rlabel polysilicon 541 -732 541 -732 0 1
rlabel polysilicon 541 -738 541 -738 0 3
rlabel polysilicon 548 -732 548 -732 0 1
rlabel polysilicon 551 -732 551 -732 0 2
rlabel polysilicon 548 -738 548 -738 0 3
rlabel polysilicon 555 -732 555 -732 0 1
rlabel polysilicon 555 -738 555 -738 0 3
rlabel polysilicon 562 -732 562 -732 0 1
rlabel polysilicon 562 -738 562 -738 0 3
rlabel polysilicon 569 -732 569 -732 0 1
rlabel polysilicon 569 -738 569 -738 0 3
rlabel polysilicon 576 -732 576 -732 0 1
rlabel polysilicon 576 -738 576 -738 0 3
rlabel polysilicon 583 -732 583 -732 0 1
rlabel polysilicon 583 -738 583 -738 0 3
rlabel polysilicon 590 -732 590 -732 0 1
rlabel polysilicon 590 -738 590 -738 0 3
rlabel polysilicon 597 -732 597 -732 0 1
rlabel polysilicon 597 -738 597 -738 0 3
rlabel polysilicon 600 -738 600 -738 0 4
rlabel polysilicon 604 -732 604 -732 0 1
rlabel polysilicon 604 -738 604 -738 0 3
rlabel polysilicon 611 -732 611 -732 0 1
rlabel polysilicon 611 -738 611 -738 0 3
rlabel polysilicon 618 -732 618 -732 0 1
rlabel polysilicon 618 -738 618 -738 0 3
rlabel polysilicon 625 -732 625 -732 0 1
rlabel polysilicon 625 -738 625 -738 0 3
rlabel polysilicon 635 -732 635 -732 0 2
rlabel polysilicon 632 -738 632 -738 0 3
rlabel polysilicon 635 -738 635 -738 0 4
rlabel polysilicon 639 -732 639 -732 0 1
rlabel polysilicon 642 -738 642 -738 0 4
rlabel polysilicon 646 -732 646 -732 0 1
rlabel polysilicon 646 -738 646 -738 0 3
rlabel polysilicon 653 -732 653 -732 0 1
rlabel polysilicon 653 -738 653 -738 0 3
rlabel polysilicon 660 -732 660 -732 0 1
rlabel polysilicon 660 -738 660 -738 0 3
rlabel polysilicon 667 -732 667 -732 0 1
rlabel polysilicon 667 -738 667 -738 0 3
rlabel polysilicon 674 -732 674 -732 0 1
rlabel polysilicon 674 -738 674 -738 0 3
rlabel polysilicon 681 -732 681 -732 0 1
rlabel polysilicon 681 -738 681 -738 0 3
rlabel polysilicon 688 -732 688 -732 0 1
rlabel polysilicon 691 -732 691 -732 0 2
rlabel polysilicon 688 -738 688 -738 0 3
rlabel polysilicon 695 -732 695 -732 0 1
rlabel polysilicon 695 -738 695 -738 0 3
rlabel polysilicon 702 -732 702 -732 0 1
rlabel polysilicon 702 -738 702 -738 0 3
rlabel polysilicon 709 -732 709 -732 0 1
rlabel polysilicon 709 -738 709 -738 0 3
rlabel polysilicon 716 -732 716 -732 0 1
rlabel polysilicon 716 -738 716 -738 0 3
rlabel polysilicon 723 -732 723 -732 0 1
rlabel polysilicon 723 -738 723 -738 0 3
rlabel polysilicon 730 -732 730 -732 0 1
rlabel polysilicon 730 -738 730 -738 0 3
rlabel polysilicon 737 -732 737 -732 0 1
rlabel polysilicon 737 -738 737 -738 0 3
rlabel polysilicon 744 -732 744 -732 0 1
rlabel polysilicon 747 -732 747 -732 0 2
rlabel polysilicon 744 -738 744 -738 0 3
rlabel polysilicon 747 -738 747 -738 0 4
rlabel polysilicon 751 -732 751 -732 0 1
rlabel polysilicon 751 -738 751 -738 0 3
rlabel polysilicon 758 -732 758 -732 0 1
rlabel polysilicon 758 -738 758 -738 0 3
rlabel polysilicon 765 -732 765 -732 0 1
rlabel polysilicon 765 -738 765 -738 0 3
rlabel polysilicon 772 -732 772 -732 0 1
rlabel polysilicon 772 -738 772 -738 0 3
rlabel polysilicon 779 -732 779 -732 0 1
rlabel polysilicon 779 -738 779 -738 0 3
rlabel polysilicon 786 -732 786 -732 0 1
rlabel polysilicon 786 -738 786 -738 0 3
rlabel polysilicon 793 -732 793 -732 0 1
rlabel polysilicon 793 -738 793 -738 0 3
rlabel polysilicon 800 -732 800 -732 0 1
rlabel polysilicon 800 -738 800 -738 0 3
rlabel polysilicon 807 -732 807 -732 0 1
rlabel polysilicon 807 -738 807 -738 0 3
rlabel polysilicon 814 -732 814 -732 0 1
rlabel polysilicon 814 -738 814 -738 0 3
rlabel polysilicon 821 -732 821 -732 0 1
rlabel polysilicon 821 -738 821 -738 0 3
rlabel polysilicon 828 -732 828 -732 0 1
rlabel polysilicon 828 -738 828 -738 0 3
rlabel polysilicon 835 -732 835 -732 0 1
rlabel polysilicon 835 -738 835 -738 0 3
rlabel polysilicon 842 -732 842 -732 0 1
rlabel polysilicon 842 -738 842 -738 0 3
rlabel polysilicon 849 -732 849 -732 0 1
rlabel polysilicon 849 -738 849 -738 0 3
rlabel polysilicon 856 -732 856 -732 0 1
rlabel polysilicon 856 -738 856 -738 0 3
rlabel polysilicon 863 -732 863 -732 0 1
rlabel polysilicon 863 -738 863 -738 0 3
rlabel polysilicon 870 -732 870 -732 0 1
rlabel polysilicon 870 -738 870 -738 0 3
rlabel polysilicon 877 -738 877 -738 0 3
rlabel polysilicon 884 -732 884 -732 0 1
rlabel polysilicon 884 -738 884 -738 0 3
rlabel polysilicon 891 -732 891 -732 0 1
rlabel polysilicon 891 -738 891 -738 0 3
rlabel polysilicon 898 -732 898 -732 0 1
rlabel polysilicon 898 -738 898 -738 0 3
rlabel polysilicon 905 -732 905 -732 0 1
rlabel polysilicon 905 -738 905 -738 0 3
rlabel polysilicon 912 -732 912 -732 0 1
rlabel polysilicon 912 -738 912 -738 0 3
rlabel polysilicon 919 -732 919 -732 0 1
rlabel polysilicon 919 -738 919 -738 0 3
rlabel polysilicon 926 -732 926 -732 0 1
rlabel polysilicon 926 -738 926 -738 0 3
rlabel polysilicon 933 -732 933 -732 0 1
rlabel polysilicon 933 -738 933 -738 0 3
rlabel polysilicon 940 -732 940 -732 0 1
rlabel polysilicon 940 -738 940 -738 0 3
rlabel polysilicon 947 -732 947 -732 0 1
rlabel polysilicon 947 -738 947 -738 0 3
rlabel polysilicon 954 -732 954 -732 0 1
rlabel polysilicon 954 -738 954 -738 0 3
rlabel polysilicon 961 -732 961 -732 0 1
rlabel polysilicon 961 -738 961 -738 0 3
rlabel polysilicon 968 -732 968 -732 0 1
rlabel polysilicon 968 -738 968 -738 0 3
rlabel polysilicon 975 -732 975 -732 0 1
rlabel polysilicon 975 -738 975 -738 0 3
rlabel polysilicon 982 -732 982 -732 0 1
rlabel polysilicon 982 -738 982 -738 0 3
rlabel polysilicon 989 -732 989 -732 0 1
rlabel polysilicon 989 -738 989 -738 0 3
rlabel polysilicon 996 -732 996 -732 0 1
rlabel polysilicon 996 -738 996 -738 0 3
rlabel polysilicon 1003 -732 1003 -732 0 1
rlabel polysilicon 1006 -732 1006 -732 0 2
rlabel polysilicon 1003 -738 1003 -738 0 3
rlabel polysilicon 1010 -732 1010 -732 0 1
rlabel polysilicon 1010 -738 1010 -738 0 3
rlabel polysilicon 1017 -732 1017 -732 0 1
rlabel polysilicon 1017 -738 1017 -738 0 3
rlabel polysilicon 1024 -732 1024 -732 0 1
rlabel polysilicon 1024 -738 1024 -738 0 3
rlabel polysilicon 1031 -732 1031 -732 0 1
rlabel polysilicon 1031 -738 1031 -738 0 3
rlabel polysilicon 1038 -732 1038 -732 0 1
rlabel polysilicon 1041 -732 1041 -732 0 2
rlabel polysilicon 1038 -738 1038 -738 0 3
rlabel polysilicon 1045 -732 1045 -732 0 1
rlabel polysilicon 1045 -738 1045 -738 0 3
rlabel polysilicon 1052 -732 1052 -732 0 1
rlabel polysilicon 1052 -738 1052 -738 0 3
rlabel polysilicon 1059 -732 1059 -732 0 1
rlabel polysilicon 1059 -738 1059 -738 0 3
rlabel polysilicon 1066 -732 1066 -732 0 1
rlabel polysilicon 1066 -738 1066 -738 0 3
rlabel polysilicon 1073 -732 1073 -732 0 1
rlabel polysilicon 1073 -738 1073 -738 0 3
rlabel polysilicon 1080 -732 1080 -732 0 1
rlabel polysilicon 1080 -738 1080 -738 0 3
rlabel polysilicon 1087 -732 1087 -732 0 1
rlabel polysilicon 1090 -732 1090 -732 0 2
rlabel polysilicon 1087 -738 1087 -738 0 3
rlabel polysilicon 1090 -738 1090 -738 0 4
rlabel polysilicon 1094 -732 1094 -732 0 1
rlabel polysilicon 1094 -738 1094 -738 0 3
rlabel polysilicon 1101 -732 1101 -732 0 1
rlabel polysilicon 1101 -738 1101 -738 0 3
rlabel polysilicon 1108 -732 1108 -732 0 1
rlabel polysilicon 1111 -732 1111 -732 0 2
rlabel polysilicon 1108 -738 1108 -738 0 3
rlabel polysilicon 1115 -732 1115 -732 0 1
rlabel polysilicon 1115 -738 1115 -738 0 3
rlabel polysilicon 1122 -732 1122 -732 0 1
rlabel polysilicon 1122 -738 1122 -738 0 3
rlabel polysilicon 1129 -732 1129 -732 0 1
rlabel polysilicon 1129 -738 1129 -738 0 3
rlabel polysilicon 1136 -732 1136 -732 0 1
rlabel polysilicon 1136 -738 1136 -738 0 3
rlabel polysilicon 1143 -732 1143 -732 0 1
rlabel polysilicon 1143 -738 1143 -738 0 3
rlabel polysilicon 1150 -732 1150 -732 0 1
rlabel polysilicon 1150 -738 1150 -738 0 3
rlabel polysilicon 1157 -738 1157 -738 0 3
rlabel polysilicon 1160 -738 1160 -738 0 4
rlabel polysilicon 1164 -732 1164 -732 0 1
rlabel polysilicon 1164 -738 1164 -738 0 3
rlabel polysilicon 1171 -732 1171 -732 0 1
rlabel polysilicon 1171 -738 1171 -738 0 3
rlabel polysilicon 1185 -732 1185 -732 0 1
rlabel polysilicon 1185 -738 1185 -738 0 3
rlabel polysilicon 9 -821 9 -821 0 1
rlabel polysilicon 9 -827 9 -827 0 3
rlabel polysilicon 16 -821 16 -821 0 1
rlabel polysilicon 16 -827 16 -827 0 3
rlabel polysilicon 23 -821 23 -821 0 1
rlabel polysilicon 23 -827 23 -827 0 3
rlabel polysilicon 30 -821 30 -821 0 1
rlabel polysilicon 30 -827 30 -827 0 3
rlabel polysilicon 37 -821 37 -821 0 1
rlabel polysilicon 37 -827 37 -827 0 3
rlabel polysilicon 44 -821 44 -821 0 1
rlabel polysilicon 44 -827 44 -827 0 3
rlabel polysilicon 51 -821 51 -821 0 1
rlabel polysilicon 51 -827 51 -827 0 3
rlabel polysilicon 58 -821 58 -821 0 1
rlabel polysilicon 58 -827 58 -827 0 3
rlabel polysilicon 65 -821 65 -821 0 1
rlabel polysilicon 65 -827 65 -827 0 3
rlabel polysilicon 72 -827 72 -827 0 3
rlabel polysilicon 79 -821 79 -821 0 1
rlabel polysilicon 79 -827 79 -827 0 3
rlabel polysilicon 86 -821 86 -821 0 1
rlabel polysilicon 86 -827 86 -827 0 3
rlabel polysilicon 93 -821 93 -821 0 1
rlabel polysilicon 93 -827 93 -827 0 3
rlabel polysilicon 100 -821 100 -821 0 1
rlabel polysilicon 107 -821 107 -821 0 1
rlabel polysilicon 107 -827 107 -827 0 3
rlabel polysilicon 117 -821 117 -821 0 2
rlabel polysilicon 114 -827 114 -827 0 3
rlabel polysilicon 117 -827 117 -827 0 4
rlabel polysilicon 121 -821 121 -821 0 1
rlabel polysilicon 121 -827 121 -827 0 3
rlabel polysilicon 124 -827 124 -827 0 4
rlabel polysilicon 131 -821 131 -821 0 2
rlabel polysilicon 128 -827 128 -827 0 3
rlabel polysilicon 135 -821 135 -821 0 1
rlabel polysilicon 138 -821 138 -821 0 2
rlabel polysilicon 142 -821 142 -821 0 1
rlabel polysilicon 142 -827 142 -827 0 3
rlabel polysilicon 149 -821 149 -821 0 1
rlabel polysilicon 149 -827 149 -827 0 3
rlabel polysilicon 156 -821 156 -821 0 1
rlabel polysilicon 156 -827 156 -827 0 3
rlabel polysilicon 163 -821 163 -821 0 1
rlabel polysilicon 163 -827 163 -827 0 3
rlabel polysilicon 170 -821 170 -821 0 1
rlabel polysilicon 173 -821 173 -821 0 2
rlabel polysilicon 177 -821 177 -821 0 1
rlabel polysilicon 177 -827 177 -827 0 3
rlabel polysilicon 184 -821 184 -821 0 1
rlabel polysilicon 184 -827 184 -827 0 3
rlabel polysilicon 191 -821 191 -821 0 1
rlabel polysilicon 191 -827 191 -827 0 3
rlabel polysilicon 198 -821 198 -821 0 1
rlabel polysilicon 198 -827 198 -827 0 3
rlabel polysilicon 205 -821 205 -821 0 1
rlabel polysilicon 205 -827 205 -827 0 3
rlabel polysilicon 212 -821 212 -821 0 1
rlabel polysilicon 212 -827 212 -827 0 3
rlabel polysilicon 219 -821 219 -821 0 1
rlabel polysilicon 219 -827 219 -827 0 3
rlabel polysilicon 226 -821 226 -821 0 1
rlabel polysilicon 226 -827 226 -827 0 3
rlabel polysilicon 233 -821 233 -821 0 1
rlabel polysilicon 233 -827 233 -827 0 3
rlabel polysilicon 240 -821 240 -821 0 1
rlabel polysilicon 240 -827 240 -827 0 3
rlabel polysilicon 247 -821 247 -821 0 1
rlabel polysilicon 247 -827 247 -827 0 3
rlabel polysilicon 254 -821 254 -821 0 1
rlabel polysilicon 254 -827 254 -827 0 3
rlabel polysilicon 268 -821 268 -821 0 1
rlabel polysilicon 268 -827 268 -827 0 3
rlabel polysilicon 275 -821 275 -821 0 1
rlabel polysilicon 275 -827 275 -827 0 3
rlabel polysilicon 282 -821 282 -821 0 1
rlabel polysilicon 282 -827 282 -827 0 3
rlabel polysilicon 289 -821 289 -821 0 1
rlabel polysilicon 289 -827 289 -827 0 3
rlabel polysilicon 296 -821 296 -821 0 1
rlabel polysilicon 296 -827 296 -827 0 3
rlabel polysilicon 303 -821 303 -821 0 1
rlabel polysilicon 303 -827 303 -827 0 3
rlabel polysilicon 310 -821 310 -821 0 1
rlabel polysilicon 310 -827 310 -827 0 3
rlabel polysilicon 317 -821 317 -821 0 1
rlabel polysilicon 317 -827 317 -827 0 3
rlabel polysilicon 324 -821 324 -821 0 1
rlabel polysilicon 324 -827 324 -827 0 3
rlabel polysilicon 331 -821 331 -821 0 1
rlabel polysilicon 331 -827 331 -827 0 3
rlabel polysilicon 338 -821 338 -821 0 1
rlabel polysilicon 338 -827 338 -827 0 3
rlabel polysilicon 345 -821 345 -821 0 1
rlabel polysilicon 345 -827 345 -827 0 3
rlabel polysilicon 352 -821 352 -821 0 1
rlabel polysilicon 352 -827 352 -827 0 3
rlabel polysilicon 355 -827 355 -827 0 4
rlabel polysilicon 362 -827 362 -827 0 4
rlabel polysilicon 366 -821 366 -821 0 1
rlabel polysilicon 366 -827 366 -827 0 3
rlabel polysilicon 373 -821 373 -821 0 1
rlabel polysilicon 373 -827 373 -827 0 3
rlabel polysilicon 380 -821 380 -821 0 1
rlabel polysilicon 383 -821 383 -821 0 2
rlabel polysilicon 380 -827 380 -827 0 3
rlabel polysilicon 383 -827 383 -827 0 4
rlabel polysilicon 387 -821 387 -821 0 1
rlabel polysilicon 387 -827 387 -827 0 3
rlabel polysilicon 394 -821 394 -821 0 1
rlabel polysilicon 394 -827 394 -827 0 3
rlabel polysilicon 401 -821 401 -821 0 1
rlabel polysilicon 401 -827 401 -827 0 3
rlabel polysilicon 408 -821 408 -821 0 1
rlabel polysilicon 408 -827 408 -827 0 3
rlabel polysilicon 415 -821 415 -821 0 1
rlabel polysilicon 415 -827 415 -827 0 3
rlabel polysilicon 425 -821 425 -821 0 2
rlabel polysilicon 422 -827 422 -827 0 3
rlabel polysilicon 425 -827 425 -827 0 4
rlabel polysilicon 429 -821 429 -821 0 1
rlabel polysilicon 429 -827 429 -827 0 3
rlabel polysilicon 436 -821 436 -821 0 1
rlabel polysilicon 436 -827 436 -827 0 3
rlabel polysilicon 443 -821 443 -821 0 1
rlabel polysilicon 443 -827 443 -827 0 3
rlabel polysilicon 450 -821 450 -821 0 1
rlabel polysilicon 450 -827 450 -827 0 3
rlabel polysilicon 457 -821 457 -821 0 1
rlabel polysilicon 457 -827 457 -827 0 3
rlabel polysilicon 464 -821 464 -821 0 1
rlabel polysilicon 464 -827 464 -827 0 3
rlabel polysilicon 471 -821 471 -821 0 1
rlabel polysilicon 471 -827 471 -827 0 3
rlabel polysilicon 478 -821 478 -821 0 1
rlabel polysilicon 485 -821 485 -821 0 1
rlabel polysilicon 485 -827 485 -827 0 3
rlabel polysilicon 495 -821 495 -821 0 2
rlabel polysilicon 492 -827 492 -827 0 3
rlabel polysilicon 495 -827 495 -827 0 4
rlabel polysilicon 499 -821 499 -821 0 1
rlabel polysilicon 502 -821 502 -821 0 2
rlabel polysilicon 502 -827 502 -827 0 4
rlabel polysilicon 506 -821 506 -821 0 1
rlabel polysilicon 506 -827 506 -827 0 3
rlabel polysilicon 513 -821 513 -821 0 1
rlabel polysilicon 513 -827 513 -827 0 3
rlabel polysilicon 520 -821 520 -821 0 1
rlabel polysilicon 523 -827 523 -827 0 4
rlabel polysilicon 527 -821 527 -821 0 1
rlabel polysilicon 527 -827 527 -827 0 3
rlabel polysilicon 534 -821 534 -821 0 1
rlabel polysilicon 534 -827 534 -827 0 3
rlabel polysilicon 541 -821 541 -821 0 1
rlabel polysilicon 541 -827 541 -827 0 3
rlabel polysilicon 548 -821 548 -821 0 1
rlabel polysilicon 548 -827 548 -827 0 3
rlabel polysilicon 555 -821 555 -821 0 1
rlabel polysilicon 555 -827 555 -827 0 3
rlabel polysilicon 558 -827 558 -827 0 4
rlabel polysilicon 562 -821 562 -821 0 1
rlabel polysilicon 565 -821 565 -821 0 2
rlabel polysilicon 569 -821 569 -821 0 1
rlabel polysilicon 572 -821 572 -821 0 2
rlabel polysilicon 569 -827 569 -827 0 3
rlabel polysilicon 576 -821 576 -821 0 1
rlabel polysilicon 576 -827 576 -827 0 3
rlabel polysilicon 583 -821 583 -821 0 1
rlabel polysilicon 583 -827 583 -827 0 3
rlabel polysilicon 590 -821 590 -821 0 1
rlabel polysilicon 590 -827 590 -827 0 3
rlabel polysilicon 597 -821 597 -821 0 1
rlabel polysilicon 597 -827 597 -827 0 3
rlabel polysilicon 604 -821 604 -821 0 1
rlabel polysilicon 604 -827 604 -827 0 3
rlabel polysilicon 611 -821 611 -821 0 1
rlabel polysilicon 611 -827 611 -827 0 3
rlabel polysilicon 621 -821 621 -821 0 2
rlabel polysilicon 618 -827 618 -827 0 3
rlabel polysilicon 621 -827 621 -827 0 4
rlabel polysilicon 625 -821 625 -821 0 1
rlabel polysilicon 632 -821 632 -821 0 1
rlabel polysilicon 632 -827 632 -827 0 3
rlabel polysilicon 639 -821 639 -821 0 1
rlabel polysilicon 642 -821 642 -821 0 2
rlabel polysilicon 646 -821 646 -821 0 1
rlabel polysilicon 646 -827 646 -827 0 3
rlabel polysilicon 656 -821 656 -821 0 2
rlabel polysilicon 656 -827 656 -827 0 4
rlabel polysilicon 660 -821 660 -821 0 1
rlabel polysilicon 663 -821 663 -821 0 2
rlabel polysilicon 663 -827 663 -827 0 4
rlabel polysilicon 667 -821 667 -821 0 1
rlabel polysilicon 667 -827 667 -827 0 3
rlabel polysilicon 674 -821 674 -821 0 1
rlabel polysilicon 674 -827 674 -827 0 3
rlabel polysilicon 681 -821 681 -821 0 1
rlabel polysilicon 681 -827 681 -827 0 3
rlabel polysilicon 688 -821 688 -821 0 1
rlabel polysilicon 688 -827 688 -827 0 3
rlabel polysilicon 695 -821 695 -821 0 1
rlabel polysilicon 698 -821 698 -821 0 2
rlabel polysilicon 695 -827 695 -827 0 3
rlabel polysilicon 698 -827 698 -827 0 4
rlabel polysilicon 702 -821 702 -821 0 1
rlabel polysilicon 702 -827 702 -827 0 3
rlabel polysilicon 709 -821 709 -821 0 1
rlabel polysilicon 709 -827 709 -827 0 3
rlabel polysilicon 716 -821 716 -821 0 1
rlabel polysilicon 716 -827 716 -827 0 3
rlabel polysilicon 723 -821 723 -821 0 1
rlabel polysilicon 726 -827 726 -827 0 4
rlabel polysilicon 730 -821 730 -821 0 1
rlabel polysilicon 730 -827 730 -827 0 3
rlabel polysilicon 737 -821 737 -821 0 1
rlabel polysilicon 737 -827 737 -827 0 3
rlabel polysilicon 744 -821 744 -821 0 1
rlabel polysilicon 744 -827 744 -827 0 3
rlabel polysilicon 751 -821 751 -821 0 1
rlabel polysilicon 751 -827 751 -827 0 3
rlabel polysilicon 758 -821 758 -821 0 1
rlabel polysilicon 758 -827 758 -827 0 3
rlabel polysilicon 765 -821 765 -821 0 1
rlabel polysilicon 765 -827 765 -827 0 3
rlabel polysilicon 772 -821 772 -821 0 1
rlabel polysilicon 772 -827 772 -827 0 3
rlabel polysilicon 779 -821 779 -821 0 1
rlabel polysilicon 782 -821 782 -821 0 2
rlabel polysilicon 786 -821 786 -821 0 1
rlabel polysilicon 786 -827 786 -827 0 3
rlabel polysilicon 793 -821 793 -821 0 1
rlabel polysilicon 793 -827 793 -827 0 3
rlabel polysilicon 800 -821 800 -821 0 1
rlabel polysilicon 800 -827 800 -827 0 3
rlabel polysilicon 807 -821 807 -821 0 1
rlabel polysilicon 807 -827 807 -827 0 3
rlabel polysilicon 817 -821 817 -821 0 2
rlabel polysilicon 814 -827 814 -827 0 3
rlabel polysilicon 817 -827 817 -827 0 4
rlabel polysilicon 821 -821 821 -821 0 1
rlabel polysilicon 821 -827 821 -827 0 3
rlabel polysilicon 828 -821 828 -821 0 1
rlabel polysilicon 828 -827 828 -827 0 3
rlabel polysilicon 835 -821 835 -821 0 1
rlabel polysilicon 835 -827 835 -827 0 3
rlabel polysilicon 842 -821 842 -821 0 1
rlabel polysilicon 842 -827 842 -827 0 3
rlabel polysilicon 849 -821 849 -821 0 1
rlabel polysilicon 852 -821 852 -821 0 2
rlabel polysilicon 856 -821 856 -821 0 1
rlabel polysilicon 856 -827 856 -827 0 3
rlabel polysilicon 863 -821 863 -821 0 1
rlabel polysilicon 863 -827 863 -827 0 3
rlabel polysilicon 870 -821 870 -821 0 1
rlabel polysilicon 870 -827 870 -827 0 3
rlabel polysilicon 877 -821 877 -821 0 1
rlabel polysilicon 877 -827 877 -827 0 3
rlabel polysilicon 884 -821 884 -821 0 1
rlabel polysilicon 884 -827 884 -827 0 3
rlabel polysilicon 891 -821 891 -821 0 1
rlabel polysilicon 891 -827 891 -827 0 3
rlabel polysilicon 898 -821 898 -821 0 1
rlabel polysilicon 898 -827 898 -827 0 3
rlabel polysilicon 905 -821 905 -821 0 1
rlabel polysilicon 905 -827 905 -827 0 3
rlabel polysilicon 912 -821 912 -821 0 1
rlabel polysilicon 912 -827 912 -827 0 3
rlabel polysilicon 919 -821 919 -821 0 1
rlabel polysilicon 919 -827 919 -827 0 3
rlabel polysilicon 926 -821 926 -821 0 1
rlabel polysilicon 926 -827 926 -827 0 3
rlabel polysilicon 933 -821 933 -821 0 1
rlabel polysilicon 933 -827 933 -827 0 3
rlabel polysilicon 940 -821 940 -821 0 1
rlabel polysilicon 940 -827 940 -827 0 3
rlabel polysilicon 947 -821 947 -821 0 1
rlabel polysilicon 947 -827 947 -827 0 3
rlabel polysilicon 954 -821 954 -821 0 1
rlabel polysilicon 954 -827 954 -827 0 3
rlabel polysilicon 961 -821 961 -821 0 1
rlabel polysilicon 961 -827 961 -827 0 3
rlabel polysilicon 968 -821 968 -821 0 1
rlabel polysilicon 968 -827 968 -827 0 3
rlabel polysilicon 975 -821 975 -821 0 1
rlabel polysilicon 975 -827 975 -827 0 3
rlabel polysilicon 982 -821 982 -821 0 1
rlabel polysilicon 982 -827 982 -827 0 3
rlabel polysilicon 989 -821 989 -821 0 1
rlabel polysilicon 989 -827 989 -827 0 3
rlabel polysilicon 996 -821 996 -821 0 1
rlabel polysilicon 996 -827 996 -827 0 3
rlabel polysilicon 999 -827 999 -827 0 4
rlabel polysilicon 1003 -821 1003 -821 0 1
rlabel polysilicon 1003 -827 1003 -827 0 3
rlabel polysilicon 1010 -821 1010 -821 0 1
rlabel polysilicon 1010 -827 1010 -827 0 3
rlabel polysilicon 1017 -821 1017 -821 0 1
rlabel polysilicon 1017 -827 1017 -827 0 3
rlabel polysilicon 1024 -821 1024 -821 0 1
rlabel polysilicon 1024 -827 1024 -827 0 3
rlabel polysilicon 1031 -821 1031 -821 0 1
rlabel polysilicon 1031 -827 1031 -827 0 3
rlabel polysilicon 1038 -821 1038 -821 0 1
rlabel polysilicon 1038 -827 1038 -827 0 3
rlabel polysilicon 1045 -821 1045 -821 0 1
rlabel polysilicon 1045 -827 1045 -827 0 3
rlabel polysilicon 1052 -821 1052 -821 0 1
rlabel polysilicon 1052 -827 1052 -827 0 3
rlabel polysilicon 1059 -821 1059 -821 0 1
rlabel polysilicon 1059 -827 1059 -827 0 3
rlabel polysilicon 1066 -821 1066 -821 0 1
rlabel polysilicon 1066 -827 1066 -827 0 3
rlabel polysilicon 1073 -821 1073 -821 0 1
rlabel polysilicon 1073 -827 1073 -827 0 3
rlabel polysilicon 1080 -821 1080 -821 0 1
rlabel polysilicon 1080 -827 1080 -827 0 3
rlabel polysilicon 1087 -821 1087 -821 0 1
rlabel polysilicon 1087 -827 1087 -827 0 3
rlabel polysilicon 1094 -821 1094 -821 0 1
rlabel polysilicon 1094 -827 1094 -827 0 3
rlabel polysilicon 1101 -821 1101 -821 0 1
rlabel polysilicon 1101 -827 1101 -827 0 3
rlabel polysilicon 1108 -821 1108 -821 0 1
rlabel polysilicon 1108 -827 1108 -827 0 3
rlabel polysilicon 1115 -821 1115 -821 0 1
rlabel polysilicon 1115 -827 1115 -827 0 3
rlabel polysilicon 1122 -821 1122 -821 0 1
rlabel polysilicon 1122 -827 1122 -827 0 3
rlabel polysilicon 1129 -821 1129 -821 0 1
rlabel polysilicon 1129 -827 1129 -827 0 3
rlabel polysilicon 1136 -821 1136 -821 0 1
rlabel polysilicon 1136 -827 1136 -827 0 3
rlabel polysilicon 1143 -821 1143 -821 0 1
rlabel polysilicon 1143 -827 1143 -827 0 3
rlabel polysilicon 1150 -821 1150 -821 0 1
rlabel polysilicon 1150 -827 1150 -827 0 3
rlabel polysilicon 1157 -821 1157 -821 0 1
rlabel polysilicon 1157 -827 1157 -827 0 3
rlabel polysilicon 1164 -821 1164 -821 0 1
rlabel polysilicon 1164 -827 1164 -827 0 3
rlabel polysilicon 1171 -821 1171 -821 0 1
rlabel polysilicon 1171 -827 1171 -827 0 3
rlabel polysilicon 1178 -821 1178 -821 0 1
rlabel polysilicon 1178 -827 1178 -827 0 3
rlabel polysilicon 1185 -821 1185 -821 0 1
rlabel polysilicon 1185 -827 1185 -827 0 3
rlabel polysilicon 1192 -821 1192 -821 0 1
rlabel polysilicon 1192 -827 1192 -827 0 3
rlabel polysilicon 1199 -821 1199 -821 0 1
rlabel polysilicon 1199 -827 1199 -827 0 3
rlabel polysilicon 1206 -821 1206 -821 0 1
rlabel polysilicon 1206 -827 1206 -827 0 3
rlabel polysilicon 1213 -821 1213 -821 0 1
rlabel polysilicon 1213 -827 1213 -827 0 3
rlabel polysilicon 1220 -821 1220 -821 0 1
rlabel polysilicon 1220 -827 1220 -827 0 3
rlabel polysilicon 5 -908 5 -908 0 2
rlabel polysilicon 9 -908 9 -908 0 1
rlabel polysilicon 9 -914 9 -914 0 3
rlabel polysilicon 19 -908 19 -908 0 2
rlabel polysilicon 19 -914 19 -914 0 4
rlabel polysilicon 23 -908 23 -908 0 1
rlabel polysilicon 23 -914 23 -914 0 3
rlabel polysilicon 33 -908 33 -908 0 2
rlabel polysilicon 33 -914 33 -914 0 4
rlabel polysilicon 37 -908 37 -908 0 1
rlabel polysilicon 40 -908 40 -908 0 2
rlabel polysilicon 37 -914 37 -914 0 3
rlabel polysilicon 40 -914 40 -914 0 4
rlabel polysilicon 44 -908 44 -908 0 1
rlabel polysilicon 44 -914 44 -914 0 3
rlabel polysilicon 51 -908 51 -908 0 1
rlabel polysilicon 51 -914 51 -914 0 3
rlabel polysilicon 58 -908 58 -908 0 1
rlabel polysilicon 58 -914 58 -914 0 3
rlabel polysilicon 65 -908 65 -908 0 1
rlabel polysilicon 65 -914 65 -914 0 3
rlabel polysilicon 72 -908 72 -908 0 1
rlabel polysilicon 72 -914 72 -914 0 3
rlabel polysilicon 79 -908 79 -908 0 1
rlabel polysilicon 79 -914 79 -914 0 3
rlabel polysilicon 86 -908 86 -908 0 1
rlabel polysilicon 86 -914 86 -914 0 3
rlabel polysilicon 93 -908 93 -908 0 1
rlabel polysilicon 93 -914 93 -914 0 3
rlabel polysilicon 100 -914 100 -914 0 3
rlabel polysilicon 107 -908 107 -908 0 1
rlabel polysilicon 107 -914 107 -914 0 3
rlabel polysilicon 117 -908 117 -908 0 2
rlabel polysilicon 114 -914 114 -914 0 3
rlabel polysilicon 117 -914 117 -914 0 4
rlabel polysilicon 121 -908 121 -908 0 1
rlabel polysilicon 121 -914 121 -914 0 3
rlabel polysilicon 128 -908 128 -908 0 1
rlabel polysilicon 128 -914 128 -914 0 3
rlabel polysilicon 135 -908 135 -908 0 1
rlabel polysilicon 135 -914 135 -914 0 3
rlabel polysilicon 142 -908 142 -908 0 1
rlabel polysilicon 142 -914 142 -914 0 3
rlabel polysilicon 149 -908 149 -908 0 1
rlabel polysilicon 152 -914 152 -914 0 4
rlabel polysilicon 156 -908 156 -908 0 1
rlabel polysilicon 156 -914 156 -914 0 3
rlabel polysilicon 163 -908 163 -908 0 1
rlabel polysilicon 163 -914 163 -914 0 3
rlabel polysilicon 170 -908 170 -908 0 1
rlabel polysilicon 170 -914 170 -914 0 3
rlabel polysilicon 177 -908 177 -908 0 1
rlabel polysilicon 177 -914 177 -914 0 3
rlabel polysilicon 184 -908 184 -908 0 1
rlabel polysilicon 184 -914 184 -914 0 3
rlabel polysilicon 191 -908 191 -908 0 1
rlabel polysilicon 191 -914 191 -914 0 3
rlabel polysilicon 198 -908 198 -908 0 1
rlabel polysilicon 198 -914 198 -914 0 3
rlabel polysilicon 205 -908 205 -908 0 1
rlabel polysilicon 208 -914 208 -914 0 4
rlabel polysilicon 212 -908 212 -908 0 1
rlabel polysilicon 212 -914 212 -914 0 3
rlabel polysilicon 219 -908 219 -908 0 1
rlabel polysilicon 219 -914 219 -914 0 3
rlabel polysilicon 226 -908 226 -908 0 1
rlabel polysilicon 226 -914 226 -914 0 3
rlabel polysilicon 233 -908 233 -908 0 1
rlabel polysilicon 233 -914 233 -914 0 3
rlabel polysilicon 240 -908 240 -908 0 1
rlabel polysilicon 240 -914 240 -914 0 3
rlabel polysilicon 247 -908 247 -908 0 1
rlabel polysilicon 247 -914 247 -914 0 3
rlabel polysilicon 254 -908 254 -908 0 1
rlabel polysilicon 254 -914 254 -914 0 3
rlabel polysilicon 264 -908 264 -908 0 2
rlabel polysilicon 261 -914 261 -914 0 3
rlabel polysilicon 264 -914 264 -914 0 4
rlabel polysilicon 268 -908 268 -908 0 1
rlabel polysilicon 268 -914 268 -914 0 3
rlabel polysilicon 278 -908 278 -908 0 2
rlabel polysilicon 275 -914 275 -914 0 3
rlabel polysilicon 282 -908 282 -908 0 1
rlabel polysilicon 282 -914 282 -914 0 3
rlabel polysilicon 289 -908 289 -908 0 1
rlabel polysilicon 292 -908 292 -908 0 2
rlabel polysilicon 289 -914 289 -914 0 3
rlabel polysilicon 296 -908 296 -908 0 1
rlabel polysilicon 296 -914 296 -914 0 3
rlabel polysilicon 303 -908 303 -908 0 1
rlabel polysilicon 303 -914 303 -914 0 3
rlabel polysilicon 310 -908 310 -908 0 1
rlabel polysilicon 313 -908 313 -908 0 2
rlabel polysilicon 317 -908 317 -908 0 1
rlabel polysilicon 317 -914 317 -914 0 3
rlabel polysilicon 324 -908 324 -908 0 1
rlabel polysilicon 324 -914 324 -914 0 3
rlabel polysilicon 331 -908 331 -908 0 1
rlabel polysilicon 331 -914 331 -914 0 3
rlabel polysilicon 338 -908 338 -908 0 1
rlabel polysilicon 338 -914 338 -914 0 3
rlabel polysilicon 348 -908 348 -908 0 2
rlabel polysilicon 348 -914 348 -914 0 4
rlabel polysilicon 352 -908 352 -908 0 1
rlabel polysilicon 352 -914 352 -914 0 3
rlabel polysilicon 359 -908 359 -908 0 1
rlabel polysilicon 359 -914 359 -914 0 3
rlabel polysilicon 366 -908 366 -908 0 1
rlabel polysilicon 366 -914 366 -914 0 3
rlabel polysilicon 373 -914 373 -914 0 3
rlabel polysilicon 380 -908 380 -908 0 1
rlabel polysilicon 380 -914 380 -914 0 3
rlabel polysilicon 387 -908 387 -908 0 1
rlabel polysilicon 387 -914 387 -914 0 3
rlabel polysilicon 394 -908 394 -908 0 1
rlabel polysilicon 394 -914 394 -914 0 3
rlabel polysilicon 401 -908 401 -908 0 1
rlabel polysilicon 401 -914 401 -914 0 3
rlabel polysilicon 408 -908 408 -908 0 1
rlabel polysilicon 408 -914 408 -914 0 3
rlabel polysilicon 415 -908 415 -908 0 1
rlabel polysilicon 415 -914 415 -914 0 3
rlabel polysilicon 425 -908 425 -908 0 2
rlabel polysilicon 422 -914 422 -914 0 3
rlabel polysilicon 429 -908 429 -908 0 1
rlabel polysilicon 429 -914 429 -914 0 3
rlabel polysilicon 436 -908 436 -908 0 1
rlabel polysilicon 436 -914 436 -914 0 3
rlabel polysilicon 439 -914 439 -914 0 4
rlabel polysilicon 443 -908 443 -908 0 1
rlabel polysilicon 443 -914 443 -914 0 3
rlabel polysilicon 450 -908 450 -908 0 1
rlabel polysilicon 450 -914 450 -914 0 3
rlabel polysilicon 457 -908 457 -908 0 1
rlabel polysilicon 457 -914 457 -914 0 3
rlabel polysilicon 464 -908 464 -908 0 1
rlabel polysilicon 464 -914 464 -914 0 3
rlabel polysilicon 471 -908 471 -908 0 1
rlabel polysilicon 471 -914 471 -914 0 3
rlabel polysilicon 478 -908 478 -908 0 1
rlabel polysilicon 485 -908 485 -908 0 1
rlabel polysilicon 485 -914 485 -914 0 3
rlabel polysilicon 492 -908 492 -908 0 1
rlabel polysilicon 492 -914 492 -914 0 3
rlabel polysilicon 499 -908 499 -908 0 1
rlabel polysilicon 499 -914 499 -914 0 3
rlabel polysilicon 506 -908 506 -908 0 1
rlabel polysilicon 506 -914 506 -914 0 3
rlabel polysilicon 513 -908 513 -908 0 1
rlabel polysilicon 513 -914 513 -914 0 3
rlabel polysilicon 520 -908 520 -908 0 1
rlabel polysilicon 520 -914 520 -914 0 3
rlabel polysilicon 527 -908 527 -908 0 1
rlabel polysilicon 527 -914 527 -914 0 3
rlabel polysilicon 534 -908 534 -908 0 1
rlabel polysilicon 534 -914 534 -914 0 3
rlabel polysilicon 541 -908 541 -908 0 1
rlabel polysilicon 544 -908 544 -908 0 2
rlabel polysilicon 548 -908 548 -908 0 1
rlabel polysilicon 548 -914 548 -914 0 3
rlabel polysilicon 555 -908 555 -908 0 1
rlabel polysilicon 555 -914 555 -914 0 3
rlabel polysilicon 558 -914 558 -914 0 4
rlabel polysilicon 562 -908 562 -908 0 1
rlabel polysilicon 562 -914 562 -914 0 3
rlabel polysilicon 569 -908 569 -908 0 1
rlabel polysilicon 569 -914 569 -914 0 3
rlabel polysilicon 576 -908 576 -908 0 1
rlabel polysilicon 576 -914 576 -914 0 3
rlabel polysilicon 583 -908 583 -908 0 1
rlabel polysilicon 583 -914 583 -914 0 3
rlabel polysilicon 590 -908 590 -908 0 1
rlabel polysilicon 590 -914 590 -914 0 3
rlabel polysilicon 597 -908 597 -908 0 1
rlabel polysilicon 600 -908 600 -908 0 2
rlabel polysilicon 597 -914 597 -914 0 3
rlabel polysilicon 604 -908 604 -908 0 1
rlabel polysilicon 604 -914 604 -914 0 3
rlabel polysilicon 611 -908 611 -908 0 1
rlabel polysilicon 614 -908 614 -908 0 2
rlabel polysilicon 614 -914 614 -914 0 4
rlabel polysilicon 621 -908 621 -908 0 2
rlabel polysilicon 625 -908 625 -908 0 1
rlabel polysilicon 625 -914 625 -914 0 3
rlabel polysilicon 632 -908 632 -908 0 1
rlabel polysilicon 632 -914 632 -914 0 3
rlabel polysilicon 639 -908 639 -908 0 1
rlabel polysilicon 639 -914 639 -914 0 3
rlabel polysilicon 646 -908 646 -908 0 1
rlabel polysilicon 646 -914 646 -914 0 3
rlabel polysilicon 653 -908 653 -908 0 1
rlabel polysilicon 656 -908 656 -908 0 2
rlabel polysilicon 653 -914 653 -914 0 3
rlabel polysilicon 656 -914 656 -914 0 4
rlabel polysilicon 660 -908 660 -908 0 1
rlabel polysilicon 660 -914 660 -914 0 3
rlabel polysilicon 667 -908 667 -908 0 1
rlabel polysilicon 670 -908 670 -908 0 2
rlabel polysilicon 674 -908 674 -908 0 1
rlabel polysilicon 677 -908 677 -908 0 2
rlabel polysilicon 681 -908 681 -908 0 1
rlabel polysilicon 684 -914 684 -914 0 4
rlabel polysilicon 688 -908 688 -908 0 1
rlabel polysilicon 688 -914 688 -914 0 3
rlabel polysilicon 695 -908 695 -908 0 1
rlabel polysilicon 695 -914 695 -914 0 3
rlabel polysilicon 702 -908 702 -908 0 1
rlabel polysilicon 702 -914 702 -914 0 3
rlabel polysilicon 709 -908 709 -908 0 1
rlabel polysilicon 709 -914 709 -914 0 3
rlabel polysilicon 716 -908 716 -908 0 1
rlabel polysilicon 716 -914 716 -914 0 3
rlabel polysilicon 723 -908 723 -908 0 1
rlabel polysilicon 723 -914 723 -914 0 3
rlabel polysilicon 730 -908 730 -908 0 1
rlabel polysilicon 730 -914 730 -914 0 3
rlabel polysilicon 737 -908 737 -908 0 1
rlabel polysilicon 737 -914 737 -914 0 3
rlabel polysilicon 744 -908 744 -908 0 1
rlabel polysilicon 744 -914 744 -914 0 3
rlabel polysilicon 751 -908 751 -908 0 1
rlabel polysilicon 751 -914 751 -914 0 3
rlabel polysilicon 758 -908 758 -908 0 1
rlabel polysilicon 758 -914 758 -914 0 3
rlabel polysilicon 765 -908 765 -908 0 1
rlabel polysilicon 765 -914 765 -914 0 3
rlabel polysilicon 772 -908 772 -908 0 1
rlabel polysilicon 772 -914 772 -914 0 3
rlabel polysilicon 779 -908 779 -908 0 1
rlabel polysilicon 779 -914 779 -914 0 3
rlabel polysilicon 786 -908 786 -908 0 1
rlabel polysilicon 786 -914 786 -914 0 3
rlabel polysilicon 793 -908 793 -908 0 1
rlabel polysilicon 793 -914 793 -914 0 3
rlabel polysilicon 800 -908 800 -908 0 1
rlabel polysilicon 800 -914 800 -914 0 3
rlabel polysilicon 807 -908 807 -908 0 1
rlabel polysilicon 807 -914 807 -914 0 3
rlabel polysilicon 814 -908 814 -908 0 1
rlabel polysilicon 814 -914 814 -914 0 3
rlabel polysilicon 821 -914 821 -914 0 3
rlabel polysilicon 824 -914 824 -914 0 4
rlabel polysilicon 828 -908 828 -908 0 1
rlabel polysilicon 828 -914 828 -914 0 3
rlabel polysilicon 835 -908 835 -908 0 1
rlabel polysilicon 835 -914 835 -914 0 3
rlabel polysilicon 842 -908 842 -908 0 1
rlabel polysilicon 842 -914 842 -914 0 3
rlabel polysilicon 849 -908 849 -908 0 1
rlabel polysilicon 849 -914 849 -914 0 3
rlabel polysilicon 856 -908 856 -908 0 1
rlabel polysilicon 856 -914 856 -914 0 3
rlabel polysilicon 863 -908 863 -908 0 1
rlabel polysilicon 863 -914 863 -914 0 3
rlabel polysilicon 870 -908 870 -908 0 1
rlabel polysilicon 870 -914 870 -914 0 3
rlabel polysilicon 877 -908 877 -908 0 1
rlabel polysilicon 877 -914 877 -914 0 3
rlabel polysilicon 884 -908 884 -908 0 1
rlabel polysilicon 884 -914 884 -914 0 3
rlabel polysilicon 891 -908 891 -908 0 1
rlabel polysilicon 891 -914 891 -914 0 3
rlabel polysilicon 898 -914 898 -914 0 3
rlabel polysilicon 901 -914 901 -914 0 4
rlabel polysilicon 905 -908 905 -908 0 1
rlabel polysilicon 905 -914 905 -914 0 3
rlabel polysilicon 912 -908 912 -908 0 1
rlabel polysilicon 912 -914 912 -914 0 3
rlabel polysilicon 919 -908 919 -908 0 1
rlabel polysilicon 919 -914 919 -914 0 3
rlabel polysilicon 926 -908 926 -908 0 1
rlabel polysilicon 926 -914 926 -914 0 3
rlabel polysilicon 933 -908 933 -908 0 1
rlabel polysilicon 933 -914 933 -914 0 3
rlabel polysilicon 940 -908 940 -908 0 1
rlabel polysilicon 940 -914 940 -914 0 3
rlabel polysilicon 947 -908 947 -908 0 1
rlabel polysilicon 947 -914 947 -914 0 3
rlabel polysilicon 954 -908 954 -908 0 1
rlabel polysilicon 954 -914 954 -914 0 3
rlabel polysilicon 961 -908 961 -908 0 1
rlabel polysilicon 961 -914 961 -914 0 3
rlabel polysilicon 968 -908 968 -908 0 1
rlabel polysilicon 968 -914 968 -914 0 3
rlabel polysilicon 975 -908 975 -908 0 1
rlabel polysilicon 975 -914 975 -914 0 3
rlabel polysilicon 982 -908 982 -908 0 1
rlabel polysilicon 982 -914 982 -914 0 3
rlabel polysilicon 989 -908 989 -908 0 1
rlabel polysilicon 989 -914 989 -914 0 3
rlabel polysilicon 996 -908 996 -908 0 1
rlabel polysilicon 999 -908 999 -908 0 2
rlabel polysilicon 996 -914 996 -914 0 3
rlabel polysilicon 1003 -908 1003 -908 0 1
rlabel polysilicon 1003 -914 1003 -914 0 3
rlabel polysilicon 1010 -908 1010 -908 0 1
rlabel polysilicon 1010 -914 1010 -914 0 3
rlabel polysilicon 1017 -908 1017 -908 0 1
rlabel polysilicon 1017 -914 1017 -914 0 3
rlabel polysilicon 1024 -908 1024 -908 0 1
rlabel polysilicon 1024 -914 1024 -914 0 3
rlabel polysilicon 1031 -908 1031 -908 0 1
rlabel polysilicon 1031 -914 1031 -914 0 3
rlabel polysilicon 1038 -908 1038 -908 0 1
rlabel polysilicon 1038 -914 1038 -914 0 3
rlabel polysilicon 1045 -908 1045 -908 0 1
rlabel polysilicon 1045 -914 1045 -914 0 3
rlabel polysilicon 1052 -908 1052 -908 0 1
rlabel polysilicon 1052 -914 1052 -914 0 3
rlabel polysilicon 1059 -908 1059 -908 0 1
rlabel polysilicon 1059 -914 1059 -914 0 3
rlabel polysilicon 1066 -908 1066 -908 0 1
rlabel polysilicon 1066 -914 1066 -914 0 3
rlabel polysilicon 1073 -908 1073 -908 0 1
rlabel polysilicon 1073 -914 1073 -914 0 3
rlabel polysilicon 1080 -908 1080 -908 0 1
rlabel polysilicon 1080 -914 1080 -914 0 3
rlabel polysilicon 1087 -908 1087 -908 0 1
rlabel polysilicon 1090 -908 1090 -908 0 2
rlabel polysilicon 1090 -914 1090 -914 0 4
rlabel polysilicon 1094 -908 1094 -908 0 1
rlabel polysilicon 1094 -914 1094 -914 0 3
rlabel polysilicon 1101 -908 1101 -908 0 1
rlabel polysilicon 1101 -914 1101 -914 0 3
rlabel polysilicon 1108 -908 1108 -908 0 1
rlabel polysilicon 1108 -914 1108 -914 0 3
rlabel polysilicon 1115 -908 1115 -908 0 1
rlabel polysilicon 1115 -914 1115 -914 0 3
rlabel polysilicon 1122 -908 1122 -908 0 1
rlabel polysilicon 1122 -914 1122 -914 0 3
rlabel polysilicon 1129 -908 1129 -908 0 1
rlabel polysilicon 1129 -914 1129 -914 0 3
rlabel polysilicon 1164 -908 1164 -908 0 1
rlabel polysilicon 1164 -914 1164 -914 0 3
rlabel polysilicon 1171 -908 1171 -908 0 1
rlabel polysilicon 1171 -914 1171 -914 0 3
rlabel polysilicon 1178 -908 1178 -908 0 1
rlabel polysilicon 1178 -914 1178 -914 0 3
rlabel polysilicon 1192 -908 1192 -908 0 1
rlabel polysilicon 1192 -914 1192 -914 0 3
rlabel polysilicon 2 -997 2 -997 0 1
rlabel polysilicon 2 -1003 2 -1003 0 3
rlabel polysilicon 9 -997 9 -997 0 1
rlabel polysilicon 9 -1003 9 -1003 0 3
rlabel polysilicon 16 -1003 16 -1003 0 3
rlabel polysilicon 23 -997 23 -997 0 1
rlabel polysilicon 23 -1003 23 -1003 0 3
rlabel polysilicon 30 -997 30 -997 0 1
rlabel polysilicon 30 -1003 30 -1003 0 3
rlabel polysilicon 40 -997 40 -997 0 2
rlabel polysilicon 40 -1003 40 -1003 0 4
rlabel polysilicon 44 -997 44 -997 0 1
rlabel polysilicon 44 -1003 44 -1003 0 3
rlabel polysilicon 51 -997 51 -997 0 1
rlabel polysilicon 51 -1003 51 -1003 0 3
rlabel polysilicon 58 -997 58 -997 0 1
rlabel polysilicon 61 -997 61 -997 0 2
rlabel polysilicon 61 -1003 61 -1003 0 4
rlabel polysilicon 65 -997 65 -997 0 1
rlabel polysilicon 65 -1003 65 -1003 0 3
rlabel polysilicon 72 -997 72 -997 0 1
rlabel polysilicon 72 -1003 72 -1003 0 3
rlabel polysilicon 79 -997 79 -997 0 1
rlabel polysilicon 79 -1003 79 -1003 0 3
rlabel polysilicon 86 -997 86 -997 0 1
rlabel polysilicon 86 -1003 86 -1003 0 3
rlabel polysilicon 93 -997 93 -997 0 1
rlabel polysilicon 96 -997 96 -997 0 2
rlabel polysilicon 96 -1003 96 -1003 0 4
rlabel polysilicon 100 -997 100 -997 0 1
rlabel polysilicon 103 -1003 103 -1003 0 4
rlabel polysilicon 107 -997 107 -997 0 1
rlabel polysilicon 107 -1003 107 -1003 0 3
rlabel polysilicon 114 -997 114 -997 0 1
rlabel polysilicon 114 -1003 114 -1003 0 3
rlabel polysilicon 121 -997 121 -997 0 1
rlabel polysilicon 124 -1003 124 -1003 0 4
rlabel polysilicon 128 -997 128 -997 0 1
rlabel polysilicon 128 -1003 128 -1003 0 3
rlabel polysilicon 135 -997 135 -997 0 1
rlabel polysilicon 135 -1003 135 -1003 0 3
rlabel polysilicon 142 -997 142 -997 0 1
rlabel polysilicon 142 -1003 142 -1003 0 3
rlabel polysilicon 149 -997 149 -997 0 1
rlabel polysilicon 149 -1003 149 -1003 0 3
rlabel polysilicon 156 -997 156 -997 0 1
rlabel polysilicon 156 -1003 156 -1003 0 3
rlabel polysilicon 163 -997 163 -997 0 1
rlabel polysilicon 163 -1003 163 -1003 0 3
rlabel polysilicon 170 -997 170 -997 0 1
rlabel polysilicon 170 -1003 170 -1003 0 3
rlabel polysilicon 177 -997 177 -997 0 1
rlabel polysilicon 177 -1003 177 -1003 0 3
rlabel polysilicon 184 -997 184 -997 0 1
rlabel polysilicon 187 -1003 187 -1003 0 4
rlabel polysilicon 191 -997 191 -997 0 1
rlabel polysilicon 191 -1003 191 -1003 0 3
rlabel polysilicon 198 -997 198 -997 0 1
rlabel polysilicon 198 -1003 198 -1003 0 3
rlabel polysilicon 201 -1003 201 -1003 0 4
rlabel polysilicon 205 -997 205 -997 0 1
rlabel polysilicon 205 -1003 205 -1003 0 3
rlabel polysilicon 212 -997 212 -997 0 1
rlabel polysilicon 212 -1003 212 -1003 0 3
rlabel polysilicon 219 -997 219 -997 0 1
rlabel polysilicon 219 -1003 219 -1003 0 3
rlabel polysilicon 226 -997 226 -997 0 1
rlabel polysilicon 226 -1003 226 -1003 0 3
rlabel polysilicon 233 -997 233 -997 0 1
rlabel polysilicon 233 -1003 233 -1003 0 3
rlabel polysilicon 240 -997 240 -997 0 1
rlabel polysilicon 240 -1003 240 -1003 0 3
rlabel polysilicon 247 -997 247 -997 0 1
rlabel polysilicon 247 -1003 247 -1003 0 3
rlabel polysilicon 254 -997 254 -997 0 1
rlabel polysilicon 254 -1003 254 -1003 0 3
rlabel polysilicon 261 -997 261 -997 0 1
rlabel polysilicon 261 -1003 261 -1003 0 3
rlabel polysilicon 268 -997 268 -997 0 1
rlabel polysilicon 268 -1003 268 -1003 0 3
rlabel polysilicon 275 -997 275 -997 0 1
rlabel polysilicon 275 -1003 275 -1003 0 3
rlabel polysilicon 282 -997 282 -997 0 1
rlabel polysilicon 282 -1003 282 -1003 0 3
rlabel polysilicon 289 -997 289 -997 0 1
rlabel polysilicon 289 -1003 289 -1003 0 3
rlabel polysilicon 296 -997 296 -997 0 1
rlabel polysilicon 296 -1003 296 -1003 0 3
rlabel polysilicon 303 -997 303 -997 0 1
rlabel polysilicon 303 -1003 303 -1003 0 3
rlabel polysilicon 310 -997 310 -997 0 1
rlabel polysilicon 310 -1003 310 -1003 0 3
rlabel polysilicon 317 -997 317 -997 0 1
rlabel polysilicon 317 -1003 317 -1003 0 3
rlabel polysilicon 324 -997 324 -997 0 1
rlabel polysilicon 324 -1003 324 -1003 0 3
rlabel polysilicon 331 -997 331 -997 0 1
rlabel polysilicon 331 -1003 331 -1003 0 3
rlabel polysilicon 338 -997 338 -997 0 1
rlabel polysilicon 338 -1003 338 -1003 0 3
rlabel polysilicon 345 -997 345 -997 0 1
rlabel polysilicon 345 -1003 345 -1003 0 3
rlabel polysilicon 352 -997 352 -997 0 1
rlabel polysilicon 352 -1003 352 -1003 0 3
rlabel polysilicon 362 -997 362 -997 0 2
rlabel polysilicon 359 -1003 359 -1003 0 3
rlabel polysilicon 362 -1003 362 -1003 0 4
rlabel polysilicon 366 -997 366 -997 0 1
rlabel polysilicon 366 -1003 366 -1003 0 3
rlabel polysilicon 376 -997 376 -997 0 2
rlabel polysilicon 373 -1003 373 -1003 0 3
rlabel polysilicon 376 -1003 376 -1003 0 4
rlabel polysilicon 380 -997 380 -997 0 1
rlabel polysilicon 380 -1003 380 -1003 0 3
rlabel polysilicon 390 -997 390 -997 0 2
rlabel polysilicon 390 -1003 390 -1003 0 4
rlabel polysilicon 394 -997 394 -997 0 1
rlabel polysilicon 394 -1003 394 -1003 0 3
rlabel polysilicon 401 -997 401 -997 0 1
rlabel polysilicon 401 -1003 401 -1003 0 3
rlabel polysilicon 408 -997 408 -997 0 1
rlabel polysilicon 408 -1003 408 -1003 0 3
rlabel polysilicon 415 -997 415 -997 0 1
rlabel polysilicon 415 -1003 415 -1003 0 3
rlabel polysilicon 422 -997 422 -997 0 1
rlabel polysilicon 422 -1003 422 -1003 0 3
rlabel polysilicon 429 -997 429 -997 0 1
rlabel polysilicon 429 -1003 429 -1003 0 3
rlabel polysilicon 439 -997 439 -997 0 2
rlabel polysilicon 436 -1003 436 -1003 0 3
rlabel polysilicon 443 -997 443 -997 0 1
rlabel polysilicon 443 -1003 443 -1003 0 3
rlabel polysilicon 450 -997 450 -997 0 1
rlabel polysilicon 450 -1003 450 -1003 0 3
rlabel polysilicon 457 -997 457 -997 0 1
rlabel polysilicon 457 -1003 457 -1003 0 3
rlabel polysilicon 464 -1003 464 -1003 0 3
rlabel polysilicon 471 -997 471 -997 0 1
rlabel polysilicon 471 -1003 471 -1003 0 3
rlabel polysilicon 478 -997 478 -997 0 1
rlabel polysilicon 478 -1003 478 -1003 0 3
rlabel polysilicon 485 -997 485 -997 0 1
rlabel polysilicon 485 -1003 485 -1003 0 3
rlabel polysilicon 492 -997 492 -997 0 1
rlabel polysilicon 492 -1003 492 -1003 0 3
rlabel polysilicon 499 -997 499 -997 0 1
rlabel polysilicon 502 -997 502 -997 0 2
rlabel polysilicon 499 -1003 499 -1003 0 3
rlabel polysilicon 502 -1003 502 -1003 0 4
rlabel polysilicon 506 -1003 506 -1003 0 3
rlabel polysilicon 509 -1003 509 -1003 0 4
rlabel polysilicon 513 -997 513 -997 0 1
rlabel polysilicon 513 -1003 513 -1003 0 3
rlabel polysilicon 520 -997 520 -997 0 1
rlabel polysilicon 520 -1003 520 -1003 0 3
rlabel polysilicon 527 -997 527 -997 0 1
rlabel polysilicon 527 -1003 527 -1003 0 3
rlabel polysilicon 534 -997 534 -997 0 1
rlabel polysilicon 534 -1003 534 -1003 0 3
rlabel polysilicon 544 -997 544 -997 0 2
rlabel polysilicon 541 -1003 541 -1003 0 3
rlabel polysilicon 544 -1003 544 -1003 0 4
rlabel polysilicon 548 -997 548 -997 0 1
rlabel polysilicon 548 -1003 548 -1003 0 3
rlabel polysilicon 555 -997 555 -997 0 1
rlabel polysilicon 555 -1003 555 -1003 0 3
rlabel polysilicon 562 -997 562 -997 0 1
rlabel polysilicon 562 -1003 562 -1003 0 3
rlabel polysilicon 569 -997 569 -997 0 1
rlabel polysilicon 569 -1003 569 -1003 0 3
rlabel polysilicon 576 -997 576 -997 0 1
rlabel polysilicon 576 -1003 576 -1003 0 3
rlabel polysilicon 583 -997 583 -997 0 1
rlabel polysilicon 583 -1003 583 -1003 0 3
rlabel polysilicon 590 -997 590 -997 0 1
rlabel polysilicon 590 -1003 590 -1003 0 3
rlabel polysilicon 597 -997 597 -997 0 1
rlabel polysilicon 597 -1003 597 -1003 0 3
rlabel polysilicon 604 -997 604 -997 0 1
rlabel polysilicon 607 -997 607 -997 0 2
rlabel polysilicon 607 -1003 607 -1003 0 4
rlabel polysilicon 611 -997 611 -997 0 1
rlabel polysilicon 611 -1003 611 -1003 0 3
rlabel polysilicon 618 -997 618 -997 0 1
rlabel polysilicon 618 -1003 618 -1003 0 3
rlabel polysilicon 628 -997 628 -997 0 2
rlabel polysilicon 632 -997 632 -997 0 1
rlabel polysilicon 632 -1003 632 -1003 0 3
rlabel polysilicon 639 -1003 639 -1003 0 3
rlabel polysilicon 642 -1003 642 -1003 0 4
rlabel polysilicon 649 -1003 649 -1003 0 4
rlabel polysilicon 653 -997 653 -997 0 1
rlabel polysilicon 653 -1003 653 -1003 0 3
rlabel polysilicon 660 -997 660 -997 0 1
rlabel polysilicon 660 -1003 660 -1003 0 3
rlabel polysilicon 667 -997 667 -997 0 1
rlabel polysilicon 667 -1003 667 -1003 0 3
rlabel polysilicon 674 -997 674 -997 0 1
rlabel polysilicon 674 -1003 674 -1003 0 3
rlabel polysilicon 681 -997 681 -997 0 1
rlabel polysilicon 681 -1003 681 -1003 0 3
rlabel polysilicon 684 -1003 684 -1003 0 4
rlabel polysilicon 688 -997 688 -997 0 1
rlabel polysilicon 688 -1003 688 -1003 0 3
rlabel polysilicon 695 -997 695 -997 0 1
rlabel polysilicon 698 -1003 698 -1003 0 4
rlabel polysilicon 702 -997 702 -997 0 1
rlabel polysilicon 702 -1003 702 -1003 0 3
rlabel polysilicon 709 -997 709 -997 0 1
rlabel polysilicon 712 -997 712 -997 0 2
rlabel polysilicon 709 -1003 709 -1003 0 3
rlabel polysilicon 716 -997 716 -997 0 1
rlabel polysilicon 716 -1003 716 -1003 0 3
rlabel polysilicon 723 -997 723 -997 0 1
rlabel polysilicon 723 -1003 723 -1003 0 3
rlabel polysilicon 730 -997 730 -997 0 1
rlabel polysilicon 733 -997 733 -997 0 2
rlabel polysilicon 730 -1003 730 -1003 0 3
rlabel polysilicon 737 -997 737 -997 0 1
rlabel polysilicon 737 -1003 737 -1003 0 3
rlabel polysilicon 744 -997 744 -997 0 1
rlabel polysilicon 744 -1003 744 -1003 0 3
rlabel polysilicon 751 -997 751 -997 0 1
rlabel polysilicon 751 -1003 751 -1003 0 3
rlabel polysilicon 758 -997 758 -997 0 1
rlabel polysilicon 758 -1003 758 -1003 0 3
rlabel polysilicon 765 -997 765 -997 0 1
rlabel polysilicon 765 -1003 765 -1003 0 3
rlabel polysilicon 772 -997 772 -997 0 1
rlabel polysilicon 772 -1003 772 -1003 0 3
rlabel polysilicon 779 -997 779 -997 0 1
rlabel polysilicon 779 -1003 779 -1003 0 3
rlabel polysilicon 786 -997 786 -997 0 1
rlabel polysilicon 786 -1003 786 -1003 0 3
rlabel polysilicon 793 -997 793 -997 0 1
rlabel polysilicon 793 -1003 793 -1003 0 3
rlabel polysilicon 800 -997 800 -997 0 1
rlabel polysilicon 800 -1003 800 -1003 0 3
rlabel polysilicon 807 -997 807 -997 0 1
rlabel polysilicon 807 -1003 807 -1003 0 3
rlabel polysilicon 814 -997 814 -997 0 1
rlabel polysilicon 814 -1003 814 -1003 0 3
rlabel polysilicon 821 -997 821 -997 0 1
rlabel polysilicon 821 -1003 821 -1003 0 3
rlabel polysilicon 828 -997 828 -997 0 1
rlabel polysilicon 828 -1003 828 -1003 0 3
rlabel polysilicon 835 -997 835 -997 0 1
rlabel polysilicon 835 -1003 835 -1003 0 3
rlabel polysilicon 842 -997 842 -997 0 1
rlabel polysilicon 842 -1003 842 -1003 0 3
rlabel polysilicon 849 -997 849 -997 0 1
rlabel polysilicon 849 -1003 849 -1003 0 3
rlabel polysilicon 859 -997 859 -997 0 2
rlabel polysilicon 856 -1003 856 -1003 0 3
rlabel polysilicon 859 -1003 859 -1003 0 4
rlabel polysilicon 863 -997 863 -997 0 1
rlabel polysilicon 863 -1003 863 -1003 0 3
rlabel polysilicon 870 -997 870 -997 0 1
rlabel polysilicon 870 -1003 870 -1003 0 3
rlabel polysilicon 877 -997 877 -997 0 1
rlabel polysilicon 877 -1003 877 -1003 0 3
rlabel polysilicon 884 -997 884 -997 0 1
rlabel polysilicon 884 -1003 884 -1003 0 3
rlabel polysilicon 891 -997 891 -997 0 1
rlabel polysilicon 891 -1003 891 -1003 0 3
rlabel polysilicon 898 -997 898 -997 0 1
rlabel polysilicon 898 -1003 898 -1003 0 3
rlabel polysilicon 905 -997 905 -997 0 1
rlabel polysilicon 905 -1003 905 -1003 0 3
rlabel polysilicon 912 -997 912 -997 0 1
rlabel polysilicon 912 -1003 912 -1003 0 3
rlabel polysilicon 919 -997 919 -997 0 1
rlabel polysilicon 919 -1003 919 -1003 0 3
rlabel polysilicon 926 -997 926 -997 0 1
rlabel polysilicon 926 -1003 926 -1003 0 3
rlabel polysilicon 933 -997 933 -997 0 1
rlabel polysilicon 933 -1003 933 -1003 0 3
rlabel polysilicon 940 -997 940 -997 0 1
rlabel polysilicon 940 -1003 940 -1003 0 3
rlabel polysilicon 947 -997 947 -997 0 1
rlabel polysilicon 947 -1003 947 -1003 0 3
rlabel polysilicon 954 -997 954 -997 0 1
rlabel polysilicon 954 -1003 954 -1003 0 3
rlabel polysilicon 961 -997 961 -997 0 1
rlabel polysilicon 961 -1003 961 -1003 0 3
rlabel polysilicon 968 -997 968 -997 0 1
rlabel polysilicon 968 -1003 968 -1003 0 3
rlabel polysilicon 975 -997 975 -997 0 1
rlabel polysilicon 975 -1003 975 -1003 0 3
rlabel polysilicon 982 -997 982 -997 0 1
rlabel polysilicon 982 -1003 982 -1003 0 3
rlabel polysilicon 989 -997 989 -997 0 1
rlabel polysilicon 989 -1003 989 -1003 0 3
rlabel polysilicon 996 -997 996 -997 0 1
rlabel polysilicon 996 -1003 996 -1003 0 3
rlabel polysilicon 1003 -997 1003 -997 0 1
rlabel polysilicon 1003 -1003 1003 -1003 0 3
rlabel polysilicon 1010 -997 1010 -997 0 1
rlabel polysilicon 1010 -1003 1010 -1003 0 3
rlabel polysilicon 1017 -997 1017 -997 0 1
rlabel polysilicon 1017 -1003 1017 -1003 0 3
rlabel polysilicon 1024 -997 1024 -997 0 1
rlabel polysilicon 1024 -1003 1024 -1003 0 3
rlabel polysilicon 1031 -997 1031 -997 0 1
rlabel polysilicon 1031 -1003 1031 -1003 0 3
rlabel polysilicon 1038 -997 1038 -997 0 1
rlabel polysilicon 1038 -1003 1038 -1003 0 3
rlabel polysilicon 1045 -997 1045 -997 0 1
rlabel polysilicon 1045 -1003 1045 -1003 0 3
rlabel polysilicon 1052 -997 1052 -997 0 1
rlabel polysilicon 1052 -1003 1052 -1003 0 3
rlabel polysilicon 1059 -997 1059 -997 0 1
rlabel polysilicon 1059 -1003 1059 -1003 0 3
rlabel polysilicon 1066 -997 1066 -997 0 1
rlabel polysilicon 1066 -1003 1066 -1003 0 3
rlabel polysilicon 1073 -997 1073 -997 0 1
rlabel polysilicon 1073 -1003 1073 -1003 0 3
rlabel polysilicon 1080 -997 1080 -997 0 1
rlabel polysilicon 1080 -1003 1080 -1003 0 3
rlabel polysilicon 1087 -997 1087 -997 0 1
rlabel polysilicon 1087 -1003 1087 -1003 0 3
rlabel polysilicon 1094 -997 1094 -997 0 1
rlabel polysilicon 1094 -1003 1094 -1003 0 3
rlabel polysilicon 1101 -997 1101 -997 0 1
rlabel polysilicon 1101 -1003 1101 -1003 0 3
rlabel polysilicon 1108 -997 1108 -997 0 1
rlabel polysilicon 1108 -1003 1108 -1003 0 3
rlabel polysilicon 1115 -997 1115 -997 0 1
rlabel polysilicon 1115 -1003 1115 -1003 0 3
rlabel polysilicon 1122 -997 1122 -997 0 1
rlabel polysilicon 1122 -1003 1122 -1003 0 3
rlabel polysilicon 1129 -997 1129 -997 0 1
rlabel polysilicon 1129 -1003 1129 -1003 0 3
rlabel polysilicon 1132 -1003 1132 -1003 0 4
rlabel polysilicon 1136 -997 1136 -997 0 1
rlabel polysilicon 1136 -1003 1136 -1003 0 3
rlabel polysilicon 1143 -997 1143 -997 0 1
rlabel polysilicon 1143 -1003 1143 -1003 0 3
rlabel polysilicon 1150 -997 1150 -997 0 1
rlabel polysilicon 1150 -1003 1150 -1003 0 3
rlabel polysilicon 1157 -997 1157 -997 0 1
rlabel polysilicon 1157 -1003 1157 -1003 0 3
rlabel polysilicon 1164 -997 1164 -997 0 1
rlabel polysilicon 1167 -1003 1167 -1003 0 4
rlabel polysilicon 1171 -997 1171 -997 0 1
rlabel polysilicon 1171 -1003 1171 -1003 0 3
rlabel polysilicon 1185 -997 1185 -997 0 1
rlabel polysilicon 1185 -1003 1185 -1003 0 3
rlabel polysilicon 1192 -997 1192 -997 0 1
rlabel polysilicon 16 -1072 16 -1072 0 1
rlabel polysilicon 16 -1078 16 -1078 0 3
rlabel polysilicon 23 -1072 23 -1072 0 1
rlabel polysilicon 23 -1078 23 -1078 0 3
rlabel polysilicon 30 -1072 30 -1072 0 1
rlabel polysilicon 30 -1078 30 -1078 0 3
rlabel polysilicon 37 -1072 37 -1072 0 1
rlabel polysilicon 37 -1078 37 -1078 0 3
rlabel polysilicon 44 -1072 44 -1072 0 1
rlabel polysilicon 44 -1078 44 -1078 0 3
rlabel polysilicon 51 -1072 51 -1072 0 1
rlabel polysilicon 51 -1078 51 -1078 0 3
rlabel polysilicon 58 -1072 58 -1072 0 1
rlabel polysilicon 61 -1072 61 -1072 0 2
rlabel polysilicon 65 -1072 65 -1072 0 1
rlabel polysilicon 68 -1078 68 -1078 0 4
rlabel polysilicon 72 -1072 72 -1072 0 1
rlabel polysilicon 72 -1078 72 -1078 0 3
rlabel polysilicon 79 -1072 79 -1072 0 1
rlabel polysilicon 79 -1078 79 -1078 0 3
rlabel polysilicon 86 -1072 86 -1072 0 1
rlabel polysilicon 89 -1072 89 -1072 0 2
rlabel polysilicon 93 -1072 93 -1072 0 1
rlabel polysilicon 96 -1072 96 -1072 0 2
rlabel polysilicon 100 -1072 100 -1072 0 1
rlabel polysilicon 100 -1078 100 -1078 0 3
rlabel polysilicon 107 -1072 107 -1072 0 1
rlabel polysilicon 107 -1078 107 -1078 0 3
rlabel polysilicon 117 -1072 117 -1072 0 2
rlabel polysilicon 121 -1072 121 -1072 0 1
rlabel polysilicon 121 -1078 121 -1078 0 3
rlabel polysilicon 128 -1072 128 -1072 0 1
rlabel polysilicon 128 -1078 128 -1078 0 3
rlabel polysilicon 135 -1072 135 -1072 0 1
rlabel polysilicon 135 -1078 135 -1078 0 3
rlabel polysilicon 142 -1072 142 -1072 0 1
rlabel polysilicon 142 -1078 142 -1078 0 3
rlabel polysilicon 152 -1072 152 -1072 0 2
rlabel polysilicon 149 -1078 149 -1078 0 3
rlabel polysilicon 156 -1072 156 -1072 0 1
rlabel polysilicon 156 -1078 156 -1078 0 3
rlabel polysilicon 163 -1072 163 -1072 0 1
rlabel polysilicon 163 -1078 163 -1078 0 3
rlabel polysilicon 173 -1072 173 -1072 0 2
rlabel polysilicon 170 -1078 170 -1078 0 3
rlabel polysilicon 177 -1072 177 -1072 0 1
rlabel polysilicon 177 -1078 177 -1078 0 3
rlabel polysilicon 184 -1072 184 -1072 0 1
rlabel polysilicon 184 -1078 184 -1078 0 3
rlabel polysilicon 191 -1072 191 -1072 0 1
rlabel polysilicon 191 -1078 191 -1078 0 3
rlabel polysilicon 198 -1072 198 -1072 0 1
rlabel polysilicon 198 -1078 198 -1078 0 3
rlabel polysilicon 205 -1072 205 -1072 0 1
rlabel polysilicon 208 -1072 208 -1072 0 2
rlabel polysilicon 205 -1078 205 -1078 0 3
rlabel polysilicon 212 -1072 212 -1072 0 1
rlabel polysilicon 212 -1078 212 -1078 0 3
rlabel polysilicon 219 -1072 219 -1072 0 1
rlabel polysilicon 219 -1078 219 -1078 0 3
rlabel polysilicon 226 -1072 226 -1072 0 1
rlabel polysilicon 226 -1078 226 -1078 0 3
rlabel polysilicon 233 -1072 233 -1072 0 1
rlabel polysilicon 233 -1078 233 -1078 0 3
rlabel polysilicon 240 -1072 240 -1072 0 1
rlabel polysilicon 240 -1078 240 -1078 0 3
rlabel polysilicon 247 -1072 247 -1072 0 1
rlabel polysilicon 247 -1078 247 -1078 0 3
rlabel polysilicon 254 -1072 254 -1072 0 1
rlabel polysilicon 254 -1078 254 -1078 0 3
rlabel polysilicon 264 -1072 264 -1072 0 2
rlabel polysilicon 261 -1078 261 -1078 0 3
rlabel polysilicon 264 -1078 264 -1078 0 4
rlabel polysilicon 268 -1072 268 -1072 0 1
rlabel polysilicon 268 -1078 268 -1078 0 3
rlabel polysilicon 275 -1072 275 -1072 0 1
rlabel polysilicon 275 -1078 275 -1078 0 3
rlabel polysilicon 282 -1072 282 -1072 0 1
rlabel polysilicon 282 -1078 282 -1078 0 3
rlabel polysilicon 289 -1072 289 -1072 0 1
rlabel polysilicon 289 -1078 289 -1078 0 3
rlabel polysilicon 296 -1078 296 -1078 0 3
rlabel polysilicon 299 -1078 299 -1078 0 4
rlabel polysilicon 303 -1072 303 -1072 0 1
rlabel polysilicon 303 -1078 303 -1078 0 3
rlabel polysilicon 310 -1072 310 -1072 0 1
rlabel polysilicon 310 -1078 310 -1078 0 3
rlabel polysilicon 317 -1072 317 -1072 0 1
rlabel polysilicon 320 -1072 320 -1072 0 2
rlabel polysilicon 317 -1078 317 -1078 0 3
rlabel polysilicon 324 -1072 324 -1072 0 1
rlabel polysilicon 324 -1078 324 -1078 0 3
rlabel polysilicon 331 -1072 331 -1072 0 1
rlabel polysilicon 331 -1078 331 -1078 0 3
rlabel polysilicon 338 -1072 338 -1072 0 1
rlabel polysilicon 338 -1078 338 -1078 0 3
rlabel polysilicon 345 -1072 345 -1072 0 1
rlabel polysilicon 345 -1078 345 -1078 0 3
rlabel polysilicon 352 -1072 352 -1072 0 1
rlabel polysilicon 355 -1072 355 -1072 0 2
rlabel polysilicon 355 -1078 355 -1078 0 4
rlabel polysilicon 359 -1072 359 -1072 0 1
rlabel polysilicon 359 -1078 359 -1078 0 3
rlabel polysilicon 366 -1072 366 -1072 0 1
rlabel polysilicon 366 -1078 366 -1078 0 3
rlabel polysilicon 373 -1072 373 -1072 0 1
rlabel polysilicon 373 -1078 373 -1078 0 3
rlabel polysilicon 380 -1072 380 -1072 0 1
rlabel polysilicon 380 -1078 380 -1078 0 3
rlabel polysilicon 387 -1072 387 -1072 0 1
rlabel polysilicon 387 -1078 387 -1078 0 3
rlabel polysilicon 394 -1072 394 -1072 0 1
rlabel polysilicon 394 -1078 394 -1078 0 3
rlabel polysilicon 401 -1072 401 -1072 0 1
rlabel polysilicon 401 -1078 401 -1078 0 3
rlabel polysilicon 408 -1072 408 -1072 0 1
rlabel polysilicon 408 -1078 408 -1078 0 3
rlabel polysilicon 415 -1072 415 -1072 0 1
rlabel polysilicon 415 -1078 415 -1078 0 3
rlabel polysilicon 422 -1072 422 -1072 0 1
rlabel polysilicon 422 -1078 422 -1078 0 3
rlabel polysilicon 429 -1072 429 -1072 0 1
rlabel polysilicon 429 -1078 429 -1078 0 3
rlabel polysilicon 436 -1072 436 -1072 0 1
rlabel polysilicon 436 -1078 436 -1078 0 3
rlabel polysilicon 443 -1072 443 -1072 0 1
rlabel polysilicon 443 -1078 443 -1078 0 3
rlabel polysilicon 450 -1072 450 -1072 0 1
rlabel polysilicon 450 -1078 450 -1078 0 3
rlabel polysilicon 457 -1072 457 -1072 0 1
rlabel polysilicon 457 -1078 457 -1078 0 3
rlabel polysilicon 464 -1078 464 -1078 0 3
rlabel polysilicon 467 -1078 467 -1078 0 4
rlabel polysilicon 471 -1072 471 -1072 0 1
rlabel polysilicon 471 -1078 471 -1078 0 3
rlabel polysilicon 478 -1072 478 -1072 0 1
rlabel polysilicon 478 -1078 478 -1078 0 3
rlabel polysilicon 485 -1072 485 -1072 0 1
rlabel polysilicon 485 -1078 485 -1078 0 3
rlabel polysilicon 492 -1072 492 -1072 0 1
rlabel polysilicon 492 -1078 492 -1078 0 3
rlabel polysilicon 499 -1072 499 -1072 0 1
rlabel polysilicon 499 -1078 499 -1078 0 3
rlabel polysilicon 506 -1078 506 -1078 0 3
rlabel polysilicon 509 -1078 509 -1078 0 4
rlabel polysilicon 513 -1072 513 -1072 0 1
rlabel polysilicon 513 -1078 513 -1078 0 3
rlabel polysilicon 520 -1072 520 -1072 0 1
rlabel polysilicon 520 -1078 520 -1078 0 3
rlabel polysilicon 527 -1072 527 -1072 0 1
rlabel polysilicon 527 -1078 527 -1078 0 3
rlabel polysilicon 534 -1072 534 -1072 0 1
rlabel polysilicon 534 -1078 534 -1078 0 3
rlabel polysilicon 537 -1078 537 -1078 0 4
rlabel polysilicon 541 -1072 541 -1072 0 1
rlabel polysilicon 541 -1078 541 -1078 0 3
rlabel polysilicon 548 -1072 548 -1072 0 1
rlabel polysilicon 548 -1078 548 -1078 0 3
rlabel polysilicon 555 -1072 555 -1072 0 1
rlabel polysilicon 555 -1078 555 -1078 0 3
rlabel polysilicon 562 -1072 562 -1072 0 1
rlabel polysilicon 562 -1078 562 -1078 0 3
rlabel polysilicon 572 -1072 572 -1072 0 2
rlabel polysilicon 569 -1078 569 -1078 0 3
rlabel polysilicon 572 -1078 572 -1078 0 4
rlabel polysilicon 576 -1072 576 -1072 0 1
rlabel polysilicon 576 -1078 576 -1078 0 3
rlabel polysilicon 583 -1072 583 -1072 0 1
rlabel polysilicon 583 -1078 583 -1078 0 3
rlabel polysilicon 590 -1072 590 -1072 0 1
rlabel polysilicon 590 -1078 590 -1078 0 3
rlabel polysilicon 597 -1072 597 -1072 0 1
rlabel polysilicon 600 -1072 600 -1072 0 2
rlabel polysilicon 600 -1078 600 -1078 0 4
rlabel polysilicon 604 -1072 604 -1072 0 1
rlabel polysilicon 604 -1078 604 -1078 0 3
rlabel polysilicon 611 -1072 611 -1072 0 1
rlabel polysilicon 611 -1078 611 -1078 0 3
rlabel polysilicon 618 -1072 618 -1072 0 1
rlabel polysilicon 621 -1072 621 -1072 0 2
rlabel polysilicon 621 -1078 621 -1078 0 4
rlabel polysilicon 625 -1072 625 -1072 0 1
rlabel polysilicon 625 -1078 625 -1078 0 3
rlabel polysilicon 632 -1078 632 -1078 0 3
rlabel polysilicon 639 -1072 639 -1072 0 1
rlabel polysilicon 639 -1078 639 -1078 0 3
rlabel polysilicon 646 -1072 646 -1072 0 1
rlabel polysilicon 646 -1078 646 -1078 0 3
rlabel polysilicon 653 -1072 653 -1072 0 1
rlabel polysilicon 653 -1078 653 -1078 0 3
rlabel polysilicon 660 -1072 660 -1072 0 1
rlabel polysilicon 660 -1078 660 -1078 0 3
rlabel polysilicon 667 -1072 667 -1072 0 1
rlabel polysilicon 667 -1078 667 -1078 0 3
rlabel polysilicon 674 -1072 674 -1072 0 1
rlabel polysilicon 674 -1078 674 -1078 0 3
rlabel polysilicon 681 -1072 681 -1072 0 1
rlabel polysilicon 681 -1078 681 -1078 0 3
rlabel polysilicon 688 -1072 688 -1072 0 1
rlabel polysilicon 691 -1072 691 -1072 0 2
rlabel polysilicon 688 -1078 688 -1078 0 3
rlabel polysilicon 695 -1072 695 -1072 0 1
rlabel polysilicon 695 -1078 695 -1078 0 3
rlabel polysilicon 702 -1072 702 -1072 0 1
rlabel polysilicon 702 -1078 702 -1078 0 3
rlabel polysilicon 709 -1072 709 -1072 0 1
rlabel polysilicon 709 -1078 709 -1078 0 3
rlabel polysilicon 716 -1072 716 -1072 0 1
rlabel polysilicon 716 -1078 716 -1078 0 3
rlabel polysilicon 723 -1072 723 -1072 0 1
rlabel polysilicon 723 -1078 723 -1078 0 3
rlabel polysilicon 733 -1072 733 -1072 0 2
rlabel polysilicon 733 -1078 733 -1078 0 4
rlabel polysilicon 737 -1072 737 -1072 0 1
rlabel polysilicon 737 -1078 737 -1078 0 3
rlabel polysilicon 744 -1072 744 -1072 0 1
rlabel polysilicon 744 -1078 744 -1078 0 3
rlabel polysilicon 751 -1072 751 -1072 0 1
rlabel polysilicon 751 -1078 751 -1078 0 3
rlabel polysilicon 758 -1078 758 -1078 0 3
rlabel polysilicon 765 -1072 765 -1072 0 1
rlabel polysilicon 765 -1078 765 -1078 0 3
rlabel polysilicon 772 -1072 772 -1072 0 1
rlabel polysilicon 772 -1078 772 -1078 0 3
rlabel polysilicon 779 -1072 779 -1072 0 1
rlabel polysilicon 779 -1078 779 -1078 0 3
rlabel polysilicon 786 -1072 786 -1072 0 1
rlabel polysilicon 786 -1078 786 -1078 0 3
rlabel polysilicon 793 -1072 793 -1072 0 1
rlabel polysilicon 793 -1078 793 -1078 0 3
rlabel polysilicon 800 -1072 800 -1072 0 1
rlabel polysilicon 800 -1078 800 -1078 0 3
rlabel polysilicon 810 -1072 810 -1072 0 2
rlabel polysilicon 810 -1078 810 -1078 0 4
rlabel polysilicon 814 -1072 814 -1072 0 1
rlabel polysilicon 814 -1078 814 -1078 0 3
rlabel polysilicon 821 -1072 821 -1072 0 1
rlabel polysilicon 821 -1078 821 -1078 0 3
rlabel polysilicon 828 -1072 828 -1072 0 1
rlabel polysilicon 828 -1078 828 -1078 0 3
rlabel polysilicon 835 -1072 835 -1072 0 1
rlabel polysilicon 835 -1078 835 -1078 0 3
rlabel polysilicon 842 -1072 842 -1072 0 1
rlabel polysilicon 842 -1078 842 -1078 0 3
rlabel polysilicon 849 -1072 849 -1072 0 1
rlabel polysilicon 849 -1078 849 -1078 0 3
rlabel polysilicon 856 -1072 856 -1072 0 1
rlabel polysilicon 856 -1078 856 -1078 0 3
rlabel polysilicon 863 -1072 863 -1072 0 1
rlabel polysilicon 863 -1078 863 -1078 0 3
rlabel polysilicon 870 -1072 870 -1072 0 1
rlabel polysilicon 870 -1078 870 -1078 0 3
rlabel polysilicon 877 -1072 877 -1072 0 1
rlabel polysilicon 877 -1078 877 -1078 0 3
rlabel polysilicon 884 -1072 884 -1072 0 1
rlabel polysilicon 884 -1078 884 -1078 0 3
rlabel polysilicon 891 -1072 891 -1072 0 1
rlabel polysilicon 891 -1078 891 -1078 0 3
rlabel polysilicon 898 -1072 898 -1072 0 1
rlabel polysilicon 898 -1078 898 -1078 0 3
rlabel polysilicon 905 -1072 905 -1072 0 1
rlabel polysilicon 905 -1078 905 -1078 0 3
rlabel polysilicon 912 -1072 912 -1072 0 1
rlabel polysilicon 912 -1078 912 -1078 0 3
rlabel polysilicon 919 -1072 919 -1072 0 1
rlabel polysilicon 919 -1078 919 -1078 0 3
rlabel polysilicon 926 -1072 926 -1072 0 1
rlabel polysilicon 926 -1078 926 -1078 0 3
rlabel polysilicon 933 -1072 933 -1072 0 1
rlabel polysilicon 933 -1078 933 -1078 0 3
rlabel polysilicon 940 -1072 940 -1072 0 1
rlabel polysilicon 940 -1078 940 -1078 0 3
rlabel polysilicon 947 -1072 947 -1072 0 1
rlabel polysilicon 947 -1078 947 -1078 0 3
rlabel polysilicon 954 -1072 954 -1072 0 1
rlabel polysilicon 957 -1078 957 -1078 0 4
rlabel polysilicon 961 -1072 961 -1072 0 1
rlabel polysilicon 961 -1078 961 -1078 0 3
rlabel polysilicon 968 -1072 968 -1072 0 1
rlabel polysilicon 968 -1078 968 -1078 0 3
rlabel polysilicon 975 -1072 975 -1072 0 1
rlabel polysilicon 975 -1078 975 -1078 0 3
rlabel polysilicon 982 -1072 982 -1072 0 1
rlabel polysilicon 982 -1078 982 -1078 0 3
rlabel polysilicon 989 -1072 989 -1072 0 1
rlabel polysilicon 989 -1078 989 -1078 0 3
rlabel polysilicon 996 -1072 996 -1072 0 1
rlabel polysilicon 996 -1078 996 -1078 0 3
rlabel polysilicon 1003 -1072 1003 -1072 0 1
rlabel polysilicon 1003 -1078 1003 -1078 0 3
rlabel polysilicon 1010 -1072 1010 -1072 0 1
rlabel polysilicon 1010 -1078 1010 -1078 0 3
rlabel polysilicon 1017 -1072 1017 -1072 0 1
rlabel polysilicon 1017 -1078 1017 -1078 0 3
rlabel polysilicon 1024 -1072 1024 -1072 0 1
rlabel polysilicon 1024 -1078 1024 -1078 0 3
rlabel polysilicon 1031 -1072 1031 -1072 0 1
rlabel polysilicon 1031 -1078 1031 -1078 0 3
rlabel polysilicon 1038 -1072 1038 -1072 0 1
rlabel polysilicon 1041 -1078 1041 -1078 0 4
rlabel polysilicon 1045 -1072 1045 -1072 0 1
rlabel polysilicon 1045 -1078 1045 -1078 0 3
rlabel polysilicon 1052 -1072 1052 -1072 0 1
rlabel polysilicon 1052 -1078 1052 -1078 0 3
rlabel polysilicon 1059 -1072 1059 -1072 0 1
rlabel polysilicon 1066 -1072 1066 -1072 0 1
rlabel polysilicon 1069 -1072 1069 -1072 0 2
rlabel polysilicon 1066 -1078 1066 -1078 0 3
rlabel polysilicon 1073 -1072 1073 -1072 0 1
rlabel polysilicon 1073 -1078 1073 -1078 0 3
rlabel polysilicon 1080 -1072 1080 -1072 0 1
rlabel polysilicon 1080 -1078 1080 -1078 0 3
rlabel polysilicon 1087 -1072 1087 -1072 0 1
rlabel polysilicon 1087 -1078 1087 -1078 0 3
rlabel polysilicon 1094 -1072 1094 -1072 0 1
rlabel polysilicon 1094 -1078 1094 -1078 0 3
rlabel polysilicon 1122 -1072 1122 -1072 0 1
rlabel polysilicon 1122 -1078 1122 -1078 0 3
rlabel polysilicon 1185 -1072 1185 -1072 0 1
rlabel polysilicon 1185 -1078 1185 -1078 0 3
rlabel polysilicon 23 -1161 23 -1161 0 3
rlabel polysilicon 30 -1155 30 -1155 0 1
rlabel polysilicon 30 -1161 30 -1161 0 3
rlabel polysilicon 37 -1155 37 -1155 0 1
rlabel polysilicon 37 -1161 37 -1161 0 3
rlabel polysilicon 44 -1155 44 -1155 0 1
rlabel polysilicon 44 -1161 44 -1161 0 3
rlabel polysilicon 51 -1155 51 -1155 0 1
rlabel polysilicon 51 -1161 51 -1161 0 3
rlabel polysilicon 58 -1155 58 -1155 0 1
rlabel polysilicon 58 -1161 58 -1161 0 3
rlabel polysilicon 65 -1155 65 -1155 0 1
rlabel polysilicon 65 -1161 65 -1161 0 3
rlabel polysilicon 72 -1155 72 -1155 0 1
rlabel polysilicon 72 -1161 72 -1161 0 3
rlabel polysilicon 82 -1155 82 -1155 0 2
rlabel polysilicon 82 -1161 82 -1161 0 4
rlabel polysilicon 89 -1161 89 -1161 0 4
rlabel polysilicon 93 -1155 93 -1155 0 1
rlabel polysilicon 93 -1161 93 -1161 0 3
rlabel polysilicon 100 -1155 100 -1155 0 1
rlabel polysilicon 100 -1161 100 -1161 0 3
rlabel polysilicon 107 -1155 107 -1155 0 1
rlabel polysilicon 107 -1161 107 -1161 0 3
rlabel polysilicon 117 -1155 117 -1155 0 2
rlabel polysilicon 114 -1161 114 -1161 0 3
rlabel polysilicon 117 -1161 117 -1161 0 4
rlabel polysilicon 121 -1155 121 -1155 0 1
rlabel polysilicon 121 -1161 121 -1161 0 3
rlabel polysilicon 128 -1155 128 -1155 0 1
rlabel polysilicon 131 -1161 131 -1161 0 4
rlabel polysilicon 135 -1155 135 -1155 0 1
rlabel polysilicon 138 -1161 138 -1161 0 4
rlabel polysilicon 142 -1155 142 -1155 0 1
rlabel polysilicon 142 -1161 142 -1161 0 3
rlabel polysilicon 149 -1155 149 -1155 0 1
rlabel polysilicon 149 -1161 149 -1161 0 3
rlabel polysilicon 156 -1155 156 -1155 0 1
rlabel polysilicon 156 -1161 156 -1161 0 3
rlabel polysilicon 166 -1155 166 -1155 0 2
rlabel polysilicon 163 -1161 163 -1161 0 3
rlabel polysilicon 166 -1161 166 -1161 0 4
rlabel polysilicon 170 -1155 170 -1155 0 1
rlabel polysilicon 170 -1161 170 -1161 0 3
rlabel polysilicon 177 -1155 177 -1155 0 1
rlabel polysilicon 177 -1161 177 -1161 0 3
rlabel polysilicon 184 -1155 184 -1155 0 1
rlabel polysilicon 187 -1155 187 -1155 0 2
rlabel polysilicon 187 -1161 187 -1161 0 4
rlabel polysilicon 191 -1155 191 -1155 0 1
rlabel polysilicon 191 -1161 191 -1161 0 3
rlabel polysilicon 198 -1161 198 -1161 0 3
rlabel polysilicon 205 -1155 205 -1155 0 1
rlabel polysilicon 205 -1161 205 -1161 0 3
rlabel polysilicon 212 -1155 212 -1155 0 1
rlabel polysilicon 212 -1161 212 -1161 0 3
rlabel polysilicon 219 -1155 219 -1155 0 1
rlabel polysilicon 219 -1161 219 -1161 0 3
rlabel polysilicon 226 -1155 226 -1155 0 1
rlabel polysilicon 229 -1161 229 -1161 0 4
rlabel polysilicon 233 -1155 233 -1155 0 1
rlabel polysilicon 233 -1161 233 -1161 0 3
rlabel polysilicon 240 -1155 240 -1155 0 1
rlabel polysilicon 240 -1161 240 -1161 0 3
rlabel polysilicon 247 -1155 247 -1155 0 1
rlabel polysilicon 247 -1161 247 -1161 0 3
rlabel polysilicon 254 -1155 254 -1155 0 1
rlabel polysilicon 254 -1161 254 -1161 0 3
rlabel polysilicon 261 -1155 261 -1155 0 1
rlabel polysilicon 261 -1161 261 -1161 0 3
rlabel polysilicon 268 -1155 268 -1155 0 1
rlabel polysilicon 268 -1161 268 -1161 0 3
rlabel polysilicon 275 -1155 275 -1155 0 1
rlabel polysilicon 275 -1161 275 -1161 0 3
rlabel polysilicon 282 -1155 282 -1155 0 1
rlabel polysilicon 285 -1161 285 -1161 0 4
rlabel polysilicon 289 -1155 289 -1155 0 1
rlabel polysilicon 289 -1161 289 -1161 0 3
rlabel polysilicon 296 -1155 296 -1155 0 1
rlabel polysilicon 296 -1161 296 -1161 0 3
rlabel polysilicon 306 -1155 306 -1155 0 2
rlabel polysilicon 306 -1161 306 -1161 0 4
rlabel polysilicon 310 -1155 310 -1155 0 1
rlabel polysilicon 310 -1161 310 -1161 0 3
rlabel polysilicon 317 -1155 317 -1155 0 1
rlabel polysilicon 317 -1161 317 -1161 0 3
rlabel polysilicon 324 -1155 324 -1155 0 1
rlabel polysilicon 324 -1161 324 -1161 0 3
rlabel polysilicon 331 -1155 331 -1155 0 1
rlabel polysilicon 338 -1155 338 -1155 0 1
rlabel polysilicon 338 -1161 338 -1161 0 3
rlabel polysilicon 345 -1155 345 -1155 0 1
rlabel polysilicon 345 -1161 345 -1161 0 3
rlabel polysilicon 352 -1155 352 -1155 0 1
rlabel polysilicon 352 -1161 352 -1161 0 3
rlabel polysilicon 359 -1155 359 -1155 0 1
rlabel polysilicon 359 -1161 359 -1161 0 3
rlabel polysilicon 366 -1155 366 -1155 0 1
rlabel polysilicon 366 -1161 366 -1161 0 3
rlabel polysilicon 373 -1155 373 -1155 0 1
rlabel polysilicon 373 -1161 373 -1161 0 3
rlabel polysilicon 380 -1155 380 -1155 0 1
rlabel polysilicon 380 -1161 380 -1161 0 3
rlabel polysilicon 387 -1155 387 -1155 0 1
rlabel polysilicon 387 -1161 387 -1161 0 3
rlabel polysilicon 394 -1155 394 -1155 0 1
rlabel polysilicon 394 -1161 394 -1161 0 3
rlabel polysilicon 401 -1155 401 -1155 0 1
rlabel polysilicon 401 -1161 401 -1161 0 3
rlabel polysilicon 408 -1155 408 -1155 0 1
rlabel polysilicon 408 -1161 408 -1161 0 3
rlabel polysilicon 415 -1155 415 -1155 0 1
rlabel polysilicon 418 -1155 418 -1155 0 2
rlabel polysilicon 415 -1161 415 -1161 0 3
rlabel polysilicon 422 -1155 422 -1155 0 1
rlabel polysilicon 422 -1161 422 -1161 0 3
rlabel polysilicon 429 -1155 429 -1155 0 1
rlabel polysilicon 429 -1161 429 -1161 0 3
rlabel polysilicon 436 -1155 436 -1155 0 1
rlabel polysilicon 436 -1161 436 -1161 0 3
rlabel polysilicon 446 -1155 446 -1155 0 2
rlabel polysilicon 446 -1161 446 -1161 0 4
rlabel polysilicon 450 -1155 450 -1155 0 1
rlabel polysilicon 450 -1161 450 -1161 0 3
rlabel polysilicon 457 -1155 457 -1155 0 1
rlabel polysilicon 457 -1161 457 -1161 0 3
rlabel polysilicon 464 -1155 464 -1155 0 1
rlabel polysilicon 464 -1161 464 -1161 0 3
rlabel polysilicon 471 -1155 471 -1155 0 1
rlabel polysilicon 471 -1161 471 -1161 0 3
rlabel polysilicon 478 -1155 478 -1155 0 1
rlabel polysilicon 478 -1161 478 -1161 0 3
rlabel polysilicon 485 -1155 485 -1155 0 1
rlabel polysilicon 485 -1161 485 -1161 0 3
rlabel polysilicon 492 -1155 492 -1155 0 1
rlabel polysilicon 492 -1161 492 -1161 0 3
rlabel polysilicon 499 -1155 499 -1155 0 1
rlabel polysilicon 499 -1161 499 -1161 0 3
rlabel polysilicon 506 -1161 506 -1161 0 3
rlabel polysilicon 509 -1161 509 -1161 0 4
rlabel polysilicon 513 -1155 513 -1155 0 1
rlabel polysilicon 513 -1161 513 -1161 0 3
rlabel polysilicon 520 -1155 520 -1155 0 1
rlabel polysilicon 520 -1161 520 -1161 0 3
rlabel polysilicon 527 -1155 527 -1155 0 1
rlabel polysilicon 527 -1161 527 -1161 0 3
rlabel polysilicon 534 -1155 534 -1155 0 1
rlabel polysilicon 534 -1161 534 -1161 0 3
rlabel polysilicon 541 -1155 541 -1155 0 1
rlabel polysilicon 541 -1161 541 -1161 0 3
rlabel polysilicon 548 -1155 548 -1155 0 1
rlabel polysilicon 551 -1155 551 -1155 0 2
rlabel polysilicon 551 -1161 551 -1161 0 4
rlabel polysilicon 555 -1155 555 -1155 0 1
rlabel polysilicon 555 -1161 555 -1161 0 3
rlabel polysilicon 562 -1155 562 -1155 0 1
rlabel polysilicon 562 -1161 562 -1161 0 3
rlabel polysilicon 569 -1155 569 -1155 0 1
rlabel polysilicon 569 -1161 569 -1161 0 3
rlabel polysilicon 576 -1155 576 -1155 0 1
rlabel polysilicon 576 -1161 576 -1161 0 3
rlabel polysilicon 583 -1155 583 -1155 0 1
rlabel polysilicon 586 -1155 586 -1155 0 2
rlabel polysilicon 583 -1161 583 -1161 0 3
rlabel polysilicon 586 -1161 586 -1161 0 4
rlabel polysilicon 590 -1155 590 -1155 0 1
rlabel polysilicon 590 -1161 590 -1161 0 3
rlabel polysilicon 597 -1155 597 -1155 0 1
rlabel polysilicon 597 -1161 597 -1161 0 3
rlabel polysilicon 607 -1155 607 -1155 0 2
rlabel polysilicon 604 -1161 604 -1161 0 3
rlabel polysilicon 607 -1161 607 -1161 0 4
rlabel polysilicon 611 -1155 611 -1155 0 1
rlabel polysilicon 611 -1161 611 -1161 0 3
rlabel polysilicon 618 -1155 618 -1155 0 1
rlabel polysilicon 618 -1161 618 -1161 0 3
rlabel polysilicon 628 -1155 628 -1155 0 2
rlabel polysilicon 625 -1161 625 -1161 0 3
rlabel polysilicon 632 -1155 632 -1155 0 1
rlabel polysilicon 632 -1161 632 -1161 0 3
rlabel polysilicon 639 -1155 639 -1155 0 1
rlabel polysilicon 639 -1161 639 -1161 0 3
rlabel polysilicon 646 -1155 646 -1155 0 1
rlabel polysilicon 646 -1161 646 -1161 0 3
rlabel polysilicon 653 -1155 653 -1155 0 1
rlabel polysilicon 656 -1161 656 -1161 0 4
rlabel polysilicon 660 -1155 660 -1155 0 1
rlabel polysilicon 660 -1161 660 -1161 0 3
rlabel polysilicon 667 -1155 667 -1155 0 1
rlabel polysilicon 670 -1155 670 -1155 0 2
rlabel polysilicon 667 -1161 667 -1161 0 3
rlabel polysilicon 674 -1155 674 -1155 0 1
rlabel polysilicon 674 -1161 674 -1161 0 3
rlabel polysilicon 681 -1155 681 -1155 0 1
rlabel polysilicon 681 -1161 681 -1161 0 3
rlabel polysilicon 688 -1155 688 -1155 0 1
rlabel polysilicon 688 -1161 688 -1161 0 3
rlabel polysilicon 695 -1155 695 -1155 0 1
rlabel polysilicon 695 -1161 695 -1161 0 3
rlabel polysilicon 702 -1155 702 -1155 0 1
rlabel polysilicon 702 -1161 702 -1161 0 3
rlabel polysilicon 709 -1155 709 -1155 0 1
rlabel polysilicon 709 -1161 709 -1161 0 3
rlabel polysilicon 716 -1155 716 -1155 0 1
rlabel polysilicon 716 -1161 716 -1161 0 3
rlabel polysilicon 723 -1155 723 -1155 0 1
rlabel polysilicon 723 -1161 723 -1161 0 3
rlabel polysilicon 730 -1155 730 -1155 0 1
rlabel polysilicon 730 -1161 730 -1161 0 3
rlabel polysilicon 737 -1155 737 -1155 0 1
rlabel polysilicon 737 -1161 737 -1161 0 3
rlabel polysilicon 744 -1155 744 -1155 0 1
rlabel polysilicon 744 -1161 744 -1161 0 3
rlabel polysilicon 751 -1155 751 -1155 0 1
rlabel polysilicon 751 -1161 751 -1161 0 3
rlabel polysilicon 758 -1155 758 -1155 0 1
rlabel polysilicon 758 -1161 758 -1161 0 3
rlabel polysilicon 765 -1155 765 -1155 0 1
rlabel polysilicon 765 -1161 765 -1161 0 3
rlabel polysilicon 772 -1155 772 -1155 0 1
rlabel polysilicon 772 -1161 772 -1161 0 3
rlabel polysilicon 779 -1155 779 -1155 0 1
rlabel polysilicon 779 -1161 779 -1161 0 3
rlabel polysilicon 786 -1155 786 -1155 0 1
rlabel polysilicon 786 -1161 786 -1161 0 3
rlabel polysilicon 793 -1155 793 -1155 0 1
rlabel polysilicon 793 -1161 793 -1161 0 3
rlabel polysilicon 800 -1155 800 -1155 0 1
rlabel polysilicon 800 -1161 800 -1161 0 3
rlabel polysilicon 807 -1155 807 -1155 0 1
rlabel polysilicon 810 -1155 810 -1155 0 2
rlabel polysilicon 810 -1161 810 -1161 0 4
rlabel polysilicon 814 -1155 814 -1155 0 1
rlabel polysilicon 814 -1161 814 -1161 0 3
rlabel polysilicon 821 -1155 821 -1155 0 1
rlabel polysilicon 821 -1161 821 -1161 0 3
rlabel polysilicon 828 -1155 828 -1155 0 1
rlabel polysilicon 828 -1161 828 -1161 0 3
rlabel polysilicon 835 -1155 835 -1155 0 1
rlabel polysilicon 835 -1161 835 -1161 0 3
rlabel polysilicon 842 -1155 842 -1155 0 1
rlabel polysilicon 842 -1161 842 -1161 0 3
rlabel polysilicon 852 -1155 852 -1155 0 2
rlabel polysilicon 856 -1155 856 -1155 0 1
rlabel polysilicon 856 -1161 856 -1161 0 3
rlabel polysilicon 863 -1155 863 -1155 0 1
rlabel polysilicon 863 -1161 863 -1161 0 3
rlabel polysilicon 870 -1155 870 -1155 0 1
rlabel polysilicon 870 -1161 870 -1161 0 3
rlabel polysilicon 877 -1155 877 -1155 0 1
rlabel polysilicon 877 -1161 877 -1161 0 3
rlabel polysilicon 884 -1155 884 -1155 0 1
rlabel polysilicon 884 -1161 884 -1161 0 3
rlabel polysilicon 891 -1155 891 -1155 0 1
rlabel polysilicon 891 -1161 891 -1161 0 3
rlabel polysilicon 898 -1155 898 -1155 0 1
rlabel polysilicon 898 -1161 898 -1161 0 3
rlabel polysilicon 905 -1155 905 -1155 0 1
rlabel polysilicon 905 -1161 905 -1161 0 3
rlabel polysilicon 912 -1155 912 -1155 0 1
rlabel polysilicon 912 -1161 912 -1161 0 3
rlabel polysilicon 919 -1155 919 -1155 0 1
rlabel polysilicon 919 -1161 919 -1161 0 3
rlabel polysilicon 926 -1155 926 -1155 0 1
rlabel polysilicon 926 -1161 926 -1161 0 3
rlabel polysilicon 933 -1155 933 -1155 0 1
rlabel polysilicon 936 -1161 936 -1161 0 4
rlabel polysilicon 940 -1155 940 -1155 0 1
rlabel polysilicon 940 -1161 940 -1161 0 3
rlabel polysilicon 947 -1155 947 -1155 0 1
rlabel polysilicon 947 -1161 947 -1161 0 3
rlabel polysilicon 954 -1155 954 -1155 0 1
rlabel polysilicon 954 -1161 954 -1161 0 3
rlabel polysilicon 961 -1155 961 -1155 0 1
rlabel polysilicon 961 -1161 961 -1161 0 3
rlabel polysilicon 968 -1155 968 -1155 0 1
rlabel polysilicon 968 -1161 968 -1161 0 3
rlabel polysilicon 978 -1155 978 -1155 0 2
rlabel polysilicon 975 -1161 975 -1161 0 3
rlabel polysilicon 978 -1161 978 -1161 0 4
rlabel polysilicon 982 -1155 982 -1155 0 1
rlabel polysilicon 982 -1161 982 -1161 0 3
rlabel polysilicon 989 -1155 989 -1155 0 1
rlabel polysilicon 989 -1161 989 -1161 0 3
rlabel polysilicon 996 -1155 996 -1155 0 1
rlabel polysilicon 996 -1161 996 -1161 0 3
rlabel polysilicon 1003 -1155 1003 -1155 0 1
rlabel polysilicon 1006 -1155 1006 -1155 0 2
rlabel polysilicon 1010 -1155 1010 -1155 0 1
rlabel polysilicon 1010 -1161 1010 -1161 0 3
rlabel polysilicon 1017 -1155 1017 -1155 0 1
rlabel polysilicon 1017 -1161 1017 -1161 0 3
rlabel polysilicon 1024 -1155 1024 -1155 0 1
rlabel polysilicon 1024 -1161 1024 -1161 0 3
rlabel polysilicon 1031 -1155 1031 -1155 0 1
rlabel polysilicon 1031 -1161 1031 -1161 0 3
rlabel polysilicon 1038 -1155 1038 -1155 0 1
rlabel polysilicon 1038 -1161 1038 -1161 0 3
rlabel polysilicon 1048 -1155 1048 -1155 0 2
rlabel polysilicon 1059 -1155 1059 -1155 0 1
rlabel polysilicon 1059 -1161 1059 -1161 0 3
rlabel polysilicon 1066 -1155 1066 -1155 0 1
rlabel polysilicon 1066 -1161 1066 -1161 0 3
rlabel polysilicon 1080 -1155 1080 -1155 0 1
rlabel polysilicon 1080 -1161 1080 -1161 0 3
rlabel polysilicon 1087 -1155 1087 -1155 0 1
rlabel polysilicon 1087 -1161 1087 -1161 0 3
rlabel polysilicon 1108 -1155 1108 -1155 0 1
rlabel polysilicon 1108 -1161 1108 -1161 0 3
rlabel polysilicon 1188 -1155 1188 -1155 0 2
rlabel polysilicon 16 -1230 16 -1230 0 1
rlabel polysilicon 16 -1236 16 -1236 0 3
rlabel polysilicon 23 -1230 23 -1230 0 1
rlabel polysilicon 26 -1230 26 -1230 0 2
rlabel polysilicon 30 -1230 30 -1230 0 1
rlabel polysilicon 30 -1236 30 -1236 0 3
rlabel polysilicon 37 -1230 37 -1230 0 1
rlabel polysilicon 37 -1236 37 -1236 0 3
rlabel polysilicon 44 -1236 44 -1236 0 3
rlabel polysilicon 47 -1236 47 -1236 0 4
rlabel polysilicon 51 -1230 51 -1230 0 1
rlabel polysilicon 51 -1236 51 -1236 0 3
rlabel polysilicon 58 -1230 58 -1230 0 1
rlabel polysilicon 61 -1230 61 -1230 0 2
rlabel polysilicon 65 -1230 65 -1230 0 1
rlabel polysilicon 68 -1236 68 -1236 0 4
rlabel polysilicon 72 -1230 72 -1230 0 1
rlabel polysilicon 72 -1236 72 -1236 0 3
rlabel polysilicon 79 -1230 79 -1230 0 1
rlabel polysilicon 79 -1236 79 -1236 0 3
rlabel polysilicon 93 -1230 93 -1230 0 1
rlabel polysilicon 93 -1236 93 -1236 0 3
rlabel polysilicon 100 -1230 100 -1230 0 1
rlabel polysilicon 100 -1236 100 -1236 0 3
rlabel polysilicon 107 -1230 107 -1230 0 1
rlabel polysilicon 107 -1236 107 -1236 0 3
rlabel polysilicon 117 -1236 117 -1236 0 4
rlabel polysilicon 121 -1230 121 -1230 0 1
rlabel polysilicon 121 -1236 121 -1236 0 3
rlabel polysilicon 128 -1230 128 -1230 0 1
rlabel polysilicon 128 -1236 128 -1236 0 3
rlabel polysilicon 135 -1230 135 -1230 0 1
rlabel polysilicon 135 -1236 135 -1236 0 3
rlabel polysilicon 142 -1230 142 -1230 0 1
rlabel polysilicon 142 -1236 142 -1236 0 3
rlabel polysilicon 152 -1230 152 -1230 0 2
rlabel polysilicon 149 -1236 149 -1236 0 3
rlabel polysilicon 152 -1236 152 -1236 0 4
rlabel polysilicon 156 -1230 156 -1230 0 1
rlabel polysilicon 156 -1236 156 -1236 0 3
rlabel polysilicon 163 -1230 163 -1230 0 1
rlabel polysilicon 163 -1236 163 -1236 0 3
rlabel polysilicon 170 -1230 170 -1230 0 1
rlabel polysilicon 170 -1236 170 -1236 0 3
rlabel polysilicon 177 -1236 177 -1236 0 3
rlabel polysilicon 180 -1236 180 -1236 0 4
rlabel polysilicon 184 -1230 184 -1230 0 1
rlabel polysilicon 184 -1236 184 -1236 0 3
rlabel polysilicon 191 -1230 191 -1230 0 1
rlabel polysilicon 191 -1236 191 -1236 0 3
rlabel polysilicon 198 -1230 198 -1230 0 1
rlabel polysilicon 198 -1236 198 -1236 0 3
rlabel polysilicon 205 -1230 205 -1230 0 1
rlabel polysilicon 205 -1236 205 -1236 0 3
rlabel polysilicon 212 -1230 212 -1230 0 1
rlabel polysilicon 212 -1236 212 -1236 0 3
rlabel polysilicon 219 -1230 219 -1230 0 1
rlabel polysilicon 219 -1236 219 -1236 0 3
rlabel polysilicon 226 -1230 226 -1230 0 1
rlabel polysilicon 226 -1236 226 -1236 0 3
rlabel polysilicon 233 -1230 233 -1230 0 1
rlabel polysilicon 233 -1236 233 -1236 0 3
rlabel polysilicon 240 -1230 240 -1230 0 1
rlabel polysilicon 240 -1236 240 -1236 0 3
rlabel polysilicon 247 -1230 247 -1230 0 1
rlabel polysilicon 247 -1236 247 -1236 0 3
rlabel polysilicon 254 -1230 254 -1230 0 1
rlabel polysilicon 254 -1236 254 -1236 0 3
rlabel polysilicon 264 -1236 264 -1236 0 4
rlabel polysilicon 268 -1230 268 -1230 0 1
rlabel polysilicon 268 -1236 268 -1236 0 3
rlabel polysilicon 275 -1230 275 -1230 0 1
rlabel polysilicon 275 -1236 275 -1236 0 3
rlabel polysilicon 282 -1230 282 -1230 0 1
rlabel polysilicon 282 -1236 282 -1236 0 3
rlabel polysilicon 289 -1230 289 -1230 0 1
rlabel polysilicon 289 -1236 289 -1236 0 3
rlabel polysilicon 296 -1230 296 -1230 0 1
rlabel polysilicon 296 -1236 296 -1236 0 3
rlabel polysilicon 303 -1230 303 -1230 0 1
rlabel polysilicon 303 -1236 303 -1236 0 3
rlabel polysilicon 310 -1230 310 -1230 0 1
rlabel polysilicon 310 -1236 310 -1236 0 3
rlabel polysilicon 317 -1230 317 -1230 0 1
rlabel polysilicon 317 -1236 317 -1236 0 3
rlabel polysilicon 320 -1236 320 -1236 0 4
rlabel polysilicon 324 -1230 324 -1230 0 1
rlabel polysilicon 324 -1236 324 -1236 0 3
rlabel polysilicon 331 -1230 331 -1230 0 1
rlabel polysilicon 331 -1236 331 -1236 0 3
rlabel polysilicon 338 -1230 338 -1230 0 1
rlabel polysilicon 338 -1236 338 -1236 0 3
rlabel polysilicon 345 -1230 345 -1230 0 1
rlabel polysilicon 345 -1236 345 -1236 0 3
rlabel polysilicon 352 -1230 352 -1230 0 1
rlabel polysilicon 352 -1236 352 -1236 0 3
rlabel polysilicon 359 -1230 359 -1230 0 1
rlabel polysilicon 359 -1236 359 -1236 0 3
rlabel polysilicon 366 -1230 366 -1230 0 1
rlabel polysilicon 366 -1236 366 -1236 0 3
rlabel polysilicon 373 -1230 373 -1230 0 1
rlabel polysilicon 376 -1236 376 -1236 0 4
rlabel polysilicon 383 -1230 383 -1230 0 2
rlabel polysilicon 380 -1236 380 -1236 0 3
rlabel polysilicon 387 -1236 387 -1236 0 3
rlabel polysilicon 390 -1236 390 -1236 0 4
rlabel polysilicon 394 -1230 394 -1230 0 1
rlabel polysilicon 394 -1236 394 -1236 0 3
rlabel polysilicon 401 -1230 401 -1230 0 1
rlabel polysilicon 401 -1236 401 -1236 0 3
rlabel polysilicon 408 -1230 408 -1230 0 1
rlabel polysilicon 408 -1236 408 -1236 0 3
rlabel polysilicon 415 -1230 415 -1230 0 1
rlabel polysilicon 415 -1236 415 -1236 0 3
rlabel polysilicon 422 -1230 422 -1230 0 1
rlabel polysilicon 422 -1236 422 -1236 0 3
rlabel polysilicon 429 -1230 429 -1230 0 1
rlabel polysilicon 429 -1236 429 -1236 0 3
rlabel polysilicon 436 -1230 436 -1230 0 1
rlabel polysilicon 436 -1236 436 -1236 0 3
rlabel polysilicon 443 -1230 443 -1230 0 1
rlabel polysilicon 446 -1236 446 -1236 0 4
rlabel polysilicon 450 -1230 450 -1230 0 1
rlabel polysilicon 450 -1236 450 -1236 0 3
rlabel polysilicon 457 -1230 457 -1230 0 1
rlabel polysilicon 457 -1236 457 -1236 0 3
rlabel polysilicon 464 -1230 464 -1230 0 1
rlabel polysilicon 464 -1236 464 -1236 0 3
rlabel polysilicon 471 -1230 471 -1230 0 1
rlabel polysilicon 471 -1236 471 -1236 0 3
rlabel polysilicon 478 -1230 478 -1230 0 1
rlabel polysilicon 478 -1236 478 -1236 0 3
rlabel polysilicon 485 -1230 485 -1230 0 1
rlabel polysilicon 485 -1236 485 -1236 0 3
rlabel polysilicon 492 -1230 492 -1230 0 1
rlabel polysilicon 492 -1236 492 -1236 0 3
rlabel polysilicon 499 -1230 499 -1230 0 1
rlabel polysilicon 499 -1236 499 -1236 0 3
rlabel polysilicon 509 -1230 509 -1230 0 2
rlabel polysilicon 506 -1236 506 -1236 0 3
rlabel polysilicon 509 -1236 509 -1236 0 4
rlabel polysilicon 513 -1230 513 -1230 0 1
rlabel polysilicon 513 -1236 513 -1236 0 3
rlabel polysilicon 520 -1230 520 -1230 0 1
rlabel polysilicon 520 -1236 520 -1236 0 3
rlabel polysilicon 527 -1230 527 -1230 0 1
rlabel polysilicon 527 -1236 527 -1236 0 3
rlabel polysilicon 534 -1230 534 -1230 0 1
rlabel polysilicon 534 -1236 534 -1236 0 3
rlabel polysilicon 544 -1230 544 -1230 0 2
rlabel polysilicon 544 -1236 544 -1236 0 4
rlabel polysilicon 548 -1230 548 -1230 0 1
rlabel polysilicon 548 -1236 548 -1236 0 3
rlabel polysilicon 555 -1230 555 -1230 0 1
rlabel polysilicon 555 -1236 555 -1236 0 3
rlabel polysilicon 562 -1230 562 -1230 0 1
rlabel polysilicon 565 -1230 565 -1230 0 2
rlabel polysilicon 562 -1236 562 -1236 0 3
rlabel polysilicon 565 -1236 565 -1236 0 4
rlabel polysilicon 569 -1230 569 -1230 0 1
rlabel polysilicon 569 -1236 569 -1236 0 3
rlabel polysilicon 572 -1236 572 -1236 0 4
rlabel polysilicon 576 -1230 576 -1230 0 1
rlabel polysilicon 576 -1236 576 -1236 0 3
rlabel polysilicon 583 -1230 583 -1230 0 1
rlabel polysilicon 583 -1236 583 -1236 0 3
rlabel polysilicon 593 -1230 593 -1230 0 2
rlabel polysilicon 590 -1236 590 -1236 0 3
rlabel polysilicon 597 -1230 597 -1230 0 1
rlabel polysilicon 597 -1236 597 -1236 0 3
rlabel polysilicon 604 -1230 604 -1230 0 1
rlabel polysilicon 604 -1236 604 -1236 0 3
rlabel polysilicon 611 -1230 611 -1230 0 1
rlabel polysilicon 611 -1236 611 -1236 0 3
rlabel polysilicon 618 -1230 618 -1230 0 1
rlabel polysilicon 618 -1236 618 -1236 0 3
rlabel polysilicon 625 -1230 625 -1230 0 1
rlabel polysilicon 625 -1236 625 -1236 0 3
rlabel polysilicon 632 -1230 632 -1230 0 1
rlabel polysilicon 632 -1236 632 -1236 0 3
rlabel polysilicon 639 -1236 639 -1236 0 3
rlabel polysilicon 642 -1236 642 -1236 0 4
rlabel polysilicon 646 -1230 646 -1230 0 1
rlabel polysilicon 646 -1236 646 -1236 0 3
rlabel polysilicon 653 -1230 653 -1230 0 1
rlabel polysilicon 656 -1230 656 -1230 0 2
rlabel polysilicon 656 -1236 656 -1236 0 4
rlabel polysilicon 660 -1236 660 -1236 0 3
rlabel polysilicon 663 -1236 663 -1236 0 4
rlabel polysilicon 667 -1230 667 -1230 0 1
rlabel polysilicon 667 -1236 667 -1236 0 3
rlabel polysilicon 674 -1230 674 -1230 0 1
rlabel polysilicon 674 -1236 674 -1236 0 3
rlabel polysilicon 681 -1230 681 -1230 0 1
rlabel polysilicon 681 -1236 681 -1236 0 3
rlabel polysilicon 688 -1230 688 -1230 0 1
rlabel polysilicon 688 -1236 688 -1236 0 3
rlabel polysilicon 695 -1230 695 -1230 0 1
rlabel polysilicon 695 -1236 695 -1236 0 3
rlabel polysilicon 702 -1230 702 -1230 0 1
rlabel polysilicon 702 -1236 702 -1236 0 3
rlabel polysilicon 709 -1230 709 -1230 0 1
rlabel polysilicon 709 -1236 709 -1236 0 3
rlabel polysilicon 716 -1230 716 -1230 0 1
rlabel polysilicon 716 -1236 716 -1236 0 3
rlabel polysilicon 723 -1230 723 -1230 0 1
rlabel polysilicon 726 -1230 726 -1230 0 2
rlabel polysilicon 723 -1236 723 -1236 0 3
rlabel polysilicon 726 -1236 726 -1236 0 4
rlabel polysilicon 730 -1230 730 -1230 0 1
rlabel polysilicon 730 -1236 730 -1236 0 3
rlabel polysilicon 737 -1230 737 -1230 0 1
rlabel polysilicon 737 -1236 737 -1236 0 3
rlabel polysilicon 744 -1230 744 -1230 0 1
rlabel polysilicon 744 -1236 744 -1236 0 3
rlabel polysilicon 751 -1230 751 -1230 0 1
rlabel polysilicon 751 -1236 751 -1236 0 3
rlabel polysilicon 758 -1230 758 -1230 0 1
rlabel polysilicon 758 -1236 758 -1236 0 3
rlabel polysilicon 765 -1230 765 -1230 0 1
rlabel polysilicon 765 -1236 765 -1236 0 3
rlabel polysilicon 772 -1230 772 -1230 0 1
rlabel polysilicon 775 -1236 775 -1236 0 4
rlabel polysilicon 779 -1230 779 -1230 0 1
rlabel polysilicon 779 -1236 779 -1236 0 3
rlabel polysilicon 786 -1230 786 -1230 0 1
rlabel polysilicon 786 -1236 786 -1236 0 3
rlabel polysilicon 793 -1230 793 -1230 0 1
rlabel polysilicon 793 -1236 793 -1236 0 3
rlabel polysilicon 800 -1230 800 -1230 0 1
rlabel polysilicon 800 -1236 800 -1236 0 3
rlabel polysilicon 807 -1230 807 -1230 0 1
rlabel polysilicon 807 -1236 807 -1236 0 3
rlabel polysilicon 814 -1230 814 -1230 0 1
rlabel polysilicon 814 -1236 814 -1236 0 3
rlabel polysilicon 821 -1230 821 -1230 0 1
rlabel polysilicon 821 -1236 821 -1236 0 3
rlabel polysilicon 828 -1230 828 -1230 0 1
rlabel polysilicon 831 -1230 831 -1230 0 2
rlabel polysilicon 828 -1236 828 -1236 0 3
rlabel polysilicon 835 -1230 835 -1230 0 1
rlabel polysilicon 835 -1236 835 -1236 0 3
rlabel polysilicon 842 -1230 842 -1230 0 1
rlabel polysilicon 842 -1236 842 -1236 0 3
rlabel polysilicon 849 -1230 849 -1230 0 1
rlabel polysilicon 849 -1236 849 -1236 0 3
rlabel polysilicon 856 -1230 856 -1230 0 1
rlabel polysilicon 856 -1236 856 -1236 0 3
rlabel polysilicon 863 -1230 863 -1230 0 1
rlabel polysilicon 863 -1236 863 -1236 0 3
rlabel polysilicon 870 -1230 870 -1230 0 1
rlabel polysilicon 870 -1236 870 -1236 0 3
rlabel polysilicon 877 -1230 877 -1230 0 1
rlabel polysilicon 877 -1236 877 -1236 0 3
rlabel polysilicon 884 -1230 884 -1230 0 1
rlabel polysilicon 884 -1236 884 -1236 0 3
rlabel polysilicon 891 -1230 891 -1230 0 1
rlabel polysilicon 891 -1236 891 -1236 0 3
rlabel polysilicon 898 -1230 898 -1230 0 1
rlabel polysilicon 898 -1236 898 -1236 0 3
rlabel polysilicon 905 -1230 905 -1230 0 1
rlabel polysilicon 905 -1236 905 -1236 0 3
rlabel polysilicon 912 -1230 912 -1230 0 1
rlabel polysilicon 912 -1236 912 -1236 0 3
rlabel polysilicon 919 -1230 919 -1230 0 1
rlabel polysilicon 919 -1236 919 -1236 0 3
rlabel polysilicon 926 -1230 926 -1230 0 1
rlabel polysilicon 926 -1236 926 -1236 0 3
rlabel polysilicon 933 -1230 933 -1230 0 1
rlabel polysilicon 933 -1236 933 -1236 0 3
rlabel polysilicon 940 -1230 940 -1230 0 1
rlabel polysilicon 940 -1236 940 -1236 0 3
rlabel polysilicon 947 -1230 947 -1230 0 1
rlabel polysilicon 947 -1236 947 -1236 0 3
rlabel polysilicon 954 -1230 954 -1230 0 1
rlabel polysilicon 954 -1236 954 -1236 0 3
rlabel polysilicon 961 -1230 961 -1230 0 1
rlabel polysilicon 961 -1236 961 -1236 0 3
rlabel polysilicon 968 -1230 968 -1230 0 1
rlabel polysilicon 968 -1236 968 -1236 0 3
rlabel polysilicon 975 -1230 975 -1230 0 1
rlabel polysilicon 975 -1236 975 -1236 0 3
rlabel polysilicon 982 -1230 982 -1230 0 1
rlabel polysilicon 982 -1236 982 -1236 0 3
rlabel polysilicon 989 -1230 989 -1230 0 1
rlabel polysilicon 989 -1236 989 -1236 0 3
rlabel polysilicon 996 -1230 996 -1230 0 1
rlabel polysilicon 996 -1236 996 -1236 0 3
rlabel polysilicon 1003 -1230 1003 -1230 0 1
rlabel polysilicon 1003 -1236 1003 -1236 0 3
rlabel polysilicon 1010 -1230 1010 -1230 0 1
rlabel polysilicon 1010 -1236 1010 -1236 0 3
rlabel polysilicon 1017 -1230 1017 -1230 0 1
rlabel polysilicon 1017 -1236 1017 -1236 0 3
rlabel polysilicon 1024 -1230 1024 -1230 0 1
rlabel polysilicon 1024 -1236 1024 -1236 0 3
rlabel polysilicon 1031 -1230 1031 -1230 0 1
rlabel polysilicon 1031 -1236 1031 -1236 0 3
rlabel polysilicon 1038 -1230 1038 -1230 0 1
rlabel polysilicon 1038 -1236 1038 -1236 0 3
rlabel polysilicon 1045 -1230 1045 -1230 0 1
rlabel polysilicon 1045 -1236 1045 -1236 0 3
rlabel polysilicon 1052 -1230 1052 -1230 0 1
rlabel polysilicon 1052 -1236 1052 -1236 0 3
rlabel polysilicon 1059 -1230 1059 -1230 0 1
rlabel polysilicon 1059 -1236 1059 -1236 0 3
rlabel polysilicon 1066 -1230 1066 -1230 0 1
rlabel polysilicon 1066 -1236 1066 -1236 0 3
rlabel polysilicon 1073 -1230 1073 -1230 0 1
rlabel polysilicon 1073 -1236 1073 -1236 0 3
rlabel polysilicon 1080 -1230 1080 -1230 0 1
rlabel polysilicon 1080 -1236 1080 -1236 0 3
rlabel polysilicon 1087 -1230 1087 -1230 0 1
rlabel polysilicon 1087 -1236 1087 -1236 0 3
rlabel polysilicon 1094 -1230 1094 -1230 0 1
rlabel polysilicon 1094 -1236 1094 -1236 0 3
rlabel polysilicon 1101 -1230 1101 -1230 0 1
rlabel polysilicon 1101 -1236 1101 -1236 0 3
rlabel polysilicon 1108 -1230 1108 -1230 0 1
rlabel polysilicon 1108 -1236 1108 -1236 0 3
rlabel polysilicon 1115 -1230 1115 -1230 0 1
rlabel polysilicon 1115 -1236 1115 -1236 0 3
rlabel polysilicon 1122 -1230 1122 -1230 0 1
rlabel polysilicon 1122 -1236 1122 -1236 0 3
rlabel polysilicon 1129 -1230 1129 -1230 0 1
rlabel polysilicon 1129 -1236 1129 -1236 0 3
rlabel polysilicon 44 -1301 44 -1301 0 1
rlabel polysilicon 44 -1307 44 -1307 0 3
rlabel polysilicon 72 -1301 72 -1301 0 1
rlabel polysilicon 72 -1307 72 -1307 0 3
rlabel polysilicon 79 -1301 79 -1301 0 1
rlabel polysilicon 79 -1307 79 -1307 0 3
rlabel polysilicon 86 -1301 86 -1301 0 1
rlabel polysilicon 86 -1307 86 -1307 0 3
rlabel polysilicon 96 -1301 96 -1301 0 2
rlabel polysilicon 93 -1307 93 -1307 0 3
rlabel polysilicon 100 -1301 100 -1301 0 1
rlabel polysilicon 100 -1307 100 -1307 0 3
rlabel polysilicon 107 -1301 107 -1301 0 1
rlabel polysilicon 107 -1307 107 -1307 0 3
rlabel polysilicon 114 -1301 114 -1301 0 1
rlabel polysilicon 114 -1307 114 -1307 0 3
rlabel polysilicon 121 -1301 121 -1301 0 1
rlabel polysilicon 121 -1307 121 -1307 0 3
rlabel polysilicon 128 -1301 128 -1301 0 1
rlabel polysilicon 128 -1307 128 -1307 0 3
rlabel polysilicon 135 -1301 135 -1301 0 1
rlabel polysilicon 135 -1307 135 -1307 0 3
rlabel polysilicon 142 -1301 142 -1301 0 1
rlabel polysilicon 142 -1307 142 -1307 0 3
rlabel polysilicon 149 -1301 149 -1301 0 1
rlabel polysilicon 149 -1307 149 -1307 0 3
rlabel polysilicon 156 -1301 156 -1301 0 1
rlabel polysilicon 156 -1307 156 -1307 0 3
rlabel polysilicon 163 -1301 163 -1301 0 1
rlabel polysilicon 163 -1307 163 -1307 0 3
rlabel polysilicon 170 -1301 170 -1301 0 1
rlabel polysilicon 170 -1307 170 -1307 0 3
rlabel polysilicon 177 -1301 177 -1301 0 1
rlabel polysilicon 177 -1307 177 -1307 0 3
rlabel polysilicon 184 -1301 184 -1301 0 1
rlabel polysilicon 184 -1307 184 -1307 0 3
rlabel polysilicon 194 -1307 194 -1307 0 4
rlabel polysilicon 198 -1301 198 -1301 0 1
rlabel polysilicon 198 -1307 198 -1307 0 3
rlabel polysilicon 205 -1301 205 -1301 0 1
rlabel polysilicon 205 -1307 205 -1307 0 3
rlabel polysilicon 212 -1301 212 -1301 0 1
rlabel polysilicon 212 -1307 212 -1307 0 3
rlabel polysilicon 219 -1301 219 -1301 0 1
rlabel polysilicon 219 -1307 219 -1307 0 3
rlabel polysilicon 226 -1301 226 -1301 0 1
rlabel polysilicon 226 -1307 226 -1307 0 3
rlabel polysilicon 233 -1301 233 -1301 0 1
rlabel polysilicon 233 -1307 233 -1307 0 3
rlabel polysilicon 240 -1301 240 -1301 0 1
rlabel polysilicon 240 -1307 240 -1307 0 3
rlabel polysilicon 247 -1301 247 -1301 0 1
rlabel polysilicon 247 -1307 247 -1307 0 3
rlabel polysilicon 254 -1301 254 -1301 0 1
rlabel polysilicon 254 -1307 254 -1307 0 3
rlabel polysilicon 261 -1301 261 -1301 0 1
rlabel polysilicon 261 -1307 261 -1307 0 3
rlabel polysilicon 268 -1301 268 -1301 0 1
rlabel polysilicon 268 -1307 268 -1307 0 3
rlabel polysilicon 275 -1301 275 -1301 0 1
rlabel polysilicon 275 -1307 275 -1307 0 3
rlabel polysilicon 282 -1301 282 -1301 0 1
rlabel polysilicon 282 -1307 282 -1307 0 3
rlabel polysilicon 289 -1301 289 -1301 0 1
rlabel polysilicon 289 -1307 289 -1307 0 3
rlabel polysilicon 296 -1301 296 -1301 0 1
rlabel polysilicon 296 -1307 296 -1307 0 3
rlabel polysilicon 303 -1301 303 -1301 0 1
rlabel polysilicon 303 -1307 303 -1307 0 3
rlabel polysilicon 306 -1307 306 -1307 0 4
rlabel polysilicon 310 -1301 310 -1301 0 1
rlabel polysilicon 310 -1307 310 -1307 0 3
rlabel polysilicon 317 -1301 317 -1301 0 1
rlabel polysilicon 317 -1307 317 -1307 0 3
rlabel polysilicon 324 -1301 324 -1301 0 1
rlabel polysilicon 324 -1307 324 -1307 0 3
rlabel polysilicon 331 -1301 331 -1301 0 1
rlabel polysilicon 331 -1307 331 -1307 0 3
rlabel polysilicon 338 -1301 338 -1301 0 1
rlabel polysilicon 341 -1301 341 -1301 0 2
rlabel polysilicon 341 -1307 341 -1307 0 4
rlabel polysilicon 345 -1301 345 -1301 0 1
rlabel polysilicon 345 -1307 345 -1307 0 3
rlabel polysilicon 352 -1301 352 -1301 0 1
rlabel polysilicon 352 -1307 352 -1307 0 3
rlabel polysilicon 359 -1301 359 -1301 0 1
rlabel polysilicon 359 -1307 359 -1307 0 3
rlabel polysilicon 366 -1301 366 -1301 0 1
rlabel polysilicon 366 -1307 366 -1307 0 3
rlabel polysilicon 373 -1301 373 -1301 0 1
rlabel polysilicon 373 -1307 373 -1307 0 3
rlabel polysilicon 380 -1301 380 -1301 0 1
rlabel polysilicon 380 -1307 380 -1307 0 3
rlabel polysilicon 387 -1301 387 -1301 0 1
rlabel polysilicon 387 -1307 387 -1307 0 3
rlabel polysilicon 394 -1301 394 -1301 0 1
rlabel polysilicon 394 -1307 394 -1307 0 3
rlabel polysilicon 401 -1301 401 -1301 0 1
rlabel polysilicon 404 -1301 404 -1301 0 2
rlabel polysilicon 404 -1307 404 -1307 0 4
rlabel polysilicon 408 -1301 408 -1301 0 1
rlabel polysilicon 408 -1307 408 -1307 0 3
rlabel polysilicon 415 -1301 415 -1301 0 1
rlabel polysilicon 415 -1307 415 -1307 0 3
rlabel polysilicon 422 -1301 422 -1301 0 1
rlabel polysilicon 422 -1307 422 -1307 0 3
rlabel polysilicon 429 -1301 429 -1301 0 1
rlabel polysilicon 429 -1307 429 -1307 0 3
rlabel polysilicon 436 -1301 436 -1301 0 1
rlabel polysilicon 436 -1307 436 -1307 0 3
rlabel polysilicon 443 -1301 443 -1301 0 1
rlabel polysilicon 443 -1307 443 -1307 0 3
rlabel polysilicon 450 -1301 450 -1301 0 1
rlabel polysilicon 450 -1307 450 -1307 0 3
rlabel polysilicon 457 -1301 457 -1301 0 1
rlabel polysilicon 457 -1307 457 -1307 0 3
rlabel polysilicon 464 -1301 464 -1301 0 1
rlabel polysilicon 467 -1301 467 -1301 0 2
rlabel polysilicon 464 -1307 464 -1307 0 3
rlabel polysilicon 467 -1307 467 -1307 0 4
rlabel polysilicon 471 -1301 471 -1301 0 1
rlabel polysilicon 471 -1307 471 -1307 0 3
rlabel polysilicon 478 -1301 478 -1301 0 1
rlabel polysilicon 481 -1301 481 -1301 0 2
rlabel polysilicon 478 -1307 478 -1307 0 3
rlabel polysilicon 481 -1307 481 -1307 0 4
rlabel polysilicon 485 -1301 485 -1301 0 1
rlabel polysilicon 485 -1307 485 -1307 0 3
rlabel polysilicon 492 -1301 492 -1301 0 1
rlabel polysilicon 492 -1307 492 -1307 0 3
rlabel polysilicon 499 -1301 499 -1301 0 1
rlabel polysilicon 502 -1301 502 -1301 0 2
rlabel polysilicon 506 -1301 506 -1301 0 1
rlabel polysilicon 506 -1307 506 -1307 0 3
rlabel polysilicon 513 -1301 513 -1301 0 1
rlabel polysilicon 513 -1307 513 -1307 0 3
rlabel polysilicon 520 -1301 520 -1301 0 1
rlabel polysilicon 520 -1307 520 -1307 0 3
rlabel polysilicon 527 -1301 527 -1301 0 1
rlabel polysilicon 527 -1307 527 -1307 0 3
rlabel polysilicon 534 -1307 534 -1307 0 3
rlabel polysilicon 537 -1307 537 -1307 0 4
rlabel polysilicon 541 -1301 541 -1301 0 1
rlabel polysilicon 541 -1307 541 -1307 0 3
rlabel polysilicon 548 -1301 548 -1301 0 1
rlabel polysilicon 548 -1307 548 -1307 0 3
rlabel polysilicon 555 -1301 555 -1301 0 1
rlabel polysilicon 555 -1307 555 -1307 0 3
rlabel polysilicon 562 -1301 562 -1301 0 1
rlabel polysilicon 562 -1307 562 -1307 0 3
rlabel polysilicon 572 -1301 572 -1301 0 2
rlabel polysilicon 569 -1307 569 -1307 0 3
rlabel polysilicon 572 -1307 572 -1307 0 4
rlabel polysilicon 579 -1301 579 -1301 0 2
rlabel polysilicon 576 -1307 576 -1307 0 3
rlabel polysilicon 583 -1301 583 -1301 0 1
rlabel polysilicon 583 -1307 583 -1307 0 3
rlabel polysilicon 590 -1301 590 -1301 0 1
rlabel polysilicon 590 -1307 590 -1307 0 3
rlabel polysilicon 597 -1307 597 -1307 0 3
rlabel polysilicon 600 -1307 600 -1307 0 4
rlabel polysilicon 604 -1301 604 -1301 0 1
rlabel polysilicon 604 -1307 604 -1307 0 3
rlabel polysilicon 611 -1301 611 -1301 0 1
rlabel polysilicon 614 -1307 614 -1307 0 4
rlabel polysilicon 618 -1301 618 -1301 0 1
rlabel polysilicon 618 -1307 618 -1307 0 3
rlabel polysilicon 625 -1301 625 -1301 0 1
rlabel polysilicon 625 -1307 625 -1307 0 3
rlabel polysilicon 635 -1307 635 -1307 0 4
rlabel polysilicon 639 -1301 639 -1301 0 1
rlabel polysilicon 639 -1307 639 -1307 0 3
rlabel polysilicon 646 -1301 646 -1301 0 1
rlabel polysilicon 646 -1307 646 -1307 0 3
rlabel polysilicon 656 -1301 656 -1301 0 2
rlabel polysilicon 660 -1301 660 -1301 0 1
rlabel polysilicon 660 -1307 660 -1307 0 3
rlabel polysilicon 667 -1301 667 -1301 0 1
rlabel polysilicon 667 -1307 667 -1307 0 3
rlabel polysilicon 674 -1301 674 -1301 0 1
rlabel polysilicon 677 -1301 677 -1301 0 2
rlabel polysilicon 674 -1307 674 -1307 0 3
rlabel polysilicon 677 -1307 677 -1307 0 4
rlabel polysilicon 681 -1301 681 -1301 0 1
rlabel polysilicon 681 -1307 681 -1307 0 3
rlabel polysilicon 688 -1301 688 -1301 0 1
rlabel polysilicon 688 -1307 688 -1307 0 3
rlabel polysilicon 695 -1301 695 -1301 0 1
rlabel polysilicon 695 -1307 695 -1307 0 3
rlabel polysilicon 702 -1301 702 -1301 0 1
rlabel polysilicon 702 -1307 702 -1307 0 3
rlabel polysilicon 709 -1301 709 -1301 0 1
rlabel polysilicon 709 -1307 709 -1307 0 3
rlabel polysilicon 716 -1301 716 -1301 0 1
rlabel polysilicon 716 -1307 716 -1307 0 3
rlabel polysilicon 723 -1301 723 -1301 0 1
rlabel polysilicon 723 -1307 723 -1307 0 3
rlabel polysilicon 730 -1301 730 -1301 0 1
rlabel polysilicon 730 -1307 730 -1307 0 3
rlabel polysilicon 737 -1301 737 -1301 0 1
rlabel polysilicon 737 -1307 737 -1307 0 3
rlabel polysilicon 744 -1301 744 -1301 0 1
rlabel polysilicon 744 -1307 744 -1307 0 3
rlabel polysilicon 751 -1301 751 -1301 0 1
rlabel polysilicon 751 -1307 751 -1307 0 3
rlabel polysilicon 758 -1301 758 -1301 0 1
rlabel polysilicon 758 -1307 758 -1307 0 3
rlabel polysilicon 765 -1301 765 -1301 0 1
rlabel polysilicon 765 -1307 765 -1307 0 3
rlabel polysilicon 772 -1301 772 -1301 0 1
rlabel polysilicon 772 -1307 772 -1307 0 3
rlabel polysilicon 779 -1301 779 -1301 0 1
rlabel polysilicon 779 -1307 779 -1307 0 3
rlabel polysilicon 786 -1301 786 -1301 0 1
rlabel polysilicon 786 -1307 786 -1307 0 3
rlabel polysilicon 793 -1301 793 -1301 0 1
rlabel polysilicon 796 -1301 796 -1301 0 2
rlabel polysilicon 793 -1307 793 -1307 0 3
rlabel polysilicon 796 -1307 796 -1307 0 4
rlabel polysilicon 800 -1301 800 -1301 0 1
rlabel polysilicon 800 -1307 800 -1307 0 3
rlabel polysilicon 807 -1301 807 -1301 0 1
rlabel polysilicon 807 -1307 807 -1307 0 3
rlabel polysilicon 814 -1301 814 -1301 0 1
rlabel polysilicon 814 -1307 814 -1307 0 3
rlabel polysilicon 821 -1301 821 -1301 0 1
rlabel polysilicon 821 -1307 821 -1307 0 3
rlabel polysilicon 828 -1301 828 -1301 0 1
rlabel polysilicon 828 -1307 828 -1307 0 3
rlabel polysilicon 835 -1301 835 -1301 0 1
rlabel polysilicon 835 -1307 835 -1307 0 3
rlabel polysilicon 842 -1301 842 -1301 0 1
rlabel polysilicon 842 -1307 842 -1307 0 3
rlabel polysilicon 849 -1301 849 -1301 0 1
rlabel polysilicon 849 -1307 849 -1307 0 3
rlabel polysilicon 856 -1301 856 -1301 0 1
rlabel polysilicon 856 -1307 856 -1307 0 3
rlabel polysilicon 866 -1301 866 -1301 0 2
rlabel polysilicon 863 -1307 863 -1307 0 3
rlabel polysilicon 870 -1301 870 -1301 0 1
rlabel polysilicon 870 -1307 870 -1307 0 3
rlabel polysilicon 877 -1301 877 -1301 0 1
rlabel polysilicon 877 -1307 877 -1307 0 3
rlabel polysilicon 884 -1301 884 -1301 0 1
rlabel polysilicon 884 -1307 884 -1307 0 3
rlabel polysilicon 891 -1301 891 -1301 0 1
rlabel polysilicon 891 -1307 891 -1307 0 3
rlabel polysilicon 898 -1301 898 -1301 0 1
rlabel polysilicon 898 -1307 898 -1307 0 3
rlabel polysilicon 905 -1301 905 -1301 0 1
rlabel polysilicon 905 -1307 905 -1307 0 3
rlabel polysilicon 912 -1301 912 -1301 0 1
rlabel polysilicon 912 -1307 912 -1307 0 3
rlabel polysilicon 922 -1307 922 -1307 0 4
rlabel polysilicon 926 -1301 926 -1301 0 1
rlabel polysilicon 926 -1307 926 -1307 0 3
rlabel polysilicon 933 -1301 933 -1301 0 1
rlabel polysilicon 933 -1307 933 -1307 0 3
rlabel polysilicon 940 -1301 940 -1301 0 1
rlabel polysilicon 940 -1307 940 -1307 0 3
rlabel polysilicon 947 -1301 947 -1301 0 1
rlabel polysilicon 947 -1307 947 -1307 0 3
rlabel polysilicon 954 -1301 954 -1301 0 1
rlabel polysilicon 954 -1307 954 -1307 0 3
rlabel polysilicon 961 -1301 961 -1301 0 1
rlabel polysilicon 961 -1307 961 -1307 0 3
rlabel polysilicon 968 -1301 968 -1301 0 1
rlabel polysilicon 968 -1307 968 -1307 0 3
rlabel polysilicon 978 -1301 978 -1301 0 2
rlabel polysilicon 975 -1307 975 -1307 0 3
rlabel polysilicon 982 -1301 982 -1301 0 1
rlabel polysilicon 982 -1307 982 -1307 0 3
rlabel polysilicon 989 -1301 989 -1301 0 1
rlabel polysilicon 989 -1307 989 -1307 0 3
rlabel polysilicon 999 -1301 999 -1301 0 2
rlabel polysilicon 1003 -1301 1003 -1301 0 1
rlabel polysilicon 1003 -1307 1003 -1307 0 3
rlabel polysilicon 1010 -1301 1010 -1301 0 1
rlabel polysilicon 1010 -1307 1010 -1307 0 3
rlabel polysilicon 1017 -1301 1017 -1301 0 1
rlabel polysilicon 1017 -1307 1017 -1307 0 3
rlabel polysilicon 1020 -1307 1020 -1307 0 4
rlabel polysilicon 1024 -1301 1024 -1301 0 1
rlabel polysilicon 1027 -1301 1027 -1301 0 2
rlabel polysilicon 1031 -1301 1031 -1301 0 1
rlabel polysilicon 1031 -1307 1031 -1307 0 3
rlabel polysilicon 1038 -1301 1038 -1301 0 1
rlabel polysilicon 1038 -1307 1038 -1307 0 3
rlabel polysilicon 1045 -1301 1045 -1301 0 1
rlabel polysilicon 1045 -1307 1045 -1307 0 3
rlabel polysilicon 1052 -1301 1052 -1301 0 1
rlabel polysilicon 1052 -1307 1052 -1307 0 3
rlabel polysilicon 1059 -1301 1059 -1301 0 1
rlabel polysilicon 1062 -1301 1062 -1301 0 2
rlabel polysilicon 1059 -1307 1059 -1307 0 3
rlabel polysilicon 1066 -1301 1066 -1301 0 1
rlabel polysilicon 1066 -1307 1066 -1307 0 3
rlabel polysilicon 1080 -1301 1080 -1301 0 1
rlabel polysilicon 1080 -1307 1080 -1307 0 3
rlabel polysilicon 1087 -1301 1087 -1301 0 1
rlabel polysilicon 1087 -1307 1087 -1307 0 3
rlabel polysilicon 1097 -1301 1097 -1301 0 2
rlabel polysilicon 1097 -1307 1097 -1307 0 4
rlabel polysilicon 1101 -1301 1101 -1301 0 1
rlabel polysilicon 1101 -1307 1101 -1307 0 3
rlabel polysilicon 2 -1378 2 -1378 0 3
rlabel polysilicon 9 -1372 9 -1372 0 1
rlabel polysilicon 16 -1372 16 -1372 0 1
rlabel polysilicon 16 -1378 16 -1378 0 3
rlabel polysilicon 23 -1372 23 -1372 0 1
rlabel polysilicon 23 -1378 23 -1378 0 3
rlabel polysilicon 30 -1372 30 -1372 0 1
rlabel polysilicon 30 -1378 30 -1378 0 3
rlabel polysilicon 37 -1372 37 -1372 0 1
rlabel polysilicon 37 -1378 37 -1378 0 3
rlabel polysilicon 44 -1372 44 -1372 0 1
rlabel polysilicon 44 -1378 44 -1378 0 3
rlabel polysilicon 51 -1372 51 -1372 0 1
rlabel polysilicon 51 -1378 51 -1378 0 3
rlabel polysilicon 58 -1372 58 -1372 0 1
rlabel polysilicon 58 -1378 58 -1378 0 3
rlabel polysilicon 65 -1372 65 -1372 0 1
rlabel polysilicon 68 -1372 68 -1372 0 2
rlabel polysilicon 72 -1372 72 -1372 0 1
rlabel polysilicon 72 -1378 72 -1378 0 3
rlabel polysilicon 79 -1372 79 -1372 0 1
rlabel polysilicon 79 -1378 79 -1378 0 3
rlabel polysilicon 86 -1372 86 -1372 0 1
rlabel polysilicon 86 -1378 86 -1378 0 3
rlabel polysilicon 93 -1372 93 -1372 0 1
rlabel polysilicon 93 -1378 93 -1378 0 3
rlabel polysilicon 100 -1372 100 -1372 0 1
rlabel polysilicon 107 -1372 107 -1372 0 1
rlabel polysilicon 107 -1378 107 -1378 0 3
rlabel polysilicon 114 -1372 114 -1372 0 1
rlabel polysilicon 114 -1378 114 -1378 0 3
rlabel polysilicon 121 -1372 121 -1372 0 1
rlabel polysilicon 121 -1378 121 -1378 0 3
rlabel polysilicon 128 -1372 128 -1372 0 1
rlabel polysilicon 128 -1378 128 -1378 0 3
rlabel polysilicon 135 -1372 135 -1372 0 1
rlabel polysilicon 138 -1378 138 -1378 0 4
rlabel polysilicon 142 -1372 142 -1372 0 1
rlabel polysilicon 142 -1378 142 -1378 0 3
rlabel polysilicon 149 -1372 149 -1372 0 1
rlabel polysilicon 149 -1378 149 -1378 0 3
rlabel polysilicon 156 -1372 156 -1372 0 1
rlabel polysilicon 156 -1378 156 -1378 0 3
rlabel polysilicon 163 -1372 163 -1372 0 1
rlabel polysilicon 163 -1378 163 -1378 0 3
rlabel polysilicon 170 -1372 170 -1372 0 1
rlabel polysilicon 170 -1378 170 -1378 0 3
rlabel polysilicon 177 -1372 177 -1372 0 1
rlabel polysilicon 180 -1372 180 -1372 0 2
rlabel polysilicon 184 -1372 184 -1372 0 1
rlabel polysilicon 184 -1378 184 -1378 0 3
rlabel polysilicon 191 -1372 191 -1372 0 1
rlabel polysilicon 191 -1378 191 -1378 0 3
rlabel polysilicon 198 -1372 198 -1372 0 1
rlabel polysilicon 201 -1372 201 -1372 0 2
rlabel polysilicon 201 -1378 201 -1378 0 4
rlabel polysilicon 205 -1372 205 -1372 0 1
rlabel polysilicon 205 -1378 205 -1378 0 3
rlabel polysilicon 212 -1372 212 -1372 0 1
rlabel polysilicon 212 -1378 212 -1378 0 3
rlabel polysilicon 219 -1372 219 -1372 0 1
rlabel polysilicon 219 -1378 219 -1378 0 3
rlabel polysilicon 226 -1372 226 -1372 0 1
rlabel polysilicon 226 -1378 226 -1378 0 3
rlabel polysilicon 233 -1372 233 -1372 0 1
rlabel polysilicon 233 -1378 233 -1378 0 3
rlabel polysilicon 240 -1372 240 -1372 0 1
rlabel polysilicon 240 -1378 240 -1378 0 3
rlabel polysilicon 247 -1378 247 -1378 0 3
rlabel polysilicon 250 -1378 250 -1378 0 4
rlabel polysilicon 254 -1372 254 -1372 0 1
rlabel polysilicon 254 -1378 254 -1378 0 3
rlabel polysilicon 261 -1372 261 -1372 0 1
rlabel polysilicon 261 -1378 261 -1378 0 3
rlabel polysilicon 268 -1372 268 -1372 0 1
rlabel polysilicon 268 -1378 268 -1378 0 3
rlabel polysilicon 275 -1372 275 -1372 0 1
rlabel polysilicon 278 -1372 278 -1372 0 2
rlabel polysilicon 275 -1378 275 -1378 0 3
rlabel polysilicon 285 -1372 285 -1372 0 2
rlabel polysilicon 285 -1378 285 -1378 0 4
rlabel polysilicon 289 -1372 289 -1372 0 1
rlabel polysilicon 289 -1378 289 -1378 0 3
rlabel polysilicon 296 -1372 296 -1372 0 1
rlabel polysilicon 296 -1378 296 -1378 0 3
rlabel polysilicon 303 -1372 303 -1372 0 1
rlabel polysilicon 303 -1378 303 -1378 0 3
rlabel polysilicon 310 -1372 310 -1372 0 1
rlabel polysilicon 310 -1378 310 -1378 0 3
rlabel polysilicon 317 -1372 317 -1372 0 1
rlabel polysilicon 317 -1378 317 -1378 0 3
rlabel polysilicon 324 -1372 324 -1372 0 1
rlabel polysilicon 324 -1378 324 -1378 0 3
rlabel polysilicon 331 -1372 331 -1372 0 1
rlabel polysilicon 331 -1378 331 -1378 0 3
rlabel polysilicon 338 -1372 338 -1372 0 1
rlabel polysilicon 338 -1378 338 -1378 0 3
rlabel polysilicon 345 -1372 345 -1372 0 1
rlabel polysilicon 348 -1372 348 -1372 0 2
rlabel polysilicon 345 -1378 345 -1378 0 3
rlabel polysilicon 348 -1378 348 -1378 0 4
rlabel polysilicon 352 -1372 352 -1372 0 1
rlabel polysilicon 352 -1378 352 -1378 0 3
rlabel polysilicon 359 -1372 359 -1372 0 1
rlabel polysilicon 359 -1378 359 -1378 0 3
rlabel polysilicon 366 -1372 366 -1372 0 1
rlabel polysilicon 369 -1372 369 -1372 0 2
rlabel polysilicon 366 -1378 366 -1378 0 3
rlabel polysilicon 369 -1378 369 -1378 0 4
rlabel polysilicon 373 -1372 373 -1372 0 1
rlabel polysilicon 373 -1378 373 -1378 0 3
rlabel polysilicon 380 -1372 380 -1372 0 1
rlabel polysilicon 380 -1378 380 -1378 0 3
rlabel polysilicon 387 -1372 387 -1372 0 1
rlabel polysilicon 387 -1378 387 -1378 0 3
rlabel polysilicon 394 -1372 394 -1372 0 1
rlabel polysilicon 394 -1378 394 -1378 0 3
rlabel polysilicon 401 -1372 401 -1372 0 1
rlabel polysilicon 401 -1378 401 -1378 0 3
rlabel polysilicon 408 -1372 408 -1372 0 1
rlabel polysilicon 411 -1372 411 -1372 0 2
rlabel polysilicon 408 -1378 408 -1378 0 3
rlabel polysilicon 415 -1372 415 -1372 0 1
rlabel polysilicon 415 -1378 415 -1378 0 3
rlabel polysilicon 422 -1372 422 -1372 0 1
rlabel polysilicon 422 -1378 422 -1378 0 3
rlabel polysilicon 429 -1372 429 -1372 0 1
rlabel polysilicon 429 -1378 429 -1378 0 3
rlabel polysilicon 436 -1372 436 -1372 0 1
rlabel polysilicon 439 -1372 439 -1372 0 2
rlabel polysilicon 436 -1378 436 -1378 0 3
rlabel polysilicon 443 -1372 443 -1372 0 1
rlabel polysilicon 443 -1378 443 -1378 0 3
rlabel polysilicon 450 -1372 450 -1372 0 1
rlabel polysilicon 450 -1378 450 -1378 0 3
rlabel polysilicon 457 -1372 457 -1372 0 1
rlabel polysilicon 457 -1378 457 -1378 0 3
rlabel polysilicon 464 -1372 464 -1372 0 1
rlabel polysilicon 464 -1378 464 -1378 0 3
rlabel polysilicon 471 -1372 471 -1372 0 1
rlabel polysilicon 471 -1378 471 -1378 0 3
rlabel polysilicon 478 -1372 478 -1372 0 1
rlabel polysilicon 481 -1372 481 -1372 0 2
rlabel polysilicon 485 -1372 485 -1372 0 1
rlabel polysilicon 485 -1378 485 -1378 0 3
rlabel polysilicon 492 -1378 492 -1378 0 3
rlabel polysilicon 495 -1378 495 -1378 0 4
rlabel polysilicon 499 -1372 499 -1372 0 1
rlabel polysilicon 499 -1378 499 -1378 0 3
rlabel polysilicon 506 -1372 506 -1372 0 1
rlabel polysilicon 509 -1378 509 -1378 0 4
rlabel polysilicon 513 -1372 513 -1372 0 1
rlabel polysilicon 513 -1378 513 -1378 0 3
rlabel polysilicon 520 -1372 520 -1372 0 1
rlabel polysilicon 520 -1378 520 -1378 0 3
rlabel polysilicon 527 -1372 527 -1372 0 1
rlabel polysilicon 527 -1378 527 -1378 0 3
rlabel polysilicon 534 -1372 534 -1372 0 1
rlabel polysilicon 534 -1378 534 -1378 0 3
rlabel polysilicon 541 -1372 541 -1372 0 1
rlabel polysilicon 544 -1372 544 -1372 0 2
rlabel polysilicon 541 -1378 541 -1378 0 3
rlabel polysilicon 544 -1378 544 -1378 0 4
rlabel polysilicon 548 -1372 548 -1372 0 1
rlabel polysilicon 548 -1378 548 -1378 0 3
rlabel polysilicon 555 -1372 555 -1372 0 1
rlabel polysilicon 555 -1378 555 -1378 0 3
rlabel polysilicon 562 -1372 562 -1372 0 1
rlabel polysilicon 562 -1378 562 -1378 0 3
rlabel polysilicon 569 -1372 569 -1372 0 1
rlabel polysilicon 572 -1372 572 -1372 0 2
rlabel polysilicon 569 -1378 569 -1378 0 3
rlabel polysilicon 576 -1372 576 -1372 0 1
rlabel polysilicon 576 -1378 576 -1378 0 3
rlabel polysilicon 583 -1372 583 -1372 0 1
rlabel polysilicon 583 -1378 583 -1378 0 3
rlabel polysilicon 590 -1372 590 -1372 0 1
rlabel polysilicon 590 -1378 590 -1378 0 3
rlabel polysilicon 597 -1372 597 -1372 0 1
rlabel polysilicon 597 -1378 597 -1378 0 3
rlabel polysilicon 604 -1372 604 -1372 0 1
rlabel polysilicon 604 -1378 604 -1378 0 3
rlabel polysilicon 611 -1372 611 -1372 0 1
rlabel polysilicon 611 -1378 611 -1378 0 3
rlabel polysilicon 618 -1372 618 -1372 0 1
rlabel polysilicon 618 -1378 618 -1378 0 3
rlabel polysilicon 625 -1372 625 -1372 0 1
rlabel polysilicon 628 -1372 628 -1372 0 2
rlabel polysilicon 628 -1378 628 -1378 0 4
rlabel polysilicon 632 -1372 632 -1372 0 1
rlabel polysilicon 632 -1378 632 -1378 0 3
rlabel polysilicon 639 -1372 639 -1372 0 1
rlabel polysilicon 639 -1378 639 -1378 0 3
rlabel polysilicon 646 -1372 646 -1372 0 1
rlabel polysilicon 646 -1378 646 -1378 0 3
rlabel polysilicon 653 -1372 653 -1372 0 1
rlabel polysilicon 653 -1378 653 -1378 0 3
rlabel polysilicon 656 -1378 656 -1378 0 4
rlabel polysilicon 660 -1372 660 -1372 0 1
rlabel polysilicon 663 -1378 663 -1378 0 4
rlabel polysilicon 667 -1372 667 -1372 0 1
rlabel polysilicon 667 -1378 667 -1378 0 3
rlabel polysilicon 674 -1372 674 -1372 0 1
rlabel polysilicon 674 -1378 674 -1378 0 3
rlabel polysilicon 681 -1372 681 -1372 0 1
rlabel polysilicon 681 -1378 681 -1378 0 3
rlabel polysilicon 688 -1372 688 -1372 0 1
rlabel polysilicon 688 -1378 688 -1378 0 3
rlabel polysilicon 695 -1372 695 -1372 0 1
rlabel polysilicon 695 -1378 695 -1378 0 3
rlabel polysilicon 702 -1372 702 -1372 0 1
rlabel polysilicon 702 -1378 702 -1378 0 3
rlabel polysilicon 709 -1372 709 -1372 0 1
rlabel polysilicon 709 -1378 709 -1378 0 3
rlabel polysilicon 716 -1372 716 -1372 0 1
rlabel polysilicon 716 -1378 716 -1378 0 3
rlabel polysilicon 723 -1372 723 -1372 0 1
rlabel polysilicon 726 -1372 726 -1372 0 2
rlabel polysilicon 723 -1378 723 -1378 0 3
rlabel polysilicon 726 -1378 726 -1378 0 4
rlabel polysilicon 730 -1372 730 -1372 0 1
rlabel polysilicon 733 -1372 733 -1372 0 2
rlabel polysilicon 737 -1372 737 -1372 0 1
rlabel polysilicon 737 -1378 737 -1378 0 3
rlabel polysilicon 744 -1372 744 -1372 0 1
rlabel polysilicon 744 -1378 744 -1378 0 3
rlabel polysilicon 751 -1372 751 -1372 0 1
rlabel polysilicon 751 -1378 751 -1378 0 3
rlabel polysilicon 758 -1372 758 -1372 0 1
rlabel polysilicon 758 -1378 758 -1378 0 3
rlabel polysilicon 765 -1372 765 -1372 0 1
rlabel polysilicon 765 -1378 765 -1378 0 3
rlabel polysilicon 772 -1372 772 -1372 0 1
rlabel polysilicon 772 -1378 772 -1378 0 3
rlabel polysilicon 779 -1372 779 -1372 0 1
rlabel polysilicon 779 -1378 779 -1378 0 3
rlabel polysilicon 786 -1372 786 -1372 0 1
rlabel polysilicon 786 -1378 786 -1378 0 3
rlabel polysilicon 793 -1372 793 -1372 0 1
rlabel polysilicon 793 -1378 793 -1378 0 3
rlabel polysilicon 800 -1372 800 -1372 0 1
rlabel polysilicon 800 -1378 800 -1378 0 3
rlabel polysilicon 807 -1372 807 -1372 0 1
rlabel polysilicon 807 -1378 807 -1378 0 3
rlabel polysilicon 814 -1372 814 -1372 0 1
rlabel polysilicon 814 -1378 814 -1378 0 3
rlabel polysilicon 821 -1372 821 -1372 0 1
rlabel polysilicon 821 -1378 821 -1378 0 3
rlabel polysilicon 828 -1372 828 -1372 0 1
rlabel polysilicon 828 -1378 828 -1378 0 3
rlabel polysilicon 835 -1372 835 -1372 0 1
rlabel polysilicon 835 -1378 835 -1378 0 3
rlabel polysilicon 842 -1372 842 -1372 0 1
rlabel polysilicon 842 -1378 842 -1378 0 3
rlabel polysilicon 849 -1372 849 -1372 0 1
rlabel polysilicon 849 -1378 849 -1378 0 3
rlabel polysilicon 856 -1372 856 -1372 0 1
rlabel polysilicon 856 -1378 856 -1378 0 3
rlabel polysilicon 863 -1372 863 -1372 0 1
rlabel polysilicon 863 -1378 863 -1378 0 3
rlabel polysilicon 870 -1372 870 -1372 0 1
rlabel polysilicon 870 -1378 870 -1378 0 3
rlabel polysilicon 877 -1372 877 -1372 0 1
rlabel polysilicon 877 -1378 877 -1378 0 3
rlabel polysilicon 884 -1372 884 -1372 0 1
rlabel polysilicon 884 -1378 884 -1378 0 3
rlabel polysilicon 891 -1372 891 -1372 0 1
rlabel polysilicon 891 -1378 891 -1378 0 3
rlabel polysilicon 898 -1372 898 -1372 0 1
rlabel polysilicon 898 -1378 898 -1378 0 3
rlabel polysilicon 905 -1372 905 -1372 0 1
rlabel polysilicon 905 -1378 905 -1378 0 3
rlabel polysilicon 912 -1372 912 -1372 0 1
rlabel polysilicon 912 -1378 912 -1378 0 3
rlabel polysilicon 919 -1372 919 -1372 0 1
rlabel polysilicon 919 -1378 919 -1378 0 3
rlabel polysilicon 926 -1372 926 -1372 0 1
rlabel polysilicon 926 -1378 926 -1378 0 3
rlabel polysilicon 933 -1372 933 -1372 0 1
rlabel polysilicon 933 -1378 933 -1378 0 3
rlabel polysilicon 940 -1372 940 -1372 0 1
rlabel polysilicon 940 -1378 940 -1378 0 3
rlabel polysilicon 947 -1372 947 -1372 0 1
rlabel polysilicon 947 -1378 947 -1378 0 3
rlabel polysilicon 954 -1372 954 -1372 0 1
rlabel polysilicon 954 -1378 954 -1378 0 3
rlabel polysilicon 961 -1372 961 -1372 0 1
rlabel polysilicon 961 -1378 961 -1378 0 3
rlabel polysilicon 968 -1372 968 -1372 0 1
rlabel polysilicon 968 -1378 968 -1378 0 3
rlabel polysilicon 975 -1372 975 -1372 0 1
rlabel polysilicon 975 -1378 975 -1378 0 3
rlabel polysilicon 982 -1372 982 -1372 0 1
rlabel polysilicon 982 -1378 982 -1378 0 3
rlabel polysilicon 989 -1372 989 -1372 0 1
rlabel polysilicon 989 -1378 989 -1378 0 3
rlabel polysilicon 996 -1372 996 -1372 0 1
rlabel polysilicon 999 -1372 999 -1372 0 2
rlabel polysilicon 996 -1378 996 -1378 0 3
rlabel polysilicon 1003 -1372 1003 -1372 0 1
rlabel polysilicon 1003 -1378 1003 -1378 0 3
rlabel polysilicon 1010 -1372 1010 -1372 0 1
rlabel polysilicon 1010 -1378 1010 -1378 0 3
rlabel polysilicon 1017 -1372 1017 -1372 0 1
rlabel polysilicon 1017 -1378 1017 -1378 0 3
rlabel polysilicon 1024 -1372 1024 -1372 0 1
rlabel polysilicon 1031 -1372 1031 -1372 0 1
rlabel polysilicon 1031 -1378 1031 -1378 0 3
rlabel polysilicon 1066 -1372 1066 -1372 0 1
rlabel polysilicon 1066 -1378 1066 -1378 0 3
rlabel polysilicon 5 -1447 5 -1447 0 2
rlabel polysilicon 9 -1447 9 -1447 0 1
rlabel polysilicon 9 -1453 9 -1453 0 3
rlabel polysilicon 19 -1453 19 -1453 0 4
rlabel polysilicon 23 -1447 23 -1447 0 1
rlabel polysilicon 23 -1453 23 -1453 0 3
rlabel polysilicon 30 -1447 30 -1447 0 1
rlabel polysilicon 30 -1453 30 -1453 0 3
rlabel polysilicon 37 -1453 37 -1453 0 3
rlabel polysilicon 40 -1453 40 -1453 0 4
rlabel polysilicon 44 -1447 44 -1447 0 1
rlabel polysilicon 44 -1453 44 -1453 0 3
rlabel polysilicon 51 -1447 51 -1447 0 1
rlabel polysilicon 51 -1453 51 -1453 0 3
rlabel polysilicon 58 -1447 58 -1447 0 1
rlabel polysilicon 58 -1453 58 -1453 0 3
rlabel polysilicon 68 -1453 68 -1453 0 4
rlabel polysilicon 72 -1447 72 -1447 0 1
rlabel polysilicon 72 -1453 72 -1453 0 3
rlabel polysilicon 79 -1447 79 -1447 0 1
rlabel polysilicon 79 -1453 79 -1453 0 3
rlabel polysilicon 86 -1447 86 -1447 0 1
rlabel polysilicon 86 -1453 86 -1453 0 3
rlabel polysilicon 93 -1447 93 -1447 0 1
rlabel polysilicon 93 -1453 93 -1453 0 3
rlabel polysilicon 100 -1447 100 -1447 0 1
rlabel polysilicon 100 -1453 100 -1453 0 3
rlabel polysilicon 107 -1447 107 -1447 0 1
rlabel polysilicon 107 -1453 107 -1453 0 3
rlabel polysilicon 114 -1447 114 -1447 0 1
rlabel polysilicon 114 -1453 114 -1453 0 3
rlabel polysilicon 121 -1447 121 -1447 0 1
rlabel polysilicon 121 -1453 121 -1453 0 3
rlabel polysilicon 128 -1447 128 -1447 0 1
rlabel polysilicon 128 -1453 128 -1453 0 3
rlabel polysilicon 135 -1447 135 -1447 0 1
rlabel polysilicon 135 -1453 135 -1453 0 3
rlabel polysilicon 138 -1453 138 -1453 0 4
rlabel polysilicon 142 -1447 142 -1447 0 1
rlabel polysilicon 142 -1453 142 -1453 0 3
rlabel polysilicon 149 -1447 149 -1447 0 1
rlabel polysilicon 149 -1453 149 -1453 0 3
rlabel polysilicon 156 -1447 156 -1447 0 1
rlabel polysilicon 156 -1453 156 -1453 0 3
rlabel polysilicon 163 -1447 163 -1447 0 1
rlabel polysilicon 163 -1453 163 -1453 0 3
rlabel polysilicon 170 -1447 170 -1447 0 1
rlabel polysilicon 170 -1453 170 -1453 0 3
rlabel polysilicon 177 -1447 177 -1447 0 1
rlabel polysilicon 177 -1453 177 -1453 0 3
rlabel polysilicon 184 -1447 184 -1447 0 1
rlabel polysilicon 184 -1453 184 -1453 0 3
rlabel polysilicon 191 -1453 191 -1453 0 3
rlabel polysilicon 194 -1453 194 -1453 0 4
rlabel polysilicon 198 -1447 198 -1447 0 1
rlabel polysilicon 198 -1453 198 -1453 0 3
rlabel polysilicon 205 -1447 205 -1447 0 1
rlabel polysilicon 208 -1447 208 -1447 0 2
rlabel polysilicon 215 -1453 215 -1453 0 4
rlabel polysilicon 219 -1447 219 -1447 0 1
rlabel polysilicon 219 -1453 219 -1453 0 3
rlabel polysilicon 226 -1447 226 -1447 0 1
rlabel polysilicon 226 -1453 226 -1453 0 3
rlabel polysilicon 233 -1447 233 -1447 0 1
rlabel polysilicon 233 -1453 233 -1453 0 3
rlabel polysilicon 240 -1447 240 -1447 0 1
rlabel polysilicon 240 -1453 240 -1453 0 3
rlabel polysilicon 247 -1447 247 -1447 0 1
rlabel polysilicon 247 -1453 247 -1453 0 3
rlabel polysilicon 254 -1447 254 -1447 0 1
rlabel polysilicon 254 -1453 254 -1453 0 3
rlabel polysilicon 261 -1447 261 -1447 0 1
rlabel polysilicon 261 -1453 261 -1453 0 3
rlabel polysilicon 268 -1447 268 -1447 0 1
rlabel polysilicon 268 -1453 268 -1453 0 3
rlabel polysilicon 275 -1453 275 -1453 0 3
rlabel polysilicon 278 -1453 278 -1453 0 4
rlabel polysilicon 285 -1453 285 -1453 0 4
rlabel polysilicon 289 -1447 289 -1447 0 1
rlabel polysilicon 289 -1453 289 -1453 0 3
rlabel polysilicon 296 -1447 296 -1447 0 1
rlabel polysilicon 296 -1453 296 -1453 0 3
rlabel polysilicon 303 -1447 303 -1447 0 1
rlabel polysilicon 303 -1453 303 -1453 0 3
rlabel polysilicon 310 -1447 310 -1447 0 1
rlabel polysilicon 310 -1453 310 -1453 0 3
rlabel polysilicon 324 -1447 324 -1447 0 1
rlabel polysilicon 324 -1453 324 -1453 0 3
rlabel polysilicon 331 -1447 331 -1447 0 1
rlabel polysilicon 331 -1453 331 -1453 0 3
rlabel polysilicon 338 -1447 338 -1447 0 1
rlabel polysilicon 338 -1453 338 -1453 0 3
rlabel polysilicon 345 -1447 345 -1447 0 1
rlabel polysilicon 345 -1453 345 -1453 0 3
rlabel polysilicon 352 -1447 352 -1447 0 1
rlabel polysilicon 352 -1453 352 -1453 0 3
rlabel polysilicon 359 -1447 359 -1447 0 1
rlabel polysilicon 359 -1453 359 -1453 0 3
rlabel polysilicon 366 -1447 366 -1447 0 1
rlabel polysilicon 369 -1447 369 -1447 0 2
rlabel polysilicon 366 -1453 366 -1453 0 3
rlabel polysilicon 373 -1447 373 -1447 0 1
rlabel polysilicon 376 -1447 376 -1447 0 2
rlabel polysilicon 373 -1453 373 -1453 0 3
rlabel polysilicon 376 -1453 376 -1453 0 4
rlabel polysilicon 380 -1447 380 -1447 0 1
rlabel polysilicon 380 -1453 380 -1453 0 3
rlabel polysilicon 387 -1447 387 -1447 0 1
rlabel polysilicon 387 -1453 387 -1453 0 3
rlabel polysilicon 394 -1447 394 -1447 0 1
rlabel polysilicon 394 -1453 394 -1453 0 3
rlabel polysilicon 401 -1447 401 -1447 0 1
rlabel polysilicon 401 -1453 401 -1453 0 3
rlabel polysilicon 408 -1447 408 -1447 0 1
rlabel polysilicon 408 -1453 408 -1453 0 3
rlabel polysilicon 415 -1447 415 -1447 0 1
rlabel polysilicon 415 -1453 415 -1453 0 3
rlabel polysilicon 422 -1447 422 -1447 0 1
rlabel polysilicon 422 -1453 422 -1453 0 3
rlabel polysilicon 425 -1453 425 -1453 0 4
rlabel polysilicon 429 -1447 429 -1447 0 1
rlabel polysilicon 429 -1453 429 -1453 0 3
rlabel polysilicon 436 -1447 436 -1447 0 1
rlabel polysilicon 439 -1447 439 -1447 0 2
rlabel polysilicon 436 -1453 436 -1453 0 3
rlabel polysilicon 443 -1447 443 -1447 0 1
rlabel polysilicon 443 -1453 443 -1453 0 3
rlabel polysilicon 450 -1447 450 -1447 0 1
rlabel polysilicon 450 -1453 450 -1453 0 3
rlabel polysilicon 460 -1447 460 -1447 0 2
rlabel polysilicon 457 -1453 457 -1453 0 3
rlabel polysilicon 460 -1453 460 -1453 0 4
rlabel polysilicon 464 -1447 464 -1447 0 1
rlabel polysilicon 464 -1453 464 -1453 0 3
rlabel polysilicon 474 -1447 474 -1447 0 2
rlabel polysilicon 471 -1453 471 -1453 0 3
rlabel polysilicon 474 -1453 474 -1453 0 4
rlabel polysilicon 478 -1447 478 -1447 0 1
rlabel polysilicon 478 -1453 478 -1453 0 3
rlabel polysilicon 485 -1447 485 -1447 0 1
rlabel polysilicon 488 -1447 488 -1447 0 2
rlabel polysilicon 488 -1453 488 -1453 0 4
rlabel polysilicon 492 -1447 492 -1447 0 1
rlabel polysilicon 492 -1453 492 -1453 0 3
rlabel polysilicon 499 -1447 499 -1447 0 1
rlabel polysilicon 499 -1453 499 -1453 0 3
rlabel polysilicon 506 -1447 506 -1447 0 1
rlabel polysilicon 506 -1453 506 -1453 0 3
rlabel polysilicon 513 -1447 513 -1447 0 1
rlabel polysilicon 513 -1453 513 -1453 0 3
rlabel polysilicon 520 -1447 520 -1447 0 1
rlabel polysilicon 523 -1447 523 -1447 0 2
rlabel polysilicon 520 -1453 520 -1453 0 3
rlabel polysilicon 527 -1447 527 -1447 0 1
rlabel polysilicon 530 -1447 530 -1447 0 2
rlabel polysilicon 527 -1453 527 -1453 0 3
rlabel polysilicon 534 -1447 534 -1447 0 1
rlabel polysilicon 537 -1447 537 -1447 0 2
rlabel polysilicon 537 -1453 537 -1453 0 4
rlabel polysilicon 541 -1447 541 -1447 0 1
rlabel polysilicon 541 -1453 541 -1453 0 3
rlabel polysilicon 548 -1447 548 -1447 0 1
rlabel polysilicon 548 -1453 548 -1453 0 3
rlabel polysilicon 555 -1447 555 -1447 0 1
rlabel polysilicon 555 -1453 555 -1453 0 3
rlabel polysilicon 562 -1447 562 -1447 0 1
rlabel polysilicon 562 -1453 562 -1453 0 3
rlabel polysilicon 569 -1447 569 -1447 0 1
rlabel polysilicon 569 -1453 569 -1453 0 3
rlabel polysilicon 576 -1447 576 -1447 0 1
rlabel polysilicon 576 -1453 576 -1453 0 3
rlabel polysilicon 583 -1447 583 -1447 0 1
rlabel polysilicon 583 -1453 583 -1453 0 3
rlabel polysilicon 590 -1447 590 -1447 0 1
rlabel polysilicon 590 -1453 590 -1453 0 3
rlabel polysilicon 597 -1447 597 -1447 0 1
rlabel polysilicon 597 -1453 597 -1453 0 3
rlabel polysilicon 607 -1453 607 -1453 0 4
rlabel polysilicon 611 -1447 611 -1447 0 1
rlabel polysilicon 611 -1453 611 -1453 0 3
rlabel polysilicon 618 -1447 618 -1447 0 1
rlabel polysilicon 618 -1453 618 -1453 0 3
rlabel polysilicon 625 -1447 625 -1447 0 1
rlabel polysilicon 625 -1453 625 -1453 0 3
rlabel polysilicon 635 -1453 635 -1453 0 4
rlabel polysilicon 639 -1447 639 -1447 0 1
rlabel polysilicon 639 -1453 639 -1453 0 3
rlabel polysilicon 642 -1453 642 -1453 0 4
rlabel polysilicon 646 -1447 646 -1447 0 1
rlabel polysilicon 646 -1453 646 -1453 0 3
rlabel polysilicon 653 -1447 653 -1447 0 1
rlabel polysilicon 653 -1453 653 -1453 0 3
rlabel polysilicon 660 -1447 660 -1447 0 1
rlabel polysilicon 660 -1453 660 -1453 0 3
rlabel polysilicon 667 -1447 667 -1447 0 1
rlabel polysilicon 667 -1453 667 -1453 0 3
rlabel polysilicon 674 -1447 674 -1447 0 1
rlabel polysilicon 674 -1453 674 -1453 0 3
rlabel polysilicon 681 -1447 681 -1447 0 1
rlabel polysilicon 681 -1453 681 -1453 0 3
rlabel polysilicon 688 -1447 688 -1447 0 1
rlabel polysilicon 688 -1453 688 -1453 0 3
rlabel polysilicon 695 -1447 695 -1447 0 1
rlabel polysilicon 695 -1453 695 -1453 0 3
rlabel polysilicon 702 -1447 702 -1447 0 1
rlabel polysilicon 702 -1453 702 -1453 0 3
rlabel polysilicon 709 -1447 709 -1447 0 1
rlabel polysilicon 709 -1453 709 -1453 0 3
rlabel polysilicon 716 -1447 716 -1447 0 1
rlabel polysilicon 723 -1447 723 -1447 0 1
rlabel polysilicon 723 -1453 723 -1453 0 3
rlabel polysilicon 730 -1447 730 -1447 0 1
rlabel polysilicon 730 -1453 730 -1453 0 3
rlabel polysilicon 737 -1447 737 -1447 0 1
rlabel polysilicon 737 -1453 737 -1453 0 3
rlabel polysilicon 744 -1447 744 -1447 0 1
rlabel polysilicon 744 -1453 744 -1453 0 3
rlabel polysilicon 747 -1453 747 -1453 0 4
rlabel polysilicon 751 -1447 751 -1447 0 1
rlabel polysilicon 751 -1453 751 -1453 0 3
rlabel polysilicon 758 -1447 758 -1447 0 1
rlabel polysilicon 758 -1453 758 -1453 0 3
rlabel polysilicon 765 -1453 765 -1453 0 3
rlabel polysilicon 768 -1453 768 -1453 0 4
rlabel polysilicon 772 -1447 772 -1447 0 1
rlabel polysilicon 772 -1453 772 -1453 0 3
rlabel polysilicon 779 -1447 779 -1447 0 1
rlabel polysilicon 779 -1453 779 -1453 0 3
rlabel polysilicon 786 -1447 786 -1447 0 1
rlabel polysilicon 786 -1453 786 -1453 0 3
rlabel polysilicon 793 -1447 793 -1447 0 1
rlabel polysilicon 796 -1447 796 -1447 0 2
rlabel polysilicon 793 -1453 793 -1453 0 3
rlabel polysilicon 796 -1453 796 -1453 0 4
rlabel polysilicon 800 -1447 800 -1447 0 1
rlabel polysilicon 800 -1453 800 -1453 0 3
rlabel polysilicon 807 -1447 807 -1447 0 1
rlabel polysilicon 807 -1453 807 -1453 0 3
rlabel polysilicon 814 -1447 814 -1447 0 1
rlabel polysilicon 814 -1453 814 -1453 0 3
rlabel polysilicon 821 -1447 821 -1447 0 1
rlabel polysilicon 824 -1453 824 -1453 0 4
rlabel polysilicon 828 -1447 828 -1447 0 1
rlabel polysilicon 828 -1453 828 -1453 0 3
rlabel polysilicon 835 -1447 835 -1447 0 1
rlabel polysilicon 835 -1453 835 -1453 0 3
rlabel polysilicon 842 -1447 842 -1447 0 1
rlabel polysilicon 842 -1453 842 -1453 0 3
rlabel polysilicon 849 -1447 849 -1447 0 1
rlabel polysilicon 849 -1453 849 -1453 0 3
rlabel polysilicon 856 -1447 856 -1447 0 1
rlabel polysilicon 856 -1453 856 -1453 0 3
rlabel polysilicon 863 -1447 863 -1447 0 1
rlabel polysilicon 863 -1453 863 -1453 0 3
rlabel polysilicon 870 -1447 870 -1447 0 1
rlabel polysilicon 870 -1453 870 -1453 0 3
rlabel polysilicon 877 -1447 877 -1447 0 1
rlabel polysilicon 877 -1453 877 -1453 0 3
rlabel polysilicon 884 -1447 884 -1447 0 1
rlabel polysilicon 884 -1453 884 -1453 0 3
rlabel polysilicon 891 -1447 891 -1447 0 1
rlabel polysilicon 891 -1453 891 -1453 0 3
rlabel polysilicon 898 -1447 898 -1447 0 1
rlabel polysilicon 898 -1453 898 -1453 0 3
rlabel polysilicon 905 -1447 905 -1447 0 1
rlabel polysilicon 905 -1453 905 -1453 0 3
rlabel polysilicon 912 -1447 912 -1447 0 1
rlabel polysilicon 912 -1453 912 -1453 0 3
rlabel polysilicon 919 -1447 919 -1447 0 1
rlabel polysilicon 919 -1453 919 -1453 0 3
rlabel polysilicon 926 -1447 926 -1447 0 1
rlabel polysilicon 926 -1453 926 -1453 0 3
rlabel polysilicon 933 -1447 933 -1447 0 1
rlabel polysilicon 933 -1453 933 -1453 0 3
rlabel polysilicon 940 -1447 940 -1447 0 1
rlabel polysilicon 940 -1453 940 -1453 0 3
rlabel polysilicon 947 -1447 947 -1447 0 1
rlabel polysilicon 947 -1453 947 -1453 0 3
rlabel polysilicon 954 -1447 954 -1447 0 1
rlabel polysilicon 954 -1453 954 -1453 0 3
rlabel polysilicon 961 -1447 961 -1447 0 1
rlabel polysilicon 961 -1453 961 -1453 0 3
rlabel polysilicon 968 -1447 968 -1447 0 1
rlabel polysilicon 968 -1453 968 -1453 0 3
rlabel polysilicon 975 -1447 975 -1447 0 1
rlabel polysilicon 975 -1453 975 -1453 0 3
rlabel polysilicon 982 -1447 982 -1447 0 1
rlabel polysilicon 982 -1453 982 -1453 0 3
rlabel polysilicon 989 -1447 989 -1447 0 1
rlabel polysilicon 989 -1453 989 -1453 0 3
rlabel polysilicon 996 -1447 996 -1447 0 1
rlabel polysilicon 996 -1453 996 -1453 0 3
rlabel polysilicon 1003 -1447 1003 -1447 0 1
rlabel polysilicon 1003 -1453 1003 -1453 0 3
rlabel polysilicon 1010 -1447 1010 -1447 0 1
rlabel polysilicon 1010 -1453 1010 -1453 0 3
rlabel polysilicon 1017 -1447 1017 -1447 0 1
rlabel polysilicon 1017 -1453 1017 -1453 0 3
rlabel polysilicon 1024 -1447 1024 -1447 0 1
rlabel polysilicon 1024 -1453 1024 -1453 0 3
rlabel polysilicon 1031 -1447 1031 -1447 0 1
rlabel polysilicon 1031 -1453 1031 -1453 0 3
rlabel polysilicon 1038 -1447 1038 -1447 0 1
rlabel polysilicon 1038 -1453 1038 -1453 0 3
rlabel polysilicon 1045 -1447 1045 -1447 0 1
rlabel polysilicon 1048 -1447 1048 -1447 0 2
rlabel polysilicon 1048 -1453 1048 -1453 0 4
rlabel polysilicon 1052 -1447 1052 -1447 0 1
rlabel polysilicon 1055 -1447 1055 -1447 0 2
rlabel polysilicon 1059 -1447 1059 -1447 0 1
rlabel polysilicon 1059 -1453 1059 -1453 0 3
rlabel polysilicon 1066 -1447 1066 -1447 0 1
rlabel polysilicon 1066 -1453 1066 -1453 0 3
rlabel polysilicon 2 -1530 2 -1530 0 1
rlabel polysilicon 2 -1536 2 -1536 0 3
rlabel polysilicon 16 -1530 16 -1530 0 1
rlabel polysilicon 16 -1536 16 -1536 0 3
rlabel polysilicon 23 -1530 23 -1530 0 1
rlabel polysilicon 23 -1536 23 -1536 0 3
rlabel polysilicon 30 -1530 30 -1530 0 1
rlabel polysilicon 30 -1536 30 -1536 0 3
rlabel polysilicon 37 -1530 37 -1530 0 1
rlabel polysilicon 37 -1536 37 -1536 0 3
rlabel polysilicon 44 -1530 44 -1530 0 1
rlabel polysilicon 44 -1536 44 -1536 0 3
rlabel polysilicon 51 -1530 51 -1530 0 1
rlabel polysilicon 51 -1536 51 -1536 0 3
rlabel polysilicon 58 -1530 58 -1530 0 1
rlabel polysilicon 58 -1536 58 -1536 0 3
rlabel polysilicon 68 -1530 68 -1530 0 2
rlabel polysilicon 68 -1536 68 -1536 0 4
rlabel polysilicon 72 -1530 72 -1530 0 1
rlabel polysilicon 72 -1536 72 -1536 0 3
rlabel polysilicon 79 -1530 79 -1530 0 1
rlabel polysilicon 79 -1536 79 -1536 0 3
rlabel polysilicon 86 -1530 86 -1530 0 1
rlabel polysilicon 86 -1536 86 -1536 0 3
rlabel polysilicon 93 -1530 93 -1530 0 1
rlabel polysilicon 96 -1530 96 -1530 0 2
rlabel polysilicon 100 -1530 100 -1530 0 1
rlabel polysilicon 100 -1536 100 -1536 0 3
rlabel polysilicon 107 -1530 107 -1530 0 1
rlabel polysilicon 107 -1536 107 -1536 0 3
rlabel polysilicon 114 -1530 114 -1530 0 1
rlabel polysilicon 114 -1536 114 -1536 0 3
rlabel polysilicon 117 -1536 117 -1536 0 4
rlabel polysilicon 121 -1530 121 -1530 0 1
rlabel polysilicon 121 -1536 121 -1536 0 3
rlabel polysilicon 128 -1530 128 -1530 0 1
rlabel polysilicon 128 -1536 128 -1536 0 3
rlabel polysilicon 135 -1530 135 -1530 0 1
rlabel polysilicon 135 -1536 135 -1536 0 3
rlabel polysilicon 142 -1530 142 -1530 0 1
rlabel polysilicon 142 -1536 142 -1536 0 3
rlabel polysilicon 149 -1530 149 -1530 0 1
rlabel polysilicon 149 -1536 149 -1536 0 3
rlabel polysilicon 156 -1530 156 -1530 0 1
rlabel polysilicon 156 -1536 156 -1536 0 3
rlabel polysilicon 163 -1530 163 -1530 0 1
rlabel polysilicon 163 -1536 163 -1536 0 3
rlabel polysilicon 170 -1530 170 -1530 0 1
rlabel polysilicon 170 -1536 170 -1536 0 3
rlabel polysilicon 177 -1530 177 -1530 0 1
rlabel polysilicon 177 -1536 177 -1536 0 3
rlabel polysilicon 184 -1530 184 -1530 0 1
rlabel polysilicon 184 -1536 184 -1536 0 3
rlabel polysilicon 191 -1530 191 -1530 0 1
rlabel polysilicon 191 -1536 191 -1536 0 3
rlabel polysilicon 198 -1530 198 -1530 0 1
rlabel polysilicon 201 -1536 201 -1536 0 4
rlabel polysilicon 205 -1530 205 -1530 0 1
rlabel polysilicon 205 -1536 205 -1536 0 3
rlabel polysilicon 212 -1530 212 -1530 0 1
rlabel polysilicon 212 -1536 212 -1536 0 3
rlabel polysilicon 219 -1530 219 -1530 0 1
rlabel polysilicon 219 -1536 219 -1536 0 3
rlabel polysilicon 226 -1530 226 -1530 0 1
rlabel polysilicon 226 -1536 226 -1536 0 3
rlabel polysilicon 233 -1530 233 -1530 0 1
rlabel polysilicon 233 -1536 233 -1536 0 3
rlabel polysilicon 240 -1530 240 -1530 0 1
rlabel polysilicon 240 -1536 240 -1536 0 3
rlabel polysilicon 247 -1530 247 -1530 0 1
rlabel polysilicon 247 -1536 247 -1536 0 3
rlabel polysilicon 254 -1530 254 -1530 0 1
rlabel polysilicon 254 -1536 254 -1536 0 3
rlabel polysilicon 261 -1530 261 -1530 0 1
rlabel polysilicon 261 -1536 261 -1536 0 3
rlabel polysilicon 268 -1530 268 -1530 0 1
rlabel polysilicon 268 -1536 268 -1536 0 3
rlabel polysilicon 275 -1530 275 -1530 0 1
rlabel polysilicon 275 -1536 275 -1536 0 3
rlabel polysilicon 282 -1530 282 -1530 0 1
rlabel polysilicon 282 -1536 282 -1536 0 3
rlabel polysilicon 289 -1530 289 -1530 0 1
rlabel polysilicon 289 -1536 289 -1536 0 3
rlabel polysilicon 296 -1530 296 -1530 0 1
rlabel polysilicon 296 -1536 296 -1536 0 3
rlabel polysilicon 303 -1530 303 -1530 0 1
rlabel polysilicon 303 -1536 303 -1536 0 3
rlabel polysilicon 310 -1530 310 -1530 0 1
rlabel polysilicon 310 -1536 310 -1536 0 3
rlabel polysilicon 317 -1530 317 -1530 0 1
rlabel polysilicon 317 -1536 317 -1536 0 3
rlabel polysilicon 324 -1530 324 -1530 0 1
rlabel polysilicon 324 -1536 324 -1536 0 3
rlabel polysilicon 331 -1530 331 -1530 0 1
rlabel polysilicon 331 -1536 331 -1536 0 3
rlabel polysilicon 338 -1530 338 -1530 0 1
rlabel polysilicon 338 -1536 338 -1536 0 3
rlabel polysilicon 348 -1530 348 -1530 0 2
rlabel polysilicon 352 -1530 352 -1530 0 1
rlabel polysilicon 355 -1536 355 -1536 0 4
rlabel polysilicon 359 -1530 359 -1530 0 1
rlabel polysilicon 359 -1536 359 -1536 0 3
rlabel polysilicon 366 -1530 366 -1530 0 1
rlabel polysilicon 366 -1536 366 -1536 0 3
rlabel polysilicon 373 -1530 373 -1530 0 1
rlabel polysilicon 373 -1536 373 -1536 0 3
rlabel polysilicon 380 -1530 380 -1530 0 1
rlabel polysilicon 380 -1536 380 -1536 0 3
rlabel polysilicon 387 -1530 387 -1530 0 1
rlabel polysilicon 387 -1536 387 -1536 0 3
rlabel polysilicon 394 -1530 394 -1530 0 1
rlabel polysilicon 394 -1536 394 -1536 0 3
rlabel polysilicon 401 -1530 401 -1530 0 1
rlabel polysilicon 401 -1536 401 -1536 0 3
rlabel polysilicon 408 -1530 408 -1530 0 1
rlabel polysilicon 408 -1536 408 -1536 0 3
rlabel polysilicon 411 -1536 411 -1536 0 4
rlabel polysilicon 415 -1530 415 -1530 0 1
rlabel polysilicon 415 -1536 415 -1536 0 3
rlabel polysilicon 422 -1530 422 -1530 0 1
rlabel polysilicon 422 -1536 422 -1536 0 3
rlabel polysilicon 429 -1530 429 -1530 0 1
rlabel polysilicon 429 -1536 429 -1536 0 3
rlabel polysilicon 436 -1530 436 -1530 0 1
rlabel polysilicon 436 -1536 436 -1536 0 3
rlabel polysilicon 443 -1530 443 -1530 0 1
rlabel polysilicon 443 -1536 443 -1536 0 3
rlabel polysilicon 450 -1530 450 -1530 0 1
rlabel polysilicon 450 -1536 450 -1536 0 3
rlabel polysilicon 457 -1530 457 -1530 0 1
rlabel polysilicon 457 -1536 457 -1536 0 3
rlabel polysilicon 464 -1530 464 -1530 0 1
rlabel polysilicon 471 -1530 471 -1530 0 1
rlabel polysilicon 471 -1536 471 -1536 0 3
rlabel polysilicon 478 -1530 478 -1530 0 1
rlabel polysilicon 478 -1536 478 -1536 0 3
rlabel polysilicon 488 -1530 488 -1530 0 2
rlabel polysilicon 488 -1536 488 -1536 0 4
rlabel polysilicon 492 -1530 492 -1530 0 1
rlabel polysilicon 492 -1536 492 -1536 0 3
rlabel polysilicon 499 -1530 499 -1530 0 1
rlabel polysilicon 499 -1536 499 -1536 0 3
rlabel polysilicon 506 -1530 506 -1530 0 1
rlabel polysilicon 509 -1530 509 -1530 0 2
rlabel polysilicon 509 -1536 509 -1536 0 4
rlabel polysilicon 516 -1530 516 -1530 0 2
rlabel polysilicon 513 -1536 513 -1536 0 3
rlabel polysilicon 520 -1530 520 -1530 0 1
rlabel polysilicon 523 -1530 523 -1530 0 2
rlabel polysilicon 520 -1536 520 -1536 0 3
rlabel polysilicon 527 -1536 527 -1536 0 3
rlabel polysilicon 534 -1530 534 -1530 0 1
rlabel polysilicon 537 -1530 537 -1530 0 2
rlabel polysilicon 537 -1536 537 -1536 0 4
rlabel polysilicon 541 -1530 541 -1530 0 1
rlabel polysilicon 544 -1530 544 -1530 0 2
rlabel polysilicon 548 -1530 548 -1530 0 1
rlabel polysilicon 548 -1536 548 -1536 0 3
rlabel polysilicon 555 -1530 555 -1530 0 1
rlabel polysilicon 555 -1536 555 -1536 0 3
rlabel polysilicon 565 -1530 565 -1530 0 2
rlabel polysilicon 565 -1536 565 -1536 0 4
rlabel polysilicon 569 -1530 569 -1530 0 1
rlabel polysilicon 569 -1536 569 -1536 0 3
rlabel polysilicon 576 -1530 576 -1530 0 1
rlabel polysilicon 576 -1536 576 -1536 0 3
rlabel polysilicon 583 -1530 583 -1530 0 1
rlabel polysilicon 583 -1536 583 -1536 0 3
rlabel polysilicon 590 -1530 590 -1530 0 1
rlabel polysilicon 593 -1530 593 -1530 0 2
rlabel polysilicon 590 -1536 590 -1536 0 3
rlabel polysilicon 597 -1530 597 -1530 0 1
rlabel polysilicon 597 -1536 597 -1536 0 3
rlabel polysilicon 604 -1530 604 -1530 0 1
rlabel polysilicon 611 -1530 611 -1530 0 1
rlabel polysilicon 611 -1536 611 -1536 0 3
rlabel polysilicon 618 -1536 618 -1536 0 3
rlabel polysilicon 625 -1530 625 -1530 0 1
rlabel polysilicon 625 -1536 625 -1536 0 3
rlabel polysilicon 632 -1530 632 -1530 0 1
rlabel polysilicon 632 -1536 632 -1536 0 3
rlabel polysilicon 639 -1530 639 -1530 0 1
rlabel polysilicon 639 -1536 639 -1536 0 3
rlabel polysilicon 646 -1530 646 -1530 0 1
rlabel polysilicon 646 -1536 646 -1536 0 3
rlabel polysilicon 653 -1530 653 -1530 0 1
rlabel polysilicon 653 -1536 653 -1536 0 3
rlabel polysilicon 660 -1530 660 -1530 0 1
rlabel polysilicon 660 -1536 660 -1536 0 3
rlabel polysilicon 663 -1536 663 -1536 0 4
rlabel polysilicon 667 -1530 667 -1530 0 1
rlabel polysilicon 667 -1536 667 -1536 0 3
rlabel polysilicon 674 -1530 674 -1530 0 1
rlabel polysilicon 674 -1536 674 -1536 0 3
rlabel polysilicon 681 -1530 681 -1530 0 1
rlabel polysilicon 684 -1530 684 -1530 0 2
rlabel polysilicon 684 -1536 684 -1536 0 4
rlabel polysilicon 688 -1530 688 -1530 0 1
rlabel polysilicon 688 -1536 688 -1536 0 3
rlabel polysilicon 695 -1530 695 -1530 0 1
rlabel polysilicon 695 -1536 695 -1536 0 3
rlabel polysilicon 702 -1530 702 -1530 0 1
rlabel polysilicon 702 -1536 702 -1536 0 3
rlabel polysilicon 709 -1530 709 -1530 0 1
rlabel polysilicon 709 -1536 709 -1536 0 3
rlabel polysilicon 716 -1536 716 -1536 0 3
rlabel polysilicon 723 -1530 723 -1530 0 1
rlabel polysilicon 726 -1530 726 -1530 0 2
rlabel polysilicon 726 -1536 726 -1536 0 4
rlabel polysilicon 730 -1530 730 -1530 0 1
rlabel polysilicon 730 -1536 730 -1536 0 3
rlabel polysilicon 740 -1530 740 -1530 0 2
rlabel polysilicon 737 -1536 737 -1536 0 3
rlabel polysilicon 740 -1536 740 -1536 0 4
rlabel polysilicon 744 -1530 744 -1530 0 1
rlabel polysilicon 747 -1530 747 -1530 0 2
rlabel polysilicon 744 -1536 744 -1536 0 3
rlabel polysilicon 751 -1530 751 -1530 0 1
rlabel polysilicon 751 -1536 751 -1536 0 3
rlabel polysilicon 758 -1530 758 -1530 0 1
rlabel polysilicon 758 -1536 758 -1536 0 3
rlabel polysilicon 765 -1530 765 -1530 0 1
rlabel polysilicon 765 -1536 765 -1536 0 3
rlabel polysilicon 772 -1530 772 -1530 0 1
rlabel polysilicon 772 -1536 772 -1536 0 3
rlabel polysilicon 779 -1530 779 -1530 0 1
rlabel polysilicon 779 -1536 779 -1536 0 3
rlabel polysilicon 786 -1530 786 -1530 0 1
rlabel polysilicon 786 -1536 786 -1536 0 3
rlabel polysilicon 793 -1530 793 -1530 0 1
rlabel polysilicon 793 -1536 793 -1536 0 3
rlabel polysilicon 800 -1530 800 -1530 0 1
rlabel polysilicon 800 -1536 800 -1536 0 3
rlabel polysilicon 807 -1530 807 -1530 0 1
rlabel polysilicon 807 -1536 807 -1536 0 3
rlabel polysilicon 814 -1530 814 -1530 0 1
rlabel polysilicon 814 -1536 814 -1536 0 3
rlabel polysilicon 821 -1530 821 -1530 0 1
rlabel polysilicon 821 -1536 821 -1536 0 3
rlabel polysilicon 828 -1530 828 -1530 0 1
rlabel polysilicon 828 -1536 828 -1536 0 3
rlabel polysilicon 835 -1530 835 -1530 0 1
rlabel polysilicon 835 -1536 835 -1536 0 3
rlabel polysilicon 842 -1530 842 -1530 0 1
rlabel polysilicon 845 -1530 845 -1530 0 2
rlabel polysilicon 849 -1530 849 -1530 0 1
rlabel polysilicon 849 -1536 849 -1536 0 3
rlabel polysilicon 856 -1530 856 -1530 0 1
rlabel polysilicon 856 -1536 856 -1536 0 3
rlabel polysilicon 863 -1530 863 -1530 0 1
rlabel polysilicon 863 -1536 863 -1536 0 3
rlabel polysilicon 870 -1530 870 -1530 0 1
rlabel polysilicon 870 -1536 870 -1536 0 3
rlabel polysilicon 877 -1530 877 -1530 0 1
rlabel polysilicon 877 -1536 877 -1536 0 3
rlabel polysilicon 884 -1530 884 -1530 0 1
rlabel polysilicon 884 -1536 884 -1536 0 3
rlabel polysilicon 891 -1530 891 -1530 0 1
rlabel polysilicon 891 -1536 891 -1536 0 3
rlabel polysilicon 898 -1530 898 -1530 0 1
rlabel polysilicon 898 -1536 898 -1536 0 3
rlabel polysilicon 905 -1530 905 -1530 0 1
rlabel polysilicon 905 -1536 905 -1536 0 3
rlabel polysilicon 912 -1530 912 -1530 0 1
rlabel polysilicon 912 -1536 912 -1536 0 3
rlabel polysilicon 919 -1530 919 -1530 0 1
rlabel polysilicon 919 -1536 919 -1536 0 3
rlabel polysilicon 926 -1530 926 -1530 0 1
rlabel polysilicon 926 -1536 926 -1536 0 3
rlabel polysilicon 933 -1530 933 -1530 0 1
rlabel polysilicon 933 -1536 933 -1536 0 3
rlabel polysilicon 940 -1530 940 -1530 0 1
rlabel polysilicon 940 -1536 940 -1536 0 3
rlabel polysilicon 947 -1530 947 -1530 0 1
rlabel polysilicon 947 -1536 947 -1536 0 3
rlabel polysilicon 954 -1530 954 -1530 0 1
rlabel polysilicon 954 -1536 954 -1536 0 3
rlabel polysilicon 961 -1530 961 -1530 0 1
rlabel polysilicon 961 -1536 961 -1536 0 3
rlabel polysilicon 968 -1530 968 -1530 0 1
rlabel polysilicon 968 -1536 968 -1536 0 3
rlabel polysilicon 975 -1530 975 -1530 0 1
rlabel polysilicon 975 -1536 975 -1536 0 3
rlabel polysilicon 982 -1530 982 -1530 0 1
rlabel polysilicon 982 -1536 982 -1536 0 3
rlabel polysilicon 989 -1530 989 -1530 0 1
rlabel polysilicon 989 -1536 989 -1536 0 3
rlabel polysilicon 996 -1530 996 -1530 0 1
rlabel polysilicon 999 -1530 999 -1530 0 2
rlabel polysilicon 996 -1536 996 -1536 0 3
rlabel polysilicon 1003 -1530 1003 -1530 0 1
rlabel polysilicon 1003 -1536 1003 -1536 0 3
rlabel polysilicon 1010 -1530 1010 -1530 0 1
rlabel polysilicon 1010 -1536 1010 -1536 0 3
rlabel polysilicon 1017 -1530 1017 -1530 0 1
rlabel polysilicon 1017 -1536 1017 -1536 0 3
rlabel polysilicon 1045 -1530 1045 -1530 0 1
rlabel polysilicon 1045 -1536 1045 -1536 0 3
rlabel polysilicon 1052 -1530 1052 -1530 0 1
rlabel polysilicon 1052 -1536 1052 -1536 0 3
rlabel polysilicon 1059 -1530 1059 -1530 0 1
rlabel polysilicon 23 -1607 23 -1607 0 1
rlabel polysilicon 23 -1613 23 -1613 0 3
rlabel polysilicon 30 -1607 30 -1607 0 1
rlabel polysilicon 30 -1613 30 -1613 0 3
rlabel polysilicon 37 -1607 37 -1607 0 1
rlabel polysilicon 37 -1613 37 -1613 0 3
rlabel polysilicon 44 -1607 44 -1607 0 1
rlabel polysilicon 44 -1613 44 -1613 0 3
rlabel polysilicon 51 -1607 51 -1607 0 1
rlabel polysilicon 51 -1613 51 -1613 0 3
rlabel polysilicon 58 -1607 58 -1607 0 1
rlabel polysilicon 58 -1613 58 -1613 0 3
rlabel polysilicon 68 -1607 68 -1607 0 2
rlabel polysilicon 68 -1613 68 -1613 0 4
rlabel polysilicon 72 -1607 72 -1607 0 1
rlabel polysilicon 79 -1607 79 -1607 0 1
rlabel polysilicon 79 -1613 79 -1613 0 3
rlabel polysilicon 86 -1607 86 -1607 0 1
rlabel polysilicon 86 -1613 86 -1613 0 3
rlabel polysilicon 93 -1607 93 -1607 0 1
rlabel polysilicon 93 -1613 93 -1613 0 3
rlabel polysilicon 100 -1607 100 -1607 0 1
rlabel polysilicon 100 -1613 100 -1613 0 3
rlabel polysilicon 107 -1607 107 -1607 0 1
rlabel polysilicon 107 -1613 107 -1613 0 3
rlabel polysilicon 110 -1613 110 -1613 0 4
rlabel polysilicon 114 -1607 114 -1607 0 1
rlabel polysilicon 114 -1613 114 -1613 0 3
rlabel polysilicon 121 -1607 121 -1607 0 1
rlabel polysilicon 121 -1613 121 -1613 0 3
rlabel polysilicon 128 -1607 128 -1607 0 1
rlabel polysilicon 128 -1613 128 -1613 0 3
rlabel polysilicon 135 -1607 135 -1607 0 1
rlabel polysilicon 135 -1613 135 -1613 0 3
rlabel polysilicon 142 -1607 142 -1607 0 1
rlabel polysilicon 142 -1613 142 -1613 0 3
rlabel polysilicon 152 -1607 152 -1607 0 2
rlabel polysilicon 152 -1613 152 -1613 0 4
rlabel polysilicon 156 -1607 156 -1607 0 1
rlabel polysilicon 156 -1613 156 -1613 0 3
rlabel polysilicon 159 -1613 159 -1613 0 4
rlabel polysilicon 163 -1607 163 -1607 0 1
rlabel polysilicon 163 -1613 163 -1613 0 3
rlabel polysilicon 173 -1607 173 -1607 0 2
rlabel polysilicon 170 -1613 170 -1613 0 3
rlabel polysilicon 177 -1607 177 -1607 0 1
rlabel polysilicon 177 -1613 177 -1613 0 3
rlabel polysilicon 184 -1607 184 -1607 0 1
rlabel polysilicon 184 -1613 184 -1613 0 3
rlabel polysilicon 191 -1607 191 -1607 0 1
rlabel polysilicon 191 -1613 191 -1613 0 3
rlabel polysilicon 198 -1613 198 -1613 0 3
rlabel polysilicon 201 -1613 201 -1613 0 4
rlabel polysilicon 205 -1607 205 -1607 0 1
rlabel polysilicon 205 -1613 205 -1613 0 3
rlabel polysilicon 212 -1607 212 -1607 0 1
rlabel polysilicon 212 -1613 212 -1613 0 3
rlabel polysilicon 219 -1607 219 -1607 0 1
rlabel polysilicon 219 -1613 219 -1613 0 3
rlabel polysilicon 226 -1613 226 -1613 0 3
rlabel polysilicon 229 -1613 229 -1613 0 4
rlabel polysilicon 233 -1607 233 -1607 0 1
rlabel polysilicon 233 -1613 233 -1613 0 3
rlabel polysilicon 240 -1607 240 -1607 0 1
rlabel polysilicon 240 -1613 240 -1613 0 3
rlabel polysilicon 247 -1607 247 -1607 0 1
rlabel polysilicon 247 -1613 247 -1613 0 3
rlabel polysilicon 254 -1607 254 -1607 0 1
rlabel polysilicon 254 -1613 254 -1613 0 3
rlabel polysilicon 261 -1607 261 -1607 0 1
rlabel polysilicon 261 -1613 261 -1613 0 3
rlabel polysilicon 268 -1607 268 -1607 0 1
rlabel polysilicon 268 -1613 268 -1613 0 3
rlabel polysilicon 275 -1607 275 -1607 0 1
rlabel polysilicon 275 -1613 275 -1613 0 3
rlabel polysilicon 282 -1607 282 -1607 0 1
rlabel polysilicon 282 -1613 282 -1613 0 3
rlabel polysilicon 289 -1607 289 -1607 0 1
rlabel polysilicon 289 -1613 289 -1613 0 3
rlabel polysilicon 296 -1607 296 -1607 0 1
rlabel polysilicon 296 -1613 296 -1613 0 3
rlabel polysilicon 306 -1607 306 -1607 0 2
rlabel polysilicon 303 -1613 303 -1613 0 3
rlabel polysilicon 306 -1613 306 -1613 0 4
rlabel polysilicon 313 -1607 313 -1607 0 2
rlabel polysilicon 310 -1613 310 -1613 0 3
rlabel polysilicon 313 -1613 313 -1613 0 4
rlabel polysilicon 317 -1607 317 -1607 0 1
rlabel polysilicon 317 -1613 317 -1613 0 3
rlabel polysilicon 324 -1607 324 -1607 0 1
rlabel polysilicon 324 -1613 324 -1613 0 3
rlabel polysilicon 331 -1607 331 -1607 0 1
rlabel polysilicon 331 -1613 331 -1613 0 3
rlabel polysilicon 338 -1607 338 -1607 0 1
rlabel polysilicon 338 -1613 338 -1613 0 3
rlabel polysilicon 345 -1607 345 -1607 0 1
rlabel polysilicon 345 -1613 345 -1613 0 3
rlabel polysilicon 355 -1607 355 -1607 0 2
rlabel polysilicon 352 -1613 352 -1613 0 3
rlabel polysilicon 355 -1613 355 -1613 0 4
rlabel polysilicon 359 -1607 359 -1607 0 1
rlabel polysilicon 359 -1613 359 -1613 0 3
rlabel polysilicon 366 -1607 366 -1607 0 1
rlabel polysilicon 366 -1613 366 -1613 0 3
rlabel polysilicon 373 -1607 373 -1607 0 1
rlabel polysilicon 373 -1613 373 -1613 0 3
rlabel polysilicon 376 -1613 376 -1613 0 4
rlabel polysilicon 380 -1607 380 -1607 0 1
rlabel polysilicon 380 -1613 380 -1613 0 3
rlabel polysilicon 387 -1607 387 -1607 0 1
rlabel polysilicon 390 -1613 390 -1613 0 4
rlabel polysilicon 394 -1607 394 -1607 0 1
rlabel polysilicon 394 -1613 394 -1613 0 3
rlabel polysilicon 401 -1607 401 -1607 0 1
rlabel polysilicon 401 -1613 401 -1613 0 3
rlabel polysilicon 408 -1607 408 -1607 0 1
rlabel polysilicon 408 -1613 408 -1613 0 3
rlabel polysilicon 415 -1607 415 -1607 0 1
rlabel polysilicon 415 -1613 415 -1613 0 3
rlabel polysilicon 425 -1607 425 -1607 0 2
rlabel polysilicon 422 -1613 422 -1613 0 3
rlabel polysilicon 425 -1613 425 -1613 0 4
rlabel polysilicon 429 -1607 429 -1607 0 1
rlabel polysilicon 429 -1613 429 -1613 0 3
rlabel polysilicon 436 -1607 436 -1607 0 1
rlabel polysilicon 436 -1613 436 -1613 0 3
rlabel polysilicon 443 -1607 443 -1607 0 1
rlabel polysilicon 443 -1613 443 -1613 0 3
rlabel polysilicon 450 -1607 450 -1607 0 1
rlabel polysilicon 450 -1613 450 -1613 0 3
rlabel polysilicon 457 -1607 457 -1607 0 1
rlabel polysilicon 457 -1613 457 -1613 0 3
rlabel polysilicon 464 -1607 464 -1607 0 1
rlabel polysilicon 464 -1613 464 -1613 0 3
rlabel polysilicon 471 -1607 471 -1607 0 1
rlabel polysilicon 471 -1613 471 -1613 0 3
rlabel polysilicon 478 -1607 478 -1607 0 1
rlabel polysilicon 478 -1613 478 -1613 0 3
rlabel polysilicon 485 -1607 485 -1607 0 1
rlabel polysilicon 485 -1613 485 -1613 0 3
rlabel polysilicon 492 -1607 492 -1607 0 1
rlabel polysilicon 492 -1613 492 -1613 0 3
rlabel polysilicon 499 -1607 499 -1607 0 1
rlabel polysilicon 499 -1613 499 -1613 0 3
rlabel polysilicon 506 -1607 506 -1607 0 1
rlabel polysilicon 506 -1613 506 -1613 0 3
rlabel polysilicon 513 -1607 513 -1607 0 1
rlabel polysilicon 513 -1613 513 -1613 0 3
rlabel polysilicon 523 -1613 523 -1613 0 4
rlabel polysilicon 530 -1607 530 -1607 0 2
rlabel polysilicon 530 -1613 530 -1613 0 4
rlabel polysilicon 534 -1607 534 -1607 0 1
rlabel polysilicon 534 -1613 534 -1613 0 3
rlabel polysilicon 541 -1607 541 -1607 0 1
rlabel polysilicon 541 -1613 541 -1613 0 3
rlabel polysilicon 548 -1607 548 -1607 0 1
rlabel polysilicon 548 -1613 548 -1613 0 3
rlabel polysilicon 555 -1607 555 -1607 0 1
rlabel polysilicon 558 -1607 558 -1607 0 2
rlabel polysilicon 555 -1613 555 -1613 0 3
rlabel polysilicon 562 -1607 562 -1607 0 1
rlabel polysilicon 565 -1607 565 -1607 0 2
rlabel polysilicon 562 -1613 562 -1613 0 3
rlabel polysilicon 565 -1613 565 -1613 0 4
rlabel polysilicon 572 -1607 572 -1607 0 2
rlabel polysilicon 569 -1613 569 -1613 0 3
rlabel polysilicon 576 -1607 576 -1607 0 1
rlabel polysilicon 576 -1613 576 -1613 0 3
rlabel polysilicon 583 -1607 583 -1607 0 1
rlabel polysilicon 583 -1613 583 -1613 0 3
rlabel polysilicon 590 -1607 590 -1607 0 1
rlabel polysilicon 590 -1613 590 -1613 0 3
rlabel polysilicon 597 -1607 597 -1607 0 1
rlabel polysilicon 597 -1613 597 -1613 0 3
rlabel polysilicon 604 -1607 604 -1607 0 1
rlabel polysilicon 604 -1613 604 -1613 0 3
rlabel polysilicon 614 -1613 614 -1613 0 4
rlabel polysilicon 618 -1607 618 -1607 0 1
rlabel polysilicon 618 -1613 618 -1613 0 3
rlabel polysilicon 628 -1607 628 -1607 0 2
rlabel polysilicon 632 -1607 632 -1607 0 1
rlabel polysilicon 632 -1613 632 -1613 0 3
rlabel polysilicon 639 -1607 639 -1607 0 1
rlabel polysilicon 639 -1613 639 -1613 0 3
rlabel polysilicon 646 -1607 646 -1607 0 1
rlabel polysilicon 646 -1613 646 -1613 0 3
rlabel polysilicon 653 -1607 653 -1607 0 1
rlabel polysilicon 653 -1613 653 -1613 0 3
rlabel polysilicon 660 -1607 660 -1607 0 1
rlabel polysilicon 660 -1613 660 -1613 0 3
rlabel polysilicon 667 -1607 667 -1607 0 1
rlabel polysilicon 667 -1613 667 -1613 0 3
rlabel polysilicon 674 -1607 674 -1607 0 1
rlabel polysilicon 674 -1613 674 -1613 0 3
rlabel polysilicon 681 -1613 681 -1613 0 3
rlabel polysilicon 684 -1613 684 -1613 0 4
rlabel polysilicon 688 -1607 688 -1607 0 1
rlabel polysilicon 688 -1613 688 -1613 0 3
rlabel polysilicon 695 -1607 695 -1607 0 1
rlabel polysilicon 695 -1613 695 -1613 0 3
rlabel polysilicon 702 -1607 702 -1607 0 1
rlabel polysilicon 702 -1613 702 -1613 0 3
rlabel polysilicon 709 -1607 709 -1607 0 1
rlabel polysilicon 709 -1613 709 -1613 0 3
rlabel polysilicon 716 -1607 716 -1607 0 1
rlabel polysilicon 716 -1613 716 -1613 0 3
rlabel polysilicon 723 -1607 723 -1607 0 1
rlabel polysilicon 723 -1613 723 -1613 0 3
rlabel polysilicon 730 -1607 730 -1607 0 1
rlabel polysilicon 730 -1613 730 -1613 0 3
rlabel polysilicon 737 -1607 737 -1607 0 1
rlabel polysilicon 737 -1613 737 -1613 0 3
rlabel polysilicon 744 -1607 744 -1607 0 1
rlabel polysilicon 744 -1613 744 -1613 0 3
rlabel polysilicon 751 -1607 751 -1607 0 1
rlabel polysilicon 751 -1613 751 -1613 0 3
rlabel polysilicon 758 -1607 758 -1607 0 1
rlabel polysilicon 758 -1613 758 -1613 0 3
rlabel polysilicon 765 -1607 765 -1607 0 1
rlabel polysilicon 765 -1613 765 -1613 0 3
rlabel polysilicon 772 -1607 772 -1607 0 1
rlabel polysilicon 772 -1613 772 -1613 0 3
rlabel polysilicon 779 -1607 779 -1607 0 1
rlabel polysilicon 779 -1613 779 -1613 0 3
rlabel polysilicon 786 -1607 786 -1607 0 1
rlabel polysilicon 786 -1613 786 -1613 0 3
rlabel polysilicon 793 -1607 793 -1607 0 1
rlabel polysilicon 793 -1613 793 -1613 0 3
rlabel polysilicon 800 -1607 800 -1607 0 1
rlabel polysilicon 800 -1613 800 -1613 0 3
rlabel polysilicon 807 -1607 807 -1607 0 1
rlabel polysilicon 807 -1613 807 -1613 0 3
rlabel polysilicon 814 -1607 814 -1607 0 1
rlabel polysilicon 814 -1613 814 -1613 0 3
rlabel polysilicon 821 -1607 821 -1607 0 1
rlabel polysilicon 821 -1613 821 -1613 0 3
rlabel polysilicon 828 -1607 828 -1607 0 1
rlabel polysilicon 828 -1613 828 -1613 0 3
rlabel polysilicon 835 -1607 835 -1607 0 1
rlabel polysilicon 835 -1613 835 -1613 0 3
rlabel polysilicon 842 -1607 842 -1607 0 1
rlabel polysilicon 842 -1613 842 -1613 0 3
rlabel polysilicon 849 -1607 849 -1607 0 1
rlabel polysilicon 849 -1613 849 -1613 0 3
rlabel polysilicon 856 -1607 856 -1607 0 1
rlabel polysilicon 859 -1613 859 -1613 0 4
rlabel polysilicon 863 -1607 863 -1607 0 1
rlabel polysilicon 863 -1613 863 -1613 0 3
rlabel polysilicon 870 -1607 870 -1607 0 1
rlabel polysilicon 870 -1613 870 -1613 0 3
rlabel polysilicon 877 -1607 877 -1607 0 1
rlabel polysilicon 877 -1613 877 -1613 0 3
rlabel polysilicon 884 -1607 884 -1607 0 1
rlabel polysilicon 884 -1613 884 -1613 0 3
rlabel polysilicon 891 -1607 891 -1607 0 1
rlabel polysilicon 891 -1613 891 -1613 0 3
rlabel polysilicon 898 -1607 898 -1607 0 1
rlabel polysilicon 898 -1613 898 -1613 0 3
rlabel polysilicon 905 -1607 905 -1607 0 1
rlabel polysilicon 905 -1613 905 -1613 0 3
rlabel polysilicon 912 -1607 912 -1607 0 1
rlabel polysilicon 912 -1613 912 -1613 0 3
rlabel polysilicon 919 -1607 919 -1607 0 1
rlabel polysilicon 919 -1613 919 -1613 0 3
rlabel polysilicon 926 -1607 926 -1607 0 1
rlabel polysilicon 926 -1613 926 -1613 0 3
rlabel polysilicon 936 -1607 936 -1607 0 2
rlabel polysilicon 936 -1613 936 -1613 0 4
rlabel polysilicon 940 -1607 940 -1607 0 1
rlabel polysilicon 940 -1613 940 -1613 0 3
rlabel polysilicon 947 -1607 947 -1607 0 1
rlabel polysilicon 947 -1613 947 -1613 0 3
rlabel polysilicon 954 -1607 954 -1607 0 1
rlabel polysilicon 954 -1613 954 -1613 0 3
rlabel polysilicon 961 -1607 961 -1607 0 1
rlabel polysilicon 961 -1613 961 -1613 0 3
rlabel polysilicon 1024 -1607 1024 -1607 0 1
rlabel polysilicon 1024 -1613 1024 -1613 0 3
rlabel polysilicon 1038 -1607 1038 -1607 0 1
rlabel polysilicon 1038 -1613 1038 -1613 0 3
rlabel polysilicon 1045 -1613 1045 -1613 0 3
rlabel polysilicon 1052 -1607 1052 -1607 0 1
rlabel polysilicon 37 -1672 37 -1672 0 1
rlabel polysilicon 40 -1672 40 -1672 0 2
rlabel polysilicon 44 -1672 44 -1672 0 1
rlabel polysilicon 47 -1678 47 -1678 0 4
rlabel polysilicon 51 -1672 51 -1672 0 1
rlabel polysilicon 51 -1678 51 -1678 0 3
rlabel polysilicon 65 -1672 65 -1672 0 1
rlabel polysilicon 65 -1678 65 -1678 0 3
rlabel polysilicon 72 -1672 72 -1672 0 1
rlabel polysilicon 75 -1678 75 -1678 0 4
rlabel polysilicon 79 -1672 79 -1672 0 1
rlabel polysilicon 86 -1672 86 -1672 0 1
rlabel polysilicon 86 -1678 86 -1678 0 3
rlabel polysilicon 93 -1672 93 -1672 0 1
rlabel polysilicon 93 -1678 93 -1678 0 3
rlabel polysilicon 100 -1672 100 -1672 0 1
rlabel polysilicon 100 -1678 100 -1678 0 3
rlabel polysilicon 107 -1672 107 -1672 0 1
rlabel polysilicon 107 -1678 107 -1678 0 3
rlabel polysilicon 114 -1672 114 -1672 0 1
rlabel polysilicon 117 -1678 117 -1678 0 4
rlabel polysilicon 121 -1672 121 -1672 0 1
rlabel polysilicon 121 -1678 121 -1678 0 3
rlabel polysilicon 128 -1672 128 -1672 0 1
rlabel polysilicon 128 -1678 128 -1678 0 3
rlabel polysilicon 135 -1672 135 -1672 0 1
rlabel polysilicon 135 -1678 135 -1678 0 3
rlabel polysilicon 142 -1672 142 -1672 0 1
rlabel polysilicon 142 -1678 142 -1678 0 3
rlabel polysilicon 149 -1672 149 -1672 0 1
rlabel polysilicon 152 -1672 152 -1672 0 2
rlabel polysilicon 156 -1672 156 -1672 0 1
rlabel polysilicon 156 -1678 156 -1678 0 3
rlabel polysilicon 163 -1672 163 -1672 0 1
rlabel polysilicon 163 -1678 163 -1678 0 3
rlabel polysilicon 170 -1672 170 -1672 0 1
rlabel polysilicon 170 -1678 170 -1678 0 3
rlabel polysilicon 177 -1678 177 -1678 0 3
rlabel polysilicon 180 -1678 180 -1678 0 4
rlabel polysilicon 184 -1672 184 -1672 0 1
rlabel polysilicon 184 -1678 184 -1678 0 3
rlabel polysilicon 191 -1672 191 -1672 0 1
rlabel polysilicon 191 -1678 191 -1678 0 3
rlabel polysilicon 198 -1678 198 -1678 0 3
rlabel polysilicon 201 -1678 201 -1678 0 4
rlabel polysilicon 205 -1672 205 -1672 0 1
rlabel polysilicon 208 -1672 208 -1672 0 2
rlabel polysilicon 212 -1672 212 -1672 0 1
rlabel polysilicon 212 -1678 212 -1678 0 3
rlabel polysilicon 219 -1672 219 -1672 0 1
rlabel polysilicon 219 -1678 219 -1678 0 3
rlabel polysilicon 226 -1672 226 -1672 0 1
rlabel polysilicon 226 -1678 226 -1678 0 3
rlabel polysilicon 233 -1672 233 -1672 0 1
rlabel polysilicon 233 -1678 233 -1678 0 3
rlabel polysilicon 240 -1672 240 -1672 0 1
rlabel polysilicon 240 -1678 240 -1678 0 3
rlabel polysilicon 247 -1672 247 -1672 0 1
rlabel polysilicon 247 -1678 247 -1678 0 3
rlabel polysilicon 257 -1672 257 -1672 0 2
rlabel polysilicon 261 -1672 261 -1672 0 1
rlabel polysilicon 261 -1678 261 -1678 0 3
rlabel polysilicon 268 -1672 268 -1672 0 1
rlabel polysilicon 268 -1678 268 -1678 0 3
rlabel polysilicon 275 -1672 275 -1672 0 1
rlabel polysilicon 275 -1678 275 -1678 0 3
rlabel polysilicon 282 -1672 282 -1672 0 1
rlabel polysilicon 282 -1678 282 -1678 0 3
rlabel polysilicon 289 -1672 289 -1672 0 1
rlabel polysilicon 289 -1678 289 -1678 0 3
rlabel polysilicon 296 -1672 296 -1672 0 1
rlabel polysilicon 303 -1672 303 -1672 0 1
rlabel polysilicon 306 -1672 306 -1672 0 2
rlabel polysilicon 306 -1678 306 -1678 0 4
rlabel polysilicon 310 -1672 310 -1672 0 1
rlabel polysilicon 310 -1678 310 -1678 0 3
rlabel polysilicon 317 -1672 317 -1672 0 1
rlabel polysilicon 317 -1678 317 -1678 0 3
rlabel polysilicon 324 -1672 324 -1672 0 1
rlabel polysilicon 324 -1678 324 -1678 0 3
rlabel polysilicon 331 -1672 331 -1672 0 1
rlabel polysilicon 334 -1672 334 -1672 0 2
rlabel polysilicon 331 -1678 331 -1678 0 3
rlabel polysilicon 334 -1678 334 -1678 0 4
rlabel polysilicon 341 -1678 341 -1678 0 4
rlabel polysilicon 345 -1672 345 -1672 0 1
rlabel polysilicon 345 -1678 345 -1678 0 3
rlabel polysilicon 352 -1672 352 -1672 0 1
rlabel polysilicon 352 -1678 352 -1678 0 3
rlabel polysilicon 359 -1672 359 -1672 0 1
rlabel polysilicon 359 -1678 359 -1678 0 3
rlabel polysilicon 366 -1672 366 -1672 0 1
rlabel polysilicon 366 -1678 366 -1678 0 3
rlabel polysilicon 373 -1672 373 -1672 0 1
rlabel polysilicon 373 -1678 373 -1678 0 3
rlabel polysilicon 380 -1672 380 -1672 0 1
rlabel polysilicon 380 -1678 380 -1678 0 3
rlabel polysilicon 387 -1672 387 -1672 0 1
rlabel polysilicon 387 -1678 387 -1678 0 3
rlabel polysilicon 394 -1672 394 -1672 0 1
rlabel polysilicon 394 -1678 394 -1678 0 3
rlabel polysilicon 401 -1672 401 -1672 0 1
rlabel polysilicon 404 -1672 404 -1672 0 2
rlabel polysilicon 401 -1678 401 -1678 0 3
rlabel polysilicon 411 -1672 411 -1672 0 2
rlabel polysilicon 408 -1678 408 -1678 0 3
rlabel polysilicon 415 -1672 415 -1672 0 1
rlabel polysilicon 415 -1678 415 -1678 0 3
rlabel polysilicon 422 -1672 422 -1672 0 1
rlabel polysilicon 422 -1678 422 -1678 0 3
rlabel polysilicon 425 -1678 425 -1678 0 4
rlabel polysilicon 429 -1672 429 -1672 0 1
rlabel polysilicon 432 -1672 432 -1672 0 2
rlabel polysilicon 432 -1678 432 -1678 0 4
rlabel polysilicon 436 -1672 436 -1672 0 1
rlabel polysilicon 436 -1678 436 -1678 0 3
rlabel polysilicon 443 -1672 443 -1672 0 1
rlabel polysilicon 443 -1678 443 -1678 0 3
rlabel polysilicon 450 -1672 450 -1672 0 1
rlabel polysilicon 450 -1678 450 -1678 0 3
rlabel polysilicon 457 -1672 457 -1672 0 1
rlabel polysilicon 457 -1678 457 -1678 0 3
rlabel polysilicon 464 -1672 464 -1672 0 1
rlabel polysilicon 464 -1678 464 -1678 0 3
rlabel polysilicon 471 -1672 471 -1672 0 1
rlabel polysilicon 471 -1678 471 -1678 0 3
rlabel polysilicon 478 -1672 478 -1672 0 1
rlabel polysilicon 478 -1678 478 -1678 0 3
rlabel polysilicon 485 -1672 485 -1672 0 1
rlabel polysilicon 485 -1678 485 -1678 0 3
rlabel polysilicon 492 -1672 492 -1672 0 1
rlabel polysilicon 492 -1678 492 -1678 0 3
rlabel polysilicon 499 -1672 499 -1672 0 1
rlabel polysilicon 499 -1678 499 -1678 0 3
rlabel polysilicon 506 -1672 506 -1672 0 1
rlabel polysilicon 506 -1678 506 -1678 0 3
rlabel polysilicon 513 -1672 513 -1672 0 1
rlabel polysilicon 516 -1672 516 -1672 0 2
rlabel polysilicon 520 -1672 520 -1672 0 1
rlabel polysilicon 523 -1672 523 -1672 0 2
rlabel polysilicon 520 -1678 520 -1678 0 3
rlabel polysilicon 523 -1678 523 -1678 0 4
rlabel polysilicon 527 -1672 527 -1672 0 1
rlabel polysilicon 527 -1678 527 -1678 0 3
rlabel polysilicon 534 -1672 534 -1672 0 1
rlabel polysilicon 534 -1678 534 -1678 0 3
rlabel polysilicon 541 -1672 541 -1672 0 1
rlabel polysilicon 544 -1672 544 -1672 0 2
rlabel polysilicon 551 -1672 551 -1672 0 2
rlabel polysilicon 548 -1678 548 -1678 0 3
rlabel polysilicon 555 -1672 555 -1672 0 1
rlabel polysilicon 555 -1678 555 -1678 0 3
rlabel polysilicon 562 -1672 562 -1672 0 1
rlabel polysilicon 562 -1678 562 -1678 0 3
rlabel polysilicon 569 -1672 569 -1672 0 1
rlabel polysilicon 569 -1678 569 -1678 0 3
rlabel polysilicon 576 -1672 576 -1672 0 1
rlabel polysilicon 576 -1678 576 -1678 0 3
rlabel polysilicon 583 -1672 583 -1672 0 1
rlabel polysilicon 583 -1678 583 -1678 0 3
rlabel polysilicon 590 -1672 590 -1672 0 1
rlabel polysilicon 590 -1678 590 -1678 0 3
rlabel polysilicon 597 -1672 597 -1672 0 1
rlabel polysilicon 597 -1678 597 -1678 0 3
rlabel polysilicon 604 -1672 604 -1672 0 1
rlabel polysilicon 604 -1678 604 -1678 0 3
rlabel polysilicon 611 -1672 611 -1672 0 1
rlabel polysilicon 611 -1678 611 -1678 0 3
rlabel polysilicon 625 -1672 625 -1672 0 1
rlabel polysilicon 625 -1678 625 -1678 0 3
rlabel polysilicon 632 -1672 632 -1672 0 1
rlabel polysilicon 632 -1678 632 -1678 0 3
rlabel polysilicon 646 -1672 646 -1672 0 1
rlabel polysilicon 646 -1678 646 -1678 0 3
rlabel polysilicon 667 -1672 667 -1672 0 1
rlabel polysilicon 667 -1678 667 -1678 0 3
rlabel polysilicon 677 -1678 677 -1678 0 4
rlabel polysilicon 681 -1672 681 -1672 0 1
rlabel polysilicon 681 -1678 681 -1678 0 3
rlabel polysilicon 688 -1672 688 -1672 0 1
rlabel polysilicon 688 -1678 688 -1678 0 3
rlabel polysilicon 691 -1678 691 -1678 0 4
rlabel polysilicon 695 -1672 695 -1672 0 1
rlabel polysilicon 695 -1678 695 -1678 0 3
rlabel polysilicon 702 -1672 702 -1672 0 1
rlabel polysilicon 702 -1678 702 -1678 0 3
rlabel polysilicon 709 -1672 709 -1672 0 1
rlabel polysilicon 709 -1678 709 -1678 0 3
rlabel polysilicon 716 -1672 716 -1672 0 1
rlabel polysilicon 716 -1678 716 -1678 0 3
rlabel polysilicon 723 -1672 723 -1672 0 1
rlabel polysilicon 723 -1678 723 -1678 0 3
rlabel polysilicon 733 -1672 733 -1672 0 2
rlabel polysilicon 737 -1672 737 -1672 0 1
rlabel polysilicon 737 -1678 737 -1678 0 3
rlabel polysilicon 744 -1672 744 -1672 0 1
rlabel polysilicon 744 -1678 744 -1678 0 3
rlabel polysilicon 751 -1672 751 -1672 0 1
rlabel polysilicon 751 -1678 751 -1678 0 3
rlabel polysilicon 758 -1672 758 -1672 0 1
rlabel polysilicon 758 -1678 758 -1678 0 3
rlabel polysilicon 765 -1672 765 -1672 0 1
rlabel polysilicon 765 -1678 765 -1678 0 3
rlabel polysilicon 775 -1672 775 -1672 0 2
rlabel polysilicon 779 -1672 779 -1672 0 1
rlabel polysilicon 782 -1678 782 -1678 0 4
rlabel polysilicon 786 -1672 786 -1672 0 1
rlabel polysilicon 786 -1678 786 -1678 0 3
rlabel polysilicon 793 -1672 793 -1672 0 1
rlabel polysilicon 793 -1678 793 -1678 0 3
rlabel polysilicon 800 -1672 800 -1672 0 1
rlabel polysilicon 803 -1672 803 -1672 0 2
rlabel polysilicon 807 -1672 807 -1672 0 1
rlabel polysilicon 807 -1678 807 -1678 0 3
rlabel polysilicon 814 -1672 814 -1672 0 1
rlabel polysilicon 814 -1678 814 -1678 0 3
rlabel polysilicon 821 -1672 821 -1672 0 1
rlabel polysilicon 821 -1678 821 -1678 0 3
rlabel polysilicon 828 -1672 828 -1672 0 1
rlabel polysilicon 828 -1678 828 -1678 0 3
rlabel polysilicon 835 -1672 835 -1672 0 1
rlabel polysilicon 838 -1672 838 -1672 0 2
rlabel polysilicon 842 -1672 842 -1672 0 1
rlabel polysilicon 842 -1678 842 -1678 0 3
rlabel polysilicon 849 -1678 849 -1678 0 3
rlabel polysilicon 852 -1678 852 -1678 0 4
rlabel polysilicon 863 -1672 863 -1672 0 1
rlabel polysilicon 863 -1678 863 -1678 0 3
rlabel polysilicon 884 -1672 884 -1672 0 1
rlabel polysilicon 884 -1678 884 -1678 0 3
rlabel polysilicon 891 -1672 891 -1672 0 1
rlabel polysilicon 891 -1678 891 -1678 0 3
rlabel polysilicon 905 -1672 905 -1672 0 1
rlabel polysilicon 905 -1678 905 -1678 0 3
rlabel polysilicon 968 -1672 968 -1672 0 1
rlabel polysilicon 968 -1678 968 -1678 0 3
rlabel polysilicon 1024 -1672 1024 -1672 0 1
rlabel polysilicon 1024 -1678 1024 -1678 0 3
rlabel polysilicon 44 -1709 44 -1709 0 1
rlabel polysilicon 44 -1715 44 -1715 0 3
rlabel polysilicon 58 -1709 58 -1709 0 1
rlabel polysilicon 58 -1715 58 -1715 0 3
rlabel polysilicon 93 -1709 93 -1709 0 1
rlabel polysilicon 93 -1715 93 -1715 0 3
rlabel polysilicon 103 -1709 103 -1709 0 2
rlabel polysilicon 100 -1715 100 -1715 0 3
rlabel polysilicon 103 -1715 103 -1715 0 4
rlabel polysilicon 114 -1709 114 -1709 0 1
rlabel polysilicon 117 -1715 117 -1715 0 4
rlabel polysilicon 128 -1709 128 -1709 0 1
rlabel polysilicon 128 -1715 128 -1715 0 3
rlabel polysilicon 142 -1709 142 -1709 0 1
rlabel polysilicon 142 -1715 142 -1715 0 3
rlabel polysilicon 149 -1709 149 -1709 0 1
rlabel polysilicon 149 -1715 149 -1715 0 3
rlabel polysilicon 156 -1709 156 -1709 0 1
rlabel polysilicon 156 -1715 156 -1715 0 3
rlabel polysilicon 163 -1709 163 -1709 0 1
rlabel polysilicon 163 -1715 163 -1715 0 3
rlabel polysilicon 170 -1709 170 -1709 0 1
rlabel polysilicon 170 -1715 170 -1715 0 3
rlabel polysilicon 177 -1709 177 -1709 0 1
rlabel polysilicon 180 -1709 180 -1709 0 2
rlabel polysilicon 184 -1715 184 -1715 0 3
rlabel polysilicon 191 -1709 191 -1709 0 1
rlabel polysilicon 191 -1715 191 -1715 0 3
rlabel polysilicon 201 -1709 201 -1709 0 2
rlabel polysilicon 208 -1709 208 -1709 0 2
rlabel polysilicon 215 -1709 215 -1709 0 2
rlabel polysilicon 212 -1715 212 -1715 0 3
rlabel polysilicon 215 -1715 215 -1715 0 4
rlabel polysilicon 219 -1709 219 -1709 0 1
rlabel polysilicon 219 -1715 219 -1715 0 3
rlabel polysilicon 226 -1709 226 -1709 0 1
rlabel polysilicon 226 -1715 226 -1715 0 3
rlabel polysilicon 233 -1709 233 -1709 0 1
rlabel polysilicon 233 -1715 233 -1715 0 3
rlabel polysilicon 240 -1709 240 -1709 0 1
rlabel polysilicon 240 -1715 240 -1715 0 3
rlabel polysilicon 254 -1709 254 -1709 0 1
rlabel polysilicon 254 -1715 254 -1715 0 3
rlabel polysilicon 264 -1709 264 -1709 0 2
rlabel polysilicon 261 -1715 261 -1715 0 3
rlabel polysilicon 268 -1709 268 -1709 0 1
rlabel polysilicon 268 -1715 268 -1715 0 3
rlabel polysilicon 275 -1709 275 -1709 0 1
rlabel polysilicon 278 -1715 278 -1715 0 4
rlabel polysilicon 282 -1709 282 -1709 0 1
rlabel polysilicon 282 -1715 282 -1715 0 3
rlabel polysilicon 289 -1709 289 -1709 0 1
rlabel polysilicon 289 -1715 289 -1715 0 3
rlabel polysilicon 296 -1715 296 -1715 0 3
rlabel polysilicon 299 -1715 299 -1715 0 4
rlabel polysilicon 303 -1709 303 -1709 0 1
rlabel polysilicon 303 -1715 303 -1715 0 3
rlabel polysilicon 310 -1709 310 -1709 0 1
rlabel polysilicon 310 -1715 310 -1715 0 3
rlabel polysilicon 317 -1709 317 -1709 0 1
rlabel polysilicon 317 -1715 317 -1715 0 3
rlabel polysilicon 324 -1709 324 -1709 0 1
rlabel polysilicon 324 -1715 324 -1715 0 3
rlabel polysilicon 331 -1709 331 -1709 0 1
rlabel polysilicon 331 -1715 331 -1715 0 3
rlabel polysilicon 341 -1709 341 -1709 0 2
rlabel polysilicon 338 -1715 338 -1715 0 3
rlabel polysilicon 345 -1709 345 -1709 0 1
rlabel polysilicon 345 -1715 345 -1715 0 3
rlabel polysilicon 355 -1709 355 -1709 0 2
rlabel polysilicon 352 -1715 352 -1715 0 3
rlabel polysilicon 359 -1709 359 -1709 0 1
rlabel polysilicon 359 -1715 359 -1715 0 3
rlabel polysilicon 366 -1709 366 -1709 0 1
rlabel polysilicon 366 -1715 366 -1715 0 3
rlabel polysilicon 373 -1709 373 -1709 0 1
rlabel polysilicon 376 -1709 376 -1709 0 2
rlabel polysilicon 373 -1715 373 -1715 0 3
rlabel polysilicon 383 -1709 383 -1709 0 2
rlabel polysilicon 383 -1715 383 -1715 0 4
rlabel polysilicon 387 -1709 387 -1709 0 1
rlabel polysilicon 394 -1709 394 -1709 0 1
rlabel polysilicon 394 -1715 394 -1715 0 3
rlabel polysilicon 404 -1709 404 -1709 0 2
rlabel polysilicon 401 -1715 401 -1715 0 3
rlabel polysilicon 408 -1709 408 -1709 0 1
rlabel polysilicon 408 -1715 408 -1715 0 3
rlabel polysilicon 415 -1709 415 -1709 0 1
rlabel polysilicon 415 -1715 415 -1715 0 3
rlabel polysilicon 422 -1709 422 -1709 0 1
rlabel polysilicon 425 -1709 425 -1709 0 2
rlabel polysilicon 422 -1715 422 -1715 0 3
rlabel polysilicon 429 -1709 429 -1709 0 1
rlabel polysilicon 429 -1715 429 -1715 0 3
rlabel polysilicon 436 -1709 436 -1709 0 1
rlabel polysilicon 436 -1715 436 -1715 0 3
rlabel polysilicon 443 -1709 443 -1709 0 1
rlabel polysilicon 443 -1715 443 -1715 0 3
rlabel polysilicon 450 -1709 450 -1709 0 1
rlabel polysilicon 450 -1715 450 -1715 0 3
rlabel polysilicon 457 -1709 457 -1709 0 1
rlabel polysilicon 457 -1715 457 -1715 0 3
rlabel polysilicon 464 -1709 464 -1709 0 1
rlabel polysilicon 464 -1715 464 -1715 0 3
rlabel polysilicon 474 -1709 474 -1709 0 2
rlabel polysilicon 471 -1715 471 -1715 0 3
rlabel polysilicon 478 -1709 478 -1709 0 1
rlabel polysilicon 478 -1715 478 -1715 0 3
rlabel polysilicon 485 -1709 485 -1709 0 1
rlabel polysilicon 485 -1715 485 -1715 0 3
rlabel polysilicon 492 -1709 492 -1709 0 1
rlabel polysilicon 492 -1715 492 -1715 0 3
rlabel polysilicon 499 -1715 499 -1715 0 3
rlabel polysilicon 506 -1709 506 -1709 0 1
rlabel polysilicon 506 -1715 506 -1715 0 3
rlabel polysilicon 513 -1709 513 -1709 0 1
rlabel polysilicon 513 -1715 513 -1715 0 3
rlabel polysilicon 520 -1709 520 -1709 0 1
rlabel polysilicon 520 -1715 520 -1715 0 3
rlabel polysilicon 527 -1709 527 -1709 0 1
rlabel polysilicon 527 -1715 527 -1715 0 3
rlabel polysilicon 534 -1709 534 -1709 0 1
rlabel polysilicon 534 -1715 534 -1715 0 3
rlabel polysilicon 541 -1709 541 -1709 0 1
rlabel polysilicon 541 -1715 541 -1715 0 3
rlabel polysilicon 548 -1709 548 -1709 0 1
rlabel polysilicon 548 -1715 548 -1715 0 3
rlabel polysilicon 555 -1709 555 -1709 0 1
rlabel polysilicon 555 -1715 555 -1715 0 3
rlabel polysilicon 562 -1709 562 -1709 0 1
rlabel polysilicon 562 -1715 562 -1715 0 3
rlabel polysilicon 569 -1709 569 -1709 0 1
rlabel polysilicon 569 -1715 569 -1715 0 3
rlabel polysilicon 576 -1709 576 -1709 0 1
rlabel polysilicon 576 -1715 576 -1715 0 3
rlabel polysilicon 583 -1709 583 -1709 0 1
rlabel polysilicon 583 -1715 583 -1715 0 3
rlabel polysilicon 590 -1709 590 -1709 0 1
rlabel polysilicon 593 -1709 593 -1709 0 2
rlabel polysilicon 593 -1715 593 -1715 0 4
rlabel polysilicon 597 -1715 597 -1715 0 3
rlabel polysilicon 604 -1709 604 -1709 0 1
rlabel polysilicon 604 -1715 604 -1715 0 3
rlabel polysilicon 611 -1709 611 -1709 0 1
rlabel polysilicon 611 -1715 611 -1715 0 3
rlabel polysilicon 618 -1709 618 -1709 0 1
rlabel polysilicon 618 -1715 618 -1715 0 3
rlabel polysilicon 639 -1709 639 -1709 0 1
rlabel polysilicon 639 -1715 639 -1715 0 3
rlabel polysilicon 646 -1709 646 -1709 0 1
rlabel polysilicon 646 -1715 646 -1715 0 3
rlabel polysilicon 653 -1709 653 -1709 0 1
rlabel polysilicon 653 -1715 653 -1715 0 3
rlabel polysilicon 674 -1709 674 -1709 0 1
rlabel polysilicon 674 -1715 674 -1715 0 3
rlabel polysilicon 681 -1715 681 -1715 0 3
rlabel polysilicon 709 -1709 709 -1709 0 1
rlabel polysilicon 709 -1715 709 -1715 0 3
rlabel polysilicon 723 -1709 723 -1709 0 1
rlabel polysilicon 723 -1715 723 -1715 0 3
rlabel polysilicon 730 -1709 730 -1709 0 1
rlabel polysilicon 730 -1715 730 -1715 0 3
rlabel polysilicon 737 -1709 737 -1709 0 1
rlabel polysilicon 737 -1715 737 -1715 0 3
rlabel polysilicon 744 -1709 744 -1709 0 1
rlabel polysilicon 744 -1715 744 -1715 0 3
rlabel polysilicon 751 -1709 751 -1709 0 1
rlabel polysilicon 751 -1715 751 -1715 0 3
rlabel polysilicon 758 -1709 758 -1709 0 1
rlabel polysilicon 758 -1715 758 -1715 0 3
rlabel polysilicon 765 -1709 765 -1709 0 1
rlabel polysilicon 765 -1715 765 -1715 0 3
rlabel polysilicon 772 -1709 772 -1709 0 1
rlabel polysilicon 772 -1715 772 -1715 0 3
rlabel polysilicon 779 -1709 779 -1709 0 1
rlabel polysilicon 779 -1715 779 -1715 0 3
rlabel polysilicon 793 -1709 793 -1709 0 1
rlabel polysilicon 793 -1715 793 -1715 0 3
rlabel polysilicon 796 -1715 796 -1715 0 4
rlabel polysilicon 800 -1709 800 -1709 0 1
rlabel polysilicon 800 -1715 800 -1715 0 3
rlabel polysilicon 807 -1709 807 -1709 0 1
rlabel polysilicon 807 -1715 807 -1715 0 3
rlabel polysilicon 817 -1709 817 -1709 0 2
rlabel polysilicon 821 -1709 821 -1709 0 1
rlabel polysilicon 821 -1715 821 -1715 0 3
rlabel polysilicon 828 -1709 828 -1709 0 1
rlabel polysilicon 828 -1715 828 -1715 0 3
rlabel polysilicon 835 -1709 835 -1709 0 1
rlabel polysilicon 835 -1715 835 -1715 0 3
rlabel polysilicon 845 -1715 845 -1715 0 4
rlabel polysilicon 849 -1709 849 -1709 0 1
rlabel polysilicon 849 -1715 849 -1715 0 3
rlabel polysilicon 856 -1709 856 -1709 0 1
rlabel polysilicon 856 -1715 856 -1715 0 3
rlabel polysilicon 863 -1709 863 -1709 0 1
rlabel polysilicon 866 -1709 866 -1709 0 2
rlabel polysilicon 866 -1715 866 -1715 0 4
rlabel polysilicon 884 -1709 884 -1709 0 1
rlabel polysilicon 884 -1715 884 -1715 0 3
rlabel polysilicon 898 -1709 898 -1709 0 1
rlabel polysilicon 898 -1715 898 -1715 0 3
rlabel polysilicon 968 -1709 968 -1709 0 1
rlabel polysilicon 968 -1715 968 -1715 0 3
rlabel polysilicon 1024 -1709 1024 -1709 0 1
rlabel polysilicon 1024 -1715 1024 -1715 0 3
rlabel polysilicon 44 -1742 44 -1742 0 1
rlabel polysilicon 44 -1748 44 -1748 0 3
rlabel polysilicon 61 -1748 61 -1748 0 4
rlabel polysilicon 65 -1742 65 -1742 0 1
rlabel polysilicon 65 -1748 65 -1748 0 3
rlabel polysilicon 100 -1742 100 -1742 0 1
rlabel polysilicon 100 -1748 100 -1748 0 3
rlabel polysilicon 107 -1742 107 -1742 0 1
rlabel polysilicon 107 -1748 107 -1748 0 3
rlabel polysilicon 114 -1742 114 -1742 0 1
rlabel polysilicon 121 -1742 121 -1742 0 1
rlabel polysilicon 121 -1748 121 -1748 0 3
rlabel polysilicon 128 -1748 128 -1748 0 3
rlabel polysilicon 131 -1748 131 -1748 0 4
rlabel polysilicon 135 -1748 135 -1748 0 3
rlabel polysilicon 138 -1748 138 -1748 0 4
rlabel polysilicon 142 -1742 142 -1742 0 1
rlabel polysilicon 145 -1742 145 -1742 0 2
rlabel polysilicon 142 -1748 142 -1748 0 3
rlabel polysilicon 145 -1748 145 -1748 0 4
rlabel polysilicon 152 -1742 152 -1742 0 2
rlabel polysilicon 156 -1742 156 -1742 0 1
rlabel polysilicon 156 -1748 156 -1748 0 3
rlabel polysilicon 159 -1748 159 -1748 0 4
rlabel polysilicon 163 -1742 163 -1742 0 1
rlabel polysilicon 163 -1748 163 -1748 0 3
rlabel polysilicon 170 -1748 170 -1748 0 3
rlabel polysilicon 173 -1748 173 -1748 0 4
rlabel polysilicon 177 -1742 177 -1742 0 1
rlabel polysilicon 177 -1748 177 -1748 0 3
rlabel polysilicon 184 -1742 184 -1742 0 1
rlabel polysilicon 184 -1748 184 -1748 0 3
rlabel polysilicon 191 -1742 191 -1742 0 1
rlabel polysilicon 191 -1748 191 -1748 0 3
rlabel polysilicon 205 -1742 205 -1742 0 1
rlabel polysilicon 205 -1748 205 -1748 0 3
rlabel polysilicon 212 -1742 212 -1742 0 1
rlabel polysilicon 219 -1748 219 -1748 0 3
rlabel polysilicon 226 -1742 226 -1742 0 1
rlabel polysilicon 233 -1742 233 -1742 0 1
rlabel polysilicon 233 -1748 233 -1748 0 3
rlabel polysilicon 240 -1742 240 -1742 0 1
rlabel polysilicon 240 -1748 240 -1748 0 3
rlabel polysilicon 247 -1742 247 -1742 0 1
rlabel polysilicon 247 -1748 247 -1748 0 3
rlabel polysilicon 275 -1742 275 -1742 0 1
rlabel polysilicon 275 -1748 275 -1748 0 3
rlabel polysilicon 296 -1742 296 -1742 0 1
rlabel polysilicon 296 -1748 296 -1748 0 3
rlabel polysilicon 303 -1742 303 -1742 0 1
rlabel polysilicon 303 -1748 303 -1748 0 3
rlabel polysilicon 310 -1742 310 -1742 0 1
rlabel polysilicon 310 -1748 310 -1748 0 3
rlabel polysilicon 317 -1742 317 -1742 0 1
rlabel polysilicon 317 -1748 317 -1748 0 3
rlabel polysilicon 324 -1742 324 -1742 0 1
rlabel polysilicon 324 -1748 324 -1748 0 3
rlabel polysilicon 331 -1742 331 -1742 0 1
rlabel polysilicon 331 -1748 331 -1748 0 3
rlabel polysilicon 338 -1742 338 -1742 0 1
rlabel polysilicon 338 -1748 338 -1748 0 3
rlabel polysilicon 345 -1742 345 -1742 0 1
rlabel polysilicon 345 -1748 345 -1748 0 3
rlabel polysilicon 352 -1742 352 -1742 0 1
rlabel polysilicon 352 -1748 352 -1748 0 3
rlabel polysilicon 359 -1742 359 -1742 0 1
rlabel polysilicon 359 -1748 359 -1748 0 3
rlabel polysilicon 366 -1742 366 -1742 0 1
rlabel polysilicon 369 -1742 369 -1742 0 2
rlabel polysilicon 366 -1748 366 -1748 0 3
rlabel polysilicon 373 -1742 373 -1742 0 1
rlabel polysilicon 373 -1748 373 -1748 0 3
rlabel polysilicon 380 -1742 380 -1742 0 1
rlabel polysilicon 380 -1748 380 -1748 0 3
rlabel polysilicon 387 -1748 387 -1748 0 3
rlabel polysilicon 394 -1742 394 -1742 0 1
rlabel polysilicon 394 -1748 394 -1748 0 3
rlabel polysilicon 404 -1748 404 -1748 0 4
rlabel polysilicon 411 -1742 411 -1742 0 2
rlabel polysilicon 411 -1748 411 -1748 0 4
rlabel polysilicon 415 -1742 415 -1742 0 1
rlabel polysilicon 415 -1748 415 -1748 0 3
rlabel polysilicon 422 -1742 422 -1742 0 1
rlabel polysilicon 422 -1748 422 -1748 0 3
rlabel polysilicon 429 -1742 429 -1742 0 1
rlabel polysilicon 429 -1748 429 -1748 0 3
rlabel polysilicon 436 -1742 436 -1742 0 1
rlabel polysilicon 436 -1748 436 -1748 0 3
rlabel polysilicon 446 -1742 446 -1742 0 2
rlabel polysilicon 450 -1742 450 -1742 0 1
rlabel polysilicon 450 -1748 450 -1748 0 3
rlabel polysilicon 457 -1742 457 -1742 0 1
rlabel polysilicon 457 -1748 457 -1748 0 3
rlabel polysilicon 464 -1742 464 -1742 0 1
rlabel polysilicon 464 -1748 464 -1748 0 3
rlabel polysilicon 471 -1748 471 -1748 0 3
rlabel polysilicon 478 -1742 478 -1742 0 1
rlabel polysilicon 478 -1748 478 -1748 0 3
rlabel polysilicon 485 -1742 485 -1742 0 1
rlabel polysilicon 488 -1748 488 -1748 0 4
rlabel polysilicon 492 -1742 492 -1742 0 1
rlabel polysilicon 492 -1748 492 -1748 0 3
rlabel polysilicon 499 -1742 499 -1742 0 1
rlabel polysilicon 499 -1748 499 -1748 0 3
rlabel polysilicon 506 -1748 506 -1748 0 3
rlabel polysilicon 509 -1748 509 -1748 0 4
rlabel polysilicon 513 -1742 513 -1742 0 1
rlabel polysilicon 513 -1748 513 -1748 0 3
rlabel polysilicon 520 -1742 520 -1742 0 1
rlabel polysilicon 520 -1748 520 -1748 0 3
rlabel polysilicon 530 -1748 530 -1748 0 4
rlabel polysilicon 534 -1742 534 -1742 0 1
rlabel polysilicon 534 -1748 534 -1748 0 3
rlabel polysilicon 541 -1742 541 -1742 0 1
rlabel polysilicon 541 -1748 541 -1748 0 3
rlabel polysilicon 548 -1742 548 -1742 0 1
rlabel polysilicon 548 -1748 548 -1748 0 3
rlabel polysilicon 555 -1742 555 -1742 0 1
rlabel polysilicon 555 -1748 555 -1748 0 3
rlabel polysilicon 562 -1748 562 -1748 0 3
rlabel polysilicon 569 -1742 569 -1742 0 1
rlabel polysilicon 569 -1748 569 -1748 0 3
rlabel polysilicon 576 -1742 576 -1742 0 1
rlabel polysilicon 576 -1748 576 -1748 0 3
rlabel polysilicon 586 -1748 586 -1748 0 4
rlabel polysilicon 590 -1742 590 -1742 0 1
rlabel polysilicon 590 -1748 590 -1748 0 3
rlabel polysilicon 597 -1742 597 -1742 0 1
rlabel polysilicon 597 -1748 597 -1748 0 3
rlabel polysilicon 646 -1742 646 -1742 0 1
rlabel polysilicon 646 -1748 646 -1748 0 3
rlabel polysilicon 656 -1742 656 -1742 0 2
rlabel polysilicon 656 -1748 656 -1748 0 4
rlabel polysilicon 702 -1742 702 -1742 0 1
rlabel polysilicon 702 -1748 702 -1748 0 3
rlabel polysilicon 709 -1742 709 -1742 0 1
rlabel polysilicon 709 -1748 709 -1748 0 3
rlabel polysilicon 716 -1748 716 -1748 0 3
rlabel polysilicon 723 -1742 723 -1742 0 1
rlabel polysilicon 723 -1748 723 -1748 0 3
rlabel polysilicon 730 -1742 730 -1742 0 1
rlabel polysilicon 730 -1748 730 -1748 0 3
rlabel polysilicon 737 -1742 737 -1742 0 1
rlabel polysilicon 737 -1748 737 -1748 0 3
rlabel polysilicon 744 -1742 744 -1742 0 1
rlabel polysilicon 744 -1748 744 -1748 0 3
rlabel polysilicon 751 -1742 751 -1742 0 1
rlabel polysilicon 751 -1748 751 -1748 0 3
rlabel polysilicon 758 -1742 758 -1742 0 1
rlabel polysilicon 758 -1748 758 -1748 0 3
rlabel polysilicon 765 -1742 765 -1742 0 1
rlabel polysilicon 765 -1748 765 -1748 0 3
rlabel polysilicon 772 -1748 772 -1748 0 3
rlabel polysilicon 782 -1742 782 -1742 0 2
rlabel polysilicon 779 -1748 779 -1748 0 3
rlabel polysilicon 782 -1748 782 -1748 0 4
rlabel polysilicon 786 -1742 786 -1742 0 1
rlabel polysilicon 786 -1748 786 -1748 0 3
rlabel polysilicon 793 -1742 793 -1742 0 1
rlabel polysilicon 796 -1742 796 -1742 0 2
rlabel polysilicon 793 -1748 793 -1748 0 3
rlabel polysilicon 800 -1742 800 -1742 0 1
rlabel polysilicon 800 -1748 800 -1748 0 3
rlabel polysilicon 807 -1742 807 -1742 0 1
rlabel polysilicon 807 -1748 807 -1748 0 3
rlabel polysilicon 828 -1742 828 -1742 0 1
rlabel polysilicon 828 -1748 828 -1748 0 3
rlabel polysilicon 842 -1742 842 -1742 0 1
rlabel polysilicon 842 -1748 842 -1748 0 3
rlabel polysilicon 856 -1742 856 -1742 0 1
rlabel polysilicon 856 -1748 856 -1748 0 3
rlabel polysilicon 884 -1742 884 -1742 0 1
rlabel polysilicon 884 -1748 884 -1748 0 3
rlabel polysilicon 898 -1742 898 -1742 0 1
rlabel polysilicon 898 -1748 898 -1748 0 3
rlabel polysilicon 968 -1742 968 -1742 0 1
rlabel polysilicon 968 -1748 968 -1748 0 3
rlabel polysilicon 975 -1748 975 -1748 0 3
rlabel polysilicon 1024 -1742 1024 -1742 0 1
rlabel polysilicon 1024 -1748 1024 -1748 0 3
rlabel polysilicon 47 -1769 47 -1769 0 2
rlabel polysilicon 58 -1769 58 -1769 0 1
rlabel polysilicon 58 -1775 58 -1775 0 3
rlabel polysilicon 65 -1769 65 -1769 0 1
rlabel polysilicon 65 -1775 65 -1775 0 3
rlabel polysilicon 72 -1769 72 -1769 0 1
rlabel polysilicon 72 -1775 72 -1775 0 3
rlabel polysilicon 79 -1769 79 -1769 0 1
rlabel polysilicon 79 -1775 79 -1775 0 3
rlabel polysilicon 93 -1769 93 -1769 0 1
rlabel polysilicon 93 -1775 93 -1775 0 3
rlabel polysilicon 100 -1769 100 -1769 0 1
rlabel polysilicon 110 -1775 110 -1775 0 4
rlabel polysilicon 117 -1769 117 -1769 0 2
rlabel polysilicon 117 -1775 117 -1775 0 4
rlabel polysilicon 121 -1769 121 -1769 0 1
rlabel polysilicon 128 -1769 128 -1769 0 1
rlabel polysilicon 128 -1775 128 -1775 0 3
rlabel polysilicon 135 -1769 135 -1769 0 1
rlabel polysilicon 135 -1775 135 -1775 0 3
rlabel polysilicon 142 -1769 142 -1769 0 1
rlabel polysilicon 142 -1775 142 -1775 0 3
rlabel polysilicon 152 -1775 152 -1775 0 4
rlabel polysilicon 156 -1769 156 -1769 0 1
rlabel polysilicon 170 -1769 170 -1769 0 1
rlabel polysilicon 170 -1775 170 -1775 0 3
rlabel polysilicon 191 -1769 191 -1769 0 1
rlabel polysilicon 191 -1775 191 -1775 0 3
rlabel polysilicon 198 -1775 198 -1775 0 3
rlabel polysilicon 205 -1769 205 -1769 0 1
rlabel polysilicon 205 -1775 205 -1775 0 3
rlabel polysilicon 212 -1769 212 -1769 0 1
rlabel polysilicon 219 -1769 219 -1769 0 1
rlabel polysilicon 219 -1775 219 -1775 0 3
rlabel polysilicon 229 -1769 229 -1769 0 2
rlabel polysilicon 226 -1775 226 -1775 0 3
rlabel polysilicon 233 -1769 233 -1769 0 1
rlabel polysilicon 233 -1775 233 -1775 0 3
rlabel polysilicon 240 -1769 240 -1769 0 1
rlabel polysilicon 240 -1775 240 -1775 0 3
rlabel polysilicon 275 -1769 275 -1769 0 1
rlabel polysilicon 275 -1775 275 -1775 0 3
rlabel polysilicon 282 -1769 282 -1769 0 1
rlabel polysilicon 282 -1775 282 -1775 0 3
rlabel polysilicon 289 -1769 289 -1769 0 1
rlabel polysilicon 289 -1775 289 -1775 0 3
rlabel polysilicon 296 -1769 296 -1769 0 1
rlabel polysilicon 296 -1775 296 -1775 0 3
rlabel polysilicon 306 -1775 306 -1775 0 4
rlabel polysilicon 310 -1769 310 -1769 0 1
rlabel polysilicon 310 -1775 310 -1775 0 3
rlabel polysilicon 317 -1769 317 -1769 0 1
rlabel polysilicon 324 -1769 324 -1769 0 1
rlabel polysilicon 324 -1775 324 -1775 0 3
rlabel polysilicon 331 -1775 331 -1775 0 3
rlabel polysilicon 338 -1769 338 -1769 0 1
rlabel polysilicon 338 -1775 338 -1775 0 3
rlabel polysilicon 345 -1769 345 -1769 0 1
rlabel polysilicon 345 -1775 345 -1775 0 3
rlabel polysilicon 352 -1769 352 -1769 0 1
rlabel polysilicon 352 -1775 352 -1775 0 3
rlabel polysilicon 359 -1769 359 -1769 0 1
rlabel polysilicon 362 -1775 362 -1775 0 4
rlabel polysilicon 369 -1769 369 -1769 0 2
rlabel polysilicon 373 -1769 373 -1769 0 1
rlabel polysilicon 373 -1775 373 -1775 0 3
rlabel polysilicon 380 -1769 380 -1769 0 1
rlabel polysilicon 380 -1775 380 -1775 0 3
rlabel polysilicon 394 -1769 394 -1769 0 1
rlabel polysilicon 394 -1775 394 -1775 0 3
rlabel polysilicon 401 -1769 401 -1769 0 1
rlabel polysilicon 401 -1775 401 -1775 0 3
rlabel polysilicon 411 -1775 411 -1775 0 4
rlabel polysilicon 415 -1769 415 -1769 0 1
rlabel polysilicon 415 -1775 415 -1775 0 3
rlabel polysilicon 422 -1769 422 -1769 0 1
rlabel polysilicon 429 -1769 429 -1769 0 1
rlabel polysilicon 443 -1769 443 -1769 0 1
rlabel polysilicon 443 -1775 443 -1775 0 3
rlabel polysilicon 450 -1769 450 -1769 0 1
rlabel polysilicon 450 -1775 450 -1775 0 3
rlabel polysilicon 457 -1769 457 -1769 0 1
rlabel polysilicon 457 -1775 457 -1775 0 3
rlabel polysilicon 464 -1769 464 -1769 0 1
rlabel polysilicon 464 -1775 464 -1775 0 3
rlabel polysilicon 471 -1769 471 -1769 0 1
rlabel polysilicon 471 -1775 471 -1775 0 3
rlabel polysilicon 478 -1769 478 -1769 0 1
rlabel polysilicon 478 -1775 478 -1775 0 3
rlabel polysilicon 506 -1769 506 -1769 0 1
rlabel polysilicon 506 -1775 506 -1775 0 3
rlabel polysilicon 513 -1769 513 -1769 0 1
rlabel polysilicon 513 -1775 513 -1775 0 3
rlabel polysilicon 527 -1769 527 -1769 0 1
rlabel polysilicon 527 -1775 527 -1775 0 3
rlabel polysilicon 562 -1769 562 -1769 0 1
rlabel polysilicon 562 -1775 562 -1775 0 3
rlabel polysilicon 709 -1769 709 -1769 0 1
rlabel polysilicon 709 -1775 709 -1775 0 3
rlabel polysilicon 716 -1775 716 -1775 0 3
rlabel polysilicon 723 -1769 723 -1769 0 1
rlabel polysilicon 723 -1775 723 -1775 0 3
rlabel polysilicon 730 -1769 730 -1769 0 1
rlabel polysilicon 730 -1775 730 -1775 0 3
rlabel polysilicon 737 -1769 737 -1769 0 1
rlabel polysilicon 737 -1775 737 -1775 0 3
rlabel polysilicon 747 -1775 747 -1775 0 4
rlabel polysilicon 751 -1769 751 -1769 0 1
rlabel polysilicon 751 -1775 751 -1775 0 3
rlabel polysilicon 758 -1769 758 -1769 0 1
rlabel polysilicon 758 -1775 758 -1775 0 3
rlabel polysilicon 772 -1769 772 -1769 0 1
rlabel polysilicon 772 -1775 772 -1775 0 3
rlabel polysilicon 779 -1775 779 -1775 0 3
rlabel polysilicon 793 -1769 793 -1769 0 1
rlabel polysilicon 793 -1775 793 -1775 0 3
rlabel polysilicon 814 -1769 814 -1769 0 1
rlabel polysilicon 814 -1775 814 -1775 0 3
rlabel polysilicon 828 -1769 828 -1769 0 1
rlabel polysilicon 828 -1775 828 -1775 0 3
rlabel polysilicon 845 -1769 845 -1769 0 2
rlabel polysilicon 856 -1769 856 -1769 0 1
rlabel polysilicon 880 -1775 880 -1775 0 4
rlabel polysilicon 884 -1769 884 -1769 0 1
rlabel polysilicon 884 -1775 884 -1775 0 3
rlabel polysilicon 898 -1769 898 -1769 0 1
rlabel polysilicon 898 -1775 898 -1775 0 3
rlabel polysilicon 1024 -1769 1024 -1769 0 1
rlabel polysilicon 1024 -1775 1024 -1775 0 3
rlabel polysilicon 68 -1796 68 -1796 0 4
rlabel polysilicon 75 -1790 75 -1790 0 2
rlabel polysilicon 79 -1790 79 -1790 0 1
rlabel polysilicon 79 -1796 79 -1796 0 3
rlabel polysilicon 142 -1790 142 -1790 0 1
rlabel polysilicon 142 -1796 142 -1796 0 3
rlabel polysilicon 152 -1790 152 -1790 0 2
rlabel polysilicon 149 -1796 149 -1796 0 3
rlabel polysilicon 156 -1790 156 -1790 0 1
rlabel polysilicon 156 -1796 156 -1796 0 3
rlabel polysilicon 173 -1790 173 -1790 0 2
rlabel polysilicon 184 -1796 184 -1796 0 3
rlabel polysilicon 205 -1790 205 -1790 0 1
rlabel polysilicon 205 -1796 205 -1796 0 3
rlabel polysilicon 226 -1790 226 -1790 0 1
rlabel polysilicon 226 -1796 226 -1796 0 3
rlabel polysilicon 240 -1790 240 -1790 0 1
rlabel polysilicon 240 -1796 240 -1796 0 3
rlabel polysilicon 247 -1790 247 -1790 0 1
rlabel polysilicon 247 -1796 247 -1796 0 3
rlabel polysilicon 261 -1790 261 -1790 0 1
rlabel polysilicon 261 -1796 261 -1796 0 3
rlabel polysilicon 282 -1790 282 -1790 0 1
rlabel polysilicon 282 -1796 282 -1796 0 3
rlabel polysilicon 296 -1790 296 -1790 0 1
rlabel polysilicon 296 -1796 296 -1796 0 3
rlabel polysilicon 303 -1790 303 -1790 0 1
rlabel polysilicon 306 -1790 306 -1790 0 2
rlabel polysilicon 313 -1790 313 -1790 0 2
rlabel polysilicon 320 -1790 320 -1790 0 2
rlabel polysilicon 324 -1790 324 -1790 0 1
rlabel polysilicon 324 -1796 324 -1796 0 3
rlabel polysilicon 331 -1790 331 -1790 0 1
rlabel polysilicon 331 -1796 331 -1796 0 3
rlabel polysilicon 338 -1790 338 -1790 0 1
rlabel polysilicon 338 -1796 338 -1796 0 3
rlabel polysilicon 345 -1796 345 -1796 0 3
rlabel polysilicon 352 -1790 352 -1790 0 1
rlabel polysilicon 352 -1796 352 -1796 0 3
rlabel polysilicon 380 -1790 380 -1790 0 1
rlabel polysilicon 380 -1796 380 -1796 0 3
rlabel polysilicon 387 -1790 387 -1790 0 1
rlabel polysilicon 387 -1796 387 -1796 0 3
rlabel polysilicon 411 -1790 411 -1790 0 2
rlabel polysilicon 415 -1790 415 -1790 0 1
rlabel polysilicon 415 -1796 415 -1796 0 3
rlabel polysilicon 422 -1790 422 -1790 0 1
rlabel polysilicon 422 -1796 422 -1796 0 3
rlabel polysilicon 429 -1796 429 -1796 0 3
rlabel polysilicon 432 -1796 432 -1796 0 4
rlabel polysilicon 439 -1796 439 -1796 0 4
rlabel polysilicon 443 -1790 443 -1790 0 1
rlabel polysilicon 443 -1796 443 -1796 0 3
rlabel polysilicon 450 -1790 450 -1790 0 1
rlabel polysilicon 450 -1796 450 -1796 0 3
rlabel polysilicon 457 -1790 457 -1790 0 1
rlabel polysilicon 457 -1796 457 -1796 0 3
rlabel polysilicon 471 -1790 471 -1790 0 1
rlabel polysilicon 471 -1796 471 -1796 0 3
rlabel polysilicon 478 -1790 478 -1790 0 1
rlabel polysilicon 478 -1796 478 -1796 0 3
rlabel polysilicon 502 -1790 502 -1790 0 2
rlabel polysilicon 506 -1796 506 -1796 0 3
rlabel polysilicon 513 -1790 513 -1790 0 1
rlabel polysilicon 513 -1796 513 -1796 0 3
rlabel polysilicon 520 -1790 520 -1790 0 1
rlabel polysilicon 520 -1796 520 -1796 0 3
rlabel polysilicon 565 -1790 565 -1790 0 2
rlabel polysilicon 737 -1790 737 -1790 0 1
rlabel polysilicon 737 -1796 737 -1796 0 3
rlabel polysilicon 744 -1796 744 -1796 0 3
rlabel polysilicon 754 -1796 754 -1796 0 4
rlabel polysilicon 758 -1790 758 -1790 0 1
rlabel polysilicon 758 -1796 758 -1796 0 3
rlabel polysilicon 765 -1790 765 -1790 0 1
rlabel polysilicon 765 -1796 765 -1796 0 3
rlabel polysilicon 772 -1790 772 -1790 0 1
rlabel polysilicon 793 -1790 793 -1790 0 1
rlabel polysilicon 793 -1796 793 -1796 0 3
rlabel polysilicon 814 -1790 814 -1790 0 1
rlabel polysilicon 838 -1790 838 -1790 0 2
rlabel polysilicon 898 -1790 898 -1790 0 1
rlabel polysilicon 898 -1796 898 -1796 0 3
rlabel polysilicon 1024 -1790 1024 -1790 0 1
rlabel polysilicon 1024 -1796 1024 -1796 0 3
rlabel polysilicon 159 -1805 159 -1805 0 2
rlabel polysilicon 187 -1811 187 -1811 0 4
rlabel polysilicon 191 -1805 191 -1805 0 1
rlabel polysilicon 191 -1811 191 -1811 0 3
rlabel polysilicon 208 -1805 208 -1805 0 2
rlabel polysilicon 222 -1811 222 -1811 0 4
rlabel polysilicon 226 -1805 226 -1805 0 1
rlabel polysilicon 226 -1811 226 -1811 0 3
rlabel polysilicon 264 -1811 264 -1811 0 4
rlabel polysilicon 268 -1805 268 -1805 0 1
rlabel polysilicon 268 -1811 268 -1811 0 3
rlabel polysilicon 282 -1805 282 -1805 0 1
rlabel polysilicon 296 -1805 296 -1805 0 1
rlabel polysilicon 296 -1811 296 -1811 0 3
rlabel polysilicon 306 -1811 306 -1811 0 4
rlabel polysilicon 324 -1811 324 -1811 0 3
rlabel polysilicon 331 -1805 331 -1805 0 1
rlabel polysilicon 331 -1811 331 -1811 0 3
rlabel polysilicon 341 -1805 341 -1805 0 2
rlabel polysilicon 352 -1805 352 -1805 0 1
rlabel polysilicon 352 -1811 352 -1811 0 3
rlabel polysilicon 359 -1811 359 -1811 0 3
rlabel polysilicon 376 -1811 376 -1811 0 4
rlabel polysilicon 383 -1805 383 -1805 0 2
rlabel polysilicon 387 -1805 387 -1805 0 1
rlabel polysilicon 387 -1811 387 -1811 0 3
rlabel polysilicon 422 -1805 422 -1805 0 1
rlabel polysilicon 422 -1811 422 -1811 0 3
rlabel polysilicon 429 -1811 429 -1811 0 3
rlabel polysilicon 464 -1805 464 -1805 0 1
rlabel polysilicon 471 -1805 471 -1805 0 1
rlabel polysilicon 481 -1805 481 -1805 0 2
rlabel polysilicon 516 -1805 516 -1805 0 2
rlabel polysilicon 747 -1811 747 -1811 0 4
rlabel polysilicon 751 -1805 751 -1805 0 1
rlabel polysilicon 751 -1811 751 -1811 0 3
rlabel polysilicon 796 -1805 796 -1805 0 2
rlabel polysilicon 901 -1811 901 -1811 0 4
rlabel polysilicon 905 -1805 905 -1805 0 1
rlabel polysilicon 905 -1811 905 -1811 0 3
rlabel polysilicon 1027 -1805 1027 -1805 0 2
rlabel metal2 177 1 177 1 0 net=3759
rlabel metal2 212 1 212 1 0 net=1983
rlabel metal2 236 1 236 1 0 net=4005
rlabel metal2 254 1 254 1 0 net=4861
rlabel metal2 285 1 285 1 0 net=2189
rlabel metal2 303 1 303 1 0 net=2651
rlabel metal2 338 1 338 1 0 net=3731
rlabel metal2 352 1 352 1 0 net=2855
rlabel metal2 366 1 366 1 0 net=2823
rlabel metal2 467 1 467 1 0 net=6401
rlabel metal2 478 1 478 1 0 net=6075
rlabel metal2 534 1 534 1 0 net=5113
rlabel metal2 576 1 576 1 0 net=6097
rlabel metal2 604 1 604 1 0 net=5489
rlabel metal2 730 1 730 1 0 net=6029
rlabel metal2 184 -1 184 -1 0 net=2045
rlabel metal2 114 -12 114 -12 0 net=1663
rlabel metal2 156 -12 156 -12 0 net=1453
rlabel metal2 170 -12 170 -12 0 net=3761
rlabel metal2 184 -12 184 -12 0 net=2047
rlabel metal2 184 -12 184 -12 0 net=2047
rlabel metal2 219 -12 219 -12 0 net=1985
rlabel metal2 240 -12 240 -12 0 net=4007
rlabel metal2 278 -12 278 -12 0 net=1037
rlabel metal2 296 -12 296 -12 0 net=1955
rlabel metal2 296 -12 296 -12 0 net=1955
rlabel metal2 303 -12 303 -12 0 net=2653
rlabel metal2 317 -12 317 -12 0 net=3233
rlabel metal2 317 -12 317 -12 0 net=3233
rlabel metal2 345 -12 345 -12 0 net=2825
rlabel metal2 408 -12 408 -12 0 net=5725
rlabel metal2 450 -12 450 -12 0 net=3021
rlabel metal2 474 -12 474 -12 0 net=5389
rlabel metal2 485 -12 485 -12 0 net=6077
rlabel metal2 527 -12 527 -12 0 net=3335
rlabel metal2 583 -12 583 -12 0 net=6099
rlabel metal2 583 -12 583 -12 0 net=6099
rlabel metal2 604 -12 604 -12 0 net=5491
rlabel metal2 618 -12 618 -12 0 net=5793
rlabel metal2 688 -12 688 -12 0 net=6331
rlabel metal2 730 -12 730 -12 0 net=6031
rlabel metal2 730 -12 730 -12 0 net=6031
rlabel metal2 215 -14 215 -14 0 net=995
rlabel metal2 247 -14 247 -14 0 net=4863
rlabel metal2 289 -14 289 -14 0 net=2191
rlabel metal2 352 -14 352 -14 0 net=2857
rlabel metal2 366 -14 366 -14 0 net=2437
rlabel metal2 415 -14 415 -14 0 net=2615
rlabel metal2 425 -14 425 -14 0 net=4011
rlabel metal2 457 -14 457 -14 0 net=3065
rlabel metal2 471 -14 471 -14 0 net=6403
rlabel metal2 541 -14 541 -14 0 net=5115
rlabel metal2 541 -14 541 -14 0 net=5115
rlabel metal2 555 -14 555 -14 0 net=4177
rlabel metal2 240 -16 240 -16 0 net=1071
rlabel metal2 278 -16 278 -16 0 net=1735
rlabel metal2 338 -16 338 -16 0 net=3733
rlabel metal2 334 -18 334 -18 0 net=4147
rlabel metal2 58 -29 58 -29 0 net=841
rlabel metal2 79 -29 79 -29 0 net=5443
rlabel metal2 79 -29 79 -29 0 net=5443
rlabel metal2 114 -29 114 -29 0 net=1249
rlabel metal2 128 -29 128 -29 0 net=545
rlabel metal2 128 -29 128 -29 0 net=545
rlabel metal2 142 -29 142 -29 0 net=3763
rlabel metal2 184 -29 184 -29 0 net=2049
rlabel metal2 212 -29 212 -29 0 net=997
rlabel metal2 226 -29 226 -29 0 net=1987
rlabel metal2 268 -29 268 -29 0 net=1957
rlabel metal2 317 -29 317 -29 0 net=3235
rlabel metal2 334 -29 334 -29 0 net=2826
rlabel metal2 352 -29 352 -29 0 net=3735
rlabel metal2 380 -29 380 -29 0 net=5445
rlabel metal2 380 -29 380 -29 0 net=5445
rlabel metal2 387 -29 387 -29 0 net=2281
rlabel metal2 408 -29 408 -29 0 net=2827
rlabel metal2 415 -29 415 -29 0 net=2616
rlabel metal2 429 -29 429 -29 0 net=4013
rlabel metal2 443 -29 443 -29 0 net=5727
rlabel metal2 478 -29 478 -29 0 net=5391
rlabel metal2 478 -29 478 -29 0 net=5391
rlabel metal2 485 -29 485 -29 0 net=6405
rlabel metal2 485 -29 485 -29 0 net=6405
rlabel metal2 492 -29 492 -29 0 net=6079
rlabel metal2 513 -29 513 -29 0 net=5971
rlabel metal2 541 -29 541 -29 0 net=5117
rlabel metal2 576 -29 576 -29 0 net=5037
rlabel metal2 583 -29 583 -29 0 net=6101
rlabel metal2 604 -29 604 -29 0 net=4179
rlabel metal2 646 -29 646 -29 0 net=4233
rlabel metal2 688 -29 688 -29 0 net=6333
rlabel metal2 688 -29 688 -29 0 net=6333
rlabel metal2 709 -29 709 -29 0 net=5309
rlabel metal2 807 -29 807 -29 0 net=4865
rlabel metal2 121 -31 121 -31 0 net=1665
rlabel metal2 152 -31 152 -31 0 net=1689
rlabel metal2 163 -31 163 -31 0 net=1454
rlabel metal2 177 -31 177 -31 0 net=1653
rlabel metal2 233 -31 233 -31 0 net=1073
rlabel metal2 254 -31 254 -31 0 net=4009
rlabel metal2 345 -31 345 -31 0 net=2439
rlabel metal2 429 -31 429 -31 0 net=6675
rlabel metal2 450 -31 450 -31 0 net=3023
rlabel metal2 450 -31 450 -31 0 net=3023
rlabel metal2 457 -31 457 -31 0 net=3067
rlabel metal2 457 -31 457 -31 0 net=3067
rlabel metal2 527 -31 527 -31 0 net=3337
rlabel metal2 572 -31 572 -31 0 net=4561
rlabel metal2 604 -31 604 -31 0 net=5493
rlabel metal2 625 -31 625 -31 0 net=5869
rlabel metal2 730 -31 730 -31 0 net=6033
rlabel metal2 730 -31 730 -31 0 net=6033
rlabel metal2 163 -33 163 -33 0 net=969
rlabel metal2 180 -33 180 -33 0 net=3051
rlabel metal2 240 -33 240 -33 0 net=1039
rlabel metal2 289 -33 289 -33 0 net=1737
rlabel metal2 289 -33 289 -33 0 net=1737
rlabel metal2 352 -33 352 -33 0 net=1915
rlabel metal2 541 -33 541 -33 0 net=5537
rlabel metal2 611 -33 611 -33 0 net=5795
rlabel metal2 247 -35 247 -35 0 net=4864
rlabel metal2 257 -35 257 -35 0 net=2401
rlabel metal2 282 -35 282 -35 0 net=2655
rlabel metal2 359 -35 359 -35 0 net=2859
rlabel metal2 247 -37 247 -37 0 net=1271
rlabel metal2 303 -37 303 -37 0 net=2193
rlabel metal2 338 -37 338 -37 0 net=4149
rlabel metal2 303 -39 303 -39 0 net=1845
rlabel metal2 317 -41 317 -41 0 net=3195
rlabel metal2 58 -52 58 -52 0 net=843
rlabel metal2 58 -52 58 -52 0 net=843
rlabel metal2 65 -52 65 -52 0 net=4331
rlabel metal2 65 -52 65 -52 0 net=4331
rlabel metal2 79 -52 79 -52 0 net=5444
rlabel metal2 79 -52 79 -52 0 net=5444
rlabel metal2 93 -52 93 -52 0 net=4805
rlabel metal2 107 -52 107 -52 0 net=943
rlabel metal2 163 -52 163 -52 0 net=971
rlabel metal2 163 -52 163 -52 0 net=971
rlabel metal2 170 -52 170 -52 0 net=3052
rlabel metal2 226 -52 226 -52 0 net=798
rlabel metal2 310 -52 310 -52 0 net=2195
rlabel metal2 338 -52 338 -52 0 net=2283
rlabel metal2 415 -52 415 -52 0 net=2349
rlabel metal2 478 -52 478 -52 0 net=5393
rlabel metal2 513 -52 513 -52 0 net=5973
rlabel metal2 534 -52 534 -52 0 net=6217
rlabel metal2 660 -52 660 -52 0 net=4235
rlabel metal2 688 -52 688 -52 0 net=6335
rlabel metal2 730 -52 730 -52 0 net=6035
rlabel metal2 730 -52 730 -52 0 net=6035
rlabel metal2 793 -52 793 -52 0 net=4867
rlabel metal2 898 -52 898 -52 0 net=6677
rlabel metal2 898 -52 898 -52 0 net=6677
rlabel metal2 1087 -52 1087 -52 0 net=6643
rlabel metal2 110 -54 110 -54 0 net=236
rlabel metal2 229 -54 229 -54 0 net=4010
rlabel metal2 345 -54 345 -54 0 net=2441
rlabel metal2 345 -54 345 -54 0 net=2441
rlabel metal2 366 -54 366 -54 0 net=2861
rlabel metal2 366 -54 366 -54 0 net=2861
rlabel metal2 373 -54 373 -54 0 net=3737
rlabel metal2 429 -54 429 -54 0 net=6676
rlabel metal2 485 -54 485 -54 0 net=6407
rlabel metal2 541 -54 541 -54 0 net=4563
rlabel metal2 611 -54 611 -54 0 net=5797
rlabel metal2 611 -54 611 -54 0 net=5797
rlabel metal2 653 -54 653 -54 0 net=3913
rlabel metal2 786 -54 786 -54 0 net=5311
rlabel metal2 114 -56 114 -56 0 net=1251
rlabel metal2 114 -56 114 -56 0 net=1251
rlabel metal2 121 -56 121 -56 0 net=1666
rlabel metal2 142 -56 142 -56 0 net=3765
rlabel metal2 142 -56 142 -56 0 net=3765
rlabel metal2 170 -56 170 -56 0 net=803
rlabel metal2 233 -56 233 -56 0 net=1075
rlabel metal2 289 -56 289 -56 0 net=1739
rlabel metal2 373 -56 373 -56 0 net=3157
rlabel metal2 474 -56 474 -56 0 net=4757
rlabel metal2 499 -56 499 -56 0 net=6081
rlabel metal2 555 -56 555 -56 0 net=3339
rlabel metal2 128 -58 128 -58 0 net=1655
rlabel metal2 184 -58 184 -58 0 net=2402
rlabel metal2 289 -58 289 -58 0 net=2017
rlabel metal2 380 -58 380 -58 0 net=5447
rlabel metal2 422 -58 422 -58 0 net=60
rlabel metal2 471 -58 471 -58 0 net=5729
rlabel metal2 527 -58 527 -58 0 net=3639
rlabel metal2 569 -58 569 -58 0 net=5871
rlabel metal2 632 -58 632 -58 0 net=4181
rlabel metal2 135 -60 135 -60 0 net=1691
rlabel metal2 191 -60 191 -60 0 net=2569
rlabel metal2 233 -60 233 -60 0 net=1989
rlabel metal2 380 -60 380 -60 0 net=2829
rlabel metal2 422 -60 422 -60 0 net=3025
rlabel metal2 495 -60 495 -60 0 net=5875
rlabel metal2 632 -60 632 -60 0 net=3125
rlabel metal2 156 -62 156 -62 0 net=2051
rlabel metal2 208 -62 208 -62 0 net=998
rlabel metal2 240 -62 240 -62 0 net=1041
rlabel metal2 240 -62 240 -62 0 net=1041
rlabel metal2 247 -62 247 -62 0 net=1273
rlabel metal2 408 -62 408 -62 0 net=3069
rlabel metal2 576 -62 576 -62 0 net=5039
rlabel metal2 198 -64 198 -64 0 net=2657
rlabel metal2 429 -64 429 -64 0 net=4143
rlabel metal2 576 -64 576 -64 0 net=5495
rlabel metal2 212 -66 212 -66 0 net=1847
rlabel metal2 436 -66 436 -66 0 net=4015
rlabel metal2 597 -66 597 -66 0 net=6103
rlabel metal2 222 -68 222 -68 0 net=1659
rlabel metal2 268 -68 268 -68 0 net=1959
rlabel metal2 439 -68 439 -68 0 net=4123
rlabel metal2 590 -68 590 -68 0 net=5529
rlabel metal2 268 -70 268 -70 0 net=4151
rlabel metal2 562 -70 562 -70 0 net=5539
rlabel metal2 282 -72 282 -72 0 net=3197
rlabel metal2 548 -72 548 -72 0 net=5119
rlabel metal2 317 -74 317 -74 0 net=1917
rlabel metal2 446 -74 446 -74 0 net=4939
rlabel metal2 324 -76 324 -76 0 net=3237
rlabel metal2 324 -78 324 -78 0 net=2115
rlabel metal2 131 -80 131 -80 0 net=570
rlabel metal2 30 -91 30 -91 0 net=5961
rlabel metal2 51 -91 51 -91 0 net=4333
rlabel metal2 89 -91 89 -91 0 net=4806
rlabel metal2 100 -91 100 -91 0 net=2053
rlabel metal2 219 -91 219 -91 0 net=4153
rlabel metal2 275 -91 275 -91 0 net=2019
rlabel metal2 299 -91 299 -91 0 net=3238
rlabel metal2 366 -91 366 -91 0 net=2863
rlabel metal2 397 -91 397 -91 0 net=230
rlabel metal2 429 -91 429 -91 0 net=4144
rlabel metal2 527 -91 527 -91 0 net=3641
rlabel metal2 583 -91 583 -91 0 net=5041
rlabel metal2 583 -91 583 -91 0 net=5041
rlabel metal2 597 -91 597 -91 0 net=5531
rlabel metal2 646 -91 646 -91 0 net=3341
rlabel metal2 730 -91 730 -91 0 net=6037
rlabel metal2 758 -91 758 -91 0 net=3521
rlabel metal2 800 -91 800 -91 0 net=5313
rlabel metal2 898 -91 898 -91 0 net=6679
rlabel metal2 975 -91 975 -91 0 net=5891
rlabel metal2 1087 -91 1087 -91 0 net=6645
rlabel metal2 1087 -91 1087 -91 0 net=6645
rlabel metal2 54 -93 54 -93 0 net=3725
rlabel metal2 93 -93 93 -93 0 net=3767
rlabel metal2 149 -93 149 -93 0 net=944
rlabel metal2 261 -93 261 -93 0 net=1275
rlabel metal2 282 -93 282 -93 0 net=3198
rlabel metal2 303 -93 303 -93 0 net=1961
rlabel metal2 331 -93 331 -93 0 net=2197
rlabel metal2 331 -93 331 -93 0 net=2197
rlabel metal2 338 -93 338 -93 0 net=2285
rlabel metal2 387 -93 387 -93 0 net=3739
rlabel metal2 401 -93 401 -93 0 net=5449
rlabel metal2 450 -93 450 -93 0 net=4017
rlabel metal2 478 -93 478 -93 0 net=4125
rlabel metal2 541 -93 541 -93 0 net=4565
rlabel metal2 604 -93 604 -93 0 net=6105
rlabel metal2 674 -93 674 -93 0 net=4237
rlabel metal2 765 -93 765 -93 0 net=4869
rlabel metal2 58 -95 58 -95 0 net=845
rlabel metal2 58 -95 58 -95 0 net=845
rlabel metal2 107 -95 107 -95 0 net=2351
rlabel metal2 450 -95 450 -95 0 net=3127
rlabel metal2 681 -95 681 -95 0 net=4367
rlabel metal2 114 -97 114 -97 0 net=1252
rlabel metal2 114 -97 114 -97 0 net=1252
rlabel metal2 121 -97 121 -97 0 net=5693
rlabel metal2 240 -97 240 -97 0 net=1043
rlabel metal2 282 -97 282 -97 0 net=1919
rlabel metal2 327 -97 327 -97 0 net=2701
rlabel metal2 373 -97 373 -97 0 net=3159
rlabel metal2 457 -97 457 -97 0 net=4759
rlabel metal2 534 -97 534 -97 0 net=6083
rlabel metal2 702 -97 702 -97 0 net=6337
rlabel metal2 124 -99 124 -99 0 net=50
rlabel metal2 240 -99 240 -99 0 net=1660
rlabel metal2 303 -99 303 -99 0 net=1741
rlabel metal2 317 -99 317 -99 0 net=2117
rlabel metal2 380 -99 380 -99 0 net=2831
rlabel metal2 408 -99 408 -99 0 net=3071
rlabel metal2 467 -99 467 -99 0 net=6501
rlabel metal2 499 -99 499 -99 0 net=5731
rlabel metal2 541 -99 541 -99 0 net=5873
rlabel metal2 590 -99 590 -99 0 net=5541
rlabel metal2 660 -99 660 -99 0 net=3915
rlabel metal2 128 -101 128 -101 0 net=1656
rlabel metal2 324 -101 324 -101 0 net=438
rlabel metal2 520 -101 520 -101 0 net=5975
rlabel metal2 593 -101 593 -101 0 net=6627
rlabel metal2 128 -103 128 -103 0 net=2443
rlabel metal2 355 -103 355 -103 0 net=6089
rlabel metal2 562 -103 562 -103 0 net=5121
rlabel metal2 611 -103 611 -103 0 net=5799
rlabel metal2 135 -105 135 -105 0 net=1692
rlabel metal2 212 -105 212 -105 0 net=1849
rlabel metal2 362 -105 362 -105 0 net=4301
rlabel metal2 506 -105 506 -105 0 net=5395
rlabel metal2 618 -105 618 -105 0 net=6219
rlabel metal2 142 -107 142 -107 0 net=2659
rlabel metal2 212 -107 212 -107 0 net=1991
rlabel metal2 373 -107 373 -107 0 net=4091
rlabel metal2 548 -107 548 -107 0 net=4941
rlabel metal2 625 -107 625 -107 0 net=5877
rlabel metal2 149 -109 149 -109 0 net=4071
rlabel metal2 233 -109 233 -109 0 net=1077
rlabel metal2 387 -109 387 -109 0 net=3027
rlabel metal2 513 -109 513 -109 0 net=6409
rlabel metal2 156 -111 156 -111 0 net=973
rlabel metal2 198 -111 198 -111 0 net=5567
rlabel metal2 390 -111 390 -111 0 net=1
rlabel metal2 576 -111 576 -111 0 net=5497
rlabel metal2 163 -113 163 -113 0 net=805
rlabel metal2 205 -113 205 -113 0 net=1693
rlabel metal2 408 -113 408 -113 0 net=4537
rlabel metal2 576 -113 576 -113 0 net=4183
rlabel metal2 170 -115 170 -115 0 net=2571
rlabel metal2 229 -115 229 -115 0 net=2625
rlabel metal2 299 -115 299 -115 0 net=2599
rlabel metal2 191 -117 191 -117 0 net=1363
rlabel metal2 23 -128 23 -128 0 net=3699
rlabel metal2 47 -128 47 -128 0 net=3726
rlabel metal2 79 -128 79 -128 0 net=1393
rlabel metal2 121 -128 121 -128 0 net=5694
rlabel metal2 219 -128 219 -128 0 net=4154
rlabel metal2 338 -128 338 -128 0 net=2703
rlabel metal2 457 -128 457 -128 0 net=4760
rlabel metal2 495 -128 495 -128 0 net=3257
rlabel metal2 541 -128 541 -128 0 net=5874
rlabel metal2 656 -128 656 -128 0 net=2871
rlabel metal2 779 -128 779 -128 0 net=3523
rlabel metal2 905 -128 905 -128 0 net=6681
rlabel metal2 975 -128 975 -128 0 net=5893
rlabel metal2 975 -128 975 -128 0 net=5893
rlabel metal2 1087 -128 1087 -128 0 net=6647
rlabel metal2 1087 -128 1087 -128 0 net=6647
rlabel metal2 30 -130 30 -130 0 net=5962
rlabel metal2 121 -130 121 -130 0 net=1695
rlabel metal2 219 -130 219 -130 0 net=1921
rlabel metal2 296 -130 296 -130 0 net=1743
rlabel metal2 324 -130 324 -130 0 net=2763
rlabel metal2 345 -130 345 -130 0 net=1850
rlabel metal2 380 -130 380 -130 0 net=5450
rlabel metal2 443 -130 443 -130 0 net=3073
rlabel metal2 509 -130 509 -130 0 net=3795
rlabel metal2 555 -130 555 -130 0 net=5878
rlabel metal2 737 -130 737 -130 0 net=6039
rlabel metal2 30 -132 30 -132 0 net=4335
rlabel metal2 149 -132 149 -132 0 net=4072
rlabel metal2 394 -132 394 -132 0 net=2865
rlabel metal2 471 -132 471 -132 0 net=4019
rlabel metal2 583 -132 583 -132 0 net=5043
rlabel metal2 667 -132 667 -132 0 net=6107
rlabel metal2 51 -134 51 -134 0 net=847
rlabel metal2 149 -134 149 -134 0 net=1599
rlabel metal2 513 -134 513 -134 0 net=4539
rlabel metal2 590 -134 590 -134 0 net=3343
rlabel metal2 695 -134 695 -134 0 net=4871
rlabel metal2 156 -136 156 -136 0 net=974
rlabel metal2 170 -136 170 -136 0 net=2573
rlabel metal2 394 -136 394 -136 0 net=3161
rlabel metal2 450 -136 450 -136 0 net=3129
rlabel metal2 520 -136 520 -136 0 net=6091
rlabel metal2 58 -138 58 -138 0 net=5963
rlabel metal2 170 -138 170 -138 0 net=857
rlabel metal2 198 -138 198 -138 0 net=5568
rlabel metal2 401 -138 401 -138 0 net=2833
rlabel metal2 450 -138 450 -138 0 net=3367
rlabel metal2 604 -138 604 -138 0 net=5123
rlabel metal2 674 -138 674 -138 0 net=6221
rlabel metal2 142 -140 142 -140 0 net=2661
rlabel metal2 499 -140 499 -140 0 net=4303
rlabel metal2 562 -140 562 -140 0 net=5397
rlabel metal2 681 -140 681 -140 0 net=6629
rlabel metal2 135 -142 135 -142 0 net=4479
rlabel metal2 527 -142 527 -142 0 net=3643
rlabel metal2 604 -142 604 -142 0 net=4369
rlabel metal2 744 -142 744 -142 0 net=5315
rlabel metal2 142 -144 142 -144 0 net=807
rlabel metal2 205 -144 205 -144 0 net=1992
rlabel metal2 226 -144 226 -144 0 net=4427
rlabel metal2 492 -144 492 -144 0 net=4127
rlabel metal2 569 -144 569 -144 0 net=5977
rlabel metal2 730 -144 730 -144 0 net=6339
rlabel metal2 212 -146 212 -146 0 net=2021
rlabel metal2 282 -146 282 -146 0 net=3833
rlabel metal2 569 -146 569 -146 0 net=3917
rlabel metal2 709 -146 709 -146 0 net=5715
rlabel metal2 229 -148 229 -148 0 net=2600
rlabel metal2 618 -148 618 -148 0 net=5499
rlabel metal2 702 -148 702 -148 0 net=5149
rlabel metal2 233 -150 233 -150 0 net=1079
rlabel metal2 359 -150 359 -150 0 net=2287
rlabel metal2 534 -150 534 -150 0 net=5733
rlabel metal2 625 -150 625 -150 0 net=6411
rlabel metal2 233 -152 233 -152 0 net=3819
rlabel metal2 250 -152 250 -152 0 net=2626
rlabel metal2 275 -152 275 -152 0 net=1493
rlabel metal2 597 -152 597 -152 0 net=4567
rlabel metal2 632 -152 632 -152 0 net=5533
rlabel metal2 240 -154 240 -154 0 net=2119
rlabel metal2 334 -154 334 -154 0 net=4789
rlabel metal2 597 -154 597 -154 0 net=4239
rlabel metal2 72 -156 72 -156 0 net=1451
rlabel metal2 345 -156 345 -156 0 net=3740
rlabel metal2 478 -156 478 -156 0 net=4705
rlabel metal2 639 -156 639 -156 0 net=6085
rlabel metal2 243 -158 243 -158 0 net=648
rlabel metal2 366 -158 366 -158 0 net=1867
rlabel metal2 422 -158 422 -158 0 net=6241
rlabel metal2 247 -160 247 -160 0 net=1045
rlabel metal2 303 -160 303 -160 0 net=2199
rlabel metal2 436 -160 436 -160 0 net=4093
rlabel metal2 646 -160 646 -160 0 net=5543
rlabel metal2 254 -162 254 -162 0 net=2135
rlabel metal2 331 -162 331 -162 0 net=3203
rlabel metal2 478 -162 478 -162 0 net=3461
rlabel metal2 107 -164 107 -164 0 net=2353
rlabel metal2 387 -164 387 -164 0 net=3029
rlabel metal2 611 -164 611 -164 0 net=4943
rlabel metal2 660 -164 660 -164 0 net=5801
rlabel metal2 107 -166 107 -166 0 net=2445
rlabel metal2 261 -166 261 -166 0 net=1277
rlabel metal2 387 -166 387 -166 0 net=6502
rlabel metal2 537 -166 537 -166 0 net=5105
rlabel metal2 128 -168 128 -168 0 net=941
rlabel metal2 268 -168 268 -168 0 net=1963
rlabel metal2 576 -168 576 -168 0 net=4185
rlabel metal2 100 -170 100 -170 0 net=2055
rlabel metal2 523 -170 523 -170 0 net=5453
rlabel metal2 93 -172 93 -172 0 net=3769
rlabel metal2 114 -172 114 -172 0 net=3199
rlabel metal2 93 -174 93 -174 0 net=1253
rlabel metal2 177 -176 177 -176 0 net=1365
rlabel metal2 191 -178 191 -178 0 net=2403
rlabel metal2 16 -189 16 -189 0 net=2201
rlabel metal2 317 -189 317 -189 0 net=5454
rlabel metal2 758 -189 758 -189 0 net=2873
rlabel metal2 919 -189 919 -189 0 net=6683
rlabel metal2 975 -189 975 -189 0 net=5895
rlabel metal2 975 -189 975 -189 0 net=5895
rlabel metal2 1087 -189 1087 -189 0 net=6649
rlabel metal2 1087 -189 1087 -189 0 net=6649
rlabel metal2 30 -191 30 -191 0 net=4336
rlabel metal2 68 -191 68 -191 0 net=422
rlabel metal2 117 -191 117 -191 0 net=737
rlabel metal2 201 -191 201 -191 0 net=3820
rlabel metal2 240 -191 240 -191 0 net=2121
rlabel metal2 338 -191 338 -191 0 net=3031
rlabel metal2 460 -191 460 -191 0 net=6412
rlabel metal2 765 -191 765 -191 0 net=6087
rlabel metal2 821 -191 821 -191 0 net=6503
rlabel metal2 23 -193 23 -193 0 net=3700
rlabel metal2 72 -193 72 -193 0 net=1452
rlabel metal2 205 -193 205 -193 0 net=1081
rlabel metal2 355 -193 355 -193 0 net=4321
rlabel metal2 485 -193 485 -193 0 net=6321
rlabel metal2 23 -195 23 -195 0 net=3771
rlabel metal2 163 -195 163 -195 0 net=1367
rlabel metal2 184 -195 184 -195 0 net=2022
rlabel metal2 233 -195 233 -195 0 net=1965
rlabel metal2 292 -195 292 -195 0 net=2639
rlabel metal2 422 -195 422 -195 0 net=4020
rlabel metal2 562 -195 562 -195 0 net=3645
rlabel metal2 562 -195 562 -195 0 net=3645
rlabel metal2 660 -195 660 -195 0 net=5107
rlabel metal2 744 -195 744 -195 0 net=5317
rlabel metal2 772 -195 772 -195 0 net=6243
rlabel metal2 30 -197 30 -197 0 net=3201
rlabel metal2 142 -197 142 -197 0 net=809
rlabel metal2 261 -197 261 -197 0 net=1279
rlabel metal2 296 -197 296 -197 0 net=1745
rlabel metal2 345 -197 345 -197 0 net=6449
rlabel metal2 37 -199 37 -199 0 net=1047
rlabel metal2 303 -199 303 -199 0 net=1857
rlabel metal2 380 -199 380 -199 0 net=2575
rlabel metal2 674 -199 674 -199 0 net=5399
rlabel metal2 786 -199 786 -199 0 net=6109
rlabel metal2 859 -199 859 -199 0 net=6619
rlabel metal2 44 -201 44 -201 0 net=3835
rlabel metal2 352 -201 352 -201 0 net=4094
rlabel metal2 702 -201 702 -201 0 net=5151
rlabel metal2 751 -201 751 -201 0 net=6041
rlabel metal2 793 -201 793 -201 0 net=6223
rlabel metal2 72 -203 72 -203 0 net=2137
rlabel metal2 170 -203 170 -203 0 net=859
rlabel metal2 187 -203 187 -203 0 net=3083
rlabel metal2 359 -203 359 -203 0 net=2289
rlabel metal2 359 -203 359 -203 0 net=2289
rlabel metal2 373 -203 373 -203 0 net=3163
rlabel metal2 408 -203 408 -203 0 net=2705
rlabel metal2 495 -203 495 -203 0 net=3229
rlabel metal2 527 -203 527 -203 0 net=4129
rlabel metal2 681 -203 681 -203 0 net=5501
rlabel metal2 800 -203 800 -203 0 net=6341
rlabel metal2 79 -205 79 -205 0 net=1395
rlabel metal2 247 -205 247 -205 0 net=1495
rlabel metal2 408 -205 408 -205 0 net=4225
rlabel metal2 541 -205 541 -205 0 net=3797
rlabel metal2 604 -205 604 -205 0 net=4371
rlabel metal2 681 -205 681 -205 0 net=5535
rlabel metal2 709 -205 709 -205 0 net=5545
rlabel metal2 800 -205 800 -205 0 net=6061
rlabel metal2 79 -207 79 -207 0 net=2411
rlabel metal2 450 -207 450 -207 0 net=3369
rlabel metal2 534 -207 534 -207 0 net=3345
rlabel metal2 625 -207 625 -207 0 net=4569
rlabel metal2 737 -207 737 -207 0 net=5717
rlabel metal2 807 -207 807 -207 0 net=6631
rlabel metal2 107 -209 107 -209 0 net=2447
rlabel metal2 429 -209 429 -209 0 net=2867
rlabel metal2 478 -209 478 -209 0 net=3463
rlabel metal2 548 -209 548 -209 0 net=4305
rlabel metal2 646 -209 646 -209 0 net=4945
rlabel metal2 716 -209 716 -209 0 net=5803
rlabel metal2 821 -209 821 -209 0 net=3525
rlabel metal2 58 -211 58 -211 0 net=5965
rlabel metal2 583 -211 583 -211 0 net=4541
rlabel metal2 667 -211 667 -211 0 net=5125
rlabel metal2 779 -211 779 -211 0 net=6093
rlabel metal2 51 -213 51 -213 0 net=848
rlabel metal2 107 -213 107 -213 0 net=2809
rlabel metal2 142 -213 142 -213 0 net=1601
rlabel metal2 187 -213 187 -213 0 net=3813
rlabel metal2 695 -213 695 -213 0 net=4873
rlabel metal2 723 -213 723 -213 0 net=5979
rlabel metal2 828 -213 828 -213 0 net=6611
rlabel metal2 51 -215 51 -215 0 net=6249
rlabel metal2 114 -215 114 -215 0 net=942
rlabel metal2 149 -215 149 -215 0 net=1923
rlabel metal2 254 -215 254 -215 0 net=2136
rlabel metal2 324 -215 324 -215 0 net=2765
rlabel metal2 464 -215 464 -215 0 net=6209
rlabel metal2 835 -215 835 -215 0 net=6431
rlabel metal2 121 -217 121 -217 0 net=1697
rlabel metal2 191 -217 191 -217 0 net=2405
rlabel metal2 275 -217 275 -217 0 net=5735
rlabel metal2 632 -217 632 -217 0 net=4707
rlabel metal2 93 -219 93 -219 0 net=1255
rlabel metal2 310 -219 310 -219 0 net=2057
rlabel metal2 345 -219 345 -219 0 net=2171
rlabel metal2 499 -219 499 -219 0 net=4481
rlabel metal2 93 -221 93 -221 0 net=6459
rlabel metal2 121 -223 121 -223 0 net=1667
rlabel metal2 467 -223 467 -223 0 net=4487
rlabel metal2 173 -225 173 -225 0 net=2423
rlabel metal2 366 -225 366 -225 0 net=1868
rlabel metal2 471 -225 471 -225 0 net=3131
rlabel metal2 513 -225 513 -225 0 net=4791
rlabel metal2 289 -227 289 -227 0 net=2355
rlabel metal2 457 -227 457 -227 0 net=3075
rlabel metal2 506 -227 506 -227 0 net=3259
rlabel metal2 593 -227 593 -227 0 net=5655
rlabel metal2 443 -229 443 -229 0 net=3205
rlabel metal2 597 -229 597 -229 0 net=4241
rlabel metal2 653 -229 653 -229 0 net=5045
rlabel metal2 415 -231 415 -231 0 net=2835
rlabel metal2 611 -231 611 -231 0 net=4187
rlabel metal2 401 -233 401 -233 0 net=2663
rlabel metal2 425 -233 425 -233 0 net=4551
rlabel metal2 100 -235 100 -235 0 net=3569
rlabel metal2 569 -235 569 -235 0 net=3919
rlabel metal2 226 -237 226 -237 0 net=4429
rlabel metal2 30 -248 30 -248 0 net=3202
rlabel metal2 170 -248 170 -248 0 net=810
rlabel metal2 233 -248 233 -248 0 net=1966
rlabel metal2 352 -248 352 -248 0 net=3207
rlabel metal2 534 -248 534 -248 0 net=3347
rlabel metal2 534 -248 534 -248 0 net=3347
rlabel metal2 579 -248 579 -248 0 net=5546
rlabel metal2 877 -248 877 -248 0 net=6245
rlabel metal2 975 -248 975 -248 0 net=5897
rlabel metal2 1087 -248 1087 -248 0 net=6651
rlabel metal2 33 -250 33 -250 0 net=6
rlabel metal2 488 -250 488 -250 0 net=5980
rlabel metal2 877 -250 877 -250 0 net=6621
rlabel metal2 947 -250 947 -250 0 net=6685
rlabel metal2 37 -252 37 -252 0 net=1049
rlabel metal2 208 -252 208 -252 0 net=2576
rlabel metal2 586 -252 586 -252 0 net=6210
rlabel metal2 905 -252 905 -252 0 net=6451
rlabel metal2 905 -252 905 -252 0 net=6451
rlabel metal2 37 -254 37 -254 0 net=2619
rlabel metal2 93 -254 93 -254 0 net=1496
rlabel metal2 254 -254 254 -254 0 net=2407
rlabel metal2 380 -254 380 -254 0 net=2448
rlabel metal2 436 -254 436 -254 0 net=4322
rlabel metal2 527 -254 527 -254 0 net=3371
rlabel metal2 593 -254 593 -254 0 net=4552
rlabel metal2 758 -254 758 -254 0 net=5401
rlabel metal2 779 -254 779 -254 0 net=5719
rlabel metal2 828 -254 828 -254 0 net=6323
rlabel metal2 44 -256 44 -256 0 net=3836
rlabel metal2 383 -256 383 -256 0 net=3709
rlabel metal2 600 -256 600 -256 0 net=4946
rlabel metal2 765 -256 765 -256 0 net=5319
rlabel metal2 884 -256 884 -256 0 net=6343
rlabel metal2 47 -258 47 -258 0 net=1717
rlabel metal2 93 -258 93 -258 0 net=1859
rlabel metal2 394 -258 394 -258 0 net=3261
rlabel metal2 520 -258 520 -258 0 net=3231
rlabel metal2 597 -258 597 -258 0 net=5737
rlabel metal2 891 -258 891 -258 0 net=5937
rlabel metal2 58 -260 58 -260 0 net=1257
rlabel metal2 205 -260 205 -260 0 net=1083
rlabel metal2 268 -260 268 -260 0 net=1281
rlabel metal2 268 -260 268 -260 0 net=1281
rlabel metal2 275 -260 275 -260 0 net=5736
rlabel metal2 495 -260 495 -260 0 net=4130
rlabel metal2 702 -260 702 -260 0 net=4793
rlabel metal2 23 -262 23 -262 0 net=3772
rlabel metal2 233 -262 233 -262 0 net=1235
rlabel metal2 464 -262 464 -262 0 net=378
rlabel metal2 653 -262 653 -262 0 net=5109
rlabel metal2 23 -264 23 -264 0 net=6251
rlabel metal2 65 -264 65 -264 0 net=5147
rlabel metal2 478 -264 478 -264 0 net=5656
rlabel metal2 79 -266 79 -266 0 net=2413
rlabel metal2 338 -266 338 -266 0 net=3033
rlabel metal2 499 -266 499 -266 0 net=3133
rlabel metal2 562 -266 562 -266 0 net=3647
rlabel metal2 604 -266 604 -266 0 net=4543
rlabel metal2 695 -266 695 -266 0 net=4709
rlabel metal2 79 -268 79 -268 0 net=5839
rlabel metal2 82 -270 82 -270 0 net=1103
rlabel metal2 103 -270 103 -270 0 net=1698
rlabel metal2 135 -270 135 -270 0 net=2811
rlabel metal2 331 -270 331 -270 0 net=2123
rlabel metal2 373 -270 373 -270 0 net=3165
rlabel metal2 541 -270 541 -270 0 net=3465
rlabel metal2 583 -270 583 -270 0 net=3815
rlabel metal2 618 -270 618 -270 0 net=4189
rlabel metal2 695 -270 695 -270 0 net=5127
rlabel metal2 107 -272 107 -272 0 net=4430
rlabel metal2 576 -272 576 -272 0 net=3799
rlabel metal2 667 -272 667 -272 0 net=4489
rlabel metal2 117 -274 117 -274 0 net=1909
rlabel metal2 359 -274 359 -274 0 net=2291
rlabel metal2 411 -274 411 -274 0 net=5743
rlabel metal2 121 -276 121 -276 0 net=1669
rlabel metal2 121 -276 121 -276 0 net=1669
rlabel metal2 128 -276 128 -276 0 net=2059
rlabel metal2 359 -276 359 -276 0 net=2665
rlabel metal2 450 -276 450 -276 0 net=2869
rlabel metal2 583 -276 583 -276 0 net=5536
rlabel metal2 702 -276 702 -276 0 net=5047
rlabel metal2 135 -278 135 -278 0 net=1643
rlabel metal2 317 -278 317 -278 0 net=1747
rlabel metal2 415 -278 415 -278 0 net=6553
rlabel metal2 142 -280 142 -280 0 net=1603
rlabel metal2 422 -280 422 -280 0 net=2707
rlabel metal2 471 -280 471 -280 0 net=3077
rlabel metal2 639 -280 639 -280 0 net=4373
rlabel metal2 681 -280 681 -280 0 net=4571
rlabel metal2 709 -280 709 -280 0 net=6095
rlabel metal2 114 -282 114 -282 0 net=4761
rlabel metal2 723 -282 723 -282 0 net=5503
rlabel metal2 849 -282 849 -282 0 net=6613
rlabel metal2 114 -284 114 -284 0 net=1369
rlabel metal2 170 -284 170 -284 0 net=3085
rlabel metal2 422 -284 422 -284 0 net=2767
rlabel metal2 471 -284 471 -284 0 net=6088
rlabel metal2 912 -284 912 -284 0 net=6461
rlabel metal2 145 -286 145 -286 0 net=5165
rlabel metal2 429 -286 429 -286 0 net=2837
rlabel metal2 474 -286 474 -286 0 net=3399
rlabel metal2 625 -286 625 -286 0 net=4307
rlabel metal2 744 -286 744 -286 0 net=5153
rlabel metal2 912 -286 912 -286 0 net=6633
rlabel metal2 156 -288 156 -288 0 net=5966
rlabel metal2 625 -288 625 -288 0 net=4483
rlabel metal2 716 -288 716 -288 0 net=4875
rlabel metal2 821 -288 821 -288 0 net=3527
rlabel metal2 156 -290 156 -290 0 net=999
rlabel metal2 219 -290 219 -290 0 net=3167
rlabel metal2 401 -290 401 -290 0 net=3571
rlabel metal2 492 -290 492 -290 0 net=6315
rlabel metal2 163 -292 163 -292 0 net=553
rlabel metal2 632 -292 632 -292 0 net=4243
rlabel metal2 786 -292 786 -292 0 net=6043
rlabel metal2 177 -294 177 -294 0 net=861
rlabel metal2 219 -294 219 -294 0 net=1397
rlabel metal2 264 -294 264 -294 0 net=2549
rlabel metal2 366 -294 366 -294 0 net=2357
rlabel metal2 492 -294 492 -294 0 net=2875
rlabel metal2 16 -296 16 -296 0 net=2203
rlabel metal2 226 -296 226 -296 0 net=1097
rlabel metal2 310 -296 310 -296 0 net=2425
rlabel metal2 611 -296 611 -296 0 net=3921
rlabel metal2 786 -296 786 -296 0 net=5805
rlabel metal2 870 -296 870 -296 0 net=6505
rlabel metal2 16 -298 16 -298 0 net=6457
rlabel metal2 807 -298 807 -298 0 net=6111
rlabel metal2 863 -298 863 -298 0 net=6225
rlabel metal2 72 -300 72 -300 0 net=2139
rlabel metal2 408 -300 408 -300 0 net=4227
rlabel metal2 842 -300 842 -300 0 net=6063
rlabel metal2 863 -300 863 -300 0 net=6433
rlabel metal2 72 -302 72 -302 0 net=2173
rlabel metal2 842 -302 842 -302 0 net=6121
rlabel metal2 149 -304 149 -304 0 net=1925
rlabel metal2 898 -304 898 -304 0 net=6345
rlabel metal2 149 -306 149 -306 0 net=2641
rlabel metal2 229 -308 229 -308 0 net=2277
rlabel metal2 9 -319 9 -319 0 net=738
rlabel metal2 156 -319 156 -319 0 net=1001
rlabel metal2 156 -319 156 -319 0 net=1001
rlabel metal2 184 -319 184 -319 0 net=863
rlabel metal2 184 -319 184 -319 0 net=863
rlabel metal2 205 -319 205 -319 0 net=677
rlabel metal2 226 -319 226 -319 0 net=1283
rlabel metal2 296 -319 296 -319 0 net=3168
rlabel metal2 436 -319 436 -319 0 net=6462
rlabel metal2 933 -319 933 -319 0 net=5899
rlabel metal2 999 -319 999 -319 0 net=3831
rlabel metal2 1094 -319 1094 -319 0 net=6653
rlabel metal2 16 -321 16 -321 0 net=6458
rlabel metal2 523 -321 523 -321 0 net=5110
rlabel metal2 681 -321 681 -321 0 net=4573
rlabel metal2 716 -321 716 -321 0 net=6452
rlabel metal2 947 -321 947 -321 0 net=6227
rlabel metal2 16 -323 16 -323 0 net=1645
rlabel metal2 208 -323 208 -323 0 net=405
rlabel metal2 317 -323 317 -323 0 net=2551
rlabel metal2 527 -323 527 -323 0 net=3232
rlabel metal2 548 -323 548 -323 0 net=6246
rlabel metal2 964 -323 964 -323 0 net=5139
rlabel metal2 23 -325 23 -325 0 net=6252
rlabel metal2 121 -325 121 -325 0 net=1671
rlabel metal2 331 -325 331 -325 0 net=1910
rlabel metal2 541 -325 541 -325 0 net=4794
rlabel metal2 23 -327 23 -327 0 net=5167
rlabel metal2 345 -327 345 -327 0 net=1926
rlabel metal2 390 -327 390 -327 0 net=3166
rlabel metal2 534 -327 534 -327 0 net=3349
rlabel metal2 548 -327 548 -327 0 net=6226
rlabel metal2 37 -329 37 -329 0 net=2621
rlabel metal2 58 -329 58 -329 0 net=1258
rlabel metal2 443 -329 443 -329 0 net=3573
rlabel metal2 632 -329 632 -329 0 net=3923
rlabel metal2 681 -329 681 -329 0 net=6344
rlabel metal2 898 -329 898 -329 0 net=6347
rlabel metal2 40 -331 40 -331 0 net=3005
rlabel metal2 65 -331 65 -331 0 net=5148
rlabel metal2 212 -331 212 -331 0 net=2415
rlabel metal2 443 -331 443 -331 0 net=2499
rlabel metal2 499 -331 499 -331 0 net=3079
rlabel metal2 579 -331 579 -331 0 net=5635
rlabel metal2 44 -333 44 -333 0 net=5561
rlabel metal2 212 -333 212 -333 0 net=815
rlabel metal2 618 -333 618 -333 0 net=3801
rlabel metal2 716 -333 716 -333 0 net=6317
rlabel metal2 821 -333 821 -333 0 net=6045
rlabel metal2 65 -335 65 -335 0 net=1427
rlabel metal2 121 -335 121 -335 0 net=1749
rlabel metal2 338 -335 338 -335 0 net=2125
rlabel metal2 352 -335 352 -335 0 net=3208
rlabel metal2 359 -335 359 -335 0 net=2667
rlabel metal2 422 -335 422 -335 0 net=2769
rlabel metal2 786 -335 786 -335 0 net=5807
rlabel metal2 901 -335 901 -335 0 net=6686
rlabel metal2 30 -337 30 -337 0 net=592
rlabel metal2 453 -337 453 -337 0 net=5402
rlabel metal2 807 -337 807 -337 0 net=6113
rlabel metal2 828 -337 828 -337 0 net=6325
rlabel metal2 93 -339 93 -339 0 net=1861
rlabel metal2 352 -339 352 -339 0 net=3263
rlabel metal2 401 -339 401 -339 0 net=2359
rlabel metal2 457 -339 457 -339 0 net=3035
rlabel metal2 702 -339 702 -339 0 net=5049
rlabel metal2 835 -339 835 -339 0 net=6555
rlabel metal2 93 -341 93 -341 0 net=2897
rlabel metal2 191 -341 191 -341 0 net=3629
rlabel metal2 639 -341 639 -341 0 net=4309
rlabel metal2 744 -341 744 -341 0 net=4877
rlabel metal2 842 -341 842 -341 0 net=6123
rlabel metal2 100 -343 100 -343 0 net=1105
rlabel metal2 135 -343 135 -343 0 net=2815
rlabel metal2 254 -343 254 -343 0 net=1085
rlabel metal2 275 -343 275 -343 0 net=1605
rlabel metal2 359 -343 359 -343 0 net=2870
rlabel metal2 506 -343 506 -343 0 net=5379
rlabel metal2 849 -343 849 -343 0 net=6615
rlabel metal2 79 -345 79 -345 0 net=2633
rlabel metal2 590 -345 590 -345 0 net=3711
rlabel metal2 723 -345 723 -345 0 net=5505
rlabel metal2 863 -345 863 -345 0 net=6435
rlabel metal2 79 -347 79 -347 0 net=3087
rlabel metal2 219 -347 219 -347 0 net=1399
rlabel metal2 261 -347 261 -347 0 net=2279
rlabel metal2 380 -347 380 -347 0 net=5947
rlabel metal2 72 -349 72 -349 0 net=2175
rlabel metal2 394 -349 394 -349 0 net=2225
rlabel metal2 474 -349 474 -349 0 net=4513
rlabel metal2 751 -349 751 -349 0 net=5155
rlabel metal2 870 -349 870 -349 0 net=6507
rlabel metal2 72 -351 72 -351 0 net=1719
rlabel metal2 100 -351 100 -351 0 net=4689
rlabel metal2 149 -351 149 -351 0 net=2643
rlabel metal2 569 -351 569 -351 0 net=3401
rlabel metal2 684 -351 684 -351 0 net=1
rlabel metal2 758 -351 758 -351 0 net=5745
rlabel metal2 870 -351 870 -351 0 net=6635
rlabel metal2 86 -353 86 -353 0 net=2427
rlabel metal2 401 -353 401 -353 0 net=5291
rlabel metal2 877 -353 877 -353 0 net=6623
rlabel metal2 149 -355 149 -355 0 net=2813
rlabel metal2 275 -355 275 -355 0 net=2708
rlabel metal2 555 -355 555 -355 0 net=3373
rlabel metal2 586 -355 586 -355 0 net=4645
rlabel metal2 765 -355 765 -355 0 net=5739
rlabel metal2 891 -355 891 -355 0 net=5939
rlabel metal2 191 -357 191 -357 0 net=1789
rlabel metal2 513 -357 513 -357 0 net=3135
rlabel metal2 730 -357 730 -357 0 net=4711
rlabel metal2 793 -357 793 -357 0 net=5841
rlabel metal2 198 -359 198 -359 0 net=1051
rlabel metal2 282 -359 282 -359 0 net=2409
rlabel metal2 366 -359 366 -359 0 net=2505
rlabel metal2 688 -359 688 -359 0 net=4763
rlabel metal2 800 -359 800 -359 0 net=5321
rlabel metal2 114 -361 114 -361 0 net=1371
rlabel metal2 404 -361 404 -361 0 net=4393
rlabel metal2 128 -363 128 -363 0 net=2061
rlabel metal2 219 -363 219 -363 0 net=1413
rlabel metal2 611 -363 611 -363 0 net=4229
rlabel metal2 695 -363 695 -363 0 net=5129
rlabel metal2 33 -365 33 -365 0 net=1879
rlabel metal2 240 -365 240 -365 0 net=1099
rlabel metal2 429 -365 429 -365 0 net=2839
rlabel metal2 492 -365 492 -365 0 net=2877
rlabel metal2 611 -365 611 -365 0 net=4545
rlabel metal2 719 -365 719 -365 0 net=5749
rlabel metal2 737 -365 737 -365 0 net=4491
rlabel metal2 240 -367 240 -367 0 net=2337
rlabel metal2 429 -369 429 -369 0 net=3677
rlabel metal2 625 -369 625 -369 0 net=4485
rlabel metal2 737 -369 737 -369 0 net=3529
rlabel metal2 492 -371 492 -371 0 net=6155
rlabel metal2 495 -373 495 -373 0 net=331
rlabel metal2 597 -373 597 -373 0 net=3649
rlabel metal2 660 -373 660 -373 0 net=4245
rlabel metal2 856 -373 856 -373 0 net=6065
rlabel metal2 562 -375 562 -375 0 net=3467
rlabel metal2 646 -375 646 -375 0 net=4191
rlabel metal2 779 -375 779 -375 0 net=5721
rlabel metal2 338 -377 338 -377 0 net=5759
rlabel metal2 779 -377 779 -377 0 net=4753
rlabel metal2 562 -379 562 -379 0 net=6096
rlabel metal2 667 -381 667 -381 0 net=4375
rlabel metal2 604 -383 604 -383 0 net=3817
rlabel metal2 387 -385 387 -385 0 net=3561
rlabel metal2 373 -387 373 -387 0 net=2293
rlabel metal2 310 -389 310 -389 0 net=2141
rlabel metal2 233 -391 233 -391 0 net=1237
rlabel metal2 177 -393 177 -393 0 net=2205
rlabel metal2 16 -404 16 -404 0 net=1646
rlabel metal2 142 -404 142 -404 0 net=2814
rlabel metal2 180 -404 180 -404 0 net=2062
rlabel metal2 233 -404 233 -404 0 net=2206
rlabel metal2 282 -404 282 -404 0 net=1373
rlabel metal2 306 -404 306 -404 0 net=2410
rlabel metal2 331 -404 331 -404 0 net=2280
rlabel metal2 422 -404 422 -404 0 net=4363
rlabel metal2 800 -404 800 -404 0 net=5131
rlabel metal2 1066 -404 1066 -404 0 net=3832
rlabel metal2 16 -406 16 -406 0 net=2623
rlabel metal2 58 -406 58 -406 0 net=3007
rlabel metal2 233 -406 233 -406 0 net=947
rlabel metal2 576 -406 576 -406 0 net=3403
rlabel metal2 600 -406 600 -406 0 net=6636
rlabel metal2 877 -406 877 -406 0 net=5741
rlabel metal2 1108 -406 1108 -406 0 net=6655
rlabel metal2 23 -408 23 -408 0 net=5168
rlabel metal2 401 -408 401 -408 0 net=4764
rlabel metal2 800 -408 800 -408 0 net=5157
rlabel metal2 863 -408 863 -408 0 net=5747
rlabel metal2 23 -410 23 -410 0 net=3837
rlabel metal2 142 -410 142 -410 0 net=2779
rlabel metal2 184 -410 184 -410 0 net=865
rlabel metal2 184 -410 184 -410 0 net=865
rlabel metal2 191 -410 191 -410 0 net=1791
rlabel metal2 247 -410 247 -410 0 net=1101
rlabel metal2 254 -410 254 -410 0 net=1400
rlabel metal2 331 -410 331 -410 0 net=2645
rlabel metal2 502 -410 502 -410 0 net=346
rlabel metal2 1003 -410 1003 -410 0 net=6509
rlabel metal2 37 -412 37 -412 0 net=817
rlabel metal2 247 -412 247 -412 0 net=1053
rlabel metal2 268 -412 268 -412 0 net=1086
rlabel metal2 282 -412 282 -412 0 net=1863
rlabel metal2 296 -412 296 -412 0 net=1673
rlabel metal2 338 -412 338 -412 0 net=3678
rlabel metal2 436 -412 436 -412 0 net=2416
rlabel metal2 509 -412 509 -412 0 net=4486
rlabel metal2 740 -412 740 -412 0 net=6389
rlabel metal2 51 -414 51 -414 0 net=1497
rlabel metal2 128 -414 128 -414 0 net=1881
rlabel metal2 219 -414 219 -414 0 net=1415
rlabel metal2 317 -414 317 -414 0 net=2585
rlabel metal2 478 -414 478 -414 0 net=2635
rlabel metal2 523 -414 523 -414 0 net=5467
rlabel metal2 919 -414 919 -414 0 net=5949
rlabel metal2 1010 -414 1010 -414 0 net=6557
rlabel metal2 58 -416 58 -416 0 net=3089
rlabel metal2 100 -416 100 -416 0 net=4691
rlabel metal2 100 -416 100 -416 0 net=4691
rlabel metal2 107 -416 107 -416 0 net=1107
rlabel metal2 128 -416 128 -416 0 net=1003
rlabel metal2 219 -416 219 -416 0 net=1607
rlabel metal2 317 -416 317 -416 0 net=2177
rlabel metal2 425 -416 425 -416 0 net=5441
rlabel metal2 65 -418 65 -418 0 net=1428
rlabel metal2 145 -418 145 -418 0 net=630
rlabel metal2 240 -418 240 -418 0 net=2339
rlabel metal2 341 -418 341 -418 0 net=2126
rlabel metal2 359 -418 359 -418 0 net=2669
rlabel metal2 429 -418 429 -418 0 net=1197
rlabel metal2 555 -418 555 -418 0 net=3137
rlabel metal2 555 -418 555 -418 0 net=3137
rlabel metal2 586 -418 586 -418 0 net=6318
rlabel metal2 730 -418 730 -418 0 net=5751
rlabel metal2 947 -418 947 -418 0 net=6125
rlabel metal2 1041 -418 1041 -418 0 net=5140
rlabel metal2 44 -420 44 -420 0 net=5563
rlabel metal2 954 -420 954 -420 0 net=6157
rlabel metal2 44 -422 44 -422 0 net=1565
rlabel metal2 285 -422 285 -422 0 net=1
rlabel metal2 345 -422 345 -422 0 net=2770
rlabel metal2 548 -422 548 -422 0 net=3385
rlabel metal2 65 -424 65 -424 0 net=3265
rlabel metal2 366 -424 366 -424 0 net=2507
rlabel metal2 485 -424 485 -424 0 net=3037
rlabel metal2 590 -424 590 -424 0 net=3469
rlabel metal2 611 -424 611 -424 0 net=4547
rlabel metal2 611 -424 611 -424 0 net=4547
rlabel metal2 646 -424 646 -424 0 net=5761
rlabel metal2 975 -424 975 -424 0 net=6327
rlabel metal2 72 -426 72 -426 0 net=1720
rlabel metal2 156 -426 156 -426 0 net=3053
rlabel metal2 478 -426 478 -426 0 net=2023
rlabel metal2 639 -426 639 -426 0 net=3713
rlabel metal2 660 -426 660 -426 0 net=4193
rlabel metal2 709 -426 709 -426 0 net=4377
rlabel metal2 744 -426 744 -426 0 net=4575
rlabel metal2 905 -426 905 -426 0 net=5637
rlabel metal2 1017 -426 1017 -426 0 net=6617
rlabel metal2 30 -428 30 -428 0 net=2935
rlabel metal2 674 -428 674 -428 0 net=4247
rlabel metal2 744 -428 744 -428 0 net=4647
rlabel metal2 772 -428 772 -428 0 net=5051
rlabel metal2 1024 -428 1024 -428 0 net=6625
rlabel metal2 72 -430 72 -430 0 net=2429
rlabel metal2 93 -430 93 -430 0 net=2899
rlabel metal2 373 -430 373 -430 0 net=2143
rlabel metal2 373 -430 373 -430 0 net=2143
rlabel metal2 380 -430 380 -430 0 net=3325
rlabel metal2 926 -430 926 -430 0 net=6047
rlabel metal2 12 -432 12 -432 0 net=561
rlabel metal2 93 -432 93 -432 0 net=1751
rlabel metal2 240 -432 240 -432 0 net=2791
rlabel metal2 653 -432 653 -432 0 net=3925
rlabel metal2 688 -432 688 -432 0 net=4231
rlabel metal2 765 -432 765 -432 0 net=4713
rlabel metal2 793 -432 793 -432 0 net=5507
rlabel metal2 870 -432 870 -432 0 net=5941
rlabel metal2 926 -432 926 -432 0 net=6437
rlabel metal2 79 -434 79 -434 0 net=2879
rlabel metal2 527 -434 527 -434 0 net=316
rlabel metal2 569 -434 569 -434 0 net=3375
rlabel metal2 779 -434 779 -434 0 net=4755
rlabel metal2 121 -436 121 -436 0 net=2817
rlabel metal2 254 -436 254 -436 0 net=2227
rlabel metal2 408 -436 408 -436 0 net=2361
rlabel metal2 457 -436 457 -436 0 net=2841
rlabel metal2 534 -436 534 -436 0 net=3081
rlabel metal2 625 -436 625 -436 0 net=3651
rlabel metal2 653 -436 653 -436 0 net=3531
rlabel metal2 807 -436 807 -436 0 net=6115
rlabel metal2 835 -436 835 -436 0 net=4395
rlabel metal2 982 -436 982 -436 0 net=6349
rlabel metal2 149 -438 149 -438 0 net=901
rlabel metal2 471 -438 471 -438 0 net=4817
rlabel metal2 814 -438 814 -438 0 net=5293
rlabel metal2 940 -438 940 -438 0 net=6067
rlabel metal2 163 -440 163 -440 0 net=2753
rlabel metal2 268 -440 268 -440 0 net=2501
rlabel metal2 520 -440 520 -440 0 net=4837
rlabel metal2 835 -440 835 -440 0 net=5809
rlabel metal2 940 -440 940 -440 0 net=4577
rlabel metal2 982 -440 982 -440 0 net=6275
rlabel metal2 170 -442 170 -442 0 net=4457
rlabel metal2 842 -442 842 -442 0 net=5323
rlabel metal2 884 -442 884 -442 0 net=6229
rlabel metal2 170 -444 170 -444 0 net=1285
rlabel metal2 303 -444 303 -444 0 net=4933
rlabel metal2 856 -444 856 -444 0 net=5723
rlabel metal2 177 -446 177 -446 0 net=1239
rlabel metal2 387 -446 387 -446 0 net=2295
rlabel metal2 408 -446 408 -446 0 net=5967
rlabel metal2 310 -448 310 -448 0 net=2433
rlabel metal2 604 -448 604 -448 0 net=3563
rlabel metal2 681 -448 681 -448 0 net=5615
rlabel metal2 933 -448 933 -448 0 net=5901
rlabel metal2 443 -450 443 -450 0 net=2553
rlabel metal2 474 -450 474 -450 0 net=5133
rlabel metal2 891 -450 891 -450 0 net=5843
rlabel metal2 464 -452 464 -452 0 net=4337
rlabel metal2 828 -452 828 -452 0 net=5381
rlabel metal2 520 -454 520 -454 0 net=3818
rlabel metal2 681 -454 681 -454 0 net=3963
rlabel metal2 534 -456 534 -456 0 net=3351
rlabel metal2 604 -456 604 -456 0 net=3631
rlabel metal2 632 -456 632 -456 0 net=3803
rlabel metal2 688 -456 688 -456 0 net=4311
rlabel metal2 723 -456 723 -456 0 net=4515
rlabel metal2 786 -456 786 -456 0 net=4879
rlabel metal2 229 -458 229 -458 0 net=2975
rlabel metal2 583 -458 583 -458 0 net=3575
rlabel metal2 723 -458 723 -458 0 net=5065
rlabel metal2 366 -460 366 -460 0 net=1889
rlabel metal2 751 -460 751 -460 0 net=4493
rlabel metal2 404 -462 404 -462 0 net=4339
rlabel metal2 9 -473 9 -473 0 net=2435
rlabel metal2 324 -473 324 -473 0 net=1675
rlabel metal2 348 -473 348 -473 0 net=727
rlabel metal2 660 -473 660 -473 0 net=5724
rlabel metal2 975 -473 975 -473 0 net=4396
rlabel metal2 1174 -473 1174 -473 0 net=4215
rlabel metal2 16 -475 16 -475 0 net=2624
rlabel metal2 135 -475 135 -475 0 net=2781
rlabel metal2 156 -475 156 -475 0 net=3054
rlabel metal2 537 -475 537 -475 0 net=5132
rlabel metal2 16 -477 16 -477 0 net=4693
rlabel metal2 107 -477 107 -477 0 net=2228
rlabel metal2 261 -477 261 -477 0 net=1102
rlabel metal2 296 -477 296 -477 0 net=1417
rlabel metal2 397 -477 397 -477 0 net=2957
rlabel metal2 527 -477 527 -477 0 net=4756
rlabel metal2 1045 -477 1045 -477 0 net=6277
rlabel metal2 37 -479 37 -479 0 net=818
rlabel metal2 401 -479 401 -479 0 net=2842
rlabel metal2 527 -479 527 -479 0 net=3353
rlabel metal2 541 -479 541 -479 0 net=2977
rlabel metal2 541 -479 541 -479 0 net=2977
rlabel metal2 555 -479 555 -479 0 net=3139
rlabel metal2 555 -479 555 -479 0 net=3139
rlabel metal2 562 -479 562 -479 0 net=6618
rlabel metal2 37 -481 37 -481 0 net=2169
rlabel metal2 205 -481 205 -481 0 net=1793
rlabel metal2 240 -481 240 -481 0 net=2793
rlabel metal2 352 -481 352 -481 0 net=2901
rlabel metal2 436 -481 436 -481 0 net=2508
rlabel metal2 632 -481 632 -481 0 net=6626
rlabel metal2 23 -483 23 -483 0 net=3839
rlabel metal2 219 -483 219 -483 0 net=1608
rlabel metal2 415 -483 415 -483 0 net=2363
rlabel metal2 450 -483 450 -483 0 net=2586
rlabel metal2 695 -483 695 -483 0 net=4195
rlabel metal2 751 -483 751 -483 0 net=5135
rlabel metal2 870 -483 870 -483 0 net=5943
rlabel metal2 975 -483 975 -483 0 net=5951
rlabel metal2 1059 -483 1059 -483 0 net=6559
rlabel metal2 1122 -483 1122 -483 0 net=6009
rlabel metal2 23 -485 23 -485 0 net=2937
rlabel metal2 72 -485 72 -485 0 net=2431
rlabel metal2 289 -485 289 -485 0 net=1375
rlabel metal2 380 -485 380 -485 0 net=3327
rlabel metal2 565 -485 565 -485 0 net=6328
rlabel metal2 58 -487 58 -487 0 net=3091
rlabel metal2 415 -487 415 -487 0 net=2025
rlabel metal2 506 -487 506 -487 0 net=4232
rlabel metal2 733 -487 733 -487 0 net=5742
rlabel metal2 58 -489 58 -489 0 net=2145
rlabel metal2 450 -489 450 -489 0 net=3039
rlabel metal2 583 -489 583 -489 0 net=3471
rlabel metal2 593 -489 593 -489 0 net=5748
rlabel metal2 79 -491 79 -491 0 net=2881
rlabel metal2 586 -491 586 -491 0 net=5052
rlabel metal2 1010 -491 1010 -491 0 net=5639
rlabel metal2 1115 -491 1115 -491 0 net=6657
rlabel metal2 86 -493 86 -493 0 net=5564
rlabel metal2 961 -493 961 -493 0 net=5903
rlabel metal2 989 -493 989 -493 0 net=6049
rlabel metal2 86 -495 86 -495 0 net=1109
rlabel metal2 142 -495 142 -495 0 net=1891
rlabel metal2 457 -495 457 -495 0 net=4935
rlabel metal2 961 -495 961 -495 0 net=5969
rlabel metal2 93 -497 93 -497 0 net=1753
rlabel metal2 166 -497 166 -497 0 net=5442
rlabel metal2 93 -499 93 -499 0 net=2819
rlabel metal2 170 -499 170 -499 0 net=1287
rlabel metal2 240 -499 240 -499 0 net=1055
rlabel metal2 261 -499 261 -499 0 net=1199
rlabel metal2 460 -499 460 -499 0 net=4578
rlabel metal2 996 -499 996 -499 0 net=6127
rlabel metal2 100 -501 100 -501 0 net=1005
rlabel metal2 149 -501 149 -501 0 net=903
rlabel metal2 177 -501 177 -501 0 net=1241
rlabel metal2 289 -501 289 -501 0 net=2477
rlabel metal2 331 -501 331 -501 0 net=2647
rlabel metal2 429 -501 429 -501 0 net=1151
rlabel metal2 611 -501 611 -501 0 net=4549
rlabel metal2 884 -501 884 -501 0 net=6231
rlabel metal2 44 -503 44 -503 0 net=1567
rlabel metal2 443 -503 443 -503 0 net=2554
rlabel metal2 548 -503 548 -503 0 net=3387
rlabel metal2 632 -503 632 -503 0 net=3533
rlabel metal2 660 -503 660 -503 0 net=6211
rlabel metal2 1003 -503 1003 -503 0 net=6159
rlabel metal2 44 -505 44 -505 0 net=2179
rlabel metal2 387 -505 387 -505 0 net=6413
rlabel metal2 110 -507 110 -507 0 net=1027
rlabel metal2 184 -507 184 -507 0 net=867
rlabel metal2 184 -507 184 -507 0 net=867
rlabel metal2 191 -507 191 -507 0 net=1883
rlabel metal2 471 -507 471 -507 0 net=3082
rlabel metal2 604 -507 604 -507 0 net=3633
rlabel metal2 723 -507 723 -507 0 net=5294
rlabel metal2 1010 -507 1010 -507 0 net=6069
rlabel metal2 33 -509 33 -509 0 net=662
rlabel metal2 730 -509 730 -509 0 net=6375
rlabel metal2 1031 -509 1031 -509 0 net=6391
rlabel metal2 114 -511 114 -511 0 net=2297
rlabel metal2 478 -511 478 -511 0 net=2637
rlabel metal2 502 -511 502 -511 0 net=4085
rlabel metal2 754 -511 754 -511 0 net=4458
rlabel metal2 828 -511 828 -511 0 net=4881
rlabel metal2 849 -511 849 -511 0 net=5067
rlabel metal2 898 -511 898 -511 0 net=5469
rlabel metal2 1017 -511 1017 -511 0 net=6351
rlabel metal2 1080 -511 1080 -511 0 net=6511
rlabel metal2 128 -513 128 -513 0 net=917
rlabel metal2 485 -513 485 -513 0 net=3609
rlabel metal2 597 -513 597 -513 0 net=2509
rlabel metal2 152 -515 152 -515 0 net=514
rlabel metal2 597 -515 597 -515 0 net=4576
rlabel metal2 926 -515 926 -515 0 net=6439
rlabel metal2 163 -517 163 -517 0 net=2755
rlabel metal2 492 -517 492 -517 0 net=2671
rlabel metal2 765 -517 765 -517 0 net=3377
rlabel metal2 191 -519 191 -519 0 net=3979
rlabel metal2 779 -519 779 -519 0 net=4819
rlabel metal2 835 -519 835 -519 0 net=5811
rlabel metal2 247 -521 247 -521 0 net=887
rlabel metal2 422 -521 422 -521 0 net=4365
rlabel metal2 877 -521 877 -521 0 net=5617
rlabel metal2 121 -523 121 -523 0 net=1429
rlabel metal2 551 -523 551 -523 0 net=5647
rlabel metal2 268 -525 268 -525 0 net=2503
rlabel metal2 688 -525 688 -525 0 net=4313
rlabel metal2 786 -525 786 -525 0 net=4495
rlabel metal2 821 -525 821 -525 0 net=4839
rlabel metal2 268 -527 268 -527 0 net=1865
rlabel metal2 317 -527 317 -527 0 net=2670
rlabel metal2 667 -527 667 -527 0 net=3805
rlabel metal2 716 -527 716 -527 0 net=4379
rlabel metal2 793 -527 793 -527 0 net=5509
rlabel metal2 891 -527 891 -527 0 net=5383
rlabel metal2 138 -529 138 -529 0 net=4033
rlabel metal2 639 -529 639 -529 0 net=3653
rlabel metal2 681 -529 681 -529 0 net=3965
rlabel metal2 744 -529 744 -529 0 net=4649
rlabel metal2 800 -529 800 -529 0 net=5159
rlabel metal2 863 -529 863 -529 0 net=5325
rlabel metal2 233 -531 233 -531 0 net=949
rlabel metal2 355 -531 355 -531 0 net=4765
rlabel metal2 807 -531 807 -531 0 net=6117
rlabel metal2 51 -533 51 -533 0 net=1499
rlabel metal2 408 -533 408 -533 0 net=4131
rlabel metal2 863 -533 863 -533 0 net=5763
rlabel metal2 51 -535 51 -535 0 net=2341
rlabel metal2 548 -535 548 -535 0 net=3747
rlabel metal2 744 -535 744 -535 0 net=4517
rlabel metal2 772 -535 772 -535 0 net=4715
rlabel metal2 933 -535 933 -535 0 net=5845
rlabel metal2 338 -537 338 -537 0 net=1587
rlabel metal2 625 -537 625 -537 0 net=3565
rlabel metal2 702 -537 702 -537 0 net=4341
rlabel metal2 919 -537 919 -537 0 net=5753
rlabel metal2 562 -539 562 -539 0 net=5597
rlabel metal2 674 -541 674 -541 0 net=3927
rlabel metal2 709 -541 709 -541 0 net=4249
rlabel metal2 646 -543 646 -543 0 net=3715
rlabel metal2 709 -543 709 -543 0 net=4145
rlabel metal2 618 -545 618 -545 0 net=3577
rlabel metal2 576 -547 576 -547 0 net=3405
rlabel metal2 65 -549 65 -549 0 net=3267
rlabel metal2 65 -551 65 -551 0 net=3009
rlabel metal2 198 -553 198 -553 0 net=4338
rlabel metal2 215 -555 215 -555 0 net=2617
rlabel metal2 194 -557 194 -557 0 net=641
rlabel metal2 2 -568 2 -568 0 net=98
rlabel metal2 534 -568 534 -568 0 net=2979
rlabel metal2 548 -568 548 -568 0 net=4146
rlabel metal2 1059 -568 1059 -568 0 net=6561
rlabel metal2 1115 -568 1115 -568 0 net=6659
rlabel metal2 1115 -568 1115 -568 0 net=6659
rlabel metal2 1122 -568 1122 -568 0 net=6011
rlabel metal2 1122 -568 1122 -568 0 net=6011
rlabel metal2 1178 -568 1178 -568 0 net=4217
rlabel metal2 1178 -568 1178 -568 0 net=4217
rlabel metal2 9 -570 9 -570 0 net=2436
rlabel metal2 82 -570 82 -570 0 net=3583
rlabel metal2 712 -570 712 -570 0 net=4840
rlabel metal2 1087 -570 1087 -570 0 net=2511
rlabel metal2 9 -572 9 -572 0 net=3093
rlabel metal2 408 -572 408 -572 0 net=4366
rlabel metal2 842 -572 842 -572 0 net=4883
rlabel metal2 1024 -572 1024 -572 0 net=6377
rlabel metal2 1101 -572 1101 -572 0 net=5641
rlabel metal2 16 -574 16 -574 0 net=4695
rlabel metal2 975 -574 975 -574 0 net=5953
rlabel metal2 16 -576 16 -576 0 net=1111
rlabel metal2 121 -576 121 -576 0 net=1430
rlabel metal2 569 -576 569 -576 0 net=6118
rlabel metal2 23 -578 23 -578 0 net=2939
rlabel metal2 548 -578 548 -578 0 net=1853
rlabel metal2 23 -580 23 -580 0 net=506
rlabel metal2 443 -580 443 -580 0 net=2504
rlabel metal2 600 -580 600 -580 0 net=5068
rlabel metal2 919 -580 919 -580 0 net=5599
rlabel metal2 30 -582 30 -582 0 net=404
rlabel metal2 86 -582 86 -582 0 net=2794
rlabel metal2 303 -582 303 -582 0 net=1377
rlabel metal2 303 -582 303 -582 0 net=1377
rlabel metal2 338 -582 338 -582 0 net=1589
rlabel metal2 464 -582 464 -582 0 net=2618
rlabel metal2 702 -582 702 -582 0 net=3929
rlabel metal2 702 -582 702 -582 0 net=3929
rlabel metal2 733 -582 733 -582 0 net=4518
rlabel metal2 751 -582 751 -582 0 net=5137
rlabel metal2 968 -582 968 -582 0 net=5945
rlabel metal2 30 -584 30 -584 0 net=1201
rlabel metal2 268 -584 268 -584 0 net=1866
rlabel metal2 380 -584 380 -584 0 net=2673
rlabel metal2 506 -584 506 -584 0 net=6513
rlabel metal2 33 -586 33 -586 0 net=599
rlabel metal2 471 -586 471 -586 0 net=2757
rlabel metal2 604 -586 604 -586 0 net=6232
rlabel metal2 37 -588 37 -588 0 net=2170
rlabel metal2 191 -588 191 -588 0 net=1795
rlabel metal2 254 -588 254 -588 0 net=1242
rlabel metal2 513 -588 513 -588 0 net=3329
rlabel metal2 604 -588 604 -588 0 net=5970
rlabel metal2 1003 -588 1003 -588 0 net=6161
rlabel metal2 37 -590 37 -590 0 net=1007
rlabel metal2 107 -590 107 -590 0 net=909
rlabel metal2 275 -590 275 -590 0 net=2432
rlabel metal2 436 -590 436 -590 0 net=2365
rlabel metal2 478 -590 478 -590 0 net=2638
rlabel metal2 551 -590 551 -590 0 net=4550
rlabel metal2 877 -590 877 -590 0 net=5619
rlabel metal2 44 -592 44 -592 0 net=2181
rlabel metal2 555 -592 555 -592 0 net=3141
rlabel metal2 625 -592 625 -592 0 net=3749
rlabel metal2 688 -592 688 -592 0 net=3807
rlabel metal2 751 -592 751 -592 0 net=4251
rlabel metal2 761 -592 761 -592 0 net=6070
rlabel metal2 44 -594 44 -594 0 net=2821
rlabel metal2 107 -594 107 -594 0 net=2579
rlabel metal2 121 -594 121 -594 0 net=1423
rlabel metal2 205 -594 205 -594 0 net=3840
rlabel metal2 415 -594 415 -594 0 net=2027
rlabel metal2 555 -594 555 -594 0 net=3567
rlabel metal2 656 -594 656 -594 0 net=6512
rlabel metal2 54 -596 54 -596 0 net=4132
rlabel metal2 807 -596 807 -596 0 net=4717
rlabel metal2 926 -596 926 -596 0 net=5649
rlabel metal2 982 -596 982 -596 0 net=5905
rlabel metal2 1017 -596 1017 -596 0 net=6353
rlabel metal2 65 -598 65 -598 0 net=3011
rlabel metal2 611 -598 611 -598 0 net=3389
rlabel metal2 660 -598 660 -598 0 net=6440
rlabel metal2 68 -600 68 -600 0 net=4936
rlabel metal2 628 -600 628 -600 0 net=5191
rlabel metal2 765 -600 765 -600 0 net=4315
rlabel metal2 926 -600 926 -600 0 net=5813
rlabel metal2 954 -600 954 -600 0 net=5847
rlabel metal2 1045 -600 1045 -600 0 net=6279
rlabel metal2 72 -602 72 -602 0 net=2649
rlabel metal2 450 -602 450 -602 0 net=3041
rlabel metal2 632 -602 632 -602 0 net=3535
rlabel metal2 723 -602 723 -602 0 net=4087
rlabel metal2 821 -602 821 -602 0 net=5161
rlabel metal2 849 -602 849 -602 0 net=5511
rlabel metal2 989 -602 989 -602 0 net=6051
rlabel metal2 79 -604 79 -604 0 net=3777
rlabel metal2 905 -604 905 -604 0 net=5471
rlabel metal2 989 -604 989 -604 0 net=6415
rlabel metal2 75 -606 75 -606 0 net=5243
rlabel metal2 933 -606 933 -606 0 net=5755
rlabel metal2 996 -606 996 -606 0 net=6129
rlabel metal2 93 -608 93 -608 0 net=2771
rlabel metal2 611 -608 611 -608 0 net=3311
rlabel metal2 646 -608 646 -608 0 net=3579
rlabel metal2 765 -608 765 -608 0 net=4381
rlabel metal2 793 -608 793 -608 0 net=4767
rlabel metal2 940 -608 940 -608 0 net=6213
rlabel metal2 114 -610 114 -610 0 net=2299
rlabel metal2 485 -610 485 -610 0 net=3611
rlabel metal2 674 -610 674 -610 0 net=3717
rlabel metal2 800 -610 800 -610 0 net=3379
rlabel metal2 128 -612 128 -612 0 net=918
rlabel metal2 537 -612 537 -612 0 net=3679
rlabel metal2 772 -612 772 -612 0 net=4343
rlabel metal2 863 -612 863 -612 0 net=5765
rlabel metal2 1031 -612 1031 -612 0 net=6393
rlabel metal2 149 -614 149 -614 0 net=929
rlabel metal2 663 -614 663 -614 0 net=5999
rlabel metal2 152 -616 152 -616 0 net=1165
rlabel metal2 331 -616 331 -616 0 net=1569
rlabel metal2 373 -616 373 -616 0 net=1527
rlabel metal2 667 -616 667 -616 0 net=3655
rlabel metal2 695 -616 695 -616 0 net=3981
rlabel metal2 814 -616 814 -616 0 net=4497
rlabel metal2 166 -618 166 -618 0 net=5384
rlabel metal2 170 -620 170 -620 0 net=905
rlabel metal2 212 -620 212 -620 0 net=66
rlabel metal2 390 -620 390 -620 0 net=4477
rlabel metal2 891 -620 891 -620 0 net=5327
rlabel metal2 51 -622 51 -622 0 net=2343
rlabel metal2 583 -622 583 -622 0 net=3473
rlabel metal2 695 -622 695 -622 0 net=3983
rlabel metal2 828 -622 828 -622 0 net=4821
rlabel metal2 170 -624 170 -624 0 net=889
rlabel metal2 289 -624 289 -624 0 net=2479
rlabel metal2 583 -624 583 -624 0 net=3407
rlabel metal2 716 -624 716 -624 0 net=3967
rlabel metal2 786 -624 786 -624 0 net=4651
rlabel metal2 177 -626 177 -626 0 net=1029
rlabel metal2 233 -626 233 -626 0 net=1501
rlabel metal2 289 -626 289 -626 0 net=1709
rlabel metal2 653 -626 653 -626 0 net=3635
rlabel metal2 737 -626 737 -626 0 net=4197
rlabel metal2 100 -628 100 -628 0 net=3701
rlabel metal2 177 -630 177 -630 0 net=869
rlabel metal2 212 -630 212 -630 0 net=1407
rlabel metal2 341 -630 341 -630 0 net=5461
rlabel metal2 142 -632 142 -632 0 net=1893
rlabel metal2 345 -632 345 -632 0 net=1677
rlabel metal2 422 -632 422 -632 0 net=667
rlabel metal2 58 -634 58 -634 0 net=2146
rlabel metal2 348 -634 348 -634 0 net=2527
rlabel metal2 576 -634 576 -634 0 net=3269
rlabel metal2 58 -636 58 -636 0 net=1057
rlabel metal2 247 -636 247 -636 0 net=951
rlabel metal2 359 -636 359 -636 0 net=4035
rlabel metal2 135 -638 135 -638 0 net=2783
rlabel metal2 282 -638 282 -638 0 net=1117
rlabel metal2 359 -638 359 -638 0 net=2903
rlabel metal2 422 -638 422 -638 0 net=1829
rlabel metal2 135 -640 135 -640 0 net=1543
rlabel metal2 184 -640 184 -640 0 net=2041
rlabel metal2 401 -640 401 -640 0 net=1153
rlabel metal2 527 -640 527 -640 0 net=3355
rlabel metal2 142 -642 142 -642 0 net=1229
rlabel metal2 163 -644 163 -644 0 net=2925
rlabel metal2 219 -644 219 -644 0 net=1289
rlabel metal2 324 -644 324 -644 0 net=1885
rlabel metal2 499 -644 499 -644 0 net=2883
rlabel metal2 156 -646 156 -646 0 net=1755
rlabel metal2 310 -646 310 -646 0 net=1419
rlabel metal2 520 -646 520 -646 0 net=2959
rlabel metal2 310 -648 310 -648 0 net=1203
rlabel metal2 9 -659 9 -659 0 net=3095
rlabel metal2 9 -659 9 -659 0 net=3095
rlabel metal2 16 -659 16 -659 0 net=1113
rlabel metal2 149 -659 149 -659 0 net=930
rlabel metal2 254 -659 254 -659 0 net=1503
rlabel metal2 425 -659 425 -659 0 net=338
rlabel metal2 611 -659 611 -659 0 net=3313
rlabel metal2 691 -659 691 -659 0 net=5946
rlabel metal2 1003 -659 1003 -659 0 net=5849
rlabel metal2 1038 -659 1038 -659 0 net=5601
rlabel metal2 1059 -659 1059 -659 0 net=1855
rlabel metal2 1178 -659 1178 -659 0 net=4219
rlabel metal2 16 -661 16 -661 0 net=2577
rlabel metal2 187 -661 187 -661 0 net=541
rlabel metal2 254 -661 254 -661 0 net=2043
rlabel metal2 324 -661 324 -661 0 net=1420
rlabel metal2 387 -661 387 -661 0 net=1591
rlabel metal2 387 -661 387 -661 0 net=1591
rlabel metal2 408 -661 408 -661 0 net=3982
rlabel metal2 807 -661 807 -661 0 net=4089
rlabel metal2 849 -661 849 -661 0 net=4499
rlabel metal2 849 -661 849 -661 0 net=4499
rlabel metal2 933 -661 933 -661 0 net=6214
rlabel metal2 1038 -661 1038 -661 0 net=6661
rlabel metal2 23 -663 23 -663 0 net=1831
rlabel metal2 439 -663 439 -663 0 net=799
rlabel metal2 737 -663 737 -663 0 net=3703
rlabel metal2 737 -663 737 -663 0 net=3703
rlabel metal2 747 -663 747 -663 0 net=3718
rlabel metal2 807 -663 807 -663 0 net=4199
rlabel metal2 933 -663 933 -663 0 net=5473
rlabel metal2 975 -663 975 -663 0 net=5955
rlabel metal2 1045 -663 1045 -663 0 net=6053
rlabel metal2 1066 -663 1066 -663 0 net=6163
rlabel metal2 1066 -663 1066 -663 0 net=6163
rlabel metal2 1087 -663 1087 -663 0 net=6379
rlabel metal2 30 -665 30 -665 0 net=1202
rlabel metal2 481 -665 481 -665 0 net=5138
rlabel metal2 947 -665 947 -665 0 net=5757
rlabel metal2 996 -665 996 -665 0 net=5767
rlabel metal2 1087 -665 1087 -665 0 net=2512
rlabel metal2 37 -667 37 -667 0 net=1008
rlabel metal2 142 -667 142 -667 0 net=1230
rlabel metal2 345 -667 345 -667 0 net=1193
rlabel metal2 513 -667 513 -667 0 net=3580
rlabel metal2 695 -667 695 -667 0 net=3985
rlabel metal2 814 -667 814 -667 0 net=4719
rlabel metal2 898 -667 898 -667 0 net=4885
rlabel metal2 968 -667 968 -667 0 net=5651
rlabel metal2 1003 -667 1003 -667 0 net=6131
rlabel metal2 1090 -667 1090 -667 0 net=5295
rlabel metal2 37 -669 37 -669 0 net=1425
rlabel metal2 142 -669 142 -669 0 net=1797
rlabel metal2 205 -669 205 -669 0 net=290
rlabel metal2 443 -669 443 -669 0 net=5817
rlabel metal2 1031 -669 1031 -669 0 net=6001
rlabel metal2 1101 -669 1101 -669 0 net=6515
rlabel metal2 44 -671 44 -671 0 net=2822
rlabel metal2 159 -671 159 -671 0 net=2758
rlabel metal2 604 -671 604 -671 0 net=6416
rlabel metal2 1010 -671 1010 -671 0 net=5907
rlabel metal2 1080 -671 1080 -671 0 net=6355
rlabel metal2 1108 -671 1108 -671 0 net=6563
rlabel metal2 44 -673 44 -673 0 net=907
rlabel metal2 208 -673 208 -673 0 net=1408
rlabel metal2 226 -673 226 -673 0 net=1031
rlabel metal2 226 -673 226 -673 0 net=1031
rlabel metal2 233 -673 233 -673 0 net=911
rlabel metal2 268 -673 268 -673 0 net=2261
rlabel metal2 758 -673 758 -673 0 net=3969
rlabel metal2 842 -673 842 -673 0 net=5163
rlabel metal2 940 -673 940 -673 0 net=5463
rlabel metal2 1073 -673 1073 -673 0 net=6281
rlabel metal2 1108 -673 1108 -673 0 net=5642
rlabel metal2 51 -675 51 -675 0 net=3435
rlabel metal2 198 -675 198 -675 0 net=1379
rlabel metal2 324 -675 324 -675 0 net=1529
rlabel metal2 380 -675 380 -675 0 net=2675
rlabel metal2 523 -675 523 -675 0 net=3317
rlabel metal2 54 -677 54 -677 0 net=96
rlabel metal2 72 -677 72 -677 0 net=2650
rlabel metal2 457 -677 457 -677 0 net=3043
rlabel metal2 457 -677 457 -677 0 net=3043
rlabel metal2 464 -677 464 -677 0 net=2182
rlabel metal2 502 -677 502 -677 0 net=4347
rlabel metal2 940 -677 940 -677 0 net=5513
rlabel metal2 961 -677 961 -677 0 net=5621
rlabel metal2 1073 -677 1073 -677 0 net=6395
rlabel metal2 1122 -677 1122 -677 0 net=6013
rlabel metal2 58 -679 58 -679 0 net=1059
rlabel metal2 303 -679 303 -679 0 net=2301
rlabel metal2 464 -679 464 -679 0 net=3584
rlabel metal2 905 -679 905 -679 0 net=5245
rlabel metal2 58 -681 58 -681 0 net=1571
rlabel metal2 366 -681 366 -681 0 net=2345
rlabel metal2 450 -681 450 -681 0 net=2367
rlabel metal2 516 -681 516 -681 0 net=6417
rlabel metal2 65 -683 65 -683 0 net=3217
rlabel metal2 551 -683 551 -683 0 net=4316
rlabel metal2 884 -683 884 -683 0 net=4769
rlabel metal2 912 -683 912 -683 0 net=5329
rlabel metal2 72 -685 72 -685 0 net=1015
rlabel metal2 317 -685 317 -685 0 net=1895
rlabel metal2 366 -685 366 -685 0 net=1535
rlabel metal2 551 -685 551 -685 0 net=3408
rlabel metal2 597 -685 597 -685 0 net=3778
rlabel metal2 891 -685 891 -685 0 net=4823
rlabel metal2 79 -687 79 -687 0 net=1465
rlabel metal2 100 -687 100 -687 0 net=1757
rlabel metal2 310 -687 310 -687 0 net=1205
rlabel metal2 345 -687 345 -687 0 net=2029
rlabel metal2 499 -687 499 -687 0 net=4671
rlabel metal2 79 -689 79 -689 0 net=2581
rlabel metal2 114 -689 114 -689 0 net=1545
rlabel metal2 152 -689 152 -689 0 net=4923
rlabel metal2 380 -689 380 -689 0 net=5305
rlabel metal2 485 -689 485 -689 0 net=2481
rlabel metal2 569 -689 569 -689 0 net=3143
rlabel metal2 604 -689 604 -689 0 net=4478
rlabel metal2 870 -689 870 -689 0 net=4697
rlabel metal2 82 -691 82 -691 0 net=345
rlabel metal2 576 -691 576 -691 0 net=3357
rlabel metal2 660 -691 660 -691 0 net=3637
rlabel metal2 765 -691 765 -691 0 net=4383
rlabel metal2 86 -693 86 -693 0 net=1131
rlabel metal2 156 -693 156 -693 0 net=6023
rlabel metal2 89 -695 89 -695 0 net=330
rlabel metal2 219 -695 219 -695 0 net=1291
rlabel metal2 506 -695 506 -695 0 net=3013
rlabel metal2 614 -695 614 -695 0 net=5814
rlabel metal2 93 -697 93 -697 0 net=2773
rlabel metal2 135 -697 135 -697 0 net=4323
rlabel metal2 93 -699 93 -699 0 net=2927
rlabel metal2 177 -699 177 -699 0 net=871
rlabel metal2 177 -699 177 -699 0 net=871
rlabel metal2 184 -699 184 -699 0 net=2229
rlabel metal2 506 -699 506 -699 0 net=3381
rlabel metal2 821 -699 821 -699 0 net=4345
rlabel metal2 103 -701 103 -701 0 net=3568
rlabel metal2 646 -701 646 -701 0 net=3613
rlabel metal2 716 -701 716 -701 0 net=4075
rlabel metal2 800 -701 800 -701 0 net=4653
rlabel metal2 156 -703 156 -703 0 net=891
rlabel metal2 240 -703 240 -703 0 net=2785
rlabel metal2 534 -703 534 -703 0 net=2981
rlabel metal2 646 -703 646 -703 0 net=3537
rlabel metal2 688 -703 688 -703 0 net=3491
rlabel metal2 702 -703 702 -703 0 net=3931
rlabel metal2 163 -705 163 -705 0 net=953
rlabel metal2 275 -705 275 -705 0 net=1119
rlabel metal2 467 -705 467 -705 0 net=5053
rlabel metal2 170 -707 170 -707 0 net=2905
rlabel metal2 527 -707 527 -707 0 net=2885
rlabel metal2 541 -707 541 -707 0 net=2941
rlabel metal2 667 -707 667 -707 0 net=3475
rlabel metal2 688 -707 688 -707 0 net=5569
rlabel metal2 1041 -707 1041 -707 0 net=1
rlabel metal2 240 -709 240 -709 0 net=1167
rlabel metal2 429 -709 429 -709 0 net=1887
rlabel metal2 639 -709 639 -709 0 net=3391
rlabel metal2 730 -709 730 -709 0 net=5193
rlabel metal2 282 -711 282 -711 0 net=1679
rlabel metal2 401 -711 401 -711 0 net=1155
rlabel metal2 527 -711 527 -711 0 net=3271
rlabel metal2 639 -711 639 -711 0 net=3501
rlabel metal2 730 -711 730 -711 0 net=4037
rlabel metal2 33 -713 33 -713 0 net=138
rlabel metal2 411 -713 411 -713 0 net=3779
rlabel metal2 289 -715 289 -715 0 net=1711
rlabel metal2 562 -715 562 -715 0 net=3331
rlabel metal2 744 -715 744 -715 0 net=3809
rlabel metal2 289 -717 289 -717 0 net=2529
rlabel metal2 562 -717 562 -717 0 net=2961
rlabel metal2 744 -717 744 -717 0 net=4579
rlabel metal2 341 -719 341 -719 0 net=3185
rlabel metal2 751 -719 751 -719 0 net=4253
rlabel metal2 492 -721 492 -721 0 net=3681
rlabel metal2 625 -723 625 -723 0 net=3751
rlabel metal2 625 -725 625 -725 0 net=1431
rlabel metal2 674 -727 674 -727 0 net=3657
rlabel metal2 656 -729 656 -729 0 net=3415
rlabel metal2 9 -740 9 -740 0 net=3096
rlabel metal2 142 -740 142 -740 0 net=1799
rlabel metal2 142 -740 142 -740 0 net=1799
rlabel metal2 149 -740 149 -740 0 net=3145
rlabel metal2 600 -740 600 -740 0 net=5514
rlabel metal2 1038 -740 1038 -740 0 net=6662
rlabel metal2 1108 -740 1108 -740 0 net=6014
rlabel metal2 1143 -740 1143 -740 0 net=6565
rlabel metal2 9 -742 9 -742 0 net=2583
rlabel metal2 86 -742 86 -742 0 net=1132
rlabel metal2 163 -742 163 -742 0 net=954
rlabel metal2 373 -742 373 -742 0 net=4924
rlabel metal2 404 -742 404 -742 0 net=2482
rlabel metal2 502 -742 502 -742 0 net=3272
rlabel metal2 583 -742 583 -742 0 net=2607
rlabel metal2 765 -742 765 -742 0 net=3811
rlabel metal2 765 -742 765 -742 0 net=3811
rlabel metal2 782 -742 782 -742 0 net=6132
rlabel metal2 1031 -742 1031 -742 0 net=5851
rlabel metal2 1045 -742 1045 -742 0 net=5909
rlabel metal2 1045 -742 1045 -742 0 net=5909
rlabel metal2 1052 -742 1052 -742 0 net=6003
rlabel metal2 1122 -742 1122 -742 0 net=6419
rlabel metal2 1185 -742 1185 -742 0 net=4221
rlabel metal2 16 -744 16 -744 0 net=2578
rlabel metal2 359 -744 359 -744 0 net=5523
rlabel metal2 1059 -744 1059 -744 0 net=6055
rlabel metal2 1129 -744 1129 -744 0 net=6517
rlabel metal2 16 -746 16 -746 0 net=1537
rlabel metal2 373 -746 373 -746 0 net=1593
rlabel metal2 408 -746 408 -746 0 net=1433
rlabel metal2 639 -746 639 -746 0 net=675
rlabel metal2 821 -746 821 -746 0 net=5054
rlabel metal2 884 -746 884 -746 0 net=4673
rlabel metal2 1059 -746 1059 -746 0 net=5981
rlabel metal2 1101 -746 1101 -746 0 net=6357
rlabel metal2 1150 -746 1150 -746 0 net=1856
rlabel metal2 1164 -746 1164 -746 0 net=3319
rlabel metal2 23 -748 23 -748 0 net=1833
rlabel metal2 411 -748 411 -748 0 net=1504
rlabel metal2 439 -748 439 -748 0 net=2457
rlabel metal2 495 -748 495 -748 0 net=5758
rlabel metal2 968 -748 968 -748 0 net=5465
rlabel metal2 1080 -748 1080 -748 0 net=6283
rlabel metal2 1171 -748 1171 -748 0 net=5297
rlabel metal2 23 -750 23 -750 0 net=2031
rlabel metal2 387 -750 387 -750 0 net=2983
rlabel metal2 572 -750 572 -750 0 net=6193
rlabel metal2 30 -752 30 -752 0 net=2907
rlabel metal2 173 -752 173 -752 0 net=3239
rlabel metal2 212 -752 212 -752 0 net=1016
rlabel metal2 464 -752 464 -752 0 net=1195
rlabel metal2 513 -752 513 -752 0 net=2676
rlabel metal2 642 -752 642 -752 0 net=4384
rlabel metal2 926 -752 926 -752 0 net=5195
rlabel metal2 947 -752 947 -752 0 net=5247
rlabel metal2 989 -752 989 -752 0 net=5623
rlabel metal2 1115 -752 1115 -752 0 net=6381
rlabel metal2 37 -754 37 -754 0 net=1426
rlabel metal2 177 -754 177 -754 0 net=873
rlabel metal2 187 -754 187 -754 0 net=1888
rlabel metal2 625 -754 625 -754 0 net=4090
rlabel metal2 954 -754 954 -754 0 net=5169
rlabel metal2 37 -756 37 -756 0 net=1721
rlabel metal2 156 -756 156 -756 0 net=893
rlabel metal2 191 -756 191 -756 0 net=2044
rlabel metal2 324 -756 324 -756 0 net=1531
rlabel metal2 324 -756 324 -756 0 net=1531
rlabel metal2 331 -756 331 -756 0 net=2231
rlabel metal2 485 -756 485 -756 0 net=2787
rlabel metal2 520 -756 520 -756 0 net=5359
rlabel metal2 982 -756 982 -756 0 net=5571
rlabel metal2 996 -756 996 -756 0 net=5653
rlabel metal2 58 -758 58 -758 0 net=1573
rlabel metal2 366 -758 366 -758 0 net=2677
rlabel metal2 523 -758 523 -758 0 net=3638
rlabel metal2 663 -758 663 -758 0 net=6235
rlabel metal2 58 -760 58 -760 0 net=2929
rlabel metal2 100 -760 100 -760 0 net=1759
rlabel metal2 338 -760 338 -760 0 net=979
rlabel metal2 604 -760 604 -760 0 net=5377
rlabel metal2 65 -762 65 -762 0 net=3219
rlabel metal2 380 -762 380 -762 0 net=5306
rlabel metal2 688 -762 688 -762 0 net=5164
rlabel metal2 933 -762 933 -762 0 net=5475
rlabel metal2 996 -762 996 -762 0 net=5819
rlabel metal2 1073 -762 1073 -762 0 net=6397
rlabel metal2 44 -764 44 -764 0 net=908
rlabel metal2 394 -764 394 -764 0 net=4535
rlabel metal2 1010 -764 1010 -764 0 net=6025
rlabel metal2 44 -766 44 -766 0 net=2263
rlabel metal2 341 -766 341 -766 0 net=5835
rlabel metal2 1073 -766 1073 -766 0 net=5603
rlabel metal2 65 -768 65 -768 0 net=3383
rlabel metal2 527 -768 527 -768 0 net=2887
rlabel metal2 541 -768 541 -768 0 net=2943
rlabel metal2 565 -768 565 -768 0 net=4841
rlabel metal2 1017 -768 1017 -768 0 net=5769
rlabel metal2 79 -770 79 -770 0 net=3307
rlabel metal2 499 -770 499 -770 0 net=2945
rlabel metal2 569 -770 569 -770 0 net=5517
rlabel metal2 1017 -770 1017 -770 0 net=6165
rlabel metal2 86 -772 86 -772 0 net=1207
rlabel metal2 394 -772 394 -772 0 net=1157
rlabel metal2 506 -772 506 -772 0 net=3015
rlabel metal2 590 -772 590 -772 0 net=3187
rlabel metal2 688 -772 688 -772 0 net=3493
rlabel metal2 698 -772 698 -772 0 net=5307
rlabel metal2 93 -774 93 -774 0 net=1169
rlabel metal2 268 -774 268 -774 0 net=1807
rlabel metal2 317 -774 317 -774 0 net=1897
rlabel metal2 415 -774 415 -774 0 net=2013
rlabel metal2 702 -774 702 -774 0 net=3503
rlabel metal2 702 -774 702 -774 0 net=3503
rlabel metal2 716 -774 716 -774 0 net=4346
rlabel metal2 870 -774 870 -774 0 net=4581
rlabel metal2 100 -776 100 -776 0 net=2183
rlabel metal2 138 -776 138 -776 0 net=1017
rlabel metal2 163 -776 163 -776 0 net=2709
rlabel metal2 429 -776 429 -776 0 net=4699
rlabel metal2 114 -778 114 -778 0 net=1546
rlabel metal2 135 -778 135 -778 0 net=2530
rlabel metal2 457 -778 457 -778 0 net=3045
rlabel metal2 590 -778 590 -778 0 net=3333
rlabel metal2 737 -778 737 -778 0 net=3705
rlabel metal2 737 -778 737 -778 0 net=3705
rlabel metal2 744 -778 744 -778 0 net=5956
rlabel metal2 170 -780 170 -780 0 net=3169
rlabel metal2 247 -780 247 -780 0 net=1467
rlabel metal2 443 -780 443 -780 0 net=2347
rlabel metal2 485 -780 485 -780 0 net=3055
rlabel metal2 786 -780 786 -780 0 net=3781
rlabel metal2 191 -782 191 -782 0 net=1713
rlabel metal2 443 -782 443 -782 0 net=2369
rlabel metal2 492 -782 492 -782 0 net=3683
rlabel metal2 786 -782 786 -782 0 net=4201
rlabel metal2 842 -782 842 -782 0 net=4349
rlabel metal2 226 -784 226 -784 0 net=1033
rlabel metal2 289 -784 289 -784 0 net=3993
rlabel metal2 548 -784 548 -784 0 net=3823
rlabel metal2 779 -784 779 -784 0 net=3987
rlabel metal2 835 -784 835 -784 0 net=4325
rlabel metal2 849 -784 849 -784 0 net=4501
rlabel metal2 891 -784 891 -784 0 net=4771
rlabel metal2 128 -786 128 -786 0 net=1115
rlabel metal2 296 -786 296 -786 0 net=3315
rlabel metal2 656 -786 656 -786 0 net=5431
rlabel metal2 303 -788 303 -788 0 net=2303
rlabel metal2 548 -788 548 -788 0 net=2963
rlabel metal2 597 -788 597 -788 0 net=3753
rlabel metal2 779 -788 779 -788 0 net=3897
rlabel metal2 198 -790 198 -790 0 net=1381
rlabel metal2 555 -790 555 -790 0 net=5579
rlabel metal2 107 -792 107 -792 0 net=2775
rlabel metal2 562 -792 562 -792 0 net=4038
rlabel metal2 751 -792 751 -792 0 net=4255
rlabel metal2 849 -792 849 -792 0 net=4209
rlabel metal2 107 -794 107 -794 0 net=1293
rlabel metal2 474 -794 474 -794 0 net=4157
rlabel metal2 856 -794 856 -794 0 net=4887
rlabel metal2 219 -796 219 -796 0 net=3359
rlabel metal2 793 -796 793 -796 0 net=4077
rlabel metal2 912 -796 912 -796 0 net=4825
rlabel metal2 611 -798 611 -798 0 net=3393
rlabel metal2 772 -798 772 -798 0 net=3933
rlabel metal2 800 -798 800 -798 0 net=4655
rlabel metal2 912 -798 912 -798 0 net=5331
rlabel metal2 478 -800 478 -800 0 net=3863
rlabel metal2 814 -800 814 -800 0 net=4721
rlabel metal2 632 -802 632 -802 0 net=5255
rlabel metal2 632 -804 632 -804 0 net=3477
rlabel metal2 758 -804 758 -804 0 net=3971
rlabel metal2 51 -806 51 -806 0 net=3437
rlabel metal2 51 -808 51 -808 0 net=1681
rlabel metal2 621 -808 621 -808 0 net=4595
rlabel metal2 233 -810 233 -810 0 net=913
rlabel metal2 667 -810 667 -810 0 net=3615
rlabel metal2 233 -812 233 -812 0 net=1121
rlabel metal2 646 -812 646 -812 0 net=3539
rlabel metal2 261 -814 261 -814 0 net=1061
rlabel metal2 646 -814 646 -814 0 net=3417
rlabel metal2 674 -816 674 -816 0 net=3659
rlabel metal2 723 -818 723 -818 0 net=3193
rlabel metal2 19 -829 19 -829 0 net=72
rlabel metal2 355 -829 355 -829 0 net=4674
rlabel metal2 30 -831 30 -831 0 net=2908
rlabel metal2 121 -831 121 -831 0 net=5308
rlabel metal2 33 -833 33 -833 0 net=2601
rlabel metal2 184 -833 184 -833 0 net=875
rlabel metal2 184 -833 184 -833 0 net=875
rlabel metal2 198 -833 198 -833 0 net=2777
rlabel metal2 523 -833 523 -833 0 net=3334
rlabel metal2 618 -833 618 -833 0 net=4656
rlabel metal2 947 -833 947 -833 0 net=5249
rlabel metal2 947 -833 947 -833 0 net=5249
rlabel metal2 975 -833 975 -833 0 net=5433
rlabel metal2 975 -833 975 -833 0 net=5433
rlabel metal2 996 -833 996 -833 0 net=5821
rlabel metal2 1003 -833 1003 -833 0 net=5853
rlabel metal2 44 -835 44 -835 0 net=2264
rlabel metal2 590 -835 590 -835 0 net=3479
rlabel metal2 639 -835 639 -835 0 net=3505
rlabel metal2 726 -835 726 -835 0 net=5580
rlabel metal2 44 -837 44 -837 0 net=3995
rlabel metal2 303 -837 303 -837 0 net=1383
rlabel metal2 303 -837 303 -837 0 net=1383
rlabel metal2 359 -837 359 -837 0 net=3841
rlabel metal2 387 -837 387 -837 0 net=2984
rlabel metal2 485 -837 485 -837 0 net=3057
rlabel metal2 541 -837 541 -837 0 net=2944
rlabel metal2 541 -837 541 -837 0 net=2944
rlabel metal2 555 -837 555 -837 0 net=3394
rlabel metal2 656 -837 656 -837 0 net=3194
rlabel metal2 758 -837 758 -837 0 net=4597
rlabel metal2 905 -837 905 -837 0 net=5573
rlabel metal2 996 -837 996 -837 0 net=5519
rlabel metal2 1017 -837 1017 -837 0 net=6167
rlabel metal2 37 -839 37 -839 0 net=1723
rlabel metal2 394 -839 394 -839 0 net=1158
rlabel metal2 558 -839 558 -839 0 net=3395
rlabel metal2 656 -839 656 -839 0 net=5624
rlabel metal2 51 -841 51 -841 0 net=1682
rlabel metal2 296 -841 296 -841 0 net=3316
rlabel metal2 562 -841 562 -841 0 net=3189
rlabel metal2 611 -841 611 -841 0 net=5770
rlabel metal2 51 -843 51 -843 0 net=1715
rlabel metal2 198 -843 198 -843 0 net=1123
rlabel metal2 296 -843 296 -843 0 net=1533
rlabel metal2 362 -843 362 -843 0 net=2348
rlabel metal2 464 -843 464 -843 0 net=1196
rlabel metal2 660 -843 660 -843 0 net=3617
rlabel metal2 695 -843 695 -843 0 net=5654
rlabel metal2 1094 -843 1094 -843 0 net=6421
rlabel metal2 16 -845 16 -845 0 net=1539
rlabel metal2 205 -845 205 -845 0 net=3241
rlabel metal2 621 -845 621 -845 0 net=3812
rlabel metal2 779 -845 779 -845 0 net=4159
rlabel metal2 968 -845 968 -845 0 net=5361
rlabel metal2 1073 -845 1073 -845 0 net=5604
rlabel metal2 1178 -845 1178 -845 0 net=5299
rlabel metal2 58 -847 58 -847 0 net=2931
rlabel metal2 72 -847 72 -847 0 net=238
rlabel metal2 72 -847 72 -847 0 net=238
rlabel metal2 86 -847 86 -847 0 net=1208
rlabel metal2 380 -847 380 -847 0 net=6441
rlabel metal2 58 -849 58 -849 0 net=3171
rlabel metal2 289 -849 289 -849 0 net=4459
rlabel metal2 968 -849 968 -849 0 net=5477
rlabel metal2 989 -849 989 -849 0 net=6237
rlabel metal2 86 -851 86 -851 0 net=3439
rlabel metal2 695 -851 695 -851 0 net=3685
rlabel metal2 730 -851 730 -851 0 net=3973
rlabel metal2 814 -851 814 -851 0 net=6566
rlabel metal2 5 -853 5 -853 0 net=4593
rlabel metal2 982 -853 982 -853 0 net=6027
rlabel metal2 1129 -853 1129 -853 0 net=6519
rlabel metal2 1192 -853 1192 -853 0 net=4223
rlabel metal2 93 -855 93 -855 0 net=1171
rlabel metal2 292 -855 292 -855 0 net=4961
rlabel metal2 1017 -855 1017 -855 0 net=5983
rlabel metal2 1073 -855 1073 -855 0 net=6285
rlabel metal2 93 -857 93 -857 0 net=2185
rlabel metal2 114 -857 114 -857 0 net=5466
rlabel metal2 1059 -857 1059 -857 0 net=6057
rlabel metal2 117 -859 117 -859 0 net=1687
rlabel metal2 401 -859 401 -859 0 net=1835
rlabel metal2 401 -859 401 -859 0 net=1835
rlabel metal2 422 -859 422 -859 0 net=3016
rlabel metal2 569 -859 569 -859 0 net=2609
rlabel metal2 663 -859 663 -859 0 net=495
rlabel metal2 681 -859 681 -859 0 net=4536
rlabel metal2 999 -859 999 -859 0 net=1
rlabel metal2 1024 -859 1024 -859 0 net=5837
rlabel metal2 1122 -859 1122 -859 0 net=6399
rlabel metal2 121 -861 121 -861 0 net=1215
rlabel metal2 698 -861 698 -861 0 net=6194
rlabel metal2 1171 -861 1171 -861 0 net=4211
rlabel metal2 124 -863 124 -863 0 net=1116
rlabel metal2 324 -863 324 -863 0 net=3221
rlabel metal2 352 -863 352 -863 0 net=2233
rlabel metal2 450 -863 450 -863 0 net=2305
rlabel metal2 464 -863 464 -863 0 net=2893
rlabel metal2 506 -863 506 -863 0 net=3047
rlabel metal2 583 -863 583 -863 0 net=3495
rlabel metal2 702 -863 702 -863 0 net=3825
rlabel metal2 751 -863 751 -863 0 net=4257
rlabel metal2 786 -863 786 -863 0 net=4203
rlabel metal2 786 -863 786 -863 0 net=4203
rlabel metal2 863 -863 863 -863 0 net=4503
rlabel metal2 1024 -863 1024 -863 0 net=6005
rlabel metal2 1164 -863 1164 -863 0 net=3321
rlabel metal2 135 -865 135 -865 0 net=1575
rlabel metal2 425 -865 425 -865 0 net=4811
rlabel metal2 674 -865 674 -865 0 net=3661
rlabel metal2 716 -865 716 -865 0 net=3865
rlabel metal2 863 -865 863 -865 0 net=4773
rlabel metal2 1031 -865 1031 -865 0 net=5911
rlabel metal2 1080 -865 1080 -865 0 net=6383
rlabel metal2 23 -867 23 -867 0 net=2032
rlabel metal2 429 -867 429 -867 0 net=4701
rlabel metal2 751 -867 751 -867 0 net=3935
rlabel metal2 856 -867 856 -867 0 net=4889
rlabel metal2 1045 -867 1045 -867 0 net=6359
rlabel metal2 23 -869 23 -869 0 net=3361
rlabel metal2 226 -869 226 -869 0 net=1009
rlabel metal2 317 -869 317 -869 0 net=1899
rlabel metal2 429 -869 429 -869 0 net=2371
rlabel metal2 471 -869 471 -869 0 net=2459
rlabel metal2 758 -869 758 -869 0 net=3989
rlabel metal2 835 -869 835 -869 0 net=4723
rlabel metal2 870 -869 870 -869 0 net=3899
rlabel metal2 107 -871 107 -871 0 net=1295
rlabel metal2 436 -871 436 -871 0 net=3754
rlabel metal2 600 -871 600 -871 0 net=4277
rlabel metal2 807 -871 807 -871 0 net=4327
rlabel metal2 870 -871 870 -871 0 net=5257
rlabel metal2 65 -873 65 -873 0 net=3384
rlabel metal2 674 -873 674 -873 0 net=5524
rlabel metal2 65 -875 65 -875 0 net=2947
rlabel metal2 576 -875 576 -875 0 net=3419
rlabel metal2 677 -875 677 -875 0 net=4951
rlabel metal2 842 -875 842 -875 0 net=4583
rlabel metal2 898 -875 898 -875 0 net=3783
rlabel metal2 79 -877 79 -877 0 net=3309
rlabel metal2 149 -877 149 -877 0 net=3147
rlabel metal2 471 -877 471 -877 0 net=3855
rlabel metal2 772 -877 772 -877 0 net=4079
rlabel metal2 877 -877 877 -877 0 net=4827
rlabel metal2 37 -879 37 -879 0 net=919
rlabel metal2 163 -879 163 -879 0 net=5378
rlabel metal2 156 -881 156 -881 0 net=1019
rlabel metal2 177 -881 177 -881 0 net=895
rlabel metal2 485 -881 485 -881 0 net=2789
rlabel metal2 534 -881 534 -881 0 net=2965
rlabel metal2 646 -881 646 -881 0 net=3541
rlabel metal2 817 -881 817 -881 0 net=5881
rlabel metal2 142 -883 142 -883 0 net=1801
rlabel metal2 205 -883 205 -883 0 net=1034
rlabel metal2 415 -883 415 -883 0 net=2015
rlabel metal2 709 -883 709 -883 0 net=3707
rlabel metal2 128 -885 128 -885 0 net=801
rlabel metal2 149 -885 149 -885 0 net=1243
rlabel metal2 348 -885 348 -885 0 net=3429
rlabel metal2 513 -885 513 -885 0 net=2889
rlabel metal2 544 -885 544 -885 0 net=5087
rlabel metal2 9 -887 9 -887 0 net=2584
rlabel metal2 156 -887 156 -887 0 net=819
rlabel metal2 527 -887 527 -887 0 net=2733
rlabel metal2 737 -887 737 -887 0 net=4843
rlabel metal2 9 -889 9 -889 0 net=2711
rlabel metal2 366 -889 366 -889 0 net=2679
rlabel metal2 933 -889 933 -889 0 net=5197
rlabel metal2 212 -891 212 -891 0 net=1761
rlabel metal2 926 -891 926 -891 0 net=4351
rlabel metal2 212 -893 212 -893 0 net=1435
rlabel metal2 926 -893 926 -893 0 net=5171
rlabel metal2 219 -895 219 -895 0 net=915
rlabel metal2 366 -895 366 -895 0 net=1595
rlabel metal2 912 -895 912 -895 0 net=5333
rlabel metal2 40 -897 40 -897 0 net=1065
rlabel metal2 912 -897 912 -897 0 net=5077
rlabel metal2 254 -899 254 -899 0 net=981
rlabel metal2 268 -901 268 -901 0 net=1809
rlabel metal2 268 -903 268 -903 0 net=1063
rlabel metal2 310 -903 310 -903 0 net=1469
rlabel metal2 310 -905 310 -905 0 net=2245
rlabel metal2 2 -916 2 -916 0 net=3441
rlabel metal2 96 -916 96 -916 0 net=2790
rlabel metal2 502 -916 502 -916 0 net=2890
rlabel metal2 548 -916 548 -916 0 net=2016
rlabel metal2 684 -916 684 -916 0 net=5838
rlabel metal2 1136 -916 1136 -916 0 net=5300
rlabel metal2 19 -918 19 -918 0 net=4594
rlabel metal2 824 -918 824 -918 0 net=6019
rlabel metal2 1101 -918 1101 -918 0 net=6443
rlabel metal2 1150 -918 1150 -918 0 net=3323
rlabel metal2 30 -920 30 -920 0 net=2603
rlabel metal2 205 -920 205 -920 0 net=3421
rlabel metal2 597 -920 597 -920 0 net=5258
rlabel metal2 898 -920 898 -920 0 net=6400
rlabel metal2 1157 -920 1157 -920 0 net=4213
rlabel metal2 33 -922 33 -922 0 net=2778
rlabel metal2 506 -922 506 -922 0 net=3049
rlabel metal2 548 -922 548 -922 0 net=3191
rlabel metal2 597 -922 597 -922 0 net=4461
rlabel metal2 1108 -922 1108 -922 0 net=3901
rlabel metal2 37 -924 37 -924 0 net=3242
rlabel metal2 618 -924 618 -924 0 net=3827
rlabel metal2 716 -924 716 -924 0 net=3867
rlabel metal2 1164 -924 1164 -924 0 net=4224
rlabel metal2 40 -926 40 -926 0 net=3222
rlabel metal2 338 -926 338 -926 0 net=1471
rlabel metal2 338 -926 338 -926 0 net=1471
rlabel metal2 345 -926 345 -926 0 net=2681
rlabel metal2 499 -926 499 -926 0 net=5205
rlabel metal2 1066 -926 1066 -926 0 net=6169
rlabel metal2 1122 -926 1122 -926 0 net=6521
rlabel metal2 1185 -926 1185 -926 0 net=5179
rlabel metal2 9 -928 9 -928 0 net=2713
rlabel metal2 348 -928 348 -928 0 net=1810
rlabel metal2 415 -928 415 -928 0 net=3431
rlabel metal2 555 -928 555 -928 0 net=6119
rlabel metal2 40 -930 40 -930 0 net=3951
rlabel metal2 628 -930 628 -930 0 net=3708
rlabel metal2 716 -930 716 -930 0 net=3975
rlabel metal2 737 -930 737 -930 0 net=4845
rlabel metal2 1052 -930 1052 -930 0 net=3784
rlabel metal2 44 -932 44 -932 0 net=3997
rlabel metal2 656 -932 656 -932 0 net=6238
rlabel metal2 1052 -932 1052 -932 0 net=6385
rlabel metal2 44 -934 44 -934 0 net=2933
rlabel metal2 117 -934 117 -934 0 net=41
rlabel metal2 394 -934 394 -934 0 net=1763
rlabel metal2 394 -934 394 -934 0 net=1763
rlabel metal2 401 -934 401 -934 0 net=1837
rlabel metal2 401 -934 401 -934 0 net=1837
rlabel metal2 408 -934 408 -934 0 net=4559
rlabel metal2 562 -934 562 -934 0 net=2611
rlabel metal2 667 -934 667 -934 0 net=3687
rlabel metal2 702 -934 702 -934 0 net=4081
rlabel metal2 975 -934 975 -934 0 net=5435
rlabel metal2 51 -936 51 -936 0 net=1716
rlabel metal2 142 -936 142 -936 0 net=802
rlabel metal2 163 -936 163 -936 0 net=1021
rlabel metal2 163 -936 163 -936 0 net=1021
rlabel metal2 170 -936 170 -936 0 net=1631
rlabel metal2 219 -936 219 -936 0 net=916
rlabel metal2 439 -936 439 -936 0 net=3396
rlabel metal2 674 -936 674 -936 0 net=4039
rlabel metal2 737 -936 737 -936 0 net=4205
rlabel metal2 975 -936 975 -936 0 net=5985
rlabel metal2 51 -938 51 -938 0 net=1401
rlabel metal2 65 -938 65 -938 0 net=2949
rlabel metal2 632 -938 632 -938 0 net=3543
rlabel metal2 695 -938 695 -938 0 net=4917
rlabel metal2 989 -938 989 -938 0 net=5913
rlabel metal2 58 -940 58 -940 0 net=3173
rlabel metal2 142 -940 142 -940 0 net=1683
rlabel metal2 268 -940 268 -940 0 net=1064
rlabel metal2 303 -940 303 -940 0 net=1385
rlabel metal2 331 -940 331 -940 0 net=1901
rlabel metal2 439 -940 439 -940 0 net=294
rlabel metal2 996 -940 996 -940 0 net=5521
rlabel metal2 58 -942 58 -942 0 net=3310
rlabel metal2 149 -942 149 -942 0 net=897
rlabel metal2 247 -942 247 -942 0 net=1245
rlabel metal2 303 -942 303 -942 0 net=1311
rlabel metal2 772 -942 772 -942 0 net=4775
rlabel metal2 961 -942 961 -942 0 net=5883
rlabel metal2 1017 -942 1017 -942 0 net=6287
rlabel metal2 72 -944 72 -944 0 net=481
rlabel metal2 786 -944 786 -944 0 net=4963
rlabel metal2 961 -944 961 -944 0 net=5823
rlabel metal2 1038 -944 1038 -944 0 net=5363
rlabel metal2 79 -946 79 -946 0 net=921
rlabel metal2 191 -946 191 -946 0 net=1541
rlabel metal2 226 -946 226 -946 0 net=1011
rlabel metal2 226 -946 226 -946 0 net=1011
rlabel metal2 233 -946 233 -946 0 net=1647
rlabel metal2 380 -946 380 -946 0 net=1688
rlabel metal2 709 -946 709 -946 0 net=6028
rlabel metal2 1010 -946 1010 -946 0 net=6423
rlabel metal2 79 -948 79 -948 0 net=1351
rlabel metal2 156 -948 156 -948 0 net=821
rlabel metal2 212 -948 212 -948 0 net=1437
rlabel metal2 261 -948 261 -948 0 net=4659
rlabel metal2 362 -948 362 -948 0 net=1993
rlabel metal2 982 -948 982 -948 0 net=5385
rlabel metal2 86 -950 86 -950 0 net=2187
rlabel metal2 121 -950 121 -950 0 net=1217
rlabel metal2 156 -950 156 -950 0 net=1125
rlabel metal2 240 -950 240 -950 0 net=1173
rlabel metal2 268 -950 268 -950 0 net=1597
rlabel metal2 373 -950 373 -950 0 net=2460
rlabel metal2 800 -950 800 -950 0 net=4725
rlabel metal2 1059 -950 1059 -950 0 net=6059
rlabel metal2 9 -952 9 -952 0 net=2397
rlabel metal2 177 -952 177 -952 0 net=1803
rlabel metal2 240 -952 240 -952 0 net=983
rlabel metal2 275 -952 275 -952 0 net=1534
rlabel metal2 352 -952 352 -952 0 net=2235
rlabel metal2 380 -952 380 -952 0 net=1725
rlabel metal2 471 -952 471 -952 0 net=3857
rlabel metal2 607 -952 607 -952 0 net=5815
rlabel metal2 23 -954 23 -954 0 net=3363
rlabel metal2 275 -954 275 -954 0 net=1067
rlabel metal2 296 -954 296 -954 0 net=1297
rlabel metal2 471 -954 471 -954 0 net=3497
rlabel metal2 625 -954 625 -954 0 net=4813
rlabel metal2 1024 -954 1024 -954 0 net=6007
rlabel metal2 23 -956 23 -956 0 net=2531
rlabel metal2 135 -956 135 -956 0 net=1577
rlabel metal2 478 -956 478 -956 0 net=3059
rlabel metal2 583 -956 583 -956 0 net=3619
rlabel metal2 723 -956 723 -956 0 net=4161
rlabel metal2 821 -956 821 -956 0 net=5487
rlabel metal2 72 -958 72 -958 0 net=4455
rlabel metal2 317 -958 317 -958 0 net=2247
rlabel metal2 485 -958 485 -958 0 net=2735
rlabel metal2 544 -958 544 -958 0 net=4135
rlabel metal2 744 -958 744 -958 0 net=4703
rlabel metal2 821 -958 821 -958 0 net=5575
rlabel metal2 93 -960 93 -960 0 net=6463
rlabel metal2 135 -962 135 -962 0 net=1339
rlabel metal2 653 -962 653 -962 0 net=3663
rlabel metal2 744 -962 744 -962 0 net=4279
rlabel metal2 905 -962 905 -962 0 net=5335
rlabel metal2 177 -964 177 -964 0 net=877
rlabel metal2 359 -964 359 -964 0 net=3843
rlabel metal2 527 -964 527 -964 0 net=2967
rlabel metal2 688 -964 688 -964 0 net=3937
rlabel metal2 793 -964 793 -964 0 net=4329
rlabel metal2 954 -964 954 -964 0 net=5479
rlabel metal2 184 -966 184 -966 0 net=2745
rlabel metal2 443 -966 443 -966 0 net=3149
rlabel metal2 751 -966 751 -966 0 net=4599
rlabel metal2 968 -966 968 -966 0 net=6361
rlabel metal2 422 -968 422 -968 0 net=6071
rlabel metal2 422 -970 422 -970 0 net=2895
rlabel metal2 807 -970 807 -970 0 net=4829
rlabel metal2 429 -972 429 -972 0 net=2373
rlabel metal2 450 -972 450 -972 0 net=3481
rlabel metal2 849 -972 849 -972 0 net=4891
rlabel metal2 429 -974 429 -974 0 net=2307
rlabel metal2 590 -974 590 -974 0 net=4953
rlabel metal2 877 -974 877 -974 0 net=5089
rlabel metal2 457 -976 457 -976 0 net=3507
rlabel metal2 765 -976 765 -976 0 net=4259
rlabel metal2 758 -978 758 -978 0 net=3991
rlabel metal2 835 -978 835 -978 0 net=5251
rlabel metal2 65 -980 65 -980 0 net=4955
rlabel metal2 884 -980 884 -980 0 net=4505
rlabel metal2 933 -980 933 -980 0 net=5199
rlabel metal2 842 -982 842 -982 0 net=4585
rlabel metal2 842 -984 842 -984 0 net=5233
rlabel metal2 884 -986 884 -986 0 net=5173
rlabel metal2 926 -988 926 -988 0 net=4353
rlabel metal2 940 -990 940 -990 0 net=5855
rlabel metal2 912 -992 912 -992 0 net=5079
rlabel metal2 604 -994 604 -994 0 net=5547
rlabel metal2 9 -1005 9 -1005 0 net=2398
rlabel metal2 100 -1005 100 -1005 0 net=923
rlabel metal2 121 -1005 121 -1005 0 net=1473
rlabel metal2 359 -1005 359 -1005 0 net=2896
rlabel metal2 464 -1005 464 -1005 0 net=3050
rlabel metal2 541 -1005 541 -1005 0 net=3992
rlabel metal2 810 -1005 810 -1005 0 net=5480
rlabel metal2 1003 -1005 1003 -1005 0 net=5081
rlabel metal2 1003 -1005 1003 -1005 0 net=5081
rlabel metal2 1129 -1005 1129 -1005 0 net=4214
rlabel metal2 1185 -1005 1185 -1005 0 net=5181
rlabel metal2 1185 -1005 1185 -1005 0 net=5181
rlabel metal2 23 -1007 23 -1007 0 net=2533
rlabel metal2 23 -1007 23 -1007 0 net=2533
rlabel metal2 37 -1007 37 -1007 0 net=1491
rlabel metal2 89 -1007 89 -1007 0 net=4814
rlabel metal2 884 -1007 884 -1007 0 net=5174
rlabel metal2 954 -1007 954 -1007 0 net=6444
rlabel metal2 1136 -1007 1136 -1007 0 net=3324
rlabel metal2 40 -1009 40 -1009 0 net=474
rlabel metal2 555 -1009 555 -1009 0 net=2951
rlabel metal2 555 -1009 555 -1009 0 net=2951
rlabel metal2 569 -1009 569 -1009 0 net=3858
rlabel metal2 625 -1009 625 -1009 0 net=4163
rlabel metal2 730 -1009 730 -1009 0 net=6060
rlabel metal2 44 -1011 44 -1011 0 net=2934
rlabel metal2 208 -1011 208 -1011 0 net=1804
rlabel metal2 219 -1011 219 -1011 0 net=1542
rlabel metal2 362 -1011 362 -1011 0 net=5816
rlabel metal2 1094 -1011 1094 -1011 0 net=3903
rlabel metal2 16 -1013 16 -1013 0 net=1905
rlabel metal2 51 -1013 51 -1013 0 net=1403
rlabel metal2 51 -1013 51 -1013 0 net=1403
rlabel metal2 58 -1013 58 -1013 0 net=4456
rlabel metal2 107 -1013 107 -1013 0 net=1765
rlabel metal2 401 -1013 401 -1013 0 net=1839
rlabel metal2 527 -1013 527 -1013 0 net=2969
rlabel metal2 597 -1013 597 -1013 0 net=4462
rlabel metal2 646 -1013 646 -1013 0 net=4041
rlabel metal2 681 -1013 681 -1013 0 net=1781
rlabel metal2 723 -1013 723 -1013 0 net=5253
rlabel metal2 856 -1013 856 -1013 0 net=5436
rlabel metal2 16 -1015 16 -1015 0 net=6149
rlabel metal2 124 -1015 124 -1015 0 net=5607
rlabel metal2 366 -1015 366 -1015 0 net=2237
rlabel metal2 366 -1015 366 -1015 0 net=2237
rlabel metal2 457 -1015 457 -1015 0 net=3509
rlabel metal2 600 -1015 600 -1015 0 net=4330
rlabel metal2 856 -1015 856 -1015 0 net=5091
rlabel metal2 884 -1015 884 -1015 0 net=5337
rlabel metal2 1024 -1015 1024 -1015 0 net=5488
rlabel metal2 1069 -1015 1069 -1015 0 net=3409
rlabel metal2 30 -1017 30 -1017 0 net=2605
rlabel metal2 254 -1017 254 -1017 0 net=3365
rlabel metal2 443 -1017 443 -1017 0 net=2375
rlabel metal2 499 -1017 499 -1017 0 net=5386
rlabel metal2 996 -1017 996 -1017 0 net=5885
rlabel metal2 30 -1019 30 -1019 0 net=1685
rlabel metal2 184 -1019 184 -1019 0 net=2747
rlabel metal2 289 -1019 289 -1019 0 net=1246
rlabel metal2 338 -1019 338 -1019 0 net=1727
rlabel metal2 429 -1019 429 -1019 0 net=2309
rlabel metal2 499 -1019 499 -1019 0 net=3621
rlabel metal2 604 -1019 604 -1019 0 net=4421
rlabel metal2 695 -1019 695 -1019 0 net=4207
rlabel metal2 751 -1019 751 -1019 0 net=4601
rlabel metal2 786 -1019 786 -1019 0 net=4965
rlabel metal2 859 -1019 859 -1019 0 net=6170
rlabel metal2 61 -1021 61 -1021 0 net=3192
rlabel metal2 632 -1021 632 -1021 0 net=3545
rlabel metal2 681 -1021 681 -1021 0 net=3939
rlabel metal2 698 -1021 698 -1021 0 net=4851
rlabel metal2 863 -1021 863 -1021 0 net=5207
rlabel metal2 905 -1021 905 -1021 0 net=6363
rlabel metal2 982 -1021 982 -1021 0 net=6425
rlabel metal2 65 -1023 65 -1023 0 net=4560
rlabel metal2 429 -1023 429 -1023 0 net=2737
rlabel metal2 502 -1023 502 -1023 0 net=6120
rlabel metal2 72 -1025 72 -1025 0 net=1069
rlabel metal2 289 -1025 289 -1025 0 net=1299
rlabel metal2 317 -1025 317 -1025 0 net=2249
rlabel metal2 471 -1025 471 -1025 0 net=3499
rlabel metal2 639 -1025 639 -1025 0 net=6020
rlabel metal2 79 -1027 79 -1027 0 net=1353
rlabel metal2 317 -1027 317 -1027 0 net=182
rlabel metal2 639 -1027 639 -1027 0 net=3665
rlabel metal2 660 -1027 660 -1027 0 net=4137
rlabel metal2 751 -1027 751 -1027 0 net=5577
rlabel metal2 968 -1027 968 -1027 0 net=5915
rlabel metal2 996 -1027 996 -1027 0 net=6289
rlabel metal2 1087 -1027 1087 -1027 0 net=6523
rlabel metal2 79 -1029 79 -1029 0 net=899
rlabel metal2 187 -1029 187 -1029 0 net=4704
rlabel metal2 786 -1029 786 -1029 0 net=4507
rlabel metal2 989 -1029 989 -1029 0 net=6465
rlabel metal2 1122 -1029 1122 -1029 0 net=6535
rlabel metal2 96 -1031 96 -1031 0 net=3727
rlabel metal2 408 -1031 408 -1031 0 net=1903
rlabel metal2 485 -1031 485 -1031 0 net=2613
rlabel metal2 649 -1031 649 -1031 0 net=4260
rlabel metal2 919 -1031 919 -1031 0 net=5364
rlabel metal2 86 -1033 86 -1033 0 net=2188
rlabel metal2 114 -1033 114 -1033 0 net=3175
rlabel metal2 191 -1033 191 -1033 0 net=823
rlabel metal2 205 -1033 205 -1033 0 net=3423
rlabel metal2 509 -1033 509 -1033 0 net=3150
rlabel metal2 653 -1033 653 -1033 0 net=4083
rlabel metal2 716 -1033 716 -1033 0 net=3977
rlabel metal2 891 -1033 891 -1033 0 net=5549
rlabel metal2 1010 -1033 1010 -1033 0 net=6525
rlabel metal2 2 -1035 2 -1035 0 net=3442
rlabel metal2 212 -1035 212 -1035 0 net=985
rlabel metal2 268 -1035 268 -1035 0 net=1598
rlabel metal2 376 -1035 376 -1035 0 net=5455
rlabel metal2 912 -1035 912 -1035 0 net=4355
rlabel metal2 1017 -1035 1017 -1035 0 net=6387
rlabel metal2 128 -1037 128 -1037 0 net=1219
rlabel metal2 128 -1037 128 -1037 0 net=1219
rlabel metal2 170 -1037 170 -1037 0 net=1633
rlabel metal2 331 -1037 331 -1037 0 net=4661
rlabel metal2 572 -1037 572 -1037 0 net=5657
rlabel metal2 177 -1039 177 -1039 0 net=879
rlabel metal2 226 -1039 226 -1039 0 net=1013
rlabel metal2 303 -1039 303 -1039 0 net=1313
rlabel metal2 373 -1039 373 -1039 0 net=3061
rlabel metal2 506 -1039 506 -1039 0 net=5261
rlabel metal2 716 -1039 716 -1039 0 net=4777
rlabel metal2 779 -1039 779 -1039 0 net=4831
rlabel metal2 821 -1039 821 -1039 0 net=4919
rlabel metal2 86 -1041 86 -1041 0 net=3209
rlabel metal2 233 -1041 233 -1041 0 net=1649
rlabel metal2 303 -1041 303 -1041 0 net=1387
rlabel metal2 380 -1041 380 -1041 0 net=3111
rlabel metal2 450 -1041 450 -1041 0 net=3483
rlabel metal2 660 -1041 660 -1041 0 net=3689
rlabel metal2 684 -1041 684 -1041 0 net=6008
rlabel metal2 117 -1043 117 -1043 0 net=1445
rlabel metal2 240 -1043 240 -1043 0 net=3223
rlabel metal2 401 -1043 401 -1043 0 net=1967
rlabel metal2 450 -1043 450 -1043 0 net=3999
rlabel metal2 667 -1043 667 -1043 0 net=4519
rlabel metal2 733 -1043 733 -1043 0 net=5522
rlabel metal2 1059 -1043 1059 -1043 0 net=5777
rlabel metal2 152 -1045 152 -1045 0 net=1811
rlabel metal2 415 -1045 415 -1045 0 net=2759
rlabel metal2 688 -1045 688 -1045 0 net=1994
rlabel metal2 842 -1045 842 -1045 0 net=5235
rlabel metal2 1031 -1045 1031 -1045 0 net=4275
rlabel metal2 156 -1047 156 -1047 0 net=1127
rlabel metal2 390 -1047 390 -1047 0 net=5259
rlabel metal2 156 -1049 156 -1049 0 net=1023
rlabel metal2 478 -1049 478 -1049 0 net=3433
rlabel metal2 534 -1049 534 -1049 0 net=4586
rlabel metal2 135 -1051 135 -1051 0 net=1341
rlabel metal2 201 -1051 201 -1051 0 net=5709
rlabel metal2 135 -1053 135 -1053 0 net=2715
rlabel metal2 345 -1053 345 -1053 0 net=2683
rlabel metal2 576 -1053 576 -1053 0 net=3953
rlabel metal2 709 -1053 709 -1053 0 net=4281
rlabel metal2 772 -1053 772 -1053 0 net=4727
rlabel metal2 814 -1053 814 -1053 0 net=4893
rlabel metal2 247 -1055 247 -1055 0 net=1439
rlabel metal2 345 -1055 345 -1055 0 net=1579
rlabel metal2 576 -1055 576 -1055 0 net=3829
rlabel metal2 744 -1055 744 -1055 0 net=4847
rlabel metal2 849 -1055 849 -1055 0 net=6073
rlabel metal2 247 -1057 247 -1057 0 net=1175
rlabel metal2 352 -1057 352 -1057 0 net=4954
rlabel metal2 618 -1057 618 -1057 0 net=5200
rlabel metal2 520 -1059 520 -1059 0 net=3845
rlabel metal2 758 -1059 758 -1059 0 net=4957
rlabel metal2 173 -1061 173 -1061 0 net=4119
rlabel metal2 800 -1061 800 -1061 0 net=3869
rlabel metal2 940 -1063 940 -1063 0 net=5857
rlabel metal2 940 -1065 940 -1065 0 net=5825
rlabel metal2 961 -1067 961 -1067 0 net=5987
rlabel metal2 61 -1069 61 -1069 0 net=6135
rlabel metal2 16 -1080 16 -1080 0 net=6150
rlabel metal2 219 -1080 219 -1080 0 net=2606
rlabel metal2 471 -1080 471 -1080 0 net=3425
rlabel metal2 632 -1080 632 -1080 0 net=4208
rlabel metal2 852 -1080 852 -1080 0 net=3978
rlabel metal2 884 -1080 884 -1080 0 net=5339
rlabel metal2 912 -1080 912 -1080 0 net=4357
rlabel metal2 912 -1080 912 -1080 0 net=4357
rlabel metal2 954 -1080 954 -1080 0 net=5989
rlabel metal2 978 -1080 978 -1080 0 net=6388
rlabel metal2 1031 -1080 1031 -1080 0 net=6199
rlabel metal2 1041 -1080 1041 -1080 0 net=4276
rlabel metal2 1108 -1080 1108 -1080 0 net=6537
rlabel metal2 1185 -1080 1185 -1080 0 net=5182
rlabel metal2 23 -1082 23 -1082 0 net=2534
rlabel metal2 170 -1082 170 -1082 0 net=3846
rlabel metal2 600 -1082 600 -1082 0 net=6543
rlabel metal2 856 -1082 856 -1082 0 net=5093
rlabel metal2 856 -1082 856 -1082 0 net=5093
rlabel metal2 877 -1082 877 -1082 0 net=5659
rlabel metal2 940 -1082 940 -1082 0 net=5827
rlabel metal2 996 -1082 996 -1082 0 net=6291
rlabel metal2 996 -1082 996 -1082 0 net=6291
rlabel metal2 1006 -1082 1006 -1082 0 net=3904
rlabel metal2 30 -1084 30 -1084 0 net=1686
rlabel metal2 268 -1084 268 -1084 0 net=1634
rlabel metal2 345 -1084 345 -1084 0 net=1581
rlabel metal2 345 -1084 345 -1084 0 net=1581
rlabel metal2 355 -1084 355 -1084 0 net=4397
rlabel metal2 607 -1084 607 -1084 0 net=5578
rlabel metal2 884 -1084 884 -1084 0 net=5457
rlabel metal2 940 -1084 940 -1084 0 net=5859
rlabel metal2 1017 -1084 1017 -1084 0 net=5887
rlabel metal2 1045 -1084 1045 -1084 0 net=1783
rlabel metal2 30 -1086 30 -1086 0 net=1907
rlabel metal2 51 -1086 51 -1086 0 net=1405
rlabel metal2 51 -1086 51 -1086 0 net=1405
rlabel metal2 58 -1086 58 -1086 0 net=935
rlabel metal2 170 -1086 170 -1086 0 net=1129
rlabel metal2 191 -1086 191 -1086 0 net=881
rlabel metal2 247 -1086 247 -1086 0 net=1177
rlabel metal2 275 -1086 275 -1086 0 net=1014
rlabel metal2 509 -1086 509 -1086 0 net=6074
rlabel metal2 891 -1086 891 -1086 0 net=5551
rlabel metal2 947 -1086 947 -1086 0 net=5083
rlabel metal2 1010 -1086 1010 -1086 0 net=6527
rlabel metal2 1048 -1086 1048 -1086 0 net=6524
rlabel metal2 37 -1088 37 -1088 0 net=1492
rlabel metal2 387 -1088 387 -1088 0 net=3366
rlabel metal2 485 -1088 485 -1088 0 net=2614
rlabel metal2 639 -1088 639 -1088 0 net=3667
rlabel metal2 639 -1088 639 -1088 0 net=3667
rlabel metal2 660 -1088 660 -1088 0 net=3691
rlabel metal2 660 -1088 660 -1088 0 net=3691
rlabel metal2 667 -1088 667 -1088 0 net=4521
rlabel metal2 989 -1088 989 -1088 0 net=6467
rlabel metal2 1080 -1088 1080 -1088 0 net=3411
rlabel metal2 37 -1090 37 -1090 0 net=1221
rlabel metal2 149 -1090 149 -1090 0 net=1025
rlabel metal2 177 -1090 177 -1090 0 net=987
rlabel metal2 254 -1090 254 -1090 0 net=1651
rlabel metal2 254 -1090 254 -1090 0 net=1651
rlabel metal2 296 -1090 296 -1090 0 net=3954
rlabel metal2 621 -1090 621 -1090 0 net=3459
rlabel metal2 667 -1090 667 -1090 0 net=5260
rlabel metal2 982 -1090 982 -1090 0 net=6427
rlabel metal2 1073 -1090 1073 -1090 0 net=5779
rlabel metal2 44 -1092 44 -1092 0 net=4001
rlabel metal2 551 -1092 551 -1092 0 net=3830
rlabel metal2 586 -1092 586 -1092 0 net=5789
rlabel metal2 968 -1092 968 -1092 0 net=5917
rlabel metal2 65 -1094 65 -1094 0 net=1231
rlabel metal2 72 -1094 72 -1094 0 net=1070
rlabel metal2 499 -1094 499 -1094 0 net=3623
rlabel metal2 590 -1094 590 -1094 0 net=4139
rlabel metal2 842 -1094 842 -1094 0 net=5237
rlabel metal2 968 -1094 968 -1094 0 net=6137
rlabel metal2 72 -1096 72 -1096 0 net=2587
rlabel metal2 93 -1096 93 -1096 0 net=925
rlabel metal2 121 -1096 121 -1096 0 net=1475
rlabel metal2 366 -1096 366 -1096 0 net=2239
rlabel metal2 499 -1096 499 -1096 0 net=2953
rlabel metal2 572 -1096 572 -1096 0 net=3500
rlabel metal2 604 -1096 604 -1096 0 net=4423
rlabel metal2 670 -1096 670 -1096 0 net=6599
rlabel metal2 79 -1098 79 -1098 0 net=900
rlabel metal2 156 -1098 156 -1098 0 net=401
rlabel metal2 583 -1098 583 -1098 0 net=4084
rlabel metal2 674 -1098 674 -1098 0 net=3547
rlabel metal2 674 -1098 674 -1098 0 net=3547
rlabel metal2 681 -1098 681 -1098 0 net=3941
rlabel metal2 702 -1098 702 -1098 0 net=5263
rlabel metal2 100 -1100 100 -1100 0 net=1145
rlabel metal2 121 -1100 121 -1100 0 net=2749
rlabel metal2 191 -1100 191 -1100 0 net=1441
rlabel metal2 359 -1100 359 -1100 0 net=5609
rlabel metal2 709 -1100 709 -1100 0 net=4283
rlabel metal2 184 -1102 184 -1102 0 net=520
rlabel metal2 422 -1102 422 -1102 0 net=2251
rlabel metal2 534 -1102 534 -1102 0 net=3251
rlabel metal2 212 -1104 212 -1104 0 net=1315
rlabel metal2 373 -1104 373 -1104 0 net=3063
rlabel metal2 646 -1104 646 -1104 0 net=4043
rlabel metal2 226 -1106 226 -1106 0 net=3211
rlabel metal2 387 -1106 387 -1106 0 net=1841
rlabel metal2 646 -1106 646 -1106 0 net=2105
rlabel metal2 226 -1108 226 -1108 0 net=2211
rlabel metal2 282 -1108 282 -1108 0 net=1355
rlabel metal2 338 -1108 338 -1108 0 net=1729
rlabel metal2 422 -1108 422 -1108 0 net=2103
rlabel metal2 688 -1108 688 -1108 0 net=5254
rlabel metal2 919 -1108 919 -1108 0 net=5711
rlabel metal2 240 -1110 240 -1110 0 net=3225
rlabel metal2 436 -1110 436 -1110 0 net=3434
rlabel metal2 513 -1110 513 -1110 0 net=3511
rlabel metal2 562 -1110 562 -1110 0 net=3485
rlabel metal2 688 -1110 688 -1110 0 net=3871
rlabel metal2 933 -1110 933 -1110 0 net=379
rlabel metal2 240 -1112 240 -1112 0 net=1091
rlabel metal2 723 -1112 723 -1112 0 net=4959
rlabel metal2 1003 -1112 1003 -1112 0 net=5185
rlabel metal2 275 -1114 275 -1114 0 net=1973
rlabel metal2 289 -1114 289 -1114 0 net=1301
rlabel metal2 317 -1114 317 -1114 0 net=1911
rlabel metal2 800 -1114 800 -1114 0 net=4895
rlabel metal2 821 -1114 821 -1114 0 net=4921
rlabel metal2 233 -1116 233 -1116 0 net=1447
rlabel metal2 303 -1116 303 -1116 0 net=1389
rlabel metal2 331 -1116 331 -1116 0 net=2555
rlabel metal2 443 -1116 443 -1116 0 net=2311
rlabel metal2 492 -1116 492 -1116 0 net=2685
rlabel metal2 744 -1116 744 -1116 0 net=4849
rlabel metal2 163 -1118 163 -1118 0 net=1343
rlabel metal2 338 -1118 338 -1118 0 net=2761
rlabel metal2 429 -1118 429 -1118 0 net=2739
rlabel metal2 527 -1118 527 -1118 0 net=2971
rlabel metal2 744 -1118 744 -1118 0 net=5209
rlabel metal2 401 -1120 401 -1120 0 net=1969
rlabel metal2 450 -1120 450 -1120 0 net=2377
rlabel metal2 478 -1120 478 -1120 0 net=3519
rlabel metal2 814 -1120 814 -1120 0 net=4967
rlabel metal2 205 -1122 205 -1122 0 net=2147
rlabel metal2 541 -1122 541 -1122 0 net=4165
rlabel metal2 653 -1122 653 -1122 0 net=5069
rlabel metal2 198 -1124 198 -1124 0 net=825
rlabel metal2 261 -1124 261 -1124 0 net=2109
rlabel metal2 408 -1124 408 -1124 0 net=1904
rlabel metal2 793 -1124 793 -1124 0 net=4853
rlabel metal2 261 -1126 261 -1126 0 net=1813
rlabel metal2 779 -1126 779 -1126 0 net=4833
rlabel metal2 310 -1128 310 -1128 0 net=1869
rlabel metal2 772 -1130 772 -1130 0 net=4729
rlabel metal2 810 -1130 810 -1130 0 net=6364
rlabel metal2 758 -1132 758 -1132 0 net=5863
rlabel metal2 786 -1132 786 -1132 0 net=4509
rlabel metal2 716 -1134 716 -1134 0 net=4779
rlabel metal2 520 -1136 520 -1136 0 net=4121
rlabel metal2 758 -1136 758 -1136 0 net=4603
rlabel metal2 520 -1138 520 -1138 0 net=1705
rlabel metal2 548 -1140 548 -1140 0 net=4663
rlabel metal2 394 -1142 394 -1142 0 net=3728
rlabel metal2 380 -1144 380 -1144 0 net=3113
rlabel metal2 107 -1146 107 -1146 0 net=1767
rlabel metal2 107 -1148 107 -1148 0 net=3177
rlabel metal2 135 -1150 135 -1150 0 net=2717
rlabel metal2 135 -1152 135 -1152 0 net=4469
rlabel metal2 16 -1163 16 -1163 0 net=2751
rlabel metal2 142 -1163 142 -1163 0 net=2719
rlabel metal2 142 -1163 142 -1163 0 net=2719
rlabel metal2 149 -1163 149 -1163 0 net=1026
rlabel metal2 170 -1163 170 -1163 0 net=1130
rlabel metal2 205 -1163 205 -1163 0 net=827
rlabel metal2 205 -1163 205 -1163 0 net=827
rlabel metal2 219 -1163 219 -1163 0 net=883
rlabel metal2 219 -1163 219 -1163 0 net=883
rlabel metal2 226 -1163 226 -1163 0 net=1179
rlabel metal2 285 -1163 285 -1163 0 net=1390
rlabel metal2 331 -1163 331 -1163 0 net=1477
rlabel metal2 422 -1163 422 -1163 0 net=2104
rlabel metal2 422 -1163 422 -1163 0 net=2104
rlabel metal2 446 -1163 446 -1163 0 net=5413
rlabel metal2 975 -1163 975 -1163 0 net=6200
rlabel metal2 1066 -1163 1066 -1163 0 net=5187
rlabel metal2 23 -1165 23 -1165 0 net=383
rlabel metal2 30 -1165 30 -1165 0 net=1908
rlabel metal2 163 -1165 163 -1165 0 net=2213
rlabel metal2 254 -1165 254 -1165 0 net=1652
rlabel metal2 695 -1165 695 -1165 0 net=3943
rlabel metal2 828 -1165 828 -1165 0 net=4922
rlabel metal2 961 -1165 961 -1165 0 net=5829
rlabel metal2 982 -1165 982 -1165 0 net=5919
rlabel metal2 982 -1165 982 -1165 0 net=5919
rlabel metal2 989 -1165 989 -1165 0 net=6429
rlabel metal2 1080 -1165 1080 -1165 0 net=5781
rlabel metal2 30 -1167 30 -1167 0 net=2955
rlabel metal2 506 -1167 506 -1167 0 net=3064
rlabel metal2 562 -1167 562 -1167 0 net=2686
rlabel metal2 618 -1167 618 -1167 0 net=3426
rlabel metal2 667 -1167 667 -1167 0 net=3873
rlabel metal2 695 -1167 695 -1167 0 net=4665
rlabel metal2 831 -1167 831 -1167 0 net=5660
rlabel metal2 884 -1167 884 -1167 0 net=5459
rlabel metal2 996 -1167 996 -1167 0 net=6293
rlabel metal2 1010 -1167 1010 -1167 0 net=6469
rlabel metal2 1087 -1167 1087 -1167 0 net=3413
rlabel metal2 37 -1169 37 -1169 0 net=1222
rlabel metal2 152 -1169 152 -1169 0 net=3520
rlabel metal2 499 -1169 499 -1169 0 net=2417
rlabel metal2 544 -1169 544 -1169 0 net=5201
rlabel metal2 905 -1169 905 -1169 0 net=4511
rlabel metal2 905 -1169 905 -1169 0 net=4511
rlabel metal2 919 -1169 919 -1169 0 net=5713
rlabel metal2 1024 -1169 1024 -1169 0 net=6529
rlabel metal2 1101 -1169 1101 -1169 0 net=6539
rlabel metal2 37 -1171 37 -1171 0 net=2513
rlabel metal2 730 -1171 730 -1171 0 net=6545
rlabel metal2 44 -1173 44 -1173 0 net=4002
rlabel metal2 117 -1173 117 -1173 0 net=1997
rlabel metal2 170 -1173 170 -1173 0 net=1975
rlabel metal2 352 -1173 352 -1173 0 net=3581
rlabel metal2 607 -1173 607 -1173 0 net=5017
rlabel metal2 926 -1173 926 -1173 0 net=5791
rlabel metal2 58 -1175 58 -1175 0 net=937
rlabel metal2 177 -1175 177 -1175 0 net=989
rlabel metal2 229 -1175 229 -1175 0 net=3226
rlabel metal2 443 -1175 443 -1175 0 net=6015
rlabel metal2 1031 -1175 1031 -1175 0 net=6601
rlabel metal2 51 -1177 51 -1177 0 net=1406
rlabel metal2 72 -1177 72 -1177 0 net=2589
rlabel metal2 184 -1177 184 -1177 0 net=1583
rlabel metal2 359 -1177 359 -1177 0 net=1769
rlabel metal2 478 -1177 478 -1177 0 net=2313
rlabel metal2 562 -1177 562 -1177 0 net=4850
rlabel metal2 842 -1177 842 -1177 0 net=5239
rlabel metal2 954 -1177 954 -1177 0 net=5991
rlabel metal2 1017 -1177 1017 -1177 0 net=5889
rlabel metal2 1059 -1177 1059 -1177 0 net=1785
rlabel metal2 65 -1179 65 -1179 0 net=1233
rlabel metal2 79 -1179 79 -1179 0 net=1209
rlabel metal2 586 -1179 586 -1179 0 net=4960
rlabel metal2 730 -1179 730 -1179 0 net=4835
rlabel metal2 814 -1179 814 -1179 0 net=4969
rlabel metal2 849 -1179 849 -1179 0 net=5341
rlabel metal2 940 -1179 940 -1179 0 net=5861
rlabel metal2 51 -1181 51 -1181 0 net=2847
rlabel metal2 82 -1181 82 -1181 0 net=2762
rlabel metal2 429 -1181 429 -1181 0 net=1971
rlabel metal2 590 -1181 590 -1181 0 net=4141
rlabel metal2 625 -1181 625 -1181 0 net=6483
rlabel metal2 89 -1183 89 -1183 0 net=2687
rlabel metal2 187 -1183 187 -1183 0 net=4609
rlabel metal2 863 -1183 863 -1183 0 net=4854
rlabel metal2 93 -1185 93 -1185 0 net=927
rlabel metal2 93 -1185 93 -1185 0 net=927
rlabel metal2 100 -1185 100 -1185 0 net=1147
rlabel metal2 100 -1185 100 -1185 0 net=1147
rlabel metal2 107 -1185 107 -1185 0 net=3179
rlabel metal2 429 -1185 429 -1185 0 net=2107
rlabel metal2 653 -1185 653 -1185 0 net=4122
rlabel metal2 765 -1185 765 -1185 0 net=5095
rlabel metal2 870 -1185 870 -1185 0 net=5265
rlabel metal2 968 -1185 968 -1185 0 net=6139
rlabel metal2 61 -1187 61 -1187 0 net=5661
rlabel metal2 107 -1189 107 -1189 0 net=2085
rlabel metal2 450 -1189 450 -1189 0 net=2379
rlabel metal2 565 -1189 565 -1189 0 net=4999
rlabel metal2 891 -1189 891 -1189 0 net=4359
rlabel metal2 233 -1191 233 -1191 0 net=1345
rlabel metal2 306 -1191 306 -1191 0 net=4431
rlabel metal2 401 -1191 401 -1191 0 net=2111
rlabel metal2 569 -1191 569 -1191 0 net=3487
rlabel metal2 625 -1191 625 -1191 0 net=3669
rlabel metal2 646 -1191 646 -1191 0 net=3549
rlabel metal2 688 -1191 688 -1191 0 net=4605
rlabel metal2 772 -1191 772 -1191 0 net=5865
rlabel metal2 131 -1193 131 -1193 0 net=4463
rlabel metal2 772 -1193 772 -1193 0 net=6687
rlabel metal2 233 -1195 233 -1195 0 net=4003
rlabel metal2 555 -1195 555 -1195 0 net=2985
rlabel metal2 611 -1195 611 -1195 0 net=4425
rlabel metal2 898 -1195 898 -1195 0 net=5553
rlabel metal2 240 -1197 240 -1197 0 net=1093
rlabel metal2 254 -1197 254 -1197 0 net=1133
rlabel metal2 898 -1197 898 -1197 0 net=5085
rlabel metal2 240 -1199 240 -1199 0 net=1449
rlabel metal2 317 -1199 317 -1199 0 net=4317
rlabel metal2 744 -1199 744 -1199 0 net=5211
rlabel metal2 261 -1201 261 -1201 0 net=1815
rlabel metal2 289 -1201 289 -1201 0 net=1303
rlabel metal2 394 -1201 394 -1201 0 net=3115
rlabel metal2 597 -1201 597 -1201 0 net=4399
rlabel metal2 779 -1201 779 -1201 0 net=4731
rlabel metal2 166 -1203 166 -1203 0 net=6239
rlabel metal2 408 -1203 408 -1203 0 net=4471
rlabel metal2 786 -1203 786 -1203 0 net=4781
rlabel metal2 800 -1203 800 -1203 0 net=4897
rlabel metal2 212 -1205 212 -1205 0 net=1317
rlabel metal2 408 -1205 408 -1205 0 net=2149
rlabel metal2 509 -1205 509 -1205 0 net=4531
rlabel metal2 191 -1207 191 -1207 0 net=1443
rlabel metal2 268 -1207 268 -1207 0 net=1871
rlabel metal2 457 -1207 457 -1207 0 net=2253
rlabel metal2 534 -1207 534 -1207 0 net=3253
rlabel metal2 611 -1207 611 -1207 0 net=3295
rlabel metal2 674 -1207 674 -1207 0 net=4285
rlabel metal2 751 -1207 751 -1207 0 net=4523
rlabel metal2 191 -1209 191 -1209 0 net=1707
rlabel metal2 527 -1209 527 -1209 0 net=2973
rlabel metal2 660 -1209 660 -1209 0 net=3693
rlabel metal2 751 -1209 751 -1209 0 net=5071
rlabel metal2 275 -1211 275 -1211 0 net=1731
rlabel metal2 464 -1211 464 -1211 0 net=2241
rlabel metal2 513 -1211 513 -1211 0 net=3513
rlabel metal2 527 -1211 527 -1211 0 net=4051
rlabel metal2 681 -1211 681 -1211 0 net=1913
rlabel metal2 23 -1213 23 -1213 0 net=2243
rlabel metal2 541 -1213 541 -1213 0 net=4167
rlabel metal2 310 -1215 310 -1215 0 net=1357
rlabel metal2 436 -1215 436 -1215 0 net=2557
rlabel metal2 681 -1215 681 -1215 0 net=4045
rlabel metal2 324 -1217 324 -1217 0 net=1843
rlabel metal2 436 -1217 436 -1217 0 net=2741
rlabel metal2 632 -1217 632 -1217 0 net=3460
rlabel metal2 492 -1219 492 -1219 0 net=2451
rlabel metal2 576 -1221 576 -1221 0 net=3625
rlabel metal2 702 -1221 702 -1221 0 net=5611
rlabel metal2 366 -1223 366 -1223 0 net=3213
rlabel metal2 366 -1225 366 -1225 0 net=4621
rlabel metal2 415 -1225 415 -1225 0 net=4095
rlabel metal2 415 -1227 415 -1227 0 net=3273
rlabel metal2 30 -1238 30 -1238 0 net=2956
rlabel metal2 569 -1238 569 -1238 0 net=210
rlabel metal2 772 -1238 772 -1238 0 net=4733
rlabel metal2 828 -1238 828 -1238 0 net=5862
rlabel metal2 1101 -1238 1101 -1238 0 net=6541
rlabel metal2 1101 -1238 1101 -1238 0 net=6541
rlabel metal2 47 -1240 47 -1240 0 net=633
rlabel metal2 180 -1240 180 -1240 0 net=2244
rlabel metal2 481 -1240 481 -1240 0 net=4426
rlabel metal2 866 -1240 866 -1240 0 net=4512
rlabel metal2 999 -1240 999 -1240 0 net=5890
rlabel metal2 68 -1242 68 -1242 0 net=1234
rlabel metal2 86 -1242 86 -1242 0 net=2215
rlabel metal2 177 -1242 177 -1242 0 net=829
rlabel metal2 212 -1242 212 -1242 0 net=1444
rlabel metal2 394 -1242 394 -1242 0 net=6240
rlabel metal2 807 -1242 807 -1242 0 net=3945
rlabel metal2 72 -1244 72 -1244 0 net=3785
rlabel metal2 394 -1244 394 -1244 0 net=5581
rlabel metal2 509 -1244 509 -1244 0 net=2974
rlabel metal2 541 -1244 541 -1244 0 net=3719
rlabel metal2 590 -1244 590 -1244 0 net=6140
rlabel metal2 93 -1246 93 -1246 0 net=928
rlabel metal2 100 -1246 100 -1246 0 net=1149
rlabel metal2 100 -1246 100 -1246 0 net=1149
rlabel metal2 114 -1246 114 -1246 0 net=2591
rlabel metal2 149 -1246 149 -1246 0 net=719
rlabel metal2 590 -1246 590 -1246 0 net=3489
rlabel metal2 625 -1246 625 -1246 0 net=3671
rlabel metal2 625 -1246 625 -1246 0 net=3671
rlabel metal2 642 -1246 642 -1246 0 net=4168
rlabel metal2 905 -1246 905 -1246 0 net=6531
rlabel metal2 1059 -1246 1059 -1246 0 net=3414
rlabel metal2 16 -1248 16 -1248 0 net=2752
rlabel metal2 163 -1248 163 -1248 0 net=1305
rlabel metal2 324 -1248 324 -1248 0 net=1844
rlabel metal2 387 -1248 387 -1248 0 net=2151
rlabel metal2 443 -1248 443 -1248 0 net=2315
rlabel metal2 544 -1248 544 -1248 0 net=1914
rlabel metal2 1017 -1248 1017 -1248 0 net=5792
rlabel metal2 117 -1250 117 -1250 0 net=1609
rlabel metal2 219 -1250 219 -1250 0 net=885
rlabel metal2 219 -1250 219 -1250 0 net=885
rlabel metal2 233 -1250 233 -1250 0 net=4004
rlabel metal2 548 -1250 548 -1250 0 net=5866
rlabel metal2 1052 -1250 1052 -1250 0 net=6715
rlabel metal2 128 -1252 128 -1252 0 net=991
rlabel metal2 205 -1252 205 -1252 0 net=1135
rlabel metal2 264 -1252 264 -1252 0 net=3582
rlabel metal2 373 -1252 373 -1252 0 net=2987
rlabel metal2 618 -1252 618 -1252 0 net=3847
rlabel metal2 656 -1252 656 -1252 0 net=5460
rlabel metal2 184 -1254 184 -1254 0 net=1585
rlabel metal2 289 -1254 289 -1254 0 net=1319
rlabel metal2 324 -1254 324 -1254 0 net=3427
rlabel metal2 478 -1254 478 -1254 0 net=4142
rlabel metal2 639 -1254 639 -1254 0 net=3875
rlabel metal2 677 -1254 677 -1254 0 net=4836
rlabel metal2 796 -1254 796 -1254 0 net=6497
rlabel metal2 961 -1254 961 -1254 0 net=6603
rlabel metal2 184 -1256 184 -1256 0 net=1181
rlabel metal2 233 -1256 233 -1256 0 net=1359
rlabel metal2 341 -1256 341 -1256 0 net=1972
rlabel metal2 604 -1256 604 -1256 0 net=3551
rlabel metal2 656 -1256 656 -1256 0 net=3694
rlabel metal2 807 -1256 807 -1256 0 net=5019
rlabel metal2 1087 -1256 1087 -1256 0 net=5189
rlabel metal2 156 -1258 156 -1258 0 net=939
rlabel metal2 240 -1258 240 -1258 0 net=1450
rlabel metal2 506 -1258 506 -1258 0 net=6247
rlabel metal2 572 -1258 572 -1258 0 net=4783
rlabel metal2 821 -1258 821 -1258 0 net=5365
rlabel metal2 152 -1260 152 -1260 0 net=955
rlabel metal2 191 -1260 191 -1260 0 net=1708
rlabel metal2 345 -1260 345 -1260 0 net=3181
rlabel metal2 404 -1260 404 -1260 0 net=2108
rlabel metal2 506 -1260 506 -1260 0 net=4053
rlabel metal2 548 -1260 548 -1260 0 net=3255
rlabel metal2 646 -1260 646 -1260 0 net=4287
rlabel metal2 709 -1260 709 -1260 0 net=5714
rlabel metal2 198 -1262 198 -1262 0 net=1927
rlabel metal2 254 -1262 254 -1262 0 net=1873
rlabel metal2 282 -1262 282 -1262 0 net=1817
rlabel metal2 352 -1262 352 -1262 0 net=3215
rlabel metal2 583 -1262 583 -1262 0 net=3443
rlabel metal2 709 -1262 709 -1262 0 net=4611
rlabel metal2 828 -1262 828 -1262 0 net=5213
rlabel metal2 121 -1264 121 -1264 0 net=1999
rlabel metal2 296 -1264 296 -1264 0 net=1347
rlabel metal2 310 -1264 310 -1264 0 net=3627
rlabel metal2 660 -1264 660 -1264 0 net=4409
rlabel metal2 723 -1264 723 -1264 0 net=6430
rlabel metal2 107 -1266 107 -1266 0 net=2087
rlabel metal2 268 -1266 268 -1266 0 net=1733
rlabel metal2 317 -1266 317 -1266 0 net=434
rlabel metal2 660 -1266 660 -1266 0 net=4047
rlabel metal2 723 -1266 723 -1266 0 net=4465
rlabel metal2 814 -1266 814 -1266 0 net=5099
rlabel metal2 1066 -1266 1066 -1266 0 net=1787
rlabel metal2 79 -1268 79 -1268 0 net=1211
rlabel metal2 366 -1268 366 -1268 0 net=4623
rlabel metal2 663 -1268 663 -1268 0 net=4782
rlabel metal2 835 -1268 835 -1268 0 net=5343
rlabel metal2 877 -1268 877 -1268 0 net=5555
rlabel metal2 79 -1270 79 -1270 0 net=2689
rlabel metal2 247 -1270 247 -1270 0 net=1095
rlabel metal2 376 -1270 376 -1270 0 net=2242
rlabel metal2 667 -1270 667 -1270 0 net=4097
rlabel metal2 730 -1270 730 -1270 0 net=4473
rlabel metal2 793 -1270 793 -1270 0 net=5086
rlabel metal2 912 -1270 912 -1270 0 net=6485
rlabel metal2 37 -1272 37 -1272 0 net=2515
rlabel metal2 247 -1272 247 -1272 0 net=1771
rlabel metal2 408 -1272 408 -1272 0 net=2113
rlabel metal2 464 -1272 464 -1272 0 net=6151
rlabel metal2 940 -1272 940 -1272 0 net=6471
rlabel metal2 1045 -1272 1045 -1272 0 net=6689
rlabel metal2 107 -1274 107 -1274 0 net=1977
rlabel metal2 359 -1274 359 -1274 0 net=2453
rlabel metal2 702 -1274 702 -1274 0 net=4319
rlabel metal2 751 -1274 751 -1274 0 net=5073
rlabel metal2 779 -1274 779 -1274 0 net=5203
rlabel metal2 142 -1276 142 -1276 0 net=2721
rlabel metal2 338 -1276 338 -1276 0 net=4433
rlabel metal2 695 -1276 695 -1276 0 net=4667
rlabel metal2 751 -1276 751 -1276 0 net=5097
rlabel metal2 849 -1276 849 -1276 0 net=5241
rlabel metal2 142 -1278 142 -1278 0 net=1479
rlabel metal2 338 -1278 338 -1278 0 net=2483
rlabel metal2 415 -1278 415 -1278 0 net=3275
rlabel metal2 695 -1278 695 -1278 0 net=4401
rlabel metal2 765 -1278 765 -1278 0 net=5613
rlabel metal2 303 -1280 303 -1280 0 net=2265
rlabel metal2 401 -1280 401 -1280 0 net=3117
rlabel metal2 429 -1280 429 -1280 0 net=2255
rlabel metal2 688 -1280 688 -1280 0 net=4607
rlabel metal2 856 -1280 856 -1280 0 net=4899
rlabel metal2 44 -1282 44 -1282 0 net=775
rlabel metal2 436 -1282 436 -1282 0 net=2743
rlabel metal2 688 -1282 688 -1282 0 net=4525
rlabel metal2 856 -1282 856 -1282 0 net=5415
rlabel metal2 954 -1282 954 -1282 0 net=5921
rlabel metal2 44 -1284 44 -1284 0 net=2849
rlabel metal2 436 -1284 436 -1284 0 net=3515
rlabel metal2 786 -1284 786 -1284 0 net=4971
rlabel metal2 884 -1284 884 -1284 0 net=5403
rlabel metal2 450 -1286 450 -1286 0 net=2381
rlabel metal2 520 -1286 520 -1286 0 net=3297
rlabel metal2 842 -1286 842 -1286 0 net=5267
rlabel metal2 933 -1286 933 -1286 0 net=6295
rlabel metal2 485 -1288 485 -1288 0 net=2559
rlabel metal2 562 -1288 562 -1288 0 net=1805
rlabel metal2 891 -1288 891 -1288 0 net=4361
rlabel metal2 1003 -1288 1003 -1288 0 net=6017
rlabel metal2 499 -1290 499 -1290 0 net=2419
rlabel metal2 800 -1290 800 -1290 0 net=4533
rlabel metal2 422 -1292 422 -1292 0 net=1505
rlabel metal2 800 -1292 800 -1292 0 net=5001
rlabel metal2 891 -1292 891 -1292 0 net=5993
rlabel metal2 870 -1294 870 -1294 0 net=5663
rlabel metal2 989 -1294 989 -1294 0 net=6547
rlabel metal2 926 -1296 926 -1296 0 net=6473
rlabel metal2 1080 -1296 1080 -1296 0 net=5783
rlabel metal2 968 -1298 968 -1298 0 net=5831
rlabel metal2 9 -1309 9 -1309 0 net=849
rlabel metal2 37 -1309 37 -1309 0 net=2593
rlabel metal2 135 -1309 135 -1309 0 net=2516
rlabel metal2 408 -1309 408 -1309 0 net=2114
rlabel metal2 499 -1309 499 -1309 0 net=2421
rlabel metal2 534 -1309 534 -1309 0 net=3490
rlabel metal2 611 -1309 611 -1309 0 net=3673
rlabel metal2 628 -1309 628 -1309 0 net=5695
rlabel metal2 922 -1309 922 -1309 0 net=5832
rlabel metal2 975 -1309 975 -1309 0 net=4362
rlabel metal2 996 -1309 996 -1309 0 net=6018
rlabel metal2 1020 -1309 1020 -1309 0 net=1788
rlabel metal2 1097 -1309 1097 -1309 0 net=6542
rlabel metal2 16 -1311 16 -1311 0 net=3787
rlabel metal2 93 -1311 93 -1311 0 net=1150
rlabel metal2 114 -1311 114 -1311 0 net=1409
rlabel metal2 212 -1311 212 -1311 0 net=1611
rlabel metal2 380 -1311 380 -1311 0 net=3183
rlabel metal2 614 -1311 614 -1311 0 net=5098
rlabel metal2 793 -1311 793 -1311 0 net=4534
rlabel metal2 1059 -1311 1059 -1311 0 net=5190
rlabel metal2 23 -1313 23 -1313 0 net=931
rlabel metal2 261 -1313 261 -1313 0 net=1586
rlabel metal2 380 -1313 380 -1313 0 net=1507
rlabel metal2 429 -1313 429 -1313 0 net=2256
rlabel metal2 471 -1313 471 -1313 0 net=3277
rlabel metal2 527 -1313 527 -1313 0 net=4625
rlabel metal2 793 -1313 793 -1313 0 net=3947
rlabel metal2 1066 -1313 1066 -1313 0 net=5785
rlabel metal2 44 -1315 44 -1315 0 net=2851
rlabel metal2 44 -1315 44 -1315 0 net=2851
rlabel metal2 51 -1315 51 -1315 0 net=1773
rlabel metal2 268 -1315 268 -1315 0 net=1734
rlabel metal2 310 -1315 310 -1315 0 net=3628
rlabel metal2 625 -1315 625 -1315 0 net=4320
rlabel metal2 726 -1315 726 -1315 0 net=266
rlabel metal2 1031 -1315 1031 -1315 0 net=6717
rlabel metal2 58 -1317 58 -1317 0 net=1259
rlabel metal2 555 -1317 555 -1317 0 net=6248
rlabel metal2 576 -1317 576 -1317 0 net=395
rlabel metal2 653 -1317 653 -1317 0 net=4608
rlabel metal2 863 -1317 863 -1317 0 net=6472
rlabel metal2 961 -1317 961 -1317 0 net=6605
rlabel metal2 68 -1319 68 -1319 0 net=467
rlabel metal2 408 -1319 408 -1319 0 net=2560
rlabel metal2 492 -1319 492 -1319 0 net=4435
rlabel metal2 541 -1319 541 -1319 0 net=3721
rlabel metal2 597 -1319 597 -1319 0 net=3553
rlabel metal2 667 -1319 667 -1319 0 net=4099
rlabel metal2 667 -1319 667 -1319 0 net=4099
rlabel metal2 677 -1319 677 -1319 0 net=4443
rlabel metal2 709 -1319 709 -1319 0 net=4613
rlabel metal2 821 -1319 821 -1319 0 net=5367
rlabel metal2 905 -1319 905 -1319 0 net=6533
rlabel metal2 999 -1319 999 -1319 0 net=6690
rlabel metal2 72 -1321 72 -1321 0 net=945
rlabel metal2 569 -1321 569 -1321 0 net=3905
rlabel metal2 681 -1321 681 -1321 0 net=4411
rlabel metal2 733 -1321 733 -1321 0 net=5614
rlabel metal2 870 -1321 870 -1321 0 net=5665
rlabel metal2 912 -1321 912 -1321 0 net=6487
rlabel metal2 93 -1323 93 -1323 0 net=486
rlabel metal2 506 -1323 506 -1323 0 net=4055
rlabel metal2 695 -1323 695 -1323 0 net=4403
rlabel metal2 695 -1323 695 -1323 0 net=4403
rlabel metal2 737 -1323 737 -1323 0 net=4785
rlabel metal2 758 -1323 758 -1323 0 net=5075
rlabel metal2 870 -1323 870 -1323 0 net=5405
rlabel metal2 891 -1323 891 -1323 0 net=5995
rlabel metal2 933 -1323 933 -1323 0 net=6297
rlabel metal2 100 -1325 100 -1325 0 net=3216
rlabel metal2 411 -1325 411 -1325 0 net=4169
rlabel metal2 723 -1325 723 -1325 0 net=4467
rlabel metal2 765 -1325 765 -1325 0 net=4973
rlabel metal2 877 -1325 877 -1325 0 net=5557
rlabel metal2 891 -1325 891 -1325 0 net=5585
rlabel metal2 128 -1327 128 -1327 0 net=993
rlabel metal2 268 -1327 268 -1327 0 net=1349
rlabel metal2 345 -1327 345 -1327 0 net=1819
rlabel metal2 422 -1327 422 -1327 0 net=2317
rlabel metal2 471 -1327 471 -1327 0 net=3299
rlabel metal2 527 -1327 527 -1327 0 net=3445
rlabel metal2 660 -1327 660 -1327 0 net=4049
rlabel metal2 86 -1329 86 -1329 0 net=2217
rlabel metal2 345 -1329 345 -1329 0 net=6571
rlabel metal2 86 -1331 86 -1331 0 net=1213
rlabel metal2 285 -1331 285 -1331 0 net=2909
rlabel metal2 506 -1331 506 -1331 0 net=6595
rlabel metal2 128 -1333 128 -1333 0 net=2455
rlabel metal2 366 -1333 366 -1333 0 net=2485
rlabel metal2 520 -1333 520 -1333 0 net=2891
rlabel metal2 716 -1333 716 -1333 0 net=4669
rlabel metal2 856 -1333 856 -1333 0 net=5417
rlabel metal2 933 -1333 933 -1333 0 net=6499
rlabel metal2 79 -1335 79 -1335 0 net=2691
rlabel metal2 366 -1335 366 -1335 0 net=2127
rlabel metal2 429 -1335 429 -1335 0 net=2383
rlabel metal2 572 -1335 572 -1335 0 net=4073
rlabel metal2 688 -1335 688 -1335 0 net=4527
rlabel metal2 723 -1335 723 -1335 0 net=5242
rlabel metal2 856 -1335 856 -1335 0 net=4901
rlabel metal2 79 -1337 79 -1337 0 net=1183
rlabel metal2 191 -1337 191 -1337 0 net=1137
rlabel metal2 212 -1337 212 -1337 0 net=2063
rlabel metal2 415 -1337 415 -1337 0 net=3119
rlabel metal2 572 -1337 572 -1337 0 net=4474
rlabel metal2 737 -1337 737 -1337 0 net=4735
rlabel metal2 835 -1337 835 -1337 0 net=5345
rlabel metal2 926 -1337 926 -1337 0 net=6475
rlabel metal2 170 -1339 170 -1339 0 net=2723
rlabel metal2 254 -1339 254 -1339 0 net=1875
rlabel metal2 310 -1339 310 -1339 0 net=2561
rlabel metal2 926 -1339 926 -1339 0 net=5923
rlabel metal2 163 -1341 163 -1341 0 net=1307
rlabel metal2 177 -1341 177 -1341 0 net=831
rlabel metal2 254 -1341 254 -1341 0 net=1509
rlabel metal2 583 -1341 583 -1341 0 net=3849
rlabel metal2 646 -1341 646 -1341 0 net=4289
rlabel metal2 954 -1341 954 -1341 0 net=6549
rlabel metal2 107 -1343 107 -1343 0 net=1979
rlabel metal2 177 -1343 177 -1343 0 net=2207
rlabel metal2 436 -1343 436 -1343 0 net=3517
rlabel metal2 478 -1343 478 -1343 0 net=3256
rlabel metal2 618 -1343 618 -1343 0 net=3877
rlabel metal2 646 -1343 646 -1343 0 net=6201
rlabel metal2 107 -1345 107 -1345 0 net=2033
rlabel metal2 180 -1345 180 -1345 0 net=940
rlabel metal2 275 -1345 275 -1345 0 net=1806
rlabel metal2 660 -1345 660 -1345 0 net=5204
rlabel metal2 898 -1345 898 -1345 0 net=6153
rlabel metal2 65 -1347 65 -1347 0 net=3729
rlabel metal2 779 -1347 779 -1347 0 net=5003
rlabel metal2 184 -1349 184 -1349 0 net=1929
rlabel metal2 226 -1349 226 -1349 0 net=1361
rlabel metal2 394 -1349 394 -1349 0 net=5583
rlabel metal2 194 -1351 194 -1351 0 net=886
rlabel metal2 233 -1351 233 -1351 0 net=1096
rlabel metal2 373 -1351 373 -1351 0 net=2989
rlabel metal2 436 -1351 436 -1351 0 net=2744
rlabel metal2 467 -1351 467 -1351 0 net=4113
rlabel metal2 800 -1351 800 -1351 0 net=5021
rlabel metal2 121 -1353 121 -1353 0 net=2089
rlabel metal2 341 -1353 341 -1353 0 net=2399
rlabel metal2 548 -1353 548 -1353 0 net=3955
rlabel metal2 807 -1353 807 -1353 0 net=5101
rlabel metal2 121 -1355 121 -1355 0 net=4807
rlabel metal2 198 -1355 198 -1355 0 net=3428
rlabel metal2 373 -1355 373 -1355 0 net=3097
rlabel metal2 814 -1355 814 -1355 0 net=5215
rlabel metal2 142 -1357 142 -1357 0 net=1481
rlabel metal2 439 -1357 439 -1357 0 net=5671
rlabel metal2 828 -1357 828 -1357 0 net=5269
rlabel metal2 142 -1359 142 -1359 0 net=5183
rlabel metal2 149 -1361 149 -1361 0 net=957
rlabel metal2 282 -1361 282 -1361 0 net=2001
rlabel metal2 635 -1361 635 -1361 0 net=5287
rlabel metal2 156 -1363 156 -1363 0 net=2153
rlabel metal2 331 -1365 331 -1365 0 net=2267
rlabel metal2 289 -1367 289 -1367 0 net=1321
rlabel metal2 289 -1369 289 -1369 0 net=6195
rlabel metal2 2 -1380 2 -1380 0 net=636
rlabel metal2 9 -1380 9 -1380 0 net=1411
rlabel metal2 142 -1380 142 -1380 0 net=2724
rlabel metal2 250 -1380 250 -1380 0 net=1350
rlabel metal2 369 -1380 369 -1380 0 net=4074
rlabel metal2 702 -1380 702 -1380 0 net=4445
rlabel metal2 737 -1380 737 -1380 0 net=4737
rlabel metal2 737 -1380 737 -1380 0 net=4737
rlabel metal2 849 -1380 849 -1380 0 net=5347
rlabel metal2 849 -1380 849 -1380 0 net=5347
rlabel metal2 996 -1380 996 -1380 0 net=6637
rlabel metal2 30 -1382 30 -1382 0 net=851
rlabel metal2 72 -1382 72 -1382 0 net=946
rlabel metal2 369 -1382 369 -1382 0 net=2892
rlabel metal2 530 -1382 530 -1382 0 net=4670
rlabel metal2 947 -1382 947 -1382 0 net=6477
rlabel metal2 1003 -1382 1003 -1382 0 net=6597
rlabel metal2 1031 -1382 1031 -1382 0 net=6719
rlabel metal2 1045 -1382 1045 -1382 0 net=5786
rlabel metal2 30 -1384 30 -1384 0 net=2853
rlabel metal2 72 -1384 72 -1384 0 net=1191
rlabel metal2 208 -1384 208 -1384 0 net=3184
rlabel metal2 611 -1384 611 -1384 0 net=3675
rlabel metal2 611 -1384 611 -1384 0 net=3675
rlabel metal2 618 -1384 618 -1384 0 net=3879
rlabel metal2 632 -1384 632 -1384 0 net=4057
rlabel metal2 681 -1384 681 -1384 0 net=4171
rlabel metal2 975 -1384 975 -1384 0 net=6489
rlabel metal2 1010 -1384 1010 -1384 0 net=6607
rlabel metal2 1055 -1384 1055 -1384 0 net=6495
rlabel metal2 79 -1386 79 -1386 0 net=1185
rlabel metal2 380 -1386 380 -1386 0 net=1508
rlabel metal2 443 -1386 443 -1386 0 net=2487
rlabel metal2 488 -1386 488 -1386 0 net=1661
rlabel metal2 509 -1386 509 -1386 0 net=3730
rlabel metal2 646 -1386 646 -1386 0 net=4468
rlabel metal2 786 -1386 786 -1386 0 net=5217
rlabel metal2 940 -1386 940 -1386 0 net=6203
rlabel metal2 982 -1386 982 -1386 0 net=6573
rlabel metal2 79 -1388 79 -1388 0 net=4809
rlabel metal2 128 -1388 128 -1388 0 net=2456
rlabel metal2 457 -1388 457 -1388 0 net=2400
rlabel metal2 499 -1388 499 -1388 0 net=2422
rlabel metal2 555 -1388 555 -1388 0 net=3723
rlabel metal2 653 -1388 653 -1388 0 net=6154
rlabel metal2 86 -1390 86 -1390 0 net=1214
rlabel metal2 513 -1390 513 -1390 0 net=3279
rlabel metal2 569 -1390 569 -1390 0 net=5879
rlabel metal2 961 -1390 961 -1390 0 net=6299
rlabel metal2 86 -1392 86 -1392 0 net=1455
rlabel metal2 366 -1392 366 -1392 0 net=4029
rlabel metal2 660 -1392 660 -1392 0 net=3949
rlabel metal2 912 -1392 912 -1392 0 net=5997
rlabel metal2 100 -1394 100 -1394 0 net=2035
rlabel metal2 114 -1394 114 -1394 0 net=2155
rlabel metal2 177 -1394 177 -1394 0 net=1139
rlabel metal2 198 -1394 198 -1394 0 net=2725
rlabel metal2 261 -1394 261 -1394 0 net=994
rlabel metal2 289 -1394 289 -1394 0 net=6197
rlabel metal2 93 -1396 93 -1396 0 net=3151
rlabel metal2 380 -1396 380 -1396 0 net=2129
rlabel metal2 408 -1396 408 -1396 0 net=3601
rlabel metal2 534 -1396 534 -1396 0 net=4437
rlabel metal2 604 -1396 604 -1396 0 net=3907
rlabel metal2 667 -1396 667 -1396 0 net=4101
rlabel metal2 702 -1396 702 -1396 0 net=4787
rlabel metal2 793 -1396 793 -1396 0 net=4133
rlabel metal2 912 -1396 912 -1396 0 net=5925
rlabel metal2 16 -1398 16 -1398 0 net=3789
rlabel metal2 121 -1398 121 -1398 0 net=811
rlabel metal2 537 -1398 537 -1398 0 net=5076
rlabel metal2 842 -1398 842 -1398 0 net=5289
rlabel metal2 128 -1400 128 -1400 0 net=5584
rlabel metal2 142 -1402 142 -1402 0 net=1309
rlabel metal2 212 -1402 212 -1402 0 net=2065
rlabel metal2 408 -1402 408 -1402 0 net=2069
rlabel metal2 667 -1402 667 -1402 0 net=4627
rlabel metal2 772 -1402 772 -1402 0 net=5023
rlabel metal2 821 -1402 821 -1402 0 net=5696
rlabel metal2 58 -1404 58 -1404 0 net=1261
rlabel metal2 219 -1404 219 -1404 0 net=2091
rlabel metal2 345 -1404 345 -1404 0 net=2995
rlabel metal2 541 -1404 541 -1404 0 net=6534
rlabel metal2 149 -1406 149 -1406 0 net=959
rlabel metal2 149 -1406 149 -1406 0 net=959
rlabel metal2 156 -1406 156 -1406 0 net=3957
rlabel metal2 569 -1406 569 -1406 0 net=3449
rlabel metal2 726 -1406 726 -1406 0 net=6500
rlabel metal2 135 -1408 135 -1408 0 net=1657
rlabel metal2 663 -1408 663 -1408 0 net=6133
rlabel metal2 205 -1410 205 -1410 0 net=833
rlabel metal2 226 -1410 226 -1410 0 net=1362
rlabel metal2 394 -1410 394 -1410 0 net=2991
rlabel metal2 394 -1410 394 -1410 0 net=2991
rlabel metal2 415 -1410 415 -1410 0 net=2209
rlabel metal2 450 -1410 450 -1410 0 net=3121
rlabel metal2 541 -1410 541 -1410 0 net=4615
rlabel metal2 751 -1410 751 -1410 0 net=4975
rlabel metal2 828 -1410 828 -1410 0 net=5271
rlabel metal2 891 -1410 891 -1410 0 net=5587
rlabel metal2 905 -1410 905 -1410 0 net=5667
rlabel metal2 107 -1412 107 -1412 0 net=1635
rlabel metal2 226 -1412 226 -1412 0 net=1511
rlabel metal2 366 -1412 366 -1412 0 net=5527
rlabel metal2 233 -1414 233 -1414 0 net=130
rlabel metal2 51 -1416 51 -1416 0 net=1775
rlabel metal2 240 -1416 240 -1416 0 net=1613
rlabel metal2 415 -1416 415 -1416 0 net=2319
rlabel metal2 429 -1416 429 -1416 0 net=2385
rlabel metal2 429 -1416 429 -1416 0 net=2385
rlabel metal2 439 -1416 439 -1416 0 net=3243
rlabel metal2 597 -1416 597 -1416 0 net=3555
rlabel metal2 796 -1416 796 -1416 0 net=6697
rlabel metal2 51 -1418 51 -1418 0 net=2269
rlabel metal2 450 -1418 450 -1418 0 net=5103
rlabel metal2 828 -1418 828 -1418 0 net=5559
rlabel metal2 58 -1420 58 -1420 0 net=1851
rlabel metal2 471 -1420 471 -1420 0 net=3301
rlabel metal2 520 -1420 520 -1420 0 net=3741
rlabel metal2 695 -1420 695 -1420 0 net=4405
rlabel metal2 779 -1420 779 -1420 0 net=5005
rlabel metal2 877 -1420 877 -1420 0 net=5419
rlabel metal2 247 -1422 247 -1422 0 net=1877
rlabel metal2 310 -1422 310 -1422 0 net=2563
rlabel metal2 387 -1422 387 -1422 0 net=3447
rlabel metal2 688 -1422 688 -1422 0 net=4291
rlabel metal2 709 -1422 709 -1422 0 net=4413
rlabel metal2 870 -1422 870 -1422 0 net=5407
rlabel metal2 254 -1424 254 -1424 0 net=2911
rlabel metal2 527 -1424 527 -1424 0 net=5184
rlabel metal2 863 -1424 863 -1424 0 net=5369
rlabel metal2 138 -1426 138 -1426 0 net=5303
rlabel metal2 303 -1428 303 -1428 0 net=1483
rlabel metal2 348 -1428 348 -1428 0 net=5111
rlabel metal2 310 -1430 310 -1430 0 net=1323
rlabel metal2 464 -1430 464 -1430 0 net=3518
rlabel metal2 628 -1430 628 -1430 0 net=5957
rlabel metal2 716 -1430 716 -1430 0 net=4529
rlabel metal2 779 -1430 779 -1430 0 net=4903
rlabel metal2 331 -1432 331 -1432 0 net=1821
rlabel metal2 359 -1432 359 -1432 0 net=2693
rlabel metal2 576 -1432 576 -1432 0 net=5673
rlabel metal2 23 -1434 23 -1434 0 net=933
rlabel metal2 460 -1434 460 -1434 0 net=4385
rlabel metal2 23 -1436 23 -1436 0 net=1981
rlabel metal2 324 -1436 324 -1436 0 net=2003
rlabel metal2 576 -1436 576 -1436 0 net=3851
rlabel metal2 639 -1436 639 -1436 0 net=4115
rlabel metal2 163 -1438 163 -1438 0 net=1931
rlabel metal2 296 -1438 296 -1438 0 net=2219
rlabel metal2 583 -1438 583 -1438 0 net=1547
rlabel metal2 37 -1440 37 -1440 0 net=2595
rlabel metal2 296 -1440 296 -1440 0 net=3099
rlabel metal2 639 -1440 639 -1440 0 net=4050
rlabel metal2 373 -1442 373 -1442 0 net=5481
rlabel metal2 954 -1442 954 -1442 0 net=6551
rlabel metal2 495 -1444 495 -1444 0 net=6171
rlabel metal2 2 -1455 2 -1455 0 net=4947
rlabel metal2 68 -1455 68 -1455 0 net=2992
rlabel metal2 415 -1455 415 -1455 0 net=2321
rlabel metal2 415 -1455 415 -1455 0 net=2321
rlabel metal2 422 -1455 422 -1455 0 net=4134
rlabel metal2 824 -1455 824 -1455 0 net=6598
rlabel metal2 1045 -1455 1045 -1455 0 net=6639
rlabel metal2 9 -1457 9 -1457 0 net=1412
rlabel metal2 142 -1457 142 -1457 0 net=1310
rlabel metal2 310 -1457 310 -1457 0 net=1325
rlabel metal2 348 -1457 348 -1457 0 net=2210
rlabel metal2 457 -1457 457 -1457 0 net=6198
rlabel metal2 999 -1457 999 -1457 0 net=6720
rlabel metal2 1048 -1457 1048 -1457 0 net=4475
rlabel metal2 1059 -1457 1059 -1457 0 net=6496
rlabel metal2 19 -1459 19 -1459 0 net=1852
rlabel metal2 72 -1459 72 -1459 0 net=1192
rlabel metal2 142 -1459 142 -1459 0 net=1141
rlabel metal2 184 -1459 184 -1459 0 net=2597
rlabel metal2 352 -1459 352 -1459 0 net=934
rlabel metal2 506 -1459 506 -1459 0 net=1662
rlabel metal2 593 -1459 593 -1459 0 net=35
rlabel metal2 982 -1459 982 -1459 0 net=6609
rlabel metal2 23 -1461 23 -1461 0 net=1982
rlabel metal2 387 -1461 387 -1461 0 net=3448
rlabel metal2 509 -1461 509 -1461 0 net=3724
rlabel metal2 625 -1461 625 -1461 0 net=3881
rlabel metal2 632 -1461 632 -1461 0 net=4103
rlabel metal2 684 -1461 684 -1461 0 net=5528
rlabel metal2 23 -1463 23 -1463 0 net=6319
rlabel metal2 429 -1463 429 -1463 0 net=2387
rlabel metal2 429 -1463 429 -1463 0 net=2387
rlabel metal2 436 -1463 436 -1463 0 net=6134
rlabel metal2 30 -1465 30 -1465 0 net=2854
rlabel metal2 72 -1465 72 -1465 0 net=3281
rlabel metal2 604 -1465 604 -1465 0 net=3676
rlabel metal2 625 -1465 625 -1465 0 net=4387
rlabel metal2 744 -1465 744 -1465 0 net=3557
rlabel metal2 751 -1465 751 -1465 0 net=4977
rlabel metal2 751 -1465 751 -1465 0 net=4977
rlabel metal2 765 -1465 765 -1465 0 net=5304
rlabel metal2 37 -1467 37 -1467 0 net=853
rlabel metal2 93 -1467 93 -1467 0 net=3791
rlabel metal2 436 -1467 436 -1467 0 net=2695
rlabel metal2 520 -1467 520 -1467 0 net=4530
rlabel metal2 765 -1467 765 -1467 0 net=5371
rlabel metal2 44 -1469 44 -1469 0 net=2071
rlabel metal2 443 -1469 443 -1469 0 net=3451
rlabel metal2 607 -1469 607 -1469 0 net=4172
rlabel metal2 58 -1471 58 -1471 0 net=1699
rlabel metal2 450 -1471 450 -1471 0 net=5104
rlabel metal2 611 -1471 611 -1471 0 net=4059
rlabel metal2 681 -1471 681 -1471 0 net=5290
rlabel metal2 93 -1473 93 -1473 0 net=2523
rlabel metal2 191 -1473 191 -1473 0 net=2488
rlabel metal2 520 -1473 520 -1473 0 net=5880
rlabel metal2 96 -1475 96 -1475 0 net=5285
rlabel metal2 768 -1475 768 -1475 0 net=5560
rlabel metal2 856 -1475 856 -1475 0 net=5675
rlabel metal2 926 -1475 926 -1475 0 net=6205
rlabel metal2 100 -1477 100 -1477 0 net=2037
rlabel metal2 100 -1477 100 -1477 0 net=2037
rlabel metal2 128 -1477 128 -1477 0 net=1485
rlabel metal2 345 -1477 345 -1477 0 net=2997
rlabel metal2 464 -1477 464 -1477 0 net=3302
rlabel metal2 534 -1477 534 -1477 0 net=1658
rlabel metal2 635 -1477 635 -1477 0 net=3950
rlabel metal2 667 -1477 667 -1477 0 net=4629
rlabel metal2 709 -1477 709 -1477 0 net=5959
rlabel metal2 975 -1477 975 -1477 0 net=6479
rlabel metal2 149 -1479 149 -1479 0 net=961
rlabel metal2 149 -1479 149 -1479 0 net=961
rlabel metal2 163 -1479 163 -1479 0 net=1933
rlabel metal2 191 -1479 191 -1479 0 net=1615
rlabel metal2 247 -1479 247 -1479 0 net=1878
rlabel metal2 387 -1479 387 -1479 0 net=4031
rlabel metal2 660 -1479 660 -1479 0 net=4261
rlabel metal2 709 -1479 709 -1479 0 net=4739
rlabel metal2 744 -1479 744 -1479 0 net=4905
rlabel metal2 786 -1479 786 -1479 0 net=5219
rlabel metal2 786 -1479 786 -1479 0 net=5219
rlabel metal2 793 -1479 793 -1479 0 net=5998
rlabel metal2 163 -1481 163 -1481 0 net=2727
rlabel metal2 215 -1481 215 -1481 0 net=6179
rlabel metal2 639 -1481 639 -1481 0 net=4788
rlabel metal2 772 -1481 772 -1481 0 net=5025
rlabel metal2 793 -1481 793 -1481 0 net=5273
rlabel metal2 856 -1481 856 -1481 0 net=5589
rlabel metal2 170 -1483 170 -1483 0 net=1263
rlabel metal2 219 -1483 219 -1483 0 net=835
rlabel metal2 219 -1483 219 -1483 0 net=835
rlabel metal2 226 -1483 226 -1483 0 net=1513
rlabel metal2 261 -1483 261 -1483 0 net=2093
rlabel metal2 261 -1483 261 -1483 0 net=2093
rlabel metal2 268 -1483 268 -1483 0 net=1186
rlabel metal2 282 -1483 282 -1483 0 net=2221
rlabel metal2 373 -1483 373 -1483 0 net=6261
rlabel metal2 107 -1485 107 -1485 0 net=1637
rlabel metal2 233 -1485 233 -1485 0 net=1777
rlabel metal2 373 -1485 373 -1485 0 net=4675
rlabel metal2 544 -1485 544 -1485 0 net=5565
rlabel metal2 107 -1487 107 -1487 0 net=2535
rlabel metal2 548 -1487 548 -1487 0 net=3853
rlabel metal2 639 -1487 639 -1487 0 net=4293
rlabel metal2 702 -1487 702 -1487 0 net=6329
rlabel metal2 772 -1487 772 -1487 0 net=5007
rlabel metal2 814 -1487 814 -1487 0 net=5421
rlabel metal2 898 -1487 898 -1487 0 net=5669
rlabel metal2 68 -1489 68 -1489 0 net=5687
rlabel metal2 114 -1491 114 -1491 0 net=2157
rlabel metal2 275 -1491 275 -1491 0 net=2005
rlabel metal2 394 -1491 394 -1491 0 net=3245
rlabel metal2 642 -1491 642 -1491 0 net=5643
rlabel metal2 79 -1493 79 -1493 0 net=4810
rlabel metal2 121 -1493 121 -1493 0 net=813
rlabel metal2 194 -1493 194 -1493 0 net=4173
rlabel metal2 233 -1493 233 -1493 0 net=1823
rlabel metal2 359 -1493 359 -1493 0 net=2067
rlabel metal2 478 -1493 478 -1493 0 net=3743
rlabel metal2 653 -1493 653 -1493 0 net=4117
rlabel metal2 695 -1493 695 -1493 0 net=4639
rlabel metal2 796 -1493 796 -1493 0 net=5301
rlabel metal2 842 -1493 842 -1493 0 net=6552
rlabel metal2 51 -1495 51 -1495 0 net=2271
rlabel metal2 240 -1495 240 -1495 0 net=1391
rlabel metal2 541 -1495 541 -1495 0 net=4617
rlabel metal2 590 -1495 590 -1495 0 net=4439
rlabel metal2 807 -1495 807 -1495 0 net=5409
rlabel metal2 989 -1495 989 -1495 0 net=6301
rlabel metal2 51 -1497 51 -1497 0 net=2913
rlabel metal2 296 -1497 296 -1497 0 net=3101
rlabel metal2 492 -1497 492 -1497 0 net=3603
rlabel metal2 79 -1499 79 -1499 0 net=3959
rlabel metal2 254 -1499 254 -1499 0 net=1549
rlabel metal2 590 -1499 590 -1499 0 net=5112
rlabel metal2 877 -1499 877 -1499 0 net=6491
rlabel metal2 86 -1501 86 -1501 0 net=1457
rlabel metal2 278 -1501 278 -1501 0 net=4795
rlabel metal2 506 -1501 506 -1501 0 net=5437
rlabel metal2 905 -1501 905 -1501 0 net=6699
rlabel metal2 86 -1503 86 -1503 0 net=4155
rlabel metal2 296 -1503 296 -1503 0 net=3017
rlabel metal2 516 -1503 516 -1503 0 net=4553
rlabel metal2 747 -1503 747 -1503 0 net=1
rlabel metal2 16 -1505 16 -1505 0 net=4937
rlabel metal2 303 -1505 303 -1505 0 net=2131
rlabel metal2 541 -1505 541 -1505 0 net=6445
rlabel metal2 331 -1507 331 -1507 0 net=3303
rlabel metal2 555 -1507 555 -1507 0 net=4021
rlabel metal2 583 -1507 583 -1507 0 net=3909
rlabel metal2 821 -1507 821 -1507 0 net=4995
rlabel metal2 338 -1509 338 -1509 0 net=2565
rlabel metal2 646 -1509 646 -1509 0 net=4447
rlabel metal2 905 -1509 905 -1509 0 net=5927
rlabel metal2 338 -1511 338 -1511 0 net=1941
rlabel metal2 499 -1511 499 -1511 0 net=3123
rlabel metal2 912 -1511 912 -1511 0 net=6173
rlabel metal2 198 -1513 198 -1513 0 net=4265
rlabel metal2 954 -1513 954 -1513 0 net=6575
rlabel metal2 366 -1515 366 -1515 0 net=4407
rlabel metal2 800 -1515 800 -1515 0 net=4415
rlabel metal2 723 -1517 723 -1517 0 net=6583
rlabel metal2 800 -1519 800 -1519 0 net=5349
rlabel metal2 849 -1521 849 -1521 0 net=5483
rlabel metal2 471 -1523 471 -1523 0 net=5697
rlabel metal2 289 -1525 289 -1525 0 net=3153
rlabel metal2 30 -1527 30 -1527 0 net=3397
rlabel metal2 23 -1538 23 -1538 0 net=6320
rlabel metal2 152 -1538 152 -1538 0 net=5566
rlabel metal2 1017 -1538 1017 -1538 0 net=6303
rlabel metal2 1038 -1538 1038 -1538 0 net=6641
rlabel metal2 1052 -1538 1052 -1538 0 net=4476
rlabel metal2 1052 -1538 1052 -1538 0 net=4476
rlabel metal2 2 -1540 2 -1540 0 net=4949
rlabel metal2 30 -1540 30 -1540 0 net=3398
rlabel metal2 436 -1540 436 -1540 0 net=2697
rlabel metal2 436 -1540 436 -1540 0 net=2697
rlabel metal2 471 -1540 471 -1540 0 net=3155
rlabel metal2 471 -1540 471 -1540 0 net=3155
rlabel metal2 488 -1540 488 -1540 0 net=586
rlabel metal2 740 -1540 740 -1540 0 net=6610
rlabel metal2 30 -1542 30 -1542 0 net=2133
rlabel metal2 306 -1542 306 -1542 0 net=3585
rlabel metal2 520 -1542 520 -1542 0 net=3604
rlabel metal2 961 -1542 961 -1542 0 net=3599
rlabel metal2 37 -1544 37 -1544 0 net=855
rlabel metal2 37 -1544 37 -1544 0 net=855
rlabel metal2 68 -1544 68 -1544 0 net=4156
rlabel metal2 93 -1544 93 -1544 0 net=2323
rlabel metal2 527 -1544 527 -1544 0 net=3854
rlabel metal2 558 -1544 558 -1544 0 net=6480
rlabel metal2 68 -1546 68 -1546 0 net=5286
rlabel metal2 842 -1546 842 -1546 0 net=5689
rlabel metal2 79 -1548 79 -1548 0 net=3961
rlabel metal2 79 -1548 79 -1548 0 net=3961
rlabel metal2 86 -1548 86 -1548 0 net=2039
rlabel metal2 135 -1548 135 -1548 0 net=2095
rlabel metal2 289 -1548 289 -1548 0 net=4262
rlabel metal2 723 -1548 723 -1548 0 net=5423
rlabel metal2 877 -1548 877 -1548 0 net=6493
rlabel metal2 100 -1550 100 -1550 0 net=1639
rlabel metal2 247 -1550 247 -1550 0 net=1515
rlabel metal2 296 -1550 296 -1550 0 net=2068
rlabel metal2 366 -1550 366 -1550 0 net=4408
rlabel metal2 646 -1550 646 -1550 0 net=4449
rlabel metal2 646 -1550 646 -1550 0 net=4449
rlabel metal2 663 -1550 663 -1550 0 net=5302
rlabel metal2 884 -1550 884 -1550 0 net=3559
rlabel metal2 128 -1552 128 -1552 0 net=1487
rlabel metal2 324 -1552 324 -1552 0 net=1779
rlabel metal2 324 -1552 324 -1552 0 net=1779
rlabel metal2 373 -1552 373 -1552 0 net=4677
rlabel metal2 499 -1552 499 -1552 0 net=4267
rlabel metal2 565 -1552 565 -1552 0 net=5960
rlabel metal2 72 -1554 72 -1554 0 net=3283
rlabel metal2 534 -1554 534 -1554 0 net=4023
rlabel metal2 583 -1554 583 -1554 0 net=3911
rlabel metal2 684 -1554 684 -1554 0 net=6365
rlabel metal2 947 -1554 947 -1554 0 net=4417
rlabel metal2 16 -1556 16 -1556 0 net=4938
rlabel metal2 121 -1556 121 -1556 0 net=2273
rlabel metal2 156 -1556 156 -1556 0 net=1458
rlabel metal2 359 -1556 359 -1556 0 net=2489
rlabel metal2 583 -1556 583 -1556 0 net=4641
rlabel metal2 726 -1556 726 -1556 0 net=5670
rlabel metal2 121 -1558 121 -1558 0 net=2007
rlabel metal2 366 -1558 366 -1558 0 net=1949
rlabel metal2 590 -1558 590 -1558 0 net=5525
rlabel metal2 898 -1558 898 -1558 0 net=6447
rlabel metal2 44 -1560 44 -1560 0 net=2073
rlabel metal2 373 -1560 373 -1560 0 net=484
rlabel metal2 541 -1560 541 -1560 0 net=4061
rlabel metal2 618 -1560 618 -1560 0 net=4118
rlabel metal2 737 -1560 737 -1560 0 net=4997
rlabel metal2 44 -1562 44 -1562 0 net=1143
rlabel metal2 156 -1562 156 -1562 0 net=1942
rlabel metal2 355 -1562 355 -1562 0 net=6253
rlabel metal2 758 -1562 758 -1562 0 net=5351
rlabel metal2 814 -1562 814 -1562 0 net=5645
rlabel metal2 107 -1564 107 -1564 0 net=2537
rlabel metal2 380 -1564 380 -1564 0 net=2567
rlabel metal2 590 -1564 590 -1564 0 net=4295
rlabel metal2 800 -1564 800 -1564 0 net=5411
rlabel metal2 821 -1564 821 -1564 0 net=5485
rlabel metal2 863 -1564 863 -1564 0 net=6175
rlabel metal2 142 -1566 142 -1566 0 net=963
rlabel metal2 170 -1566 170 -1566 0 net=814
rlabel metal2 807 -1566 807 -1566 0 net=5677
rlabel metal2 912 -1566 912 -1566 0 net=6701
rlabel metal2 177 -1568 177 -1568 0 net=2525
rlabel metal2 387 -1568 387 -1568 0 net=4032
rlabel metal2 576 -1568 576 -1568 0 net=4619
rlabel metal2 660 -1568 660 -1568 0 net=5833
rlabel metal2 870 -1568 870 -1568 0 net=6207
rlabel metal2 177 -1570 177 -1570 0 net=1617
rlabel metal2 201 -1570 201 -1570 0 net=2598
rlabel metal2 401 -1570 401 -1570 0 net=3103
rlabel metal2 478 -1570 478 -1570 0 net=3745
rlabel metal2 562 -1570 562 -1570 0 net=6669
rlabel metal2 184 -1572 184 -1572 0 net=1935
rlabel metal2 184 -1572 184 -1572 0 net=1935
rlabel metal2 191 -1572 191 -1572 0 net=1265
rlabel metal2 212 -1572 212 -1572 0 net=4175
rlabel metal2 394 -1572 394 -1572 0 net=3247
rlabel metal2 576 -1572 576 -1572 0 net=4105
rlabel metal2 660 -1572 660 -1572 0 net=4555
rlabel metal2 205 -1574 205 -1574 0 net=1825
rlabel metal2 240 -1574 240 -1574 0 net=1392
rlabel metal2 401 -1574 401 -1574 0 net=2389
rlabel metal2 569 -1574 569 -1574 0 net=6181
rlabel metal2 688 -1574 688 -1574 0 net=4741
rlabel metal2 163 -1576 163 -1576 0 net=2729
rlabel metal2 240 -1576 240 -1576 0 net=3793
rlabel metal2 429 -1576 429 -1576 0 net=3019
rlabel metal2 604 -1576 604 -1576 0 net=4389
rlabel metal2 709 -1576 709 -1576 0 net=4907
rlabel metal2 58 -1578 58 -1578 0 net=1701
rlabel metal2 212 -1578 212 -1578 0 net=837
rlabel metal2 247 -1578 247 -1578 0 net=2223
rlabel metal2 345 -1578 345 -1578 0 net=2083
rlabel metal2 408 -1578 408 -1578 0 net=6330
rlabel metal2 744 -1578 744 -1578 0 net=5027
rlabel metal2 58 -1580 58 -1580 0 net=5387
rlabel metal2 408 -1580 408 -1580 0 net=3453
rlabel metal2 450 -1580 450 -1580 0 net=2999
rlabel metal2 597 -1580 597 -1580 0 net=4441
rlabel metal2 51 -1582 51 -1582 0 net=2915
rlabel metal2 618 -1582 618 -1582 0 net=4631
rlabel metal2 702 -1582 702 -1582 0 net=6263
rlabel metal2 51 -1584 51 -1584 0 net=2843
rlabel metal2 716 -1584 716 -1584 0 net=3883
rlabel metal2 114 -1586 114 -1586 0 net=3773
rlabel metal2 387 -1586 387 -1586 0 net=5175
rlabel metal2 716 -1586 716 -1586 0 net=4979
rlabel metal2 107 -1588 107 -1588 0 net=6567
rlabel metal2 117 -1588 117 -1588 0 net=3227
rlabel metal2 411 -1588 411 -1588 0 net=3124
rlabel metal2 751 -1588 751 -1588 0 net=5221
rlabel metal2 443 -1590 443 -1590 0 net=3859
rlabel metal2 730 -1590 730 -1590 0 net=5009
rlabel metal2 786 -1590 786 -1590 0 net=5591
rlabel metal2 492 -1592 492 -1592 0 net=4797
rlabel metal2 765 -1592 765 -1592 0 net=5373
rlabel metal2 856 -1592 856 -1592 0 net=283
rlabel metal2 331 -1594 331 -1594 0 net=3305
rlabel metal2 765 -1594 765 -1594 0 net=5275
rlabel metal2 317 -1596 317 -1596 0 net=1327
rlabel metal2 793 -1596 793 -1596 0 net=5439
rlabel metal2 268 -1598 268 -1598 0 net=2159
rlabel metal2 835 -1598 835 -1598 0 net=5699
rlabel metal2 254 -1600 254 -1600 0 net=1551
rlabel metal2 891 -1600 891 -1600 0 net=6577
rlabel metal2 254 -1602 254 -1602 0 net=2009
rlabel metal2 905 -1602 905 -1602 0 net=5929
rlabel metal2 905 -1604 905 -1604 0 net=6585
rlabel metal2 30 -1615 30 -1615 0 net=2134
rlabel metal2 366 -1615 366 -1615 0 net=1951
rlabel metal2 530 -1615 530 -1615 0 net=4442
rlabel metal2 926 -1615 926 -1615 0 net=6670
rlabel metal2 954 -1615 954 -1615 0 net=5931
rlabel metal2 1024 -1615 1024 -1615 0 net=6305
rlabel metal2 1024 -1615 1024 -1615 0 net=6305
rlabel metal2 1038 -1615 1038 -1615 0 net=6642
rlabel metal2 37 -1617 37 -1617 0 net=856
rlabel metal2 37 -1617 37 -1617 0 net=856
rlabel metal2 58 -1617 58 -1617 0 net=5388
rlabel metal2 310 -1617 310 -1617 0 net=3156
rlabel metal2 523 -1617 523 -1617 0 net=3912
rlabel metal2 681 -1617 681 -1617 0 net=4998
rlabel metal2 775 -1617 775 -1617 0 net=5834
rlabel metal2 65 -1619 65 -1619 0 net=6021
rlabel metal2 121 -1619 121 -1619 0 net=2008
rlabel metal2 310 -1619 310 -1619 0 net=5685
rlabel metal2 366 -1619 366 -1619 0 net=2391
rlabel metal2 425 -1619 425 -1619 0 net=6663
rlabel metal2 534 -1619 534 -1619 0 net=4025
rlabel metal2 534 -1619 534 -1619 0 net=4025
rlabel metal2 544 -1619 544 -1619 0 net=5440
rlabel metal2 68 -1621 68 -1621 0 net=3794
rlabel metal2 257 -1621 257 -1621 0 net=1780
rlabel metal2 352 -1621 352 -1621 0 net=3455
rlabel metal2 429 -1621 429 -1621 0 net=3020
rlabel metal2 551 -1621 551 -1621 0 net=4620
rlabel metal2 646 -1621 646 -1621 0 net=4451
rlabel metal2 681 -1621 681 -1621 0 net=5691
rlabel metal2 695 -1621 695 -1621 0 net=6494
rlabel metal2 72 -1623 72 -1623 0 net=40
rlabel metal2 562 -1623 562 -1623 0 net=360
rlabel metal2 79 -1625 79 -1625 0 net=3962
rlabel metal2 562 -1625 562 -1625 0 net=6265
rlabel metal2 723 -1625 723 -1625 0 net=5425
rlabel metal2 751 -1625 751 -1625 0 net=5223
rlabel metal2 79 -1627 79 -1627 0 net=220
rlabel metal2 261 -1627 261 -1627 0 net=1517
rlabel metal2 261 -1627 261 -1627 0 net=1517
rlabel metal2 268 -1627 268 -1627 0 net=1552
rlabel metal2 565 -1627 565 -1627 0 net=4632
rlabel metal2 688 -1627 688 -1627 0 net=4743
rlabel metal2 779 -1627 779 -1627 0 net=5486
rlabel metal2 107 -1629 107 -1629 0 net=3746
rlabel metal2 569 -1629 569 -1629 0 net=5646
rlabel metal2 93 -1631 93 -1631 0 net=2325
rlabel metal2 121 -1631 121 -1631 0 net=5451
rlabel metal2 163 -1631 163 -1631 0 net=1703
rlabel metal2 268 -1631 268 -1631 0 net=1553
rlabel metal2 513 -1631 513 -1631 0 net=711
rlabel metal2 93 -1633 93 -1633 0 net=2011
rlabel metal2 282 -1633 282 -1633 0 net=3228
rlabel metal2 569 -1633 569 -1633 0 net=6183
rlabel metal2 688 -1633 688 -1633 0 net=6208
rlabel metal2 128 -1635 128 -1635 0 net=2275
rlabel metal2 198 -1635 198 -1635 0 net=2084
rlabel metal2 376 -1635 376 -1635 0 net=2526
rlabel metal2 387 -1635 387 -1635 0 net=3861
rlabel metal2 576 -1635 576 -1635 0 net=4107
rlabel metal2 695 -1635 695 -1635 0 net=975
rlabel metal2 814 -1635 814 -1635 0 net=3885
rlabel metal2 114 -1637 114 -1637 0 net=6569
rlabel metal2 142 -1637 142 -1637 0 net=965
rlabel metal2 142 -1637 142 -1637 0 net=965
rlabel metal2 149 -1637 149 -1637 0 net=546
rlabel metal2 208 -1637 208 -1637 0 net=6141
rlabel metal2 443 -1637 443 -1637 0 net=3105
rlabel metal2 478 -1637 478 -1637 0 net=3249
rlabel metal2 590 -1637 590 -1637 0 net=4297
rlabel metal2 702 -1637 702 -1637 0 net=5277
rlabel metal2 86 -1639 86 -1639 0 net=2040
rlabel metal2 152 -1639 152 -1639 0 net=2224
rlabel metal2 275 -1639 275 -1639 0 net=2075
rlabel metal2 296 -1639 296 -1639 0 net=4176
rlabel metal2 478 -1639 478 -1639 0 net=3285
rlabel metal2 590 -1639 590 -1639 0 net=4557
rlabel metal2 709 -1639 709 -1639 0 net=4909
rlabel metal2 86 -1641 86 -1641 0 net=1827
rlabel metal2 212 -1641 212 -1641 0 net=838
rlabel metal2 247 -1641 247 -1641 0 net=1489
rlabel metal2 296 -1641 296 -1641 0 net=1329
rlabel metal2 359 -1641 359 -1641 0 net=2491
rlabel metal2 390 -1641 390 -1641 0 net=3306
rlabel metal2 499 -1641 499 -1641 0 net=5867
rlabel metal2 597 -1641 597 -1641 0 net=5177
rlabel metal2 597 -1641 597 -1641 0 net=5177
rlabel metal2 604 -1641 604 -1641 0 net=4391
rlabel metal2 709 -1641 709 -1641 0 net=5029
rlabel metal2 758 -1641 758 -1641 0 net=5353
rlabel metal2 44 -1643 44 -1643 0 net=1144
rlabel metal2 212 -1643 212 -1643 0 net=3775
rlabel metal2 226 -1643 226 -1643 0 net=2731
rlabel metal2 289 -1643 289 -1643 0 net=2699
rlabel metal2 485 -1643 485 -1643 0 net=4679
rlabel metal2 583 -1643 583 -1643 0 net=4643
rlabel metal2 611 -1643 611 -1643 0 net=6255
rlabel metal2 716 -1643 716 -1643 0 net=4981
rlabel metal2 730 -1643 730 -1643 0 net=5011
rlabel metal2 23 -1645 23 -1645 0 net=4950
rlabel metal2 135 -1645 135 -1645 0 net=2097
rlabel metal2 317 -1645 317 -1645 0 net=2161
rlabel metal2 373 -1645 373 -1645 0 net=5787
rlabel metal2 485 -1645 485 -1645 0 net=3587
rlabel metal2 541 -1645 541 -1645 0 net=4063
rlabel metal2 614 -1645 614 -1645 0 net=5690
rlabel metal2 135 -1647 135 -1647 0 net=4633
rlabel metal2 156 -1647 156 -1647 0 net=6448
rlabel metal2 100 -1649 100 -1649 0 net=1641
rlabel metal2 170 -1649 170 -1649 0 net=1559
rlabel metal2 306 -1649 306 -1649 0 net=2797
rlabel metal2 394 -1649 394 -1649 0 net=5526
rlabel metal2 842 -1649 842 -1649 0 net=6367
rlabel metal2 51 -1651 51 -1651 0 net=2845
rlabel metal2 177 -1651 177 -1651 0 net=1619
rlabel metal2 317 -1651 317 -1651 0 net=1159
rlabel metal2 716 -1651 716 -1651 0 net=5701
rlabel metal2 40 -1653 40 -1653 0 net=1459
rlabel metal2 184 -1653 184 -1653 0 net=1937
rlabel metal2 324 -1653 324 -1653 0 net=4657
rlabel metal2 555 -1653 555 -1653 0 net=4799
rlabel metal2 733 -1653 733 -1653 0 net=3560
rlabel metal2 184 -1655 184 -1655 0 net=1267
rlabel metal2 331 -1655 331 -1655 0 net=2568
rlabel metal2 436 -1655 436 -1655 0 net=3001
rlabel metal2 506 -1655 506 -1655 0 net=4269
rlabel metal2 744 -1655 744 -1655 0 net=5679
rlabel metal2 884 -1655 884 -1655 0 net=4419
rlabel metal2 191 -1657 191 -1657 0 net=5141
rlabel metal2 338 -1657 338 -1657 0 net=2539
rlabel metal2 394 -1657 394 -1657 0 net=2917
rlabel metal2 786 -1657 786 -1657 0 net=5593
rlabel metal2 303 -1659 303 -1659 0 net=5771
rlabel metal2 772 -1659 772 -1659 0 net=5375
rlabel metal2 800 -1659 800 -1659 0 net=5412
rlabel metal2 313 -1661 313 -1661 0 net=5055
rlabel metal2 429 -1661 429 -1661 0 net=5605
rlabel metal2 800 -1661 800 -1661 0 net=3600
rlabel metal2 807 -1663 807 -1663 0 net=6177
rlabel metal2 863 -1665 863 -1665 0 net=6579
rlabel metal2 891 -1667 891 -1667 0 net=6587
rlabel metal2 905 -1669 905 -1669 0 net=6703
rlabel metal2 44 -1680 44 -1680 0 net=1461
rlabel metal2 65 -1680 65 -1680 0 net=6022
rlabel metal2 107 -1680 107 -1680 0 net=2327
rlabel metal2 264 -1680 264 -1680 0 net=4658
rlabel metal2 359 -1680 359 -1680 0 net=2541
rlabel metal2 359 -1680 359 -1680 0 net=2541
rlabel metal2 366 -1680 366 -1680 0 net=2393
rlabel metal2 366 -1680 366 -1680 0 net=2393
rlabel metal2 383 -1680 383 -1680 0 net=3862
rlabel metal2 408 -1680 408 -1680 0 net=5868
rlabel metal2 513 -1680 513 -1680 0 net=4991
rlabel metal2 541 -1680 541 -1680 0 net=6185
rlabel metal2 593 -1680 593 -1680 0 net=5178
rlabel metal2 611 -1680 611 -1680 0 net=6257
rlabel metal2 625 -1680 625 -1680 0 net=4299
rlabel metal2 646 -1680 646 -1680 0 net=4392
rlabel metal2 723 -1680 723 -1680 0 net=4983
rlabel metal2 758 -1680 758 -1680 0 net=5013
rlabel metal2 779 -1680 779 -1680 0 net=5625
rlabel metal2 856 -1680 856 -1680 0 net=6581
rlabel metal2 898 -1680 898 -1680 0 net=6705
rlabel metal2 968 -1680 968 -1680 0 net=5933
rlabel metal2 968 -1680 968 -1680 0 net=5933
rlabel metal2 1024 -1680 1024 -1680 0 net=6307
rlabel metal2 1024 -1680 1024 -1680 0 net=6307
rlabel metal2 47 -1682 47 -1682 0 net=2461
rlabel metal2 86 -1682 86 -1682 0 net=1828
rlabel metal2 310 -1682 310 -1682 0 net=5686
rlabel metal2 380 -1682 380 -1682 0 net=2493
rlabel metal2 422 -1682 422 -1682 0 net=6143
rlabel metal2 429 -1682 429 -1682 0 net=3107
rlabel metal2 450 -1682 450 -1682 0 net=5606
rlabel metal2 520 -1682 520 -1682 0 net=4558
rlabel metal2 604 -1682 604 -1682 0 net=4644
rlabel metal2 632 -1682 632 -1682 0 net=4109
rlabel metal2 653 -1682 653 -1682 0 net=977
rlabel metal2 709 -1682 709 -1682 0 net=5031
rlabel metal2 737 -1682 737 -1682 0 net=5427
rlabel metal2 782 -1682 782 -1682 0 net=6178
rlabel metal2 817 -1682 817 -1682 0 net=4420
rlabel metal2 93 -1684 93 -1684 0 net=2012
rlabel metal2 212 -1684 212 -1684 0 net=3776
rlabel metal2 373 -1684 373 -1684 0 net=2799
rlabel metal2 422 -1684 422 -1684 0 net=3003
rlabel metal2 450 -1684 450 -1684 0 net=3589
rlabel metal2 569 -1684 569 -1684 0 net=1421
rlabel metal2 709 -1684 709 -1684 0 net=5703
rlabel metal2 737 -1684 737 -1684 0 net=5681
rlabel metal2 786 -1684 786 -1684 0 net=5376
rlabel metal2 884 -1684 884 -1684 0 net=6589
rlabel metal2 75 -1686 75 -1686 0 net=6695
rlabel metal2 100 -1686 100 -1686 0 net=2846
rlabel metal2 201 -1686 201 -1686 0 net=2732
rlabel metal2 233 -1686 233 -1686 0 net=2099
rlabel metal2 233 -1686 233 -1686 0 net=2099
rlabel metal2 240 -1686 240 -1686 0 net=1704
rlabel metal2 282 -1686 282 -1686 0 net=2077
rlabel metal2 310 -1686 310 -1686 0 net=2163
rlabel metal2 373 -1686 373 -1686 0 net=5788
rlabel metal2 576 -1686 576 -1686 0 net=3250
rlabel metal2 667 -1686 667 -1686 0 net=4453
rlabel metal2 677 -1686 677 -1686 0 net=5692
rlabel metal2 744 -1686 744 -1686 0 net=4745
rlabel metal2 793 -1686 793 -1686 0 net=5225
rlabel metal2 807 -1686 807 -1686 0 net=6369
rlabel metal2 849 -1686 849 -1686 0 net=2257
rlabel metal2 114 -1688 114 -1688 0 net=5631
rlabel metal2 156 -1688 156 -1688 0 net=1642
rlabel metal2 219 -1688 219 -1688 0 net=1621
rlabel metal2 240 -1688 240 -1688 0 net=1939
rlabel metal2 324 -1688 324 -1688 0 net=1995
rlabel metal2 345 -1688 345 -1688 0 net=3457
rlabel metal2 401 -1688 401 -1688 0 net=4263
rlabel metal2 527 -1688 527 -1688 0 net=1953
rlabel metal2 702 -1688 702 -1688 0 net=5279
rlabel metal2 765 -1688 765 -1688 0 net=4911
rlabel metal2 821 -1688 821 -1688 0 net=5355
rlabel metal2 117 -1690 117 -1690 0 net=5452
rlabel metal2 128 -1690 128 -1690 0 net=6570
rlabel metal2 184 -1690 184 -1690 0 net=1269
rlabel metal2 247 -1690 247 -1690 0 net=1490
rlabel metal2 404 -1690 404 -1690 0 net=6671
rlabel metal2 464 -1690 464 -1690 0 net=4027
rlabel metal2 765 -1690 765 -1690 0 net=3887
rlabel metal2 821 -1690 821 -1690 0 net=2517
rlabel metal2 128 -1692 128 -1692 0 net=4635
rlabel metal2 142 -1692 142 -1692 0 net=967
rlabel metal2 142 -1692 142 -1692 0 net=967
rlabel metal2 156 -1692 156 -1692 0 net=1247
rlabel metal2 268 -1692 268 -1692 0 net=1555
rlabel metal2 415 -1692 415 -1692 0 net=5057
rlabel metal2 527 -1692 527 -1692 0 net=4801
rlabel metal2 828 -1692 828 -1692 0 net=5595
rlabel metal2 828 -1692 828 -1692 0 net=5595
rlabel metal2 163 -1694 163 -1694 0 net=2276
rlabel metal2 261 -1694 261 -1694 0 net=1519
rlabel metal2 275 -1694 275 -1694 0 net=2700
rlabel metal2 394 -1694 394 -1694 0 net=2919
rlabel metal2 436 -1694 436 -1694 0 net=3287
rlabel metal2 163 -1696 163 -1696 0 net=5143
rlabel metal2 289 -1696 289 -1696 0 net=1161
rlabel metal2 394 -1696 394 -1696 0 net=4815
rlabel metal2 457 -1696 457 -1696 0 net=5773
rlabel metal2 170 -1698 170 -1698 0 net=1561
rlabel metal2 170 -1698 170 -1698 0 net=1561
rlabel metal2 177 -1698 177 -1698 0 net=741
rlabel metal2 457 -1698 457 -1698 0 net=2469
rlabel metal2 191 -1700 191 -1700 0 net=1223
rlabel metal2 317 -1700 317 -1700 0 net=1943
rlabel metal2 471 -1700 471 -1700 0 net=6665
rlabel metal2 478 -1702 478 -1702 0 net=4271
rlabel metal2 548 -1702 548 -1702 0 net=6267
rlabel metal2 492 -1704 492 -1704 0 net=4681
rlabel metal2 562 -1704 562 -1704 0 net=4065
rlabel metal2 425 -1706 425 -1706 0 net=1
rlabel metal2 583 -1706 583 -1706 0 net=6373
rlabel metal2 44 -1717 44 -1717 0 net=1463
rlabel metal2 44 -1717 44 -1717 0 net=1463
rlabel metal2 58 -1717 58 -1717 0 net=2463
rlabel metal2 93 -1717 93 -1717 0 net=6696
rlabel metal2 121 -1717 121 -1717 0 net=4637
rlabel metal2 142 -1717 142 -1717 0 net=968
rlabel metal2 156 -1717 156 -1717 0 net=1248
rlabel metal2 191 -1717 191 -1717 0 net=1225
rlabel metal2 191 -1717 191 -1717 0 net=1225
rlabel metal2 212 -1717 212 -1717 0 net=1940
rlabel metal2 268 -1717 268 -1717 0 net=1521
rlabel metal2 289 -1717 289 -1717 0 net=1162
rlabel metal2 411 -1717 411 -1717 0 net=4264
rlabel metal2 541 -1717 541 -1717 0 net=6187
rlabel metal2 541 -1717 541 -1717 0 net=6187
rlabel metal2 562 -1717 562 -1717 0 net=4067
rlabel metal2 593 -1717 593 -1717 0 net=426
rlabel metal2 793 -1717 793 -1717 0 net=4913
rlabel metal2 800 -1717 800 -1717 0 net=5227
rlabel metal2 800 -1717 800 -1717 0 net=5227
rlabel metal2 828 -1717 828 -1717 0 net=5596
rlabel metal2 884 -1717 884 -1717 0 net=6591
rlabel metal2 884 -1717 884 -1717 0 net=6591
rlabel metal2 898 -1717 898 -1717 0 net=6707
rlabel metal2 898 -1717 898 -1717 0 net=6707
rlabel metal2 968 -1717 968 -1717 0 net=5935
rlabel metal2 968 -1717 968 -1717 0 net=5935
rlabel metal2 1024 -1717 1024 -1717 0 net=6309
rlabel metal2 1024 -1717 1024 -1717 0 net=6309
rlabel metal2 100 -1719 100 -1719 0 net=4069
rlabel metal2 100 -1719 100 -1719 0 net=4069
rlabel metal2 103 -1719 103 -1719 0 net=272
rlabel metal2 149 -1719 149 -1719 0 net=5633
rlabel metal2 205 -1719 205 -1719 0 net=4855
rlabel metal2 215 -1719 215 -1719 0 net=571
rlabel metal2 299 -1719 299 -1719 0 net=1422
rlabel metal2 583 -1719 583 -1719 0 net=6374
rlabel metal2 604 -1719 604 -1719 0 net=978
rlabel metal2 674 -1719 674 -1719 0 net=4454
rlabel metal2 702 -1719 702 -1719 0 net=5705
rlabel metal2 723 -1719 723 -1719 0 net=5033
rlabel metal2 723 -1719 723 -1719 0 net=5033
rlabel metal2 730 -1719 730 -1719 0 net=4985
rlabel metal2 772 -1719 772 -1719 0 net=5015
rlabel metal2 793 -1719 793 -1719 0 net=6371
rlabel metal2 821 -1719 821 -1719 0 net=2519
rlabel metal2 835 -1719 835 -1719 0 net=5357
rlabel metal2 845 -1719 845 -1719 0 net=6582
rlabel metal2 107 -1721 107 -1721 0 net=3821
rlabel metal2 142 -1721 142 -1721 0 net=44
rlabel metal2 163 -1721 163 -1721 0 net=5145
rlabel metal2 219 -1721 219 -1721 0 net=1270
rlabel metal2 303 -1721 303 -1721 0 net=2079
rlabel metal2 303 -1721 303 -1721 0 net=2079
rlabel metal2 310 -1721 310 -1721 0 net=2165
rlabel metal2 310 -1721 310 -1721 0 net=2165
rlabel metal2 324 -1721 324 -1721 0 net=1996
rlabel metal2 380 -1721 380 -1721 0 net=2801
rlabel metal2 422 -1721 422 -1721 0 net=3004
rlabel metal2 464 -1721 464 -1721 0 net=4028
rlabel metal2 597 -1721 597 -1721 0 net=6259
rlabel metal2 639 -1721 639 -1721 0 net=4300
rlabel metal2 709 -1721 709 -1721 0 net=5627
rlabel metal2 849 -1721 849 -1721 0 net=2259
rlabel metal2 163 -1723 163 -1723 0 net=1563
rlabel metal2 226 -1723 226 -1723 0 net=1623
rlabel metal2 296 -1723 296 -1723 0 net=4925
rlabel metal2 338 -1723 338 -1723 0 net=3458
rlabel metal2 352 -1723 352 -1723 0 net=465
rlabel metal2 646 -1723 646 -1723 0 net=4111
rlabel metal2 646 -1723 646 -1723 0 net=4111
rlabel metal2 730 -1723 730 -1723 0 net=5683
rlabel metal2 233 -1725 233 -1725 0 net=2101
rlabel metal2 282 -1725 282 -1725 0 net=1557
rlabel metal2 338 -1725 338 -1725 0 net=2627
rlabel metal2 422 -1725 422 -1725 0 net=3109
rlabel metal2 464 -1725 464 -1725 0 net=4273
rlabel metal2 492 -1725 492 -1725 0 net=6145
rlabel metal2 737 -1725 737 -1725 0 net=4747
rlabel metal2 226 -1727 226 -1727 0 net=3695
rlabel metal2 331 -1727 331 -1727 0 net=1333
rlabel metal2 429 -1727 429 -1727 0 net=2471
rlabel metal2 471 -1727 471 -1727 0 net=1954
rlabel metal2 744 -1727 744 -1727 0 net=3889
rlabel metal2 317 -1729 317 -1729 0 net=1945
rlabel metal2 345 -1729 345 -1729 0 net=2543
rlabel metal2 366 -1729 366 -1729 0 net=2395
rlabel metal2 457 -1729 457 -1729 0 net=6269
rlabel metal2 555 -1729 555 -1729 0 net=6667
rlabel metal2 758 -1729 758 -1729 0 net=5429
rlabel metal2 254 -1731 254 -1731 0 net=2329
rlabel metal2 352 -1731 352 -1731 0 net=2449
rlabel metal2 478 -1731 478 -1731 0 net=4683
rlabel metal2 534 -1731 534 -1731 0 net=5775
rlabel metal2 555 -1731 555 -1731 0 net=6691
rlabel metal2 751 -1731 751 -1731 0 net=5281
rlabel metal2 359 -1733 359 -1733 0 net=2921
rlabel metal2 485 -1733 485 -1733 0 net=5059
rlabel metal2 499 -1733 499 -1733 0 net=4803
rlabel metal2 366 -1735 366 -1735 0 net=4816
rlabel metal2 415 -1735 415 -1735 0 net=3591
rlabel metal2 513 -1735 513 -1735 0 net=4993
rlabel metal2 436 -1737 436 -1737 0 net=3289
rlabel metal2 485 -1737 485 -1737 0 net=4587
rlabel metal2 436 -1739 436 -1739 0 net=6673
rlabel metal2 796 -1739 796 -1739 0 net=1
rlabel metal2 44 -1750 44 -1750 0 net=1464
rlabel metal2 58 -1750 58 -1750 0 net=6233
rlabel metal2 65 -1750 65 -1750 0 net=2465
rlabel metal2 93 -1750 93 -1750 0 net=6215
rlabel metal2 121 -1750 121 -1750 0 net=4638
rlabel metal2 156 -1750 156 -1750 0 net=161
rlabel metal2 156 -1750 156 -1750 0 net=161
rlabel metal2 159 -1750 159 -1750 0 net=5634
rlabel metal2 184 -1750 184 -1750 0 net=5146
rlabel metal2 219 -1750 219 -1750 0 net=2102
rlabel metal2 275 -1750 275 -1750 0 net=1523
rlabel metal2 275 -1750 275 -1750 0 net=1523
rlabel metal2 282 -1750 282 -1750 0 net=2081
rlabel metal2 352 -1750 352 -1750 0 net=2450
rlabel metal2 373 -1750 373 -1750 0 net=1335
rlabel metal2 415 -1750 415 -1750 0 net=3593
rlabel metal2 415 -1750 415 -1750 0 net=3593
rlabel metal2 422 -1750 422 -1750 0 net=3110
rlabel metal2 422 -1750 422 -1750 0 net=3110
rlabel metal2 443 -1750 443 -1750 0 net=6271
rlabel metal2 464 -1750 464 -1750 0 net=4274
rlabel metal2 478 -1750 478 -1750 0 net=4685
rlabel metal2 478 -1750 478 -1750 0 net=4685
rlabel metal2 488 -1750 488 -1750 0 net=6668
rlabel metal2 586 -1750 586 -1750 0 net=4068
rlabel metal2 646 -1750 646 -1750 0 net=4112
rlabel metal2 716 -1750 716 -1750 0 net=5684
rlabel metal2 765 -1750 765 -1750 0 net=5430
rlabel metal2 807 -1750 807 -1750 0 net=4915
rlabel metal2 828 -1750 828 -1750 0 net=2521
rlabel metal2 828 -1750 828 -1750 0 net=2521
rlabel metal2 842 -1750 842 -1750 0 net=5358
rlabel metal2 856 -1750 856 -1750 0 net=2260
rlabel metal2 856 -1750 856 -1750 0 net=2260
rlabel metal2 884 -1750 884 -1750 0 net=6593
rlabel metal2 884 -1750 884 -1750 0 net=6593
rlabel metal2 898 -1750 898 -1750 0 net=6709
rlabel metal2 898 -1750 898 -1750 0 net=6709
rlabel metal2 968 -1750 968 -1750 0 net=5936
rlabel metal2 1024 -1750 1024 -1750 0 net=6311
rlabel metal2 1024 -1750 1024 -1750 0 net=6311
rlabel metal2 65 -1752 65 -1752 0 net=2795
rlabel metal2 100 -1752 100 -1752 0 net=4070
rlabel metal2 100 -1752 100 -1752 0 net=4070
rlabel metal2 107 -1752 107 -1752 0 net=3822
rlabel metal2 128 -1752 128 -1752 0 net=759
rlabel metal2 163 -1752 163 -1752 0 net=1564
rlabel metal2 191 -1752 191 -1752 0 net=1227
rlabel metal2 191 -1752 191 -1752 0 net=1227
rlabel metal2 205 -1752 205 -1752 0 net=4857
rlabel metal2 205 -1752 205 -1752 0 net=4857
rlabel metal2 219 -1752 219 -1752 0 net=3697
rlabel metal2 289 -1752 289 -1752 0 net=2167
rlabel metal2 317 -1752 317 -1752 0 net=2331
rlabel metal2 366 -1752 366 -1752 0 net=6453
rlabel metal2 380 -1752 380 -1752 0 net=2803
rlabel metal2 380 -1752 380 -1752 0 net=2803
rlabel metal2 387 -1752 387 -1752 0 net=2396
rlabel metal2 450 -1752 450 -1752 0 net=3291
rlabel metal2 471 -1752 471 -1752 0 net=5061
rlabel metal2 499 -1752 499 -1752 0 net=4804
rlabel metal2 513 -1752 513 -1752 0 net=4589
rlabel metal2 513 -1752 513 -1752 0 net=4589
rlabel metal2 527 -1752 527 -1752 0 net=6189
rlabel metal2 548 -1752 548 -1752 0 net=5776
rlabel metal2 562 -1752 562 -1752 0 net=6260
rlabel metal2 709 -1752 709 -1752 0 net=5629
rlabel metal2 772 -1752 772 -1752 0 net=5016
rlabel metal2 128 -1754 128 -1754 0 net=1163
rlabel metal2 135 -1754 135 -1754 0 net=2993
rlabel metal2 170 -1754 170 -1754 0 net=839
rlabel metal2 170 -1754 170 -1754 0 net=839
rlabel metal2 233 -1754 233 -1754 0 net=1625
rlabel metal2 296 -1754 296 -1754 0 net=1558
rlabel metal2 394 -1754 394 -1754 0 net=2497
rlabel metal2 394 -1754 394 -1754 0 net=2497
rlabel metal2 429 -1754 429 -1754 0 net=2473
rlabel metal2 457 -1754 457 -1754 0 net=6147
rlabel metal2 530 -1754 530 -1754 0 net=4994
rlabel metal2 562 -1754 562 -1754 0 net=6693
rlabel metal2 702 -1754 702 -1754 0 net=5707
rlabel metal2 723 -1754 723 -1754 0 net=5035
rlabel metal2 723 -1754 723 -1754 0 net=5035
rlabel metal2 758 -1754 758 -1754 0 net=5283
rlabel metal2 779 -1754 779 -1754 0 net=6372
rlabel metal2 138 -1756 138 -1756 0 net=3755
rlabel metal2 229 -1756 229 -1756 0 net=3605
rlabel metal2 296 -1756 296 -1756 0 net=1947
rlabel metal2 429 -1756 429 -1756 0 net=6674
rlabel metal2 506 -1756 506 -1756 0 net=6481
rlabel metal2 506 -1756 506 -1756 0 net=6481
rlabel metal2 751 -1756 751 -1756 0 net=4987
rlabel metal2 793 -1756 793 -1756 0 net=5229
rlabel metal2 310 -1758 310 -1758 0 net=2629
rlabel metal2 737 -1758 737 -1758 0 net=4749
rlabel metal2 324 -1760 324 -1760 0 net=4927
rlabel metal2 737 -1760 737 -1760 0 net=3891
rlabel metal2 324 -1762 324 -1762 0 net=2545
rlabel metal2 345 -1764 345 -1764 0 net=2923
rlabel metal2 359 -1766 359 -1766 0 net=200
rlabel metal2 58 -1777 58 -1777 0 net=6234
rlabel metal2 75 -1777 75 -1777 0 net=2796
rlabel metal2 93 -1777 93 -1777 0 net=6216
rlabel metal2 117 -1777 117 -1777 0 net=1164
rlabel metal2 135 -1777 135 -1777 0 net=2994
rlabel metal2 170 -1777 170 -1777 0 net=840
rlabel metal2 191 -1777 191 -1777 0 net=1228
rlabel metal2 205 -1777 205 -1777 0 net=4859
rlabel metal2 205 -1777 205 -1777 0 net=4859
rlabel metal2 219 -1777 219 -1777 0 net=3698
rlabel metal2 240 -1777 240 -1777 0 net=3607
rlabel metal2 240 -1777 240 -1777 0 net=3607
rlabel metal2 247 -1777 247 -1777 0 net=1187
rlabel metal2 282 -1777 282 -1777 0 net=2082
rlabel metal2 331 -1777 331 -1777 0 net=2924
rlabel metal2 352 -1777 352 -1777 0 net=2333
rlabel metal2 352 -1777 352 -1777 0 net=2333
rlabel metal2 380 -1777 380 -1777 0 net=2805
rlabel metal2 394 -1777 394 -1777 0 net=2498
rlabel metal2 415 -1777 415 -1777 0 net=3595
rlabel metal2 415 -1777 415 -1777 0 net=3595
rlabel metal2 443 -1777 443 -1777 0 net=6273
rlabel metal2 443 -1777 443 -1777 0 net=6273
rlabel metal2 478 -1777 478 -1777 0 net=4687
rlabel metal2 478 -1777 478 -1777 0 net=4687
rlabel metal2 502 -1777 502 -1777 0 net=6482
rlabel metal2 513 -1777 513 -1777 0 net=4591
rlabel metal2 513 -1777 513 -1777 0 net=4591
rlabel metal2 520 -1777 520 -1777 0 net=6191
rlabel metal2 562 -1777 562 -1777 0 net=6694
rlabel metal2 709 -1777 709 -1777 0 net=5708
rlabel metal2 723 -1777 723 -1777 0 net=5036
rlabel metal2 751 -1777 751 -1777 0 net=4751
rlabel metal2 772 -1777 772 -1777 0 net=5284
rlabel metal2 793 -1777 793 -1777 0 net=5231
rlabel metal2 793 -1777 793 -1777 0 net=5231
rlabel metal2 814 -1777 814 -1777 0 net=4916
rlabel metal2 814 -1777 814 -1777 0 net=4916
rlabel metal2 828 -1777 828 -1777 0 net=2522
rlabel metal2 880 -1777 880 -1777 0 net=6594
rlabel metal2 898 -1777 898 -1777 0 net=6711
rlabel metal2 898 -1777 898 -1777 0 net=6711
rlabel metal2 1024 -1777 1024 -1777 0 net=6313
rlabel metal2 1024 -1777 1024 -1777 0 net=6313
rlabel metal2 72 -1779 72 -1779 0 net=2467
rlabel metal2 142 -1779 142 -1779 0 net=3757
rlabel metal2 142 -1779 142 -1779 0 net=3757
rlabel metal2 152 -1779 152 -1779 0 net=5515
rlabel metal2 226 -1779 226 -1779 0 net=1627
rlabel metal2 275 -1779 275 -1779 0 net=1525
rlabel metal2 289 -1779 289 -1779 0 net=2168
rlabel metal2 324 -1779 324 -1779 0 net=2547
rlabel metal2 338 -1779 338 -1779 0 net=4929
rlabel metal2 338 -1779 338 -1779 0 net=4929
rlabel metal2 373 -1779 373 -1779 0 net=6455
rlabel metal2 401 -1779 401 -1779 0 net=1337
rlabel metal2 730 -1779 730 -1779 0 net=5630
rlabel metal2 296 -1781 296 -1781 0 net=1948
rlabel metal2 411 -1781 411 -1781 0 net=6148
rlabel metal2 737 -1781 737 -1781 0 net=3893
rlabel metal2 737 -1781 737 -1781 0 net=3893
rlabel metal2 758 -1781 758 -1781 0 net=4989
rlabel metal2 758 -1781 758 -1781 0 net=4989
rlabel metal2 296 -1783 296 -1783 0 net=1087
rlabel metal2 306 -1783 306 -1783 0 net=280
rlabel metal2 450 -1783 450 -1783 0 net=2475
rlabel metal2 310 -1785 310 -1785 0 net=2631
rlabel metal2 450 -1785 450 -1785 0 net=5063
rlabel metal2 464 -1787 464 -1787 0 net=3293
rlabel metal2 68 -1798 68 -1798 0 net=2468
rlabel metal2 142 -1798 142 -1798 0 net=3758
rlabel metal2 156 -1798 156 -1798 0 net=5516
rlabel metal2 184 -1798 184 -1798 0 net=1035
rlabel metal2 205 -1798 205 -1798 0 net=4860
rlabel metal2 226 -1798 226 -1798 0 net=1629
rlabel metal2 226 -1798 226 -1798 0 net=1629
rlabel metal2 240 -1798 240 -1798 0 net=3608
rlabel metal2 261 -1798 261 -1798 0 net=1189
rlabel metal2 282 -1798 282 -1798 0 net=1526
rlabel metal2 282 -1798 282 -1798 0 net=1526
rlabel metal2 296 -1798 296 -1798 0 net=1089
rlabel metal2 296 -1798 296 -1798 0 net=1089
rlabel metal2 324 -1798 324 -1798 0 net=2632
rlabel metal2 352 -1798 352 -1798 0 net=2335
rlabel metal2 352 -1798 352 -1798 0 net=2335
rlabel metal2 380 -1798 380 -1798 0 net=6456
rlabel metal2 387 -1798 387 -1798 0 net=2807
rlabel metal2 387 -1798 387 -1798 0 net=2807
rlabel metal2 422 -1798 422 -1798 0 net=1338
rlabel metal2 432 -1798 432 -1798 0 net=6274
rlabel metal2 457 -1798 457 -1798 0 net=2476
rlabel metal2 471 -1798 471 -1798 0 net=3294
rlabel metal2 506 -1798 506 -1798 0 net=4592
rlabel metal2 516 -1798 516 -1798 0 net=6192
rlabel metal2 737 -1798 737 -1798 0 net=3895
rlabel metal2 754 -1798 754 -1798 0 net=4752
rlabel metal2 793 -1798 793 -1798 0 net=5232
rlabel metal2 898 -1798 898 -1798 0 net=6713
rlabel metal2 1024 -1798 1024 -1798 0 net=6314
rlabel metal2 331 -1800 331 -1800 0 net=2548
rlabel metal2 415 -1800 415 -1800 0 net=3597
rlabel metal2 439 -1800 439 -1800 0 net=5064
rlabel metal2 471 -1800 471 -1800 0 net=4688
rlabel metal2 744 -1800 744 -1800 0 net=4990
rlabel metal2 331 -1802 331 -1802 0 net=4931
rlabel metal2 187 -1813 187 -1813 0 net=1036
rlabel metal2 222 -1813 222 -1813 0 net=1630
rlabel metal2 264 -1813 264 -1813 0 net=1190
rlabel metal2 296 -1813 296 -1813 0 net=1090
rlabel metal2 324 -1813 324 -1813 0 net=4932
rlabel metal2 352 -1813 352 -1813 0 net=2336
rlabel metal2 376 -1813 376 -1813 0 net=2808
rlabel metal2 422 -1813 422 -1813 0 net=3598
rlabel metal2 747 -1813 747 -1813 0 net=3896
rlabel metal2 901 -1813 901 -1813 0 net=6714
<< end >>
