magic
tech scmos
timestamp 1555071769 
<< pdiffusion >>
rect 1 -8 7 -2
rect 8 -8 14 -2
rect 15 -8 21 -2
rect 78 -8 84 -2
rect 85 -8 91 -2
rect 92 -8 98 -2
rect 99 -8 105 -2
rect 106 -8 109 -2
rect 148 -8 154 -2
rect 1 -25 7 -19
rect 8 -25 14 -19
rect 29 -25 35 -19
rect 50 -25 56 -19
rect 57 -25 60 -19
rect 64 -25 67 -19
rect 71 -25 77 -19
rect 78 -25 84 -19
rect 85 -25 88 -19
rect 92 -25 95 -19
rect 99 -25 105 -19
rect 106 -25 109 -19
rect 113 -25 116 -19
rect 120 -25 126 -19
rect 127 -25 130 -19
rect 134 -25 137 -19
rect 141 -25 144 -19
rect 148 -25 154 -19
rect 1 -46 7 -40
rect 22 -46 25 -40
rect 29 -46 32 -40
rect 36 -46 39 -40
rect 43 -46 49 -40
rect 50 -46 53 -40
rect 57 -46 63 -40
rect 64 -46 70 -40
rect 71 -46 74 -40
rect 78 -46 84 -40
rect 85 -46 91 -40
rect 92 -46 95 -40
rect 99 -46 105 -40
rect 106 -46 112 -40
rect 113 -46 119 -40
rect 120 -46 123 -40
rect 127 -46 130 -40
rect 134 -46 137 -40
rect 141 -46 144 -40
rect 148 -46 151 -40
rect 155 -46 161 -40
rect 162 -46 165 -40
rect 169 -46 172 -40
rect 176 -46 179 -40
rect 183 -46 186 -40
rect 190 -46 193 -40
rect 1 -75 7 -69
rect 15 -75 18 -69
rect 22 -75 25 -69
rect 29 -75 32 -69
rect 36 -75 42 -69
rect 43 -75 46 -69
rect 50 -75 53 -69
rect 57 -75 63 -69
rect 64 -75 70 -69
rect 71 -75 77 -69
rect 78 -75 84 -69
rect 85 -75 91 -69
rect 92 -75 98 -69
rect 99 -75 102 -69
rect 106 -75 109 -69
rect 113 -75 119 -69
rect 120 -75 123 -69
rect 127 -75 130 -69
rect 134 -75 137 -69
rect 141 -75 144 -69
rect 148 -75 151 -69
rect 155 -75 158 -69
rect 162 -75 165 -69
rect 169 -75 175 -69
rect 183 -75 186 -69
rect 190 -75 196 -69
rect 29 -102 32 -96
rect 36 -102 42 -96
rect 43 -102 49 -96
rect 50 -102 53 -96
rect 57 -102 63 -96
rect 64 -102 70 -96
rect 71 -102 74 -96
rect 78 -102 84 -96
rect 85 -102 91 -96
rect 92 -102 95 -96
rect 99 -102 105 -96
rect 106 -102 109 -96
rect 113 -102 116 -96
rect 120 -102 126 -96
rect 127 -102 130 -96
rect 134 -102 137 -96
rect 141 -102 144 -96
rect 148 -102 151 -96
rect 155 -102 161 -96
rect 183 -102 189 -96
rect 1 -129 4 -123
rect 8 -129 11 -123
rect 15 -129 18 -123
rect 22 -129 25 -123
rect 29 -129 35 -123
rect 36 -129 39 -123
rect 43 -129 49 -123
rect 50 -129 53 -123
rect 57 -129 60 -123
rect 64 -129 70 -123
rect 71 -129 74 -123
rect 78 -129 84 -123
rect 85 -129 91 -123
rect 92 -129 98 -123
rect 99 -129 102 -123
rect 106 -129 109 -123
rect 113 -129 119 -123
rect 120 -129 123 -123
rect 127 -129 133 -123
rect 134 -129 140 -123
rect 141 -129 147 -123
rect 148 -129 151 -123
rect 155 -129 158 -123
rect 162 -129 165 -123
rect 169 -129 172 -123
rect 176 -129 179 -123
rect 183 -129 186 -123
rect 15 -160 18 -154
rect 22 -160 25 -154
rect 29 -160 35 -154
rect 36 -160 39 -154
rect 43 -160 49 -154
rect 50 -160 56 -154
rect 57 -160 60 -154
rect 64 -160 67 -154
rect 71 -160 74 -154
rect 78 -160 84 -154
rect 85 -160 91 -154
rect 92 -160 98 -154
rect 99 -160 105 -154
rect 106 -160 109 -154
rect 113 -160 119 -154
rect 120 -160 123 -154
rect 127 -160 133 -154
rect 134 -160 140 -154
rect 141 -160 144 -154
rect 148 -160 151 -154
rect 155 -160 158 -154
rect 162 -160 165 -154
rect 169 -160 172 -154
rect 176 -160 179 -154
rect 183 -160 186 -154
rect 29 -193 35 -187
rect 36 -193 42 -187
rect 43 -193 49 -187
rect 50 -193 53 -187
rect 57 -193 63 -187
rect 64 -193 67 -187
rect 71 -193 77 -187
rect 78 -193 81 -187
rect 85 -193 91 -187
rect 92 -193 98 -187
rect 99 -193 102 -187
rect 106 -193 109 -187
rect 113 -193 116 -187
rect 120 -193 126 -187
rect 127 -193 130 -187
rect 134 -193 137 -187
rect 141 -193 147 -187
rect 148 -193 151 -187
rect 155 -193 158 -187
rect 162 -193 165 -187
rect 169 -193 172 -187
rect 176 -193 179 -187
rect 183 -193 186 -187
rect 50 -212 53 -206
rect 57 -212 60 -206
rect 64 -212 70 -206
rect 71 -212 74 -206
rect 78 -212 84 -206
rect 85 -212 88 -206
rect 92 -212 95 -206
rect 99 -212 102 -206
rect 106 -212 112 -206
rect 113 -212 119 -206
rect 120 -212 123 -206
rect 127 -212 130 -206
rect 134 -212 137 -206
rect 141 -212 147 -206
rect 148 -212 154 -206
rect 155 -212 161 -206
rect 57 -229 60 -223
rect 64 -229 70 -223
rect 71 -229 77 -223
rect 78 -229 84 -223
rect 85 -229 88 -223
rect 120 -229 126 -223
rect 134 -229 137 -223
rect 155 -229 161 -223
rect 155 -240 161 -234
rect 162 -240 165 -234
<< polysilicon >>
rect 79 -9 80 -7
rect 86 -3 87 -1
rect 86 -9 87 -7
rect 96 -9 97 -7
rect 100 -9 101 -7
rect 107 -3 108 -1
rect 107 -9 108 -7
rect 152 -9 153 -7
rect 33 -26 34 -24
rect 51 -20 52 -18
rect 58 -20 59 -18
rect 58 -26 59 -24
rect 65 -20 66 -18
rect 65 -26 66 -24
rect 72 -20 73 -18
rect 79 -20 80 -18
rect 82 -20 83 -18
rect 79 -26 80 -24
rect 86 -20 87 -18
rect 86 -26 87 -24
rect 93 -20 94 -18
rect 93 -26 94 -24
rect 100 -20 101 -18
rect 103 -20 104 -18
rect 100 -26 101 -24
rect 107 -20 108 -18
rect 107 -26 108 -24
rect 114 -20 115 -18
rect 114 -26 115 -24
rect 121 -20 122 -18
rect 128 -20 129 -18
rect 128 -26 129 -24
rect 135 -20 136 -18
rect 135 -26 136 -24
rect 142 -20 143 -18
rect 142 -26 143 -24
rect 149 -20 150 -18
rect 152 -20 153 -18
rect 149 -26 150 -24
rect 23 -41 24 -39
rect 23 -47 24 -45
rect 30 -41 31 -39
rect 30 -47 31 -45
rect 37 -41 38 -39
rect 37 -47 38 -45
rect 44 -47 45 -45
rect 51 -41 52 -39
rect 51 -47 52 -45
rect 58 -47 59 -45
rect 68 -41 69 -39
rect 65 -47 66 -45
rect 68 -47 69 -45
rect 72 -41 73 -39
rect 72 -47 73 -45
rect 79 -41 80 -39
rect 82 -47 83 -45
rect 86 -41 87 -39
rect 89 -41 90 -39
rect 86 -47 87 -45
rect 89 -47 90 -45
rect 93 -41 94 -39
rect 93 -47 94 -45
rect 100 -41 101 -39
rect 103 -41 104 -39
rect 100 -47 101 -45
rect 103 -47 104 -45
rect 107 -41 108 -39
rect 110 -41 111 -39
rect 107 -47 108 -45
rect 114 -47 115 -45
rect 117 -47 118 -45
rect 121 -41 122 -39
rect 121 -47 122 -45
rect 128 -41 129 -39
rect 128 -47 129 -45
rect 135 -41 136 -39
rect 135 -47 136 -45
rect 142 -41 143 -39
rect 142 -47 143 -45
rect 149 -41 150 -39
rect 149 -47 150 -45
rect 159 -41 160 -39
rect 163 -41 164 -39
rect 163 -47 164 -45
rect 170 -41 171 -39
rect 170 -47 171 -45
rect 177 -41 178 -39
rect 177 -47 178 -45
rect 184 -41 185 -39
rect 184 -47 185 -45
rect 191 -41 192 -39
rect 191 -47 192 -45
rect 16 -70 17 -68
rect 16 -76 17 -74
rect 23 -70 24 -68
rect 23 -76 24 -74
rect 30 -70 31 -68
rect 30 -76 31 -74
rect 37 -70 38 -68
rect 40 -70 41 -68
rect 40 -76 41 -74
rect 44 -70 45 -68
rect 44 -76 45 -74
rect 51 -70 52 -68
rect 51 -76 52 -74
rect 58 -70 59 -68
rect 61 -70 62 -68
rect 65 -70 66 -68
rect 68 -70 69 -68
rect 65 -76 66 -74
rect 72 -70 73 -68
rect 75 -70 76 -68
rect 72 -76 73 -74
rect 75 -76 76 -74
rect 82 -70 83 -68
rect 79 -76 80 -74
rect 86 -70 87 -68
rect 86 -76 87 -74
rect 93 -70 94 -68
rect 96 -70 97 -68
rect 96 -76 97 -74
rect 100 -70 101 -68
rect 100 -76 101 -74
rect 107 -70 108 -68
rect 107 -76 108 -74
rect 117 -70 118 -68
rect 114 -76 115 -74
rect 117 -76 118 -74
rect 121 -70 122 -68
rect 121 -76 122 -74
rect 128 -70 129 -68
rect 128 -76 129 -74
rect 135 -70 136 -68
rect 135 -76 136 -74
rect 142 -70 143 -68
rect 142 -76 143 -74
rect 149 -70 150 -68
rect 149 -76 150 -74
rect 156 -70 157 -68
rect 156 -76 157 -74
rect 163 -70 164 -68
rect 163 -76 164 -74
rect 173 -70 174 -68
rect 184 -70 185 -68
rect 184 -76 185 -74
rect 191 -70 192 -68
rect 30 -97 31 -95
rect 30 -103 31 -101
rect 37 -97 38 -95
rect 40 -97 41 -95
rect 40 -103 41 -101
rect 44 -97 45 -95
rect 47 -103 48 -101
rect 51 -97 52 -95
rect 51 -103 52 -101
rect 58 -97 59 -95
rect 58 -103 59 -101
rect 65 -97 66 -95
rect 65 -103 66 -101
rect 72 -97 73 -95
rect 72 -103 73 -101
rect 82 -97 83 -95
rect 79 -103 80 -101
rect 86 -97 87 -95
rect 89 -97 90 -95
rect 86 -103 87 -101
rect 89 -103 90 -101
rect 93 -97 94 -95
rect 93 -103 94 -101
rect 100 -97 101 -95
rect 103 -97 104 -95
rect 100 -103 101 -101
rect 107 -97 108 -95
rect 107 -103 108 -101
rect 114 -97 115 -95
rect 114 -103 115 -101
rect 121 -103 122 -101
rect 124 -103 125 -101
rect 128 -97 129 -95
rect 128 -103 129 -101
rect 135 -97 136 -95
rect 135 -103 136 -101
rect 142 -97 143 -95
rect 142 -103 143 -101
rect 149 -97 150 -95
rect 149 -103 150 -101
rect 156 -97 157 -95
rect 156 -103 157 -101
rect 184 -97 185 -95
rect 2 -124 3 -122
rect 2 -130 3 -128
rect 9 -124 10 -122
rect 9 -130 10 -128
rect 16 -124 17 -122
rect 16 -130 17 -128
rect 23 -124 24 -122
rect 23 -130 24 -128
rect 30 -124 31 -122
rect 33 -124 34 -122
rect 37 -124 38 -122
rect 37 -130 38 -128
rect 44 -124 45 -122
rect 47 -124 48 -122
rect 44 -130 45 -128
rect 47 -130 48 -128
rect 51 -124 52 -122
rect 51 -130 52 -128
rect 58 -124 59 -122
rect 58 -130 59 -128
rect 65 -124 66 -122
rect 68 -124 69 -122
rect 72 -124 73 -122
rect 72 -130 73 -128
rect 82 -124 83 -122
rect 82 -130 83 -128
rect 86 -124 87 -122
rect 89 -124 90 -122
rect 89 -130 90 -128
rect 93 -124 94 -122
rect 96 -124 97 -122
rect 93 -130 94 -128
rect 100 -124 101 -122
rect 100 -130 101 -128
rect 107 -124 108 -122
rect 107 -130 108 -128
rect 114 -124 115 -122
rect 117 -124 118 -122
rect 117 -130 118 -128
rect 121 -124 122 -122
rect 121 -130 122 -128
rect 131 -124 132 -122
rect 131 -130 132 -128
rect 135 -124 136 -122
rect 138 -124 139 -122
rect 145 -130 146 -128
rect 149 -124 150 -122
rect 149 -130 150 -128
rect 156 -124 157 -122
rect 156 -130 157 -128
rect 163 -124 164 -122
rect 163 -130 164 -128
rect 170 -124 171 -122
rect 170 -130 171 -128
rect 177 -124 178 -122
rect 177 -130 178 -128
rect 184 -124 185 -122
rect 184 -130 185 -128
rect 16 -155 17 -153
rect 16 -161 17 -159
rect 23 -155 24 -153
rect 23 -161 24 -159
rect 33 -155 34 -153
rect 33 -161 34 -159
rect 37 -155 38 -153
rect 37 -161 38 -159
rect 44 -155 45 -153
rect 47 -161 48 -159
rect 51 -155 52 -153
rect 54 -155 55 -153
rect 54 -161 55 -159
rect 58 -155 59 -153
rect 58 -161 59 -159
rect 65 -155 66 -153
rect 65 -161 66 -159
rect 72 -155 73 -153
rect 72 -161 73 -159
rect 79 -155 80 -153
rect 79 -161 80 -159
rect 86 -155 87 -153
rect 89 -155 90 -153
rect 86 -161 87 -159
rect 89 -161 90 -159
rect 93 -155 94 -153
rect 96 -155 97 -153
rect 93 -161 94 -159
rect 96 -161 97 -159
rect 100 -155 101 -153
rect 103 -155 104 -153
rect 100 -161 101 -159
rect 103 -161 104 -159
rect 107 -155 108 -153
rect 107 -161 108 -159
rect 114 -155 115 -153
rect 117 -155 118 -153
rect 114 -161 115 -159
rect 117 -161 118 -159
rect 121 -155 122 -153
rect 121 -161 122 -159
rect 131 -155 132 -153
rect 128 -161 129 -159
rect 135 -161 136 -159
rect 138 -161 139 -159
rect 142 -155 143 -153
rect 142 -161 143 -159
rect 149 -155 150 -153
rect 149 -161 150 -159
rect 156 -155 157 -153
rect 156 -161 157 -159
rect 163 -155 164 -153
rect 163 -161 164 -159
rect 170 -155 171 -153
rect 170 -161 171 -159
rect 177 -155 178 -153
rect 177 -161 178 -159
rect 184 -155 185 -153
rect 184 -161 185 -159
rect 33 -188 34 -186
rect 40 -188 41 -186
rect 44 -188 45 -186
rect 47 -194 48 -192
rect 51 -188 52 -186
rect 51 -194 52 -192
rect 61 -188 62 -186
rect 65 -188 66 -186
rect 65 -194 66 -192
rect 75 -188 76 -186
rect 72 -194 73 -192
rect 79 -188 80 -186
rect 79 -194 80 -192
rect 86 -194 87 -192
rect 89 -194 90 -192
rect 96 -188 97 -186
rect 93 -194 94 -192
rect 96 -194 97 -192
rect 100 -188 101 -186
rect 100 -194 101 -192
rect 107 -188 108 -186
rect 107 -194 108 -192
rect 114 -188 115 -186
rect 114 -194 115 -192
rect 121 -188 122 -186
rect 124 -188 125 -186
rect 121 -194 122 -192
rect 128 -188 129 -186
rect 128 -194 129 -192
rect 135 -188 136 -186
rect 135 -194 136 -192
rect 145 -194 146 -192
rect 149 -188 150 -186
rect 149 -194 150 -192
rect 156 -188 157 -186
rect 156 -194 157 -192
rect 163 -188 164 -186
rect 163 -194 164 -192
rect 170 -188 171 -186
rect 170 -194 171 -192
rect 177 -188 178 -186
rect 177 -194 178 -192
rect 184 -188 185 -186
rect 184 -194 185 -192
rect 51 -207 52 -205
rect 51 -213 52 -211
rect 58 -207 59 -205
rect 58 -213 59 -211
rect 68 -207 69 -205
rect 65 -213 66 -211
rect 68 -213 69 -211
rect 72 -207 73 -205
rect 72 -213 73 -211
rect 79 -207 80 -205
rect 79 -213 80 -211
rect 82 -213 83 -211
rect 86 -207 87 -205
rect 86 -213 87 -211
rect 93 -207 94 -205
rect 93 -213 94 -211
rect 100 -207 101 -205
rect 100 -213 101 -211
rect 110 -207 111 -205
rect 117 -207 118 -205
rect 114 -213 115 -211
rect 121 -207 122 -205
rect 121 -213 122 -211
rect 128 -207 129 -205
rect 128 -213 129 -211
rect 135 -207 136 -205
rect 135 -213 136 -211
rect 142 -207 143 -205
rect 142 -213 143 -211
rect 145 -213 146 -211
rect 152 -207 153 -205
rect 149 -213 150 -211
rect 152 -213 153 -211
rect 156 -207 157 -205
rect 58 -224 59 -222
rect 58 -230 59 -228
rect 68 -230 69 -228
rect 75 -224 76 -222
rect 79 -230 80 -228
rect 86 -224 87 -222
rect 86 -230 87 -228
rect 124 -224 125 -222
rect 124 -230 125 -228
rect 135 -224 136 -222
rect 135 -230 136 -228
rect 159 -224 160 -222
rect 156 -230 157 -228
rect 156 -241 157 -239
rect 163 -235 164 -233
rect 163 -241 164 -239
<< metal1 >>
rect 86 0 108 1
rect 51 -11 59 -10
rect 65 -11 73 -10
rect 82 -11 87 -10
rect 93 -11 97 -10
rect 100 -11 108 -10
rect 121 -11 129 -10
rect 149 -11 153 -10
rect 79 -13 87 -12
rect 100 -13 108 -12
rect 142 -13 153 -12
rect 79 -15 136 -14
rect 103 -17 115 -16
rect 30 -28 34 -27
rect 37 -28 66 -27
rect 68 -28 73 -27
rect 79 -28 104 -27
rect 107 -28 164 -27
rect 23 -30 108 -29
rect 110 -30 178 -29
rect 51 -32 59 -31
rect 79 -32 122 -31
rect 135 -32 171 -31
rect 86 -34 90 -33
rect 93 -34 101 -33
rect 128 -34 136 -33
rect 149 -34 185 -33
rect 86 -36 94 -35
rect 100 -36 129 -35
rect 142 -36 150 -35
rect 159 -36 192 -35
rect 114 -38 143 -37
rect 16 -49 31 -48
rect 37 -49 83 -48
rect 86 -49 164 -48
rect 173 -49 185 -48
rect 23 -51 66 -50
rect 72 -51 87 -50
rect 100 -51 143 -50
rect 163 -51 171 -50
rect 23 -53 76 -52
rect 96 -53 143 -52
rect 40 -55 69 -54
rect 103 -55 150 -54
rect 44 -57 90 -56
rect 107 -57 178 -56
rect 37 -59 45 -58
rect 51 -59 83 -58
rect 93 -59 108 -58
rect 114 -59 192 -58
rect 51 -61 62 -60
rect 72 -61 94 -60
rect 117 -61 150 -60
rect 184 -61 192 -60
rect 58 -63 66 -62
rect 100 -63 118 -62
rect 135 -63 157 -62
rect 30 -65 59 -64
rect 121 -65 136 -64
rect 68 -67 122 -66
rect 16 -78 41 -77
rect 51 -78 73 -77
rect 75 -78 108 -77
rect 114 -78 164 -77
rect 23 -80 59 -79
rect 82 -80 122 -79
rect 30 -82 66 -81
rect 86 -82 94 -81
rect 96 -82 136 -81
rect 30 -84 38 -83
rect 40 -84 45 -83
rect 65 -84 73 -83
rect 86 -84 108 -83
rect 117 -84 157 -83
rect 44 -86 52 -85
rect 89 -86 115 -85
rect 142 -86 157 -85
rect 79 -88 143 -87
rect 100 -90 136 -89
rect 103 -92 150 -91
rect 100 -94 150 -93
rect 2 -105 34 -104
rect 37 -105 52 -104
rect 58 -105 83 -104
rect 86 -105 136 -104
rect 142 -105 164 -104
rect 9 -107 101 -106
rect 121 -107 129 -106
rect 131 -107 178 -106
rect 16 -109 31 -108
rect 40 -109 48 -108
rect 51 -109 157 -108
rect 23 -111 31 -110
rect 44 -111 118 -110
rect 124 -111 139 -110
rect 149 -111 171 -110
rect 47 -113 69 -112
rect 72 -113 80 -112
rect 89 -113 108 -112
rect 114 -113 150 -112
rect 58 -115 97 -114
rect 107 -115 115 -114
rect 135 -115 185 -114
rect 65 -117 87 -116
rect 89 -117 122 -116
rect 65 -119 73 -118
rect 93 -119 157 -118
rect 93 -121 101 -120
rect 2 -132 48 -131
rect 58 -132 80 -131
rect 82 -132 115 -131
rect 117 -132 150 -131
rect 16 -134 45 -133
rect 65 -134 104 -133
rect 131 -134 150 -133
rect 16 -136 34 -135
rect 37 -136 45 -135
rect 72 -136 90 -135
rect 93 -136 164 -135
rect 9 -138 90 -137
rect 93 -138 143 -137
rect 145 -138 171 -137
rect 51 -140 73 -139
rect 86 -140 101 -139
rect 163 -140 178 -139
rect 37 -142 101 -141
rect 121 -142 178 -141
rect 51 -144 59 -143
rect 96 -144 157 -143
rect 170 -144 185 -143
rect 54 -146 157 -145
rect 107 -148 122 -147
rect 107 -150 132 -149
rect 117 -152 185 -151
rect 16 -163 45 -162
rect 51 -163 104 -162
rect 114 -163 157 -162
rect 23 -165 34 -164
rect 37 -165 55 -164
rect 58 -165 118 -164
rect 121 -165 157 -164
rect 33 -167 48 -166
rect 61 -167 108 -166
rect 114 -167 143 -166
rect 40 -169 87 -168
rect 100 -169 171 -168
rect 65 -171 101 -170
rect 121 -171 171 -170
rect 65 -173 76 -172
rect 128 -173 164 -172
rect 72 -175 94 -174
rect 96 -175 164 -174
rect 96 -177 108 -176
rect 128 -177 139 -176
rect 135 -179 178 -178
rect 135 -181 150 -180
rect 177 -181 185 -180
rect 89 -183 150 -182
rect 124 -185 185 -184
rect 51 -196 73 -195
rect 79 -196 94 -195
rect 96 -196 115 -195
rect 121 -196 136 -195
rect 142 -196 164 -195
rect 47 -198 52 -197
rect 58 -198 80 -197
rect 86 -198 157 -197
rect 65 -200 73 -199
rect 89 -200 101 -199
rect 110 -200 136 -199
rect 145 -200 171 -199
rect 68 -202 87 -201
rect 93 -202 118 -201
rect 121 -202 129 -201
rect 152 -202 178 -201
rect 100 -204 108 -203
rect 128 -204 150 -203
rect 156 -204 185 -203
rect 51 -215 69 -214
rect 72 -215 76 -214
rect 79 -215 101 -214
rect 114 -215 136 -214
rect 149 -215 160 -214
rect 65 -217 83 -216
rect 93 -217 125 -216
rect 128 -217 146 -216
rect 121 -219 143 -218
rect 135 -221 153 -220
rect 58 -232 69 -231
rect 79 -232 87 -231
rect 124 -232 136 -231
rect 156 -232 164 -231
rect 156 -243 164 -242
<< m2contact >>
rect 86 0 87 1
rect 107 0 108 1
rect 51 -11 52 -10
rect 58 -11 59 -10
rect 65 -11 66 -10
rect 72 -11 73 -10
rect 82 -11 83 -10
rect 86 -11 87 -10
rect 93 -11 94 -10
rect 96 -11 97 -10
rect 100 -11 101 -10
rect 107 -11 108 -10
rect 121 -11 122 -10
rect 128 -11 129 -10
rect 149 -11 150 -10
rect 152 -11 153 -10
rect 79 -13 80 -12
rect 86 -13 87 -12
rect 100 -13 101 -12
rect 107 -13 108 -12
rect 142 -13 143 -12
rect 152 -13 153 -12
rect 79 -15 80 -14
rect 135 -15 136 -14
rect 103 -17 104 -16
rect 114 -17 115 -16
rect 30 -28 31 -27
rect 33 -28 34 -27
rect 37 -28 38 -27
rect 65 -28 66 -27
rect 68 -28 69 -27
rect 72 -28 73 -27
rect 79 -28 80 -27
rect 103 -28 104 -27
rect 107 -28 108 -27
rect 163 -28 164 -27
rect 23 -30 24 -29
rect 107 -30 108 -29
rect 110 -30 111 -29
rect 177 -30 178 -29
rect 51 -32 52 -31
rect 58 -32 59 -31
rect 79 -32 80 -31
rect 121 -32 122 -31
rect 135 -32 136 -31
rect 170 -32 171 -31
rect 86 -34 87 -33
rect 89 -34 90 -33
rect 93 -34 94 -33
rect 100 -34 101 -33
rect 128 -34 129 -33
rect 135 -34 136 -33
rect 149 -34 150 -33
rect 184 -34 185 -33
rect 86 -36 87 -35
rect 93 -36 94 -35
rect 100 -36 101 -35
rect 128 -36 129 -35
rect 142 -36 143 -35
rect 149 -36 150 -35
rect 159 -36 160 -35
rect 191 -36 192 -35
rect 114 -38 115 -37
rect 142 -38 143 -37
rect 16 -49 17 -48
rect 30 -49 31 -48
rect 37 -49 38 -48
rect 82 -49 83 -48
rect 86 -49 87 -48
rect 163 -49 164 -48
rect 173 -49 174 -48
rect 184 -49 185 -48
rect 23 -51 24 -50
rect 65 -51 66 -50
rect 72 -51 73 -50
rect 86 -51 87 -50
rect 100 -51 101 -50
rect 142 -51 143 -50
rect 163 -51 164 -50
rect 170 -51 171 -50
rect 23 -53 24 -52
rect 75 -53 76 -52
rect 96 -53 97 -52
rect 142 -53 143 -52
rect 40 -55 41 -54
rect 68 -55 69 -54
rect 103 -55 104 -54
rect 149 -55 150 -54
rect 44 -57 45 -56
rect 89 -57 90 -56
rect 107 -57 108 -56
rect 177 -57 178 -56
rect 37 -59 38 -58
rect 44 -59 45 -58
rect 51 -59 52 -58
rect 82 -59 83 -58
rect 93 -59 94 -58
rect 107 -59 108 -58
rect 114 -59 115 -58
rect 191 -59 192 -58
rect 51 -61 52 -60
rect 61 -61 62 -60
rect 72 -61 73 -60
rect 93 -61 94 -60
rect 117 -61 118 -60
rect 149 -61 150 -60
rect 184 -61 185 -60
rect 191 -61 192 -60
rect 58 -63 59 -62
rect 65 -63 66 -62
rect 100 -63 101 -62
rect 117 -63 118 -62
rect 135 -63 136 -62
rect 156 -63 157 -62
rect 30 -65 31 -64
rect 58 -65 59 -64
rect 121 -65 122 -64
rect 135 -65 136 -64
rect 68 -67 69 -66
rect 121 -67 122 -66
rect 16 -78 17 -77
rect 40 -78 41 -77
rect 51 -78 52 -77
rect 72 -78 73 -77
rect 75 -78 76 -77
rect 107 -78 108 -77
rect 114 -78 115 -77
rect 163 -78 164 -77
rect 23 -80 24 -79
rect 58 -80 59 -79
rect 82 -80 83 -79
rect 121 -80 122 -79
rect 30 -82 31 -81
rect 65 -82 66 -81
rect 86 -82 87 -81
rect 93 -82 94 -81
rect 96 -82 97 -81
rect 135 -82 136 -81
rect 30 -84 31 -83
rect 37 -84 38 -83
rect 40 -84 41 -83
rect 44 -84 45 -83
rect 65 -84 66 -83
rect 72 -84 73 -83
rect 86 -84 87 -83
rect 107 -84 108 -83
rect 117 -84 118 -83
rect 156 -84 157 -83
rect 44 -86 45 -85
rect 51 -86 52 -85
rect 89 -86 90 -85
rect 114 -86 115 -85
rect 142 -86 143 -85
rect 156 -86 157 -85
rect 79 -88 80 -87
rect 142 -88 143 -87
rect 100 -90 101 -89
rect 135 -90 136 -89
rect 103 -92 104 -91
rect 149 -92 150 -91
rect 100 -94 101 -93
rect 149 -94 150 -93
rect 2 -105 3 -104
rect 33 -105 34 -104
rect 37 -105 38 -104
rect 51 -105 52 -104
rect 58 -105 59 -104
rect 82 -105 83 -104
rect 86 -105 87 -104
rect 135 -105 136 -104
rect 142 -105 143 -104
rect 163 -105 164 -104
rect 9 -107 10 -106
rect 100 -107 101 -106
rect 121 -107 122 -106
rect 128 -107 129 -106
rect 131 -107 132 -106
rect 177 -107 178 -106
rect 16 -109 17 -108
rect 30 -109 31 -108
rect 40 -109 41 -108
rect 47 -109 48 -108
rect 51 -109 52 -108
rect 156 -109 157 -108
rect 23 -111 24 -110
rect 30 -111 31 -110
rect 44 -111 45 -110
rect 117 -111 118 -110
rect 124 -111 125 -110
rect 138 -111 139 -110
rect 149 -111 150 -110
rect 170 -111 171 -110
rect 47 -113 48 -112
rect 68 -113 69 -112
rect 72 -113 73 -112
rect 79 -113 80 -112
rect 89 -113 90 -112
rect 107 -113 108 -112
rect 114 -113 115 -112
rect 149 -113 150 -112
rect 58 -115 59 -114
rect 96 -115 97 -114
rect 107 -115 108 -114
rect 114 -115 115 -114
rect 135 -115 136 -114
rect 184 -115 185 -114
rect 65 -117 66 -116
rect 86 -117 87 -116
rect 89 -117 90 -116
rect 121 -117 122 -116
rect 65 -119 66 -118
rect 72 -119 73 -118
rect 93 -119 94 -118
rect 156 -119 157 -118
rect 93 -121 94 -120
rect 100 -121 101 -120
rect 2 -132 3 -131
rect 47 -132 48 -131
rect 58 -132 59 -131
rect 79 -132 80 -131
rect 82 -132 83 -131
rect 114 -132 115 -131
rect 117 -132 118 -131
rect 149 -132 150 -131
rect 16 -134 17 -133
rect 44 -134 45 -133
rect 65 -134 66 -133
rect 103 -134 104 -133
rect 131 -134 132 -133
rect 149 -134 150 -133
rect 16 -136 17 -135
rect 33 -136 34 -135
rect 37 -136 38 -135
rect 44 -136 45 -135
rect 72 -136 73 -135
rect 89 -136 90 -135
rect 93 -136 94 -135
rect 163 -136 164 -135
rect 9 -138 10 -137
rect 89 -138 90 -137
rect 93 -138 94 -137
rect 142 -138 143 -137
rect 145 -138 146 -137
rect 170 -138 171 -137
rect 51 -140 52 -139
rect 72 -140 73 -139
rect 86 -140 87 -139
rect 100 -140 101 -139
rect 163 -140 164 -139
rect 177 -140 178 -139
rect 37 -142 38 -141
rect 100 -142 101 -141
rect 121 -142 122 -141
rect 177 -142 178 -141
rect 51 -144 52 -143
rect 58 -144 59 -143
rect 96 -144 97 -143
rect 156 -144 157 -143
rect 170 -144 171 -143
rect 184 -144 185 -143
rect 54 -146 55 -145
rect 156 -146 157 -145
rect 107 -148 108 -147
rect 121 -148 122 -147
rect 107 -150 108 -149
rect 131 -150 132 -149
rect 117 -152 118 -151
rect 184 -152 185 -151
rect 16 -163 17 -162
rect 44 -163 45 -162
rect 51 -163 52 -162
rect 103 -163 104 -162
rect 114 -163 115 -162
rect 156 -163 157 -162
rect 23 -165 24 -164
rect 33 -165 34 -164
rect 37 -165 38 -164
rect 54 -165 55 -164
rect 58 -165 59 -164
rect 117 -165 118 -164
rect 121 -165 122 -164
rect 156 -165 157 -164
rect 33 -167 34 -166
rect 47 -167 48 -166
rect 61 -167 62 -166
rect 107 -167 108 -166
rect 114 -167 115 -166
rect 142 -167 143 -166
rect 40 -169 41 -168
rect 86 -169 87 -168
rect 100 -169 101 -168
rect 170 -169 171 -168
rect 65 -171 66 -170
rect 100 -171 101 -170
rect 121 -171 122 -170
rect 170 -171 171 -170
rect 65 -173 66 -172
rect 75 -173 76 -172
rect 128 -173 129 -172
rect 163 -173 164 -172
rect 72 -175 73 -174
rect 93 -175 94 -174
rect 96 -175 97 -174
rect 163 -175 164 -174
rect 96 -177 97 -176
rect 107 -177 108 -176
rect 128 -177 129 -176
rect 138 -177 139 -176
rect 135 -179 136 -178
rect 177 -179 178 -178
rect 135 -181 136 -180
rect 149 -181 150 -180
rect 177 -181 178 -180
rect 184 -181 185 -180
rect 89 -183 90 -182
rect 149 -183 150 -182
rect 124 -185 125 -184
rect 184 -185 185 -184
rect 51 -196 52 -195
rect 72 -196 73 -195
rect 79 -196 80 -195
rect 93 -196 94 -195
rect 96 -196 97 -195
rect 114 -196 115 -195
rect 121 -196 122 -195
rect 135 -196 136 -195
rect 142 -196 143 -195
rect 163 -196 164 -195
rect 47 -198 48 -197
rect 51 -198 52 -197
rect 58 -198 59 -197
rect 79 -198 80 -197
rect 86 -198 87 -197
rect 156 -198 157 -197
rect 65 -200 66 -199
rect 72 -200 73 -199
rect 89 -200 90 -199
rect 100 -200 101 -199
rect 110 -200 111 -199
rect 135 -200 136 -199
rect 145 -200 146 -199
rect 170 -200 171 -199
rect 68 -202 69 -201
rect 86 -202 87 -201
rect 93 -202 94 -201
rect 117 -202 118 -201
rect 121 -202 122 -201
rect 128 -202 129 -201
rect 152 -202 153 -201
rect 177 -202 178 -201
rect 100 -204 101 -203
rect 107 -204 108 -203
rect 128 -204 129 -203
rect 149 -204 150 -203
rect 156 -204 157 -203
rect 184 -204 185 -203
rect 51 -215 52 -214
rect 68 -215 69 -214
rect 72 -215 73 -214
rect 75 -215 76 -214
rect 79 -215 80 -214
rect 100 -215 101 -214
rect 114 -215 115 -214
rect 135 -215 136 -214
rect 149 -215 150 -214
rect 159 -215 160 -214
rect 65 -217 66 -216
rect 82 -217 83 -216
rect 93 -217 94 -216
rect 124 -217 125 -216
rect 128 -217 129 -216
rect 145 -217 146 -216
rect 121 -219 122 -218
rect 142 -219 143 -218
rect 135 -221 136 -220
rect 152 -221 153 -220
rect 58 -232 59 -231
rect 68 -232 69 -231
rect 79 -232 80 -231
rect 86 -232 87 -231
rect 124 -232 125 -231
rect 135 -232 136 -231
rect 156 -232 157 -231
rect 163 -232 164 -231
rect 156 -243 157 -242
rect 163 -243 164 -242
<< metal2 >>
rect 86 -1 87 1
rect 107 -1 108 1
rect 51 -18 52 -10
rect 58 -18 59 -10
rect 65 -18 66 -10
rect 72 -18 73 -10
rect 82 -18 83 -10
rect 86 -11 87 -9
rect 93 -18 94 -10
rect 96 -11 97 -9
rect 100 -11 101 -9
rect 107 -11 108 -9
rect 121 -18 122 -10
rect 128 -18 129 -10
rect 149 -18 150 -10
rect 152 -11 153 -9
rect 79 -13 80 -9
rect 86 -18 87 -12
rect 100 -18 101 -12
rect 107 -18 108 -12
rect 142 -18 143 -12
rect 152 -18 153 -12
rect 79 -18 80 -14
rect 135 -18 136 -14
rect 103 -18 104 -16
rect 114 -18 115 -16
rect 30 -39 31 -27
rect 33 -28 34 -26
rect 37 -39 38 -27
rect 65 -28 66 -26
rect 68 -39 69 -27
rect 72 -39 73 -27
rect 79 -28 80 -26
rect 103 -39 104 -27
rect 107 -28 108 -26
rect 163 -39 164 -27
rect 23 -39 24 -29
rect 107 -39 108 -29
rect 110 -39 111 -29
rect 177 -39 178 -29
rect 51 -39 52 -31
rect 58 -32 59 -26
rect 79 -39 80 -31
rect 121 -39 122 -31
rect 135 -32 136 -26
rect 170 -39 171 -31
rect 86 -34 87 -26
rect 89 -39 90 -33
rect 93 -34 94 -26
rect 100 -34 101 -26
rect 128 -34 129 -26
rect 135 -39 136 -33
rect 149 -34 150 -26
rect 184 -39 185 -33
rect 86 -39 87 -35
rect 93 -39 94 -35
rect 100 -39 101 -35
rect 128 -39 129 -35
rect 142 -36 143 -26
rect 149 -39 150 -35
rect 159 -39 160 -35
rect 191 -39 192 -35
rect 114 -38 115 -26
rect 142 -39 143 -37
rect 16 -68 17 -48
rect 30 -49 31 -47
rect 37 -49 38 -47
rect 82 -49 83 -47
rect 86 -49 87 -47
rect 163 -49 164 -47
rect 173 -68 174 -48
rect 184 -49 185 -47
rect 23 -51 24 -47
rect 65 -51 66 -47
rect 72 -51 73 -47
rect 86 -68 87 -50
rect 100 -51 101 -47
rect 142 -51 143 -47
rect 163 -68 164 -50
rect 170 -51 171 -47
rect 23 -68 24 -52
rect 75 -68 76 -52
rect 96 -68 97 -52
rect 142 -68 143 -52
rect 40 -68 41 -54
rect 68 -55 69 -47
rect 103 -55 104 -47
rect 149 -55 150 -47
rect 44 -57 45 -47
rect 89 -57 90 -47
rect 107 -57 108 -47
rect 177 -57 178 -47
rect 37 -68 38 -58
rect 44 -68 45 -58
rect 51 -59 52 -47
rect 82 -68 83 -58
rect 93 -59 94 -47
rect 107 -68 108 -58
rect 114 -59 115 -47
rect 191 -59 192 -47
rect 51 -68 52 -60
rect 61 -68 62 -60
rect 72 -68 73 -60
rect 93 -68 94 -60
rect 117 -61 118 -47
rect 149 -68 150 -60
rect 184 -68 185 -60
rect 191 -68 192 -60
rect 58 -63 59 -47
rect 65 -68 66 -62
rect 100 -68 101 -62
rect 117 -68 118 -62
rect 128 -63 129 -47
rect 128 -68 129 -62
rect 128 -63 129 -47
rect 128 -68 129 -62
rect 135 -63 136 -47
rect 156 -68 157 -62
rect 30 -68 31 -64
rect 58 -68 59 -64
rect 121 -65 122 -47
rect 135 -68 136 -64
rect 68 -68 69 -66
rect 121 -68 122 -66
rect 16 -78 17 -76
rect 40 -78 41 -76
rect 51 -78 52 -76
rect 72 -78 73 -76
rect 75 -78 76 -76
rect 107 -78 108 -76
rect 114 -78 115 -76
rect 163 -78 164 -76
rect 184 -78 185 -76
rect 184 -95 185 -77
rect 184 -78 185 -76
rect 184 -95 185 -77
rect 23 -80 24 -76
rect 58 -95 59 -79
rect 82 -95 83 -79
rect 121 -80 122 -76
rect 128 -80 129 -76
rect 128 -95 129 -79
rect 128 -80 129 -76
rect 128 -95 129 -79
rect 30 -82 31 -76
rect 65 -82 66 -76
rect 86 -82 87 -76
rect 93 -95 94 -81
rect 96 -82 97 -76
rect 135 -82 136 -76
rect 30 -95 31 -83
rect 37 -95 38 -83
rect 40 -95 41 -83
rect 44 -84 45 -76
rect 65 -95 66 -83
rect 72 -95 73 -83
rect 86 -95 87 -83
rect 107 -95 108 -83
rect 117 -84 118 -76
rect 156 -84 157 -76
rect 44 -95 45 -85
rect 51 -95 52 -85
rect 89 -95 90 -85
rect 114 -95 115 -85
rect 142 -86 143 -76
rect 156 -95 157 -85
rect 79 -88 80 -76
rect 142 -95 143 -87
rect 100 -90 101 -76
rect 135 -95 136 -89
rect 103 -95 104 -91
rect 149 -92 150 -76
rect 100 -95 101 -93
rect 149 -95 150 -93
rect 2 -122 3 -104
rect 33 -122 34 -104
rect 37 -122 38 -104
rect 51 -105 52 -103
rect 58 -105 59 -103
rect 82 -122 83 -104
rect 86 -105 87 -103
rect 135 -105 136 -103
rect 142 -105 143 -103
rect 163 -122 164 -104
rect 9 -122 10 -106
rect 100 -107 101 -103
rect 121 -107 122 -103
rect 128 -107 129 -103
rect 131 -122 132 -106
rect 177 -122 178 -106
rect 16 -122 17 -108
rect 30 -109 31 -103
rect 40 -109 41 -103
rect 47 -109 48 -103
rect 51 -122 52 -108
rect 156 -109 157 -103
rect 23 -122 24 -110
rect 30 -122 31 -110
rect 44 -122 45 -110
rect 117 -122 118 -110
rect 124 -111 125 -103
rect 138 -122 139 -110
rect 149 -111 150 -103
rect 170 -122 171 -110
rect 47 -122 48 -112
rect 68 -122 69 -112
rect 72 -113 73 -103
rect 79 -113 80 -103
rect 89 -113 90 -103
rect 107 -113 108 -103
rect 114 -113 115 -103
rect 149 -122 150 -112
rect 58 -122 59 -114
rect 96 -122 97 -114
rect 107 -122 108 -114
rect 114 -122 115 -114
rect 135 -122 136 -114
rect 184 -122 185 -114
rect 65 -117 66 -103
rect 86 -122 87 -116
rect 89 -122 90 -116
rect 121 -122 122 -116
rect 65 -122 66 -118
rect 72 -122 73 -118
rect 93 -119 94 -103
rect 156 -122 157 -118
rect 93 -122 94 -120
rect 100 -122 101 -120
rect 2 -132 3 -130
rect 47 -132 48 -130
rect 58 -132 59 -130
rect 79 -153 80 -131
rect 82 -132 83 -130
rect 114 -153 115 -131
rect 117 -132 118 -130
rect 149 -132 150 -130
rect 16 -134 17 -130
rect 44 -134 45 -130
rect 65 -153 66 -133
rect 103 -153 104 -133
rect 131 -134 132 -130
rect 149 -153 150 -133
rect 16 -153 17 -135
rect 33 -153 34 -135
rect 37 -136 38 -130
rect 44 -153 45 -135
rect 72 -136 73 -130
rect 89 -136 90 -130
rect 93 -136 94 -130
rect 163 -136 164 -130
rect 9 -138 10 -130
rect 89 -153 90 -137
rect 93 -153 94 -137
rect 142 -153 143 -137
rect 145 -138 146 -130
rect 170 -138 171 -130
rect 23 -140 24 -130
rect 23 -153 24 -139
rect 23 -140 24 -130
rect 23 -153 24 -139
rect 51 -140 52 -130
rect 72 -153 73 -139
rect 86 -153 87 -139
rect 100 -140 101 -130
rect 163 -153 164 -139
rect 177 -140 178 -130
rect 37 -153 38 -141
rect 100 -153 101 -141
rect 121 -142 122 -130
rect 177 -153 178 -141
rect 51 -153 52 -143
rect 58 -153 59 -143
rect 96 -153 97 -143
rect 156 -144 157 -130
rect 170 -153 171 -143
rect 184 -144 185 -130
rect 54 -153 55 -145
rect 156 -153 157 -145
rect 107 -148 108 -130
rect 121 -153 122 -147
rect 107 -153 108 -149
rect 131 -153 132 -149
rect 117 -153 118 -151
rect 184 -153 185 -151
rect 16 -163 17 -161
rect 44 -186 45 -162
rect 51 -186 52 -162
rect 103 -163 104 -161
rect 114 -163 115 -161
rect 156 -163 157 -161
rect 23 -165 24 -161
rect 33 -165 34 -161
rect 37 -165 38 -161
rect 54 -165 55 -161
rect 58 -165 59 -161
rect 117 -165 118 -161
rect 121 -165 122 -161
rect 156 -186 157 -164
rect 33 -186 34 -166
rect 47 -167 48 -161
rect 61 -186 62 -166
rect 107 -167 108 -161
rect 114 -186 115 -166
rect 142 -167 143 -161
rect 40 -186 41 -168
rect 86 -169 87 -161
rect 100 -169 101 -161
rect 170 -169 171 -161
rect 65 -171 66 -161
rect 100 -186 101 -170
rect 121 -186 122 -170
rect 170 -186 171 -170
rect 65 -186 66 -172
rect 75 -186 76 -172
rect 79 -173 80 -161
rect 79 -186 80 -172
rect 79 -173 80 -161
rect 79 -186 80 -172
rect 128 -173 129 -161
rect 163 -173 164 -161
rect 72 -175 73 -161
rect 93 -175 94 -161
rect 96 -175 97 -161
rect 163 -186 164 -174
rect 96 -186 97 -176
rect 107 -186 108 -176
rect 128 -186 129 -176
rect 138 -177 139 -161
rect 135 -179 136 -161
rect 177 -179 178 -161
rect 135 -186 136 -180
rect 149 -181 150 -161
rect 177 -186 178 -180
rect 184 -181 185 -161
rect 89 -183 90 -161
rect 149 -186 150 -182
rect 124 -186 125 -184
rect 184 -186 185 -184
rect 51 -196 52 -194
rect 72 -196 73 -194
rect 79 -196 80 -194
rect 93 -196 94 -194
rect 96 -196 97 -194
rect 114 -196 115 -194
rect 121 -196 122 -194
rect 135 -196 136 -194
rect 142 -205 143 -195
rect 163 -196 164 -194
rect 47 -198 48 -194
rect 51 -205 52 -197
rect 58 -205 59 -197
rect 79 -205 80 -197
rect 86 -198 87 -194
rect 156 -198 157 -194
rect 65 -200 66 -194
rect 72 -205 73 -199
rect 89 -200 90 -194
rect 100 -200 101 -194
rect 110 -205 111 -199
rect 135 -205 136 -199
rect 145 -200 146 -194
rect 170 -200 171 -194
rect 68 -205 69 -201
rect 86 -205 87 -201
rect 93 -205 94 -201
rect 117 -205 118 -201
rect 121 -205 122 -201
rect 128 -202 129 -194
rect 152 -205 153 -201
rect 177 -202 178 -194
rect 100 -205 101 -203
rect 107 -204 108 -194
rect 128 -205 129 -203
rect 149 -204 150 -194
rect 156 -205 157 -203
rect 184 -204 185 -194
rect 51 -215 52 -213
rect 68 -215 69 -213
rect 72 -215 73 -213
rect 75 -222 76 -214
rect 79 -215 80 -213
rect 100 -215 101 -213
rect 114 -215 115 -213
rect 135 -215 136 -213
rect 149 -215 150 -213
rect 159 -222 160 -214
rect 58 -217 59 -213
rect 58 -222 59 -216
rect 58 -217 59 -213
rect 58 -222 59 -216
rect 65 -217 66 -213
rect 82 -217 83 -213
rect 86 -217 87 -213
rect 86 -222 87 -216
rect 86 -217 87 -213
rect 86 -222 87 -216
rect 93 -217 94 -213
rect 124 -222 125 -216
rect 128 -217 129 -213
rect 145 -217 146 -213
rect 121 -219 122 -213
rect 142 -219 143 -213
rect 135 -222 136 -220
rect 152 -221 153 -213
rect 58 -232 59 -230
rect 68 -232 69 -230
rect 79 -232 80 -230
rect 86 -232 87 -230
rect 124 -232 125 -230
rect 135 -232 136 -230
rect 156 -232 157 -230
rect 163 -233 164 -231
rect 156 -243 157 -241
rect 163 -243 164 -241
<< labels >>
rlabel pdiffusion 3 -6 3 -6 0 cellNo=1
rlabel pdiffusion 10 -6 10 -6 0 cellNo=18
rlabel pdiffusion 17 -6 17 -6 0 cellNo=55
rlabel pdiffusion 80 -6 80 -6 0 cellNo=13
rlabel pdiffusion 87 -6 87 -6 0 cellNo=24
rlabel pdiffusion 94 -6 94 -6 0 cellNo=56
rlabel pdiffusion 101 -6 101 -6 0 cellNo=6
rlabel pdiffusion 108 -6 108 -6 0 feedthrough
rlabel pdiffusion 150 -6 150 -6 0 cellNo=9
rlabel pdiffusion 3 -23 3 -23 0 cellNo=19
rlabel pdiffusion 10 -23 10 -23 0 cellNo=57
rlabel pdiffusion 31 -23 31 -23 0 cellNo=3
rlabel pdiffusion 52 -23 52 -23 0 cellNo=47
rlabel pdiffusion 59 -23 59 -23 0 feedthrough
rlabel pdiffusion 66 -23 66 -23 0 feedthrough
rlabel pdiffusion 73 -23 73 -23 0 cellNo=35
rlabel pdiffusion 80 -23 80 -23 0 cellNo=11
rlabel pdiffusion 87 -23 87 -23 0 feedthrough
rlabel pdiffusion 94 -23 94 -23 0 feedthrough
rlabel pdiffusion 101 -23 101 -23 0 cellNo=36
rlabel pdiffusion 108 -23 108 -23 0 feedthrough
rlabel pdiffusion 115 -23 115 -23 0 feedthrough
rlabel pdiffusion 122 -23 122 -23 0 cellNo=70
rlabel pdiffusion 129 -23 129 -23 0 feedthrough
rlabel pdiffusion 136 -23 136 -23 0 feedthrough
rlabel pdiffusion 143 -23 143 -23 0 feedthrough
rlabel pdiffusion 150 -23 150 -23 0 cellNo=43
rlabel pdiffusion 3 -44 3 -44 0 cellNo=32
rlabel pdiffusion 24 -44 24 -44 0 feedthrough
rlabel pdiffusion 31 -44 31 -44 0 feedthrough
rlabel pdiffusion 38 -44 38 -44 0 feedthrough
rlabel pdiffusion 45 -44 45 -44 0 cellNo=72
rlabel pdiffusion 52 -44 52 -44 0 feedthrough
rlabel pdiffusion 59 -44 59 -44 0 cellNo=64
rlabel pdiffusion 66 -44 66 -44 0 cellNo=31
rlabel pdiffusion 73 -44 73 -44 0 feedthrough
rlabel pdiffusion 80 -44 80 -44 0 cellNo=58
rlabel pdiffusion 87 -44 87 -44 0 cellNo=44
rlabel pdiffusion 94 -44 94 -44 0 feedthrough
rlabel pdiffusion 101 -44 101 -44 0 cellNo=68
rlabel pdiffusion 108 -44 108 -44 0 cellNo=22
rlabel pdiffusion 115 -44 115 -44 0 cellNo=30
rlabel pdiffusion 122 -44 122 -44 0 feedthrough
rlabel pdiffusion 129 -44 129 -44 0 feedthrough
rlabel pdiffusion 136 -44 136 -44 0 feedthrough
rlabel pdiffusion 143 -44 143 -44 0 feedthrough
rlabel pdiffusion 150 -44 150 -44 0 feedthrough
rlabel pdiffusion 157 -44 157 -44 0 cellNo=12
rlabel pdiffusion 164 -44 164 -44 0 feedthrough
rlabel pdiffusion 171 -44 171 -44 0 feedthrough
rlabel pdiffusion 178 -44 178 -44 0 feedthrough
rlabel pdiffusion 185 -44 185 -44 0 feedthrough
rlabel pdiffusion 192 -44 192 -44 0 feedthrough
rlabel pdiffusion 3 -73 3 -73 0 cellNo=67
rlabel pdiffusion 17 -73 17 -73 0 feedthrough
rlabel pdiffusion 24 -73 24 -73 0 feedthrough
rlabel pdiffusion 31 -73 31 -73 0 feedthrough
rlabel pdiffusion 38 -73 38 -73 0 cellNo=28
rlabel pdiffusion 45 -73 45 -73 0 feedthrough
rlabel pdiffusion 52 -73 52 -73 0 feedthrough
rlabel pdiffusion 59 -73 59 -73 0 cellNo=26
rlabel pdiffusion 66 -73 66 -73 0 cellNo=65
rlabel pdiffusion 73 -73 73 -73 0 cellNo=84
rlabel pdiffusion 80 -73 80 -73 0 cellNo=14
rlabel pdiffusion 87 -73 87 -73 0 cellNo=85
rlabel pdiffusion 94 -73 94 -73 0 cellNo=7
rlabel pdiffusion 101 -73 101 -73 0 feedthrough
rlabel pdiffusion 108 -73 108 -73 0 feedthrough
rlabel pdiffusion 115 -73 115 -73 0 cellNo=37
rlabel pdiffusion 122 -73 122 -73 0 feedthrough
rlabel pdiffusion 129 -73 129 -73 0 feedthrough
rlabel pdiffusion 136 -73 136 -73 0 feedthrough
rlabel pdiffusion 143 -73 143 -73 0 feedthrough
rlabel pdiffusion 150 -73 150 -73 0 feedthrough
rlabel pdiffusion 157 -73 157 -73 0 feedthrough
rlabel pdiffusion 164 -73 164 -73 0 feedthrough
rlabel pdiffusion 171 -73 171 -73 0 cellNo=21
rlabel pdiffusion 185 -73 185 -73 0 feedthrough
rlabel pdiffusion 192 -73 192 -73 0 cellNo=15
rlabel pdiffusion 31 -100 31 -100 0 feedthrough
rlabel pdiffusion 38 -100 38 -100 0 cellNo=59
rlabel pdiffusion 45 -100 45 -100 0 cellNo=60
rlabel pdiffusion 52 -100 52 -100 0 feedthrough
rlabel pdiffusion 59 -100 59 -100 0 cellNo=40
rlabel pdiffusion 66 -100 66 -100 0 cellNo=78
rlabel pdiffusion 73 -100 73 -100 0 feedthrough
rlabel pdiffusion 80 -100 80 -100 0 cellNo=82
rlabel pdiffusion 87 -100 87 -100 0 cellNo=48
rlabel pdiffusion 94 -100 94 -100 0 feedthrough
rlabel pdiffusion 101 -100 101 -100 0 cellNo=80
rlabel pdiffusion 108 -100 108 -100 0 feedthrough
rlabel pdiffusion 115 -100 115 -100 0 feedthrough
rlabel pdiffusion 122 -100 122 -100 0 cellNo=2
rlabel pdiffusion 129 -100 129 -100 0 feedthrough
rlabel pdiffusion 136 -100 136 -100 0 feedthrough
rlabel pdiffusion 143 -100 143 -100 0 feedthrough
rlabel pdiffusion 150 -100 150 -100 0 feedthrough
rlabel pdiffusion 157 -100 157 -100 0 cellNo=4
rlabel pdiffusion 185 -100 185 -100 0 cellNo=10
rlabel pdiffusion 3 -127 3 -127 0 feedthrough
rlabel pdiffusion 10 -127 10 -127 0 feedthrough
rlabel pdiffusion 17 -127 17 -127 0 feedthrough
rlabel pdiffusion 24 -127 24 -127 0 feedthrough
rlabel pdiffusion 31 -127 31 -127 0 cellNo=29
rlabel pdiffusion 38 -127 38 -127 0 feedthrough
rlabel pdiffusion 45 -127 45 -127 0 cellNo=87
rlabel pdiffusion 52 -127 52 -127 0 feedthrough
rlabel pdiffusion 59 -127 59 -127 0 feedthrough
rlabel pdiffusion 66 -127 66 -127 0 cellNo=42
rlabel pdiffusion 73 -127 73 -127 0 feedthrough
rlabel pdiffusion 80 -127 80 -127 0 cellNo=86
rlabel pdiffusion 87 -127 87 -127 0 cellNo=90
rlabel pdiffusion 94 -127 94 -127 0 cellNo=46
rlabel pdiffusion 101 -127 101 -127 0 feedthrough
rlabel pdiffusion 108 -127 108 -127 0 feedthrough
rlabel pdiffusion 115 -127 115 -127 0 cellNo=69
rlabel pdiffusion 122 -127 122 -127 0 feedthrough
rlabel pdiffusion 129 -127 129 -127 0 cellNo=61
rlabel pdiffusion 136 -127 136 -127 0 cellNo=52
rlabel pdiffusion 143 -127 143 -127 0 cellNo=41
rlabel pdiffusion 150 -127 150 -127 0 feedthrough
rlabel pdiffusion 157 -127 157 -127 0 feedthrough
rlabel pdiffusion 164 -127 164 -127 0 feedthrough
rlabel pdiffusion 171 -127 171 -127 0 feedthrough
rlabel pdiffusion 178 -127 178 -127 0 feedthrough
rlabel pdiffusion 185 -127 185 -127 0 feedthrough
rlabel pdiffusion 17 -158 17 -158 0 feedthrough
rlabel pdiffusion 24 -158 24 -158 0 feedthrough
rlabel pdiffusion 31 -158 31 -158 0 cellNo=25
rlabel pdiffusion 38 -158 38 -158 0 feedthrough
rlabel pdiffusion 45 -158 45 -158 0 cellNo=27
rlabel pdiffusion 52 -158 52 -158 0 cellNo=89
rlabel pdiffusion 59 -158 59 -158 0 feedthrough
rlabel pdiffusion 66 -158 66 -158 0 feedthrough
rlabel pdiffusion 73 -158 73 -158 0 feedthrough
rlabel pdiffusion 80 -158 80 -158 0 cellNo=33
rlabel pdiffusion 87 -158 87 -158 0 cellNo=38
rlabel pdiffusion 94 -158 94 -158 0 cellNo=53
rlabel pdiffusion 101 -158 101 -158 0 cellNo=76
rlabel pdiffusion 108 -158 108 -158 0 feedthrough
rlabel pdiffusion 115 -158 115 -158 0 cellNo=5
rlabel pdiffusion 122 -158 122 -158 0 feedthrough
rlabel pdiffusion 129 -158 129 -158 0 cellNo=49
rlabel pdiffusion 136 -158 136 -158 0 cellNo=39
rlabel pdiffusion 143 -158 143 -158 0 feedthrough
rlabel pdiffusion 150 -158 150 -158 0 feedthrough
rlabel pdiffusion 157 -158 157 -158 0 feedthrough
rlabel pdiffusion 164 -158 164 -158 0 feedthrough
rlabel pdiffusion 171 -158 171 -158 0 feedthrough
rlabel pdiffusion 178 -158 178 -158 0 feedthrough
rlabel pdiffusion 185 -158 185 -158 0 feedthrough
rlabel pdiffusion 31 -191 31 -191 0 cellNo=50
rlabel pdiffusion 38 -191 38 -191 0 cellNo=74
rlabel pdiffusion 45 -191 45 -191 0 cellNo=79
rlabel pdiffusion 52 -191 52 -191 0 feedthrough
rlabel pdiffusion 59 -191 59 -191 0 cellNo=63
rlabel pdiffusion 66 -191 66 -191 0 feedthrough
rlabel pdiffusion 73 -191 73 -191 0 cellNo=8
rlabel pdiffusion 80 -191 80 -191 0 feedthrough
rlabel pdiffusion 87 -191 87 -191 0 cellNo=83
rlabel pdiffusion 94 -191 94 -191 0 cellNo=34
rlabel pdiffusion 101 -191 101 -191 0 feedthrough
rlabel pdiffusion 108 -191 108 -191 0 feedthrough
rlabel pdiffusion 115 -191 115 -191 0 feedthrough
rlabel pdiffusion 122 -191 122 -191 0 cellNo=17
rlabel pdiffusion 129 -191 129 -191 0 feedthrough
rlabel pdiffusion 136 -191 136 -191 0 feedthrough
rlabel pdiffusion 143 -191 143 -191 0 cellNo=51
rlabel pdiffusion 150 -191 150 -191 0 feedthrough
rlabel pdiffusion 157 -191 157 -191 0 feedthrough
rlabel pdiffusion 164 -191 164 -191 0 feedthrough
rlabel pdiffusion 171 -191 171 -191 0 feedthrough
rlabel pdiffusion 178 -191 178 -191 0 feedthrough
rlabel pdiffusion 185 -191 185 -191 0 feedthrough
rlabel pdiffusion 52 -210 52 -210 0 feedthrough
rlabel pdiffusion 59 -210 59 -210 0 feedthrough
rlabel pdiffusion 66 -210 66 -210 0 cellNo=16
rlabel pdiffusion 73 -210 73 -210 0 feedthrough
rlabel pdiffusion 80 -210 80 -210 0 cellNo=77
rlabel pdiffusion 87 -210 87 -210 0 feedthrough
rlabel pdiffusion 94 -210 94 -210 0 feedthrough
rlabel pdiffusion 101 -210 101 -210 0 feedthrough
rlabel pdiffusion 108 -210 108 -210 0 cellNo=88
rlabel pdiffusion 115 -210 115 -210 0 cellNo=45
rlabel pdiffusion 122 -210 122 -210 0 feedthrough
rlabel pdiffusion 129 -210 129 -210 0 feedthrough
rlabel pdiffusion 136 -210 136 -210 0 feedthrough
rlabel pdiffusion 143 -210 143 -210 0 cellNo=54
rlabel pdiffusion 150 -210 150 -210 0 cellNo=62
rlabel pdiffusion 157 -210 157 -210 0 cellNo=20
rlabel pdiffusion 59 -227 59 -227 0 feedthrough
rlabel pdiffusion 66 -227 66 -227 0 cellNo=81
rlabel pdiffusion 73 -227 73 -227 0 cellNo=66
rlabel pdiffusion 80 -227 80 -227 0 cellNo=23
rlabel pdiffusion 87 -227 87 -227 0 feedthrough
rlabel pdiffusion 122 -227 122 -227 0 cellNo=73
rlabel pdiffusion 136 -227 136 -227 0 feedthrough
rlabel pdiffusion 157 -227 157 -227 0 cellNo=75
rlabel pdiffusion 157 -238 157 -238 0 cellNo=71
rlabel pdiffusion 164 -238 164 -238 0 feedthrough
rlabel polysilicon 79 -8 79 -8 0 3
rlabel polysilicon 86 -2 86 -2 0 1
rlabel polysilicon 86 -8 86 -8 0 3
rlabel polysilicon 96 -8 96 -8 0 4
rlabel polysilicon 100 -8 100 -8 0 3
rlabel polysilicon 107 -2 107 -2 0 1
rlabel polysilicon 107 -8 107 -8 0 3
rlabel polysilicon 152 -8 152 -8 0 4
rlabel polysilicon 33 -25 33 -25 0 4
rlabel polysilicon 51 -19 51 -19 0 1
rlabel polysilicon 58 -19 58 -19 0 1
rlabel polysilicon 58 -25 58 -25 0 3
rlabel polysilicon 65 -19 65 -19 0 1
rlabel polysilicon 65 -25 65 -25 0 3
rlabel polysilicon 72 -19 72 -19 0 1
rlabel polysilicon 79 -19 79 -19 0 1
rlabel polysilicon 82 -19 82 -19 0 2
rlabel polysilicon 79 -25 79 -25 0 3
rlabel polysilicon 86 -19 86 -19 0 1
rlabel polysilicon 86 -25 86 -25 0 3
rlabel polysilicon 93 -19 93 -19 0 1
rlabel polysilicon 93 -25 93 -25 0 3
rlabel polysilicon 100 -19 100 -19 0 1
rlabel polysilicon 103 -19 103 -19 0 2
rlabel polysilicon 100 -25 100 -25 0 3
rlabel polysilicon 107 -19 107 -19 0 1
rlabel polysilicon 107 -25 107 -25 0 3
rlabel polysilicon 114 -19 114 -19 0 1
rlabel polysilicon 114 -25 114 -25 0 3
rlabel polysilicon 121 -19 121 -19 0 1
rlabel polysilicon 128 -19 128 -19 0 1
rlabel polysilicon 128 -25 128 -25 0 3
rlabel polysilicon 135 -19 135 -19 0 1
rlabel polysilicon 135 -25 135 -25 0 3
rlabel polysilicon 142 -19 142 -19 0 1
rlabel polysilicon 142 -25 142 -25 0 3
rlabel polysilicon 149 -19 149 -19 0 1
rlabel polysilicon 152 -19 152 -19 0 2
rlabel polysilicon 149 -25 149 -25 0 3
rlabel polysilicon 23 -40 23 -40 0 1
rlabel polysilicon 23 -46 23 -46 0 3
rlabel polysilicon 30 -40 30 -40 0 1
rlabel polysilicon 30 -46 30 -46 0 3
rlabel polysilicon 37 -40 37 -40 0 1
rlabel polysilicon 37 -46 37 -46 0 3
rlabel polysilicon 44 -46 44 -46 0 3
rlabel polysilicon 51 -40 51 -40 0 1
rlabel polysilicon 51 -46 51 -46 0 3
rlabel polysilicon 58 -46 58 -46 0 3
rlabel polysilicon 68 -40 68 -40 0 2
rlabel polysilicon 65 -46 65 -46 0 3
rlabel polysilicon 68 -46 68 -46 0 4
rlabel polysilicon 72 -40 72 -40 0 1
rlabel polysilicon 72 -46 72 -46 0 3
rlabel polysilicon 79 -40 79 -40 0 1
rlabel polysilicon 82 -46 82 -46 0 4
rlabel polysilicon 86 -40 86 -40 0 1
rlabel polysilicon 89 -40 89 -40 0 2
rlabel polysilicon 86 -46 86 -46 0 3
rlabel polysilicon 89 -46 89 -46 0 4
rlabel polysilicon 93 -40 93 -40 0 1
rlabel polysilicon 93 -46 93 -46 0 3
rlabel polysilicon 100 -40 100 -40 0 1
rlabel polysilicon 103 -40 103 -40 0 2
rlabel polysilicon 100 -46 100 -46 0 3
rlabel polysilicon 103 -46 103 -46 0 4
rlabel polysilicon 107 -40 107 -40 0 1
rlabel polysilicon 110 -40 110 -40 0 2
rlabel polysilicon 107 -46 107 -46 0 3
rlabel polysilicon 114 -46 114 -46 0 3
rlabel polysilicon 117 -46 117 -46 0 4
rlabel polysilicon 121 -40 121 -40 0 1
rlabel polysilicon 121 -46 121 -46 0 3
rlabel polysilicon 128 -40 128 -40 0 1
rlabel polysilicon 128 -46 128 -46 0 3
rlabel polysilicon 135 -40 135 -40 0 1
rlabel polysilicon 135 -46 135 -46 0 3
rlabel polysilicon 142 -40 142 -40 0 1
rlabel polysilicon 142 -46 142 -46 0 3
rlabel polysilicon 149 -40 149 -40 0 1
rlabel polysilicon 149 -46 149 -46 0 3
rlabel polysilicon 159 -40 159 -40 0 2
rlabel polysilicon 163 -40 163 -40 0 1
rlabel polysilicon 163 -46 163 -46 0 3
rlabel polysilicon 170 -40 170 -40 0 1
rlabel polysilicon 170 -46 170 -46 0 3
rlabel polysilicon 177 -40 177 -40 0 1
rlabel polysilicon 177 -46 177 -46 0 3
rlabel polysilicon 184 -40 184 -40 0 1
rlabel polysilicon 184 -46 184 -46 0 3
rlabel polysilicon 191 -40 191 -40 0 1
rlabel polysilicon 191 -46 191 -46 0 3
rlabel polysilicon 16 -69 16 -69 0 1
rlabel polysilicon 16 -75 16 -75 0 3
rlabel polysilicon 23 -69 23 -69 0 1
rlabel polysilicon 23 -75 23 -75 0 3
rlabel polysilicon 30 -69 30 -69 0 1
rlabel polysilicon 30 -75 30 -75 0 3
rlabel polysilicon 37 -69 37 -69 0 1
rlabel polysilicon 40 -69 40 -69 0 2
rlabel polysilicon 40 -75 40 -75 0 4
rlabel polysilicon 44 -69 44 -69 0 1
rlabel polysilicon 44 -75 44 -75 0 3
rlabel polysilicon 51 -69 51 -69 0 1
rlabel polysilicon 51 -75 51 -75 0 3
rlabel polysilicon 58 -69 58 -69 0 1
rlabel polysilicon 61 -69 61 -69 0 2
rlabel polysilicon 65 -69 65 -69 0 1
rlabel polysilicon 68 -69 68 -69 0 2
rlabel polysilicon 65 -75 65 -75 0 3
rlabel polysilicon 72 -69 72 -69 0 1
rlabel polysilicon 75 -69 75 -69 0 2
rlabel polysilicon 72 -75 72 -75 0 3
rlabel polysilicon 75 -75 75 -75 0 4
rlabel polysilicon 82 -69 82 -69 0 2
rlabel polysilicon 79 -75 79 -75 0 3
rlabel polysilicon 86 -69 86 -69 0 1
rlabel polysilicon 86 -75 86 -75 0 3
rlabel polysilicon 93 -69 93 -69 0 1
rlabel polysilicon 96 -69 96 -69 0 2
rlabel polysilicon 96 -75 96 -75 0 4
rlabel polysilicon 100 -69 100 -69 0 1
rlabel polysilicon 100 -75 100 -75 0 3
rlabel polysilicon 107 -69 107 -69 0 1
rlabel polysilicon 107 -75 107 -75 0 3
rlabel polysilicon 117 -69 117 -69 0 2
rlabel polysilicon 114 -75 114 -75 0 3
rlabel polysilicon 117 -75 117 -75 0 4
rlabel polysilicon 121 -69 121 -69 0 1
rlabel polysilicon 121 -75 121 -75 0 3
rlabel polysilicon 128 -69 128 -69 0 1
rlabel polysilicon 128 -75 128 -75 0 3
rlabel polysilicon 135 -69 135 -69 0 1
rlabel polysilicon 135 -75 135 -75 0 3
rlabel polysilicon 142 -69 142 -69 0 1
rlabel polysilicon 142 -75 142 -75 0 3
rlabel polysilicon 149 -69 149 -69 0 1
rlabel polysilicon 149 -75 149 -75 0 3
rlabel polysilicon 156 -69 156 -69 0 1
rlabel polysilicon 156 -75 156 -75 0 3
rlabel polysilicon 163 -69 163 -69 0 1
rlabel polysilicon 163 -75 163 -75 0 3
rlabel polysilicon 173 -69 173 -69 0 2
rlabel polysilicon 184 -69 184 -69 0 1
rlabel polysilicon 184 -75 184 -75 0 3
rlabel polysilicon 191 -69 191 -69 0 1
rlabel polysilicon 30 -96 30 -96 0 1
rlabel polysilicon 30 -102 30 -102 0 3
rlabel polysilicon 37 -96 37 -96 0 1
rlabel polysilicon 40 -96 40 -96 0 2
rlabel polysilicon 40 -102 40 -102 0 4
rlabel polysilicon 44 -96 44 -96 0 1
rlabel polysilicon 47 -102 47 -102 0 4
rlabel polysilicon 51 -96 51 -96 0 1
rlabel polysilicon 51 -102 51 -102 0 3
rlabel polysilicon 58 -96 58 -96 0 1
rlabel polysilicon 58 -102 58 -102 0 3
rlabel polysilicon 65 -96 65 -96 0 1
rlabel polysilicon 65 -102 65 -102 0 3
rlabel polysilicon 72 -96 72 -96 0 1
rlabel polysilicon 72 -102 72 -102 0 3
rlabel polysilicon 82 -96 82 -96 0 2
rlabel polysilicon 79 -102 79 -102 0 3
rlabel polysilicon 86 -96 86 -96 0 1
rlabel polysilicon 89 -96 89 -96 0 2
rlabel polysilicon 86 -102 86 -102 0 3
rlabel polysilicon 89 -102 89 -102 0 4
rlabel polysilicon 93 -96 93 -96 0 1
rlabel polysilicon 93 -102 93 -102 0 3
rlabel polysilicon 100 -96 100 -96 0 1
rlabel polysilicon 103 -96 103 -96 0 2
rlabel polysilicon 100 -102 100 -102 0 3
rlabel polysilicon 107 -96 107 -96 0 1
rlabel polysilicon 107 -102 107 -102 0 3
rlabel polysilicon 114 -96 114 -96 0 1
rlabel polysilicon 114 -102 114 -102 0 3
rlabel polysilicon 121 -102 121 -102 0 3
rlabel polysilicon 124 -102 124 -102 0 4
rlabel polysilicon 128 -96 128 -96 0 1
rlabel polysilicon 128 -102 128 -102 0 3
rlabel polysilicon 135 -96 135 -96 0 1
rlabel polysilicon 135 -102 135 -102 0 3
rlabel polysilicon 142 -96 142 -96 0 1
rlabel polysilicon 142 -102 142 -102 0 3
rlabel polysilicon 149 -96 149 -96 0 1
rlabel polysilicon 149 -102 149 -102 0 3
rlabel polysilicon 156 -96 156 -96 0 1
rlabel polysilicon 156 -102 156 -102 0 3
rlabel polysilicon 184 -96 184 -96 0 1
rlabel polysilicon 2 -123 2 -123 0 1
rlabel polysilicon 2 -129 2 -129 0 3
rlabel polysilicon 9 -123 9 -123 0 1
rlabel polysilicon 9 -129 9 -129 0 3
rlabel polysilicon 16 -123 16 -123 0 1
rlabel polysilicon 16 -129 16 -129 0 3
rlabel polysilicon 23 -123 23 -123 0 1
rlabel polysilicon 23 -129 23 -129 0 3
rlabel polysilicon 30 -123 30 -123 0 1
rlabel polysilicon 33 -123 33 -123 0 2
rlabel polysilicon 37 -123 37 -123 0 1
rlabel polysilicon 37 -129 37 -129 0 3
rlabel polysilicon 44 -123 44 -123 0 1
rlabel polysilicon 47 -123 47 -123 0 2
rlabel polysilicon 44 -129 44 -129 0 3
rlabel polysilicon 47 -129 47 -129 0 4
rlabel polysilicon 51 -123 51 -123 0 1
rlabel polysilicon 51 -129 51 -129 0 3
rlabel polysilicon 58 -123 58 -123 0 1
rlabel polysilicon 58 -129 58 -129 0 3
rlabel polysilicon 65 -123 65 -123 0 1
rlabel polysilicon 68 -123 68 -123 0 2
rlabel polysilicon 72 -123 72 -123 0 1
rlabel polysilicon 72 -129 72 -129 0 3
rlabel polysilicon 82 -123 82 -123 0 2
rlabel polysilicon 82 -129 82 -129 0 4
rlabel polysilicon 86 -123 86 -123 0 1
rlabel polysilicon 89 -123 89 -123 0 2
rlabel polysilicon 89 -129 89 -129 0 4
rlabel polysilicon 93 -123 93 -123 0 1
rlabel polysilicon 96 -123 96 -123 0 2
rlabel polysilicon 93 -129 93 -129 0 3
rlabel polysilicon 100 -123 100 -123 0 1
rlabel polysilicon 100 -129 100 -129 0 3
rlabel polysilicon 107 -123 107 -123 0 1
rlabel polysilicon 107 -129 107 -129 0 3
rlabel polysilicon 114 -123 114 -123 0 1
rlabel polysilicon 117 -123 117 -123 0 2
rlabel polysilicon 117 -129 117 -129 0 4
rlabel polysilicon 121 -123 121 -123 0 1
rlabel polysilicon 121 -129 121 -129 0 3
rlabel polysilicon 131 -123 131 -123 0 2
rlabel polysilicon 131 -129 131 -129 0 4
rlabel polysilicon 135 -123 135 -123 0 1
rlabel polysilicon 138 -123 138 -123 0 2
rlabel polysilicon 145 -129 145 -129 0 4
rlabel polysilicon 149 -123 149 -123 0 1
rlabel polysilicon 149 -129 149 -129 0 3
rlabel polysilicon 156 -123 156 -123 0 1
rlabel polysilicon 156 -129 156 -129 0 3
rlabel polysilicon 163 -123 163 -123 0 1
rlabel polysilicon 163 -129 163 -129 0 3
rlabel polysilicon 170 -123 170 -123 0 1
rlabel polysilicon 170 -129 170 -129 0 3
rlabel polysilicon 177 -123 177 -123 0 1
rlabel polysilicon 177 -129 177 -129 0 3
rlabel polysilicon 184 -123 184 -123 0 1
rlabel polysilicon 184 -129 184 -129 0 3
rlabel polysilicon 16 -154 16 -154 0 1
rlabel polysilicon 16 -160 16 -160 0 3
rlabel polysilicon 23 -154 23 -154 0 1
rlabel polysilicon 23 -160 23 -160 0 3
rlabel polysilicon 33 -154 33 -154 0 2
rlabel polysilicon 33 -160 33 -160 0 4
rlabel polysilicon 37 -154 37 -154 0 1
rlabel polysilicon 37 -160 37 -160 0 3
rlabel polysilicon 44 -154 44 -154 0 1
rlabel polysilicon 47 -160 47 -160 0 4
rlabel polysilicon 51 -154 51 -154 0 1
rlabel polysilicon 54 -154 54 -154 0 2
rlabel polysilicon 54 -160 54 -160 0 4
rlabel polysilicon 58 -154 58 -154 0 1
rlabel polysilicon 58 -160 58 -160 0 3
rlabel polysilicon 65 -154 65 -154 0 1
rlabel polysilicon 65 -160 65 -160 0 3
rlabel polysilicon 72 -154 72 -154 0 1
rlabel polysilicon 72 -160 72 -160 0 3
rlabel polysilicon 79 -154 79 -154 0 1
rlabel polysilicon 79 -160 79 -160 0 3
rlabel polysilicon 86 -154 86 -154 0 1
rlabel polysilicon 89 -154 89 -154 0 2
rlabel polysilicon 86 -160 86 -160 0 3
rlabel polysilicon 89 -160 89 -160 0 4
rlabel polysilicon 93 -154 93 -154 0 1
rlabel polysilicon 96 -154 96 -154 0 2
rlabel polysilicon 93 -160 93 -160 0 3
rlabel polysilicon 96 -160 96 -160 0 4
rlabel polysilicon 100 -154 100 -154 0 1
rlabel polysilicon 103 -154 103 -154 0 2
rlabel polysilicon 100 -160 100 -160 0 3
rlabel polysilicon 103 -160 103 -160 0 4
rlabel polysilicon 107 -154 107 -154 0 1
rlabel polysilicon 107 -160 107 -160 0 3
rlabel polysilicon 114 -154 114 -154 0 1
rlabel polysilicon 117 -154 117 -154 0 2
rlabel polysilicon 114 -160 114 -160 0 3
rlabel polysilicon 117 -160 117 -160 0 4
rlabel polysilicon 121 -154 121 -154 0 1
rlabel polysilicon 121 -160 121 -160 0 3
rlabel polysilicon 131 -154 131 -154 0 2
rlabel polysilicon 128 -160 128 -160 0 3
rlabel polysilicon 135 -160 135 -160 0 3
rlabel polysilicon 138 -160 138 -160 0 4
rlabel polysilicon 142 -154 142 -154 0 1
rlabel polysilicon 142 -160 142 -160 0 3
rlabel polysilicon 149 -154 149 -154 0 1
rlabel polysilicon 149 -160 149 -160 0 3
rlabel polysilicon 156 -154 156 -154 0 1
rlabel polysilicon 156 -160 156 -160 0 3
rlabel polysilicon 163 -154 163 -154 0 1
rlabel polysilicon 163 -160 163 -160 0 3
rlabel polysilicon 170 -154 170 -154 0 1
rlabel polysilicon 170 -160 170 -160 0 3
rlabel polysilicon 177 -154 177 -154 0 1
rlabel polysilicon 177 -160 177 -160 0 3
rlabel polysilicon 184 -154 184 -154 0 1
rlabel polysilicon 184 -160 184 -160 0 3
rlabel polysilicon 33 -187 33 -187 0 2
rlabel polysilicon 40 -187 40 -187 0 2
rlabel polysilicon 44 -187 44 -187 0 1
rlabel polysilicon 47 -193 47 -193 0 4
rlabel polysilicon 51 -187 51 -187 0 1
rlabel polysilicon 51 -193 51 -193 0 3
rlabel polysilicon 61 -187 61 -187 0 2
rlabel polysilicon 65 -187 65 -187 0 1
rlabel polysilicon 65 -193 65 -193 0 3
rlabel polysilicon 75 -187 75 -187 0 2
rlabel polysilicon 72 -193 72 -193 0 3
rlabel polysilicon 79 -187 79 -187 0 1
rlabel polysilicon 79 -193 79 -193 0 3
rlabel polysilicon 86 -193 86 -193 0 3
rlabel polysilicon 89 -193 89 -193 0 4
rlabel polysilicon 96 -187 96 -187 0 2
rlabel polysilicon 93 -193 93 -193 0 3
rlabel polysilicon 96 -193 96 -193 0 4
rlabel polysilicon 100 -187 100 -187 0 1
rlabel polysilicon 100 -193 100 -193 0 3
rlabel polysilicon 107 -187 107 -187 0 1
rlabel polysilicon 107 -193 107 -193 0 3
rlabel polysilicon 114 -187 114 -187 0 1
rlabel polysilicon 114 -193 114 -193 0 3
rlabel polysilicon 121 -187 121 -187 0 1
rlabel polysilicon 124 -187 124 -187 0 2
rlabel polysilicon 121 -193 121 -193 0 3
rlabel polysilicon 128 -187 128 -187 0 1
rlabel polysilicon 128 -193 128 -193 0 3
rlabel polysilicon 135 -187 135 -187 0 1
rlabel polysilicon 135 -193 135 -193 0 3
rlabel polysilicon 145 -193 145 -193 0 4
rlabel polysilicon 149 -187 149 -187 0 1
rlabel polysilicon 149 -193 149 -193 0 3
rlabel polysilicon 156 -187 156 -187 0 1
rlabel polysilicon 156 -193 156 -193 0 3
rlabel polysilicon 163 -187 163 -187 0 1
rlabel polysilicon 163 -193 163 -193 0 3
rlabel polysilicon 170 -187 170 -187 0 1
rlabel polysilicon 170 -193 170 -193 0 3
rlabel polysilicon 177 -187 177 -187 0 1
rlabel polysilicon 177 -193 177 -193 0 3
rlabel polysilicon 184 -187 184 -187 0 1
rlabel polysilicon 184 -193 184 -193 0 3
rlabel polysilicon 51 -206 51 -206 0 1
rlabel polysilicon 51 -212 51 -212 0 3
rlabel polysilicon 58 -206 58 -206 0 1
rlabel polysilicon 58 -212 58 -212 0 3
rlabel polysilicon 68 -206 68 -206 0 2
rlabel polysilicon 65 -212 65 -212 0 3
rlabel polysilicon 68 -212 68 -212 0 4
rlabel polysilicon 72 -206 72 -206 0 1
rlabel polysilicon 72 -212 72 -212 0 3
rlabel polysilicon 79 -206 79 -206 0 1
rlabel polysilicon 79 -212 79 -212 0 3
rlabel polysilicon 82 -212 82 -212 0 4
rlabel polysilicon 86 -206 86 -206 0 1
rlabel polysilicon 86 -212 86 -212 0 3
rlabel polysilicon 93 -206 93 -206 0 1
rlabel polysilicon 93 -212 93 -212 0 3
rlabel polysilicon 100 -206 100 -206 0 1
rlabel polysilicon 100 -212 100 -212 0 3
rlabel polysilicon 110 -206 110 -206 0 2
rlabel polysilicon 117 -206 117 -206 0 2
rlabel polysilicon 114 -212 114 -212 0 3
rlabel polysilicon 121 -206 121 -206 0 1
rlabel polysilicon 121 -212 121 -212 0 3
rlabel polysilicon 128 -206 128 -206 0 1
rlabel polysilicon 128 -212 128 -212 0 3
rlabel polysilicon 135 -206 135 -206 0 1
rlabel polysilicon 135 -212 135 -212 0 3
rlabel polysilicon 142 -206 142 -206 0 1
rlabel polysilicon 142 -212 142 -212 0 3
rlabel polysilicon 145 -212 145 -212 0 4
rlabel polysilicon 152 -206 152 -206 0 2
rlabel polysilicon 149 -212 149 -212 0 3
rlabel polysilicon 152 -212 152 -212 0 4
rlabel polysilicon 156 -206 156 -206 0 1
rlabel polysilicon 58 -223 58 -223 0 1
rlabel polysilicon 58 -229 58 -229 0 3
rlabel polysilicon 68 -229 68 -229 0 4
rlabel polysilicon 75 -223 75 -223 0 2
rlabel polysilicon 79 -229 79 -229 0 3
rlabel polysilicon 86 -223 86 -223 0 1
rlabel polysilicon 86 -229 86 -229 0 3
rlabel polysilicon 124 -223 124 -223 0 2
rlabel polysilicon 124 -229 124 -229 0 4
rlabel polysilicon 135 -223 135 -223 0 1
rlabel polysilicon 135 -229 135 -229 0 3
rlabel polysilicon 159 -223 159 -223 0 2
rlabel polysilicon 156 -229 156 -229 0 3
rlabel polysilicon 156 -240 156 -240 0 3
rlabel polysilicon 163 -234 163 -234 0 1
rlabel polysilicon 163 -240 163 -240 0 3
rlabel metal2 86 1 86 1 0 net=223
rlabel metal2 51 -10 51 -10 0 net=139
rlabel metal2 65 -10 65 -10 0 net=129
rlabel metal2 82 -10 82 -10 0 net=36
rlabel metal2 93 -10 93 -10 0 net=169
rlabel metal2 100 -10 100 -10 0 net=224
rlabel metal2 121 -10 121 -10 0 net=177
rlabel metal2 149 -10 149 -10 0 net=32
rlabel metal2 79 -12 79 -12 0 net=227
rlabel metal2 100 -12 100 -12 0 net=155
rlabel metal2 142 -12 142 -12 0 net=183
rlabel metal2 79 -14 79 -14 0 net=231
rlabel metal2 103 -16 103 -16 0 net=161
rlabel metal2 30 -27 30 -27 0 net=219
rlabel metal2 37 -27 37 -27 0 net=131
rlabel metal2 68 -27 68 -27 0 net=125
rlabel metal2 79 -27 79 -27 0 net=18
rlabel metal2 107 -27 107 -27 0 net=157
rlabel metal2 23 -29 23 -29 0 net=249
rlabel metal2 110 -29 110 -29 0 net=189
rlabel metal2 51 -31 51 -31 0 net=141
rlabel metal2 79 -31 79 -31 0 net=143
rlabel metal2 135 -31 135 -31 0 net=233
rlabel metal2 86 -33 86 -33 0 net=228
rlabel metal2 93 -33 93 -33 0 net=170
rlabel metal2 128 -33 128 -33 0 net=179
rlabel metal2 149 -33 149 -33 0 net=281
rlabel metal2 86 -35 86 -35 0 net=113
rlabel metal2 100 -35 100 -35 0 net=197
rlabel metal2 142 -35 142 -35 0 net=185
rlabel metal2 159 -35 159 -35 0 net=309
rlabel metal2 114 -37 114 -37 0 net=163
rlabel metal2 16 -48 16 -48 0 net=221
rlabel metal2 37 -48 37 -48 0 net=132
rlabel metal2 86 -48 86 -48 0 net=158
rlabel metal2 173 -48 173 -48 0 net=282
rlabel metal2 23 -50 23 -50 0 net=250
rlabel metal2 72 -50 72 -50 0 net=126
rlabel metal2 100 -50 100 -50 0 net=164
rlabel metal2 163 -50 163 -50 0 net=235
rlabel metal2 23 -52 23 -52 0 net=127
rlabel metal2 96 -52 96 -52 0 net=149
rlabel metal2 40 -54 40 -54 0 net=28
rlabel metal2 103 -54 103 -54 0 net=186
rlabel metal2 44 -56 44 -56 0 net=82
rlabel metal2 107 -56 107 -56 0 net=190
rlabel metal2 37 -58 37 -58 0 net=225
rlabel metal2 51 -58 51 -58 0 net=142
rlabel metal2 93 -58 93 -58 0 net=115
rlabel metal2 114 -58 114 -58 0 net=310
rlabel metal2 51 -60 51 -60 0 net=111
rlabel metal2 72 -60 72 -60 0 net=84
rlabel metal2 117 -60 117 -60 0 net=159
rlabel metal2 184 -60 184 -60 0 net=283
rlabel metal2 58 -62 58 -62 0 net=85
rlabel metal2 100 -62 100 -62 0 net=93
rlabel metal2 128 -62 128 -62 0 net=199
rlabel metal2 128 -62 128 -62 0 net=199
rlabel metal2 135 -62 135 -62 0 net=181
rlabel metal2 30 -64 30 -64 0 net=107
rlabel metal2 121 -64 121 -64 0 net=145
rlabel metal2 68 -66 68 -66 0 net=123
rlabel metal2 16 -77 16 -77 0 net=222
rlabel metal2 51 -77 51 -77 0 net=112
rlabel metal2 75 -77 75 -77 0 net=116
rlabel metal2 114 -77 114 -77 0 net=236
rlabel metal2 184 -77 184 -77 0 net=284
rlabel metal2 184 -77 184 -77 0 net=284
rlabel metal2 23 -79 23 -79 0 net=128
rlabel metal2 82 -79 82 -79 0 net=124
rlabel metal2 128 -79 128 -79 0 net=201
rlabel metal2 128 -79 128 -79 0 net=201
rlabel metal2 30 -81 30 -81 0 net=108
rlabel metal2 86 -81 86 -81 0 net=251
rlabel metal2 96 -81 96 -81 0 net=146
rlabel metal2 30 -83 30 -83 0 net=165
rlabel metal2 40 -83 40 -83 0 net=226
rlabel metal2 65 -83 65 -83 0 net=121
rlabel metal2 86 -83 86 -83 0 net=147
rlabel metal2 117 -83 117 -83 0 net=182
rlabel metal2 44 -85 44 -85 0 net=133
rlabel metal2 89 -85 89 -85 0 net=245
rlabel metal2 142 -85 142 -85 0 net=150
rlabel metal2 79 -87 79 -87 0 net=257
rlabel metal2 100 -89 100 -89 0 net=95
rlabel metal2 103 -91 103 -91 0 net=160
rlabel metal2 100 -93 100 -93 0 net=261
rlabel metal2 2 -104 2 -104 0 net=303
rlabel metal2 37 -104 37 -104 0 net=135
rlabel metal2 58 -104 58 -104 0 net=56
rlabel metal2 86 -104 86 -104 0 net=96
rlabel metal2 142 -104 142 -104 0 net=259
rlabel metal2 9 -106 9 -106 0 net=295
rlabel metal2 121 -106 121 -106 0 net=202
rlabel metal2 131 -106 131 -106 0 net=265
rlabel metal2 16 -108 16 -108 0 net=167
rlabel metal2 40 -108 40 -108 0 net=27
rlabel metal2 51 -108 51 -108 0 net=151
rlabel metal2 23 -110 23 -110 0 net=193
rlabel metal2 44 -110 44 -110 0 net=15
rlabel metal2 124 -110 124 -110 0 net=47
rlabel metal2 149 -110 149 -110 0 net=263
rlabel metal2 47 -112 47 -112 0 net=81
rlabel metal2 72 -112 72 -112 0 net=122
rlabel metal2 89 -112 89 -112 0 net=148
rlabel metal2 114 -112 114 -112 0 net=247
rlabel metal2 58 -114 58 -114 0 net=187
rlabel metal2 107 -114 107 -114 0 net=205
rlabel metal2 135 -114 135 -114 0 net=269
rlabel metal2 65 -116 65 -116 0 net=88
rlabel metal2 89 -116 89 -116 0 net=285
rlabel metal2 65 -118 65 -118 0 net=91
rlabel metal2 93 -118 93 -118 0 net=253
rlabel metal2 93 -120 93 -120 0 net=101
rlabel metal2 2 -131 2 -131 0 net=304
rlabel metal2 58 -131 58 -131 0 net=188
rlabel metal2 82 -131 82 -131 0 net=2
rlabel metal2 117 -131 117 -131 0 net=248
rlabel metal2 16 -133 16 -133 0 net=168
rlabel metal2 65 -133 65 -133 0 net=97
rlabel metal2 131 -133 131 -133 0 net=239
rlabel metal2 16 -135 16 -135 0 net=293
rlabel metal2 37 -135 37 -135 0 net=136
rlabel metal2 72 -135 72 -135 0 net=92
rlabel metal2 93 -135 93 -135 0 net=260
rlabel metal2 9 -137 9 -137 0 net=296
rlabel metal2 93 -137 93 -137 0 net=211
rlabel metal2 145 -137 145 -137 0 net=264
rlabel metal2 23 -139 23 -139 0 net=195
rlabel metal2 23 -139 23 -139 0 net=195
rlabel metal2 51 -139 51 -139 0 net=153
rlabel metal2 86 -139 86 -139 0 net=102
rlabel metal2 163 -139 163 -139 0 net=267
rlabel metal2 37 -141 37 -141 0 net=191
rlabel metal2 121 -141 121 -141 0 net=287
rlabel metal2 51 -143 51 -143 0 net=203
rlabel metal2 96 -143 96 -143 0 net=254
rlabel metal2 170 -143 170 -143 0 net=271
rlabel metal2 54 -145 54 -145 0 net=243
rlabel metal2 107 -147 107 -147 0 net=207
rlabel metal2 107 -149 107 -149 0 net=171
rlabel metal2 117 -151 117 -151 0 net=299
rlabel metal2 16 -162 16 -162 0 net=294
rlabel metal2 51 -162 51 -162 0 net=109
rlabel metal2 114 -162 114 -162 0 net=244
rlabel metal2 23 -164 23 -164 0 net=196
rlabel metal2 37 -164 37 -164 0 net=192
rlabel metal2 58 -164 58 -164 0 net=204
rlabel metal2 121 -164 121 -164 0 net=209
rlabel metal2 33 -166 33 -166 0 net=6
rlabel metal2 61 -166 61 -166 0 net=172
rlabel metal2 114 -166 114 -166 0 net=213
rlabel metal2 40 -168 40 -168 0 net=37
rlabel metal2 100 -168 100 -168 0 net=272
rlabel metal2 65 -170 65 -170 0 net=99
rlabel metal2 121 -170 121 -170 0 net=297
rlabel metal2 65 -172 65 -172 0 net=173
rlabel metal2 79 -172 79 -172 0 net=137
rlabel metal2 79 -172 79 -172 0 net=137
rlabel metal2 128 -172 128 -172 0 net=268
rlabel metal2 72 -174 72 -174 0 net=154
rlabel metal2 96 -174 96 -174 0 net=291
rlabel metal2 96 -176 96 -176 0 net=117
rlabel metal2 128 -176 128 -176 0 net=277
rlabel metal2 135 -178 135 -178 0 net=288
rlabel metal2 135 -180 135 -180 0 net=241
rlabel metal2 177 -180 177 -180 0 net=301
rlabel metal2 89 -182 89 -182 0 net=273
rlabel metal2 124 -184 124 -184 0 net=307
rlabel metal2 51 -195 51 -195 0 net=110
rlabel metal2 79 -195 79 -195 0 net=138
rlabel metal2 96 -195 96 -195 0 net=214
rlabel metal2 121 -195 121 -195 0 net=242
rlabel metal2 142 -195 142 -195 0 net=292
rlabel metal2 47 -197 47 -197 0 net=255
rlabel metal2 58 -197 58 -197 0 net=215
rlabel metal2 86 -197 86 -197 0 net=210
rlabel metal2 65 -199 65 -199 0 net=175
rlabel metal2 89 -199 89 -199 0 net=100
rlabel metal2 110 -199 110 -199 0 net=289
rlabel metal2 145 -199 145 -199 0 net=298
rlabel metal2 68 -201 68 -201 0 net=103
rlabel metal2 93 -201 93 -201 0 net=229
rlabel metal2 121 -201 121 -201 0 net=279
rlabel metal2 152 -201 152 -201 0 net=302
rlabel metal2 100 -203 100 -203 0 net=119
rlabel metal2 128 -203 128 -203 0 net=275
rlabel metal2 156 -203 156 -203 0 net=308
rlabel metal2 51 -214 51 -214 0 net=256
rlabel metal2 72 -214 72 -214 0 net=176
rlabel metal2 79 -214 79 -214 0 net=120
rlabel metal2 114 -214 114 -214 0 net=290
rlabel metal2 149 -214 149 -214 0 net=67
rlabel metal2 58 -216 58 -216 0 net=217
rlabel metal2 58 -216 58 -216 0 net=217
rlabel metal2 65 -216 65 -216 0 net=49
rlabel metal2 86 -216 86 -216 0 net=105
rlabel metal2 86 -216 86 -216 0 net=105
rlabel metal2 93 -216 93 -216 0 net=230
rlabel metal2 128 -216 128 -216 0 net=276
rlabel metal2 121 -218 121 -218 0 net=280
rlabel metal2 135 -220 135 -220 0 net=237
rlabel metal2 58 -231 58 -231 0 net=218
rlabel metal2 79 -231 79 -231 0 net=106
rlabel metal2 124 -231 124 -231 0 net=238
rlabel metal2 156 -231 156 -231 0 net=305
rlabel metal2 156 -242 156 -242 0 net=306
<< end >>
