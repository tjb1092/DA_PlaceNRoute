magic
tech scmos
timestamp 1555016718 
<< pdiffusion >>
rect 1 -8 7 -2
rect 8 -8 14 -2
rect 15 -8 21 -2
rect 43 -8 46 -2
rect 50 -8 56 -2
rect 57 -8 63 -2
rect 64 -8 67 -2
rect 71 -8 77 -2
rect 78 -8 84 -2
rect 1 -23 7 -17
rect 15 -23 21 -17
rect 22 -23 28 -17
rect 29 -23 32 -17
rect 36 -23 39 -17
rect 43 -23 49 -17
rect 50 -23 53 -17
rect 57 -23 63 -17
rect 64 -23 67 -17
rect 71 -23 77 -17
rect 78 -23 81 -17
rect 85 -23 91 -17
rect 92 -23 95 -17
rect 106 -23 112 -17
rect 113 -23 119 -17
rect 1 -46 7 -40
rect 8 -46 11 -40
rect 15 -46 18 -40
rect 22 -46 25 -40
rect 29 -46 35 -40
rect 36 -46 42 -40
rect 43 -46 49 -40
rect 50 -46 56 -40
rect 57 -46 60 -40
rect 64 -46 70 -40
rect 71 -46 77 -40
rect 78 -46 81 -40
rect 85 -46 91 -40
rect 92 -46 95 -40
rect 99 -46 105 -40
rect 106 -46 109 -40
rect 113 -46 116 -40
rect 120 -46 123 -40
rect 127 -46 130 -40
rect 134 -46 137 -40
rect 141 -46 144 -40
rect 1 -73 7 -67
rect 8 -73 11 -67
rect 15 -73 18 -67
rect 22 -73 28 -67
rect 29 -73 35 -67
rect 36 -73 39 -67
rect 43 -73 49 -67
rect 50 -73 53 -67
rect 57 -73 60 -67
rect 64 -73 70 -67
rect 71 -73 74 -67
rect 78 -73 84 -67
rect 85 -73 91 -67
rect 92 -73 95 -67
rect 99 -73 102 -67
rect 106 -73 109 -67
rect 113 -73 116 -67
rect 120 -73 126 -67
rect 127 -73 133 -67
rect 134 -73 137 -67
rect 1 -96 4 -90
rect 8 -96 14 -90
rect 15 -96 21 -90
rect 22 -96 25 -90
rect 29 -96 32 -90
rect 36 -96 39 -90
rect 43 -96 46 -90
rect 50 -96 56 -90
rect 57 -96 63 -90
rect 64 -96 70 -90
rect 71 -96 74 -90
rect 78 -96 81 -90
rect 85 -96 91 -90
rect 92 -96 95 -90
rect 99 -96 105 -90
rect 106 -96 109 -90
rect 113 -96 116 -90
rect 120 -96 126 -90
rect 127 -96 130 -90
rect 134 -96 137 -90
rect 141 -96 144 -90
rect 148 -96 154 -90
rect 15 -129 21 -123
rect 22 -129 25 -123
rect 29 -129 35 -123
rect 36 -129 39 -123
rect 43 -129 49 -123
rect 50 -129 53 -123
rect 57 -129 60 -123
rect 64 -129 70 -123
rect 71 -129 74 -123
rect 78 -129 84 -123
rect 85 -129 91 -123
rect 92 -129 95 -123
rect 99 -129 105 -123
rect 106 -129 109 -123
rect 113 -129 116 -123
rect 120 -129 123 -123
rect 127 -129 133 -123
rect 134 -129 137 -123
rect 141 -129 144 -123
rect 148 -129 151 -123
rect 155 -129 158 -123
rect 162 -129 165 -123
rect 169 -129 175 -123
rect 1 -156 4 -150
rect 8 -156 11 -150
rect 15 -156 18 -150
rect 22 -156 25 -150
rect 29 -156 32 -150
rect 36 -156 42 -150
rect 43 -156 49 -150
rect 50 -156 56 -150
rect 57 -156 63 -150
rect 64 -156 70 -150
rect 71 -156 77 -150
rect 78 -156 81 -150
rect 85 -156 88 -150
rect 92 -156 98 -150
rect 99 -156 102 -150
rect 106 -156 112 -150
rect 113 -156 116 -150
rect 120 -156 126 -150
rect 127 -156 130 -150
rect 134 -156 137 -150
rect 141 -156 144 -150
rect 148 -156 151 -150
rect 155 -156 158 -150
rect 162 -156 165 -150
rect 169 -156 172 -150
rect 176 -156 179 -150
rect 183 -156 186 -150
rect 190 -156 193 -150
rect 197 -156 203 -150
rect 204 -156 207 -150
rect 8 -187 14 -181
rect 22 -187 25 -181
rect 36 -187 42 -181
rect 43 -187 49 -181
rect 57 -187 60 -181
rect 64 -187 70 -181
rect 71 -187 77 -181
rect 78 -187 81 -181
rect 85 -187 91 -181
rect 92 -187 98 -181
rect 106 -187 112 -181
rect 113 -187 116 -181
rect 127 -187 130 -181
rect 134 -187 137 -181
rect 141 -187 147 -181
rect 162 -187 168 -181
rect 169 -187 172 -181
rect 1 -212 4 -206
rect 8 -212 11 -206
rect 15 -212 18 -206
rect 22 -212 25 -206
rect 29 -212 32 -206
rect 36 -212 42 -206
rect 43 -212 49 -206
rect 50 -212 56 -206
rect 57 -212 63 -206
rect 64 -212 70 -206
rect 71 -212 74 -206
rect 78 -212 84 -206
rect 85 -212 88 -206
rect 92 -212 95 -206
rect 99 -212 102 -206
rect 106 -212 109 -206
rect 113 -212 119 -206
rect 120 -212 123 -206
rect 127 -212 133 -206
rect 134 -212 137 -206
rect 141 -212 144 -206
rect 148 -212 151 -206
rect 155 -212 161 -206
rect 15 -237 18 -231
rect 22 -237 28 -231
rect 29 -237 35 -231
rect 36 -237 42 -231
rect 43 -237 46 -231
rect 50 -237 56 -231
rect 57 -237 63 -231
rect 64 -237 70 -231
rect 71 -237 74 -231
rect 78 -237 84 -231
rect 85 -237 91 -231
rect 99 -237 105 -231
<< polysilicon >>
rect 44 -3 45 -1
rect 44 -9 45 -7
rect 51 -9 52 -7
rect 58 -3 59 -1
rect 58 -9 59 -7
rect 65 -3 66 -1
rect 65 -9 66 -7
rect 75 -9 76 -7
rect 79 -3 80 -1
rect 26 -24 27 -22
rect 30 -18 31 -16
rect 30 -24 31 -22
rect 37 -18 38 -16
rect 37 -24 38 -22
rect 44 -18 45 -16
rect 44 -24 45 -22
rect 47 -24 48 -22
rect 51 -18 52 -16
rect 51 -24 52 -22
rect 61 -18 62 -16
rect 58 -24 59 -22
rect 61 -24 62 -22
rect 65 -18 66 -16
rect 65 -24 66 -22
rect 72 -18 73 -16
rect 79 -18 80 -16
rect 79 -24 80 -22
rect 86 -18 87 -16
rect 86 -24 87 -22
rect 93 -18 94 -16
rect 93 -24 94 -22
rect 110 -18 111 -16
rect 114 -24 115 -22
rect 9 -41 10 -39
rect 9 -47 10 -45
rect 16 -41 17 -39
rect 16 -47 17 -45
rect 23 -41 24 -39
rect 23 -47 24 -45
rect 30 -41 31 -39
rect 37 -41 38 -39
rect 37 -47 38 -45
rect 44 -41 45 -39
rect 47 -47 48 -45
rect 54 -47 55 -45
rect 58 -41 59 -39
rect 58 -47 59 -45
rect 68 -41 69 -39
rect 65 -47 66 -45
rect 68 -47 69 -45
rect 72 -41 73 -39
rect 75 -41 76 -39
rect 72 -47 73 -45
rect 75 -47 76 -45
rect 79 -41 80 -39
rect 79 -47 80 -45
rect 86 -41 87 -39
rect 89 -41 90 -39
rect 86 -47 87 -45
rect 93 -41 94 -39
rect 93 -47 94 -45
rect 100 -41 101 -39
rect 103 -47 104 -45
rect 107 -41 108 -39
rect 107 -47 108 -45
rect 114 -41 115 -39
rect 114 -47 115 -45
rect 121 -41 122 -39
rect 121 -47 122 -45
rect 128 -41 129 -39
rect 128 -47 129 -45
rect 135 -41 136 -39
rect 135 -47 136 -45
rect 142 -41 143 -39
rect 142 -47 143 -45
rect 9 -68 10 -66
rect 9 -74 10 -72
rect 16 -68 17 -66
rect 16 -74 17 -72
rect 23 -68 24 -66
rect 26 -68 27 -66
rect 23 -74 24 -72
rect 30 -68 31 -66
rect 33 -68 34 -66
rect 30 -74 31 -72
rect 37 -68 38 -66
rect 37 -74 38 -72
rect 47 -68 48 -66
rect 44 -74 45 -72
rect 47 -74 48 -72
rect 51 -68 52 -66
rect 51 -74 52 -72
rect 58 -68 59 -66
rect 58 -74 59 -72
rect 65 -68 66 -66
rect 68 -68 69 -66
rect 68 -74 69 -72
rect 72 -68 73 -66
rect 72 -74 73 -72
rect 79 -68 80 -66
rect 82 -68 83 -66
rect 79 -74 80 -72
rect 86 -68 87 -66
rect 89 -68 90 -66
rect 89 -74 90 -72
rect 93 -68 94 -66
rect 93 -74 94 -72
rect 100 -68 101 -66
rect 100 -74 101 -72
rect 107 -68 108 -66
rect 107 -74 108 -72
rect 114 -68 115 -66
rect 114 -74 115 -72
rect 124 -74 125 -72
rect 131 -68 132 -66
rect 131 -74 132 -72
rect 135 -68 136 -66
rect 135 -74 136 -72
rect 2 -91 3 -89
rect 2 -97 3 -95
rect 9 -91 10 -89
rect 19 -91 20 -89
rect 16 -97 17 -95
rect 23 -91 24 -89
rect 23 -97 24 -95
rect 30 -91 31 -89
rect 30 -97 31 -95
rect 37 -91 38 -89
rect 37 -97 38 -95
rect 44 -91 45 -89
rect 44 -97 45 -95
rect 51 -91 52 -89
rect 54 -91 55 -89
rect 58 -91 59 -89
rect 61 -91 62 -89
rect 58 -97 59 -95
rect 61 -97 62 -95
rect 65 -91 66 -89
rect 68 -91 69 -89
rect 65 -97 66 -95
rect 68 -97 69 -95
rect 72 -91 73 -89
rect 72 -97 73 -95
rect 79 -91 80 -89
rect 79 -97 80 -95
rect 86 -91 87 -89
rect 89 -91 90 -89
rect 86 -97 87 -95
rect 93 -91 94 -89
rect 93 -97 94 -95
rect 100 -97 101 -95
rect 107 -91 108 -89
rect 107 -97 108 -95
rect 114 -91 115 -89
rect 114 -97 115 -95
rect 121 -91 122 -89
rect 124 -91 125 -89
rect 128 -91 129 -89
rect 128 -97 129 -95
rect 135 -91 136 -89
rect 135 -97 136 -95
rect 142 -91 143 -89
rect 142 -97 143 -95
rect 149 -91 150 -89
rect 149 -97 150 -95
rect 152 -97 153 -95
rect 19 -124 20 -122
rect 23 -124 24 -122
rect 23 -130 24 -128
rect 30 -130 31 -128
rect 33 -130 34 -128
rect 37 -124 38 -122
rect 37 -130 38 -128
rect 44 -124 45 -122
rect 47 -124 48 -122
rect 47 -130 48 -128
rect 51 -124 52 -122
rect 51 -130 52 -128
rect 58 -124 59 -122
rect 58 -130 59 -128
rect 65 -124 66 -122
rect 68 -124 69 -122
rect 65 -130 66 -128
rect 72 -124 73 -122
rect 72 -130 73 -128
rect 79 -124 80 -122
rect 82 -124 83 -122
rect 79 -130 80 -128
rect 82 -130 83 -128
rect 89 -124 90 -122
rect 86 -130 87 -128
rect 93 -124 94 -122
rect 93 -130 94 -128
rect 100 -124 101 -122
rect 103 -124 104 -122
rect 100 -130 101 -128
rect 103 -130 104 -128
rect 107 -124 108 -122
rect 107 -130 108 -128
rect 114 -124 115 -122
rect 114 -130 115 -128
rect 121 -124 122 -122
rect 121 -130 122 -128
rect 128 -124 129 -122
rect 131 -124 132 -122
rect 128 -130 129 -128
rect 135 -124 136 -122
rect 135 -130 136 -128
rect 142 -124 143 -122
rect 142 -130 143 -128
rect 149 -124 150 -122
rect 149 -130 150 -128
rect 156 -124 157 -122
rect 156 -130 157 -128
rect 163 -124 164 -122
rect 163 -130 164 -128
rect 170 -130 171 -128
rect 173 -130 174 -128
rect 2 -151 3 -149
rect 2 -157 3 -155
rect 9 -151 10 -149
rect 9 -157 10 -155
rect 16 -151 17 -149
rect 16 -157 17 -155
rect 23 -151 24 -149
rect 23 -157 24 -155
rect 30 -151 31 -149
rect 30 -157 31 -155
rect 40 -151 41 -149
rect 37 -157 38 -155
rect 40 -157 41 -155
rect 44 -151 45 -149
rect 47 -151 48 -149
rect 44 -157 45 -155
rect 47 -157 48 -155
rect 54 -157 55 -155
rect 58 -157 59 -155
rect 61 -157 62 -155
rect 65 -151 66 -149
rect 68 -157 69 -155
rect 75 -151 76 -149
rect 79 -151 80 -149
rect 79 -157 80 -155
rect 86 -151 87 -149
rect 86 -157 87 -155
rect 93 -151 94 -149
rect 93 -157 94 -155
rect 100 -151 101 -149
rect 100 -157 101 -155
rect 107 -151 108 -149
rect 110 -151 111 -149
rect 107 -157 108 -155
rect 110 -157 111 -155
rect 114 -151 115 -149
rect 114 -157 115 -155
rect 121 -157 122 -155
rect 128 -151 129 -149
rect 128 -157 129 -155
rect 135 -151 136 -149
rect 135 -157 136 -155
rect 142 -151 143 -149
rect 142 -157 143 -155
rect 149 -151 150 -149
rect 149 -157 150 -155
rect 156 -151 157 -149
rect 156 -157 157 -155
rect 163 -151 164 -149
rect 163 -157 164 -155
rect 170 -151 171 -149
rect 170 -157 171 -155
rect 177 -151 178 -149
rect 177 -157 178 -155
rect 184 -151 185 -149
rect 184 -157 185 -155
rect 191 -151 192 -149
rect 191 -157 192 -155
rect 198 -151 199 -149
rect 201 -151 202 -149
rect 201 -157 202 -155
rect 205 -151 206 -149
rect 205 -157 206 -155
rect 12 -188 13 -186
rect 23 -182 24 -180
rect 23 -188 24 -186
rect 37 -182 38 -180
rect 40 -188 41 -186
rect 47 -182 48 -180
rect 47 -188 48 -186
rect 58 -182 59 -180
rect 58 -188 59 -186
rect 65 -182 66 -180
rect 65 -188 66 -186
rect 72 -182 73 -180
rect 79 -182 80 -180
rect 79 -188 80 -186
rect 86 -182 87 -180
rect 89 -182 90 -180
rect 89 -188 90 -186
rect 96 -182 97 -180
rect 107 -182 108 -180
rect 110 -182 111 -180
rect 114 -182 115 -180
rect 114 -188 115 -186
rect 128 -182 129 -180
rect 128 -188 129 -186
rect 135 -182 136 -180
rect 135 -188 136 -186
rect 142 -182 143 -180
rect 142 -188 143 -186
rect 163 -182 164 -180
rect 166 -182 167 -180
rect 170 -182 171 -180
rect 170 -188 171 -186
rect 2 -207 3 -205
rect 2 -213 3 -211
rect 9 -207 10 -205
rect 9 -213 10 -211
rect 16 -207 17 -205
rect 16 -213 17 -211
rect 23 -207 24 -205
rect 23 -213 24 -211
rect 30 -207 31 -205
rect 30 -213 31 -211
rect 37 -207 38 -205
rect 40 -207 41 -205
rect 40 -213 41 -211
rect 44 -213 45 -211
rect 47 -213 48 -211
rect 54 -207 55 -205
rect 51 -213 52 -211
rect 58 -207 59 -205
rect 61 -207 62 -205
rect 58 -213 59 -211
rect 65 -207 66 -205
rect 68 -207 69 -205
rect 65 -213 66 -211
rect 68 -213 69 -211
rect 72 -207 73 -205
rect 72 -213 73 -211
rect 79 -207 80 -205
rect 82 -207 83 -205
rect 79 -213 80 -211
rect 82 -213 83 -211
rect 86 -207 87 -205
rect 86 -213 87 -211
rect 93 -207 94 -205
rect 93 -213 94 -211
rect 100 -207 101 -205
rect 100 -213 101 -211
rect 107 -207 108 -205
rect 107 -213 108 -211
rect 117 -207 118 -205
rect 114 -213 115 -211
rect 121 -207 122 -205
rect 121 -213 122 -211
rect 128 -213 129 -211
rect 135 -207 136 -205
rect 135 -213 136 -211
rect 142 -207 143 -205
rect 142 -213 143 -211
rect 149 -207 150 -205
rect 149 -213 150 -211
rect 159 -207 160 -205
rect 16 -232 17 -230
rect 16 -238 17 -236
rect 26 -232 27 -230
rect 33 -232 34 -230
rect 30 -238 31 -236
rect 40 -232 41 -230
rect 44 -232 45 -230
rect 44 -238 45 -236
rect 54 -232 55 -230
rect 54 -238 55 -236
rect 61 -232 62 -230
rect 61 -238 62 -236
rect 68 -232 69 -230
rect 65 -238 66 -236
rect 72 -232 73 -230
rect 72 -238 73 -236
rect 82 -232 83 -230
rect 79 -238 80 -236
rect 82 -238 83 -236
rect 86 -238 87 -236
rect 100 -232 101 -230
<< metal1 >>
rect 44 0 59 1
rect 65 0 80 1
rect 37 -11 45 -10
rect 51 -11 62 -10
rect 65 -11 73 -10
rect 79 -11 87 -10
rect 93 -11 111 -10
rect 30 -13 45 -12
rect 51 -13 76 -12
rect 58 -15 66 -14
rect 16 -26 38 -25
rect 44 -26 69 -25
rect 89 -26 108 -25
rect 114 -26 143 -25
rect 9 -28 38 -27
rect 47 -28 59 -27
rect 61 -28 122 -27
rect 26 -30 31 -29
rect 44 -30 59 -29
rect 65 -30 76 -29
rect 93 -30 129 -29
rect 23 -32 31 -31
rect 72 -32 115 -31
rect 79 -34 94 -33
rect 100 -34 136 -33
rect 79 -36 87 -35
rect 51 -38 87 -37
rect 9 -49 34 -48
rect 37 -49 66 -48
rect 68 -49 115 -48
rect 131 -49 136 -48
rect 23 -51 48 -50
rect 51 -51 90 -50
rect 103 -51 122 -50
rect 9 -53 24 -52
rect 30 -53 38 -52
rect 68 -53 94 -52
rect 107 -53 136 -52
rect 16 -55 48 -54
rect 54 -55 94 -54
rect 16 -57 27 -56
rect 65 -57 108 -56
rect 72 -59 80 -58
rect 86 -59 129 -58
rect 72 -61 83 -60
rect 86 -61 101 -60
rect 75 -63 115 -62
rect 79 -65 143 -64
rect 2 -76 31 -75
rect 47 -76 52 -75
rect 58 -76 69 -75
rect 89 -76 94 -75
rect 100 -76 143 -75
rect 9 -78 45 -77
rect 51 -78 80 -77
rect 86 -78 94 -77
rect 107 -78 111 -77
rect 114 -78 150 -77
rect 9 -80 20 -79
rect 30 -80 90 -79
rect 107 -80 136 -79
rect 16 -82 24 -81
rect 37 -82 59 -81
rect 68 -82 80 -81
rect 110 -82 136 -81
rect 23 -84 55 -83
rect 114 -84 125 -83
rect 37 -86 62 -85
rect 121 -86 132 -85
rect 44 -88 66 -87
rect 124 -88 129 -87
rect 2 -99 17 -98
rect 19 -99 59 -98
rect 61 -99 153 -98
rect 23 -101 52 -100
rect 58 -101 83 -100
rect 86 -101 115 -100
rect 149 -101 157 -100
rect 23 -103 38 -102
rect 47 -103 143 -102
rect 30 -105 66 -104
rect 68 -105 108 -104
rect 114 -105 132 -104
rect 37 -107 45 -106
rect 65 -107 122 -106
rect 128 -107 143 -106
rect 68 -109 150 -108
rect 72 -111 90 -110
rect 100 -111 104 -110
rect 128 -111 164 -110
rect 72 -113 101 -112
rect 79 -115 108 -114
rect 79 -117 136 -116
rect 93 -119 136 -118
rect 44 -121 94 -120
rect 9 -132 48 -131
rect 51 -132 80 -131
rect 100 -132 136 -131
rect 142 -132 185 -131
rect 198 -132 206 -131
rect 16 -134 45 -133
rect 72 -134 83 -133
rect 107 -134 129 -133
rect 149 -134 192 -133
rect 23 -136 66 -135
rect 75 -136 80 -135
rect 100 -136 108 -135
rect 110 -136 178 -135
rect 2 -138 66 -137
rect 103 -138 129 -137
rect 149 -138 164 -137
rect 170 -138 202 -137
rect 23 -140 59 -139
rect 86 -140 171 -139
rect 30 -142 38 -141
rect 47 -142 87 -141
rect 114 -142 136 -141
rect 156 -142 174 -141
rect 30 -144 41 -143
rect 93 -144 115 -143
rect 121 -144 164 -143
rect 33 -146 143 -145
rect 93 -148 157 -147
rect 16 -159 48 -158
rect 54 -159 164 -158
rect 166 -159 178 -158
rect 23 -161 66 -160
rect 68 -161 80 -160
rect 89 -161 101 -160
rect 107 -161 115 -160
rect 121 -161 157 -160
rect 163 -161 202 -160
rect 9 -163 80 -162
rect 93 -163 136 -162
rect 30 -165 45 -164
rect 58 -165 97 -164
rect 107 -165 115 -164
rect 128 -165 136 -164
rect 37 -167 150 -166
rect 2 -169 38 -168
rect 40 -169 73 -168
rect 86 -169 129 -168
rect 23 -171 87 -170
rect 110 -171 185 -170
rect 47 -173 59 -172
rect 61 -173 192 -172
rect 110 -175 143 -174
rect 142 -177 171 -176
rect 170 -179 206 -178
rect 2 -190 24 -189
rect 30 -190 83 -189
rect 89 -190 129 -189
rect 142 -190 171 -189
rect 9 -192 38 -191
rect 40 -192 80 -191
rect 114 -192 122 -191
rect 16 -194 55 -193
rect 58 -194 108 -193
rect 117 -194 160 -193
rect 12 -196 59 -195
rect 61 -196 150 -195
rect 23 -198 48 -197
rect 65 -198 101 -197
rect 40 -200 87 -199
rect 65 -202 73 -201
rect 79 -202 94 -201
rect 68 -204 143 -203
rect 2 -215 45 -214
rect 51 -215 108 -214
rect 128 -215 136 -214
rect 9 -217 69 -216
rect 79 -217 122 -216
rect 23 -219 59 -218
rect 61 -219 101 -218
rect 30 -221 48 -220
rect 65 -221 87 -220
rect 100 -221 150 -220
rect 33 -223 55 -222
rect 82 -223 115 -222
rect 40 -225 94 -224
rect 16 -227 41 -226
rect 44 -227 69 -226
rect 82 -227 143 -226
rect 16 -229 27 -228
rect 16 -240 31 -239
rect 44 -240 80 -239
rect 54 -242 83 -241
rect 61 -244 73 -243
rect 65 -246 87 -245
<< m2contact >>
rect 44 0 45 1
rect 58 0 59 1
rect 65 0 66 1
rect 79 0 80 1
rect 37 -11 38 -10
rect 44 -11 45 -10
rect 51 -11 52 -10
rect 61 -11 62 -10
rect 65 -11 66 -10
rect 72 -11 73 -10
rect 79 -11 80 -10
rect 86 -11 87 -10
rect 93 -11 94 -10
rect 110 -11 111 -10
rect 30 -13 31 -12
rect 44 -13 45 -12
rect 51 -13 52 -12
rect 75 -13 76 -12
rect 58 -15 59 -14
rect 65 -15 66 -14
rect 16 -26 17 -25
rect 37 -26 38 -25
rect 44 -26 45 -25
rect 68 -26 69 -25
rect 89 -26 90 -25
rect 107 -26 108 -25
rect 114 -26 115 -25
rect 142 -26 143 -25
rect 9 -28 10 -27
rect 37 -28 38 -27
rect 47 -28 48 -27
rect 58 -28 59 -27
rect 61 -28 62 -27
rect 121 -28 122 -27
rect 26 -30 27 -29
rect 30 -30 31 -29
rect 44 -30 45 -29
rect 58 -30 59 -29
rect 65 -30 66 -29
rect 75 -30 76 -29
rect 93 -30 94 -29
rect 128 -30 129 -29
rect 23 -32 24 -31
rect 30 -32 31 -31
rect 72 -32 73 -31
rect 114 -32 115 -31
rect 79 -34 80 -33
rect 93 -34 94 -33
rect 100 -34 101 -33
rect 135 -34 136 -33
rect 79 -36 80 -35
rect 86 -36 87 -35
rect 51 -38 52 -37
rect 86 -38 87 -37
rect 9 -49 10 -48
rect 33 -49 34 -48
rect 37 -49 38 -48
rect 65 -49 66 -48
rect 68 -49 69 -48
rect 114 -49 115 -48
rect 131 -49 132 -48
rect 135 -49 136 -48
rect 23 -51 24 -50
rect 47 -51 48 -50
rect 51 -51 52 -50
rect 89 -51 90 -50
rect 103 -51 104 -50
rect 121 -51 122 -50
rect 9 -53 10 -52
rect 23 -53 24 -52
rect 30 -53 31 -52
rect 37 -53 38 -52
rect 68 -53 69 -52
rect 93 -53 94 -52
rect 107 -53 108 -52
rect 135 -53 136 -52
rect 16 -55 17 -54
rect 47 -55 48 -54
rect 54 -55 55 -54
rect 93 -55 94 -54
rect 16 -57 17 -56
rect 26 -57 27 -56
rect 65 -57 66 -56
rect 107 -57 108 -56
rect 72 -59 73 -58
rect 79 -59 80 -58
rect 86 -59 87 -58
rect 128 -59 129 -58
rect 72 -61 73 -60
rect 82 -61 83 -60
rect 86 -61 87 -60
rect 100 -61 101 -60
rect 75 -63 76 -62
rect 114 -63 115 -62
rect 79 -65 80 -64
rect 142 -65 143 -64
rect 2 -76 3 -75
rect 30 -76 31 -75
rect 47 -76 48 -75
rect 51 -76 52 -75
rect 58 -76 59 -75
rect 68 -76 69 -75
rect 89 -76 90 -75
rect 93 -76 94 -75
rect 100 -76 101 -75
rect 142 -76 143 -75
rect 9 -78 10 -77
rect 44 -78 45 -77
rect 51 -78 52 -77
rect 79 -78 80 -77
rect 86 -78 87 -77
rect 93 -78 94 -77
rect 107 -78 108 -77
rect 110 -78 111 -77
rect 114 -78 115 -77
rect 149 -78 150 -77
rect 9 -80 10 -79
rect 19 -80 20 -79
rect 30 -80 31 -79
rect 89 -80 90 -79
rect 107 -80 108 -79
rect 135 -80 136 -79
rect 16 -82 17 -81
rect 23 -82 24 -81
rect 37 -82 38 -81
rect 58 -82 59 -81
rect 68 -82 69 -81
rect 79 -82 80 -81
rect 110 -82 111 -81
rect 135 -82 136 -81
rect 23 -84 24 -83
rect 54 -84 55 -83
rect 114 -84 115 -83
rect 124 -84 125 -83
rect 37 -86 38 -85
rect 61 -86 62 -85
rect 121 -86 122 -85
rect 131 -86 132 -85
rect 44 -88 45 -87
rect 65 -88 66 -87
rect 124 -88 125 -87
rect 128 -88 129 -87
rect 2 -99 3 -98
rect 16 -99 17 -98
rect 19 -99 20 -98
rect 58 -99 59 -98
rect 61 -99 62 -98
rect 152 -99 153 -98
rect 23 -101 24 -100
rect 51 -101 52 -100
rect 58 -101 59 -100
rect 82 -101 83 -100
rect 86 -101 87 -100
rect 114 -101 115 -100
rect 149 -101 150 -100
rect 156 -101 157 -100
rect 23 -103 24 -102
rect 37 -103 38 -102
rect 47 -103 48 -102
rect 142 -103 143 -102
rect 30 -105 31 -104
rect 65 -105 66 -104
rect 68 -105 69 -104
rect 107 -105 108 -104
rect 114 -105 115 -104
rect 131 -105 132 -104
rect 37 -107 38 -106
rect 44 -107 45 -106
rect 65 -107 66 -106
rect 121 -107 122 -106
rect 128 -107 129 -106
rect 142 -107 143 -106
rect 68 -109 69 -108
rect 149 -109 150 -108
rect 72 -111 73 -110
rect 89 -111 90 -110
rect 100 -111 101 -110
rect 103 -111 104 -110
rect 128 -111 129 -110
rect 163 -111 164 -110
rect 72 -113 73 -112
rect 100 -113 101 -112
rect 79 -115 80 -114
rect 107 -115 108 -114
rect 79 -117 80 -116
rect 135 -117 136 -116
rect 93 -119 94 -118
rect 135 -119 136 -118
rect 44 -121 45 -120
rect 93 -121 94 -120
rect 9 -132 10 -131
rect 47 -132 48 -131
rect 51 -132 52 -131
rect 79 -132 80 -131
rect 100 -132 101 -131
rect 135 -132 136 -131
rect 142 -132 143 -131
rect 184 -132 185 -131
rect 198 -132 199 -131
rect 205 -132 206 -131
rect 16 -134 17 -133
rect 44 -134 45 -133
rect 72 -134 73 -133
rect 82 -134 83 -133
rect 107 -134 108 -133
rect 128 -134 129 -133
rect 149 -134 150 -133
rect 191 -134 192 -133
rect 23 -136 24 -135
rect 65 -136 66 -135
rect 75 -136 76 -135
rect 79 -136 80 -135
rect 100 -136 101 -135
rect 107 -136 108 -135
rect 110 -136 111 -135
rect 177 -136 178 -135
rect 2 -138 3 -137
rect 65 -138 66 -137
rect 103 -138 104 -137
rect 128 -138 129 -137
rect 149 -138 150 -137
rect 163 -138 164 -137
rect 170 -138 171 -137
rect 201 -138 202 -137
rect 23 -140 24 -139
rect 58 -140 59 -139
rect 86 -140 87 -139
rect 170 -140 171 -139
rect 30 -142 31 -141
rect 37 -142 38 -141
rect 47 -142 48 -141
rect 86 -142 87 -141
rect 114 -142 115 -141
rect 135 -142 136 -141
rect 156 -142 157 -141
rect 173 -142 174 -141
rect 30 -144 31 -143
rect 40 -144 41 -143
rect 93 -144 94 -143
rect 114 -144 115 -143
rect 121 -144 122 -143
rect 163 -144 164 -143
rect 33 -146 34 -145
rect 142 -146 143 -145
rect 93 -148 94 -147
rect 156 -148 157 -147
rect 16 -159 17 -158
rect 47 -159 48 -158
rect 54 -159 55 -158
rect 163 -159 164 -158
rect 166 -159 167 -158
rect 177 -159 178 -158
rect 23 -161 24 -160
rect 65 -161 66 -160
rect 68 -161 69 -160
rect 79 -161 80 -160
rect 89 -161 90 -160
rect 100 -161 101 -160
rect 107 -161 108 -160
rect 114 -161 115 -160
rect 121 -161 122 -160
rect 156 -161 157 -160
rect 163 -161 164 -160
rect 201 -161 202 -160
rect 9 -163 10 -162
rect 79 -163 80 -162
rect 93 -163 94 -162
rect 135 -163 136 -162
rect 30 -165 31 -164
rect 44 -165 45 -164
rect 58 -165 59 -164
rect 96 -165 97 -164
rect 107 -165 108 -164
rect 114 -165 115 -164
rect 128 -165 129 -164
rect 135 -165 136 -164
rect 37 -167 38 -166
rect 149 -167 150 -166
rect 2 -169 3 -168
rect 37 -169 38 -168
rect 40 -169 41 -168
rect 72 -169 73 -168
rect 86 -169 87 -168
rect 128 -169 129 -168
rect 23 -171 24 -170
rect 86 -171 87 -170
rect 110 -171 111 -170
rect 184 -171 185 -170
rect 47 -173 48 -172
rect 58 -173 59 -172
rect 61 -173 62 -172
rect 191 -173 192 -172
rect 110 -175 111 -174
rect 142 -175 143 -174
rect 142 -177 143 -176
rect 170 -177 171 -176
rect 170 -179 171 -178
rect 205 -179 206 -178
rect 2 -190 3 -189
rect 23 -190 24 -189
rect 30 -190 31 -189
rect 82 -190 83 -189
rect 89 -190 90 -189
rect 128 -190 129 -189
rect 142 -190 143 -189
rect 170 -190 171 -189
rect 9 -192 10 -191
rect 37 -192 38 -191
rect 40 -192 41 -191
rect 79 -192 80 -191
rect 114 -192 115 -191
rect 121 -192 122 -191
rect 16 -194 17 -193
rect 54 -194 55 -193
rect 58 -194 59 -193
rect 107 -194 108 -193
rect 117 -194 118 -193
rect 159 -194 160 -193
rect 12 -196 13 -195
rect 58 -196 59 -195
rect 61 -196 62 -195
rect 149 -196 150 -195
rect 23 -198 24 -197
rect 47 -198 48 -197
rect 65 -198 66 -197
rect 100 -198 101 -197
rect 40 -200 41 -199
rect 86 -200 87 -199
rect 65 -202 66 -201
rect 72 -202 73 -201
rect 79 -202 80 -201
rect 93 -202 94 -201
rect 68 -204 69 -203
rect 142 -204 143 -203
rect 2 -215 3 -214
rect 44 -215 45 -214
rect 51 -215 52 -214
rect 107 -215 108 -214
rect 128 -215 129 -214
rect 135 -215 136 -214
rect 9 -217 10 -216
rect 68 -217 69 -216
rect 79 -217 80 -216
rect 121 -217 122 -216
rect 23 -219 24 -218
rect 58 -219 59 -218
rect 61 -219 62 -218
rect 100 -219 101 -218
rect 30 -221 31 -220
rect 47 -221 48 -220
rect 65 -221 66 -220
rect 86 -221 87 -220
rect 100 -221 101 -220
rect 149 -221 150 -220
rect 33 -223 34 -222
rect 54 -223 55 -222
rect 82 -223 83 -222
rect 114 -223 115 -222
rect 40 -225 41 -224
rect 93 -225 94 -224
rect 16 -227 17 -226
rect 40 -227 41 -226
rect 44 -227 45 -226
rect 68 -227 69 -226
rect 82 -227 83 -226
rect 142 -227 143 -226
rect 16 -229 17 -228
rect 26 -229 27 -228
rect 16 -240 17 -239
rect 30 -240 31 -239
rect 44 -240 45 -239
rect 79 -240 80 -239
rect 54 -242 55 -241
rect 82 -242 83 -241
rect 61 -244 62 -243
rect 72 -244 73 -243
rect 65 -246 66 -245
rect 86 -246 87 -245
<< metal2 >>
rect 44 -1 45 1
rect 58 -1 59 1
rect 65 -1 66 1
rect 79 -1 80 1
rect 37 -16 38 -10
rect 44 -11 45 -9
rect 51 -11 52 -9
rect 61 -16 62 -10
rect 65 -11 66 -9
rect 72 -16 73 -10
rect 79 -16 80 -10
rect 86 -16 87 -10
rect 93 -16 94 -10
rect 110 -16 111 -10
rect 30 -16 31 -12
rect 44 -16 45 -12
rect 51 -16 52 -12
rect 75 -13 76 -9
rect 58 -15 59 -9
rect 65 -16 66 -14
rect 16 -39 17 -25
rect 37 -26 38 -24
rect 44 -26 45 -24
rect 68 -39 69 -25
rect 89 -39 90 -25
rect 107 -39 108 -25
rect 114 -26 115 -24
rect 142 -39 143 -25
rect 9 -39 10 -27
rect 37 -39 38 -27
rect 47 -28 48 -24
rect 58 -28 59 -24
rect 61 -28 62 -24
rect 121 -39 122 -27
rect 26 -30 27 -24
rect 30 -30 31 -24
rect 44 -39 45 -29
rect 58 -39 59 -29
rect 65 -30 66 -24
rect 75 -39 76 -29
rect 93 -30 94 -24
rect 128 -39 129 -29
rect 23 -39 24 -31
rect 30 -39 31 -31
rect 72 -39 73 -31
rect 114 -39 115 -31
rect 79 -34 80 -24
rect 93 -39 94 -33
rect 100 -39 101 -33
rect 135 -39 136 -33
rect 79 -39 80 -35
rect 86 -36 87 -24
rect 51 -38 52 -24
rect 86 -39 87 -37
rect 9 -49 10 -47
rect 33 -66 34 -48
rect 37 -49 38 -47
rect 65 -49 66 -47
rect 68 -49 69 -47
rect 114 -49 115 -47
rect 131 -66 132 -48
rect 135 -49 136 -47
rect 23 -51 24 -47
rect 47 -51 48 -47
rect 51 -66 52 -50
rect 89 -66 90 -50
rect 103 -51 104 -47
rect 121 -51 122 -47
rect 9 -66 10 -52
rect 23 -66 24 -52
rect 30 -66 31 -52
rect 37 -66 38 -52
rect 58 -53 59 -47
rect 58 -66 59 -52
rect 58 -53 59 -47
rect 58 -66 59 -52
rect 68 -66 69 -52
rect 93 -53 94 -47
rect 107 -53 108 -47
rect 135 -66 136 -52
rect 16 -55 17 -47
rect 47 -66 48 -54
rect 54 -55 55 -47
rect 93 -66 94 -54
rect 16 -66 17 -56
rect 26 -66 27 -56
rect 65 -66 66 -56
rect 107 -66 108 -56
rect 72 -59 73 -47
rect 79 -59 80 -47
rect 86 -59 87 -47
rect 128 -59 129 -47
rect 72 -66 73 -60
rect 82 -66 83 -60
rect 86 -66 87 -60
rect 100 -66 101 -60
rect 75 -63 76 -47
rect 114 -66 115 -62
rect 79 -66 80 -64
rect 142 -65 143 -47
rect 2 -89 3 -75
rect 30 -76 31 -74
rect 47 -76 48 -74
rect 51 -76 52 -74
rect 58 -76 59 -74
rect 68 -76 69 -74
rect 72 -76 73 -74
rect 72 -89 73 -75
rect 72 -76 73 -74
rect 72 -89 73 -75
rect 89 -76 90 -74
rect 93 -76 94 -74
rect 100 -76 101 -74
rect 142 -89 143 -75
rect 9 -78 10 -74
rect 44 -78 45 -74
rect 51 -89 52 -77
rect 79 -78 80 -74
rect 86 -89 87 -77
rect 93 -89 94 -77
rect 107 -78 108 -74
rect 110 -82 111 -77
rect 114 -78 115 -74
rect 149 -89 150 -77
rect 9 -89 10 -79
rect 19 -89 20 -79
rect 30 -89 31 -79
rect 89 -89 90 -79
rect 107 -89 108 -79
rect 135 -80 136 -74
rect 16 -82 17 -74
rect 23 -82 24 -74
rect 37 -82 38 -74
rect 58 -89 59 -81
rect 68 -89 69 -81
rect 79 -89 80 -81
rect 135 -89 136 -81
rect 23 -89 24 -83
rect 54 -89 55 -83
rect 114 -89 115 -83
rect 124 -84 125 -74
rect 37 -89 38 -85
rect 61 -89 62 -85
rect 121 -89 122 -85
rect 131 -86 132 -74
rect 44 -89 45 -87
rect 65 -89 66 -87
rect 124 -89 125 -87
rect 128 -89 129 -87
rect 2 -99 3 -97
rect 16 -99 17 -97
rect 19 -122 20 -98
rect 58 -99 59 -97
rect 61 -99 62 -97
rect 152 -99 153 -97
rect 23 -101 24 -97
rect 51 -122 52 -100
rect 58 -122 59 -100
rect 82 -122 83 -100
rect 86 -101 87 -97
rect 114 -101 115 -97
rect 149 -101 150 -97
rect 156 -122 157 -100
rect 23 -122 24 -102
rect 37 -103 38 -97
rect 47 -122 48 -102
rect 142 -103 143 -97
rect 30 -105 31 -97
rect 65 -105 66 -97
rect 68 -105 69 -97
rect 107 -105 108 -97
rect 114 -122 115 -104
rect 131 -122 132 -104
rect 37 -122 38 -106
rect 44 -107 45 -97
rect 65 -122 66 -106
rect 121 -122 122 -106
rect 128 -107 129 -97
rect 142 -122 143 -106
rect 68 -122 69 -108
rect 149 -122 150 -108
rect 72 -111 73 -97
rect 89 -122 90 -110
rect 100 -111 101 -97
rect 103 -122 104 -110
rect 128 -122 129 -110
rect 163 -122 164 -110
rect 72 -122 73 -112
rect 100 -122 101 -112
rect 79 -115 80 -97
rect 107 -122 108 -114
rect 79 -122 80 -116
rect 135 -117 136 -97
rect 93 -119 94 -97
rect 135 -122 136 -118
rect 44 -122 45 -120
rect 93 -122 94 -120
rect 9 -149 10 -131
rect 47 -132 48 -130
rect 51 -132 52 -130
rect 79 -132 80 -130
rect 100 -132 101 -130
rect 135 -132 136 -130
rect 142 -132 143 -130
rect 184 -149 185 -131
rect 198 -149 199 -131
rect 205 -149 206 -131
rect 16 -149 17 -133
rect 44 -149 45 -133
rect 72 -134 73 -130
rect 82 -134 83 -130
rect 107 -134 108 -130
rect 128 -134 129 -130
rect 149 -134 150 -130
rect 191 -149 192 -133
rect 23 -136 24 -130
rect 65 -136 66 -130
rect 75 -149 76 -135
rect 79 -149 80 -135
rect 100 -149 101 -135
rect 107 -149 108 -135
rect 110 -149 111 -135
rect 177 -149 178 -135
rect 2 -149 3 -137
rect 65 -149 66 -137
rect 103 -138 104 -130
rect 128 -149 129 -137
rect 149 -149 150 -137
rect 163 -138 164 -130
rect 170 -138 171 -130
rect 201 -149 202 -137
rect 23 -149 24 -139
rect 58 -140 59 -130
rect 86 -140 87 -130
rect 170 -149 171 -139
rect 30 -142 31 -130
rect 37 -142 38 -130
rect 47 -149 48 -141
rect 86 -149 87 -141
rect 114 -142 115 -130
rect 135 -149 136 -141
rect 156 -142 157 -130
rect 173 -142 174 -130
rect 30 -149 31 -143
rect 40 -149 41 -143
rect 93 -144 94 -130
rect 114 -149 115 -143
rect 121 -144 122 -130
rect 163 -149 164 -143
rect 33 -146 34 -130
rect 142 -149 143 -145
rect 93 -149 94 -147
rect 156 -149 157 -147
rect 16 -159 17 -157
rect 47 -159 48 -157
rect 54 -159 55 -157
rect 163 -159 164 -157
rect 166 -180 167 -158
rect 177 -159 178 -157
rect 23 -161 24 -157
rect 65 -180 66 -160
rect 68 -161 69 -157
rect 79 -161 80 -157
rect 89 -180 90 -160
rect 100 -161 101 -157
rect 107 -161 108 -157
rect 114 -161 115 -157
rect 121 -161 122 -157
rect 156 -161 157 -157
rect 163 -180 164 -160
rect 201 -161 202 -157
rect 9 -163 10 -157
rect 79 -180 80 -162
rect 93 -163 94 -157
rect 135 -163 136 -157
rect 30 -165 31 -157
rect 44 -165 45 -157
rect 58 -165 59 -157
rect 96 -180 97 -164
rect 107 -180 108 -164
rect 114 -180 115 -164
rect 128 -165 129 -157
rect 135 -180 136 -164
rect 37 -167 38 -157
rect 149 -167 150 -157
rect 2 -169 3 -157
rect 37 -180 38 -168
rect 40 -169 41 -157
rect 72 -180 73 -168
rect 86 -169 87 -157
rect 128 -180 129 -168
rect 23 -180 24 -170
rect 86 -180 87 -170
rect 110 -171 111 -157
rect 184 -171 185 -157
rect 47 -180 48 -172
rect 58 -180 59 -172
rect 61 -173 62 -157
rect 191 -173 192 -157
rect 110 -180 111 -174
rect 142 -175 143 -157
rect 142 -180 143 -176
rect 170 -177 171 -157
rect 170 -180 171 -178
rect 205 -179 206 -157
rect 2 -205 3 -189
rect 23 -190 24 -188
rect 30 -205 31 -189
rect 82 -205 83 -189
rect 89 -190 90 -188
rect 128 -190 129 -188
rect 135 -190 136 -188
rect 135 -205 136 -189
rect 135 -190 136 -188
rect 135 -205 136 -189
rect 142 -190 143 -188
rect 170 -190 171 -188
rect 9 -205 10 -191
rect 37 -205 38 -191
rect 40 -192 41 -188
rect 79 -192 80 -188
rect 114 -192 115 -188
rect 121 -205 122 -191
rect 16 -205 17 -193
rect 54 -205 55 -193
rect 58 -194 59 -188
rect 107 -205 108 -193
rect 117 -205 118 -193
rect 159 -205 160 -193
rect 12 -196 13 -188
rect 58 -205 59 -195
rect 61 -205 62 -195
rect 149 -205 150 -195
rect 23 -205 24 -197
rect 47 -198 48 -188
rect 65 -198 66 -188
rect 100 -205 101 -197
rect 40 -205 41 -199
rect 86 -205 87 -199
rect 65 -205 66 -201
rect 72 -205 73 -201
rect 79 -205 80 -201
rect 93 -205 94 -201
rect 68 -205 69 -203
rect 142 -205 143 -203
rect 2 -215 3 -213
rect 44 -215 45 -213
rect 51 -215 52 -213
rect 107 -215 108 -213
rect 128 -215 129 -213
rect 135 -215 136 -213
rect 9 -217 10 -213
rect 68 -217 69 -213
rect 72 -217 73 -213
rect 72 -230 73 -216
rect 72 -217 73 -213
rect 72 -230 73 -216
rect 79 -217 80 -213
rect 121 -217 122 -213
rect 23 -219 24 -213
rect 58 -219 59 -213
rect 61 -230 62 -218
rect 100 -219 101 -213
rect 30 -221 31 -213
rect 47 -221 48 -213
rect 65 -221 66 -213
rect 86 -221 87 -213
rect 100 -230 101 -220
rect 149 -221 150 -213
rect 33 -230 34 -222
rect 54 -230 55 -222
rect 82 -223 83 -213
rect 114 -223 115 -213
rect 40 -225 41 -213
rect 93 -225 94 -213
rect 16 -227 17 -213
rect 40 -230 41 -226
rect 44 -230 45 -226
rect 68 -230 69 -226
rect 82 -230 83 -226
rect 142 -227 143 -213
rect 16 -230 17 -228
rect 26 -230 27 -228
rect 16 -240 17 -238
rect 30 -240 31 -238
rect 44 -240 45 -238
rect 79 -240 80 -238
rect 54 -242 55 -238
rect 82 -242 83 -238
rect 61 -244 62 -238
rect 72 -244 73 -238
rect 65 -246 66 -238
rect 86 -246 87 -238
<< labels >>
rlabel pdiffusion 3 -6 3 -6 0 cellNo=1
rlabel pdiffusion 10 -6 10 -6 0 cellNo=55
rlabel pdiffusion 17 -6 17 -6 0 cellNo=32
rlabel pdiffusion 45 -6 45 -6 0 feedthrough
rlabel pdiffusion 52 -6 52 -6 0 cellNo=23
rlabel pdiffusion 59 -6 59 -6 0 cellNo=85
rlabel pdiffusion 66 -6 66 -6 0 feedthrough
rlabel pdiffusion 73 -6 73 -6 0 cellNo=9
rlabel pdiffusion 80 -6 80 -6 0 cellNo=10
rlabel pdiffusion 3 -21 3 -21 0 cellNo=19
rlabel pdiffusion 17 -21 17 -21 0 cellNo=67
rlabel pdiffusion 24 -21 24 -21 0 cellNo=81
rlabel pdiffusion 31 -21 31 -21 0 feedthrough
rlabel pdiffusion 38 -21 38 -21 0 feedthrough
rlabel pdiffusion 45 -21 45 -21 0 cellNo=77
rlabel pdiffusion 52 -21 52 -21 0 feedthrough
rlabel pdiffusion 59 -21 59 -21 0 cellNo=16
rlabel pdiffusion 66 -21 66 -21 0 feedthrough
rlabel pdiffusion 73 -21 73 -21 0 cellNo=15
rlabel pdiffusion 80 -21 80 -21 0 feedthrough
rlabel pdiffusion 87 -21 87 -21 0 cellNo=4
rlabel pdiffusion 94 -21 94 -21 0 feedthrough
rlabel pdiffusion 108 -21 108 -21 0 cellNo=21
rlabel pdiffusion 115 -21 115 -21 0 cellNo=64
rlabel pdiffusion 3 -44 3 -44 0 cellNo=18
rlabel pdiffusion 10 -44 10 -44 0 feedthrough
rlabel pdiffusion 17 -44 17 -44 0 feedthrough
rlabel pdiffusion 24 -44 24 -44 0 feedthrough
rlabel pdiffusion 31 -44 31 -44 0 cellNo=35
rlabel pdiffusion 38 -44 38 -44 0 cellNo=33
rlabel pdiffusion 45 -44 45 -44 0 cellNo=58
rlabel pdiffusion 52 -44 52 -44 0 cellNo=3
rlabel pdiffusion 59 -44 59 -44 0 feedthrough
rlabel pdiffusion 66 -44 66 -44 0 cellNo=34
rlabel pdiffusion 73 -44 73 -44 0 cellNo=53
rlabel pdiffusion 80 -44 80 -44 0 feedthrough
rlabel pdiffusion 87 -44 87 -44 0 cellNo=43
rlabel pdiffusion 94 -44 94 -44 0 feedthrough
rlabel pdiffusion 101 -44 101 -44 0 cellNo=79
rlabel pdiffusion 108 -44 108 -44 0 feedthrough
rlabel pdiffusion 115 -44 115 -44 0 feedthrough
rlabel pdiffusion 122 -44 122 -44 0 feedthrough
rlabel pdiffusion 129 -44 129 -44 0 feedthrough
rlabel pdiffusion 136 -44 136 -44 0 feedthrough
rlabel pdiffusion 143 -44 143 -44 0 feedthrough
rlabel pdiffusion 3 -71 3 -71 0 cellNo=57
rlabel pdiffusion 10 -71 10 -71 0 feedthrough
rlabel pdiffusion 17 -71 17 -71 0 feedthrough
rlabel pdiffusion 24 -71 24 -71 0 cellNo=22
rlabel pdiffusion 31 -71 31 -71 0 cellNo=46
rlabel pdiffusion 38 -71 38 -71 0 feedthrough
rlabel pdiffusion 45 -71 45 -71 0 cellNo=31
rlabel pdiffusion 52 -71 52 -71 0 feedthrough
rlabel pdiffusion 59 -71 59 -71 0 feedthrough
rlabel pdiffusion 66 -71 66 -71 0 cellNo=7
rlabel pdiffusion 73 -71 73 -71 0 feedthrough
rlabel pdiffusion 80 -71 80 -71 0 cellNo=65
rlabel pdiffusion 87 -71 87 -71 0 cellNo=28
rlabel pdiffusion 94 -71 94 -71 0 feedthrough
rlabel pdiffusion 101 -71 101 -71 0 feedthrough
rlabel pdiffusion 108 -71 108 -71 0 feedthrough
rlabel pdiffusion 115 -71 115 -71 0 feedthrough
rlabel pdiffusion 122 -71 122 -71 0 cellNo=56
rlabel pdiffusion 129 -71 129 -71 0 cellNo=25
rlabel pdiffusion 136 -71 136 -71 0 feedthrough
rlabel pdiffusion 3 -94 3 -94 0 feedthrough
rlabel pdiffusion 10 -94 10 -94 0 cellNo=47
rlabel pdiffusion 17 -94 17 -94 0 cellNo=14
rlabel pdiffusion 24 -94 24 -94 0 feedthrough
rlabel pdiffusion 31 -94 31 -94 0 feedthrough
rlabel pdiffusion 38 -94 38 -94 0 feedthrough
rlabel pdiffusion 45 -94 45 -94 0 feedthrough
rlabel pdiffusion 52 -94 52 -94 0 cellNo=26
rlabel pdiffusion 59 -94 59 -94 0 cellNo=38
rlabel pdiffusion 66 -94 66 -94 0 cellNo=68
rlabel pdiffusion 73 -94 73 -94 0 feedthrough
rlabel pdiffusion 80 -94 80 -94 0 feedthrough
rlabel pdiffusion 87 -94 87 -94 0 cellNo=36
rlabel pdiffusion 94 -94 94 -94 0 feedthrough
rlabel pdiffusion 101 -94 101 -94 0 cellNo=13
rlabel pdiffusion 108 -94 108 -94 0 feedthrough
rlabel pdiffusion 115 -94 115 -94 0 feedthrough
rlabel pdiffusion 122 -94 122 -94 0 cellNo=29
rlabel pdiffusion 129 -94 129 -94 0 feedthrough
rlabel pdiffusion 136 -94 136 -94 0 feedthrough
rlabel pdiffusion 143 -94 143 -94 0 feedthrough
rlabel pdiffusion 150 -94 150 -94 0 cellNo=54
rlabel pdiffusion 17 -127 17 -127 0 cellNo=74
rlabel pdiffusion 24 -127 24 -127 0 feedthrough
rlabel pdiffusion 31 -127 31 -127 0 cellNo=2
rlabel pdiffusion 38 -127 38 -127 0 feedthrough
rlabel pdiffusion 45 -127 45 -127 0 cellNo=59
rlabel pdiffusion 52 -127 52 -127 0 feedthrough
rlabel pdiffusion 59 -127 59 -127 0 feedthrough
rlabel pdiffusion 66 -127 66 -127 0 cellNo=80
rlabel pdiffusion 73 -127 73 -127 0 feedthrough
rlabel pdiffusion 80 -127 80 -127 0 cellNo=84
rlabel pdiffusion 87 -127 87 -127 0 cellNo=82
rlabel pdiffusion 94 -127 94 -127 0 feedthrough
rlabel pdiffusion 101 -127 101 -127 0 cellNo=44
rlabel pdiffusion 108 -127 108 -127 0 feedthrough
rlabel pdiffusion 115 -127 115 -127 0 feedthrough
rlabel pdiffusion 122 -127 122 -127 0 feedthrough
rlabel pdiffusion 129 -127 129 -127 0 cellNo=11
rlabel pdiffusion 136 -127 136 -127 0 feedthrough
rlabel pdiffusion 143 -127 143 -127 0 feedthrough
rlabel pdiffusion 150 -127 150 -127 0 feedthrough
rlabel pdiffusion 157 -127 157 -127 0 feedthrough
rlabel pdiffusion 164 -127 164 -127 0 feedthrough
rlabel pdiffusion 171 -127 171 -127 0 cellNo=39
rlabel pdiffusion 3 -154 3 -154 0 feedthrough
rlabel pdiffusion 10 -154 10 -154 0 feedthrough
rlabel pdiffusion 17 -154 17 -154 0 feedthrough
rlabel pdiffusion 24 -154 24 -154 0 feedthrough
rlabel pdiffusion 31 -154 31 -154 0 feedthrough
rlabel pdiffusion 38 -154 38 -154 0 cellNo=37
rlabel pdiffusion 45 -154 45 -154 0 cellNo=48
rlabel pdiffusion 52 -154 52 -154 0 cellNo=41
rlabel pdiffusion 59 -154 59 -154 0 cellNo=30
rlabel pdiffusion 66 -154 66 -154 0 cellNo=27
rlabel pdiffusion 73 -154 73 -154 0 cellNo=50
rlabel pdiffusion 80 -154 80 -154 0 feedthrough
rlabel pdiffusion 87 -154 87 -154 0 feedthrough
rlabel pdiffusion 94 -154 94 -154 0 cellNo=24
rlabel pdiffusion 101 -154 101 -154 0 feedthrough
rlabel pdiffusion 108 -154 108 -154 0 cellNo=87
rlabel pdiffusion 115 -154 115 -154 0 feedthrough
rlabel pdiffusion 122 -154 122 -154 0 cellNo=6
rlabel pdiffusion 129 -154 129 -154 0 feedthrough
rlabel pdiffusion 136 -154 136 -154 0 feedthrough
rlabel pdiffusion 143 -154 143 -154 0 feedthrough
rlabel pdiffusion 150 -154 150 -154 0 feedthrough
rlabel pdiffusion 157 -154 157 -154 0 feedthrough
rlabel pdiffusion 164 -154 164 -154 0 feedthrough
rlabel pdiffusion 171 -154 171 -154 0 feedthrough
rlabel pdiffusion 178 -154 178 -154 0 feedthrough
rlabel pdiffusion 185 -154 185 -154 0 feedthrough
rlabel pdiffusion 192 -154 192 -154 0 feedthrough
rlabel pdiffusion 199 -154 199 -154 0 cellNo=90
rlabel pdiffusion 206 -154 206 -154 0 feedthrough
rlabel pdiffusion 10 -185 10 -185 0 cellNo=51
rlabel pdiffusion 24 -185 24 -185 0 feedthrough
rlabel pdiffusion 38 -185 38 -185 0 cellNo=60
rlabel pdiffusion 45 -185 45 -185 0 cellNo=61
rlabel pdiffusion 59 -185 59 -185 0 feedthrough
rlabel pdiffusion 66 -185 66 -185 0 cellNo=40
rlabel pdiffusion 73 -185 73 -185 0 cellNo=70
rlabel pdiffusion 80 -185 80 -185 0 feedthrough
rlabel pdiffusion 87 -185 87 -185 0 cellNo=69
rlabel pdiffusion 94 -185 94 -185 0 cellNo=12
rlabel pdiffusion 108 -185 108 -185 0 cellNo=52
rlabel pdiffusion 115 -185 115 -185 0 feedthrough
rlabel pdiffusion 129 -185 129 -185 0 feedthrough
rlabel pdiffusion 136 -185 136 -185 0 feedthrough
rlabel pdiffusion 143 -185 143 -185 0 cellNo=78
rlabel pdiffusion 164 -185 164 -185 0 cellNo=42
rlabel pdiffusion 171 -185 171 -185 0 feedthrough
rlabel pdiffusion 3 -210 3 -210 0 feedthrough
rlabel pdiffusion 10 -210 10 -210 0 feedthrough
rlabel pdiffusion 17 -210 17 -210 0 feedthrough
rlabel pdiffusion 24 -210 24 -210 0 feedthrough
rlabel pdiffusion 31 -210 31 -210 0 feedthrough
rlabel pdiffusion 38 -210 38 -210 0 cellNo=89
rlabel pdiffusion 45 -210 45 -210 0 cellNo=83
rlabel pdiffusion 52 -210 52 -210 0 cellNo=49
rlabel pdiffusion 59 -210 59 -210 0 cellNo=17
rlabel pdiffusion 66 -210 66 -210 0 cellNo=5
rlabel pdiffusion 73 -210 73 -210 0 feedthrough
rlabel pdiffusion 80 -210 80 -210 0 cellNo=76
rlabel pdiffusion 87 -210 87 -210 0 feedthrough
rlabel pdiffusion 94 -210 94 -210 0 feedthrough
rlabel pdiffusion 101 -210 101 -210 0 feedthrough
rlabel pdiffusion 108 -210 108 -210 0 feedthrough
rlabel pdiffusion 115 -210 115 -210 0 cellNo=8
rlabel pdiffusion 122 -210 122 -210 0 feedthrough
rlabel pdiffusion 129 -210 129 -210 0 cellNo=72
rlabel pdiffusion 136 -210 136 -210 0 feedthrough
rlabel pdiffusion 143 -210 143 -210 0 feedthrough
rlabel pdiffusion 150 -210 150 -210 0 feedthrough
rlabel pdiffusion 157 -210 157 -210 0 cellNo=66
rlabel pdiffusion 17 -235 17 -235 0 feedthrough
rlabel pdiffusion 24 -235 24 -235 0 cellNo=88
rlabel pdiffusion 31 -235 31 -235 0 cellNo=45
rlabel pdiffusion 38 -235 38 -235 0 cellNo=63
rlabel pdiffusion 45 -235 45 -235 0 feedthrough
rlabel pdiffusion 52 -235 52 -235 0 cellNo=73
rlabel pdiffusion 59 -235 59 -235 0 cellNo=86
rlabel pdiffusion 66 -235 66 -235 0 cellNo=75
rlabel pdiffusion 73 -235 73 -235 0 feedthrough
rlabel pdiffusion 80 -235 80 -235 0 cellNo=62
rlabel pdiffusion 87 -235 87 -235 0 cellNo=71
rlabel pdiffusion 101 -235 101 -235 0 cellNo=20
rlabel polysilicon 44 -2 44 -2 0 1
rlabel polysilicon 44 -8 44 -8 0 3
rlabel polysilicon 51 -8 51 -8 0 3
rlabel polysilicon 58 -2 58 -2 0 1
rlabel polysilicon 58 -8 58 -8 0 3
rlabel polysilicon 65 -2 65 -2 0 1
rlabel polysilicon 65 -8 65 -8 0 3
rlabel polysilicon 75 -8 75 -8 0 4
rlabel polysilicon 79 -2 79 -2 0 1
rlabel polysilicon 26 -23 26 -23 0 4
rlabel polysilicon 30 -17 30 -17 0 1
rlabel polysilicon 30 -23 30 -23 0 3
rlabel polysilicon 37 -17 37 -17 0 1
rlabel polysilicon 37 -23 37 -23 0 3
rlabel polysilicon 44 -17 44 -17 0 1
rlabel polysilicon 44 -23 44 -23 0 3
rlabel polysilicon 47 -23 47 -23 0 4
rlabel polysilicon 51 -17 51 -17 0 1
rlabel polysilicon 51 -23 51 -23 0 3
rlabel polysilicon 61 -17 61 -17 0 2
rlabel polysilicon 58 -23 58 -23 0 3
rlabel polysilicon 61 -23 61 -23 0 4
rlabel polysilicon 65 -17 65 -17 0 1
rlabel polysilicon 65 -23 65 -23 0 3
rlabel polysilicon 72 -17 72 -17 0 1
rlabel polysilicon 79 -17 79 -17 0 1
rlabel polysilicon 79 -23 79 -23 0 3
rlabel polysilicon 86 -17 86 -17 0 1
rlabel polysilicon 86 -23 86 -23 0 3
rlabel polysilicon 93 -17 93 -17 0 1
rlabel polysilicon 93 -23 93 -23 0 3
rlabel polysilicon 110 -17 110 -17 0 2
rlabel polysilicon 114 -23 114 -23 0 3
rlabel polysilicon 9 -40 9 -40 0 1
rlabel polysilicon 9 -46 9 -46 0 3
rlabel polysilicon 16 -40 16 -40 0 1
rlabel polysilicon 16 -46 16 -46 0 3
rlabel polysilicon 23 -40 23 -40 0 1
rlabel polysilicon 23 -46 23 -46 0 3
rlabel polysilicon 30 -40 30 -40 0 1
rlabel polysilicon 37 -40 37 -40 0 1
rlabel polysilicon 37 -46 37 -46 0 3
rlabel polysilicon 44 -40 44 -40 0 1
rlabel polysilicon 47 -46 47 -46 0 4
rlabel polysilicon 54 -46 54 -46 0 4
rlabel polysilicon 58 -40 58 -40 0 1
rlabel polysilicon 58 -46 58 -46 0 3
rlabel polysilicon 68 -40 68 -40 0 2
rlabel polysilicon 65 -46 65 -46 0 3
rlabel polysilicon 68 -46 68 -46 0 4
rlabel polysilicon 72 -40 72 -40 0 1
rlabel polysilicon 75 -40 75 -40 0 2
rlabel polysilicon 72 -46 72 -46 0 3
rlabel polysilicon 75 -46 75 -46 0 4
rlabel polysilicon 79 -40 79 -40 0 1
rlabel polysilicon 79 -46 79 -46 0 3
rlabel polysilicon 86 -40 86 -40 0 1
rlabel polysilicon 89 -40 89 -40 0 2
rlabel polysilicon 86 -46 86 -46 0 3
rlabel polysilicon 93 -40 93 -40 0 1
rlabel polysilicon 93 -46 93 -46 0 3
rlabel polysilicon 100 -40 100 -40 0 1
rlabel polysilicon 103 -46 103 -46 0 4
rlabel polysilicon 107 -40 107 -40 0 1
rlabel polysilicon 107 -46 107 -46 0 3
rlabel polysilicon 114 -40 114 -40 0 1
rlabel polysilicon 114 -46 114 -46 0 3
rlabel polysilicon 121 -40 121 -40 0 1
rlabel polysilicon 121 -46 121 -46 0 3
rlabel polysilicon 128 -40 128 -40 0 1
rlabel polysilicon 128 -46 128 -46 0 3
rlabel polysilicon 135 -40 135 -40 0 1
rlabel polysilicon 135 -46 135 -46 0 3
rlabel polysilicon 142 -40 142 -40 0 1
rlabel polysilicon 142 -46 142 -46 0 3
rlabel polysilicon 9 -67 9 -67 0 1
rlabel polysilicon 9 -73 9 -73 0 3
rlabel polysilicon 16 -67 16 -67 0 1
rlabel polysilicon 16 -73 16 -73 0 3
rlabel polysilicon 23 -67 23 -67 0 1
rlabel polysilicon 26 -67 26 -67 0 2
rlabel polysilicon 23 -73 23 -73 0 3
rlabel polysilicon 30 -67 30 -67 0 1
rlabel polysilicon 33 -67 33 -67 0 2
rlabel polysilicon 30 -73 30 -73 0 3
rlabel polysilicon 37 -67 37 -67 0 1
rlabel polysilicon 37 -73 37 -73 0 3
rlabel polysilicon 47 -67 47 -67 0 2
rlabel polysilicon 44 -73 44 -73 0 3
rlabel polysilicon 47 -73 47 -73 0 4
rlabel polysilicon 51 -67 51 -67 0 1
rlabel polysilicon 51 -73 51 -73 0 3
rlabel polysilicon 58 -67 58 -67 0 1
rlabel polysilicon 58 -73 58 -73 0 3
rlabel polysilicon 65 -67 65 -67 0 1
rlabel polysilicon 68 -67 68 -67 0 2
rlabel polysilicon 68 -73 68 -73 0 4
rlabel polysilicon 72 -67 72 -67 0 1
rlabel polysilicon 72 -73 72 -73 0 3
rlabel polysilicon 79 -67 79 -67 0 1
rlabel polysilicon 82 -67 82 -67 0 2
rlabel polysilicon 79 -73 79 -73 0 3
rlabel polysilicon 86 -67 86 -67 0 1
rlabel polysilicon 89 -67 89 -67 0 2
rlabel polysilicon 89 -73 89 -73 0 4
rlabel polysilicon 93 -67 93 -67 0 1
rlabel polysilicon 93 -73 93 -73 0 3
rlabel polysilicon 100 -67 100 -67 0 1
rlabel polysilicon 100 -73 100 -73 0 3
rlabel polysilicon 107 -67 107 -67 0 1
rlabel polysilicon 107 -73 107 -73 0 3
rlabel polysilicon 114 -67 114 -67 0 1
rlabel polysilicon 114 -73 114 -73 0 3
rlabel polysilicon 124 -73 124 -73 0 4
rlabel polysilicon 131 -67 131 -67 0 2
rlabel polysilicon 131 -73 131 -73 0 4
rlabel polysilicon 135 -67 135 -67 0 1
rlabel polysilicon 135 -73 135 -73 0 3
rlabel polysilicon 2 -90 2 -90 0 1
rlabel polysilicon 2 -96 2 -96 0 3
rlabel polysilicon 9 -90 9 -90 0 1
rlabel polysilicon 19 -90 19 -90 0 2
rlabel polysilicon 16 -96 16 -96 0 3
rlabel polysilicon 23 -90 23 -90 0 1
rlabel polysilicon 23 -96 23 -96 0 3
rlabel polysilicon 30 -90 30 -90 0 1
rlabel polysilicon 30 -96 30 -96 0 3
rlabel polysilicon 37 -90 37 -90 0 1
rlabel polysilicon 37 -96 37 -96 0 3
rlabel polysilicon 44 -90 44 -90 0 1
rlabel polysilicon 44 -96 44 -96 0 3
rlabel polysilicon 51 -90 51 -90 0 1
rlabel polysilicon 54 -90 54 -90 0 2
rlabel polysilicon 58 -90 58 -90 0 1
rlabel polysilicon 61 -90 61 -90 0 2
rlabel polysilicon 58 -96 58 -96 0 3
rlabel polysilicon 61 -96 61 -96 0 4
rlabel polysilicon 65 -90 65 -90 0 1
rlabel polysilicon 68 -90 68 -90 0 2
rlabel polysilicon 65 -96 65 -96 0 3
rlabel polysilicon 68 -96 68 -96 0 4
rlabel polysilicon 72 -90 72 -90 0 1
rlabel polysilicon 72 -96 72 -96 0 3
rlabel polysilicon 79 -90 79 -90 0 1
rlabel polysilicon 79 -96 79 -96 0 3
rlabel polysilicon 86 -90 86 -90 0 1
rlabel polysilicon 89 -90 89 -90 0 2
rlabel polysilicon 86 -96 86 -96 0 3
rlabel polysilicon 93 -90 93 -90 0 1
rlabel polysilicon 93 -96 93 -96 0 3
rlabel polysilicon 100 -96 100 -96 0 3
rlabel polysilicon 107 -90 107 -90 0 1
rlabel polysilicon 107 -96 107 -96 0 3
rlabel polysilicon 114 -90 114 -90 0 1
rlabel polysilicon 114 -96 114 -96 0 3
rlabel polysilicon 121 -90 121 -90 0 1
rlabel polysilicon 124 -90 124 -90 0 2
rlabel polysilicon 128 -90 128 -90 0 1
rlabel polysilicon 128 -96 128 -96 0 3
rlabel polysilicon 135 -90 135 -90 0 1
rlabel polysilicon 135 -96 135 -96 0 3
rlabel polysilicon 142 -90 142 -90 0 1
rlabel polysilicon 142 -96 142 -96 0 3
rlabel polysilicon 149 -90 149 -90 0 1
rlabel polysilicon 149 -96 149 -96 0 3
rlabel polysilicon 152 -96 152 -96 0 4
rlabel polysilicon 19 -123 19 -123 0 2
rlabel polysilicon 23 -123 23 -123 0 1
rlabel polysilicon 23 -129 23 -129 0 3
rlabel polysilicon 30 -129 30 -129 0 3
rlabel polysilicon 33 -129 33 -129 0 4
rlabel polysilicon 37 -123 37 -123 0 1
rlabel polysilicon 37 -129 37 -129 0 3
rlabel polysilicon 44 -123 44 -123 0 1
rlabel polysilicon 47 -123 47 -123 0 2
rlabel polysilicon 47 -129 47 -129 0 4
rlabel polysilicon 51 -123 51 -123 0 1
rlabel polysilicon 51 -129 51 -129 0 3
rlabel polysilicon 58 -123 58 -123 0 1
rlabel polysilicon 58 -129 58 -129 0 3
rlabel polysilicon 65 -123 65 -123 0 1
rlabel polysilicon 68 -123 68 -123 0 2
rlabel polysilicon 65 -129 65 -129 0 3
rlabel polysilicon 72 -123 72 -123 0 1
rlabel polysilicon 72 -129 72 -129 0 3
rlabel polysilicon 79 -123 79 -123 0 1
rlabel polysilicon 82 -123 82 -123 0 2
rlabel polysilicon 79 -129 79 -129 0 3
rlabel polysilicon 82 -129 82 -129 0 4
rlabel polysilicon 89 -123 89 -123 0 2
rlabel polysilicon 86 -129 86 -129 0 3
rlabel polysilicon 93 -123 93 -123 0 1
rlabel polysilicon 93 -129 93 -129 0 3
rlabel polysilicon 100 -123 100 -123 0 1
rlabel polysilicon 103 -123 103 -123 0 2
rlabel polysilicon 100 -129 100 -129 0 3
rlabel polysilicon 103 -129 103 -129 0 4
rlabel polysilicon 107 -123 107 -123 0 1
rlabel polysilicon 107 -129 107 -129 0 3
rlabel polysilicon 114 -123 114 -123 0 1
rlabel polysilicon 114 -129 114 -129 0 3
rlabel polysilicon 121 -123 121 -123 0 1
rlabel polysilicon 121 -129 121 -129 0 3
rlabel polysilicon 128 -123 128 -123 0 1
rlabel polysilicon 131 -123 131 -123 0 2
rlabel polysilicon 128 -129 128 -129 0 3
rlabel polysilicon 135 -123 135 -123 0 1
rlabel polysilicon 135 -129 135 -129 0 3
rlabel polysilicon 142 -123 142 -123 0 1
rlabel polysilicon 142 -129 142 -129 0 3
rlabel polysilicon 149 -123 149 -123 0 1
rlabel polysilicon 149 -129 149 -129 0 3
rlabel polysilicon 156 -123 156 -123 0 1
rlabel polysilicon 156 -129 156 -129 0 3
rlabel polysilicon 163 -123 163 -123 0 1
rlabel polysilicon 163 -129 163 -129 0 3
rlabel polysilicon 170 -129 170 -129 0 3
rlabel polysilicon 173 -129 173 -129 0 4
rlabel polysilicon 2 -150 2 -150 0 1
rlabel polysilicon 2 -156 2 -156 0 3
rlabel polysilicon 9 -150 9 -150 0 1
rlabel polysilicon 9 -156 9 -156 0 3
rlabel polysilicon 16 -150 16 -150 0 1
rlabel polysilicon 16 -156 16 -156 0 3
rlabel polysilicon 23 -150 23 -150 0 1
rlabel polysilicon 23 -156 23 -156 0 3
rlabel polysilicon 30 -150 30 -150 0 1
rlabel polysilicon 30 -156 30 -156 0 3
rlabel polysilicon 40 -150 40 -150 0 2
rlabel polysilicon 37 -156 37 -156 0 3
rlabel polysilicon 40 -156 40 -156 0 4
rlabel polysilicon 44 -150 44 -150 0 1
rlabel polysilicon 47 -150 47 -150 0 2
rlabel polysilicon 44 -156 44 -156 0 3
rlabel polysilicon 47 -156 47 -156 0 4
rlabel polysilicon 54 -156 54 -156 0 4
rlabel polysilicon 58 -156 58 -156 0 3
rlabel polysilicon 61 -156 61 -156 0 4
rlabel polysilicon 65 -150 65 -150 0 1
rlabel polysilicon 68 -156 68 -156 0 4
rlabel polysilicon 75 -150 75 -150 0 2
rlabel polysilicon 79 -150 79 -150 0 1
rlabel polysilicon 79 -156 79 -156 0 3
rlabel polysilicon 86 -150 86 -150 0 1
rlabel polysilicon 86 -156 86 -156 0 3
rlabel polysilicon 93 -150 93 -150 0 1
rlabel polysilicon 93 -156 93 -156 0 3
rlabel polysilicon 100 -150 100 -150 0 1
rlabel polysilicon 100 -156 100 -156 0 3
rlabel polysilicon 107 -150 107 -150 0 1
rlabel polysilicon 110 -150 110 -150 0 2
rlabel polysilicon 107 -156 107 -156 0 3
rlabel polysilicon 110 -156 110 -156 0 4
rlabel polysilicon 114 -150 114 -150 0 1
rlabel polysilicon 114 -156 114 -156 0 3
rlabel polysilicon 121 -156 121 -156 0 3
rlabel polysilicon 128 -150 128 -150 0 1
rlabel polysilicon 128 -156 128 -156 0 3
rlabel polysilicon 135 -150 135 -150 0 1
rlabel polysilicon 135 -156 135 -156 0 3
rlabel polysilicon 142 -150 142 -150 0 1
rlabel polysilicon 142 -156 142 -156 0 3
rlabel polysilicon 149 -150 149 -150 0 1
rlabel polysilicon 149 -156 149 -156 0 3
rlabel polysilicon 156 -150 156 -150 0 1
rlabel polysilicon 156 -156 156 -156 0 3
rlabel polysilicon 163 -150 163 -150 0 1
rlabel polysilicon 163 -156 163 -156 0 3
rlabel polysilicon 170 -150 170 -150 0 1
rlabel polysilicon 170 -156 170 -156 0 3
rlabel polysilicon 177 -150 177 -150 0 1
rlabel polysilicon 177 -156 177 -156 0 3
rlabel polysilicon 184 -150 184 -150 0 1
rlabel polysilicon 184 -156 184 -156 0 3
rlabel polysilicon 191 -150 191 -150 0 1
rlabel polysilicon 191 -156 191 -156 0 3
rlabel polysilicon 198 -150 198 -150 0 1
rlabel polysilicon 201 -150 201 -150 0 2
rlabel polysilicon 201 -156 201 -156 0 4
rlabel polysilicon 205 -150 205 -150 0 1
rlabel polysilicon 205 -156 205 -156 0 3
rlabel polysilicon 12 -187 12 -187 0 4
rlabel polysilicon 23 -181 23 -181 0 1
rlabel polysilicon 23 -187 23 -187 0 3
rlabel polysilicon 37 -181 37 -181 0 1
rlabel polysilicon 40 -187 40 -187 0 4
rlabel polysilicon 47 -181 47 -181 0 2
rlabel polysilicon 47 -187 47 -187 0 4
rlabel polysilicon 58 -181 58 -181 0 1
rlabel polysilicon 58 -187 58 -187 0 3
rlabel polysilicon 65 -181 65 -181 0 1
rlabel polysilicon 65 -187 65 -187 0 3
rlabel polysilicon 72 -181 72 -181 0 1
rlabel polysilicon 79 -181 79 -181 0 1
rlabel polysilicon 79 -187 79 -187 0 3
rlabel polysilicon 86 -181 86 -181 0 1
rlabel polysilicon 89 -181 89 -181 0 2
rlabel polysilicon 89 -187 89 -187 0 4
rlabel polysilicon 96 -181 96 -181 0 2
rlabel polysilicon 107 -181 107 -181 0 1
rlabel polysilicon 110 -181 110 -181 0 2
rlabel polysilicon 114 -181 114 -181 0 1
rlabel polysilicon 114 -187 114 -187 0 3
rlabel polysilicon 128 -181 128 -181 0 1
rlabel polysilicon 128 -187 128 -187 0 3
rlabel polysilicon 135 -181 135 -181 0 1
rlabel polysilicon 135 -187 135 -187 0 3
rlabel polysilicon 142 -181 142 -181 0 1
rlabel polysilicon 142 -187 142 -187 0 3
rlabel polysilicon 163 -181 163 -181 0 1
rlabel polysilicon 166 -181 166 -181 0 2
rlabel polysilicon 170 -181 170 -181 0 1
rlabel polysilicon 170 -187 170 -187 0 3
rlabel polysilicon 2 -206 2 -206 0 1
rlabel polysilicon 2 -212 2 -212 0 3
rlabel polysilicon 9 -206 9 -206 0 1
rlabel polysilicon 9 -212 9 -212 0 3
rlabel polysilicon 16 -206 16 -206 0 1
rlabel polysilicon 16 -212 16 -212 0 3
rlabel polysilicon 23 -206 23 -206 0 1
rlabel polysilicon 23 -212 23 -212 0 3
rlabel polysilicon 30 -206 30 -206 0 1
rlabel polysilicon 30 -212 30 -212 0 3
rlabel polysilicon 37 -206 37 -206 0 1
rlabel polysilicon 40 -206 40 -206 0 2
rlabel polysilicon 40 -212 40 -212 0 4
rlabel polysilicon 44 -212 44 -212 0 3
rlabel polysilicon 47 -212 47 -212 0 4
rlabel polysilicon 54 -206 54 -206 0 2
rlabel polysilicon 51 -212 51 -212 0 3
rlabel polysilicon 58 -206 58 -206 0 1
rlabel polysilicon 61 -206 61 -206 0 2
rlabel polysilicon 58 -212 58 -212 0 3
rlabel polysilicon 65 -206 65 -206 0 1
rlabel polysilicon 68 -206 68 -206 0 2
rlabel polysilicon 65 -212 65 -212 0 3
rlabel polysilicon 68 -212 68 -212 0 4
rlabel polysilicon 72 -206 72 -206 0 1
rlabel polysilicon 72 -212 72 -212 0 3
rlabel polysilicon 79 -206 79 -206 0 1
rlabel polysilicon 82 -206 82 -206 0 2
rlabel polysilicon 79 -212 79 -212 0 3
rlabel polysilicon 82 -212 82 -212 0 4
rlabel polysilicon 86 -206 86 -206 0 1
rlabel polysilicon 86 -212 86 -212 0 3
rlabel polysilicon 93 -206 93 -206 0 1
rlabel polysilicon 93 -212 93 -212 0 3
rlabel polysilicon 100 -206 100 -206 0 1
rlabel polysilicon 100 -212 100 -212 0 3
rlabel polysilicon 107 -206 107 -206 0 1
rlabel polysilicon 107 -212 107 -212 0 3
rlabel polysilicon 117 -206 117 -206 0 2
rlabel polysilicon 114 -212 114 -212 0 3
rlabel polysilicon 121 -206 121 -206 0 1
rlabel polysilicon 121 -212 121 -212 0 3
rlabel polysilicon 128 -212 128 -212 0 3
rlabel polysilicon 135 -206 135 -206 0 1
rlabel polysilicon 135 -212 135 -212 0 3
rlabel polysilicon 142 -206 142 -206 0 1
rlabel polysilicon 142 -212 142 -212 0 3
rlabel polysilicon 149 -206 149 -206 0 1
rlabel polysilicon 149 -212 149 -212 0 3
rlabel polysilicon 159 -206 159 -206 0 2
rlabel polysilicon 16 -231 16 -231 0 1
rlabel polysilicon 16 -237 16 -237 0 3
rlabel polysilicon 26 -231 26 -231 0 2
rlabel polysilicon 33 -231 33 -231 0 2
rlabel polysilicon 30 -237 30 -237 0 3
rlabel polysilicon 40 -231 40 -231 0 2
rlabel polysilicon 44 -231 44 -231 0 1
rlabel polysilicon 44 -237 44 -237 0 3
rlabel polysilicon 54 -231 54 -231 0 2
rlabel polysilicon 54 -237 54 -237 0 4
rlabel polysilicon 61 -231 61 -231 0 2
rlabel polysilicon 61 -237 61 -237 0 4
rlabel polysilicon 68 -231 68 -231 0 2
rlabel polysilicon 65 -237 65 -237 0 3
rlabel polysilicon 72 -231 72 -231 0 1
rlabel polysilicon 72 -237 72 -237 0 3
rlabel polysilicon 82 -231 82 -231 0 2
rlabel polysilicon 79 -237 79 -237 0 3
rlabel polysilicon 82 -237 82 -237 0 4
rlabel polysilicon 86 -237 86 -237 0 3
rlabel polysilicon 100 -231 100 -231 0 1
rlabel metal2 44 1 44 1 0 net=117
rlabel metal2 65 1 65 1 0 net=255
rlabel metal2 37 -10 37 -10 0 net=119
rlabel metal2 51 -10 51 -10 0 net=7
rlabel metal2 65 -10 65 -10 0 net=256
rlabel metal2 79 -10 79 -10 0 net=141
rlabel metal2 93 -10 93 -10 0 net=251
rlabel metal2 30 -12 30 -12 0 net=203
rlabel metal2 51 -12 51 -12 0 net=163
rlabel metal2 58 -14 58 -14 0 net=229
rlabel metal2 16 -25 16 -25 0 net=121
rlabel metal2 44 -25 44 -25 0 net=12
rlabel metal2 89 -25 89 -25 0 net=177
rlabel metal2 114 -25 114 -25 0 net=281
rlabel metal2 9 -27 9 -27 0 net=183
rlabel metal2 47 -27 47 -27 0 net=49
rlabel metal2 61 -27 61 -27 0 net=231
rlabel metal2 26 -29 26 -29 0 net=204
rlabel metal2 44 -29 44 -29 0 net=135
rlabel metal2 65 -29 65 -29 0 net=230
rlabel metal2 93 -29 93 -29 0 net=253
rlabel metal2 23 -31 23 -31 0 net=131
rlabel metal2 72 -31 72 -31 0 net=201
rlabel metal2 79 -33 79 -33 0 net=143
rlabel metal2 100 -33 100 -33 0 net=261
rlabel metal2 79 -35 79 -35 0 net=145
rlabel metal2 51 -37 51 -37 0 net=164
rlabel metal2 9 -48 9 -48 0 net=184
rlabel metal2 37 -48 37 -48 0 net=21
rlabel metal2 68 -48 68 -48 0 net=202
rlabel metal2 131 -48 131 -48 0 net=262
rlabel metal2 23 -50 23 -50 0 net=132
rlabel metal2 51 -50 51 -50 0 net=151
rlabel metal2 103 -50 103 -50 0 net=232
rlabel metal2 9 -52 9 -52 0 net=227
rlabel metal2 30 -52 30 -52 0 net=99
rlabel metal2 58 -52 58 -52 0 net=137
rlabel metal2 58 -52 58 -52 0 net=137
rlabel metal2 68 -52 68 -52 0 net=144
rlabel metal2 107 -52 107 -52 0 net=179
rlabel metal2 16 -54 16 -54 0 net=122
rlabel metal2 54 -54 54 -54 0 net=205
rlabel metal2 16 -56 16 -56 0 net=185
rlabel metal2 65 -56 65 -56 0 net=277
rlabel metal2 72 -58 72 -58 0 net=146
rlabel metal2 86 -58 86 -58 0 net=254
rlabel metal2 72 -60 72 -60 0 net=111
rlabel metal2 86 -60 86 -60 0 net=209
rlabel metal2 75 -62 75 -62 0 net=259
rlabel metal2 79 -64 79 -64 0 net=282
rlabel metal2 2 -75 2 -75 0 net=233
rlabel metal2 47 -75 47 -75 0 net=152
rlabel metal2 58 -75 58 -75 0 net=138
rlabel metal2 72 -75 72 -75 0 net=113
rlabel metal2 72 -75 72 -75 0 net=113
rlabel metal2 89 -75 89 -75 0 net=206
rlabel metal2 100 -75 100 -75 0 net=211
rlabel metal2 9 -77 9 -77 0 net=228
rlabel metal2 51 -77 51 -77 0 net=8
rlabel metal2 86 -77 86 -77 0 net=153
rlabel metal2 107 -77 107 -77 0 net=279
rlabel metal2 114 -77 114 -77 0 net=260
rlabel metal2 9 -79 9 -79 0 net=22
rlabel metal2 30 -79 30 -79 0 net=161
rlabel metal2 107 -79 107 -79 0 net=181
rlabel metal2 16 -81 16 -81 0 net=186
rlabel metal2 37 -81 37 -81 0 net=100
rlabel metal2 68 -81 68 -81 0 net=127
rlabel metal2 23 -83 23 -83 0 net=103
rlabel metal2 114 -83 114 -83 0 net=169
rlabel metal2 37 -85 37 -85 0 net=263
rlabel metal2 121 -85 121 -85 0 net=44
rlabel metal2 44 -87 44 -87 0 net=189
rlabel metal2 124 -87 124 -87 0 net=283
rlabel metal2 2 -98 2 -98 0 net=234
rlabel metal2 19 -98 19 -98 0 net=37
rlabel metal2 61 -98 61 -98 0 net=71
rlabel metal2 23 -100 23 -100 0 net=105
rlabel metal2 58 -100 58 -100 0 net=123
rlabel metal2 86 -100 86 -100 0 net=170
rlabel metal2 149 -100 149 -100 0 net=249
rlabel metal2 23 -102 23 -102 0 net=265
rlabel metal2 47 -102 47 -102 0 net=212
rlabel metal2 30 -104 30 -104 0 net=162
rlabel metal2 68 -104 68 -104 0 net=182
rlabel metal2 114 -104 114 -104 0 net=173
rlabel metal2 37 -106 37 -106 0 net=191
rlabel metal2 65 -106 65 -106 0 net=237
rlabel metal2 128 -106 128 -106 0 net=285
rlabel metal2 68 -108 68 -108 0 net=157
rlabel metal2 72 -110 72 -110 0 net=114
rlabel metal2 100 -110 100 -110 0 net=55
rlabel metal2 128 -110 128 -110 0 net=215
rlabel metal2 72 -112 72 -112 0 net=107
rlabel metal2 79 -114 79 -114 0 net=129
rlabel metal2 79 -116 79 -116 0 net=280
rlabel metal2 93 -118 93 -118 0 net=155
rlabel metal2 44 -120 44 -120 0 net=165
rlabel metal2 9 -131 9 -131 0 net=147
rlabel metal2 51 -131 51 -131 0 net=106
rlabel metal2 100 -131 100 -131 0 net=156
rlabel metal2 142 -131 142 -131 0 net=287
rlabel metal2 198 -131 198 -131 0 net=289
rlabel metal2 16 -133 16 -133 0 net=139
rlabel metal2 72 -133 72 -133 0 net=108
rlabel metal2 107 -133 107 -133 0 net=130
rlabel metal2 149 -133 149 -133 0 net=159
rlabel metal2 23 -135 23 -135 0 net=266
rlabel metal2 75 -135 75 -135 0 net=101
rlabel metal2 100 -135 100 -135 0 net=115
rlabel metal2 110 -135 110 -135 0 net=267
rlabel metal2 2 -137 2 -137 0 net=133
rlabel metal2 103 -137 103 -137 0 net=269
rlabel metal2 149 -137 149 -137 0 net=217
rlabel metal2 170 -137 170 -137 0 net=75
rlabel metal2 23 -139 23 -139 0 net=125
rlabel metal2 86 -139 86 -139 0 net=109
rlabel metal2 30 -141 30 -141 0 net=192
rlabel metal2 47 -141 47 -141 0 net=223
rlabel metal2 114 -141 114 -141 0 net=175
rlabel metal2 156 -141 156 -141 0 net=250
rlabel metal2 30 -143 30 -143 0 net=95
rlabel metal2 93 -143 93 -143 0 net=167
rlabel metal2 121 -143 121 -143 0 net=239
rlabel metal2 33 -145 33 -145 0 net=195
rlabel metal2 93 -147 93 -147 0 net=207
rlabel metal2 16 -158 16 -158 0 net=140
rlabel metal2 54 -158 54 -158 0 net=240
rlabel metal2 166 -158 166 -158 0 net=268
rlabel metal2 23 -160 23 -160 0 net=126
rlabel metal2 68 -160 68 -160 0 net=102
rlabel metal2 89 -160 89 -160 0 net=116
rlabel metal2 107 -160 107 -160 0 net=168
rlabel metal2 121 -160 121 -160 0 net=208
rlabel metal2 163 -160 163 -160 0 net=1
rlabel metal2 9 -162 9 -162 0 net=149
rlabel metal2 93 -162 93 -162 0 net=176
rlabel metal2 30 -164 30 -164 0 net=96
rlabel metal2 58 -164 58 -164 0 net=90
rlabel metal2 107 -164 107 -164 0 net=245
rlabel metal2 128 -164 128 -164 0 net=271
rlabel metal2 37 -166 37 -166 0 net=218
rlabel metal2 2 -168 2 -168 0 net=134
rlabel metal2 40 -168 40 -168 0 net=39
rlabel metal2 86 -168 86 -168 0 net=225
rlabel metal2 23 -170 23 -170 0 net=197
rlabel metal2 110 -170 110 -170 0 net=288
rlabel metal2 47 -172 47 -172 0 net=241
rlabel metal2 61 -172 61 -172 0 net=160
rlabel metal2 110 -174 110 -174 0 net=196
rlabel metal2 142 -176 142 -176 0 net=110
rlabel metal2 170 -178 170 -178 0 net=291
rlabel metal2 2 -189 2 -189 0 net=199
rlabel metal2 30 -189 30 -189 0 net=97
rlabel metal2 89 -189 89 -189 0 net=226
rlabel metal2 135 -189 135 -189 0 net=273
rlabel metal2 135 -189 135 -189 0 net=273
rlabel metal2 142 -189 142 -189 0 net=292
rlabel metal2 9 -191 9 -191 0 net=193
rlabel metal2 40 -191 40 -191 0 net=150
rlabel metal2 114 -191 114 -191 0 net=247
rlabel metal2 16 -193 16 -193 0 net=171
rlabel metal2 58 -193 58 -193 0 net=243
rlabel metal2 117 -193 117 -193 0 net=38
rlabel metal2 12 -195 12 -195 0 net=80
rlabel metal2 61 -195 61 -195 0 net=293
rlabel metal2 23 -197 23 -197 0 net=219
rlabel metal2 65 -197 65 -197 0 net=213
rlabel metal2 40 -199 40 -199 0 net=221
rlabel metal2 65 -201 65 -201 0 net=91
rlabel metal2 79 -201 79 -201 0 net=187
rlabel metal2 68 -203 68 -203 0 net=275
rlabel metal2 2 -214 2 -214 0 net=200
rlabel metal2 51 -214 51 -214 0 net=244
rlabel metal2 128 -214 128 -214 0 net=274
rlabel metal2 9 -216 9 -216 0 net=194
rlabel metal2 72 -216 72 -216 0 net=93
rlabel metal2 72 -216 72 -216 0 net=93
rlabel metal2 79 -216 79 -216 0 net=248
rlabel metal2 23 -218 23 -218 0 net=220
rlabel metal2 61 -218 61 -218 0 net=214
rlabel metal2 30 -220 30 -220 0 net=98
rlabel metal2 65 -220 65 -220 0 net=222
rlabel metal2 100 -220 100 -220 0 net=294
rlabel metal2 33 -222 33 -222 0 net=57
rlabel metal2 82 -222 82 -222 0 net=9
rlabel metal2 40 -224 40 -224 0 net=188
rlabel metal2 16 -226 16 -226 0 net=172
rlabel metal2 44 -226 44 -226 0 net=235
rlabel metal2 82 -226 82 -226 0 net=276
rlabel metal2 16 -228 16 -228 0 net=257
rlabel metal2 16 -239 16 -239 0 net=258
rlabel metal2 44 -239 44 -239 0 net=236
rlabel metal2 54 -241 54 -241 0 net=59
rlabel metal2 61 -243 61 -243 0 net=94
rlabel metal2 65 -245 65 -245 0 net=87
<< end >>
