magic
tech scmos
timestamp 1555016725 
<< pdiffusion >>
rect 1 -8 7 -2
rect 8 -8 14 -2
rect 15 -8 21 -2
rect 22 -8 28 -2
rect 71 -8 77 -2
rect 78 -8 81 -2
rect 99 -8 105 -2
rect 106 -8 109 -2
rect 113 -8 119 -2
rect 120 -8 126 -2
rect 127 -8 130 -2
rect 1 -29 7 -23
rect 8 -29 14 -23
rect 43 -29 46 -23
rect 50 -29 53 -23
rect 57 -29 63 -23
rect 64 -29 70 -23
rect 71 -29 74 -23
rect 78 -29 84 -23
rect 85 -29 88 -23
rect 92 -29 98 -23
rect 99 -29 102 -23
rect 106 -29 112 -23
rect 113 -29 119 -23
rect 120 -29 123 -23
rect 127 -29 130 -23
rect 134 -29 137 -23
rect 141 -29 144 -23
rect 155 -29 161 -23
rect 260 -29 266 -23
rect 1 -50 7 -44
rect 8 -50 14 -44
rect 29 -50 35 -44
rect 36 -50 42 -44
rect 43 -50 46 -44
rect 50 -50 53 -44
rect 57 -50 63 -44
rect 64 -50 70 -44
rect 71 -50 77 -44
rect 78 -50 81 -44
rect 85 -50 91 -44
rect 92 -50 95 -44
rect 99 -50 102 -44
rect 106 -50 109 -44
rect 113 -50 119 -44
rect 127 -50 133 -44
rect 134 -50 137 -44
rect 141 -50 144 -44
rect 148 -50 154 -44
rect 162 -50 168 -44
rect 169 -50 172 -44
rect 176 -50 179 -44
rect 232 -50 238 -44
rect 246 -50 249 -44
rect 1 -73 4 -67
rect 8 -73 14 -67
rect 15 -73 21 -67
rect 22 -73 25 -67
rect 29 -73 35 -67
rect 36 -73 42 -67
rect 43 -73 46 -67
rect 50 -73 53 -67
rect 57 -73 60 -67
rect 64 -73 67 -67
rect 71 -73 77 -67
rect 78 -73 84 -67
rect 85 -73 91 -67
rect 92 -73 98 -67
rect 99 -73 102 -67
rect 106 -73 109 -67
rect 113 -73 119 -67
rect 120 -73 123 -67
rect 127 -73 130 -67
rect 134 -73 140 -67
rect 141 -73 144 -67
rect 148 -73 151 -67
rect 155 -73 158 -67
rect 162 -73 165 -67
rect 169 -73 175 -67
rect 176 -73 179 -67
rect 183 -73 186 -67
rect 190 -73 196 -67
rect 197 -73 200 -67
rect 204 -73 207 -67
rect 211 -73 217 -67
rect 218 -73 221 -67
rect 225 -73 231 -67
rect 232 -73 235 -67
rect 8 -102 11 -96
rect 15 -102 18 -96
rect 22 -102 25 -96
rect 29 -102 35 -96
rect 36 -102 39 -96
rect 43 -102 49 -96
rect 50 -102 56 -96
rect 57 -102 60 -96
rect 64 -102 70 -96
rect 71 -102 74 -96
rect 78 -102 84 -96
rect 85 -102 88 -96
rect 92 -102 98 -96
rect 99 -102 102 -96
rect 106 -102 109 -96
rect 113 -102 116 -96
rect 120 -102 126 -96
rect 127 -102 133 -96
rect 134 -102 140 -96
rect 141 -102 147 -96
rect 148 -102 154 -96
rect 155 -102 158 -96
rect 162 -102 168 -96
rect 169 -102 172 -96
rect 176 -102 179 -96
rect 183 -102 186 -96
rect 190 -102 193 -96
rect 197 -102 200 -96
rect 204 -102 207 -96
rect 211 -102 214 -96
rect 218 -102 221 -96
rect 225 -102 228 -96
rect 232 -102 235 -96
rect 239 -102 242 -96
rect 246 -102 249 -96
rect 253 -102 256 -96
rect 260 -102 266 -96
rect 267 -102 273 -96
rect 281 -102 284 -96
rect 8 -135 11 -129
rect 15 -135 18 -129
rect 22 -135 25 -129
rect 29 -135 35 -129
rect 36 -135 42 -129
rect 43 -135 49 -129
rect 50 -135 53 -129
rect 57 -135 60 -129
rect 64 -135 67 -129
rect 71 -135 77 -129
rect 78 -135 81 -129
rect 85 -135 88 -129
rect 92 -135 98 -129
rect 99 -135 102 -129
rect 106 -135 112 -129
rect 113 -135 119 -129
rect 120 -135 123 -129
rect 127 -135 130 -129
rect 134 -135 140 -129
rect 141 -135 144 -129
rect 148 -135 154 -129
rect 155 -135 161 -129
rect 162 -135 165 -129
rect 169 -135 175 -129
rect 176 -135 182 -129
rect 183 -135 189 -129
rect 190 -135 193 -129
rect 197 -135 200 -129
rect 204 -135 210 -129
rect 211 -135 214 -129
rect 218 -135 221 -129
rect 225 -135 228 -129
rect 232 -135 235 -129
rect 295 -135 298 -129
rect 1 -178 4 -172
rect 8 -178 11 -172
rect 15 -178 18 -172
rect 22 -178 25 -172
rect 29 -178 35 -172
rect 36 -178 39 -172
rect 43 -178 46 -172
rect 50 -178 56 -172
rect 57 -178 60 -172
rect 64 -178 70 -172
rect 71 -178 74 -172
rect 78 -178 81 -172
rect 85 -178 91 -172
rect 92 -178 98 -172
rect 99 -178 105 -172
rect 106 -178 112 -172
rect 113 -178 119 -172
rect 120 -178 126 -172
rect 127 -178 133 -172
rect 134 -178 140 -172
rect 141 -178 144 -172
rect 148 -178 154 -172
rect 155 -178 158 -172
rect 162 -178 168 -172
rect 169 -178 172 -172
rect 176 -178 179 -172
rect 183 -178 186 -172
rect 190 -178 193 -172
rect 197 -178 200 -172
rect 204 -178 207 -172
rect 211 -178 214 -172
rect 218 -178 221 -172
rect 225 -178 228 -172
rect 232 -178 235 -172
rect 239 -178 242 -172
rect 246 -178 249 -172
rect 253 -178 256 -172
rect 260 -178 263 -172
rect 267 -178 270 -172
rect 274 -178 277 -172
rect 281 -178 284 -172
rect 29 -217 32 -211
rect 36 -217 39 -211
rect 43 -217 49 -211
rect 50 -217 56 -211
rect 57 -217 63 -211
rect 64 -217 67 -211
rect 71 -217 77 -211
rect 78 -217 81 -211
rect 85 -217 91 -211
rect 92 -217 98 -211
rect 99 -217 102 -211
rect 106 -217 112 -211
rect 113 -217 116 -211
rect 120 -217 123 -211
rect 127 -217 133 -211
rect 134 -217 137 -211
rect 141 -217 147 -211
rect 148 -217 154 -211
rect 155 -217 158 -211
rect 162 -217 168 -211
rect 169 -217 175 -211
rect 176 -217 179 -211
rect 183 -217 186 -211
rect 190 -217 193 -211
rect 197 -217 200 -211
rect 204 -217 207 -211
rect 218 -217 224 -211
rect 225 -217 228 -211
rect 8 -254 11 -248
rect 15 -254 18 -248
rect 22 -254 25 -248
rect 29 -254 35 -248
rect 36 -254 39 -248
rect 43 -254 49 -248
rect 50 -254 56 -248
rect 57 -254 63 -248
rect 64 -254 67 -248
rect 71 -254 74 -248
rect 78 -254 84 -248
rect 85 -254 91 -248
rect 92 -254 95 -248
rect 99 -254 102 -248
rect 106 -254 112 -248
rect 113 -254 116 -248
rect 120 -254 126 -248
rect 127 -254 130 -248
rect 134 -254 140 -248
rect 141 -254 147 -248
rect 148 -254 154 -248
rect 155 -254 158 -248
rect 162 -254 165 -248
rect 169 -254 172 -248
rect 176 -254 179 -248
rect 183 -254 186 -248
rect 190 -254 193 -248
rect 197 -254 200 -248
rect 204 -254 207 -248
rect 211 -254 214 -248
rect 218 -254 221 -248
rect 225 -254 228 -248
rect 232 -254 238 -248
rect 239 -254 242 -248
rect 246 -254 249 -248
rect 253 -254 256 -248
rect 260 -254 263 -248
rect 267 -254 273 -248
rect 274 -254 280 -248
rect 295 -254 298 -248
rect 1 -293 7 -287
rect 8 -293 11 -287
rect 15 -293 18 -287
rect 22 -293 28 -287
rect 29 -293 35 -287
rect 36 -293 42 -287
rect 43 -293 46 -287
rect 50 -293 56 -287
rect 57 -293 60 -287
rect 64 -293 67 -287
rect 71 -293 77 -287
rect 78 -293 84 -287
rect 85 -293 91 -287
rect 92 -293 98 -287
rect 99 -293 102 -287
rect 106 -293 109 -287
rect 113 -293 116 -287
rect 120 -293 123 -287
rect 127 -293 130 -287
rect 134 -293 137 -287
rect 141 -293 147 -287
rect 148 -293 151 -287
rect 155 -293 158 -287
rect 162 -293 165 -287
rect 169 -293 172 -287
rect 176 -293 182 -287
rect 183 -293 186 -287
rect 190 -293 193 -287
rect 197 -293 203 -287
rect 204 -293 207 -287
rect 211 -293 214 -287
rect 218 -293 221 -287
rect 225 -293 228 -287
rect 232 -293 235 -287
rect 239 -293 242 -287
rect 246 -293 252 -287
rect 253 -293 256 -287
rect 260 -293 263 -287
rect 267 -293 273 -287
rect 274 -293 277 -287
rect 1 -330 7 -324
rect 8 -330 11 -324
rect 15 -330 18 -324
rect 22 -330 25 -324
rect 29 -330 32 -324
rect 36 -330 42 -324
rect 43 -330 49 -324
rect 50 -330 53 -324
rect 57 -330 60 -324
rect 64 -330 67 -324
rect 71 -330 77 -324
rect 78 -330 81 -324
rect 85 -330 91 -324
rect 92 -330 98 -324
rect 99 -330 105 -324
rect 106 -330 109 -324
rect 113 -330 119 -324
rect 120 -330 123 -324
rect 127 -330 133 -324
rect 134 -330 137 -324
rect 141 -330 147 -324
rect 148 -330 154 -324
rect 155 -330 161 -324
rect 162 -330 165 -324
rect 169 -330 172 -324
rect 176 -330 179 -324
rect 183 -330 186 -324
rect 190 -330 193 -324
rect 197 -330 200 -324
rect 204 -330 207 -324
rect 211 -330 214 -324
rect 218 -330 224 -324
rect 225 -330 228 -324
rect 1 -361 7 -355
rect 22 -361 25 -355
rect 29 -361 32 -355
rect 36 -361 39 -355
rect 43 -361 49 -355
rect 50 -361 56 -355
rect 57 -361 63 -355
rect 64 -361 70 -355
rect 71 -361 74 -355
rect 78 -361 81 -355
rect 85 -361 91 -355
rect 92 -361 98 -355
rect 99 -361 102 -355
rect 106 -361 109 -355
rect 113 -361 119 -355
rect 120 -361 123 -355
rect 127 -361 130 -355
rect 134 -361 137 -355
rect 141 -361 144 -355
rect 148 -361 151 -355
rect 155 -361 161 -355
rect 162 -361 165 -355
rect 169 -361 175 -355
rect 176 -361 179 -355
rect 183 -361 186 -355
rect 190 -361 193 -355
rect 197 -361 200 -355
rect 204 -361 210 -355
rect 211 -361 217 -355
rect 8 -394 14 -388
rect 15 -394 18 -388
rect 22 -394 25 -388
rect 29 -394 32 -388
rect 36 -394 42 -388
rect 43 -394 49 -388
rect 50 -394 56 -388
rect 57 -394 60 -388
rect 64 -394 67 -388
rect 71 -394 74 -388
rect 78 -394 81 -388
rect 85 -394 91 -388
rect 92 -394 98 -388
rect 99 -394 102 -388
rect 106 -394 112 -388
rect 113 -394 119 -388
rect 120 -394 123 -388
rect 127 -394 133 -388
rect 134 -394 140 -388
rect 141 -394 144 -388
rect 148 -394 154 -388
rect 155 -394 158 -388
rect 162 -394 165 -388
rect 169 -394 172 -388
rect 176 -394 179 -388
rect 183 -394 189 -388
rect 190 -394 193 -388
rect 197 -394 203 -388
rect 204 -394 207 -388
rect 211 -394 214 -388
rect 218 -394 224 -388
rect 225 -394 228 -388
rect 8 -427 14 -421
rect 15 -427 21 -421
rect 22 -427 28 -421
rect 29 -427 32 -421
rect 43 -427 49 -421
rect 50 -427 56 -421
rect 57 -427 63 -421
rect 64 -427 67 -421
rect 71 -427 77 -421
rect 78 -427 84 -421
rect 85 -427 91 -421
rect 92 -427 98 -421
rect 99 -427 102 -421
rect 106 -427 109 -421
rect 113 -427 116 -421
rect 120 -427 126 -421
rect 127 -427 130 -421
rect 134 -427 140 -421
rect 141 -427 144 -421
rect 148 -427 151 -421
rect 155 -427 158 -421
rect 183 -427 189 -421
rect 197 -427 203 -421
<< polysilicon >>
rect 72 -3 73 -1
rect 75 -9 76 -7
rect 79 -3 80 -1
rect 79 -9 80 -7
rect 100 -3 101 -1
rect 107 -3 108 -1
rect 107 -9 108 -7
rect 114 -9 115 -7
rect 121 -3 122 -1
rect 128 -3 129 -1
rect 128 -9 129 -7
rect 44 -24 45 -22
rect 44 -30 45 -28
rect 51 -24 52 -22
rect 51 -30 52 -28
rect 61 -24 62 -22
rect 68 -24 69 -22
rect 72 -24 73 -22
rect 72 -30 73 -28
rect 79 -24 80 -22
rect 82 -24 83 -22
rect 86 -24 87 -22
rect 86 -30 87 -28
rect 96 -24 97 -22
rect 93 -30 94 -28
rect 100 -24 101 -22
rect 100 -30 101 -28
rect 107 -24 108 -22
rect 110 -24 111 -22
rect 117 -24 118 -22
rect 121 -24 122 -22
rect 121 -30 122 -28
rect 128 -24 129 -22
rect 128 -30 129 -28
rect 135 -24 136 -22
rect 135 -30 136 -28
rect 142 -24 143 -22
rect 142 -30 143 -28
rect 159 -30 160 -28
rect 264 -30 265 -28
rect 30 -51 31 -49
rect 40 -51 41 -49
rect 44 -45 45 -43
rect 44 -51 45 -49
rect 51 -45 52 -43
rect 51 -51 52 -49
rect 58 -45 59 -43
rect 61 -45 62 -43
rect 58 -51 59 -49
rect 61 -51 62 -49
rect 65 -45 66 -43
rect 65 -51 66 -49
rect 72 -45 73 -43
rect 75 -45 76 -43
rect 79 -45 80 -43
rect 79 -51 80 -49
rect 86 -45 87 -43
rect 86 -51 87 -49
rect 89 -51 90 -49
rect 93 -45 94 -43
rect 93 -51 94 -49
rect 100 -45 101 -43
rect 100 -51 101 -49
rect 107 -45 108 -43
rect 107 -51 108 -49
rect 114 -51 115 -49
rect 128 -45 129 -43
rect 131 -45 132 -43
rect 135 -45 136 -43
rect 135 -51 136 -49
rect 142 -45 143 -43
rect 142 -51 143 -49
rect 149 -45 150 -43
rect 152 -51 153 -49
rect 163 -45 164 -43
rect 166 -45 167 -43
rect 163 -51 164 -49
rect 170 -45 171 -43
rect 170 -51 171 -49
rect 177 -45 178 -43
rect 177 -51 178 -49
rect 233 -51 234 -49
rect 236 -51 237 -49
rect 247 -45 248 -43
rect 247 -51 248 -49
rect 2 -68 3 -66
rect 2 -74 3 -72
rect 19 -74 20 -72
rect 23 -68 24 -66
rect 23 -74 24 -72
rect 33 -68 34 -66
rect 30 -74 31 -72
rect 37 -68 38 -66
rect 44 -68 45 -66
rect 44 -74 45 -72
rect 51 -68 52 -66
rect 51 -74 52 -72
rect 58 -68 59 -66
rect 58 -74 59 -72
rect 65 -68 66 -66
rect 65 -74 66 -72
rect 72 -68 73 -66
rect 75 -68 76 -66
rect 72 -74 73 -72
rect 79 -74 80 -72
rect 86 -68 87 -66
rect 93 -68 94 -66
rect 96 -68 97 -66
rect 93 -74 94 -72
rect 100 -68 101 -66
rect 100 -74 101 -72
rect 107 -68 108 -66
rect 107 -74 108 -72
rect 117 -68 118 -66
rect 117 -74 118 -72
rect 121 -68 122 -66
rect 121 -74 122 -72
rect 128 -68 129 -66
rect 128 -74 129 -72
rect 135 -68 136 -66
rect 138 -68 139 -66
rect 135 -74 136 -72
rect 142 -68 143 -66
rect 142 -74 143 -72
rect 149 -68 150 -66
rect 149 -74 150 -72
rect 156 -68 157 -66
rect 156 -74 157 -72
rect 163 -68 164 -66
rect 163 -74 164 -72
rect 170 -68 171 -66
rect 173 -74 174 -72
rect 177 -68 178 -66
rect 177 -74 178 -72
rect 184 -68 185 -66
rect 184 -74 185 -72
rect 191 -68 192 -66
rect 194 -68 195 -66
rect 191 -74 192 -72
rect 198 -68 199 -66
rect 198 -74 199 -72
rect 205 -68 206 -66
rect 205 -74 206 -72
rect 212 -68 213 -66
rect 212 -74 213 -72
rect 219 -68 220 -66
rect 219 -74 220 -72
rect 229 -68 230 -66
rect 233 -68 234 -66
rect 233 -74 234 -72
rect 9 -97 10 -95
rect 9 -103 10 -101
rect 16 -97 17 -95
rect 16 -103 17 -101
rect 23 -97 24 -95
rect 23 -103 24 -101
rect 30 -97 31 -95
rect 30 -103 31 -101
rect 37 -97 38 -95
rect 37 -103 38 -101
rect 44 -97 45 -95
rect 44 -103 45 -101
rect 51 -97 52 -95
rect 54 -97 55 -95
rect 58 -97 59 -95
rect 58 -103 59 -101
rect 68 -97 69 -95
rect 65 -103 66 -101
rect 68 -103 69 -101
rect 72 -97 73 -95
rect 72 -103 73 -101
rect 79 -97 80 -95
rect 79 -103 80 -101
rect 86 -97 87 -95
rect 86 -103 87 -101
rect 93 -97 94 -95
rect 96 -97 97 -95
rect 96 -103 97 -101
rect 100 -97 101 -95
rect 100 -103 101 -101
rect 107 -97 108 -95
rect 107 -103 108 -101
rect 114 -97 115 -95
rect 114 -103 115 -101
rect 124 -97 125 -95
rect 121 -103 122 -101
rect 124 -103 125 -101
rect 128 -97 129 -95
rect 131 -97 132 -95
rect 135 -97 136 -95
rect 135 -103 136 -101
rect 138 -103 139 -101
rect 145 -97 146 -95
rect 142 -103 143 -101
rect 149 -97 150 -95
rect 149 -103 150 -101
rect 152 -103 153 -101
rect 156 -97 157 -95
rect 156 -103 157 -101
rect 163 -103 164 -101
rect 166 -103 167 -101
rect 170 -97 171 -95
rect 170 -103 171 -101
rect 177 -97 178 -95
rect 177 -103 178 -101
rect 184 -97 185 -95
rect 184 -103 185 -101
rect 191 -97 192 -95
rect 191 -103 192 -101
rect 198 -97 199 -95
rect 198 -103 199 -101
rect 205 -97 206 -95
rect 205 -103 206 -101
rect 212 -97 213 -95
rect 212 -103 213 -101
rect 219 -97 220 -95
rect 219 -103 220 -101
rect 226 -97 227 -95
rect 226 -103 227 -101
rect 233 -97 234 -95
rect 233 -103 234 -101
rect 240 -97 241 -95
rect 240 -103 241 -101
rect 247 -97 248 -95
rect 247 -103 248 -101
rect 254 -97 255 -95
rect 254 -103 255 -101
rect 264 -97 265 -95
rect 261 -103 262 -101
rect 268 -103 269 -101
rect 282 -97 283 -95
rect 282 -103 283 -101
rect 9 -130 10 -128
rect 9 -136 10 -134
rect 16 -130 17 -128
rect 16 -136 17 -134
rect 23 -130 24 -128
rect 23 -136 24 -134
rect 33 -130 34 -128
rect 30 -136 31 -134
rect 33 -136 34 -134
rect 37 -130 38 -128
rect 37 -136 38 -134
rect 40 -136 41 -134
rect 47 -130 48 -128
rect 51 -130 52 -128
rect 51 -136 52 -134
rect 58 -130 59 -128
rect 58 -136 59 -134
rect 65 -130 66 -128
rect 65 -136 66 -134
rect 72 -136 73 -134
rect 79 -130 80 -128
rect 79 -136 80 -134
rect 86 -130 87 -128
rect 86 -136 87 -134
rect 93 -130 94 -128
rect 93 -136 94 -134
rect 96 -136 97 -134
rect 100 -130 101 -128
rect 100 -136 101 -134
rect 110 -130 111 -128
rect 107 -136 108 -134
rect 110 -136 111 -134
rect 114 -130 115 -128
rect 117 -130 118 -128
rect 114 -136 115 -134
rect 117 -136 118 -134
rect 121 -130 122 -128
rect 121 -136 122 -134
rect 128 -130 129 -128
rect 128 -136 129 -134
rect 135 -130 136 -128
rect 135 -136 136 -134
rect 138 -136 139 -134
rect 142 -130 143 -128
rect 142 -136 143 -134
rect 149 -136 150 -134
rect 159 -136 160 -134
rect 163 -130 164 -128
rect 163 -136 164 -134
rect 173 -130 174 -128
rect 177 -130 178 -128
rect 180 -136 181 -134
rect 187 -130 188 -128
rect 184 -136 185 -134
rect 191 -130 192 -128
rect 191 -136 192 -134
rect 198 -130 199 -128
rect 198 -136 199 -134
rect 208 -130 209 -128
rect 208 -136 209 -134
rect 212 -130 213 -128
rect 212 -136 213 -134
rect 219 -130 220 -128
rect 219 -136 220 -134
rect 226 -130 227 -128
rect 226 -136 227 -134
rect 233 -130 234 -128
rect 233 -136 234 -134
rect 296 -130 297 -128
rect 296 -136 297 -134
rect 2 -173 3 -171
rect 2 -179 3 -177
rect 9 -173 10 -171
rect 9 -179 10 -177
rect 16 -173 17 -171
rect 16 -179 17 -177
rect 23 -173 24 -171
rect 23 -179 24 -177
rect 33 -179 34 -177
rect 37 -173 38 -171
rect 37 -179 38 -177
rect 44 -173 45 -171
rect 44 -179 45 -177
rect 51 -173 52 -171
rect 54 -173 55 -171
rect 58 -173 59 -171
rect 58 -179 59 -177
rect 65 -179 66 -177
rect 68 -179 69 -177
rect 72 -173 73 -171
rect 72 -179 73 -177
rect 79 -173 80 -171
rect 79 -179 80 -177
rect 86 -173 87 -171
rect 89 -173 90 -171
rect 86 -179 87 -177
rect 89 -179 90 -177
rect 93 -173 94 -171
rect 93 -179 94 -177
rect 96 -179 97 -177
rect 100 -173 101 -171
rect 103 -173 104 -171
rect 100 -179 101 -177
rect 103 -179 104 -177
rect 107 -173 108 -171
rect 107 -179 108 -177
rect 110 -179 111 -177
rect 114 -173 115 -171
rect 117 -173 118 -171
rect 114 -179 115 -177
rect 117 -179 118 -177
rect 124 -173 125 -171
rect 121 -179 122 -177
rect 128 -173 129 -171
rect 131 -173 132 -171
rect 128 -179 129 -177
rect 131 -179 132 -177
rect 135 -173 136 -171
rect 138 -173 139 -171
rect 135 -179 136 -177
rect 142 -173 143 -171
rect 142 -179 143 -177
rect 149 -173 150 -171
rect 152 -173 153 -171
rect 152 -179 153 -177
rect 156 -173 157 -171
rect 156 -179 157 -177
rect 163 -173 164 -171
rect 163 -179 164 -177
rect 170 -173 171 -171
rect 170 -179 171 -177
rect 177 -173 178 -171
rect 177 -179 178 -177
rect 184 -173 185 -171
rect 184 -179 185 -177
rect 191 -173 192 -171
rect 191 -179 192 -177
rect 198 -173 199 -171
rect 198 -179 199 -177
rect 205 -173 206 -171
rect 205 -179 206 -177
rect 212 -173 213 -171
rect 212 -179 213 -177
rect 219 -173 220 -171
rect 219 -179 220 -177
rect 226 -173 227 -171
rect 226 -179 227 -177
rect 233 -173 234 -171
rect 233 -179 234 -177
rect 240 -173 241 -171
rect 240 -179 241 -177
rect 247 -173 248 -171
rect 247 -179 248 -177
rect 254 -173 255 -171
rect 254 -179 255 -177
rect 261 -173 262 -171
rect 261 -179 262 -177
rect 268 -173 269 -171
rect 268 -179 269 -177
rect 275 -173 276 -171
rect 275 -179 276 -177
rect 282 -173 283 -171
rect 282 -179 283 -177
rect 30 -212 31 -210
rect 30 -218 31 -216
rect 37 -212 38 -210
rect 37 -218 38 -216
rect 44 -212 45 -210
rect 44 -218 45 -216
rect 54 -212 55 -210
rect 51 -218 52 -216
rect 61 -212 62 -210
rect 61 -218 62 -216
rect 65 -212 66 -210
rect 65 -218 66 -216
rect 75 -218 76 -216
rect 79 -212 80 -210
rect 79 -218 80 -216
rect 86 -212 87 -210
rect 89 -212 90 -210
rect 86 -218 87 -216
rect 96 -212 97 -210
rect 93 -218 94 -216
rect 100 -212 101 -210
rect 100 -218 101 -216
rect 110 -212 111 -210
rect 107 -218 108 -216
rect 110 -218 111 -216
rect 114 -212 115 -210
rect 114 -218 115 -216
rect 121 -212 122 -210
rect 121 -218 122 -216
rect 128 -212 129 -210
rect 131 -218 132 -216
rect 135 -212 136 -210
rect 135 -218 136 -216
rect 142 -212 143 -210
rect 145 -212 146 -210
rect 149 -212 150 -210
rect 152 -212 153 -210
rect 152 -218 153 -216
rect 156 -212 157 -210
rect 156 -218 157 -216
rect 163 -212 164 -210
rect 166 -212 167 -210
rect 166 -218 167 -216
rect 170 -218 171 -216
rect 173 -218 174 -216
rect 177 -212 178 -210
rect 177 -218 178 -216
rect 184 -212 185 -210
rect 184 -218 185 -216
rect 191 -212 192 -210
rect 191 -218 192 -216
rect 198 -212 199 -210
rect 198 -218 199 -216
rect 205 -212 206 -210
rect 205 -218 206 -216
rect 219 -212 220 -210
rect 222 -212 223 -210
rect 219 -218 220 -216
rect 222 -218 223 -216
rect 226 -212 227 -210
rect 226 -218 227 -216
rect 9 -249 10 -247
rect 9 -255 10 -253
rect 16 -249 17 -247
rect 16 -255 17 -253
rect 23 -249 24 -247
rect 23 -255 24 -253
rect 30 -249 31 -247
rect 33 -249 34 -247
rect 37 -249 38 -247
rect 37 -255 38 -253
rect 47 -249 48 -247
rect 47 -255 48 -253
rect 54 -249 55 -247
rect 51 -255 52 -253
rect 61 -249 62 -247
rect 58 -255 59 -253
rect 65 -249 66 -247
rect 65 -255 66 -253
rect 72 -249 73 -247
rect 72 -255 73 -253
rect 79 -249 80 -247
rect 79 -255 80 -253
rect 89 -249 90 -247
rect 86 -255 87 -253
rect 89 -255 90 -253
rect 93 -249 94 -247
rect 93 -255 94 -253
rect 100 -249 101 -247
rect 100 -255 101 -253
rect 110 -249 111 -247
rect 110 -255 111 -253
rect 114 -249 115 -247
rect 114 -255 115 -253
rect 121 -249 122 -247
rect 121 -255 122 -253
rect 128 -249 129 -247
rect 128 -255 129 -253
rect 135 -249 136 -247
rect 138 -249 139 -247
rect 135 -255 136 -253
rect 138 -255 139 -253
rect 145 -249 146 -247
rect 142 -255 143 -253
rect 149 -249 150 -247
rect 152 -249 153 -247
rect 149 -255 150 -253
rect 152 -255 153 -253
rect 156 -249 157 -247
rect 156 -255 157 -253
rect 163 -249 164 -247
rect 163 -255 164 -253
rect 170 -249 171 -247
rect 170 -255 171 -253
rect 177 -249 178 -247
rect 177 -255 178 -253
rect 184 -249 185 -247
rect 184 -255 185 -253
rect 191 -249 192 -247
rect 191 -255 192 -253
rect 198 -249 199 -247
rect 198 -255 199 -253
rect 205 -249 206 -247
rect 205 -255 206 -253
rect 212 -249 213 -247
rect 212 -255 213 -253
rect 219 -249 220 -247
rect 219 -255 220 -253
rect 226 -249 227 -247
rect 226 -255 227 -253
rect 233 -249 234 -247
rect 236 -255 237 -253
rect 240 -249 241 -247
rect 240 -255 241 -253
rect 247 -249 248 -247
rect 247 -255 248 -253
rect 254 -249 255 -247
rect 254 -255 255 -253
rect 261 -249 262 -247
rect 261 -255 262 -253
rect 268 -249 269 -247
rect 275 -249 276 -247
rect 278 -249 279 -247
rect 296 -249 297 -247
rect 296 -255 297 -253
rect 2 -294 3 -292
rect 9 -288 10 -286
rect 9 -294 10 -292
rect 16 -288 17 -286
rect 16 -294 17 -292
rect 23 -288 24 -286
rect 26 -288 27 -286
rect 33 -288 34 -286
rect 37 -294 38 -292
rect 44 -288 45 -286
rect 44 -294 45 -292
rect 51 -288 52 -286
rect 58 -288 59 -286
rect 58 -294 59 -292
rect 65 -288 66 -286
rect 65 -294 66 -292
rect 75 -288 76 -286
rect 72 -294 73 -292
rect 75 -294 76 -292
rect 79 -288 80 -286
rect 79 -294 80 -292
rect 82 -294 83 -292
rect 86 -288 87 -286
rect 89 -288 90 -286
rect 89 -294 90 -292
rect 93 -294 94 -292
rect 96 -294 97 -292
rect 100 -288 101 -286
rect 100 -294 101 -292
rect 107 -288 108 -286
rect 107 -294 108 -292
rect 114 -288 115 -286
rect 114 -294 115 -292
rect 121 -288 122 -286
rect 121 -294 122 -292
rect 128 -288 129 -286
rect 128 -294 129 -292
rect 135 -288 136 -286
rect 135 -294 136 -292
rect 142 -288 143 -286
rect 145 -288 146 -286
rect 142 -294 143 -292
rect 145 -294 146 -292
rect 149 -288 150 -286
rect 149 -294 150 -292
rect 156 -288 157 -286
rect 156 -294 157 -292
rect 163 -288 164 -286
rect 163 -294 164 -292
rect 170 -288 171 -286
rect 170 -294 171 -292
rect 177 -288 178 -286
rect 180 -288 181 -286
rect 177 -294 178 -292
rect 184 -288 185 -286
rect 184 -294 185 -292
rect 191 -288 192 -286
rect 191 -294 192 -292
rect 201 -288 202 -286
rect 205 -288 206 -286
rect 205 -294 206 -292
rect 212 -288 213 -286
rect 212 -294 213 -292
rect 219 -288 220 -286
rect 219 -294 220 -292
rect 226 -288 227 -286
rect 226 -294 227 -292
rect 233 -288 234 -286
rect 233 -294 234 -292
rect 240 -288 241 -286
rect 240 -294 241 -292
rect 247 -294 248 -292
rect 250 -294 251 -292
rect 254 -288 255 -286
rect 254 -294 255 -292
rect 261 -288 262 -286
rect 261 -294 262 -292
rect 271 -288 272 -286
rect 271 -294 272 -292
rect 275 -288 276 -286
rect 275 -294 276 -292
rect 2 -325 3 -323
rect 5 -325 6 -323
rect 9 -325 10 -323
rect 9 -331 10 -329
rect 16 -325 17 -323
rect 16 -331 17 -329
rect 23 -325 24 -323
rect 23 -331 24 -329
rect 30 -325 31 -323
rect 30 -331 31 -329
rect 37 -325 38 -323
rect 40 -325 41 -323
rect 40 -331 41 -329
rect 47 -325 48 -323
rect 44 -331 45 -329
rect 51 -325 52 -323
rect 51 -331 52 -329
rect 58 -325 59 -323
rect 58 -331 59 -329
rect 65 -325 66 -323
rect 65 -331 66 -329
rect 75 -325 76 -323
rect 72 -331 73 -329
rect 75 -331 76 -329
rect 79 -325 80 -323
rect 79 -331 80 -329
rect 89 -325 90 -323
rect 86 -331 87 -329
rect 93 -325 94 -323
rect 93 -331 94 -329
rect 96 -331 97 -329
rect 100 -325 101 -323
rect 103 -325 104 -323
rect 100 -331 101 -329
rect 103 -331 104 -329
rect 107 -325 108 -323
rect 107 -331 108 -329
rect 114 -325 115 -323
rect 117 -325 118 -323
rect 114 -331 115 -329
rect 117 -331 118 -329
rect 121 -325 122 -323
rect 121 -331 122 -329
rect 128 -325 129 -323
rect 131 -325 132 -323
rect 128 -331 129 -329
rect 131 -331 132 -329
rect 135 -325 136 -323
rect 135 -331 136 -329
rect 142 -325 143 -323
rect 145 -325 146 -323
rect 149 -325 150 -323
rect 149 -331 150 -329
rect 156 -325 157 -323
rect 156 -331 157 -329
rect 163 -325 164 -323
rect 163 -331 164 -329
rect 170 -325 171 -323
rect 170 -331 171 -329
rect 177 -325 178 -323
rect 177 -331 178 -329
rect 184 -325 185 -323
rect 184 -331 185 -329
rect 191 -325 192 -323
rect 191 -331 192 -329
rect 198 -325 199 -323
rect 198 -331 199 -329
rect 205 -325 206 -323
rect 205 -331 206 -329
rect 212 -325 213 -323
rect 212 -331 213 -329
rect 222 -325 223 -323
rect 219 -331 220 -329
rect 226 -325 227 -323
rect 226 -331 227 -329
rect 2 -356 3 -354
rect 23 -356 24 -354
rect 23 -362 24 -360
rect 30 -356 31 -354
rect 30 -362 31 -360
rect 37 -356 38 -354
rect 37 -362 38 -360
rect 44 -356 45 -354
rect 51 -356 52 -354
rect 58 -356 59 -354
rect 61 -356 62 -354
rect 58 -362 59 -360
rect 68 -356 69 -354
rect 68 -362 69 -360
rect 72 -356 73 -354
rect 72 -362 73 -360
rect 79 -356 80 -354
rect 79 -362 80 -360
rect 86 -362 87 -360
rect 96 -356 97 -354
rect 96 -362 97 -360
rect 100 -356 101 -354
rect 100 -362 101 -360
rect 107 -356 108 -354
rect 107 -362 108 -360
rect 114 -356 115 -354
rect 114 -362 115 -360
rect 117 -362 118 -360
rect 121 -356 122 -354
rect 121 -362 122 -360
rect 128 -356 129 -354
rect 128 -362 129 -360
rect 135 -356 136 -354
rect 135 -362 136 -360
rect 142 -356 143 -354
rect 142 -362 143 -360
rect 149 -356 150 -354
rect 149 -362 150 -360
rect 159 -356 160 -354
rect 156 -362 157 -360
rect 159 -362 160 -360
rect 163 -356 164 -354
rect 163 -362 164 -360
rect 170 -356 171 -354
rect 170 -362 171 -360
rect 177 -356 178 -354
rect 177 -362 178 -360
rect 184 -356 185 -354
rect 184 -362 185 -360
rect 191 -356 192 -354
rect 191 -362 192 -360
rect 198 -356 199 -354
rect 198 -362 199 -360
rect 208 -362 209 -360
rect 215 -356 216 -354
rect 212 -362 213 -360
rect 12 -389 13 -387
rect 16 -389 17 -387
rect 16 -395 17 -393
rect 23 -389 24 -387
rect 23 -395 24 -393
rect 30 -389 31 -387
rect 30 -395 31 -393
rect 37 -395 38 -393
rect 40 -395 41 -393
rect 44 -389 45 -387
rect 47 -389 48 -387
rect 51 -389 52 -387
rect 54 -395 55 -393
rect 58 -389 59 -387
rect 58 -395 59 -393
rect 65 -389 66 -387
rect 65 -395 66 -393
rect 72 -389 73 -387
rect 72 -395 73 -393
rect 79 -389 80 -387
rect 79 -395 80 -393
rect 86 -395 87 -393
rect 89 -395 90 -393
rect 96 -389 97 -387
rect 96 -395 97 -393
rect 100 -389 101 -387
rect 100 -395 101 -393
rect 107 -389 108 -387
rect 110 -395 111 -393
rect 114 -389 115 -387
rect 114 -395 115 -393
rect 117 -395 118 -393
rect 121 -389 122 -387
rect 121 -395 122 -393
rect 128 -395 129 -393
rect 131 -395 132 -393
rect 138 -389 139 -387
rect 138 -395 139 -393
rect 142 -389 143 -387
rect 142 -395 143 -393
rect 152 -395 153 -393
rect 156 -389 157 -387
rect 156 -395 157 -393
rect 163 -389 164 -387
rect 163 -395 164 -393
rect 170 -389 171 -387
rect 170 -395 171 -393
rect 177 -389 178 -387
rect 177 -395 178 -393
rect 184 -389 185 -387
rect 184 -395 185 -393
rect 187 -395 188 -393
rect 191 -389 192 -387
rect 191 -395 192 -393
rect 198 -395 199 -393
rect 205 -389 206 -387
rect 205 -395 206 -393
rect 212 -389 213 -387
rect 212 -395 213 -393
rect 222 -389 223 -387
rect 226 -389 227 -387
rect 226 -395 227 -393
rect 12 -428 13 -426
rect 19 -428 20 -426
rect 26 -422 27 -420
rect 30 -422 31 -420
rect 30 -428 31 -426
rect 44 -422 45 -420
rect 47 -428 48 -426
rect 54 -422 55 -420
rect 61 -422 62 -420
rect 61 -428 62 -426
rect 65 -422 66 -420
rect 65 -428 66 -426
rect 72 -428 73 -426
rect 75 -428 76 -426
rect 79 -422 80 -420
rect 82 -422 83 -420
rect 79 -428 80 -426
rect 89 -428 90 -426
rect 93 -422 94 -420
rect 96 -422 97 -420
rect 96 -428 97 -426
rect 100 -422 101 -420
rect 100 -428 101 -426
rect 107 -422 108 -420
rect 107 -428 108 -426
rect 114 -422 115 -420
rect 114 -428 115 -426
rect 121 -428 122 -426
rect 124 -428 125 -426
rect 128 -422 129 -420
rect 128 -428 129 -426
rect 135 -422 136 -420
rect 142 -422 143 -420
rect 142 -428 143 -426
rect 149 -422 150 -420
rect 149 -428 150 -426
rect 156 -422 157 -420
rect 156 -428 157 -426
rect 187 -422 188 -420
rect 198 -422 199 -420
<< metal1 >>
rect 72 0 80 1
rect 100 0 108 1
rect 121 0 129 1
rect 51 -11 62 -10
rect 68 -11 73 -10
rect 75 -11 80 -10
rect 82 -11 122 -10
rect 44 -13 80 -12
rect 86 -13 118 -12
rect 96 -15 136 -14
rect 100 -17 111 -16
rect 107 -19 143 -18
rect 107 -21 115 -20
rect 44 -32 76 -31
rect 93 -32 143 -31
rect 159 -32 164 -31
rect 247 -32 265 -31
rect 44 -34 62 -33
rect 86 -34 94 -33
rect 107 -34 122 -33
rect 128 -34 143 -33
rect 51 -36 66 -35
rect 86 -36 178 -35
rect 51 -38 59 -37
rect 100 -38 129 -37
rect 131 -38 171 -37
rect 72 -40 101 -39
rect 135 -40 150 -39
rect 72 -42 80 -41
rect 135 -42 167 -41
rect 2 -53 62 -52
rect 75 -53 108 -52
rect 121 -53 195 -52
rect 212 -53 230 -52
rect 233 -53 248 -52
rect 23 -55 34 -54
rect 37 -55 41 -54
rect 51 -55 129 -54
rect 135 -55 157 -54
rect 170 -55 199 -54
rect 233 -55 237 -54
rect 30 -57 45 -56
rect 51 -57 80 -56
rect 89 -57 94 -56
rect 96 -57 108 -56
rect 135 -57 206 -56
rect 44 -59 73 -58
rect 93 -59 115 -58
rect 138 -59 164 -58
rect 177 -59 185 -58
rect 58 -61 101 -60
rect 142 -61 150 -60
rect 152 -61 220 -60
rect 86 -63 143 -62
rect 163 -63 192 -62
rect 58 -65 87 -64
rect 100 -65 118 -64
rect 170 -65 178 -64
rect 2 -76 55 -75
rect 58 -76 115 -75
rect 117 -76 157 -75
rect 173 -76 227 -75
rect 264 -76 283 -75
rect 9 -78 80 -77
rect 86 -78 101 -77
rect 107 -78 146 -77
rect 149 -78 171 -77
rect 184 -78 213 -77
rect 219 -78 248 -77
rect 16 -80 73 -79
rect 100 -80 122 -79
rect 128 -80 136 -79
rect 156 -80 192 -79
rect 198 -80 255 -79
rect 37 -82 69 -81
rect 72 -82 150 -81
rect 177 -82 213 -81
rect 44 -84 97 -83
rect 107 -84 125 -83
rect 128 -84 220 -83
rect 30 -86 45 -85
rect 51 -86 94 -85
rect 131 -86 185 -85
rect 198 -86 234 -85
rect 23 -88 31 -87
rect 51 -88 192 -87
rect 205 -88 241 -87
rect 19 -90 24 -89
rect 58 -90 66 -89
rect 79 -90 206 -89
rect 93 -92 143 -91
rect 163 -92 234 -91
rect 135 -94 178 -93
rect 9 -105 136 -104
rect 149 -105 248 -104
rect 268 -105 283 -104
rect 16 -107 48 -106
rect 58 -107 66 -106
rect 79 -107 115 -106
rect 121 -107 157 -106
rect 163 -107 255 -106
rect 16 -109 24 -108
rect 33 -109 52 -108
rect 58 -109 73 -108
rect 79 -109 108 -108
rect 117 -109 122 -108
rect 124 -109 227 -108
rect 23 -111 31 -110
rect 37 -111 45 -110
rect 65 -111 111 -110
rect 135 -111 171 -110
rect 173 -111 227 -110
rect 9 -113 38 -112
rect 86 -113 115 -112
rect 152 -113 213 -112
rect 68 -115 87 -114
rect 93 -115 101 -114
rect 163 -115 192 -114
rect 208 -115 220 -114
rect 96 -117 129 -116
rect 142 -117 192 -116
rect 219 -117 241 -116
rect 100 -119 262 -118
rect 142 -121 167 -120
rect 177 -121 213 -120
rect 138 -123 178 -122
rect 184 -123 297 -122
rect 187 -125 234 -124
rect 205 -127 234 -126
rect 9 -138 31 -137
rect 40 -138 108 -137
rect 121 -138 153 -137
rect 159 -138 206 -137
rect 212 -138 276 -137
rect 9 -140 94 -139
rect 96 -140 115 -139
rect 117 -140 213 -139
rect 219 -140 269 -139
rect 16 -142 34 -141
rect 44 -142 80 -141
rect 86 -142 108 -141
rect 117 -142 255 -141
rect 16 -144 90 -143
rect 103 -144 129 -143
rect 131 -144 220 -143
rect 226 -144 283 -143
rect 23 -146 38 -145
rect 51 -146 55 -145
rect 72 -146 101 -145
rect 124 -146 262 -145
rect 2 -148 52 -147
rect 72 -148 101 -147
rect 138 -148 248 -147
rect 23 -150 94 -149
rect 138 -150 297 -149
rect 37 -152 129 -151
rect 149 -152 234 -151
rect 79 -154 136 -153
rect 149 -154 157 -153
rect 163 -154 227 -153
rect 86 -156 143 -155
rect 163 -156 199 -155
rect 110 -158 234 -157
rect 114 -160 143 -159
rect 170 -160 209 -159
rect 135 -162 199 -161
rect 177 -164 192 -163
rect 180 -166 241 -165
rect 184 -168 192 -167
rect 65 -170 185 -169
rect 2 -181 118 -180
rect 131 -181 220 -180
rect 222 -181 241 -180
rect 9 -183 129 -182
rect 145 -183 227 -182
rect 16 -185 55 -184
rect 58 -185 115 -184
rect 149 -185 206 -184
rect 219 -185 255 -184
rect 23 -187 69 -186
rect 96 -187 185 -186
rect 191 -187 206 -186
rect 226 -187 276 -186
rect 30 -189 97 -188
rect 100 -189 262 -188
rect 33 -191 38 -190
rect 44 -191 129 -190
rect 142 -191 185 -190
rect 37 -193 73 -192
rect 107 -193 192 -192
rect 44 -195 122 -194
rect 152 -195 269 -194
rect 61 -197 157 -196
rect 166 -197 171 -196
rect 65 -199 90 -198
rect 103 -199 122 -198
rect 152 -199 213 -198
rect 65 -201 87 -200
rect 89 -201 199 -200
rect 86 -203 164 -202
rect 177 -203 199 -202
rect 100 -205 164 -204
rect 177 -205 234 -204
rect 110 -207 283 -206
rect 93 -209 111 -208
rect 114 -209 143 -208
rect 156 -209 248 -208
rect 23 -220 153 -219
rect 173 -220 227 -219
rect 233 -220 241 -219
rect 275 -220 297 -219
rect 16 -222 153 -221
rect 198 -222 227 -221
rect 30 -224 34 -223
rect 37 -224 76 -223
rect 89 -224 136 -223
rect 138 -224 167 -223
rect 184 -224 199 -223
rect 205 -224 248 -223
rect 30 -226 262 -225
rect 37 -228 62 -227
rect 72 -228 87 -227
rect 93 -228 178 -227
rect 184 -228 279 -227
rect 44 -230 52 -229
rect 54 -230 171 -229
rect 212 -230 220 -229
rect 222 -230 269 -229
rect 47 -232 178 -231
rect 191 -232 220 -231
rect 93 -234 111 -233
rect 114 -234 129 -233
rect 131 -234 255 -233
rect 100 -236 115 -235
rect 121 -236 192 -235
rect 61 -238 101 -237
rect 107 -238 157 -237
rect 65 -240 122 -239
rect 135 -240 171 -239
rect 65 -242 80 -241
rect 110 -242 164 -241
rect 9 -244 80 -243
rect 145 -244 206 -243
rect 149 -246 157 -245
rect 9 -257 59 -256
rect 79 -257 202 -256
rect 219 -257 237 -256
rect 240 -257 244 -256
rect 275 -257 297 -256
rect 9 -259 34 -258
rect 44 -259 73 -258
rect 110 -259 129 -258
rect 135 -259 206 -258
rect 219 -259 255 -258
rect 16 -261 87 -260
rect 138 -261 199 -260
rect 240 -261 262 -260
rect 16 -263 90 -262
rect 142 -263 178 -262
rect 243 -263 262 -262
rect 23 -265 87 -264
rect 89 -265 129 -264
rect 135 -265 143 -264
rect 145 -265 213 -264
rect 247 -265 255 -264
rect 23 -267 52 -266
rect 58 -267 66 -266
rect 107 -267 178 -266
rect 26 -269 234 -268
rect 47 -271 80 -270
rect 152 -271 227 -270
rect 51 -273 101 -272
rect 156 -273 206 -272
rect 65 -275 76 -274
rect 93 -275 101 -274
rect 114 -275 157 -274
rect 170 -275 213 -274
rect 114 -277 150 -276
rect 170 -277 272 -276
rect 149 -279 181 -278
rect 191 -279 227 -278
rect 121 -281 192 -280
rect 121 -283 164 -282
rect 37 -285 164 -284
rect 2 -296 6 -295
rect 23 -296 115 -295
rect 121 -296 132 -295
rect 142 -296 213 -295
rect 222 -296 241 -295
rect 247 -296 255 -295
rect 261 -296 272 -295
rect 30 -298 108 -297
rect 142 -298 199 -297
rect 205 -298 213 -297
rect 250 -298 276 -297
rect 16 -300 108 -299
rect 156 -300 178 -299
rect 205 -300 220 -299
rect 37 -302 146 -301
rect 156 -302 192 -301
rect 9 -304 38 -303
rect 40 -304 48 -303
rect 51 -304 118 -303
rect 145 -304 192 -303
rect 2 -306 10 -305
rect 44 -306 97 -305
rect 100 -306 115 -305
rect 177 -306 185 -305
rect 58 -308 80 -307
rect 82 -308 90 -307
rect 93 -308 234 -307
rect 58 -310 129 -309
rect 163 -310 185 -309
rect 16 -312 129 -311
rect 149 -312 164 -311
rect 65 -314 122 -313
rect 65 -316 94 -315
rect 103 -316 150 -315
rect 72 -318 227 -317
rect 75 -320 90 -319
rect 100 -320 227 -319
rect 75 -322 80 -321
rect 2 -333 10 -332
rect 16 -333 69 -332
rect 72 -333 108 -332
rect 114 -333 199 -332
rect 23 -335 87 -334
rect 96 -335 185 -334
rect 198 -335 227 -334
rect 30 -337 104 -336
rect 107 -337 132 -336
rect 135 -337 143 -336
rect 149 -337 171 -336
rect 184 -337 220 -336
rect 30 -339 59 -338
rect 96 -339 129 -338
rect 135 -339 160 -338
rect 170 -339 206 -338
rect 23 -341 59 -340
rect 93 -341 129 -340
rect 156 -341 192 -340
rect 37 -343 118 -342
rect 191 -343 213 -342
rect 40 -345 76 -344
rect 100 -345 122 -344
rect 44 -347 62 -346
rect 79 -347 101 -346
rect 114 -347 150 -346
rect 44 -349 66 -348
rect 121 -349 216 -348
rect 51 -351 73 -350
rect 51 -353 80 -352
rect 12 -364 17 -363
rect 23 -364 45 -363
rect 65 -364 80 -363
rect 86 -364 164 -363
rect 184 -364 209 -363
rect 23 -366 48 -365
rect 114 -366 206 -365
rect 30 -368 59 -367
rect 117 -368 122 -367
rect 138 -368 223 -367
rect 30 -370 52 -369
rect 58 -370 69 -369
rect 121 -370 136 -369
rect 142 -370 164 -369
rect 184 -370 199 -369
rect 37 -372 171 -371
rect 191 -372 213 -371
rect 96 -374 192 -373
rect 79 -376 97 -375
rect 114 -376 171 -375
rect 149 -378 227 -377
rect 156 -380 213 -379
rect 128 -382 157 -381
rect 159 -382 178 -381
rect 107 -384 178 -383
rect 107 -386 143 -385
rect 23 -397 150 -396
rect 152 -397 185 -396
rect 26 -399 129 -398
rect 131 -399 178 -398
rect 30 -401 45 -400
rect 54 -401 59 -400
rect 79 -401 108 -400
rect 110 -401 192 -400
rect 16 -403 31 -402
rect 40 -403 171 -402
rect 54 -405 157 -404
rect 37 -407 157 -406
rect 61 -409 80 -408
rect 82 -409 129 -408
rect 135 -409 188 -408
rect 86 -411 101 -410
rect 117 -411 206 -410
rect 89 -413 97 -412
rect 100 -413 143 -412
rect 187 -413 213 -412
rect 65 -415 97 -414
rect 138 -415 227 -414
rect 65 -417 73 -416
rect 93 -417 115 -416
rect 142 -417 164 -416
rect 114 -419 122 -418
rect 12 -430 129 -429
rect 19 -432 31 -431
rect 47 -432 62 -431
rect 65 -432 76 -431
rect 79 -432 157 -431
rect 72 -434 150 -433
rect 89 -436 108 -435
rect 114 -436 125 -435
rect 96 -438 101 -437
rect 121 -438 143 -437
<< m2contact >>
rect 72 0 73 1
rect 79 0 80 1
rect 100 0 101 1
rect 107 0 108 1
rect 121 0 122 1
rect 128 0 129 1
rect 51 -11 52 -10
rect 61 -11 62 -10
rect 68 -11 69 -10
rect 72 -11 73 -10
rect 75 -11 76 -10
rect 79 -11 80 -10
rect 82 -11 83 -10
rect 121 -11 122 -10
rect 44 -13 45 -12
rect 79 -13 80 -12
rect 86 -13 87 -12
rect 117 -13 118 -12
rect 96 -15 97 -14
rect 135 -15 136 -14
rect 100 -17 101 -16
rect 110 -17 111 -16
rect 107 -19 108 -18
rect 142 -19 143 -18
rect 107 -21 108 -20
rect 114 -21 115 -20
rect 44 -32 45 -31
rect 75 -32 76 -31
rect 93 -32 94 -31
rect 142 -32 143 -31
rect 159 -32 160 -31
rect 163 -32 164 -31
rect 247 -32 248 -31
rect 264 -32 265 -31
rect 44 -34 45 -33
rect 61 -34 62 -33
rect 86 -34 87 -33
rect 93 -34 94 -33
rect 107 -34 108 -33
rect 121 -34 122 -33
rect 128 -34 129 -33
rect 142 -34 143 -33
rect 51 -36 52 -35
rect 65 -36 66 -35
rect 86 -36 87 -35
rect 177 -36 178 -35
rect 51 -38 52 -37
rect 58 -38 59 -37
rect 100 -38 101 -37
rect 128 -38 129 -37
rect 131 -38 132 -37
rect 170 -38 171 -37
rect 72 -40 73 -39
rect 100 -40 101 -39
rect 135 -40 136 -39
rect 149 -40 150 -39
rect 72 -42 73 -41
rect 79 -42 80 -41
rect 135 -42 136 -41
rect 166 -42 167 -41
rect 2 -53 3 -52
rect 61 -53 62 -52
rect 75 -53 76 -52
rect 107 -53 108 -52
rect 121 -53 122 -52
rect 194 -53 195 -52
rect 212 -53 213 -52
rect 229 -53 230 -52
rect 233 -53 234 -52
rect 247 -53 248 -52
rect 23 -55 24 -54
rect 33 -55 34 -54
rect 37 -55 38 -54
rect 40 -55 41 -54
rect 51 -55 52 -54
rect 128 -55 129 -54
rect 135 -55 136 -54
rect 156 -55 157 -54
rect 170 -55 171 -54
rect 198 -55 199 -54
rect 233 -55 234 -54
rect 236 -55 237 -54
rect 30 -57 31 -56
rect 44 -57 45 -56
rect 51 -57 52 -56
rect 79 -57 80 -56
rect 89 -57 90 -56
rect 93 -57 94 -56
rect 96 -57 97 -56
rect 107 -57 108 -56
rect 135 -57 136 -56
rect 205 -57 206 -56
rect 44 -59 45 -58
rect 72 -59 73 -58
rect 93 -59 94 -58
rect 114 -59 115 -58
rect 138 -59 139 -58
rect 163 -59 164 -58
rect 177 -59 178 -58
rect 184 -59 185 -58
rect 58 -61 59 -60
rect 100 -61 101 -60
rect 142 -61 143 -60
rect 149 -61 150 -60
rect 152 -61 153 -60
rect 219 -61 220 -60
rect 86 -63 87 -62
rect 142 -63 143 -62
rect 163 -63 164 -62
rect 191 -63 192 -62
rect 58 -65 59 -64
rect 86 -65 87 -64
rect 100 -65 101 -64
rect 117 -65 118 -64
rect 170 -65 171 -64
rect 177 -65 178 -64
rect 2 -76 3 -75
rect 54 -76 55 -75
rect 58 -76 59 -75
rect 114 -76 115 -75
rect 117 -76 118 -75
rect 156 -76 157 -75
rect 173 -76 174 -75
rect 226 -76 227 -75
rect 264 -76 265 -75
rect 282 -76 283 -75
rect 9 -78 10 -77
rect 79 -78 80 -77
rect 86 -78 87 -77
rect 100 -78 101 -77
rect 107 -78 108 -77
rect 145 -78 146 -77
rect 149 -78 150 -77
rect 170 -78 171 -77
rect 184 -78 185 -77
rect 212 -78 213 -77
rect 219 -78 220 -77
rect 247 -78 248 -77
rect 16 -80 17 -79
rect 72 -80 73 -79
rect 100 -80 101 -79
rect 121 -80 122 -79
rect 128 -80 129 -79
rect 135 -80 136 -79
rect 156 -80 157 -79
rect 191 -80 192 -79
rect 198 -80 199 -79
rect 254 -80 255 -79
rect 37 -82 38 -81
rect 68 -82 69 -81
rect 72 -82 73 -81
rect 149 -82 150 -81
rect 177 -82 178 -81
rect 212 -82 213 -81
rect 44 -84 45 -83
rect 96 -84 97 -83
rect 107 -84 108 -83
rect 124 -84 125 -83
rect 128 -84 129 -83
rect 219 -84 220 -83
rect 30 -86 31 -85
rect 44 -86 45 -85
rect 51 -86 52 -85
rect 93 -86 94 -85
rect 131 -86 132 -85
rect 184 -86 185 -85
rect 198 -86 199 -85
rect 233 -86 234 -85
rect 23 -88 24 -87
rect 30 -88 31 -87
rect 51 -88 52 -87
rect 191 -88 192 -87
rect 205 -88 206 -87
rect 240 -88 241 -87
rect 19 -90 20 -89
rect 23 -90 24 -89
rect 58 -90 59 -89
rect 65 -90 66 -89
rect 79 -90 80 -89
rect 205 -90 206 -89
rect 93 -92 94 -91
rect 142 -92 143 -91
rect 163 -92 164 -91
rect 233 -92 234 -91
rect 135 -94 136 -93
rect 177 -94 178 -93
rect 9 -105 10 -104
rect 135 -105 136 -104
rect 149 -105 150 -104
rect 247 -105 248 -104
rect 268 -105 269 -104
rect 282 -105 283 -104
rect 16 -107 17 -106
rect 47 -107 48 -106
rect 58 -107 59 -106
rect 65 -107 66 -106
rect 79 -107 80 -106
rect 114 -107 115 -106
rect 121 -107 122 -106
rect 156 -107 157 -106
rect 163 -107 164 -106
rect 254 -107 255 -106
rect 16 -109 17 -108
rect 23 -109 24 -108
rect 33 -109 34 -108
rect 51 -109 52 -108
rect 58 -109 59 -108
rect 72 -109 73 -108
rect 79 -109 80 -108
rect 107 -109 108 -108
rect 117 -109 118 -108
rect 121 -109 122 -108
rect 124 -109 125 -108
rect 226 -109 227 -108
rect 23 -111 24 -110
rect 30 -111 31 -110
rect 37 -111 38 -110
rect 44 -111 45 -110
rect 65 -111 66 -110
rect 110 -111 111 -110
rect 135 -111 136 -110
rect 170 -111 171 -110
rect 173 -111 174 -110
rect 226 -111 227 -110
rect 9 -113 10 -112
rect 37 -113 38 -112
rect 86 -113 87 -112
rect 114 -113 115 -112
rect 152 -113 153 -112
rect 212 -113 213 -112
rect 68 -115 69 -114
rect 86 -115 87 -114
rect 93 -115 94 -114
rect 100 -115 101 -114
rect 163 -115 164 -114
rect 191 -115 192 -114
rect 208 -115 209 -114
rect 219 -115 220 -114
rect 96 -117 97 -116
rect 128 -117 129 -116
rect 142 -117 143 -116
rect 191 -117 192 -116
rect 219 -117 220 -116
rect 240 -117 241 -116
rect 100 -119 101 -118
rect 261 -119 262 -118
rect 142 -121 143 -120
rect 166 -121 167 -120
rect 177 -121 178 -120
rect 212 -121 213 -120
rect 138 -123 139 -122
rect 177 -123 178 -122
rect 184 -123 185 -122
rect 296 -123 297 -122
rect 187 -125 188 -124
rect 233 -125 234 -124
rect 205 -127 206 -126
rect 233 -127 234 -126
rect 9 -138 10 -137
rect 30 -138 31 -137
rect 40 -138 41 -137
rect 107 -138 108 -137
rect 121 -138 122 -137
rect 152 -138 153 -137
rect 159 -138 160 -137
rect 205 -138 206 -137
rect 212 -138 213 -137
rect 275 -138 276 -137
rect 9 -140 10 -139
rect 93 -140 94 -139
rect 96 -140 97 -139
rect 114 -140 115 -139
rect 117 -140 118 -139
rect 212 -140 213 -139
rect 219 -140 220 -139
rect 268 -140 269 -139
rect 16 -142 17 -141
rect 33 -142 34 -141
rect 44 -142 45 -141
rect 79 -142 80 -141
rect 86 -142 87 -141
rect 107 -142 108 -141
rect 117 -142 118 -141
rect 254 -142 255 -141
rect 16 -144 17 -143
rect 89 -144 90 -143
rect 103 -144 104 -143
rect 128 -144 129 -143
rect 131 -144 132 -143
rect 219 -144 220 -143
rect 226 -144 227 -143
rect 282 -144 283 -143
rect 23 -146 24 -145
rect 37 -146 38 -145
rect 51 -146 52 -145
rect 54 -146 55 -145
rect 72 -146 73 -145
rect 100 -146 101 -145
rect 124 -146 125 -145
rect 261 -146 262 -145
rect 2 -148 3 -147
rect 51 -148 52 -147
rect 72 -148 73 -147
rect 100 -148 101 -147
rect 138 -148 139 -147
rect 247 -148 248 -147
rect 23 -150 24 -149
rect 93 -150 94 -149
rect 138 -150 139 -149
rect 296 -150 297 -149
rect 37 -152 38 -151
rect 128 -152 129 -151
rect 149 -152 150 -151
rect 233 -152 234 -151
rect 79 -154 80 -153
rect 135 -154 136 -153
rect 149 -154 150 -153
rect 156 -154 157 -153
rect 163 -154 164 -153
rect 226 -154 227 -153
rect 86 -156 87 -155
rect 142 -156 143 -155
rect 163 -156 164 -155
rect 198 -156 199 -155
rect 110 -158 111 -157
rect 233 -158 234 -157
rect 114 -160 115 -159
rect 142 -160 143 -159
rect 170 -160 171 -159
rect 208 -160 209 -159
rect 135 -162 136 -161
rect 198 -162 199 -161
rect 177 -164 178 -163
rect 191 -164 192 -163
rect 180 -166 181 -165
rect 240 -166 241 -165
rect 184 -168 185 -167
rect 191 -168 192 -167
rect 65 -170 66 -169
rect 184 -170 185 -169
rect 2 -181 3 -180
rect 117 -181 118 -180
rect 131 -181 132 -180
rect 219 -181 220 -180
rect 222 -181 223 -180
rect 240 -181 241 -180
rect 9 -183 10 -182
rect 128 -183 129 -182
rect 145 -183 146 -182
rect 226 -183 227 -182
rect 16 -185 17 -184
rect 54 -185 55 -184
rect 58 -185 59 -184
rect 114 -185 115 -184
rect 149 -185 150 -184
rect 205 -185 206 -184
rect 219 -185 220 -184
rect 254 -185 255 -184
rect 23 -187 24 -186
rect 68 -187 69 -186
rect 96 -187 97 -186
rect 184 -187 185 -186
rect 191 -187 192 -186
rect 205 -187 206 -186
rect 226 -187 227 -186
rect 275 -187 276 -186
rect 30 -189 31 -188
rect 96 -189 97 -188
rect 100 -189 101 -188
rect 261 -189 262 -188
rect 33 -191 34 -190
rect 37 -191 38 -190
rect 44 -191 45 -190
rect 128 -191 129 -190
rect 142 -191 143 -190
rect 184 -191 185 -190
rect 37 -193 38 -192
rect 72 -193 73 -192
rect 107 -193 108 -192
rect 191 -193 192 -192
rect 44 -195 45 -194
rect 121 -195 122 -194
rect 152 -195 153 -194
rect 268 -195 269 -194
rect 61 -197 62 -196
rect 156 -197 157 -196
rect 166 -197 167 -196
rect 170 -197 171 -196
rect 65 -199 66 -198
rect 89 -199 90 -198
rect 103 -199 104 -198
rect 121 -199 122 -198
rect 152 -199 153 -198
rect 212 -199 213 -198
rect 65 -201 66 -200
rect 86 -201 87 -200
rect 89 -201 90 -200
rect 198 -201 199 -200
rect 86 -203 87 -202
rect 163 -203 164 -202
rect 177 -203 178 -202
rect 198 -203 199 -202
rect 100 -205 101 -204
rect 163 -205 164 -204
rect 177 -205 178 -204
rect 233 -205 234 -204
rect 110 -207 111 -206
rect 282 -207 283 -206
rect 93 -209 94 -208
rect 110 -209 111 -208
rect 114 -209 115 -208
rect 142 -209 143 -208
rect 156 -209 157 -208
rect 247 -209 248 -208
rect 23 -220 24 -219
rect 152 -220 153 -219
rect 173 -220 174 -219
rect 226 -220 227 -219
rect 233 -220 234 -219
rect 240 -220 241 -219
rect 275 -220 276 -219
rect 296 -220 297 -219
rect 16 -222 17 -221
rect 152 -222 153 -221
rect 198 -222 199 -221
rect 226 -222 227 -221
rect 30 -224 31 -223
rect 33 -224 34 -223
rect 37 -224 38 -223
rect 75 -224 76 -223
rect 89 -224 90 -223
rect 135 -224 136 -223
rect 138 -224 139 -223
rect 166 -224 167 -223
rect 184 -224 185 -223
rect 198 -224 199 -223
rect 205 -224 206 -223
rect 247 -224 248 -223
rect 30 -226 31 -225
rect 261 -226 262 -225
rect 37 -228 38 -227
rect 61 -228 62 -227
rect 72 -228 73 -227
rect 86 -228 87 -227
rect 93 -228 94 -227
rect 177 -228 178 -227
rect 184 -228 185 -227
rect 278 -228 279 -227
rect 44 -230 45 -229
rect 51 -230 52 -229
rect 54 -230 55 -229
rect 170 -230 171 -229
rect 212 -230 213 -229
rect 219 -230 220 -229
rect 222 -230 223 -229
rect 268 -230 269 -229
rect 47 -232 48 -231
rect 177 -232 178 -231
rect 191 -232 192 -231
rect 219 -232 220 -231
rect 93 -234 94 -233
rect 110 -234 111 -233
rect 114 -234 115 -233
rect 128 -234 129 -233
rect 131 -234 132 -233
rect 254 -234 255 -233
rect 100 -236 101 -235
rect 114 -236 115 -235
rect 121 -236 122 -235
rect 191 -236 192 -235
rect 61 -238 62 -237
rect 100 -238 101 -237
rect 107 -238 108 -237
rect 156 -238 157 -237
rect 65 -240 66 -239
rect 121 -240 122 -239
rect 135 -240 136 -239
rect 170 -240 171 -239
rect 65 -242 66 -241
rect 79 -242 80 -241
rect 110 -242 111 -241
rect 163 -242 164 -241
rect 9 -244 10 -243
rect 79 -244 80 -243
rect 145 -244 146 -243
rect 205 -244 206 -243
rect 149 -246 150 -245
rect 156 -246 157 -245
rect 9 -257 10 -256
rect 58 -257 59 -256
rect 79 -257 80 -256
rect 201 -257 202 -256
rect 219 -257 220 -256
rect 236 -257 237 -256
rect 240 -257 241 -256
rect 243 -257 244 -256
rect 275 -257 276 -256
rect 296 -257 297 -256
rect 9 -259 10 -258
rect 33 -259 34 -258
rect 44 -259 45 -258
rect 72 -259 73 -258
rect 110 -259 111 -258
rect 128 -259 129 -258
rect 135 -259 136 -258
rect 205 -259 206 -258
rect 219 -259 220 -258
rect 254 -259 255 -258
rect 16 -261 17 -260
rect 86 -261 87 -260
rect 138 -261 139 -260
rect 198 -261 199 -260
rect 240 -261 241 -260
rect 261 -261 262 -260
rect 16 -263 17 -262
rect 89 -263 90 -262
rect 142 -263 143 -262
rect 177 -263 178 -262
rect 243 -263 244 -262
rect 261 -263 262 -262
rect 23 -265 24 -264
rect 86 -265 87 -264
rect 89 -265 90 -264
rect 128 -265 129 -264
rect 135 -265 136 -264
rect 142 -265 143 -264
rect 145 -265 146 -264
rect 212 -265 213 -264
rect 247 -265 248 -264
rect 254 -265 255 -264
rect 23 -267 24 -266
rect 51 -267 52 -266
rect 58 -267 59 -266
rect 65 -267 66 -266
rect 107 -267 108 -266
rect 177 -267 178 -266
rect 26 -269 27 -268
rect 233 -269 234 -268
rect 47 -271 48 -270
rect 79 -271 80 -270
rect 152 -271 153 -270
rect 226 -271 227 -270
rect 51 -273 52 -272
rect 100 -273 101 -272
rect 156 -273 157 -272
rect 205 -273 206 -272
rect 65 -275 66 -274
rect 75 -275 76 -274
rect 93 -275 94 -274
rect 100 -275 101 -274
rect 114 -275 115 -274
rect 156 -275 157 -274
rect 170 -275 171 -274
rect 212 -275 213 -274
rect 114 -277 115 -276
rect 149 -277 150 -276
rect 170 -277 171 -276
rect 271 -277 272 -276
rect 149 -279 150 -278
rect 180 -279 181 -278
rect 191 -279 192 -278
rect 226 -279 227 -278
rect 121 -281 122 -280
rect 191 -281 192 -280
rect 121 -283 122 -282
rect 163 -283 164 -282
rect 37 -285 38 -284
rect 163 -285 164 -284
rect 2 -296 3 -295
rect 5 -296 6 -295
rect 23 -296 24 -295
rect 114 -296 115 -295
rect 121 -296 122 -295
rect 131 -296 132 -295
rect 142 -296 143 -295
rect 212 -296 213 -295
rect 222 -296 223 -295
rect 240 -296 241 -295
rect 247 -296 248 -295
rect 254 -296 255 -295
rect 261 -296 262 -295
rect 271 -296 272 -295
rect 30 -298 31 -297
rect 107 -298 108 -297
rect 142 -298 143 -297
rect 198 -298 199 -297
rect 205 -298 206 -297
rect 212 -298 213 -297
rect 250 -298 251 -297
rect 275 -298 276 -297
rect 16 -300 17 -299
rect 107 -300 108 -299
rect 156 -300 157 -299
rect 177 -300 178 -299
rect 205 -300 206 -299
rect 219 -300 220 -299
rect 37 -302 38 -301
rect 145 -302 146 -301
rect 156 -302 157 -301
rect 191 -302 192 -301
rect 9 -304 10 -303
rect 37 -304 38 -303
rect 40 -304 41 -303
rect 47 -304 48 -303
rect 51 -304 52 -303
rect 117 -304 118 -303
rect 145 -304 146 -303
rect 191 -304 192 -303
rect 2 -306 3 -305
rect 9 -306 10 -305
rect 44 -306 45 -305
rect 96 -306 97 -305
rect 100 -306 101 -305
rect 114 -306 115 -305
rect 177 -306 178 -305
rect 184 -306 185 -305
rect 58 -308 59 -307
rect 79 -308 80 -307
rect 82 -308 83 -307
rect 89 -308 90 -307
rect 93 -308 94 -307
rect 233 -308 234 -307
rect 58 -310 59 -309
rect 128 -310 129 -309
rect 163 -310 164 -309
rect 184 -310 185 -309
rect 16 -312 17 -311
rect 128 -312 129 -311
rect 149 -312 150 -311
rect 163 -312 164 -311
rect 65 -314 66 -313
rect 121 -314 122 -313
rect 65 -316 66 -315
rect 93 -316 94 -315
rect 103 -316 104 -315
rect 149 -316 150 -315
rect 72 -318 73 -317
rect 226 -318 227 -317
rect 75 -320 76 -319
rect 89 -320 90 -319
rect 100 -320 101 -319
rect 226 -320 227 -319
rect 75 -322 76 -321
rect 79 -322 80 -321
rect 2 -333 3 -332
rect 9 -333 10 -332
rect 16 -333 17 -332
rect 68 -333 69 -332
rect 72 -333 73 -332
rect 107 -333 108 -332
rect 114 -333 115 -332
rect 198 -333 199 -332
rect 23 -335 24 -334
rect 86 -335 87 -334
rect 96 -335 97 -334
rect 184 -335 185 -334
rect 198 -335 199 -334
rect 226 -335 227 -334
rect 30 -337 31 -336
rect 103 -337 104 -336
rect 107 -337 108 -336
rect 131 -337 132 -336
rect 135 -337 136 -336
rect 142 -337 143 -336
rect 149 -337 150 -336
rect 170 -337 171 -336
rect 184 -337 185 -336
rect 219 -337 220 -336
rect 30 -339 31 -338
rect 58 -339 59 -338
rect 96 -339 97 -338
rect 128 -339 129 -338
rect 135 -339 136 -338
rect 159 -339 160 -338
rect 170 -339 171 -338
rect 205 -339 206 -338
rect 23 -341 24 -340
rect 58 -341 59 -340
rect 93 -341 94 -340
rect 128 -341 129 -340
rect 156 -341 157 -340
rect 191 -341 192 -340
rect 37 -343 38 -342
rect 117 -343 118 -342
rect 191 -343 192 -342
rect 212 -343 213 -342
rect 40 -345 41 -344
rect 75 -345 76 -344
rect 100 -345 101 -344
rect 121 -345 122 -344
rect 44 -347 45 -346
rect 61 -347 62 -346
rect 79 -347 80 -346
rect 100 -347 101 -346
rect 114 -347 115 -346
rect 149 -347 150 -346
rect 44 -349 45 -348
rect 65 -349 66 -348
rect 121 -349 122 -348
rect 215 -349 216 -348
rect 51 -351 52 -350
rect 72 -351 73 -350
rect 51 -353 52 -352
rect 79 -353 80 -352
rect 12 -364 13 -363
rect 16 -364 17 -363
rect 23 -364 24 -363
rect 44 -364 45 -363
rect 65 -364 66 -363
rect 79 -364 80 -363
rect 86 -364 87 -363
rect 163 -364 164 -363
rect 184 -364 185 -363
rect 208 -364 209 -363
rect 23 -366 24 -365
rect 47 -366 48 -365
rect 114 -366 115 -365
rect 205 -366 206 -365
rect 30 -368 31 -367
rect 58 -368 59 -367
rect 117 -368 118 -367
rect 121 -368 122 -367
rect 138 -368 139 -367
rect 222 -368 223 -367
rect 30 -370 31 -369
rect 51 -370 52 -369
rect 58 -370 59 -369
rect 68 -370 69 -369
rect 121 -370 122 -369
rect 135 -370 136 -369
rect 142 -370 143 -369
rect 163 -370 164 -369
rect 184 -370 185 -369
rect 198 -370 199 -369
rect 37 -372 38 -371
rect 170 -372 171 -371
rect 191 -372 192 -371
rect 212 -372 213 -371
rect 96 -374 97 -373
rect 191 -374 192 -373
rect 79 -376 80 -375
rect 96 -376 97 -375
rect 114 -376 115 -375
rect 170 -376 171 -375
rect 149 -378 150 -377
rect 226 -378 227 -377
rect 156 -380 157 -379
rect 212 -380 213 -379
rect 128 -382 129 -381
rect 156 -382 157 -381
rect 159 -382 160 -381
rect 177 -382 178 -381
rect 107 -384 108 -383
rect 177 -384 178 -383
rect 107 -386 108 -385
rect 142 -386 143 -385
rect 23 -397 24 -396
rect 149 -397 150 -396
rect 152 -397 153 -396
rect 184 -397 185 -396
rect 26 -399 27 -398
rect 128 -399 129 -398
rect 131 -399 132 -398
rect 177 -399 178 -398
rect 30 -401 31 -400
rect 44 -401 45 -400
rect 54 -401 55 -400
rect 58 -401 59 -400
rect 79 -401 80 -400
rect 107 -401 108 -400
rect 110 -401 111 -400
rect 191 -401 192 -400
rect 16 -403 17 -402
rect 30 -403 31 -402
rect 40 -403 41 -402
rect 170 -403 171 -402
rect 54 -405 55 -404
rect 156 -405 157 -404
rect 37 -407 38 -406
rect 156 -407 157 -406
rect 61 -409 62 -408
rect 79 -409 80 -408
rect 82 -409 83 -408
rect 128 -409 129 -408
rect 135 -409 136 -408
rect 187 -409 188 -408
rect 86 -411 87 -410
rect 100 -411 101 -410
rect 117 -411 118 -410
rect 205 -411 206 -410
rect 89 -413 90 -412
rect 96 -413 97 -412
rect 100 -413 101 -412
rect 142 -413 143 -412
rect 187 -413 188 -412
rect 212 -413 213 -412
rect 65 -415 66 -414
rect 96 -415 97 -414
rect 138 -415 139 -414
rect 226 -415 227 -414
rect 65 -417 66 -416
rect 72 -417 73 -416
rect 93 -417 94 -416
rect 114 -417 115 -416
rect 142 -417 143 -416
rect 163 -417 164 -416
rect 114 -419 115 -418
rect 121 -419 122 -418
rect 12 -430 13 -429
rect 128 -430 129 -429
rect 19 -432 20 -431
rect 30 -432 31 -431
rect 47 -432 48 -431
rect 61 -432 62 -431
rect 65 -432 66 -431
rect 75 -432 76 -431
rect 79 -432 80 -431
rect 156 -432 157 -431
rect 72 -434 73 -433
rect 149 -434 150 -433
rect 89 -436 90 -435
rect 107 -436 108 -435
rect 114 -436 115 -435
rect 124 -436 125 -435
rect 96 -438 97 -437
rect 100 -438 101 -437
rect 121 -438 122 -437
rect 142 -438 143 -437
<< metal2 >>
rect 72 -1 73 1
rect 79 -1 80 1
rect 100 -1 101 1
rect 107 -1 108 1
rect 121 -1 122 1
rect 128 -1 129 1
rect 51 -22 52 -10
rect 61 -22 62 -10
rect 68 -22 69 -10
rect 72 -22 73 -10
rect 75 -11 76 -9
rect 79 -11 80 -9
rect 82 -22 83 -10
rect 121 -22 122 -10
rect 128 -11 129 -9
rect 128 -22 129 -10
rect 128 -11 129 -9
rect 128 -22 129 -10
rect 44 -22 45 -12
rect 79 -22 80 -12
rect 86 -22 87 -12
rect 117 -22 118 -12
rect 96 -22 97 -14
rect 135 -22 136 -14
rect 100 -22 101 -16
rect 110 -22 111 -16
rect 107 -19 108 -9
rect 142 -22 143 -18
rect 107 -22 108 -20
rect 114 -21 115 -9
rect 44 -32 45 -30
rect 75 -43 76 -31
rect 93 -32 94 -30
rect 142 -32 143 -30
rect 159 -32 160 -30
rect 163 -43 164 -31
rect 247 -43 248 -31
rect 264 -32 265 -30
rect 44 -43 45 -33
rect 61 -43 62 -33
rect 86 -34 87 -30
rect 93 -43 94 -33
rect 107 -43 108 -33
rect 121 -34 122 -30
rect 128 -34 129 -30
rect 142 -43 143 -33
rect 51 -36 52 -30
rect 65 -43 66 -35
rect 86 -43 87 -35
rect 177 -43 178 -35
rect 51 -43 52 -37
rect 58 -43 59 -37
rect 100 -38 101 -30
rect 128 -43 129 -37
rect 131 -43 132 -37
rect 170 -43 171 -37
rect 72 -40 73 -30
rect 100 -43 101 -39
rect 135 -40 136 -30
rect 149 -43 150 -39
rect 72 -43 73 -41
rect 79 -43 80 -41
rect 135 -43 136 -41
rect 166 -43 167 -41
rect 2 -66 3 -52
rect 61 -53 62 -51
rect 65 -53 66 -51
rect 65 -66 66 -52
rect 65 -53 66 -51
rect 65 -66 66 -52
rect 75 -66 76 -52
rect 107 -53 108 -51
rect 121 -66 122 -52
rect 194 -66 195 -52
rect 212 -66 213 -52
rect 229 -66 230 -52
rect 233 -53 234 -51
rect 247 -53 248 -51
rect 23 -66 24 -54
rect 33 -66 34 -54
rect 37 -66 38 -54
rect 40 -55 41 -51
rect 51 -55 52 -51
rect 128 -66 129 -54
rect 135 -55 136 -51
rect 156 -66 157 -54
rect 170 -55 171 -51
rect 198 -66 199 -54
rect 233 -66 234 -54
rect 236 -55 237 -51
rect 30 -57 31 -51
rect 44 -57 45 -51
rect 51 -66 52 -56
rect 79 -57 80 -51
rect 89 -57 90 -51
rect 93 -57 94 -51
rect 96 -66 97 -56
rect 107 -66 108 -56
rect 135 -66 136 -56
rect 205 -66 206 -56
rect 44 -66 45 -58
rect 72 -66 73 -58
rect 93 -66 94 -58
rect 114 -59 115 -51
rect 138 -66 139 -58
rect 163 -59 164 -51
rect 177 -59 178 -51
rect 184 -66 185 -58
rect 58 -61 59 -51
rect 100 -61 101 -51
rect 142 -61 143 -51
rect 149 -66 150 -60
rect 152 -61 153 -51
rect 219 -66 220 -60
rect 86 -63 87 -51
rect 142 -66 143 -62
rect 163 -66 164 -62
rect 191 -66 192 -62
rect 58 -66 59 -64
rect 86 -66 87 -64
rect 100 -66 101 -64
rect 117 -66 118 -64
rect 170 -66 171 -64
rect 177 -66 178 -64
rect 2 -76 3 -74
rect 54 -95 55 -75
rect 58 -76 59 -74
rect 114 -95 115 -75
rect 117 -76 118 -74
rect 156 -76 157 -74
rect 173 -76 174 -74
rect 226 -95 227 -75
rect 264 -95 265 -75
rect 282 -95 283 -75
rect 9 -95 10 -77
rect 79 -78 80 -74
rect 86 -95 87 -77
rect 100 -78 101 -74
rect 107 -78 108 -74
rect 145 -95 146 -77
rect 149 -78 150 -74
rect 170 -95 171 -77
rect 184 -78 185 -74
rect 212 -78 213 -74
rect 219 -78 220 -74
rect 247 -95 248 -77
rect 16 -95 17 -79
rect 72 -80 73 -74
rect 100 -95 101 -79
rect 121 -80 122 -74
rect 128 -80 129 -74
rect 135 -80 136 -74
rect 156 -95 157 -79
rect 191 -80 192 -74
rect 198 -80 199 -74
rect 254 -95 255 -79
rect 37 -95 38 -81
rect 68 -95 69 -81
rect 72 -95 73 -81
rect 149 -95 150 -81
rect 177 -82 178 -74
rect 212 -95 213 -81
rect 44 -84 45 -74
rect 96 -95 97 -83
rect 107 -95 108 -83
rect 124 -95 125 -83
rect 128 -95 129 -83
rect 219 -95 220 -83
rect 30 -86 31 -74
rect 44 -95 45 -85
rect 51 -86 52 -74
rect 93 -86 94 -74
rect 131 -95 132 -85
rect 184 -95 185 -85
rect 198 -95 199 -85
rect 233 -86 234 -74
rect 23 -88 24 -74
rect 30 -95 31 -87
rect 51 -95 52 -87
rect 191 -95 192 -87
rect 205 -88 206 -74
rect 240 -95 241 -87
rect 19 -90 20 -74
rect 23 -95 24 -89
rect 58 -95 59 -89
rect 65 -90 66 -74
rect 79 -95 80 -89
rect 205 -95 206 -89
rect 93 -95 94 -91
rect 142 -92 143 -74
rect 163 -92 164 -74
rect 233 -95 234 -91
rect 135 -95 136 -93
rect 177 -95 178 -93
rect 9 -105 10 -103
rect 135 -105 136 -103
rect 149 -105 150 -103
rect 247 -105 248 -103
rect 268 -105 269 -103
rect 282 -105 283 -103
rect 16 -107 17 -103
rect 47 -128 48 -106
rect 58 -107 59 -103
rect 65 -107 66 -103
rect 79 -107 80 -103
rect 114 -107 115 -103
rect 121 -107 122 -103
rect 156 -107 157 -103
rect 163 -107 164 -103
rect 254 -107 255 -103
rect 16 -128 17 -108
rect 23 -109 24 -103
rect 33 -128 34 -108
rect 51 -128 52 -108
rect 58 -128 59 -108
rect 72 -109 73 -103
rect 79 -128 80 -108
rect 107 -109 108 -103
rect 117 -128 118 -108
rect 121 -128 122 -108
rect 124 -109 125 -103
rect 226 -109 227 -103
rect 23 -128 24 -110
rect 30 -111 31 -103
rect 37 -111 38 -103
rect 44 -111 45 -103
rect 65 -128 66 -110
rect 110 -128 111 -110
rect 135 -128 136 -110
rect 170 -111 171 -103
rect 173 -128 174 -110
rect 226 -128 227 -110
rect 9 -128 10 -112
rect 37 -128 38 -112
rect 86 -113 87 -103
rect 114 -128 115 -112
rect 152 -113 153 -103
rect 212 -113 213 -103
rect 68 -115 69 -103
rect 86 -128 87 -114
rect 93 -128 94 -114
rect 100 -115 101 -103
rect 163 -128 164 -114
rect 191 -115 192 -103
rect 198 -115 199 -103
rect 198 -128 199 -114
rect 198 -115 199 -103
rect 198 -128 199 -114
rect 208 -128 209 -114
rect 219 -115 220 -103
rect 96 -117 97 -103
rect 128 -128 129 -116
rect 142 -117 143 -103
rect 191 -128 192 -116
rect 219 -128 220 -116
rect 240 -117 241 -103
rect 100 -128 101 -118
rect 261 -119 262 -103
rect 142 -128 143 -120
rect 166 -121 167 -103
rect 177 -121 178 -103
rect 212 -128 213 -120
rect 138 -123 139 -103
rect 177 -128 178 -122
rect 184 -123 185 -103
rect 296 -128 297 -122
rect 187 -128 188 -124
rect 233 -125 234 -103
rect 205 -127 206 -103
rect 233 -128 234 -126
rect 9 -138 10 -136
rect 30 -138 31 -136
rect 40 -138 41 -136
rect 107 -138 108 -136
rect 121 -138 122 -136
rect 152 -171 153 -137
rect 159 -138 160 -136
rect 205 -171 206 -137
rect 212 -138 213 -136
rect 275 -171 276 -137
rect 9 -171 10 -139
rect 93 -140 94 -136
rect 96 -140 97 -136
rect 114 -140 115 -136
rect 117 -140 118 -136
rect 212 -171 213 -139
rect 219 -140 220 -136
rect 268 -171 269 -139
rect 16 -142 17 -136
rect 33 -142 34 -136
rect 44 -171 45 -141
rect 79 -142 80 -136
rect 86 -142 87 -136
rect 107 -171 108 -141
rect 117 -171 118 -141
rect 254 -171 255 -141
rect 16 -171 17 -143
rect 89 -171 90 -143
rect 103 -171 104 -143
rect 128 -144 129 -136
rect 131 -171 132 -143
rect 219 -171 220 -143
rect 226 -144 227 -136
rect 282 -171 283 -143
rect 23 -146 24 -136
rect 37 -146 38 -136
rect 51 -146 52 -136
rect 54 -171 55 -145
rect 58 -146 59 -136
rect 58 -171 59 -145
rect 58 -146 59 -136
rect 58 -171 59 -145
rect 72 -146 73 -136
rect 100 -146 101 -136
rect 124 -171 125 -145
rect 261 -171 262 -145
rect 2 -171 3 -147
rect 51 -171 52 -147
rect 72 -171 73 -147
rect 100 -171 101 -147
rect 138 -148 139 -136
rect 247 -171 248 -147
rect 23 -171 24 -149
rect 93 -171 94 -149
rect 138 -171 139 -149
rect 296 -150 297 -136
rect 37 -171 38 -151
rect 128 -171 129 -151
rect 149 -152 150 -136
rect 233 -152 234 -136
rect 79 -171 80 -153
rect 135 -154 136 -136
rect 149 -171 150 -153
rect 156 -171 157 -153
rect 163 -154 164 -136
rect 226 -171 227 -153
rect 86 -171 87 -155
rect 142 -156 143 -136
rect 163 -171 164 -155
rect 198 -156 199 -136
rect 110 -158 111 -136
rect 233 -171 234 -157
rect 114 -171 115 -159
rect 142 -171 143 -159
rect 170 -171 171 -159
rect 208 -160 209 -136
rect 135 -171 136 -161
rect 198 -171 199 -161
rect 177 -171 178 -163
rect 191 -164 192 -136
rect 180 -166 181 -136
rect 240 -171 241 -165
rect 184 -168 185 -136
rect 191 -171 192 -167
rect 65 -170 66 -136
rect 184 -171 185 -169
rect 2 -181 3 -179
rect 117 -181 118 -179
rect 131 -181 132 -179
rect 219 -181 220 -179
rect 222 -210 223 -180
rect 240 -181 241 -179
rect 9 -183 10 -179
rect 128 -183 129 -179
rect 135 -183 136 -179
rect 135 -210 136 -182
rect 135 -183 136 -179
rect 135 -210 136 -182
rect 145 -210 146 -182
rect 226 -183 227 -179
rect 16 -185 17 -179
rect 54 -210 55 -184
rect 58 -185 59 -179
rect 114 -185 115 -179
rect 149 -210 150 -184
rect 205 -185 206 -179
rect 219 -210 220 -184
rect 254 -185 255 -179
rect 23 -187 24 -179
rect 68 -187 69 -179
rect 79 -187 80 -179
rect 79 -210 80 -186
rect 79 -187 80 -179
rect 79 -210 80 -186
rect 96 -187 97 -179
rect 184 -187 185 -179
rect 191 -187 192 -179
rect 205 -210 206 -186
rect 226 -210 227 -186
rect 275 -187 276 -179
rect 30 -210 31 -188
rect 96 -210 97 -188
rect 100 -189 101 -179
rect 261 -189 262 -179
rect 33 -191 34 -179
rect 37 -191 38 -179
rect 44 -191 45 -179
rect 128 -210 129 -190
rect 142 -191 143 -179
rect 184 -210 185 -190
rect 37 -210 38 -192
rect 72 -193 73 -179
rect 107 -193 108 -179
rect 191 -210 192 -192
rect 44 -210 45 -194
rect 121 -195 122 -179
rect 152 -195 153 -179
rect 268 -195 269 -179
rect 61 -210 62 -196
rect 156 -197 157 -179
rect 166 -210 167 -196
rect 170 -197 171 -179
rect 65 -199 66 -179
rect 89 -199 90 -179
rect 103 -199 104 -179
rect 121 -210 122 -198
rect 152 -210 153 -198
rect 212 -199 213 -179
rect 65 -210 66 -200
rect 86 -201 87 -179
rect 89 -210 90 -200
rect 198 -201 199 -179
rect 86 -210 87 -202
rect 163 -203 164 -179
rect 177 -203 178 -179
rect 198 -210 199 -202
rect 100 -210 101 -204
rect 163 -210 164 -204
rect 177 -210 178 -204
rect 233 -205 234 -179
rect 110 -207 111 -179
rect 282 -207 283 -179
rect 93 -209 94 -179
rect 110 -210 111 -208
rect 114 -210 115 -208
rect 142 -210 143 -208
rect 156 -210 157 -208
rect 247 -209 248 -179
rect 23 -247 24 -219
rect 152 -220 153 -218
rect 173 -220 174 -218
rect 226 -220 227 -218
rect 233 -247 234 -219
rect 240 -247 241 -219
rect 275 -247 276 -219
rect 296 -247 297 -219
rect 16 -247 17 -221
rect 152 -247 153 -221
rect 198 -222 199 -218
rect 226 -247 227 -221
rect 30 -224 31 -218
rect 33 -247 34 -223
rect 37 -224 38 -218
rect 75 -224 76 -218
rect 89 -247 90 -223
rect 135 -224 136 -218
rect 138 -247 139 -223
rect 166 -224 167 -218
rect 184 -224 185 -218
rect 198 -247 199 -223
rect 205 -224 206 -218
rect 247 -247 248 -223
rect 30 -247 31 -225
rect 261 -247 262 -225
rect 37 -247 38 -227
rect 61 -228 62 -218
rect 72 -247 73 -227
rect 86 -228 87 -218
rect 93 -228 94 -218
rect 177 -228 178 -218
rect 184 -247 185 -227
rect 278 -247 279 -227
rect 44 -230 45 -218
rect 51 -230 52 -218
rect 54 -247 55 -229
rect 170 -230 171 -218
rect 212 -247 213 -229
rect 219 -230 220 -218
rect 222 -230 223 -218
rect 268 -247 269 -229
rect 47 -247 48 -231
rect 177 -247 178 -231
rect 191 -232 192 -218
rect 219 -247 220 -231
rect 93 -247 94 -233
rect 110 -234 111 -218
rect 114 -234 115 -218
rect 128 -247 129 -233
rect 131 -234 132 -218
rect 254 -247 255 -233
rect 100 -236 101 -218
rect 114 -247 115 -235
rect 121 -236 122 -218
rect 191 -247 192 -235
rect 61 -247 62 -237
rect 100 -247 101 -237
rect 107 -238 108 -218
rect 156 -238 157 -218
rect 65 -240 66 -218
rect 121 -247 122 -239
rect 135 -247 136 -239
rect 170 -247 171 -239
rect 65 -247 66 -241
rect 79 -242 80 -218
rect 110 -247 111 -241
rect 163 -247 164 -241
rect 9 -247 10 -243
rect 79 -247 80 -243
rect 145 -247 146 -243
rect 205 -247 206 -243
rect 149 -247 150 -245
rect 156 -247 157 -245
rect 9 -257 10 -255
rect 58 -257 59 -255
rect 79 -257 80 -255
rect 201 -286 202 -256
rect 219 -257 220 -255
rect 236 -257 237 -255
rect 240 -257 241 -255
rect 243 -263 244 -256
rect 275 -286 276 -256
rect 296 -257 297 -255
rect 9 -286 10 -258
rect 33 -286 34 -258
rect 44 -286 45 -258
rect 72 -259 73 -255
rect 110 -259 111 -255
rect 128 -259 129 -255
rect 135 -259 136 -255
rect 205 -259 206 -255
rect 219 -286 220 -258
rect 254 -259 255 -255
rect 16 -261 17 -255
rect 86 -261 87 -255
rect 138 -261 139 -255
rect 198 -261 199 -255
rect 240 -286 241 -260
rect 261 -261 262 -255
rect 16 -286 17 -262
rect 89 -263 90 -255
rect 142 -263 143 -255
rect 177 -263 178 -255
rect 184 -263 185 -255
rect 184 -286 185 -262
rect 184 -263 185 -255
rect 184 -286 185 -262
rect 261 -286 262 -262
rect 23 -265 24 -255
rect 86 -286 87 -264
rect 89 -286 90 -264
rect 128 -286 129 -264
rect 135 -286 136 -264
rect 142 -286 143 -264
rect 145 -286 146 -264
rect 212 -265 213 -255
rect 247 -265 248 -255
rect 254 -286 255 -264
rect 23 -286 24 -266
rect 51 -267 52 -255
rect 58 -286 59 -266
rect 65 -267 66 -255
rect 107 -286 108 -266
rect 177 -286 178 -266
rect 26 -286 27 -268
rect 233 -286 234 -268
rect 47 -271 48 -255
rect 79 -286 80 -270
rect 152 -271 153 -255
rect 226 -271 227 -255
rect 51 -286 52 -272
rect 100 -273 101 -255
rect 156 -273 157 -255
rect 205 -286 206 -272
rect 65 -286 66 -274
rect 75 -286 76 -274
rect 93 -275 94 -255
rect 100 -286 101 -274
rect 114 -275 115 -255
rect 156 -286 157 -274
rect 170 -275 171 -255
rect 212 -286 213 -274
rect 114 -286 115 -276
rect 149 -277 150 -255
rect 170 -286 171 -276
rect 271 -286 272 -276
rect 149 -286 150 -278
rect 180 -286 181 -278
rect 191 -279 192 -255
rect 226 -286 227 -278
rect 121 -281 122 -255
rect 191 -286 192 -280
rect 121 -286 122 -282
rect 163 -283 164 -255
rect 37 -285 38 -255
rect 163 -286 164 -284
rect 2 -296 3 -294
rect 5 -323 6 -295
rect 23 -323 24 -295
rect 114 -296 115 -294
rect 121 -296 122 -294
rect 131 -323 132 -295
rect 135 -296 136 -294
rect 135 -323 136 -295
rect 135 -296 136 -294
rect 135 -323 136 -295
rect 142 -296 143 -294
rect 212 -296 213 -294
rect 222 -323 223 -295
rect 240 -296 241 -294
rect 247 -296 248 -294
rect 254 -296 255 -294
rect 261 -296 262 -294
rect 271 -296 272 -294
rect 30 -323 31 -297
rect 107 -298 108 -294
rect 142 -323 143 -297
rect 198 -323 199 -297
rect 205 -298 206 -294
rect 212 -323 213 -297
rect 250 -298 251 -294
rect 275 -298 276 -294
rect 16 -300 17 -294
rect 107 -323 108 -299
rect 156 -300 157 -294
rect 177 -300 178 -294
rect 205 -323 206 -299
rect 219 -300 220 -294
rect 37 -302 38 -294
rect 145 -302 146 -294
rect 156 -323 157 -301
rect 191 -302 192 -294
rect 9 -304 10 -294
rect 37 -323 38 -303
rect 40 -323 41 -303
rect 47 -323 48 -303
rect 51 -323 52 -303
rect 117 -323 118 -303
rect 145 -323 146 -303
rect 191 -323 192 -303
rect 2 -323 3 -305
rect 9 -323 10 -305
rect 44 -306 45 -294
rect 96 -306 97 -294
rect 100 -306 101 -294
rect 114 -323 115 -305
rect 170 -306 171 -294
rect 170 -323 171 -305
rect 170 -306 171 -294
rect 170 -323 171 -305
rect 177 -323 178 -305
rect 184 -306 185 -294
rect 58 -308 59 -294
rect 79 -308 80 -294
rect 82 -308 83 -294
rect 89 -308 90 -294
rect 93 -308 94 -294
rect 233 -308 234 -294
rect 58 -323 59 -309
rect 128 -310 129 -294
rect 163 -310 164 -294
rect 184 -323 185 -309
rect 16 -323 17 -311
rect 128 -323 129 -311
rect 149 -312 150 -294
rect 163 -323 164 -311
rect 65 -314 66 -294
rect 121 -323 122 -313
rect 65 -323 66 -315
rect 93 -323 94 -315
rect 103 -323 104 -315
rect 149 -323 150 -315
rect 72 -318 73 -294
rect 226 -318 227 -294
rect 75 -320 76 -294
rect 89 -323 90 -319
rect 100 -323 101 -319
rect 226 -323 227 -319
rect 75 -323 76 -321
rect 79 -323 80 -321
rect 2 -354 3 -332
rect 9 -333 10 -331
rect 16 -333 17 -331
rect 68 -354 69 -332
rect 72 -333 73 -331
rect 107 -333 108 -331
rect 114 -333 115 -331
rect 198 -333 199 -331
rect 23 -335 24 -331
rect 86 -335 87 -331
rect 96 -335 97 -331
rect 184 -335 185 -331
rect 198 -354 199 -334
rect 226 -335 227 -331
rect 30 -337 31 -331
rect 103 -337 104 -331
rect 107 -354 108 -336
rect 131 -337 132 -331
rect 135 -337 136 -331
rect 142 -354 143 -336
rect 149 -337 150 -331
rect 170 -337 171 -331
rect 177 -337 178 -331
rect 177 -354 178 -336
rect 177 -337 178 -331
rect 177 -354 178 -336
rect 184 -354 185 -336
rect 219 -337 220 -331
rect 30 -354 31 -338
rect 58 -339 59 -331
rect 96 -354 97 -338
rect 128 -339 129 -331
rect 135 -354 136 -338
rect 159 -354 160 -338
rect 163 -339 164 -331
rect 163 -354 164 -338
rect 163 -339 164 -331
rect 163 -354 164 -338
rect 170 -354 171 -338
rect 205 -339 206 -331
rect 23 -354 24 -340
rect 58 -354 59 -340
rect 93 -341 94 -331
rect 128 -354 129 -340
rect 156 -341 157 -331
rect 191 -341 192 -331
rect 37 -354 38 -342
rect 117 -343 118 -331
rect 191 -354 192 -342
rect 212 -343 213 -331
rect 40 -345 41 -331
rect 75 -345 76 -331
rect 100 -345 101 -331
rect 121 -345 122 -331
rect 44 -347 45 -331
rect 61 -354 62 -346
rect 79 -347 80 -331
rect 100 -354 101 -346
rect 114 -354 115 -346
rect 149 -354 150 -346
rect 44 -354 45 -348
rect 65 -349 66 -331
rect 121 -354 122 -348
rect 215 -354 216 -348
rect 51 -351 52 -331
rect 72 -354 73 -350
rect 51 -354 52 -352
rect 79 -354 80 -352
rect 12 -387 13 -363
rect 16 -387 17 -363
rect 23 -364 24 -362
rect 44 -387 45 -363
rect 65 -387 66 -363
rect 79 -364 80 -362
rect 86 -364 87 -362
rect 163 -364 164 -362
rect 184 -364 185 -362
rect 208 -364 209 -362
rect 23 -387 24 -365
rect 47 -387 48 -365
rect 72 -366 73 -362
rect 72 -387 73 -365
rect 72 -366 73 -362
rect 72 -387 73 -365
rect 100 -366 101 -362
rect 100 -387 101 -365
rect 100 -366 101 -362
rect 100 -387 101 -365
rect 114 -366 115 -362
rect 205 -387 206 -365
rect 30 -368 31 -362
rect 58 -368 59 -362
rect 117 -368 118 -362
rect 121 -368 122 -362
rect 138 -387 139 -367
rect 222 -387 223 -367
rect 30 -387 31 -369
rect 51 -387 52 -369
rect 58 -387 59 -369
rect 68 -370 69 -362
rect 121 -387 122 -369
rect 135 -370 136 -362
rect 142 -370 143 -362
rect 163 -387 164 -369
rect 184 -387 185 -369
rect 198 -370 199 -362
rect 37 -372 38 -362
rect 170 -372 171 -362
rect 191 -372 192 -362
rect 212 -372 213 -362
rect 96 -374 97 -362
rect 191 -387 192 -373
rect 79 -387 80 -375
rect 96 -387 97 -375
rect 114 -387 115 -375
rect 170 -387 171 -375
rect 149 -378 150 -362
rect 226 -387 227 -377
rect 156 -380 157 -362
rect 212 -387 213 -379
rect 128 -382 129 -362
rect 156 -387 157 -381
rect 159 -382 160 -362
rect 177 -382 178 -362
rect 107 -384 108 -362
rect 177 -387 178 -383
rect 107 -387 108 -385
rect 142 -387 143 -385
rect 23 -397 24 -395
rect 149 -420 150 -396
rect 152 -397 153 -395
rect 184 -397 185 -395
rect 198 -397 199 -395
rect 198 -420 199 -396
rect 198 -397 199 -395
rect 198 -420 199 -396
rect 26 -420 27 -398
rect 128 -399 129 -395
rect 131 -399 132 -395
rect 177 -399 178 -395
rect 30 -401 31 -395
rect 44 -420 45 -400
rect 54 -401 55 -395
rect 58 -401 59 -395
rect 79 -401 80 -395
rect 107 -420 108 -400
rect 110 -401 111 -395
rect 191 -401 192 -395
rect 16 -403 17 -395
rect 30 -420 31 -402
rect 40 -403 41 -395
rect 170 -403 171 -395
rect 54 -420 55 -404
rect 156 -405 157 -395
rect 37 -407 38 -395
rect 156 -420 157 -406
rect 61 -420 62 -408
rect 79 -420 80 -408
rect 82 -420 83 -408
rect 128 -420 129 -408
rect 135 -420 136 -408
rect 187 -409 188 -395
rect 86 -411 87 -395
rect 100 -411 101 -395
rect 117 -411 118 -395
rect 205 -411 206 -395
rect 89 -413 90 -395
rect 96 -413 97 -395
rect 100 -420 101 -412
rect 142 -413 143 -395
rect 187 -420 188 -412
rect 212 -413 213 -395
rect 65 -415 66 -395
rect 96 -420 97 -414
rect 138 -415 139 -395
rect 226 -415 227 -395
rect 65 -420 66 -416
rect 72 -417 73 -395
rect 93 -420 94 -416
rect 114 -417 115 -395
rect 142 -420 143 -416
rect 163 -417 164 -395
rect 114 -420 115 -418
rect 121 -419 122 -395
rect 12 -430 13 -428
rect 128 -430 129 -428
rect 19 -432 20 -428
rect 30 -432 31 -428
rect 47 -432 48 -428
rect 61 -432 62 -428
rect 65 -432 66 -428
rect 75 -432 76 -428
rect 79 -432 80 -428
rect 156 -432 157 -428
rect 72 -434 73 -428
rect 149 -434 150 -428
rect 89 -436 90 -428
rect 107 -436 108 -428
rect 114 -436 115 -428
rect 124 -436 125 -428
rect 96 -438 97 -428
rect 100 -438 101 -428
rect 121 -438 122 -428
rect 142 -438 143 -428
<< labels >>
rlabel pdiffusion 3 -6 3 -6 0 cellNo=35
rlabel pdiffusion 10 -6 10 -6 0 cellNo=64
rlabel pdiffusion 17 -6 17 -6 0 cellNo=106
rlabel pdiffusion 24 -6 24 -6 0 cellNo=109
rlabel pdiffusion 73 -6 73 -6 0 cellNo=48
rlabel pdiffusion 80 -6 80 -6 0 feedthrough
rlabel pdiffusion 101 -6 101 -6 0 cellNo=110
rlabel pdiffusion 108 -6 108 -6 0 feedthrough
rlabel pdiffusion 115 -6 115 -6 0 cellNo=32
rlabel pdiffusion 122 -6 122 -6 0 cellNo=174
rlabel pdiffusion 129 -6 129 -6 0 feedthrough
rlabel pdiffusion 3 -27 3 -27 0 cellNo=67
rlabel pdiffusion 10 -27 10 -27 0 cellNo=108
rlabel pdiffusion 45 -27 45 -27 0 feedthrough
rlabel pdiffusion 52 -27 52 -27 0 feedthrough
rlabel pdiffusion 59 -27 59 -27 0 cellNo=63
rlabel pdiffusion 66 -27 66 -27 0 cellNo=23
rlabel pdiffusion 73 -27 73 -27 0 feedthrough
rlabel pdiffusion 80 -27 80 -27 0 cellNo=73
rlabel pdiffusion 87 -27 87 -27 0 feedthrough
rlabel pdiffusion 94 -27 94 -27 0 cellNo=131
rlabel pdiffusion 101 -27 101 -27 0 feedthrough
rlabel pdiffusion 108 -27 108 -27 0 cellNo=76
rlabel pdiffusion 115 -27 115 -27 0 cellNo=52
rlabel pdiffusion 122 -27 122 -27 0 feedthrough
rlabel pdiffusion 129 -27 129 -27 0 feedthrough
rlabel pdiffusion 136 -27 136 -27 0 feedthrough
rlabel pdiffusion 143 -27 143 -27 0 feedthrough
rlabel pdiffusion 157 -27 157 -27 0 cellNo=79
rlabel pdiffusion 262 -27 262 -27 0 cellNo=21
rlabel pdiffusion 3 -48 3 -48 0 cellNo=62
rlabel pdiffusion 10 -48 10 -48 0 cellNo=157
rlabel pdiffusion 31 -48 31 -48 0 cellNo=24
rlabel pdiffusion 38 -48 38 -48 0 cellNo=58
rlabel pdiffusion 45 -48 45 -48 0 feedthrough
rlabel pdiffusion 52 -48 52 -48 0 feedthrough
rlabel pdiffusion 59 -48 59 -48 0 cellNo=101
rlabel pdiffusion 66 -48 66 -48 0 cellNo=4
rlabel pdiffusion 73 -48 73 -48 0 cellNo=26
rlabel pdiffusion 80 -48 80 -48 0 feedthrough
rlabel pdiffusion 87 -48 87 -48 0 cellNo=92
rlabel pdiffusion 94 -48 94 -48 0 feedthrough
rlabel pdiffusion 101 -48 101 -48 0 feedthrough
rlabel pdiffusion 108 -48 108 -48 0 feedthrough
rlabel pdiffusion 115 -48 115 -48 0 cellNo=154
rlabel pdiffusion 129 -48 129 -48 0 cellNo=15
rlabel pdiffusion 136 -48 136 -48 0 feedthrough
rlabel pdiffusion 143 -48 143 -48 0 feedthrough
rlabel pdiffusion 150 -48 150 -48 0 cellNo=45
rlabel pdiffusion 164 -48 164 -48 0 cellNo=138
rlabel pdiffusion 171 -48 171 -48 0 feedthrough
rlabel pdiffusion 178 -48 178 -48 0 feedthrough
rlabel pdiffusion 234 -48 234 -48 0 cellNo=71
rlabel pdiffusion 248 -48 248 -48 0 feedthrough
rlabel pdiffusion 3 -71 3 -71 0 feedthrough
rlabel pdiffusion 10 -71 10 -71 0 cellNo=147
rlabel pdiffusion 17 -71 17 -71 0 cellNo=28
rlabel pdiffusion 24 -71 24 -71 0 feedthrough
rlabel pdiffusion 31 -71 31 -71 0 cellNo=88
rlabel pdiffusion 38 -71 38 -71 0 cellNo=125
rlabel pdiffusion 45 -71 45 -71 0 feedthrough
rlabel pdiffusion 52 -71 52 -71 0 feedthrough
rlabel pdiffusion 59 -71 59 -71 0 feedthrough
rlabel pdiffusion 66 -71 66 -71 0 feedthrough
rlabel pdiffusion 73 -71 73 -71 0 cellNo=135
rlabel pdiffusion 80 -71 80 -71 0 cellNo=6
rlabel pdiffusion 87 -71 87 -71 0 cellNo=59
rlabel pdiffusion 94 -71 94 -71 0 cellNo=65
rlabel pdiffusion 101 -71 101 -71 0 feedthrough
rlabel pdiffusion 108 -71 108 -71 0 feedthrough
rlabel pdiffusion 115 -71 115 -71 0 cellNo=69
rlabel pdiffusion 122 -71 122 -71 0 feedthrough
rlabel pdiffusion 129 -71 129 -71 0 feedthrough
rlabel pdiffusion 136 -71 136 -71 0 cellNo=37
rlabel pdiffusion 143 -71 143 -71 0 feedthrough
rlabel pdiffusion 150 -71 150 -71 0 feedthrough
rlabel pdiffusion 157 -71 157 -71 0 feedthrough
rlabel pdiffusion 164 -71 164 -71 0 feedthrough
rlabel pdiffusion 171 -71 171 -71 0 cellNo=170
rlabel pdiffusion 178 -71 178 -71 0 feedthrough
rlabel pdiffusion 185 -71 185 -71 0 feedthrough
rlabel pdiffusion 192 -71 192 -71 0 cellNo=136
rlabel pdiffusion 199 -71 199 -71 0 feedthrough
rlabel pdiffusion 206 -71 206 -71 0 feedthrough
rlabel pdiffusion 213 -71 213 -71 0 cellNo=49
rlabel pdiffusion 220 -71 220 -71 0 feedthrough
rlabel pdiffusion 227 -71 227 -71 0 cellNo=66
rlabel pdiffusion 234 -71 234 -71 0 feedthrough
rlabel pdiffusion 10 -100 10 -100 0 feedthrough
rlabel pdiffusion 17 -100 17 -100 0 feedthrough
rlabel pdiffusion 24 -100 24 -100 0 feedthrough
rlabel pdiffusion 31 -100 31 -100 0 cellNo=122
rlabel pdiffusion 38 -100 38 -100 0 feedthrough
rlabel pdiffusion 45 -100 45 -100 0 cellNo=85
rlabel pdiffusion 52 -100 52 -100 0 cellNo=1
rlabel pdiffusion 59 -100 59 -100 0 feedthrough
rlabel pdiffusion 66 -100 66 -100 0 cellNo=143
rlabel pdiffusion 73 -100 73 -100 0 feedthrough
rlabel pdiffusion 80 -100 80 -100 0 cellNo=177
rlabel pdiffusion 87 -100 87 -100 0 feedthrough
rlabel pdiffusion 94 -100 94 -100 0 cellNo=68
rlabel pdiffusion 101 -100 101 -100 0 feedthrough
rlabel pdiffusion 108 -100 108 -100 0 feedthrough
rlabel pdiffusion 115 -100 115 -100 0 feedthrough
rlabel pdiffusion 122 -100 122 -100 0 cellNo=104
rlabel pdiffusion 129 -100 129 -100 0 cellNo=55
rlabel pdiffusion 136 -100 136 -100 0 cellNo=51
rlabel pdiffusion 143 -100 143 -100 0 cellNo=82
rlabel pdiffusion 150 -100 150 -100 0 cellNo=60
rlabel pdiffusion 157 -100 157 -100 0 feedthrough
rlabel pdiffusion 164 -100 164 -100 0 cellNo=50
rlabel pdiffusion 171 -100 171 -100 0 feedthrough
rlabel pdiffusion 178 -100 178 -100 0 feedthrough
rlabel pdiffusion 185 -100 185 -100 0 feedthrough
rlabel pdiffusion 192 -100 192 -100 0 feedthrough
rlabel pdiffusion 199 -100 199 -100 0 feedthrough
rlabel pdiffusion 206 -100 206 -100 0 feedthrough
rlabel pdiffusion 213 -100 213 -100 0 feedthrough
rlabel pdiffusion 220 -100 220 -100 0 feedthrough
rlabel pdiffusion 227 -100 227 -100 0 feedthrough
rlabel pdiffusion 234 -100 234 -100 0 feedthrough
rlabel pdiffusion 241 -100 241 -100 0 feedthrough
rlabel pdiffusion 248 -100 248 -100 0 feedthrough
rlabel pdiffusion 255 -100 255 -100 0 feedthrough
rlabel pdiffusion 262 -100 262 -100 0 cellNo=12
rlabel pdiffusion 269 -100 269 -100 0 cellNo=120
rlabel pdiffusion 283 -100 283 -100 0 feedthrough
rlabel pdiffusion 10 -133 10 -133 0 feedthrough
rlabel pdiffusion 17 -133 17 -133 0 feedthrough
rlabel pdiffusion 24 -133 24 -133 0 feedthrough
rlabel pdiffusion 31 -133 31 -133 0 cellNo=93
rlabel pdiffusion 38 -133 38 -133 0 cellNo=44
rlabel pdiffusion 45 -133 45 -133 0 cellNo=178
rlabel pdiffusion 52 -133 52 -133 0 feedthrough
rlabel pdiffusion 59 -133 59 -133 0 feedthrough
rlabel pdiffusion 66 -133 66 -133 0 feedthrough
rlabel pdiffusion 73 -133 73 -133 0 cellNo=91
rlabel pdiffusion 80 -133 80 -133 0 feedthrough
rlabel pdiffusion 87 -133 87 -133 0 feedthrough
rlabel pdiffusion 94 -133 94 -133 0 cellNo=33
rlabel pdiffusion 101 -133 101 -133 0 feedthrough
rlabel pdiffusion 108 -133 108 -133 0 cellNo=162
rlabel pdiffusion 115 -133 115 -133 0 cellNo=87
rlabel pdiffusion 122 -133 122 -133 0 feedthrough
rlabel pdiffusion 129 -133 129 -133 0 feedthrough
rlabel pdiffusion 136 -133 136 -133 0 cellNo=7
rlabel pdiffusion 143 -133 143 -133 0 feedthrough
rlabel pdiffusion 150 -133 150 -133 0 cellNo=29
rlabel pdiffusion 157 -133 157 -133 0 cellNo=25
rlabel pdiffusion 164 -133 164 -133 0 feedthrough
rlabel pdiffusion 171 -133 171 -133 0 cellNo=2
rlabel pdiffusion 178 -133 178 -133 0 cellNo=107
rlabel pdiffusion 185 -133 185 -133 0 cellNo=3
rlabel pdiffusion 192 -133 192 -133 0 feedthrough
rlabel pdiffusion 199 -133 199 -133 0 feedthrough
rlabel pdiffusion 206 -133 206 -133 0 cellNo=160
rlabel pdiffusion 213 -133 213 -133 0 feedthrough
rlabel pdiffusion 220 -133 220 -133 0 feedthrough
rlabel pdiffusion 227 -133 227 -133 0 feedthrough
rlabel pdiffusion 234 -133 234 -133 0 feedthrough
rlabel pdiffusion 297 -133 297 -133 0 feedthrough
rlabel pdiffusion 3 -176 3 -176 0 feedthrough
rlabel pdiffusion 10 -176 10 -176 0 feedthrough
rlabel pdiffusion 17 -176 17 -176 0 feedthrough
rlabel pdiffusion 24 -176 24 -176 0 feedthrough
rlabel pdiffusion 31 -176 31 -176 0 cellNo=127
rlabel pdiffusion 38 -176 38 -176 0 feedthrough
rlabel pdiffusion 45 -176 45 -176 0 feedthrough
rlabel pdiffusion 52 -176 52 -176 0 cellNo=43
rlabel pdiffusion 59 -176 59 -176 0 feedthrough
rlabel pdiffusion 66 -176 66 -176 0 cellNo=86
rlabel pdiffusion 73 -176 73 -176 0 feedthrough
rlabel pdiffusion 80 -176 80 -176 0 feedthrough
rlabel pdiffusion 87 -176 87 -176 0 cellNo=153
rlabel pdiffusion 94 -176 94 -176 0 cellNo=5
rlabel pdiffusion 101 -176 101 -176 0 cellNo=133
rlabel pdiffusion 108 -176 108 -176 0 cellNo=54
rlabel pdiffusion 115 -176 115 -176 0 cellNo=9
rlabel pdiffusion 122 -176 122 -176 0 cellNo=111
rlabel pdiffusion 129 -176 129 -176 0 cellNo=70
rlabel pdiffusion 136 -176 136 -176 0 cellNo=20
rlabel pdiffusion 143 -176 143 -176 0 feedthrough
rlabel pdiffusion 150 -176 150 -176 0 cellNo=42
rlabel pdiffusion 157 -176 157 -176 0 feedthrough
rlabel pdiffusion 164 -176 164 -176 0 cellNo=57
rlabel pdiffusion 171 -176 171 -176 0 feedthrough
rlabel pdiffusion 178 -176 178 -176 0 feedthrough
rlabel pdiffusion 185 -176 185 -176 0 feedthrough
rlabel pdiffusion 192 -176 192 -176 0 feedthrough
rlabel pdiffusion 199 -176 199 -176 0 feedthrough
rlabel pdiffusion 206 -176 206 -176 0 feedthrough
rlabel pdiffusion 213 -176 213 -176 0 feedthrough
rlabel pdiffusion 220 -176 220 -176 0 feedthrough
rlabel pdiffusion 227 -176 227 -176 0 feedthrough
rlabel pdiffusion 234 -176 234 -176 0 feedthrough
rlabel pdiffusion 241 -176 241 -176 0 feedthrough
rlabel pdiffusion 248 -176 248 -176 0 feedthrough
rlabel pdiffusion 255 -176 255 -176 0 feedthrough
rlabel pdiffusion 262 -176 262 -176 0 feedthrough
rlabel pdiffusion 269 -176 269 -176 0 feedthrough
rlabel pdiffusion 276 -176 276 -176 0 feedthrough
rlabel pdiffusion 283 -176 283 -176 0 feedthrough
rlabel pdiffusion 31 -215 31 -215 0 feedthrough
rlabel pdiffusion 38 -215 38 -215 0 feedthrough
rlabel pdiffusion 45 -215 45 -215 0 cellNo=130
rlabel pdiffusion 52 -215 52 -215 0 cellNo=139
rlabel pdiffusion 59 -215 59 -215 0 cellNo=144
rlabel pdiffusion 66 -215 66 -215 0 feedthrough
rlabel pdiffusion 73 -215 73 -215 0 cellNo=41
rlabel pdiffusion 80 -215 80 -215 0 feedthrough
rlabel pdiffusion 87 -215 87 -215 0 cellNo=17
rlabel pdiffusion 94 -215 94 -215 0 cellNo=102
rlabel pdiffusion 101 -215 101 -215 0 feedthrough
rlabel pdiffusion 108 -215 108 -215 0 cellNo=179
rlabel pdiffusion 115 -215 115 -215 0 feedthrough
rlabel pdiffusion 122 -215 122 -215 0 feedthrough
rlabel pdiffusion 129 -215 129 -215 0 cellNo=47
rlabel pdiffusion 136 -215 136 -215 0 feedthrough
rlabel pdiffusion 143 -215 143 -215 0 cellNo=89
rlabel pdiffusion 150 -215 150 -215 0 cellNo=119
rlabel pdiffusion 157 -215 157 -215 0 feedthrough
rlabel pdiffusion 164 -215 164 -215 0 cellNo=36
rlabel pdiffusion 171 -215 171 -215 0 cellNo=145
rlabel pdiffusion 178 -215 178 -215 0 feedthrough
rlabel pdiffusion 185 -215 185 -215 0 feedthrough
rlabel pdiffusion 192 -215 192 -215 0 feedthrough
rlabel pdiffusion 199 -215 199 -215 0 feedthrough
rlabel pdiffusion 206 -215 206 -215 0 feedthrough
rlabel pdiffusion 220 -215 220 -215 0 cellNo=146
rlabel pdiffusion 227 -215 227 -215 0 feedthrough
rlabel pdiffusion 10 -252 10 -252 0 feedthrough
rlabel pdiffusion 17 -252 17 -252 0 feedthrough
rlabel pdiffusion 24 -252 24 -252 0 feedthrough
rlabel pdiffusion 31 -252 31 -252 0 cellNo=141
rlabel pdiffusion 38 -252 38 -252 0 feedthrough
rlabel pdiffusion 45 -252 45 -252 0 cellNo=90
rlabel pdiffusion 52 -252 52 -252 0 cellNo=172
rlabel pdiffusion 59 -252 59 -252 0 cellNo=121
rlabel pdiffusion 66 -252 66 -252 0 feedthrough
rlabel pdiffusion 73 -252 73 -252 0 feedthrough
rlabel pdiffusion 80 -252 80 -252 0 cellNo=112
rlabel pdiffusion 87 -252 87 -252 0 cellNo=77
rlabel pdiffusion 94 -252 94 -252 0 feedthrough
rlabel pdiffusion 101 -252 101 -252 0 feedthrough
rlabel pdiffusion 108 -252 108 -252 0 cellNo=95
rlabel pdiffusion 115 -252 115 -252 0 feedthrough
rlabel pdiffusion 122 -252 122 -252 0 cellNo=78
rlabel pdiffusion 129 -252 129 -252 0 feedthrough
rlabel pdiffusion 136 -252 136 -252 0 cellNo=137
rlabel pdiffusion 143 -252 143 -252 0 cellNo=129
rlabel pdiffusion 150 -252 150 -252 0 cellNo=124
rlabel pdiffusion 157 -252 157 -252 0 feedthrough
rlabel pdiffusion 164 -252 164 -252 0 feedthrough
rlabel pdiffusion 171 -252 171 -252 0 feedthrough
rlabel pdiffusion 178 -252 178 -252 0 feedthrough
rlabel pdiffusion 185 -252 185 -252 0 feedthrough
rlabel pdiffusion 192 -252 192 -252 0 feedthrough
rlabel pdiffusion 199 -252 199 -252 0 feedthrough
rlabel pdiffusion 206 -252 206 -252 0 feedthrough
rlabel pdiffusion 213 -252 213 -252 0 feedthrough
rlabel pdiffusion 220 -252 220 -252 0 feedthrough
rlabel pdiffusion 227 -252 227 -252 0 feedthrough
rlabel pdiffusion 234 -252 234 -252 0 cellNo=39
rlabel pdiffusion 241 -252 241 -252 0 feedthrough
rlabel pdiffusion 248 -252 248 -252 0 feedthrough
rlabel pdiffusion 255 -252 255 -252 0 feedthrough
rlabel pdiffusion 262 -252 262 -252 0 feedthrough
rlabel pdiffusion 269 -252 269 -252 0 cellNo=74
rlabel pdiffusion 276 -252 276 -252 0 cellNo=14
rlabel pdiffusion 297 -252 297 -252 0 feedthrough
rlabel pdiffusion 3 -291 3 -291 0 cellNo=155
rlabel pdiffusion 10 -291 10 -291 0 feedthrough
rlabel pdiffusion 17 -291 17 -291 0 feedthrough
rlabel pdiffusion 24 -291 24 -291 0 cellNo=168
rlabel pdiffusion 31 -291 31 -291 0 cellNo=115
rlabel pdiffusion 38 -291 38 -291 0 cellNo=161
rlabel pdiffusion 45 -291 45 -291 0 feedthrough
rlabel pdiffusion 52 -291 52 -291 0 cellNo=175
rlabel pdiffusion 59 -291 59 -291 0 feedthrough
rlabel pdiffusion 66 -291 66 -291 0 feedthrough
rlabel pdiffusion 73 -291 73 -291 0 cellNo=116
rlabel pdiffusion 80 -291 80 -291 0 cellNo=132
rlabel pdiffusion 87 -291 87 -291 0 cellNo=126
rlabel pdiffusion 94 -291 94 -291 0 cellNo=151
rlabel pdiffusion 101 -291 101 -291 0 feedthrough
rlabel pdiffusion 108 -291 108 -291 0 feedthrough
rlabel pdiffusion 115 -291 115 -291 0 feedthrough
rlabel pdiffusion 122 -291 122 -291 0 feedthrough
rlabel pdiffusion 129 -291 129 -291 0 feedthrough
rlabel pdiffusion 136 -291 136 -291 0 feedthrough
rlabel pdiffusion 143 -291 143 -291 0 cellNo=159
rlabel pdiffusion 150 -291 150 -291 0 feedthrough
rlabel pdiffusion 157 -291 157 -291 0 feedthrough
rlabel pdiffusion 164 -291 164 -291 0 feedthrough
rlabel pdiffusion 171 -291 171 -291 0 feedthrough
rlabel pdiffusion 178 -291 178 -291 0 cellNo=134
rlabel pdiffusion 185 -291 185 -291 0 feedthrough
rlabel pdiffusion 192 -291 192 -291 0 feedthrough
rlabel pdiffusion 199 -291 199 -291 0 cellNo=22
rlabel pdiffusion 206 -291 206 -291 0 feedthrough
rlabel pdiffusion 213 -291 213 -291 0 feedthrough
rlabel pdiffusion 220 -291 220 -291 0 feedthrough
rlabel pdiffusion 227 -291 227 -291 0 feedthrough
rlabel pdiffusion 234 -291 234 -291 0 feedthrough
rlabel pdiffusion 241 -291 241 -291 0 feedthrough
rlabel pdiffusion 248 -291 248 -291 0 cellNo=81
rlabel pdiffusion 255 -291 255 -291 0 feedthrough
rlabel pdiffusion 262 -291 262 -291 0 feedthrough
rlabel pdiffusion 269 -291 269 -291 0 cellNo=176
rlabel pdiffusion 276 -291 276 -291 0 feedthrough
rlabel pdiffusion 3 -328 3 -328 0 cellNo=105
rlabel pdiffusion 10 -328 10 -328 0 feedthrough
rlabel pdiffusion 17 -328 17 -328 0 feedthrough
rlabel pdiffusion 24 -328 24 -328 0 feedthrough
rlabel pdiffusion 31 -328 31 -328 0 feedthrough
rlabel pdiffusion 38 -328 38 -328 0 cellNo=169
rlabel pdiffusion 45 -328 45 -328 0 cellNo=11
rlabel pdiffusion 52 -328 52 -328 0 feedthrough
rlabel pdiffusion 59 -328 59 -328 0 feedthrough
rlabel pdiffusion 66 -328 66 -328 0 feedthrough
rlabel pdiffusion 73 -328 73 -328 0 cellNo=16
rlabel pdiffusion 80 -328 80 -328 0 feedthrough
rlabel pdiffusion 87 -328 87 -328 0 cellNo=123
rlabel pdiffusion 94 -328 94 -328 0 cellNo=38
rlabel pdiffusion 101 -328 101 -328 0 cellNo=84
rlabel pdiffusion 108 -328 108 -328 0 feedthrough
rlabel pdiffusion 115 -328 115 -328 0 cellNo=166
rlabel pdiffusion 122 -328 122 -328 0 feedthrough
rlabel pdiffusion 129 -328 129 -328 0 cellNo=152
rlabel pdiffusion 136 -328 136 -328 0 feedthrough
rlabel pdiffusion 143 -328 143 -328 0 cellNo=142
rlabel pdiffusion 150 -328 150 -328 0 cellNo=40
rlabel pdiffusion 157 -328 157 -328 0 cellNo=180
rlabel pdiffusion 164 -328 164 -328 0 feedthrough
rlabel pdiffusion 171 -328 171 -328 0 feedthrough
rlabel pdiffusion 178 -328 178 -328 0 feedthrough
rlabel pdiffusion 185 -328 185 -328 0 feedthrough
rlabel pdiffusion 192 -328 192 -328 0 feedthrough
rlabel pdiffusion 199 -328 199 -328 0 feedthrough
rlabel pdiffusion 206 -328 206 -328 0 feedthrough
rlabel pdiffusion 213 -328 213 -328 0 feedthrough
rlabel pdiffusion 220 -328 220 -328 0 cellNo=19
rlabel pdiffusion 227 -328 227 -328 0 feedthrough
rlabel pdiffusion 3 -359 3 -359 0 cellNo=10
rlabel pdiffusion 24 -359 24 -359 0 feedthrough
rlabel pdiffusion 31 -359 31 -359 0 feedthrough
rlabel pdiffusion 38 -359 38 -359 0 feedthrough
rlabel pdiffusion 45 -359 45 -359 0 cellNo=46
rlabel pdiffusion 52 -359 52 -359 0 cellNo=94
rlabel pdiffusion 59 -359 59 -359 0 cellNo=158
rlabel pdiffusion 66 -359 66 -359 0 cellNo=56
rlabel pdiffusion 73 -359 73 -359 0 feedthrough
rlabel pdiffusion 80 -359 80 -359 0 feedthrough
rlabel pdiffusion 87 -359 87 -359 0 cellNo=13
rlabel pdiffusion 94 -359 94 -359 0 cellNo=75
rlabel pdiffusion 101 -359 101 -359 0 feedthrough
rlabel pdiffusion 108 -359 108 -359 0 feedthrough
rlabel pdiffusion 115 -359 115 -359 0 cellNo=30
rlabel pdiffusion 122 -359 122 -359 0 feedthrough
rlabel pdiffusion 129 -359 129 -359 0 feedthrough
rlabel pdiffusion 136 -359 136 -359 0 feedthrough
rlabel pdiffusion 143 -359 143 -359 0 feedthrough
rlabel pdiffusion 150 -359 150 -359 0 feedthrough
rlabel pdiffusion 157 -359 157 -359 0 cellNo=165
rlabel pdiffusion 164 -359 164 -359 0 feedthrough
rlabel pdiffusion 171 -359 171 -359 0 cellNo=98
rlabel pdiffusion 178 -359 178 -359 0 feedthrough
rlabel pdiffusion 185 -359 185 -359 0 feedthrough
rlabel pdiffusion 192 -359 192 -359 0 feedthrough
rlabel pdiffusion 199 -359 199 -359 0 feedthrough
rlabel pdiffusion 206 -359 206 -359 0 cellNo=99
rlabel pdiffusion 213 -359 213 -359 0 cellNo=80
rlabel pdiffusion 10 -392 10 -392 0 cellNo=128
rlabel pdiffusion 17 -392 17 -392 0 feedthrough
rlabel pdiffusion 24 -392 24 -392 0 feedthrough
rlabel pdiffusion 31 -392 31 -392 0 feedthrough
rlabel pdiffusion 38 -392 38 -392 0 cellNo=34
rlabel pdiffusion 45 -392 45 -392 0 cellNo=103
rlabel pdiffusion 52 -392 52 -392 0 cellNo=27
rlabel pdiffusion 59 -392 59 -392 0 feedthrough
rlabel pdiffusion 66 -392 66 -392 0 feedthrough
rlabel pdiffusion 73 -392 73 -392 0 feedthrough
rlabel pdiffusion 80 -392 80 -392 0 feedthrough
rlabel pdiffusion 87 -392 87 -392 0 cellNo=113
rlabel pdiffusion 94 -392 94 -392 0 cellNo=140
rlabel pdiffusion 101 -392 101 -392 0 feedthrough
rlabel pdiffusion 108 -392 108 -392 0 cellNo=148
rlabel pdiffusion 115 -392 115 -392 0 cellNo=53
rlabel pdiffusion 122 -392 122 -392 0 feedthrough
rlabel pdiffusion 129 -392 129 -392 0 cellNo=163
rlabel pdiffusion 136 -392 136 -392 0 cellNo=8
rlabel pdiffusion 143 -392 143 -392 0 feedthrough
rlabel pdiffusion 150 -392 150 -392 0 cellNo=18
rlabel pdiffusion 157 -392 157 -392 0 feedthrough
rlabel pdiffusion 164 -392 164 -392 0 feedthrough
rlabel pdiffusion 171 -392 171 -392 0 feedthrough
rlabel pdiffusion 178 -392 178 -392 0 feedthrough
rlabel pdiffusion 185 -392 185 -392 0 cellNo=171
rlabel pdiffusion 192 -392 192 -392 0 feedthrough
rlabel pdiffusion 199 -392 199 -392 0 cellNo=96
rlabel pdiffusion 206 -392 206 -392 0 feedthrough
rlabel pdiffusion 213 -392 213 -392 0 feedthrough
rlabel pdiffusion 220 -392 220 -392 0 cellNo=156
rlabel pdiffusion 227 -392 227 -392 0 feedthrough
rlabel pdiffusion 10 -425 10 -425 0 cellNo=31
rlabel pdiffusion 17 -425 17 -425 0 cellNo=61
rlabel pdiffusion 24 -425 24 -425 0 cellNo=72
rlabel pdiffusion 31 -425 31 -425 0 feedthrough
rlabel pdiffusion 45 -425 45 -425 0 cellNo=150
rlabel pdiffusion 52 -425 52 -425 0 cellNo=164
rlabel pdiffusion 59 -425 59 -425 0 cellNo=149
rlabel pdiffusion 66 -425 66 -425 0 feedthrough
rlabel pdiffusion 73 -425 73 -425 0 cellNo=173
rlabel pdiffusion 80 -425 80 -425 0 cellNo=118
rlabel pdiffusion 87 -425 87 -425 0 cellNo=117
rlabel pdiffusion 94 -425 94 -425 0 cellNo=97
rlabel pdiffusion 101 -425 101 -425 0 feedthrough
rlabel pdiffusion 108 -425 108 -425 0 feedthrough
rlabel pdiffusion 115 -425 115 -425 0 feedthrough
rlabel pdiffusion 122 -425 122 -425 0 cellNo=83
rlabel pdiffusion 129 -425 129 -425 0 feedthrough
rlabel pdiffusion 136 -425 136 -425 0 cellNo=167
rlabel pdiffusion 143 -425 143 -425 0 feedthrough
rlabel pdiffusion 150 -425 150 -425 0 feedthrough
rlabel pdiffusion 157 -425 157 -425 0 feedthrough
rlabel pdiffusion 185 -425 185 -425 0 cellNo=100
rlabel pdiffusion 199 -425 199 -425 0 cellNo=114
rlabel polysilicon 72 -2 72 -2 0 1
rlabel polysilicon 75 -8 75 -8 0 4
rlabel polysilicon 79 -2 79 -2 0 1
rlabel polysilicon 79 -8 79 -8 0 3
rlabel polysilicon 100 -2 100 -2 0 1
rlabel polysilicon 107 -2 107 -2 0 1
rlabel polysilicon 107 -8 107 -8 0 3
rlabel polysilicon 114 -8 114 -8 0 3
rlabel polysilicon 121 -2 121 -2 0 1
rlabel polysilicon 128 -2 128 -2 0 1
rlabel polysilicon 128 -8 128 -8 0 3
rlabel polysilicon 44 -23 44 -23 0 1
rlabel polysilicon 44 -29 44 -29 0 3
rlabel polysilicon 51 -23 51 -23 0 1
rlabel polysilicon 51 -29 51 -29 0 3
rlabel polysilicon 61 -23 61 -23 0 2
rlabel polysilicon 68 -23 68 -23 0 2
rlabel polysilicon 72 -23 72 -23 0 1
rlabel polysilicon 72 -29 72 -29 0 3
rlabel polysilicon 79 -23 79 -23 0 1
rlabel polysilicon 82 -23 82 -23 0 2
rlabel polysilicon 86 -23 86 -23 0 1
rlabel polysilicon 86 -29 86 -29 0 3
rlabel polysilicon 96 -23 96 -23 0 2
rlabel polysilicon 93 -29 93 -29 0 3
rlabel polysilicon 100 -23 100 -23 0 1
rlabel polysilicon 100 -29 100 -29 0 3
rlabel polysilicon 107 -23 107 -23 0 1
rlabel polysilicon 110 -23 110 -23 0 2
rlabel polysilicon 117 -23 117 -23 0 2
rlabel polysilicon 121 -23 121 -23 0 1
rlabel polysilicon 121 -29 121 -29 0 3
rlabel polysilicon 128 -23 128 -23 0 1
rlabel polysilicon 128 -29 128 -29 0 3
rlabel polysilicon 135 -23 135 -23 0 1
rlabel polysilicon 135 -29 135 -29 0 3
rlabel polysilicon 142 -23 142 -23 0 1
rlabel polysilicon 142 -29 142 -29 0 3
rlabel polysilicon 159 -29 159 -29 0 4
rlabel polysilicon 264 -29 264 -29 0 4
rlabel polysilicon 30 -50 30 -50 0 3
rlabel polysilicon 40 -50 40 -50 0 4
rlabel polysilicon 44 -44 44 -44 0 1
rlabel polysilicon 44 -50 44 -50 0 3
rlabel polysilicon 51 -44 51 -44 0 1
rlabel polysilicon 51 -50 51 -50 0 3
rlabel polysilicon 58 -44 58 -44 0 1
rlabel polysilicon 61 -44 61 -44 0 2
rlabel polysilicon 58 -50 58 -50 0 3
rlabel polysilicon 61 -50 61 -50 0 4
rlabel polysilicon 65 -44 65 -44 0 1
rlabel polysilicon 65 -50 65 -50 0 3
rlabel polysilicon 72 -44 72 -44 0 1
rlabel polysilicon 75 -44 75 -44 0 2
rlabel polysilicon 79 -44 79 -44 0 1
rlabel polysilicon 79 -50 79 -50 0 3
rlabel polysilicon 86 -44 86 -44 0 1
rlabel polysilicon 86 -50 86 -50 0 3
rlabel polysilicon 89 -50 89 -50 0 4
rlabel polysilicon 93 -44 93 -44 0 1
rlabel polysilicon 93 -50 93 -50 0 3
rlabel polysilicon 100 -44 100 -44 0 1
rlabel polysilicon 100 -50 100 -50 0 3
rlabel polysilicon 107 -44 107 -44 0 1
rlabel polysilicon 107 -50 107 -50 0 3
rlabel polysilicon 114 -50 114 -50 0 3
rlabel polysilicon 128 -44 128 -44 0 1
rlabel polysilicon 131 -44 131 -44 0 2
rlabel polysilicon 135 -44 135 -44 0 1
rlabel polysilicon 135 -50 135 -50 0 3
rlabel polysilicon 142 -44 142 -44 0 1
rlabel polysilicon 142 -50 142 -50 0 3
rlabel polysilicon 149 -44 149 -44 0 1
rlabel polysilicon 152 -50 152 -50 0 4
rlabel polysilicon 163 -44 163 -44 0 1
rlabel polysilicon 166 -44 166 -44 0 2
rlabel polysilicon 163 -50 163 -50 0 3
rlabel polysilicon 170 -44 170 -44 0 1
rlabel polysilicon 170 -50 170 -50 0 3
rlabel polysilicon 177 -44 177 -44 0 1
rlabel polysilicon 177 -50 177 -50 0 3
rlabel polysilicon 233 -50 233 -50 0 3
rlabel polysilicon 236 -50 236 -50 0 4
rlabel polysilicon 247 -44 247 -44 0 1
rlabel polysilicon 247 -50 247 -50 0 3
rlabel polysilicon 2 -67 2 -67 0 1
rlabel polysilicon 2 -73 2 -73 0 3
rlabel polysilicon 19 -73 19 -73 0 4
rlabel polysilicon 23 -67 23 -67 0 1
rlabel polysilicon 23 -73 23 -73 0 3
rlabel polysilicon 33 -67 33 -67 0 2
rlabel polysilicon 30 -73 30 -73 0 3
rlabel polysilicon 37 -67 37 -67 0 1
rlabel polysilicon 44 -67 44 -67 0 1
rlabel polysilicon 44 -73 44 -73 0 3
rlabel polysilicon 51 -67 51 -67 0 1
rlabel polysilicon 51 -73 51 -73 0 3
rlabel polysilicon 58 -67 58 -67 0 1
rlabel polysilicon 58 -73 58 -73 0 3
rlabel polysilicon 65 -67 65 -67 0 1
rlabel polysilicon 65 -73 65 -73 0 3
rlabel polysilicon 72 -67 72 -67 0 1
rlabel polysilicon 75 -67 75 -67 0 2
rlabel polysilicon 72 -73 72 -73 0 3
rlabel polysilicon 79 -73 79 -73 0 3
rlabel polysilicon 86 -67 86 -67 0 1
rlabel polysilicon 93 -67 93 -67 0 1
rlabel polysilicon 96 -67 96 -67 0 2
rlabel polysilicon 93 -73 93 -73 0 3
rlabel polysilicon 100 -67 100 -67 0 1
rlabel polysilicon 100 -73 100 -73 0 3
rlabel polysilicon 107 -67 107 -67 0 1
rlabel polysilicon 107 -73 107 -73 0 3
rlabel polysilicon 117 -67 117 -67 0 2
rlabel polysilicon 117 -73 117 -73 0 4
rlabel polysilicon 121 -67 121 -67 0 1
rlabel polysilicon 121 -73 121 -73 0 3
rlabel polysilicon 128 -67 128 -67 0 1
rlabel polysilicon 128 -73 128 -73 0 3
rlabel polysilicon 135 -67 135 -67 0 1
rlabel polysilicon 138 -67 138 -67 0 2
rlabel polysilicon 135 -73 135 -73 0 3
rlabel polysilicon 142 -67 142 -67 0 1
rlabel polysilicon 142 -73 142 -73 0 3
rlabel polysilicon 149 -67 149 -67 0 1
rlabel polysilicon 149 -73 149 -73 0 3
rlabel polysilicon 156 -67 156 -67 0 1
rlabel polysilicon 156 -73 156 -73 0 3
rlabel polysilicon 163 -67 163 -67 0 1
rlabel polysilicon 163 -73 163 -73 0 3
rlabel polysilicon 170 -67 170 -67 0 1
rlabel polysilicon 173 -73 173 -73 0 4
rlabel polysilicon 177 -67 177 -67 0 1
rlabel polysilicon 177 -73 177 -73 0 3
rlabel polysilicon 184 -67 184 -67 0 1
rlabel polysilicon 184 -73 184 -73 0 3
rlabel polysilicon 191 -67 191 -67 0 1
rlabel polysilicon 194 -67 194 -67 0 2
rlabel polysilicon 191 -73 191 -73 0 3
rlabel polysilicon 198 -67 198 -67 0 1
rlabel polysilicon 198 -73 198 -73 0 3
rlabel polysilicon 205 -67 205 -67 0 1
rlabel polysilicon 205 -73 205 -73 0 3
rlabel polysilicon 212 -67 212 -67 0 1
rlabel polysilicon 212 -73 212 -73 0 3
rlabel polysilicon 219 -67 219 -67 0 1
rlabel polysilicon 219 -73 219 -73 0 3
rlabel polysilicon 229 -67 229 -67 0 2
rlabel polysilicon 233 -67 233 -67 0 1
rlabel polysilicon 233 -73 233 -73 0 3
rlabel polysilicon 9 -96 9 -96 0 1
rlabel polysilicon 9 -102 9 -102 0 3
rlabel polysilicon 16 -96 16 -96 0 1
rlabel polysilicon 16 -102 16 -102 0 3
rlabel polysilicon 23 -96 23 -96 0 1
rlabel polysilicon 23 -102 23 -102 0 3
rlabel polysilicon 30 -96 30 -96 0 1
rlabel polysilicon 30 -102 30 -102 0 3
rlabel polysilicon 37 -96 37 -96 0 1
rlabel polysilicon 37 -102 37 -102 0 3
rlabel polysilicon 44 -96 44 -96 0 1
rlabel polysilicon 44 -102 44 -102 0 3
rlabel polysilicon 51 -96 51 -96 0 1
rlabel polysilicon 54 -96 54 -96 0 2
rlabel polysilicon 58 -96 58 -96 0 1
rlabel polysilicon 58 -102 58 -102 0 3
rlabel polysilicon 68 -96 68 -96 0 2
rlabel polysilicon 65 -102 65 -102 0 3
rlabel polysilicon 68 -102 68 -102 0 4
rlabel polysilicon 72 -96 72 -96 0 1
rlabel polysilicon 72 -102 72 -102 0 3
rlabel polysilicon 79 -96 79 -96 0 1
rlabel polysilicon 79 -102 79 -102 0 3
rlabel polysilicon 86 -96 86 -96 0 1
rlabel polysilicon 86 -102 86 -102 0 3
rlabel polysilicon 93 -96 93 -96 0 1
rlabel polysilicon 96 -96 96 -96 0 2
rlabel polysilicon 96 -102 96 -102 0 4
rlabel polysilicon 100 -96 100 -96 0 1
rlabel polysilicon 100 -102 100 -102 0 3
rlabel polysilicon 107 -96 107 -96 0 1
rlabel polysilicon 107 -102 107 -102 0 3
rlabel polysilicon 114 -96 114 -96 0 1
rlabel polysilicon 114 -102 114 -102 0 3
rlabel polysilicon 124 -96 124 -96 0 2
rlabel polysilicon 121 -102 121 -102 0 3
rlabel polysilicon 124 -102 124 -102 0 4
rlabel polysilicon 128 -96 128 -96 0 1
rlabel polysilicon 131 -96 131 -96 0 2
rlabel polysilicon 135 -96 135 -96 0 1
rlabel polysilicon 135 -102 135 -102 0 3
rlabel polysilicon 138 -102 138 -102 0 4
rlabel polysilicon 145 -96 145 -96 0 2
rlabel polysilicon 142 -102 142 -102 0 3
rlabel polysilicon 149 -96 149 -96 0 1
rlabel polysilicon 149 -102 149 -102 0 3
rlabel polysilicon 152 -102 152 -102 0 4
rlabel polysilicon 156 -96 156 -96 0 1
rlabel polysilicon 156 -102 156 -102 0 3
rlabel polysilicon 163 -102 163 -102 0 3
rlabel polysilicon 166 -102 166 -102 0 4
rlabel polysilicon 170 -96 170 -96 0 1
rlabel polysilicon 170 -102 170 -102 0 3
rlabel polysilicon 177 -96 177 -96 0 1
rlabel polysilicon 177 -102 177 -102 0 3
rlabel polysilicon 184 -96 184 -96 0 1
rlabel polysilicon 184 -102 184 -102 0 3
rlabel polysilicon 191 -96 191 -96 0 1
rlabel polysilicon 191 -102 191 -102 0 3
rlabel polysilicon 198 -96 198 -96 0 1
rlabel polysilicon 198 -102 198 -102 0 3
rlabel polysilicon 205 -96 205 -96 0 1
rlabel polysilicon 205 -102 205 -102 0 3
rlabel polysilicon 212 -96 212 -96 0 1
rlabel polysilicon 212 -102 212 -102 0 3
rlabel polysilicon 219 -96 219 -96 0 1
rlabel polysilicon 219 -102 219 -102 0 3
rlabel polysilicon 226 -96 226 -96 0 1
rlabel polysilicon 226 -102 226 -102 0 3
rlabel polysilicon 233 -96 233 -96 0 1
rlabel polysilicon 233 -102 233 -102 0 3
rlabel polysilicon 240 -96 240 -96 0 1
rlabel polysilicon 240 -102 240 -102 0 3
rlabel polysilicon 247 -96 247 -96 0 1
rlabel polysilicon 247 -102 247 -102 0 3
rlabel polysilicon 254 -96 254 -96 0 1
rlabel polysilicon 254 -102 254 -102 0 3
rlabel polysilicon 264 -96 264 -96 0 2
rlabel polysilicon 261 -102 261 -102 0 3
rlabel polysilicon 268 -102 268 -102 0 3
rlabel polysilicon 282 -96 282 -96 0 1
rlabel polysilicon 282 -102 282 -102 0 3
rlabel polysilicon 9 -129 9 -129 0 1
rlabel polysilicon 9 -135 9 -135 0 3
rlabel polysilicon 16 -129 16 -129 0 1
rlabel polysilicon 16 -135 16 -135 0 3
rlabel polysilicon 23 -129 23 -129 0 1
rlabel polysilicon 23 -135 23 -135 0 3
rlabel polysilicon 33 -129 33 -129 0 2
rlabel polysilicon 30 -135 30 -135 0 3
rlabel polysilicon 33 -135 33 -135 0 4
rlabel polysilicon 37 -129 37 -129 0 1
rlabel polysilicon 37 -135 37 -135 0 3
rlabel polysilicon 40 -135 40 -135 0 4
rlabel polysilicon 47 -129 47 -129 0 2
rlabel polysilicon 51 -129 51 -129 0 1
rlabel polysilicon 51 -135 51 -135 0 3
rlabel polysilicon 58 -129 58 -129 0 1
rlabel polysilicon 58 -135 58 -135 0 3
rlabel polysilicon 65 -129 65 -129 0 1
rlabel polysilicon 65 -135 65 -135 0 3
rlabel polysilicon 72 -135 72 -135 0 3
rlabel polysilicon 79 -129 79 -129 0 1
rlabel polysilicon 79 -135 79 -135 0 3
rlabel polysilicon 86 -129 86 -129 0 1
rlabel polysilicon 86 -135 86 -135 0 3
rlabel polysilicon 93 -129 93 -129 0 1
rlabel polysilicon 93 -135 93 -135 0 3
rlabel polysilicon 96 -135 96 -135 0 4
rlabel polysilicon 100 -129 100 -129 0 1
rlabel polysilicon 100 -135 100 -135 0 3
rlabel polysilicon 110 -129 110 -129 0 2
rlabel polysilicon 107 -135 107 -135 0 3
rlabel polysilicon 110 -135 110 -135 0 4
rlabel polysilicon 114 -129 114 -129 0 1
rlabel polysilicon 117 -129 117 -129 0 2
rlabel polysilicon 114 -135 114 -135 0 3
rlabel polysilicon 117 -135 117 -135 0 4
rlabel polysilicon 121 -129 121 -129 0 1
rlabel polysilicon 121 -135 121 -135 0 3
rlabel polysilicon 128 -129 128 -129 0 1
rlabel polysilicon 128 -135 128 -135 0 3
rlabel polysilicon 135 -129 135 -129 0 1
rlabel polysilicon 135 -135 135 -135 0 3
rlabel polysilicon 138 -135 138 -135 0 4
rlabel polysilicon 142 -129 142 -129 0 1
rlabel polysilicon 142 -135 142 -135 0 3
rlabel polysilicon 149 -135 149 -135 0 3
rlabel polysilicon 159 -135 159 -135 0 4
rlabel polysilicon 163 -129 163 -129 0 1
rlabel polysilicon 163 -135 163 -135 0 3
rlabel polysilicon 173 -129 173 -129 0 2
rlabel polysilicon 177 -129 177 -129 0 1
rlabel polysilicon 180 -135 180 -135 0 4
rlabel polysilicon 187 -129 187 -129 0 2
rlabel polysilicon 184 -135 184 -135 0 3
rlabel polysilicon 191 -129 191 -129 0 1
rlabel polysilicon 191 -135 191 -135 0 3
rlabel polysilicon 198 -129 198 -129 0 1
rlabel polysilicon 198 -135 198 -135 0 3
rlabel polysilicon 208 -129 208 -129 0 2
rlabel polysilicon 208 -135 208 -135 0 4
rlabel polysilicon 212 -129 212 -129 0 1
rlabel polysilicon 212 -135 212 -135 0 3
rlabel polysilicon 219 -129 219 -129 0 1
rlabel polysilicon 219 -135 219 -135 0 3
rlabel polysilicon 226 -129 226 -129 0 1
rlabel polysilicon 226 -135 226 -135 0 3
rlabel polysilicon 233 -129 233 -129 0 1
rlabel polysilicon 233 -135 233 -135 0 3
rlabel polysilicon 296 -129 296 -129 0 1
rlabel polysilicon 296 -135 296 -135 0 3
rlabel polysilicon 2 -172 2 -172 0 1
rlabel polysilicon 2 -178 2 -178 0 3
rlabel polysilicon 9 -172 9 -172 0 1
rlabel polysilicon 9 -178 9 -178 0 3
rlabel polysilicon 16 -172 16 -172 0 1
rlabel polysilicon 16 -178 16 -178 0 3
rlabel polysilicon 23 -172 23 -172 0 1
rlabel polysilicon 23 -178 23 -178 0 3
rlabel polysilicon 33 -178 33 -178 0 4
rlabel polysilicon 37 -172 37 -172 0 1
rlabel polysilicon 37 -178 37 -178 0 3
rlabel polysilicon 44 -172 44 -172 0 1
rlabel polysilicon 44 -178 44 -178 0 3
rlabel polysilicon 51 -172 51 -172 0 1
rlabel polysilicon 54 -172 54 -172 0 2
rlabel polysilicon 58 -172 58 -172 0 1
rlabel polysilicon 58 -178 58 -178 0 3
rlabel polysilicon 65 -178 65 -178 0 3
rlabel polysilicon 68 -178 68 -178 0 4
rlabel polysilicon 72 -172 72 -172 0 1
rlabel polysilicon 72 -178 72 -178 0 3
rlabel polysilicon 79 -172 79 -172 0 1
rlabel polysilicon 79 -178 79 -178 0 3
rlabel polysilicon 86 -172 86 -172 0 1
rlabel polysilicon 89 -172 89 -172 0 2
rlabel polysilicon 86 -178 86 -178 0 3
rlabel polysilicon 89 -178 89 -178 0 4
rlabel polysilicon 93 -172 93 -172 0 1
rlabel polysilicon 93 -178 93 -178 0 3
rlabel polysilicon 96 -178 96 -178 0 4
rlabel polysilicon 100 -172 100 -172 0 1
rlabel polysilicon 103 -172 103 -172 0 2
rlabel polysilicon 100 -178 100 -178 0 3
rlabel polysilicon 103 -178 103 -178 0 4
rlabel polysilicon 107 -172 107 -172 0 1
rlabel polysilicon 107 -178 107 -178 0 3
rlabel polysilicon 110 -178 110 -178 0 4
rlabel polysilicon 114 -172 114 -172 0 1
rlabel polysilicon 117 -172 117 -172 0 2
rlabel polysilicon 114 -178 114 -178 0 3
rlabel polysilicon 117 -178 117 -178 0 4
rlabel polysilicon 124 -172 124 -172 0 2
rlabel polysilicon 121 -178 121 -178 0 3
rlabel polysilicon 128 -172 128 -172 0 1
rlabel polysilicon 131 -172 131 -172 0 2
rlabel polysilicon 128 -178 128 -178 0 3
rlabel polysilicon 131 -178 131 -178 0 4
rlabel polysilicon 135 -172 135 -172 0 1
rlabel polysilicon 138 -172 138 -172 0 2
rlabel polysilicon 135 -178 135 -178 0 3
rlabel polysilicon 142 -172 142 -172 0 1
rlabel polysilicon 142 -178 142 -178 0 3
rlabel polysilicon 149 -172 149 -172 0 1
rlabel polysilicon 152 -172 152 -172 0 2
rlabel polysilicon 152 -178 152 -178 0 4
rlabel polysilicon 156 -172 156 -172 0 1
rlabel polysilicon 156 -178 156 -178 0 3
rlabel polysilicon 163 -172 163 -172 0 1
rlabel polysilicon 163 -178 163 -178 0 3
rlabel polysilicon 170 -172 170 -172 0 1
rlabel polysilicon 170 -178 170 -178 0 3
rlabel polysilicon 177 -172 177 -172 0 1
rlabel polysilicon 177 -178 177 -178 0 3
rlabel polysilicon 184 -172 184 -172 0 1
rlabel polysilicon 184 -178 184 -178 0 3
rlabel polysilicon 191 -172 191 -172 0 1
rlabel polysilicon 191 -178 191 -178 0 3
rlabel polysilicon 198 -172 198 -172 0 1
rlabel polysilicon 198 -178 198 -178 0 3
rlabel polysilicon 205 -172 205 -172 0 1
rlabel polysilicon 205 -178 205 -178 0 3
rlabel polysilicon 212 -172 212 -172 0 1
rlabel polysilicon 212 -178 212 -178 0 3
rlabel polysilicon 219 -172 219 -172 0 1
rlabel polysilicon 219 -178 219 -178 0 3
rlabel polysilicon 226 -172 226 -172 0 1
rlabel polysilicon 226 -178 226 -178 0 3
rlabel polysilicon 233 -172 233 -172 0 1
rlabel polysilicon 233 -178 233 -178 0 3
rlabel polysilicon 240 -172 240 -172 0 1
rlabel polysilicon 240 -178 240 -178 0 3
rlabel polysilicon 247 -172 247 -172 0 1
rlabel polysilicon 247 -178 247 -178 0 3
rlabel polysilicon 254 -172 254 -172 0 1
rlabel polysilicon 254 -178 254 -178 0 3
rlabel polysilicon 261 -172 261 -172 0 1
rlabel polysilicon 261 -178 261 -178 0 3
rlabel polysilicon 268 -172 268 -172 0 1
rlabel polysilicon 268 -178 268 -178 0 3
rlabel polysilicon 275 -172 275 -172 0 1
rlabel polysilicon 275 -178 275 -178 0 3
rlabel polysilicon 282 -172 282 -172 0 1
rlabel polysilicon 282 -178 282 -178 0 3
rlabel polysilicon 30 -211 30 -211 0 1
rlabel polysilicon 30 -217 30 -217 0 3
rlabel polysilicon 37 -211 37 -211 0 1
rlabel polysilicon 37 -217 37 -217 0 3
rlabel polysilicon 44 -211 44 -211 0 1
rlabel polysilicon 44 -217 44 -217 0 3
rlabel polysilicon 54 -211 54 -211 0 2
rlabel polysilicon 51 -217 51 -217 0 3
rlabel polysilicon 61 -211 61 -211 0 2
rlabel polysilicon 61 -217 61 -217 0 4
rlabel polysilicon 65 -211 65 -211 0 1
rlabel polysilicon 65 -217 65 -217 0 3
rlabel polysilicon 75 -217 75 -217 0 4
rlabel polysilicon 79 -211 79 -211 0 1
rlabel polysilicon 79 -217 79 -217 0 3
rlabel polysilicon 86 -211 86 -211 0 1
rlabel polysilicon 89 -211 89 -211 0 2
rlabel polysilicon 86 -217 86 -217 0 3
rlabel polysilicon 96 -211 96 -211 0 2
rlabel polysilicon 93 -217 93 -217 0 3
rlabel polysilicon 100 -211 100 -211 0 1
rlabel polysilicon 100 -217 100 -217 0 3
rlabel polysilicon 110 -211 110 -211 0 2
rlabel polysilicon 107 -217 107 -217 0 3
rlabel polysilicon 110 -217 110 -217 0 4
rlabel polysilicon 114 -211 114 -211 0 1
rlabel polysilicon 114 -217 114 -217 0 3
rlabel polysilicon 121 -211 121 -211 0 1
rlabel polysilicon 121 -217 121 -217 0 3
rlabel polysilicon 128 -211 128 -211 0 1
rlabel polysilicon 131 -217 131 -217 0 4
rlabel polysilicon 135 -211 135 -211 0 1
rlabel polysilicon 135 -217 135 -217 0 3
rlabel polysilicon 142 -211 142 -211 0 1
rlabel polysilicon 145 -211 145 -211 0 2
rlabel polysilicon 149 -211 149 -211 0 1
rlabel polysilicon 152 -211 152 -211 0 2
rlabel polysilicon 152 -217 152 -217 0 4
rlabel polysilicon 156 -211 156 -211 0 1
rlabel polysilicon 156 -217 156 -217 0 3
rlabel polysilicon 163 -211 163 -211 0 1
rlabel polysilicon 166 -211 166 -211 0 2
rlabel polysilicon 166 -217 166 -217 0 4
rlabel polysilicon 170 -217 170 -217 0 3
rlabel polysilicon 173 -217 173 -217 0 4
rlabel polysilicon 177 -211 177 -211 0 1
rlabel polysilicon 177 -217 177 -217 0 3
rlabel polysilicon 184 -211 184 -211 0 1
rlabel polysilicon 184 -217 184 -217 0 3
rlabel polysilicon 191 -211 191 -211 0 1
rlabel polysilicon 191 -217 191 -217 0 3
rlabel polysilicon 198 -211 198 -211 0 1
rlabel polysilicon 198 -217 198 -217 0 3
rlabel polysilicon 205 -211 205 -211 0 1
rlabel polysilicon 205 -217 205 -217 0 3
rlabel polysilicon 219 -211 219 -211 0 1
rlabel polysilicon 222 -211 222 -211 0 2
rlabel polysilicon 219 -217 219 -217 0 3
rlabel polysilicon 222 -217 222 -217 0 4
rlabel polysilicon 226 -211 226 -211 0 1
rlabel polysilicon 226 -217 226 -217 0 3
rlabel polysilicon 9 -248 9 -248 0 1
rlabel polysilicon 9 -254 9 -254 0 3
rlabel polysilicon 16 -248 16 -248 0 1
rlabel polysilicon 16 -254 16 -254 0 3
rlabel polysilicon 23 -248 23 -248 0 1
rlabel polysilicon 23 -254 23 -254 0 3
rlabel polysilicon 30 -248 30 -248 0 1
rlabel polysilicon 33 -248 33 -248 0 2
rlabel polysilicon 37 -248 37 -248 0 1
rlabel polysilicon 37 -254 37 -254 0 3
rlabel polysilicon 47 -248 47 -248 0 2
rlabel polysilicon 47 -254 47 -254 0 4
rlabel polysilicon 54 -248 54 -248 0 2
rlabel polysilicon 51 -254 51 -254 0 3
rlabel polysilicon 61 -248 61 -248 0 2
rlabel polysilicon 58 -254 58 -254 0 3
rlabel polysilicon 65 -248 65 -248 0 1
rlabel polysilicon 65 -254 65 -254 0 3
rlabel polysilicon 72 -248 72 -248 0 1
rlabel polysilicon 72 -254 72 -254 0 3
rlabel polysilicon 79 -248 79 -248 0 1
rlabel polysilicon 79 -254 79 -254 0 3
rlabel polysilicon 89 -248 89 -248 0 2
rlabel polysilicon 86 -254 86 -254 0 3
rlabel polysilicon 89 -254 89 -254 0 4
rlabel polysilicon 93 -248 93 -248 0 1
rlabel polysilicon 93 -254 93 -254 0 3
rlabel polysilicon 100 -248 100 -248 0 1
rlabel polysilicon 100 -254 100 -254 0 3
rlabel polysilicon 110 -248 110 -248 0 2
rlabel polysilicon 110 -254 110 -254 0 4
rlabel polysilicon 114 -248 114 -248 0 1
rlabel polysilicon 114 -254 114 -254 0 3
rlabel polysilicon 121 -248 121 -248 0 1
rlabel polysilicon 121 -254 121 -254 0 3
rlabel polysilicon 128 -248 128 -248 0 1
rlabel polysilicon 128 -254 128 -254 0 3
rlabel polysilicon 135 -248 135 -248 0 1
rlabel polysilicon 138 -248 138 -248 0 2
rlabel polysilicon 135 -254 135 -254 0 3
rlabel polysilicon 138 -254 138 -254 0 4
rlabel polysilicon 145 -248 145 -248 0 2
rlabel polysilicon 142 -254 142 -254 0 3
rlabel polysilicon 149 -248 149 -248 0 1
rlabel polysilicon 152 -248 152 -248 0 2
rlabel polysilicon 149 -254 149 -254 0 3
rlabel polysilicon 152 -254 152 -254 0 4
rlabel polysilicon 156 -248 156 -248 0 1
rlabel polysilicon 156 -254 156 -254 0 3
rlabel polysilicon 163 -248 163 -248 0 1
rlabel polysilicon 163 -254 163 -254 0 3
rlabel polysilicon 170 -248 170 -248 0 1
rlabel polysilicon 170 -254 170 -254 0 3
rlabel polysilicon 177 -248 177 -248 0 1
rlabel polysilicon 177 -254 177 -254 0 3
rlabel polysilicon 184 -248 184 -248 0 1
rlabel polysilicon 184 -254 184 -254 0 3
rlabel polysilicon 191 -248 191 -248 0 1
rlabel polysilicon 191 -254 191 -254 0 3
rlabel polysilicon 198 -248 198 -248 0 1
rlabel polysilicon 198 -254 198 -254 0 3
rlabel polysilicon 205 -248 205 -248 0 1
rlabel polysilicon 205 -254 205 -254 0 3
rlabel polysilicon 212 -248 212 -248 0 1
rlabel polysilicon 212 -254 212 -254 0 3
rlabel polysilicon 219 -248 219 -248 0 1
rlabel polysilicon 219 -254 219 -254 0 3
rlabel polysilicon 226 -248 226 -248 0 1
rlabel polysilicon 226 -254 226 -254 0 3
rlabel polysilicon 233 -248 233 -248 0 1
rlabel polysilicon 236 -254 236 -254 0 4
rlabel polysilicon 240 -248 240 -248 0 1
rlabel polysilicon 240 -254 240 -254 0 3
rlabel polysilicon 247 -248 247 -248 0 1
rlabel polysilicon 247 -254 247 -254 0 3
rlabel polysilicon 254 -248 254 -248 0 1
rlabel polysilicon 254 -254 254 -254 0 3
rlabel polysilicon 261 -248 261 -248 0 1
rlabel polysilicon 261 -254 261 -254 0 3
rlabel polysilicon 268 -248 268 -248 0 1
rlabel polysilicon 275 -248 275 -248 0 1
rlabel polysilicon 278 -248 278 -248 0 2
rlabel polysilicon 296 -248 296 -248 0 1
rlabel polysilicon 296 -254 296 -254 0 3
rlabel polysilicon 2 -293 2 -293 0 3
rlabel polysilicon 9 -287 9 -287 0 1
rlabel polysilicon 9 -293 9 -293 0 3
rlabel polysilicon 16 -287 16 -287 0 1
rlabel polysilicon 16 -293 16 -293 0 3
rlabel polysilicon 23 -287 23 -287 0 1
rlabel polysilicon 26 -287 26 -287 0 2
rlabel polysilicon 33 -287 33 -287 0 2
rlabel polysilicon 37 -293 37 -293 0 3
rlabel polysilicon 44 -287 44 -287 0 1
rlabel polysilicon 44 -293 44 -293 0 3
rlabel polysilicon 51 -287 51 -287 0 1
rlabel polysilicon 58 -287 58 -287 0 1
rlabel polysilicon 58 -293 58 -293 0 3
rlabel polysilicon 65 -287 65 -287 0 1
rlabel polysilicon 65 -293 65 -293 0 3
rlabel polysilicon 75 -287 75 -287 0 2
rlabel polysilicon 72 -293 72 -293 0 3
rlabel polysilicon 75 -293 75 -293 0 4
rlabel polysilicon 79 -287 79 -287 0 1
rlabel polysilicon 79 -293 79 -293 0 3
rlabel polysilicon 82 -293 82 -293 0 4
rlabel polysilicon 86 -287 86 -287 0 1
rlabel polysilicon 89 -287 89 -287 0 2
rlabel polysilicon 89 -293 89 -293 0 4
rlabel polysilicon 93 -293 93 -293 0 3
rlabel polysilicon 96 -293 96 -293 0 4
rlabel polysilicon 100 -287 100 -287 0 1
rlabel polysilicon 100 -293 100 -293 0 3
rlabel polysilicon 107 -287 107 -287 0 1
rlabel polysilicon 107 -293 107 -293 0 3
rlabel polysilicon 114 -287 114 -287 0 1
rlabel polysilicon 114 -293 114 -293 0 3
rlabel polysilicon 121 -287 121 -287 0 1
rlabel polysilicon 121 -293 121 -293 0 3
rlabel polysilicon 128 -287 128 -287 0 1
rlabel polysilicon 128 -293 128 -293 0 3
rlabel polysilicon 135 -287 135 -287 0 1
rlabel polysilicon 135 -293 135 -293 0 3
rlabel polysilicon 142 -287 142 -287 0 1
rlabel polysilicon 145 -287 145 -287 0 2
rlabel polysilicon 142 -293 142 -293 0 3
rlabel polysilicon 145 -293 145 -293 0 4
rlabel polysilicon 149 -287 149 -287 0 1
rlabel polysilicon 149 -293 149 -293 0 3
rlabel polysilicon 156 -287 156 -287 0 1
rlabel polysilicon 156 -293 156 -293 0 3
rlabel polysilicon 163 -287 163 -287 0 1
rlabel polysilicon 163 -293 163 -293 0 3
rlabel polysilicon 170 -287 170 -287 0 1
rlabel polysilicon 170 -293 170 -293 0 3
rlabel polysilicon 177 -287 177 -287 0 1
rlabel polysilicon 180 -287 180 -287 0 2
rlabel polysilicon 177 -293 177 -293 0 3
rlabel polysilicon 184 -287 184 -287 0 1
rlabel polysilicon 184 -293 184 -293 0 3
rlabel polysilicon 191 -287 191 -287 0 1
rlabel polysilicon 191 -293 191 -293 0 3
rlabel polysilicon 201 -287 201 -287 0 2
rlabel polysilicon 205 -287 205 -287 0 1
rlabel polysilicon 205 -293 205 -293 0 3
rlabel polysilicon 212 -287 212 -287 0 1
rlabel polysilicon 212 -293 212 -293 0 3
rlabel polysilicon 219 -287 219 -287 0 1
rlabel polysilicon 219 -293 219 -293 0 3
rlabel polysilicon 226 -287 226 -287 0 1
rlabel polysilicon 226 -293 226 -293 0 3
rlabel polysilicon 233 -287 233 -287 0 1
rlabel polysilicon 233 -293 233 -293 0 3
rlabel polysilicon 240 -287 240 -287 0 1
rlabel polysilicon 240 -293 240 -293 0 3
rlabel polysilicon 247 -293 247 -293 0 3
rlabel polysilicon 250 -293 250 -293 0 4
rlabel polysilicon 254 -287 254 -287 0 1
rlabel polysilicon 254 -293 254 -293 0 3
rlabel polysilicon 261 -287 261 -287 0 1
rlabel polysilicon 261 -293 261 -293 0 3
rlabel polysilicon 271 -287 271 -287 0 2
rlabel polysilicon 271 -293 271 -293 0 4
rlabel polysilicon 275 -287 275 -287 0 1
rlabel polysilicon 275 -293 275 -293 0 3
rlabel polysilicon 2 -324 2 -324 0 1
rlabel polysilicon 5 -324 5 -324 0 2
rlabel polysilicon 9 -324 9 -324 0 1
rlabel polysilicon 9 -330 9 -330 0 3
rlabel polysilicon 16 -324 16 -324 0 1
rlabel polysilicon 16 -330 16 -330 0 3
rlabel polysilicon 23 -324 23 -324 0 1
rlabel polysilicon 23 -330 23 -330 0 3
rlabel polysilicon 30 -324 30 -324 0 1
rlabel polysilicon 30 -330 30 -330 0 3
rlabel polysilicon 37 -324 37 -324 0 1
rlabel polysilicon 40 -324 40 -324 0 2
rlabel polysilicon 40 -330 40 -330 0 4
rlabel polysilicon 47 -324 47 -324 0 2
rlabel polysilicon 44 -330 44 -330 0 3
rlabel polysilicon 51 -324 51 -324 0 1
rlabel polysilicon 51 -330 51 -330 0 3
rlabel polysilicon 58 -324 58 -324 0 1
rlabel polysilicon 58 -330 58 -330 0 3
rlabel polysilicon 65 -324 65 -324 0 1
rlabel polysilicon 65 -330 65 -330 0 3
rlabel polysilicon 75 -324 75 -324 0 2
rlabel polysilicon 72 -330 72 -330 0 3
rlabel polysilicon 75 -330 75 -330 0 4
rlabel polysilicon 79 -324 79 -324 0 1
rlabel polysilicon 79 -330 79 -330 0 3
rlabel polysilicon 89 -324 89 -324 0 2
rlabel polysilicon 86 -330 86 -330 0 3
rlabel polysilicon 93 -324 93 -324 0 1
rlabel polysilicon 93 -330 93 -330 0 3
rlabel polysilicon 96 -330 96 -330 0 4
rlabel polysilicon 100 -324 100 -324 0 1
rlabel polysilicon 103 -324 103 -324 0 2
rlabel polysilicon 100 -330 100 -330 0 3
rlabel polysilicon 103 -330 103 -330 0 4
rlabel polysilicon 107 -324 107 -324 0 1
rlabel polysilicon 107 -330 107 -330 0 3
rlabel polysilicon 114 -324 114 -324 0 1
rlabel polysilicon 117 -324 117 -324 0 2
rlabel polysilicon 114 -330 114 -330 0 3
rlabel polysilicon 117 -330 117 -330 0 4
rlabel polysilicon 121 -324 121 -324 0 1
rlabel polysilicon 121 -330 121 -330 0 3
rlabel polysilicon 128 -324 128 -324 0 1
rlabel polysilicon 131 -324 131 -324 0 2
rlabel polysilicon 128 -330 128 -330 0 3
rlabel polysilicon 131 -330 131 -330 0 4
rlabel polysilicon 135 -324 135 -324 0 1
rlabel polysilicon 135 -330 135 -330 0 3
rlabel polysilicon 142 -324 142 -324 0 1
rlabel polysilicon 145 -324 145 -324 0 2
rlabel polysilicon 149 -324 149 -324 0 1
rlabel polysilicon 149 -330 149 -330 0 3
rlabel polysilicon 156 -324 156 -324 0 1
rlabel polysilicon 156 -330 156 -330 0 3
rlabel polysilicon 163 -324 163 -324 0 1
rlabel polysilicon 163 -330 163 -330 0 3
rlabel polysilicon 170 -324 170 -324 0 1
rlabel polysilicon 170 -330 170 -330 0 3
rlabel polysilicon 177 -324 177 -324 0 1
rlabel polysilicon 177 -330 177 -330 0 3
rlabel polysilicon 184 -324 184 -324 0 1
rlabel polysilicon 184 -330 184 -330 0 3
rlabel polysilicon 191 -324 191 -324 0 1
rlabel polysilicon 191 -330 191 -330 0 3
rlabel polysilicon 198 -324 198 -324 0 1
rlabel polysilicon 198 -330 198 -330 0 3
rlabel polysilicon 205 -324 205 -324 0 1
rlabel polysilicon 205 -330 205 -330 0 3
rlabel polysilicon 212 -324 212 -324 0 1
rlabel polysilicon 212 -330 212 -330 0 3
rlabel polysilicon 222 -324 222 -324 0 2
rlabel polysilicon 219 -330 219 -330 0 3
rlabel polysilicon 226 -324 226 -324 0 1
rlabel polysilicon 226 -330 226 -330 0 3
rlabel polysilicon 2 -355 2 -355 0 1
rlabel polysilicon 23 -355 23 -355 0 1
rlabel polysilicon 23 -361 23 -361 0 3
rlabel polysilicon 30 -355 30 -355 0 1
rlabel polysilicon 30 -361 30 -361 0 3
rlabel polysilicon 37 -355 37 -355 0 1
rlabel polysilicon 37 -361 37 -361 0 3
rlabel polysilicon 44 -355 44 -355 0 1
rlabel polysilicon 51 -355 51 -355 0 1
rlabel polysilicon 58 -355 58 -355 0 1
rlabel polysilicon 61 -355 61 -355 0 2
rlabel polysilicon 58 -361 58 -361 0 3
rlabel polysilicon 68 -355 68 -355 0 2
rlabel polysilicon 68 -361 68 -361 0 4
rlabel polysilicon 72 -355 72 -355 0 1
rlabel polysilicon 72 -361 72 -361 0 3
rlabel polysilicon 79 -355 79 -355 0 1
rlabel polysilicon 79 -361 79 -361 0 3
rlabel polysilicon 86 -361 86 -361 0 3
rlabel polysilicon 96 -355 96 -355 0 2
rlabel polysilicon 96 -361 96 -361 0 4
rlabel polysilicon 100 -355 100 -355 0 1
rlabel polysilicon 100 -361 100 -361 0 3
rlabel polysilicon 107 -355 107 -355 0 1
rlabel polysilicon 107 -361 107 -361 0 3
rlabel polysilicon 114 -355 114 -355 0 1
rlabel polysilicon 114 -361 114 -361 0 3
rlabel polysilicon 117 -361 117 -361 0 4
rlabel polysilicon 121 -355 121 -355 0 1
rlabel polysilicon 121 -361 121 -361 0 3
rlabel polysilicon 128 -355 128 -355 0 1
rlabel polysilicon 128 -361 128 -361 0 3
rlabel polysilicon 135 -355 135 -355 0 1
rlabel polysilicon 135 -361 135 -361 0 3
rlabel polysilicon 142 -355 142 -355 0 1
rlabel polysilicon 142 -361 142 -361 0 3
rlabel polysilicon 149 -355 149 -355 0 1
rlabel polysilicon 149 -361 149 -361 0 3
rlabel polysilicon 159 -355 159 -355 0 2
rlabel polysilicon 156 -361 156 -361 0 3
rlabel polysilicon 159 -361 159 -361 0 4
rlabel polysilicon 163 -355 163 -355 0 1
rlabel polysilicon 163 -361 163 -361 0 3
rlabel polysilicon 170 -355 170 -355 0 1
rlabel polysilicon 170 -361 170 -361 0 3
rlabel polysilicon 177 -355 177 -355 0 1
rlabel polysilicon 177 -361 177 -361 0 3
rlabel polysilicon 184 -355 184 -355 0 1
rlabel polysilicon 184 -361 184 -361 0 3
rlabel polysilicon 191 -355 191 -355 0 1
rlabel polysilicon 191 -361 191 -361 0 3
rlabel polysilicon 198 -355 198 -355 0 1
rlabel polysilicon 198 -361 198 -361 0 3
rlabel polysilicon 208 -361 208 -361 0 4
rlabel polysilicon 215 -355 215 -355 0 2
rlabel polysilicon 212 -361 212 -361 0 3
rlabel polysilicon 12 -388 12 -388 0 2
rlabel polysilicon 16 -388 16 -388 0 1
rlabel polysilicon 16 -394 16 -394 0 3
rlabel polysilicon 23 -388 23 -388 0 1
rlabel polysilicon 23 -394 23 -394 0 3
rlabel polysilicon 30 -388 30 -388 0 1
rlabel polysilicon 30 -394 30 -394 0 3
rlabel polysilicon 37 -394 37 -394 0 3
rlabel polysilicon 40 -394 40 -394 0 4
rlabel polysilicon 44 -388 44 -388 0 1
rlabel polysilicon 47 -388 47 -388 0 2
rlabel polysilicon 51 -388 51 -388 0 1
rlabel polysilicon 54 -394 54 -394 0 4
rlabel polysilicon 58 -388 58 -388 0 1
rlabel polysilicon 58 -394 58 -394 0 3
rlabel polysilicon 65 -388 65 -388 0 1
rlabel polysilicon 65 -394 65 -394 0 3
rlabel polysilicon 72 -388 72 -388 0 1
rlabel polysilicon 72 -394 72 -394 0 3
rlabel polysilicon 79 -388 79 -388 0 1
rlabel polysilicon 79 -394 79 -394 0 3
rlabel polysilicon 86 -394 86 -394 0 3
rlabel polysilicon 89 -394 89 -394 0 4
rlabel polysilicon 96 -388 96 -388 0 2
rlabel polysilicon 96 -394 96 -394 0 4
rlabel polysilicon 100 -388 100 -388 0 1
rlabel polysilicon 100 -394 100 -394 0 3
rlabel polysilicon 107 -388 107 -388 0 1
rlabel polysilicon 110 -394 110 -394 0 4
rlabel polysilicon 114 -388 114 -388 0 1
rlabel polysilicon 114 -394 114 -394 0 3
rlabel polysilicon 117 -394 117 -394 0 4
rlabel polysilicon 121 -388 121 -388 0 1
rlabel polysilicon 121 -394 121 -394 0 3
rlabel polysilicon 128 -394 128 -394 0 3
rlabel polysilicon 131 -394 131 -394 0 4
rlabel polysilicon 138 -388 138 -388 0 2
rlabel polysilicon 138 -394 138 -394 0 4
rlabel polysilicon 142 -388 142 -388 0 1
rlabel polysilicon 142 -394 142 -394 0 3
rlabel polysilicon 152 -394 152 -394 0 4
rlabel polysilicon 156 -388 156 -388 0 1
rlabel polysilicon 156 -394 156 -394 0 3
rlabel polysilicon 163 -388 163 -388 0 1
rlabel polysilicon 163 -394 163 -394 0 3
rlabel polysilicon 170 -388 170 -388 0 1
rlabel polysilicon 170 -394 170 -394 0 3
rlabel polysilicon 177 -388 177 -388 0 1
rlabel polysilicon 177 -394 177 -394 0 3
rlabel polysilicon 184 -388 184 -388 0 1
rlabel polysilicon 184 -394 184 -394 0 3
rlabel polysilicon 187 -394 187 -394 0 4
rlabel polysilicon 191 -388 191 -388 0 1
rlabel polysilicon 191 -394 191 -394 0 3
rlabel polysilicon 198 -394 198 -394 0 3
rlabel polysilicon 205 -388 205 -388 0 1
rlabel polysilicon 205 -394 205 -394 0 3
rlabel polysilicon 212 -388 212 -388 0 1
rlabel polysilicon 212 -394 212 -394 0 3
rlabel polysilicon 222 -388 222 -388 0 2
rlabel polysilicon 226 -388 226 -388 0 1
rlabel polysilicon 226 -394 226 -394 0 3
rlabel polysilicon 12 -427 12 -427 0 4
rlabel polysilicon 19 -427 19 -427 0 4
rlabel polysilicon 26 -421 26 -421 0 2
rlabel polysilicon 30 -421 30 -421 0 1
rlabel polysilicon 30 -427 30 -427 0 3
rlabel polysilicon 44 -421 44 -421 0 1
rlabel polysilicon 47 -427 47 -427 0 4
rlabel polysilicon 54 -421 54 -421 0 2
rlabel polysilicon 61 -421 61 -421 0 2
rlabel polysilicon 61 -427 61 -427 0 4
rlabel polysilicon 65 -421 65 -421 0 1
rlabel polysilicon 65 -427 65 -427 0 3
rlabel polysilicon 72 -427 72 -427 0 3
rlabel polysilicon 75 -427 75 -427 0 4
rlabel polysilicon 79 -421 79 -421 0 1
rlabel polysilicon 82 -421 82 -421 0 2
rlabel polysilicon 79 -427 79 -427 0 3
rlabel polysilicon 89 -427 89 -427 0 4
rlabel polysilicon 93 -421 93 -421 0 1
rlabel polysilicon 96 -421 96 -421 0 2
rlabel polysilicon 96 -427 96 -427 0 4
rlabel polysilicon 100 -421 100 -421 0 1
rlabel polysilicon 100 -427 100 -427 0 3
rlabel polysilicon 107 -421 107 -421 0 1
rlabel polysilicon 107 -427 107 -427 0 3
rlabel polysilicon 114 -421 114 -421 0 1
rlabel polysilicon 114 -427 114 -427 0 3
rlabel polysilicon 121 -427 121 -427 0 3
rlabel polysilicon 124 -427 124 -427 0 4
rlabel polysilicon 128 -421 128 -421 0 1
rlabel polysilicon 128 -427 128 -427 0 3
rlabel polysilicon 135 -421 135 -421 0 1
rlabel polysilicon 142 -421 142 -421 0 1
rlabel polysilicon 142 -427 142 -427 0 3
rlabel polysilicon 149 -421 149 -421 0 1
rlabel polysilicon 149 -427 149 -427 0 3
rlabel polysilicon 156 -421 156 -421 0 1
rlabel polysilicon 156 -427 156 -427 0 3
rlabel polysilicon 187 -421 187 -421 0 2
rlabel polysilicon 198 -421 198 -421 0 1
rlabel metal2 72 1 72 1 0 net=251
rlabel metal2 100 1 100 1 0 net=593
rlabel metal2 121 1 121 1 0 net=445
rlabel metal2 51 -10 51 -10 0 net=563
rlabel metal2 68 -10 68 -10 0 net=437
rlabel metal2 75 -10 75 -10 0 net=252
rlabel metal2 82 -10 82 -10 0 net=361
rlabel metal2 128 -10 128 -10 0 net=447
rlabel metal2 128 -10 128 -10 0 net=447
rlabel metal2 44 -12 44 -12 0 net=485
rlabel metal2 86 -12 86 -12 0 net=317
rlabel metal2 96 -14 96 -14 0 net=533
rlabel metal2 100 -16 100 -16 0 net=591
rlabel metal2 107 -18 107 -18 0 net=595
rlabel metal2 107 -20 107 -20 0 net=172
rlabel metal2 44 -31 44 -31 0 net=486
rlabel metal2 93 -31 93 -31 0 net=596
rlabel metal2 159 -31 159 -31 0 net=121
rlabel metal2 247 -31 247 -31 0 net=667
rlabel metal2 44 -33 44 -33 0 net=285
rlabel metal2 86 -33 86 -33 0 net=319
rlabel metal2 107 -33 107 -33 0 net=363
rlabel metal2 128 -33 128 -33 0 net=449
rlabel metal2 51 -35 51 -35 0 net=564
rlabel metal2 86 -35 86 -35 0 net=605
rlabel metal2 51 -37 51 -37 0 net=367
rlabel metal2 100 -37 100 -37 0 net=592
rlabel metal2 131 -37 131 -37 0 net=633
rlabel metal2 72 -39 72 -39 0 net=439
rlabel metal2 135 -39 135 -39 0 net=534
rlabel metal2 72 -41 72 -41 0 net=203
rlabel metal2 135 -41 135 -41 0 net=379
rlabel metal2 2 -52 2 -52 0 net=627
rlabel metal2 65 -52 65 -52 0 net=257
rlabel metal2 65 -52 65 -52 0 net=257
rlabel metal2 75 -52 75 -52 0 net=364
rlabel metal2 121 -52 121 -52 0 net=299
rlabel metal2 212 -52 212 -52 0 net=162
rlabel metal2 233 -52 233 -52 0 net=668
rlabel metal2 23 -54 23 -54 0 net=483
rlabel metal2 37 -54 37 -54 0 net=20
rlabel metal2 51 -54 51 -54 0 net=369
rlabel metal2 135 -54 135 -54 0 net=381
rlabel metal2 170 -54 170 -54 0 net=635
rlabel metal2 233 -54 233 -54 0 net=639
rlabel metal2 30 -56 30 -56 0 net=286
rlabel metal2 51 -56 51 -56 0 net=205
rlabel metal2 89 -56 89 -56 0 net=320
rlabel metal2 96 -56 96 -56 0 net=225
rlabel metal2 135 -56 135 -56 0 net=619
rlabel metal2 44 -58 44 -58 0 net=423
rlabel metal2 93 -58 93 -58 0 net=102
rlabel metal2 138 -58 138 -58 0 net=3
rlabel metal2 177 -58 177 -58 0 net=607
rlabel metal2 58 -60 58 -60 0 net=440
rlabel metal2 142 -60 142 -60 0 net=451
rlabel metal2 152 -60 152 -60 0 net=629
rlabel metal2 86 -62 86 -62 0 net=309
rlabel metal2 163 -62 163 -62 0 net=585
rlabel metal2 58 -64 58 -64 0 net=279
rlabel metal2 100 -64 100 -64 0 net=227
rlabel metal2 170 -64 170 -64 0 net=529
rlabel metal2 2 -75 2 -75 0 net=628
rlabel metal2 58 -75 58 -75 0 net=281
rlabel metal2 117 -75 117 -75 0 net=382
rlabel metal2 173 -75 173 -75 0 net=553
rlabel metal2 264 -75 264 -75 0 net=471
rlabel metal2 9 -77 9 -77 0 net=495
rlabel metal2 86 -77 86 -77 0 net=229
rlabel metal2 107 -77 107 -77 0 net=226
rlabel metal2 149 -77 149 -77 0 net=453
rlabel metal2 184 -77 184 -77 0 net=608
rlabel metal2 219 -77 219 -77 0 net=631
rlabel metal2 16 -79 16 -79 0 net=415
rlabel metal2 100 -79 100 -79 0 net=301
rlabel metal2 128 -79 128 -79 0 net=370
rlabel metal2 156 -79 156 -79 0 net=389
rlabel metal2 198 -79 198 -79 0 net=637
rlabel metal2 37 -81 37 -81 0 net=387
rlabel metal2 72 -81 72 -81 0 net=321
rlabel metal2 177 -81 177 -81 0 net=531
rlabel metal2 44 -83 44 -83 0 net=424
rlabel metal2 107 -83 107 -83 0 net=241
rlabel metal2 128 -83 128 -83 0 net=507
rlabel metal2 30 -85 30 -85 0 net=26
rlabel metal2 51 -85 51 -85 0 net=206
rlabel metal2 131 -85 131 -85 0 net=535
rlabel metal2 198 -85 198 -85 0 net=641
rlabel metal2 23 -87 23 -87 0 net=484
rlabel metal2 51 -87 51 -87 0 net=501
rlabel metal2 205 -87 205 -87 0 net=621
rlabel metal2 19 -89 19 -89 0 net=343
rlabel metal2 58 -89 58 -89 0 net=259
rlabel metal2 79 -89 79 -89 0 net=509
rlabel metal2 93 -91 93 -91 0 net=310
rlabel metal2 163 -91 163 -91 0 net=587
rlabel metal2 135 -93 135 -93 0 net=657
rlabel metal2 9 -104 9 -104 0 net=496
rlabel metal2 149 -104 149 -104 0 net=632
rlabel metal2 268 -104 268 -104 0 net=472
rlabel metal2 16 -106 16 -106 0 net=416
rlabel metal2 58 -106 58 -106 0 net=260
rlabel metal2 79 -106 79 -106 0 net=282
rlabel metal2 121 -106 121 -106 0 net=390
rlabel metal2 163 -106 163 -106 0 net=638
rlabel metal2 16 -108 16 -108 0 net=345
rlabel metal2 33 -108 33 -108 0 net=429
rlabel metal2 58 -108 58 -108 0 net=323
rlabel metal2 79 -108 79 -108 0 net=243
rlabel metal2 117 -108 117 -108 0 net=427
rlabel metal2 124 -108 124 -108 0 net=554
rlabel metal2 23 -110 23 -110 0 net=467
rlabel metal2 37 -110 37 -110 0 net=388
rlabel metal2 65 -110 65 -110 0 net=409
rlabel metal2 135 -110 135 -110 0 net=454
rlabel metal2 173 -110 173 -110 0 net=669
rlabel metal2 9 -112 9 -112 0 net=645
rlabel metal2 86 -112 86 -112 0 net=230
rlabel metal2 152 -112 152 -112 0 net=532
rlabel metal2 68 -114 68 -114 0 net=417
rlabel metal2 93 -114 93 -114 0 net=302
rlabel metal2 163 -114 163 -114 0 net=503
rlabel metal2 198 -114 198 -114 0 net=643
rlabel metal2 198 -114 198 -114 0 net=643
rlabel metal2 208 -114 208 -114 0 net=508
rlabel metal2 96 -116 96 -116 0 net=297
rlabel metal2 142 -116 142 -116 0 net=647
rlabel metal2 219 -116 219 -116 0 net=623
rlabel metal2 100 -118 100 -118 0 net=611
rlabel metal2 142 -120 142 -120 0 net=655
rlabel metal2 177 -120 177 -120 0 net=659
rlabel metal2 138 -122 138 -122 0 net=92
rlabel metal2 184 -122 184 -122 0 net=537
rlabel metal2 187 -124 187 -124 0 net=588
rlabel metal2 205 -126 205 -126 0 net=511
rlabel metal2 9 -137 9 -137 0 net=646
rlabel metal2 40 -137 40 -137 0 net=95
rlabel metal2 121 -137 121 -137 0 net=428
rlabel metal2 159 -137 159 -137 0 net=307
rlabel metal2 212 -137 212 -137 0 net=661
rlabel metal2 9 -139 9 -139 0 net=385
rlabel metal2 96 -139 96 -139 0 net=78
rlabel metal2 117 -139 117 -139 0 net=463
rlabel metal2 219 -139 219 -139 0 net=625
rlabel metal2 16 -141 16 -141 0 net=346
rlabel metal2 44 -141 44 -141 0 net=245
rlabel metal2 86 -141 86 -141 0 net=418
rlabel metal2 117 -141 117 -141 0 net=613
rlabel metal2 16 -143 16 -143 0 net=283
rlabel metal2 103 -143 103 -143 0 net=298
rlabel metal2 131 -143 131 -143 0 net=499
rlabel metal2 226 -143 226 -143 0 net=671
rlabel metal2 23 -145 23 -145 0 net=468
rlabel metal2 51 -145 51 -145 0 net=430
rlabel metal2 58 -145 58 -145 0 net=325
rlabel metal2 58 -145 58 -145 0 net=325
rlabel metal2 72 -145 72 -145 0 net=612
rlabel metal2 124 -145 124 -145 0 net=405
rlabel metal2 2 -147 2 -147 0 net=277
rlabel metal2 72 -147 72 -147 0 net=291
rlabel metal2 138 -147 138 -147 0 net=615
rlabel metal2 23 -149 23 -149 0 net=181
rlabel metal2 138 -149 138 -149 0 net=538
rlabel metal2 37 -151 37 -151 0 net=295
rlabel metal2 149 -151 149 -151 0 net=512
rlabel metal2 79 -153 79 -153 0 net=473
rlabel metal2 149 -153 149 -153 0 net=365
rlabel metal2 163 -153 163 -153 0 net=505
rlabel metal2 86 -155 86 -155 0 net=656
rlabel metal2 163 -155 163 -155 0 net=644
rlabel metal2 110 -157 110 -157 0 net=601
rlabel metal2 114 -159 114 -159 0 net=489
rlabel metal2 170 -159 170 -159 0 net=393
rlabel metal2 135 -161 135 -161 0 net=469
rlabel metal2 177 -163 177 -163 0 net=649
rlabel metal2 180 -165 180 -165 0 net=579
rlabel metal2 184 -167 184 -167 0 net=565
rlabel metal2 65 -169 65 -169 0 net=411
rlabel metal2 2 -180 2 -180 0 net=278
rlabel metal2 131 -180 131 -180 0 net=500
rlabel metal2 222 -180 222 -180 0 net=580
rlabel metal2 9 -182 9 -182 0 net=386
rlabel metal2 135 -182 135 -182 0 net=555
rlabel metal2 135 -182 135 -182 0 net=555
rlabel metal2 145 -182 145 -182 0 net=506
rlabel metal2 16 -184 16 -184 0 net=284
rlabel metal2 58 -184 58 -184 0 net=326
rlabel metal2 149 -184 149 -184 0 net=308
rlabel metal2 219 -184 219 -184 0 net=614
rlabel metal2 23 -186 23 -186 0 net=182
rlabel metal2 79 -186 79 -186 0 net=475
rlabel metal2 79 -186 79 -186 0 net=475
rlabel metal2 96 -186 96 -186 0 net=412
rlabel metal2 191 -186 191 -186 0 net=567
rlabel metal2 226 -186 226 -186 0 net=663
rlabel metal2 30 -188 30 -188 0 net=513
rlabel metal2 100 -188 100 -188 0 net=406
rlabel metal2 33 -190 33 -190 0 net=296
rlabel metal2 44 -190 44 -190 0 net=246
rlabel metal2 142 -190 142 -190 0 net=491
rlabel metal2 37 -192 37 -192 0 net=293
rlabel metal2 107 -192 107 -192 0 net=401
rlabel metal2 44 -194 44 -194 0 net=130
rlabel metal2 152 -194 152 -194 0 net=626
rlabel metal2 61 -196 61 -196 0 net=366
rlabel metal2 166 -196 166 -196 0 net=394
rlabel metal2 65 -198 65 -198 0 net=115
rlabel metal2 103 -198 103 -198 0 net=541
rlabel metal2 152 -198 152 -198 0 net=464
rlabel metal2 65 -200 65 -200 0 net=557
rlabel metal2 89 -200 89 -200 0 net=470
rlabel metal2 86 -202 86 -202 0 net=149
rlabel metal2 177 -202 177 -202 0 net=651
rlabel metal2 100 -204 100 -204 0 net=263
rlabel metal2 177 -204 177 -204 0 net=603
rlabel metal2 110 -206 110 -206 0 net=672
rlabel metal2 93 -208 93 -208 0 net=68
rlabel metal2 114 -208 114 -208 0 net=311
rlabel metal2 156 -208 156 -208 0 net=617
rlabel metal2 23 -219 23 -219 0 net=315
rlabel metal2 173 -219 173 -219 0 net=664
rlabel metal2 233 -219 233 -219 0 net=549
rlabel metal2 275 -219 275 -219 0 net=347
rlabel metal2 16 -221 16 -221 0 net=217
rlabel metal2 198 -221 198 -221 0 net=653
rlabel metal2 30 -223 30 -223 0 net=514
rlabel metal2 37 -223 37 -223 0 net=294
rlabel metal2 89 -223 89 -223 0 net=556
rlabel metal2 138 -223 138 -223 0 net=150
rlabel metal2 184 -223 184 -223 0 net=493
rlabel metal2 205 -223 205 -223 0 net=569
rlabel metal2 30 -225 30 -225 0 net=581
rlabel metal2 37 -227 37 -227 0 net=395
rlabel metal2 72 -227 72 -227 0 net=375
rlabel metal2 93 -227 93 -227 0 net=604
rlabel metal2 184 -227 184 -227 0 net=455
rlabel metal2 44 -229 44 -229 0 net=70
rlabel metal2 54 -229 54 -229 0 net=135
rlabel metal2 212 -229 212 -229 0 net=539
rlabel metal2 222 -229 222 -229 0 net=133
rlabel metal2 47 -231 47 -231 0 net=413
rlabel metal2 191 -231 191 -231 0 net=403
rlabel metal2 93 -233 93 -233 0 net=303
rlabel metal2 114 -233 114 -233 0 net=313
rlabel metal2 131 -233 131 -233 0 net=573
rlabel metal2 100 -235 100 -235 0 net=265
rlabel metal2 121 -235 121 -235 0 net=543
rlabel metal2 61 -237 61 -237 0 net=231
rlabel metal2 107 -237 107 -237 0 net=618
rlabel metal2 65 -239 65 -239 0 net=558
rlabel metal2 135 -239 135 -239 0 net=517
rlabel metal2 65 -241 65 -241 0 net=477
rlabel metal2 110 -241 110 -241 0 net=441
rlabel metal2 9 -243 9 -243 0 net=383
rlabel metal2 145 -243 145 -243 0 net=497
rlabel metal2 149 -245 149 -245 0 net=521
rlabel metal2 9 -256 9 -256 0 net=384
rlabel metal2 79 -256 79 -256 0 net=45
rlabel metal2 219 -256 219 -256 0 net=404
rlabel metal2 240 -256 240 -256 0 net=551
rlabel metal2 275 -256 275 -256 0 net=349
rlabel metal2 9 -258 9 -258 0 net=425
rlabel metal2 44 -258 44 -258 0 net=377
rlabel metal2 110 -258 110 -258 0 net=314
rlabel metal2 135 -258 135 -258 0 net=498
rlabel metal2 219 -258 219 -258 0 net=575
rlabel metal2 16 -260 16 -260 0 net=218
rlabel metal2 138 -260 138 -260 0 net=494
rlabel metal2 240 -260 240 -260 0 net=583
rlabel metal2 16 -262 16 -262 0 net=337
rlabel metal2 142 -262 142 -262 0 net=414
rlabel metal2 184 -262 184 -262 0 net=457
rlabel metal2 184 -262 184 -262 0 net=457
rlabel metal2 23 -264 23 -264 0 net=316
rlabel metal2 89 -264 89 -264 0 net=271
rlabel metal2 135 -264 135 -264 0 net=327
rlabel metal2 145 -264 145 -264 0 net=540
rlabel metal2 247 -264 247 -264 0 net=571
rlabel metal2 23 -266 23 -266 0 net=14
rlabel metal2 58 -266 58 -266 0 net=479
rlabel metal2 107 -266 107 -266 0 net=213
rlabel metal2 26 -268 26 -268 0 net=589
rlabel metal2 47 -270 47 -270 0 net=1
rlabel metal2 152 -270 152 -270 0 net=654
rlabel metal2 51 -272 51 -272 0 net=232
rlabel metal2 156 -272 156 -272 0 net=523
rlabel metal2 65 -274 65 -274 0 net=209
rlabel metal2 93 -274 93 -274 0 net=305
rlabel metal2 114 -274 114 -274 0 net=267
rlabel metal2 170 -274 170 -274 0 net=519
rlabel metal2 114 -276 114 -276 0 net=235
rlabel metal2 170 -276 170 -276 0 net=357
rlabel metal2 149 -278 149 -278 0 net=351
rlabel metal2 191 -278 191 -278 0 net=545
rlabel metal2 121 -280 121 -280 0 net=465
rlabel metal2 121 -282 121 -282 0 net=443
rlabel metal2 37 -284 37 -284 0 net=397
rlabel metal2 2 -295 2 -295 0 net=127
rlabel metal2 23 -295 23 -295 0 net=237
rlabel metal2 121 -295 121 -295 0 net=444
rlabel metal2 135 -295 135 -295 0 net=329
rlabel metal2 135 -295 135 -295 0 net=329
rlabel metal2 142 -295 142 -295 0 net=520
rlabel metal2 222 -295 222 -295 0 net=584
rlabel metal2 247 -295 247 -295 0 net=572
rlabel metal2 261 -295 261 -295 0 net=552
rlabel metal2 30 -297 30 -297 0 net=215
rlabel metal2 142 -297 142 -297 0 net=391
rlabel metal2 205 -297 205 -297 0 net=525
rlabel metal2 250 -297 250 -297 0 net=350
rlabel metal2 16 -299 16 -299 0 net=339
rlabel metal2 156 -299 156 -299 0 net=268
rlabel metal2 205 -299 205 -299 0 net=577
rlabel metal2 37 -301 37 -301 0 net=91
rlabel metal2 156 -301 156 -301 0 net=466
rlabel metal2 9 -303 9 -303 0 net=426
rlabel metal2 40 -303 40 -303 0 net=147
rlabel metal2 51 -303 51 -303 0 net=183
rlabel metal2 145 -303 145 -303 0 net=665
rlabel metal2 2 -305 2 -305 0 net=407
rlabel metal2 44 -305 44 -305 0 net=378
rlabel metal2 100 -305 100 -305 0 net=306
rlabel metal2 170 -305 170 -305 0 net=359
rlabel metal2 170 -305 170 -305 0 net=359
rlabel metal2 177 -305 177 -305 0 net=459
rlabel metal2 58 -307 58 -307 0 net=480
rlabel metal2 82 -307 82 -307 0 net=178
rlabel metal2 93 -307 93 -307 0 net=590
rlabel metal2 58 -309 58 -309 0 net=273
rlabel metal2 163 -309 163 -309 0 net=399
rlabel metal2 16 -311 16 -311 0 net=481
rlabel metal2 149 -311 149 -311 0 net=353
rlabel metal2 65 -313 65 -313 0 net=211
rlabel metal2 65 -315 65 -315 0 net=191
rlabel metal2 103 -315 103 -315 0 net=18
rlabel metal2 72 -317 72 -317 0 net=546
rlabel metal2 75 -319 75 -319 0 net=156
rlabel metal2 100 -319 100 -319 0 net=597
rlabel metal2 75 -321 75 -321 0 net=197
rlabel metal2 2 -332 2 -332 0 net=408
rlabel metal2 16 -332 16 -332 0 net=482
rlabel metal2 72 -332 72 -332 0 net=340
rlabel metal2 114 -332 114 -332 0 net=392
rlabel metal2 23 -334 23 -334 0 net=238
rlabel metal2 96 -334 96 -334 0 net=400
rlabel metal2 198 -334 198 -334 0 net=599
rlabel metal2 30 -336 30 -336 0 net=216
rlabel metal2 107 -336 107 -336 0 net=371
rlabel metal2 135 -336 135 -336 0 net=331
rlabel metal2 149 -336 149 -336 0 net=360
rlabel metal2 177 -336 177 -336 0 net=461
rlabel metal2 177 -336 177 -336 0 net=461
rlabel metal2 184 -336 184 -336 0 net=487
rlabel metal2 30 -338 30 -338 0 net=275
rlabel metal2 96 -338 96 -338 0 net=76
rlabel metal2 135 -338 135 -338 0 net=219
rlabel metal2 163 -338 163 -338 0 net=355
rlabel metal2 163 -338 163 -338 0 net=355
rlabel metal2 170 -338 170 -338 0 net=578
rlabel metal2 23 -340 23 -340 0 net=515
rlabel metal2 93 -340 93 -340 0 net=287
rlabel metal2 156 -340 156 -340 0 net=666
rlabel metal2 37 -342 37 -342 0 net=207
rlabel metal2 191 -342 191 -342 0 net=527
rlabel metal2 40 -344 40 -344 0 net=74
rlabel metal2 100 -344 100 -344 0 net=212
rlabel metal2 44 -346 44 -346 0 net=19
rlabel metal2 79 -346 79 -346 0 net=199
rlabel metal2 114 -346 114 -346 0 net=559
rlabel metal2 44 -348 44 -348 0 net=192
rlabel metal2 121 -348 121 -348 0 net=269
rlabel metal2 51 -350 51 -350 0 net=185
rlabel metal2 51 -352 51 -352 0 net=253
rlabel metal2 12 -363 12 -363 0 net=419
rlabel metal2 23 -363 23 -363 0 net=516
rlabel metal2 65 -363 65 -363 0 net=255
rlabel metal2 86 -363 86 -363 0 net=356
rlabel metal2 184 -363 184 -363 0 net=488
rlabel metal2 23 -365 23 -365 0 net=431
rlabel metal2 72 -365 72 -365 0 net=187
rlabel metal2 72 -365 72 -365 0 net=187
rlabel metal2 100 -365 100 -365 0 net=201
rlabel metal2 100 -365 100 -365 0 net=201
rlabel metal2 114 -365 114 -365 0 net=609
rlabel metal2 30 -367 30 -367 0 net=276
rlabel metal2 117 -367 117 -367 0 net=270
rlabel metal2 138 -367 138 -367 0 net=40
rlabel metal2 30 -369 30 -369 0 net=233
rlabel metal2 58 -369 58 -369 0 net=239
rlabel metal2 121 -369 121 -369 0 net=221
rlabel metal2 142 -369 142 -369 0 net=333
rlabel metal2 184 -369 184 -369 0 net=600
rlabel metal2 37 -371 37 -371 0 net=208
rlabel metal2 191 -371 191 -371 0 net=528
rlabel metal2 96 -373 96 -373 0 net=435
rlabel metal2 79 -375 79 -375 0 net=193
rlabel metal2 114 -375 114 -375 0 net=341
rlabel metal2 149 -377 149 -377 0 net=561
rlabel metal2 156 -379 156 -379 0 net=673
rlabel metal2 128 -381 128 -381 0 net=289
rlabel metal2 159 -381 159 -381 0 net=462
rlabel metal2 107 -383 107 -383 0 net=373
rlabel metal2 107 -385 107 -385 0 net=247
rlabel metal2 23 -396 23 -396 0 net=433
rlabel metal2 152 -396 152 -396 0 net=122
rlabel metal2 198 -396 198 -396 0 net=59
rlabel metal2 198 -396 198 -396 0 net=59
rlabel metal2 26 -398 26 -398 0 net=169
rlabel metal2 131 -398 131 -398 0 net=374
rlabel metal2 30 -400 30 -400 0 net=234
rlabel metal2 54 -400 54 -400 0 net=240
rlabel metal2 79 -400 79 -400 0 net=195
rlabel metal2 110 -400 110 -400 0 net=436
rlabel metal2 16 -402 16 -402 0 net=421
rlabel metal2 40 -402 40 -402 0 net=342
rlabel metal2 54 -404 54 -404 0 net=290
rlabel metal2 37 -406 37 -406 0 net=547
rlabel metal2 61 -408 61 -408 0 net=60
rlabel metal2 82 -408 82 -408 0 net=261
rlabel metal2 135 -408 135 -408 0 net=56
rlabel metal2 86 -410 86 -410 0 net=202
rlabel metal2 117 -410 117 -410 0 net=610
rlabel metal2 89 -412 89 -412 0 net=173
rlabel metal2 100 -412 100 -412 0 net=249
rlabel metal2 187 -412 187 -412 0 net=674
rlabel metal2 65 -414 65 -414 0 net=256
rlabel metal2 138 -414 138 -414 0 net=562
rlabel metal2 65 -416 65 -416 0 net=189
rlabel metal2 93 -416 93 -416 0 net=124
rlabel metal2 142 -416 142 -416 0 net=335
rlabel metal2 114 -418 114 -418 0 net=223
rlabel metal2 12 -429 12 -429 0 net=262
rlabel metal2 19 -431 19 -431 0 net=422
rlabel metal2 47 -431 47 -431 0 net=30
rlabel metal2 65 -431 65 -431 0 net=190
rlabel metal2 79 -431 79 -431 0 net=548
rlabel metal2 72 -433 72 -433 0 net=434
rlabel metal2 89 -435 89 -435 0 net=196
rlabel metal2 114 -435 114 -435 0 net=224
rlabel metal2 96 -437 96 -437 0 net=250
rlabel metal2 121 -437 121 -437 0 net=336
<< end >>
