magic
tech scmos
timestamp 1555017055 
<< pdiffusion >>
rect 1 -10 7 -4
rect 8 -10 14 -4
rect 57 -10 63 -4
rect 71 -10 77 -4
rect 78 -10 84 -4
rect 99 -10 105 -4
rect 106 -10 112 -4
rect 113 -10 116 -4
rect 120 -10 126 -4
rect 127 -10 130 -4
rect 134 -10 140 -4
rect 141 -10 147 -4
rect 1 -29 7 -23
rect 8 -29 11 -23
rect 15 -29 21 -23
rect 22 -29 28 -23
rect 29 -29 32 -23
rect 36 -29 42 -23
rect 43 -29 46 -23
rect 50 -29 56 -23
rect 57 -29 63 -23
rect 64 -29 67 -23
rect 71 -29 74 -23
rect 78 -29 81 -23
rect 85 -29 91 -23
rect 92 -29 95 -23
rect 99 -29 105 -23
rect 106 -29 112 -23
rect 113 -29 116 -23
rect 120 -29 123 -23
rect 127 -29 130 -23
rect 134 -29 137 -23
rect 141 -29 144 -23
rect 148 -29 151 -23
rect 155 -29 158 -23
rect 162 -29 165 -23
rect 169 -29 175 -23
rect 8 -56 14 -50
rect 15 -56 18 -50
rect 22 -56 25 -50
rect 29 -56 35 -50
rect 36 -56 42 -50
rect 43 -56 49 -50
rect 50 -56 56 -50
rect 57 -56 60 -50
rect 64 -56 70 -50
rect 71 -56 77 -50
rect 78 -56 81 -50
rect 85 -56 91 -50
rect 92 -56 98 -50
rect 99 -56 102 -50
rect 106 -56 109 -50
rect 113 -56 116 -50
rect 120 -56 123 -50
rect 127 -56 130 -50
rect 134 -56 137 -50
rect 141 -56 144 -50
rect 148 -56 151 -50
rect 155 -56 158 -50
rect 162 -56 165 -50
rect 169 -56 172 -50
rect 176 -56 179 -50
rect 183 -56 189 -50
rect 1 -85 4 -79
rect 8 -85 14 -79
rect 15 -85 18 -79
rect 22 -85 28 -79
rect 29 -85 35 -79
rect 36 -85 39 -79
rect 43 -85 49 -79
rect 50 -85 56 -79
rect 57 -85 60 -79
rect 64 -85 67 -79
rect 71 -85 74 -79
rect 78 -85 84 -79
rect 85 -85 91 -79
rect 92 -85 95 -79
rect 99 -85 102 -79
rect 106 -85 109 -79
rect 113 -85 119 -79
rect 120 -85 126 -79
rect 127 -85 133 -79
rect 134 -85 137 -79
rect 141 -85 144 -79
rect 148 -85 151 -79
rect 155 -85 158 -79
rect 162 -85 165 -79
rect 169 -85 172 -79
rect 176 -85 179 -79
rect 183 -85 186 -79
rect 190 -85 193 -79
rect 197 -85 200 -79
rect 1 -124 7 -118
rect 8 -124 14 -118
rect 15 -124 18 -118
rect 22 -124 25 -118
rect 29 -124 35 -118
rect 36 -124 39 -118
rect 43 -124 46 -118
rect 50 -124 53 -118
rect 57 -124 63 -118
rect 64 -124 70 -118
rect 71 -124 74 -118
rect 78 -124 81 -118
rect 85 -124 88 -118
rect 92 -124 98 -118
rect 99 -124 102 -118
rect 106 -124 109 -118
rect 113 -124 119 -118
rect 120 -124 126 -118
rect 127 -124 133 -118
rect 134 -124 137 -118
rect 141 -124 144 -118
rect 148 -124 151 -118
rect 155 -124 158 -118
rect 162 -124 165 -118
rect 169 -124 175 -118
rect 176 -124 179 -118
rect 183 -124 186 -118
rect 190 -124 193 -118
rect 197 -124 200 -118
rect 204 -124 207 -118
rect 211 -124 214 -118
rect 1 -157 4 -151
rect 8 -157 14 -151
rect 15 -157 18 -151
rect 22 -157 28 -151
rect 29 -157 35 -151
rect 36 -157 39 -151
rect 43 -157 49 -151
rect 50 -157 53 -151
rect 57 -157 60 -151
rect 64 -157 67 -151
rect 71 -157 74 -151
rect 78 -157 81 -151
rect 85 -157 88 -151
rect 92 -157 98 -151
rect 99 -157 102 -151
rect 106 -157 109 -151
rect 113 -157 119 -151
rect 120 -157 126 -151
rect 127 -157 130 -151
rect 134 -157 140 -151
rect 141 -157 147 -151
rect 148 -157 154 -151
rect 155 -157 158 -151
rect 162 -157 165 -151
rect 169 -157 172 -151
rect 176 -157 179 -151
rect 183 -157 186 -151
rect 190 -157 193 -151
rect 197 -157 200 -151
rect 204 -157 207 -151
rect 211 -157 214 -151
rect 218 -157 221 -151
rect 225 -157 228 -151
rect 232 -157 235 -151
rect 239 -157 242 -151
rect 246 -157 249 -151
rect 1 -200 7 -194
rect 8 -200 14 -194
rect 15 -200 18 -194
rect 22 -200 25 -194
rect 29 -200 32 -194
rect 36 -200 39 -194
rect 43 -200 46 -194
rect 50 -200 56 -194
rect 57 -200 63 -194
rect 64 -200 70 -194
rect 71 -200 77 -194
rect 78 -200 81 -194
rect 85 -200 91 -194
rect 92 -200 95 -194
rect 99 -200 102 -194
rect 106 -200 112 -194
rect 113 -200 119 -194
rect 120 -200 123 -194
rect 127 -200 130 -194
rect 134 -200 137 -194
rect 141 -200 144 -194
rect 148 -200 151 -194
rect 155 -200 161 -194
rect 162 -200 165 -194
rect 169 -200 172 -194
rect 176 -200 179 -194
rect 183 -200 186 -194
rect 190 -200 193 -194
rect 197 -200 200 -194
rect 204 -200 207 -194
rect 211 -200 214 -194
rect 218 -200 221 -194
rect 225 -200 228 -194
rect 232 -200 235 -194
rect 239 -200 242 -194
rect 246 -200 249 -194
rect 253 -200 256 -194
rect 260 -200 263 -194
rect 267 -200 270 -194
rect 274 -200 277 -194
rect 281 -200 284 -194
rect 8 -241 11 -235
rect 15 -241 18 -235
rect 22 -241 25 -235
rect 29 -241 32 -235
rect 36 -241 42 -235
rect 43 -241 49 -235
rect 50 -241 56 -235
rect 57 -241 63 -235
rect 64 -241 70 -235
rect 71 -241 74 -235
rect 78 -241 81 -235
rect 85 -241 88 -235
rect 92 -241 98 -235
rect 99 -241 102 -235
rect 106 -241 109 -235
rect 113 -241 116 -235
rect 120 -241 123 -235
rect 127 -241 133 -235
rect 134 -241 137 -235
rect 141 -241 144 -235
rect 148 -241 151 -235
rect 155 -241 158 -235
rect 162 -241 165 -235
rect 169 -241 172 -235
rect 176 -241 182 -235
rect 183 -241 186 -235
rect 190 -241 196 -235
rect 197 -241 200 -235
rect 204 -241 207 -235
rect 211 -241 214 -235
rect 218 -241 221 -235
rect 225 -241 228 -235
rect 232 -241 238 -235
rect 239 -241 242 -235
rect 246 -241 249 -235
rect 1 -266 7 -260
rect 43 -266 46 -260
rect 57 -266 60 -260
rect 64 -266 70 -260
rect 71 -266 77 -260
rect 78 -266 81 -260
rect 85 -266 88 -260
rect 92 -266 95 -260
rect 99 -266 102 -260
rect 106 -266 109 -260
rect 113 -266 116 -260
rect 120 -266 126 -260
rect 127 -266 130 -260
rect 134 -266 137 -260
rect 141 -266 147 -260
rect 148 -266 151 -260
rect 155 -266 161 -260
rect 162 -266 165 -260
rect 169 -266 175 -260
rect 176 -266 179 -260
rect 183 -266 186 -260
rect 190 -266 196 -260
rect 197 -266 200 -260
rect 204 -266 210 -260
rect 211 -266 217 -260
rect 218 -266 221 -260
rect 225 -266 228 -260
rect 232 -266 235 -260
rect 239 -266 242 -260
rect 1 -283 7 -277
rect 43 -283 49 -277
rect 64 -283 70 -277
rect 71 -283 74 -277
rect 78 -283 84 -277
rect 99 -283 105 -277
rect 120 -283 123 -277
rect 127 -283 133 -277
rect 134 -283 140 -277
rect 141 -283 144 -277
rect 148 -283 154 -277
rect 197 -283 203 -277
rect 204 -283 210 -277
<< polysilicon >>
rect 61 -11 62 -9
rect 72 -11 73 -9
rect 79 -11 80 -9
rect 103 -11 104 -9
rect 107 -5 108 -3
rect 110 -11 111 -9
rect 114 -5 115 -3
rect 114 -11 115 -9
rect 124 -5 125 -3
rect 128 -5 129 -3
rect 128 -11 129 -9
rect 138 -11 139 -9
rect 145 -11 146 -9
rect 9 -24 10 -22
rect 9 -30 10 -28
rect 19 -30 20 -28
rect 23 -30 24 -28
rect 26 -30 27 -28
rect 30 -24 31 -22
rect 30 -30 31 -28
rect 40 -24 41 -22
rect 44 -24 45 -22
rect 44 -30 45 -28
rect 54 -24 55 -22
rect 54 -30 55 -28
rect 61 -24 62 -22
rect 58 -30 59 -28
rect 61 -30 62 -28
rect 65 -24 66 -22
rect 65 -30 66 -28
rect 72 -24 73 -22
rect 72 -30 73 -28
rect 79 -24 80 -22
rect 79 -30 80 -28
rect 86 -30 87 -28
rect 89 -30 90 -28
rect 93 -24 94 -22
rect 93 -30 94 -28
rect 103 -24 104 -22
rect 110 -24 111 -22
rect 110 -30 111 -28
rect 114 -24 115 -22
rect 114 -30 115 -28
rect 121 -24 122 -22
rect 121 -30 122 -28
rect 128 -24 129 -22
rect 128 -30 129 -28
rect 135 -24 136 -22
rect 135 -30 136 -28
rect 142 -24 143 -22
rect 142 -30 143 -28
rect 149 -24 150 -22
rect 149 -30 150 -28
rect 156 -24 157 -22
rect 156 -30 157 -28
rect 163 -24 164 -22
rect 163 -30 164 -28
rect 170 -24 171 -22
rect 9 -57 10 -55
rect 16 -51 17 -49
rect 16 -57 17 -55
rect 23 -51 24 -49
rect 23 -57 24 -55
rect 30 -51 31 -49
rect 33 -57 34 -55
rect 37 -51 38 -49
rect 40 -51 41 -49
rect 47 -51 48 -49
rect 44 -57 45 -55
rect 54 -51 55 -49
rect 51 -57 52 -55
rect 54 -57 55 -55
rect 58 -51 59 -49
rect 58 -57 59 -55
rect 65 -51 66 -49
rect 68 -51 69 -49
rect 65 -57 66 -55
rect 72 -51 73 -49
rect 75 -57 76 -55
rect 79 -51 80 -49
rect 79 -57 80 -55
rect 86 -51 87 -49
rect 89 -57 90 -55
rect 93 -51 94 -49
rect 93 -57 94 -55
rect 100 -51 101 -49
rect 100 -57 101 -55
rect 107 -51 108 -49
rect 107 -57 108 -55
rect 114 -51 115 -49
rect 114 -57 115 -55
rect 121 -51 122 -49
rect 121 -57 122 -55
rect 128 -51 129 -49
rect 128 -57 129 -55
rect 135 -51 136 -49
rect 135 -57 136 -55
rect 142 -51 143 -49
rect 142 -57 143 -55
rect 149 -51 150 -49
rect 149 -57 150 -55
rect 156 -51 157 -49
rect 156 -57 157 -55
rect 163 -51 164 -49
rect 163 -57 164 -55
rect 170 -51 171 -49
rect 170 -57 171 -55
rect 177 -51 178 -49
rect 177 -57 178 -55
rect 184 -57 185 -55
rect 2 -80 3 -78
rect 2 -86 3 -84
rect 16 -80 17 -78
rect 16 -86 17 -84
rect 26 -80 27 -78
rect 26 -86 27 -84
rect 33 -80 34 -78
rect 30 -86 31 -84
rect 37 -80 38 -78
rect 37 -86 38 -84
rect 44 -80 45 -78
rect 47 -80 48 -78
rect 51 -80 52 -78
rect 54 -86 55 -84
rect 58 -80 59 -78
rect 58 -86 59 -84
rect 65 -80 66 -78
rect 65 -86 66 -84
rect 72 -80 73 -78
rect 72 -86 73 -84
rect 79 -80 80 -78
rect 82 -80 83 -78
rect 79 -86 80 -84
rect 89 -86 90 -84
rect 93 -80 94 -78
rect 93 -86 94 -84
rect 100 -80 101 -78
rect 100 -86 101 -84
rect 107 -80 108 -78
rect 107 -86 108 -84
rect 114 -80 115 -78
rect 114 -86 115 -84
rect 117 -86 118 -84
rect 124 -80 125 -78
rect 124 -86 125 -84
rect 131 -86 132 -84
rect 135 -80 136 -78
rect 135 -86 136 -84
rect 142 -80 143 -78
rect 142 -86 143 -84
rect 149 -80 150 -78
rect 149 -86 150 -84
rect 156 -80 157 -78
rect 156 -86 157 -84
rect 163 -80 164 -78
rect 163 -86 164 -84
rect 170 -80 171 -78
rect 170 -86 171 -84
rect 177 -80 178 -78
rect 177 -86 178 -84
rect 184 -80 185 -78
rect 184 -86 185 -84
rect 191 -80 192 -78
rect 191 -86 192 -84
rect 198 -80 199 -78
rect 198 -86 199 -84
rect 2 -119 3 -117
rect 2 -125 3 -123
rect 9 -125 10 -123
rect 16 -119 17 -117
rect 16 -125 17 -123
rect 23 -119 24 -117
rect 23 -125 24 -123
rect 33 -119 34 -117
rect 30 -125 31 -123
rect 33 -125 34 -123
rect 37 -119 38 -117
rect 37 -125 38 -123
rect 44 -119 45 -117
rect 44 -125 45 -123
rect 51 -119 52 -117
rect 51 -125 52 -123
rect 58 -119 59 -117
rect 58 -125 59 -123
rect 61 -125 62 -123
rect 68 -119 69 -117
rect 68 -125 69 -123
rect 72 -119 73 -117
rect 72 -125 73 -123
rect 79 -119 80 -117
rect 79 -125 80 -123
rect 86 -119 87 -117
rect 86 -125 87 -123
rect 93 -119 94 -117
rect 96 -119 97 -117
rect 93 -125 94 -123
rect 96 -125 97 -123
rect 100 -119 101 -117
rect 100 -125 101 -123
rect 107 -119 108 -117
rect 107 -125 108 -123
rect 117 -119 118 -117
rect 114 -125 115 -123
rect 117 -125 118 -123
rect 121 -119 122 -117
rect 124 -119 125 -117
rect 121 -125 122 -123
rect 124 -125 125 -123
rect 128 -119 129 -117
rect 131 -119 132 -117
rect 135 -119 136 -117
rect 135 -125 136 -123
rect 142 -119 143 -117
rect 142 -125 143 -123
rect 149 -119 150 -117
rect 149 -125 150 -123
rect 156 -119 157 -117
rect 156 -125 157 -123
rect 163 -119 164 -117
rect 163 -125 164 -123
rect 170 -125 171 -123
rect 173 -125 174 -123
rect 177 -119 178 -117
rect 177 -125 178 -123
rect 184 -119 185 -117
rect 184 -125 185 -123
rect 191 -119 192 -117
rect 191 -125 192 -123
rect 198 -119 199 -117
rect 198 -125 199 -123
rect 205 -119 206 -117
rect 205 -125 206 -123
rect 212 -119 213 -117
rect 212 -125 213 -123
rect 2 -152 3 -150
rect 2 -158 3 -156
rect 12 -152 13 -150
rect 9 -158 10 -156
rect 16 -152 17 -150
rect 16 -158 17 -156
rect 23 -158 24 -156
rect 26 -158 27 -156
rect 33 -152 34 -150
rect 30 -158 31 -156
rect 33 -158 34 -156
rect 37 -152 38 -150
rect 37 -158 38 -156
rect 44 -152 45 -150
rect 47 -152 48 -150
rect 44 -158 45 -156
rect 51 -152 52 -150
rect 51 -158 52 -156
rect 58 -152 59 -150
rect 58 -158 59 -156
rect 65 -152 66 -150
rect 65 -158 66 -156
rect 72 -152 73 -150
rect 72 -158 73 -156
rect 79 -152 80 -150
rect 79 -158 80 -156
rect 86 -152 87 -150
rect 86 -158 87 -156
rect 93 -152 94 -150
rect 93 -158 94 -156
rect 96 -158 97 -156
rect 100 -152 101 -150
rect 100 -158 101 -156
rect 107 -152 108 -150
rect 107 -158 108 -156
rect 114 -152 115 -150
rect 117 -152 118 -150
rect 114 -158 115 -156
rect 117 -158 118 -156
rect 121 -152 122 -150
rect 124 -158 125 -156
rect 128 -152 129 -150
rect 128 -158 129 -156
rect 135 -152 136 -150
rect 145 -152 146 -150
rect 142 -158 143 -156
rect 149 -152 150 -150
rect 152 -152 153 -150
rect 152 -158 153 -156
rect 156 -152 157 -150
rect 156 -158 157 -156
rect 163 -152 164 -150
rect 163 -158 164 -156
rect 170 -152 171 -150
rect 170 -158 171 -156
rect 177 -152 178 -150
rect 177 -158 178 -156
rect 184 -152 185 -150
rect 184 -158 185 -156
rect 191 -152 192 -150
rect 191 -158 192 -156
rect 198 -152 199 -150
rect 198 -158 199 -156
rect 205 -152 206 -150
rect 205 -158 206 -156
rect 212 -152 213 -150
rect 212 -158 213 -156
rect 219 -152 220 -150
rect 219 -158 220 -156
rect 226 -152 227 -150
rect 226 -158 227 -156
rect 233 -152 234 -150
rect 233 -158 234 -156
rect 240 -152 241 -150
rect 240 -158 241 -156
rect 247 -152 248 -150
rect 247 -158 248 -156
rect 2 -195 3 -193
rect 5 -195 6 -193
rect 9 -195 10 -193
rect 9 -201 10 -199
rect 16 -195 17 -193
rect 16 -201 17 -199
rect 23 -195 24 -193
rect 23 -201 24 -199
rect 30 -195 31 -193
rect 30 -201 31 -199
rect 37 -195 38 -193
rect 37 -201 38 -199
rect 44 -195 45 -193
rect 44 -201 45 -199
rect 51 -195 52 -193
rect 54 -195 55 -193
rect 54 -201 55 -199
rect 61 -195 62 -193
rect 58 -201 59 -199
rect 61 -201 62 -199
rect 65 -195 66 -193
rect 68 -201 69 -199
rect 72 -195 73 -193
rect 75 -195 76 -193
rect 75 -201 76 -199
rect 79 -195 80 -193
rect 79 -201 80 -199
rect 86 -195 87 -193
rect 89 -195 90 -193
rect 86 -201 87 -199
rect 89 -201 90 -199
rect 93 -195 94 -193
rect 93 -201 94 -199
rect 100 -195 101 -193
rect 100 -201 101 -199
rect 107 -195 108 -193
rect 110 -195 111 -193
rect 107 -201 108 -199
rect 110 -201 111 -199
rect 114 -195 115 -193
rect 117 -195 118 -193
rect 114 -201 115 -199
rect 117 -201 118 -199
rect 121 -195 122 -193
rect 121 -201 122 -199
rect 128 -195 129 -193
rect 128 -201 129 -199
rect 135 -195 136 -193
rect 135 -201 136 -199
rect 142 -195 143 -193
rect 142 -201 143 -199
rect 149 -195 150 -193
rect 149 -201 150 -199
rect 159 -195 160 -193
rect 156 -201 157 -199
rect 159 -201 160 -199
rect 163 -195 164 -193
rect 163 -201 164 -199
rect 170 -195 171 -193
rect 170 -201 171 -199
rect 177 -195 178 -193
rect 177 -201 178 -199
rect 184 -195 185 -193
rect 184 -201 185 -199
rect 191 -195 192 -193
rect 191 -201 192 -199
rect 198 -195 199 -193
rect 198 -201 199 -199
rect 205 -195 206 -193
rect 205 -201 206 -199
rect 212 -195 213 -193
rect 212 -201 213 -199
rect 219 -195 220 -193
rect 219 -201 220 -199
rect 226 -195 227 -193
rect 226 -201 227 -199
rect 233 -195 234 -193
rect 233 -201 234 -199
rect 240 -195 241 -193
rect 240 -201 241 -199
rect 247 -195 248 -193
rect 247 -201 248 -199
rect 254 -195 255 -193
rect 254 -201 255 -199
rect 261 -195 262 -193
rect 261 -201 262 -199
rect 268 -195 269 -193
rect 268 -201 269 -199
rect 275 -195 276 -193
rect 275 -201 276 -199
rect 282 -195 283 -193
rect 282 -201 283 -199
rect 9 -236 10 -234
rect 9 -242 10 -240
rect 16 -236 17 -234
rect 16 -242 17 -240
rect 23 -236 24 -234
rect 23 -242 24 -240
rect 30 -236 31 -234
rect 30 -242 31 -240
rect 37 -236 38 -234
rect 40 -236 41 -234
rect 47 -236 48 -234
rect 44 -242 45 -240
rect 47 -242 48 -240
rect 51 -236 52 -234
rect 54 -242 55 -240
rect 58 -236 59 -234
rect 58 -242 59 -240
rect 61 -242 62 -240
rect 65 -242 66 -240
rect 68 -242 69 -240
rect 72 -236 73 -234
rect 72 -242 73 -240
rect 79 -236 80 -234
rect 79 -242 80 -240
rect 86 -236 87 -234
rect 86 -242 87 -240
rect 93 -236 94 -234
rect 93 -242 94 -240
rect 96 -242 97 -240
rect 100 -236 101 -234
rect 100 -242 101 -240
rect 107 -236 108 -234
rect 107 -242 108 -240
rect 114 -236 115 -234
rect 114 -242 115 -240
rect 121 -236 122 -234
rect 121 -242 122 -240
rect 128 -236 129 -234
rect 131 -236 132 -234
rect 128 -242 129 -240
rect 131 -242 132 -240
rect 135 -236 136 -234
rect 135 -242 136 -240
rect 142 -236 143 -234
rect 142 -242 143 -240
rect 149 -236 150 -234
rect 149 -242 150 -240
rect 156 -236 157 -234
rect 156 -242 157 -240
rect 163 -236 164 -234
rect 163 -242 164 -240
rect 170 -236 171 -234
rect 170 -242 171 -240
rect 177 -236 178 -234
rect 180 -236 181 -234
rect 177 -242 178 -240
rect 184 -236 185 -234
rect 184 -242 185 -240
rect 194 -236 195 -234
rect 194 -242 195 -240
rect 198 -236 199 -234
rect 198 -242 199 -240
rect 205 -236 206 -234
rect 205 -242 206 -240
rect 212 -236 213 -234
rect 212 -242 213 -240
rect 219 -236 220 -234
rect 219 -242 220 -240
rect 226 -236 227 -234
rect 226 -242 227 -240
rect 233 -236 234 -234
rect 240 -236 241 -234
rect 240 -242 241 -240
rect 247 -236 248 -234
rect 247 -242 248 -240
rect 44 -261 45 -259
rect 44 -267 45 -265
rect 58 -261 59 -259
rect 58 -267 59 -265
rect 65 -261 66 -259
rect 65 -267 66 -265
rect 72 -267 73 -265
rect 75 -267 76 -265
rect 79 -261 80 -259
rect 79 -267 80 -265
rect 86 -261 87 -259
rect 86 -267 87 -265
rect 93 -261 94 -259
rect 93 -267 94 -265
rect 100 -261 101 -259
rect 100 -267 101 -265
rect 107 -261 108 -259
rect 107 -267 108 -265
rect 114 -261 115 -259
rect 114 -267 115 -265
rect 121 -267 122 -265
rect 124 -267 125 -265
rect 128 -261 129 -259
rect 128 -267 129 -265
rect 135 -261 136 -259
rect 135 -267 136 -265
rect 142 -267 143 -265
rect 145 -267 146 -265
rect 149 -261 150 -259
rect 149 -267 150 -265
rect 159 -261 160 -259
rect 156 -267 157 -265
rect 159 -267 160 -265
rect 163 -261 164 -259
rect 163 -267 164 -265
rect 170 -261 171 -259
rect 173 -267 174 -265
rect 177 -261 178 -259
rect 177 -267 178 -265
rect 184 -261 185 -259
rect 184 -267 185 -265
rect 191 -261 192 -259
rect 191 -267 192 -265
rect 194 -267 195 -265
rect 198 -261 199 -259
rect 198 -267 199 -265
rect 208 -261 209 -259
rect 205 -267 206 -265
rect 212 -261 213 -259
rect 215 -261 216 -259
rect 219 -261 220 -259
rect 219 -267 220 -265
rect 226 -261 227 -259
rect 226 -267 227 -265
rect 233 -261 234 -259
rect 233 -267 234 -265
rect 240 -261 241 -259
rect 240 -267 241 -265
rect 47 -278 48 -276
rect 65 -284 66 -282
rect 72 -278 73 -276
rect 72 -284 73 -282
rect 79 -278 80 -276
rect 100 -278 101 -276
rect 103 -278 104 -276
rect 121 -278 122 -276
rect 121 -284 122 -282
rect 128 -278 129 -276
rect 131 -284 132 -282
rect 138 -278 139 -276
rect 142 -278 143 -276
rect 142 -284 143 -282
rect 149 -284 150 -282
rect 201 -278 202 -276
rect 205 -278 206 -276
rect 208 -278 209 -276
<< metal1 >>
rect 107 0 129 1
rect 114 -2 125 -1
rect 30 -13 41 -12
rect 44 -13 62 -12
rect 65 -13 73 -12
rect 103 -13 136 -12
rect 138 -13 150 -12
rect 156 -13 171 -12
rect 9 -15 62 -14
rect 72 -15 80 -14
rect 93 -15 104 -14
rect 128 -15 143 -14
rect 145 -15 164 -14
rect 54 -17 80 -16
rect 114 -17 129 -16
rect 110 -19 115 -18
rect 110 -21 122 -20
rect 9 -32 55 -31
rect 58 -32 101 -31
rect 110 -32 150 -31
rect 16 -34 66 -33
rect 68 -34 80 -33
rect 121 -34 150 -33
rect 23 -36 27 -35
rect 30 -36 41 -35
rect 44 -36 80 -35
rect 114 -36 122 -35
rect 128 -36 171 -35
rect 19 -38 24 -37
rect 30 -38 48 -37
rect 54 -38 66 -37
rect 72 -38 87 -37
rect 89 -38 115 -37
rect 37 -40 59 -39
rect 61 -40 136 -39
rect 72 -42 129 -41
rect 86 -44 108 -43
rect 93 -46 136 -45
rect 93 -48 178 -47
rect 2 -59 48 -58
rect 51 -59 101 -58
rect 142 -59 199 -58
rect 16 -61 76 -60
rect 82 -61 136 -60
rect 156 -61 192 -60
rect 16 -63 125 -62
rect 135 -63 178 -62
rect 26 -65 101 -64
rect 121 -65 157 -64
rect 37 -67 45 -66
rect 51 -67 143 -66
rect 149 -67 178 -66
rect 9 -69 45 -68
rect 54 -69 73 -68
rect 93 -69 115 -68
rect 23 -71 94 -70
rect 107 -71 150 -70
rect 65 -73 90 -72
rect 114 -73 171 -72
rect 58 -75 66 -74
rect 79 -75 108 -74
rect 128 -75 171 -74
rect 58 -77 80 -76
rect 23 -88 31 -87
rect 37 -88 45 -87
rect 51 -88 59 -87
rect 68 -88 108 -87
rect 114 -88 178 -87
rect 26 -90 66 -89
rect 79 -90 150 -89
rect 163 -90 213 -89
rect 16 -92 80 -91
rect 86 -92 118 -91
rect 124 -92 192 -91
rect 16 -94 94 -93
rect 96 -94 108 -93
rect 128 -94 199 -93
rect 33 -96 150 -95
rect 170 -96 178 -95
rect 184 -96 192 -95
rect 37 -98 122 -97
rect 142 -98 164 -97
rect 58 -100 132 -99
rect 89 -102 136 -101
rect 54 -104 136 -103
rect 93 -106 157 -105
rect 100 -108 157 -107
rect 72 -110 101 -109
rect 117 -110 199 -109
rect 2 -112 73 -111
rect 124 -112 143 -111
rect 2 -114 206 -113
rect 131 -116 185 -115
rect 2 -127 17 -126
rect 23 -127 31 -126
rect 33 -127 125 -126
rect 149 -127 248 -126
rect 2 -129 59 -128
rect 61 -129 101 -128
rect 117 -129 129 -128
rect 149 -129 234 -128
rect 9 -131 13 -130
rect 16 -131 48 -130
rect 51 -131 66 -130
rect 72 -131 118 -130
rect 121 -131 213 -130
rect 33 -133 52 -132
rect 58 -133 94 -132
rect 96 -133 199 -132
rect 37 -135 73 -134
rect 79 -135 115 -134
rect 121 -135 220 -134
rect 37 -137 45 -136
rect 68 -137 80 -136
rect 86 -137 101 -136
rect 114 -137 227 -136
rect 86 -139 136 -138
rect 152 -139 171 -138
rect 173 -139 213 -138
rect 93 -141 146 -140
rect 163 -141 171 -140
rect 191 -141 199 -140
rect 135 -143 241 -142
rect 142 -145 164 -144
rect 184 -145 192 -144
rect 177 -147 185 -146
rect 44 -149 178 -148
rect 5 -160 10 -159
rect 23 -160 52 -159
rect 61 -160 220 -159
rect 233 -160 283 -159
rect 9 -162 17 -161
rect 23 -162 90 -161
rect 117 -162 185 -161
rect 191 -162 234 -161
rect 16 -164 59 -163
rect 75 -164 122 -163
rect 124 -164 150 -163
rect 177 -164 276 -163
rect 26 -166 241 -165
rect 30 -168 269 -167
rect 30 -170 66 -169
rect 79 -170 178 -169
rect 198 -170 241 -169
rect 33 -172 87 -171
rect 117 -172 136 -171
rect 142 -172 164 -171
rect 198 -172 248 -171
rect 2 -174 164 -173
rect 205 -174 255 -173
rect 2 -176 227 -175
rect 44 -178 192 -177
rect 212 -178 262 -177
rect 44 -180 111 -179
rect 114 -180 143 -179
rect 152 -180 248 -179
rect 51 -182 185 -181
rect 54 -184 80 -183
rect 96 -184 227 -183
rect 65 -186 94 -185
rect 128 -186 220 -185
rect 72 -188 87 -187
rect 100 -188 129 -187
rect 156 -188 206 -187
rect 72 -190 94 -189
rect 100 -190 108 -189
rect 170 -190 213 -189
rect 107 -192 115 -191
rect 159 -192 171 -191
rect 9 -203 164 -202
rect 180 -203 192 -202
rect 9 -205 69 -204
rect 72 -205 122 -204
rect 135 -205 164 -204
rect 30 -207 34 -206
rect 47 -207 269 -206
rect 30 -209 38 -208
rect 51 -209 132 -208
rect 156 -209 255 -208
rect 33 -211 38 -210
rect 54 -211 248 -210
rect 58 -213 90 -212
rect 107 -213 136 -212
rect 156 -213 171 -212
rect 198 -213 248 -212
rect 44 -215 59 -214
rect 75 -215 118 -214
rect 121 -215 143 -214
rect 159 -215 283 -214
rect 86 -217 101 -216
rect 107 -217 150 -216
rect 170 -217 213 -216
rect 23 -219 101 -218
rect 110 -219 220 -218
rect 16 -221 24 -220
rect 40 -221 87 -220
rect 114 -221 206 -220
rect 212 -221 234 -220
rect 16 -223 62 -222
rect 79 -223 115 -222
rect 142 -223 178 -222
rect 198 -223 227 -222
rect 79 -225 94 -224
rect 149 -225 185 -224
rect 205 -225 234 -224
rect 93 -227 129 -226
rect 177 -227 220 -226
rect 226 -227 262 -226
rect 128 -229 276 -228
rect 184 -231 241 -230
rect 194 -233 241 -232
rect 9 -244 94 -243
rect 131 -244 150 -243
rect 159 -244 206 -243
rect 233 -244 241 -243
rect 16 -246 62 -245
rect 68 -246 80 -245
rect 86 -246 94 -245
rect 135 -246 192 -245
rect 194 -246 227 -245
rect 23 -248 66 -247
rect 79 -248 143 -247
rect 149 -248 164 -247
rect 177 -248 248 -247
rect 30 -250 55 -249
rect 65 -250 97 -249
rect 128 -250 136 -249
rect 163 -250 185 -249
rect 212 -250 241 -249
rect 44 -252 73 -251
rect 86 -252 115 -251
rect 128 -252 171 -251
rect 177 -252 199 -251
rect 208 -252 213 -251
rect 44 -254 48 -253
rect 114 -254 122 -253
rect 156 -254 185 -253
rect 198 -254 220 -253
rect 170 -256 227 -255
rect 215 -258 220 -257
rect 44 -269 48 -268
rect 58 -269 66 -268
rect 75 -269 80 -268
rect 86 -269 125 -268
rect 135 -269 139 -268
rect 142 -269 150 -268
rect 163 -269 174 -268
rect 177 -269 195 -268
rect 201 -269 227 -268
rect 79 -271 94 -270
rect 100 -271 104 -270
rect 121 -271 185 -270
rect 191 -271 199 -270
rect 205 -271 234 -270
rect 100 -273 108 -272
rect 114 -273 122 -272
rect 128 -273 143 -272
rect 145 -273 157 -272
rect 205 -273 220 -272
rect 128 -275 160 -274
rect 208 -275 241 -274
rect 65 -286 73 -285
rect 121 -286 132 -285
rect 142 -286 150 -285
<< m2contact >>
rect 107 0 108 1
rect 128 0 129 1
rect 114 -2 115 -1
rect 124 -2 125 -1
rect 30 -13 31 -12
rect 40 -13 41 -12
rect 44 -13 45 -12
rect 61 -13 62 -12
rect 65 -13 66 -12
rect 72 -13 73 -12
rect 103 -13 104 -12
rect 135 -13 136 -12
rect 138 -13 139 -12
rect 149 -13 150 -12
rect 156 -13 157 -12
rect 170 -13 171 -12
rect 9 -15 10 -14
rect 61 -15 62 -14
rect 72 -15 73 -14
rect 79 -15 80 -14
rect 93 -15 94 -14
rect 103 -15 104 -14
rect 128 -15 129 -14
rect 142 -15 143 -14
rect 145 -15 146 -14
rect 163 -15 164 -14
rect 54 -17 55 -16
rect 79 -17 80 -16
rect 114 -17 115 -16
rect 128 -17 129 -16
rect 110 -19 111 -18
rect 114 -19 115 -18
rect 110 -21 111 -20
rect 121 -21 122 -20
rect 9 -32 10 -31
rect 54 -32 55 -31
rect 58 -32 59 -31
rect 100 -32 101 -31
rect 110 -32 111 -31
rect 149 -32 150 -31
rect 16 -34 17 -33
rect 65 -34 66 -33
rect 68 -34 69 -33
rect 79 -34 80 -33
rect 121 -34 122 -33
rect 149 -34 150 -33
rect 23 -36 24 -35
rect 26 -36 27 -35
rect 30 -36 31 -35
rect 40 -36 41 -35
rect 44 -36 45 -35
rect 79 -36 80 -35
rect 114 -36 115 -35
rect 121 -36 122 -35
rect 128 -36 129 -35
rect 170 -36 171 -35
rect 19 -38 20 -37
rect 23 -38 24 -37
rect 30 -38 31 -37
rect 47 -38 48 -37
rect 54 -38 55 -37
rect 65 -38 66 -37
rect 72 -38 73 -37
rect 86 -38 87 -37
rect 89 -38 90 -37
rect 114 -38 115 -37
rect 37 -40 38 -39
rect 58 -40 59 -39
rect 61 -40 62 -39
rect 135 -40 136 -39
rect 72 -42 73 -41
rect 128 -42 129 -41
rect 86 -44 87 -43
rect 107 -44 108 -43
rect 93 -46 94 -45
rect 135 -46 136 -45
rect 93 -48 94 -47
rect 177 -48 178 -47
rect 2 -59 3 -58
rect 47 -59 48 -58
rect 51 -59 52 -58
rect 100 -59 101 -58
rect 142 -59 143 -58
rect 198 -59 199 -58
rect 16 -61 17 -60
rect 75 -61 76 -60
rect 82 -61 83 -60
rect 135 -61 136 -60
rect 156 -61 157 -60
rect 191 -61 192 -60
rect 16 -63 17 -62
rect 124 -63 125 -62
rect 135 -63 136 -62
rect 177 -63 178 -62
rect 26 -65 27 -64
rect 100 -65 101 -64
rect 121 -65 122 -64
rect 156 -65 157 -64
rect 37 -67 38 -66
rect 44 -67 45 -66
rect 51 -67 52 -66
rect 142 -67 143 -66
rect 149 -67 150 -66
rect 177 -67 178 -66
rect 9 -69 10 -68
rect 44 -69 45 -68
rect 54 -69 55 -68
rect 72 -69 73 -68
rect 93 -69 94 -68
rect 114 -69 115 -68
rect 23 -71 24 -70
rect 93 -71 94 -70
rect 107 -71 108 -70
rect 149 -71 150 -70
rect 65 -73 66 -72
rect 89 -73 90 -72
rect 114 -73 115 -72
rect 170 -73 171 -72
rect 58 -75 59 -74
rect 65 -75 66 -74
rect 79 -75 80 -74
rect 107 -75 108 -74
rect 128 -75 129 -74
rect 170 -75 171 -74
rect 58 -77 59 -76
rect 79 -77 80 -76
rect 23 -88 24 -87
rect 30 -88 31 -87
rect 37 -88 38 -87
rect 44 -88 45 -87
rect 51 -88 52 -87
rect 58 -88 59 -87
rect 68 -88 69 -87
rect 107 -88 108 -87
rect 114 -88 115 -87
rect 177 -88 178 -87
rect 26 -90 27 -89
rect 65 -90 66 -89
rect 79 -90 80 -89
rect 149 -90 150 -89
rect 163 -90 164 -89
rect 212 -90 213 -89
rect 16 -92 17 -91
rect 79 -92 80 -91
rect 86 -92 87 -91
rect 117 -92 118 -91
rect 124 -92 125 -91
rect 191 -92 192 -91
rect 16 -94 17 -93
rect 93 -94 94 -93
rect 96 -94 97 -93
rect 107 -94 108 -93
rect 128 -94 129 -93
rect 198 -94 199 -93
rect 33 -96 34 -95
rect 149 -96 150 -95
rect 170 -96 171 -95
rect 177 -96 178 -95
rect 184 -96 185 -95
rect 191 -96 192 -95
rect 37 -98 38 -97
rect 121 -98 122 -97
rect 142 -98 143 -97
rect 163 -98 164 -97
rect 58 -100 59 -99
rect 131 -100 132 -99
rect 89 -102 90 -101
rect 135 -102 136 -101
rect 54 -104 55 -103
rect 135 -104 136 -103
rect 93 -106 94 -105
rect 156 -106 157 -105
rect 100 -108 101 -107
rect 156 -108 157 -107
rect 72 -110 73 -109
rect 100 -110 101 -109
rect 117 -110 118 -109
rect 198 -110 199 -109
rect 2 -112 3 -111
rect 72 -112 73 -111
rect 124 -112 125 -111
rect 142 -112 143 -111
rect 2 -114 3 -113
rect 205 -114 206 -113
rect 131 -116 132 -115
rect 184 -116 185 -115
rect 2 -127 3 -126
rect 16 -127 17 -126
rect 23 -127 24 -126
rect 30 -127 31 -126
rect 33 -127 34 -126
rect 124 -127 125 -126
rect 149 -127 150 -126
rect 247 -127 248 -126
rect 2 -129 3 -128
rect 58 -129 59 -128
rect 61 -129 62 -128
rect 100 -129 101 -128
rect 117 -129 118 -128
rect 128 -129 129 -128
rect 149 -129 150 -128
rect 233 -129 234 -128
rect 9 -131 10 -130
rect 12 -131 13 -130
rect 16 -131 17 -130
rect 47 -131 48 -130
rect 51 -131 52 -130
rect 65 -131 66 -130
rect 72 -131 73 -130
rect 117 -131 118 -130
rect 121 -131 122 -130
rect 212 -131 213 -130
rect 33 -133 34 -132
rect 51 -133 52 -132
rect 58 -133 59 -132
rect 93 -133 94 -132
rect 96 -133 97 -132
rect 198 -133 199 -132
rect 37 -135 38 -134
rect 72 -135 73 -134
rect 79 -135 80 -134
rect 114 -135 115 -134
rect 121 -135 122 -134
rect 219 -135 220 -134
rect 37 -137 38 -136
rect 44 -137 45 -136
rect 68 -137 69 -136
rect 79 -137 80 -136
rect 86 -137 87 -136
rect 100 -137 101 -136
rect 114 -137 115 -136
rect 226 -137 227 -136
rect 86 -139 87 -138
rect 135 -139 136 -138
rect 152 -139 153 -138
rect 170 -139 171 -138
rect 173 -139 174 -138
rect 212 -139 213 -138
rect 93 -141 94 -140
rect 145 -141 146 -140
rect 163 -141 164 -140
rect 170 -141 171 -140
rect 191 -141 192 -140
rect 198 -141 199 -140
rect 135 -143 136 -142
rect 240 -143 241 -142
rect 142 -145 143 -144
rect 163 -145 164 -144
rect 184 -145 185 -144
rect 191 -145 192 -144
rect 177 -147 178 -146
rect 184 -147 185 -146
rect 44 -149 45 -148
rect 177 -149 178 -148
rect 5 -160 6 -159
rect 9 -160 10 -159
rect 23 -160 24 -159
rect 51 -160 52 -159
rect 61 -160 62 -159
rect 219 -160 220 -159
rect 233 -160 234 -159
rect 282 -160 283 -159
rect 9 -162 10 -161
rect 16 -162 17 -161
rect 23 -162 24 -161
rect 89 -162 90 -161
rect 117 -162 118 -161
rect 184 -162 185 -161
rect 191 -162 192 -161
rect 233 -162 234 -161
rect 16 -164 17 -163
rect 58 -164 59 -163
rect 75 -164 76 -163
rect 121 -164 122 -163
rect 124 -164 125 -163
rect 149 -164 150 -163
rect 177 -164 178 -163
rect 275 -164 276 -163
rect 26 -166 27 -165
rect 240 -166 241 -165
rect 30 -168 31 -167
rect 268 -168 269 -167
rect 30 -170 31 -169
rect 65 -170 66 -169
rect 79 -170 80 -169
rect 177 -170 178 -169
rect 198 -170 199 -169
rect 240 -170 241 -169
rect 33 -172 34 -171
rect 86 -172 87 -171
rect 117 -172 118 -171
rect 135 -172 136 -171
rect 142 -172 143 -171
rect 163 -172 164 -171
rect 198 -172 199 -171
rect 247 -172 248 -171
rect 2 -174 3 -173
rect 163 -174 164 -173
rect 205 -174 206 -173
rect 254 -174 255 -173
rect 2 -176 3 -175
rect 226 -176 227 -175
rect 44 -178 45 -177
rect 191 -178 192 -177
rect 212 -178 213 -177
rect 261 -178 262 -177
rect 44 -180 45 -179
rect 110 -180 111 -179
rect 114 -180 115 -179
rect 142 -180 143 -179
rect 152 -180 153 -179
rect 247 -180 248 -179
rect 51 -182 52 -181
rect 184 -182 185 -181
rect 54 -184 55 -183
rect 79 -184 80 -183
rect 96 -184 97 -183
rect 226 -184 227 -183
rect 65 -186 66 -185
rect 93 -186 94 -185
rect 128 -186 129 -185
rect 219 -186 220 -185
rect 72 -188 73 -187
rect 86 -188 87 -187
rect 100 -188 101 -187
rect 128 -188 129 -187
rect 156 -188 157 -187
rect 205 -188 206 -187
rect 72 -190 73 -189
rect 93 -190 94 -189
rect 100 -190 101 -189
rect 107 -190 108 -189
rect 170 -190 171 -189
rect 212 -190 213 -189
rect 107 -192 108 -191
rect 114 -192 115 -191
rect 159 -192 160 -191
rect 170 -192 171 -191
rect 9 -203 10 -202
rect 163 -203 164 -202
rect 180 -203 181 -202
rect 191 -203 192 -202
rect 9 -205 10 -204
rect 68 -205 69 -204
rect 72 -205 73 -204
rect 121 -205 122 -204
rect 135 -205 136 -204
rect 163 -205 164 -204
rect 30 -207 31 -206
rect 33 -207 34 -206
rect 47 -207 48 -206
rect 268 -207 269 -206
rect 30 -209 31 -208
rect 37 -209 38 -208
rect 51 -209 52 -208
rect 131 -209 132 -208
rect 156 -209 157 -208
rect 254 -209 255 -208
rect 33 -211 34 -210
rect 37 -211 38 -210
rect 54 -211 55 -210
rect 247 -211 248 -210
rect 58 -213 59 -212
rect 89 -213 90 -212
rect 107 -213 108 -212
rect 135 -213 136 -212
rect 156 -213 157 -212
rect 170 -213 171 -212
rect 198 -213 199 -212
rect 247 -213 248 -212
rect 44 -215 45 -214
rect 58 -215 59 -214
rect 75 -215 76 -214
rect 117 -215 118 -214
rect 121 -215 122 -214
rect 142 -215 143 -214
rect 159 -215 160 -214
rect 282 -215 283 -214
rect 86 -217 87 -216
rect 100 -217 101 -216
rect 107 -217 108 -216
rect 149 -217 150 -216
rect 170 -217 171 -216
rect 212 -217 213 -216
rect 23 -219 24 -218
rect 100 -219 101 -218
rect 110 -219 111 -218
rect 219 -219 220 -218
rect 16 -221 17 -220
rect 23 -221 24 -220
rect 40 -221 41 -220
rect 86 -221 87 -220
rect 114 -221 115 -220
rect 205 -221 206 -220
rect 212 -221 213 -220
rect 233 -221 234 -220
rect 16 -223 17 -222
rect 61 -223 62 -222
rect 79 -223 80 -222
rect 114 -223 115 -222
rect 142 -223 143 -222
rect 177 -223 178 -222
rect 198 -223 199 -222
rect 226 -223 227 -222
rect 79 -225 80 -224
rect 93 -225 94 -224
rect 149 -225 150 -224
rect 184 -225 185 -224
rect 205 -225 206 -224
rect 233 -225 234 -224
rect 93 -227 94 -226
rect 128 -227 129 -226
rect 177 -227 178 -226
rect 219 -227 220 -226
rect 226 -227 227 -226
rect 261 -227 262 -226
rect 128 -229 129 -228
rect 275 -229 276 -228
rect 184 -231 185 -230
rect 240 -231 241 -230
rect 194 -233 195 -232
rect 240 -233 241 -232
rect 9 -244 10 -243
rect 93 -244 94 -243
rect 131 -244 132 -243
rect 149 -244 150 -243
rect 159 -244 160 -243
rect 205 -244 206 -243
rect 233 -244 234 -243
rect 240 -244 241 -243
rect 16 -246 17 -245
rect 61 -246 62 -245
rect 68 -246 69 -245
rect 79 -246 80 -245
rect 86 -246 87 -245
rect 93 -246 94 -245
rect 135 -246 136 -245
rect 191 -246 192 -245
rect 194 -246 195 -245
rect 226 -246 227 -245
rect 23 -248 24 -247
rect 65 -248 66 -247
rect 79 -248 80 -247
rect 142 -248 143 -247
rect 149 -248 150 -247
rect 163 -248 164 -247
rect 177 -248 178 -247
rect 247 -248 248 -247
rect 30 -250 31 -249
rect 54 -250 55 -249
rect 65 -250 66 -249
rect 96 -250 97 -249
rect 128 -250 129 -249
rect 135 -250 136 -249
rect 163 -250 164 -249
rect 184 -250 185 -249
rect 212 -250 213 -249
rect 240 -250 241 -249
rect 44 -252 45 -251
rect 72 -252 73 -251
rect 86 -252 87 -251
rect 114 -252 115 -251
rect 128 -252 129 -251
rect 170 -252 171 -251
rect 177 -252 178 -251
rect 198 -252 199 -251
rect 208 -252 209 -251
rect 212 -252 213 -251
rect 44 -254 45 -253
rect 47 -254 48 -253
rect 114 -254 115 -253
rect 121 -254 122 -253
rect 156 -254 157 -253
rect 184 -254 185 -253
rect 198 -254 199 -253
rect 219 -254 220 -253
rect 170 -256 171 -255
rect 226 -256 227 -255
rect 215 -258 216 -257
rect 219 -258 220 -257
rect 44 -269 45 -268
rect 47 -269 48 -268
rect 58 -269 59 -268
rect 65 -269 66 -268
rect 75 -269 76 -268
rect 79 -269 80 -268
rect 86 -269 87 -268
rect 124 -269 125 -268
rect 135 -269 136 -268
rect 138 -269 139 -268
rect 142 -269 143 -268
rect 149 -269 150 -268
rect 163 -269 164 -268
rect 173 -269 174 -268
rect 177 -269 178 -268
rect 194 -269 195 -268
rect 201 -269 202 -268
rect 226 -269 227 -268
rect 79 -271 80 -270
rect 93 -271 94 -270
rect 100 -271 101 -270
rect 103 -271 104 -270
rect 121 -271 122 -270
rect 184 -271 185 -270
rect 191 -271 192 -270
rect 198 -271 199 -270
rect 205 -271 206 -270
rect 233 -271 234 -270
rect 100 -273 101 -272
rect 107 -273 108 -272
rect 114 -273 115 -272
rect 121 -273 122 -272
rect 128 -273 129 -272
rect 142 -273 143 -272
rect 145 -273 146 -272
rect 156 -273 157 -272
rect 205 -273 206 -272
rect 219 -273 220 -272
rect 128 -275 129 -274
rect 159 -275 160 -274
rect 208 -275 209 -274
rect 240 -275 241 -274
rect 65 -286 66 -285
rect 72 -286 73 -285
rect 121 -286 122 -285
rect 131 -286 132 -285
rect 142 -286 143 -285
rect 149 -286 150 -285
<< metal2 >>
rect 107 -3 108 1
rect 128 -3 129 1
rect 114 -3 115 -1
rect 124 -3 125 -1
rect 30 -22 31 -12
rect 40 -22 41 -12
rect 44 -22 45 -12
rect 61 -13 62 -11
rect 65 -22 66 -12
rect 72 -13 73 -11
rect 103 -13 104 -11
rect 135 -22 136 -12
rect 138 -13 139 -11
rect 149 -22 150 -12
rect 156 -22 157 -12
rect 170 -22 171 -12
rect 9 -22 10 -14
rect 61 -22 62 -14
rect 72 -22 73 -14
rect 79 -15 80 -11
rect 93 -22 94 -14
rect 103 -22 104 -14
rect 128 -15 129 -11
rect 142 -22 143 -14
rect 145 -15 146 -11
rect 163 -22 164 -14
rect 54 -22 55 -16
rect 79 -22 80 -16
rect 114 -17 115 -11
rect 128 -22 129 -16
rect 110 -19 111 -11
rect 114 -22 115 -18
rect 110 -22 111 -20
rect 121 -22 122 -20
rect 9 -32 10 -30
rect 54 -32 55 -30
rect 58 -32 59 -30
rect 100 -49 101 -31
rect 110 -32 111 -30
rect 149 -32 150 -30
rect 156 -32 157 -30
rect 156 -49 157 -31
rect 156 -32 157 -30
rect 156 -49 157 -31
rect 163 -32 164 -30
rect 163 -49 164 -31
rect 163 -32 164 -30
rect 163 -49 164 -31
rect 16 -49 17 -33
rect 65 -34 66 -30
rect 68 -49 69 -33
rect 79 -34 80 -30
rect 121 -34 122 -30
rect 149 -49 150 -33
rect 23 -36 24 -30
rect 26 -36 27 -30
rect 30 -36 31 -30
rect 40 -49 41 -35
rect 44 -36 45 -30
rect 79 -49 80 -35
rect 114 -36 115 -30
rect 121 -49 122 -35
rect 128 -36 129 -30
rect 170 -49 171 -35
rect 19 -38 20 -30
rect 23 -49 24 -37
rect 30 -49 31 -37
rect 47 -49 48 -37
rect 54 -49 55 -37
rect 65 -49 66 -37
rect 72 -38 73 -30
rect 86 -38 87 -30
rect 89 -38 90 -30
rect 114 -49 115 -37
rect 142 -38 143 -30
rect 142 -49 143 -37
rect 142 -38 143 -30
rect 142 -49 143 -37
rect 37 -49 38 -39
rect 58 -49 59 -39
rect 61 -40 62 -30
rect 135 -40 136 -30
rect 72 -49 73 -41
rect 128 -49 129 -41
rect 86 -49 87 -43
rect 107 -49 108 -43
rect 93 -46 94 -30
rect 135 -49 136 -45
rect 93 -49 94 -47
rect 177 -49 178 -47
rect 2 -78 3 -58
rect 47 -78 48 -58
rect 51 -59 52 -57
rect 100 -59 101 -57
rect 142 -59 143 -57
rect 198 -78 199 -58
rect 16 -61 17 -57
rect 75 -61 76 -57
rect 82 -78 83 -60
rect 135 -61 136 -57
rect 156 -61 157 -57
rect 191 -78 192 -60
rect 16 -78 17 -62
rect 124 -78 125 -62
rect 135 -78 136 -62
rect 177 -63 178 -57
rect 184 -63 185 -57
rect 184 -78 185 -62
rect 184 -63 185 -57
rect 184 -78 185 -62
rect 26 -78 27 -64
rect 100 -78 101 -64
rect 121 -65 122 -57
rect 156 -78 157 -64
rect 163 -65 164 -57
rect 163 -78 164 -64
rect 163 -65 164 -57
rect 163 -78 164 -64
rect 33 -67 34 -57
rect 33 -78 34 -66
rect 33 -67 34 -57
rect 33 -78 34 -66
rect 37 -78 38 -66
rect 44 -67 45 -57
rect 51 -78 52 -66
rect 142 -78 143 -66
rect 149 -67 150 -57
rect 177 -78 178 -66
rect 9 -69 10 -57
rect 44 -78 45 -68
rect 54 -69 55 -57
rect 72 -78 73 -68
rect 93 -69 94 -57
rect 114 -69 115 -57
rect 23 -71 24 -57
rect 93 -78 94 -70
rect 107 -71 108 -57
rect 149 -78 150 -70
rect 65 -73 66 -57
rect 89 -73 90 -57
rect 114 -78 115 -72
rect 170 -73 171 -57
rect 58 -75 59 -57
rect 65 -78 66 -74
rect 79 -75 80 -57
rect 107 -78 108 -74
rect 128 -75 129 -57
rect 170 -78 171 -74
rect 58 -78 59 -76
rect 79 -78 80 -76
rect 23 -117 24 -87
rect 30 -88 31 -86
rect 37 -88 38 -86
rect 44 -117 45 -87
rect 51 -117 52 -87
rect 58 -88 59 -86
rect 68 -117 69 -87
rect 107 -88 108 -86
rect 114 -88 115 -86
rect 177 -88 178 -86
rect 26 -90 27 -86
rect 65 -90 66 -86
rect 79 -90 80 -86
rect 149 -90 150 -86
rect 163 -90 164 -86
rect 212 -117 213 -89
rect 16 -92 17 -86
rect 79 -117 80 -91
rect 86 -117 87 -91
rect 117 -92 118 -86
rect 124 -92 125 -86
rect 191 -92 192 -86
rect 16 -117 17 -93
rect 93 -94 94 -86
rect 96 -117 97 -93
rect 107 -117 108 -93
rect 128 -117 129 -93
rect 198 -94 199 -86
rect 33 -117 34 -95
rect 149 -117 150 -95
rect 170 -96 171 -86
rect 177 -117 178 -95
rect 184 -96 185 -86
rect 191 -117 192 -95
rect 37 -117 38 -97
rect 121 -117 122 -97
rect 142 -98 143 -86
rect 163 -117 164 -97
rect 58 -117 59 -99
rect 131 -100 132 -86
rect 89 -102 90 -86
rect 135 -102 136 -86
rect 54 -104 55 -86
rect 135 -117 136 -103
rect 93 -117 94 -105
rect 156 -106 157 -86
rect 100 -108 101 -86
rect 156 -117 157 -107
rect 72 -110 73 -86
rect 100 -117 101 -109
rect 117 -117 118 -109
rect 198 -117 199 -109
rect 2 -112 3 -86
rect 72 -117 73 -111
rect 124 -117 125 -111
rect 142 -117 143 -111
rect 2 -117 3 -113
rect 205 -117 206 -113
rect 131 -117 132 -115
rect 184 -117 185 -115
rect 2 -127 3 -125
rect 16 -127 17 -125
rect 23 -127 24 -125
rect 30 -127 31 -125
rect 33 -127 34 -125
rect 124 -127 125 -125
rect 149 -127 150 -125
rect 247 -150 248 -126
rect 2 -150 3 -128
rect 58 -129 59 -125
rect 61 -129 62 -125
rect 100 -129 101 -125
rect 107 -129 108 -125
rect 107 -150 108 -128
rect 107 -129 108 -125
rect 107 -150 108 -128
rect 117 -129 118 -125
rect 128 -150 129 -128
rect 149 -150 150 -128
rect 233 -150 234 -128
rect 9 -131 10 -125
rect 12 -150 13 -130
rect 16 -150 17 -130
rect 47 -150 48 -130
rect 51 -131 52 -125
rect 65 -150 66 -130
rect 72 -131 73 -125
rect 117 -150 118 -130
rect 121 -131 122 -125
rect 212 -131 213 -125
rect 33 -150 34 -132
rect 51 -150 52 -132
rect 58 -150 59 -132
rect 93 -133 94 -125
rect 96 -133 97 -125
rect 198 -133 199 -125
rect 205 -133 206 -125
rect 205 -150 206 -132
rect 205 -133 206 -125
rect 205 -150 206 -132
rect 37 -135 38 -125
rect 72 -150 73 -134
rect 79 -135 80 -125
rect 114 -135 115 -125
rect 121 -150 122 -134
rect 219 -150 220 -134
rect 37 -150 38 -136
rect 44 -137 45 -125
rect 68 -137 69 -125
rect 79 -150 80 -136
rect 86 -137 87 -125
rect 100 -150 101 -136
rect 114 -150 115 -136
rect 226 -150 227 -136
rect 86 -150 87 -138
rect 135 -139 136 -125
rect 152 -150 153 -138
rect 170 -139 171 -125
rect 173 -139 174 -125
rect 212 -150 213 -138
rect 93 -150 94 -140
rect 145 -150 146 -140
rect 156 -141 157 -125
rect 156 -150 157 -140
rect 156 -141 157 -125
rect 156 -150 157 -140
rect 163 -141 164 -125
rect 170 -150 171 -140
rect 191 -141 192 -125
rect 198 -150 199 -140
rect 135 -150 136 -142
rect 240 -150 241 -142
rect 142 -145 143 -125
rect 163 -150 164 -144
rect 184 -145 185 -125
rect 191 -150 192 -144
rect 177 -147 178 -125
rect 184 -150 185 -146
rect 44 -150 45 -148
rect 177 -150 178 -148
rect 5 -193 6 -159
rect 9 -160 10 -158
rect 23 -160 24 -158
rect 51 -160 52 -158
rect 61 -193 62 -159
rect 219 -160 220 -158
rect 233 -160 234 -158
rect 282 -193 283 -159
rect 9 -193 10 -161
rect 16 -162 17 -158
rect 23 -193 24 -161
rect 89 -193 90 -161
rect 117 -162 118 -158
rect 184 -162 185 -158
rect 191 -162 192 -158
rect 233 -193 234 -161
rect 16 -193 17 -163
rect 58 -164 59 -158
rect 75 -193 76 -163
rect 121 -193 122 -163
rect 124 -164 125 -158
rect 149 -193 150 -163
rect 177 -164 178 -158
rect 275 -193 276 -163
rect 26 -166 27 -158
rect 240 -166 241 -158
rect 30 -168 31 -158
rect 268 -193 269 -167
rect 30 -193 31 -169
rect 65 -170 66 -158
rect 79 -170 80 -158
rect 177 -193 178 -169
rect 198 -170 199 -158
rect 240 -193 241 -169
rect 33 -172 34 -158
rect 86 -172 87 -158
rect 117 -193 118 -171
rect 135 -193 136 -171
rect 142 -172 143 -158
rect 163 -172 164 -158
rect 198 -193 199 -171
rect 247 -172 248 -158
rect 2 -174 3 -158
rect 163 -193 164 -173
rect 205 -174 206 -158
rect 254 -193 255 -173
rect 2 -193 3 -175
rect 226 -176 227 -158
rect 37 -178 38 -158
rect 37 -193 38 -177
rect 37 -178 38 -158
rect 37 -193 38 -177
rect 44 -178 45 -158
rect 191 -193 192 -177
rect 212 -178 213 -158
rect 261 -193 262 -177
rect 44 -193 45 -179
rect 110 -193 111 -179
rect 114 -180 115 -158
rect 142 -193 143 -179
rect 152 -180 153 -158
rect 247 -193 248 -179
rect 51 -193 52 -181
rect 184 -193 185 -181
rect 54 -193 55 -183
rect 79 -193 80 -183
rect 96 -184 97 -158
rect 226 -193 227 -183
rect 65 -193 66 -185
rect 93 -186 94 -158
rect 128 -186 129 -158
rect 219 -193 220 -185
rect 72 -188 73 -158
rect 86 -193 87 -187
rect 100 -188 101 -158
rect 128 -193 129 -187
rect 156 -188 157 -158
rect 205 -193 206 -187
rect 72 -193 73 -189
rect 93 -193 94 -189
rect 100 -193 101 -189
rect 107 -190 108 -158
rect 170 -190 171 -158
rect 212 -193 213 -189
rect 107 -193 108 -191
rect 114 -193 115 -191
rect 159 -193 160 -191
rect 170 -193 171 -191
rect 9 -203 10 -201
rect 163 -203 164 -201
rect 180 -234 181 -202
rect 191 -203 192 -201
rect 9 -234 10 -204
rect 68 -205 69 -201
rect 72 -234 73 -204
rect 121 -205 122 -201
rect 135 -205 136 -201
rect 163 -234 164 -204
rect 30 -207 31 -201
rect 33 -211 34 -206
rect 47 -234 48 -206
rect 268 -207 269 -201
rect 30 -234 31 -208
rect 37 -209 38 -201
rect 51 -234 52 -208
rect 131 -234 132 -208
rect 156 -209 157 -201
rect 254 -209 255 -201
rect 37 -234 38 -210
rect 54 -211 55 -201
rect 247 -211 248 -201
rect 58 -213 59 -201
rect 89 -213 90 -201
rect 107 -213 108 -201
rect 135 -234 136 -212
rect 156 -234 157 -212
rect 170 -213 171 -201
rect 198 -213 199 -201
rect 247 -234 248 -212
rect 44 -215 45 -201
rect 58 -234 59 -214
rect 75 -215 76 -201
rect 117 -215 118 -201
rect 121 -234 122 -214
rect 142 -215 143 -201
rect 159 -215 160 -201
rect 282 -215 283 -201
rect 86 -217 87 -201
rect 100 -217 101 -201
rect 107 -234 108 -216
rect 149 -217 150 -201
rect 170 -234 171 -216
rect 212 -217 213 -201
rect 23 -219 24 -201
rect 100 -234 101 -218
rect 110 -219 111 -201
rect 219 -219 220 -201
rect 16 -221 17 -201
rect 23 -234 24 -220
rect 40 -234 41 -220
rect 86 -234 87 -220
rect 114 -221 115 -201
rect 205 -221 206 -201
rect 212 -234 213 -220
rect 233 -221 234 -201
rect 16 -234 17 -222
rect 61 -223 62 -201
rect 79 -223 80 -201
rect 114 -234 115 -222
rect 142 -234 143 -222
rect 177 -223 178 -201
rect 198 -234 199 -222
rect 226 -223 227 -201
rect 79 -234 80 -224
rect 93 -225 94 -201
rect 149 -234 150 -224
rect 184 -225 185 -201
rect 205 -234 206 -224
rect 233 -234 234 -224
rect 93 -234 94 -226
rect 128 -227 129 -201
rect 177 -234 178 -226
rect 219 -234 220 -226
rect 226 -234 227 -226
rect 261 -227 262 -201
rect 128 -234 129 -228
rect 275 -229 276 -201
rect 184 -234 185 -230
rect 240 -231 241 -201
rect 194 -234 195 -232
rect 240 -234 241 -232
rect 9 -244 10 -242
rect 93 -244 94 -242
rect 100 -244 101 -242
rect 100 -259 101 -243
rect 100 -244 101 -242
rect 100 -259 101 -243
rect 107 -244 108 -242
rect 107 -259 108 -243
rect 107 -244 108 -242
rect 107 -259 108 -243
rect 131 -244 132 -242
rect 149 -244 150 -242
rect 159 -259 160 -243
rect 205 -244 206 -242
rect 233 -259 234 -243
rect 240 -244 241 -242
rect 16 -246 17 -242
rect 61 -246 62 -242
rect 68 -246 69 -242
rect 79 -246 80 -242
rect 86 -246 87 -242
rect 93 -259 94 -245
rect 135 -246 136 -242
rect 191 -259 192 -245
rect 194 -246 195 -242
rect 226 -246 227 -242
rect 23 -248 24 -242
rect 65 -248 66 -242
rect 79 -259 80 -247
rect 142 -248 143 -242
rect 149 -259 150 -247
rect 163 -248 164 -242
rect 177 -248 178 -242
rect 247 -248 248 -242
rect 30 -250 31 -242
rect 54 -250 55 -242
rect 58 -250 59 -242
rect 58 -259 59 -249
rect 58 -250 59 -242
rect 58 -259 59 -249
rect 65 -259 66 -249
rect 96 -250 97 -242
rect 128 -250 129 -242
rect 135 -259 136 -249
rect 163 -259 164 -249
rect 184 -250 185 -242
rect 212 -250 213 -242
rect 240 -259 241 -249
rect 44 -252 45 -242
rect 72 -252 73 -242
rect 86 -259 87 -251
rect 114 -252 115 -242
rect 128 -259 129 -251
rect 170 -252 171 -242
rect 177 -259 178 -251
rect 198 -252 199 -242
rect 208 -259 209 -251
rect 212 -259 213 -251
rect 44 -259 45 -253
rect 47 -254 48 -242
rect 114 -259 115 -253
rect 121 -254 122 -242
rect 156 -254 157 -242
rect 184 -259 185 -253
rect 198 -259 199 -253
rect 219 -254 220 -242
rect 170 -259 171 -255
rect 226 -259 227 -255
rect 215 -259 216 -257
rect 219 -259 220 -257
rect 44 -269 45 -267
rect 47 -276 48 -268
rect 58 -269 59 -267
rect 65 -269 66 -267
rect 72 -269 73 -267
rect 72 -276 73 -268
rect 72 -269 73 -267
rect 72 -276 73 -268
rect 75 -269 76 -267
rect 79 -269 80 -267
rect 86 -269 87 -267
rect 124 -269 125 -267
rect 135 -269 136 -267
rect 138 -276 139 -268
rect 142 -269 143 -267
rect 149 -269 150 -267
rect 163 -269 164 -267
rect 173 -269 174 -267
rect 177 -269 178 -267
rect 194 -269 195 -267
rect 201 -276 202 -268
rect 226 -269 227 -267
rect 79 -276 80 -270
rect 93 -271 94 -267
rect 100 -271 101 -267
rect 103 -276 104 -270
rect 121 -271 122 -267
rect 184 -271 185 -267
rect 191 -271 192 -267
rect 198 -271 199 -267
rect 205 -271 206 -267
rect 233 -271 234 -267
rect 100 -276 101 -272
rect 107 -273 108 -267
rect 114 -273 115 -267
rect 121 -276 122 -272
rect 128 -273 129 -267
rect 142 -276 143 -272
rect 145 -273 146 -267
rect 156 -273 157 -267
rect 205 -276 206 -272
rect 219 -273 220 -267
rect 128 -276 129 -274
rect 159 -275 160 -267
rect 208 -276 209 -274
rect 240 -275 241 -267
rect 65 -286 66 -284
rect 72 -286 73 -284
rect 121 -286 122 -284
rect 131 -286 132 -284
rect 142 -286 143 -284
rect 149 -286 150 -284
<< labels >>
rlabel pdiffusion 3 -8 3 -8 0 cellNo=35
rlabel pdiffusion 10 -8 10 -8 0 cellNo=48
rlabel pdiffusion 59 -8 59 -8 0 cellNo=2
rlabel pdiffusion 73 -8 73 -8 0 cellNo=57
rlabel pdiffusion 80 -8 80 -8 0 cellNo=63
rlabel pdiffusion 101 -8 101 -8 0 cellNo=17
rlabel pdiffusion 108 -8 108 -8 0 cellNo=3
rlabel pdiffusion 115 -8 115 -8 0 feedthrough
rlabel pdiffusion 122 -8 122 -8 0 cellNo=62
rlabel pdiffusion 129 -8 129 -8 0 feedthrough
rlabel pdiffusion 136 -8 136 -8 0 cellNo=77
rlabel pdiffusion 143 -8 143 -8 0 cellNo=8
rlabel pdiffusion 3 -27 3 -27 0 cellNo=41
rlabel pdiffusion 10 -27 10 -27 0 feedthrough
rlabel pdiffusion 17 -27 17 -27 0 cellNo=73
rlabel pdiffusion 24 -27 24 -27 0 cellNo=15
rlabel pdiffusion 31 -27 31 -27 0 feedthrough
rlabel pdiffusion 38 -27 38 -27 0 cellNo=31
rlabel pdiffusion 45 -27 45 -27 0 feedthrough
rlabel pdiffusion 52 -27 52 -27 0 cellNo=16
rlabel pdiffusion 59 -27 59 -27 0 cellNo=37
rlabel pdiffusion 66 -27 66 -27 0 feedthrough
rlabel pdiffusion 73 -27 73 -27 0 feedthrough
rlabel pdiffusion 80 -27 80 -27 0 feedthrough
rlabel pdiffusion 87 -27 87 -27 0 cellNo=51
rlabel pdiffusion 94 -27 94 -27 0 feedthrough
rlabel pdiffusion 101 -27 101 -27 0 cellNo=12
rlabel pdiffusion 108 -27 108 -27 0 cellNo=6
rlabel pdiffusion 115 -27 115 -27 0 feedthrough
rlabel pdiffusion 122 -27 122 -27 0 feedthrough
rlabel pdiffusion 129 -27 129 -27 0 feedthrough
rlabel pdiffusion 136 -27 136 -27 0 feedthrough
rlabel pdiffusion 143 -27 143 -27 0 feedthrough
rlabel pdiffusion 150 -27 150 -27 0 feedthrough
rlabel pdiffusion 157 -27 157 -27 0 feedthrough
rlabel pdiffusion 164 -27 164 -27 0 feedthrough
rlabel pdiffusion 171 -27 171 -27 0 cellNo=19
rlabel pdiffusion 10 -54 10 -54 0 cellNo=20
rlabel pdiffusion 17 -54 17 -54 0 feedthrough
rlabel pdiffusion 24 -54 24 -54 0 feedthrough
rlabel pdiffusion 31 -54 31 -54 0 cellNo=22
rlabel pdiffusion 38 -54 38 -54 0 cellNo=47
rlabel pdiffusion 45 -54 45 -54 0 cellNo=81
rlabel pdiffusion 52 -54 52 -54 0 cellNo=4
rlabel pdiffusion 59 -54 59 -54 0 feedthrough
rlabel pdiffusion 66 -54 66 -54 0 cellNo=26
rlabel pdiffusion 73 -54 73 -54 0 cellNo=46
rlabel pdiffusion 80 -54 80 -54 0 feedthrough
rlabel pdiffusion 87 -54 87 -54 0 cellNo=85
rlabel pdiffusion 94 -54 94 -54 0 cellNo=40
rlabel pdiffusion 101 -54 101 -54 0 feedthrough
rlabel pdiffusion 108 -54 108 -54 0 feedthrough
rlabel pdiffusion 115 -54 115 -54 0 feedthrough
rlabel pdiffusion 122 -54 122 -54 0 feedthrough
rlabel pdiffusion 129 -54 129 -54 0 feedthrough
rlabel pdiffusion 136 -54 136 -54 0 feedthrough
rlabel pdiffusion 143 -54 143 -54 0 feedthrough
rlabel pdiffusion 150 -54 150 -54 0 feedthrough
rlabel pdiffusion 157 -54 157 -54 0 feedthrough
rlabel pdiffusion 164 -54 164 -54 0 feedthrough
rlabel pdiffusion 171 -54 171 -54 0 feedthrough
rlabel pdiffusion 178 -54 178 -54 0 feedthrough
rlabel pdiffusion 185 -54 185 -54 0 cellNo=90
rlabel pdiffusion 3 -83 3 -83 0 feedthrough
rlabel pdiffusion 10 -83 10 -83 0 cellNo=69
rlabel pdiffusion 17 -83 17 -83 0 feedthrough
rlabel pdiffusion 24 -83 24 -83 0 cellNo=53
rlabel pdiffusion 31 -83 31 -83 0 cellNo=28
rlabel pdiffusion 38 -83 38 -83 0 feedthrough
rlabel pdiffusion 45 -83 45 -83 0 cellNo=64
rlabel pdiffusion 52 -83 52 -83 0 cellNo=18
rlabel pdiffusion 59 -83 59 -83 0 feedthrough
rlabel pdiffusion 66 -83 66 -83 0 feedthrough
rlabel pdiffusion 73 -83 73 -83 0 feedthrough
rlabel pdiffusion 80 -83 80 -83 0 cellNo=33
rlabel pdiffusion 87 -83 87 -83 0 cellNo=68
rlabel pdiffusion 94 -83 94 -83 0 feedthrough
rlabel pdiffusion 101 -83 101 -83 0 feedthrough
rlabel pdiffusion 108 -83 108 -83 0 feedthrough
rlabel pdiffusion 115 -83 115 -83 0 cellNo=1
rlabel pdiffusion 122 -83 122 -83 0 cellNo=58
rlabel pdiffusion 129 -83 129 -83 0 cellNo=45
rlabel pdiffusion 136 -83 136 -83 0 feedthrough
rlabel pdiffusion 143 -83 143 -83 0 feedthrough
rlabel pdiffusion 150 -83 150 -83 0 feedthrough
rlabel pdiffusion 157 -83 157 -83 0 feedthrough
rlabel pdiffusion 164 -83 164 -83 0 feedthrough
rlabel pdiffusion 171 -83 171 -83 0 feedthrough
rlabel pdiffusion 178 -83 178 -83 0 feedthrough
rlabel pdiffusion 185 -83 185 -83 0 feedthrough
rlabel pdiffusion 192 -83 192 -83 0 feedthrough
rlabel pdiffusion 199 -83 199 -83 0 feedthrough
rlabel pdiffusion 3 -122 3 -122 0 cellNo=11
rlabel pdiffusion 10 -122 10 -122 0 cellNo=21
rlabel pdiffusion 17 -122 17 -122 0 feedthrough
rlabel pdiffusion 24 -122 24 -122 0 feedthrough
rlabel pdiffusion 31 -122 31 -122 0 cellNo=67
rlabel pdiffusion 38 -122 38 -122 0 feedthrough
rlabel pdiffusion 45 -122 45 -122 0 feedthrough
rlabel pdiffusion 52 -122 52 -122 0 feedthrough
rlabel pdiffusion 59 -122 59 -122 0 cellNo=39
rlabel pdiffusion 66 -122 66 -122 0 cellNo=9
rlabel pdiffusion 73 -122 73 -122 0 feedthrough
rlabel pdiffusion 80 -122 80 -122 0 feedthrough
rlabel pdiffusion 87 -122 87 -122 0 feedthrough
rlabel pdiffusion 94 -122 94 -122 0 cellNo=44
rlabel pdiffusion 101 -122 101 -122 0 feedthrough
rlabel pdiffusion 108 -122 108 -122 0 feedthrough
rlabel pdiffusion 115 -122 115 -122 0 cellNo=52
rlabel pdiffusion 122 -122 122 -122 0 cellNo=100
rlabel pdiffusion 129 -122 129 -122 0 cellNo=54
rlabel pdiffusion 136 -122 136 -122 0 feedthrough
rlabel pdiffusion 143 -122 143 -122 0 feedthrough
rlabel pdiffusion 150 -122 150 -122 0 feedthrough
rlabel pdiffusion 157 -122 157 -122 0 feedthrough
rlabel pdiffusion 164 -122 164 -122 0 feedthrough
rlabel pdiffusion 171 -122 171 -122 0 cellNo=86
rlabel pdiffusion 178 -122 178 -122 0 feedthrough
rlabel pdiffusion 185 -122 185 -122 0 feedthrough
rlabel pdiffusion 192 -122 192 -122 0 feedthrough
rlabel pdiffusion 199 -122 199 -122 0 feedthrough
rlabel pdiffusion 206 -122 206 -122 0 feedthrough
rlabel pdiffusion 213 -122 213 -122 0 feedthrough
rlabel pdiffusion 3 -155 3 -155 0 feedthrough
rlabel pdiffusion 10 -155 10 -155 0 cellNo=72
rlabel pdiffusion 17 -155 17 -155 0 feedthrough
rlabel pdiffusion 24 -155 24 -155 0 cellNo=30
rlabel pdiffusion 31 -155 31 -155 0 cellNo=5
rlabel pdiffusion 38 -155 38 -155 0 feedthrough
rlabel pdiffusion 45 -155 45 -155 0 cellNo=74
rlabel pdiffusion 52 -155 52 -155 0 feedthrough
rlabel pdiffusion 59 -155 59 -155 0 feedthrough
rlabel pdiffusion 66 -155 66 -155 0 feedthrough
rlabel pdiffusion 73 -155 73 -155 0 feedthrough
rlabel pdiffusion 80 -155 80 -155 0 feedthrough
rlabel pdiffusion 87 -155 87 -155 0 feedthrough
rlabel pdiffusion 94 -155 94 -155 0 cellNo=7
rlabel pdiffusion 101 -155 101 -155 0 feedthrough
rlabel pdiffusion 108 -155 108 -155 0 feedthrough
rlabel pdiffusion 115 -155 115 -155 0 cellNo=87
rlabel pdiffusion 122 -155 122 -155 0 cellNo=60
rlabel pdiffusion 129 -155 129 -155 0 feedthrough
rlabel pdiffusion 136 -155 136 -155 0 cellNo=34
rlabel pdiffusion 143 -155 143 -155 0 cellNo=56
rlabel pdiffusion 150 -155 150 -155 0 cellNo=10
rlabel pdiffusion 157 -155 157 -155 0 feedthrough
rlabel pdiffusion 164 -155 164 -155 0 feedthrough
rlabel pdiffusion 171 -155 171 -155 0 feedthrough
rlabel pdiffusion 178 -155 178 -155 0 feedthrough
rlabel pdiffusion 185 -155 185 -155 0 feedthrough
rlabel pdiffusion 192 -155 192 -155 0 feedthrough
rlabel pdiffusion 199 -155 199 -155 0 feedthrough
rlabel pdiffusion 206 -155 206 -155 0 feedthrough
rlabel pdiffusion 213 -155 213 -155 0 feedthrough
rlabel pdiffusion 220 -155 220 -155 0 feedthrough
rlabel pdiffusion 227 -155 227 -155 0 feedthrough
rlabel pdiffusion 234 -155 234 -155 0 feedthrough
rlabel pdiffusion 241 -155 241 -155 0 feedthrough
rlabel pdiffusion 248 -155 248 -155 0 feedthrough
rlabel pdiffusion 3 -198 3 -198 0 cellNo=25
rlabel pdiffusion 10 -198 10 -198 0 cellNo=66
rlabel pdiffusion 17 -198 17 -198 0 feedthrough
rlabel pdiffusion 24 -198 24 -198 0 feedthrough
rlabel pdiffusion 31 -198 31 -198 0 feedthrough
rlabel pdiffusion 38 -198 38 -198 0 feedthrough
rlabel pdiffusion 45 -198 45 -198 0 feedthrough
rlabel pdiffusion 52 -198 52 -198 0 cellNo=76
rlabel pdiffusion 59 -198 59 -198 0 cellNo=43
rlabel pdiffusion 66 -198 66 -198 0 cellNo=78
rlabel pdiffusion 73 -198 73 -198 0 cellNo=61
rlabel pdiffusion 80 -198 80 -198 0 feedthrough
rlabel pdiffusion 87 -198 87 -198 0 cellNo=55
rlabel pdiffusion 94 -198 94 -198 0 feedthrough
rlabel pdiffusion 101 -198 101 -198 0 feedthrough
rlabel pdiffusion 108 -198 108 -198 0 cellNo=84
rlabel pdiffusion 115 -198 115 -198 0 cellNo=14
rlabel pdiffusion 122 -198 122 -198 0 feedthrough
rlabel pdiffusion 129 -198 129 -198 0 feedthrough
rlabel pdiffusion 136 -198 136 -198 0 feedthrough
rlabel pdiffusion 143 -198 143 -198 0 feedthrough
rlabel pdiffusion 150 -198 150 -198 0 feedthrough
rlabel pdiffusion 157 -198 157 -198 0 cellNo=82
rlabel pdiffusion 164 -198 164 -198 0 feedthrough
rlabel pdiffusion 171 -198 171 -198 0 feedthrough
rlabel pdiffusion 178 -198 178 -198 0 feedthrough
rlabel pdiffusion 185 -198 185 -198 0 feedthrough
rlabel pdiffusion 192 -198 192 -198 0 feedthrough
rlabel pdiffusion 199 -198 199 -198 0 feedthrough
rlabel pdiffusion 206 -198 206 -198 0 feedthrough
rlabel pdiffusion 213 -198 213 -198 0 feedthrough
rlabel pdiffusion 220 -198 220 -198 0 feedthrough
rlabel pdiffusion 227 -198 227 -198 0 feedthrough
rlabel pdiffusion 234 -198 234 -198 0 feedthrough
rlabel pdiffusion 241 -198 241 -198 0 feedthrough
rlabel pdiffusion 248 -198 248 -198 0 feedthrough
rlabel pdiffusion 255 -198 255 -198 0 feedthrough
rlabel pdiffusion 262 -198 262 -198 0 feedthrough
rlabel pdiffusion 269 -198 269 -198 0 feedthrough
rlabel pdiffusion 276 -198 276 -198 0 feedthrough
rlabel pdiffusion 283 -198 283 -198 0 feedthrough
rlabel pdiffusion 10 -239 10 -239 0 feedthrough
rlabel pdiffusion 17 -239 17 -239 0 feedthrough
rlabel pdiffusion 24 -239 24 -239 0 feedthrough
rlabel pdiffusion 31 -239 31 -239 0 feedthrough
rlabel pdiffusion 38 -239 38 -239 0 cellNo=71
rlabel pdiffusion 45 -239 45 -239 0 cellNo=98
rlabel pdiffusion 52 -239 52 -239 0 cellNo=65
rlabel pdiffusion 59 -239 59 -239 0 cellNo=94
rlabel pdiffusion 66 -239 66 -239 0 cellNo=42
rlabel pdiffusion 73 -239 73 -239 0 feedthrough
rlabel pdiffusion 80 -239 80 -239 0 feedthrough
rlabel pdiffusion 87 -239 87 -239 0 feedthrough
rlabel pdiffusion 94 -239 94 -239 0 cellNo=70
rlabel pdiffusion 101 -239 101 -239 0 feedthrough
rlabel pdiffusion 108 -239 108 -239 0 feedthrough
rlabel pdiffusion 115 -239 115 -239 0 feedthrough
rlabel pdiffusion 122 -239 122 -239 0 feedthrough
rlabel pdiffusion 129 -239 129 -239 0 cellNo=13
rlabel pdiffusion 136 -239 136 -239 0 feedthrough
rlabel pdiffusion 143 -239 143 -239 0 feedthrough
rlabel pdiffusion 150 -239 150 -239 0 feedthrough
rlabel pdiffusion 157 -239 157 -239 0 feedthrough
rlabel pdiffusion 164 -239 164 -239 0 feedthrough
rlabel pdiffusion 171 -239 171 -239 0 feedthrough
rlabel pdiffusion 178 -239 178 -239 0 cellNo=36
rlabel pdiffusion 185 -239 185 -239 0 feedthrough
rlabel pdiffusion 192 -239 192 -239 0 cellNo=23
rlabel pdiffusion 199 -239 199 -239 0 feedthrough
rlabel pdiffusion 206 -239 206 -239 0 feedthrough
rlabel pdiffusion 213 -239 213 -239 0 feedthrough
rlabel pdiffusion 220 -239 220 -239 0 feedthrough
rlabel pdiffusion 227 -239 227 -239 0 feedthrough
rlabel pdiffusion 234 -239 234 -239 0 cellNo=80
rlabel pdiffusion 241 -239 241 -239 0 feedthrough
rlabel pdiffusion 248 -239 248 -239 0 feedthrough
rlabel pdiffusion 3 -264 3 -264 0 cellNo=75
rlabel pdiffusion 45 -264 45 -264 0 feedthrough
rlabel pdiffusion 59 -264 59 -264 0 feedthrough
rlabel pdiffusion 66 -264 66 -264 0 cellNo=29
rlabel pdiffusion 73 -264 73 -264 0 cellNo=59
rlabel pdiffusion 80 -264 80 -264 0 feedthrough
rlabel pdiffusion 87 -264 87 -264 0 feedthrough
rlabel pdiffusion 94 -264 94 -264 0 feedthrough
rlabel pdiffusion 101 -264 101 -264 0 feedthrough
rlabel pdiffusion 108 -264 108 -264 0 feedthrough
rlabel pdiffusion 115 -264 115 -264 0 feedthrough
rlabel pdiffusion 122 -264 122 -264 0 cellNo=93
rlabel pdiffusion 129 -264 129 -264 0 feedthrough
rlabel pdiffusion 136 -264 136 -264 0 feedthrough
rlabel pdiffusion 143 -264 143 -264 0 cellNo=83
rlabel pdiffusion 150 -264 150 -264 0 feedthrough
rlabel pdiffusion 157 -264 157 -264 0 cellNo=38
rlabel pdiffusion 164 -264 164 -264 0 feedthrough
rlabel pdiffusion 171 -264 171 -264 0 cellNo=99
rlabel pdiffusion 178 -264 178 -264 0 feedthrough
rlabel pdiffusion 185 -264 185 -264 0 feedthrough
rlabel pdiffusion 192 -264 192 -264 0 cellNo=88
rlabel pdiffusion 199 -264 199 -264 0 feedthrough
rlabel pdiffusion 206 -264 206 -264 0 cellNo=79
rlabel pdiffusion 213 -264 213 -264 0 cellNo=50
rlabel pdiffusion 220 -264 220 -264 0 feedthrough
rlabel pdiffusion 227 -264 227 -264 0 feedthrough
rlabel pdiffusion 234 -264 234 -264 0 feedthrough
rlabel pdiffusion 241 -264 241 -264 0 feedthrough
rlabel pdiffusion 3 -281 3 -281 0 cellNo=92
rlabel pdiffusion 45 -281 45 -281 0 cellNo=27
rlabel pdiffusion 66 -281 66 -281 0 cellNo=96
rlabel pdiffusion 73 -281 73 -281 0 feedthrough
rlabel pdiffusion 80 -281 80 -281 0 cellNo=97
rlabel pdiffusion 101 -281 101 -281 0 cellNo=32
rlabel pdiffusion 122 -281 122 -281 0 feedthrough
rlabel pdiffusion 129 -281 129 -281 0 cellNo=91
rlabel pdiffusion 136 -281 136 -281 0 cellNo=49
rlabel pdiffusion 143 -281 143 -281 0 feedthrough
rlabel pdiffusion 150 -281 150 -281 0 cellNo=95
rlabel pdiffusion 199 -281 199 -281 0 cellNo=89
rlabel pdiffusion 206 -281 206 -281 0 cellNo=24
rlabel polysilicon 61 -10 61 -10 0 4
rlabel polysilicon 72 -10 72 -10 0 3
rlabel polysilicon 79 -10 79 -10 0 3
rlabel polysilicon 103 -10 103 -10 0 4
rlabel polysilicon 107 -4 107 -4 0 1
rlabel polysilicon 110 -10 110 -10 0 4
rlabel polysilicon 114 -4 114 -4 0 1
rlabel polysilicon 114 -10 114 -10 0 3
rlabel polysilicon 124 -4 124 -4 0 2
rlabel polysilicon 128 -4 128 -4 0 1
rlabel polysilicon 128 -10 128 -10 0 3
rlabel polysilicon 138 -10 138 -10 0 4
rlabel polysilicon 145 -10 145 -10 0 4
rlabel polysilicon 9 -23 9 -23 0 1
rlabel polysilicon 9 -29 9 -29 0 3
rlabel polysilicon 19 -29 19 -29 0 4
rlabel polysilicon 23 -29 23 -29 0 3
rlabel polysilicon 26 -29 26 -29 0 4
rlabel polysilicon 30 -23 30 -23 0 1
rlabel polysilicon 30 -29 30 -29 0 3
rlabel polysilicon 40 -23 40 -23 0 2
rlabel polysilicon 44 -23 44 -23 0 1
rlabel polysilicon 44 -29 44 -29 0 3
rlabel polysilicon 54 -23 54 -23 0 2
rlabel polysilicon 54 -29 54 -29 0 4
rlabel polysilicon 61 -23 61 -23 0 2
rlabel polysilicon 58 -29 58 -29 0 3
rlabel polysilicon 61 -29 61 -29 0 4
rlabel polysilicon 65 -23 65 -23 0 1
rlabel polysilicon 65 -29 65 -29 0 3
rlabel polysilicon 72 -23 72 -23 0 1
rlabel polysilicon 72 -29 72 -29 0 3
rlabel polysilicon 79 -23 79 -23 0 1
rlabel polysilicon 79 -29 79 -29 0 3
rlabel polysilicon 86 -29 86 -29 0 3
rlabel polysilicon 89 -29 89 -29 0 4
rlabel polysilicon 93 -23 93 -23 0 1
rlabel polysilicon 93 -29 93 -29 0 3
rlabel polysilicon 103 -23 103 -23 0 2
rlabel polysilicon 110 -23 110 -23 0 2
rlabel polysilicon 110 -29 110 -29 0 4
rlabel polysilicon 114 -23 114 -23 0 1
rlabel polysilicon 114 -29 114 -29 0 3
rlabel polysilicon 121 -23 121 -23 0 1
rlabel polysilicon 121 -29 121 -29 0 3
rlabel polysilicon 128 -23 128 -23 0 1
rlabel polysilicon 128 -29 128 -29 0 3
rlabel polysilicon 135 -23 135 -23 0 1
rlabel polysilicon 135 -29 135 -29 0 3
rlabel polysilicon 142 -23 142 -23 0 1
rlabel polysilicon 142 -29 142 -29 0 3
rlabel polysilicon 149 -23 149 -23 0 1
rlabel polysilicon 149 -29 149 -29 0 3
rlabel polysilicon 156 -23 156 -23 0 1
rlabel polysilicon 156 -29 156 -29 0 3
rlabel polysilicon 163 -23 163 -23 0 1
rlabel polysilicon 163 -29 163 -29 0 3
rlabel polysilicon 170 -23 170 -23 0 1
rlabel polysilicon 9 -56 9 -56 0 3
rlabel polysilicon 16 -50 16 -50 0 1
rlabel polysilicon 16 -56 16 -56 0 3
rlabel polysilicon 23 -50 23 -50 0 1
rlabel polysilicon 23 -56 23 -56 0 3
rlabel polysilicon 30 -50 30 -50 0 1
rlabel polysilicon 33 -56 33 -56 0 4
rlabel polysilicon 37 -50 37 -50 0 1
rlabel polysilicon 40 -50 40 -50 0 2
rlabel polysilicon 47 -50 47 -50 0 2
rlabel polysilicon 44 -56 44 -56 0 3
rlabel polysilicon 54 -50 54 -50 0 2
rlabel polysilicon 51 -56 51 -56 0 3
rlabel polysilicon 54 -56 54 -56 0 4
rlabel polysilicon 58 -50 58 -50 0 1
rlabel polysilicon 58 -56 58 -56 0 3
rlabel polysilicon 65 -50 65 -50 0 1
rlabel polysilicon 68 -50 68 -50 0 2
rlabel polysilicon 65 -56 65 -56 0 3
rlabel polysilicon 72 -50 72 -50 0 1
rlabel polysilicon 75 -56 75 -56 0 4
rlabel polysilicon 79 -50 79 -50 0 1
rlabel polysilicon 79 -56 79 -56 0 3
rlabel polysilicon 86 -50 86 -50 0 1
rlabel polysilicon 89 -56 89 -56 0 4
rlabel polysilicon 93 -50 93 -50 0 1
rlabel polysilicon 93 -56 93 -56 0 3
rlabel polysilicon 100 -50 100 -50 0 1
rlabel polysilicon 100 -56 100 -56 0 3
rlabel polysilicon 107 -50 107 -50 0 1
rlabel polysilicon 107 -56 107 -56 0 3
rlabel polysilicon 114 -50 114 -50 0 1
rlabel polysilicon 114 -56 114 -56 0 3
rlabel polysilicon 121 -50 121 -50 0 1
rlabel polysilicon 121 -56 121 -56 0 3
rlabel polysilicon 128 -50 128 -50 0 1
rlabel polysilicon 128 -56 128 -56 0 3
rlabel polysilicon 135 -50 135 -50 0 1
rlabel polysilicon 135 -56 135 -56 0 3
rlabel polysilicon 142 -50 142 -50 0 1
rlabel polysilicon 142 -56 142 -56 0 3
rlabel polysilicon 149 -50 149 -50 0 1
rlabel polysilicon 149 -56 149 -56 0 3
rlabel polysilicon 156 -50 156 -50 0 1
rlabel polysilicon 156 -56 156 -56 0 3
rlabel polysilicon 163 -50 163 -50 0 1
rlabel polysilicon 163 -56 163 -56 0 3
rlabel polysilicon 170 -50 170 -50 0 1
rlabel polysilicon 170 -56 170 -56 0 3
rlabel polysilicon 177 -50 177 -50 0 1
rlabel polysilicon 177 -56 177 -56 0 3
rlabel polysilicon 184 -56 184 -56 0 3
rlabel polysilicon 2 -79 2 -79 0 1
rlabel polysilicon 2 -85 2 -85 0 3
rlabel polysilicon 16 -79 16 -79 0 1
rlabel polysilicon 16 -85 16 -85 0 3
rlabel polysilicon 26 -79 26 -79 0 2
rlabel polysilicon 26 -85 26 -85 0 4
rlabel polysilicon 33 -79 33 -79 0 2
rlabel polysilicon 30 -85 30 -85 0 3
rlabel polysilicon 37 -79 37 -79 0 1
rlabel polysilicon 37 -85 37 -85 0 3
rlabel polysilicon 44 -79 44 -79 0 1
rlabel polysilicon 47 -79 47 -79 0 2
rlabel polysilicon 51 -79 51 -79 0 1
rlabel polysilicon 54 -85 54 -85 0 4
rlabel polysilicon 58 -79 58 -79 0 1
rlabel polysilicon 58 -85 58 -85 0 3
rlabel polysilicon 65 -79 65 -79 0 1
rlabel polysilicon 65 -85 65 -85 0 3
rlabel polysilicon 72 -79 72 -79 0 1
rlabel polysilicon 72 -85 72 -85 0 3
rlabel polysilicon 79 -79 79 -79 0 1
rlabel polysilicon 82 -79 82 -79 0 2
rlabel polysilicon 79 -85 79 -85 0 3
rlabel polysilicon 89 -85 89 -85 0 4
rlabel polysilicon 93 -79 93 -79 0 1
rlabel polysilicon 93 -85 93 -85 0 3
rlabel polysilicon 100 -79 100 -79 0 1
rlabel polysilicon 100 -85 100 -85 0 3
rlabel polysilicon 107 -79 107 -79 0 1
rlabel polysilicon 107 -85 107 -85 0 3
rlabel polysilicon 114 -79 114 -79 0 1
rlabel polysilicon 114 -85 114 -85 0 3
rlabel polysilicon 117 -85 117 -85 0 4
rlabel polysilicon 124 -79 124 -79 0 2
rlabel polysilicon 124 -85 124 -85 0 4
rlabel polysilicon 131 -85 131 -85 0 4
rlabel polysilicon 135 -79 135 -79 0 1
rlabel polysilicon 135 -85 135 -85 0 3
rlabel polysilicon 142 -79 142 -79 0 1
rlabel polysilicon 142 -85 142 -85 0 3
rlabel polysilicon 149 -79 149 -79 0 1
rlabel polysilicon 149 -85 149 -85 0 3
rlabel polysilicon 156 -79 156 -79 0 1
rlabel polysilicon 156 -85 156 -85 0 3
rlabel polysilicon 163 -79 163 -79 0 1
rlabel polysilicon 163 -85 163 -85 0 3
rlabel polysilicon 170 -79 170 -79 0 1
rlabel polysilicon 170 -85 170 -85 0 3
rlabel polysilicon 177 -79 177 -79 0 1
rlabel polysilicon 177 -85 177 -85 0 3
rlabel polysilicon 184 -79 184 -79 0 1
rlabel polysilicon 184 -85 184 -85 0 3
rlabel polysilicon 191 -79 191 -79 0 1
rlabel polysilicon 191 -85 191 -85 0 3
rlabel polysilicon 198 -79 198 -79 0 1
rlabel polysilicon 198 -85 198 -85 0 3
rlabel polysilicon 2 -118 2 -118 0 1
rlabel polysilicon 2 -124 2 -124 0 3
rlabel polysilicon 9 -124 9 -124 0 3
rlabel polysilicon 16 -118 16 -118 0 1
rlabel polysilicon 16 -124 16 -124 0 3
rlabel polysilicon 23 -118 23 -118 0 1
rlabel polysilicon 23 -124 23 -124 0 3
rlabel polysilicon 33 -118 33 -118 0 2
rlabel polysilicon 30 -124 30 -124 0 3
rlabel polysilicon 33 -124 33 -124 0 4
rlabel polysilicon 37 -118 37 -118 0 1
rlabel polysilicon 37 -124 37 -124 0 3
rlabel polysilicon 44 -118 44 -118 0 1
rlabel polysilicon 44 -124 44 -124 0 3
rlabel polysilicon 51 -118 51 -118 0 1
rlabel polysilicon 51 -124 51 -124 0 3
rlabel polysilicon 58 -118 58 -118 0 1
rlabel polysilicon 58 -124 58 -124 0 3
rlabel polysilicon 61 -124 61 -124 0 4
rlabel polysilicon 68 -118 68 -118 0 2
rlabel polysilicon 68 -124 68 -124 0 4
rlabel polysilicon 72 -118 72 -118 0 1
rlabel polysilicon 72 -124 72 -124 0 3
rlabel polysilicon 79 -118 79 -118 0 1
rlabel polysilicon 79 -124 79 -124 0 3
rlabel polysilicon 86 -118 86 -118 0 1
rlabel polysilicon 86 -124 86 -124 0 3
rlabel polysilicon 93 -118 93 -118 0 1
rlabel polysilicon 96 -118 96 -118 0 2
rlabel polysilicon 93 -124 93 -124 0 3
rlabel polysilicon 96 -124 96 -124 0 4
rlabel polysilicon 100 -118 100 -118 0 1
rlabel polysilicon 100 -124 100 -124 0 3
rlabel polysilicon 107 -118 107 -118 0 1
rlabel polysilicon 107 -124 107 -124 0 3
rlabel polysilicon 117 -118 117 -118 0 2
rlabel polysilicon 114 -124 114 -124 0 3
rlabel polysilicon 117 -124 117 -124 0 4
rlabel polysilicon 121 -118 121 -118 0 1
rlabel polysilicon 124 -118 124 -118 0 2
rlabel polysilicon 121 -124 121 -124 0 3
rlabel polysilicon 124 -124 124 -124 0 4
rlabel polysilicon 128 -118 128 -118 0 1
rlabel polysilicon 131 -118 131 -118 0 2
rlabel polysilicon 135 -118 135 -118 0 1
rlabel polysilicon 135 -124 135 -124 0 3
rlabel polysilicon 142 -118 142 -118 0 1
rlabel polysilicon 142 -124 142 -124 0 3
rlabel polysilicon 149 -118 149 -118 0 1
rlabel polysilicon 149 -124 149 -124 0 3
rlabel polysilicon 156 -118 156 -118 0 1
rlabel polysilicon 156 -124 156 -124 0 3
rlabel polysilicon 163 -118 163 -118 0 1
rlabel polysilicon 163 -124 163 -124 0 3
rlabel polysilicon 170 -124 170 -124 0 3
rlabel polysilicon 173 -124 173 -124 0 4
rlabel polysilicon 177 -118 177 -118 0 1
rlabel polysilicon 177 -124 177 -124 0 3
rlabel polysilicon 184 -118 184 -118 0 1
rlabel polysilicon 184 -124 184 -124 0 3
rlabel polysilicon 191 -118 191 -118 0 1
rlabel polysilicon 191 -124 191 -124 0 3
rlabel polysilicon 198 -118 198 -118 0 1
rlabel polysilicon 198 -124 198 -124 0 3
rlabel polysilicon 205 -118 205 -118 0 1
rlabel polysilicon 205 -124 205 -124 0 3
rlabel polysilicon 212 -118 212 -118 0 1
rlabel polysilicon 212 -124 212 -124 0 3
rlabel polysilicon 2 -151 2 -151 0 1
rlabel polysilicon 2 -157 2 -157 0 3
rlabel polysilicon 12 -151 12 -151 0 2
rlabel polysilicon 9 -157 9 -157 0 3
rlabel polysilicon 16 -151 16 -151 0 1
rlabel polysilicon 16 -157 16 -157 0 3
rlabel polysilicon 23 -157 23 -157 0 3
rlabel polysilicon 26 -157 26 -157 0 4
rlabel polysilicon 33 -151 33 -151 0 2
rlabel polysilicon 30 -157 30 -157 0 3
rlabel polysilicon 33 -157 33 -157 0 4
rlabel polysilicon 37 -151 37 -151 0 1
rlabel polysilicon 37 -157 37 -157 0 3
rlabel polysilicon 44 -151 44 -151 0 1
rlabel polysilicon 47 -151 47 -151 0 2
rlabel polysilicon 44 -157 44 -157 0 3
rlabel polysilicon 51 -151 51 -151 0 1
rlabel polysilicon 51 -157 51 -157 0 3
rlabel polysilicon 58 -151 58 -151 0 1
rlabel polysilicon 58 -157 58 -157 0 3
rlabel polysilicon 65 -151 65 -151 0 1
rlabel polysilicon 65 -157 65 -157 0 3
rlabel polysilicon 72 -151 72 -151 0 1
rlabel polysilicon 72 -157 72 -157 0 3
rlabel polysilicon 79 -151 79 -151 0 1
rlabel polysilicon 79 -157 79 -157 0 3
rlabel polysilicon 86 -151 86 -151 0 1
rlabel polysilicon 86 -157 86 -157 0 3
rlabel polysilicon 93 -151 93 -151 0 1
rlabel polysilicon 93 -157 93 -157 0 3
rlabel polysilicon 96 -157 96 -157 0 4
rlabel polysilicon 100 -151 100 -151 0 1
rlabel polysilicon 100 -157 100 -157 0 3
rlabel polysilicon 107 -151 107 -151 0 1
rlabel polysilicon 107 -157 107 -157 0 3
rlabel polysilicon 114 -151 114 -151 0 1
rlabel polysilicon 117 -151 117 -151 0 2
rlabel polysilicon 114 -157 114 -157 0 3
rlabel polysilicon 117 -157 117 -157 0 4
rlabel polysilicon 121 -151 121 -151 0 1
rlabel polysilicon 124 -157 124 -157 0 4
rlabel polysilicon 128 -151 128 -151 0 1
rlabel polysilicon 128 -157 128 -157 0 3
rlabel polysilicon 135 -151 135 -151 0 1
rlabel polysilicon 145 -151 145 -151 0 2
rlabel polysilicon 142 -157 142 -157 0 3
rlabel polysilicon 149 -151 149 -151 0 1
rlabel polysilicon 152 -151 152 -151 0 2
rlabel polysilicon 152 -157 152 -157 0 4
rlabel polysilicon 156 -151 156 -151 0 1
rlabel polysilicon 156 -157 156 -157 0 3
rlabel polysilicon 163 -151 163 -151 0 1
rlabel polysilicon 163 -157 163 -157 0 3
rlabel polysilicon 170 -151 170 -151 0 1
rlabel polysilicon 170 -157 170 -157 0 3
rlabel polysilicon 177 -151 177 -151 0 1
rlabel polysilicon 177 -157 177 -157 0 3
rlabel polysilicon 184 -151 184 -151 0 1
rlabel polysilicon 184 -157 184 -157 0 3
rlabel polysilicon 191 -151 191 -151 0 1
rlabel polysilicon 191 -157 191 -157 0 3
rlabel polysilicon 198 -151 198 -151 0 1
rlabel polysilicon 198 -157 198 -157 0 3
rlabel polysilicon 205 -151 205 -151 0 1
rlabel polysilicon 205 -157 205 -157 0 3
rlabel polysilicon 212 -151 212 -151 0 1
rlabel polysilicon 212 -157 212 -157 0 3
rlabel polysilicon 219 -151 219 -151 0 1
rlabel polysilicon 219 -157 219 -157 0 3
rlabel polysilicon 226 -151 226 -151 0 1
rlabel polysilicon 226 -157 226 -157 0 3
rlabel polysilicon 233 -151 233 -151 0 1
rlabel polysilicon 233 -157 233 -157 0 3
rlabel polysilicon 240 -151 240 -151 0 1
rlabel polysilicon 240 -157 240 -157 0 3
rlabel polysilicon 247 -151 247 -151 0 1
rlabel polysilicon 247 -157 247 -157 0 3
rlabel polysilicon 2 -194 2 -194 0 1
rlabel polysilicon 5 -194 5 -194 0 2
rlabel polysilicon 9 -194 9 -194 0 1
rlabel polysilicon 9 -200 9 -200 0 3
rlabel polysilicon 16 -194 16 -194 0 1
rlabel polysilicon 16 -200 16 -200 0 3
rlabel polysilicon 23 -194 23 -194 0 1
rlabel polysilicon 23 -200 23 -200 0 3
rlabel polysilicon 30 -194 30 -194 0 1
rlabel polysilicon 30 -200 30 -200 0 3
rlabel polysilicon 37 -194 37 -194 0 1
rlabel polysilicon 37 -200 37 -200 0 3
rlabel polysilicon 44 -194 44 -194 0 1
rlabel polysilicon 44 -200 44 -200 0 3
rlabel polysilicon 51 -194 51 -194 0 1
rlabel polysilicon 54 -194 54 -194 0 2
rlabel polysilicon 54 -200 54 -200 0 4
rlabel polysilicon 61 -194 61 -194 0 2
rlabel polysilicon 58 -200 58 -200 0 3
rlabel polysilicon 61 -200 61 -200 0 4
rlabel polysilicon 65 -194 65 -194 0 1
rlabel polysilicon 68 -200 68 -200 0 4
rlabel polysilicon 72 -194 72 -194 0 1
rlabel polysilicon 75 -194 75 -194 0 2
rlabel polysilicon 75 -200 75 -200 0 4
rlabel polysilicon 79 -194 79 -194 0 1
rlabel polysilicon 79 -200 79 -200 0 3
rlabel polysilicon 86 -194 86 -194 0 1
rlabel polysilicon 89 -194 89 -194 0 2
rlabel polysilicon 86 -200 86 -200 0 3
rlabel polysilicon 89 -200 89 -200 0 4
rlabel polysilicon 93 -194 93 -194 0 1
rlabel polysilicon 93 -200 93 -200 0 3
rlabel polysilicon 100 -194 100 -194 0 1
rlabel polysilicon 100 -200 100 -200 0 3
rlabel polysilicon 107 -194 107 -194 0 1
rlabel polysilicon 110 -194 110 -194 0 2
rlabel polysilicon 107 -200 107 -200 0 3
rlabel polysilicon 110 -200 110 -200 0 4
rlabel polysilicon 114 -194 114 -194 0 1
rlabel polysilicon 117 -194 117 -194 0 2
rlabel polysilicon 114 -200 114 -200 0 3
rlabel polysilicon 117 -200 117 -200 0 4
rlabel polysilicon 121 -194 121 -194 0 1
rlabel polysilicon 121 -200 121 -200 0 3
rlabel polysilicon 128 -194 128 -194 0 1
rlabel polysilicon 128 -200 128 -200 0 3
rlabel polysilicon 135 -194 135 -194 0 1
rlabel polysilicon 135 -200 135 -200 0 3
rlabel polysilicon 142 -194 142 -194 0 1
rlabel polysilicon 142 -200 142 -200 0 3
rlabel polysilicon 149 -194 149 -194 0 1
rlabel polysilicon 149 -200 149 -200 0 3
rlabel polysilicon 159 -194 159 -194 0 2
rlabel polysilicon 156 -200 156 -200 0 3
rlabel polysilicon 159 -200 159 -200 0 4
rlabel polysilicon 163 -194 163 -194 0 1
rlabel polysilicon 163 -200 163 -200 0 3
rlabel polysilicon 170 -194 170 -194 0 1
rlabel polysilicon 170 -200 170 -200 0 3
rlabel polysilicon 177 -194 177 -194 0 1
rlabel polysilicon 177 -200 177 -200 0 3
rlabel polysilicon 184 -194 184 -194 0 1
rlabel polysilicon 184 -200 184 -200 0 3
rlabel polysilicon 191 -194 191 -194 0 1
rlabel polysilicon 191 -200 191 -200 0 3
rlabel polysilicon 198 -194 198 -194 0 1
rlabel polysilicon 198 -200 198 -200 0 3
rlabel polysilicon 205 -194 205 -194 0 1
rlabel polysilicon 205 -200 205 -200 0 3
rlabel polysilicon 212 -194 212 -194 0 1
rlabel polysilicon 212 -200 212 -200 0 3
rlabel polysilicon 219 -194 219 -194 0 1
rlabel polysilicon 219 -200 219 -200 0 3
rlabel polysilicon 226 -194 226 -194 0 1
rlabel polysilicon 226 -200 226 -200 0 3
rlabel polysilicon 233 -194 233 -194 0 1
rlabel polysilicon 233 -200 233 -200 0 3
rlabel polysilicon 240 -194 240 -194 0 1
rlabel polysilicon 240 -200 240 -200 0 3
rlabel polysilicon 247 -194 247 -194 0 1
rlabel polysilicon 247 -200 247 -200 0 3
rlabel polysilicon 254 -194 254 -194 0 1
rlabel polysilicon 254 -200 254 -200 0 3
rlabel polysilicon 261 -194 261 -194 0 1
rlabel polysilicon 261 -200 261 -200 0 3
rlabel polysilicon 268 -194 268 -194 0 1
rlabel polysilicon 268 -200 268 -200 0 3
rlabel polysilicon 275 -194 275 -194 0 1
rlabel polysilicon 275 -200 275 -200 0 3
rlabel polysilicon 282 -194 282 -194 0 1
rlabel polysilicon 282 -200 282 -200 0 3
rlabel polysilicon 9 -235 9 -235 0 1
rlabel polysilicon 9 -241 9 -241 0 3
rlabel polysilicon 16 -235 16 -235 0 1
rlabel polysilicon 16 -241 16 -241 0 3
rlabel polysilicon 23 -235 23 -235 0 1
rlabel polysilicon 23 -241 23 -241 0 3
rlabel polysilicon 30 -235 30 -235 0 1
rlabel polysilicon 30 -241 30 -241 0 3
rlabel polysilicon 37 -235 37 -235 0 1
rlabel polysilicon 40 -235 40 -235 0 2
rlabel polysilicon 47 -235 47 -235 0 2
rlabel polysilicon 44 -241 44 -241 0 3
rlabel polysilicon 47 -241 47 -241 0 4
rlabel polysilicon 51 -235 51 -235 0 1
rlabel polysilicon 54 -241 54 -241 0 4
rlabel polysilicon 58 -235 58 -235 0 1
rlabel polysilicon 58 -241 58 -241 0 3
rlabel polysilicon 61 -241 61 -241 0 4
rlabel polysilicon 65 -241 65 -241 0 3
rlabel polysilicon 68 -241 68 -241 0 4
rlabel polysilicon 72 -235 72 -235 0 1
rlabel polysilicon 72 -241 72 -241 0 3
rlabel polysilicon 79 -235 79 -235 0 1
rlabel polysilicon 79 -241 79 -241 0 3
rlabel polysilicon 86 -235 86 -235 0 1
rlabel polysilicon 86 -241 86 -241 0 3
rlabel polysilicon 93 -235 93 -235 0 1
rlabel polysilicon 93 -241 93 -241 0 3
rlabel polysilicon 96 -241 96 -241 0 4
rlabel polysilicon 100 -235 100 -235 0 1
rlabel polysilicon 100 -241 100 -241 0 3
rlabel polysilicon 107 -235 107 -235 0 1
rlabel polysilicon 107 -241 107 -241 0 3
rlabel polysilicon 114 -235 114 -235 0 1
rlabel polysilicon 114 -241 114 -241 0 3
rlabel polysilicon 121 -235 121 -235 0 1
rlabel polysilicon 121 -241 121 -241 0 3
rlabel polysilicon 128 -235 128 -235 0 1
rlabel polysilicon 131 -235 131 -235 0 2
rlabel polysilicon 128 -241 128 -241 0 3
rlabel polysilicon 131 -241 131 -241 0 4
rlabel polysilicon 135 -235 135 -235 0 1
rlabel polysilicon 135 -241 135 -241 0 3
rlabel polysilicon 142 -235 142 -235 0 1
rlabel polysilicon 142 -241 142 -241 0 3
rlabel polysilicon 149 -235 149 -235 0 1
rlabel polysilicon 149 -241 149 -241 0 3
rlabel polysilicon 156 -235 156 -235 0 1
rlabel polysilicon 156 -241 156 -241 0 3
rlabel polysilicon 163 -235 163 -235 0 1
rlabel polysilicon 163 -241 163 -241 0 3
rlabel polysilicon 170 -235 170 -235 0 1
rlabel polysilicon 170 -241 170 -241 0 3
rlabel polysilicon 177 -235 177 -235 0 1
rlabel polysilicon 180 -235 180 -235 0 2
rlabel polysilicon 177 -241 177 -241 0 3
rlabel polysilicon 184 -235 184 -235 0 1
rlabel polysilicon 184 -241 184 -241 0 3
rlabel polysilicon 194 -235 194 -235 0 2
rlabel polysilicon 194 -241 194 -241 0 4
rlabel polysilicon 198 -235 198 -235 0 1
rlabel polysilicon 198 -241 198 -241 0 3
rlabel polysilicon 205 -235 205 -235 0 1
rlabel polysilicon 205 -241 205 -241 0 3
rlabel polysilicon 212 -235 212 -235 0 1
rlabel polysilicon 212 -241 212 -241 0 3
rlabel polysilicon 219 -235 219 -235 0 1
rlabel polysilicon 219 -241 219 -241 0 3
rlabel polysilicon 226 -235 226 -235 0 1
rlabel polysilicon 226 -241 226 -241 0 3
rlabel polysilicon 233 -235 233 -235 0 1
rlabel polysilicon 240 -235 240 -235 0 1
rlabel polysilicon 240 -241 240 -241 0 3
rlabel polysilicon 247 -235 247 -235 0 1
rlabel polysilicon 247 -241 247 -241 0 3
rlabel polysilicon 44 -260 44 -260 0 1
rlabel polysilicon 44 -266 44 -266 0 3
rlabel polysilicon 58 -260 58 -260 0 1
rlabel polysilicon 58 -266 58 -266 0 3
rlabel polysilicon 65 -260 65 -260 0 1
rlabel polysilicon 65 -266 65 -266 0 3
rlabel polysilicon 72 -266 72 -266 0 3
rlabel polysilicon 75 -266 75 -266 0 4
rlabel polysilicon 79 -260 79 -260 0 1
rlabel polysilicon 79 -266 79 -266 0 3
rlabel polysilicon 86 -260 86 -260 0 1
rlabel polysilicon 86 -266 86 -266 0 3
rlabel polysilicon 93 -260 93 -260 0 1
rlabel polysilicon 93 -266 93 -266 0 3
rlabel polysilicon 100 -260 100 -260 0 1
rlabel polysilicon 100 -266 100 -266 0 3
rlabel polysilicon 107 -260 107 -260 0 1
rlabel polysilicon 107 -266 107 -266 0 3
rlabel polysilicon 114 -260 114 -260 0 1
rlabel polysilicon 114 -266 114 -266 0 3
rlabel polysilicon 121 -266 121 -266 0 3
rlabel polysilicon 124 -266 124 -266 0 4
rlabel polysilicon 128 -260 128 -260 0 1
rlabel polysilicon 128 -266 128 -266 0 3
rlabel polysilicon 135 -260 135 -260 0 1
rlabel polysilicon 135 -266 135 -266 0 3
rlabel polysilicon 142 -266 142 -266 0 3
rlabel polysilicon 145 -266 145 -266 0 4
rlabel polysilicon 149 -260 149 -260 0 1
rlabel polysilicon 149 -266 149 -266 0 3
rlabel polysilicon 159 -260 159 -260 0 2
rlabel polysilicon 156 -266 156 -266 0 3
rlabel polysilicon 159 -266 159 -266 0 4
rlabel polysilicon 163 -260 163 -260 0 1
rlabel polysilicon 163 -266 163 -266 0 3
rlabel polysilicon 170 -260 170 -260 0 1
rlabel polysilicon 173 -266 173 -266 0 4
rlabel polysilicon 177 -260 177 -260 0 1
rlabel polysilicon 177 -266 177 -266 0 3
rlabel polysilicon 184 -260 184 -260 0 1
rlabel polysilicon 184 -266 184 -266 0 3
rlabel polysilicon 191 -260 191 -260 0 1
rlabel polysilicon 191 -266 191 -266 0 3
rlabel polysilicon 194 -266 194 -266 0 4
rlabel polysilicon 198 -260 198 -260 0 1
rlabel polysilicon 198 -266 198 -266 0 3
rlabel polysilicon 208 -260 208 -260 0 2
rlabel polysilicon 205 -266 205 -266 0 3
rlabel polysilicon 212 -260 212 -260 0 1
rlabel polysilicon 215 -260 215 -260 0 2
rlabel polysilicon 219 -260 219 -260 0 1
rlabel polysilicon 219 -266 219 -266 0 3
rlabel polysilicon 226 -260 226 -260 0 1
rlabel polysilicon 226 -266 226 -266 0 3
rlabel polysilicon 233 -260 233 -260 0 1
rlabel polysilicon 233 -266 233 -266 0 3
rlabel polysilicon 240 -260 240 -260 0 1
rlabel polysilicon 240 -266 240 -266 0 3
rlabel polysilicon 47 -277 47 -277 0 2
rlabel polysilicon 65 -283 65 -283 0 3
rlabel polysilicon 72 -277 72 -277 0 1
rlabel polysilicon 72 -283 72 -283 0 3
rlabel polysilicon 79 -277 79 -277 0 1
rlabel polysilicon 100 -277 100 -277 0 1
rlabel polysilicon 103 -277 103 -277 0 2
rlabel polysilicon 121 -277 121 -277 0 1
rlabel polysilicon 121 -283 121 -283 0 3
rlabel polysilicon 128 -277 128 -277 0 1
rlabel polysilicon 131 -283 131 -283 0 4
rlabel polysilicon 138 -277 138 -277 0 2
rlabel polysilicon 142 -277 142 -277 0 1
rlabel polysilicon 142 -283 142 -283 0 3
rlabel polysilicon 149 -283 149 -283 0 3
rlabel polysilicon 201 -277 201 -277 0 2
rlabel polysilicon 205 -277 205 -277 0 1
rlabel polysilicon 208 -277 208 -277 0 2
rlabel metal2 107 1 107 1 0 net=349
rlabel metal2 114 -1 114 -1 0 net=393
rlabel metal2 30 -12 30 -12 0 net=185
rlabel metal2 44 -12 44 -12 0 net=179
rlabel metal2 65 -12 65 -12 0 net=171
rlabel metal2 103 -12 103 -12 0 net=269
rlabel metal2 138 -12 138 -12 0 net=289
rlabel metal2 156 -12 156 -12 0 net=399
rlabel metal2 9 -14 9 -14 0 net=237
rlabel metal2 72 -14 72 -14 0 net=251
rlabel metal2 93 -14 93 -14 0 net=299
rlabel metal2 128 -14 128 -14 0 net=351
rlabel metal2 145 -14 145 -14 0 net=437
rlabel metal2 54 -16 54 -16 0 net=197
rlabel metal2 114 -16 114 -16 0 net=395
rlabel metal2 110 -18 110 -18 0 net=343
rlabel metal2 110 -20 110 -20 0 net=365
rlabel metal2 9 -31 9 -31 0 net=238
rlabel metal2 58 -31 58 -31 0 net=121
rlabel metal2 110 -31 110 -31 0 net=290
rlabel metal2 156 -31 156 -31 0 net=401
rlabel metal2 156 -31 156 -31 0 net=401
rlabel metal2 163 -31 163 -31 0 net=439
rlabel metal2 163 -31 163 -31 0 net=439
rlabel metal2 16 -33 16 -33 0 net=173
rlabel metal2 68 -33 68 -33 0 net=198
rlabel metal2 121 -33 121 -33 0 net=367
rlabel metal2 23 -35 23 -35 0 net=23
rlabel metal2 30 -35 30 -35 0 net=186
rlabel metal2 44 -35 44 -35 0 net=181
rlabel metal2 114 -35 114 -35 0 net=345
rlabel metal2 128 -35 128 -35 0 net=397
rlabel metal2 19 -37 19 -37 0 net=155
rlabel metal2 30 -37 30 -37 0 net=37
rlabel metal2 54 -37 54 -37 0 net=76
rlabel metal2 72 -37 72 -37 0 net=252
rlabel metal2 89 -37 89 -37 0 net=255
rlabel metal2 142 -37 142 -37 0 net=353
rlabel metal2 142 -37 142 -37 0 net=353
rlabel metal2 37 -39 37 -39 0 net=221
rlabel metal2 61 -39 61 -39 0 net=270
rlabel metal2 72 -41 72 -41 0 net=357
rlabel metal2 86 -43 86 -43 0 net=339
rlabel metal2 93 -45 93 -45 0 net=301
rlabel metal2 93 -47 93 -47 0 net=167
rlabel metal2 2 -58 2 -58 0 net=257
rlabel metal2 51 -58 51 -58 0 net=122
rlabel metal2 142 -58 142 -58 0 net=355
rlabel metal2 16 -60 16 -60 0 net=174
rlabel metal2 82 -60 82 -60 0 net=302
rlabel metal2 156 -60 156 -60 0 net=403
rlabel metal2 16 -62 16 -62 0 net=125
rlabel metal2 135 -62 135 -62 0 net=169
rlabel metal2 184 -62 184 -62 0 net=381
rlabel metal2 184 -62 184 -62 0 net=381
rlabel metal2 26 -64 26 -64 0 net=303
rlabel metal2 121 -64 121 -64 0 net=347
rlabel metal2 163 -64 163 -64 0 net=441
rlabel metal2 163 -64 163 -64 0 net=441
rlabel metal2 33 -66 33 -66 0 net=22
rlabel metal2 33 -66 33 -66 0 net=22
rlabel metal2 37 -66 37 -66 0 net=101
rlabel metal2 51 -66 51 -66 0 net=311
rlabel metal2 149 -66 149 -66 0 net=369
rlabel metal2 9 -68 9 -68 0 net=45
rlabel metal2 54 -68 54 -68 0 net=229
rlabel metal2 93 -68 93 -68 0 net=256
rlabel metal2 23 -70 23 -70 0 net=157
rlabel metal2 107 -70 107 -70 0 net=341
rlabel metal2 65 -72 65 -72 0 net=78
rlabel metal2 114 -72 114 -72 0 net=398
rlabel metal2 58 -74 58 -74 0 net=223
rlabel metal2 79 -74 79 -74 0 net=183
rlabel metal2 128 -74 128 -74 0 net=359
rlabel metal2 58 -76 58 -76 0 net=133
rlabel metal2 23 -87 23 -87 0 net=147
rlabel metal2 37 -87 37 -87 0 net=103
rlabel metal2 51 -87 51 -87 0 net=135
rlabel metal2 68 -87 68 -87 0 net=184
rlabel metal2 114 -87 114 -87 0 net=370
rlabel metal2 26 -89 26 -89 0 net=224
rlabel metal2 79 -89 79 -89 0 net=342
rlabel metal2 163 -89 163 -89 0 net=443
rlabel metal2 16 -91 16 -91 0 net=127
rlabel metal2 86 -91 86 -91 0 net=187
rlabel metal2 124 -91 124 -91 0 net=404
rlabel metal2 16 -93 16 -93 0 net=159
rlabel metal2 96 -93 96 -93 0 net=149
rlabel metal2 128 -93 128 -93 0 net=356
rlabel metal2 33 -95 33 -95 0 net=281
rlabel metal2 170 -95 170 -95 0 net=361
rlabel metal2 184 -95 184 -95 0 net=383
rlabel metal2 37 -97 37 -97 0 net=143
rlabel metal2 142 -97 142 -97 0 net=313
rlabel metal2 58 -99 58 -99 0 net=11
rlabel metal2 89 -101 89 -101 0 net=170
rlabel metal2 54 -103 54 -103 0 net=245
rlabel metal2 93 -105 93 -105 0 net=348
rlabel metal2 100 -107 100 -107 0 net=305
rlabel metal2 72 -109 72 -109 0 net=231
rlabel metal2 117 -109 117 -109 0 net=405
rlabel metal2 2 -111 2 -111 0 net=259
rlabel metal2 124 -111 124 -111 0 net=325
rlabel metal2 2 -113 2 -113 0 net=409
rlabel metal2 131 -115 131 -115 0 net=371
rlabel metal2 2 -126 2 -126 0 net=160
rlabel metal2 23 -126 23 -126 0 net=148
rlabel metal2 33 -126 33 -126 0 net=42
rlabel metal2 149 -126 149 -126 0 net=283
rlabel metal2 2 -128 2 -128 0 net=233
rlabel metal2 61 -128 61 -128 0 net=232
rlabel metal2 107 -128 107 -128 0 net=151
rlabel metal2 107 -128 107 -128 0 net=151
rlabel metal2 117 -128 117 -128 0 net=329
rlabel metal2 149 -128 149 -128 0 net=449
rlabel metal2 9 -130 9 -130 0 net=85
rlabel metal2 16 -130 16 -130 0 net=253
rlabel metal2 51 -130 51 -130 0 net=137
rlabel metal2 72 -130 72 -130 0 net=260
rlabel metal2 121 -130 121 -130 0 net=444
rlabel metal2 33 -132 33 -132 0 net=123
rlabel metal2 58 -132 58 -132 0 net=111
rlabel metal2 96 -132 96 -132 0 net=406
rlabel metal2 205 -132 205 -132 0 net=411
rlabel metal2 205 -132 205 -132 0 net=411
rlabel metal2 37 -134 37 -134 0 net=145
rlabel metal2 79 -134 79 -134 0 net=128
rlabel metal2 121 -134 121 -134 0 net=425
rlabel metal2 37 -136 37 -136 0 net=105
rlabel metal2 68 -136 68 -136 0 net=261
rlabel metal2 86 -136 86 -136 0 net=189
rlabel metal2 114 -136 114 -136 0 net=427
rlabel metal2 86 -138 86 -138 0 net=247
rlabel metal2 152 -138 152 -138 0 net=55
rlabel metal2 173 -138 173 -138 0 net=419
rlabel metal2 93 -140 93 -140 0 net=90
rlabel metal2 156 -140 156 -140 0 net=307
rlabel metal2 156 -140 156 -140 0 net=307
rlabel metal2 163 -140 163 -140 0 net=315
rlabel metal2 191 -140 191 -140 0 net=385
rlabel metal2 135 -142 135 -142 0 net=453
rlabel metal2 142 -144 142 -144 0 net=327
rlabel metal2 184 -144 184 -144 0 net=373
rlabel metal2 177 -146 177 -146 0 net=363
rlabel metal2 44 -148 44 -148 0 net=445
rlabel metal2 5 -159 5 -159 0 net=95
rlabel metal2 23 -159 23 -159 0 net=124
rlabel metal2 61 -159 61 -159 0 net=426
rlabel metal2 233 -159 233 -159 0 net=451
rlabel metal2 9 -161 9 -161 0 net=254
rlabel metal2 23 -161 23 -161 0 net=161
rlabel metal2 117 -161 117 -161 0 net=364
rlabel metal2 191 -161 191 -161 0 net=375
rlabel metal2 16 -163 16 -163 0 net=113
rlabel metal2 75 -163 75 -163 0 net=175
rlabel metal2 124 -163 124 -163 0 net=209
rlabel metal2 177 -163 177 -163 0 net=447
rlabel metal2 26 -165 26 -165 0 net=454
rlabel metal2 30 -167 30 -167 0 net=433
rlabel metal2 30 -169 30 -169 0 net=139
rlabel metal2 79 -169 79 -169 0 net=263
rlabel metal2 198 -169 198 -169 0 net=387
rlabel metal2 33 -171 33 -171 0 net=248
rlabel metal2 117 -171 117 -171 0 net=275
rlabel metal2 142 -171 142 -171 0 net=328
rlabel metal2 198 -171 198 -171 0 net=285
rlabel metal2 2 -173 2 -173 0 net=235
rlabel metal2 205 -173 205 -173 0 net=413
rlabel metal2 2 -175 2 -175 0 net=428
rlabel metal2 37 -177 37 -177 0 net=107
rlabel metal2 37 -177 37 -177 0 net=107
rlabel metal2 44 -177 44 -177 0 net=193
rlabel metal2 212 -177 212 -177 0 net=421
rlabel metal2 44 -179 44 -179 0 net=117
rlabel metal2 114 -179 114 -179 0 net=201
rlabel metal2 152 -179 152 -179 0 net=407
rlabel metal2 51 -181 51 -181 0 net=271
rlabel metal2 54 -183 54 -183 0 net=215
rlabel metal2 96 -183 96 -183 0 net=333
rlabel metal2 65 -185 65 -185 0 net=60
rlabel metal2 128 -185 128 -185 0 net=331
rlabel metal2 72 -187 72 -187 0 net=146
rlabel metal2 100 -187 100 -187 0 net=191
rlabel metal2 156 -187 156 -187 0 net=309
rlabel metal2 72 -189 72 -189 0 net=129
rlabel metal2 100 -189 100 -189 0 net=153
rlabel metal2 170 -189 170 -189 0 net=317
rlabel metal2 107 -191 107 -191 0 net=35
rlabel metal2 159 -191 159 -191 0 net=239
rlabel metal2 9 -202 9 -202 0 net=236
rlabel metal2 180 -202 180 -202 0 net=194
rlabel metal2 9 -204 9 -204 0 net=195
rlabel metal2 72 -204 72 -204 0 net=177
rlabel metal2 135 -204 135 -204 0 net=277
rlabel metal2 30 -206 30 -206 0 net=140
rlabel metal2 47 -206 47 -206 0 net=434
rlabel metal2 30 -208 30 -208 0 net=109
rlabel metal2 51 -208 51 -208 0 net=48
rlabel metal2 156 -208 156 -208 0 net=414
rlabel metal2 54 -210 54 -210 0 net=408
rlabel metal2 58 -212 58 -212 0 net=74
rlabel metal2 107 -212 107 -212 0 net=435
rlabel metal2 156 -212 156 -212 0 net=241
rlabel metal2 198 -212 198 -212 0 net=287
rlabel metal2 44 -214 44 -214 0 net=118
rlabel metal2 75 -214 75 -214 0 net=100
rlabel metal2 121 -214 121 -214 0 net=203
rlabel metal2 159 -214 159 -214 0 net=452
rlabel metal2 86 -216 86 -216 0 net=154
rlabel metal2 107 -216 107 -216 0 net=211
rlabel metal2 170 -216 170 -216 0 net=319
rlabel metal2 23 -218 23 -218 0 net=163
rlabel metal2 110 -218 110 -218 0 net=332
rlabel metal2 16 -220 16 -220 0 net=115
rlabel metal2 40 -220 40 -220 0 net=293
rlabel metal2 114 -220 114 -220 0 net=310
rlabel metal2 212 -220 212 -220 0 net=377
rlabel metal2 16 -222 16 -222 0 net=141
rlabel metal2 79 -222 79 -222 0 net=217
rlabel metal2 142 -222 142 -222 0 net=265
rlabel metal2 198 -222 198 -222 0 net=335
rlabel metal2 79 -224 79 -224 0 net=131
rlabel metal2 149 -224 149 -224 0 net=273
rlabel metal2 205 -224 205 -224 0 net=291
rlabel metal2 93 -226 93 -226 0 net=192
rlabel metal2 177 -226 177 -226 0 net=429
rlabel metal2 226 -226 226 -226 0 net=423
rlabel metal2 128 -228 128 -228 0 net=448
rlabel metal2 184 -230 184 -230 0 net=389
rlabel metal2 194 -232 194 -232 0 net=225
rlabel metal2 9 -243 9 -243 0 net=196
rlabel metal2 100 -243 100 -243 0 net=165
rlabel metal2 100 -243 100 -243 0 net=165
rlabel metal2 107 -243 107 -243 0 net=213
rlabel metal2 107 -243 107 -243 0 net=213
rlabel metal2 131 -243 131 -243 0 net=274
rlabel metal2 159 -243 159 -243 0 net=292
rlabel metal2 233 -243 233 -243 0 net=227
rlabel metal2 16 -245 16 -245 0 net=142
rlabel metal2 68 -245 68 -245 0 net=132
rlabel metal2 86 -245 86 -245 0 net=295
rlabel metal2 135 -245 135 -245 0 net=436
rlabel metal2 194 -245 194 -245 0 net=424
rlabel metal2 23 -247 23 -247 0 net=116
rlabel metal2 79 -247 79 -247 0 net=267
rlabel metal2 149 -247 149 -247 0 net=279
rlabel metal2 177 -247 177 -247 0 net=288
rlabel metal2 30 -249 30 -249 0 net=110
rlabel metal2 58 -249 58 -249 0 net=119
rlabel metal2 58 -249 58 -249 0 net=119
rlabel metal2 65 -249 65 -249 0 net=30
rlabel metal2 128 -249 128 -249 0 net=297
rlabel metal2 163 -249 163 -249 0 net=391
rlabel metal2 212 -249 212 -249 0 net=379
rlabel metal2 44 -251 44 -251 0 net=178
rlabel metal2 86 -251 86 -251 0 net=219
rlabel metal2 128 -251 128 -251 0 net=321
rlabel metal2 177 -251 177 -251 0 net=337
rlabel metal2 208 -251 208 -251 0 net=15
rlabel metal2 44 -253 44 -253 0 net=417
rlabel metal2 114 -253 114 -253 0 net=205
rlabel metal2 156 -253 156 -253 0 net=243
rlabel metal2 198 -253 198 -253 0 net=431
rlabel metal2 170 -255 170 -255 0 net=199
rlabel metal2 215 -257 215 -257 0 net=415
rlabel metal2 44 -268 44 -268 0 net=418
rlabel metal2 58 -268 58 -268 0 net=120
rlabel metal2 72 -268 72 -268 0 net=249
rlabel metal2 72 -268 72 -268 0 net=249
rlabel metal2 75 -268 75 -268 0 net=268
rlabel metal2 86 -268 86 -268 0 net=220
rlabel metal2 135 -268 135 -268 0 net=298
rlabel metal2 142 -268 142 -268 0 net=280
rlabel metal2 163 -268 163 -268 0 net=392
rlabel metal2 177 -268 177 -268 0 net=338
rlabel metal2 201 -268 201 -268 0 net=200
rlabel metal2 79 -270 79 -270 0 net=296
rlabel metal2 100 -270 100 -270 0 net=166
rlabel metal2 121 -270 121 -270 0 net=244
rlabel metal2 191 -270 191 -270 0 net=432
rlabel metal2 205 -270 205 -270 0 net=228
rlabel metal2 100 -272 100 -272 0 net=214
rlabel metal2 114 -272 114 -272 0 net=207
rlabel metal2 128 -272 128 -272 0 net=323
rlabel metal2 145 -272 145 -272 0 net=36
rlabel metal2 205 -272 205 -272 0 net=416
rlabel metal2 128 -274 128 -274 0 net=27
rlabel metal2 208 -274 208 -274 0 net=380
rlabel metal2 65 -285 65 -285 0 net=250
rlabel metal2 121 -285 121 -285 0 net=208
rlabel metal2 142 -285 142 -285 0 net=324
<< end >>
