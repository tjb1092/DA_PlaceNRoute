magic
tech scmos
timestamp 1555016740 
<< pdiffusion >>
rect 1 -12 7 -6
rect 8 -12 14 -6
rect 15 -12 21 -6
rect 22 -12 28 -6
rect 29 -12 35 -6
rect 36 -12 42 -6
rect 43 -12 49 -6
rect 50 -12 56 -6
rect 57 -12 63 -6
rect 64 -12 67 -6
rect 71 -12 77 -6
rect 78 -12 84 -6
rect 85 -12 91 -6
rect 92 -12 98 -6
rect 99 -12 105 -6
rect 106 -12 109 -6
rect 113 -12 119 -6
rect 120 -12 126 -6
rect 127 -12 130 -6
rect 134 -12 140 -6
rect 141 -12 147 -6
rect 148 -12 151 -6
rect 155 -12 161 -6
rect 162 -12 165 -6
rect 1 -31 7 -25
rect 8 -31 14 -25
rect 15 -31 21 -25
rect 22 -31 28 -25
rect 29 -31 35 -25
rect 36 -31 42 -25
rect 43 -31 49 -25
rect 50 -31 56 -25
rect 71 -31 74 -25
rect 78 -31 84 -25
rect 92 -31 98 -25
rect 99 -31 105 -25
rect 106 -31 112 -25
rect 113 -31 119 -25
rect 120 -31 126 -25
rect 127 -31 130 -25
rect 141 -31 144 -25
rect 148 -31 151 -25
rect 162 -31 165 -25
rect 169 -31 175 -25
rect 176 -31 179 -25
rect 183 -31 189 -25
rect 190 -31 196 -25
rect 197 -31 203 -25
rect 1 -62 7 -56
rect 8 -62 14 -56
rect 15 -62 21 -56
rect 22 -62 28 -56
rect 29 -62 35 -56
rect 36 -62 42 -56
rect 43 -62 49 -56
rect 50 -62 53 -56
rect 57 -62 60 -56
rect 64 -62 67 -56
rect 71 -62 74 -56
rect 78 -62 84 -56
rect 85 -62 91 -56
rect 92 -62 98 -56
rect 99 -62 102 -56
rect 106 -62 112 -56
rect 113 -62 119 -56
rect 120 -62 126 -56
rect 127 -62 133 -56
rect 134 -62 140 -56
rect 141 -62 147 -56
rect 148 -62 154 -56
rect 155 -62 158 -56
rect 162 -62 165 -56
rect 169 -62 172 -56
rect 176 -62 179 -56
rect 183 -62 186 -56
rect 190 -62 196 -56
rect 197 -62 200 -56
rect 204 -62 207 -56
rect 211 -62 214 -56
rect 218 -62 221 -56
rect 225 -62 228 -56
rect 232 -62 235 -56
rect 239 -62 245 -56
rect 246 -62 249 -56
rect 253 -62 256 -56
rect 8 -95 14 -89
rect 15 -95 21 -89
rect 22 -95 28 -89
rect 29 -95 32 -89
rect 36 -95 42 -89
rect 43 -95 46 -89
rect 50 -95 53 -89
rect 57 -95 60 -89
rect 64 -95 67 -89
rect 71 -95 74 -89
rect 78 -95 84 -89
rect 85 -95 88 -89
rect 92 -95 98 -89
rect 99 -95 105 -89
rect 106 -95 112 -89
rect 113 -95 119 -89
rect 120 -95 123 -89
rect 127 -95 133 -89
rect 134 -95 140 -89
rect 141 -95 147 -89
rect 148 -95 154 -89
rect 155 -95 161 -89
rect 162 -95 168 -89
rect 169 -95 175 -89
rect 176 -95 179 -89
rect 183 -95 189 -89
rect 190 -95 193 -89
rect 197 -95 203 -89
rect 204 -95 207 -89
rect 211 -95 214 -89
rect 218 -95 221 -89
rect 225 -95 228 -89
rect 232 -95 235 -89
rect 239 -95 242 -89
rect 246 -95 249 -89
rect 253 -95 256 -89
rect 260 -95 263 -89
rect 267 -95 270 -89
rect 274 -95 277 -89
rect 281 -95 284 -89
rect 288 -95 291 -89
rect 295 -95 298 -89
rect 302 -95 308 -89
rect 330 -95 333 -89
rect 1 -150 7 -144
rect 8 -150 14 -144
rect 15 -150 21 -144
rect 22 -150 28 -144
rect 29 -150 35 -144
rect 36 -150 42 -144
rect 43 -150 46 -144
rect 50 -150 53 -144
rect 57 -150 63 -144
rect 64 -150 67 -144
rect 71 -150 74 -144
rect 78 -150 84 -144
rect 85 -150 91 -144
rect 92 -150 95 -144
rect 99 -150 102 -144
rect 106 -150 109 -144
rect 113 -150 119 -144
rect 120 -150 126 -144
rect 127 -150 133 -144
rect 134 -150 140 -144
rect 141 -150 144 -144
rect 148 -150 154 -144
rect 155 -150 158 -144
rect 162 -150 168 -144
rect 169 -150 172 -144
rect 176 -150 179 -144
rect 183 -150 186 -144
rect 190 -150 196 -144
rect 197 -150 203 -144
rect 204 -150 210 -144
rect 211 -150 214 -144
rect 218 -150 221 -144
rect 225 -150 228 -144
rect 232 -150 235 -144
rect 239 -150 242 -144
rect 246 -150 249 -144
rect 253 -150 256 -144
rect 260 -150 263 -144
rect 267 -150 273 -144
rect 274 -150 277 -144
rect 281 -150 284 -144
rect 288 -150 291 -144
rect 295 -150 298 -144
rect 302 -150 305 -144
rect 309 -150 312 -144
rect 316 -150 319 -144
rect 323 -150 326 -144
rect 330 -150 333 -144
rect 337 -150 340 -144
rect 344 -150 347 -144
rect 351 -150 354 -144
rect 358 -150 361 -144
rect 365 -150 368 -144
rect 372 -150 375 -144
rect 1 -201 7 -195
rect 8 -201 11 -195
rect 15 -201 18 -195
rect 22 -201 28 -195
rect 29 -201 32 -195
rect 36 -201 39 -195
rect 43 -201 49 -195
rect 50 -201 53 -195
rect 57 -201 63 -195
rect 64 -201 67 -195
rect 71 -201 77 -195
rect 78 -201 84 -195
rect 85 -201 88 -195
rect 92 -201 98 -195
rect 99 -201 105 -195
rect 106 -201 109 -195
rect 113 -201 116 -195
rect 120 -201 123 -195
rect 127 -201 133 -195
rect 134 -201 140 -195
rect 141 -201 144 -195
rect 148 -201 154 -195
rect 155 -201 158 -195
rect 162 -201 168 -195
rect 169 -201 175 -195
rect 176 -201 179 -195
rect 183 -201 189 -195
rect 190 -201 193 -195
rect 197 -201 203 -195
rect 204 -201 210 -195
rect 211 -201 214 -195
rect 218 -201 224 -195
rect 225 -201 228 -195
rect 232 -201 235 -195
rect 239 -201 242 -195
rect 246 -201 249 -195
rect 253 -201 256 -195
rect 260 -201 263 -195
rect 267 -201 270 -195
rect 274 -201 277 -195
rect 281 -201 284 -195
rect 288 -201 291 -195
rect 295 -201 298 -195
rect 302 -201 305 -195
rect 309 -201 312 -195
rect 316 -201 322 -195
rect 323 -201 326 -195
rect 330 -201 333 -195
rect 337 -201 340 -195
rect 344 -201 347 -195
rect 351 -201 354 -195
rect 358 -201 361 -195
rect 365 -201 368 -195
rect 372 -201 375 -195
rect 379 -201 382 -195
rect 386 -201 389 -195
rect 393 -201 396 -195
rect 400 -201 403 -195
rect 407 -201 413 -195
rect 414 -201 417 -195
rect 1 -260 7 -254
rect 8 -260 14 -254
rect 15 -260 18 -254
rect 22 -260 25 -254
rect 29 -260 35 -254
rect 36 -260 39 -254
rect 43 -260 46 -254
rect 50 -260 56 -254
rect 57 -260 60 -254
rect 64 -260 67 -254
rect 71 -260 77 -254
rect 78 -260 84 -254
rect 85 -260 88 -254
rect 92 -260 98 -254
rect 99 -260 105 -254
rect 106 -260 112 -254
rect 113 -260 119 -254
rect 120 -260 126 -254
rect 127 -260 130 -254
rect 134 -260 140 -254
rect 141 -260 144 -254
rect 148 -260 151 -254
rect 155 -260 158 -254
rect 162 -260 165 -254
rect 169 -260 172 -254
rect 176 -260 182 -254
rect 183 -260 189 -254
rect 190 -260 193 -254
rect 197 -260 203 -254
rect 204 -260 207 -254
rect 211 -260 214 -254
rect 218 -260 224 -254
rect 225 -260 228 -254
rect 232 -260 235 -254
rect 239 -260 245 -254
rect 246 -260 249 -254
rect 253 -260 259 -254
rect 260 -260 263 -254
rect 267 -260 270 -254
rect 274 -260 277 -254
rect 281 -260 287 -254
rect 288 -260 291 -254
rect 295 -260 298 -254
rect 302 -260 305 -254
rect 309 -260 312 -254
rect 316 -260 319 -254
rect 323 -260 326 -254
rect 330 -260 333 -254
rect 337 -260 340 -254
rect 344 -260 347 -254
rect 351 -260 354 -254
rect 358 -260 361 -254
rect 365 -260 368 -254
rect 372 -260 375 -254
rect 379 -260 382 -254
rect 386 -260 389 -254
rect 393 -260 396 -254
rect 400 -260 403 -254
rect 407 -260 410 -254
rect 414 -260 417 -254
rect 1 -309 7 -303
rect 8 -309 14 -303
rect 15 -309 18 -303
rect 22 -309 25 -303
rect 29 -309 32 -303
rect 36 -309 39 -303
rect 43 -309 46 -303
rect 50 -309 53 -303
rect 57 -309 63 -303
rect 64 -309 67 -303
rect 71 -309 77 -303
rect 78 -309 81 -303
rect 85 -309 88 -303
rect 92 -309 98 -303
rect 99 -309 105 -303
rect 106 -309 112 -303
rect 113 -309 119 -303
rect 120 -309 126 -303
rect 127 -309 130 -303
rect 134 -309 137 -303
rect 141 -309 144 -303
rect 148 -309 151 -303
rect 155 -309 158 -303
rect 162 -309 168 -303
rect 169 -309 175 -303
rect 176 -309 179 -303
rect 183 -309 186 -303
rect 190 -309 193 -303
rect 197 -309 203 -303
rect 204 -309 210 -303
rect 211 -309 217 -303
rect 218 -309 221 -303
rect 225 -309 228 -303
rect 232 -309 235 -303
rect 239 -309 245 -303
rect 246 -309 252 -303
rect 253 -309 256 -303
rect 260 -309 266 -303
rect 267 -309 270 -303
rect 274 -309 277 -303
rect 281 -309 284 -303
rect 288 -309 291 -303
rect 295 -309 298 -303
rect 302 -309 305 -303
rect 309 -309 312 -303
rect 316 -309 319 -303
rect 323 -309 326 -303
rect 330 -309 333 -303
rect 337 -309 340 -303
rect 344 -309 347 -303
rect 351 -309 354 -303
rect 358 -309 361 -303
rect 365 -309 368 -303
rect 372 -309 375 -303
rect 379 -309 382 -303
rect 386 -309 389 -303
rect 393 -309 396 -303
rect 400 -309 403 -303
rect 407 -309 410 -303
rect 414 -309 417 -303
rect 421 -309 427 -303
rect 428 -309 434 -303
rect 435 -309 438 -303
rect 1 -370 4 -364
rect 8 -370 14 -364
rect 15 -370 18 -364
rect 22 -370 28 -364
rect 29 -370 35 -364
rect 36 -370 42 -364
rect 43 -370 49 -364
rect 50 -370 56 -364
rect 57 -370 60 -364
rect 64 -370 70 -364
rect 71 -370 77 -364
rect 78 -370 84 -364
rect 85 -370 91 -364
rect 92 -370 95 -364
rect 99 -370 102 -364
rect 106 -370 112 -364
rect 113 -370 119 -364
rect 120 -370 123 -364
rect 127 -370 130 -364
rect 134 -370 137 -364
rect 141 -370 144 -364
rect 148 -370 151 -364
rect 155 -370 161 -364
rect 162 -370 165 -364
rect 169 -370 175 -364
rect 176 -370 179 -364
rect 183 -370 189 -364
rect 190 -370 193 -364
rect 197 -370 200 -364
rect 204 -370 207 -364
rect 211 -370 214 -364
rect 218 -370 224 -364
rect 225 -370 228 -364
rect 232 -370 238 -364
rect 239 -370 242 -364
rect 246 -370 249 -364
rect 253 -370 259 -364
rect 260 -370 263 -364
rect 267 -370 273 -364
rect 274 -370 277 -364
rect 281 -370 284 -364
rect 288 -370 291 -364
rect 295 -370 298 -364
rect 302 -370 305 -364
rect 309 -370 312 -364
rect 316 -370 319 -364
rect 323 -370 326 -364
rect 330 -370 333 -364
rect 337 -370 340 -364
rect 344 -370 347 -364
rect 351 -370 354 -364
rect 358 -370 361 -364
rect 365 -370 368 -364
rect 372 -370 375 -364
rect 379 -370 382 -364
rect 386 -370 389 -364
rect 393 -370 396 -364
rect 400 -370 403 -364
rect 407 -370 410 -364
rect 414 -370 417 -364
rect 421 -370 424 -364
rect 428 -370 431 -364
rect 435 -370 438 -364
rect 8 -419 11 -413
rect 15 -419 18 -413
rect 22 -419 28 -413
rect 29 -419 32 -413
rect 36 -419 39 -413
rect 43 -419 49 -413
rect 50 -419 56 -413
rect 57 -419 63 -413
rect 64 -419 67 -413
rect 71 -419 74 -413
rect 78 -419 81 -413
rect 85 -419 88 -413
rect 92 -419 95 -413
rect 99 -419 105 -413
rect 106 -419 112 -413
rect 113 -419 119 -413
rect 120 -419 123 -413
rect 127 -419 133 -413
rect 134 -419 137 -413
rect 141 -419 144 -413
rect 148 -419 151 -413
rect 155 -419 158 -413
rect 162 -419 168 -413
rect 169 -419 172 -413
rect 176 -419 179 -413
rect 183 -419 186 -413
rect 190 -419 193 -413
rect 197 -419 203 -413
rect 204 -419 207 -413
rect 211 -419 214 -413
rect 218 -419 221 -413
rect 225 -419 231 -413
rect 232 -419 235 -413
rect 239 -419 245 -413
rect 246 -419 252 -413
rect 253 -419 256 -413
rect 260 -419 266 -413
rect 267 -419 273 -413
rect 274 -419 277 -413
rect 281 -419 284 -413
rect 288 -419 291 -413
rect 295 -419 298 -413
rect 302 -419 305 -413
rect 309 -419 312 -413
rect 316 -419 319 -413
rect 323 -419 329 -413
rect 330 -419 336 -413
rect 337 -419 340 -413
rect 344 -419 347 -413
rect 351 -419 354 -413
rect 358 -419 361 -413
rect 365 -419 368 -413
rect 372 -419 375 -413
rect 379 -419 382 -413
rect 386 -419 389 -413
rect 393 -419 396 -413
rect 400 -419 403 -413
rect 407 -419 410 -413
rect 414 -419 417 -413
rect 421 -419 424 -413
rect 428 -419 434 -413
rect 435 -419 438 -413
rect 442 -419 448 -413
rect 15 -474 18 -468
rect 22 -474 28 -468
rect 29 -474 35 -468
rect 36 -474 39 -468
rect 50 -474 53 -468
rect 57 -474 60 -468
rect 64 -474 67 -468
rect 71 -474 77 -468
rect 78 -474 81 -468
rect 85 -474 88 -468
rect 92 -474 95 -468
rect 99 -474 102 -468
rect 106 -474 112 -468
rect 113 -474 116 -468
rect 120 -474 123 -468
rect 127 -474 133 -468
rect 134 -474 137 -468
rect 141 -474 144 -468
rect 148 -474 151 -468
rect 155 -474 158 -468
rect 162 -474 165 -468
rect 169 -474 172 -468
rect 176 -474 182 -468
rect 183 -474 186 -468
rect 190 -474 196 -468
rect 197 -474 203 -468
rect 204 -474 207 -468
rect 211 -474 217 -468
rect 218 -474 224 -468
rect 225 -474 231 -468
rect 232 -474 238 -468
rect 239 -474 245 -468
rect 246 -474 252 -468
rect 253 -474 259 -468
rect 260 -474 266 -468
rect 267 -474 270 -468
rect 274 -474 277 -468
rect 281 -474 287 -468
rect 288 -474 291 -468
rect 295 -474 298 -468
rect 302 -474 305 -468
rect 309 -474 312 -468
rect 316 -474 319 -468
rect 323 -474 326 -468
rect 330 -474 333 -468
rect 337 -474 340 -468
rect 344 -474 347 -468
rect 351 -474 354 -468
rect 358 -474 361 -468
rect 365 -474 368 -468
rect 372 -474 375 -468
rect 379 -474 382 -468
rect 386 -474 389 -468
rect 393 -474 396 -468
rect 414 -474 417 -468
rect 421 -474 424 -468
rect 428 -474 434 -468
rect 435 -474 438 -468
rect 442 -474 448 -468
rect 449 -474 452 -468
rect 456 -474 459 -468
rect 463 -474 466 -468
rect 8 -515 11 -509
rect 15 -515 18 -509
rect 22 -515 28 -509
rect 29 -515 35 -509
rect 36 -515 42 -509
rect 43 -515 46 -509
rect 50 -515 53 -509
rect 57 -515 60 -509
rect 64 -515 67 -509
rect 71 -515 77 -509
rect 78 -515 84 -509
rect 85 -515 88 -509
rect 92 -515 95 -509
rect 99 -515 105 -509
rect 106 -515 109 -509
rect 113 -515 116 -509
rect 120 -515 126 -509
rect 127 -515 130 -509
rect 134 -515 140 -509
rect 141 -515 144 -509
rect 148 -515 151 -509
rect 155 -515 158 -509
rect 162 -515 165 -509
rect 169 -515 175 -509
rect 176 -515 179 -509
rect 183 -515 186 -509
rect 190 -515 193 -509
rect 197 -515 200 -509
rect 204 -515 210 -509
rect 211 -515 217 -509
rect 218 -515 221 -509
rect 225 -515 228 -509
rect 232 -515 235 -509
rect 239 -515 245 -509
rect 246 -515 249 -509
rect 253 -515 256 -509
rect 260 -515 263 -509
rect 267 -515 270 -509
rect 274 -515 280 -509
rect 281 -515 287 -509
rect 288 -515 291 -509
rect 295 -515 298 -509
rect 302 -515 308 -509
rect 309 -515 312 -509
rect 316 -515 319 -509
rect 323 -515 326 -509
rect 330 -515 333 -509
rect 337 -515 340 -509
rect 344 -515 347 -509
rect 351 -515 354 -509
rect 358 -515 361 -509
rect 365 -515 371 -509
rect 372 -515 375 -509
rect 379 -515 382 -509
rect 386 -515 389 -509
rect 400 -515 403 -509
rect 407 -515 410 -509
rect 414 -515 420 -509
rect 428 -515 434 -509
rect 435 -515 438 -509
rect 442 -515 448 -509
rect 449 -515 452 -509
rect 456 -515 459 -509
rect 463 -515 466 -509
rect 8 -568 11 -562
rect 15 -568 21 -562
rect 22 -568 28 -562
rect 29 -568 32 -562
rect 36 -568 39 -562
rect 43 -568 46 -562
rect 50 -568 53 -562
rect 57 -568 60 -562
rect 64 -568 70 -562
rect 71 -568 74 -562
rect 78 -568 84 -562
rect 85 -568 88 -562
rect 92 -568 98 -562
rect 99 -568 105 -562
rect 106 -568 109 -562
rect 113 -568 119 -562
rect 120 -568 126 -562
rect 127 -568 130 -562
rect 134 -568 137 -562
rect 141 -568 144 -562
rect 148 -568 151 -562
rect 155 -568 158 -562
rect 162 -568 168 -562
rect 169 -568 175 -562
rect 176 -568 182 -562
rect 183 -568 189 -562
rect 190 -568 193 -562
rect 197 -568 200 -562
rect 204 -568 210 -562
rect 211 -568 214 -562
rect 218 -568 221 -562
rect 225 -568 228 -562
rect 232 -568 238 -562
rect 239 -568 245 -562
rect 246 -568 249 -562
rect 253 -568 256 -562
rect 260 -568 263 -562
rect 267 -568 270 -562
rect 274 -568 277 -562
rect 281 -568 287 -562
rect 288 -568 291 -562
rect 295 -568 298 -562
rect 302 -568 308 -562
rect 309 -568 312 -562
rect 316 -568 319 -562
rect 323 -568 326 -562
rect 330 -568 333 -562
rect 337 -568 343 -562
rect 344 -568 347 -562
rect 351 -568 354 -562
rect 358 -568 361 -562
rect 365 -568 368 -562
rect 372 -568 375 -562
rect 379 -568 382 -562
rect 386 -568 389 -562
rect 393 -568 396 -562
rect 400 -568 403 -562
rect 407 -568 410 -562
rect 414 -568 417 -562
rect 421 -568 424 -562
rect 428 -568 431 -562
rect 435 -568 438 -562
rect 442 -568 445 -562
rect 456 -568 462 -562
rect 463 -568 466 -562
rect 8 -621 11 -615
rect 15 -621 18 -615
rect 22 -621 25 -615
rect 29 -621 35 -615
rect 36 -621 42 -615
rect 43 -621 46 -615
rect 50 -621 53 -615
rect 57 -621 60 -615
rect 64 -621 67 -615
rect 71 -621 74 -615
rect 78 -621 81 -615
rect 85 -621 91 -615
rect 92 -621 95 -615
rect 99 -621 105 -615
rect 106 -621 109 -615
rect 113 -621 119 -615
rect 120 -621 123 -615
rect 127 -621 133 -615
rect 134 -621 140 -615
rect 141 -621 144 -615
rect 148 -621 151 -615
rect 155 -621 158 -615
rect 162 -621 165 -615
rect 169 -621 175 -615
rect 176 -621 179 -615
rect 183 -621 186 -615
rect 190 -621 196 -615
rect 197 -621 200 -615
rect 204 -621 210 -615
rect 211 -621 217 -615
rect 218 -621 221 -615
rect 225 -621 228 -615
rect 232 -621 235 -615
rect 239 -621 242 -615
rect 246 -621 252 -615
rect 253 -621 259 -615
rect 260 -621 266 -615
rect 267 -621 270 -615
rect 274 -621 277 -615
rect 281 -621 284 -615
rect 288 -621 291 -615
rect 295 -621 301 -615
rect 302 -621 305 -615
rect 309 -621 312 -615
rect 316 -621 319 -615
rect 323 -621 326 -615
rect 330 -621 336 -615
rect 337 -621 340 -615
rect 344 -621 347 -615
rect 351 -621 354 -615
rect 358 -621 361 -615
rect 365 -621 368 -615
rect 372 -621 375 -615
rect 379 -621 382 -615
rect 386 -621 389 -615
rect 393 -621 396 -615
rect 400 -621 403 -615
rect 407 -621 410 -615
rect 414 -621 417 -615
rect 421 -621 424 -615
rect 428 -621 431 -615
rect 435 -621 438 -615
rect 442 -621 448 -615
rect 449 -621 455 -615
rect 456 -621 459 -615
rect 463 -621 469 -615
rect 470 -621 473 -615
rect 1 -672 4 -666
rect 8 -672 11 -666
rect 15 -672 18 -666
rect 22 -672 25 -666
rect 29 -672 32 -666
rect 36 -672 39 -666
rect 43 -672 49 -666
rect 50 -672 56 -666
rect 57 -672 60 -666
rect 64 -672 67 -666
rect 71 -672 77 -666
rect 78 -672 81 -666
rect 85 -672 88 -666
rect 92 -672 95 -666
rect 99 -672 105 -666
rect 106 -672 109 -666
rect 113 -672 119 -666
rect 120 -672 123 -666
rect 127 -672 133 -666
rect 134 -672 137 -666
rect 141 -672 144 -666
rect 148 -672 151 -666
rect 155 -672 158 -666
rect 162 -672 165 -666
rect 169 -672 172 -666
rect 176 -672 182 -666
rect 183 -672 189 -666
rect 190 -672 196 -666
rect 197 -672 200 -666
rect 204 -672 210 -666
rect 211 -672 217 -666
rect 218 -672 224 -666
rect 225 -672 228 -666
rect 232 -672 235 -666
rect 239 -672 245 -666
rect 246 -672 252 -666
rect 253 -672 256 -666
rect 260 -672 263 -666
rect 267 -672 273 -666
rect 274 -672 277 -666
rect 281 -672 284 -666
rect 288 -672 291 -666
rect 295 -672 301 -666
rect 302 -672 305 -666
rect 309 -672 312 -666
rect 316 -672 319 -666
rect 323 -672 326 -666
rect 330 -672 336 -666
rect 337 -672 340 -666
rect 344 -672 347 -666
rect 351 -672 354 -666
rect 358 -672 361 -666
rect 365 -672 368 -666
rect 372 -672 375 -666
rect 379 -672 382 -666
rect 386 -672 389 -666
rect 393 -672 396 -666
rect 400 -672 403 -666
rect 407 -672 410 -666
rect 414 -672 417 -666
rect 421 -672 424 -666
rect 428 -672 431 -666
rect 435 -672 438 -666
rect 442 -672 445 -666
rect 449 -672 452 -666
rect 456 -672 462 -666
rect 463 -672 469 -666
rect 470 -672 473 -666
rect 1 -723 4 -717
rect 8 -723 11 -717
rect 15 -723 18 -717
rect 22 -723 25 -717
rect 29 -723 32 -717
rect 36 -723 42 -717
rect 43 -723 46 -717
rect 50 -723 56 -717
rect 57 -723 60 -717
rect 64 -723 67 -717
rect 71 -723 77 -717
rect 78 -723 84 -717
rect 85 -723 88 -717
rect 92 -723 95 -717
rect 99 -723 102 -717
rect 106 -723 109 -717
rect 113 -723 116 -717
rect 120 -723 126 -717
rect 127 -723 133 -717
rect 134 -723 137 -717
rect 141 -723 144 -717
rect 148 -723 151 -717
rect 155 -723 158 -717
rect 162 -723 165 -717
rect 169 -723 175 -717
rect 176 -723 182 -717
rect 183 -723 189 -717
rect 190 -723 193 -717
rect 197 -723 203 -717
rect 204 -723 210 -717
rect 211 -723 214 -717
rect 218 -723 221 -717
rect 225 -723 231 -717
rect 232 -723 235 -717
rect 239 -723 245 -717
rect 246 -723 252 -717
rect 253 -723 256 -717
rect 260 -723 263 -717
rect 267 -723 270 -717
rect 274 -723 280 -717
rect 281 -723 284 -717
rect 288 -723 291 -717
rect 295 -723 301 -717
rect 309 -723 312 -717
rect 316 -723 319 -717
rect 323 -723 326 -717
rect 330 -723 333 -717
rect 337 -723 343 -717
rect 344 -723 347 -717
rect 351 -723 354 -717
rect 358 -723 361 -717
rect 365 -723 368 -717
rect 372 -723 378 -717
rect 379 -723 382 -717
rect 386 -723 389 -717
rect 393 -723 396 -717
rect 400 -723 403 -717
rect 407 -723 413 -717
rect 428 -723 431 -717
rect 15 -776 21 -770
rect 22 -776 25 -770
rect 29 -776 35 -770
rect 36 -776 42 -770
rect 43 -776 49 -770
rect 50 -776 53 -770
rect 57 -776 60 -770
rect 64 -776 67 -770
rect 71 -776 77 -770
rect 78 -776 84 -770
rect 85 -776 88 -770
rect 92 -776 98 -770
rect 99 -776 105 -770
rect 106 -776 112 -770
rect 113 -776 119 -770
rect 120 -776 126 -770
rect 127 -776 130 -770
rect 134 -776 137 -770
rect 141 -776 144 -770
rect 148 -776 151 -770
rect 155 -776 158 -770
rect 162 -776 165 -770
rect 169 -776 172 -770
rect 176 -776 182 -770
rect 183 -776 186 -770
rect 190 -776 193 -770
rect 197 -776 203 -770
rect 204 -776 210 -770
rect 211 -776 217 -770
rect 218 -776 221 -770
rect 225 -776 228 -770
rect 232 -776 238 -770
rect 239 -776 242 -770
rect 246 -776 249 -770
rect 253 -776 256 -770
rect 260 -776 263 -770
rect 267 -776 270 -770
rect 274 -776 280 -770
rect 281 -776 284 -770
rect 288 -776 291 -770
rect 302 -776 305 -770
rect 309 -776 312 -770
rect 323 -776 326 -770
rect 330 -776 336 -770
rect 337 -776 340 -770
rect 344 -776 347 -770
rect 407 -776 413 -770
rect 8 -821 11 -815
rect 15 -821 21 -815
rect 22 -821 25 -815
rect 29 -821 35 -815
rect 36 -821 39 -815
rect 43 -821 49 -815
rect 50 -821 56 -815
rect 57 -821 63 -815
rect 64 -821 70 -815
rect 71 -821 74 -815
rect 78 -821 84 -815
rect 85 -821 91 -815
rect 92 -821 98 -815
rect 99 -821 102 -815
rect 106 -821 112 -815
rect 113 -821 119 -815
rect 120 -821 126 -815
rect 127 -821 133 -815
rect 134 -821 137 -815
rect 141 -821 147 -815
rect 148 -821 154 -815
rect 155 -821 158 -815
rect 162 -821 165 -815
rect 169 -821 172 -815
rect 176 -821 182 -815
rect 183 -821 186 -815
rect 190 -821 193 -815
rect 197 -821 200 -815
rect 204 -821 207 -815
rect 211 -821 214 -815
rect 218 -821 224 -815
rect 225 -821 228 -815
rect 232 -821 235 -815
rect 239 -821 245 -815
rect 246 -821 249 -815
rect 253 -821 256 -815
rect 260 -821 263 -815
rect 267 -821 270 -815
rect 281 -821 284 -815
rect 288 -821 291 -815
rect 302 -821 305 -815
rect 309 -821 312 -815
rect 316 -821 319 -815
rect 323 -821 326 -815
rect 344 -821 350 -815
rect 15 -854 21 -848
rect 22 -854 25 -848
rect 29 -854 35 -848
rect 36 -854 39 -848
rect 43 -854 49 -848
rect 50 -854 56 -848
rect 57 -854 60 -848
rect 64 -854 70 -848
rect 71 -854 74 -848
rect 78 -854 84 -848
rect 85 -854 88 -848
rect 92 -854 95 -848
rect 99 -854 105 -848
rect 106 -854 112 -848
rect 113 -854 119 -848
rect 120 -854 126 -848
rect 127 -854 133 -848
rect 134 -854 140 -848
rect 141 -854 147 -848
rect 148 -854 151 -848
rect 155 -854 158 -848
rect 162 -854 165 -848
rect 169 -854 172 -848
rect 183 -854 189 -848
rect 190 -854 193 -848
rect 211 -854 217 -848
rect 225 -854 231 -848
rect 267 -854 270 -848
rect 281 -854 287 -848
rect 288 -854 294 -848
rect 323 -854 329 -848
<< polysilicon >>
rect 12 -7 13 -5
rect 26 -7 27 -5
rect 37 -7 38 -5
rect 51 -7 52 -5
rect 58 -7 59 -5
rect 65 -7 66 -5
rect 65 -13 66 -11
rect 72 -7 73 -5
rect 72 -13 73 -11
rect 89 -7 90 -5
rect 93 -7 94 -5
rect 96 -13 97 -11
rect 100 -13 101 -11
rect 107 -7 108 -5
rect 107 -13 108 -11
rect 114 -13 115 -11
rect 121 -7 122 -5
rect 128 -7 129 -5
rect 128 -13 129 -11
rect 135 -7 136 -5
rect 138 -7 139 -5
rect 145 -13 146 -11
rect 149 -7 150 -5
rect 149 -13 150 -11
rect 156 -13 157 -11
rect 159 -13 160 -11
rect 163 -7 164 -5
rect 163 -13 164 -11
rect 5 -32 6 -30
rect 30 -32 31 -30
rect 37 -32 38 -30
rect 72 -26 73 -24
rect 72 -32 73 -30
rect 79 -26 80 -24
rect 93 -32 94 -30
rect 100 -26 101 -24
rect 107 -26 108 -24
rect 114 -26 115 -24
rect 117 -32 118 -30
rect 124 -32 125 -30
rect 128 -26 129 -24
rect 128 -32 129 -30
rect 142 -26 143 -24
rect 142 -32 143 -30
rect 149 -26 150 -24
rect 149 -32 150 -30
rect 163 -26 164 -24
rect 163 -32 164 -30
rect 173 -26 174 -24
rect 177 -26 178 -24
rect 177 -32 178 -30
rect 187 -26 188 -24
rect 191 -26 192 -24
rect 191 -32 192 -30
rect 201 -26 202 -24
rect 198 -32 199 -30
rect 5 -57 6 -55
rect 16 -57 17 -55
rect 30 -57 31 -55
rect 30 -63 31 -61
rect 40 -63 41 -61
rect 47 -57 48 -55
rect 51 -57 52 -55
rect 51 -63 52 -61
rect 58 -57 59 -55
rect 58 -63 59 -61
rect 65 -57 66 -55
rect 65 -63 66 -61
rect 72 -57 73 -55
rect 72 -63 73 -61
rect 79 -57 80 -55
rect 82 -63 83 -61
rect 86 -57 87 -55
rect 89 -63 90 -61
rect 93 -57 94 -55
rect 96 -57 97 -55
rect 100 -57 101 -55
rect 100 -63 101 -61
rect 107 -63 108 -61
rect 110 -63 111 -61
rect 114 -63 115 -61
rect 121 -57 122 -55
rect 124 -57 125 -55
rect 128 -57 129 -55
rect 128 -63 129 -61
rect 131 -63 132 -61
rect 135 -63 136 -61
rect 145 -57 146 -55
rect 149 -57 150 -55
rect 152 -57 153 -55
rect 156 -57 157 -55
rect 156 -63 157 -61
rect 163 -57 164 -55
rect 163 -63 164 -61
rect 170 -57 171 -55
rect 170 -63 171 -61
rect 177 -57 178 -55
rect 177 -63 178 -61
rect 184 -57 185 -55
rect 184 -63 185 -61
rect 191 -63 192 -61
rect 198 -57 199 -55
rect 198 -63 199 -61
rect 205 -57 206 -55
rect 205 -63 206 -61
rect 212 -57 213 -55
rect 212 -63 213 -61
rect 219 -57 220 -55
rect 219 -63 220 -61
rect 226 -57 227 -55
rect 226 -63 227 -61
rect 233 -57 234 -55
rect 233 -63 234 -61
rect 243 -63 244 -61
rect 247 -57 248 -55
rect 247 -63 248 -61
rect 254 -57 255 -55
rect 254 -63 255 -61
rect 9 -96 10 -94
rect 19 -90 20 -88
rect 23 -96 24 -94
rect 30 -90 31 -88
rect 30 -96 31 -94
rect 40 -90 41 -88
rect 44 -90 45 -88
rect 44 -96 45 -94
rect 51 -90 52 -88
rect 51 -96 52 -94
rect 58 -90 59 -88
rect 58 -96 59 -94
rect 65 -90 66 -88
rect 65 -96 66 -94
rect 72 -90 73 -88
rect 72 -96 73 -94
rect 79 -90 80 -88
rect 86 -90 87 -88
rect 86 -96 87 -94
rect 96 -90 97 -88
rect 96 -96 97 -94
rect 100 -90 101 -88
rect 110 -90 111 -88
rect 117 -96 118 -94
rect 121 -90 122 -88
rect 121 -96 122 -94
rect 131 -90 132 -88
rect 128 -96 129 -94
rect 131 -96 132 -94
rect 138 -90 139 -88
rect 135 -96 136 -94
rect 138 -96 139 -94
rect 142 -90 143 -88
rect 145 -96 146 -94
rect 149 -90 150 -88
rect 149 -96 150 -94
rect 159 -90 160 -88
rect 156 -96 157 -94
rect 163 -96 164 -94
rect 166 -96 167 -94
rect 170 -90 171 -88
rect 173 -96 174 -94
rect 177 -90 178 -88
rect 177 -96 178 -94
rect 184 -90 185 -88
rect 191 -90 192 -88
rect 191 -96 192 -94
rect 198 -96 199 -94
rect 201 -96 202 -94
rect 205 -90 206 -88
rect 205 -96 206 -94
rect 212 -90 213 -88
rect 212 -96 213 -94
rect 219 -90 220 -88
rect 219 -96 220 -94
rect 226 -90 227 -88
rect 226 -96 227 -94
rect 233 -90 234 -88
rect 233 -96 234 -94
rect 240 -90 241 -88
rect 240 -96 241 -94
rect 247 -90 248 -88
rect 247 -96 248 -94
rect 254 -90 255 -88
rect 254 -96 255 -94
rect 261 -90 262 -88
rect 261 -96 262 -94
rect 268 -90 269 -88
rect 268 -96 269 -94
rect 275 -90 276 -88
rect 275 -96 276 -94
rect 282 -90 283 -88
rect 282 -96 283 -94
rect 289 -90 290 -88
rect 289 -96 290 -94
rect 296 -90 297 -88
rect 296 -96 297 -94
rect 303 -96 304 -94
rect 331 -90 332 -88
rect 331 -96 332 -94
rect 16 -151 17 -149
rect 19 -151 20 -149
rect 26 -145 27 -143
rect 23 -151 24 -149
rect 30 -145 31 -143
rect 30 -151 31 -149
rect 37 -145 38 -143
rect 37 -151 38 -149
rect 44 -145 45 -143
rect 44 -151 45 -149
rect 51 -145 52 -143
rect 51 -151 52 -149
rect 58 -145 59 -143
rect 58 -151 59 -149
rect 61 -151 62 -149
rect 65 -145 66 -143
rect 65 -151 66 -149
rect 72 -145 73 -143
rect 72 -151 73 -149
rect 79 -151 80 -149
rect 82 -151 83 -149
rect 86 -145 87 -143
rect 86 -151 87 -149
rect 89 -151 90 -149
rect 93 -145 94 -143
rect 93 -151 94 -149
rect 100 -145 101 -143
rect 100 -151 101 -149
rect 107 -145 108 -143
rect 107 -151 108 -149
rect 114 -151 115 -149
rect 121 -145 122 -143
rect 124 -145 125 -143
rect 121 -151 122 -149
rect 128 -145 129 -143
rect 128 -151 129 -149
rect 138 -145 139 -143
rect 135 -151 136 -149
rect 142 -145 143 -143
rect 142 -151 143 -149
rect 149 -145 150 -143
rect 152 -145 153 -143
rect 149 -151 150 -149
rect 152 -151 153 -149
rect 156 -145 157 -143
rect 156 -151 157 -149
rect 163 -145 164 -143
rect 166 -145 167 -143
rect 163 -151 164 -149
rect 170 -145 171 -143
rect 170 -151 171 -149
rect 177 -145 178 -143
rect 177 -151 178 -149
rect 184 -145 185 -143
rect 184 -151 185 -149
rect 194 -145 195 -143
rect 191 -151 192 -149
rect 194 -151 195 -149
rect 201 -145 202 -143
rect 198 -151 199 -149
rect 208 -145 209 -143
rect 205 -151 206 -149
rect 208 -151 209 -149
rect 212 -145 213 -143
rect 212 -151 213 -149
rect 219 -145 220 -143
rect 219 -151 220 -149
rect 226 -145 227 -143
rect 226 -151 227 -149
rect 233 -145 234 -143
rect 233 -151 234 -149
rect 240 -145 241 -143
rect 240 -151 241 -149
rect 247 -145 248 -143
rect 247 -151 248 -149
rect 254 -145 255 -143
rect 254 -151 255 -149
rect 261 -145 262 -143
rect 261 -151 262 -149
rect 271 -145 272 -143
rect 268 -151 269 -149
rect 275 -145 276 -143
rect 275 -151 276 -149
rect 282 -145 283 -143
rect 282 -151 283 -149
rect 289 -145 290 -143
rect 289 -151 290 -149
rect 296 -145 297 -143
rect 296 -151 297 -149
rect 303 -145 304 -143
rect 303 -151 304 -149
rect 310 -145 311 -143
rect 310 -151 311 -149
rect 317 -145 318 -143
rect 317 -151 318 -149
rect 324 -145 325 -143
rect 324 -151 325 -149
rect 331 -145 332 -143
rect 331 -151 332 -149
rect 338 -145 339 -143
rect 338 -151 339 -149
rect 345 -145 346 -143
rect 345 -151 346 -149
rect 352 -145 353 -143
rect 352 -151 353 -149
rect 359 -145 360 -143
rect 359 -151 360 -149
rect 366 -145 367 -143
rect 366 -151 367 -149
rect 373 -145 374 -143
rect 373 -151 374 -149
rect 5 -196 6 -194
rect 9 -196 10 -194
rect 9 -202 10 -200
rect 16 -196 17 -194
rect 16 -202 17 -200
rect 23 -196 24 -194
rect 26 -196 27 -194
rect 30 -196 31 -194
rect 30 -202 31 -200
rect 37 -196 38 -194
rect 37 -202 38 -200
rect 47 -196 48 -194
rect 44 -202 45 -200
rect 51 -196 52 -194
rect 51 -202 52 -200
rect 61 -196 62 -194
rect 58 -202 59 -200
rect 65 -196 66 -194
rect 65 -202 66 -200
rect 72 -196 73 -194
rect 75 -196 76 -194
rect 75 -202 76 -200
rect 79 -196 80 -194
rect 82 -196 83 -194
rect 82 -202 83 -200
rect 86 -196 87 -194
rect 86 -202 87 -200
rect 96 -196 97 -194
rect 100 -196 101 -194
rect 103 -196 104 -194
rect 100 -202 101 -200
rect 107 -196 108 -194
rect 107 -202 108 -200
rect 114 -196 115 -194
rect 114 -202 115 -200
rect 121 -196 122 -194
rect 121 -202 122 -200
rect 128 -196 129 -194
rect 128 -202 129 -200
rect 135 -202 136 -200
rect 142 -196 143 -194
rect 142 -202 143 -200
rect 149 -196 150 -194
rect 152 -196 153 -194
rect 149 -202 150 -200
rect 156 -196 157 -194
rect 156 -202 157 -200
rect 163 -196 164 -194
rect 166 -196 167 -194
rect 166 -202 167 -200
rect 173 -196 174 -194
rect 177 -196 178 -194
rect 177 -202 178 -200
rect 184 -196 185 -194
rect 187 -202 188 -200
rect 191 -196 192 -194
rect 191 -202 192 -200
rect 198 -196 199 -194
rect 198 -202 199 -200
rect 201 -202 202 -200
rect 205 -196 206 -194
rect 208 -196 209 -194
rect 205 -202 206 -200
rect 212 -196 213 -194
rect 212 -202 213 -200
rect 219 -196 220 -194
rect 222 -196 223 -194
rect 219 -202 220 -200
rect 222 -202 223 -200
rect 226 -196 227 -194
rect 226 -202 227 -200
rect 233 -196 234 -194
rect 233 -202 234 -200
rect 240 -196 241 -194
rect 240 -202 241 -200
rect 247 -196 248 -194
rect 247 -202 248 -200
rect 254 -196 255 -194
rect 254 -202 255 -200
rect 261 -196 262 -194
rect 261 -202 262 -200
rect 268 -196 269 -194
rect 268 -202 269 -200
rect 275 -196 276 -194
rect 275 -202 276 -200
rect 282 -196 283 -194
rect 282 -202 283 -200
rect 289 -196 290 -194
rect 289 -202 290 -200
rect 296 -196 297 -194
rect 296 -202 297 -200
rect 303 -196 304 -194
rect 303 -202 304 -200
rect 310 -196 311 -194
rect 310 -202 311 -200
rect 320 -196 321 -194
rect 324 -196 325 -194
rect 324 -202 325 -200
rect 331 -196 332 -194
rect 331 -202 332 -200
rect 338 -196 339 -194
rect 338 -202 339 -200
rect 345 -196 346 -194
rect 345 -202 346 -200
rect 352 -196 353 -194
rect 352 -202 353 -200
rect 359 -196 360 -194
rect 359 -202 360 -200
rect 366 -196 367 -194
rect 366 -202 367 -200
rect 373 -196 374 -194
rect 373 -202 374 -200
rect 380 -196 381 -194
rect 380 -202 381 -200
rect 387 -196 388 -194
rect 387 -202 388 -200
rect 394 -196 395 -194
rect 394 -202 395 -200
rect 401 -196 402 -194
rect 401 -202 402 -200
rect 408 -196 409 -194
rect 415 -196 416 -194
rect 415 -202 416 -200
rect 9 -255 10 -253
rect 12 -261 13 -259
rect 16 -255 17 -253
rect 16 -261 17 -259
rect 23 -255 24 -253
rect 23 -261 24 -259
rect 30 -255 31 -253
rect 33 -261 34 -259
rect 37 -255 38 -253
rect 37 -261 38 -259
rect 44 -255 45 -253
rect 44 -261 45 -259
rect 54 -255 55 -253
rect 54 -261 55 -259
rect 58 -255 59 -253
rect 58 -261 59 -259
rect 65 -255 66 -253
rect 65 -261 66 -259
rect 72 -255 73 -253
rect 75 -261 76 -259
rect 79 -255 80 -253
rect 82 -255 83 -253
rect 79 -261 80 -259
rect 86 -255 87 -253
rect 86 -261 87 -259
rect 93 -255 94 -253
rect 96 -255 97 -253
rect 96 -261 97 -259
rect 100 -261 101 -259
rect 103 -261 104 -259
rect 107 -255 108 -253
rect 110 -255 111 -253
rect 110 -261 111 -259
rect 114 -255 115 -253
rect 117 -255 118 -253
rect 117 -261 118 -259
rect 121 -255 122 -253
rect 124 -255 125 -253
rect 128 -255 129 -253
rect 128 -261 129 -259
rect 138 -255 139 -253
rect 135 -261 136 -259
rect 138 -261 139 -259
rect 142 -255 143 -253
rect 142 -261 143 -259
rect 149 -255 150 -253
rect 149 -261 150 -259
rect 156 -255 157 -253
rect 156 -261 157 -259
rect 163 -255 164 -253
rect 163 -261 164 -259
rect 170 -255 171 -253
rect 170 -261 171 -259
rect 177 -255 178 -253
rect 180 -255 181 -253
rect 180 -261 181 -259
rect 184 -255 185 -253
rect 187 -255 188 -253
rect 184 -261 185 -259
rect 191 -255 192 -253
rect 191 -261 192 -259
rect 198 -255 199 -253
rect 201 -255 202 -253
rect 198 -261 199 -259
rect 201 -261 202 -259
rect 205 -255 206 -253
rect 205 -261 206 -259
rect 212 -255 213 -253
rect 212 -261 213 -259
rect 222 -255 223 -253
rect 222 -261 223 -259
rect 226 -255 227 -253
rect 226 -261 227 -259
rect 233 -255 234 -253
rect 233 -261 234 -259
rect 240 -255 241 -253
rect 240 -261 241 -259
rect 243 -261 244 -259
rect 247 -255 248 -253
rect 247 -261 248 -259
rect 254 -255 255 -253
rect 254 -261 255 -259
rect 261 -255 262 -253
rect 261 -261 262 -259
rect 268 -255 269 -253
rect 268 -261 269 -259
rect 275 -255 276 -253
rect 275 -261 276 -259
rect 282 -255 283 -253
rect 289 -255 290 -253
rect 289 -261 290 -259
rect 296 -255 297 -253
rect 296 -261 297 -259
rect 303 -255 304 -253
rect 303 -261 304 -259
rect 310 -255 311 -253
rect 310 -261 311 -259
rect 317 -255 318 -253
rect 317 -261 318 -259
rect 324 -255 325 -253
rect 324 -261 325 -259
rect 331 -255 332 -253
rect 331 -261 332 -259
rect 338 -255 339 -253
rect 338 -261 339 -259
rect 345 -255 346 -253
rect 345 -261 346 -259
rect 352 -255 353 -253
rect 352 -261 353 -259
rect 359 -255 360 -253
rect 359 -261 360 -259
rect 366 -255 367 -253
rect 366 -261 367 -259
rect 373 -255 374 -253
rect 373 -261 374 -259
rect 380 -255 381 -253
rect 380 -261 381 -259
rect 387 -255 388 -253
rect 387 -261 388 -259
rect 394 -255 395 -253
rect 394 -261 395 -259
rect 401 -255 402 -253
rect 401 -261 402 -259
rect 408 -255 409 -253
rect 408 -261 409 -259
rect 415 -255 416 -253
rect 415 -261 416 -259
rect 16 -304 17 -302
rect 16 -310 17 -308
rect 23 -304 24 -302
rect 23 -310 24 -308
rect 30 -304 31 -302
rect 30 -310 31 -308
rect 37 -304 38 -302
rect 37 -310 38 -308
rect 44 -304 45 -302
rect 44 -310 45 -308
rect 51 -304 52 -302
rect 51 -310 52 -308
rect 61 -304 62 -302
rect 61 -310 62 -308
rect 65 -304 66 -302
rect 65 -310 66 -308
rect 72 -304 73 -302
rect 72 -310 73 -308
rect 79 -304 80 -302
rect 79 -310 80 -308
rect 86 -304 87 -302
rect 86 -310 87 -308
rect 93 -304 94 -302
rect 93 -310 94 -308
rect 100 -304 101 -302
rect 103 -310 104 -308
rect 107 -304 108 -302
rect 110 -310 111 -308
rect 114 -304 115 -302
rect 117 -310 118 -308
rect 124 -304 125 -302
rect 121 -310 122 -308
rect 124 -310 125 -308
rect 128 -304 129 -302
rect 128 -310 129 -308
rect 135 -304 136 -302
rect 135 -310 136 -308
rect 142 -304 143 -302
rect 142 -310 143 -308
rect 149 -304 150 -302
rect 149 -310 150 -308
rect 156 -304 157 -302
rect 156 -310 157 -308
rect 163 -304 164 -302
rect 166 -304 167 -302
rect 170 -304 171 -302
rect 173 -304 174 -302
rect 170 -310 171 -308
rect 173 -310 174 -308
rect 177 -304 178 -302
rect 177 -310 178 -308
rect 184 -304 185 -302
rect 184 -310 185 -308
rect 191 -304 192 -302
rect 191 -310 192 -308
rect 198 -304 199 -302
rect 201 -304 202 -302
rect 198 -310 199 -308
rect 205 -304 206 -302
rect 205 -310 206 -308
rect 212 -304 213 -302
rect 212 -310 213 -308
rect 219 -304 220 -302
rect 219 -310 220 -308
rect 226 -304 227 -302
rect 226 -310 227 -308
rect 233 -304 234 -302
rect 233 -310 234 -308
rect 240 -304 241 -302
rect 243 -310 244 -308
rect 247 -304 248 -302
rect 250 -304 251 -302
rect 250 -310 251 -308
rect 254 -304 255 -302
rect 254 -310 255 -308
rect 261 -304 262 -302
rect 264 -304 265 -302
rect 264 -310 265 -308
rect 268 -304 269 -302
rect 268 -310 269 -308
rect 275 -304 276 -302
rect 275 -310 276 -308
rect 282 -304 283 -302
rect 282 -310 283 -308
rect 289 -304 290 -302
rect 289 -310 290 -308
rect 296 -304 297 -302
rect 296 -310 297 -308
rect 303 -304 304 -302
rect 303 -310 304 -308
rect 310 -304 311 -302
rect 310 -310 311 -308
rect 317 -304 318 -302
rect 317 -310 318 -308
rect 324 -304 325 -302
rect 324 -310 325 -308
rect 331 -304 332 -302
rect 331 -310 332 -308
rect 338 -304 339 -302
rect 338 -310 339 -308
rect 345 -304 346 -302
rect 345 -310 346 -308
rect 352 -304 353 -302
rect 352 -310 353 -308
rect 359 -304 360 -302
rect 359 -310 360 -308
rect 366 -304 367 -302
rect 366 -310 367 -308
rect 373 -304 374 -302
rect 373 -310 374 -308
rect 380 -304 381 -302
rect 380 -310 381 -308
rect 387 -304 388 -302
rect 387 -310 388 -308
rect 394 -304 395 -302
rect 394 -310 395 -308
rect 401 -304 402 -302
rect 401 -310 402 -308
rect 408 -304 409 -302
rect 408 -310 409 -308
rect 415 -304 416 -302
rect 415 -310 416 -308
rect 422 -304 423 -302
rect 425 -304 426 -302
rect 425 -310 426 -308
rect 432 -304 433 -302
rect 436 -304 437 -302
rect 436 -310 437 -308
rect 2 -365 3 -363
rect 2 -371 3 -369
rect 16 -365 17 -363
rect 16 -371 17 -369
rect 23 -365 24 -363
rect 26 -365 27 -363
rect 26 -371 27 -369
rect 30 -365 31 -363
rect 33 -365 34 -363
rect 30 -371 31 -369
rect 37 -365 38 -363
rect 40 -365 41 -363
rect 37 -371 38 -369
rect 47 -371 48 -369
rect 51 -365 52 -363
rect 54 -365 55 -363
rect 58 -365 59 -363
rect 58 -371 59 -369
rect 65 -365 66 -363
rect 68 -365 69 -363
rect 68 -371 69 -369
rect 72 -371 73 -369
rect 79 -365 80 -363
rect 79 -371 80 -369
rect 82 -371 83 -369
rect 86 -371 87 -369
rect 89 -371 90 -369
rect 93 -365 94 -363
rect 93 -371 94 -369
rect 100 -365 101 -363
rect 100 -371 101 -369
rect 107 -365 108 -363
rect 110 -365 111 -363
rect 110 -371 111 -369
rect 114 -365 115 -363
rect 117 -365 118 -363
rect 117 -371 118 -369
rect 121 -365 122 -363
rect 121 -371 122 -369
rect 128 -365 129 -363
rect 128 -371 129 -369
rect 135 -365 136 -363
rect 135 -371 136 -369
rect 142 -365 143 -363
rect 142 -371 143 -369
rect 149 -365 150 -363
rect 149 -371 150 -369
rect 156 -365 157 -363
rect 159 -365 160 -363
rect 156 -371 157 -369
rect 159 -371 160 -369
rect 163 -365 164 -363
rect 163 -371 164 -369
rect 170 -371 171 -369
rect 173 -371 174 -369
rect 177 -365 178 -363
rect 177 -371 178 -369
rect 187 -365 188 -363
rect 184 -371 185 -369
rect 191 -365 192 -363
rect 191 -371 192 -369
rect 198 -365 199 -363
rect 198 -371 199 -369
rect 205 -365 206 -363
rect 205 -371 206 -369
rect 212 -365 213 -363
rect 212 -371 213 -369
rect 222 -365 223 -363
rect 219 -371 220 -369
rect 222 -371 223 -369
rect 226 -365 227 -363
rect 226 -371 227 -369
rect 233 -365 234 -363
rect 236 -371 237 -369
rect 240 -365 241 -363
rect 240 -371 241 -369
rect 247 -365 248 -363
rect 247 -371 248 -369
rect 254 -365 255 -363
rect 254 -371 255 -369
rect 257 -371 258 -369
rect 261 -365 262 -363
rect 261 -371 262 -369
rect 268 -365 269 -363
rect 271 -365 272 -363
rect 271 -371 272 -369
rect 275 -365 276 -363
rect 275 -371 276 -369
rect 282 -365 283 -363
rect 282 -371 283 -369
rect 289 -365 290 -363
rect 289 -371 290 -369
rect 296 -365 297 -363
rect 296 -371 297 -369
rect 303 -365 304 -363
rect 303 -371 304 -369
rect 310 -365 311 -363
rect 310 -371 311 -369
rect 317 -365 318 -363
rect 317 -371 318 -369
rect 324 -365 325 -363
rect 324 -371 325 -369
rect 331 -365 332 -363
rect 331 -371 332 -369
rect 338 -365 339 -363
rect 338 -371 339 -369
rect 345 -365 346 -363
rect 345 -371 346 -369
rect 352 -365 353 -363
rect 352 -371 353 -369
rect 359 -365 360 -363
rect 359 -371 360 -369
rect 366 -365 367 -363
rect 366 -371 367 -369
rect 373 -365 374 -363
rect 373 -371 374 -369
rect 380 -365 381 -363
rect 380 -371 381 -369
rect 387 -365 388 -363
rect 387 -371 388 -369
rect 394 -365 395 -363
rect 394 -371 395 -369
rect 401 -365 402 -363
rect 401 -371 402 -369
rect 408 -365 409 -363
rect 408 -371 409 -369
rect 415 -365 416 -363
rect 415 -371 416 -369
rect 422 -365 423 -363
rect 422 -371 423 -369
rect 429 -365 430 -363
rect 429 -371 430 -369
rect 436 -365 437 -363
rect 436 -371 437 -369
rect 9 -414 10 -412
rect 9 -420 10 -418
rect 16 -414 17 -412
rect 16 -420 17 -418
rect 23 -414 24 -412
rect 30 -414 31 -412
rect 30 -420 31 -418
rect 37 -414 38 -412
rect 37 -420 38 -418
rect 47 -414 48 -412
rect 44 -420 45 -418
rect 47 -420 48 -418
rect 51 -414 52 -412
rect 54 -414 55 -412
rect 51 -420 52 -418
rect 58 -414 59 -412
rect 61 -414 62 -412
rect 65 -414 66 -412
rect 65 -420 66 -418
rect 72 -414 73 -412
rect 72 -420 73 -418
rect 79 -414 80 -412
rect 79 -420 80 -418
rect 86 -414 87 -412
rect 86 -420 87 -418
rect 93 -414 94 -412
rect 93 -420 94 -418
rect 100 -414 101 -412
rect 100 -420 101 -418
rect 110 -414 111 -412
rect 107 -420 108 -418
rect 114 -414 115 -412
rect 117 -414 118 -412
rect 117 -420 118 -418
rect 121 -414 122 -412
rect 121 -420 122 -418
rect 128 -420 129 -418
rect 131 -420 132 -418
rect 135 -414 136 -412
rect 135 -420 136 -418
rect 142 -414 143 -412
rect 142 -420 143 -418
rect 149 -414 150 -412
rect 149 -420 150 -418
rect 156 -414 157 -412
rect 156 -420 157 -418
rect 163 -414 164 -412
rect 166 -414 167 -412
rect 163 -420 164 -418
rect 166 -420 167 -418
rect 170 -414 171 -412
rect 170 -420 171 -418
rect 177 -414 178 -412
rect 177 -420 178 -418
rect 184 -414 185 -412
rect 184 -420 185 -418
rect 191 -414 192 -412
rect 191 -420 192 -418
rect 201 -414 202 -412
rect 205 -414 206 -412
rect 205 -420 206 -418
rect 212 -414 213 -412
rect 212 -420 213 -418
rect 219 -414 220 -412
rect 219 -420 220 -418
rect 229 -414 230 -412
rect 226 -420 227 -418
rect 233 -414 234 -412
rect 233 -420 234 -418
rect 240 -414 241 -412
rect 240 -420 241 -418
rect 250 -414 251 -412
rect 247 -420 248 -418
rect 250 -420 251 -418
rect 254 -414 255 -412
rect 254 -420 255 -418
rect 261 -414 262 -412
rect 264 -414 265 -412
rect 261 -420 262 -418
rect 268 -414 269 -412
rect 271 -414 272 -412
rect 268 -420 269 -418
rect 275 -414 276 -412
rect 275 -420 276 -418
rect 282 -414 283 -412
rect 282 -420 283 -418
rect 289 -414 290 -412
rect 289 -420 290 -418
rect 296 -414 297 -412
rect 296 -420 297 -418
rect 303 -414 304 -412
rect 303 -420 304 -418
rect 310 -414 311 -412
rect 310 -420 311 -418
rect 317 -414 318 -412
rect 317 -420 318 -418
rect 327 -414 328 -412
rect 324 -420 325 -418
rect 327 -420 328 -418
rect 334 -420 335 -418
rect 338 -414 339 -412
rect 338 -420 339 -418
rect 345 -414 346 -412
rect 345 -420 346 -418
rect 352 -414 353 -412
rect 352 -420 353 -418
rect 359 -414 360 -412
rect 359 -420 360 -418
rect 366 -414 367 -412
rect 366 -420 367 -418
rect 373 -414 374 -412
rect 373 -420 374 -418
rect 380 -414 381 -412
rect 380 -420 381 -418
rect 387 -414 388 -412
rect 387 -420 388 -418
rect 394 -414 395 -412
rect 394 -420 395 -418
rect 401 -414 402 -412
rect 401 -420 402 -418
rect 408 -414 409 -412
rect 408 -420 409 -418
rect 415 -414 416 -412
rect 415 -420 416 -418
rect 422 -414 423 -412
rect 422 -420 423 -418
rect 429 -414 430 -412
rect 432 -414 433 -412
rect 432 -420 433 -418
rect 436 -414 437 -412
rect 436 -420 437 -418
rect 443 -420 444 -418
rect 16 -469 17 -467
rect 16 -475 17 -473
rect 26 -469 27 -467
rect 33 -469 34 -467
rect 37 -469 38 -467
rect 37 -475 38 -473
rect 51 -469 52 -467
rect 51 -475 52 -473
rect 58 -469 59 -467
rect 58 -475 59 -473
rect 65 -469 66 -467
rect 65 -475 66 -473
rect 72 -469 73 -467
rect 75 -469 76 -467
rect 72 -475 73 -473
rect 79 -469 80 -467
rect 79 -475 80 -473
rect 86 -469 87 -467
rect 86 -475 87 -473
rect 93 -469 94 -467
rect 93 -475 94 -473
rect 100 -469 101 -467
rect 100 -475 101 -473
rect 107 -469 108 -467
rect 107 -475 108 -473
rect 110 -475 111 -473
rect 114 -469 115 -467
rect 114 -475 115 -473
rect 121 -469 122 -467
rect 121 -475 122 -473
rect 128 -469 129 -467
rect 128 -475 129 -473
rect 131 -475 132 -473
rect 135 -469 136 -467
rect 135 -475 136 -473
rect 142 -469 143 -467
rect 142 -475 143 -473
rect 149 -469 150 -467
rect 149 -475 150 -473
rect 156 -469 157 -467
rect 156 -475 157 -473
rect 163 -469 164 -467
rect 163 -475 164 -473
rect 170 -469 171 -467
rect 170 -475 171 -473
rect 177 -469 178 -467
rect 180 -469 181 -467
rect 180 -475 181 -473
rect 184 -469 185 -467
rect 184 -475 185 -473
rect 191 -469 192 -467
rect 194 -469 195 -467
rect 191 -475 192 -473
rect 194 -475 195 -473
rect 198 -469 199 -467
rect 201 -469 202 -467
rect 205 -469 206 -467
rect 205 -475 206 -473
rect 212 -469 213 -467
rect 215 -469 216 -467
rect 212 -475 213 -473
rect 222 -469 223 -467
rect 222 -475 223 -473
rect 226 -469 227 -467
rect 229 -469 230 -467
rect 236 -469 237 -467
rect 236 -475 237 -473
rect 243 -469 244 -467
rect 250 -469 251 -467
rect 247 -475 248 -473
rect 250 -475 251 -473
rect 254 -469 255 -467
rect 257 -469 258 -467
rect 261 -469 262 -467
rect 261 -475 262 -473
rect 264 -475 265 -473
rect 268 -469 269 -467
rect 268 -475 269 -473
rect 275 -469 276 -467
rect 275 -475 276 -473
rect 282 -469 283 -467
rect 282 -475 283 -473
rect 285 -475 286 -473
rect 289 -469 290 -467
rect 289 -475 290 -473
rect 296 -469 297 -467
rect 296 -475 297 -473
rect 303 -469 304 -467
rect 303 -475 304 -473
rect 310 -469 311 -467
rect 310 -475 311 -473
rect 317 -469 318 -467
rect 317 -475 318 -473
rect 324 -469 325 -467
rect 324 -475 325 -473
rect 331 -469 332 -467
rect 331 -475 332 -473
rect 338 -469 339 -467
rect 338 -475 339 -473
rect 345 -469 346 -467
rect 345 -475 346 -473
rect 352 -469 353 -467
rect 352 -475 353 -473
rect 359 -469 360 -467
rect 359 -475 360 -473
rect 366 -469 367 -467
rect 366 -475 367 -473
rect 373 -469 374 -467
rect 373 -475 374 -473
rect 380 -469 381 -467
rect 380 -475 381 -473
rect 387 -469 388 -467
rect 387 -475 388 -473
rect 394 -469 395 -467
rect 394 -475 395 -473
rect 415 -469 416 -467
rect 415 -475 416 -473
rect 422 -469 423 -467
rect 422 -475 423 -473
rect 432 -469 433 -467
rect 429 -475 430 -473
rect 436 -469 437 -467
rect 436 -475 437 -473
rect 446 -469 447 -467
rect 446 -475 447 -473
rect 450 -469 451 -467
rect 450 -475 451 -473
rect 457 -469 458 -467
rect 457 -475 458 -473
rect 464 -469 465 -467
rect 464 -475 465 -473
rect 9 -510 10 -508
rect 9 -516 10 -514
rect 16 -510 17 -508
rect 16 -516 17 -514
rect 23 -510 24 -508
rect 30 -510 31 -508
rect 33 -510 34 -508
rect 30 -516 31 -514
rect 37 -510 38 -508
rect 40 -510 41 -508
rect 37 -516 38 -514
rect 40 -516 41 -514
rect 44 -510 45 -508
rect 44 -516 45 -514
rect 51 -510 52 -508
rect 51 -516 52 -514
rect 58 -510 59 -508
rect 58 -516 59 -514
rect 65 -510 66 -508
rect 65 -516 66 -514
rect 72 -510 73 -508
rect 72 -516 73 -514
rect 79 -510 80 -508
rect 82 -510 83 -508
rect 82 -516 83 -514
rect 86 -510 87 -508
rect 86 -516 87 -514
rect 93 -510 94 -508
rect 93 -516 94 -514
rect 103 -510 104 -508
rect 103 -516 104 -514
rect 107 -510 108 -508
rect 107 -516 108 -514
rect 114 -510 115 -508
rect 114 -516 115 -514
rect 121 -510 122 -508
rect 124 -510 125 -508
rect 121 -516 122 -514
rect 124 -516 125 -514
rect 128 -510 129 -508
rect 128 -516 129 -514
rect 138 -510 139 -508
rect 138 -516 139 -514
rect 142 -510 143 -508
rect 142 -516 143 -514
rect 149 -510 150 -508
rect 149 -516 150 -514
rect 156 -510 157 -508
rect 156 -516 157 -514
rect 163 -510 164 -508
rect 163 -516 164 -514
rect 173 -510 174 -508
rect 173 -516 174 -514
rect 177 -510 178 -508
rect 177 -516 178 -514
rect 184 -510 185 -508
rect 184 -516 185 -514
rect 191 -510 192 -508
rect 191 -516 192 -514
rect 198 -510 199 -508
rect 198 -516 199 -514
rect 205 -510 206 -508
rect 205 -516 206 -514
rect 208 -516 209 -514
rect 215 -510 216 -508
rect 212 -516 213 -514
rect 215 -516 216 -514
rect 219 -510 220 -508
rect 219 -516 220 -514
rect 226 -510 227 -508
rect 226 -516 227 -514
rect 233 -510 234 -508
rect 233 -516 234 -514
rect 240 -510 241 -508
rect 243 -510 244 -508
rect 243 -516 244 -514
rect 247 -510 248 -508
rect 247 -516 248 -514
rect 254 -510 255 -508
rect 254 -516 255 -514
rect 261 -510 262 -508
rect 261 -516 262 -514
rect 268 -510 269 -508
rect 268 -516 269 -514
rect 275 -516 276 -514
rect 278 -516 279 -514
rect 282 -516 283 -514
rect 289 -510 290 -508
rect 289 -516 290 -514
rect 296 -510 297 -508
rect 296 -516 297 -514
rect 303 -510 304 -508
rect 303 -516 304 -514
rect 306 -516 307 -514
rect 310 -510 311 -508
rect 310 -516 311 -514
rect 317 -510 318 -508
rect 317 -516 318 -514
rect 324 -510 325 -508
rect 324 -516 325 -514
rect 331 -510 332 -508
rect 331 -516 332 -514
rect 338 -510 339 -508
rect 338 -516 339 -514
rect 345 -510 346 -508
rect 345 -516 346 -514
rect 352 -510 353 -508
rect 352 -516 353 -514
rect 359 -510 360 -508
rect 359 -516 360 -514
rect 366 -516 367 -514
rect 373 -510 374 -508
rect 373 -516 374 -514
rect 380 -510 381 -508
rect 380 -516 381 -514
rect 387 -510 388 -508
rect 387 -516 388 -514
rect 401 -510 402 -508
rect 401 -516 402 -514
rect 408 -510 409 -508
rect 408 -516 409 -514
rect 415 -510 416 -508
rect 418 -510 419 -508
rect 415 -516 416 -514
rect 429 -510 430 -508
rect 432 -510 433 -508
rect 432 -516 433 -514
rect 436 -510 437 -508
rect 436 -516 437 -514
rect 443 -510 444 -508
rect 443 -516 444 -514
rect 450 -510 451 -508
rect 450 -516 451 -514
rect 457 -510 458 -508
rect 457 -516 458 -514
rect 464 -510 465 -508
rect 464 -516 465 -514
rect 9 -563 10 -561
rect 9 -569 10 -567
rect 19 -563 20 -561
rect 16 -569 17 -567
rect 23 -563 24 -561
rect 26 -563 27 -561
rect 30 -563 31 -561
rect 30 -569 31 -567
rect 37 -563 38 -561
rect 37 -569 38 -567
rect 44 -563 45 -561
rect 44 -569 45 -567
rect 51 -563 52 -561
rect 51 -569 52 -567
rect 58 -563 59 -561
rect 58 -569 59 -567
rect 65 -563 66 -561
rect 68 -563 69 -561
rect 68 -569 69 -567
rect 72 -563 73 -561
rect 72 -569 73 -567
rect 82 -563 83 -561
rect 79 -569 80 -567
rect 86 -563 87 -561
rect 86 -569 87 -567
rect 93 -563 94 -561
rect 96 -563 97 -561
rect 93 -569 94 -567
rect 103 -563 104 -561
rect 103 -569 104 -567
rect 107 -563 108 -561
rect 107 -569 108 -567
rect 114 -563 115 -561
rect 117 -563 118 -561
rect 124 -563 125 -561
rect 121 -569 122 -567
rect 128 -563 129 -561
rect 128 -569 129 -567
rect 135 -563 136 -561
rect 135 -569 136 -567
rect 142 -563 143 -561
rect 142 -569 143 -567
rect 149 -563 150 -561
rect 149 -569 150 -567
rect 156 -563 157 -561
rect 156 -569 157 -567
rect 163 -563 164 -561
rect 166 -563 167 -561
rect 163 -569 164 -567
rect 170 -563 171 -561
rect 173 -563 174 -561
rect 170 -569 171 -567
rect 173 -569 174 -567
rect 177 -563 178 -561
rect 180 -569 181 -567
rect 184 -563 185 -561
rect 187 -563 188 -561
rect 191 -563 192 -561
rect 191 -569 192 -567
rect 198 -563 199 -561
rect 198 -569 199 -567
rect 205 -563 206 -561
rect 205 -569 206 -567
rect 208 -569 209 -567
rect 212 -563 213 -561
rect 212 -569 213 -567
rect 219 -563 220 -561
rect 219 -569 220 -567
rect 226 -563 227 -561
rect 226 -569 227 -567
rect 233 -563 234 -561
rect 236 -563 237 -561
rect 233 -569 234 -567
rect 236 -569 237 -567
rect 240 -563 241 -561
rect 240 -569 241 -567
rect 243 -569 244 -567
rect 247 -563 248 -561
rect 247 -569 248 -567
rect 254 -563 255 -561
rect 254 -569 255 -567
rect 261 -563 262 -561
rect 261 -569 262 -567
rect 268 -563 269 -561
rect 268 -569 269 -567
rect 275 -563 276 -561
rect 275 -569 276 -567
rect 282 -563 283 -561
rect 285 -563 286 -561
rect 282 -569 283 -567
rect 289 -563 290 -561
rect 289 -569 290 -567
rect 296 -563 297 -561
rect 296 -569 297 -567
rect 303 -569 304 -567
rect 306 -569 307 -567
rect 310 -563 311 -561
rect 310 -569 311 -567
rect 317 -563 318 -561
rect 317 -569 318 -567
rect 324 -563 325 -561
rect 324 -569 325 -567
rect 331 -563 332 -561
rect 331 -569 332 -567
rect 341 -563 342 -561
rect 338 -569 339 -567
rect 341 -569 342 -567
rect 345 -563 346 -561
rect 345 -569 346 -567
rect 352 -563 353 -561
rect 352 -569 353 -567
rect 359 -563 360 -561
rect 359 -569 360 -567
rect 366 -563 367 -561
rect 366 -569 367 -567
rect 373 -563 374 -561
rect 373 -569 374 -567
rect 380 -563 381 -561
rect 380 -569 381 -567
rect 387 -563 388 -561
rect 387 -569 388 -567
rect 394 -563 395 -561
rect 394 -569 395 -567
rect 401 -563 402 -561
rect 401 -569 402 -567
rect 408 -563 409 -561
rect 408 -569 409 -567
rect 415 -563 416 -561
rect 415 -569 416 -567
rect 422 -563 423 -561
rect 422 -569 423 -567
rect 429 -563 430 -561
rect 429 -569 430 -567
rect 436 -563 437 -561
rect 436 -569 437 -567
rect 443 -563 444 -561
rect 443 -569 444 -567
rect 457 -563 458 -561
rect 464 -563 465 -561
rect 464 -569 465 -567
rect 9 -616 10 -614
rect 9 -622 10 -620
rect 16 -616 17 -614
rect 16 -622 17 -620
rect 23 -616 24 -614
rect 23 -622 24 -620
rect 30 -616 31 -614
rect 33 -616 34 -614
rect 33 -622 34 -620
rect 40 -616 41 -614
rect 37 -622 38 -620
rect 40 -622 41 -620
rect 44 -616 45 -614
rect 44 -622 45 -620
rect 51 -616 52 -614
rect 51 -622 52 -620
rect 58 -616 59 -614
rect 58 -622 59 -620
rect 65 -616 66 -614
rect 65 -622 66 -620
rect 72 -616 73 -614
rect 72 -622 73 -620
rect 79 -616 80 -614
rect 79 -622 80 -620
rect 86 -616 87 -614
rect 89 -616 90 -614
rect 89 -622 90 -620
rect 93 -616 94 -614
rect 93 -622 94 -620
rect 100 -616 101 -614
rect 100 -622 101 -620
rect 103 -622 104 -620
rect 107 -616 108 -614
rect 107 -622 108 -620
rect 114 -616 115 -614
rect 114 -622 115 -620
rect 117 -622 118 -620
rect 121 -616 122 -614
rect 121 -622 122 -620
rect 128 -622 129 -620
rect 131 -622 132 -620
rect 138 -616 139 -614
rect 135 -622 136 -620
rect 142 -616 143 -614
rect 142 -622 143 -620
rect 149 -616 150 -614
rect 149 -622 150 -620
rect 156 -616 157 -614
rect 156 -622 157 -620
rect 163 -616 164 -614
rect 163 -622 164 -620
rect 170 -616 171 -614
rect 173 -616 174 -614
rect 170 -622 171 -620
rect 177 -616 178 -614
rect 177 -622 178 -620
rect 184 -616 185 -614
rect 184 -622 185 -620
rect 194 -616 195 -614
rect 191 -622 192 -620
rect 194 -622 195 -620
rect 198 -616 199 -614
rect 198 -622 199 -620
rect 208 -616 209 -614
rect 208 -622 209 -620
rect 212 -622 213 -620
rect 215 -622 216 -620
rect 219 -616 220 -614
rect 219 -622 220 -620
rect 226 -616 227 -614
rect 226 -622 227 -620
rect 233 -616 234 -614
rect 233 -622 234 -620
rect 240 -616 241 -614
rect 240 -622 241 -620
rect 247 -616 248 -614
rect 250 -622 251 -620
rect 257 -616 258 -614
rect 254 -622 255 -620
rect 264 -616 265 -614
rect 261 -622 262 -620
rect 268 -616 269 -614
rect 268 -622 269 -620
rect 275 -616 276 -614
rect 275 -622 276 -620
rect 282 -616 283 -614
rect 282 -622 283 -620
rect 289 -616 290 -614
rect 289 -622 290 -620
rect 296 -616 297 -614
rect 299 -622 300 -620
rect 303 -616 304 -614
rect 303 -622 304 -620
rect 310 -616 311 -614
rect 310 -622 311 -620
rect 317 -616 318 -614
rect 317 -622 318 -620
rect 324 -616 325 -614
rect 324 -622 325 -620
rect 331 -616 332 -614
rect 331 -622 332 -620
rect 334 -622 335 -620
rect 338 -616 339 -614
rect 338 -622 339 -620
rect 345 -616 346 -614
rect 345 -622 346 -620
rect 352 -616 353 -614
rect 352 -622 353 -620
rect 359 -616 360 -614
rect 359 -622 360 -620
rect 366 -616 367 -614
rect 366 -622 367 -620
rect 373 -616 374 -614
rect 373 -622 374 -620
rect 380 -616 381 -614
rect 380 -622 381 -620
rect 387 -616 388 -614
rect 387 -622 388 -620
rect 394 -616 395 -614
rect 394 -622 395 -620
rect 401 -616 402 -614
rect 401 -622 402 -620
rect 408 -616 409 -614
rect 408 -622 409 -620
rect 415 -616 416 -614
rect 415 -622 416 -620
rect 422 -616 423 -614
rect 422 -622 423 -620
rect 429 -616 430 -614
rect 429 -622 430 -620
rect 436 -616 437 -614
rect 436 -622 437 -620
rect 443 -616 444 -614
rect 446 -616 447 -614
rect 446 -622 447 -620
rect 453 -616 454 -614
rect 450 -622 451 -620
rect 457 -616 458 -614
rect 457 -622 458 -620
rect 464 -616 465 -614
rect 471 -616 472 -614
rect 471 -622 472 -620
rect 2 -667 3 -665
rect 2 -673 3 -671
rect 9 -667 10 -665
rect 9 -673 10 -671
rect 16 -667 17 -665
rect 16 -673 17 -671
rect 23 -667 24 -665
rect 23 -673 24 -671
rect 30 -667 31 -665
rect 30 -673 31 -671
rect 37 -667 38 -665
rect 37 -673 38 -671
rect 44 -667 45 -665
rect 51 -667 52 -665
rect 54 -667 55 -665
rect 54 -673 55 -671
rect 58 -667 59 -665
rect 58 -673 59 -671
rect 65 -667 66 -665
rect 65 -673 66 -671
rect 75 -667 76 -665
rect 72 -673 73 -671
rect 79 -667 80 -665
rect 79 -673 80 -671
rect 86 -667 87 -665
rect 86 -673 87 -671
rect 93 -667 94 -665
rect 93 -673 94 -671
rect 100 -667 101 -665
rect 103 -667 104 -665
rect 100 -673 101 -671
rect 107 -667 108 -665
rect 107 -673 108 -671
rect 114 -667 115 -665
rect 114 -673 115 -671
rect 117 -673 118 -671
rect 121 -667 122 -665
rect 121 -673 122 -671
rect 128 -667 129 -665
rect 128 -673 129 -671
rect 131 -673 132 -671
rect 135 -667 136 -665
rect 135 -673 136 -671
rect 142 -667 143 -665
rect 142 -673 143 -671
rect 149 -667 150 -665
rect 149 -673 150 -671
rect 156 -667 157 -665
rect 156 -673 157 -671
rect 163 -667 164 -665
rect 163 -673 164 -671
rect 170 -667 171 -665
rect 170 -673 171 -671
rect 177 -667 178 -665
rect 180 -667 181 -665
rect 177 -673 178 -671
rect 180 -673 181 -671
rect 184 -667 185 -665
rect 187 -667 188 -665
rect 184 -673 185 -671
rect 194 -667 195 -665
rect 191 -673 192 -671
rect 194 -673 195 -671
rect 198 -667 199 -665
rect 198 -673 199 -671
rect 205 -667 206 -665
rect 208 -667 209 -665
rect 215 -667 216 -665
rect 212 -673 213 -671
rect 215 -673 216 -671
rect 222 -667 223 -665
rect 219 -673 220 -671
rect 226 -667 227 -665
rect 226 -673 227 -671
rect 233 -667 234 -665
rect 233 -673 234 -671
rect 240 -667 241 -665
rect 243 -667 244 -665
rect 240 -673 241 -671
rect 247 -667 248 -665
rect 250 -667 251 -665
rect 250 -673 251 -671
rect 254 -667 255 -665
rect 254 -673 255 -671
rect 261 -667 262 -665
rect 261 -673 262 -671
rect 271 -667 272 -665
rect 268 -673 269 -671
rect 275 -667 276 -665
rect 275 -673 276 -671
rect 282 -667 283 -665
rect 282 -673 283 -671
rect 289 -667 290 -665
rect 289 -673 290 -671
rect 296 -667 297 -665
rect 299 -667 300 -665
rect 299 -673 300 -671
rect 303 -667 304 -665
rect 303 -673 304 -671
rect 310 -667 311 -665
rect 310 -673 311 -671
rect 317 -667 318 -665
rect 317 -673 318 -671
rect 324 -667 325 -665
rect 324 -673 325 -671
rect 331 -667 332 -665
rect 334 -673 335 -671
rect 338 -667 339 -665
rect 338 -673 339 -671
rect 345 -667 346 -665
rect 345 -673 346 -671
rect 352 -667 353 -665
rect 352 -673 353 -671
rect 359 -667 360 -665
rect 359 -673 360 -671
rect 366 -667 367 -665
rect 366 -673 367 -671
rect 373 -667 374 -665
rect 373 -673 374 -671
rect 380 -667 381 -665
rect 380 -673 381 -671
rect 387 -667 388 -665
rect 387 -673 388 -671
rect 394 -667 395 -665
rect 394 -673 395 -671
rect 401 -667 402 -665
rect 401 -673 402 -671
rect 408 -667 409 -665
rect 408 -673 409 -671
rect 415 -667 416 -665
rect 415 -673 416 -671
rect 422 -667 423 -665
rect 422 -673 423 -671
rect 429 -667 430 -665
rect 429 -673 430 -671
rect 436 -667 437 -665
rect 436 -673 437 -671
rect 443 -667 444 -665
rect 443 -673 444 -671
rect 450 -667 451 -665
rect 450 -673 451 -671
rect 457 -667 458 -665
rect 460 -667 461 -665
rect 457 -673 458 -671
rect 464 -667 465 -665
rect 464 -673 465 -671
rect 471 -667 472 -665
rect 471 -673 472 -671
rect 2 -718 3 -716
rect 2 -724 3 -722
rect 9 -718 10 -716
rect 9 -724 10 -722
rect 16 -718 17 -716
rect 16 -724 17 -722
rect 23 -718 24 -716
rect 23 -724 24 -722
rect 30 -718 31 -716
rect 30 -724 31 -722
rect 37 -718 38 -716
rect 40 -718 41 -716
rect 37 -724 38 -722
rect 44 -718 45 -716
rect 44 -724 45 -722
rect 51 -718 52 -716
rect 54 -724 55 -722
rect 58 -718 59 -716
rect 58 -724 59 -722
rect 65 -718 66 -716
rect 65 -724 66 -722
rect 72 -718 73 -716
rect 75 -718 76 -716
rect 75 -724 76 -722
rect 82 -718 83 -716
rect 82 -724 83 -722
rect 86 -718 87 -716
rect 86 -724 87 -722
rect 93 -718 94 -716
rect 93 -724 94 -722
rect 100 -718 101 -716
rect 100 -724 101 -722
rect 107 -718 108 -716
rect 107 -724 108 -722
rect 114 -718 115 -716
rect 114 -724 115 -722
rect 121 -718 122 -716
rect 124 -718 125 -716
rect 131 -718 132 -716
rect 128 -724 129 -722
rect 135 -718 136 -716
rect 135 -724 136 -722
rect 142 -718 143 -716
rect 142 -724 143 -722
rect 149 -718 150 -716
rect 149 -724 150 -722
rect 156 -718 157 -716
rect 156 -724 157 -722
rect 163 -718 164 -716
rect 163 -724 164 -722
rect 170 -718 171 -716
rect 173 -718 174 -716
rect 177 -718 178 -716
rect 180 -724 181 -722
rect 184 -718 185 -716
rect 187 -718 188 -716
rect 184 -724 185 -722
rect 191 -718 192 -716
rect 191 -724 192 -722
rect 198 -718 199 -716
rect 198 -724 199 -722
rect 201 -724 202 -722
rect 205 -718 206 -716
rect 205 -724 206 -722
rect 208 -724 209 -722
rect 212 -718 213 -716
rect 212 -724 213 -722
rect 219 -718 220 -716
rect 219 -724 220 -722
rect 229 -718 230 -716
rect 226 -724 227 -722
rect 233 -718 234 -716
rect 233 -724 234 -722
rect 240 -718 241 -716
rect 243 -724 244 -722
rect 250 -718 251 -716
rect 250 -724 251 -722
rect 254 -718 255 -716
rect 254 -724 255 -722
rect 261 -718 262 -716
rect 261 -724 262 -722
rect 268 -718 269 -716
rect 268 -724 269 -722
rect 278 -724 279 -722
rect 282 -718 283 -716
rect 282 -724 283 -722
rect 289 -718 290 -716
rect 289 -724 290 -722
rect 296 -718 297 -716
rect 296 -724 297 -722
rect 310 -718 311 -716
rect 310 -724 311 -722
rect 317 -718 318 -716
rect 317 -724 318 -722
rect 324 -718 325 -716
rect 324 -724 325 -722
rect 331 -718 332 -716
rect 331 -724 332 -722
rect 341 -724 342 -722
rect 345 -718 346 -716
rect 345 -724 346 -722
rect 352 -718 353 -716
rect 352 -724 353 -722
rect 359 -718 360 -716
rect 359 -724 360 -722
rect 366 -718 367 -716
rect 366 -724 367 -722
rect 373 -718 374 -716
rect 376 -724 377 -722
rect 380 -718 381 -716
rect 380 -724 381 -722
rect 387 -718 388 -716
rect 387 -724 388 -722
rect 394 -718 395 -716
rect 394 -724 395 -722
rect 401 -718 402 -716
rect 401 -724 402 -722
rect 411 -724 412 -722
rect 429 -718 430 -716
rect 429 -724 430 -722
rect 16 -771 17 -769
rect 23 -771 24 -769
rect 23 -777 24 -775
rect 30 -777 31 -775
rect 33 -777 34 -775
rect 37 -771 38 -769
rect 40 -771 41 -769
rect 37 -777 38 -775
rect 44 -771 45 -769
rect 47 -777 48 -775
rect 51 -771 52 -769
rect 51 -777 52 -775
rect 58 -771 59 -769
rect 58 -777 59 -775
rect 65 -771 66 -769
rect 65 -777 66 -775
rect 72 -771 73 -769
rect 75 -771 76 -769
rect 75 -777 76 -775
rect 79 -771 80 -769
rect 82 -771 83 -769
rect 86 -771 87 -769
rect 86 -777 87 -775
rect 96 -771 97 -769
rect 93 -777 94 -775
rect 96 -777 97 -775
rect 100 -771 101 -769
rect 103 -771 104 -769
rect 103 -777 104 -775
rect 110 -771 111 -769
rect 107 -777 108 -775
rect 114 -771 115 -769
rect 117 -777 118 -775
rect 121 -771 122 -769
rect 124 -777 125 -775
rect 128 -771 129 -769
rect 128 -777 129 -775
rect 135 -771 136 -769
rect 135 -777 136 -775
rect 142 -771 143 -769
rect 142 -777 143 -775
rect 149 -771 150 -769
rect 149 -777 150 -775
rect 156 -771 157 -769
rect 156 -777 157 -775
rect 163 -771 164 -769
rect 163 -777 164 -775
rect 170 -771 171 -769
rect 170 -777 171 -775
rect 180 -771 181 -769
rect 177 -777 178 -775
rect 184 -771 185 -769
rect 184 -777 185 -775
rect 191 -771 192 -769
rect 191 -777 192 -775
rect 198 -771 199 -769
rect 198 -777 199 -775
rect 208 -771 209 -769
rect 212 -771 213 -769
rect 215 -771 216 -769
rect 212 -777 213 -775
rect 219 -771 220 -769
rect 219 -777 220 -775
rect 226 -771 227 -769
rect 226 -777 227 -775
rect 233 -771 234 -769
rect 236 -771 237 -769
rect 236 -777 237 -775
rect 240 -771 241 -769
rect 240 -777 241 -775
rect 247 -771 248 -769
rect 247 -777 248 -775
rect 254 -771 255 -769
rect 254 -777 255 -775
rect 261 -771 262 -769
rect 261 -777 262 -775
rect 268 -771 269 -769
rect 268 -777 269 -775
rect 275 -777 276 -775
rect 282 -771 283 -769
rect 282 -777 283 -775
rect 289 -771 290 -769
rect 289 -777 290 -775
rect 303 -771 304 -769
rect 303 -777 304 -775
rect 310 -771 311 -769
rect 310 -777 311 -775
rect 324 -771 325 -769
rect 324 -777 325 -775
rect 331 -771 332 -769
rect 338 -771 339 -769
rect 338 -777 339 -775
rect 345 -771 346 -769
rect 345 -777 346 -775
rect 408 -771 409 -769
rect 9 -816 10 -814
rect 9 -822 10 -820
rect 16 -822 17 -820
rect 23 -816 24 -814
rect 23 -822 24 -820
rect 30 -816 31 -814
rect 33 -816 34 -814
rect 33 -822 34 -820
rect 37 -816 38 -814
rect 37 -822 38 -820
rect 44 -822 45 -820
rect 47 -822 48 -820
rect 51 -816 52 -814
rect 51 -822 52 -820
rect 61 -816 62 -814
rect 65 -822 66 -820
rect 72 -816 73 -814
rect 72 -822 73 -820
rect 79 -816 80 -814
rect 82 -816 83 -814
rect 89 -822 90 -820
rect 96 -822 97 -820
rect 100 -816 101 -814
rect 100 -822 101 -820
rect 107 -816 108 -814
rect 110 -816 111 -814
rect 114 -816 115 -814
rect 117 -816 118 -814
rect 114 -822 115 -820
rect 117 -822 118 -820
rect 124 -816 125 -814
rect 131 -816 132 -814
rect 128 -822 129 -820
rect 135 -816 136 -814
rect 135 -822 136 -820
rect 145 -822 146 -820
rect 152 -816 153 -814
rect 152 -822 153 -820
rect 156 -816 157 -814
rect 156 -822 157 -820
rect 163 -816 164 -814
rect 163 -822 164 -820
rect 170 -816 171 -814
rect 170 -822 171 -820
rect 177 -816 178 -814
rect 180 -822 181 -820
rect 184 -816 185 -814
rect 184 -822 185 -820
rect 191 -816 192 -814
rect 191 -822 192 -820
rect 198 -816 199 -814
rect 198 -822 199 -820
rect 205 -816 206 -814
rect 205 -822 206 -820
rect 212 -816 213 -814
rect 212 -822 213 -820
rect 222 -822 223 -820
rect 226 -816 227 -814
rect 226 -822 227 -820
rect 233 -816 234 -814
rect 233 -822 234 -820
rect 240 -822 241 -820
rect 247 -816 248 -814
rect 247 -822 248 -820
rect 254 -816 255 -814
rect 254 -822 255 -820
rect 261 -816 262 -814
rect 261 -822 262 -820
rect 268 -816 269 -814
rect 268 -822 269 -820
rect 282 -816 283 -814
rect 282 -822 283 -820
rect 289 -816 290 -814
rect 289 -822 290 -820
rect 303 -816 304 -814
rect 303 -822 304 -820
rect 310 -816 311 -814
rect 310 -822 311 -820
rect 317 -816 318 -814
rect 317 -822 318 -820
rect 324 -816 325 -814
rect 324 -822 325 -820
rect 345 -822 346 -820
rect 19 -849 20 -847
rect 23 -849 24 -847
rect 23 -855 24 -853
rect 33 -849 34 -847
rect 37 -849 38 -847
rect 37 -855 38 -853
rect 44 -849 45 -847
rect 44 -855 45 -853
rect 47 -855 48 -853
rect 51 -849 52 -847
rect 54 -855 55 -853
rect 58 -849 59 -847
rect 58 -855 59 -853
rect 65 -855 66 -853
rect 72 -849 73 -847
rect 72 -855 73 -853
rect 79 -849 80 -847
rect 82 -855 83 -853
rect 86 -849 87 -847
rect 86 -855 87 -853
rect 93 -849 94 -847
rect 93 -855 94 -853
rect 103 -855 104 -853
rect 107 -855 108 -853
rect 117 -849 118 -847
rect 114 -855 115 -853
rect 124 -849 125 -847
rect 131 -855 132 -853
rect 135 -849 136 -847
rect 142 -855 143 -853
rect 149 -849 150 -847
rect 149 -855 150 -853
rect 156 -849 157 -847
rect 156 -855 157 -853
rect 163 -849 164 -847
rect 163 -855 164 -853
rect 170 -849 171 -847
rect 170 -855 171 -853
rect 184 -849 185 -847
rect 187 -855 188 -853
rect 191 -849 192 -847
rect 191 -855 192 -853
rect 212 -849 213 -847
rect 226 -849 227 -847
rect 268 -849 269 -847
rect 268 -855 269 -853
rect 282 -849 283 -847
rect 285 -855 286 -853
rect 289 -849 290 -847
rect 292 -849 293 -847
rect 327 -849 328 -847
<< metal1 >>
rect 12 0 27 1
rect 37 0 66 1
rect 93 0 108 1
rect 121 0 129 1
rect 135 0 164 1
rect 51 -2 90 -1
rect 138 -2 150 -1
rect 58 -4 73 -3
rect 72 -15 97 -14
rect 100 -15 108 -14
rect 114 -15 157 -14
rect 159 -15 192 -14
rect 65 -17 73 -16
rect 79 -17 101 -16
rect 107 -17 143 -16
rect 145 -17 150 -16
rect 163 -17 174 -16
rect 114 -19 178 -18
rect 149 -21 202 -20
rect 163 -23 188 -22
rect 47 -34 213 -33
rect 51 -36 150 -35
rect 163 -36 220 -35
rect 58 -38 73 -37
rect 86 -38 164 -37
rect 177 -38 234 -37
rect 16 -40 178 -39
rect 191 -40 255 -39
rect 65 -42 118 -41
rect 121 -42 171 -41
rect 198 -42 248 -41
rect 72 -44 80 -43
rect 93 -44 185 -43
rect 37 -46 94 -45
rect 96 -46 199 -45
rect 124 -48 153 -47
rect 100 -50 125 -49
rect 142 -50 227 -49
rect 145 -52 157 -51
rect 149 -54 206 -53
rect 19 -65 213 -64
rect 219 -65 276 -64
rect 40 -67 80 -66
rect 82 -67 111 -66
rect 121 -67 160 -66
rect 177 -67 220 -66
rect 226 -67 332 -66
rect 40 -69 178 -68
rect 191 -69 255 -68
rect 44 -71 52 -70
rect 58 -71 90 -70
rect 100 -71 129 -70
rect 131 -71 262 -70
rect 30 -73 132 -72
rect 138 -73 143 -72
rect 149 -73 213 -72
rect 233 -73 283 -72
rect 30 -75 115 -74
rect 163 -75 227 -74
rect 243 -75 255 -74
rect 51 -77 97 -76
rect 107 -77 136 -76
rect 184 -77 192 -76
rect 205 -77 241 -76
rect 247 -77 269 -76
rect 58 -79 66 -78
rect 86 -79 157 -78
rect 170 -79 206 -78
rect 65 -81 73 -80
rect 110 -81 297 -80
rect 72 -83 101 -82
rect 170 -83 290 -82
rect 184 -85 234 -84
rect 198 -87 248 -86
rect 23 -98 87 -97
rect 93 -98 132 -97
rect 135 -98 227 -97
rect 268 -98 360 -97
rect 26 -100 353 -99
rect 30 -102 199 -101
rect 201 -102 318 -101
rect 51 -104 101 -103
rect 107 -104 118 -103
rect 121 -104 143 -103
rect 145 -104 311 -103
rect 51 -106 66 -105
rect 96 -106 262 -105
rect 271 -106 367 -105
rect 65 -108 174 -107
rect 194 -108 227 -107
rect 254 -108 262 -107
rect 275 -108 346 -107
rect 30 -110 276 -109
rect 289 -110 374 -109
rect 86 -112 255 -111
rect 303 -112 325 -111
rect 128 -114 248 -113
rect 138 -116 304 -115
rect 138 -118 202 -117
rect 233 -118 290 -117
rect 149 -120 206 -119
rect 233 -120 297 -119
rect 149 -122 209 -121
rect 240 -122 297 -121
rect 152 -124 171 -123
rect 191 -124 248 -123
rect 156 -126 339 -125
rect 44 -128 157 -127
rect 163 -128 283 -127
rect 9 -130 45 -129
rect 124 -130 164 -129
rect 166 -130 220 -129
rect 37 -132 283 -131
rect 166 -134 185 -133
rect 212 -134 241 -133
rect 128 -136 213 -135
rect 177 -138 220 -137
rect 72 -140 178 -139
rect 72 -142 122 -141
rect 5 -153 20 -152
rect 23 -153 311 -152
rect 345 -153 381 -152
rect 9 -155 27 -154
rect 61 -155 339 -154
rect 345 -155 353 -154
rect 373 -155 402 -154
rect 16 -157 38 -156
rect 65 -157 104 -156
rect 128 -157 290 -156
rect 338 -157 367 -156
rect 16 -159 52 -158
rect 86 -159 304 -158
rect 320 -159 367 -158
rect 23 -161 31 -160
rect 37 -161 108 -160
rect 128 -161 199 -160
rect 208 -161 360 -160
rect 30 -163 174 -162
rect 191 -163 374 -162
rect 51 -165 97 -164
rect 107 -165 206 -164
rect 222 -165 388 -164
rect 79 -167 206 -166
rect 226 -167 304 -166
rect 359 -167 409 -166
rect 65 -169 80 -168
rect 86 -169 94 -168
rect 149 -169 185 -168
rect 194 -169 297 -168
rect 89 -171 143 -170
rect 149 -171 297 -170
rect 72 -173 143 -172
rect 152 -173 248 -172
rect 261 -173 416 -172
rect 47 -175 73 -174
rect 156 -175 185 -174
rect 198 -175 311 -174
rect 100 -177 157 -176
rect 163 -177 241 -176
rect 261 -177 283 -176
rect 75 -179 164 -178
rect 166 -179 395 -178
rect 82 -181 241 -180
rect 254 -181 283 -180
rect 82 -183 122 -182
rect 177 -183 192 -182
rect 208 -183 227 -182
rect 233 -183 248 -182
rect 268 -183 318 -182
rect 100 -185 136 -184
rect 152 -185 269 -184
rect 275 -185 290 -184
rect 61 -187 276 -186
rect 114 -189 122 -188
rect 170 -189 178 -188
rect 212 -189 234 -188
rect 44 -191 115 -190
rect 219 -191 255 -190
rect 58 -193 213 -192
rect 219 -193 353 -192
rect 16 -204 73 -203
rect 86 -204 150 -203
rect 166 -204 304 -203
rect 16 -206 181 -205
rect 184 -206 388 -205
rect 23 -208 108 -207
rect 110 -208 199 -207
rect 205 -208 374 -207
rect 44 -210 115 -209
rect 117 -210 276 -209
rect 338 -210 374 -209
rect 44 -212 101 -211
rect 107 -212 304 -211
rect 338 -212 346 -211
rect 54 -214 199 -213
rect 219 -214 416 -213
rect 65 -216 83 -215
rect 86 -216 115 -215
rect 124 -216 129 -215
rect 138 -216 192 -215
rect 240 -216 388 -215
rect 30 -218 129 -217
rect 142 -218 164 -217
rect 170 -218 234 -217
rect 275 -218 290 -217
rect 310 -218 416 -217
rect 9 -220 31 -219
rect 37 -220 143 -219
rect 177 -220 234 -219
rect 289 -220 297 -219
rect 345 -220 353 -219
rect 9 -222 76 -221
rect 93 -222 157 -221
rect 187 -222 318 -221
rect 352 -222 360 -221
rect 37 -224 83 -223
rect 96 -224 395 -223
rect 65 -226 80 -225
rect 121 -226 157 -225
rect 187 -226 206 -225
rect 222 -226 241 -225
rect 261 -226 297 -225
rect 359 -226 367 -225
rect 51 -228 223 -227
rect 121 -230 367 -229
rect 135 -232 395 -231
rect 149 -234 178 -233
rect 191 -234 213 -233
rect 201 -236 262 -235
rect 201 -238 381 -237
rect 58 -240 381 -239
rect 58 -242 227 -241
rect 212 -244 255 -243
rect 226 -246 269 -245
rect 254 -248 409 -247
rect 268 -250 283 -249
rect 282 -252 311 -251
rect 12 -263 339 -262
rect 380 -263 437 -262
rect 33 -265 55 -264
rect 61 -265 66 -264
rect 72 -265 108 -264
rect 110 -265 269 -264
rect 282 -265 433 -264
rect 37 -267 66 -266
rect 75 -267 139 -266
rect 163 -267 185 -266
rect 226 -267 423 -266
rect 30 -269 164 -268
rect 173 -269 213 -268
rect 240 -269 290 -268
rect 338 -269 346 -268
rect 380 -269 426 -268
rect 37 -271 59 -270
rect 86 -271 115 -270
rect 117 -271 143 -270
rect 177 -271 202 -270
rect 205 -271 227 -270
rect 247 -271 255 -270
rect 268 -271 318 -270
rect 345 -271 374 -270
rect 394 -271 398 -270
rect 51 -273 199 -272
rect 212 -273 297 -272
rect 317 -273 332 -272
rect 366 -273 374 -272
rect 394 -273 416 -272
rect 79 -275 87 -274
rect 96 -275 290 -274
rect 331 -275 353 -274
rect 359 -275 367 -274
rect 401 -275 416 -274
rect 23 -277 80 -276
rect 100 -277 143 -276
rect 180 -277 234 -276
rect 250 -277 388 -276
rect 401 -277 409 -276
rect 23 -279 45 -278
rect 100 -279 157 -278
rect 184 -279 276 -278
rect 397 -279 409 -278
rect 44 -281 202 -280
rect 205 -281 353 -280
rect 103 -283 171 -282
rect 198 -283 297 -282
rect 128 -285 241 -284
rect 254 -285 262 -284
rect 275 -285 311 -284
rect 16 -287 262 -286
rect 264 -287 311 -286
rect 16 -289 244 -288
rect 128 -291 171 -290
rect 219 -291 248 -290
rect 135 -293 388 -292
rect 93 -295 136 -294
rect 156 -295 192 -294
rect 222 -295 360 -294
rect 166 -297 192 -296
rect 233 -297 304 -296
rect 303 -299 325 -298
rect 124 -301 325 -300
rect 2 -312 174 -311
rect 184 -312 241 -311
rect 243 -312 339 -311
rect 401 -312 430 -311
rect 23 -314 94 -313
rect 100 -314 129 -313
rect 142 -314 206 -313
rect 233 -314 262 -313
rect 264 -314 416 -313
rect 26 -316 104 -315
rect 107 -316 416 -315
rect 30 -318 188 -317
rect 191 -318 223 -317
rect 247 -318 255 -317
rect 317 -318 339 -317
rect 23 -320 192 -319
rect 198 -320 304 -319
rect 317 -320 325 -319
rect 30 -322 374 -321
rect 37 -324 171 -323
rect 198 -324 220 -323
rect 250 -324 381 -323
rect 33 -326 38 -325
rect 40 -326 402 -325
rect 44 -328 125 -327
rect 142 -328 213 -327
rect 254 -328 423 -327
rect 54 -330 304 -329
rect 345 -330 381 -329
rect 58 -332 87 -331
rect 110 -332 129 -331
rect 159 -332 178 -331
rect 296 -332 325 -331
rect 373 -332 388 -331
rect 61 -334 94 -333
rect 110 -334 346 -333
rect 65 -336 206 -335
rect 233 -336 388 -335
rect 65 -338 297 -337
rect 72 -340 437 -339
rect 79 -342 164 -341
rect 394 -342 437 -341
rect 16 -344 80 -343
rect 114 -344 213 -343
rect 366 -344 395 -343
rect 16 -346 69 -345
rect 121 -346 150 -345
rect 359 -346 367 -345
rect 117 -348 122 -347
rect 135 -348 178 -347
rect 352 -348 360 -347
rect 117 -350 409 -349
rect 51 -352 409 -351
rect 51 -354 150 -353
rect 289 -354 353 -353
rect 135 -356 157 -355
rect 289 -356 311 -355
rect 156 -358 269 -357
rect 282 -358 311 -357
rect 268 -360 426 -359
rect 271 -362 283 -361
rect 2 -373 174 -372
rect 201 -373 220 -372
rect 222 -373 360 -372
rect 9 -375 31 -374
rect 37 -375 90 -374
rect 110 -375 367 -374
rect 16 -377 24 -376
rect 26 -377 237 -376
rect 247 -377 258 -376
rect 268 -377 311 -376
rect 317 -377 367 -376
rect 16 -379 52 -378
rect 65 -379 199 -378
rect 226 -379 234 -378
rect 271 -379 395 -378
rect 30 -381 48 -380
rect 68 -381 192 -380
rect 271 -381 290 -380
rect 317 -381 325 -380
rect 338 -381 360 -380
rect 387 -381 395 -380
rect 37 -383 59 -382
rect 79 -383 328 -382
rect 61 -385 80 -384
rect 82 -385 297 -384
rect 86 -387 206 -386
rect 212 -387 290 -386
rect 72 -389 87 -388
rect 110 -389 346 -388
rect 72 -391 101 -390
rect 114 -391 409 -390
rect 100 -393 164 -392
rect 184 -393 220 -392
rect 229 -393 388 -392
rect 408 -393 430 -392
rect 117 -395 416 -394
rect 135 -397 167 -396
rect 205 -397 251 -396
rect 261 -397 339 -396
rect 352 -397 430 -396
rect 135 -399 160 -398
rect 163 -399 311 -398
rect 331 -399 353 -398
rect 415 -399 423 -398
rect 142 -401 192 -400
rect 212 -401 241 -400
rect 261 -401 402 -400
rect 422 -401 437 -400
rect 93 -403 143 -402
rect 149 -403 157 -402
rect 184 -403 241 -402
rect 275 -403 297 -402
rect 303 -403 346 -402
rect 373 -403 402 -402
rect 432 -403 437 -402
rect 54 -405 94 -404
rect 121 -405 150 -404
rect 170 -405 304 -404
rect 373 -405 381 -404
rect 47 -407 122 -406
rect 128 -407 157 -406
rect 170 -407 178 -406
rect 254 -407 276 -406
rect 58 -409 178 -408
rect 264 -409 381 -408
rect 117 -411 255 -410
rect 9 -422 52 -421
rect 79 -422 83 -421
rect 107 -422 216 -421
rect 226 -422 346 -421
rect 432 -422 458 -421
rect 16 -424 34 -423
rect 44 -424 143 -423
rect 166 -424 171 -423
rect 194 -424 213 -423
rect 229 -424 290 -423
rect 317 -424 346 -423
rect 359 -424 433 -423
rect 443 -424 451 -423
rect 16 -426 27 -425
rect 30 -426 76 -425
rect 79 -426 87 -425
rect 93 -426 108 -425
rect 121 -426 143 -425
rect 163 -426 290 -425
rect 327 -426 423 -425
rect 446 -426 465 -425
rect 51 -428 73 -427
rect 86 -428 101 -427
rect 121 -428 136 -427
rect 156 -428 164 -427
rect 177 -428 318 -427
rect 334 -428 402 -427
rect 58 -430 73 -429
rect 82 -430 101 -429
rect 114 -430 178 -429
rect 201 -430 339 -429
rect 352 -430 360 -429
rect 93 -432 181 -431
rect 212 -432 234 -431
rect 236 -432 339 -431
rect 128 -434 220 -433
rect 240 -434 423 -433
rect 117 -436 129 -435
rect 131 -436 150 -435
rect 156 -436 192 -435
rect 243 -436 304 -435
rect 135 -438 185 -437
rect 191 -438 437 -437
rect 149 -440 199 -439
rect 247 -440 297 -439
rect 387 -440 437 -439
rect 226 -442 297 -441
rect 387 -442 409 -441
rect 250 -444 395 -443
rect 250 -446 416 -445
rect 254 -448 304 -447
rect 310 -448 416 -447
rect 254 -450 353 -449
rect 373 -450 395 -449
rect 257 -452 367 -451
rect 373 -452 381 -451
rect 261 -454 332 -453
rect 170 -456 262 -455
rect 268 -456 381 -455
rect 65 -458 269 -457
rect 275 -458 311 -457
rect 324 -458 367 -457
rect 47 -460 276 -459
rect 282 -460 325 -459
rect 65 -462 206 -461
rect 184 -464 283 -463
rect 205 -466 223 -465
rect 9 -477 125 -476
rect 142 -477 234 -476
rect 247 -477 255 -476
rect 261 -477 318 -476
rect 352 -477 402 -476
rect 418 -477 451 -476
rect 30 -479 237 -478
rect 250 -479 339 -478
rect 345 -479 353 -478
rect 387 -479 409 -478
rect 422 -479 447 -478
rect 33 -481 216 -480
rect 222 -481 416 -480
rect 432 -481 437 -480
rect 37 -483 129 -482
rect 131 -483 346 -482
rect 380 -483 388 -482
rect 415 -483 451 -482
rect 16 -485 38 -484
rect 40 -485 59 -484
rect 72 -485 94 -484
rect 100 -485 143 -484
rect 173 -485 199 -484
rect 205 -485 262 -484
rect 264 -485 311 -484
rect 359 -485 381 -484
rect 16 -487 24 -486
rect 44 -487 139 -486
rect 180 -487 430 -486
rect 51 -489 104 -488
rect 107 -489 227 -488
rect 240 -489 437 -488
rect 51 -491 73 -490
rect 82 -491 178 -490
rect 191 -491 220 -490
rect 275 -491 283 -490
rect 285 -491 395 -490
rect 429 -491 458 -490
rect 58 -493 80 -492
rect 93 -493 111 -492
rect 128 -493 136 -492
rect 184 -493 192 -492
rect 212 -493 248 -492
rect 296 -493 318 -492
rect 359 -493 367 -492
rect 443 -493 458 -492
rect 79 -495 332 -494
rect 107 -497 122 -496
rect 156 -497 185 -496
rect 268 -497 332 -496
rect 121 -499 164 -498
rect 170 -499 269 -498
rect 289 -499 297 -498
rect 303 -499 339 -498
rect 65 -501 290 -500
rect 310 -501 325 -500
rect 65 -503 87 -502
rect 156 -503 195 -502
rect 243 -503 325 -502
rect 86 -505 150 -504
rect 163 -505 304 -504
rect 149 -507 206 -506
rect 9 -518 69 -517
rect 72 -518 94 -517
rect 117 -518 125 -517
rect 138 -518 437 -517
rect 9 -520 104 -519
rect 121 -520 227 -519
rect 243 -520 255 -519
rect 278 -520 353 -519
rect 366 -520 423 -519
rect 429 -520 444 -519
rect 16 -522 38 -521
rect 44 -522 206 -521
rect 208 -522 339 -521
rect 401 -522 416 -521
rect 443 -522 458 -521
rect 19 -524 276 -523
rect 285 -524 381 -523
rect 457 -524 465 -523
rect 37 -526 157 -525
rect 166 -526 255 -525
rect 303 -526 409 -525
rect 450 -526 465 -525
rect 44 -528 52 -527
rect 58 -528 97 -527
rect 124 -528 174 -527
rect 184 -528 206 -527
rect 212 -528 332 -527
rect 359 -528 381 -527
rect 30 -530 59 -529
rect 72 -530 171 -529
rect 173 -530 437 -529
rect 30 -532 94 -531
rect 149 -532 188 -531
rect 212 -532 269 -531
rect 306 -532 342 -531
rect 373 -532 416 -531
rect 26 -534 269 -533
rect 310 -534 353 -533
rect 373 -534 433 -533
rect 51 -536 66 -535
rect 82 -536 367 -535
rect 40 -538 66 -537
rect 82 -538 283 -537
rect 324 -538 395 -537
rect 86 -540 157 -539
rect 184 -540 360 -539
rect 86 -542 108 -541
rect 149 -542 164 -541
rect 198 -542 311 -541
rect 331 -542 346 -541
rect 107 -544 129 -543
rect 163 -544 178 -543
rect 219 -544 227 -543
rect 233 -544 409 -543
rect 103 -546 129 -545
rect 135 -546 178 -545
rect 191 -546 220 -545
rect 233 -546 388 -545
rect 114 -548 199 -547
rect 240 -548 388 -547
rect 191 -550 216 -549
rect 247 -550 276 -549
rect 282 -550 402 -549
rect 247 -552 262 -551
rect 296 -552 325 -551
rect 23 -554 297 -553
rect 317 -554 346 -553
rect 236 -556 262 -555
rect 289 -556 318 -555
rect 142 -558 290 -557
rect 114 -560 143 -559
rect 9 -571 185 -570
rect 212 -571 265 -570
rect 303 -571 346 -570
rect 464 -571 472 -570
rect 16 -573 101 -572
rect 138 -573 304 -572
rect 341 -573 395 -572
rect 457 -573 465 -572
rect 16 -575 115 -574
rect 163 -575 447 -574
rect 23 -577 129 -576
rect 163 -577 209 -576
rect 233 -577 248 -576
rect 257 -577 402 -576
rect 9 -579 209 -578
rect 236 -579 367 -578
rect 394 -579 430 -578
rect 30 -581 104 -580
rect 170 -581 283 -580
rect 33 -583 45 -582
rect 58 -583 90 -582
rect 93 -583 244 -582
rect 247 -583 318 -582
rect 40 -585 430 -584
rect 44 -587 52 -586
rect 58 -587 108 -586
rect 149 -587 283 -586
rect 317 -587 332 -586
rect 37 -589 52 -588
rect 65 -589 157 -588
rect 173 -589 220 -588
rect 240 -589 353 -588
rect 68 -591 346 -590
rect 352 -591 360 -590
rect 79 -593 290 -592
rect 331 -593 367 -592
rect 72 -595 80 -594
rect 93 -595 437 -594
rect 30 -597 437 -596
rect 72 -599 87 -598
rect 107 -599 195 -598
rect 205 -599 234 -598
rect 240 -599 269 -598
rect 289 -599 325 -598
rect 359 -599 381 -598
rect 86 -601 143 -600
rect 156 -601 174 -600
rect 177 -601 192 -600
rect 219 -601 276 -600
rect 306 -601 381 -600
rect 135 -603 150 -602
rect 180 -603 409 -602
rect 142 -605 171 -604
rect 254 -605 402 -604
rect 268 -607 311 -606
rect 338 -607 409 -606
rect 261 -609 311 -608
rect 338 -609 374 -608
rect 275 -611 297 -610
rect 373 -611 388 -610
rect 296 -613 325 -612
rect 387 -613 454 -612
rect 2 -624 52 -623
rect 72 -624 115 -623
rect 117 -624 213 -623
rect 222 -624 269 -623
rect 299 -624 423 -623
rect 436 -624 444 -623
rect 450 -624 458 -623
rect 460 -624 465 -623
rect 9 -626 104 -625
rect 170 -626 185 -625
rect 187 -626 283 -625
rect 299 -626 416 -625
rect 429 -626 437 -625
rect 9 -628 76 -627
rect 79 -628 132 -627
rect 142 -628 171 -627
rect 191 -628 216 -627
rect 233 -628 423 -627
rect 23 -630 136 -629
rect 142 -630 227 -629
rect 240 -630 255 -629
rect 261 -630 353 -629
rect 380 -630 430 -629
rect 16 -632 24 -631
rect 30 -632 164 -631
rect 194 -632 402 -631
rect 415 -632 447 -631
rect 16 -634 66 -633
rect 93 -634 97 -633
rect 128 -634 195 -633
rect 205 -634 304 -633
rect 331 -634 360 -633
rect 33 -636 66 -635
rect 86 -636 129 -635
rect 135 -636 150 -635
rect 208 -636 388 -635
rect 37 -638 199 -637
rect 215 -638 283 -637
rect 289 -638 304 -637
rect 331 -638 353 -637
rect 387 -638 395 -637
rect 37 -640 178 -639
rect 180 -640 395 -639
rect 40 -642 272 -641
rect 334 -642 409 -641
rect 44 -644 52 -643
rect 54 -644 451 -643
rect 44 -646 276 -645
rect 345 -646 381 -645
rect 58 -648 80 -647
rect 93 -648 122 -647
rect 156 -648 199 -647
rect 219 -648 234 -647
rect 243 -648 360 -647
rect 366 -648 409 -647
rect 58 -650 90 -649
rect 96 -650 122 -649
rect 163 -650 209 -649
rect 226 -650 248 -649
rect 254 -650 458 -649
rect 107 -652 150 -651
rect 184 -652 290 -651
rect 324 -652 367 -651
rect 100 -654 108 -653
rect 114 -654 178 -653
rect 240 -654 325 -653
rect 338 -654 346 -653
rect 100 -656 157 -655
rect 261 -656 318 -655
rect 103 -658 339 -657
rect 250 -660 318 -659
rect 250 -662 402 -661
rect 275 -664 297 -663
rect 2 -675 132 -674
rect 135 -675 181 -674
rect 187 -675 220 -674
rect 233 -675 241 -674
rect 250 -675 304 -674
rect 331 -675 339 -674
rect 443 -675 458 -674
rect 464 -675 472 -674
rect 16 -677 101 -676
rect 114 -677 150 -676
rect 170 -677 174 -676
rect 191 -677 318 -676
rect 334 -677 430 -676
rect 9 -679 17 -678
rect 37 -679 178 -678
rect 191 -679 227 -678
rect 250 -679 437 -678
rect 9 -681 94 -680
rect 128 -681 402 -680
rect 23 -683 94 -682
rect 149 -683 241 -682
rect 268 -683 318 -682
rect 380 -683 430 -682
rect 23 -685 290 -684
rect 296 -685 367 -684
rect 380 -685 409 -684
rect 37 -687 206 -686
rect 212 -687 423 -686
rect 40 -689 132 -688
rect 170 -689 213 -688
rect 229 -689 290 -688
rect 299 -689 346 -688
rect 359 -689 367 -688
rect 401 -689 416 -688
rect 44 -691 87 -690
rect 177 -691 283 -690
rect 345 -691 353 -690
rect 359 -691 374 -690
rect 51 -693 353 -692
rect 58 -695 136 -694
rect 194 -695 220 -694
rect 268 -695 311 -694
rect 58 -697 255 -696
rect 261 -697 311 -696
rect 72 -699 101 -698
rect 198 -699 216 -698
rect 254 -699 276 -698
rect 282 -699 325 -698
rect 2 -701 73 -700
rect 75 -701 185 -700
rect 261 -701 374 -700
rect 79 -703 115 -702
rect 142 -703 199 -702
rect 324 -703 395 -702
rect 82 -705 108 -704
rect 142 -705 157 -704
rect 184 -705 234 -704
rect 394 -705 451 -704
rect 65 -707 108 -706
rect 156 -707 164 -706
rect 54 -709 66 -708
rect 86 -709 125 -708
rect 121 -711 164 -710
rect 30 -713 122 -712
rect 30 -715 118 -714
rect 9 -726 73 -725
rect 96 -726 185 -725
rect 198 -726 353 -725
rect 376 -726 402 -725
rect 411 -726 430 -725
rect 16 -728 76 -727
rect 110 -728 251 -727
rect 254 -728 279 -727
rect 289 -728 297 -727
rect 338 -728 381 -727
rect 387 -728 409 -727
rect 23 -730 199 -729
rect 215 -730 234 -729
rect 243 -730 311 -729
rect 341 -730 346 -729
rect 2 -732 311 -731
rect 345 -732 360 -731
rect 23 -734 87 -733
rect 121 -734 304 -733
rect 37 -736 80 -735
rect 86 -736 192 -735
rect 233 -736 269 -735
rect 289 -736 325 -735
rect 37 -738 181 -737
rect 205 -738 269 -737
rect 324 -738 395 -737
rect 40 -740 59 -739
rect 65 -740 76 -739
rect 128 -740 255 -739
rect 16 -742 59 -741
rect 114 -742 129 -741
rect 135 -742 185 -741
rect 247 -742 283 -741
rect 44 -744 192 -743
rect 236 -744 283 -743
rect 44 -746 66 -745
rect 93 -746 136 -745
rect 142 -746 209 -745
rect 51 -748 83 -747
rect 100 -748 143 -747
rect 156 -748 202 -747
rect 54 -750 241 -749
rect 82 -752 115 -751
rect 163 -752 171 -751
rect 180 -752 318 -751
rect 100 -754 262 -753
rect 30 -756 262 -755
rect 103 -758 209 -757
rect 107 -760 157 -759
rect 163 -760 227 -759
rect 219 -762 227 -761
rect 212 -764 220 -763
rect 212 -766 332 -765
rect 331 -768 367 -767
rect 9 -779 48 -778
rect 58 -779 108 -778
rect 110 -779 157 -778
rect 177 -779 304 -778
rect 317 -779 339 -778
rect 30 -781 52 -780
rect 65 -781 76 -780
rect 93 -781 143 -780
rect 177 -781 227 -780
rect 233 -781 262 -780
rect 51 -783 80 -782
rect 96 -783 255 -782
rect 72 -785 83 -784
rect 100 -785 153 -784
rect 163 -785 262 -784
rect 103 -787 304 -786
rect 107 -789 241 -788
rect 247 -789 276 -788
rect 30 -791 248 -790
rect 254 -791 283 -790
rect 117 -793 171 -792
rect 205 -793 213 -792
rect 219 -793 227 -792
rect 282 -793 290 -792
rect 23 -795 171 -794
rect 212 -795 237 -794
rect 23 -797 62 -796
rect 124 -797 136 -796
rect 163 -797 192 -796
rect 33 -799 136 -798
rect 149 -799 192 -798
rect 33 -801 118 -800
rect 124 -801 185 -800
rect 37 -803 290 -802
rect 37 -805 115 -804
rect 128 -805 157 -804
rect 86 -807 185 -806
rect 131 -809 311 -808
rect 310 -811 325 -810
rect 324 -813 346 -812
rect 9 -824 17 -823
rect 23 -824 66 -823
rect 72 -824 94 -823
rect 96 -824 234 -823
rect 240 -824 269 -823
rect 292 -824 318 -823
rect 324 -824 346 -823
rect 23 -826 262 -825
rect 310 -826 328 -825
rect 33 -828 48 -827
rect 58 -828 80 -827
rect 86 -828 115 -827
rect 117 -828 192 -827
rect 222 -828 227 -827
rect 254 -828 269 -827
rect 37 -830 90 -829
rect 117 -830 290 -829
rect 33 -832 38 -831
rect 72 -832 101 -831
rect 124 -832 164 -831
rect 191 -832 248 -831
rect 51 -834 164 -833
rect 212 -834 227 -833
rect 44 -836 52 -835
rect 128 -836 157 -835
rect 205 -836 213 -835
rect 19 -838 45 -837
rect 135 -838 181 -837
rect 135 -840 146 -839
rect 149 -840 199 -839
rect 152 -842 304 -841
rect 156 -844 171 -843
rect 170 -846 290 -845
rect 23 -857 143 -856
rect 187 -857 192 -856
rect 268 -857 286 -856
rect 37 -859 45 -858
rect 47 -859 59 -858
rect 65 -859 87 -858
rect 93 -859 115 -858
rect 131 -859 150 -858
rect 54 -861 171 -860
rect 72 -863 104 -862
rect 107 -863 157 -862
rect 82 -865 164 -864
<< m2contact >>
rect 12 0 13 1
rect 26 0 27 1
rect 37 0 38 1
rect 65 0 66 1
rect 93 0 94 1
rect 107 0 108 1
rect 121 0 122 1
rect 128 0 129 1
rect 135 0 136 1
rect 163 0 164 1
rect 51 -2 52 -1
rect 89 -2 90 -1
rect 138 -2 139 -1
rect 149 -2 150 -1
rect 58 -4 59 -3
rect 72 -4 73 -3
rect 72 -15 73 -14
rect 96 -15 97 -14
rect 100 -15 101 -14
rect 107 -15 108 -14
rect 114 -15 115 -14
rect 156 -15 157 -14
rect 159 -15 160 -14
rect 191 -15 192 -14
rect 65 -17 66 -16
rect 72 -17 73 -16
rect 79 -17 80 -16
rect 100 -17 101 -16
rect 107 -17 108 -16
rect 142 -17 143 -16
rect 145 -17 146 -16
rect 149 -17 150 -16
rect 163 -17 164 -16
rect 173 -17 174 -16
rect 114 -19 115 -18
rect 177 -19 178 -18
rect 149 -21 150 -20
rect 201 -21 202 -20
rect 163 -23 164 -22
rect 187 -23 188 -22
rect 47 -34 48 -33
rect 212 -34 213 -33
rect 51 -36 52 -35
rect 149 -36 150 -35
rect 163 -36 164 -35
rect 219 -36 220 -35
rect 58 -38 59 -37
rect 72 -38 73 -37
rect 86 -38 87 -37
rect 163 -38 164 -37
rect 177 -38 178 -37
rect 233 -38 234 -37
rect 16 -40 17 -39
rect 177 -40 178 -39
rect 191 -40 192 -39
rect 254 -40 255 -39
rect 65 -42 66 -41
rect 117 -42 118 -41
rect 121 -42 122 -41
rect 170 -42 171 -41
rect 198 -42 199 -41
rect 247 -42 248 -41
rect 72 -44 73 -43
rect 79 -44 80 -43
rect 93 -44 94 -43
rect 184 -44 185 -43
rect 37 -46 38 -45
rect 93 -46 94 -45
rect 96 -46 97 -45
rect 198 -46 199 -45
rect 124 -48 125 -47
rect 152 -48 153 -47
rect 100 -50 101 -49
rect 124 -50 125 -49
rect 142 -50 143 -49
rect 226 -50 227 -49
rect 145 -52 146 -51
rect 156 -52 157 -51
rect 149 -54 150 -53
rect 205 -54 206 -53
rect 19 -65 20 -64
rect 212 -65 213 -64
rect 219 -65 220 -64
rect 275 -65 276 -64
rect 40 -67 41 -66
rect 79 -67 80 -66
rect 82 -67 83 -66
rect 110 -67 111 -66
rect 121 -67 122 -66
rect 159 -67 160 -66
rect 177 -67 178 -66
rect 219 -67 220 -66
rect 226 -67 227 -66
rect 331 -67 332 -66
rect 40 -69 41 -68
rect 177 -69 178 -68
rect 191 -69 192 -68
rect 254 -69 255 -68
rect 44 -71 45 -70
rect 51 -71 52 -70
rect 58 -71 59 -70
rect 89 -71 90 -70
rect 100 -71 101 -70
rect 128 -71 129 -70
rect 131 -71 132 -70
rect 261 -71 262 -70
rect 30 -73 31 -72
rect 131 -73 132 -72
rect 138 -73 139 -72
rect 142 -73 143 -72
rect 149 -73 150 -72
rect 212 -73 213 -72
rect 233 -73 234 -72
rect 282 -73 283 -72
rect 30 -75 31 -74
rect 114 -75 115 -74
rect 163 -75 164 -74
rect 226 -75 227 -74
rect 243 -75 244 -74
rect 254 -75 255 -74
rect 51 -77 52 -76
rect 96 -77 97 -76
rect 107 -77 108 -76
rect 135 -77 136 -76
rect 184 -77 185 -76
rect 191 -77 192 -76
rect 205 -77 206 -76
rect 240 -77 241 -76
rect 247 -77 248 -76
rect 268 -77 269 -76
rect 58 -79 59 -78
rect 65 -79 66 -78
rect 86 -79 87 -78
rect 156 -79 157 -78
rect 170 -79 171 -78
rect 205 -79 206 -78
rect 65 -81 66 -80
rect 72 -81 73 -80
rect 110 -81 111 -80
rect 296 -81 297 -80
rect 72 -83 73 -82
rect 100 -83 101 -82
rect 170 -83 171 -82
rect 289 -83 290 -82
rect 184 -85 185 -84
rect 233 -85 234 -84
rect 198 -87 199 -86
rect 247 -87 248 -86
rect 23 -98 24 -97
rect 86 -98 87 -97
rect 93 -98 94 -97
rect 131 -98 132 -97
rect 135 -98 136 -97
rect 226 -98 227 -97
rect 268 -98 269 -97
rect 359 -98 360 -97
rect 26 -100 27 -99
rect 352 -100 353 -99
rect 30 -102 31 -101
rect 198 -102 199 -101
rect 201 -102 202 -101
rect 317 -102 318 -101
rect 51 -104 52 -103
rect 100 -104 101 -103
rect 107 -104 108 -103
rect 117 -104 118 -103
rect 121 -104 122 -103
rect 142 -104 143 -103
rect 145 -104 146 -103
rect 310 -104 311 -103
rect 51 -106 52 -105
rect 65 -106 66 -105
rect 96 -106 97 -105
rect 261 -106 262 -105
rect 271 -106 272 -105
rect 366 -106 367 -105
rect 65 -108 66 -107
rect 173 -108 174 -107
rect 194 -108 195 -107
rect 226 -108 227 -107
rect 254 -108 255 -107
rect 261 -108 262 -107
rect 275 -108 276 -107
rect 345 -108 346 -107
rect 30 -110 31 -109
rect 275 -110 276 -109
rect 289 -110 290 -109
rect 373 -110 374 -109
rect 86 -112 87 -111
rect 254 -112 255 -111
rect 303 -112 304 -111
rect 324 -112 325 -111
rect 128 -114 129 -113
rect 247 -114 248 -113
rect 138 -116 139 -115
rect 303 -116 304 -115
rect 138 -118 139 -117
rect 201 -118 202 -117
rect 233 -118 234 -117
rect 289 -118 290 -117
rect 149 -120 150 -119
rect 205 -120 206 -119
rect 233 -120 234 -119
rect 296 -120 297 -119
rect 149 -122 150 -121
rect 208 -122 209 -121
rect 240 -122 241 -121
rect 296 -122 297 -121
rect 152 -124 153 -123
rect 170 -124 171 -123
rect 191 -124 192 -123
rect 247 -124 248 -123
rect 156 -126 157 -125
rect 338 -126 339 -125
rect 44 -128 45 -127
rect 156 -128 157 -127
rect 163 -128 164 -127
rect 282 -128 283 -127
rect 9 -130 10 -129
rect 44 -130 45 -129
rect 124 -130 125 -129
rect 163 -130 164 -129
rect 166 -130 167 -129
rect 219 -130 220 -129
rect 37 -132 38 -131
rect 282 -132 283 -131
rect 166 -134 167 -133
rect 184 -134 185 -133
rect 212 -134 213 -133
rect 240 -134 241 -133
rect 128 -136 129 -135
rect 212 -136 213 -135
rect 177 -138 178 -137
rect 219 -138 220 -137
rect 72 -140 73 -139
rect 177 -140 178 -139
rect 72 -142 73 -141
rect 121 -142 122 -141
rect 5 -153 6 -152
rect 19 -153 20 -152
rect 23 -153 24 -152
rect 310 -153 311 -152
rect 345 -153 346 -152
rect 380 -153 381 -152
rect 9 -155 10 -154
rect 26 -155 27 -154
rect 61 -155 62 -154
rect 338 -155 339 -154
rect 345 -155 346 -154
rect 352 -155 353 -154
rect 373 -155 374 -154
rect 401 -155 402 -154
rect 16 -157 17 -156
rect 37 -157 38 -156
rect 65 -157 66 -156
rect 103 -157 104 -156
rect 128 -157 129 -156
rect 289 -157 290 -156
rect 338 -157 339 -156
rect 366 -157 367 -156
rect 16 -159 17 -158
rect 51 -159 52 -158
rect 86 -159 87 -158
rect 303 -159 304 -158
rect 320 -159 321 -158
rect 366 -159 367 -158
rect 23 -161 24 -160
rect 30 -161 31 -160
rect 37 -161 38 -160
rect 107 -161 108 -160
rect 128 -161 129 -160
rect 198 -161 199 -160
rect 208 -161 209 -160
rect 359 -161 360 -160
rect 30 -163 31 -162
rect 173 -163 174 -162
rect 191 -163 192 -162
rect 373 -163 374 -162
rect 51 -165 52 -164
rect 96 -165 97 -164
rect 107 -165 108 -164
rect 205 -165 206 -164
rect 222 -165 223 -164
rect 387 -165 388 -164
rect 79 -167 80 -166
rect 205 -167 206 -166
rect 226 -167 227 -166
rect 303 -167 304 -166
rect 359 -167 360 -166
rect 408 -167 409 -166
rect 65 -169 66 -168
rect 79 -169 80 -168
rect 86 -169 87 -168
rect 93 -169 94 -168
rect 149 -169 150 -168
rect 184 -169 185 -168
rect 194 -169 195 -168
rect 296 -169 297 -168
rect 89 -171 90 -170
rect 142 -171 143 -170
rect 149 -171 150 -170
rect 296 -171 297 -170
rect 72 -173 73 -172
rect 142 -173 143 -172
rect 152 -173 153 -172
rect 247 -173 248 -172
rect 261 -173 262 -172
rect 415 -173 416 -172
rect 47 -175 48 -174
rect 72 -175 73 -174
rect 156 -175 157 -174
rect 184 -175 185 -174
rect 198 -175 199 -174
rect 310 -175 311 -174
rect 100 -177 101 -176
rect 156 -177 157 -176
rect 163 -177 164 -176
rect 240 -177 241 -176
rect 261 -177 262 -176
rect 282 -177 283 -176
rect 75 -179 76 -178
rect 163 -179 164 -178
rect 166 -179 167 -178
rect 394 -179 395 -178
rect 82 -181 83 -180
rect 240 -181 241 -180
rect 254 -181 255 -180
rect 282 -181 283 -180
rect 82 -183 83 -182
rect 121 -183 122 -182
rect 177 -183 178 -182
rect 191 -183 192 -182
rect 208 -183 209 -182
rect 226 -183 227 -182
rect 233 -183 234 -182
rect 247 -183 248 -182
rect 268 -183 269 -182
rect 317 -183 318 -182
rect 100 -185 101 -184
rect 135 -185 136 -184
rect 152 -185 153 -184
rect 268 -185 269 -184
rect 275 -185 276 -184
rect 289 -185 290 -184
rect 61 -187 62 -186
rect 275 -187 276 -186
rect 114 -189 115 -188
rect 121 -189 122 -188
rect 170 -189 171 -188
rect 177 -189 178 -188
rect 212 -189 213 -188
rect 233 -189 234 -188
rect 44 -191 45 -190
rect 114 -191 115 -190
rect 219 -191 220 -190
rect 254 -191 255 -190
rect 58 -193 59 -192
rect 212 -193 213 -192
rect 219 -193 220 -192
rect 352 -193 353 -192
rect 16 -204 17 -203
rect 72 -204 73 -203
rect 86 -204 87 -203
rect 149 -204 150 -203
rect 166 -204 167 -203
rect 303 -204 304 -203
rect 16 -206 17 -205
rect 180 -206 181 -205
rect 184 -206 185 -205
rect 387 -206 388 -205
rect 23 -208 24 -207
rect 107 -208 108 -207
rect 110 -208 111 -207
rect 198 -208 199 -207
rect 205 -208 206 -207
rect 373 -208 374 -207
rect 44 -210 45 -209
rect 114 -210 115 -209
rect 117 -210 118 -209
rect 275 -210 276 -209
rect 338 -210 339 -209
rect 373 -210 374 -209
rect 44 -212 45 -211
rect 100 -212 101 -211
rect 107 -212 108 -211
rect 303 -212 304 -211
rect 338 -212 339 -211
rect 345 -212 346 -211
rect 54 -214 55 -213
rect 198 -214 199 -213
rect 219 -214 220 -213
rect 415 -214 416 -213
rect 65 -216 66 -215
rect 82 -216 83 -215
rect 86 -216 87 -215
rect 114 -216 115 -215
rect 124 -216 125 -215
rect 128 -216 129 -215
rect 138 -216 139 -215
rect 191 -216 192 -215
rect 240 -216 241 -215
rect 387 -216 388 -215
rect 30 -218 31 -217
rect 128 -218 129 -217
rect 142 -218 143 -217
rect 163 -218 164 -217
rect 170 -218 171 -217
rect 233 -218 234 -217
rect 275 -218 276 -217
rect 289 -218 290 -217
rect 310 -218 311 -217
rect 415 -218 416 -217
rect 9 -220 10 -219
rect 30 -220 31 -219
rect 37 -220 38 -219
rect 142 -220 143 -219
rect 177 -220 178 -219
rect 233 -220 234 -219
rect 289 -220 290 -219
rect 296 -220 297 -219
rect 345 -220 346 -219
rect 352 -220 353 -219
rect 9 -222 10 -221
rect 75 -222 76 -221
rect 93 -222 94 -221
rect 156 -222 157 -221
rect 187 -222 188 -221
rect 317 -222 318 -221
rect 352 -222 353 -221
rect 359 -222 360 -221
rect 37 -224 38 -223
rect 82 -224 83 -223
rect 96 -224 97 -223
rect 394 -224 395 -223
rect 65 -226 66 -225
rect 79 -226 80 -225
rect 121 -226 122 -225
rect 156 -226 157 -225
rect 187 -226 188 -225
rect 205 -226 206 -225
rect 222 -226 223 -225
rect 240 -226 241 -225
rect 261 -226 262 -225
rect 296 -226 297 -225
rect 359 -226 360 -225
rect 366 -226 367 -225
rect 51 -228 52 -227
rect 222 -228 223 -227
rect 121 -230 122 -229
rect 366 -230 367 -229
rect 135 -232 136 -231
rect 394 -232 395 -231
rect 149 -234 150 -233
rect 177 -234 178 -233
rect 191 -234 192 -233
rect 212 -234 213 -233
rect 201 -236 202 -235
rect 261 -236 262 -235
rect 201 -238 202 -237
rect 380 -238 381 -237
rect 58 -240 59 -239
rect 380 -240 381 -239
rect 58 -242 59 -241
rect 226 -242 227 -241
rect 212 -244 213 -243
rect 254 -244 255 -243
rect 226 -246 227 -245
rect 268 -246 269 -245
rect 254 -248 255 -247
rect 408 -248 409 -247
rect 268 -250 269 -249
rect 282 -250 283 -249
rect 282 -252 283 -251
rect 310 -252 311 -251
rect 12 -263 13 -262
rect 338 -263 339 -262
rect 380 -263 381 -262
rect 436 -263 437 -262
rect 33 -265 34 -264
rect 54 -265 55 -264
rect 61 -265 62 -264
rect 65 -265 66 -264
rect 72 -265 73 -264
rect 107 -265 108 -264
rect 110 -265 111 -264
rect 268 -265 269 -264
rect 282 -265 283 -264
rect 432 -265 433 -264
rect 37 -267 38 -266
rect 65 -267 66 -266
rect 75 -267 76 -266
rect 138 -267 139 -266
rect 163 -267 164 -266
rect 184 -267 185 -266
rect 226 -267 227 -266
rect 422 -267 423 -266
rect 30 -269 31 -268
rect 163 -269 164 -268
rect 173 -269 174 -268
rect 212 -269 213 -268
rect 240 -269 241 -268
rect 289 -269 290 -268
rect 338 -269 339 -268
rect 345 -269 346 -268
rect 380 -269 381 -268
rect 425 -269 426 -268
rect 37 -271 38 -270
rect 58 -271 59 -270
rect 86 -271 87 -270
rect 114 -271 115 -270
rect 117 -271 118 -270
rect 142 -271 143 -270
rect 177 -271 178 -270
rect 201 -271 202 -270
rect 205 -271 206 -270
rect 226 -271 227 -270
rect 247 -271 248 -270
rect 254 -271 255 -270
rect 268 -271 269 -270
rect 317 -271 318 -270
rect 345 -271 346 -270
rect 373 -271 374 -270
rect 394 -271 395 -270
rect 397 -271 398 -270
rect 51 -273 52 -272
rect 198 -273 199 -272
rect 212 -273 213 -272
rect 296 -273 297 -272
rect 317 -273 318 -272
rect 331 -273 332 -272
rect 366 -273 367 -272
rect 373 -273 374 -272
rect 394 -273 395 -272
rect 415 -273 416 -272
rect 79 -275 80 -274
rect 86 -275 87 -274
rect 96 -275 97 -274
rect 289 -275 290 -274
rect 331 -275 332 -274
rect 352 -275 353 -274
rect 359 -275 360 -274
rect 366 -275 367 -274
rect 401 -275 402 -274
rect 415 -275 416 -274
rect 23 -277 24 -276
rect 79 -277 80 -276
rect 100 -277 101 -276
rect 142 -277 143 -276
rect 180 -277 181 -276
rect 233 -277 234 -276
rect 250 -277 251 -276
rect 387 -277 388 -276
rect 401 -277 402 -276
rect 408 -277 409 -276
rect 23 -279 24 -278
rect 44 -279 45 -278
rect 100 -279 101 -278
rect 156 -279 157 -278
rect 184 -279 185 -278
rect 275 -279 276 -278
rect 397 -279 398 -278
rect 408 -279 409 -278
rect 44 -281 45 -280
rect 201 -281 202 -280
rect 205 -281 206 -280
rect 352 -281 353 -280
rect 103 -283 104 -282
rect 170 -283 171 -282
rect 198 -283 199 -282
rect 296 -283 297 -282
rect 128 -285 129 -284
rect 240 -285 241 -284
rect 254 -285 255 -284
rect 261 -285 262 -284
rect 275 -285 276 -284
rect 310 -285 311 -284
rect 16 -287 17 -286
rect 261 -287 262 -286
rect 264 -287 265 -286
rect 310 -287 311 -286
rect 16 -289 17 -288
rect 243 -289 244 -288
rect 128 -291 129 -290
rect 170 -291 171 -290
rect 219 -291 220 -290
rect 247 -291 248 -290
rect 135 -293 136 -292
rect 387 -293 388 -292
rect 93 -295 94 -294
rect 135 -295 136 -294
rect 156 -295 157 -294
rect 191 -295 192 -294
rect 222 -295 223 -294
rect 359 -295 360 -294
rect 166 -297 167 -296
rect 191 -297 192 -296
rect 233 -297 234 -296
rect 303 -297 304 -296
rect 303 -299 304 -298
rect 324 -299 325 -298
rect 124 -301 125 -300
rect 324 -301 325 -300
rect 2 -312 3 -311
rect 173 -312 174 -311
rect 184 -312 185 -311
rect 240 -312 241 -311
rect 243 -312 244 -311
rect 338 -312 339 -311
rect 401 -312 402 -311
rect 429 -312 430 -311
rect 23 -314 24 -313
rect 93 -314 94 -313
rect 100 -314 101 -313
rect 128 -314 129 -313
rect 142 -314 143 -313
rect 205 -314 206 -313
rect 233 -314 234 -313
rect 261 -314 262 -313
rect 264 -314 265 -313
rect 415 -314 416 -313
rect 26 -316 27 -315
rect 103 -316 104 -315
rect 107 -316 108 -315
rect 415 -316 416 -315
rect 30 -318 31 -317
rect 187 -318 188 -317
rect 191 -318 192 -317
rect 222 -318 223 -317
rect 247 -318 248 -317
rect 254 -318 255 -317
rect 317 -318 318 -317
rect 338 -318 339 -317
rect 23 -320 24 -319
rect 191 -320 192 -319
rect 198 -320 199 -319
rect 303 -320 304 -319
rect 317 -320 318 -319
rect 324 -320 325 -319
rect 30 -322 31 -321
rect 373 -322 374 -321
rect 37 -324 38 -323
rect 170 -324 171 -323
rect 198 -324 199 -323
rect 219 -324 220 -323
rect 250 -324 251 -323
rect 380 -324 381 -323
rect 33 -326 34 -325
rect 37 -326 38 -325
rect 40 -326 41 -325
rect 401 -326 402 -325
rect 44 -328 45 -327
rect 124 -328 125 -327
rect 142 -328 143 -327
rect 212 -328 213 -327
rect 254 -328 255 -327
rect 422 -328 423 -327
rect 54 -330 55 -329
rect 303 -330 304 -329
rect 345 -330 346 -329
rect 380 -330 381 -329
rect 58 -332 59 -331
rect 86 -332 87 -331
rect 110 -332 111 -331
rect 128 -332 129 -331
rect 159 -332 160 -331
rect 177 -332 178 -331
rect 296 -332 297 -331
rect 324 -332 325 -331
rect 373 -332 374 -331
rect 387 -332 388 -331
rect 61 -334 62 -333
rect 93 -334 94 -333
rect 110 -334 111 -333
rect 345 -334 346 -333
rect 65 -336 66 -335
rect 205 -336 206 -335
rect 233 -336 234 -335
rect 387 -336 388 -335
rect 65 -338 66 -337
rect 296 -338 297 -337
rect 72 -340 73 -339
rect 436 -340 437 -339
rect 79 -342 80 -341
rect 163 -342 164 -341
rect 394 -342 395 -341
rect 436 -342 437 -341
rect 16 -344 17 -343
rect 79 -344 80 -343
rect 114 -344 115 -343
rect 212 -344 213 -343
rect 366 -344 367 -343
rect 394 -344 395 -343
rect 16 -346 17 -345
rect 68 -346 69 -345
rect 121 -346 122 -345
rect 149 -346 150 -345
rect 359 -346 360 -345
rect 366 -346 367 -345
rect 117 -348 118 -347
rect 121 -348 122 -347
rect 135 -348 136 -347
rect 177 -348 178 -347
rect 352 -348 353 -347
rect 359 -348 360 -347
rect 117 -350 118 -349
rect 408 -350 409 -349
rect 51 -352 52 -351
rect 408 -352 409 -351
rect 51 -354 52 -353
rect 149 -354 150 -353
rect 289 -354 290 -353
rect 352 -354 353 -353
rect 135 -356 136 -355
rect 156 -356 157 -355
rect 289 -356 290 -355
rect 310 -356 311 -355
rect 156 -358 157 -357
rect 268 -358 269 -357
rect 282 -358 283 -357
rect 310 -358 311 -357
rect 268 -360 269 -359
rect 425 -360 426 -359
rect 271 -362 272 -361
rect 282 -362 283 -361
rect 2 -373 3 -372
rect 173 -373 174 -372
rect 201 -373 202 -372
rect 219 -373 220 -372
rect 222 -373 223 -372
rect 359 -373 360 -372
rect 9 -375 10 -374
rect 30 -375 31 -374
rect 37 -375 38 -374
rect 89 -375 90 -374
rect 110 -375 111 -374
rect 366 -375 367 -374
rect 16 -377 17 -376
rect 23 -377 24 -376
rect 26 -377 27 -376
rect 236 -377 237 -376
rect 247 -377 248 -376
rect 257 -377 258 -376
rect 268 -377 269 -376
rect 310 -377 311 -376
rect 317 -377 318 -376
rect 366 -377 367 -376
rect 16 -379 17 -378
rect 51 -379 52 -378
rect 65 -379 66 -378
rect 198 -379 199 -378
rect 226 -379 227 -378
rect 233 -379 234 -378
rect 271 -379 272 -378
rect 394 -379 395 -378
rect 30 -381 31 -380
rect 47 -381 48 -380
rect 68 -381 69 -380
rect 191 -381 192 -380
rect 271 -381 272 -380
rect 289 -381 290 -380
rect 317 -381 318 -380
rect 324 -381 325 -380
rect 338 -381 339 -380
rect 359 -381 360 -380
rect 387 -381 388 -380
rect 394 -381 395 -380
rect 37 -383 38 -382
rect 58 -383 59 -382
rect 79 -383 80 -382
rect 327 -383 328 -382
rect 61 -385 62 -384
rect 79 -385 80 -384
rect 82 -385 83 -384
rect 296 -385 297 -384
rect 86 -387 87 -386
rect 205 -387 206 -386
rect 212 -387 213 -386
rect 289 -387 290 -386
rect 72 -389 73 -388
rect 86 -389 87 -388
rect 110 -389 111 -388
rect 345 -389 346 -388
rect 72 -391 73 -390
rect 100 -391 101 -390
rect 114 -391 115 -390
rect 408 -391 409 -390
rect 100 -393 101 -392
rect 163 -393 164 -392
rect 184 -393 185 -392
rect 219 -393 220 -392
rect 229 -393 230 -392
rect 387 -393 388 -392
rect 408 -393 409 -392
rect 429 -393 430 -392
rect 117 -395 118 -394
rect 415 -395 416 -394
rect 135 -397 136 -396
rect 166 -397 167 -396
rect 205 -397 206 -396
rect 250 -397 251 -396
rect 261 -397 262 -396
rect 338 -397 339 -396
rect 352 -397 353 -396
rect 429 -397 430 -396
rect 135 -399 136 -398
rect 159 -399 160 -398
rect 163 -399 164 -398
rect 310 -399 311 -398
rect 331 -399 332 -398
rect 352 -399 353 -398
rect 415 -399 416 -398
rect 422 -399 423 -398
rect 142 -401 143 -400
rect 191 -401 192 -400
rect 212 -401 213 -400
rect 240 -401 241 -400
rect 261 -401 262 -400
rect 401 -401 402 -400
rect 422 -401 423 -400
rect 436 -401 437 -400
rect 93 -403 94 -402
rect 142 -403 143 -402
rect 149 -403 150 -402
rect 156 -403 157 -402
rect 184 -403 185 -402
rect 240 -403 241 -402
rect 275 -403 276 -402
rect 296 -403 297 -402
rect 303 -403 304 -402
rect 345 -403 346 -402
rect 373 -403 374 -402
rect 401 -403 402 -402
rect 432 -403 433 -402
rect 436 -403 437 -402
rect 54 -405 55 -404
rect 93 -405 94 -404
rect 121 -405 122 -404
rect 149 -405 150 -404
rect 170 -405 171 -404
rect 303 -405 304 -404
rect 373 -405 374 -404
rect 380 -405 381 -404
rect 47 -407 48 -406
rect 121 -407 122 -406
rect 128 -407 129 -406
rect 156 -407 157 -406
rect 170 -407 171 -406
rect 177 -407 178 -406
rect 254 -407 255 -406
rect 275 -407 276 -406
rect 58 -409 59 -408
rect 177 -409 178 -408
rect 264 -409 265 -408
rect 380 -409 381 -408
rect 117 -411 118 -410
rect 254 -411 255 -410
rect 9 -422 10 -421
rect 51 -422 52 -421
rect 79 -422 80 -421
rect 82 -422 83 -421
rect 107 -422 108 -421
rect 215 -422 216 -421
rect 226 -422 227 -421
rect 345 -422 346 -421
rect 432 -422 433 -421
rect 457 -422 458 -421
rect 16 -424 17 -423
rect 33 -424 34 -423
rect 44 -424 45 -423
rect 142 -424 143 -423
rect 166 -424 167 -423
rect 170 -424 171 -423
rect 194 -424 195 -423
rect 212 -424 213 -423
rect 229 -424 230 -423
rect 289 -424 290 -423
rect 317 -424 318 -423
rect 345 -424 346 -423
rect 359 -424 360 -423
rect 432 -424 433 -423
rect 443 -424 444 -423
rect 450 -424 451 -423
rect 16 -426 17 -425
rect 26 -426 27 -425
rect 30 -426 31 -425
rect 75 -426 76 -425
rect 79 -426 80 -425
rect 86 -426 87 -425
rect 93 -426 94 -425
rect 107 -426 108 -425
rect 121 -426 122 -425
rect 142 -426 143 -425
rect 163 -426 164 -425
rect 289 -426 290 -425
rect 327 -426 328 -425
rect 422 -426 423 -425
rect 446 -426 447 -425
rect 464 -426 465 -425
rect 51 -428 52 -427
rect 72 -428 73 -427
rect 86 -428 87 -427
rect 100 -428 101 -427
rect 121 -428 122 -427
rect 135 -428 136 -427
rect 156 -428 157 -427
rect 163 -428 164 -427
rect 177 -428 178 -427
rect 317 -428 318 -427
rect 334 -428 335 -427
rect 401 -428 402 -427
rect 58 -430 59 -429
rect 72 -430 73 -429
rect 82 -430 83 -429
rect 100 -430 101 -429
rect 114 -430 115 -429
rect 177 -430 178 -429
rect 201 -430 202 -429
rect 338 -430 339 -429
rect 352 -430 353 -429
rect 359 -430 360 -429
rect 93 -432 94 -431
rect 180 -432 181 -431
rect 212 -432 213 -431
rect 233 -432 234 -431
rect 236 -432 237 -431
rect 338 -432 339 -431
rect 128 -434 129 -433
rect 219 -434 220 -433
rect 240 -434 241 -433
rect 422 -434 423 -433
rect 117 -436 118 -435
rect 128 -436 129 -435
rect 131 -436 132 -435
rect 149 -436 150 -435
rect 156 -436 157 -435
rect 191 -436 192 -435
rect 243 -436 244 -435
rect 303 -436 304 -435
rect 135 -438 136 -437
rect 184 -438 185 -437
rect 191 -438 192 -437
rect 436 -438 437 -437
rect 149 -440 150 -439
rect 198 -440 199 -439
rect 247 -440 248 -439
rect 296 -440 297 -439
rect 387 -440 388 -439
rect 436 -440 437 -439
rect 226 -442 227 -441
rect 296 -442 297 -441
rect 387 -442 388 -441
rect 408 -442 409 -441
rect 250 -444 251 -443
rect 394 -444 395 -443
rect 250 -446 251 -445
rect 415 -446 416 -445
rect 254 -448 255 -447
rect 303 -448 304 -447
rect 310 -448 311 -447
rect 415 -448 416 -447
rect 254 -450 255 -449
rect 352 -450 353 -449
rect 373 -450 374 -449
rect 394 -450 395 -449
rect 257 -452 258 -451
rect 366 -452 367 -451
rect 373 -452 374 -451
rect 380 -452 381 -451
rect 261 -454 262 -453
rect 331 -454 332 -453
rect 170 -456 171 -455
rect 261 -456 262 -455
rect 268 -456 269 -455
rect 380 -456 381 -455
rect 65 -458 66 -457
rect 268 -458 269 -457
rect 275 -458 276 -457
rect 310 -458 311 -457
rect 324 -458 325 -457
rect 366 -458 367 -457
rect 47 -460 48 -459
rect 275 -460 276 -459
rect 282 -460 283 -459
rect 324 -460 325 -459
rect 65 -462 66 -461
rect 205 -462 206 -461
rect 184 -464 185 -463
rect 282 -464 283 -463
rect 205 -466 206 -465
rect 222 -466 223 -465
rect 9 -477 10 -476
rect 124 -477 125 -476
rect 142 -477 143 -476
rect 233 -477 234 -476
rect 247 -477 248 -476
rect 254 -477 255 -476
rect 261 -477 262 -476
rect 317 -477 318 -476
rect 352 -477 353 -476
rect 401 -477 402 -476
rect 418 -477 419 -476
rect 450 -477 451 -476
rect 30 -479 31 -478
rect 236 -479 237 -478
rect 250 -479 251 -478
rect 338 -479 339 -478
rect 345 -479 346 -478
rect 352 -479 353 -478
rect 387 -479 388 -478
rect 408 -479 409 -478
rect 422 -479 423 -478
rect 446 -479 447 -478
rect 33 -481 34 -480
rect 215 -481 216 -480
rect 222 -481 223 -480
rect 415 -481 416 -480
rect 432 -481 433 -480
rect 436 -481 437 -480
rect 37 -483 38 -482
rect 128 -483 129 -482
rect 131 -483 132 -482
rect 345 -483 346 -482
rect 380 -483 381 -482
rect 387 -483 388 -482
rect 415 -483 416 -482
rect 450 -483 451 -482
rect 16 -485 17 -484
rect 37 -485 38 -484
rect 40 -485 41 -484
rect 58 -485 59 -484
rect 72 -485 73 -484
rect 93 -485 94 -484
rect 100 -485 101 -484
rect 142 -485 143 -484
rect 173 -485 174 -484
rect 198 -485 199 -484
rect 205 -485 206 -484
rect 261 -485 262 -484
rect 264 -485 265 -484
rect 310 -485 311 -484
rect 359 -485 360 -484
rect 380 -485 381 -484
rect 16 -487 17 -486
rect 23 -487 24 -486
rect 44 -487 45 -486
rect 138 -487 139 -486
rect 180 -487 181 -486
rect 429 -487 430 -486
rect 51 -489 52 -488
rect 103 -489 104 -488
rect 107 -489 108 -488
rect 226 -489 227 -488
rect 240 -489 241 -488
rect 436 -489 437 -488
rect 51 -491 52 -490
rect 72 -491 73 -490
rect 82 -491 83 -490
rect 177 -491 178 -490
rect 191 -491 192 -490
rect 219 -491 220 -490
rect 275 -491 276 -490
rect 282 -491 283 -490
rect 285 -491 286 -490
rect 394 -491 395 -490
rect 429 -491 430 -490
rect 457 -491 458 -490
rect 58 -493 59 -492
rect 79 -493 80 -492
rect 93 -493 94 -492
rect 110 -493 111 -492
rect 128 -493 129 -492
rect 135 -493 136 -492
rect 184 -493 185 -492
rect 191 -493 192 -492
rect 212 -493 213 -492
rect 247 -493 248 -492
rect 296 -493 297 -492
rect 317 -493 318 -492
rect 359 -493 360 -492
rect 366 -493 367 -492
rect 443 -493 444 -492
rect 457 -493 458 -492
rect 79 -495 80 -494
rect 331 -495 332 -494
rect 107 -497 108 -496
rect 121 -497 122 -496
rect 156 -497 157 -496
rect 184 -497 185 -496
rect 268 -497 269 -496
rect 331 -497 332 -496
rect 121 -499 122 -498
rect 163 -499 164 -498
rect 170 -499 171 -498
rect 268 -499 269 -498
rect 289 -499 290 -498
rect 296 -499 297 -498
rect 303 -499 304 -498
rect 338 -499 339 -498
rect 65 -501 66 -500
rect 289 -501 290 -500
rect 310 -501 311 -500
rect 324 -501 325 -500
rect 65 -503 66 -502
rect 86 -503 87 -502
rect 156 -503 157 -502
rect 194 -503 195 -502
rect 243 -503 244 -502
rect 324 -503 325 -502
rect 86 -505 87 -504
rect 149 -505 150 -504
rect 163 -505 164 -504
rect 303 -505 304 -504
rect 149 -507 150 -506
rect 205 -507 206 -506
rect 9 -518 10 -517
rect 68 -518 69 -517
rect 72 -518 73 -517
rect 93 -518 94 -517
rect 117 -518 118 -517
rect 124 -518 125 -517
rect 138 -518 139 -517
rect 436 -518 437 -517
rect 9 -520 10 -519
rect 103 -520 104 -519
rect 121 -520 122 -519
rect 226 -520 227 -519
rect 243 -520 244 -519
rect 254 -520 255 -519
rect 278 -520 279 -519
rect 352 -520 353 -519
rect 366 -520 367 -519
rect 422 -520 423 -519
rect 429 -520 430 -519
rect 443 -520 444 -519
rect 16 -522 17 -521
rect 37 -522 38 -521
rect 44 -522 45 -521
rect 205 -522 206 -521
rect 208 -522 209 -521
rect 338 -522 339 -521
rect 401 -522 402 -521
rect 415 -522 416 -521
rect 443 -522 444 -521
rect 457 -522 458 -521
rect 19 -524 20 -523
rect 275 -524 276 -523
rect 285 -524 286 -523
rect 380 -524 381 -523
rect 457 -524 458 -523
rect 464 -524 465 -523
rect 37 -526 38 -525
rect 156 -526 157 -525
rect 166 -526 167 -525
rect 254 -526 255 -525
rect 303 -526 304 -525
rect 408 -526 409 -525
rect 450 -526 451 -525
rect 464 -526 465 -525
rect 44 -528 45 -527
rect 51 -528 52 -527
rect 58 -528 59 -527
rect 96 -528 97 -527
rect 124 -528 125 -527
rect 173 -528 174 -527
rect 184 -528 185 -527
rect 205 -528 206 -527
rect 212 -528 213 -527
rect 331 -528 332 -527
rect 359 -528 360 -527
rect 380 -528 381 -527
rect 30 -530 31 -529
rect 58 -530 59 -529
rect 72 -530 73 -529
rect 170 -530 171 -529
rect 173 -530 174 -529
rect 436 -530 437 -529
rect 30 -532 31 -531
rect 93 -532 94 -531
rect 149 -532 150 -531
rect 187 -532 188 -531
rect 212 -532 213 -531
rect 268 -532 269 -531
rect 306 -532 307 -531
rect 341 -532 342 -531
rect 373 -532 374 -531
rect 415 -532 416 -531
rect 26 -534 27 -533
rect 268 -534 269 -533
rect 310 -534 311 -533
rect 352 -534 353 -533
rect 373 -534 374 -533
rect 432 -534 433 -533
rect 51 -536 52 -535
rect 65 -536 66 -535
rect 82 -536 83 -535
rect 366 -536 367 -535
rect 40 -538 41 -537
rect 65 -538 66 -537
rect 82 -538 83 -537
rect 282 -538 283 -537
rect 324 -538 325 -537
rect 394 -538 395 -537
rect 86 -540 87 -539
rect 156 -540 157 -539
rect 184 -540 185 -539
rect 359 -540 360 -539
rect 86 -542 87 -541
rect 107 -542 108 -541
rect 149 -542 150 -541
rect 163 -542 164 -541
rect 198 -542 199 -541
rect 310 -542 311 -541
rect 331 -542 332 -541
rect 345 -542 346 -541
rect 107 -544 108 -543
rect 128 -544 129 -543
rect 163 -544 164 -543
rect 177 -544 178 -543
rect 219 -544 220 -543
rect 226 -544 227 -543
rect 233 -544 234 -543
rect 408 -544 409 -543
rect 103 -546 104 -545
rect 128 -546 129 -545
rect 135 -546 136 -545
rect 177 -546 178 -545
rect 191 -546 192 -545
rect 219 -546 220 -545
rect 233 -546 234 -545
rect 387 -546 388 -545
rect 114 -548 115 -547
rect 198 -548 199 -547
rect 240 -548 241 -547
rect 387 -548 388 -547
rect 191 -550 192 -549
rect 215 -550 216 -549
rect 247 -550 248 -549
rect 275 -550 276 -549
rect 282 -550 283 -549
rect 401 -550 402 -549
rect 247 -552 248 -551
rect 261 -552 262 -551
rect 296 -552 297 -551
rect 324 -552 325 -551
rect 23 -554 24 -553
rect 296 -554 297 -553
rect 317 -554 318 -553
rect 345 -554 346 -553
rect 236 -556 237 -555
rect 261 -556 262 -555
rect 289 -556 290 -555
rect 317 -556 318 -555
rect 142 -558 143 -557
rect 289 -558 290 -557
rect 114 -560 115 -559
rect 142 -560 143 -559
rect 9 -571 10 -570
rect 184 -571 185 -570
rect 212 -571 213 -570
rect 264 -571 265 -570
rect 303 -571 304 -570
rect 345 -571 346 -570
rect 464 -571 465 -570
rect 471 -571 472 -570
rect 16 -573 17 -572
rect 100 -573 101 -572
rect 138 -573 139 -572
rect 303 -573 304 -572
rect 341 -573 342 -572
rect 394 -573 395 -572
rect 457 -573 458 -572
rect 464 -573 465 -572
rect 16 -575 17 -574
rect 114 -575 115 -574
rect 163 -575 164 -574
rect 446 -575 447 -574
rect 23 -577 24 -576
rect 128 -577 129 -576
rect 163 -577 164 -576
rect 208 -577 209 -576
rect 233 -577 234 -576
rect 247 -577 248 -576
rect 257 -577 258 -576
rect 401 -577 402 -576
rect 9 -579 10 -578
rect 208 -579 209 -578
rect 236 -579 237 -578
rect 366 -579 367 -578
rect 394 -579 395 -578
rect 429 -579 430 -578
rect 30 -581 31 -580
rect 103 -581 104 -580
rect 170 -581 171 -580
rect 282 -581 283 -580
rect 33 -583 34 -582
rect 44 -583 45 -582
rect 58 -583 59 -582
rect 89 -583 90 -582
rect 93 -583 94 -582
rect 243 -583 244 -582
rect 247 -583 248 -582
rect 317 -583 318 -582
rect 40 -585 41 -584
rect 429 -585 430 -584
rect 44 -587 45 -586
rect 51 -587 52 -586
rect 58 -587 59 -586
rect 107 -587 108 -586
rect 149 -587 150 -586
rect 282 -587 283 -586
rect 317 -587 318 -586
rect 331 -587 332 -586
rect 37 -589 38 -588
rect 51 -589 52 -588
rect 65 -589 66 -588
rect 156 -589 157 -588
rect 173 -589 174 -588
rect 219 -589 220 -588
rect 240 -589 241 -588
rect 352 -589 353 -588
rect 68 -591 69 -590
rect 345 -591 346 -590
rect 352 -591 353 -590
rect 359 -591 360 -590
rect 79 -593 80 -592
rect 289 -593 290 -592
rect 331 -593 332 -592
rect 366 -593 367 -592
rect 72 -595 73 -594
rect 79 -595 80 -594
rect 93 -595 94 -594
rect 436 -595 437 -594
rect 30 -597 31 -596
rect 436 -597 437 -596
rect 72 -599 73 -598
rect 86 -599 87 -598
rect 107 -599 108 -598
rect 194 -599 195 -598
rect 205 -599 206 -598
rect 233 -599 234 -598
rect 240 -599 241 -598
rect 268 -599 269 -598
rect 289 -599 290 -598
rect 324 -599 325 -598
rect 359 -599 360 -598
rect 380 -599 381 -598
rect 86 -601 87 -600
rect 142 -601 143 -600
rect 156 -601 157 -600
rect 173 -601 174 -600
rect 177 -601 178 -600
rect 191 -601 192 -600
rect 219 -601 220 -600
rect 275 -601 276 -600
rect 306 -601 307 -600
rect 380 -601 381 -600
rect 135 -603 136 -602
rect 149 -603 150 -602
rect 180 -603 181 -602
rect 408 -603 409 -602
rect 142 -605 143 -604
rect 170 -605 171 -604
rect 254 -605 255 -604
rect 401 -605 402 -604
rect 268 -607 269 -606
rect 310 -607 311 -606
rect 338 -607 339 -606
rect 408 -607 409 -606
rect 261 -609 262 -608
rect 310 -609 311 -608
rect 338 -609 339 -608
rect 373 -609 374 -608
rect 275 -611 276 -610
rect 296 -611 297 -610
rect 373 -611 374 -610
rect 387 -611 388 -610
rect 296 -613 297 -612
rect 324 -613 325 -612
rect 387 -613 388 -612
rect 453 -613 454 -612
rect 2 -624 3 -623
rect 51 -624 52 -623
rect 72 -624 73 -623
rect 114 -624 115 -623
rect 117 -624 118 -623
rect 212 -624 213 -623
rect 222 -624 223 -623
rect 268 -624 269 -623
rect 299 -624 300 -623
rect 422 -624 423 -623
rect 436 -624 437 -623
rect 443 -624 444 -623
rect 450 -624 451 -623
rect 457 -624 458 -623
rect 460 -624 461 -623
rect 464 -624 465 -623
rect 9 -626 10 -625
rect 103 -626 104 -625
rect 170 -626 171 -625
rect 184 -626 185 -625
rect 187 -626 188 -625
rect 282 -626 283 -625
rect 299 -626 300 -625
rect 415 -626 416 -625
rect 429 -626 430 -625
rect 436 -626 437 -625
rect 9 -628 10 -627
rect 75 -628 76 -627
rect 79 -628 80 -627
rect 131 -628 132 -627
rect 142 -628 143 -627
rect 170 -628 171 -627
rect 191 -628 192 -627
rect 215 -628 216 -627
rect 233 -628 234 -627
rect 422 -628 423 -627
rect 23 -630 24 -629
rect 135 -630 136 -629
rect 142 -630 143 -629
rect 226 -630 227 -629
rect 240 -630 241 -629
rect 254 -630 255 -629
rect 261 -630 262 -629
rect 352 -630 353 -629
rect 380 -630 381 -629
rect 429 -630 430 -629
rect 16 -632 17 -631
rect 23 -632 24 -631
rect 30 -632 31 -631
rect 163 -632 164 -631
rect 194 -632 195 -631
rect 401 -632 402 -631
rect 415 -632 416 -631
rect 446 -632 447 -631
rect 16 -634 17 -633
rect 65 -634 66 -633
rect 93 -634 94 -633
rect 96 -634 97 -633
rect 128 -634 129 -633
rect 194 -634 195 -633
rect 205 -634 206 -633
rect 303 -634 304 -633
rect 331 -634 332 -633
rect 359 -634 360 -633
rect 33 -636 34 -635
rect 65 -636 66 -635
rect 86 -636 87 -635
rect 128 -636 129 -635
rect 135 -636 136 -635
rect 149 -636 150 -635
rect 208 -636 209 -635
rect 387 -636 388 -635
rect 37 -638 38 -637
rect 198 -638 199 -637
rect 215 -638 216 -637
rect 282 -638 283 -637
rect 289 -638 290 -637
rect 303 -638 304 -637
rect 331 -638 332 -637
rect 352 -638 353 -637
rect 387 -638 388 -637
rect 394 -638 395 -637
rect 37 -640 38 -639
rect 177 -640 178 -639
rect 180 -640 181 -639
rect 394 -640 395 -639
rect 40 -642 41 -641
rect 271 -642 272 -641
rect 334 -642 335 -641
rect 408 -642 409 -641
rect 44 -644 45 -643
rect 51 -644 52 -643
rect 54 -644 55 -643
rect 450 -644 451 -643
rect 44 -646 45 -645
rect 275 -646 276 -645
rect 345 -646 346 -645
rect 380 -646 381 -645
rect 58 -648 59 -647
rect 79 -648 80 -647
rect 93 -648 94 -647
rect 121 -648 122 -647
rect 156 -648 157 -647
rect 198 -648 199 -647
rect 219 -648 220 -647
rect 233 -648 234 -647
rect 243 -648 244 -647
rect 359 -648 360 -647
rect 366 -648 367 -647
rect 408 -648 409 -647
rect 58 -650 59 -649
rect 89 -650 90 -649
rect 96 -650 97 -649
rect 121 -650 122 -649
rect 163 -650 164 -649
rect 208 -650 209 -649
rect 226 -650 227 -649
rect 247 -650 248 -649
rect 254 -650 255 -649
rect 457 -650 458 -649
rect 107 -652 108 -651
rect 149 -652 150 -651
rect 184 -652 185 -651
rect 289 -652 290 -651
rect 324 -652 325 -651
rect 366 -652 367 -651
rect 100 -654 101 -653
rect 107 -654 108 -653
rect 114 -654 115 -653
rect 177 -654 178 -653
rect 240 -654 241 -653
rect 324 -654 325 -653
rect 338 -654 339 -653
rect 345 -654 346 -653
rect 100 -656 101 -655
rect 156 -656 157 -655
rect 261 -656 262 -655
rect 317 -656 318 -655
rect 103 -658 104 -657
rect 338 -658 339 -657
rect 250 -660 251 -659
rect 317 -660 318 -659
rect 250 -662 251 -661
rect 401 -662 402 -661
rect 275 -664 276 -663
rect 296 -664 297 -663
rect 2 -675 3 -674
rect 131 -675 132 -674
rect 135 -675 136 -674
rect 180 -675 181 -674
rect 187 -675 188 -674
rect 219 -675 220 -674
rect 233 -675 234 -674
rect 240 -675 241 -674
rect 250 -675 251 -674
rect 303 -675 304 -674
rect 331 -675 332 -674
rect 338 -675 339 -674
rect 443 -675 444 -674
rect 457 -675 458 -674
rect 464 -675 465 -674
rect 471 -675 472 -674
rect 16 -677 17 -676
rect 100 -677 101 -676
rect 114 -677 115 -676
rect 149 -677 150 -676
rect 170 -677 171 -676
rect 173 -677 174 -676
rect 191 -677 192 -676
rect 317 -677 318 -676
rect 334 -677 335 -676
rect 429 -677 430 -676
rect 9 -679 10 -678
rect 16 -679 17 -678
rect 37 -679 38 -678
rect 177 -679 178 -678
rect 191 -679 192 -678
rect 226 -679 227 -678
rect 250 -679 251 -678
rect 436 -679 437 -678
rect 9 -681 10 -680
rect 93 -681 94 -680
rect 128 -681 129 -680
rect 401 -681 402 -680
rect 23 -683 24 -682
rect 93 -683 94 -682
rect 149 -683 150 -682
rect 240 -683 241 -682
rect 268 -683 269 -682
rect 317 -683 318 -682
rect 380 -683 381 -682
rect 429 -683 430 -682
rect 23 -685 24 -684
rect 289 -685 290 -684
rect 296 -685 297 -684
rect 366 -685 367 -684
rect 380 -685 381 -684
rect 408 -685 409 -684
rect 37 -687 38 -686
rect 205 -687 206 -686
rect 212 -687 213 -686
rect 422 -687 423 -686
rect 40 -689 41 -688
rect 131 -689 132 -688
rect 170 -689 171 -688
rect 212 -689 213 -688
rect 229 -689 230 -688
rect 289 -689 290 -688
rect 299 -689 300 -688
rect 345 -689 346 -688
rect 359 -689 360 -688
rect 366 -689 367 -688
rect 401 -689 402 -688
rect 415 -689 416 -688
rect 44 -691 45 -690
rect 86 -691 87 -690
rect 177 -691 178 -690
rect 282 -691 283 -690
rect 345 -691 346 -690
rect 352 -691 353 -690
rect 359 -691 360 -690
rect 373 -691 374 -690
rect 51 -693 52 -692
rect 352 -693 353 -692
rect 58 -695 59 -694
rect 135 -695 136 -694
rect 194 -695 195 -694
rect 219 -695 220 -694
rect 268 -695 269 -694
rect 310 -695 311 -694
rect 58 -697 59 -696
rect 254 -697 255 -696
rect 261 -697 262 -696
rect 310 -697 311 -696
rect 72 -699 73 -698
rect 100 -699 101 -698
rect 198 -699 199 -698
rect 215 -699 216 -698
rect 254 -699 255 -698
rect 275 -699 276 -698
rect 282 -699 283 -698
rect 324 -699 325 -698
rect 2 -701 3 -700
rect 72 -701 73 -700
rect 75 -701 76 -700
rect 184 -701 185 -700
rect 261 -701 262 -700
rect 373 -701 374 -700
rect 79 -703 80 -702
rect 114 -703 115 -702
rect 142 -703 143 -702
rect 198 -703 199 -702
rect 324 -703 325 -702
rect 394 -703 395 -702
rect 82 -705 83 -704
rect 107 -705 108 -704
rect 142 -705 143 -704
rect 156 -705 157 -704
rect 184 -705 185 -704
rect 233 -705 234 -704
rect 394 -705 395 -704
rect 450 -705 451 -704
rect 65 -707 66 -706
rect 107 -707 108 -706
rect 156 -707 157 -706
rect 163 -707 164 -706
rect 54 -709 55 -708
rect 65 -709 66 -708
rect 86 -709 87 -708
rect 124 -709 125 -708
rect 121 -711 122 -710
rect 163 -711 164 -710
rect 30 -713 31 -712
rect 121 -713 122 -712
rect 30 -715 31 -714
rect 117 -715 118 -714
rect 9 -726 10 -725
rect 72 -726 73 -725
rect 96 -726 97 -725
rect 184 -726 185 -725
rect 198 -726 199 -725
rect 352 -726 353 -725
rect 376 -726 377 -725
rect 401 -726 402 -725
rect 411 -726 412 -725
rect 429 -726 430 -725
rect 16 -728 17 -727
rect 75 -728 76 -727
rect 110 -728 111 -727
rect 250 -728 251 -727
rect 254 -728 255 -727
rect 278 -728 279 -727
rect 289 -728 290 -727
rect 296 -728 297 -727
rect 338 -728 339 -727
rect 380 -728 381 -727
rect 387 -728 388 -727
rect 408 -728 409 -727
rect 23 -730 24 -729
rect 198 -730 199 -729
rect 215 -730 216 -729
rect 233 -730 234 -729
rect 243 -730 244 -729
rect 310 -730 311 -729
rect 341 -730 342 -729
rect 345 -730 346 -729
rect 2 -732 3 -731
rect 310 -732 311 -731
rect 345 -732 346 -731
rect 359 -732 360 -731
rect 23 -734 24 -733
rect 86 -734 87 -733
rect 121 -734 122 -733
rect 303 -734 304 -733
rect 37 -736 38 -735
rect 79 -736 80 -735
rect 86 -736 87 -735
rect 191 -736 192 -735
rect 233 -736 234 -735
rect 268 -736 269 -735
rect 289 -736 290 -735
rect 324 -736 325 -735
rect 37 -738 38 -737
rect 180 -738 181 -737
rect 205 -738 206 -737
rect 268 -738 269 -737
rect 324 -738 325 -737
rect 394 -738 395 -737
rect 40 -740 41 -739
rect 58 -740 59 -739
rect 65 -740 66 -739
rect 75 -740 76 -739
rect 128 -740 129 -739
rect 254 -740 255 -739
rect 16 -742 17 -741
rect 58 -742 59 -741
rect 114 -742 115 -741
rect 128 -742 129 -741
rect 135 -742 136 -741
rect 184 -742 185 -741
rect 247 -742 248 -741
rect 282 -742 283 -741
rect 44 -744 45 -743
rect 191 -744 192 -743
rect 236 -744 237 -743
rect 282 -744 283 -743
rect 44 -746 45 -745
rect 65 -746 66 -745
rect 93 -746 94 -745
rect 135 -746 136 -745
rect 142 -746 143 -745
rect 208 -746 209 -745
rect 51 -748 52 -747
rect 82 -748 83 -747
rect 100 -748 101 -747
rect 142 -748 143 -747
rect 156 -748 157 -747
rect 201 -748 202 -747
rect 54 -750 55 -749
rect 240 -750 241 -749
rect 82 -752 83 -751
rect 114 -752 115 -751
rect 163 -752 164 -751
rect 170 -752 171 -751
rect 180 -752 181 -751
rect 317 -752 318 -751
rect 100 -754 101 -753
rect 261 -754 262 -753
rect 30 -756 31 -755
rect 261 -756 262 -755
rect 103 -758 104 -757
rect 208 -758 209 -757
rect 107 -760 108 -759
rect 156 -760 157 -759
rect 163 -760 164 -759
rect 226 -760 227 -759
rect 219 -762 220 -761
rect 226 -762 227 -761
rect 212 -764 213 -763
rect 219 -764 220 -763
rect 212 -766 213 -765
rect 331 -766 332 -765
rect 331 -768 332 -767
rect 366 -768 367 -767
rect 9 -779 10 -778
rect 47 -779 48 -778
rect 58 -779 59 -778
rect 107 -779 108 -778
rect 110 -779 111 -778
rect 156 -779 157 -778
rect 177 -779 178 -778
rect 303 -779 304 -778
rect 317 -779 318 -778
rect 338 -779 339 -778
rect 30 -781 31 -780
rect 51 -781 52 -780
rect 65 -781 66 -780
rect 75 -781 76 -780
rect 93 -781 94 -780
rect 142 -781 143 -780
rect 177 -781 178 -780
rect 226 -781 227 -780
rect 233 -781 234 -780
rect 261 -781 262 -780
rect 51 -783 52 -782
rect 79 -783 80 -782
rect 96 -783 97 -782
rect 254 -783 255 -782
rect 72 -785 73 -784
rect 82 -785 83 -784
rect 100 -785 101 -784
rect 152 -785 153 -784
rect 163 -785 164 -784
rect 261 -785 262 -784
rect 103 -787 104 -786
rect 303 -787 304 -786
rect 107 -789 108 -788
rect 240 -789 241 -788
rect 247 -789 248 -788
rect 275 -789 276 -788
rect 30 -791 31 -790
rect 247 -791 248 -790
rect 254 -791 255 -790
rect 282 -791 283 -790
rect 117 -793 118 -792
rect 170 -793 171 -792
rect 205 -793 206 -792
rect 212 -793 213 -792
rect 219 -793 220 -792
rect 226 -793 227 -792
rect 282 -793 283 -792
rect 289 -793 290 -792
rect 23 -795 24 -794
rect 170 -795 171 -794
rect 212 -795 213 -794
rect 236 -795 237 -794
rect 23 -797 24 -796
rect 61 -797 62 -796
rect 124 -797 125 -796
rect 135 -797 136 -796
rect 163 -797 164 -796
rect 191 -797 192 -796
rect 33 -799 34 -798
rect 135 -799 136 -798
rect 149 -799 150 -798
rect 191 -799 192 -798
rect 33 -801 34 -800
rect 117 -801 118 -800
rect 124 -801 125 -800
rect 184 -801 185 -800
rect 37 -803 38 -802
rect 289 -803 290 -802
rect 37 -805 38 -804
rect 114 -805 115 -804
rect 128 -805 129 -804
rect 156 -805 157 -804
rect 86 -807 87 -806
rect 184 -807 185 -806
rect 131 -809 132 -808
rect 310 -809 311 -808
rect 310 -811 311 -810
rect 324 -811 325 -810
rect 324 -813 325 -812
rect 345 -813 346 -812
rect 9 -824 10 -823
rect 16 -824 17 -823
rect 23 -824 24 -823
rect 65 -824 66 -823
rect 72 -824 73 -823
rect 93 -824 94 -823
rect 96 -824 97 -823
rect 233 -824 234 -823
rect 240 -824 241 -823
rect 268 -824 269 -823
rect 292 -824 293 -823
rect 317 -824 318 -823
rect 324 -824 325 -823
rect 345 -824 346 -823
rect 23 -826 24 -825
rect 261 -826 262 -825
rect 310 -826 311 -825
rect 327 -826 328 -825
rect 33 -828 34 -827
rect 47 -828 48 -827
rect 58 -828 59 -827
rect 79 -828 80 -827
rect 86 -828 87 -827
rect 114 -828 115 -827
rect 117 -828 118 -827
rect 191 -828 192 -827
rect 222 -828 223 -827
rect 226 -828 227 -827
rect 254 -828 255 -827
rect 268 -828 269 -827
rect 37 -830 38 -829
rect 89 -830 90 -829
rect 117 -830 118 -829
rect 289 -830 290 -829
rect 33 -832 34 -831
rect 37 -832 38 -831
rect 72 -832 73 -831
rect 100 -832 101 -831
rect 124 -832 125 -831
rect 163 -832 164 -831
rect 191 -832 192 -831
rect 247 -832 248 -831
rect 51 -834 52 -833
rect 163 -834 164 -833
rect 212 -834 213 -833
rect 226 -834 227 -833
rect 44 -836 45 -835
rect 51 -836 52 -835
rect 128 -836 129 -835
rect 156 -836 157 -835
rect 205 -836 206 -835
rect 212 -836 213 -835
rect 19 -838 20 -837
rect 44 -838 45 -837
rect 135 -838 136 -837
rect 180 -838 181 -837
rect 135 -840 136 -839
rect 145 -840 146 -839
rect 149 -840 150 -839
rect 198 -840 199 -839
rect 152 -842 153 -841
rect 303 -842 304 -841
rect 156 -844 157 -843
rect 170 -844 171 -843
rect 170 -846 171 -845
rect 289 -846 290 -845
rect 23 -857 24 -856
rect 142 -857 143 -856
rect 187 -857 188 -856
rect 191 -857 192 -856
rect 268 -857 269 -856
rect 285 -857 286 -856
rect 37 -859 38 -858
rect 44 -859 45 -858
rect 47 -859 48 -858
rect 58 -859 59 -858
rect 65 -859 66 -858
rect 86 -859 87 -858
rect 93 -859 94 -858
rect 114 -859 115 -858
rect 131 -859 132 -858
rect 149 -859 150 -858
rect 54 -861 55 -860
rect 170 -861 171 -860
rect 72 -863 73 -862
rect 103 -863 104 -862
rect 107 -863 108 -862
rect 156 -863 157 -862
rect 82 -865 83 -864
rect 163 -865 164 -864
<< metal2 >>
rect 12 -5 13 1
rect 26 -5 27 1
rect 37 -5 38 1
rect 65 -5 66 1
rect 93 -5 94 1
rect 107 -5 108 1
rect 121 -5 122 1
rect 128 -5 129 1
rect 135 -5 136 1
rect 163 -5 164 1
rect 51 -5 52 -1
rect 89 -5 90 -1
rect 138 -5 139 -1
rect 149 -5 150 -1
rect 58 -5 59 -3
rect 72 -5 73 -3
rect 72 -15 73 -13
rect 96 -15 97 -13
rect 100 -15 101 -13
rect 107 -15 108 -13
rect 114 -15 115 -13
rect 156 -15 157 -13
rect 159 -15 160 -13
rect 191 -24 192 -14
rect 65 -17 66 -13
rect 72 -24 73 -16
rect 79 -24 80 -16
rect 100 -24 101 -16
rect 107 -24 108 -16
rect 142 -24 143 -16
rect 145 -17 146 -13
rect 149 -17 150 -13
rect 163 -17 164 -13
rect 173 -24 174 -16
rect 114 -24 115 -18
rect 177 -24 178 -18
rect 128 -21 129 -13
rect 128 -24 129 -20
rect 128 -21 129 -13
rect 128 -24 129 -20
rect 149 -24 150 -20
rect 201 -24 202 -20
rect 163 -24 164 -22
rect 187 -24 188 -22
rect 5 -34 6 -32
rect 5 -55 6 -33
rect 5 -34 6 -32
rect 5 -55 6 -33
rect 30 -34 31 -32
rect 30 -55 31 -33
rect 30 -34 31 -32
rect 30 -55 31 -33
rect 47 -55 48 -33
rect 212 -55 213 -33
rect 51 -55 52 -35
rect 149 -36 150 -32
rect 163 -36 164 -32
rect 219 -55 220 -35
rect 58 -55 59 -37
rect 72 -38 73 -32
rect 86 -55 87 -37
rect 163 -55 164 -37
rect 177 -38 178 -32
rect 233 -55 234 -37
rect 16 -55 17 -39
rect 177 -55 178 -39
rect 191 -40 192 -32
rect 254 -55 255 -39
rect 65 -55 66 -41
rect 117 -42 118 -32
rect 121 -55 122 -41
rect 170 -55 171 -41
rect 198 -42 199 -32
rect 247 -55 248 -41
rect 72 -55 73 -43
rect 79 -55 80 -43
rect 93 -44 94 -32
rect 184 -55 185 -43
rect 37 -46 38 -32
rect 93 -55 94 -45
rect 96 -55 97 -45
rect 198 -55 199 -45
rect 124 -48 125 -32
rect 152 -55 153 -47
rect 100 -55 101 -49
rect 124 -55 125 -49
rect 128 -50 129 -32
rect 128 -55 129 -49
rect 128 -50 129 -32
rect 128 -55 129 -49
rect 142 -50 143 -32
rect 226 -55 227 -49
rect 145 -55 146 -51
rect 156 -55 157 -51
rect 149 -55 150 -53
rect 205 -55 206 -53
rect 19 -88 20 -64
rect 212 -65 213 -63
rect 219 -65 220 -63
rect 275 -88 276 -64
rect 40 -67 41 -63
rect 79 -88 80 -66
rect 82 -67 83 -63
rect 110 -67 111 -63
rect 121 -88 122 -66
rect 159 -88 160 -66
rect 177 -67 178 -63
rect 219 -88 220 -66
rect 226 -67 227 -63
rect 331 -88 332 -66
rect 40 -88 41 -68
rect 177 -88 178 -68
rect 191 -69 192 -63
rect 254 -69 255 -63
rect 44 -88 45 -70
rect 51 -71 52 -63
rect 58 -71 59 -63
rect 89 -71 90 -63
rect 100 -71 101 -63
rect 128 -71 129 -63
rect 131 -71 132 -63
rect 261 -88 262 -70
rect 30 -73 31 -63
rect 131 -88 132 -72
rect 138 -88 139 -72
rect 142 -88 143 -72
rect 149 -88 150 -72
rect 212 -88 213 -72
rect 233 -73 234 -63
rect 282 -88 283 -72
rect 30 -88 31 -74
rect 114 -75 115 -63
rect 163 -75 164 -63
rect 226 -88 227 -74
rect 243 -75 244 -63
rect 254 -88 255 -74
rect 51 -88 52 -76
rect 96 -88 97 -76
rect 107 -77 108 -63
rect 135 -77 136 -63
rect 184 -77 185 -63
rect 191 -88 192 -76
rect 205 -77 206 -63
rect 240 -88 241 -76
rect 247 -77 248 -63
rect 268 -88 269 -76
rect 58 -88 59 -78
rect 65 -79 66 -63
rect 86 -88 87 -78
rect 156 -79 157 -63
rect 170 -79 171 -63
rect 205 -88 206 -78
rect 65 -88 66 -80
rect 72 -81 73 -63
rect 110 -88 111 -80
rect 296 -88 297 -80
rect 72 -88 73 -82
rect 100 -88 101 -82
rect 170 -88 171 -82
rect 289 -88 290 -82
rect 184 -88 185 -84
rect 233 -88 234 -84
rect 198 -87 199 -63
rect 247 -88 248 -86
rect 23 -98 24 -96
rect 86 -98 87 -96
rect 93 -143 94 -97
rect 131 -98 132 -96
rect 135 -98 136 -96
rect 226 -98 227 -96
rect 268 -98 269 -96
rect 359 -143 360 -97
rect 26 -143 27 -99
rect 352 -143 353 -99
rect 30 -102 31 -96
rect 198 -102 199 -96
rect 201 -102 202 -96
rect 317 -143 318 -101
rect 331 -102 332 -96
rect 331 -143 332 -101
rect 331 -102 332 -96
rect 331 -143 332 -101
rect 51 -104 52 -96
rect 100 -143 101 -103
rect 107 -143 108 -103
rect 117 -104 118 -96
rect 121 -104 122 -96
rect 142 -143 143 -103
rect 145 -104 146 -96
rect 310 -143 311 -103
rect 51 -143 52 -105
rect 65 -106 66 -96
rect 96 -106 97 -96
rect 261 -106 262 -96
rect 271 -143 272 -105
rect 366 -143 367 -105
rect 58 -108 59 -96
rect 58 -143 59 -107
rect 58 -108 59 -96
rect 58 -143 59 -107
rect 65 -143 66 -107
rect 173 -108 174 -96
rect 194 -143 195 -107
rect 226 -143 227 -107
rect 254 -108 255 -96
rect 261 -143 262 -107
rect 275 -108 276 -96
rect 345 -143 346 -107
rect 30 -143 31 -109
rect 275 -143 276 -109
rect 289 -110 290 -96
rect 373 -143 374 -109
rect 86 -143 87 -111
rect 254 -143 255 -111
rect 303 -112 304 -96
rect 324 -143 325 -111
rect 128 -114 129 -96
rect 247 -114 248 -96
rect 138 -116 139 -96
rect 303 -143 304 -115
rect 138 -143 139 -117
rect 201 -143 202 -117
rect 233 -118 234 -96
rect 289 -143 290 -117
rect 149 -120 150 -96
rect 205 -120 206 -96
rect 233 -143 234 -119
rect 296 -120 297 -96
rect 149 -143 150 -121
rect 208 -143 209 -121
rect 240 -122 241 -96
rect 296 -143 297 -121
rect 152 -143 153 -123
rect 170 -143 171 -123
rect 191 -124 192 -96
rect 247 -143 248 -123
rect 156 -126 157 -96
rect 338 -143 339 -125
rect 44 -128 45 -96
rect 156 -143 157 -127
rect 163 -128 164 -96
rect 282 -128 283 -96
rect 9 -130 10 -96
rect 44 -143 45 -129
rect 124 -143 125 -129
rect 163 -143 164 -129
rect 166 -130 167 -96
rect 219 -130 220 -96
rect 37 -143 38 -131
rect 282 -143 283 -131
rect 166 -143 167 -133
rect 184 -143 185 -133
rect 212 -134 213 -96
rect 240 -143 241 -133
rect 128 -143 129 -135
rect 212 -143 213 -135
rect 177 -138 178 -96
rect 219 -143 220 -137
rect 72 -140 73 -96
rect 177 -143 178 -139
rect 72 -143 73 -141
rect 121 -143 122 -141
rect 5 -194 6 -152
rect 19 -153 20 -151
rect 23 -153 24 -151
rect 310 -153 311 -151
rect 324 -153 325 -151
rect 324 -194 325 -152
rect 324 -153 325 -151
rect 324 -194 325 -152
rect 331 -153 332 -151
rect 331 -194 332 -152
rect 331 -153 332 -151
rect 331 -194 332 -152
rect 345 -153 346 -151
rect 380 -194 381 -152
rect 9 -194 10 -154
rect 26 -194 27 -154
rect 61 -155 62 -151
rect 338 -155 339 -151
rect 345 -194 346 -154
rect 352 -155 353 -151
rect 373 -155 374 -151
rect 401 -194 402 -154
rect 16 -157 17 -151
rect 37 -157 38 -151
rect 65 -157 66 -151
rect 103 -194 104 -156
rect 128 -157 129 -151
rect 289 -157 290 -151
rect 338 -194 339 -156
rect 366 -157 367 -151
rect 16 -194 17 -158
rect 51 -159 52 -151
rect 86 -159 87 -151
rect 303 -159 304 -151
rect 320 -194 321 -158
rect 366 -194 367 -158
rect 23 -194 24 -160
rect 30 -161 31 -151
rect 37 -194 38 -160
rect 107 -161 108 -151
rect 128 -194 129 -160
rect 198 -161 199 -151
rect 208 -161 209 -151
rect 359 -161 360 -151
rect 30 -194 31 -162
rect 173 -194 174 -162
rect 191 -163 192 -151
rect 373 -194 374 -162
rect 51 -194 52 -164
rect 96 -194 97 -164
rect 107 -194 108 -164
rect 205 -165 206 -151
rect 222 -194 223 -164
rect 387 -194 388 -164
rect 79 -167 80 -151
rect 205 -194 206 -166
rect 226 -167 227 -151
rect 303 -194 304 -166
rect 359 -194 360 -166
rect 408 -194 409 -166
rect 65 -194 66 -168
rect 79 -194 80 -168
rect 86 -194 87 -168
rect 93 -169 94 -151
rect 149 -169 150 -151
rect 184 -169 185 -151
rect 194 -169 195 -151
rect 296 -169 297 -151
rect 89 -171 90 -151
rect 142 -171 143 -151
rect 149 -194 150 -170
rect 296 -194 297 -170
rect 72 -173 73 -151
rect 142 -194 143 -172
rect 152 -173 153 -151
rect 247 -173 248 -151
rect 261 -173 262 -151
rect 415 -194 416 -172
rect 47 -194 48 -174
rect 72 -194 73 -174
rect 156 -175 157 -151
rect 184 -194 185 -174
rect 198 -194 199 -174
rect 310 -194 311 -174
rect 100 -177 101 -151
rect 156 -194 157 -176
rect 163 -177 164 -151
rect 240 -177 241 -151
rect 261 -194 262 -176
rect 282 -177 283 -151
rect 75 -194 76 -178
rect 163 -194 164 -178
rect 166 -194 167 -178
rect 394 -194 395 -178
rect 82 -181 83 -151
rect 240 -194 241 -180
rect 254 -181 255 -151
rect 282 -194 283 -180
rect 82 -194 83 -182
rect 121 -183 122 -151
rect 177 -183 178 -151
rect 191 -194 192 -182
rect 208 -194 209 -182
rect 226 -194 227 -182
rect 233 -183 234 -151
rect 247 -194 248 -182
rect 268 -183 269 -151
rect 317 -183 318 -151
rect 100 -194 101 -184
rect 135 -185 136 -151
rect 152 -194 153 -184
rect 268 -194 269 -184
rect 275 -185 276 -151
rect 289 -194 290 -184
rect 61 -194 62 -186
rect 275 -194 276 -186
rect 114 -189 115 -151
rect 121 -194 122 -188
rect 170 -189 171 -151
rect 177 -194 178 -188
rect 212 -189 213 -151
rect 233 -194 234 -188
rect 44 -191 45 -151
rect 114 -194 115 -190
rect 219 -191 220 -151
rect 254 -194 255 -190
rect 58 -193 59 -151
rect 212 -194 213 -192
rect 219 -194 220 -192
rect 352 -194 353 -192
rect 16 -204 17 -202
rect 72 -253 73 -203
rect 86 -204 87 -202
rect 149 -204 150 -202
rect 166 -204 167 -202
rect 303 -204 304 -202
rect 324 -204 325 -202
rect 324 -253 325 -203
rect 324 -204 325 -202
rect 324 -253 325 -203
rect 331 -204 332 -202
rect 331 -253 332 -203
rect 331 -204 332 -202
rect 331 -253 332 -203
rect 401 -204 402 -202
rect 401 -253 402 -203
rect 401 -204 402 -202
rect 401 -253 402 -203
rect 16 -253 17 -205
rect 180 -253 181 -205
rect 184 -253 185 -205
rect 387 -206 388 -202
rect 23 -253 24 -207
rect 107 -208 108 -202
rect 110 -253 111 -207
rect 198 -208 199 -202
rect 205 -208 206 -202
rect 373 -208 374 -202
rect 44 -210 45 -202
rect 114 -210 115 -202
rect 117 -253 118 -209
rect 275 -210 276 -202
rect 338 -210 339 -202
rect 373 -253 374 -209
rect 44 -253 45 -211
rect 100 -212 101 -202
rect 107 -253 108 -211
rect 303 -253 304 -211
rect 338 -253 339 -211
rect 345 -212 346 -202
rect 54 -253 55 -213
rect 198 -253 199 -213
rect 219 -214 220 -202
rect 415 -214 416 -202
rect 65 -216 66 -202
rect 82 -216 83 -202
rect 86 -253 87 -215
rect 114 -253 115 -215
rect 124 -253 125 -215
rect 128 -216 129 -202
rect 138 -253 139 -215
rect 191 -216 192 -202
rect 240 -216 241 -202
rect 387 -253 388 -215
rect 30 -218 31 -202
rect 128 -253 129 -217
rect 142 -218 143 -202
rect 163 -253 164 -217
rect 170 -253 171 -217
rect 233 -218 234 -202
rect 247 -218 248 -202
rect 247 -253 248 -217
rect 247 -218 248 -202
rect 247 -253 248 -217
rect 275 -253 276 -217
rect 289 -218 290 -202
rect 310 -218 311 -202
rect 415 -253 416 -217
rect 9 -220 10 -202
rect 30 -253 31 -219
rect 37 -220 38 -202
rect 142 -253 143 -219
rect 177 -220 178 -202
rect 233 -253 234 -219
rect 289 -253 290 -219
rect 296 -220 297 -202
rect 345 -253 346 -219
rect 352 -220 353 -202
rect 9 -253 10 -221
rect 75 -222 76 -202
rect 93 -253 94 -221
rect 156 -222 157 -202
rect 187 -222 188 -202
rect 317 -253 318 -221
rect 352 -253 353 -221
rect 359 -222 360 -202
rect 37 -253 38 -223
rect 82 -253 83 -223
rect 96 -253 97 -223
rect 394 -224 395 -202
rect 65 -253 66 -225
rect 79 -253 80 -225
rect 121 -226 122 -202
rect 156 -253 157 -225
rect 187 -253 188 -225
rect 205 -253 206 -225
rect 222 -226 223 -202
rect 240 -253 241 -225
rect 261 -226 262 -202
rect 296 -253 297 -225
rect 359 -253 360 -225
rect 366 -226 367 -202
rect 51 -228 52 -202
rect 222 -253 223 -227
rect 121 -253 122 -229
rect 366 -253 367 -229
rect 135 -232 136 -202
rect 394 -253 395 -231
rect 149 -253 150 -233
rect 177 -253 178 -233
rect 191 -253 192 -233
rect 212 -234 213 -202
rect 201 -236 202 -202
rect 261 -253 262 -235
rect 201 -253 202 -237
rect 380 -238 381 -202
rect 58 -240 59 -202
rect 380 -253 381 -239
rect 58 -253 59 -241
rect 226 -242 227 -202
rect 212 -253 213 -243
rect 254 -244 255 -202
rect 226 -253 227 -245
rect 268 -246 269 -202
rect 254 -253 255 -247
rect 408 -253 409 -247
rect 268 -253 269 -249
rect 282 -250 283 -202
rect 282 -253 283 -251
rect 310 -253 311 -251
rect 12 -263 13 -261
rect 338 -263 339 -261
rect 380 -263 381 -261
rect 436 -302 437 -262
rect 33 -265 34 -261
rect 54 -265 55 -261
rect 61 -302 62 -264
rect 65 -265 66 -261
rect 72 -302 73 -264
rect 107 -302 108 -264
rect 110 -265 111 -261
rect 268 -265 269 -261
rect 282 -302 283 -264
rect 432 -302 433 -264
rect 37 -267 38 -261
rect 65 -302 66 -266
rect 75 -267 76 -261
rect 138 -267 139 -261
rect 149 -267 150 -261
rect 149 -302 150 -266
rect 149 -267 150 -261
rect 149 -302 150 -266
rect 163 -267 164 -261
rect 184 -267 185 -261
rect 226 -267 227 -261
rect 422 -302 423 -266
rect 30 -302 31 -268
rect 163 -302 164 -268
rect 173 -302 174 -268
rect 212 -269 213 -261
rect 240 -269 241 -261
rect 289 -269 290 -261
rect 338 -302 339 -268
rect 345 -269 346 -261
rect 380 -302 381 -268
rect 425 -302 426 -268
rect 37 -302 38 -270
rect 58 -271 59 -261
rect 86 -271 87 -261
rect 114 -302 115 -270
rect 117 -271 118 -261
rect 142 -271 143 -261
rect 177 -302 178 -270
rect 201 -271 202 -261
rect 205 -271 206 -261
rect 226 -302 227 -270
rect 247 -271 248 -261
rect 254 -271 255 -261
rect 268 -302 269 -270
rect 317 -271 318 -261
rect 345 -302 346 -270
rect 373 -271 374 -261
rect 394 -271 395 -261
rect 397 -279 398 -270
rect 51 -302 52 -272
rect 198 -273 199 -261
rect 212 -302 213 -272
rect 296 -273 297 -261
rect 317 -302 318 -272
rect 331 -273 332 -261
rect 366 -273 367 -261
rect 373 -302 374 -272
rect 394 -302 395 -272
rect 415 -273 416 -261
rect 79 -275 80 -261
rect 86 -302 87 -274
rect 96 -275 97 -261
rect 289 -302 290 -274
rect 331 -302 332 -274
rect 352 -275 353 -261
rect 359 -275 360 -261
rect 366 -302 367 -274
rect 401 -275 402 -261
rect 415 -302 416 -274
rect 23 -277 24 -261
rect 79 -302 80 -276
rect 100 -277 101 -261
rect 142 -302 143 -276
rect 180 -277 181 -261
rect 233 -277 234 -261
rect 250 -302 251 -276
rect 387 -277 388 -261
rect 401 -302 402 -276
rect 408 -277 409 -261
rect 23 -302 24 -278
rect 44 -279 45 -261
rect 100 -302 101 -278
rect 156 -279 157 -261
rect 184 -302 185 -278
rect 275 -279 276 -261
rect 408 -302 409 -278
rect 44 -302 45 -280
rect 201 -302 202 -280
rect 205 -302 206 -280
rect 352 -302 353 -280
rect 103 -283 104 -261
rect 170 -283 171 -261
rect 198 -302 199 -282
rect 296 -302 297 -282
rect 128 -285 129 -261
rect 240 -302 241 -284
rect 254 -302 255 -284
rect 261 -285 262 -261
rect 275 -302 276 -284
rect 310 -285 311 -261
rect 16 -287 17 -261
rect 261 -302 262 -286
rect 264 -302 265 -286
rect 310 -302 311 -286
rect 16 -302 17 -288
rect 243 -289 244 -261
rect 128 -302 129 -290
rect 170 -302 171 -290
rect 219 -302 220 -290
rect 247 -302 248 -290
rect 135 -293 136 -261
rect 387 -302 388 -292
rect 93 -302 94 -294
rect 135 -302 136 -294
rect 156 -302 157 -294
rect 191 -295 192 -261
rect 222 -295 223 -261
rect 359 -302 360 -294
rect 166 -302 167 -296
rect 191 -302 192 -296
rect 233 -302 234 -296
rect 303 -297 304 -261
rect 303 -302 304 -298
rect 324 -299 325 -261
rect 124 -302 125 -300
rect 324 -302 325 -300
rect 2 -363 3 -311
rect 173 -312 174 -310
rect 184 -312 185 -310
rect 240 -363 241 -311
rect 243 -312 244 -310
rect 338 -312 339 -310
rect 401 -312 402 -310
rect 429 -363 430 -311
rect 23 -314 24 -310
rect 93 -314 94 -310
rect 100 -363 101 -313
rect 128 -314 129 -310
rect 142 -314 143 -310
rect 205 -314 206 -310
rect 226 -314 227 -310
rect 226 -363 227 -313
rect 226 -314 227 -310
rect 226 -363 227 -313
rect 233 -314 234 -310
rect 261 -363 262 -313
rect 264 -314 265 -310
rect 415 -314 416 -310
rect 26 -363 27 -315
rect 103 -316 104 -310
rect 107 -363 108 -315
rect 415 -363 416 -315
rect 30 -318 31 -310
rect 187 -363 188 -317
rect 191 -318 192 -310
rect 222 -363 223 -317
rect 247 -363 248 -317
rect 254 -318 255 -310
rect 275 -318 276 -310
rect 275 -363 276 -317
rect 275 -318 276 -310
rect 275 -363 276 -317
rect 317 -318 318 -310
rect 338 -363 339 -317
rect 23 -363 24 -319
rect 191 -363 192 -319
rect 198 -320 199 -310
rect 303 -320 304 -310
rect 317 -363 318 -319
rect 324 -320 325 -310
rect 331 -320 332 -310
rect 331 -363 332 -319
rect 331 -320 332 -310
rect 331 -363 332 -319
rect 30 -363 31 -321
rect 373 -322 374 -310
rect 37 -324 38 -310
rect 170 -324 171 -310
rect 198 -363 199 -323
rect 219 -324 220 -310
rect 250 -324 251 -310
rect 380 -324 381 -310
rect 33 -363 34 -325
rect 37 -363 38 -325
rect 40 -363 41 -325
rect 401 -363 402 -325
rect 44 -328 45 -310
rect 124 -328 125 -310
rect 142 -363 143 -327
rect 212 -328 213 -310
rect 254 -363 255 -327
rect 422 -363 423 -327
rect 54 -363 55 -329
rect 303 -363 304 -329
rect 345 -330 346 -310
rect 380 -363 381 -329
rect 58 -363 59 -331
rect 86 -332 87 -310
rect 110 -332 111 -310
rect 128 -363 129 -331
rect 159 -363 160 -331
rect 177 -332 178 -310
rect 296 -332 297 -310
rect 324 -363 325 -331
rect 373 -363 374 -331
rect 387 -332 388 -310
rect 61 -334 62 -310
rect 93 -363 94 -333
rect 110 -363 111 -333
rect 345 -363 346 -333
rect 65 -336 66 -310
rect 205 -363 206 -335
rect 233 -363 234 -335
rect 387 -363 388 -335
rect 65 -363 66 -337
rect 296 -363 297 -337
rect 72 -340 73 -310
rect 436 -340 437 -310
rect 79 -342 80 -310
rect 163 -363 164 -341
rect 394 -342 395 -310
rect 436 -363 437 -341
rect 16 -344 17 -310
rect 79 -363 80 -343
rect 114 -363 115 -343
rect 212 -363 213 -343
rect 366 -344 367 -310
rect 394 -363 395 -343
rect 16 -363 17 -345
rect 68 -363 69 -345
rect 121 -346 122 -310
rect 149 -346 150 -310
rect 359 -346 360 -310
rect 366 -363 367 -345
rect 117 -348 118 -310
rect 121 -363 122 -347
rect 135 -348 136 -310
rect 177 -363 178 -347
rect 352 -348 353 -310
rect 359 -363 360 -347
rect 117 -363 118 -349
rect 408 -350 409 -310
rect 51 -352 52 -310
rect 408 -363 409 -351
rect 51 -363 52 -353
rect 149 -363 150 -353
rect 289 -354 290 -310
rect 352 -363 353 -353
rect 135 -363 136 -355
rect 156 -356 157 -310
rect 289 -363 290 -355
rect 310 -356 311 -310
rect 156 -363 157 -357
rect 268 -358 269 -310
rect 282 -358 283 -310
rect 310 -363 311 -357
rect 268 -363 269 -359
rect 425 -360 426 -310
rect 271 -363 272 -361
rect 282 -363 283 -361
rect 2 -373 3 -371
rect 173 -373 174 -371
rect 201 -412 202 -372
rect 219 -373 220 -371
rect 222 -373 223 -371
rect 359 -373 360 -371
rect 9 -412 10 -374
rect 30 -375 31 -371
rect 37 -375 38 -371
rect 89 -375 90 -371
rect 110 -375 111 -371
rect 366 -375 367 -371
rect 16 -377 17 -371
rect 23 -412 24 -376
rect 26 -377 27 -371
rect 236 -377 237 -371
rect 247 -377 248 -371
rect 257 -377 258 -371
rect 268 -412 269 -376
rect 310 -377 311 -371
rect 317 -377 318 -371
rect 366 -412 367 -376
rect 16 -412 17 -378
rect 51 -412 52 -378
rect 65 -412 66 -378
rect 198 -379 199 -371
rect 226 -379 227 -371
rect 233 -412 234 -378
rect 271 -379 272 -371
rect 394 -379 395 -371
rect 30 -412 31 -380
rect 47 -381 48 -371
rect 68 -381 69 -371
rect 191 -381 192 -371
rect 271 -412 272 -380
rect 289 -381 290 -371
rect 317 -412 318 -380
rect 324 -381 325 -371
rect 338 -381 339 -371
rect 359 -412 360 -380
rect 387 -381 388 -371
rect 394 -412 395 -380
rect 37 -412 38 -382
rect 58 -383 59 -371
rect 79 -383 80 -371
rect 327 -412 328 -382
rect 61 -412 62 -384
rect 79 -412 80 -384
rect 82 -385 83 -371
rect 296 -385 297 -371
rect 86 -387 87 -371
rect 205 -387 206 -371
rect 212 -387 213 -371
rect 289 -412 290 -386
rect 72 -389 73 -371
rect 86 -412 87 -388
rect 110 -412 111 -388
rect 345 -389 346 -371
rect 72 -412 73 -390
rect 100 -391 101 -371
rect 114 -412 115 -390
rect 408 -391 409 -371
rect 100 -412 101 -392
rect 163 -393 164 -371
rect 184 -393 185 -371
rect 219 -412 220 -392
rect 229 -412 230 -392
rect 387 -412 388 -392
rect 408 -412 409 -392
rect 429 -393 430 -371
rect 117 -395 118 -371
rect 415 -395 416 -371
rect 135 -397 136 -371
rect 166 -412 167 -396
rect 205 -412 206 -396
rect 250 -412 251 -396
rect 261 -397 262 -371
rect 338 -412 339 -396
rect 352 -397 353 -371
rect 429 -412 430 -396
rect 135 -412 136 -398
rect 159 -399 160 -371
rect 163 -412 164 -398
rect 310 -412 311 -398
rect 331 -399 332 -371
rect 352 -412 353 -398
rect 415 -412 416 -398
rect 422 -399 423 -371
rect 142 -401 143 -371
rect 191 -412 192 -400
rect 212 -412 213 -400
rect 240 -401 241 -371
rect 261 -412 262 -400
rect 401 -401 402 -371
rect 422 -412 423 -400
rect 436 -401 437 -371
rect 93 -403 94 -371
rect 142 -412 143 -402
rect 149 -403 150 -371
rect 156 -403 157 -371
rect 184 -412 185 -402
rect 240 -412 241 -402
rect 275 -403 276 -371
rect 296 -412 297 -402
rect 303 -403 304 -371
rect 345 -412 346 -402
rect 373 -403 374 -371
rect 401 -412 402 -402
rect 432 -412 433 -402
rect 436 -412 437 -402
rect 54 -412 55 -404
rect 93 -412 94 -404
rect 121 -405 122 -371
rect 149 -412 150 -404
rect 170 -405 171 -371
rect 303 -412 304 -404
rect 373 -412 374 -404
rect 380 -405 381 -371
rect 47 -412 48 -406
rect 121 -412 122 -406
rect 128 -407 129 -371
rect 156 -412 157 -406
rect 170 -412 171 -406
rect 177 -407 178 -371
rect 254 -407 255 -371
rect 275 -412 276 -406
rect 282 -407 283 -371
rect 282 -412 283 -406
rect 282 -407 283 -371
rect 282 -412 283 -406
rect 58 -412 59 -408
rect 177 -412 178 -408
rect 264 -412 265 -408
rect 380 -412 381 -408
rect 117 -412 118 -410
rect 254 -412 255 -410
rect 9 -422 10 -420
rect 51 -422 52 -420
rect 79 -422 80 -420
rect 82 -430 83 -421
rect 107 -422 108 -420
rect 215 -467 216 -421
rect 226 -422 227 -420
rect 345 -422 346 -420
rect 432 -422 433 -420
rect 457 -467 458 -421
rect 16 -424 17 -420
rect 33 -467 34 -423
rect 37 -424 38 -420
rect 37 -467 38 -423
rect 37 -424 38 -420
rect 37 -467 38 -423
rect 44 -424 45 -420
rect 142 -424 143 -420
rect 166 -424 167 -420
rect 170 -424 171 -420
rect 194 -467 195 -423
rect 212 -424 213 -420
rect 229 -467 230 -423
rect 289 -424 290 -420
rect 317 -424 318 -420
rect 345 -467 346 -423
rect 359 -424 360 -420
rect 432 -467 433 -423
rect 443 -424 444 -420
rect 450 -467 451 -423
rect 16 -467 17 -425
rect 26 -467 27 -425
rect 30 -426 31 -420
rect 75 -467 76 -425
rect 79 -467 80 -425
rect 86 -426 87 -420
rect 93 -426 94 -420
rect 107 -467 108 -425
rect 121 -426 122 -420
rect 142 -467 143 -425
rect 163 -426 164 -420
rect 289 -467 290 -425
rect 327 -426 328 -420
rect 422 -426 423 -420
rect 446 -467 447 -425
rect 464 -467 465 -425
rect 51 -467 52 -427
rect 72 -428 73 -420
rect 86 -467 87 -427
rect 100 -428 101 -420
rect 121 -467 122 -427
rect 135 -428 136 -420
rect 156 -428 157 -420
rect 163 -467 164 -427
rect 177 -428 178 -420
rect 317 -467 318 -427
rect 334 -428 335 -420
rect 401 -428 402 -420
rect 58 -467 59 -429
rect 72 -467 73 -429
rect 100 -467 101 -429
rect 114 -467 115 -429
rect 177 -467 178 -429
rect 201 -467 202 -429
rect 338 -430 339 -420
rect 352 -430 353 -420
rect 359 -467 360 -429
rect 93 -467 94 -431
rect 180 -467 181 -431
rect 212 -467 213 -431
rect 233 -432 234 -420
rect 236 -467 237 -431
rect 338 -467 339 -431
rect 128 -434 129 -420
rect 219 -434 220 -420
rect 240 -434 241 -420
rect 422 -467 423 -433
rect 117 -436 118 -420
rect 128 -467 129 -435
rect 131 -436 132 -420
rect 149 -436 150 -420
rect 156 -467 157 -435
rect 191 -436 192 -420
rect 243 -467 244 -435
rect 303 -436 304 -420
rect 135 -467 136 -437
rect 184 -438 185 -420
rect 191 -467 192 -437
rect 436 -438 437 -420
rect 149 -467 150 -439
rect 198 -467 199 -439
rect 247 -440 248 -420
rect 296 -440 297 -420
rect 387 -440 388 -420
rect 436 -467 437 -439
rect 226 -467 227 -441
rect 296 -467 297 -441
rect 387 -467 388 -441
rect 408 -442 409 -420
rect 250 -444 251 -420
rect 394 -444 395 -420
rect 250 -467 251 -445
rect 415 -446 416 -420
rect 254 -448 255 -420
rect 303 -467 304 -447
rect 310 -448 311 -420
rect 415 -467 416 -447
rect 254 -467 255 -449
rect 352 -467 353 -449
rect 373 -450 374 -420
rect 394 -467 395 -449
rect 257 -467 258 -451
rect 366 -452 367 -420
rect 373 -467 374 -451
rect 380 -452 381 -420
rect 261 -454 262 -420
rect 331 -467 332 -453
rect 170 -467 171 -455
rect 261 -467 262 -455
rect 268 -456 269 -420
rect 380 -467 381 -455
rect 65 -458 66 -420
rect 268 -467 269 -457
rect 275 -458 276 -420
rect 310 -467 311 -457
rect 324 -458 325 -420
rect 366 -467 367 -457
rect 47 -460 48 -420
rect 275 -467 276 -459
rect 282 -460 283 -420
rect 324 -467 325 -459
rect 65 -467 66 -461
rect 205 -462 206 -420
rect 184 -467 185 -463
rect 282 -467 283 -463
rect 205 -467 206 -465
rect 222 -467 223 -465
rect 9 -508 10 -476
rect 124 -508 125 -476
rect 142 -477 143 -475
rect 233 -508 234 -476
rect 247 -477 248 -475
rect 254 -508 255 -476
rect 261 -477 262 -475
rect 317 -477 318 -475
rect 352 -477 353 -475
rect 401 -508 402 -476
rect 418 -508 419 -476
rect 450 -477 451 -475
rect 464 -477 465 -475
rect 464 -508 465 -476
rect 464 -477 465 -475
rect 464 -508 465 -476
rect 30 -508 31 -478
rect 236 -479 237 -475
rect 250 -479 251 -475
rect 338 -479 339 -475
rect 345 -479 346 -475
rect 352 -508 353 -478
rect 373 -479 374 -475
rect 373 -508 374 -478
rect 373 -479 374 -475
rect 373 -508 374 -478
rect 387 -479 388 -475
rect 408 -508 409 -478
rect 422 -479 423 -475
rect 446 -479 447 -475
rect 33 -508 34 -480
rect 215 -508 216 -480
rect 222 -481 223 -475
rect 415 -481 416 -475
rect 432 -508 433 -480
rect 436 -481 437 -475
rect 37 -483 38 -475
rect 128 -483 129 -475
rect 131 -483 132 -475
rect 345 -508 346 -482
rect 380 -483 381 -475
rect 387 -508 388 -482
rect 415 -508 416 -482
rect 450 -508 451 -482
rect 16 -485 17 -475
rect 37 -508 38 -484
rect 40 -508 41 -484
rect 58 -485 59 -475
rect 72 -485 73 -475
rect 93 -485 94 -475
rect 100 -485 101 -475
rect 142 -508 143 -484
rect 173 -508 174 -484
rect 198 -508 199 -484
rect 205 -485 206 -475
rect 261 -508 262 -484
rect 264 -485 265 -475
rect 310 -485 311 -475
rect 359 -485 360 -475
rect 380 -508 381 -484
rect 16 -508 17 -486
rect 23 -508 24 -486
rect 44 -508 45 -486
rect 138 -508 139 -486
rect 180 -487 181 -475
rect 429 -487 430 -475
rect 51 -489 52 -475
rect 103 -508 104 -488
rect 107 -489 108 -475
rect 226 -508 227 -488
rect 240 -508 241 -488
rect 436 -508 437 -488
rect 51 -508 52 -490
rect 72 -508 73 -490
rect 82 -508 83 -490
rect 177 -508 178 -490
rect 191 -491 192 -475
rect 219 -508 220 -490
rect 275 -491 276 -475
rect 282 -491 283 -475
rect 285 -491 286 -475
rect 394 -491 395 -475
rect 429 -508 430 -490
rect 457 -491 458 -475
rect 58 -508 59 -492
rect 79 -493 80 -475
rect 93 -508 94 -492
rect 110 -493 111 -475
rect 114 -493 115 -475
rect 114 -508 115 -492
rect 114 -493 115 -475
rect 114 -508 115 -492
rect 128 -508 129 -492
rect 135 -493 136 -475
rect 184 -493 185 -475
rect 191 -508 192 -492
rect 212 -493 213 -475
rect 247 -508 248 -492
rect 296 -493 297 -475
rect 317 -508 318 -492
rect 359 -508 360 -492
rect 366 -493 367 -475
rect 443 -508 444 -492
rect 457 -508 458 -492
rect 79 -508 80 -494
rect 331 -495 332 -475
rect 107 -508 108 -496
rect 121 -497 122 -475
rect 156 -497 157 -475
rect 184 -508 185 -496
rect 268 -497 269 -475
rect 331 -508 332 -496
rect 121 -508 122 -498
rect 163 -499 164 -475
rect 170 -499 171 -475
rect 268 -508 269 -498
rect 289 -499 290 -475
rect 296 -508 297 -498
rect 303 -499 304 -475
rect 338 -508 339 -498
rect 65 -501 66 -475
rect 289 -508 290 -500
rect 310 -508 311 -500
rect 324 -501 325 -475
rect 65 -508 66 -502
rect 86 -503 87 -475
rect 156 -508 157 -502
rect 194 -503 195 -475
rect 243 -508 244 -502
rect 324 -508 325 -502
rect 86 -508 87 -504
rect 149 -505 150 -475
rect 163 -508 164 -504
rect 303 -508 304 -504
rect 149 -508 150 -506
rect 205 -508 206 -506
rect 9 -518 10 -516
rect 68 -561 69 -517
rect 72 -518 73 -516
rect 93 -518 94 -516
rect 117 -561 118 -517
rect 124 -518 125 -516
rect 138 -518 139 -516
rect 436 -518 437 -516
rect 9 -561 10 -519
rect 103 -520 104 -516
rect 121 -520 122 -516
rect 226 -520 227 -516
rect 243 -520 244 -516
rect 254 -520 255 -516
rect 278 -520 279 -516
rect 352 -520 353 -516
rect 366 -520 367 -516
rect 422 -561 423 -519
rect 429 -561 430 -519
rect 443 -520 444 -516
rect 16 -522 17 -516
rect 37 -522 38 -516
rect 44 -522 45 -516
rect 205 -522 206 -516
rect 208 -522 209 -516
rect 338 -522 339 -516
rect 401 -522 402 -516
rect 415 -522 416 -516
rect 443 -561 444 -521
rect 457 -522 458 -516
rect 19 -561 20 -523
rect 275 -524 276 -516
rect 285 -561 286 -523
rect 380 -524 381 -516
rect 457 -561 458 -523
rect 464 -524 465 -516
rect 37 -561 38 -525
rect 156 -526 157 -516
rect 166 -561 167 -525
rect 254 -561 255 -525
rect 303 -526 304 -516
rect 408 -526 409 -516
rect 450 -526 451 -516
rect 464 -561 465 -525
rect 44 -561 45 -527
rect 51 -528 52 -516
rect 58 -528 59 -516
rect 96 -561 97 -527
rect 124 -561 125 -527
rect 173 -528 174 -516
rect 184 -528 185 -516
rect 205 -561 206 -527
rect 212 -528 213 -516
rect 331 -528 332 -516
rect 359 -528 360 -516
rect 380 -561 381 -527
rect 30 -530 31 -516
rect 58 -561 59 -529
rect 72 -561 73 -529
rect 170 -561 171 -529
rect 173 -561 174 -529
rect 436 -561 437 -529
rect 30 -561 31 -531
rect 93 -561 94 -531
rect 149 -532 150 -516
rect 187 -561 188 -531
rect 212 -561 213 -531
rect 268 -532 269 -516
rect 306 -532 307 -516
rect 341 -561 342 -531
rect 373 -532 374 -516
rect 415 -561 416 -531
rect 26 -561 27 -533
rect 268 -561 269 -533
rect 310 -534 311 -516
rect 352 -561 353 -533
rect 373 -561 374 -533
rect 432 -534 433 -516
rect 51 -561 52 -535
rect 65 -536 66 -516
rect 82 -536 83 -516
rect 366 -561 367 -535
rect 40 -538 41 -516
rect 65 -561 66 -537
rect 82 -561 83 -537
rect 282 -538 283 -516
rect 324 -538 325 -516
rect 394 -561 395 -537
rect 86 -540 87 -516
rect 156 -561 157 -539
rect 184 -561 185 -539
rect 359 -561 360 -539
rect 86 -561 87 -541
rect 107 -542 108 -516
rect 149 -561 150 -541
rect 163 -542 164 -516
rect 198 -542 199 -516
rect 310 -561 311 -541
rect 331 -561 332 -541
rect 345 -542 346 -516
rect 107 -561 108 -543
rect 128 -544 129 -516
rect 163 -561 164 -543
rect 177 -544 178 -516
rect 219 -544 220 -516
rect 226 -561 227 -543
rect 233 -544 234 -516
rect 408 -561 409 -543
rect 103 -561 104 -545
rect 128 -561 129 -545
rect 135 -561 136 -545
rect 177 -561 178 -545
rect 191 -546 192 -516
rect 219 -561 220 -545
rect 233 -561 234 -545
rect 387 -546 388 -516
rect 114 -548 115 -516
rect 198 -561 199 -547
rect 240 -561 241 -547
rect 387 -561 388 -547
rect 191 -561 192 -549
rect 215 -550 216 -516
rect 247 -550 248 -516
rect 275 -561 276 -549
rect 282 -561 283 -549
rect 401 -561 402 -549
rect 247 -561 248 -551
rect 261 -552 262 -516
rect 296 -552 297 -516
rect 324 -561 325 -551
rect 23 -561 24 -553
rect 296 -561 297 -553
rect 317 -554 318 -516
rect 345 -561 346 -553
rect 236 -561 237 -555
rect 261 -561 262 -555
rect 289 -556 290 -516
rect 317 -561 318 -555
rect 142 -558 143 -516
rect 289 -561 290 -557
rect 114 -561 115 -559
rect 142 -561 143 -559
rect 9 -571 10 -569
rect 184 -614 185 -570
rect 198 -571 199 -569
rect 198 -614 199 -570
rect 198 -571 199 -569
rect 198 -614 199 -570
rect 212 -571 213 -569
rect 264 -614 265 -570
rect 303 -571 304 -569
rect 345 -571 346 -569
rect 415 -571 416 -569
rect 415 -614 416 -570
rect 415 -571 416 -569
rect 415 -614 416 -570
rect 422 -571 423 -569
rect 422 -614 423 -570
rect 422 -571 423 -569
rect 422 -614 423 -570
rect 443 -571 444 -569
rect 443 -614 444 -570
rect 443 -571 444 -569
rect 443 -614 444 -570
rect 464 -571 465 -569
rect 471 -614 472 -570
rect 16 -573 17 -569
rect 100 -614 101 -572
rect 121 -573 122 -569
rect 121 -614 122 -572
rect 121 -573 122 -569
rect 121 -614 122 -572
rect 138 -614 139 -572
rect 303 -614 304 -572
rect 341 -573 342 -569
rect 394 -573 395 -569
rect 457 -614 458 -572
rect 464 -614 465 -572
rect 16 -614 17 -574
rect 114 -614 115 -574
rect 163 -575 164 -569
rect 446 -614 447 -574
rect 23 -614 24 -576
rect 128 -577 129 -569
rect 163 -614 164 -576
rect 208 -577 209 -569
rect 226 -577 227 -569
rect 226 -614 227 -576
rect 226 -577 227 -569
rect 226 -614 227 -576
rect 233 -577 234 -569
rect 247 -577 248 -569
rect 257 -614 258 -576
rect 401 -577 402 -569
rect 9 -614 10 -578
rect 208 -614 209 -578
rect 236 -579 237 -569
rect 366 -579 367 -569
rect 394 -614 395 -578
rect 429 -579 430 -569
rect 30 -581 31 -569
rect 103 -581 104 -569
rect 170 -581 171 -569
rect 282 -581 283 -569
rect 33 -614 34 -582
rect 44 -583 45 -569
rect 58 -583 59 -569
rect 89 -614 90 -582
rect 93 -583 94 -569
rect 243 -583 244 -569
rect 247 -614 248 -582
rect 317 -583 318 -569
rect 40 -614 41 -584
rect 429 -614 430 -584
rect 44 -614 45 -586
rect 51 -587 52 -569
rect 58 -614 59 -586
rect 107 -587 108 -569
rect 149 -587 150 -569
rect 282 -614 283 -586
rect 317 -614 318 -586
rect 331 -587 332 -569
rect 37 -589 38 -569
rect 51 -614 52 -588
rect 65 -614 66 -588
rect 156 -589 157 -569
rect 173 -589 174 -569
rect 219 -589 220 -569
rect 240 -589 241 -569
rect 352 -589 353 -569
rect 68 -591 69 -569
rect 345 -614 346 -590
rect 352 -614 353 -590
rect 359 -591 360 -569
rect 79 -593 80 -569
rect 289 -593 290 -569
rect 331 -614 332 -592
rect 366 -614 367 -592
rect 72 -595 73 -569
rect 79 -614 80 -594
rect 93 -614 94 -594
rect 436 -595 437 -569
rect 30 -614 31 -596
rect 436 -614 437 -596
rect 72 -614 73 -598
rect 86 -599 87 -569
rect 107 -614 108 -598
rect 194 -614 195 -598
rect 205 -599 206 -569
rect 233 -614 234 -598
rect 240 -614 241 -598
rect 268 -599 269 -569
rect 289 -614 290 -598
rect 324 -599 325 -569
rect 359 -614 360 -598
rect 380 -599 381 -569
rect 86 -614 87 -600
rect 142 -601 143 -569
rect 156 -614 157 -600
rect 173 -614 174 -600
rect 177 -614 178 -600
rect 191 -601 192 -569
rect 219 -614 220 -600
rect 275 -601 276 -569
rect 306 -601 307 -569
rect 380 -614 381 -600
rect 135 -603 136 -569
rect 149 -614 150 -602
rect 180 -603 181 -569
rect 408 -603 409 -569
rect 142 -614 143 -604
rect 170 -614 171 -604
rect 254 -605 255 -569
rect 401 -614 402 -604
rect 268 -614 269 -606
rect 310 -607 311 -569
rect 338 -607 339 -569
rect 408 -614 409 -606
rect 261 -609 262 -569
rect 310 -614 311 -608
rect 338 -614 339 -608
rect 373 -609 374 -569
rect 275 -614 276 -610
rect 296 -611 297 -569
rect 373 -614 374 -610
rect 387 -611 388 -569
rect 296 -614 297 -612
rect 324 -614 325 -612
rect 387 -614 388 -612
rect 453 -614 454 -612
rect 2 -665 3 -623
rect 51 -624 52 -622
rect 72 -624 73 -622
rect 114 -624 115 -622
rect 117 -624 118 -622
rect 212 -624 213 -622
rect 222 -665 223 -623
rect 268 -624 269 -622
rect 299 -624 300 -622
rect 422 -624 423 -622
rect 436 -624 437 -622
rect 443 -665 444 -623
rect 450 -624 451 -622
rect 457 -624 458 -622
rect 460 -665 461 -623
rect 464 -665 465 -623
rect 471 -624 472 -622
rect 471 -665 472 -623
rect 471 -624 472 -622
rect 471 -665 472 -623
rect 9 -626 10 -622
rect 103 -626 104 -622
rect 170 -626 171 -622
rect 184 -626 185 -622
rect 187 -665 188 -625
rect 282 -626 283 -622
rect 299 -665 300 -625
rect 415 -626 416 -622
rect 429 -626 430 -622
rect 436 -665 437 -625
rect 9 -665 10 -627
rect 75 -665 76 -627
rect 79 -628 80 -622
rect 131 -628 132 -622
rect 142 -628 143 -622
rect 170 -665 171 -627
rect 191 -628 192 -622
rect 215 -628 216 -622
rect 233 -628 234 -622
rect 422 -665 423 -627
rect 23 -630 24 -622
rect 135 -630 136 -622
rect 142 -665 143 -629
rect 226 -630 227 -622
rect 240 -630 241 -622
rect 254 -630 255 -622
rect 261 -630 262 -622
rect 352 -630 353 -622
rect 373 -630 374 -622
rect 373 -665 374 -629
rect 373 -630 374 -622
rect 373 -665 374 -629
rect 380 -630 381 -622
rect 429 -665 430 -629
rect 16 -632 17 -622
rect 23 -665 24 -631
rect 30 -665 31 -631
rect 163 -632 164 -622
rect 194 -632 195 -622
rect 401 -632 402 -622
rect 415 -665 416 -631
rect 446 -632 447 -622
rect 16 -665 17 -633
rect 65 -634 66 -622
rect 93 -634 94 -622
rect 96 -650 97 -633
rect 128 -634 129 -622
rect 194 -665 195 -633
rect 205 -665 206 -633
rect 303 -634 304 -622
rect 310 -634 311 -622
rect 310 -665 311 -633
rect 310 -634 311 -622
rect 310 -665 311 -633
rect 331 -634 332 -622
rect 359 -634 360 -622
rect 33 -636 34 -622
rect 65 -665 66 -635
rect 86 -665 87 -635
rect 128 -665 129 -635
rect 135 -665 136 -635
rect 149 -636 150 -622
rect 208 -636 209 -622
rect 387 -636 388 -622
rect 37 -638 38 -622
rect 198 -638 199 -622
rect 215 -665 216 -637
rect 282 -665 283 -637
rect 289 -638 290 -622
rect 303 -665 304 -637
rect 331 -665 332 -637
rect 352 -665 353 -637
rect 387 -665 388 -637
rect 394 -638 395 -622
rect 37 -665 38 -639
rect 177 -640 178 -622
rect 180 -665 181 -639
rect 394 -665 395 -639
rect 40 -642 41 -622
rect 271 -665 272 -641
rect 334 -642 335 -622
rect 408 -642 409 -622
rect 44 -644 45 -622
rect 51 -665 52 -643
rect 54 -665 55 -643
rect 450 -665 451 -643
rect 44 -665 45 -645
rect 275 -646 276 -622
rect 345 -646 346 -622
rect 380 -665 381 -645
rect 58 -648 59 -622
rect 79 -665 80 -647
rect 93 -665 94 -647
rect 121 -648 122 -622
rect 156 -648 157 -622
rect 198 -665 199 -647
rect 219 -648 220 -622
rect 233 -665 234 -647
rect 243 -665 244 -647
rect 359 -665 360 -647
rect 366 -648 367 -622
rect 408 -665 409 -647
rect 58 -665 59 -649
rect 89 -650 90 -622
rect 121 -665 122 -649
rect 163 -665 164 -649
rect 208 -665 209 -649
rect 226 -665 227 -649
rect 247 -665 248 -649
rect 254 -665 255 -649
rect 457 -665 458 -649
rect 107 -652 108 -622
rect 149 -665 150 -651
rect 184 -665 185 -651
rect 289 -665 290 -651
rect 324 -652 325 -622
rect 366 -665 367 -651
rect 100 -654 101 -622
rect 107 -665 108 -653
rect 114 -665 115 -653
rect 177 -665 178 -653
rect 240 -665 241 -653
rect 324 -665 325 -653
rect 338 -654 339 -622
rect 345 -665 346 -653
rect 100 -665 101 -655
rect 156 -665 157 -655
rect 261 -665 262 -655
rect 317 -656 318 -622
rect 103 -665 104 -657
rect 338 -665 339 -657
rect 250 -660 251 -622
rect 317 -665 318 -659
rect 250 -665 251 -661
rect 401 -665 402 -661
rect 275 -665 276 -663
rect 296 -665 297 -663
rect 2 -675 3 -673
rect 131 -675 132 -673
rect 135 -675 136 -673
rect 180 -675 181 -673
rect 187 -716 188 -674
rect 219 -675 220 -673
rect 233 -675 234 -673
rect 240 -675 241 -673
rect 250 -675 251 -673
rect 303 -675 304 -673
rect 331 -716 332 -674
rect 338 -675 339 -673
rect 387 -675 388 -673
rect 387 -716 388 -674
rect 387 -675 388 -673
rect 387 -716 388 -674
rect 443 -675 444 -673
rect 457 -675 458 -673
rect 464 -675 465 -673
rect 471 -675 472 -673
rect 16 -677 17 -673
rect 100 -677 101 -673
rect 114 -677 115 -673
rect 149 -677 150 -673
rect 170 -677 171 -673
rect 173 -716 174 -676
rect 191 -677 192 -673
rect 317 -677 318 -673
rect 334 -677 335 -673
rect 429 -677 430 -673
rect 9 -679 10 -673
rect 16 -716 17 -678
rect 37 -679 38 -673
rect 177 -679 178 -673
rect 191 -716 192 -678
rect 226 -679 227 -673
rect 250 -716 251 -678
rect 436 -679 437 -673
rect 9 -716 10 -680
rect 93 -681 94 -673
rect 128 -681 129 -673
rect 401 -681 402 -673
rect 23 -683 24 -673
rect 93 -716 94 -682
rect 149 -716 150 -682
rect 240 -716 241 -682
rect 268 -683 269 -673
rect 317 -716 318 -682
rect 380 -683 381 -673
rect 429 -716 430 -682
rect 23 -716 24 -684
rect 289 -685 290 -673
rect 296 -716 297 -684
rect 366 -685 367 -673
rect 380 -716 381 -684
rect 408 -685 409 -673
rect 37 -716 38 -686
rect 205 -716 206 -686
rect 212 -687 213 -673
rect 422 -687 423 -673
rect 40 -716 41 -688
rect 131 -716 132 -688
rect 170 -716 171 -688
rect 212 -716 213 -688
rect 229 -716 230 -688
rect 289 -716 290 -688
rect 299 -689 300 -673
rect 345 -689 346 -673
rect 359 -689 360 -673
rect 366 -716 367 -688
rect 401 -716 402 -688
rect 415 -689 416 -673
rect 44 -716 45 -690
rect 86 -691 87 -673
rect 177 -716 178 -690
rect 282 -691 283 -673
rect 345 -716 346 -690
rect 352 -691 353 -673
rect 359 -716 360 -690
rect 373 -691 374 -673
rect 51 -716 52 -692
rect 352 -716 353 -692
rect 58 -695 59 -673
rect 135 -716 136 -694
rect 194 -695 195 -673
rect 219 -716 220 -694
rect 268 -716 269 -694
rect 310 -695 311 -673
rect 58 -716 59 -696
rect 254 -697 255 -673
rect 261 -697 262 -673
rect 310 -716 311 -696
rect 72 -699 73 -673
rect 100 -716 101 -698
rect 198 -699 199 -673
rect 215 -699 216 -673
rect 254 -716 255 -698
rect 275 -699 276 -673
rect 282 -716 283 -698
rect 324 -699 325 -673
rect 2 -716 3 -700
rect 72 -716 73 -700
rect 75 -716 76 -700
rect 184 -701 185 -673
rect 261 -716 262 -700
rect 373 -716 374 -700
rect 79 -703 80 -673
rect 114 -716 115 -702
rect 142 -703 143 -673
rect 198 -716 199 -702
rect 324 -716 325 -702
rect 394 -703 395 -673
rect 82 -716 83 -704
rect 107 -705 108 -673
rect 142 -716 143 -704
rect 156 -705 157 -673
rect 184 -716 185 -704
rect 233 -716 234 -704
rect 394 -716 395 -704
rect 450 -705 451 -673
rect 65 -707 66 -673
rect 107 -716 108 -706
rect 156 -716 157 -706
rect 163 -707 164 -673
rect 54 -709 55 -673
rect 65 -716 66 -708
rect 86 -716 87 -708
rect 124 -716 125 -708
rect 121 -711 122 -673
rect 163 -716 164 -710
rect 30 -713 31 -673
rect 121 -716 122 -712
rect 30 -716 31 -714
rect 117 -715 118 -673
rect 9 -726 10 -724
rect 72 -769 73 -725
rect 96 -769 97 -725
rect 184 -726 185 -724
rect 198 -726 199 -724
rect 352 -726 353 -724
rect 376 -726 377 -724
rect 401 -726 402 -724
rect 411 -726 412 -724
rect 429 -726 430 -724
rect 16 -728 17 -724
rect 75 -728 76 -724
rect 110 -769 111 -727
rect 250 -728 251 -724
rect 254 -728 255 -724
rect 278 -728 279 -724
rect 289 -728 290 -724
rect 296 -728 297 -724
rect 338 -769 339 -727
rect 380 -728 381 -724
rect 387 -728 388 -724
rect 408 -769 409 -727
rect 23 -730 24 -724
rect 198 -769 199 -729
rect 215 -769 216 -729
rect 233 -730 234 -724
rect 243 -730 244 -724
rect 310 -730 311 -724
rect 341 -730 342 -724
rect 345 -730 346 -724
rect 2 -732 3 -724
rect 310 -769 311 -731
rect 345 -769 346 -731
rect 359 -732 360 -724
rect 23 -769 24 -733
rect 86 -734 87 -724
rect 121 -769 122 -733
rect 303 -769 304 -733
rect 37 -736 38 -724
rect 79 -769 80 -735
rect 86 -769 87 -735
rect 191 -736 192 -724
rect 233 -769 234 -735
rect 268 -736 269 -724
rect 289 -769 290 -735
rect 324 -736 325 -724
rect 37 -769 38 -737
rect 180 -738 181 -724
rect 205 -738 206 -724
rect 268 -769 269 -737
rect 324 -769 325 -737
rect 394 -738 395 -724
rect 40 -769 41 -739
rect 58 -740 59 -724
rect 65 -740 66 -724
rect 75 -769 76 -739
rect 128 -740 129 -724
rect 254 -769 255 -739
rect 16 -769 17 -741
rect 58 -769 59 -741
rect 114 -742 115 -724
rect 128 -769 129 -741
rect 135 -742 136 -724
rect 184 -769 185 -741
rect 247 -769 248 -741
rect 282 -742 283 -724
rect 44 -744 45 -724
rect 191 -769 192 -743
rect 236 -769 237 -743
rect 282 -769 283 -743
rect 44 -769 45 -745
rect 65 -769 66 -745
rect 93 -746 94 -724
rect 135 -769 136 -745
rect 142 -746 143 -724
rect 208 -746 209 -724
rect 51 -769 52 -747
rect 82 -748 83 -724
rect 100 -748 101 -724
rect 142 -769 143 -747
rect 149 -748 150 -724
rect 149 -769 150 -747
rect 149 -748 150 -724
rect 149 -769 150 -747
rect 156 -748 157 -724
rect 201 -748 202 -724
rect 54 -750 55 -724
rect 240 -769 241 -749
rect 82 -769 83 -751
rect 114 -769 115 -751
rect 163 -752 164 -724
rect 170 -769 171 -751
rect 180 -769 181 -751
rect 317 -752 318 -724
rect 100 -769 101 -753
rect 261 -754 262 -724
rect 30 -756 31 -724
rect 261 -769 262 -755
rect 103 -769 104 -757
rect 208 -769 209 -757
rect 107 -760 108 -724
rect 156 -769 157 -759
rect 163 -769 164 -759
rect 226 -760 227 -724
rect 219 -762 220 -724
rect 226 -769 227 -761
rect 212 -764 213 -724
rect 219 -769 220 -763
rect 212 -769 213 -765
rect 331 -766 332 -724
rect 331 -769 332 -767
rect 366 -768 367 -724
rect 9 -814 10 -778
rect 47 -779 48 -777
rect 58 -779 59 -777
rect 107 -779 108 -777
rect 110 -814 111 -778
rect 156 -779 157 -777
rect 177 -779 178 -777
rect 303 -779 304 -777
rect 317 -814 318 -778
rect 338 -779 339 -777
rect 30 -781 31 -777
rect 51 -781 52 -777
rect 65 -781 66 -777
rect 75 -781 76 -777
rect 93 -781 94 -777
rect 142 -781 143 -777
rect 177 -814 178 -780
rect 226 -781 227 -777
rect 233 -814 234 -780
rect 261 -781 262 -777
rect 268 -781 269 -777
rect 268 -814 269 -780
rect 268 -781 269 -777
rect 268 -814 269 -780
rect 51 -814 52 -782
rect 79 -814 80 -782
rect 96 -783 97 -777
rect 254 -783 255 -777
rect 72 -814 73 -784
rect 82 -814 83 -784
rect 100 -814 101 -784
rect 152 -814 153 -784
rect 163 -785 164 -777
rect 261 -814 262 -784
rect 103 -787 104 -777
rect 303 -814 304 -786
rect 107 -814 108 -788
rect 240 -789 241 -777
rect 247 -789 248 -777
rect 275 -789 276 -777
rect 30 -814 31 -790
rect 247 -814 248 -790
rect 254 -814 255 -790
rect 282 -791 283 -777
rect 117 -793 118 -777
rect 170 -793 171 -777
rect 198 -793 199 -777
rect 198 -814 199 -792
rect 198 -793 199 -777
rect 198 -814 199 -792
rect 205 -814 206 -792
rect 212 -793 213 -777
rect 219 -793 220 -777
rect 226 -814 227 -792
rect 282 -814 283 -792
rect 289 -793 290 -777
rect 23 -795 24 -777
rect 170 -814 171 -794
rect 212 -814 213 -794
rect 236 -795 237 -777
rect 23 -814 24 -796
rect 61 -814 62 -796
rect 124 -797 125 -777
rect 135 -797 136 -777
rect 163 -814 164 -796
rect 191 -797 192 -777
rect 33 -799 34 -777
rect 135 -814 136 -798
rect 149 -799 150 -777
rect 191 -814 192 -798
rect 33 -814 34 -800
rect 117 -814 118 -800
rect 124 -814 125 -800
rect 184 -801 185 -777
rect 37 -803 38 -777
rect 289 -814 290 -802
rect 37 -814 38 -804
rect 114 -814 115 -804
rect 128 -805 129 -777
rect 156 -814 157 -804
rect 86 -807 87 -777
rect 184 -814 185 -806
rect 131 -814 132 -808
rect 310 -809 311 -777
rect 310 -814 311 -810
rect 324 -811 325 -777
rect 324 -814 325 -812
rect 345 -813 346 -777
rect 9 -824 10 -822
rect 16 -824 17 -822
rect 23 -824 24 -822
rect 65 -824 66 -822
rect 72 -824 73 -822
rect 93 -847 94 -823
rect 96 -824 97 -822
rect 233 -824 234 -822
rect 240 -824 241 -822
rect 268 -824 269 -822
rect 282 -824 283 -822
rect 282 -847 283 -823
rect 282 -824 283 -822
rect 282 -847 283 -823
rect 292 -847 293 -823
rect 317 -824 318 -822
rect 324 -824 325 -822
rect 345 -824 346 -822
rect 23 -847 24 -825
rect 261 -826 262 -822
rect 310 -826 311 -822
rect 327 -847 328 -825
rect 33 -828 34 -822
rect 47 -828 48 -822
rect 58 -847 59 -827
rect 79 -847 80 -827
rect 86 -847 87 -827
rect 114 -828 115 -822
rect 117 -828 118 -822
rect 191 -828 192 -822
rect 222 -828 223 -822
rect 226 -828 227 -822
rect 254 -828 255 -822
rect 268 -847 269 -827
rect 37 -830 38 -822
rect 89 -830 90 -822
rect 117 -847 118 -829
rect 289 -830 290 -822
rect 33 -847 34 -831
rect 37 -847 38 -831
rect 72 -847 73 -831
rect 100 -832 101 -822
rect 124 -847 125 -831
rect 163 -832 164 -822
rect 184 -832 185 -822
rect 184 -847 185 -831
rect 184 -832 185 -822
rect 184 -847 185 -831
rect 191 -847 192 -831
rect 247 -832 248 -822
rect 51 -834 52 -822
rect 163 -847 164 -833
rect 212 -834 213 -822
rect 226 -847 227 -833
rect 44 -836 45 -822
rect 51 -847 52 -835
rect 128 -836 129 -822
rect 156 -836 157 -822
rect 205 -836 206 -822
rect 212 -847 213 -835
rect 19 -847 20 -837
rect 44 -847 45 -837
rect 135 -838 136 -822
rect 180 -838 181 -822
rect 135 -847 136 -839
rect 145 -840 146 -822
rect 149 -847 150 -839
rect 198 -840 199 -822
rect 152 -842 153 -822
rect 303 -842 304 -822
rect 156 -847 157 -843
rect 170 -844 171 -822
rect 170 -847 171 -845
rect 289 -847 290 -845
rect 23 -857 24 -855
rect 142 -857 143 -855
rect 187 -857 188 -855
rect 191 -857 192 -855
rect 268 -857 269 -855
rect 285 -857 286 -855
rect 37 -859 38 -855
rect 44 -859 45 -855
rect 47 -859 48 -855
rect 58 -859 59 -855
rect 65 -859 66 -855
rect 86 -859 87 -855
rect 93 -859 94 -855
rect 114 -859 115 -855
rect 131 -859 132 -855
rect 149 -859 150 -855
rect 54 -861 55 -855
rect 170 -861 171 -855
rect 72 -863 73 -855
rect 103 -863 104 -855
rect 107 -863 108 -855
rect 156 -863 157 -855
rect 82 -865 83 -855
rect 163 -865 164 -855
<< labels >>
rlabel pdiffusion 3 -10 3 -10 0 cellNo=17
rlabel pdiffusion 10 -10 10 -10 0 cellNo=8
rlabel pdiffusion 17 -10 17 -10 0 cellNo=25
rlabel pdiffusion 24 -10 24 -10 0 cellNo=156
rlabel pdiffusion 31 -10 31 -10 0 cellNo=63
rlabel pdiffusion 38 -10 38 -10 0 cellNo=328
rlabel pdiffusion 45 -10 45 -10 0 cellNo=114
rlabel pdiffusion 52 -10 52 -10 0 cellNo=226
rlabel pdiffusion 59 -10 59 -10 0 cellNo=208
rlabel pdiffusion 66 -10 66 -10 0 feedthrough
rlabel pdiffusion 73 -10 73 -10 0 cellNo=199
rlabel pdiffusion 80 -10 80 -10 0 cellNo=355
rlabel pdiffusion 87 -10 87 -10 0 cellNo=102
rlabel pdiffusion 94 -10 94 -10 0 cellNo=99
rlabel pdiffusion 101 -10 101 -10 0 cellNo=154
rlabel pdiffusion 108 -10 108 -10 0 feedthrough
rlabel pdiffusion 115 -10 115 -10 0 cellNo=183
rlabel pdiffusion 122 -10 122 -10 0 cellNo=46
rlabel pdiffusion 129 -10 129 -10 0 feedthrough
rlabel pdiffusion 136 -10 136 -10 0 cellNo=274
rlabel pdiffusion 143 -10 143 -10 0 cellNo=325
rlabel pdiffusion 150 -10 150 -10 0 feedthrough
rlabel pdiffusion 157 -10 157 -10 0 cellNo=261
rlabel pdiffusion 164 -10 164 -10 0 feedthrough
rlabel pdiffusion 3 -29 3 -29 0 cellNo=35
rlabel pdiffusion 10 -29 10 -29 0 cellNo=21
rlabel pdiffusion 17 -29 17 -29 0 cellNo=221
rlabel pdiffusion 24 -29 24 -29 0 cellNo=69
rlabel pdiffusion 31 -29 31 -29 0 cellNo=96
rlabel pdiffusion 38 -29 38 -29 0 cellNo=91
rlabel pdiffusion 45 -29 45 -29 0 cellNo=82
rlabel pdiffusion 52 -29 52 -29 0 cellNo=190
rlabel pdiffusion 73 -29 73 -29 0 feedthrough
rlabel pdiffusion 80 -29 80 -29 0 cellNo=105
rlabel pdiffusion 94 -29 94 -29 0 cellNo=296
rlabel pdiffusion 101 -29 101 -29 0 cellNo=10
rlabel pdiffusion 108 -29 108 -29 0 cellNo=286
rlabel pdiffusion 115 -29 115 -29 0 cellNo=193
rlabel pdiffusion 122 -29 122 -29 0 cellNo=52
rlabel pdiffusion 129 -29 129 -29 0 feedthrough
rlabel pdiffusion 143 -29 143 -29 0 feedthrough
rlabel pdiffusion 150 -29 150 -29 0 feedthrough
rlabel pdiffusion 164 -29 164 -29 0 feedthrough
rlabel pdiffusion 171 -29 171 -29 0 cellNo=297
rlabel pdiffusion 178 -29 178 -29 0 feedthrough
rlabel pdiffusion 185 -29 185 -29 0 cellNo=109
rlabel pdiffusion 192 -29 192 -29 0 cellNo=194
rlabel pdiffusion 199 -29 199 -29 0 cellNo=243
rlabel pdiffusion 3 -60 3 -60 0 cellNo=198
rlabel pdiffusion 10 -60 10 -60 0 cellNo=42
rlabel pdiffusion 17 -60 17 -60 0 cellNo=254
rlabel pdiffusion 24 -60 24 -60 0 cellNo=64
rlabel pdiffusion 31 -60 31 -60 0 cellNo=294
rlabel pdiffusion 38 -60 38 -60 0 cellNo=214
rlabel pdiffusion 45 -60 45 -60 0 cellNo=244
rlabel pdiffusion 52 -60 52 -60 0 feedthrough
rlabel pdiffusion 59 -60 59 -60 0 feedthrough
rlabel pdiffusion 66 -60 66 -60 0 feedthrough
rlabel pdiffusion 73 -60 73 -60 0 feedthrough
rlabel pdiffusion 80 -60 80 -60 0 cellNo=207
rlabel pdiffusion 87 -60 87 -60 0 cellNo=97
rlabel pdiffusion 94 -60 94 -60 0 cellNo=348
rlabel pdiffusion 101 -60 101 -60 0 feedthrough
rlabel pdiffusion 108 -60 108 -60 0 cellNo=236
rlabel pdiffusion 115 -60 115 -60 0 cellNo=51
rlabel pdiffusion 122 -60 122 -60 0 cellNo=164
rlabel pdiffusion 129 -60 129 -60 0 cellNo=38
rlabel pdiffusion 136 -60 136 -60 0 cellNo=268
rlabel pdiffusion 143 -60 143 -60 0 cellNo=128
rlabel pdiffusion 150 -60 150 -60 0 cellNo=120
rlabel pdiffusion 157 -60 157 -60 0 feedthrough
rlabel pdiffusion 164 -60 164 -60 0 feedthrough
rlabel pdiffusion 171 -60 171 -60 0 feedthrough
rlabel pdiffusion 178 -60 178 -60 0 feedthrough
rlabel pdiffusion 185 -60 185 -60 0 feedthrough
rlabel pdiffusion 192 -60 192 -60 0 cellNo=32
rlabel pdiffusion 199 -60 199 -60 0 feedthrough
rlabel pdiffusion 206 -60 206 -60 0 feedthrough
rlabel pdiffusion 213 -60 213 -60 0 feedthrough
rlabel pdiffusion 220 -60 220 -60 0 feedthrough
rlabel pdiffusion 227 -60 227 -60 0 feedthrough
rlabel pdiffusion 234 -60 234 -60 0 feedthrough
rlabel pdiffusion 241 -60 241 -60 0 cellNo=201
rlabel pdiffusion 248 -60 248 -60 0 feedthrough
rlabel pdiffusion 255 -60 255 -60 0 feedthrough
rlabel pdiffusion 10 -93 10 -93 0 cellNo=310
rlabel pdiffusion 17 -93 17 -93 0 cellNo=251
rlabel pdiffusion 24 -93 24 -93 0 cellNo=170
rlabel pdiffusion 31 -93 31 -93 0 feedthrough
rlabel pdiffusion 38 -93 38 -93 0 cellNo=95
rlabel pdiffusion 45 -93 45 -93 0 feedthrough
rlabel pdiffusion 52 -93 52 -93 0 feedthrough
rlabel pdiffusion 59 -93 59 -93 0 feedthrough
rlabel pdiffusion 66 -93 66 -93 0 feedthrough
rlabel pdiffusion 73 -93 73 -93 0 feedthrough
rlabel pdiffusion 80 -93 80 -93 0 cellNo=53
rlabel pdiffusion 87 -93 87 -93 0 feedthrough
rlabel pdiffusion 94 -93 94 -93 0 cellNo=324
rlabel pdiffusion 101 -93 101 -93 0 cellNo=118
rlabel pdiffusion 108 -93 108 -93 0 cellNo=285
rlabel pdiffusion 115 -93 115 -93 0 cellNo=28
rlabel pdiffusion 122 -93 122 -93 0 feedthrough
rlabel pdiffusion 129 -93 129 -93 0 cellNo=151
rlabel pdiffusion 136 -93 136 -93 0 cellNo=233
rlabel pdiffusion 143 -93 143 -93 0 cellNo=210
rlabel pdiffusion 150 -93 150 -93 0 cellNo=130
rlabel pdiffusion 157 -93 157 -93 0 cellNo=80
rlabel pdiffusion 164 -93 164 -93 0 cellNo=326
rlabel pdiffusion 171 -93 171 -93 0 cellNo=211
rlabel pdiffusion 178 -93 178 -93 0 feedthrough
rlabel pdiffusion 185 -93 185 -93 0 cellNo=311
rlabel pdiffusion 192 -93 192 -93 0 feedthrough
rlabel pdiffusion 199 -93 199 -93 0 cellNo=6
rlabel pdiffusion 206 -93 206 -93 0 feedthrough
rlabel pdiffusion 213 -93 213 -93 0 feedthrough
rlabel pdiffusion 220 -93 220 -93 0 feedthrough
rlabel pdiffusion 227 -93 227 -93 0 feedthrough
rlabel pdiffusion 234 -93 234 -93 0 feedthrough
rlabel pdiffusion 241 -93 241 -93 0 feedthrough
rlabel pdiffusion 248 -93 248 -93 0 feedthrough
rlabel pdiffusion 255 -93 255 -93 0 feedthrough
rlabel pdiffusion 262 -93 262 -93 0 feedthrough
rlabel pdiffusion 269 -93 269 -93 0 feedthrough
rlabel pdiffusion 276 -93 276 -93 0 feedthrough
rlabel pdiffusion 283 -93 283 -93 0 feedthrough
rlabel pdiffusion 290 -93 290 -93 0 feedthrough
rlabel pdiffusion 297 -93 297 -93 0 feedthrough
rlabel pdiffusion 304 -93 304 -93 0 cellNo=24
rlabel pdiffusion 332 -93 332 -93 0 feedthrough
rlabel pdiffusion 3 -148 3 -148 0 cellNo=45
rlabel pdiffusion 10 -148 10 -148 0 cellNo=100
rlabel pdiffusion 17 -148 17 -148 0 cellNo=132
rlabel pdiffusion 24 -148 24 -148 0 cellNo=49
rlabel pdiffusion 31 -148 31 -148 0 cellNo=115
rlabel pdiffusion 38 -148 38 -148 0 cellNo=7
rlabel pdiffusion 45 -148 45 -148 0 feedthrough
rlabel pdiffusion 52 -148 52 -148 0 feedthrough
rlabel pdiffusion 59 -148 59 -148 0 cellNo=5
rlabel pdiffusion 66 -148 66 -148 0 feedthrough
rlabel pdiffusion 73 -148 73 -148 0 feedthrough
rlabel pdiffusion 80 -148 80 -148 0 cellNo=259
rlabel pdiffusion 87 -148 87 -148 0 cellNo=30
rlabel pdiffusion 94 -148 94 -148 0 feedthrough
rlabel pdiffusion 101 -148 101 -148 0 feedthrough
rlabel pdiffusion 108 -148 108 -148 0 feedthrough
rlabel pdiffusion 115 -148 115 -148 0 cellNo=357
rlabel pdiffusion 122 -148 122 -148 0 cellNo=265
rlabel pdiffusion 129 -148 129 -148 0 cellNo=234
rlabel pdiffusion 136 -148 136 -148 0 cellNo=122
rlabel pdiffusion 143 -148 143 -148 0 feedthrough
rlabel pdiffusion 150 -148 150 -148 0 cellNo=133
rlabel pdiffusion 157 -148 157 -148 0 feedthrough
rlabel pdiffusion 164 -148 164 -148 0 cellNo=111
rlabel pdiffusion 171 -148 171 -148 0 feedthrough
rlabel pdiffusion 178 -148 178 -148 0 feedthrough
rlabel pdiffusion 185 -148 185 -148 0 feedthrough
rlabel pdiffusion 192 -148 192 -148 0 cellNo=119
rlabel pdiffusion 199 -148 199 -148 0 cellNo=27
rlabel pdiffusion 206 -148 206 -148 0 cellNo=125
rlabel pdiffusion 213 -148 213 -148 0 feedthrough
rlabel pdiffusion 220 -148 220 -148 0 feedthrough
rlabel pdiffusion 227 -148 227 -148 0 feedthrough
rlabel pdiffusion 234 -148 234 -148 0 feedthrough
rlabel pdiffusion 241 -148 241 -148 0 feedthrough
rlabel pdiffusion 248 -148 248 -148 0 feedthrough
rlabel pdiffusion 255 -148 255 -148 0 feedthrough
rlabel pdiffusion 262 -148 262 -148 0 feedthrough
rlabel pdiffusion 269 -148 269 -148 0 cellNo=67
rlabel pdiffusion 276 -148 276 -148 0 feedthrough
rlabel pdiffusion 283 -148 283 -148 0 feedthrough
rlabel pdiffusion 290 -148 290 -148 0 feedthrough
rlabel pdiffusion 297 -148 297 -148 0 feedthrough
rlabel pdiffusion 304 -148 304 -148 0 feedthrough
rlabel pdiffusion 311 -148 311 -148 0 feedthrough
rlabel pdiffusion 318 -148 318 -148 0 feedthrough
rlabel pdiffusion 325 -148 325 -148 0 feedthrough
rlabel pdiffusion 332 -148 332 -148 0 feedthrough
rlabel pdiffusion 339 -148 339 -148 0 feedthrough
rlabel pdiffusion 346 -148 346 -148 0 feedthrough
rlabel pdiffusion 353 -148 353 -148 0 feedthrough
rlabel pdiffusion 360 -148 360 -148 0 feedthrough
rlabel pdiffusion 367 -148 367 -148 0 feedthrough
rlabel pdiffusion 374 -148 374 -148 0 feedthrough
rlabel pdiffusion 3 -199 3 -199 0 cellNo=136
rlabel pdiffusion 10 -199 10 -199 0 feedthrough
rlabel pdiffusion 17 -199 17 -199 0 feedthrough
rlabel pdiffusion 24 -199 24 -199 0 cellNo=186
rlabel pdiffusion 31 -199 31 -199 0 feedthrough
rlabel pdiffusion 38 -199 38 -199 0 feedthrough
rlabel pdiffusion 45 -199 45 -199 0 cellNo=139
rlabel pdiffusion 52 -199 52 -199 0 feedthrough
rlabel pdiffusion 59 -199 59 -199 0 cellNo=43
rlabel pdiffusion 66 -199 66 -199 0 feedthrough
rlabel pdiffusion 73 -199 73 -199 0 cellNo=41
rlabel pdiffusion 80 -199 80 -199 0 cellNo=48
rlabel pdiffusion 87 -199 87 -199 0 feedthrough
rlabel pdiffusion 94 -199 94 -199 0 cellNo=289
rlabel pdiffusion 101 -199 101 -199 0 cellNo=298
rlabel pdiffusion 108 -199 108 -199 0 feedthrough
rlabel pdiffusion 115 -199 115 -199 0 feedthrough
rlabel pdiffusion 122 -199 122 -199 0 feedthrough
rlabel pdiffusion 129 -199 129 -199 0 cellNo=112
rlabel pdiffusion 136 -199 136 -199 0 cellNo=174
rlabel pdiffusion 143 -199 143 -199 0 feedthrough
rlabel pdiffusion 150 -199 150 -199 0 cellNo=197
rlabel pdiffusion 157 -199 157 -199 0 feedthrough
rlabel pdiffusion 164 -199 164 -199 0 cellNo=267
rlabel pdiffusion 171 -199 171 -199 0 cellNo=277
rlabel pdiffusion 178 -199 178 -199 0 feedthrough
rlabel pdiffusion 185 -199 185 -199 0 cellNo=4
rlabel pdiffusion 192 -199 192 -199 0 feedthrough
rlabel pdiffusion 199 -199 199 -199 0 cellNo=266
rlabel pdiffusion 206 -199 206 -199 0 cellNo=75
rlabel pdiffusion 213 -199 213 -199 0 feedthrough
rlabel pdiffusion 220 -199 220 -199 0 cellNo=71
rlabel pdiffusion 227 -199 227 -199 0 feedthrough
rlabel pdiffusion 234 -199 234 -199 0 feedthrough
rlabel pdiffusion 241 -199 241 -199 0 feedthrough
rlabel pdiffusion 248 -199 248 -199 0 feedthrough
rlabel pdiffusion 255 -199 255 -199 0 feedthrough
rlabel pdiffusion 262 -199 262 -199 0 feedthrough
rlabel pdiffusion 269 -199 269 -199 0 feedthrough
rlabel pdiffusion 276 -199 276 -199 0 feedthrough
rlabel pdiffusion 283 -199 283 -199 0 feedthrough
rlabel pdiffusion 290 -199 290 -199 0 feedthrough
rlabel pdiffusion 297 -199 297 -199 0 feedthrough
rlabel pdiffusion 304 -199 304 -199 0 feedthrough
rlabel pdiffusion 311 -199 311 -199 0 feedthrough
rlabel pdiffusion 318 -199 318 -199 0 cellNo=202
rlabel pdiffusion 325 -199 325 -199 0 feedthrough
rlabel pdiffusion 332 -199 332 -199 0 feedthrough
rlabel pdiffusion 339 -199 339 -199 0 feedthrough
rlabel pdiffusion 346 -199 346 -199 0 feedthrough
rlabel pdiffusion 353 -199 353 -199 0 feedthrough
rlabel pdiffusion 360 -199 360 -199 0 feedthrough
rlabel pdiffusion 367 -199 367 -199 0 feedthrough
rlabel pdiffusion 374 -199 374 -199 0 feedthrough
rlabel pdiffusion 381 -199 381 -199 0 feedthrough
rlabel pdiffusion 388 -199 388 -199 0 feedthrough
rlabel pdiffusion 395 -199 395 -199 0 feedthrough
rlabel pdiffusion 402 -199 402 -199 0 feedthrough
rlabel pdiffusion 409 -199 409 -199 0 cellNo=74
rlabel pdiffusion 416 -199 416 -199 0 feedthrough
rlabel pdiffusion 3 -258 3 -258 0 cellNo=81
rlabel pdiffusion 10 -258 10 -258 0 cellNo=313
rlabel pdiffusion 17 -258 17 -258 0 feedthrough
rlabel pdiffusion 24 -258 24 -258 0 feedthrough
rlabel pdiffusion 31 -258 31 -258 0 cellNo=141
rlabel pdiffusion 38 -258 38 -258 0 feedthrough
rlabel pdiffusion 45 -258 45 -258 0 feedthrough
rlabel pdiffusion 52 -258 52 -258 0 cellNo=110
rlabel pdiffusion 59 -258 59 -258 0 feedthrough
rlabel pdiffusion 66 -258 66 -258 0 feedthrough
rlabel pdiffusion 73 -258 73 -258 0 cellNo=330
rlabel pdiffusion 80 -258 80 -258 0 cellNo=281
rlabel pdiffusion 87 -258 87 -258 0 feedthrough
rlabel pdiffusion 94 -258 94 -258 0 cellNo=222
rlabel pdiffusion 101 -258 101 -258 0 cellNo=143
rlabel pdiffusion 108 -258 108 -258 0 cellNo=188
rlabel pdiffusion 115 -258 115 -258 0 cellNo=93
rlabel pdiffusion 122 -258 122 -258 0 cellNo=22
rlabel pdiffusion 129 -258 129 -258 0 feedthrough
rlabel pdiffusion 136 -258 136 -258 0 cellNo=149
rlabel pdiffusion 143 -258 143 -258 0 feedthrough
rlabel pdiffusion 150 -258 150 -258 0 feedthrough
rlabel pdiffusion 157 -258 157 -258 0 feedthrough
rlabel pdiffusion 164 -258 164 -258 0 feedthrough
rlabel pdiffusion 171 -258 171 -258 0 feedthrough
rlabel pdiffusion 178 -258 178 -258 0 cellNo=68
rlabel pdiffusion 185 -258 185 -258 0 cellNo=88
rlabel pdiffusion 192 -258 192 -258 0 feedthrough
rlabel pdiffusion 199 -258 199 -258 0 cellNo=353
rlabel pdiffusion 206 -258 206 -258 0 feedthrough
rlabel pdiffusion 213 -258 213 -258 0 feedthrough
rlabel pdiffusion 220 -258 220 -258 0 cellNo=246
rlabel pdiffusion 227 -258 227 -258 0 feedthrough
rlabel pdiffusion 234 -258 234 -258 0 feedthrough
rlabel pdiffusion 241 -258 241 -258 0 cellNo=57
rlabel pdiffusion 248 -258 248 -258 0 feedthrough
rlabel pdiffusion 255 -258 255 -258 0 cellNo=155
rlabel pdiffusion 262 -258 262 -258 0 feedthrough
rlabel pdiffusion 269 -258 269 -258 0 feedthrough
rlabel pdiffusion 276 -258 276 -258 0 feedthrough
rlabel pdiffusion 283 -258 283 -258 0 cellNo=290
rlabel pdiffusion 290 -258 290 -258 0 feedthrough
rlabel pdiffusion 297 -258 297 -258 0 feedthrough
rlabel pdiffusion 304 -258 304 -258 0 feedthrough
rlabel pdiffusion 311 -258 311 -258 0 feedthrough
rlabel pdiffusion 318 -258 318 -258 0 feedthrough
rlabel pdiffusion 325 -258 325 -258 0 feedthrough
rlabel pdiffusion 332 -258 332 -258 0 feedthrough
rlabel pdiffusion 339 -258 339 -258 0 feedthrough
rlabel pdiffusion 346 -258 346 -258 0 feedthrough
rlabel pdiffusion 353 -258 353 -258 0 feedthrough
rlabel pdiffusion 360 -258 360 -258 0 feedthrough
rlabel pdiffusion 367 -258 367 -258 0 feedthrough
rlabel pdiffusion 374 -258 374 -258 0 feedthrough
rlabel pdiffusion 381 -258 381 -258 0 feedthrough
rlabel pdiffusion 388 -258 388 -258 0 feedthrough
rlabel pdiffusion 395 -258 395 -258 0 feedthrough
rlabel pdiffusion 402 -258 402 -258 0 feedthrough
rlabel pdiffusion 409 -258 409 -258 0 feedthrough
rlabel pdiffusion 416 -258 416 -258 0 feedthrough
rlabel pdiffusion 3 -307 3 -307 0 cellNo=152
rlabel pdiffusion 10 -307 10 -307 0 cellNo=276
rlabel pdiffusion 17 -307 17 -307 0 feedthrough
rlabel pdiffusion 24 -307 24 -307 0 feedthrough
rlabel pdiffusion 31 -307 31 -307 0 feedthrough
rlabel pdiffusion 38 -307 38 -307 0 feedthrough
rlabel pdiffusion 45 -307 45 -307 0 feedthrough
rlabel pdiffusion 52 -307 52 -307 0 feedthrough
rlabel pdiffusion 59 -307 59 -307 0 cellNo=44
rlabel pdiffusion 66 -307 66 -307 0 feedthrough
rlabel pdiffusion 73 -307 73 -307 0 cellNo=31
rlabel pdiffusion 80 -307 80 -307 0 feedthrough
rlabel pdiffusion 87 -307 87 -307 0 feedthrough
rlabel pdiffusion 94 -307 94 -307 0 cellNo=34
rlabel pdiffusion 101 -307 101 -307 0 cellNo=239
rlabel pdiffusion 108 -307 108 -307 0 cellNo=127
rlabel pdiffusion 115 -307 115 -307 0 cellNo=148
rlabel pdiffusion 122 -307 122 -307 0 cellNo=272
rlabel pdiffusion 129 -307 129 -307 0 feedthrough
rlabel pdiffusion 136 -307 136 -307 0 feedthrough
rlabel pdiffusion 143 -307 143 -307 0 feedthrough
rlabel pdiffusion 150 -307 150 -307 0 feedthrough
rlabel pdiffusion 157 -307 157 -307 0 feedthrough
rlabel pdiffusion 164 -307 164 -307 0 cellNo=253
rlabel pdiffusion 171 -307 171 -307 0 cellNo=332
rlabel pdiffusion 178 -307 178 -307 0 feedthrough
rlabel pdiffusion 185 -307 185 -307 0 feedthrough
rlabel pdiffusion 192 -307 192 -307 0 feedthrough
rlabel pdiffusion 199 -307 199 -307 0 cellNo=232
rlabel pdiffusion 206 -307 206 -307 0 cellNo=184
rlabel pdiffusion 213 -307 213 -307 0 cellNo=218
rlabel pdiffusion 220 -307 220 -307 0 feedthrough
rlabel pdiffusion 227 -307 227 -307 0 feedthrough
rlabel pdiffusion 234 -307 234 -307 0 feedthrough
rlabel pdiffusion 241 -307 241 -307 0 cellNo=94
rlabel pdiffusion 248 -307 248 -307 0 cellNo=78
rlabel pdiffusion 255 -307 255 -307 0 feedthrough
rlabel pdiffusion 262 -307 262 -307 0 cellNo=135
rlabel pdiffusion 269 -307 269 -307 0 feedthrough
rlabel pdiffusion 276 -307 276 -307 0 feedthrough
rlabel pdiffusion 283 -307 283 -307 0 feedthrough
rlabel pdiffusion 290 -307 290 -307 0 feedthrough
rlabel pdiffusion 297 -307 297 -307 0 feedthrough
rlabel pdiffusion 304 -307 304 -307 0 feedthrough
rlabel pdiffusion 311 -307 311 -307 0 feedthrough
rlabel pdiffusion 318 -307 318 -307 0 feedthrough
rlabel pdiffusion 325 -307 325 -307 0 feedthrough
rlabel pdiffusion 332 -307 332 -307 0 feedthrough
rlabel pdiffusion 339 -307 339 -307 0 feedthrough
rlabel pdiffusion 346 -307 346 -307 0 feedthrough
rlabel pdiffusion 353 -307 353 -307 0 feedthrough
rlabel pdiffusion 360 -307 360 -307 0 feedthrough
rlabel pdiffusion 367 -307 367 -307 0 feedthrough
rlabel pdiffusion 374 -307 374 -307 0 feedthrough
rlabel pdiffusion 381 -307 381 -307 0 feedthrough
rlabel pdiffusion 388 -307 388 -307 0 feedthrough
rlabel pdiffusion 395 -307 395 -307 0 feedthrough
rlabel pdiffusion 402 -307 402 -307 0 feedthrough
rlabel pdiffusion 409 -307 409 -307 0 feedthrough
rlabel pdiffusion 416 -307 416 -307 0 feedthrough
rlabel pdiffusion 423 -307 423 -307 0 cellNo=200
rlabel pdiffusion 430 -307 430 -307 0 cellNo=66
rlabel pdiffusion 437 -307 437 -307 0 feedthrough
rlabel pdiffusion 3 -368 3 -368 0 feedthrough
rlabel pdiffusion 10 -368 10 -368 0 cellNo=335
rlabel pdiffusion 17 -368 17 -368 0 feedthrough
rlabel pdiffusion 24 -368 24 -368 0 cellNo=107
rlabel pdiffusion 31 -368 31 -368 0 cellNo=284
rlabel pdiffusion 38 -368 38 -368 0 cellNo=47
rlabel pdiffusion 45 -368 45 -368 0 cellNo=287
rlabel pdiffusion 52 -368 52 -368 0 cellNo=142
rlabel pdiffusion 59 -368 59 -368 0 feedthrough
rlabel pdiffusion 66 -368 66 -368 0 cellNo=231
rlabel pdiffusion 73 -368 73 -368 0 cellNo=13
rlabel pdiffusion 80 -368 80 -368 0 cellNo=145
rlabel pdiffusion 87 -368 87 -368 0 cellNo=204
rlabel pdiffusion 94 -368 94 -368 0 feedthrough
rlabel pdiffusion 101 -368 101 -368 0 feedthrough
rlabel pdiffusion 108 -368 108 -368 0 cellNo=98
rlabel pdiffusion 115 -368 115 -368 0 cellNo=15
rlabel pdiffusion 122 -368 122 -368 0 feedthrough
rlabel pdiffusion 129 -368 129 -368 0 feedthrough
rlabel pdiffusion 136 -368 136 -368 0 feedthrough
rlabel pdiffusion 143 -368 143 -368 0 feedthrough
rlabel pdiffusion 150 -368 150 -368 0 feedthrough
rlabel pdiffusion 157 -368 157 -368 0 cellNo=166
rlabel pdiffusion 164 -368 164 -368 0 feedthrough
rlabel pdiffusion 171 -368 171 -368 0 cellNo=163
rlabel pdiffusion 178 -368 178 -368 0 feedthrough
rlabel pdiffusion 185 -368 185 -368 0 cellNo=161
rlabel pdiffusion 192 -368 192 -368 0 feedthrough
rlabel pdiffusion 199 -368 199 -368 0 feedthrough
rlabel pdiffusion 206 -368 206 -368 0 feedthrough
rlabel pdiffusion 213 -368 213 -368 0 feedthrough
rlabel pdiffusion 220 -368 220 -368 0 cellNo=315
rlabel pdiffusion 227 -368 227 -368 0 feedthrough
rlabel pdiffusion 234 -368 234 -368 0 cellNo=227
rlabel pdiffusion 241 -368 241 -368 0 feedthrough
rlabel pdiffusion 248 -368 248 -368 0 feedthrough
rlabel pdiffusion 255 -368 255 -368 0 cellNo=39
rlabel pdiffusion 262 -368 262 -368 0 feedthrough
rlabel pdiffusion 269 -368 269 -368 0 cellNo=150
rlabel pdiffusion 276 -368 276 -368 0 feedthrough
rlabel pdiffusion 283 -368 283 -368 0 feedthrough
rlabel pdiffusion 290 -368 290 -368 0 feedthrough
rlabel pdiffusion 297 -368 297 -368 0 feedthrough
rlabel pdiffusion 304 -368 304 -368 0 feedthrough
rlabel pdiffusion 311 -368 311 -368 0 feedthrough
rlabel pdiffusion 318 -368 318 -368 0 feedthrough
rlabel pdiffusion 325 -368 325 -368 0 feedthrough
rlabel pdiffusion 332 -368 332 -368 0 feedthrough
rlabel pdiffusion 339 -368 339 -368 0 feedthrough
rlabel pdiffusion 346 -368 346 -368 0 feedthrough
rlabel pdiffusion 353 -368 353 -368 0 feedthrough
rlabel pdiffusion 360 -368 360 -368 0 feedthrough
rlabel pdiffusion 367 -368 367 -368 0 feedthrough
rlabel pdiffusion 374 -368 374 -368 0 feedthrough
rlabel pdiffusion 381 -368 381 -368 0 feedthrough
rlabel pdiffusion 388 -368 388 -368 0 feedthrough
rlabel pdiffusion 395 -368 395 -368 0 feedthrough
rlabel pdiffusion 402 -368 402 -368 0 feedthrough
rlabel pdiffusion 409 -368 409 -368 0 feedthrough
rlabel pdiffusion 416 -368 416 -368 0 feedthrough
rlabel pdiffusion 423 -368 423 -368 0 feedthrough
rlabel pdiffusion 430 -368 430 -368 0 feedthrough
rlabel pdiffusion 437 -368 437 -368 0 feedthrough
rlabel pdiffusion 10 -417 10 -417 0 feedthrough
rlabel pdiffusion 17 -417 17 -417 0 feedthrough
rlabel pdiffusion 24 -417 24 -417 0 cellNo=89
rlabel pdiffusion 31 -417 31 -417 0 feedthrough
rlabel pdiffusion 38 -417 38 -417 0 feedthrough
rlabel pdiffusion 45 -417 45 -417 0 cellNo=162
rlabel pdiffusion 52 -417 52 -417 0 cellNo=316
rlabel pdiffusion 59 -417 59 -417 0 cellNo=126
rlabel pdiffusion 66 -417 66 -417 0 feedthrough
rlabel pdiffusion 73 -417 73 -417 0 feedthrough
rlabel pdiffusion 80 -417 80 -417 0 feedthrough
rlabel pdiffusion 87 -417 87 -417 0 feedthrough
rlabel pdiffusion 94 -417 94 -417 0 feedthrough
rlabel pdiffusion 101 -417 101 -417 0 cellNo=314
rlabel pdiffusion 108 -417 108 -417 0 cellNo=62
rlabel pdiffusion 115 -417 115 -417 0 cellNo=270
rlabel pdiffusion 122 -417 122 -417 0 feedthrough
rlabel pdiffusion 129 -417 129 -417 0 cellNo=255
rlabel pdiffusion 136 -417 136 -417 0 feedthrough
rlabel pdiffusion 143 -417 143 -417 0 feedthrough
rlabel pdiffusion 150 -417 150 -417 0 feedthrough
rlabel pdiffusion 157 -417 157 -417 0 feedthrough
rlabel pdiffusion 164 -417 164 -417 0 cellNo=359
rlabel pdiffusion 171 -417 171 -417 0 feedthrough
rlabel pdiffusion 178 -417 178 -417 0 feedthrough
rlabel pdiffusion 185 -417 185 -417 0 feedthrough
rlabel pdiffusion 192 -417 192 -417 0 feedthrough
rlabel pdiffusion 199 -417 199 -417 0 cellNo=358
rlabel pdiffusion 206 -417 206 -417 0 feedthrough
rlabel pdiffusion 213 -417 213 -417 0 feedthrough
rlabel pdiffusion 220 -417 220 -417 0 feedthrough
rlabel pdiffusion 227 -417 227 -417 0 cellNo=180
rlabel pdiffusion 234 -417 234 -417 0 feedthrough
rlabel pdiffusion 241 -417 241 -417 0 cellNo=168
rlabel pdiffusion 248 -417 248 -417 0 cellNo=131
rlabel pdiffusion 255 -417 255 -417 0 feedthrough
rlabel pdiffusion 262 -417 262 -417 0 cellNo=343
rlabel pdiffusion 269 -417 269 -417 0 cellNo=229
rlabel pdiffusion 276 -417 276 -417 0 feedthrough
rlabel pdiffusion 283 -417 283 -417 0 feedthrough
rlabel pdiffusion 290 -417 290 -417 0 feedthrough
rlabel pdiffusion 297 -417 297 -417 0 feedthrough
rlabel pdiffusion 304 -417 304 -417 0 feedthrough
rlabel pdiffusion 311 -417 311 -417 0 feedthrough
rlabel pdiffusion 318 -417 318 -417 0 feedthrough
rlabel pdiffusion 325 -417 325 -417 0 cellNo=172
rlabel pdiffusion 332 -417 332 -417 0 cellNo=238
rlabel pdiffusion 339 -417 339 -417 0 feedthrough
rlabel pdiffusion 346 -417 346 -417 0 feedthrough
rlabel pdiffusion 353 -417 353 -417 0 feedthrough
rlabel pdiffusion 360 -417 360 -417 0 feedthrough
rlabel pdiffusion 367 -417 367 -417 0 feedthrough
rlabel pdiffusion 374 -417 374 -417 0 feedthrough
rlabel pdiffusion 381 -417 381 -417 0 feedthrough
rlabel pdiffusion 388 -417 388 -417 0 feedthrough
rlabel pdiffusion 395 -417 395 -417 0 feedthrough
rlabel pdiffusion 402 -417 402 -417 0 feedthrough
rlabel pdiffusion 409 -417 409 -417 0 feedthrough
rlabel pdiffusion 416 -417 416 -417 0 feedthrough
rlabel pdiffusion 423 -417 423 -417 0 feedthrough
rlabel pdiffusion 430 -417 430 -417 0 cellNo=217
rlabel pdiffusion 437 -417 437 -417 0 feedthrough
rlabel pdiffusion 444 -417 444 -417 0 cellNo=300
rlabel pdiffusion 17 -472 17 -472 0 feedthrough
rlabel pdiffusion 24 -472 24 -472 0 cellNo=256
rlabel pdiffusion 31 -472 31 -472 0 cellNo=3
rlabel pdiffusion 38 -472 38 -472 0 feedthrough
rlabel pdiffusion 52 -472 52 -472 0 feedthrough
rlabel pdiffusion 59 -472 59 -472 0 feedthrough
rlabel pdiffusion 66 -472 66 -472 0 feedthrough
rlabel pdiffusion 73 -472 73 -472 0 cellNo=146
rlabel pdiffusion 80 -472 80 -472 0 feedthrough
rlabel pdiffusion 87 -472 87 -472 0 feedthrough
rlabel pdiffusion 94 -472 94 -472 0 feedthrough
rlabel pdiffusion 101 -472 101 -472 0 feedthrough
rlabel pdiffusion 108 -472 108 -472 0 cellNo=33
rlabel pdiffusion 115 -472 115 -472 0 feedthrough
rlabel pdiffusion 122 -472 122 -472 0 feedthrough
rlabel pdiffusion 129 -472 129 -472 0 cellNo=312
rlabel pdiffusion 136 -472 136 -472 0 feedthrough
rlabel pdiffusion 143 -472 143 -472 0 feedthrough
rlabel pdiffusion 150 -472 150 -472 0 feedthrough
rlabel pdiffusion 157 -472 157 -472 0 feedthrough
rlabel pdiffusion 164 -472 164 -472 0 feedthrough
rlabel pdiffusion 171 -472 171 -472 0 feedthrough
rlabel pdiffusion 178 -472 178 -472 0 cellNo=159
rlabel pdiffusion 185 -472 185 -472 0 feedthrough
rlabel pdiffusion 192 -472 192 -472 0 cellNo=16
rlabel pdiffusion 199 -472 199 -472 0 cellNo=245
rlabel pdiffusion 206 -472 206 -472 0 feedthrough
rlabel pdiffusion 213 -472 213 -472 0 cellNo=302
rlabel pdiffusion 220 -472 220 -472 0 cellNo=90
rlabel pdiffusion 227 -472 227 -472 0 cellNo=76
rlabel pdiffusion 234 -472 234 -472 0 cellNo=2
rlabel pdiffusion 241 -472 241 -472 0 cellNo=252
rlabel pdiffusion 248 -472 248 -472 0 cellNo=54
rlabel pdiffusion 255 -472 255 -472 0 cellNo=288
rlabel pdiffusion 262 -472 262 -472 0 cellNo=55
rlabel pdiffusion 269 -472 269 -472 0 feedthrough
rlabel pdiffusion 276 -472 276 -472 0 feedthrough
rlabel pdiffusion 283 -472 283 -472 0 cellNo=282
rlabel pdiffusion 290 -472 290 -472 0 feedthrough
rlabel pdiffusion 297 -472 297 -472 0 feedthrough
rlabel pdiffusion 304 -472 304 -472 0 feedthrough
rlabel pdiffusion 311 -472 311 -472 0 feedthrough
rlabel pdiffusion 318 -472 318 -472 0 feedthrough
rlabel pdiffusion 325 -472 325 -472 0 feedthrough
rlabel pdiffusion 332 -472 332 -472 0 feedthrough
rlabel pdiffusion 339 -472 339 -472 0 feedthrough
rlabel pdiffusion 346 -472 346 -472 0 feedthrough
rlabel pdiffusion 353 -472 353 -472 0 feedthrough
rlabel pdiffusion 360 -472 360 -472 0 feedthrough
rlabel pdiffusion 367 -472 367 -472 0 feedthrough
rlabel pdiffusion 374 -472 374 -472 0 feedthrough
rlabel pdiffusion 381 -472 381 -472 0 feedthrough
rlabel pdiffusion 388 -472 388 -472 0 feedthrough
rlabel pdiffusion 395 -472 395 -472 0 feedthrough
rlabel pdiffusion 416 -472 416 -472 0 feedthrough
rlabel pdiffusion 423 -472 423 -472 0 feedthrough
rlabel pdiffusion 430 -472 430 -472 0 cellNo=341
rlabel pdiffusion 437 -472 437 -472 0 feedthrough
rlabel pdiffusion 444 -472 444 -472 0 cellNo=19
rlabel pdiffusion 451 -472 451 -472 0 feedthrough
rlabel pdiffusion 458 -472 458 -472 0 feedthrough
rlabel pdiffusion 465 -472 465 -472 0 feedthrough
rlabel pdiffusion 10 -513 10 -513 0 feedthrough
rlabel pdiffusion 17 -513 17 -513 0 feedthrough
rlabel pdiffusion 24 -513 24 -513 0 cellNo=240
rlabel pdiffusion 31 -513 31 -513 0 cellNo=319
rlabel pdiffusion 38 -513 38 -513 0 cellNo=9
rlabel pdiffusion 45 -513 45 -513 0 feedthrough
rlabel pdiffusion 52 -513 52 -513 0 feedthrough
rlabel pdiffusion 59 -513 59 -513 0 feedthrough
rlabel pdiffusion 66 -513 66 -513 0 feedthrough
rlabel pdiffusion 73 -513 73 -513 0 cellNo=87
rlabel pdiffusion 80 -513 80 -513 0 cellNo=121
rlabel pdiffusion 87 -513 87 -513 0 feedthrough
rlabel pdiffusion 94 -513 94 -513 0 feedthrough
rlabel pdiffusion 101 -513 101 -513 0 cellNo=56
rlabel pdiffusion 108 -513 108 -513 0 feedthrough
rlabel pdiffusion 115 -513 115 -513 0 feedthrough
rlabel pdiffusion 122 -513 122 -513 0 cellNo=250
rlabel pdiffusion 129 -513 129 -513 0 feedthrough
rlabel pdiffusion 136 -513 136 -513 0 cellNo=176
rlabel pdiffusion 143 -513 143 -513 0 feedthrough
rlabel pdiffusion 150 -513 150 -513 0 feedthrough
rlabel pdiffusion 157 -513 157 -513 0 feedthrough
rlabel pdiffusion 164 -513 164 -513 0 feedthrough
rlabel pdiffusion 171 -513 171 -513 0 cellNo=235
rlabel pdiffusion 178 -513 178 -513 0 feedthrough
rlabel pdiffusion 185 -513 185 -513 0 feedthrough
rlabel pdiffusion 192 -513 192 -513 0 feedthrough
rlabel pdiffusion 199 -513 199 -513 0 feedthrough
rlabel pdiffusion 206 -513 206 -513 0 cellNo=40
rlabel pdiffusion 213 -513 213 -513 0 cellNo=333
rlabel pdiffusion 220 -513 220 -513 0 feedthrough
rlabel pdiffusion 227 -513 227 -513 0 feedthrough
rlabel pdiffusion 234 -513 234 -513 0 feedthrough
rlabel pdiffusion 241 -513 241 -513 0 cellNo=219
rlabel pdiffusion 248 -513 248 -513 0 feedthrough
rlabel pdiffusion 255 -513 255 -513 0 feedthrough
rlabel pdiffusion 262 -513 262 -513 0 feedthrough
rlabel pdiffusion 269 -513 269 -513 0 feedthrough
rlabel pdiffusion 276 -513 276 -513 0 cellNo=318
rlabel pdiffusion 283 -513 283 -513 0 cellNo=11
rlabel pdiffusion 290 -513 290 -513 0 feedthrough
rlabel pdiffusion 297 -513 297 -513 0 feedthrough
rlabel pdiffusion 304 -513 304 -513 0 cellNo=220
rlabel pdiffusion 311 -513 311 -513 0 feedthrough
rlabel pdiffusion 318 -513 318 -513 0 feedthrough
rlabel pdiffusion 325 -513 325 -513 0 feedthrough
rlabel pdiffusion 332 -513 332 -513 0 feedthrough
rlabel pdiffusion 339 -513 339 -513 0 feedthrough
rlabel pdiffusion 346 -513 346 -513 0 feedthrough
rlabel pdiffusion 353 -513 353 -513 0 feedthrough
rlabel pdiffusion 360 -513 360 -513 0 feedthrough
rlabel pdiffusion 367 -513 367 -513 0 cellNo=50
rlabel pdiffusion 374 -513 374 -513 0 feedthrough
rlabel pdiffusion 381 -513 381 -513 0 feedthrough
rlabel pdiffusion 388 -513 388 -513 0 feedthrough
rlabel pdiffusion 402 -513 402 -513 0 feedthrough
rlabel pdiffusion 409 -513 409 -513 0 feedthrough
rlabel pdiffusion 416 -513 416 -513 0 cellNo=12
rlabel pdiffusion 430 -513 430 -513 0 cellNo=242
rlabel pdiffusion 437 -513 437 -513 0 feedthrough
rlabel pdiffusion 444 -513 444 -513 0 cellNo=213
rlabel pdiffusion 451 -513 451 -513 0 feedthrough
rlabel pdiffusion 458 -513 458 -513 0 feedthrough
rlabel pdiffusion 465 -513 465 -513 0 feedthrough
rlabel pdiffusion 10 -566 10 -566 0 feedthrough
rlabel pdiffusion 17 -566 17 -566 0 cellNo=37
rlabel pdiffusion 24 -566 24 -566 0 cellNo=103
rlabel pdiffusion 31 -566 31 -566 0 feedthrough
rlabel pdiffusion 38 -566 38 -566 0 feedthrough
rlabel pdiffusion 45 -566 45 -566 0 feedthrough
rlabel pdiffusion 52 -566 52 -566 0 feedthrough
rlabel pdiffusion 59 -566 59 -566 0 feedthrough
rlabel pdiffusion 66 -566 66 -566 0 cellNo=223
rlabel pdiffusion 73 -566 73 -566 0 feedthrough
rlabel pdiffusion 80 -566 80 -566 0 cellNo=158
rlabel pdiffusion 87 -566 87 -566 0 feedthrough
rlabel pdiffusion 94 -566 94 -566 0 cellNo=134
rlabel pdiffusion 101 -566 101 -566 0 cellNo=264
rlabel pdiffusion 108 -566 108 -566 0 feedthrough
rlabel pdiffusion 115 -566 115 -566 0 cellNo=70
rlabel pdiffusion 122 -566 122 -566 0 cellNo=339
rlabel pdiffusion 129 -566 129 -566 0 feedthrough
rlabel pdiffusion 136 -566 136 -566 0 feedthrough
rlabel pdiffusion 143 -566 143 -566 0 feedthrough
rlabel pdiffusion 150 -566 150 -566 0 feedthrough
rlabel pdiffusion 157 -566 157 -566 0 feedthrough
rlabel pdiffusion 164 -566 164 -566 0 cellNo=175
rlabel pdiffusion 171 -566 171 -566 0 cellNo=346
rlabel pdiffusion 178 -566 178 -566 0 cellNo=185
rlabel pdiffusion 185 -566 185 -566 0 cellNo=113
rlabel pdiffusion 192 -566 192 -566 0 feedthrough
rlabel pdiffusion 199 -566 199 -566 0 feedthrough
rlabel pdiffusion 206 -566 206 -566 0 cellNo=108
rlabel pdiffusion 213 -566 213 -566 0 feedthrough
rlabel pdiffusion 220 -566 220 -566 0 feedthrough
rlabel pdiffusion 227 -566 227 -566 0 feedthrough
rlabel pdiffusion 234 -566 234 -566 0 cellNo=129
rlabel pdiffusion 241 -566 241 -566 0 cellNo=263
rlabel pdiffusion 248 -566 248 -566 0 feedthrough
rlabel pdiffusion 255 -566 255 -566 0 feedthrough
rlabel pdiffusion 262 -566 262 -566 0 feedthrough
rlabel pdiffusion 269 -566 269 -566 0 feedthrough
rlabel pdiffusion 276 -566 276 -566 0 feedthrough
rlabel pdiffusion 283 -566 283 -566 0 cellNo=337
rlabel pdiffusion 290 -566 290 -566 0 feedthrough
rlabel pdiffusion 297 -566 297 -566 0 feedthrough
rlabel pdiffusion 304 -566 304 -566 0 cellNo=212
rlabel pdiffusion 311 -566 311 -566 0 feedthrough
rlabel pdiffusion 318 -566 318 -566 0 feedthrough
rlabel pdiffusion 325 -566 325 -566 0 feedthrough
rlabel pdiffusion 332 -566 332 -566 0 feedthrough
rlabel pdiffusion 339 -566 339 -566 0 cellNo=347
rlabel pdiffusion 346 -566 346 -566 0 feedthrough
rlabel pdiffusion 353 -566 353 -566 0 feedthrough
rlabel pdiffusion 360 -566 360 -566 0 feedthrough
rlabel pdiffusion 367 -566 367 -566 0 feedthrough
rlabel pdiffusion 374 -566 374 -566 0 feedthrough
rlabel pdiffusion 381 -566 381 -566 0 feedthrough
rlabel pdiffusion 388 -566 388 -566 0 feedthrough
rlabel pdiffusion 395 -566 395 -566 0 feedthrough
rlabel pdiffusion 402 -566 402 -566 0 feedthrough
rlabel pdiffusion 409 -566 409 -566 0 feedthrough
rlabel pdiffusion 416 -566 416 -566 0 feedthrough
rlabel pdiffusion 423 -566 423 -566 0 feedthrough
rlabel pdiffusion 430 -566 430 -566 0 feedthrough
rlabel pdiffusion 437 -566 437 -566 0 feedthrough
rlabel pdiffusion 444 -566 444 -566 0 feedthrough
rlabel pdiffusion 458 -566 458 -566 0 cellNo=321
rlabel pdiffusion 465 -566 465 -566 0 feedthrough
rlabel pdiffusion 10 -619 10 -619 0 feedthrough
rlabel pdiffusion 17 -619 17 -619 0 feedthrough
rlabel pdiffusion 24 -619 24 -619 0 feedthrough
rlabel pdiffusion 31 -619 31 -619 0 cellNo=249
rlabel pdiffusion 38 -619 38 -619 0 cellNo=83
rlabel pdiffusion 45 -619 45 -619 0 feedthrough
rlabel pdiffusion 52 -619 52 -619 0 feedthrough
rlabel pdiffusion 59 -619 59 -619 0 feedthrough
rlabel pdiffusion 66 -619 66 -619 0 feedthrough
rlabel pdiffusion 73 -619 73 -619 0 feedthrough
rlabel pdiffusion 80 -619 80 -619 0 feedthrough
rlabel pdiffusion 87 -619 87 -619 0 cellNo=241
rlabel pdiffusion 94 -619 94 -619 0 feedthrough
rlabel pdiffusion 101 -619 101 -619 0 cellNo=101
rlabel pdiffusion 108 -619 108 -619 0 feedthrough
rlabel pdiffusion 115 -619 115 -619 0 cellNo=278
rlabel pdiffusion 122 -619 122 -619 0 feedthrough
rlabel pdiffusion 129 -619 129 -619 0 cellNo=179
rlabel pdiffusion 136 -619 136 -619 0 cellNo=329
rlabel pdiffusion 143 -619 143 -619 0 feedthrough
rlabel pdiffusion 150 -619 150 -619 0 feedthrough
rlabel pdiffusion 157 -619 157 -619 0 feedthrough
rlabel pdiffusion 164 -619 164 -619 0 feedthrough
rlabel pdiffusion 171 -619 171 -619 0 cellNo=36
rlabel pdiffusion 178 -619 178 -619 0 feedthrough
rlabel pdiffusion 185 -619 185 -619 0 feedthrough
rlabel pdiffusion 192 -619 192 -619 0 cellNo=196
rlabel pdiffusion 199 -619 199 -619 0 feedthrough
rlabel pdiffusion 206 -619 206 -619 0 cellNo=181
rlabel pdiffusion 213 -619 213 -619 0 cellNo=257
rlabel pdiffusion 220 -619 220 -619 0 feedthrough
rlabel pdiffusion 227 -619 227 -619 0 feedthrough
rlabel pdiffusion 234 -619 234 -619 0 feedthrough
rlabel pdiffusion 241 -619 241 -619 0 feedthrough
rlabel pdiffusion 248 -619 248 -619 0 cellNo=225
rlabel pdiffusion 255 -619 255 -619 0 cellNo=173
rlabel pdiffusion 262 -619 262 -619 0 cellNo=340
rlabel pdiffusion 269 -619 269 -619 0 feedthrough
rlabel pdiffusion 276 -619 276 -619 0 feedthrough
rlabel pdiffusion 283 -619 283 -619 0 feedthrough
rlabel pdiffusion 290 -619 290 -619 0 feedthrough
rlabel pdiffusion 297 -619 297 -619 0 cellNo=92
rlabel pdiffusion 304 -619 304 -619 0 feedthrough
rlabel pdiffusion 311 -619 311 -619 0 feedthrough
rlabel pdiffusion 318 -619 318 -619 0 feedthrough
rlabel pdiffusion 325 -619 325 -619 0 feedthrough
rlabel pdiffusion 332 -619 332 -619 0 cellNo=192
rlabel pdiffusion 339 -619 339 -619 0 feedthrough
rlabel pdiffusion 346 -619 346 -619 0 feedthrough
rlabel pdiffusion 353 -619 353 -619 0 feedthrough
rlabel pdiffusion 360 -619 360 -619 0 feedthrough
rlabel pdiffusion 367 -619 367 -619 0 feedthrough
rlabel pdiffusion 374 -619 374 -619 0 feedthrough
rlabel pdiffusion 381 -619 381 -619 0 feedthrough
rlabel pdiffusion 388 -619 388 -619 0 feedthrough
rlabel pdiffusion 395 -619 395 -619 0 feedthrough
rlabel pdiffusion 402 -619 402 -619 0 feedthrough
rlabel pdiffusion 409 -619 409 -619 0 feedthrough
rlabel pdiffusion 416 -619 416 -619 0 feedthrough
rlabel pdiffusion 423 -619 423 -619 0 feedthrough
rlabel pdiffusion 430 -619 430 -619 0 feedthrough
rlabel pdiffusion 437 -619 437 -619 0 feedthrough
rlabel pdiffusion 444 -619 444 -619 0 cellNo=147
rlabel pdiffusion 451 -619 451 -619 0 cellNo=29
rlabel pdiffusion 458 -619 458 -619 0 feedthrough
rlabel pdiffusion 465 -619 465 -619 0 cellNo=177
rlabel pdiffusion 472 -619 472 -619 0 feedthrough
rlabel pdiffusion 3 -670 3 -670 0 feedthrough
rlabel pdiffusion 10 -670 10 -670 0 feedthrough
rlabel pdiffusion 17 -670 17 -670 0 feedthrough
rlabel pdiffusion 24 -670 24 -670 0 feedthrough
rlabel pdiffusion 31 -670 31 -670 0 feedthrough
rlabel pdiffusion 38 -670 38 -670 0 feedthrough
rlabel pdiffusion 45 -670 45 -670 0 cellNo=338
rlabel pdiffusion 52 -670 52 -670 0 cellNo=216
rlabel pdiffusion 59 -670 59 -670 0 feedthrough
rlabel pdiffusion 66 -670 66 -670 0 feedthrough
rlabel pdiffusion 73 -670 73 -670 0 cellNo=123
rlabel pdiffusion 80 -670 80 -670 0 feedthrough
rlabel pdiffusion 87 -670 87 -670 0 feedthrough
rlabel pdiffusion 94 -670 94 -670 0 feedthrough
rlabel pdiffusion 101 -670 101 -670 0 cellNo=334
rlabel pdiffusion 108 -670 108 -670 0 feedthrough
rlabel pdiffusion 115 -670 115 -670 0 cellNo=293
rlabel pdiffusion 122 -670 122 -670 0 feedthrough
rlabel pdiffusion 129 -670 129 -670 0 cellNo=169
rlabel pdiffusion 136 -670 136 -670 0 feedthrough
rlabel pdiffusion 143 -670 143 -670 0 feedthrough
rlabel pdiffusion 150 -670 150 -670 0 feedthrough
rlabel pdiffusion 157 -670 157 -670 0 feedthrough
rlabel pdiffusion 164 -670 164 -670 0 feedthrough
rlabel pdiffusion 171 -670 171 -670 0 feedthrough
rlabel pdiffusion 178 -670 178 -670 0 cellNo=86
rlabel pdiffusion 185 -670 185 -670 0 cellNo=84
rlabel pdiffusion 192 -670 192 -670 0 cellNo=60
rlabel pdiffusion 199 -670 199 -670 0 feedthrough
rlabel pdiffusion 206 -670 206 -670 0 cellNo=178
rlabel pdiffusion 213 -670 213 -670 0 cellNo=160
rlabel pdiffusion 220 -670 220 -670 0 cellNo=20
rlabel pdiffusion 227 -670 227 -670 0 feedthrough
rlabel pdiffusion 234 -670 234 -670 0 feedthrough
rlabel pdiffusion 241 -670 241 -670 0 cellNo=224
rlabel pdiffusion 248 -670 248 -670 0 cellNo=187
rlabel pdiffusion 255 -670 255 -670 0 feedthrough
rlabel pdiffusion 262 -670 262 -670 0 feedthrough
rlabel pdiffusion 269 -670 269 -670 0 cellNo=165
rlabel pdiffusion 276 -670 276 -670 0 feedthrough
rlabel pdiffusion 283 -670 283 -670 0 feedthrough
rlabel pdiffusion 290 -670 290 -670 0 feedthrough
rlabel pdiffusion 297 -670 297 -670 0 cellNo=271
rlabel pdiffusion 304 -670 304 -670 0 feedthrough
rlabel pdiffusion 311 -670 311 -670 0 feedthrough
rlabel pdiffusion 318 -670 318 -670 0 feedthrough
rlabel pdiffusion 325 -670 325 -670 0 feedthrough
rlabel pdiffusion 332 -670 332 -670 0 cellNo=336
rlabel pdiffusion 339 -670 339 -670 0 feedthrough
rlabel pdiffusion 346 -670 346 -670 0 feedthrough
rlabel pdiffusion 353 -670 353 -670 0 feedthrough
rlabel pdiffusion 360 -670 360 -670 0 feedthrough
rlabel pdiffusion 367 -670 367 -670 0 feedthrough
rlabel pdiffusion 374 -670 374 -670 0 feedthrough
rlabel pdiffusion 381 -670 381 -670 0 feedthrough
rlabel pdiffusion 388 -670 388 -670 0 feedthrough
rlabel pdiffusion 395 -670 395 -670 0 feedthrough
rlabel pdiffusion 402 -670 402 -670 0 feedthrough
rlabel pdiffusion 409 -670 409 -670 0 feedthrough
rlabel pdiffusion 416 -670 416 -670 0 feedthrough
rlabel pdiffusion 423 -670 423 -670 0 feedthrough
rlabel pdiffusion 430 -670 430 -670 0 feedthrough
rlabel pdiffusion 437 -670 437 -670 0 feedthrough
rlabel pdiffusion 444 -670 444 -670 0 feedthrough
rlabel pdiffusion 451 -670 451 -670 0 feedthrough
rlabel pdiffusion 458 -670 458 -670 0 cellNo=1
rlabel pdiffusion 465 -670 465 -670 0 cellNo=228
rlabel pdiffusion 472 -670 472 -670 0 feedthrough
rlabel pdiffusion 3 -721 3 -721 0 feedthrough
rlabel pdiffusion 10 -721 10 -721 0 feedthrough
rlabel pdiffusion 17 -721 17 -721 0 feedthrough
rlabel pdiffusion 24 -721 24 -721 0 feedthrough
rlabel pdiffusion 31 -721 31 -721 0 feedthrough
rlabel pdiffusion 38 -721 38 -721 0 cellNo=65
rlabel pdiffusion 45 -721 45 -721 0 feedthrough
rlabel pdiffusion 52 -721 52 -721 0 cellNo=79
rlabel pdiffusion 59 -721 59 -721 0 feedthrough
rlabel pdiffusion 66 -721 66 -721 0 feedthrough
rlabel pdiffusion 73 -721 73 -721 0 cellNo=116
rlabel pdiffusion 80 -721 80 -721 0 cellNo=203
rlabel pdiffusion 87 -721 87 -721 0 feedthrough
rlabel pdiffusion 94 -721 94 -721 0 feedthrough
rlabel pdiffusion 101 -721 101 -721 0 feedthrough
rlabel pdiffusion 108 -721 108 -721 0 feedthrough
rlabel pdiffusion 115 -721 115 -721 0 feedthrough
rlabel pdiffusion 122 -721 122 -721 0 cellNo=309
rlabel pdiffusion 129 -721 129 -721 0 cellNo=262
rlabel pdiffusion 136 -721 136 -721 0 feedthrough
rlabel pdiffusion 143 -721 143 -721 0 feedthrough
rlabel pdiffusion 150 -721 150 -721 0 feedthrough
rlabel pdiffusion 157 -721 157 -721 0 feedthrough
rlabel pdiffusion 164 -721 164 -721 0 feedthrough
rlabel pdiffusion 171 -721 171 -721 0 cellNo=283
rlabel pdiffusion 178 -721 178 -721 0 cellNo=275
rlabel pdiffusion 185 -721 185 -721 0 cellNo=77
rlabel pdiffusion 192 -721 192 -721 0 feedthrough
rlabel pdiffusion 199 -721 199 -721 0 cellNo=345
rlabel pdiffusion 206 -721 206 -721 0 cellNo=72
rlabel pdiffusion 213 -721 213 -721 0 feedthrough
rlabel pdiffusion 220 -721 220 -721 0 feedthrough
rlabel pdiffusion 227 -721 227 -721 0 cellNo=342
rlabel pdiffusion 234 -721 234 -721 0 feedthrough
rlabel pdiffusion 241 -721 241 -721 0 cellNo=306
rlabel pdiffusion 248 -721 248 -721 0 cellNo=327
rlabel pdiffusion 255 -721 255 -721 0 feedthrough
rlabel pdiffusion 262 -721 262 -721 0 feedthrough
rlabel pdiffusion 269 -721 269 -721 0 feedthrough
rlabel pdiffusion 276 -721 276 -721 0 cellNo=307
rlabel pdiffusion 283 -721 283 -721 0 feedthrough
rlabel pdiffusion 290 -721 290 -721 0 feedthrough
rlabel pdiffusion 297 -721 297 -721 0 cellNo=247
rlabel pdiffusion 311 -721 311 -721 0 feedthrough
rlabel pdiffusion 318 -721 318 -721 0 feedthrough
rlabel pdiffusion 325 -721 325 -721 0 feedthrough
rlabel pdiffusion 332 -721 332 -721 0 feedthrough
rlabel pdiffusion 339 -721 339 -721 0 cellNo=182
rlabel pdiffusion 346 -721 346 -721 0 feedthrough
rlabel pdiffusion 353 -721 353 -721 0 feedthrough
rlabel pdiffusion 360 -721 360 -721 0 feedthrough
rlabel pdiffusion 367 -721 367 -721 0 feedthrough
rlabel pdiffusion 374 -721 374 -721 0 cellNo=144
rlabel pdiffusion 381 -721 381 -721 0 feedthrough
rlabel pdiffusion 388 -721 388 -721 0 feedthrough
rlabel pdiffusion 395 -721 395 -721 0 feedthrough
rlabel pdiffusion 402 -721 402 -721 0 feedthrough
rlabel pdiffusion 409 -721 409 -721 0 cellNo=14
rlabel pdiffusion 430 -721 430 -721 0 feedthrough
rlabel pdiffusion 17 -774 17 -774 0 cellNo=292
rlabel pdiffusion 24 -774 24 -774 0 feedthrough
rlabel pdiffusion 31 -774 31 -774 0 cellNo=104
rlabel pdiffusion 38 -774 38 -774 0 cellNo=269
rlabel pdiffusion 45 -774 45 -774 0 cellNo=189
rlabel pdiffusion 52 -774 52 -774 0 feedthrough
rlabel pdiffusion 59 -774 59 -774 0 feedthrough
rlabel pdiffusion 66 -774 66 -774 0 feedthrough
rlabel pdiffusion 73 -774 73 -774 0 cellNo=317
rlabel pdiffusion 80 -774 80 -774 0 cellNo=26
rlabel pdiffusion 87 -774 87 -774 0 feedthrough
rlabel pdiffusion 94 -774 94 -774 0 cellNo=124
rlabel pdiffusion 101 -774 101 -774 0 cellNo=349
rlabel pdiffusion 108 -774 108 -774 0 cellNo=301
rlabel pdiffusion 115 -774 115 -774 0 cellNo=73
rlabel pdiffusion 122 -774 122 -774 0 cellNo=331
rlabel pdiffusion 129 -774 129 -774 0 feedthrough
rlabel pdiffusion 136 -774 136 -774 0 feedthrough
rlabel pdiffusion 143 -774 143 -774 0 feedthrough
rlabel pdiffusion 150 -774 150 -774 0 feedthrough
rlabel pdiffusion 157 -774 157 -774 0 feedthrough
rlabel pdiffusion 164 -774 164 -774 0 feedthrough
rlabel pdiffusion 171 -774 171 -774 0 feedthrough
rlabel pdiffusion 178 -774 178 -774 0 cellNo=280
rlabel pdiffusion 185 -774 185 -774 0 feedthrough
rlabel pdiffusion 192 -774 192 -774 0 feedthrough
rlabel pdiffusion 199 -774 199 -774 0 cellNo=351
rlabel pdiffusion 206 -774 206 -774 0 cellNo=191
rlabel pdiffusion 213 -774 213 -774 0 cellNo=260
rlabel pdiffusion 220 -774 220 -774 0 feedthrough
rlabel pdiffusion 227 -774 227 -774 0 feedthrough
rlabel pdiffusion 234 -774 234 -774 0 cellNo=171
rlabel pdiffusion 241 -774 241 -774 0 feedthrough
rlabel pdiffusion 248 -774 248 -774 0 feedthrough
rlabel pdiffusion 255 -774 255 -774 0 feedthrough
rlabel pdiffusion 262 -774 262 -774 0 feedthrough
rlabel pdiffusion 269 -774 269 -774 0 feedthrough
rlabel pdiffusion 276 -774 276 -774 0 cellNo=273
rlabel pdiffusion 283 -774 283 -774 0 feedthrough
rlabel pdiffusion 290 -774 290 -774 0 feedthrough
rlabel pdiffusion 304 -774 304 -774 0 feedthrough
rlabel pdiffusion 311 -774 311 -774 0 feedthrough
rlabel pdiffusion 325 -774 325 -774 0 feedthrough
rlabel pdiffusion 332 -774 332 -774 0 cellNo=344
rlabel pdiffusion 339 -774 339 -774 0 feedthrough
rlabel pdiffusion 346 -774 346 -774 0 feedthrough
rlabel pdiffusion 409 -774 409 -774 0 cellNo=303
rlabel pdiffusion 10 -819 10 -819 0 feedthrough
rlabel pdiffusion 17 -819 17 -819 0 cellNo=157
rlabel pdiffusion 24 -819 24 -819 0 feedthrough
rlabel pdiffusion 31 -819 31 -819 0 cellNo=248
rlabel pdiffusion 38 -819 38 -819 0 feedthrough
rlabel pdiffusion 45 -819 45 -819 0 cellNo=258
rlabel pdiffusion 52 -819 52 -819 0 cellNo=322
rlabel pdiffusion 59 -819 59 -819 0 cellNo=291
rlabel pdiffusion 66 -819 66 -819 0 cellNo=279
rlabel pdiffusion 73 -819 73 -819 0 feedthrough
rlabel pdiffusion 80 -819 80 -819 0 cellNo=323
rlabel pdiffusion 87 -819 87 -819 0 cellNo=205
rlabel pdiffusion 94 -819 94 -819 0 cellNo=140
rlabel pdiffusion 101 -819 101 -819 0 feedthrough
rlabel pdiffusion 108 -819 108 -819 0 cellNo=138
rlabel pdiffusion 115 -819 115 -819 0 cellNo=299
rlabel pdiffusion 122 -819 122 -819 0 cellNo=308
rlabel pdiffusion 129 -819 129 -819 0 cellNo=352
rlabel pdiffusion 136 -819 136 -819 0 feedthrough
rlabel pdiffusion 143 -819 143 -819 0 cellNo=58
rlabel pdiffusion 150 -819 150 -819 0 cellNo=320
rlabel pdiffusion 157 -819 157 -819 0 feedthrough
rlabel pdiffusion 164 -819 164 -819 0 feedthrough
rlabel pdiffusion 171 -819 171 -819 0 feedthrough
rlabel pdiffusion 178 -819 178 -819 0 cellNo=350
rlabel pdiffusion 185 -819 185 -819 0 feedthrough
rlabel pdiffusion 192 -819 192 -819 0 feedthrough
rlabel pdiffusion 199 -819 199 -819 0 feedthrough
rlabel pdiffusion 206 -819 206 -819 0 feedthrough
rlabel pdiffusion 213 -819 213 -819 0 feedthrough
rlabel pdiffusion 220 -819 220 -819 0 cellNo=106
rlabel pdiffusion 227 -819 227 -819 0 feedthrough
rlabel pdiffusion 234 -819 234 -819 0 feedthrough
rlabel pdiffusion 241 -819 241 -819 0 cellNo=215
rlabel pdiffusion 248 -819 248 -819 0 feedthrough
rlabel pdiffusion 255 -819 255 -819 0 feedthrough
rlabel pdiffusion 262 -819 262 -819 0 feedthrough
rlabel pdiffusion 269 -819 269 -819 0 feedthrough
rlabel pdiffusion 283 -819 283 -819 0 feedthrough
rlabel pdiffusion 290 -819 290 -819 0 feedthrough
rlabel pdiffusion 304 -819 304 -819 0 feedthrough
rlabel pdiffusion 311 -819 311 -819 0 feedthrough
rlabel pdiffusion 318 -819 318 -819 0 feedthrough
rlabel pdiffusion 325 -819 325 -819 0 feedthrough
rlabel pdiffusion 346 -819 346 -819 0 cellNo=23
rlabel pdiffusion 17 -852 17 -852 0 cellNo=206
rlabel pdiffusion 24 -852 24 -852 0 feedthrough
rlabel pdiffusion 31 -852 31 -852 0 cellNo=195
rlabel pdiffusion 38 -852 38 -852 0 feedthrough
rlabel pdiffusion 45 -852 45 -852 0 cellNo=230
rlabel pdiffusion 52 -852 52 -852 0 cellNo=360
rlabel pdiffusion 59 -852 59 -852 0 feedthrough
rlabel pdiffusion 66 -852 66 -852 0 cellNo=209
rlabel pdiffusion 73 -852 73 -852 0 feedthrough
rlabel pdiffusion 80 -852 80 -852 0 cellNo=153
rlabel pdiffusion 87 -852 87 -852 0 feedthrough
rlabel pdiffusion 94 -852 94 -852 0 feedthrough
rlabel pdiffusion 101 -852 101 -852 0 cellNo=117
rlabel pdiffusion 108 -852 108 -852 0 cellNo=137
rlabel pdiffusion 115 -852 115 -852 0 cellNo=85
rlabel pdiffusion 122 -852 122 -852 0 cellNo=295
rlabel pdiffusion 129 -852 129 -852 0 cellNo=18
rlabel pdiffusion 136 -852 136 -852 0 cellNo=305
rlabel pdiffusion 143 -852 143 -852 0 cellNo=59
rlabel pdiffusion 150 -852 150 -852 0 feedthrough
rlabel pdiffusion 157 -852 157 -852 0 feedthrough
rlabel pdiffusion 164 -852 164 -852 0 feedthrough
rlabel pdiffusion 171 -852 171 -852 0 feedthrough
rlabel pdiffusion 185 -852 185 -852 0 cellNo=354
rlabel pdiffusion 192 -852 192 -852 0 feedthrough
rlabel pdiffusion 213 -852 213 -852 0 cellNo=304
rlabel pdiffusion 227 -852 227 -852 0 cellNo=167
rlabel pdiffusion 269 -852 269 -852 0 feedthrough
rlabel pdiffusion 283 -852 283 -852 0 cellNo=237
rlabel pdiffusion 290 -852 290 -852 0 cellNo=356
rlabel pdiffusion 325 -852 325 -852 0 cellNo=61
rlabel polysilicon 12 -6 12 -6 0 2
rlabel polysilicon 26 -6 26 -6 0 2
rlabel polysilicon 37 -6 37 -6 0 1
rlabel polysilicon 51 -6 51 -6 0 1
rlabel polysilicon 58 -6 58 -6 0 1
rlabel polysilicon 65 -6 65 -6 0 1
rlabel polysilicon 65 -12 65 -12 0 3
rlabel polysilicon 72 -6 72 -6 0 1
rlabel polysilicon 72 -12 72 -12 0 3
rlabel polysilicon 89 -6 89 -6 0 2
rlabel polysilicon 93 -6 93 -6 0 1
rlabel polysilicon 96 -12 96 -12 0 4
rlabel polysilicon 100 -12 100 -12 0 3
rlabel polysilicon 107 -6 107 -6 0 1
rlabel polysilicon 107 -12 107 -12 0 3
rlabel polysilicon 114 -12 114 -12 0 3
rlabel polysilicon 121 -6 121 -6 0 1
rlabel polysilicon 128 -6 128 -6 0 1
rlabel polysilicon 128 -12 128 -12 0 3
rlabel polysilicon 135 -6 135 -6 0 1
rlabel polysilicon 138 -6 138 -6 0 2
rlabel polysilicon 145 -12 145 -12 0 4
rlabel polysilicon 149 -6 149 -6 0 1
rlabel polysilicon 149 -12 149 -12 0 3
rlabel polysilicon 156 -12 156 -12 0 3
rlabel polysilicon 159 -12 159 -12 0 4
rlabel polysilicon 163 -6 163 -6 0 1
rlabel polysilicon 163 -12 163 -12 0 3
rlabel polysilicon 5 -31 5 -31 0 4
rlabel polysilicon 30 -31 30 -31 0 3
rlabel polysilicon 37 -31 37 -31 0 3
rlabel polysilicon 72 -25 72 -25 0 1
rlabel polysilicon 72 -31 72 -31 0 3
rlabel polysilicon 79 -25 79 -25 0 1
rlabel polysilicon 93 -31 93 -31 0 3
rlabel polysilicon 100 -25 100 -25 0 1
rlabel polysilicon 107 -25 107 -25 0 1
rlabel polysilicon 114 -25 114 -25 0 1
rlabel polysilicon 117 -31 117 -31 0 4
rlabel polysilicon 124 -31 124 -31 0 4
rlabel polysilicon 128 -25 128 -25 0 1
rlabel polysilicon 128 -31 128 -31 0 3
rlabel polysilicon 142 -25 142 -25 0 1
rlabel polysilicon 142 -31 142 -31 0 3
rlabel polysilicon 149 -25 149 -25 0 1
rlabel polysilicon 149 -31 149 -31 0 3
rlabel polysilicon 163 -25 163 -25 0 1
rlabel polysilicon 163 -31 163 -31 0 3
rlabel polysilicon 173 -25 173 -25 0 2
rlabel polysilicon 177 -25 177 -25 0 1
rlabel polysilicon 177 -31 177 -31 0 3
rlabel polysilicon 187 -25 187 -25 0 2
rlabel polysilicon 191 -25 191 -25 0 1
rlabel polysilicon 191 -31 191 -31 0 3
rlabel polysilicon 201 -25 201 -25 0 2
rlabel polysilicon 198 -31 198 -31 0 3
rlabel polysilicon 5 -56 5 -56 0 2
rlabel polysilicon 16 -56 16 -56 0 1
rlabel polysilicon 30 -56 30 -56 0 1
rlabel polysilicon 30 -62 30 -62 0 3
rlabel polysilicon 40 -62 40 -62 0 4
rlabel polysilicon 47 -56 47 -56 0 2
rlabel polysilicon 51 -56 51 -56 0 1
rlabel polysilicon 51 -62 51 -62 0 3
rlabel polysilicon 58 -56 58 -56 0 1
rlabel polysilicon 58 -62 58 -62 0 3
rlabel polysilicon 65 -56 65 -56 0 1
rlabel polysilicon 65 -62 65 -62 0 3
rlabel polysilicon 72 -56 72 -56 0 1
rlabel polysilicon 72 -62 72 -62 0 3
rlabel polysilicon 79 -56 79 -56 0 1
rlabel polysilicon 82 -62 82 -62 0 4
rlabel polysilicon 86 -56 86 -56 0 1
rlabel polysilicon 89 -62 89 -62 0 4
rlabel polysilicon 93 -56 93 -56 0 1
rlabel polysilicon 96 -56 96 -56 0 2
rlabel polysilicon 100 -56 100 -56 0 1
rlabel polysilicon 100 -62 100 -62 0 3
rlabel polysilicon 107 -62 107 -62 0 3
rlabel polysilicon 110 -62 110 -62 0 4
rlabel polysilicon 114 -62 114 -62 0 3
rlabel polysilicon 121 -56 121 -56 0 1
rlabel polysilicon 124 -56 124 -56 0 2
rlabel polysilicon 128 -56 128 -56 0 1
rlabel polysilicon 128 -62 128 -62 0 3
rlabel polysilicon 131 -62 131 -62 0 4
rlabel polysilicon 135 -62 135 -62 0 3
rlabel polysilicon 145 -56 145 -56 0 2
rlabel polysilicon 149 -56 149 -56 0 1
rlabel polysilicon 152 -56 152 -56 0 2
rlabel polysilicon 156 -56 156 -56 0 1
rlabel polysilicon 156 -62 156 -62 0 3
rlabel polysilicon 163 -56 163 -56 0 1
rlabel polysilicon 163 -62 163 -62 0 3
rlabel polysilicon 170 -56 170 -56 0 1
rlabel polysilicon 170 -62 170 -62 0 3
rlabel polysilicon 177 -56 177 -56 0 1
rlabel polysilicon 177 -62 177 -62 0 3
rlabel polysilicon 184 -56 184 -56 0 1
rlabel polysilicon 184 -62 184 -62 0 3
rlabel polysilicon 191 -62 191 -62 0 3
rlabel polysilicon 198 -56 198 -56 0 1
rlabel polysilicon 198 -62 198 -62 0 3
rlabel polysilicon 205 -56 205 -56 0 1
rlabel polysilicon 205 -62 205 -62 0 3
rlabel polysilicon 212 -56 212 -56 0 1
rlabel polysilicon 212 -62 212 -62 0 3
rlabel polysilicon 219 -56 219 -56 0 1
rlabel polysilicon 219 -62 219 -62 0 3
rlabel polysilicon 226 -56 226 -56 0 1
rlabel polysilicon 226 -62 226 -62 0 3
rlabel polysilicon 233 -56 233 -56 0 1
rlabel polysilicon 233 -62 233 -62 0 3
rlabel polysilicon 243 -62 243 -62 0 4
rlabel polysilicon 247 -56 247 -56 0 1
rlabel polysilicon 247 -62 247 -62 0 3
rlabel polysilicon 254 -56 254 -56 0 1
rlabel polysilicon 254 -62 254 -62 0 3
rlabel polysilicon 9 -95 9 -95 0 3
rlabel polysilicon 19 -89 19 -89 0 2
rlabel polysilicon 23 -95 23 -95 0 3
rlabel polysilicon 30 -89 30 -89 0 1
rlabel polysilicon 30 -95 30 -95 0 3
rlabel polysilicon 40 -89 40 -89 0 2
rlabel polysilicon 44 -89 44 -89 0 1
rlabel polysilicon 44 -95 44 -95 0 3
rlabel polysilicon 51 -89 51 -89 0 1
rlabel polysilicon 51 -95 51 -95 0 3
rlabel polysilicon 58 -89 58 -89 0 1
rlabel polysilicon 58 -95 58 -95 0 3
rlabel polysilicon 65 -89 65 -89 0 1
rlabel polysilicon 65 -95 65 -95 0 3
rlabel polysilicon 72 -89 72 -89 0 1
rlabel polysilicon 72 -95 72 -95 0 3
rlabel polysilicon 79 -89 79 -89 0 1
rlabel polysilicon 86 -89 86 -89 0 1
rlabel polysilicon 86 -95 86 -95 0 3
rlabel polysilicon 96 -89 96 -89 0 2
rlabel polysilicon 96 -95 96 -95 0 4
rlabel polysilicon 100 -89 100 -89 0 1
rlabel polysilicon 110 -89 110 -89 0 2
rlabel polysilicon 117 -95 117 -95 0 4
rlabel polysilicon 121 -89 121 -89 0 1
rlabel polysilicon 121 -95 121 -95 0 3
rlabel polysilicon 131 -89 131 -89 0 2
rlabel polysilicon 128 -95 128 -95 0 3
rlabel polysilicon 131 -95 131 -95 0 4
rlabel polysilicon 138 -89 138 -89 0 2
rlabel polysilicon 135 -95 135 -95 0 3
rlabel polysilicon 138 -95 138 -95 0 4
rlabel polysilicon 142 -89 142 -89 0 1
rlabel polysilicon 145 -95 145 -95 0 4
rlabel polysilicon 149 -89 149 -89 0 1
rlabel polysilicon 149 -95 149 -95 0 3
rlabel polysilicon 159 -89 159 -89 0 2
rlabel polysilicon 156 -95 156 -95 0 3
rlabel polysilicon 163 -95 163 -95 0 3
rlabel polysilicon 166 -95 166 -95 0 4
rlabel polysilicon 170 -89 170 -89 0 1
rlabel polysilicon 173 -95 173 -95 0 4
rlabel polysilicon 177 -89 177 -89 0 1
rlabel polysilicon 177 -95 177 -95 0 3
rlabel polysilicon 184 -89 184 -89 0 1
rlabel polysilicon 191 -89 191 -89 0 1
rlabel polysilicon 191 -95 191 -95 0 3
rlabel polysilicon 198 -95 198 -95 0 3
rlabel polysilicon 201 -95 201 -95 0 4
rlabel polysilicon 205 -89 205 -89 0 1
rlabel polysilicon 205 -95 205 -95 0 3
rlabel polysilicon 212 -89 212 -89 0 1
rlabel polysilicon 212 -95 212 -95 0 3
rlabel polysilicon 219 -89 219 -89 0 1
rlabel polysilicon 219 -95 219 -95 0 3
rlabel polysilicon 226 -89 226 -89 0 1
rlabel polysilicon 226 -95 226 -95 0 3
rlabel polysilicon 233 -89 233 -89 0 1
rlabel polysilicon 233 -95 233 -95 0 3
rlabel polysilicon 240 -89 240 -89 0 1
rlabel polysilicon 240 -95 240 -95 0 3
rlabel polysilicon 247 -89 247 -89 0 1
rlabel polysilicon 247 -95 247 -95 0 3
rlabel polysilicon 254 -89 254 -89 0 1
rlabel polysilicon 254 -95 254 -95 0 3
rlabel polysilicon 261 -89 261 -89 0 1
rlabel polysilicon 261 -95 261 -95 0 3
rlabel polysilicon 268 -89 268 -89 0 1
rlabel polysilicon 268 -95 268 -95 0 3
rlabel polysilicon 275 -89 275 -89 0 1
rlabel polysilicon 275 -95 275 -95 0 3
rlabel polysilicon 282 -89 282 -89 0 1
rlabel polysilicon 282 -95 282 -95 0 3
rlabel polysilicon 289 -89 289 -89 0 1
rlabel polysilicon 289 -95 289 -95 0 3
rlabel polysilicon 296 -89 296 -89 0 1
rlabel polysilicon 296 -95 296 -95 0 3
rlabel polysilicon 303 -95 303 -95 0 3
rlabel polysilicon 331 -89 331 -89 0 1
rlabel polysilicon 331 -95 331 -95 0 3
rlabel polysilicon 16 -150 16 -150 0 3
rlabel polysilicon 19 -150 19 -150 0 4
rlabel polysilicon 26 -144 26 -144 0 2
rlabel polysilicon 23 -150 23 -150 0 3
rlabel polysilicon 30 -144 30 -144 0 1
rlabel polysilicon 30 -150 30 -150 0 3
rlabel polysilicon 37 -144 37 -144 0 1
rlabel polysilicon 37 -150 37 -150 0 3
rlabel polysilicon 44 -144 44 -144 0 1
rlabel polysilicon 44 -150 44 -150 0 3
rlabel polysilicon 51 -144 51 -144 0 1
rlabel polysilicon 51 -150 51 -150 0 3
rlabel polysilicon 58 -144 58 -144 0 1
rlabel polysilicon 58 -150 58 -150 0 3
rlabel polysilicon 61 -150 61 -150 0 4
rlabel polysilicon 65 -144 65 -144 0 1
rlabel polysilicon 65 -150 65 -150 0 3
rlabel polysilicon 72 -144 72 -144 0 1
rlabel polysilicon 72 -150 72 -150 0 3
rlabel polysilicon 79 -150 79 -150 0 3
rlabel polysilicon 82 -150 82 -150 0 4
rlabel polysilicon 86 -144 86 -144 0 1
rlabel polysilicon 86 -150 86 -150 0 3
rlabel polysilicon 89 -150 89 -150 0 4
rlabel polysilicon 93 -144 93 -144 0 1
rlabel polysilicon 93 -150 93 -150 0 3
rlabel polysilicon 100 -144 100 -144 0 1
rlabel polysilicon 100 -150 100 -150 0 3
rlabel polysilicon 107 -144 107 -144 0 1
rlabel polysilicon 107 -150 107 -150 0 3
rlabel polysilicon 114 -150 114 -150 0 3
rlabel polysilicon 121 -144 121 -144 0 1
rlabel polysilicon 124 -144 124 -144 0 2
rlabel polysilicon 121 -150 121 -150 0 3
rlabel polysilicon 128 -144 128 -144 0 1
rlabel polysilicon 128 -150 128 -150 0 3
rlabel polysilicon 138 -144 138 -144 0 2
rlabel polysilicon 135 -150 135 -150 0 3
rlabel polysilicon 142 -144 142 -144 0 1
rlabel polysilicon 142 -150 142 -150 0 3
rlabel polysilicon 149 -144 149 -144 0 1
rlabel polysilicon 152 -144 152 -144 0 2
rlabel polysilicon 149 -150 149 -150 0 3
rlabel polysilicon 152 -150 152 -150 0 4
rlabel polysilicon 156 -144 156 -144 0 1
rlabel polysilicon 156 -150 156 -150 0 3
rlabel polysilicon 163 -144 163 -144 0 1
rlabel polysilicon 166 -144 166 -144 0 2
rlabel polysilicon 163 -150 163 -150 0 3
rlabel polysilicon 170 -144 170 -144 0 1
rlabel polysilicon 170 -150 170 -150 0 3
rlabel polysilicon 177 -144 177 -144 0 1
rlabel polysilicon 177 -150 177 -150 0 3
rlabel polysilicon 184 -144 184 -144 0 1
rlabel polysilicon 184 -150 184 -150 0 3
rlabel polysilicon 194 -144 194 -144 0 2
rlabel polysilicon 191 -150 191 -150 0 3
rlabel polysilicon 194 -150 194 -150 0 4
rlabel polysilicon 201 -144 201 -144 0 2
rlabel polysilicon 198 -150 198 -150 0 3
rlabel polysilicon 208 -144 208 -144 0 2
rlabel polysilicon 205 -150 205 -150 0 3
rlabel polysilicon 208 -150 208 -150 0 4
rlabel polysilicon 212 -144 212 -144 0 1
rlabel polysilicon 212 -150 212 -150 0 3
rlabel polysilicon 219 -144 219 -144 0 1
rlabel polysilicon 219 -150 219 -150 0 3
rlabel polysilicon 226 -144 226 -144 0 1
rlabel polysilicon 226 -150 226 -150 0 3
rlabel polysilicon 233 -144 233 -144 0 1
rlabel polysilicon 233 -150 233 -150 0 3
rlabel polysilicon 240 -144 240 -144 0 1
rlabel polysilicon 240 -150 240 -150 0 3
rlabel polysilicon 247 -144 247 -144 0 1
rlabel polysilicon 247 -150 247 -150 0 3
rlabel polysilicon 254 -144 254 -144 0 1
rlabel polysilicon 254 -150 254 -150 0 3
rlabel polysilicon 261 -144 261 -144 0 1
rlabel polysilicon 261 -150 261 -150 0 3
rlabel polysilicon 271 -144 271 -144 0 2
rlabel polysilicon 268 -150 268 -150 0 3
rlabel polysilicon 275 -144 275 -144 0 1
rlabel polysilicon 275 -150 275 -150 0 3
rlabel polysilicon 282 -144 282 -144 0 1
rlabel polysilicon 282 -150 282 -150 0 3
rlabel polysilicon 289 -144 289 -144 0 1
rlabel polysilicon 289 -150 289 -150 0 3
rlabel polysilicon 296 -144 296 -144 0 1
rlabel polysilicon 296 -150 296 -150 0 3
rlabel polysilicon 303 -144 303 -144 0 1
rlabel polysilicon 303 -150 303 -150 0 3
rlabel polysilicon 310 -144 310 -144 0 1
rlabel polysilicon 310 -150 310 -150 0 3
rlabel polysilicon 317 -144 317 -144 0 1
rlabel polysilicon 317 -150 317 -150 0 3
rlabel polysilicon 324 -144 324 -144 0 1
rlabel polysilicon 324 -150 324 -150 0 3
rlabel polysilicon 331 -144 331 -144 0 1
rlabel polysilicon 331 -150 331 -150 0 3
rlabel polysilicon 338 -144 338 -144 0 1
rlabel polysilicon 338 -150 338 -150 0 3
rlabel polysilicon 345 -144 345 -144 0 1
rlabel polysilicon 345 -150 345 -150 0 3
rlabel polysilicon 352 -144 352 -144 0 1
rlabel polysilicon 352 -150 352 -150 0 3
rlabel polysilicon 359 -144 359 -144 0 1
rlabel polysilicon 359 -150 359 -150 0 3
rlabel polysilicon 366 -144 366 -144 0 1
rlabel polysilicon 366 -150 366 -150 0 3
rlabel polysilicon 373 -144 373 -144 0 1
rlabel polysilicon 373 -150 373 -150 0 3
rlabel polysilicon 5 -195 5 -195 0 2
rlabel polysilicon 9 -195 9 -195 0 1
rlabel polysilicon 9 -201 9 -201 0 3
rlabel polysilicon 16 -195 16 -195 0 1
rlabel polysilicon 16 -201 16 -201 0 3
rlabel polysilicon 23 -195 23 -195 0 1
rlabel polysilicon 26 -195 26 -195 0 2
rlabel polysilicon 30 -195 30 -195 0 1
rlabel polysilicon 30 -201 30 -201 0 3
rlabel polysilicon 37 -195 37 -195 0 1
rlabel polysilicon 37 -201 37 -201 0 3
rlabel polysilicon 47 -195 47 -195 0 2
rlabel polysilicon 44 -201 44 -201 0 3
rlabel polysilicon 51 -195 51 -195 0 1
rlabel polysilicon 51 -201 51 -201 0 3
rlabel polysilicon 61 -195 61 -195 0 2
rlabel polysilicon 58 -201 58 -201 0 3
rlabel polysilicon 65 -195 65 -195 0 1
rlabel polysilicon 65 -201 65 -201 0 3
rlabel polysilicon 72 -195 72 -195 0 1
rlabel polysilicon 75 -195 75 -195 0 2
rlabel polysilicon 75 -201 75 -201 0 4
rlabel polysilicon 79 -195 79 -195 0 1
rlabel polysilicon 82 -195 82 -195 0 2
rlabel polysilicon 82 -201 82 -201 0 4
rlabel polysilicon 86 -195 86 -195 0 1
rlabel polysilicon 86 -201 86 -201 0 3
rlabel polysilicon 96 -195 96 -195 0 2
rlabel polysilicon 100 -195 100 -195 0 1
rlabel polysilicon 103 -195 103 -195 0 2
rlabel polysilicon 100 -201 100 -201 0 3
rlabel polysilicon 107 -195 107 -195 0 1
rlabel polysilicon 107 -201 107 -201 0 3
rlabel polysilicon 114 -195 114 -195 0 1
rlabel polysilicon 114 -201 114 -201 0 3
rlabel polysilicon 121 -195 121 -195 0 1
rlabel polysilicon 121 -201 121 -201 0 3
rlabel polysilicon 128 -195 128 -195 0 1
rlabel polysilicon 128 -201 128 -201 0 3
rlabel polysilicon 135 -201 135 -201 0 3
rlabel polysilicon 142 -195 142 -195 0 1
rlabel polysilicon 142 -201 142 -201 0 3
rlabel polysilicon 149 -195 149 -195 0 1
rlabel polysilicon 152 -195 152 -195 0 2
rlabel polysilicon 149 -201 149 -201 0 3
rlabel polysilicon 156 -195 156 -195 0 1
rlabel polysilicon 156 -201 156 -201 0 3
rlabel polysilicon 163 -195 163 -195 0 1
rlabel polysilicon 166 -195 166 -195 0 2
rlabel polysilicon 166 -201 166 -201 0 4
rlabel polysilicon 173 -195 173 -195 0 2
rlabel polysilicon 177 -195 177 -195 0 1
rlabel polysilicon 177 -201 177 -201 0 3
rlabel polysilicon 184 -195 184 -195 0 1
rlabel polysilicon 187 -201 187 -201 0 4
rlabel polysilicon 191 -195 191 -195 0 1
rlabel polysilicon 191 -201 191 -201 0 3
rlabel polysilicon 198 -195 198 -195 0 1
rlabel polysilicon 198 -201 198 -201 0 3
rlabel polysilicon 201 -201 201 -201 0 4
rlabel polysilicon 205 -195 205 -195 0 1
rlabel polysilicon 208 -195 208 -195 0 2
rlabel polysilicon 205 -201 205 -201 0 3
rlabel polysilicon 212 -195 212 -195 0 1
rlabel polysilicon 212 -201 212 -201 0 3
rlabel polysilicon 219 -195 219 -195 0 1
rlabel polysilicon 222 -195 222 -195 0 2
rlabel polysilicon 219 -201 219 -201 0 3
rlabel polysilicon 222 -201 222 -201 0 4
rlabel polysilicon 226 -195 226 -195 0 1
rlabel polysilicon 226 -201 226 -201 0 3
rlabel polysilicon 233 -195 233 -195 0 1
rlabel polysilicon 233 -201 233 -201 0 3
rlabel polysilicon 240 -195 240 -195 0 1
rlabel polysilicon 240 -201 240 -201 0 3
rlabel polysilicon 247 -195 247 -195 0 1
rlabel polysilicon 247 -201 247 -201 0 3
rlabel polysilicon 254 -195 254 -195 0 1
rlabel polysilicon 254 -201 254 -201 0 3
rlabel polysilicon 261 -195 261 -195 0 1
rlabel polysilicon 261 -201 261 -201 0 3
rlabel polysilicon 268 -195 268 -195 0 1
rlabel polysilicon 268 -201 268 -201 0 3
rlabel polysilicon 275 -195 275 -195 0 1
rlabel polysilicon 275 -201 275 -201 0 3
rlabel polysilicon 282 -195 282 -195 0 1
rlabel polysilicon 282 -201 282 -201 0 3
rlabel polysilicon 289 -195 289 -195 0 1
rlabel polysilicon 289 -201 289 -201 0 3
rlabel polysilicon 296 -195 296 -195 0 1
rlabel polysilicon 296 -201 296 -201 0 3
rlabel polysilicon 303 -195 303 -195 0 1
rlabel polysilicon 303 -201 303 -201 0 3
rlabel polysilicon 310 -195 310 -195 0 1
rlabel polysilicon 310 -201 310 -201 0 3
rlabel polysilicon 320 -195 320 -195 0 2
rlabel polysilicon 324 -195 324 -195 0 1
rlabel polysilicon 324 -201 324 -201 0 3
rlabel polysilicon 331 -195 331 -195 0 1
rlabel polysilicon 331 -201 331 -201 0 3
rlabel polysilicon 338 -195 338 -195 0 1
rlabel polysilicon 338 -201 338 -201 0 3
rlabel polysilicon 345 -195 345 -195 0 1
rlabel polysilicon 345 -201 345 -201 0 3
rlabel polysilicon 352 -195 352 -195 0 1
rlabel polysilicon 352 -201 352 -201 0 3
rlabel polysilicon 359 -195 359 -195 0 1
rlabel polysilicon 359 -201 359 -201 0 3
rlabel polysilicon 366 -195 366 -195 0 1
rlabel polysilicon 366 -201 366 -201 0 3
rlabel polysilicon 373 -195 373 -195 0 1
rlabel polysilicon 373 -201 373 -201 0 3
rlabel polysilicon 380 -195 380 -195 0 1
rlabel polysilicon 380 -201 380 -201 0 3
rlabel polysilicon 387 -195 387 -195 0 1
rlabel polysilicon 387 -201 387 -201 0 3
rlabel polysilicon 394 -195 394 -195 0 1
rlabel polysilicon 394 -201 394 -201 0 3
rlabel polysilicon 401 -195 401 -195 0 1
rlabel polysilicon 401 -201 401 -201 0 3
rlabel polysilicon 408 -195 408 -195 0 1
rlabel polysilicon 415 -195 415 -195 0 1
rlabel polysilicon 415 -201 415 -201 0 3
rlabel polysilicon 9 -254 9 -254 0 1
rlabel polysilicon 12 -260 12 -260 0 4
rlabel polysilicon 16 -254 16 -254 0 1
rlabel polysilicon 16 -260 16 -260 0 3
rlabel polysilicon 23 -254 23 -254 0 1
rlabel polysilicon 23 -260 23 -260 0 3
rlabel polysilicon 30 -254 30 -254 0 1
rlabel polysilicon 33 -260 33 -260 0 4
rlabel polysilicon 37 -254 37 -254 0 1
rlabel polysilicon 37 -260 37 -260 0 3
rlabel polysilicon 44 -254 44 -254 0 1
rlabel polysilicon 44 -260 44 -260 0 3
rlabel polysilicon 54 -254 54 -254 0 2
rlabel polysilicon 54 -260 54 -260 0 4
rlabel polysilicon 58 -254 58 -254 0 1
rlabel polysilicon 58 -260 58 -260 0 3
rlabel polysilicon 65 -254 65 -254 0 1
rlabel polysilicon 65 -260 65 -260 0 3
rlabel polysilicon 72 -254 72 -254 0 1
rlabel polysilicon 75 -260 75 -260 0 4
rlabel polysilicon 79 -254 79 -254 0 1
rlabel polysilicon 82 -254 82 -254 0 2
rlabel polysilicon 79 -260 79 -260 0 3
rlabel polysilicon 86 -254 86 -254 0 1
rlabel polysilicon 86 -260 86 -260 0 3
rlabel polysilicon 93 -254 93 -254 0 1
rlabel polysilicon 96 -254 96 -254 0 2
rlabel polysilicon 96 -260 96 -260 0 4
rlabel polysilicon 100 -260 100 -260 0 3
rlabel polysilicon 103 -260 103 -260 0 4
rlabel polysilicon 107 -254 107 -254 0 1
rlabel polysilicon 110 -254 110 -254 0 2
rlabel polysilicon 110 -260 110 -260 0 4
rlabel polysilicon 114 -254 114 -254 0 1
rlabel polysilicon 117 -254 117 -254 0 2
rlabel polysilicon 117 -260 117 -260 0 4
rlabel polysilicon 121 -254 121 -254 0 1
rlabel polysilicon 124 -254 124 -254 0 2
rlabel polysilicon 128 -254 128 -254 0 1
rlabel polysilicon 128 -260 128 -260 0 3
rlabel polysilicon 138 -254 138 -254 0 2
rlabel polysilicon 135 -260 135 -260 0 3
rlabel polysilicon 138 -260 138 -260 0 4
rlabel polysilicon 142 -254 142 -254 0 1
rlabel polysilicon 142 -260 142 -260 0 3
rlabel polysilicon 149 -254 149 -254 0 1
rlabel polysilicon 149 -260 149 -260 0 3
rlabel polysilicon 156 -254 156 -254 0 1
rlabel polysilicon 156 -260 156 -260 0 3
rlabel polysilicon 163 -254 163 -254 0 1
rlabel polysilicon 163 -260 163 -260 0 3
rlabel polysilicon 170 -254 170 -254 0 1
rlabel polysilicon 170 -260 170 -260 0 3
rlabel polysilicon 177 -254 177 -254 0 1
rlabel polysilicon 180 -254 180 -254 0 2
rlabel polysilicon 180 -260 180 -260 0 4
rlabel polysilicon 184 -254 184 -254 0 1
rlabel polysilicon 187 -254 187 -254 0 2
rlabel polysilicon 184 -260 184 -260 0 3
rlabel polysilicon 191 -254 191 -254 0 1
rlabel polysilicon 191 -260 191 -260 0 3
rlabel polysilicon 198 -254 198 -254 0 1
rlabel polysilicon 201 -254 201 -254 0 2
rlabel polysilicon 198 -260 198 -260 0 3
rlabel polysilicon 201 -260 201 -260 0 4
rlabel polysilicon 205 -254 205 -254 0 1
rlabel polysilicon 205 -260 205 -260 0 3
rlabel polysilicon 212 -254 212 -254 0 1
rlabel polysilicon 212 -260 212 -260 0 3
rlabel polysilicon 222 -254 222 -254 0 2
rlabel polysilicon 222 -260 222 -260 0 4
rlabel polysilicon 226 -254 226 -254 0 1
rlabel polysilicon 226 -260 226 -260 0 3
rlabel polysilicon 233 -254 233 -254 0 1
rlabel polysilicon 233 -260 233 -260 0 3
rlabel polysilicon 240 -254 240 -254 0 1
rlabel polysilicon 240 -260 240 -260 0 3
rlabel polysilicon 243 -260 243 -260 0 4
rlabel polysilicon 247 -254 247 -254 0 1
rlabel polysilicon 247 -260 247 -260 0 3
rlabel polysilicon 254 -254 254 -254 0 1
rlabel polysilicon 254 -260 254 -260 0 3
rlabel polysilicon 261 -254 261 -254 0 1
rlabel polysilicon 261 -260 261 -260 0 3
rlabel polysilicon 268 -254 268 -254 0 1
rlabel polysilicon 268 -260 268 -260 0 3
rlabel polysilicon 275 -254 275 -254 0 1
rlabel polysilicon 275 -260 275 -260 0 3
rlabel polysilicon 282 -254 282 -254 0 1
rlabel polysilicon 289 -254 289 -254 0 1
rlabel polysilicon 289 -260 289 -260 0 3
rlabel polysilicon 296 -254 296 -254 0 1
rlabel polysilicon 296 -260 296 -260 0 3
rlabel polysilicon 303 -254 303 -254 0 1
rlabel polysilicon 303 -260 303 -260 0 3
rlabel polysilicon 310 -254 310 -254 0 1
rlabel polysilicon 310 -260 310 -260 0 3
rlabel polysilicon 317 -254 317 -254 0 1
rlabel polysilicon 317 -260 317 -260 0 3
rlabel polysilicon 324 -254 324 -254 0 1
rlabel polysilicon 324 -260 324 -260 0 3
rlabel polysilicon 331 -254 331 -254 0 1
rlabel polysilicon 331 -260 331 -260 0 3
rlabel polysilicon 338 -254 338 -254 0 1
rlabel polysilicon 338 -260 338 -260 0 3
rlabel polysilicon 345 -254 345 -254 0 1
rlabel polysilicon 345 -260 345 -260 0 3
rlabel polysilicon 352 -254 352 -254 0 1
rlabel polysilicon 352 -260 352 -260 0 3
rlabel polysilicon 359 -254 359 -254 0 1
rlabel polysilicon 359 -260 359 -260 0 3
rlabel polysilicon 366 -254 366 -254 0 1
rlabel polysilicon 366 -260 366 -260 0 3
rlabel polysilicon 373 -254 373 -254 0 1
rlabel polysilicon 373 -260 373 -260 0 3
rlabel polysilicon 380 -254 380 -254 0 1
rlabel polysilicon 380 -260 380 -260 0 3
rlabel polysilicon 387 -254 387 -254 0 1
rlabel polysilicon 387 -260 387 -260 0 3
rlabel polysilicon 394 -254 394 -254 0 1
rlabel polysilicon 394 -260 394 -260 0 3
rlabel polysilicon 401 -254 401 -254 0 1
rlabel polysilicon 401 -260 401 -260 0 3
rlabel polysilicon 408 -254 408 -254 0 1
rlabel polysilicon 408 -260 408 -260 0 3
rlabel polysilicon 415 -254 415 -254 0 1
rlabel polysilicon 415 -260 415 -260 0 3
rlabel polysilicon 16 -303 16 -303 0 1
rlabel polysilicon 16 -309 16 -309 0 3
rlabel polysilicon 23 -303 23 -303 0 1
rlabel polysilicon 23 -309 23 -309 0 3
rlabel polysilicon 30 -303 30 -303 0 1
rlabel polysilicon 30 -309 30 -309 0 3
rlabel polysilicon 37 -303 37 -303 0 1
rlabel polysilicon 37 -309 37 -309 0 3
rlabel polysilicon 44 -303 44 -303 0 1
rlabel polysilicon 44 -309 44 -309 0 3
rlabel polysilicon 51 -303 51 -303 0 1
rlabel polysilicon 51 -309 51 -309 0 3
rlabel polysilicon 61 -303 61 -303 0 2
rlabel polysilicon 61 -309 61 -309 0 4
rlabel polysilicon 65 -303 65 -303 0 1
rlabel polysilicon 65 -309 65 -309 0 3
rlabel polysilicon 72 -303 72 -303 0 1
rlabel polysilicon 72 -309 72 -309 0 3
rlabel polysilicon 79 -303 79 -303 0 1
rlabel polysilicon 79 -309 79 -309 0 3
rlabel polysilicon 86 -303 86 -303 0 1
rlabel polysilicon 86 -309 86 -309 0 3
rlabel polysilicon 93 -303 93 -303 0 1
rlabel polysilicon 93 -309 93 -309 0 3
rlabel polysilicon 100 -303 100 -303 0 1
rlabel polysilicon 103 -309 103 -309 0 4
rlabel polysilicon 107 -303 107 -303 0 1
rlabel polysilicon 110 -309 110 -309 0 4
rlabel polysilicon 114 -303 114 -303 0 1
rlabel polysilicon 117 -309 117 -309 0 4
rlabel polysilicon 124 -303 124 -303 0 2
rlabel polysilicon 121 -309 121 -309 0 3
rlabel polysilicon 124 -309 124 -309 0 4
rlabel polysilicon 128 -303 128 -303 0 1
rlabel polysilicon 128 -309 128 -309 0 3
rlabel polysilicon 135 -303 135 -303 0 1
rlabel polysilicon 135 -309 135 -309 0 3
rlabel polysilicon 142 -303 142 -303 0 1
rlabel polysilicon 142 -309 142 -309 0 3
rlabel polysilicon 149 -303 149 -303 0 1
rlabel polysilicon 149 -309 149 -309 0 3
rlabel polysilicon 156 -303 156 -303 0 1
rlabel polysilicon 156 -309 156 -309 0 3
rlabel polysilicon 163 -303 163 -303 0 1
rlabel polysilicon 166 -303 166 -303 0 2
rlabel polysilicon 170 -303 170 -303 0 1
rlabel polysilicon 173 -303 173 -303 0 2
rlabel polysilicon 170 -309 170 -309 0 3
rlabel polysilicon 173 -309 173 -309 0 4
rlabel polysilicon 177 -303 177 -303 0 1
rlabel polysilicon 177 -309 177 -309 0 3
rlabel polysilicon 184 -303 184 -303 0 1
rlabel polysilicon 184 -309 184 -309 0 3
rlabel polysilicon 191 -303 191 -303 0 1
rlabel polysilicon 191 -309 191 -309 0 3
rlabel polysilicon 198 -303 198 -303 0 1
rlabel polysilicon 201 -303 201 -303 0 2
rlabel polysilicon 198 -309 198 -309 0 3
rlabel polysilicon 205 -303 205 -303 0 1
rlabel polysilicon 205 -309 205 -309 0 3
rlabel polysilicon 212 -303 212 -303 0 1
rlabel polysilicon 212 -309 212 -309 0 3
rlabel polysilicon 219 -303 219 -303 0 1
rlabel polysilicon 219 -309 219 -309 0 3
rlabel polysilicon 226 -303 226 -303 0 1
rlabel polysilicon 226 -309 226 -309 0 3
rlabel polysilicon 233 -303 233 -303 0 1
rlabel polysilicon 233 -309 233 -309 0 3
rlabel polysilicon 240 -303 240 -303 0 1
rlabel polysilicon 243 -309 243 -309 0 4
rlabel polysilicon 247 -303 247 -303 0 1
rlabel polysilicon 250 -303 250 -303 0 2
rlabel polysilicon 250 -309 250 -309 0 4
rlabel polysilicon 254 -303 254 -303 0 1
rlabel polysilicon 254 -309 254 -309 0 3
rlabel polysilicon 261 -303 261 -303 0 1
rlabel polysilicon 264 -303 264 -303 0 2
rlabel polysilicon 264 -309 264 -309 0 4
rlabel polysilicon 268 -303 268 -303 0 1
rlabel polysilicon 268 -309 268 -309 0 3
rlabel polysilicon 275 -303 275 -303 0 1
rlabel polysilicon 275 -309 275 -309 0 3
rlabel polysilicon 282 -303 282 -303 0 1
rlabel polysilicon 282 -309 282 -309 0 3
rlabel polysilicon 289 -303 289 -303 0 1
rlabel polysilicon 289 -309 289 -309 0 3
rlabel polysilicon 296 -303 296 -303 0 1
rlabel polysilicon 296 -309 296 -309 0 3
rlabel polysilicon 303 -303 303 -303 0 1
rlabel polysilicon 303 -309 303 -309 0 3
rlabel polysilicon 310 -303 310 -303 0 1
rlabel polysilicon 310 -309 310 -309 0 3
rlabel polysilicon 317 -303 317 -303 0 1
rlabel polysilicon 317 -309 317 -309 0 3
rlabel polysilicon 324 -303 324 -303 0 1
rlabel polysilicon 324 -309 324 -309 0 3
rlabel polysilicon 331 -303 331 -303 0 1
rlabel polysilicon 331 -309 331 -309 0 3
rlabel polysilicon 338 -303 338 -303 0 1
rlabel polysilicon 338 -309 338 -309 0 3
rlabel polysilicon 345 -303 345 -303 0 1
rlabel polysilicon 345 -309 345 -309 0 3
rlabel polysilicon 352 -303 352 -303 0 1
rlabel polysilicon 352 -309 352 -309 0 3
rlabel polysilicon 359 -303 359 -303 0 1
rlabel polysilicon 359 -309 359 -309 0 3
rlabel polysilicon 366 -303 366 -303 0 1
rlabel polysilicon 366 -309 366 -309 0 3
rlabel polysilicon 373 -303 373 -303 0 1
rlabel polysilicon 373 -309 373 -309 0 3
rlabel polysilicon 380 -303 380 -303 0 1
rlabel polysilicon 380 -309 380 -309 0 3
rlabel polysilicon 387 -303 387 -303 0 1
rlabel polysilicon 387 -309 387 -309 0 3
rlabel polysilicon 394 -303 394 -303 0 1
rlabel polysilicon 394 -309 394 -309 0 3
rlabel polysilicon 401 -303 401 -303 0 1
rlabel polysilicon 401 -309 401 -309 0 3
rlabel polysilicon 408 -303 408 -303 0 1
rlabel polysilicon 408 -309 408 -309 0 3
rlabel polysilicon 415 -303 415 -303 0 1
rlabel polysilicon 415 -309 415 -309 0 3
rlabel polysilicon 422 -303 422 -303 0 1
rlabel polysilicon 425 -303 425 -303 0 2
rlabel polysilicon 425 -309 425 -309 0 4
rlabel polysilicon 432 -303 432 -303 0 2
rlabel polysilicon 436 -303 436 -303 0 1
rlabel polysilicon 436 -309 436 -309 0 3
rlabel polysilicon 2 -364 2 -364 0 1
rlabel polysilicon 2 -370 2 -370 0 3
rlabel polysilicon 16 -364 16 -364 0 1
rlabel polysilicon 16 -370 16 -370 0 3
rlabel polysilicon 23 -364 23 -364 0 1
rlabel polysilicon 26 -364 26 -364 0 2
rlabel polysilicon 26 -370 26 -370 0 4
rlabel polysilicon 30 -364 30 -364 0 1
rlabel polysilicon 33 -364 33 -364 0 2
rlabel polysilicon 30 -370 30 -370 0 3
rlabel polysilicon 37 -364 37 -364 0 1
rlabel polysilicon 40 -364 40 -364 0 2
rlabel polysilicon 37 -370 37 -370 0 3
rlabel polysilicon 47 -370 47 -370 0 4
rlabel polysilicon 51 -364 51 -364 0 1
rlabel polysilicon 54 -364 54 -364 0 2
rlabel polysilicon 58 -364 58 -364 0 1
rlabel polysilicon 58 -370 58 -370 0 3
rlabel polysilicon 65 -364 65 -364 0 1
rlabel polysilicon 68 -364 68 -364 0 2
rlabel polysilicon 68 -370 68 -370 0 4
rlabel polysilicon 72 -370 72 -370 0 3
rlabel polysilicon 79 -364 79 -364 0 1
rlabel polysilicon 79 -370 79 -370 0 3
rlabel polysilicon 82 -370 82 -370 0 4
rlabel polysilicon 86 -370 86 -370 0 3
rlabel polysilicon 89 -370 89 -370 0 4
rlabel polysilicon 93 -364 93 -364 0 1
rlabel polysilicon 93 -370 93 -370 0 3
rlabel polysilicon 100 -364 100 -364 0 1
rlabel polysilicon 100 -370 100 -370 0 3
rlabel polysilicon 107 -364 107 -364 0 1
rlabel polysilicon 110 -364 110 -364 0 2
rlabel polysilicon 110 -370 110 -370 0 4
rlabel polysilicon 114 -364 114 -364 0 1
rlabel polysilicon 117 -364 117 -364 0 2
rlabel polysilicon 117 -370 117 -370 0 4
rlabel polysilicon 121 -364 121 -364 0 1
rlabel polysilicon 121 -370 121 -370 0 3
rlabel polysilicon 128 -364 128 -364 0 1
rlabel polysilicon 128 -370 128 -370 0 3
rlabel polysilicon 135 -364 135 -364 0 1
rlabel polysilicon 135 -370 135 -370 0 3
rlabel polysilicon 142 -364 142 -364 0 1
rlabel polysilicon 142 -370 142 -370 0 3
rlabel polysilicon 149 -364 149 -364 0 1
rlabel polysilicon 149 -370 149 -370 0 3
rlabel polysilicon 156 -364 156 -364 0 1
rlabel polysilicon 159 -364 159 -364 0 2
rlabel polysilicon 156 -370 156 -370 0 3
rlabel polysilicon 159 -370 159 -370 0 4
rlabel polysilicon 163 -364 163 -364 0 1
rlabel polysilicon 163 -370 163 -370 0 3
rlabel polysilicon 170 -370 170 -370 0 3
rlabel polysilicon 173 -370 173 -370 0 4
rlabel polysilicon 177 -364 177 -364 0 1
rlabel polysilicon 177 -370 177 -370 0 3
rlabel polysilicon 187 -364 187 -364 0 2
rlabel polysilicon 184 -370 184 -370 0 3
rlabel polysilicon 191 -364 191 -364 0 1
rlabel polysilicon 191 -370 191 -370 0 3
rlabel polysilicon 198 -364 198 -364 0 1
rlabel polysilicon 198 -370 198 -370 0 3
rlabel polysilicon 205 -364 205 -364 0 1
rlabel polysilicon 205 -370 205 -370 0 3
rlabel polysilicon 212 -364 212 -364 0 1
rlabel polysilicon 212 -370 212 -370 0 3
rlabel polysilicon 222 -364 222 -364 0 2
rlabel polysilicon 219 -370 219 -370 0 3
rlabel polysilicon 222 -370 222 -370 0 4
rlabel polysilicon 226 -364 226 -364 0 1
rlabel polysilicon 226 -370 226 -370 0 3
rlabel polysilicon 233 -364 233 -364 0 1
rlabel polysilicon 236 -370 236 -370 0 4
rlabel polysilicon 240 -364 240 -364 0 1
rlabel polysilicon 240 -370 240 -370 0 3
rlabel polysilicon 247 -364 247 -364 0 1
rlabel polysilicon 247 -370 247 -370 0 3
rlabel polysilicon 254 -364 254 -364 0 1
rlabel polysilicon 254 -370 254 -370 0 3
rlabel polysilicon 257 -370 257 -370 0 4
rlabel polysilicon 261 -364 261 -364 0 1
rlabel polysilicon 261 -370 261 -370 0 3
rlabel polysilicon 268 -364 268 -364 0 1
rlabel polysilicon 271 -364 271 -364 0 2
rlabel polysilicon 271 -370 271 -370 0 4
rlabel polysilicon 275 -364 275 -364 0 1
rlabel polysilicon 275 -370 275 -370 0 3
rlabel polysilicon 282 -364 282 -364 0 1
rlabel polysilicon 282 -370 282 -370 0 3
rlabel polysilicon 289 -364 289 -364 0 1
rlabel polysilicon 289 -370 289 -370 0 3
rlabel polysilicon 296 -364 296 -364 0 1
rlabel polysilicon 296 -370 296 -370 0 3
rlabel polysilicon 303 -364 303 -364 0 1
rlabel polysilicon 303 -370 303 -370 0 3
rlabel polysilicon 310 -364 310 -364 0 1
rlabel polysilicon 310 -370 310 -370 0 3
rlabel polysilicon 317 -364 317 -364 0 1
rlabel polysilicon 317 -370 317 -370 0 3
rlabel polysilicon 324 -364 324 -364 0 1
rlabel polysilicon 324 -370 324 -370 0 3
rlabel polysilicon 331 -364 331 -364 0 1
rlabel polysilicon 331 -370 331 -370 0 3
rlabel polysilicon 338 -364 338 -364 0 1
rlabel polysilicon 338 -370 338 -370 0 3
rlabel polysilicon 345 -364 345 -364 0 1
rlabel polysilicon 345 -370 345 -370 0 3
rlabel polysilicon 352 -364 352 -364 0 1
rlabel polysilicon 352 -370 352 -370 0 3
rlabel polysilicon 359 -364 359 -364 0 1
rlabel polysilicon 359 -370 359 -370 0 3
rlabel polysilicon 366 -364 366 -364 0 1
rlabel polysilicon 366 -370 366 -370 0 3
rlabel polysilicon 373 -364 373 -364 0 1
rlabel polysilicon 373 -370 373 -370 0 3
rlabel polysilicon 380 -364 380 -364 0 1
rlabel polysilicon 380 -370 380 -370 0 3
rlabel polysilicon 387 -364 387 -364 0 1
rlabel polysilicon 387 -370 387 -370 0 3
rlabel polysilicon 394 -364 394 -364 0 1
rlabel polysilicon 394 -370 394 -370 0 3
rlabel polysilicon 401 -364 401 -364 0 1
rlabel polysilicon 401 -370 401 -370 0 3
rlabel polysilicon 408 -364 408 -364 0 1
rlabel polysilicon 408 -370 408 -370 0 3
rlabel polysilicon 415 -364 415 -364 0 1
rlabel polysilicon 415 -370 415 -370 0 3
rlabel polysilicon 422 -364 422 -364 0 1
rlabel polysilicon 422 -370 422 -370 0 3
rlabel polysilicon 429 -364 429 -364 0 1
rlabel polysilicon 429 -370 429 -370 0 3
rlabel polysilicon 436 -364 436 -364 0 1
rlabel polysilicon 436 -370 436 -370 0 3
rlabel polysilicon 9 -413 9 -413 0 1
rlabel polysilicon 9 -419 9 -419 0 3
rlabel polysilicon 16 -413 16 -413 0 1
rlabel polysilicon 16 -419 16 -419 0 3
rlabel polysilicon 23 -413 23 -413 0 1
rlabel polysilicon 30 -413 30 -413 0 1
rlabel polysilicon 30 -419 30 -419 0 3
rlabel polysilicon 37 -413 37 -413 0 1
rlabel polysilicon 37 -419 37 -419 0 3
rlabel polysilicon 47 -413 47 -413 0 2
rlabel polysilicon 44 -419 44 -419 0 3
rlabel polysilicon 47 -419 47 -419 0 4
rlabel polysilicon 51 -413 51 -413 0 1
rlabel polysilicon 54 -413 54 -413 0 2
rlabel polysilicon 51 -419 51 -419 0 3
rlabel polysilicon 58 -413 58 -413 0 1
rlabel polysilicon 61 -413 61 -413 0 2
rlabel polysilicon 65 -413 65 -413 0 1
rlabel polysilicon 65 -419 65 -419 0 3
rlabel polysilicon 72 -413 72 -413 0 1
rlabel polysilicon 72 -419 72 -419 0 3
rlabel polysilicon 79 -413 79 -413 0 1
rlabel polysilicon 79 -419 79 -419 0 3
rlabel polysilicon 86 -413 86 -413 0 1
rlabel polysilicon 86 -419 86 -419 0 3
rlabel polysilicon 93 -413 93 -413 0 1
rlabel polysilicon 93 -419 93 -419 0 3
rlabel polysilicon 100 -413 100 -413 0 1
rlabel polysilicon 100 -419 100 -419 0 3
rlabel polysilicon 110 -413 110 -413 0 2
rlabel polysilicon 107 -419 107 -419 0 3
rlabel polysilicon 114 -413 114 -413 0 1
rlabel polysilicon 117 -413 117 -413 0 2
rlabel polysilicon 117 -419 117 -419 0 4
rlabel polysilicon 121 -413 121 -413 0 1
rlabel polysilicon 121 -419 121 -419 0 3
rlabel polysilicon 128 -419 128 -419 0 3
rlabel polysilicon 131 -419 131 -419 0 4
rlabel polysilicon 135 -413 135 -413 0 1
rlabel polysilicon 135 -419 135 -419 0 3
rlabel polysilicon 142 -413 142 -413 0 1
rlabel polysilicon 142 -419 142 -419 0 3
rlabel polysilicon 149 -413 149 -413 0 1
rlabel polysilicon 149 -419 149 -419 0 3
rlabel polysilicon 156 -413 156 -413 0 1
rlabel polysilicon 156 -419 156 -419 0 3
rlabel polysilicon 163 -413 163 -413 0 1
rlabel polysilicon 166 -413 166 -413 0 2
rlabel polysilicon 163 -419 163 -419 0 3
rlabel polysilicon 166 -419 166 -419 0 4
rlabel polysilicon 170 -413 170 -413 0 1
rlabel polysilicon 170 -419 170 -419 0 3
rlabel polysilicon 177 -413 177 -413 0 1
rlabel polysilicon 177 -419 177 -419 0 3
rlabel polysilicon 184 -413 184 -413 0 1
rlabel polysilicon 184 -419 184 -419 0 3
rlabel polysilicon 191 -413 191 -413 0 1
rlabel polysilicon 191 -419 191 -419 0 3
rlabel polysilicon 201 -413 201 -413 0 2
rlabel polysilicon 205 -413 205 -413 0 1
rlabel polysilicon 205 -419 205 -419 0 3
rlabel polysilicon 212 -413 212 -413 0 1
rlabel polysilicon 212 -419 212 -419 0 3
rlabel polysilicon 219 -413 219 -413 0 1
rlabel polysilicon 219 -419 219 -419 0 3
rlabel polysilicon 229 -413 229 -413 0 2
rlabel polysilicon 226 -419 226 -419 0 3
rlabel polysilicon 233 -413 233 -413 0 1
rlabel polysilicon 233 -419 233 -419 0 3
rlabel polysilicon 240 -413 240 -413 0 1
rlabel polysilicon 240 -419 240 -419 0 3
rlabel polysilicon 250 -413 250 -413 0 2
rlabel polysilicon 247 -419 247 -419 0 3
rlabel polysilicon 250 -419 250 -419 0 4
rlabel polysilicon 254 -413 254 -413 0 1
rlabel polysilicon 254 -419 254 -419 0 3
rlabel polysilicon 261 -413 261 -413 0 1
rlabel polysilicon 264 -413 264 -413 0 2
rlabel polysilicon 261 -419 261 -419 0 3
rlabel polysilicon 268 -413 268 -413 0 1
rlabel polysilicon 271 -413 271 -413 0 2
rlabel polysilicon 268 -419 268 -419 0 3
rlabel polysilicon 275 -413 275 -413 0 1
rlabel polysilicon 275 -419 275 -419 0 3
rlabel polysilicon 282 -413 282 -413 0 1
rlabel polysilicon 282 -419 282 -419 0 3
rlabel polysilicon 289 -413 289 -413 0 1
rlabel polysilicon 289 -419 289 -419 0 3
rlabel polysilicon 296 -413 296 -413 0 1
rlabel polysilicon 296 -419 296 -419 0 3
rlabel polysilicon 303 -413 303 -413 0 1
rlabel polysilicon 303 -419 303 -419 0 3
rlabel polysilicon 310 -413 310 -413 0 1
rlabel polysilicon 310 -419 310 -419 0 3
rlabel polysilicon 317 -413 317 -413 0 1
rlabel polysilicon 317 -419 317 -419 0 3
rlabel polysilicon 327 -413 327 -413 0 2
rlabel polysilicon 324 -419 324 -419 0 3
rlabel polysilicon 327 -419 327 -419 0 4
rlabel polysilicon 334 -419 334 -419 0 4
rlabel polysilicon 338 -413 338 -413 0 1
rlabel polysilicon 338 -419 338 -419 0 3
rlabel polysilicon 345 -413 345 -413 0 1
rlabel polysilicon 345 -419 345 -419 0 3
rlabel polysilicon 352 -413 352 -413 0 1
rlabel polysilicon 352 -419 352 -419 0 3
rlabel polysilicon 359 -413 359 -413 0 1
rlabel polysilicon 359 -419 359 -419 0 3
rlabel polysilicon 366 -413 366 -413 0 1
rlabel polysilicon 366 -419 366 -419 0 3
rlabel polysilicon 373 -413 373 -413 0 1
rlabel polysilicon 373 -419 373 -419 0 3
rlabel polysilicon 380 -413 380 -413 0 1
rlabel polysilicon 380 -419 380 -419 0 3
rlabel polysilicon 387 -413 387 -413 0 1
rlabel polysilicon 387 -419 387 -419 0 3
rlabel polysilicon 394 -413 394 -413 0 1
rlabel polysilicon 394 -419 394 -419 0 3
rlabel polysilicon 401 -413 401 -413 0 1
rlabel polysilicon 401 -419 401 -419 0 3
rlabel polysilicon 408 -413 408 -413 0 1
rlabel polysilicon 408 -419 408 -419 0 3
rlabel polysilicon 415 -413 415 -413 0 1
rlabel polysilicon 415 -419 415 -419 0 3
rlabel polysilicon 422 -413 422 -413 0 1
rlabel polysilicon 422 -419 422 -419 0 3
rlabel polysilicon 429 -413 429 -413 0 1
rlabel polysilicon 432 -413 432 -413 0 2
rlabel polysilicon 432 -419 432 -419 0 4
rlabel polysilicon 436 -413 436 -413 0 1
rlabel polysilicon 436 -419 436 -419 0 3
rlabel polysilicon 443 -419 443 -419 0 3
rlabel polysilicon 16 -468 16 -468 0 1
rlabel polysilicon 16 -474 16 -474 0 3
rlabel polysilicon 26 -468 26 -468 0 2
rlabel polysilicon 33 -468 33 -468 0 2
rlabel polysilicon 37 -468 37 -468 0 1
rlabel polysilicon 37 -474 37 -474 0 3
rlabel polysilicon 51 -468 51 -468 0 1
rlabel polysilicon 51 -474 51 -474 0 3
rlabel polysilicon 58 -468 58 -468 0 1
rlabel polysilicon 58 -474 58 -474 0 3
rlabel polysilicon 65 -468 65 -468 0 1
rlabel polysilicon 65 -474 65 -474 0 3
rlabel polysilicon 72 -468 72 -468 0 1
rlabel polysilicon 75 -468 75 -468 0 2
rlabel polysilicon 72 -474 72 -474 0 3
rlabel polysilicon 79 -468 79 -468 0 1
rlabel polysilicon 79 -474 79 -474 0 3
rlabel polysilicon 86 -468 86 -468 0 1
rlabel polysilicon 86 -474 86 -474 0 3
rlabel polysilicon 93 -468 93 -468 0 1
rlabel polysilicon 93 -474 93 -474 0 3
rlabel polysilicon 100 -468 100 -468 0 1
rlabel polysilicon 100 -474 100 -474 0 3
rlabel polysilicon 107 -468 107 -468 0 1
rlabel polysilicon 107 -474 107 -474 0 3
rlabel polysilicon 110 -474 110 -474 0 4
rlabel polysilicon 114 -468 114 -468 0 1
rlabel polysilicon 114 -474 114 -474 0 3
rlabel polysilicon 121 -468 121 -468 0 1
rlabel polysilicon 121 -474 121 -474 0 3
rlabel polysilicon 128 -468 128 -468 0 1
rlabel polysilicon 128 -474 128 -474 0 3
rlabel polysilicon 131 -474 131 -474 0 4
rlabel polysilicon 135 -468 135 -468 0 1
rlabel polysilicon 135 -474 135 -474 0 3
rlabel polysilicon 142 -468 142 -468 0 1
rlabel polysilicon 142 -474 142 -474 0 3
rlabel polysilicon 149 -468 149 -468 0 1
rlabel polysilicon 149 -474 149 -474 0 3
rlabel polysilicon 156 -468 156 -468 0 1
rlabel polysilicon 156 -474 156 -474 0 3
rlabel polysilicon 163 -468 163 -468 0 1
rlabel polysilicon 163 -474 163 -474 0 3
rlabel polysilicon 170 -468 170 -468 0 1
rlabel polysilicon 170 -474 170 -474 0 3
rlabel polysilicon 177 -468 177 -468 0 1
rlabel polysilicon 180 -468 180 -468 0 2
rlabel polysilicon 180 -474 180 -474 0 4
rlabel polysilicon 184 -468 184 -468 0 1
rlabel polysilicon 184 -474 184 -474 0 3
rlabel polysilicon 191 -468 191 -468 0 1
rlabel polysilicon 194 -468 194 -468 0 2
rlabel polysilicon 191 -474 191 -474 0 3
rlabel polysilicon 194 -474 194 -474 0 4
rlabel polysilicon 198 -468 198 -468 0 1
rlabel polysilicon 201 -468 201 -468 0 2
rlabel polysilicon 205 -468 205 -468 0 1
rlabel polysilicon 205 -474 205 -474 0 3
rlabel polysilicon 212 -468 212 -468 0 1
rlabel polysilicon 215 -468 215 -468 0 2
rlabel polysilicon 212 -474 212 -474 0 3
rlabel polysilicon 222 -468 222 -468 0 2
rlabel polysilicon 222 -474 222 -474 0 4
rlabel polysilicon 226 -468 226 -468 0 1
rlabel polysilicon 229 -468 229 -468 0 2
rlabel polysilicon 236 -468 236 -468 0 2
rlabel polysilicon 236 -474 236 -474 0 4
rlabel polysilicon 243 -468 243 -468 0 2
rlabel polysilicon 250 -468 250 -468 0 2
rlabel polysilicon 247 -474 247 -474 0 3
rlabel polysilicon 250 -474 250 -474 0 4
rlabel polysilicon 254 -468 254 -468 0 1
rlabel polysilicon 257 -468 257 -468 0 2
rlabel polysilicon 261 -468 261 -468 0 1
rlabel polysilicon 261 -474 261 -474 0 3
rlabel polysilicon 264 -474 264 -474 0 4
rlabel polysilicon 268 -468 268 -468 0 1
rlabel polysilicon 268 -474 268 -474 0 3
rlabel polysilicon 275 -468 275 -468 0 1
rlabel polysilicon 275 -474 275 -474 0 3
rlabel polysilicon 282 -468 282 -468 0 1
rlabel polysilicon 282 -474 282 -474 0 3
rlabel polysilicon 285 -474 285 -474 0 4
rlabel polysilicon 289 -468 289 -468 0 1
rlabel polysilicon 289 -474 289 -474 0 3
rlabel polysilicon 296 -468 296 -468 0 1
rlabel polysilicon 296 -474 296 -474 0 3
rlabel polysilicon 303 -468 303 -468 0 1
rlabel polysilicon 303 -474 303 -474 0 3
rlabel polysilicon 310 -468 310 -468 0 1
rlabel polysilicon 310 -474 310 -474 0 3
rlabel polysilicon 317 -468 317 -468 0 1
rlabel polysilicon 317 -474 317 -474 0 3
rlabel polysilicon 324 -468 324 -468 0 1
rlabel polysilicon 324 -474 324 -474 0 3
rlabel polysilicon 331 -468 331 -468 0 1
rlabel polysilicon 331 -474 331 -474 0 3
rlabel polysilicon 338 -468 338 -468 0 1
rlabel polysilicon 338 -474 338 -474 0 3
rlabel polysilicon 345 -468 345 -468 0 1
rlabel polysilicon 345 -474 345 -474 0 3
rlabel polysilicon 352 -468 352 -468 0 1
rlabel polysilicon 352 -474 352 -474 0 3
rlabel polysilicon 359 -468 359 -468 0 1
rlabel polysilicon 359 -474 359 -474 0 3
rlabel polysilicon 366 -468 366 -468 0 1
rlabel polysilicon 366 -474 366 -474 0 3
rlabel polysilicon 373 -468 373 -468 0 1
rlabel polysilicon 373 -474 373 -474 0 3
rlabel polysilicon 380 -468 380 -468 0 1
rlabel polysilicon 380 -474 380 -474 0 3
rlabel polysilicon 387 -468 387 -468 0 1
rlabel polysilicon 387 -474 387 -474 0 3
rlabel polysilicon 394 -468 394 -468 0 1
rlabel polysilicon 394 -474 394 -474 0 3
rlabel polysilicon 415 -468 415 -468 0 1
rlabel polysilicon 415 -474 415 -474 0 3
rlabel polysilicon 422 -468 422 -468 0 1
rlabel polysilicon 422 -474 422 -474 0 3
rlabel polysilicon 432 -468 432 -468 0 2
rlabel polysilicon 429 -474 429 -474 0 3
rlabel polysilicon 436 -468 436 -468 0 1
rlabel polysilicon 436 -474 436 -474 0 3
rlabel polysilicon 446 -468 446 -468 0 2
rlabel polysilicon 446 -474 446 -474 0 4
rlabel polysilicon 450 -468 450 -468 0 1
rlabel polysilicon 450 -474 450 -474 0 3
rlabel polysilicon 457 -468 457 -468 0 1
rlabel polysilicon 457 -474 457 -474 0 3
rlabel polysilicon 464 -468 464 -468 0 1
rlabel polysilicon 464 -474 464 -474 0 3
rlabel polysilicon 9 -509 9 -509 0 1
rlabel polysilicon 9 -515 9 -515 0 3
rlabel polysilicon 16 -509 16 -509 0 1
rlabel polysilicon 16 -515 16 -515 0 3
rlabel polysilicon 23 -509 23 -509 0 1
rlabel polysilicon 30 -509 30 -509 0 1
rlabel polysilicon 33 -509 33 -509 0 2
rlabel polysilicon 30 -515 30 -515 0 3
rlabel polysilicon 37 -509 37 -509 0 1
rlabel polysilicon 40 -509 40 -509 0 2
rlabel polysilicon 37 -515 37 -515 0 3
rlabel polysilicon 40 -515 40 -515 0 4
rlabel polysilicon 44 -509 44 -509 0 1
rlabel polysilicon 44 -515 44 -515 0 3
rlabel polysilicon 51 -509 51 -509 0 1
rlabel polysilicon 51 -515 51 -515 0 3
rlabel polysilicon 58 -509 58 -509 0 1
rlabel polysilicon 58 -515 58 -515 0 3
rlabel polysilicon 65 -509 65 -509 0 1
rlabel polysilicon 65 -515 65 -515 0 3
rlabel polysilicon 72 -509 72 -509 0 1
rlabel polysilicon 72 -515 72 -515 0 3
rlabel polysilicon 79 -509 79 -509 0 1
rlabel polysilicon 82 -509 82 -509 0 2
rlabel polysilicon 82 -515 82 -515 0 4
rlabel polysilicon 86 -509 86 -509 0 1
rlabel polysilicon 86 -515 86 -515 0 3
rlabel polysilicon 93 -509 93 -509 0 1
rlabel polysilicon 93 -515 93 -515 0 3
rlabel polysilicon 103 -509 103 -509 0 2
rlabel polysilicon 103 -515 103 -515 0 4
rlabel polysilicon 107 -509 107 -509 0 1
rlabel polysilicon 107 -515 107 -515 0 3
rlabel polysilicon 114 -509 114 -509 0 1
rlabel polysilicon 114 -515 114 -515 0 3
rlabel polysilicon 121 -509 121 -509 0 1
rlabel polysilicon 124 -509 124 -509 0 2
rlabel polysilicon 121 -515 121 -515 0 3
rlabel polysilicon 124 -515 124 -515 0 4
rlabel polysilicon 128 -509 128 -509 0 1
rlabel polysilicon 128 -515 128 -515 0 3
rlabel polysilicon 138 -509 138 -509 0 2
rlabel polysilicon 138 -515 138 -515 0 4
rlabel polysilicon 142 -509 142 -509 0 1
rlabel polysilicon 142 -515 142 -515 0 3
rlabel polysilicon 149 -509 149 -509 0 1
rlabel polysilicon 149 -515 149 -515 0 3
rlabel polysilicon 156 -509 156 -509 0 1
rlabel polysilicon 156 -515 156 -515 0 3
rlabel polysilicon 163 -509 163 -509 0 1
rlabel polysilicon 163 -515 163 -515 0 3
rlabel polysilicon 173 -509 173 -509 0 2
rlabel polysilicon 173 -515 173 -515 0 4
rlabel polysilicon 177 -509 177 -509 0 1
rlabel polysilicon 177 -515 177 -515 0 3
rlabel polysilicon 184 -509 184 -509 0 1
rlabel polysilicon 184 -515 184 -515 0 3
rlabel polysilicon 191 -509 191 -509 0 1
rlabel polysilicon 191 -515 191 -515 0 3
rlabel polysilicon 198 -509 198 -509 0 1
rlabel polysilicon 198 -515 198 -515 0 3
rlabel polysilicon 205 -509 205 -509 0 1
rlabel polysilicon 205 -515 205 -515 0 3
rlabel polysilicon 208 -515 208 -515 0 4
rlabel polysilicon 215 -509 215 -509 0 2
rlabel polysilicon 212 -515 212 -515 0 3
rlabel polysilicon 215 -515 215 -515 0 4
rlabel polysilicon 219 -509 219 -509 0 1
rlabel polysilicon 219 -515 219 -515 0 3
rlabel polysilicon 226 -509 226 -509 0 1
rlabel polysilicon 226 -515 226 -515 0 3
rlabel polysilicon 233 -509 233 -509 0 1
rlabel polysilicon 233 -515 233 -515 0 3
rlabel polysilicon 240 -509 240 -509 0 1
rlabel polysilicon 243 -509 243 -509 0 2
rlabel polysilicon 243 -515 243 -515 0 4
rlabel polysilicon 247 -509 247 -509 0 1
rlabel polysilicon 247 -515 247 -515 0 3
rlabel polysilicon 254 -509 254 -509 0 1
rlabel polysilicon 254 -515 254 -515 0 3
rlabel polysilicon 261 -509 261 -509 0 1
rlabel polysilicon 261 -515 261 -515 0 3
rlabel polysilicon 268 -509 268 -509 0 1
rlabel polysilicon 268 -515 268 -515 0 3
rlabel polysilicon 275 -515 275 -515 0 3
rlabel polysilicon 278 -515 278 -515 0 4
rlabel polysilicon 282 -515 282 -515 0 3
rlabel polysilicon 289 -509 289 -509 0 1
rlabel polysilicon 289 -515 289 -515 0 3
rlabel polysilicon 296 -509 296 -509 0 1
rlabel polysilicon 296 -515 296 -515 0 3
rlabel polysilicon 303 -509 303 -509 0 1
rlabel polysilicon 303 -515 303 -515 0 3
rlabel polysilicon 306 -515 306 -515 0 4
rlabel polysilicon 310 -509 310 -509 0 1
rlabel polysilicon 310 -515 310 -515 0 3
rlabel polysilicon 317 -509 317 -509 0 1
rlabel polysilicon 317 -515 317 -515 0 3
rlabel polysilicon 324 -509 324 -509 0 1
rlabel polysilicon 324 -515 324 -515 0 3
rlabel polysilicon 331 -509 331 -509 0 1
rlabel polysilicon 331 -515 331 -515 0 3
rlabel polysilicon 338 -509 338 -509 0 1
rlabel polysilicon 338 -515 338 -515 0 3
rlabel polysilicon 345 -509 345 -509 0 1
rlabel polysilicon 345 -515 345 -515 0 3
rlabel polysilicon 352 -509 352 -509 0 1
rlabel polysilicon 352 -515 352 -515 0 3
rlabel polysilicon 359 -509 359 -509 0 1
rlabel polysilicon 359 -515 359 -515 0 3
rlabel polysilicon 366 -515 366 -515 0 3
rlabel polysilicon 373 -509 373 -509 0 1
rlabel polysilicon 373 -515 373 -515 0 3
rlabel polysilicon 380 -509 380 -509 0 1
rlabel polysilicon 380 -515 380 -515 0 3
rlabel polysilicon 387 -509 387 -509 0 1
rlabel polysilicon 387 -515 387 -515 0 3
rlabel polysilicon 401 -509 401 -509 0 1
rlabel polysilicon 401 -515 401 -515 0 3
rlabel polysilicon 408 -509 408 -509 0 1
rlabel polysilicon 408 -515 408 -515 0 3
rlabel polysilicon 415 -509 415 -509 0 1
rlabel polysilicon 418 -509 418 -509 0 2
rlabel polysilicon 415 -515 415 -515 0 3
rlabel polysilicon 429 -509 429 -509 0 1
rlabel polysilicon 432 -509 432 -509 0 2
rlabel polysilicon 432 -515 432 -515 0 4
rlabel polysilicon 436 -509 436 -509 0 1
rlabel polysilicon 436 -515 436 -515 0 3
rlabel polysilicon 443 -509 443 -509 0 1
rlabel polysilicon 443 -515 443 -515 0 3
rlabel polysilicon 450 -509 450 -509 0 1
rlabel polysilicon 450 -515 450 -515 0 3
rlabel polysilicon 457 -509 457 -509 0 1
rlabel polysilicon 457 -515 457 -515 0 3
rlabel polysilicon 464 -509 464 -509 0 1
rlabel polysilicon 464 -515 464 -515 0 3
rlabel polysilicon 9 -562 9 -562 0 1
rlabel polysilicon 9 -568 9 -568 0 3
rlabel polysilicon 19 -562 19 -562 0 2
rlabel polysilicon 16 -568 16 -568 0 3
rlabel polysilicon 23 -562 23 -562 0 1
rlabel polysilicon 26 -562 26 -562 0 2
rlabel polysilicon 30 -562 30 -562 0 1
rlabel polysilicon 30 -568 30 -568 0 3
rlabel polysilicon 37 -562 37 -562 0 1
rlabel polysilicon 37 -568 37 -568 0 3
rlabel polysilicon 44 -562 44 -562 0 1
rlabel polysilicon 44 -568 44 -568 0 3
rlabel polysilicon 51 -562 51 -562 0 1
rlabel polysilicon 51 -568 51 -568 0 3
rlabel polysilicon 58 -562 58 -562 0 1
rlabel polysilicon 58 -568 58 -568 0 3
rlabel polysilicon 65 -562 65 -562 0 1
rlabel polysilicon 68 -562 68 -562 0 2
rlabel polysilicon 68 -568 68 -568 0 4
rlabel polysilicon 72 -562 72 -562 0 1
rlabel polysilicon 72 -568 72 -568 0 3
rlabel polysilicon 82 -562 82 -562 0 2
rlabel polysilicon 79 -568 79 -568 0 3
rlabel polysilicon 86 -562 86 -562 0 1
rlabel polysilicon 86 -568 86 -568 0 3
rlabel polysilicon 93 -562 93 -562 0 1
rlabel polysilicon 96 -562 96 -562 0 2
rlabel polysilicon 93 -568 93 -568 0 3
rlabel polysilicon 103 -562 103 -562 0 2
rlabel polysilicon 103 -568 103 -568 0 4
rlabel polysilicon 107 -562 107 -562 0 1
rlabel polysilicon 107 -568 107 -568 0 3
rlabel polysilicon 114 -562 114 -562 0 1
rlabel polysilicon 117 -562 117 -562 0 2
rlabel polysilicon 124 -562 124 -562 0 2
rlabel polysilicon 121 -568 121 -568 0 3
rlabel polysilicon 128 -562 128 -562 0 1
rlabel polysilicon 128 -568 128 -568 0 3
rlabel polysilicon 135 -562 135 -562 0 1
rlabel polysilicon 135 -568 135 -568 0 3
rlabel polysilicon 142 -562 142 -562 0 1
rlabel polysilicon 142 -568 142 -568 0 3
rlabel polysilicon 149 -562 149 -562 0 1
rlabel polysilicon 149 -568 149 -568 0 3
rlabel polysilicon 156 -562 156 -562 0 1
rlabel polysilicon 156 -568 156 -568 0 3
rlabel polysilicon 163 -562 163 -562 0 1
rlabel polysilicon 166 -562 166 -562 0 2
rlabel polysilicon 163 -568 163 -568 0 3
rlabel polysilicon 170 -562 170 -562 0 1
rlabel polysilicon 173 -562 173 -562 0 2
rlabel polysilicon 170 -568 170 -568 0 3
rlabel polysilicon 173 -568 173 -568 0 4
rlabel polysilicon 177 -562 177 -562 0 1
rlabel polysilicon 180 -568 180 -568 0 4
rlabel polysilicon 184 -562 184 -562 0 1
rlabel polysilicon 187 -562 187 -562 0 2
rlabel polysilicon 191 -562 191 -562 0 1
rlabel polysilicon 191 -568 191 -568 0 3
rlabel polysilicon 198 -562 198 -562 0 1
rlabel polysilicon 198 -568 198 -568 0 3
rlabel polysilicon 205 -562 205 -562 0 1
rlabel polysilicon 205 -568 205 -568 0 3
rlabel polysilicon 208 -568 208 -568 0 4
rlabel polysilicon 212 -562 212 -562 0 1
rlabel polysilicon 212 -568 212 -568 0 3
rlabel polysilicon 219 -562 219 -562 0 1
rlabel polysilicon 219 -568 219 -568 0 3
rlabel polysilicon 226 -562 226 -562 0 1
rlabel polysilicon 226 -568 226 -568 0 3
rlabel polysilicon 233 -562 233 -562 0 1
rlabel polysilicon 236 -562 236 -562 0 2
rlabel polysilicon 233 -568 233 -568 0 3
rlabel polysilicon 236 -568 236 -568 0 4
rlabel polysilicon 240 -562 240 -562 0 1
rlabel polysilicon 240 -568 240 -568 0 3
rlabel polysilicon 243 -568 243 -568 0 4
rlabel polysilicon 247 -562 247 -562 0 1
rlabel polysilicon 247 -568 247 -568 0 3
rlabel polysilicon 254 -562 254 -562 0 1
rlabel polysilicon 254 -568 254 -568 0 3
rlabel polysilicon 261 -562 261 -562 0 1
rlabel polysilicon 261 -568 261 -568 0 3
rlabel polysilicon 268 -562 268 -562 0 1
rlabel polysilicon 268 -568 268 -568 0 3
rlabel polysilicon 275 -562 275 -562 0 1
rlabel polysilicon 275 -568 275 -568 0 3
rlabel polysilicon 282 -562 282 -562 0 1
rlabel polysilicon 285 -562 285 -562 0 2
rlabel polysilicon 282 -568 282 -568 0 3
rlabel polysilicon 289 -562 289 -562 0 1
rlabel polysilicon 289 -568 289 -568 0 3
rlabel polysilicon 296 -562 296 -562 0 1
rlabel polysilicon 296 -568 296 -568 0 3
rlabel polysilicon 303 -568 303 -568 0 3
rlabel polysilicon 306 -568 306 -568 0 4
rlabel polysilicon 310 -562 310 -562 0 1
rlabel polysilicon 310 -568 310 -568 0 3
rlabel polysilicon 317 -562 317 -562 0 1
rlabel polysilicon 317 -568 317 -568 0 3
rlabel polysilicon 324 -562 324 -562 0 1
rlabel polysilicon 324 -568 324 -568 0 3
rlabel polysilicon 331 -562 331 -562 0 1
rlabel polysilicon 331 -568 331 -568 0 3
rlabel polysilicon 341 -562 341 -562 0 2
rlabel polysilicon 338 -568 338 -568 0 3
rlabel polysilicon 341 -568 341 -568 0 4
rlabel polysilicon 345 -562 345 -562 0 1
rlabel polysilicon 345 -568 345 -568 0 3
rlabel polysilicon 352 -562 352 -562 0 1
rlabel polysilicon 352 -568 352 -568 0 3
rlabel polysilicon 359 -562 359 -562 0 1
rlabel polysilicon 359 -568 359 -568 0 3
rlabel polysilicon 366 -562 366 -562 0 1
rlabel polysilicon 366 -568 366 -568 0 3
rlabel polysilicon 373 -562 373 -562 0 1
rlabel polysilicon 373 -568 373 -568 0 3
rlabel polysilicon 380 -562 380 -562 0 1
rlabel polysilicon 380 -568 380 -568 0 3
rlabel polysilicon 387 -562 387 -562 0 1
rlabel polysilicon 387 -568 387 -568 0 3
rlabel polysilicon 394 -562 394 -562 0 1
rlabel polysilicon 394 -568 394 -568 0 3
rlabel polysilicon 401 -562 401 -562 0 1
rlabel polysilicon 401 -568 401 -568 0 3
rlabel polysilicon 408 -562 408 -562 0 1
rlabel polysilicon 408 -568 408 -568 0 3
rlabel polysilicon 415 -562 415 -562 0 1
rlabel polysilicon 415 -568 415 -568 0 3
rlabel polysilicon 422 -562 422 -562 0 1
rlabel polysilicon 422 -568 422 -568 0 3
rlabel polysilicon 429 -562 429 -562 0 1
rlabel polysilicon 429 -568 429 -568 0 3
rlabel polysilicon 436 -562 436 -562 0 1
rlabel polysilicon 436 -568 436 -568 0 3
rlabel polysilicon 443 -562 443 -562 0 1
rlabel polysilicon 443 -568 443 -568 0 3
rlabel polysilicon 457 -562 457 -562 0 1
rlabel polysilicon 464 -562 464 -562 0 1
rlabel polysilicon 464 -568 464 -568 0 3
rlabel polysilicon 9 -615 9 -615 0 1
rlabel polysilicon 9 -621 9 -621 0 3
rlabel polysilicon 16 -615 16 -615 0 1
rlabel polysilicon 16 -621 16 -621 0 3
rlabel polysilicon 23 -615 23 -615 0 1
rlabel polysilicon 23 -621 23 -621 0 3
rlabel polysilicon 30 -615 30 -615 0 1
rlabel polysilicon 33 -615 33 -615 0 2
rlabel polysilicon 33 -621 33 -621 0 4
rlabel polysilicon 40 -615 40 -615 0 2
rlabel polysilicon 37 -621 37 -621 0 3
rlabel polysilicon 40 -621 40 -621 0 4
rlabel polysilicon 44 -615 44 -615 0 1
rlabel polysilicon 44 -621 44 -621 0 3
rlabel polysilicon 51 -615 51 -615 0 1
rlabel polysilicon 51 -621 51 -621 0 3
rlabel polysilicon 58 -615 58 -615 0 1
rlabel polysilicon 58 -621 58 -621 0 3
rlabel polysilicon 65 -615 65 -615 0 1
rlabel polysilicon 65 -621 65 -621 0 3
rlabel polysilicon 72 -615 72 -615 0 1
rlabel polysilicon 72 -621 72 -621 0 3
rlabel polysilicon 79 -615 79 -615 0 1
rlabel polysilicon 79 -621 79 -621 0 3
rlabel polysilicon 86 -615 86 -615 0 1
rlabel polysilicon 89 -615 89 -615 0 2
rlabel polysilicon 89 -621 89 -621 0 4
rlabel polysilicon 93 -615 93 -615 0 1
rlabel polysilicon 93 -621 93 -621 0 3
rlabel polysilicon 100 -615 100 -615 0 1
rlabel polysilicon 100 -621 100 -621 0 3
rlabel polysilicon 103 -621 103 -621 0 4
rlabel polysilicon 107 -615 107 -615 0 1
rlabel polysilicon 107 -621 107 -621 0 3
rlabel polysilicon 114 -615 114 -615 0 1
rlabel polysilicon 114 -621 114 -621 0 3
rlabel polysilicon 117 -621 117 -621 0 4
rlabel polysilicon 121 -615 121 -615 0 1
rlabel polysilicon 121 -621 121 -621 0 3
rlabel polysilicon 128 -621 128 -621 0 3
rlabel polysilicon 131 -621 131 -621 0 4
rlabel polysilicon 138 -615 138 -615 0 2
rlabel polysilicon 135 -621 135 -621 0 3
rlabel polysilicon 142 -615 142 -615 0 1
rlabel polysilicon 142 -621 142 -621 0 3
rlabel polysilicon 149 -615 149 -615 0 1
rlabel polysilicon 149 -621 149 -621 0 3
rlabel polysilicon 156 -615 156 -615 0 1
rlabel polysilicon 156 -621 156 -621 0 3
rlabel polysilicon 163 -615 163 -615 0 1
rlabel polysilicon 163 -621 163 -621 0 3
rlabel polysilicon 170 -615 170 -615 0 1
rlabel polysilicon 173 -615 173 -615 0 2
rlabel polysilicon 170 -621 170 -621 0 3
rlabel polysilicon 177 -615 177 -615 0 1
rlabel polysilicon 177 -621 177 -621 0 3
rlabel polysilicon 184 -615 184 -615 0 1
rlabel polysilicon 184 -621 184 -621 0 3
rlabel polysilicon 194 -615 194 -615 0 2
rlabel polysilicon 191 -621 191 -621 0 3
rlabel polysilicon 194 -621 194 -621 0 4
rlabel polysilicon 198 -615 198 -615 0 1
rlabel polysilicon 198 -621 198 -621 0 3
rlabel polysilicon 208 -615 208 -615 0 2
rlabel polysilicon 208 -621 208 -621 0 4
rlabel polysilicon 212 -621 212 -621 0 3
rlabel polysilicon 215 -621 215 -621 0 4
rlabel polysilicon 219 -615 219 -615 0 1
rlabel polysilicon 219 -621 219 -621 0 3
rlabel polysilicon 226 -615 226 -615 0 1
rlabel polysilicon 226 -621 226 -621 0 3
rlabel polysilicon 233 -615 233 -615 0 1
rlabel polysilicon 233 -621 233 -621 0 3
rlabel polysilicon 240 -615 240 -615 0 1
rlabel polysilicon 240 -621 240 -621 0 3
rlabel polysilicon 247 -615 247 -615 0 1
rlabel polysilicon 250 -621 250 -621 0 4
rlabel polysilicon 257 -615 257 -615 0 2
rlabel polysilicon 254 -621 254 -621 0 3
rlabel polysilicon 264 -615 264 -615 0 2
rlabel polysilicon 261 -621 261 -621 0 3
rlabel polysilicon 268 -615 268 -615 0 1
rlabel polysilicon 268 -621 268 -621 0 3
rlabel polysilicon 275 -615 275 -615 0 1
rlabel polysilicon 275 -621 275 -621 0 3
rlabel polysilicon 282 -615 282 -615 0 1
rlabel polysilicon 282 -621 282 -621 0 3
rlabel polysilicon 289 -615 289 -615 0 1
rlabel polysilicon 289 -621 289 -621 0 3
rlabel polysilicon 296 -615 296 -615 0 1
rlabel polysilicon 299 -621 299 -621 0 4
rlabel polysilicon 303 -615 303 -615 0 1
rlabel polysilicon 303 -621 303 -621 0 3
rlabel polysilicon 310 -615 310 -615 0 1
rlabel polysilicon 310 -621 310 -621 0 3
rlabel polysilicon 317 -615 317 -615 0 1
rlabel polysilicon 317 -621 317 -621 0 3
rlabel polysilicon 324 -615 324 -615 0 1
rlabel polysilicon 324 -621 324 -621 0 3
rlabel polysilicon 331 -615 331 -615 0 1
rlabel polysilicon 331 -621 331 -621 0 3
rlabel polysilicon 334 -621 334 -621 0 4
rlabel polysilicon 338 -615 338 -615 0 1
rlabel polysilicon 338 -621 338 -621 0 3
rlabel polysilicon 345 -615 345 -615 0 1
rlabel polysilicon 345 -621 345 -621 0 3
rlabel polysilicon 352 -615 352 -615 0 1
rlabel polysilicon 352 -621 352 -621 0 3
rlabel polysilicon 359 -615 359 -615 0 1
rlabel polysilicon 359 -621 359 -621 0 3
rlabel polysilicon 366 -615 366 -615 0 1
rlabel polysilicon 366 -621 366 -621 0 3
rlabel polysilicon 373 -615 373 -615 0 1
rlabel polysilicon 373 -621 373 -621 0 3
rlabel polysilicon 380 -615 380 -615 0 1
rlabel polysilicon 380 -621 380 -621 0 3
rlabel polysilicon 387 -615 387 -615 0 1
rlabel polysilicon 387 -621 387 -621 0 3
rlabel polysilicon 394 -615 394 -615 0 1
rlabel polysilicon 394 -621 394 -621 0 3
rlabel polysilicon 401 -615 401 -615 0 1
rlabel polysilicon 401 -621 401 -621 0 3
rlabel polysilicon 408 -615 408 -615 0 1
rlabel polysilicon 408 -621 408 -621 0 3
rlabel polysilicon 415 -615 415 -615 0 1
rlabel polysilicon 415 -621 415 -621 0 3
rlabel polysilicon 422 -615 422 -615 0 1
rlabel polysilicon 422 -621 422 -621 0 3
rlabel polysilicon 429 -615 429 -615 0 1
rlabel polysilicon 429 -621 429 -621 0 3
rlabel polysilicon 436 -615 436 -615 0 1
rlabel polysilicon 436 -621 436 -621 0 3
rlabel polysilicon 443 -615 443 -615 0 1
rlabel polysilicon 446 -615 446 -615 0 2
rlabel polysilicon 446 -621 446 -621 0 4
rlabel polysilicon 453 -615 453 -615 0 2
rlabel polysilicon 450 -621 450 -621 0 3
rlabel polysilicon 457 -615 457 -615 0 1
rlabel polysilicon 457 -621 457 -621 0 3
rlabel polysilicon 464 -615 464 -615 0 1
rlabel polysilicon 471 -615 471 -615 0 1
rlabel polysilicon 471 -621 471 -621 0 3
rlabel polysilicon 2 -666 2 -666 0 1
rlabel polysilicon 2 -672 2 -672 0 3
rlabel polysilicon 9 -666 9 -666 0 1
rlabel polysilicon 9 -672 9 -672 0 3
rlabel polysilicon 16 -666 16 -666 0 1
rlabel polysilicon 16 -672 16 -672 0 3
rlabel polysilicon 23 -666 23 -666 0 1
rlabel polysilicon 23 -672 23 -672 0 3
rlabel polysilicon 30 -666 30 -666 0 1
rlabel polysilicon 30 -672 30 -672 0 3
rlabel polysilicon 37 -666 37 -666 0 1
rlabel polysilicon 37 -672 37 -672 0 3
rlabel polysilicon 44 -666 44 -666 0 1
rlabel polysilicon 51 -666 51 -666 0 1
rlabel polysilicon 54 -666 54 -666 0 2
rlabel polysilicon 54 -672 54 -672 0 4
rlabel polysilicon 58 -666 58 -666 0 1
rlabel polysilicon 58 -672 58 -672 0 3
rlabel polysilicon 65 -666 65 -666 0 1
rlabel polysilicon 65 -672 65 -672 0 3
rlabel polysilicon 75 -666 75 -666 0 2
rlabel polysilicon 72 -672 72 -672 0 3
rlabel polysilicon 79 -666 79 -666 0 1
rlabel polysilicon 79 -672 79 -672 0 3
rlabel polysilicon 86 -666 86 -666 0 1
rlabel polysilicon 86 -672 86 -672 0 3
rlabel polysilicon 93 -666 93 -666 0 1
rlabel polysilicon 93 -672 93 -672 0 3
rlabel polysilicon 100 -666 100 -666 0 1
rlabel polysilicon 103 -666 103 -666 0 2
rlabel polysilicon 100 -672 100 -672 0 3
rlabel polysilicon 107 -666 107 -666 0 1
rlabel polysilicon 107 -672 107 -672 0 3
rlabel polysilicon 114 -666 114 -666 0 1
rlabel polysilicon 114 -672 114 -672 0 3
rlabel polysilicon 117 -672 117 -672 0 4
rlabel polysilicon 121 -666 121 -666 0 1
rlabel polysilicon 121 -672 121 -672 0 3
rlabel polysilicon 128 -666 128 -666 0 1
rlabel polysilicon 128 -672 128 -672 0 3
rlabel polysilicon 131 -672 131 -672 0 4
rlabel polysilicon 135 -666 135 -666 0 1
rlabel polysilicon 135 -672 135 -672 0 3
rlabel polysilicon 142 -666 142 -666 0 1
rlabel polysilicon 142 -672 142 -672 0 3
rlabel polysilicon 149 -666 149 -666 0 1
rlabel polysilicon 149 -672 149 -672 0 3
rlabel polysilicon 156 -666 156 -666 0 1
rlabel polysilicon 156 -672 156 -672 0 3
rlabel polysilicon 163 -666 163 -666 0 1
rlabel polysilicon 163 -672 163 -672 0 3
rlabel polysilicon 170 -666 170 -666 0 1
rlabel polysilicon 170 -672 170 -672 0 3
rlabel polysilicon 177 -666 177 -666 0 1
rlabel polysilicon 180 -666 180 -666 0 2
rlabel polysilicon 177 -672 177 -672 0 3
rlabel polysilicon 180 -672 180 -672 0 4
rlabel polysilicon 184 -666 184 -666 0 1
rlabel polysilicon 187 -666 187 -666 0 2
rlabel polysilicon 184 -672 184 -672 0 3
rlabel polysilicon 194 -666 194 -666 0 2
rlabel polysilicon 191 -672 191 -672 0 3
rlabel polysilicon 194 -672 194 -672 0 4
rlabel polysilicon 198 -666 198 -666 0 1
rlabel polysilicon 198 -672 198 -672 0 3
rlabel polysilicon 205 -666 205 -666 0 1
rlabel polysilicon 208 -666 208 -666 0 2
rlabel polysilicon 215 -666 215 -666 0 2
rlabel polysilicon 212 -672 212 -672 0 3
rlabel polysilicon 215 -672 215 -672 0 4
rlabel polysilicon 222 -666 222 -666 0 2
rlabel polysilicon 219 -672 219 -672 0 3
rlabel polysilicon 226 -666 226 -666 0 1
rlabel polysilicon 226 -672 226 -672 0 3
rlabel polysilicon 233 -666 233 -666 0 1
rlabel polysilicon 233 -672 233 -672 0 3
rlabel polysilicon 240 -666 240 -666 0 1
rlabel polysilicon 243 -666 243 -666 0 2
rlabel polysilicon 240 -672 240 -672 0 3
rlabel polysilicon 247 -666 247 -666 0 1
rlabel polysilicon 250 -666 250 -666 0 2
rlabel polysilicon 250 -672 250 -672 0 4
rlabel polysilicon 254 -666 254 -666 0 1
rlabel polysilicon 254 -672 254 -672 0 3
rlabel polysilicon 261 -666 261 -666 0 1
rlabel polysilicon 261 -672 261 -672 0 3
rlabel polysilicon 271 -666 271 -666 0 2
rlabel polysilicon 268 -672 268 -672 0 3
rlabel polysilicon 275 -666 275 -666 0 1
rlabel polysilicon 275 -672 275 -672 0 3
rlabel polysilicon 282 -666 282 -666 0 1
rlabel polysilicon 282 -672 282 -672 0 3
rlabel polysilicon 289 -666 289 -666 0 1
rlabel polysilicon 289 -672 289 -672 0 3
rlabel polysilicon 296 -666 296 -666 0 1
rlabel polysilicon 299 -666 299 -666 0 2
rlabel polysilicon 299 -672 299 -672 0 4
rlabel polysilicon 303 -666 303 -666 0 1
rlabel polysilicon 303 -672 303 -672 0 3
rlabel polysilicon 310 -666 310 -666 0 1
rlabel polysilicon 310 -672 310 -672 0 3
rlabel polysilicon 317 -666 317 -666 0 1
rlabel polysilicon 317 -672 317 -672 0 3
rlabel polysilicon 324 -666 324 -666 0 1
rlabel polysilicon 324 -672 324 -672 0 3
rlabel polysilicon 331 -666 331 -666 0 1
rlabel polysilicon 334 -672 334 -672 0 4
rlabel polysilicon 338 -666 338 -666 0 1
rlabel polysilicon 338 -672 338 -672 0 3
rlabel polysilicon 345 -666 345 -666 0 1
rlabel polysilicon 345 -672 345 -672 0 3
rlabel polysilicon 352 -666 352 -666 0 1
rlabel polysilicon 352 -672 352 -672 0 3
rlabel polysilicon 359 -666 359 -666 0 1
rlabel polysilicon 359 -672 359 -672 0 3
rlabel polysilicon 366 -666 366 -666 0 1
rlabel polysilicon 366 -672 366 -672 0 3
rlabel polysilicon 373 -666 373 -666 0 1
rlabel polysilicon 373 -672 373 -672 0 3
rlabel polysilicon 380 -666 380 -666 0 1
rlabel polysilicon 380 -672 380 -672 0 3
rlabel polysilicon 387 -666 387 -666 0 1
rlabel polysilicon 387 -672 387 -672 0 3
rlabel polysilicon 394 -666 394 -666 0 1
rlabel polysilicon 394 -672 394 -672 0 3
rlabel polysilicon 401 -666 401 -666 0 1
rlabel polysilicon 401 -672 401 -672 0 3
rlabel polysilicon 408 -666 408 -666 0 1
rlabel polysilicon 408 -672 408 -672 0 3
rlabel polysilicon 415 -666 415 -666 0 1
rlabel polysilicon 415 -672 415 -672 0 3
rlabel polysilicon 422 -666 422 -666 0 1
rlabel polysilicon 422 -672 422 -672 0 3
rlabel polysilicon 429 -666 429 -666 0 1
rlabel polysilicon 429 -672 429 -672 0 3
rlabel polysilicon 436 -666 436 -666 0 1
rlabel polysilicon 436 -672 436 -672 0 3
rlabel polysilicon 443 -666 443 -666 0 1
rlabel polysilicon 443 -672 443 -672 0 3
rlabel polysilicon 450 -666 450 -666 0 1
rlabel polysilicon 450 -672 450 -672 0 3
rlabel polysilicon 457 -666 457 -666 0 1
rlabel polysilicon 460 -666 460 -666 0 2
rlabel polysilicon 457 -672 457 -672 0 3
rlabel polysilicon 464 -666 464 -666 0 1
rlabel polysilicon 464 -672 464 -672 0 3
rlabel polysilicon 471 -666 471 -666 0 1
rlabel polysilicon 471 -672 471 -672 0 3
rlabel polysilicon 2 -717 2 -717 0 1
rlabel polysilicon 2 -723 2 -723 0 3
rlabel polysilicon 9 -717 9 -717 0 1
rlabel polysilicon 9 -723 9 -723 0 3
rlabel polysilicon 16 -717 16 -717 0 1
rlabel polysilicon 16 -723 16 -723 0 3
rlabel polysilicon 23 -717 23 -717 0 1
rlabel polysilicon 23 -723 23 -723 0 3
rlabel polysilicon 30 -717 30 -717 0 1
rlabel polysilicon 30 -723 30 -723 0 3
rlabel polysilicon 37 -717 37 -717 0 1
rlabel polysilicon 40 -717 40 -717 0 2
rlabel polysilicon 37 -723 37 -723 0 3
rlabel polysilicon 44 -717 44 -717 0 1
rlabel polysilicon 44 -723 44 -723 0 3
rlabel polysilicon 51 -717 51 -717 0 1
rlabel polysilicon 54 -723 54 -723 0 4
rlabel polysilicon 58 -717 58 -717 0 1
rlabel polysilicon 58 -723 58 -723 0 3
rlabel polysilicon 65 -717 65 -717 0 1
rlabel polysilicon 65 -723 65 -723 0 3
rlabel polysilicon 72 -717 72 -717 0 1
rlabel polysilicon 75 -717 75 -717 0 2
rlabel polysilicon 75 -723 75 -723 0 4
rlabel polysilicon 82 -717 82 -717 0 2
rlabel polysilicon 82 -723 82 -723 0 4
rlabel polysilicon 86 -717 86 -717 0 1
rlabel polysilicon 86 -723 86 -723 0 3
rlabel polysilicon 93 -717 93 -717 0 1
rlabel polysilicon 93 -723 93 -723 0 3
rlabel polysilicon 100 -717 100 -717 0 1
rlabel polysilicon 100 -723 100 -723 0 3
rlabel polysilicon 107 -717 107 -717 0 1
rlabel polysilicon 107 -723 107 -723 0 3
rlabel polysilicon 114 -717 114 -717 0 1
rlabel polysilicon 114 -723 114 -723 0 3
rlabel polysilicon 121 -717 121 -717 0 1
rlabel polysilicon 124 -717 124 -717 0 2
rlabel polysilicon 131 -717 131 -717 0 2
rlabel polysilicon 128 -723 128 -723 0 3
rlabel polysilicon 135 -717 135 -717 0 1
rlabel polysilicon 135 -723 135 -723 0 3
rlabel polysilicon 142 -717 142 -717 0 1
rlabel polysilicon 142 -723 142 -723 0 3
rlabel polysilicon 149 -717 149 -717 0 1
rlabel polysilicon 149 -723 149 -723 0 3
rlabel polysilicon 156 -717 156 -717 0 1
rlabel polysilicon 156 -723 156 -723 0 3
rlabel polysilicon 163 -717 163 -717 0 1
rlabel polysilicon 163 -723 163 -723 0 3
rlabel polysilicon 170 -717 170 -717 0 1
rlabel polysilicon 173 -717 173 -717 0 2
rlabel polysilicon 177 -717 177 -717 0 1
rlabel polysilicon 180 -723 180 -723 0 4
rlabel polysilicon 184 -717 184 -717 0 1
rlabel polysilicon 187 -717 187 -717 0 2
rlabel polysilicon 184 -723 184 -723 0 3
rlabel polysilicon 191 -717 191 -717 0 1
rlabel polysilicon 191 -723 191 -723 0 3
rlabel polysilicon 198 -717 198 -717 0 1
rlabel polysilicon 198 -723 198 -723 0 3
rlabel polysilicon 201 -723 201 -723 0 4
rlabel polysilicon 205 -717 205 -717 0 1
rlabel polysilicon 205 -723 205 -723 0 3
rlabel polysilicon 208 -723 208 -723 0 4
rlabel polysilicon 212 -717 212 -717 0 1
rlabel polysilicon 212 -723 212 -723 0 3
rlabel polysilicon 219 -717 219 -717 0 1
rlabel polysilicon 219 -723 219 -723 0 3
rlabel polysilicon 229 -717 229 -717 0 2
rlabel polysilicon 226 -723 226 -723 0 3
rlabel polysilicon 233 -717 233 -717 0 1
rlabel polysilicon 233 -723 233 -723 0 3
rlabel polysilicon 240 -717 240 -717 0 1
rlabel polysilicon 243 -723 243 -723 0 4
rlabel polysilicon 250 -717 250 -717 0 2
rlabel polysilicon 250 -723 250 -723 0 4
rlabel polysilicon 254 -717 254 -717 0 1
rlabel polysilicon 254 -723 254 -723 0 3
rlabel polysilicon 261 -717 261 -717 0 1
rlabel polysilicon 261 -723 261 -723 0 3
rlabel polysilicon 268 -717 268 -717 0 1
rlabel polysilicon 268 -723 268 -723 0 3
rlabel polysilicon 278 -723 278 -723 0 4
rlabel polysilicon 282 -717 282 -717 0 1
rlabel polysilicon 282 -723 282 -723 0 3
rlabel polysilicon 289 -717 289 -717 0 1
rlabel polysilicon 289 -723 289 -723 0 3
rlabel polysilicon 296 -717 296 -717 0 1
rlabel polysilicon 296 -723 296 -723 0 3
rlabel polysilicon 310 -717 310 -717 0 1
rlabel polysilicon 310 -723 310 -723 0 3
rlabel polysilicon 317 -717 317 -717 0 1
rlabel polysilicon 317 -723 317 -723 0 3
rlabel polysilicon 324 -717 324 -717 0 1
rlabel polysilicon 324 -723 324 -723 0 3
rlabel polysilicon 331 -717 331 -717 0 1
rlabel polysilicon 331 -723 331 -723 0 3
rlabel polysilicon 341 -723 341 -723 0 4
rlabel polysilicon 345 -717 345 -717 0 1
rlabel polysilicon 345 -723 345 -723 0 3
rlabel polysilicon 352 -717 352 -717 0 1
rlabel polysilicon 352 -723 352 -723 0 3
rlabel polysilicon 359 -717 359 -717 0 1
rlabel polysilicon 359 -723 359 -723 0 3
rlabel polysilicon 366 -717 366 -717 0 1
rlabel polysilicon 366 -723 366 -723 0 3
rlabel polysilicon 373 -717 373 -717 0 1
rlabel polysilicon 376 -723 376 -723 0 4
rlabel polysilicon 380 -717 380 -717 0 1
rlabel polysilicon 380 -723 380 -723 0 3
rlabel polysilicon 387 -717 387 -717 0 1
rlabel polysilicon 387 -723 387 -723 0 3
rlabel polysilicon 394 -717 394 -717 0 1
rlabel polysilicon 394 -723 394 -723 0 3
rlabel polysilicon 401 -717 401 -717 0 1
rlabel polysilicon 401 -723 401 -723 0 3
rlabel polysilicon 411 -723 411 -723 0 4
rlabel polysilicon 429 -717 429 -717 0 1
rlabel polysilicon 429 -723 429 -723 0 3
rlabel polysilicon 16 -770 16 -770 0 1
rlabel polysilicon 23 -770 23 -770 0 1
rlabel polysilicon 23 -776 23 -776 0 3
rlabel polysilicon 30 -776 30 -776 0 3
rlabel polysilicon 33 -776 33 -776 0 4
rlabel polysilicon 37 -770 37 -770 0 1
rlabel polysilicon 40 -770 40 -770 0 2
rlabel polysilicon 37 -776 37 -776 0 3
rlabel polysilicon 44 -770 44 -770 0 1
rlabel polysilicon 47 -776 47 -776 0 4
rlabel polysilicon 51 -770 51 -770 0 1
rlabel polysilicon 51 -776 51 -776 0 3
rlabel polysilicon 58 -770 58 -770 0 1
rlabel polysilicon 58 -776 58 -776 0 3
rlabel polysilicon 65 -770 65 -770 0 1
rlabel polysilicon 65 -776 65 -776 0 3
rlabel polysilicon 72 -770 72 -770 0 1
rlabel polysilicon 75 -770 75 -770 0 2
rlabel polysilicon 75 -776 75 -776 0 4
rlabel polysilicon 79 -770 79 -770 0 1
rlabel polysilicon 82 -770 82 -770 0 2
rlabel polysilicon 86 -770 86 -770 0 1
rlabel polysilicon 86 -776 86 -776 0 3
rlabel polysilicon 96 -770 96 -770 0 2
rlabel polysilicon 93 -776 93 -776 0 3
rlabel polysilicon 96 -776 96 -776 0 4
rlabel polysilicon 100 -770 100 -770 0 1
rlabel polysilicon 103 -770 103 -770 0 2
rlabel polysilicon 103 -776 103 -776 0 4
rlabel polysilicon 110 -770 110 -770 0 2
rlabel polysilicon 107 -776 107 -776 0 3
rlabel polysilicon 114 -770 114 -770 0 1
rlabel polysilicon 117 -776 117 -776 0 4
rlabel polysilicon 121 -770 121 -770 0 1
rlabel polysilicon 124 -776 124 -776 0 4
rlabel polysilicon 128 -770 128 -770 0 1
rlabel polysilicon 128 -776 128 -776 0 3
rlabel polysilicon 135 -770 135 -770 0 1
rlabel polysilicon 135 -776 135 -776 0 3
rlabel polysilicon 142 -770 142 -770 0 1
rlabel polysilicon 142 -776 142 -776 0 3
rlabel polysilicon 149 -770 149 -770 0 1
rlabel polysilicon 149 -776 149 -776 0 3
rlabel polysilicon 156 -770 156 -770 0 1
rlabel polysilicon 156 -776 156 -776 0 3
rlabel polysilicon 163 -770 163 -770 0 1
rlabel polysilicon 163 -776 163 -776 0 3
rlabel polysilicon 170 -770 170 -770 0 1
rlabel polysilicon 170 -776 170 -776 0 3
rlabel polysilicon 180 -770 180 -770 0 2
rlabel polysilicon 177 -776 177 -776 0 3
rlabel polysilicon 184 -770 184 -770 0 1
rlabel polysilicon 184 -776 184 -776 0 3
rlabel polysilicon 191 -770 191 -770 0 1
rlabel polysilicon 191 -776 191 -776 0 3
rlabel polysilicon 198 -770 198 -770 0 1
rlabel polysilicon 198 -776 198 -776 0 3
rlabel polysilicon 208 -770 208 -770 0 2
rlabel polysilicon 212 -770 212 -770 0 1
rlabel polysilicon 215 -770 215 -770 0 2
rlabel polysilicon 212 -776 212 -776 0 3
rlabel polysilicon 219 -770 219 -770 0 1
rlabel polysilicon 219 -776 219 -776 0 3
rlabel polysilicon 226 -770 226 -770 0 1
rlabel polysilicon 226 -776 226 -776 0 3
rlabel polysilicon 233 -770 233 -770 0 1
rlabel polysilicon 236 -770 236 -770 0 2
rlabel polysilicon 236 -776 236 -776 0 4
rlabel polysilicon 240 -770 240 -770 0 1
rlabel polysilicon 240 -776 240 -776 0 3
rlabel polysilicon 247 -770 247 -770 0 1
rlabel polysilicon 247 -776 247 -776 0 3
rlabel polysilicon 254 -770 254 -770 0 1
rlabel polysilicon 254 -776 254 -776 0 3
rlabel polysilicon 261 -770 261 -770 0 1
rlabel polysilicon 261 -776 261 -776 0 3
rlabel polysilicon 268 -770 268 -770 0 1
rlabel polysilicon 268 -776 268 -776 0 3
rlabel polysilicon 275 -776 275 -776 0 3
rlabel polysilicon 282 -770 282 -770 0 1
rlabel polysilicon 282 -776 282 -776 0 3
rlabel polysilicon 289 -770 289 -770 0 1
rlabel polysilicon 289 -776 289 -776 0 3
rlabel polysilicon 303 -770 303 -770 0 1
rlabel polysilicon 303 -776 303 -776 0 3
rlabel polysilicon 310 -770 310 -770 0 1
rlabel polysilicon 310 -776 310 -776 0 3
rlabel polysilicon 324 -770 324 -770 0 1
rlabel polysilicon 324 -776 324 -776 0 3
rlabel polysilicon 331 -770 331 -770 0 1
rlabel polysilicon 338 -770 338 -770 0 1
rlabel polysilicon 338 -776 338 -776 0 3
rlabel polysilicon 345 -770 345 -770 0 1
rlabel polysilicon 345 -776 345 -776 0 3
rlabel polysilicon 408 -770 408 -770 0 1
rlabel polysilicon 9 -815 9 -815 0 1
rlabel polysilicon 9 -821 9 -821 0 3
rlabel polysilicon 16 -821 16 -821 0 3
rlabel polysilicon 23 -815 23 -815 0 1
rlabel polysilicon 23 -821 23 -821 0 3
rlabel polysilicon 30 -815 30 -815 0 1
rlabel polysilicon 33 -815 33 -815 0 2
rlabel polysilicon 33 -821 33 -821 0 4
rlabel polysilicon 37 -815 37 -815 0 1
rlabel polysilicon 37 -821 37 -821 0 3
rlabel polysilicon 44 -821 44 -821 0 3
rlabel polysilicon 47 -821 47 -821 0 4
rlabel polysilicon 51 -815 51 -815 0 1
rlabel polysilicon 51 -821 51 -821 0 3
rlabel polysilicon 61 -815 61 -815 0 2
rlabel polysilicon 65 -821 65 -821 0 3
rlabel polysilicon 72 -815 72 -815 0 1
rlabel polysilicon 72 -821 72 -821 0 3
rlabel polysilicon 79 -815 79 -815 0 1
rlabel polysilicon 82 -815 82 -815 0 2
rlabel polysilicon 89 -821 89 -821 0 4
rlabel polysilicon 96 -821 96 -821 0 4
rlabel polysilicon 100 -815 100 -815 0 1
rlabel polysilicon 100 -821 100 -821 0 3
rlabel polysilicon 107 -815 107 -815 0 1
rlabel polysilicon 110 -815 110 -815 0 2
rlabel polysilicon 114 -815 114 -815 0 1
rlabel polysilicon 117 -815 117 -815 0 2
rlabel polysilicon 114 -821 114 -821 0 3
rlabel polysilicon 117 -821 117 -821 0 4
rlabel polysilicon 124 -815 124 -815 0 2
rlabel polysilicon 131 -815 131 -815 0 2
rlabel polysilicon 128 -821 128 -821 0 3
rlabel polysilicon 135 -815 135 -815 0 1
rlabel polysilicon 135 -821 135 -821 0 3
rlabel polysilicon 145 -821 145 -821 0 4
rlabel polysilicon 152 -815 152 -815 0 2
rlabel polysilicon 152 -821 152 -821 0 4
rlabel polysilicon 156 -815 156 -815 0 1
rlabel polysilicon 156 -821 156 -821 0 3
rlabel polysilicon 163 -815 163 -815 0 1
rlabel polysilicon 163 -821 163 -821 0 3
rlabel polysilicon 170 -815 170 -815 0 1
rlabel polysilicon 170 -821 170 -821 0 3
rlabel polysilicon 177 -815 177 -815 0 1
rlabel polysilicon 180 -821 180 -821 0 4
rlabel polysilicon 184 -815 184 -815 0 1
rlabel polysilicon 184 -821 184 -821 0 3
rlabel polysilicon 191 -815 191 -815 0 1
rlabel polysilicon 191 -821 191 -821 0 3
rlabel polysilicon 198 -815 198 -815 0 1
rlabel polysilicon 198 -821 198 -821 0 3
rlabel polysilicon 205 -815 205 -815 0 1
rlabel polysilicon 205 -821 205 -821 0 3
rlabel polysilicon 212 -815 212 -815 0 1
rlabel polysilicon 212 -821 212 -821 0 3
rlabel polysilicon 222 -821 222 -821 0 4
rlabel polysilicon 226 -815 226 -815 0 1
rlabel polysilicon 226 -821 226 -821 0 3
rlabel polysilicon 233 -815 233 -815 0 1
rlabel polysilicon 233 -821 233 -821 0 3
rlabel polysilicon 240 -821 240 -821 0 3
rlabel polysilicon 247 -815 247 -815 0 1
rlabel polysilicon 247 -821 247 -821 0 3
rlabel polysilicon 254 -815 254 -815 0 1
rlabel polysilicon 254 -821 254 -821 0 3
rlabel polysilicon 261 -815 261 -815 0 1
rlabel polysilicon 261 -821 261 -821 0 3
rlabel polysilicon 268 -815 268 -815 0 1
rlabel polysilicon 268 -821 268 -821 0 3
rlabel polysilicon 282 -815 282 -815 0 1
rlabel polysilicon 282 -821 282 -821 0 3
rlabel polysilicon 289 -815 289 -815 0 1
rlabel polysilicon 289 -821 289 -821 0 3
rlabel polysilicon 303 -815 303 -815 0 1
rlabel polysilicon 303 -821 303 -821 0 3
rlabel polysilicon 310 -815 310 -815 0 1
rlabel polysilicon 310 -821 310 -821 0 3
rlabel polysilicon 317 -815 317 -815 0 1
rlabel polysilicon 317 -821 317 -821 0 3
rlabel polysilicon 324 -815 324 -815 0 1
rlabel polysilicon 324 -821 324 -821 0 3
rlabel polysilicon 345 -821 345 -821 0 3
rlabel polysilicon 19 -848 19 -848 0 2
rlabel polysilicon 23 -848 23 -848 0 1
rlabel polysilicon 23 -854 23 -854 0 3
rlabel polysilicon 33 -848 33 -848 0 2
rlabel polysilicon 37 -848 37 -848 0 1
rlabel polysilicon 37 -854 37 -854 0 3
rlabel polysilicon 44 -848 44 -848 0 1
rlabel polysilicon 44 -854 44 -854 0 3
rlabel polysilicon 47 -854 47 -854 0 4
rlabel polysilicon 51 -848 51 -848 0 1
rlabel polysilicon 54 -854 54 -854 0 4
rlabel polysilicon 58 -848 58 -848 0 1
rlabel polysilicon 58 -854 58 -854 0 3
rlabel polysilicon 65 -854 65 -854 0 3
rlabel polysilicon 72 -848 72 -848 0 1
rlabel polysilicon 72 -854 72 -854 0 3
rlabel polysilicon 79 -848 79 -848 0 1
rlabel polysilicon 82 -854 82 -854 0 4
rlabel polysilicon 86 -848 86 -848 0 1
rlabel polysilicon 86 -854 86 -854 0 3
rlabel polysilicon 93 -848 93 -848 0 1
rlabel polysilicon 93 -854 93 -854 0 3
rlabel polysilicon 103 -854 103 -854 0 4
rlabel polysilicon 107 -854 107 -854 0 3
rlabel polysilicon 117 -848 117 -848 0 2
rlabel polysilicon 114 -854 114 -854 0 3
rlabel polysilicon 124 -848 124 -848 0 2
rlabel polysilicon 131 -854 131 -854 0 4
rlabel polysilicon 135 -848 135 -848 0 1
rlabel polysilicon 142 -854 142 -854 0 3
rlabel polysilicon 149 -848 149 -848 0 1
rlabel polysilicon 149 -854 149 -854 0 3
rlabel polysilicon 156 -848 156 -848 0 1
rlabel polysilicon 156 -854 156 -854 0 3
rlabel polysilicon 163 -848 163 -848 0 1
rlabel polysilicon 163 -854 163 -854 0 3
rlabel polysilicon 170 -848 170 -848 0 1
rlabel polysilicon 170 -854 170 -854 0 3
rlabel polysilicon 184 -848 184 -848 0 1
rlabel polysilicon 187 -854 187 -854 0 4
rlabel polysilicon 191 -848 191 -848 0 1
rlabel polysilicon 191 -854 191 -854 0 3
rlabel polysilicon 212 -848 212 -848 0 1
rlabel polysilicon 226 -848 226 -848 0 1
rlabel polysilicon 268 -848 268 -848 0 1
rlabel polysilicon 268 -854 268 -854 0 3
rlabel polysilicon 282 -848 282 -848 0 1
rlabel polysilicon 285 -854 285 -854 0 4
rlabel polysilicon 289 -848 289 -848 0 1
rlabel polysilicon 292 -848 292 -848 0 2
rlabel polysilicon 327 -848 327 -848 0 2
rlabel metal2 12 1 12 1 0 net=45
rlabel metal2 37 1 37 1 0 net=435
rlabel metal2 93 1 93 1 0 net=1637
rlabel metal2 121 1 121 1 0 net=369
rlabel metal2 135 1 135 1 0 net=1639
rlabel metal2 51 -1 51 -1 0 net=87
rlabel metal2 138 -1 138 -1 0 net=1183
rlabel metal2 58 -3 58 -3 0 net=307
rlabel metal2 72 -14 72 -14 0 net=132
rlabel metal2 100 -14 100 -14 0 net=1638
rlabel metal2 114 -14 114 -14 0 net=177
rlabel metal2 159 -14 159 -14 0 net=63
rlabel metal2 65 -16 65 -16 0 net=437
rlabel metal2 79 -16 79 -16 0 net=95
rlabel metal2 107 -16 107 -16 0 net=1265
rlabel metal2 145 -16 145 -16 0 net=1184
rlabel metal2 163 -16 163 -16 0 net=1640
rlabel metal2 114 -18 114 -18 0 net=1313
rlabel metal2 128 -20 128 -20 0 net=371
rlabel metal2 128 -20 128 -20 0 net=371
rlabel metal2 149 -20 149 -20 0 net=973
rlabel metal2 163 -22 163 -22 0 net=1319
rlabel metal2 5 -33 5 -33 0 net=295
rlabel metal2 5 -33 5 -33 0 net=295
rlabel metal2 30 -33 30 -33 0 net=64
rlabel metal2 30 -33 30 -33 0 net=64
rlabel metal2 47 -33 47 -33 0 net=1205
rlabel metal2 51 -35 51 -35 0 net=975
rlabel metal2 163 -35 163 -35 0 net=1321
rlabel metal2 58 -37 58 -37 0 net=439
rlabel metal2 86 -37 86 -37 0 net=859
rlabel metal2 177 -37 177 -37 0 net=1315
rlabel metal2 16 -39 16 -39 0 net=921
rlabel metal2 191 -39 191 -39 0 net=1619
rlabel metal2 65 -41 65 -41 0 net=1229
rlabel metal2 121 -41 121 -41 0 net=887
rlabel metal2 198 -41 198 -41 0 net=1353
rlabel metal2 72 -43 72 -43 0 net=423
rlabel metal2 93 -43 93 -43 0 net=927
rlabel metal2 37 -45 37 -45 0 net=17
rlabel metal2 96 -45 96 -45 0 net=1045
rlabel metal2 124 -47 124 -47 0 net=319
rlabel metal2 100 -49 100 -49 0 net=505
rlabel metal2 128 -49 128 -49 0 net=372
rlabel metal2 128 -49 128 -49 0 net=372
rlabel metal2 142 -49 142 -49 0 net=1267
rlabel metal2 145 -51 145 -51 0 net=727
rlabel metal2 149 -53 149 -53 0 net=1049
rlabel metal2 19 -64 19 -64 0 net=1206
rlabel metal2 219 -64 219 -64 0 net=1323
rlabel metal2 40 -66 40 -66 0 net=60
rlabel metal2 82 -66 82 -66 0 net=24
rlabel metal2 121 -66 121 -66 0 net=471
rlabel metal2 177 -66 177 -66 0 net=923
rlabel metal2 226 -66 226 -66 0 net=1269
rlabel metal2 40 -68 40 -68 0 net=755
rlabel metal2 191 -68 191 -68 0 net=1620
rlabel metal2 44 -70 44 -70 0 net=977
rlabel metal2 58 -70 58 -70 0 net=440
rlabel metal2 100 -70 100 -70 0 net=506
rlabel metal2 131 -70 131 -70 0 net=667
rlabel metal2 30 -72 30 -72 0 net=277
rlabel metal2 138 -72 138 -72 0 net=250
rlabel metal2 149 -72 149 -72 0 net=891
rlabel metal2 233 -72 233 -72 0 net=1317
rlabel metal2 30 -74 30 -74 0 net=819
rlabel metal2 163 -74 163 -74 0 net=861
rlabel metal2 243 -74 243 -74 0 net=1185
rlabel metal2 51 -76 51 -76 0 net=573
rlabel metal2 107 -76 107 -76 0 net=353
rlabel metal2 184 -76 184 -76 0 net=929
rlabel metal2 205 -76 205 -76 0 net=1051
rlabel metal2 247 -76 247 -76 0 net=1355
rlabel metal2 58 -78 58 -78 0 net=1231
rlabel metal2 86 -78 86 -78 0 net=729
rlabel metal2 170 -78 170 -78 0 net=889
rlabel metal2 65 -80 65 -80 0 net=425
rlabel metal2 110 -80 110 -80 0 net=873
rlabel metal2 72 -82 72 -82 0 net=557
rlabel metal2 170 -82 170 -82 0 net=1555
rlabel metal2 184 -84 184 -84 0 net=1029
rlabel metal2 198 -86 198 -86 0 net=1047
rlabel metal2 23 -97 23 -97 0 net=730
rlabel metal2 93 -97 93 -97 0 net=581
rlabel metal2 135 -97 135 -97 0 net=862
rlabel metal2 268 -97 268 -97 0 net=1357
rlabel metal2 26 -99 26 -99 0 net=1341
rlabel metal2 30 -101 30 -101 0 net=820
rlabel metal2 201 -101 201 -101 0 net=1215
rlabel metal2 331 -101 331 -101 0 net=1271
rlabel metal2 331 -101 331 -101 0 net=1271
rlabel metal2 51 -103 51 -103 0 net=575
rlabel metal2 107 -103 107 -103 0 net=551
rlabel metal2 121 -103 121 -103 0 net=473
rlabel metal2 145 -103 145 -103 0 net=971
rlabel metal2 51 -105 51 -105 0 net=427
rlabel metal2 96 -105 96 -105 0 net=668
rlabel metal2 271 -105 271 -105 0 net=1447
rlabel metal2 58 -107 58 -107 0 net=1232
rlabel metal2 58 -107 58 -107 0 net=1232
rlabel metal2 65 -107 65 -107 0 net=461
rlabel metal2 194 -107 194 -107 0 net=781
rlabel metal2 254 -107 254 -107 0 net=1187
rlabel metal2 275 -107 275 -107 0 net=1325
rlabel metal2 30 -109 30 -109 0 net=983
rlabel metal2 289 -109 289 -109 0 net=1557
rlabel metal2 86 -111 86 -111 0 net=965
rlabel metal2 303 -111 303 -111 0 net=1243
rlabel metal2 128 -113 128 -113 0 net=1048
rlabel metal2 138 -115 138 -115 0 net=1081
rlabel metal2 138 -117 138 -117 0 net=268
rlabel metal2 233 -117 233 -117 0 net=1031
rlabel metal2 149 -119 149 -119 0 net=890
rlabel metal2 233 -119 233 -119 0 net=875
rlabel metal2 149 -121 149 -121 0 net=252
rlabel metal2 240 -121 240 -121 0 net=1053
rlabel metal2 152 -123 152 -123 0 net=513
rlabel metal2 191 -123 191 -123 0 net=931
rlabel metal2 156 -125 156 -125 0 net=1295
rlabel metal2 44 -127 44 -127 0 net=979
rlabel metal2 163 -127 163 -127 0 net=1318
rlabel metal2 9 -129 9 -129 0 net=599
rlabel metal2 124 -129 124 -129 0 net=334
rlabel metal2 166 -129 166 -129 0 net=924
rlabel metal2 37 -131 37 -131 0 net=1015
rlabel metal2 166 -133 166 -133 0 net=671
rlabel metal2 212 -133 212 -133 0 net=893
rlabel metal2 128 -135 128 -135 0 net=689
rlabel metal2 177 -137 177 -137 0 net=757
rlabel metal2 72 -139 72 -139 0 net=559
rlabel metal2 72 -141 72 -141 0 net=441
rlabel metal2 5 -152 5 -152 0 net=331
rlabel metal2 23 -152 23 -152 0 net=972
rlabel metal2 324 -152 324 -152 0 net=1245
rlabel metal2 324 -152 324 -152 0 net=1245
rlabel metal2 331 -152 331 -152 0 net=1273
rlabel metal2 331 -152 331 -152 0 net=1273
rlabel metal2 345 -152 345 -152 0 net=1327
rlabel metal2 9 -154 9 -154 0 net=1595
rlabel metal2 61 -154 61 -154 0 net=1296
rlabel metal2 345 -154 345 -154 0 net=1343
rlabel metal2 373 -154 373 -154 0 net=1559
rlabel metal2 16 -156 16 -156 0 net=127
rlabel metal2 65 -156 65 -156 0 net=462
rlabel metal2 128 -156 128 -156 0 net=1032
rlabel metal2 338 -156 338 -156 0 net=1449
rlabel metal2 16 -158 16 -158 0 net=429
rlabel metal2 86 -158 86 -158 0 net=1082
rlabel metal2 320 -158 320 -158 0 net=1403
rlabel metal2 23 -160 23 -160 0 net=287
rlabel metal2 37 -160 37 -160 0 net=553
rlabel metal2 128 -160 128 -160 0 net=280
rlabel metal2 208 -160 208 -160 0 net=1358
rlabel metal2 30 -162 30 -162 0 net=451
rlabel metal2 191 -162 191 -162 0 net=1445
rlabel metal2 51 -164 51 -164 0 net=1227
rlabel metal2 107 -164 107 -164 0 net=483
rlabel metal2 222 -164 222 -164 0 net=1529
rlabel metal2 79 -166 79 -166 0 net=249
rlabel metal2 226 -166 226 -166 0 net=783
rlabel metal2 359 -166 359 -166 0 net=1365
rlabel metal2 65 -168 65 -168 0 net=447
rlabel metal2 86 -168 86 -168 0 net=583
rlabel metal2 149 -168 149 -168 0 net=672
rlabel metal2 194 -168 194 -168 0 net=1054
rlabel metal2 89 -170 89 -170 0 net=474
rlabel metal2 149 -170 149 -170 0 net=1005
rlabel metal2 72 -172 72 -172 0 net=443
rlabel metal2 152 -172 152 -172 0 net=932
rlabel metal2 261 -172 261 -172 0 net=1189
rlabel metal2 47 -174 47 -174 0 net=79
rlabel metal2 156 -174 156 -174 0 net=980
rlabel metal2 198 -174 198 -174 0 net=1621
rlabel metal2 100 -176 100 -176 0 net=577
rlabel metal2 163 -176 163 -176 0 net=894
rlabel metal2 261 -176 261 -176 0 net=1017
rlabel metal2 75 -178 75 -178 0 net=346
rlabel metal2 166 -178 166 -178 0 net=733
rlabel metal2 82 -180 82 -180 0 net=1535
rlabel metal2 254 -180 254 -180 0 net=967
rlabel metal2 82 -182 82 -182 0 net=211
rlabel metal2 177 -182 177 -182 0 net=561
rlabel metal2 208 -182 208 -182 0 net=633
rlabel metal2 233 -182 233 -182 0 net=877
rlabel metal2 268 -182 268 -182 0 net=1216
rlabel metal2 100 -184 100 -184 0 net=199
rlabel metal2 152 -184 152 -184 0 net=795
rlabel metal2 275 -184 275 -184 0 net=985
rlabel metal2 61 -186 61 -186 0 net=735
rlabel metal2 114 -188 114 -188 0 net=491
rlabel metal2 170 -188 170 -188 0 net=515
rlabel metal2 212 -188 212 -188 0 net=691
rlabel metal2 44 -190 44 -190 0 net=601
rlabel metal2 219 -190 219 -190 0 net=759
rlabel metal2 58 -192 58 -192 0 net=585
rlabel metal2 219 -192 219 -192 0 net=1359
rlabel metal2 16 -203 16 -203 0 net=430
rlabel metal2 86 -203 86 -203 0 net=584
rlabel metal2 166 -203 166 -203 0 net=784
rlabel metal2 324 -203 324 -203 0 net=1247
rlabel metal2 324 -203 324 -203 0 net=1247
rlabel metal2 331 -203 331 -203 0 net=1275
rlabel metal2 331 -203 331 -203 0 net=1275
rlabel metal2 401 -203 401 -203 0 net=1561
rlabel metal2 401 -203 401 -203 0 net=1561
rlabel metal2 16 -205 16 -205 0 net=703
rlabel metal2 184 -205 184 -205 0 net=1530
rlabel metal2 23 -207 23 -207 0 net=485
rlabel metal2 110 -207 110 -207 0 net=281
rlabel metal2 205 -207 205 -207 0 net=1446
rlabel metal2 44 -209 44 -209 0 net=602
rlabel metal2 117 -209 117 -209 0 net=736
rlabel metal2 338 -209 338 -209 0 net=1451
rlabel metal2 44 -211 44 -211 0 net=933
rlabel metal2 107 -211 107 -211 0 net=1035
rlabel metal2 338 -211 338 -211 0 net=1345
rlabel metal2 54 -213 54 -213 0 net=283
rlabel metal2 219 -213 219 -213 0 net=1190
rlabel metal2 65 -215 65 -215 0 net=448
rlabel metal2 86 -215 86 -215 0 net=857
rlabel metal2 124 -215 124 -215 0 net=50
rlabel metal2 138 -215 138 -215 0 net=562
rlabel metal2 240 -215 240 -215 0 net=1537
rlabel metal2 30 -217 30 -217 0 net=453
rlabel metal2 142 -217 142 -217 0 net=445
rlabel metal2 170 -217 170 -217 0 net=693
rlabel metal2 247 -217 247 -217 0 net=879
rlabel metal2 247 -217 247 -217 0 net=879
rlabel metal2 275 -217 275 -217 0 net=987
rlabel metal2 310 -217 310 -217 0 net=1623
rlabel metal2 9 -219 9 -219 0 net=1596
rlabel metal2 37 -219 37 -219 0 net=555
rlabel metal2 177 -219 177 -219 0 net=517
rlabel metal2 289 -219 289 -219 0 net=1007
rlabel metal2 345 -219 345 -219 0 net=1361
rlabel metal2 9 -221 9 -221 0 net=46
rlabel metal2 93 -221 93 -221 0 net=578
rlabel metal2 187 -221 187 -221 0 net=1077
rlabel metal2 352 -221 352 -221 0 net=1367
rlabel metal2 37 -223 37 -223 0 net=499
rlabel metal2 96 -223 96 -223 0 net=734
rlabel metal2 65 -225 65 -225 0 net=995
rlabel metal2 121 -225 121 -225 0 net=493
rlabel metal2 187 -225 187 -225 0 net=809
rlabel metal2 222 -225 222 -225 0 net=218
rlabel metal2 261 -225 261 -225 0 net=1019
rlabel metal2 359 -225 359 -225 0 net=1405
rlabel metal2 51 -227 51 -227 0 net=1228
rlabel metal2 121 -229 121 -229 0 net=1419
rlabel metal2 135 -231 135 -231 0 net=1545
rlabel metal2 149 -233 149 -233 0 net=527
rlabel metal2 191 -233 191 -233 0 net=587
rlabel metal2 201 -235 201 -235 0 net=949
rlabel metal2 201 -237 201 -237 0 net=1328
rlabel metal2 58 -239 58 -239 0 net=1495
rlabel metal2 58 -241 58 -241 0 net=635
rlabel metal2 212 -243 212 -243 0 net=761
rlabel metal2 226 -245 226 -245 0 net=797
rlabel metal2 254 -247 254 -247 0 net=1607
rlabel metal2 268 -249 268 -249 0 net=969
rlabel metal2 282 -251 282 -251 0 net=1059
rlabel metal2 12 -262 12 -262 0 net=1346
rlabel metal2 380 -262 380 -262 0 net=1497
rlabel metal2 33 -264 33 -264 0 net=339
rlabel metal2 61 -264 61 -264 0 net=996
rlabel metal2 72 -264 72 -264 0 net=306
rlabel metal2 110 -264 110 -264 0 net=970
rlabel metal2 282 -264 282 -264 0 net=1087
rlabel metal2 37 -266 37 -266 0 net=501
rlabel metal2 75 -266 75 -266 0 net=33
rlabel metal2 149 -266 149 -266 0 net=529
rlabel metal2 149 -266 149 -266 0 net=529
rlabel metal2 163 -266 163 -266 0 net=446
rlabel metal2 226 -266 226 -266 0 net=798
rlabel metal2 30 -268 30 -268 0 net=853
rlabel metal2 173 -268 173 -268 0 net=762
rlabel metal2 240 -268 240 -268 0 net=1008
rlabel metal2 338 -268 338 -268 0 net=1363
rlabel metal2 380 -268 380 -268 0 net=1379
rlabel metal2 37 -270 37 -270 0 net=637
rlabel metal2 86 -270 86 -270 0 net=858
rlabel metal2 117 -270 117 -270 0 net=556
rlabel metal2 177 -270 177 -270 0 net=367
rlabel metal2 205 -270 205 -270 0 net=811
rlabel metal2 247 -270 247 -270 0 net=880
rlabel metal2 268 -270 268 -270 0 net=1079
rlabel metal2 345 -270 345 -270 0 net=1453
rlabel metal2 394 -270 394 -270 0 net=1547
rlabel metal2 51 -272 51 -272 0 net=1531
rlabel metal2 212 -272 212 -272 0 net=1020
rlabel metal2 317 -272 317 -272 0 net=1277
rlabel metal2 366 -272 366 -272 0 net=1421
rlabel metal2 394 -272 394 -272 0 net=1625
rlabel metal2 79 -274 79 -274 0 net=937
rlabel metal2 96 -274 96 -274 0 net=1111
rlabel metal2 331 -274 331 -274 0 net=1369
rlabel metal2 359 -274 359 -274 0 net=1407
rlabel metal2 401 -274 401 -274 0 net=1563
rlabel metal2 23 -276 23 -276 0 net=487
rlabel metal2 100 -276 100 -276 0 net=459
rlabel metal2 180 -276 180 -276 0 net=518
rlabel metal2 250 -276 250 -276 0 net=1538
rlabel metal2 401 -276 401 -276 0 net=1609
rlabel metal2 23 -278 23 -278 0 net=935
rlabel metal2 100 -278 100 -278 0 net=494
rlabel metal2 184 -278 184 -278 0 net=989
rlabel metal2 44 -280 44 -280 0 net=537
rlabel metal2 205 -280 205 -280 0 net=1381
rlabel metal2 103 -282 103 -282 0 net=694
rlabel metal2 198 -282 198 -282 0 net=1217
rlabel metal2 128 -284 128 -284 0 net=454
rlabel metal2 254 -284 254 -284 0 net=951
rlabel metal2 275 -284 275 -284 0 net=1061
rlabel metal2 16 -286 16 -286 0 net=704
rlabel metal2 264 -286 264 -286 0 net=1257
rlabel metal2 16 -288 16 -288 0 net=1589
rlabel metal2 128 -290 128 -290 0 net=801
rlabel metal2 219 -290 219 -290 0 net=955
rlabel metal2 135 -292 135 -292 0 net=1489
rlabel metal2 93 -294 93 -294 0 net=613
rlabel metal2 156 -294 156 -294 0 net=589
rlabel metal2 222 -294 222 -294 0 net=1385
rlabel metal2 166 -296 166 -296 0 net=571
rlabel metal2 233 -296 233 -296 0 net=1037
rlabel metal2 303 -298 303 -298 0 net=1249
rlabel metal2 124 -300 124 -300 0 net=1287
rlabel metal2 2 -311 2 -311 0 net=579
rlabel metal2 184 -311 184 -311 0 net=991
rlabel metal2 243 -311 243 -311 0 net=1364
rlabel metal2 401 -311 401 -311 0 net=1611
rlabel metal2 23 -313 23 -313 0 net=936
rlabel metal2 100 -313 100 -313 0 net=803
rlabel metal2 142 -313 142 -313 0 net=460
rlabel metal2 226 -313 226 -313 0 net=813
rlabel metal2 226 -313 226 -313 0 net=813
rlabel metal2 233 -313 233 -313 0 net=1039
rlabel metal2 264 -313 264 -313 0 net=1564
rlabel metal2 26 -315 26 -315 0 net=272
rlabel metal2 107 -315 107 -315 0 net=1579
rlabel metal2 30 -317 30 -317 0 net=854
rlabel metal2 191 -317 191 -317 0 net=572
rlabel metal2 247 -317 247 -317 0 net=953
rlabel metal2 275 -317 275 -317 0 net=1063
rlabel metal2 275 -317 275 -317 0 net=1063
rlabel metal2 317 -317 317 -317 0 net=1279
rlabel metal2 23 -319 23 -319 0 net=731
rlabel metal2 198 -319 198 -319 0 net=1250
rlabel metal2 317 -319 317 -319 0 net=1289
rlabel metal2 331 -319 331 -319 0 net=1371
rlabel metal2 331 -319 331 -319 0 net=1371
rlabel metal2 30 -321 30 -321 0 net=1422
rlabel metal2 37 -323 37 -323 0 net=638
rlabel metal2 198 -323 198 -323 0 net=957
rlabel metal2 250 -323 250 -323 0 net=1380
rlabel metal2 33 -325 33 -325 0 net=25
rlabel metal2 40 -325 40 -325 0 net=1499
rlabel metal2 44 -327 44 -327 0 net=538
rlabel metal2 142 -327 142 -327 0 net=639
rlabel metal2 254 -327 254 -327 0 net=1591
rlabel metal2 54 -329 54 -329 0 net=1161
rlabel metal2 345 -329 345 -329 0 net=1455
rlabel metal2 58 -331 58 -331 0 net=939
rlabel metal2 110 -331 110 -331 0 net=507
rlabel metal2 159 -331 159 -331 0 net=368
rlabel metal2 296 -331 296 -331 0 net=1219
rlabel metal2 373 -331 373 -331 0 net=1491
rlabel metal2 61 -333 61 -333 0 net=741
rlabel metal2 110 -333 110 -333 0 net=1213
rlabel metal2 65 -335 65 -335 0 net=503
rlabel metal2 233 -335 233 -335 0 net=1465
rlabel metal2 65 -337 65 -337 0 net=1155
rlabel metal2 72 -339 72 -339 0 net=1498
rlabel metal2 79 -341 79 -341 0 net=489
rlabel metal2 394 -341 394 -341 0 net=1627
rlabel metal2 16 -343 16 -343 0 net=1590
rlabel metal2 114 -343 114 -343 0 net=1055
rlabel metal2 366 -343 366 -343 0 net=1409
rlabel metal2 16 -345 16 -345 0 net=687
rlabel metal2 121 -345 121 -345 0 net=530
rlabel metal2 359 -345 359 -345 0 net=1387
rlabel metal2 117 -347 117 -347 0 net=749
rlabel metal2 135 -347 135 -347 0 net=615
rlabel metal2 352 -347 352 -347 0 net=1383
rlabel metal2 117 -349 117 -349 0 net=1548
rlabel metal2 51 -351 51 -351 0 net=1533
rlabel metal2 51 -353 51 -353 0 net=649
rlabel metal2 289 -353 289 -353 0 net=1113
rlabel metal2 135 -355 135 -355 0 net=591
rlabel metal2 289 -355 289 -355 0 net=1259
rlabel metal2 156 -357 156 -357 0 net=1080
rlabel metal2 282 -357 282 -357 0 net=1089
rlabel metal2 268 -359 268 -359 0 net=259
rlabel metal2 271 -361 271 -361 0 net=1165
rlabel metal2 2 -372 2 -372 0 net=580
rlabel metal2 201 -372 201 -372 0 net=98
rlabel metal2 222 -372 222 -372 0 net=1384
rlabel metal2 9 -374 9 -374 0 net=631
rlabel metal2 37 -374 37 -374 0 net=264
rlabel metal2 110 -374 110 -374 0 net=1388
rlabel metal2 16 -376 16 -376 0 net=688
rlabel metal2 26 -376 26 -376 0 net=301
rlabel metal2 247 -376 247 -376 0 net=954
rlabel metal2 268 -376 268 -376 0 net=1090
rlabel metal2 317 -376 317 -376 0 net=1291
rlabel metal2 16 -378 16 -378 0 net=1043
rlabel metal2 65 -378 65 -378 0 net=959
rlabel metal2 226 -378 226 -378 0 net=815
rlabel metal2 271 -378 271 -378 0 net=1410
rlabel metal2 30 -380 30 -380 0 net=997
rlabel metal2 68 -380 68 -380 0 net=732
rlabel metal2 271 -380 271 -380 0 net=1260
rlabel metal2 317 -380 317 -380 0 net=1221
rlabel metal2 338 -380 338 -380 0 net=1281
rlabel metal2 387 -380 387 -380 0 net=1467
rlabel metal2 37 -382 37 -382 0 net=941
rlabel metal2 79 -382 79 -382 0 net=161
rlabel metal2 61 -384 61 -384 0 net=475
rlabel metal2 82 -384 82 -384 0 net=1156
rlabel metal2 86 -386 86 -386 0 net=504
rlabel metal2 212 -386 212 -386 0 net=1057
rlabel metal2 72 -388 72 -388 0 net=563
rlabel metal2 110 -388 110 -388 0 net=1214
rlabel metal2 72 -390 72 -390 0 net=805
rlabel metal2 114 -390 114 -390 0 net=1534
rlabel metal2 100 -392 100 -392 0 net=490
rlabel metal2 184 -392 184 -392 0 net=785
rlabel metal2 229 -392 229 -392 0 net=1575
rlabel metal2 408 -392 408 -392 0 net=1613
rlabel metal2 117 -394 117 -394 0 net=1580
rlabel metal2 135 -396 135 -396 0 net=592
rlabel metal2 205 -396 205 -396 0 net=899
rlabel metal2 261 -396 261 -396 0 net=1041
rlabel metal2 352 -396 352 -396 0 net=1114
rlabel metal2 135 -398 135 -398 0 net=381
rlabel metal2 163 -398 163 -398 0 net=1157
rlabel metal2 331 -398 331 -398 0 net=1373
rlabel metal2 415 -398 415 -398 0 net=1593
rlabel metal2 142 -400 142 -400 0 net=641
rlabel metal2 212 -400 212 -400 0 net=993
rlabel metal2 261 -400 261 -400 0 net=1500
rlabel metal2 422 -400 422 -400 0 net=1629
rlabel metal2 93 -402 93 -402 0 net=743
rlabel metal2 149 -402 149 -402 0 net=650
rlabel metal2 184 -402 184 -402 0 net=393
rlabel metal2 275 -402 275 -402 0 net=1065
rlabel metal2 303 -402 303 -402 0 net=1163
rlabel metal2 373 -402 373 -402 0 net=1493
rlabel metal2 432 -402 432 -402 0 net=897
rlabel metal2 54 -404 54 -404 0 net=519
rlabel metal2 121 -404 121 -404 0 net=751
rlabel metal2 170 -404 170 -404 0 net=1129
rlabel metal2 373 -404 373 -404 0 net=1457
rlabel metal2 47 -406 47 -406 0 net=673
rlabel metal2 128 -406 128 -406 0 net=509
rlabel metal2 170 -406 170 -406 0 net=617
rlabel metal2 254 -406 254 -406 0 net=1261
rlabel metal2 282 -406 282 -406 0 net=1167
rlabel metal2 282 -406 282 -406 0 net=1167
rlabel metal2 58 -408 58 -408 0 net=1441
rlabel metal2 264 -408 264 -408 0 net=1501
rlabel metal2 117 -410 117 -410 0 net=1119
rlabel metal2 9 -421 9 -421 0 net=632
rlabel metal2 79 -421 79 -421 0 net=477
rlabel metal2 107 -421 107 -421 0 net=342
rlabel metal2 226 -421 226 -421 0 net=1164
rlabel metal2 432 -421 432 -421 0 net=1393
rlabel metal2 16 -423 16 -423 0 net=1044
rlabel metal2 37 -423 37 -423 0 net=943
rlabel metal2 37 -423 37 -423 0 net=943
rlabel metal2 44 -423 44 -423 0 net=744
rlabel metal2 166 -423 166 -423 0 net=618
rlabel metal2 194 -423 194 -423 0 net=994
rlabel metal2 229 -423 229 -423 0 net=1058
rlabel metal2 317 -423 317 -423 0 net=1223
rlabel metal2 359 -423 359 -423 0 net=1282
rlabel metal2 443 -423 443 -423 0 net=799
rlabel metal2 16 -425 16 -425 0 net=1101
rlabel metal2 30 -425 30 -425 0 net=998
rlabel metal2 79 -425 79 -425 0 net=565
rlabel metal2 93 -425 93 -425 0 net=520
rlabel metal2 121 -425 121 -425 0 net=675
rlabel metal2 163 -425 163 -425 0 net=1091
rlabel metal2 327 -425 327 -425 0 net=1630
rlabel metal2 446 -425 446 -425 0 net=1001
rlabel metal2 51 -427 51 -427 0 net=807
rlabel metal2 86 -427 86 -427 0 net=463
rlabel metal2 121 -427 121 -427 0 net=383
rlabel metal2 156 -427 156 -427 0 net=511
rlabel metal2 177 -427 177 -427 0 net=1443
rlabel metal2 334 -427 334 -427 0 net=1494
rlabel metal2 58 -429 58 -429 0 net=1085
rlabel metal2 114 -429 114 -429 0 net=541
rlabel metal2 201 -429 201 -429 0 net=1042
rlabel metal2 352 -429 352 -429 0 net=1375
rlabel metal2 93 -431 93 -431 0 net=925
rlabel metal2 212 -431 212 -431 0 net=816
rlabel metal2 236 -431 236 -431 0 net=1201
rlabel metal2 128 -433 128 -433 0 net=786
rlabel metal2 240 -433 240 -433 0 net=1631
rlabel metal2 117 -435 117 -435 0 net=1
rlabel metal2 131 -435 131 -435 0 net=752
rlabel metal2 156 -435 156 -435 0 net=643
rlabel metal2 243 -435 243 -435 0 net=1130
rlabel metal2 135 -437 135 -437 0 net=395
rlabel metal2 191 -437 191 -437 0 net=898
rlabel metal2 149 -439 149 -439 0 net=771
rlabel metal2 247 -439 247 -439 0 net=1066
rlabel metal2 387 -439 387 -439 0 net=1577
rlabel metal2 226 -441 226 -441 0 net=1139
rlabel metal2 387 -441 387 -441 0 net=1615
rlabel metal2 250 -443 250 -443 0 net=1468
rlabel metal2 250 -445 250 -445 0 net=1594
rlabel metal2 254 -447 254 -447 0 net=1121
rlabel metal2 310 -447 310 -447 0 net=1159
rlabel metal2 254 -449 254 -449 0 net=1297
rlabel metal2 373 -449 373 -449 0 net=1459
rlabel metal2 257 -451 257 -451 0 net=1292
rlabel metal2 373 -451 373 -451 0 net=1503
rlabel metal2 261 -453 261 -453 0 net=1175
rlabel metal2 170 -455 170 -455 0 net=839
rlabel metal2 268 -455 268 -455 0 net=1597
rlabel metal2 65 -457 65 -457 0 net=961
rlabel metal2 275 -457 275 -457 0 net=1263
rlabel metal2 324 -457 324 -457 0 net=1433
rlabel metal2 47 -459 47 -459 0 net=1075
rlabel metal2 282 -459 282 -459 0 net=1169
rlabel metal2 65 -461 65 -461 0 net=901
rlabel metal2 184 -463 184 -463 0 net=605
rlabel metal2 205 -465 205 -465 0 net=681
rlabel metal2 9 -476 9 -476 0 net=855
rlabel metal2 142 -476 142 -476 0 net=677
rlabel metal2 247 -476 247 -476 0 net=669
rlabel metal2 261 -476 261 -476 0 net=1444
rlabel metal2 352 -476 352 -476 0 net=1299
rlabel metal2 418 -476 418 -476 0 net=800
rlabel metal2 464 -476 464 -476 0 net=1003
rlabel metal2 464 -476 464 -476 0 net=1003
rlabel metal2 30 -478 30 -478 0 net=246
rlabel metal2 250 -478 250 -478 0 net=1202
rlabel metal2 345 -478 345 -478 0 net=1225
rlabel metal2 373 -478 373 -478 0 net=1505
rlabel metal2 373 -478 373 -478 0 net=1505
rlabel metal2 387 -478 387 -478 0 net=1617
rlabel metal2 422 -478 422 -478 0 net=1632
rlabel metal2 33 -480 33 -480 0 net=42
rlabel metal2 222 -480 222 -480 0 net=1160
rlabel metal2 432 -480 432 -480 0 net=1578
rlabel metal2 37 -482 37 -482 0 net=944
rlabel metal2 131 -482 131 -482 0 net=1191
rlabel metal2 380 -482 380 -482 0 net=1599
rlabel metal2 415 -482 415 -482 0 net=1329
rlabel metal2 16 -484 16 -484 0 net=1102
rlabel metal2 40 -484 40 -484 0 net=1086
rlabel metal2 72 -484 72 -484 0 net=926
rlabel metal2 100 -484 100 -484 0 net=479
rlabel metal2 173 -484 173 -484 0 net=915
rlabel metal2 205 -484 205 -484 0 net=683
rlabel metal2 264 -484 264 -484 0 net=1264
rlabel metal2 359 -484 359 -484 0 net=1377
rlabel metal2 16 -486 16 -486 0 net=539
rlabel metal2 44 -486 44 -486 0 net=569
rlabel metal2 180 -486 180 -486 0 net=109
rlabel metal2 51 -488 51 -488 0 net=808
rlabel metal2 107 -488 107 -488 0 net=611
rlabel metal2 240 -488 240 -488 0 net=945
rlabel metal2 51 -490 51 -490 0 net=411
rlabel metal2 82 -490 82 -490 0 net=415
rlabel metal2 191 -490 191 -490 0 net=719
rlabel metal2 275 -490 275 -490 0 net=1076
rlabel metal2 285 -490 285 -490 0 net=1460
rlabel metal2 429 -490 429 -490 0 net=1394
rlabel metal2 58 -492 58 -492 0 net=567
rlabel metal2 93 -492 93 -492 0 net=651
rlabel metal2 114 -492 114 -492 0 net=543
rlabel metal2 114 -492 114 -492 0 net=543
rlabel metal2 128 -492 128 -492 0 net=397
rlabel metal2 184 -492 184 -492 0 net=607
rlabel metal2 212 -492 212 -492 0 net=787
rlabel metal2 296 -492 296 -492 0 net=1141
rlabel metal2 359 -492 359 -492 0 net=1435
rlabel metal2 443 -492 443 -492 0 net=1399
rlabel metal2 79 -494 79 -494 0 net=1176
rlabel metal2 107 -496 107 -496 0 net=385
rlabel metal2 156 -496 156 -496 0 net=645
rlabel metal2 268 -496 268 -496 0 net=963
rlabel metal2 121 -498 121 -498 0 net=512
rlabel metal2 170 -498 170 -498 0 net=841
rlabel metal2 289 -498 289 -498 0 net=1093
rlabel metal2 303 -498 303 -498 0 net=1123
rlabel metal2 65 -500 65 -500 0 net=903
rlabel metal2 310 -500 310 -500 0 net=1171
rlabel metal2 65 -502 65 -502 0 net=465
rlabel metal2 156 -502 156 -502 0 net=623
rlabel metal2 243 -502 243 -502 0 net=1337
rlabel metal2 86 -504 86 -504 0 net=773
rlabel metal2 163 -504 163 -504 0 net=417
rlabel metal2 149 -506 149 -506 0 net=449
rlabel metal2 9 -517 9 -517 0 net=856
rlabel metal2 72 -517 72 -517 0 net=652
rlabel metal2 117 -517 117 -517 0 net=137
rlabel metal2 138 -517 138 -517 0 net=946
rlabel metal2 9 -519 9 -519 0 net=495
rlabel metal2 121 -519 121 -519 0 net=612
rlabel metal2 243 -519 243 -519 0 net=670
rlabel metal2 278 -519 278 -519 0 net=1226
rlabel metal2 366 -519 366 -519 0 net=1511
rlabel metal2 429 -519 429 -519 0 net=1515
rlabel metal2 16 -521 16 -521 0 net=540
rlabel metal2 44 -521 44 -521 0 net=570
rlabel metal2 208 -521 208 -521 0 net=1124
rlabel metal2 401 -521 401 -521 0 net=1300
rlabel metal2 443 -521 443 -521 0 net=1401
rlabel metal2 19 -523 19 -523 0 net=3
rlabel metal2 285 -523 285 -523 0 net=1378
rlabel metal2 457 -523 457 -523 0 net=1004
rlabel metal2 37 -525 37 -525 0 net=625
rlabel metal2 166 -525 166 -525 0 net=1461
rlabel metal2 303 -525 303 -525 0 net=1618
rlabel metal2 450 -525 450 -525 0 net=1331
rlabel metal2 44 -527 44 -527 0 net=413
rlabel metal2 58 -527 58 -527 0 net=568
rlabel metal2 124 -527 124 -527 0 net=238
rlabel metal2 184 -527 184 -527 0 net=646
rlabel metal2 212 -527 212 -527 0 net=964
rlabel metal2 359 -527 359 -527 0 net=1437
rlabel metal2 30 -529 30 -529 0 net=647
rlabel metal2 72 -529 72 -529 0 net=521
rlabel metal2 173 -529 173 -529 0 net=653
rlabel metal2 30 -531 30 -531 0 net=391
rlabel metal2 149 -531 149 -531 0 net=450
rlabel metal2 212 -531 212 -531 0 net=843
rlabel metal2 306 -531 306 -531 0 net=261
rlabel metal2 373 -531 373 -531 0 net=1507
rlabel metal2 26 -533 26 -533 0 net=745
rlabel metal2 310 -533 310 -533 0 net=1173
rlabel metal2 373 -533 373 -533 0 net=1251
rlabel metal2 51 -535 51 -535 0 net=467
rlabel metal2 82 -535 82 -535 0 net=1211
rlabel metal2 40 -537 40 -537 0 net=39
rlabel metal2 82 -537 82 -537 0 net=20
rlabel metal2 324 -537 324 -537 0 net=1339
rlabel metal2 86 -539 86 -539 0 net=775
rlabel metal2 184 -539 184 -539 0 net=1207
rlabel metal2 86 -541 86 -541 0 net=387
rlabel metal2 149 -541 149 -541 0 net=419
rlabel metal2 198 -541 198 -541 0 net=917
rlabel metal2 331 -541 331 -541 0 net=1193
rlabel metal2 107 -543 107 -543 0 net=399
rlabel metal2 163 -543 163 -543 0 net=416
rlabel metal2 219 -543 219 -543 0 net=721
rlabel metal2 233 -543 233 -543 0 net=679
rlabel metal2 103 -545 103 -545 0 net=455
rlabel metal2 135 -545 135 -545 0 net=361
rlabel metal2 191 -545 191 -545 0 net=609
rlabel metal2 233 -545 233 -545 0 net=1600
rlabel metal2 114 -547 114 -547 0 net=545
rlabel metal2 240 -547 240 -547 0 net=1475
rlabel metal2 191 -549 191 -549 0 net=821
rlabel metal2 247 -549 247 -549 0 net=789
rlabel metal2 282 -549 282 -549 0 net=1553
rlabel metal2 247 -551 247 -551 0 net=685
rlabel metal2 296 -551 296 -551 0 net=1095
rlabel metal2 23 -553 23 -553 0 net=863
rlabel metal2 317 -553 317 -553 0 net=1143
rlabel metal2 236 -555 236 -555 0 net=1103
rlabel metal2 289 -555 289 -555 0 net=905
rlabel metal2 142 -557 142 -557 0 net=481
rlabel metal2 114 -559 114 -559 0 net=713
rlabel metal2 9 -570 9 -570 0 net=497
rlabel metal2 198 -570 198 -570 0 net=547
rlabel metal2 198 -570 198 -570 0 net=547
rlabel metal2 212 -570 212 -570 0 net=844
rlabel metal2 303 -570 303 -570 0 net=1144
rlabel metal2 415 -570 415 -570 0 net=1509
rlabel metal2 415 -570 415 -570 0 net=1509
rlabel metal2 422 -570 422 -570 0 net=1513
rlabel metal2 422 -570 422 -570 0 net=1513
rlabel metal2 443 -570 443 -570 0 net=1402
rlabel metal2 443 -570 443 -570 0 net=1402
rlabel metal2 464 -570 464 -570 0 net=1333
rlabel metal2 16 -572 16 -572 0 net=70
rlabel metal2 121 -572 121 -572 0 net=867
rlabel metal2 121 -572 121 -572 0 net=867
rlabel metal2 138 -572 138 -572 0 net=1083
rlabel metal2 341 -572 341 -572 0 net=1340
rlabel metal2 457 -572 457 -572 0 net=845
rlabel metal2 16 -574 16 -574 0 net=907
rlabel metal2 163 -574 163 -574 0 net=269
rlabel metal2 23 -576 23 -576 0 net=457
rlabel metal2 163 -576 163 -576 0 net=1389
rlabel metal2 226 -576 226 -576 0 net=723
rlabel metal2 226 -576 226 -576 0 net=723
rlabel metal2 233 -576 233 -576 0 net=686
rlabel metal2 257 -576 257 -576 0 net=1554
rlabel metal2 9 -578 9 -578 0 net=1115
rlabel metal2 236 -578 236 -578 0 net=1212
rlabel metal2 394 -578 394 -578 0 net=1517
rlabel metal2 30 -580 30 -580 0 net=392
rlabel metal2 170 -580 170 -580 0 net=183
rlabel metal2 33 -582 33 -582 0 net=414
rlabel metal2 58 -582 58 -582 0 net=648
rlabel metal2 93 -582 93 -582 0 net=317
rlabel metal2 247 -582 247 -582 0 net=906
rlabel metal2 40 -584 40 -584 0 net=1601
rlabel metal2 44 -586 44 -586 0 net=469
rlabel metal2 58 -586 58 -586 0 net=401
rlabel metal2 149 -586 149 -586 0 net=421
rlabel metal2 317 -586 317 -586 0 net=1195
rlabel metal2 37 -588 37 -588 0 net=627
rlabel metal2 65 -588 65 -588 0 net=777
rlabel metal2 173 -588 173 -588 0 net=610
rlabel metal2 240 -588 240 -588 0 net=1174
rlabel metal2 68 -590 68 -590 0 net=1233
rlabel metal2 352 -590 352 -590 0 net=1209
rlabel metal2 79 -592 79 -592 0 net=482
rlabel metal2 331 -592 331 -592 0 net=1565
rlabel metal2 72 -594 72 -594 0 net=523
rlabel metal2 93 -594 93 -594 0 net=655
rlabel metal2 30 -596 30 -596 0 net=1633
rlabel metal2 72 -598 72 -598 0 net=389
rlabel metal2 107 -598 107 -598 0 net=377
rlabel metal2 205 -598 205 -598 0 net=1523
rlabel metal2 240 -598 240 -598 0 net=747
rlabel metal2 289 -598 289 -598 0 net=1097
rlabel metal2 359 -598 359 -598 0 net=1439
rlabel metal2 86 -600 86 -600 0 net=714
rlabel metal2 156 -600 156 -600 0 net=663
rlabel metal2 177 -600 177 -600 0 net=823
rlabel metal2 219 -600 219 -600 0 net=791
rlabel metal2 306 -600 306 -600 0 net=1549
rlabel metal2 135 -602 135 -602 0 net=363
rlabel metal2 180 -602 180 -602 0 net=680
rlabel metal2 142 -604 142 -604 0 net=737
rlabel metal2 254 -604 254 -604 0 net=1463
rlabel metal2 268 -606 268 -606 0 net=919
rlabel metal2 338 -606 338 -606 0 net=1301
rlabel metal2 261 -608 261 -608 0 net=1105
rlabel metal2 338 -608 338 -608 0 net=1253
rlabel metal2 275 -610 275 -610 0 net=865
rlabel metal2 373 -610 373 -610 0 net=1477
rlabel metal2 296 -612 296 -612 0 net=1411
rlabel metal2 387 -612 387 -612 0 net=1293
rlabel metal2 2 -623 2 -623 0 net=629
rlabel metal2 72 -623 72 -623 0 net=390
rlabel metal2 117 -623 117 -623 0 net=215
rlabel metal2 222 -623 222 -623 0 net=920
rlabel metal2 299 -623 299 -623 0 net=1514
rlabel metal2 436 -623 436 -623 0 net=1635
rlabel metal2 450 -623 450 -623 0 net=846
rlabel metal2 460 -623 460 -623 0 net=278
rlabel metal2 471 -623 471 -623 0 net=1335
rlabel metal2 471 -623 471 -623 0 net=1335
rlabel metal2 9 -625 9 -625 0 net=1116
rlabel metal2 170 -625 170 -625 0 net=498
rlabel metal2 187 -625 187 -625 0 net=422
rlabel metal2 299 -625 299 -625 0 net=1510
rlabel metal2 429 -625 429 -625 0 net=1603
rlabel metal2 9 -627 9 -627 0 net=1071
rlabel metal2 79 -627 79 -627 0 net=524
rlabel metal2 142 -627 142 -627 0 net=739
rlabel metal2 191 -627 191 -627 0 net=59
rlabel metal2 233 -627 233 -627 0 net=1525
rlabel metal2 23 -629 23 -629 0 net=458
rlabel metal2 142 -629 142 -629 0 net=725
rlabel metal2 240 -629 240 -629 0 net=748
rlabel metal2 261 -629 261 -629 0 net=1210
rlabel metal2 373 -629 373 -629 0 net=1479
rlabel metal2 373 -629 373 -629 0 net=1479
rlabel metal2 380 -629 380 -629 0 net=1551
rlabel metal2 16 -631 16 -631 0 net=909
rlabel metal2 30 -631 30 -631 0 net=1391
rlabel metal2 194 -631 194 -631 0 net=1464
rlabel metal2 415 -631 415 -631 0 net=1471
rlabel metal2 16 -633 16 -633 0 net=779
rlabel metal2 93 -633 93 -633 0 net=657
rlabel metal2 128 -633 128 -633 0 net=248
rlabel metal2 205 -633 205 -633 0 net=1084
rlabel metal2 310 -633 310 -633 0 net=1107
rlabel metal2 310 -633 310 -633 0 net=1107
rlabel metal2 331 -633 331 -633 0 net=1440
rlabel metal2 33 -635 33 -635 0 net=593
rlabel metal2 86 -635 86 -635 0 net=705
rlabel metal2 135 -635 135 -635 0 net=365
rlabel metal2 208 -635 208 -635 0 net=1294
rlabel metal2 37 -637 37 -637 0 net=548
rlabel metal2 215 -637 215 -637 0 net=1033
rlabel metal2 289 -637 289 -637 0 net=1099
rlabel metal2 331 -637 331 -637 0 net=1283
rlabel metal2 387 -637 387 -637 0 net=1519
rlabel metal2 37 -639 37 -639 0 net=825
rlabel metal2 180 -639 180 -639 0 net=1425
rlabel metal2 40 -641 40 -641 0 net=13
rlabel metal2 334 -641 334 -641 0 net=1302
rlabel metal2 44 -643 44 -643 0 net=470
rlabel metal2 54 -643 54 -643 0 net=1581
rlabel metal2 44 -645 44 -645 0 net=866
rlabel metal2 345 -645 345 -645 0 net=1235
rlabel metal2 58 -647 58 -647 0 net=403
rlabel metal2 93 -647 93 -647 0 net=869
rlabel metal2 156 -647 156 -647 0 net=665
rlabel metal2 219 -647 219 -647 0 net=793
rlabel metal2 243 -647 243 -647 0 net=1415
rlabel metal2 366 -647 366 -647 0 net=1567
rlabel metal2 58 -649 58 -649 0 net=697
rlabel metal2 163 -649 163 -649 0 net=715
rlabel metal2 226 -649 226 -649 0 net=763
rlabel metal2 254 -649 254 -649 0 net=835
rlabel metal2 107 -651 107 -651 0 net=379
rlabel metal2 184 -651 184 -651 0 net=1067
rlabel metal2 324 -651 324 -651 0 net=1413
rlabel metal2 100 -653 100 -653 0 net=753
rlabel metal2 114 -653 114 -653 0 net=285
rlabel metal2 240 -653 240 -653 0 net=1131
rlabel metal2 338 -653 338 -653 0 net=1255
rlabel metal2 100 -655 100 -655 0 net=1309
rlabel metal2 261 -655 261 -655 0 net=1197
rlabel metal2 103 -657 103 -657 0 net=1395
rlabel metal2 250 -659 250 -659 0 net=1125
rlabel metal2 250 -661 250 -661 0 net=1423
rlabel metal2 275 -663 275 -663 0 net=1023
rlabel metal2 2 -674 2 -674 0 net=630
rlabel metal2 135 -674 135 -674 0 net=366
rlabel metal2 187 -674 187 -674 0 net=167
rlabel metal2 233 -674 233 -674 0 net=794
rlabel metal2 250 -674 250 -674 0 net=1100
rlabel metal2 331 -674 331 -674 0 net=1397
rlabel metal2 387 -674 387 -674 0 net=1521
rlabel metal2 387 -674 387 -674 0 net=1521
rlabel metal2 443 -674 443 -674 0 net=1636
rlabel metal2 464 -674 464 -674 0 net=1336
rlabel metal2 16 -676 16 -676 0 net=780
rlabel metal2 114 -676 114 -676 0 net=380
rlabel metal2 170 -676 170 -676 0 net=740
rlabel metal2 191 -676 191 -676 0 net=1126
rlabel metal2 334 -676 334 -676 0 net=1552
rlabel metal2 9 -678 9 -678 0 net=1073
rlabel metal2 37 -678 37 -678 0 net=826
rlabel metal2 191 -678 191 -678 0 net=765
rlabel metal2 250 -678 250 -678 0 net=1604
rlabel metal2 9 -680 9 -680 0 net=871
rlabel metal2 128 -680 128 -680 0 net=1424
rlabel metal2 23 -682 23 -682 0 net=911
rlabel metal2 149 -682 149 -682 0 net=531
rlabel metal2 268 -682 268 -682 0 net=1203
rlabel metal2 380 -682 380 -682 0 net=1237
rlabel metal2 23 -684 23 -684 0 net=1069
rlabel metal2 296 -684 296 -684 0 net=1414
rlabel metal2 380 -684 380 -684 0 net=1569
rlabel metal2 37 -686 37 -686 0 net=172
rlabel metal2 212 -686 212 -686 0 net=1526
rlabel metal2 40 -688 40 -688 0 net=15
rlabel metal2 170 -688 170 -688 0 net=1009
rlabel metal2 229 -688 229 -688 0 net=1117
rlabel metal2 299 -688 299 -688 0 net=1256
rlabel metal2 359 -688 359 -688 0 net=1417
rlabel metal2 401 -688 401 -688 0 net=1473
rlabel metal2 44 -690 44 -690 0 net=707
rlabel metal2 177 -690 177 -690 0 net=1034
rlabel metal2 345 -690 345 -690 0 net=1285
rlabel metal2 359 -690 359 -690 0 net=1481
rlabel metal2 51 -692 51 -692 0 net=1469
rlabel metal2 58 -694 58 -694 0 net=699
rlabel metal2 194 -694 194 -694 0 net=883
rlabel metal2 268 -694 268 -694 0 net=1109
rlabel metal2 58 -696 58 -696 0 net=837
rlabel metal2 261 -696 261 -696 0 net=1199
rlabel metal2 72 -698 72 -698 0 net=431
rlabel metal2 198 -698 198 -698 0 net=666
rlabel metal2 254 -698 254 -698 0 net=1025
rlabel metal2 282 -698 282 -698 0 net=1133
rlabel metal2 2 -700 2 -700 0 net=1539
rlabel metal2 75 -700 75 -700 0 net=10
rlabel metal2 261 -700 261 -700 0 net=1027
rlabel metal2 79 -702 79 -702 0 net=405
rlabel metal2 142 -702 142 -702 0 net=726
rlabel metal2 324 -702 324 -702 0 net=1427
rlabel metal2 82 -704 82 -704 0 net=754
rlabel metal2 142 -704 142 -704 0 net=1311
rlabel metal2 184 -704 184 -704 0 net=999
rlabel metal2 394 -704 394 -704 0 net=1583
rlabel metal2 65 -706 65 -706 0 net=595
rlabel metal2 156 -706 156 -706 0 net=717
rlabel metal2 54 -708 54 -708 0 net=1021
rlabel metal2 86 -708 86 -708 0 net=827
rlabel metal2 121 -710 121 -710 0 net=659
rlabel metal2 30 -712 30 -712 0 net=1392
rlabel metal2 30 -714 30 -714 0 net=1147
rlabel metal2 9 -725 9 -725 0 net=872
rlabel metal2 96 -725 96 -725 0 net=12
rlabel metal2 198 -725 198 -725 0 net=1470
rlabel metal2 376 -725 376 -725 0 net=1474
rlabel metal2 411 -725 411 -725 0 net=1238
rlabel metal2 16 -727 16 -727 0 net=1074
rlabel metal2 110 -727 110 -727 0 net=176
rlabel metal2 254 -727 254 -727 0 net=1026
rlabel metal2 289 -727 289 -727 0 net=1118
rlabel metal2 338 -727 338 -727 0 net=1571
rlabel metal2 387 -727 387 -727 0 net=1522
rlabel metal2 23 -729 23 -729 0 net=1070
rlabel metal2 215 -729 215 -729 0 net=1000
rlabel metal2 243 -729 243 -729 0 net=1200
rlabel metal2 341 -729 341 -729 0 net=1286
rlabel metal2 2 -731 2 -731 0 net=1541
rlabel metal2 345 -731 345 -731 0 net=1483
rlabel metal2 23 -733 23 -733 0 net=829
rlabel metal2 121 -733 121 -733 0 net=1527
rlabel metal2 37 -735 37 -735 0 net=8
rlabel metal2 86 -735 86 -735 0 net=767
rlabel metal2 233 -735 233 -735 0 net=1110
rlabel metal2 289 -735 289 -735 0 net=1429
rlabel metal2 37 -737 37 -737 0 net=54
rlabel metal2 205 -737 205 -737 0 net=1239
rlabel metal2 324 -737 324 -737 0 net=1585
rlabel metal2 40 -739 40 -739 0 net=838
rlabel metal2 65 -739 65 -739 0 net=1022
rlabel metal2 128 -739 128 -739 0 net=1137
rlabel metal2 16 -741 16 -741 0 net=603
rlabel metal2 114 -741 114 -741 0 net=407
rlabel metal2 135 -741 135 -741 0 net=701
rlabel metal2 247 -741 247 -741 0 net=1135
rlabel metal2 44 -743 44 -743 0 net=709
rlabel metal2 236 -743 236 -743 0 net=1347
rlabel metal2 44 -745 44 -745 0 net=817
rlabel metal2 93 -745 93 -745 0 net=913
rlabel metal2 142 -745 142 -745 0 net=1312
rlabel metal2 51 -747 51 -747 0 net=695
rlabel metal2 100 -747 100 -747 0 net=433
rlabel metal2 149 -747 149 -747 0 net=533
rlabel metal2 149 -747 149 -747 0 net=533
rlabel metal2 156 -747 156 -747 0 net=718
rlabel metal2 54 -749 54 -749 0 net=847
rlabel metal2 82 -751 82 -751 0 net=131
rlabel metal2 163 -751 163 -751 0 net=661
rlabel metal2 180 -751 180 -751 0 net=1204
rlabel metal2 100 -753 100 -753 0 net=1028
rlabel metal2 30 -755 30 -755 0 net=1149
rlabel metal2 103 -757 103 -757 0 net=181
rlabel metal2 107 -759 107 -759 0 net=597
rlabel metal2 163 -759 163 -759 0 net=1303
rlabel metal2 219 -761 219 -761 0 net=885
rlabel metal2 212 -763 212 -763 0 net=1011
rlabel metal2 212 -765 212 -765 0 net=1398
rlabel metal2 331 -767 331 -767 0 net=1418
rlabel metal2 9 -778 9 -778 0 net=1177
rlabel metal2 58 -778 58 -778 0 net=604
rlabel metal2 110 -778 110 -778 0 net=598
rlabel metal2 177 -778 177 -778 0 net=1528
rlabel metal2 317 -778 317 -778 0 net=1573
rlabel metal2 30 -780 30 -780 0 net=696
rlabel metal2 65 -780 65 -780 0 net=818
rlabel metal2 93 -780 93 -780 0 net=434
rlabel metal2 177 -780 177 -780 0 net=886
rlabel metal2 233 -780 233 -780 0 net=1151
rlabel metal2 268 -780 268 -780 0 net=1241
rlabel metal2 268 -780 268 -780 0 net=1241
rlabel metal2 51 -782 51 -782 0 net=128
rlabel metal2 96 -782 96 -782 0 net=1138
rlabel metal2 72 -784 72 -784 0 net=619
rlabel metal2 100 -784 100 -784 0 net=373
rlabel metal2 163 -784 163 -784 0 net=1305
rlabel metal2 103 -786 103 -786 0 net=1605
rlabel metal2 107 -788 107 -788 0 net=848
rlabel metal2 247 -788 247 -788 0 net=1136
rlabel metal2 30 -790 30 -790 0 net=1179
rlabel metal2 254 -790 254 -790 0 net=1349
rlabel metal2 117 -792 117 -792 0 net=662
rlabel metal2 198 -792 198 -792 0 net=849
rlabel metal2 198 -792 198 -792 0 net=849
rlabel metal2 205 -792 205 -792 0 net=881
rlabel metal2 219 -792 219 -792 0 net=1013
rlabel metal2 282 -792 282 -792 0 net=1431
rlabel metal2 23 -794 23 -794 0 net=831
rlabel metal2 212 -794 212 -794 0 net=549
rlabel metal2 23 -796 23 -796 0 net=1145
rlabel metal2 124 -796 124 -796 0 net=914
rlabel metal2 163 -796 163 -796 0 net=711
rlabel metal2 33 -798 33 -798 0 net=947
rlabel metal2 149 -798 149 -798 0 net=535
rlabel metal2 33 -800 33 -800 0 net=340
rlabel metal2 124 -800 124 -800 0 net=702
rlabel metal2 37 -802 37 -802 0 net=1543
rlabel metal2 37 -804 37 -804 0 net=525
rlabel metal2 128 -804 128 -804 0 net=409
rlabel metal2 86 -806 86 -806 0 net=769
rlabel metal2 131 -808 131 -808 0 net=1542
rlabel metal2 310 -810 310 -810 0 net=1587
rlabel metal2 324 -812 324 -812 0 net=1485
rlabel metal2 9 -823 9 -823 0 net=1178
rlabel metal2 23 -823 23 -823 0 net=1146
rlabel metal2 72 -823 72 -823 0 net=621
rlabel metal2 96 -823 96 -823 0 net=1152
rlabel metal2 240 -823 240 -823 0 net=1242
rlabel metal2 282 -823 282 -823 0 net=1432
rlabel metal2 282 -823 282 -823 0 net=1432
rlabel metal2 292 -823 292 -823 0 net=1574
rlabel metal2 324 -823 324 -823 0 net=1486
rlabel metal2 23 -825 23 -825 0 net=1307
rlabel metal2 310 -825 310 -825 0 net=1588
rlabel metal2 33 -827 33 -827 0 net=298
rlabel metal2 58 -827 58 -827 0 net=1153
rlabel metal2 86 -827 86 -827 0 net=981
rlabel metal2 117 -827 117 -827 0 net=536
rlabel metal2 222 -827 222 -827 0 net=1014
rlabel metal2 254 -827 254 -827 0 net=1351
rlabel metal2 37 -829 37 -829 0 net=526
rlabel metal2 117 -829 117 -829 0 net=1544
rlabel metal2 33 -831 33 -831 0 net=1127
rlabel metal2 72 -831 72 -831 0 net=375
rlabel metal2 124 -831 124 -831 0 net=712
rlabel metal2 184 -831 184 -831 0 net=770
rlabel metal2 184 -831 184 -831 0 net=770
rlabel metal2 191 -831 191 -831 0 net=1181
rlabel metal2 51 -833 51 -833 0 net=895
rlabel metal2 212 -833 212 -833 0 net=550
rlabel metal2 44 -835 44 -835 0 net=123
rlabel metal2 128 -835 128 -835 0 net=410
rlabel metal2 205 -835 205 -835 0 net=882
rlabel metal2 19 -837 19 -837 0 net=223
rlabel metal2 135 -837 135 -837 0 net=948
rlabel metal2 135 -839 135 -839 0 net=21
rlabel metal2 149 -839 149 -839 0 net=851
rlabel metal2 152 -841 152 -841 0 net=1606
rlabel metal2 156 -843 156 -843 0 net=833
rlabel metal2 170 -845 170 -845 0 net=1487
rlabel metal2 23 -856 23 -856 0 net=1308
rlabel metal2 187 -856 187 -856 0 net=1182
rlabel metal2 268 -856 268 -856 0 net=1352
rlabel metal2 37 -858 37 -858 0 net=1128
rlabel metal2 47 -858 47 -858 0 net=1154
rlabel metal2 65 -858 65 -858 0 net=982
rlabel metal2 93 -858 93 -858 0 net=622
rlabel metal2 131 -858 131 -858 0 net=852
rlabel metal2 54 -860 54 -860 0 net=1488
rlabel metal2 72 -862 72 -862 0 net=376
rlabel metal2 107 -862 107 -862 0 net=834
rlabel metal2 82 -864 82 -864 0 net=896
<< end >>
